

module b21_C_2inp_gates_syn ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, 
        P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, 
        P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, 
        P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, 
        P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, 
        P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, 
        P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, 
        P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, 
        P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, 
        P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, 
        P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, 
        P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, 
        P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, 
        P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, 
        P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, 
        P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, 
        P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, 
        P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, 
        P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, 
        P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, 
        P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, 
        P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, 
        P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, 
        P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, 
        P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, 
        ADD_1071_U57, ADD_1071_U58, ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, 
        ADD_1071_U62, ADD_1071_U63, ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, 
        ADD_1071_U50, ADD_1071_U51, ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, 
        ADD_1071_U5, ADD_1071_U46, U126, U123, P1_U3353, P1_U3352, P1_U3351, 
        P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, 
        P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, 
        P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, 
        P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, 
        P1_U3322, P1_U3440, P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, 
        P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, 
        P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, 
        P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, 
        P1_U3296, P1_U3295, P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, 
        P1_U3460, P1_U3463, P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, 
        P1_U3481, P1_U3484, P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, 
        P1_U3502, P1_U3505, P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, 
        P1_U3514, P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, 
        P1_U3521, P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, 
        P1_U3528, P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, 
        P1_U3535, P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, 
        P1_U3542, P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, 
        P1_U3549, P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, 
        P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, 
        P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, 
        P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, 
        P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, 
        P1_U3355, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, 
        P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, 
        P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, 
        P1_U3242, P1_U3241, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, 
        P1_U3560, P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, 
        P1_U3567, P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, 
        P1_U3574, P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, 
        P1_U3581, P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, 
        P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, 
        P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, 
        P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, 
        P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, 
        P1_U3211, P1_U3084, P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, 
        P2_U3355, P2_U3354, P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, 
        P2_U3348, P2_U3347, P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, 
        P2_U3341, P2_U3340, P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, 
        P2_U3334, P2_U3333, P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, 
        P2_U3327, P2_U3437, P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, 
        P2_U3322, P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, 
        P2_U3315, P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, 
        P2_U3308, P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, 
        P2_U3301, P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, 
        P2_U3457, P2_U3460, P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, 
        P2_U3478, P2_U3481, P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, 
        P2_U3499, P2_U3502, P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, 
        P2_U3511, P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, 
        P2_U3518, P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, 
        P2_U3525, P2_U3526, P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, 
        P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, 
        P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, 
        P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, 
        P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, 
        P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, 
        P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, 
        P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, 
        P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, 
        P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, 
        P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, 
        P2_U3246, P2_U3245, P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, 
        P2_U3557, P2_U3558, P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, 
        P2_U3564, P2_U3565, P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, 
        P2_U3571, P2_U3572, P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, 
        P2_U3578, P2_U3579, P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, 
        P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, 
        P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, 
        P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, 
        P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, 
        P2_U3215, P2_U3152, P2_U3151, P2_U3966, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, 
        keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, 
        keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, 
        keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, 
        keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, 
        keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, 
        keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, 
        keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, 
        keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, 
        keyinput113, keyinput114, keyinput115, keyinput116, keyinput117, 
        keyinput118, keyinput119, keyinput120, keyinput121, keyinput122, 
        keyinput123, keyinput124, keyinput125, keyinput126, keyinput127 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN,
         P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN,
         P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN,
         P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN,
         P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN,
         P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN,
         P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN,
         P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN,
         P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN,
         P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN,
         P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN,
         P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN,
         P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN,
         P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN,
         P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN,
         P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN,
         P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN,
         P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN,
         P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN,
         P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN,
         P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN,
         P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
         keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
         keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
         keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
         keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
         keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
         keyinput90, keyinput91, keyinput92, keyinput93, keyinput94,
         keyinput95, keyinput96, keyinput97, keyinput98, keyinput99,
         keyinput100, keyinput101, keyinput102, keyinput103, keyinput104,
         keyinput105, keyinput106, keyinput107, keyinput108, keyinput109,
         keyinput110, keyinput111, keyinput112, keyinput113, keyinput114,
         keyinput115, keyinput116, keyinput117, keyinput118, keyinput119,
         keyinput120, keyinput121, keyinput122, keyinput123, keyinput124,
         keyinput125, keyinput126, keyinput127;
  output ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, ADD_1071_U57, ADD_1071_U58,
         ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, ADD_1071_U62, ADD_1071_U63,
         ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, ADD_1071_U50, ADD_1071_U51,
         ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, ADD_1071_U5, ADD_1071_U46,
         U126, U123, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349,
         P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342,
         P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335,
         P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328,
         P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, P1_U3322, P1_U3440,
         P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316,
         P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309,
         P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302,
         P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295,
         P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, P1_U3460, P1_U3463,
         P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, P1_U3481, P1_U3484,
         P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, P1_U3502, P1_U3505,
         P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515,
         P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522,
         P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529,
         P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536,
         P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543,
         P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550,
         P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, P1_U3290, P1_U3289,
         P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282,
         P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275,
         P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268,
         P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, P1_U3355, P1_U3262,
         P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255,
         P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248,
         P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3242, P1_U3241,
         P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561,
         P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568,
         P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575,
         P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582,
         P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, P1_U3239, P1_U3238,
         P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231,
         P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224,
         P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217,
         P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, P1_U3084,
         P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, P2_U3355, P2_U3354,
         P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, P2_U3348, P2_U3347,
         P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, P2_U3341, P2_U3340,
         P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, P2_U3334, P2_U3333,
         P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, P2_U3327, P2_U3437,
         P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321,
         P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314,
         P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307,
         P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300,
         P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, P2_U3457, P2_U3460,
         P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481,
         P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, P2_U3499, P2_U3502,
         P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512,
         P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519,
         P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526,
         P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, P2_U3532, P2_U3533,
         P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540,
         P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547,
         P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, P2_U3295, P2_U3294,
         P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287,
         P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280,
         P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273,
         P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266,
         P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259,
         P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252,
         P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245,
         P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558,
         P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, P2_U3564, P2_U3565,
         P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, P2_U3571, P2_U3572,
         P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, P2_U3578, P2_U3579,
         P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, P2_U3243, P2_U3242,
         P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235,
         P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228,
         P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221,
         P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3152,
         P2_U3151, P2_U3966;
  wire   n4391, n4392, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401,
         n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411,
         n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421,
         n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431,
         n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441,
         n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451,
         n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461,
         n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471,
         n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481,
         n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491,
         n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501,
         n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511,
         n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521,
         n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531,
         n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541,
         n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551,
         n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561,
         n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571,
         n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581,
         n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591,
         n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601,
         n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611,
         n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621,
         n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631,
         n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641,
         n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651,
         n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661,
         n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671,
         n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681,
         n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691,
         n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701,
         n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711,
         n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721,
         n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731,
         n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741,
         n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751,
         n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761,
         n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771,
         n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781,
         n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791,
         n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801,
         n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811,
         n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821,
         n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831,
         n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841,
         n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851,
         n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861,
         n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871,
         n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881,
         n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891,
         n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901,
         n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911,
         n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921,
         n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931,
         n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941,
         n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951,
         n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961,
         n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971,
         n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981,
         n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991,
         n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001,
         n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011,
         n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021,
         n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031,
         n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041,
         n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051,
         n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061,
         n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071,
         n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081,
         n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091,
         n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101,
         n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111,
         n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121,
         n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131,
         n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141,
         n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151,
         n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161,
         n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171,
         n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181,
         n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191,
         n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201,
         n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211,
         n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221,
         n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231,
         n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241,
         n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251,
         n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261,
         n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271,
         n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281,
         n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291,
         n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301,
         n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311,
         n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321,
         n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331,
         n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341,
         n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351,
         n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361,
         n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371,
         n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381,
         n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391,
         n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401,
         n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411,
         n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421,
         n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431,
         n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441,
         n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451,
         n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461,
         n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471,
         n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481,
         n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491,
         n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501,
         n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511,
         n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521,
         n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531,
         n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541,
         n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551,
         n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561,
         n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571,
         n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581,
         n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591,
         n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601,
         n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611,
         n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621,
         n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631,
         n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641,
         n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651,
         n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661,
         n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671,
         n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681,
         n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691,
         n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701,
         n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711,
         n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721,
         n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731,
         n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741,
         n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751,
         n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761,
         n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771,
         n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781,
         n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791,
         n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801,
         n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811,
         n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821,
         n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831,
         n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841,
         n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851,
         n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861,
         n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871,
         n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881,
         n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891,
         n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901,
         n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911,
         n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921,
         n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931,
         n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941,
         n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951,
         n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961,
         n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971,
         n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981,
         n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991,
         n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001,
         n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011,
         n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021,
         n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031,
         n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041,
         n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051,
         n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061,
         n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071,
         n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081,
         n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091,
         n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101,
         n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111,
         n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121,
         n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131,
         n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141,
         n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151,
         n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161,
         n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171,
         n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181,
         n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191,
         n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201,
         n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211,
         n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221,
         n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231,
         n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241,
         n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251,
         n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261,
         n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271,
         n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281,
         n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291,
         n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301,
         n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311,
         n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321,
         n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331,
         n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341,
         n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351,
         n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361,
         n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371,
         n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381,
         n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391,
         n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401,
         n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411,
         n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421,
         n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431,
         n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441,
         n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451,
         n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461,
         n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471,
         n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481,
         n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491,
         n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501,
         n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511,
         n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521,
         n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531,
         n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541,
         n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551,
         n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561,
         n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571,
         n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581,
         n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591,
         n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601,
         n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611,
         n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621,
         n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631,
         n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641,
         n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651,
         n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661,
         n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671,
         n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681,
         n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691,
         n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701,
         n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711,
         n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721,
         n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731,
         n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741,
         n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751,
         n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761,
         n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771,
         n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781,
         n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791,
         n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801,
         n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811,
         n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821,
         n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831,
         n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841,
         n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851,
         n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861,
         n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871,
         n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881,
         n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891,
         n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901,
         n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911,
         n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921,
         n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931,
         n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941,
         n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951,
         n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961,
         n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971,
         n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981,
         n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991,
         n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001,
         n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011,
         n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021,
         n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031,
         n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041,
         n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051,
         n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061,
         n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071,
         n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081,
         n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091,
         n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101,
         n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111,
         n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121,
         n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131,
         n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141,
         n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151,
         n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161,
         n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171,
         n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181,
         n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191,
         n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201,
         n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211,
         n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221,
         n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231,
         n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241,
         n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251,
         n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261,
         n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271,
         n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281,
         n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291,
         n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301,
         n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311,
         n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321,
         n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331,
         n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341,
         n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351,
         n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361,
         n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371,
         n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381,
         n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391,
         n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401,
         n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411,
         n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421,
         n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431,
         n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441,
         n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451,
         n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461,
         n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471,
         n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481,
         n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491,
         n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501,
         n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511,
         n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521,
         n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531,
         n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541,
         n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551,
         n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561,
         n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571,
         n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581,
         n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591,
         n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601,
         n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611,
         n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621,
         n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631,
         n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641,
         n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651,
         n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661,
         n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671,
         n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681,
         n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691,
         n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701,
         n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711,
         n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721,
         n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731,
         n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741,
         n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751,
         n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761,
         n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771,
         n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781,
         n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791,
         n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801,
         n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811,
         n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821,
         n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831,
         n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841,
         n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851,
         n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861,
         n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871,
         n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881,
         n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891,
         n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901,
         n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911,
         n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921,
         n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931,
         n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941,
         n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951,
         n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961,
         n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971,
         n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981,
         n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991,
         n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001,
         n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011,
         n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021,
         n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031,
         n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041,
         n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051,
         n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061,
         n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071,
         n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081,
         n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091,
         n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101,
         n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111,
         n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121,
         n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131,
         n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141,
         n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151,
         n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161,
         n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171,
         n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181,
         n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191,
         n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201,
         n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211,
         n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221,
         n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231,
         n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241,
         n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251,
         n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261,
         n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271,
         n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281,
         n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291,
         n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301,
         n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311,
         n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321,
         n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331,
         n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341,
         n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351,
         n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361,
         n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371,
         n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381,
         n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391,
         n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401,
         n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411,
         n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421,
         n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431,
         n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441,
         n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451,
         n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461,
         n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471,
         n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481,
         n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491,
         n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501,
         n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511,
         n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521,
         n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531,
         n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541,
         n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551,
         n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561,
         n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571,
         n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581,
         n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591,
         n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601,
         n8602, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612,
         n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622,
         n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632,
         n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642,
         n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652,
         n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662,
         n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672,
         n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682,
         n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692,
         n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702,
         n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712,
         n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722,
         n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732,
         n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742,
         n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752,
         n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762,
         n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772,
         n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782,
         n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792,
         n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802,
         n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812,
         n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822,
         n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832,
         n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842,
         n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852,
         n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862,
         n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872,
         n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882,
         n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892,
         n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902,
         n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912,
         n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922,
         n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932,
         n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942,
         n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952,
         n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962,
         n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972,
         n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982,
         n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992,
         n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002,
         n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012,
         n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022,
         n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032,
         n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042,
         n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052,
         n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062,
         n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072,
         n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082,
         n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092,
         n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102,
         n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112,
         n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122,
         n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132,
         n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142,
         n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152,
         n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162,
         n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172,
         n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182,
         n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192,
         n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202,
         n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212,
         n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222,
         n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232,
         n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242,
         n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252,
         n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262,
         n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272,
         n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282,
         n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292,
         n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302,
         n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312,
         n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322,
         n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332,
         n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342,
         n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352,
         n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362,
         n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372,
         n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382,
         n9383, n9384, n9385, n9387, n9388, n9389, n9390, n9391, n9392, n9393,
         n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403,
         n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413,
         n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423,
         n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433,
         n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443,
         n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453,
         n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463,
         n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473,
         n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483,
         n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493,
         n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503,
         n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513,
         n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523,
         n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533,
         n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543,
         n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553,
         n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563,
         n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573,
         n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583,
         n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593,
         n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603,
         n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613,
         n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623,
         n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633,
         n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643,
         n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653,
         n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663,
         n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673,
         n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683,
         n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693,
         n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703,
         n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713,
         n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723,
         n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733,
         n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743,
         n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753,
         n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763,
         n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773,
         n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783,
         n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793,
         n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803,
         n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813,
         n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823,
         n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833,
         n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843,
         n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853,
         n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863,
         n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873,
         n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883,
         n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893,
         n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903,
         n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913,
         n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923,
         n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933,
         n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943,
         n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953,
         n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963,
         n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973,
         n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983,
         n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993,
         n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001, n10002,
         n10003, n10004, n10005, n10006, n10007, n10008, n10009, n10010,
         n10011, n10012, n10013, n10014, n10015, n10016, n10017, n10018,
         n10019, n10020, n10021, n10022, n10023, n10024, n10025, n10026,
         n10027, n10028, n10029, n10030, n10031, n10032, n10033, n10034,
         n10035, n10036, n10037, n10038, n10039, n10040, n10041, n10042,
         n10043, n10044, n10045, n10046, n10047, n10048, n10049, n10050,
         n10051, n10052, n10053, n10054, n10055, n10056, n10057, n10058,
         n10059, n10060, n10061, n10062, n10063, n10064, n10065, n10066,
         n10067, n10068, n10069, n10070, n10071, n10072, n10073, n10074,
         n10075, n10076, n10077, n10078, n10079, n10080, n10081, n10082,
         n10083, n10084, n10085, n10086, n10087, n10088, n10089, n10090,
         n10091, n10092, n10093, n10094, n10095, n10096, n10097, n10098,
         n10099, n10100, n10101, n10102, n10103, n10104, n10105, n10106,
         n10107, n10108, n10109, n10110, n10111, n10112, n10113, n10114,
         n10115, n10116, n10117, n10118, n10119, n10120, n10121, n10122,
         n10123, n10124, n10125, n10126, n10127, n10128, n10129, n10130,
         n10131, n10132, n10133, n10134, n10135, n10136, n10137, n10138,
         n10139, n10140, n10141, n10142, n10143, n10144, n10145, n10146,
         n10147, n10148, n10149, n10150, n10151, n10152, n10153, n10154,
         n10155, n10156, n10157, n10158, n10159, n10160, n10161, n10162,
         n10163, n10164, n10165, n10166, n10167, n10168, n10169, n10170,
         n10171, n10172, n10173, n10174, n10175, n10176, n10177, n10178,
         n10179, n10180, n10181, n10182, n10183, n10184, n10185, n10186,
         n10187, n10188, n10189, n10190, n10191, n10192, n10193, n10194,
         n10195, n10196, n10197, n10198, n10199, n10200, n10201, n10202,
         n10203, n10204, n10205, n10206, n10207, n10208, n10209, n10210,
         n10211, n10212, n10213, n10214, n10215, n10216, n10217, n10218,
         n10219, n10220, n10221, n10222, n10223, n10224, n10225, n10226,
         n10227, n10228, n10229, n10230, n10231, n10232, n10233, n10234,
         n10235, n10236, n10237, n10238, n10239, n10240, n10241, n10242,
         n10243, n10244, n10245, n10246, n10247, n10248, n10249, n10250,
         n10251, n10252, n10253, n10254, n10255, n10256, n10257, n10258,
         n10259, n10260, n10261, n10262, n10263, n10264, n10265, n10266,
         n10267, n10268, n10269, n10270, n10271, n10272, n10273, n10274,
         n10275, n10276, n10277, n10278, n10279, n10280, n10281, n10282,
         n10283, n10284, n10285, n10286, n10287, n10288, n10290, n10291,
         n10292, n10293, n10294, n10295, n10296, n10297, n10298, n10299,
         n10300, n10301, n10302, n10303, n10304, n10305, n10306, n10307,
         n10308, n10309, n10310, n10311, n10312, n10313, n10314, n10315,
         n10316, n10317, n10318, n10319, n10320, n10321, n10322, n10323,
         n10324, n10325, n10326, n10327, n10328, n10329, n10330, n10331,
         n10332, n10333, n10334, n10335, n10336, n10337, n10338, n10339,
         n10340, n10341, n10342, n10343, n10344, n10345, n10346, n10347,
         n10348, n10349, n10350, n10351, n10352, n10353, n10354, n10355,
         n10356, n10357, n10358, n10359, n10360, n10361, n10362, n10363,
         n10364, n10365, n10366, n10367, n10368, n10369, n10370, n10371,
         n10372, n10373, n10374, n10375, n10376, n10377, n10378, n10379,
         n10380, n10381, n10382, n10383, n10384, n10385, n10386, n10387,
         n10388, n10389, n10390, n10391, n10392, n10393, n10394, n10395,
         n10396, n10397, n10398, n10399, n10400, n10401, n10402, n10403,
         n10404, n10405, n10406, n10407, n10408, n10409, n10410, n10411,
         n10412, n10413, n10414, n10415, n10416, n10417, n10418, n10419,
         n10420, n10421, n10422, n10423, n10424, n10425, n10426, n10427,
         n10428, n10429, n10430, n10431, n10432, n10433, n10434, n10435,
         n10436, n10437, n10438, n10439, n10440, n10441, n10442, n10443,
         n10444, n10445, n10446, n10447, n10448, n10449, n10450, n10451,
         n10452, n10453, n10454, n10455, n10456, n10457, n10458, n10459,
         n10460, n10461, n10462, n10463, n10464, n10465, n10466, n10467,
         n10468, n10469, n10470, n10471, n10472, n10473, n10474, n10475,
         n10476, n10477, n10478, n10479, n10480, n10481, n10482, n10483,
         n10484, n10485, n10486, n10487, n10488, n10489, n10490, n10491,
         n10492, n10493, n10494, n10495, n10496, n10497, n10498, n10499,
         n10500, n10501, n10502, n10503, n10504, n10505, n10506, n10507,
         n10508, n10509, n10510, n10511, n10512, n10513, n10514, n10515,
         n10516, n10517, n10518, n10519, n10520, n10521, n10522, n10523,
         n10524, n10525, n10526, n10527, n10528, n10529, n10530, n10531,
         n10532, n10533, n10534, n10535, n10536, n10537, n10538, n10539,
         n10540, n10541, n10542, n10543, n10544, n10545, n10546, n10547,
         n10548, n10549, n10550, n10551, n10552, n10553, n10554, n10555,
         n10556, n10557, n10558, n10559, n10560, n10561, n10562, n10563,
         n10564, n10565, n10566, n10567, n10568, n10569, n10570, n10571,
         n10572, n10573, n10574, n10575, n10576, n10577, n10578, n10579,
         n10580, n10581, n10582, n10583, n10584, n10585, n10586, n10587,
         n10588, n10589, n10590, n10591, n10592, n10593, n10594, n10595,
         n10596, n10597, n10598, n10599, n10600, n10601, n10602, n10603,
         n10604, n10605, n10606, n10607, n10608, n10609, n10610, n10611,
         n10612, n10613, n10614, n10615, n10616, n10617, n10618, n10619,
         n10620, n10621, n10622, n10623, n10624, n10625, n10626, n10627,
         n10628, n10629, n10630, n10631, n10632, n10633, n10634, n10635,
         n10636, n10637, n10638, n10639, n10640, n10641, n10642, n10643,
         n10644, n10645, n10646, n10647, n10648, n10649, n10650, n10651,
         n10652, n10653, n10654, n10655, n10656, n10657, n10658, n10659;

  NAND2_X1 U4896 ( .A1(n9682), .A2(n5890), .ZN(n9697) );
  AND2_X1 U4897 ( .A1(n5312), .A2(n5311), .ZN(n9699) );
  AND2_X1 U4898 ( .A1(n5326), .A2(n5325), .ZN(n9722) );
  AND2_X1 U4899 ( .A1(n5335), .A2(n5334), .ZN(n10025) );
  INV_X1 U4900 ( .A(n10050), .ZN(n10048) );
  CLKBUF_X3 U4901 ( .A(n7425), .Z(n8592) );
  INV_X2 U4902 ( .A(n8599), .ZN(n8496) );
  NAND2_X4 U4903 ( .A1(n7424), .A2(n7423), .ZN(n8476) );
  BUF_X1 U4904 ( .A(n6705), .Z(n6821) );
  NAND2_X1 U4905 ( .A1(n6511), .A2(n6513), .ZN(n7578) );
  NAND2_X1 U4906 ( .A1(n6507), .A2(n6517), .ZN(n7540) );
  NAND2_X1 U4907 ( .A1(n5913), .A2(n5855), .ZN(n7889) );
  XNOR2_X1 U4908 ( .A(n5945), .B(n5944), .ZN(n6067) );
  INV_X1 U4909 ( .A(n6966), .ZN(n5678) );
  AND2_X1 U4910 ( .A1(n5504), .A2(n5640), .ZN(n4623) );
  NOR2_X1 U4911 ( .A1(P1_IR_REG_12__SCAN_IN), .A2(P1_IR_REG_6__SCAN_IN), .ZN(
        n5253) );
  NOR2_X1 U4912 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(P1_IR_REG_21__SCAN_IN), .ZN(
        n5258) );
  NAND3_X1 U4913 ( .A1(n9635), .A2(n4706), .A3(n4705), .ZN(n4883) );
  NAND2_X1 U4914 ( .A1(n5346), .A2(n10042), .ZN(n5991) );
  BUF_X1 U4915 ( .A(n5612), .Z(n5716) );
  NAND3_X1 U4916 ( .A1(n4882), .A2(P1_ADDR_REG_19__SCAN_IN), .A3(
        P2_ADDR_REG_19__SCAN_IN), .ZN(n4881) );
  AND2_X1 U4918 ( .A1(n6136), .A2(n6122), .ZN(n6199) );
  OR2_X1 U4919 ( .A1(n8930), .A2(n9003), .ZN(n8978) );
  NAND2_X1 U4920 ( .A1(n8427), .A2(n5783), .ZN(n10050) );
  AND2_X1 U4921 ( .A1(n5973), .A2(n5974), .ZN(n8139) );
  NAND2_X1 U4922 ( .A1(n9733), .A2(n7806), .ZN(n6951) );
  AND3_X1 U4923 ( .A1(n5597), .A2(n5596), .A3(n5595), .ZN(n7979) );
  OR2_X1 U4924 ( .A1(n5269), .A2(P1_IR_REG_28__SCAN_IN), .ZN(n5268) );
  INV_X1 U4925 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n5640) );
  AND4_X1 U4926 ( .A1(n6254), .A2(n6253), .A3(n6252), .A4(n6251), .ZN(n8115)
         );
  AND4_X1 U4927 ( .A1(n6144), .A2(n6143), .A3(n6142), .A4(n6141), .ZN(n7325)
         );
  NAND2_X1 U4928 ( .A1(n6640), .A2(n6639), .ZN(n8290) );
  AND3_X1 U4929 ( .A1(n4523), .A2(n9645), .A3(n10418), .ZN(n10174) );
  AND2_X1 U4930 ( .A1(n5272), .A2(n5271), .ZN(n5289) );
  NOR2_X1 U4931 ( .A1(n5594), .A2(n5456), .ZN(n7284) );
  AOI21_X1 U4932 ( .B1(n9099), .B2(n9098), .A(n4507), .ZN(n9083) );
  AND2_X2 U4933 ( .A1(n7601), .A2(n7603), .ZN(n4441) );
  AND2_X2 U4934 ( .A1(n6859), .A2(n6858), .ZN(n6871) );
  NOR2_X2 U4935 ( .A1(P2_IR_REG_7__SCAN_IN), .A2(P2_IR_REG_14__SCAN_IN), .ZN(
        n6091) );
  OAI21_X2 U4936 ( .B1(n8923), .B2(n4854), .A(n4852), .ZN(n8954) );
  NOR2_X2 U4937 ( .A1(P2_IR_REG_16__SCAN_IN), .A2(P2_IR_REG_13__SCAN_IN), .ZN(
        n6090) );
  OR2_X1 U4938 ( .A1(n5484), .A2(n5483), .ZN(n4893) );
  OAI21_X2 U4939 ( .B1(n6463), .B2(n5073), .A(n5072), .ZN(n6477) );
  NAND2_X2 U4940 ( .A1(n8961), .A2(n6449), .ZN(n6463) );
  BUF_X1 U4941 ( .A(n7946), .Z(n4391) );
  NAND2_X2 U4942 ( .A1(n6110), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5065) );
  NAND2_X2 U4943 ( .A1(n5390), .A2(n5389), .ZN(n10114) );
  NAND2_X2 U4944 ( .A1(n6429), .A2(n6428), .ZN(n9268) );
  NAND2_X2 U4945 ( .A1(n5490), .A2(n5489), .ZN(n8329) );
  NAND2_X2 U4946 ( .A1(n7611), .A2(n6718), .ZN(n7603) );
  NAND2_X2 U4947 ( .A1(n5283), .A2(n5282), .ZN(n8619) );
  OR2_X1 U4948 ( .A1(n6697), .A2(n6624), .ZN(n6696) );
  XNOR2_X2 U4949 ( .A(n4997), .B(P2_IR_REG_22__SCAN_IN), .ZN(n6624) );
  BUF_X4 U4950 ( .A(n6192), .Z(n6351) );
  NAND2_X1 U4951 ( .A1(n6047), .A2(n9697), .ZN(n9709) );
  NAND2_X1 U4952 ( .A1(n9088), .A2(n9087), .ZN(n9090) );
  NAND2_X1 U4953 ( .A1(n8194), .A2(n4419), .ZN(n8318) );
  NAND2_X1 U4954 ( .A1(n7750), .A2(n5002), .ZN(n7931) );
  INV_X1 U4955 ( .A(n9117), .ZN(n9307) );
  INV_X1 U4956 ( .A(n9184), .ZN(n5064) );
  NAND2_X1 U4957 ( .A1(n10401), .A2(n6013), .ZN(n5744) );
  NAND2_X1 U4958 ( .A1(n7946), .A2(n9589), .ZN(n5863) );
  INV_X1 U4959 ( .A(n8837), .ZN(n7988) );
  NAND2_X1 U4960 ( .A1(n8843), .A2(n10524), .ZN(n6517) );
  NAND2_X2 U4961 ( .A1(n7498), .A2(n7423), .ZN(n7865) );
  OR2_X1 U4962 ( .A1(n7360), .A2(n4910), .ZN(n7424) );
  INV_X2 U4963 ( .A(n6455), .ZN(n6469) );
  XNOR2_X1 U4964 ( .A(n7671), .B(n6705), .ZN(n6703) );
  INV_X1 U4965 ( .A(n6161), .ZN(n6411) );
  NAND2_X1 U4966 ( .A1(n6134), .A2(n4678), .ZN(n6161) );
  CLKBUF_X2 U4967 ( .A(n6199), .Z(n6437) );
  CLKBUF_X1 U4968 ( .A(n6196), .Z(n6464) );
  INV_X1 U4969 ( .A(n6136), .ZN(n4678) );
  CLKBUF_X2 U4970 ( .A(n6698), .Z(n4396) );
  INV_X1 U4971 ( .A(n6697), .ZN(n8533) );
  NAND3_X1 U4972 ( .A1(n4922), .A2(n4921), .A3(n5570), .ZN(n5730) );
  INV_X1 U4973 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n4918) );
  INV_X1 U4974 ( .A(P1_RD_REG_SCAN_IN), .ZN(n4705) );
  INV_X2 U4975 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3152) );
  AND2_X2 U4976 ( .A1(n5052), .A2(n5050), .ZN(n8644) );
  AOI21_X1 U4977 ( .B1(n5806), .B2(n4763), .A(n4762), .ZN(n4761) );
  NAND2_X1 U4978 ( .A1(n9489), .A2(n8577), .ZN(n9457) );
  NAND2_X1 U4979 ( .A1(n9709), .A2(n6048), .ZN(n9678) );
  NOR2_X2 U4980 ( .A1(n9020), .A2(n9268), .ZN(n9007) );
  NAND2_X1 U4981 ( .A1(n6780), .A2(n6779), .ZN(n8717) );
  OR2_X1 U4982 ( .A1(n8926), .A2(n9051), .ZN(n5105) );
  AND2_X1 U4983 ( .A1(n9052), .A2(n9044), .ZN(n9051) );
  NAND2_X1 U4984 ( .A1(n6593), .A2(n6583), .ZN(n9044) );
  NAND2_X1 U4985 ( .A1(n6397), .A2(n6396), .ZN(n9286) );
  NAND2_X1 U4986 ( .A1(n5350), .A2(n5349), .ZN(n10201) );
  NAND2_X1 U4987 ( .A1(n5304), .A2(n5303), .ZN(n9690) );
  XNOR2_X1 U4988 ( .A(n5281), .B(n5280), .ZN(n10288) );
  NAND2_X1 U4989 ( .A1(n6419), .A2(n6418), .ZN(n9275) );
  NAND2_X1 U4990 ( .A1(n6386), .A2(n6385), .ZN(n9291) );
  NAND2_X1 U4991 ( .A1(n5316), .A2(n5315), .ZN(n10190) );
  NAND2_X1 U4992 ( .A1(n5338), .A2(n5337), .ZN(n5346) );
  NOR2_X1 U4993 ( .A1(n9307), .A2(n9312), .ZN(n4991) );
  OR2_X1 U4994 ( .A1(n10114), .A2(n10133), .ZN(n10087) );
  XNOR2_X1 U4995 ( .A(n5293), .B(n5294), .ZN(n8420) );
  AOI21_X1 U4996 ( .B1(n4975), .B2(n4971), .A(n4974), .ZN(n4970) );
  XNOR2_X1 U4997 ( .A(n4606), .B(n5336), .ZN(n7993) );
  NAND2_X1 U4998 ( .A1(n8293), .A2(n8292), .ZN(n8295) );
  AND2_X1 U4999 ( .A1(n6562), .A2(n6347), .ZN(n6348) );
  NAND2_X1 U5000 ( .A1(n5362), .A2(n5361), .ZN(n10061) );
  AOI21_X1 U5001 ( .B1(n5069), .B2(n5071), .A(n5067), .ZN(n4506) );
  OR2_X1 U5002 ( .A1(n4840), .A2(n8112), .ZN(n4837) );
  NAND2_X1 U5003 ( .A1(n5417), .A2(n5416), .ZN(n10226) );
  AND2_X1 U5004 ( .A1(n9142), .A2(n6554), .ZN(n9184) );
  NAND2_X1 U5005 ( .A1(n5429), .A2(n5428), .ZN(n10230) );
  NAND2_X1 U5006 ( .A1(n6312), .A2(n6311), .ZN(n9327) );
  NAND2_X1 U5007 ( .A1(n4886), .A2(n5180), .ZN(n5414) );
  NAND2_X1 U5008 ( .A1(n4627), .A2(n4753), .ZN(n7963) );
  NAND2_X1 U5009 ( .A1(n5476), .A2(n5475), .ZN(n8287) );
  OAI211_X1 U5010 ( .C1(n5744), .C2(n4810), .A(n4808), .B(n5964), .ZN(n5967)
         );
  NAND2_X1 U5011 ( .A1(n6295), .A2(n6294), .ZN(n9342) );
  NAND2_X2 U5012 ( .A1(n4546), .A2(n6259), .ZN(n9347) );
  NAND2_X1 U5013 ( .A1(n6538), .A2(n8089), .ZN(n8047) );
  NAND2_X1 U5014 ( .A1(n5521), .A2(n5520), .ZN(n10239) );
  NAND2_X1 U5015 ( .A1(n5509), .A2(n5508), .ZN(n8066) );
  AND2_X1 U5016 ( .A1(n6228), .A2(n8043), .ZN(n6924) );
  OR2_X1 U5017 ( .A1(n10475), .A2(n8008), .ZN(n7900) );
  INV_X2 U5018 ( .A(n9060), .ZN(n4392) );
  AND2_X1 U5019 ( .A1(n6528), .A2(n6527), .ZN(n7817) );
  AND2_X1 U5020 ( .A1(n6013), .A2(n6012), .ZN(n10415) );
  NAND2_X1 U5021 ( .A1(n4758), .A2(n4756), .ZN(n5913) );
  NAND2_X1 U5022 ( .A1(n7348), .A2(n5739), .ZN(n4785) );
  NAND2_X1 U5023 ( .A1(n4760), .A2(n4759), .ZN(n7894) );
  AND2_X2 U5024 ( .A1(n6965), .A2(P1_STATE_REG_SCAN_IN), .ZN(P1_U4006) );
  NAND2_X2 U5025 ( .A1(n7425), .A2(n6952), .ZN(n8599) );
  NAND2_X1 U5026 ( .A1(n7795), .A2(n5738), .ZN(n7348) );
  INV_X1 U5027 ( .A(n7850), .ZN(n4756) );
  AND3_X1 U5028 ( .A1(n6166), .A2(n6164), .A3(n4543), .ZN(n7715) );
  NAND2_X1 U5029 ( .A1(n6720), .A2(n8763), .ZN(n7600) );
  NAND2_X1 U5030 ( .A1(n4430), .A2(n4402), .ZN(n8844) );
  NAND4_X2 U5031 ( .A1(n6191), .A2(n6190), .A3(n6189), .A4(n6188), .ZN(n8840)
         );
  CLKBUF_X1 U5032 ( .A(n7498), .Z(n4520) );
  NAND2_X2 U5033 ( .A1(n7498), .A2(n6953), .ZN(n8593) );
  AND4_X1 U5034 ( .A1(n6151), .A2(n6150), .A3(n6149), .A4(n6148), .ZN(n7580)
         );
  INV_X1 U5035 ( .A(n6941), .ZN(n8800) );
  AND2_X1 U5036 ( .A1(n4911), .A2(n7367), .ZN(n7360) );
  AND2_X1 U5037 ( .A1(n4980), .A2(n4979), .ZN(n6941) );
  NAND2_X2 U5038 ( .A1(n6657), .A2(n4995), .ZN(n6812) );
  NAND2_X1 U5039 ( .A1(n6133), .A2(n6132), .ZN(n7671) );
  BUF_X4 U5040 ( .A(n6187), .Z(n6452) );
  AND2_X2 U5041 ( .A1(n6134), .A2(n6136), .ZN(n6175) );
  NAND2_X1 U5042 ( .A1(n5948), .A2(n5949), .ZN(n8405) );
  AND2_X2 U5043 ( .A1(n6122), .A2(n8642), .ZN(n6187) );
  NAND2_X1 U5044 ( .A1(n5949), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5945) );
  XNOR2_X1 U5045 ( .A(n5833), .B(n5832), .ZN(n7806) );
  AND2_X1 U5046 ( .A1(n5142), .A2(n5136), .ZN(n4896) );
  INV_X1 U5047 ( .A(n6131), .ZN(n6192) );
  AND3_X2 U5048 ( .A1(n5942), .A2(n5736), .A3(n5735), .ZN(n6950) );
  NOR2_X1 U5049 ( .A1(n4440), .A2(n4885), .ZN(n4884) );
  INV_X1 U5050 ( .A(n6136), .ZN(n8642) );
  INV_X1 U5051 ( .A(n6122), .ZN(n6134) );
  BUF_X2 U5052 ( .A(n5617), .Z(n10290) );
  INV_X2 U5053 ( .A(n4397), .ZN(n4394) );
  NAND2_X1 U5054 ( .A1(n4914), .A2(n4913), .ZN(n5404) );
  CLKBUF_X1 U5055 ( .A(n6110), .Z(n9385) );
  MUX2_X1 U5056 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5262), .S(
        P1_IR_REG_28__SCAN_IN), .Z(n5263) );
  XNOR2_X1 U5057 ( .A(n6496), .B(n6495), .ZN(n6698) );
  NAND2_X1 U5058 ( .A1(n5721), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5415) );
  NAND2_X1 U5059 ( .A1(n6494), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6496) );
  NAND2_X1 U5060 ( .A1(n6668), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4997) );
  NAND2_X1 U5061 ( .A1(n4537), .A2(n4536), .ZN(n5942) );
  OR2_X1 U5062 ( .A1(n5273), .A2(n4918), .ZN(n5275) );
  NAND2_X2 U5063 ( .A1(n4545), .A2(P1_U3084), .ZN(n10294) );
  NAND2_X1 U5064 ( .A1(n4621), .A2(n4620), .ZN(n5269) );
  NAND2_X1 U5065 ( .A1(n6488), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6493) );
  NAND4_X1 U5066 ( .A1(n4618), .A2(n4619), .A3(n4435), .A4(n4405), .ZN(n4625)
         );
  AOI21_X1 U5067 ( .B1(n4916), .B2(n4918), .A(n4918), .ZN(n4913) );
  INV_X1 U5068 ( .A(n6119), .ZN(n6490) );
  AND4_X2 U5069 ( .A1(n5251), .A2(n5252), .A3(n5255), .A4(n5458), .ZN(n4617)
         );
  NAND2_X1 U5070 ( .A1(n6495), .A2(n6492), .ZN(n6119) );
  AND4_X1 U5071 ( .A1(n6666), .A2(n6118), .A3(n6489), .A4(n6098), .ZN(n5092)
         );
  AND2_X1 U5072 ( .A1(n4624), .A2(n5568), .ZN(n4619) );
  INV_X1 U5073 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n5458) );
  INV_X1 U5074 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n5504) );
  INV_X1 U5075 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n5274) );
  NOR2_X1 U5076 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(P1_IR_REG_11__SCAN_IN), .ZN(
        n4624) );
  INV_X1 U5077 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n5946) );
  INV_X1 U5078 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n4706) );
  INV_X1 U5079 ( .A(P2_RD_REG_SCAN_IN), .ZN(n4882) );
  INV_X1 U5080 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n6269) );
  INV_X1 U5081 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n6666) );
  INV_X1 U5082 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n6495) );
  INV_X1 U5083 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n6098) );
  NOR2_X1 U5084 ( .A1(P2_IR_REG_12__SCAN_IN), .A2(P2_IR_REG_11__SCAN_IN), .ZN(
        n6092) );
  INV_X1 U5085 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n6329) );
  AOI21_X1 U5086 ( .B1(n9384), .B2(n5591), .A(n5096), .ZN(n10248) );
  NAND2_X2 U5087 ( .A1(n7746), .A2(n6743), .ZN(n7750) );
  AND2_X2 U5088 ( .A1(n8220), .A2(n9423), .ZN(n8221) );
  NAND3_X1 U5089 ( .A1(n6171), .A2(n6097), .A3(n5031), .ZN(n6488) );
  AND2_X4 U5090 ( .A1(n6168), .A2(n6089), .ZN(n6171) );
  AND2_X2 U5091 ( .A1(n6145), .A2(n6088), .ZN(n6168) );
  INV_X2 U5092 ( .A(n7802), .ZN(n6054) );
  OAI222_X1 U5093 ( .A1(n10317), .A2(P1_U3084), .B1(n10283), .B2(n7029), .C1(
        n7028), .C2(n10294), .ZN(P1_U3352) );
  OAI222_X1 U5094 ( .A1(n9395), .A2(n5620), .B1(n9399), .B2(n7029), .C1(
        P2_U3152), .C2(n7272), .ZN(P2_U3357) );
  OAI21_X2 U5095 ( .B1(n8644), .B2(n6827), .A(n8643), .ZN(n8648) );
  INV_X1 U5096 ( .A(n6812), .ZN(n4395) );
  NAND2_X2 U5097 ( .A1(n6673), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6683) );
  NAND2_X1 U5098 ( .A1(n4510), .A2(n4509), .ZN(n4754) );
  NAND2_X1 U5099 ( .A1(n7963), .A2(n6950), .ZN(n4626) );
  OR2_X1 U5100 ( .A1(n9275), .A2(n9036), .ZN(n6595) );
  NAND2_X1 U5101 ( .A1(n5196), .A2(n9816), .ZN(n5199) );
  INV_X1 U5102 ( .A(SI_10_), .ZN(n5145) );
  OR2_X1 U5103 ( .A1(n9278), .A2(n9049), .ZN(n8927) );
  OR2_X1 U5104 ( .A1(n9261), .A2(n8928), .ZN(n8962) );
  AND2_X1 U5105 ( .A1(n6949), .A2(n6950), .ZN(n7367) );
  INV_X1 U5106 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n5250) );
  NAND2_X1 U5107 ( .A1(n4605), .A2(n4887), .ZN(n5439) );
  AND2_X1 U5108 ( .A1(n4888), .A2(n5169), .ZN(n4887) );
  OAI21_X1 U5109 ( .B1(n6518), .B2(n4394), .A(n4828), .ZN(n6519) );
  NAND2_X1 U5110 ( .A1(n6506), .A2(n4394), .ZN(n4828) );
  NAND2_X1 U5111 ( .A1(n5747), .A2(n4766), .ZN(n4765) );
  NOR2_X1 U5112 ( .A1(n4767), .A2(n7994), .ZN(n4766) );
  INV_X1 U5113 ( .A(n5851), .ZN(n4767) );
  AOI21_X1 U5114 ( .B1(n5771), .B2(n5770), .A(n5769), .ZN(n5775) );
  NOR2_X1 U5115 ( .A1(n4976), .A2(n5085), .ZN(n4975) );
  INV_X1 U5116 ( .A(n8439), .ZN(n4976) );
  AND2_X1 U5117 ( .A1(n5399), .A2(n5193), .ZN(n5194) );
  NAND2_X1 U5118 ( .A1(n4884), .A2(n4600), .ZN(n4599) );
  INV_X1 U5119 ( .A(n4884), .ZN(n4601) );
  INV_X1 U5120 ( .A(n5385), .ZN(n5182) );
  INV_X1 U5121 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n5175) );
  INV_X1 U5122 ( .A(n5058), .ZN(n5057) );
  OAI21_X1 U5123 ( .B1(n6818), .B2(n5061), .A(n5060), .ZN(n5058) );
  AND2_X1 U5124 ( .A1(n6818), .A2(n5061), .ZN(n5055) );
  OR2_X1 U5125 ( .A1(n7308), .A2(n4417), .ZN(n4657) );
  INV_X1 U5126 ( .A(n7331), .ZN(n4656) );
  NOR2_X1 U5127 ( .A1(n6230), .A2(P2_IR_REG_8__SCAN_IN), .ZN(n6271) );
  AOI21_X1 U5128 ( .B1(n4655), .B2(n4653), .A(n4651), .ZN(n4650) );
  INV_X1 U5129 ( .A(n7474), .ZN(n4651) );
  INV_X1 U5130 ( .A(n4653), .ZN(n4652) );
  OR2_X1 U5131 ( .A1(n9245), .A2(n8969), .ZN(n6612) );
  NAND2_X1 U5132 ( .A1(n4991), .A2(n4990), .ZN(n4989) );
  NOR2_X1 U5133 ( .A1(n4668), .A2(n4667), .ZN(n4666) );
  NAND2_X1 U5134 ( .A1(n6552), .A2(n6632), .ZN(n4668) );
  OR2_X1 U5135 ( .A1(n9347), .A2(n8088), .ZN(n6640) );
  NAND2_X1 U5136 ( .A1(n6589), .A2(n6595), .ZN(n8953) );
  AOI21_X1 U5137 ( .B1(n4672), .B2(n4674), .A(n4671), .ZN(n4670) );
  INV_X1 U5138 ( .A(n6595), .ZN(n4671) );
  NAND2_X1 U5139 ( .A1(n9500), .A2(n4945), .ZN(n4944) );
  OAI21_X1 U5140 ( .B1(n4948), .B2(n4950), .A(n4947), .ZN(n4945) );
  INV_X1 U5141 ( .A(n4954), .ZN(n4947) );
  INV_X1 U5142 ( .A(n4953), .ZN(n4948) );
  INV_X1 U5143 ( .A(n8476), .ZN(n8563) );
  NOR2_X1 U5144 ( .A1(n5085), .A2(n4973), .ZN(n4969) );
  INV_X1 U5145 ( .A(n8440), .ZN(n4973) );
  INV_X1 U5146 ( .A(n8629), .ZN(n5288) );
  OR2_X1 U5147 ( .A1(n10061), .A2(n10074), .ZN(n8427) );
  AOI21_X1 U5148 ( .B1(n5020), .B2(n4449), .A(n6036), .ZN(n4687) );
  OR2_X1 U5149 ( .A1(n10075), .A2(n10091), .ZN(n8426) );
  NOR2_X1 U5150 ( .A1(n10230), .A2(n8454), .ZN(n4909) );
  NAND2_X1 U5151 ( .A1(n4809), .A2(n5855), .ZN(n4808) );
  AOI22_X1 U5152 ( .A1(n6949), .A2(n4911), .B1(n6950), .B2(n9733), .ZN(n4910)
         );
  AND2_X1 U5153 ( .A1(n6966), .A2(n4545), .ZN(n5567) );
  NOR2_X1 U5154 ( .A1(n9590), .A2(n7794), .ZN(n7796) );
  NAND2_X1 U5155 ( .A1(n7796), .A2(n4784), .ZN(n7795) );
  OR3_X2 U5156 ( .A1(n6067), .A2(n8405), .A3(n8334), .ZN(n7498) );
  INV_X1 U5157 ( .A(n4732), .ZN(n4731) );
  AOI21_X1 U5158 ( .B1(n4732), .B2(n4734), .A(SI_29_), .ZN(n4730) );
  NOR2_X1 U5159 ( .A1(n5729), .A2(n5254), .ZN(n4620) );
  INV_X1 U5160 ( .A(n4625), .ZN(n4621) );
  NAND2_X1 U5161 ( .A1(n4720), .A2(n4718), .ZN(n5328) );
  AND2_X1 U5162 ( .A1(n4719), .A2(n4724), .ZN(n4718) );
  AOI21_X1 U5163 ( .B1(n5347), .B2(n4726), .A(n4725), .ZN(n4724) );
  INV_X1 U5164 ( .A(n5729), .ZN(n4536) );
  INV_X1 U5165 ( .A(n5730), .ZN(n4537) );
  INV_X1 U5166 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n5387) );
  INV_X1 U5167 ( .A(n5441), .ZN(n5388) );
  NAND2_X1 U5168 ( .A1(n5426), .A2(n5100), .ZN(n4886) );
  NAND2_X1 U5169 ( .A1(n5153), .A2(n5152), .ZN(n5517) );
  NOR2_X1 U5170 ( .A1(n5503), .A2(P1_IR_REG_10__SCAN_IN), .ZN(n5518) );
  INV_X1 U5171 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n5457) );
  OR2_X1 U5172 ( .A1(n6287), .A2(n9890), .ZN(n6340) );
  OR2_X1 U5173 ( .A1(n6862), .A2(n10530), .ZN(n6860) );
  AND2_X1 U5174 ( .A1(n6448), .A2(n6447), .ZN(n8928) );
  OR2_X1 U5175 ( .A1(n8984), .A2(n6467), .ZN(n6448) );
  OR2_X1 U5176 ( .A1(n6679), .A2(n8256), .ZN(n7099) );
  INV_X1 U5177 ( .A(n6437), .ZN(n6467) );
  NAND2_X1 U5178 ( .A1(n6105), .A2(n6104), .ZN(n8901) );
  AOI21_X1 U5179 ( .B1(n4855), .B2(n4860), .A(n4853), .ZN(n4852) );
  INV_X1 U5180 ( .A(n4855), .ZN(n4854) );
  INV_X1 U5181 ( .A(n8927), .ZN(n4853) );
  OAI21_X1 U5182 ( .B1(n9076), .B2(n9086), .A(n9083), .ZN(n8923) );
  AND2_X1 U5183 ( .A1(n4858), .A2(n4856), .ZN(n4855) );
  OR2_X1 U5184 ( .A1(n9317), .A2(n9175), .ZN(n8916) );
  NAND2_X1 U5185 ( .A1(n4848), .A2(n4416), .ZN(n4847) );
  NOR2_X1 U5186 ( .A1(n6100), .A2(P2_IR_REG_28__SCAN_IN), .ZN(n6101) );
  NAND2_X1 U5187 ( .A1(n8954), .A2(n8953), .ZN(n9000) );
  NAND2_X1 U5188 ( .A1(n6657), .A2(n4396), .ZN(n10590) );
  AND2_X1 U5189 ( .A1(n6111), .A2(n5098), .ZN(n5066) );
  INV_X1 U5190 ( .A(n7367), .ZN(n6904) );
  INV_X1 U5191 ( .A(n5705), .ZN(n5434) );
  INV_X1 U5192 ( .A(n5715), .ZN(n5422) );
  NAND2_X1 U5193 ( .A1(n5305), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n5307) );
  AND2_X1 U5194 ( .A1(n9540), .A2(n4930), .ZN(n4929) );
  AOI21_X1 U5195 ( .B1(n5899), .B2(n5900), .A(n5937), .ZN(n5901) );
  NOR2_X1 U5196 ( .A1(n5937), .A2(n4707), .ZN(n5728) );
  AND2_X1 U5197 ( .A1(n6875), .A2(n4459), .ZN(n4708) );
  AND2_X1 U5198 ( .A1(n5289), .A2(n8629), .ZN(n5611) );
  AOI21_X1 U5199 ( .B1(n9678), .B2(n5029), .A(n5027), .ZN(n6873) );
  NOR2_X1 U5200 ( .A1(n5695), .A2(n5030), .ZN(n5029) );
  INV_X1 U5201 ( .A(n6050), .ZN(n5030) );
  OR2_X1 U5202 ( .A1(n8450), .A2(n8441), .ZN(n8338) );
  OR2_X1 U5203 ( .A1(n6904), .A2(n10290), .ZN(n10403) );
  INV_X1 U5204 ( .A(n10403), .ZN(n10103) );
  OR2_X1 U5205 ( .A1(n6904), .A2(n7366), .ZN(n10405) );
  NAND2_X1 U5206 ( .A1(n6873), .A2(n4786), .ZN(n9653) );
  INV_X1 U5207 ( .A(n6902), .ZN(n7497) );
  NAND2_X1 U5208 ( .A1(n4593), .A2(n4591), .ZN(n9651) );
  INV_X1 U5209 ( .A(n4592), .ZN(n4591) );
  NAND2_X1 U5210 ( .A1(n4594), .A2(n10101), .ZN(n4593) );
  OAI22_X1 U5211 ( .A1(n9671), .A2(n10403), .B1(n9639), .B2(n6002), .ZN(n4592)
         );
  AND3_X1 U5212 ( .A1(n4827), .A2(n4826), .A3(n6160), .ZN(n6516) );
  NAND2_X1 U5213 ( .A1(n6504), .A2(n6505), .ZN(n4826) );
  AOI21_X1 U5214 ( .B1(n5763), .B2(n5856), .A(n4781), .ZN(n4780) );
  INV_X1 U5215 ( .A(n8338), .ZN(n4781) );
  NOR2_X1 U5216 ( .A1(n4805), .A2(n4397), .ZN(n4804) );
  INV_X1 U5217 ( .A(n6632), .ZN(n4805) );
  OAI21_X1 U5218 ( .B1(n4806), .B2(n6546), .A(n4802), .ZN(n4801) );
  AND2_X1 U5219 ( .A1(n8298), .A2(n4397), .ZN(n4802) );
  NAND2_X1 U5220 ( .A1(n4629), .A2(n5755), .ZN(n5761) );
  AOI21_X1 U5221 ( .B1(n4780), .B2(n5978), .A(n4776), .ZN(n4775) );
  INV_X1 U5222 ( .A(n5850), .ZN(n4776) );
  AOI21_X1 U5223 ( .B1(n5758), .B2(n5759), .A(n4457), .ZN(n4778) );
  AOI21_X1 U5224 ( .B1(n4775), .B2(n4777), .A(n7994), .ZN(n4773) );
  INV_X1 U5225 ( .A(n4780), .ZN(n4777) );
  NOR2_X1 U5226 ( .A1(n4800), .A2(n4797), .ZN(n6557) );
  NAND2_X1 U5227 ( .A1(n4799), .A2(n4798), .ZN(n4797) );
  AND3_X1 U5228 ( .A1(n4801), .A2(n4803), .A3(n8299), .ZN(n4800) );
  INV_X1 U5229 ( .A(n6550), .ZN(n4799) );
  NOR2_X1 U5230 ( .A1(n10226), .A2(n7994), .ZN(n4751) );
  AOI21_X1 U5231 ( .B1(n5775), .B2(n5774), .A(n5773), .ZN(n5786) );
  AOI21_X1 U5232 ( .B1(n6570), .B2(n4817), .A(n6582), .ZN(n4816) );
  NOR2_X1 U5233 ( .A1(n4819), .A2(n4818), .ZN(n4817) );
  NAND2_X1 U5234 ( .A1(n5781), .A2(n4752), .ZN(n5782) );
  AND2_X1 U5235 ( .A1(n10087), .A2(n10107), .ZN(n4752) );
  AND2_X1 U5236 ( .A1(n8980), .A2(n6600), .ZN(n4796) );
  INV_X1 U5237 ( .A(n6611), .ZN(n5075) );
  NOR2_X1 U5238 ( .A1(n5960), .A2(n5961), .ZN(n5963) );
  OR2_X1 U5239 ( .A1(n6597), .A2(n4397), .ZN(n4513) );
  AND2_X1 U5240 ( .A1(n4512), .A2(n4791), .ZN(n4511) );
  NAND2_X1 U5241 ( .A1(n4957), .A2(n8566), .ZN(n4954) );
  INV_X1 U5242 ( .A(n8523), .ZN(n4950) );
  NAND2_X1 U5243 ( .A1(n4942), .A2(n8486), .ZN(n4941) );
  INV_X1 U5244 ( .A(n8472), .ZN(n4942) );
  NOR2_X1 U5245 ( .A1(n4406), .A2(n9683), .ZN(n4764) );
  NAND2_X1 U5246 ( .A1(n4538), .A2(n9682), .ZN(n5806) );
  NAND2_X1 U5247 ( .A1(n5816), .A2(n4539), .ZN(n4538) );
  NOR2_X1 U5248 ( .A1(n4445), .A2(n4540), .ZN(n4539) );
  NOR2_X1 U5249 ( .A1(n5805), .A2(n5923), .ZN(n4540) );
  AND2_X1 U5250 ( .A1(n10230), .A2(n10132), .ZN(n5848) );
  NOR2_X1 U5251 ( .A1(n4823), .A2(n4604), .ZN(n4603) );
  INV_X1 U5252 ( .A(n5988), .ZN(n4821) );
  INV_X1 U5253 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n5259) );
  NAND2_X1 U5254 ( .A1(n5177), .A2(n5176), .ZN(n5180) );
  AND2_X1 U5255 ( .A1(n4895), .A2(n5099), .ZN(n4894) );
  NAND2_X1 U5256 ( .A1(n5483), .A2(n5161), .ZN(n4895) );
  NOR2_X1 U5257 ( .A1(n5648), .A2(n5121), .ZN(n5126) );
  NOR2_X1 U5258 ( .A1(n6365), .A2(n6364), .ZN(n4526) );
  INV_X1 U5259 ( .A(n6787), .ZN(n5036) );
  OR2_X1 U5260 ( .A1(n8735), .A2(n5035), .ZN(n5034) );
  NAND2_X1 U5261 ( .A1(n8720), .A2(n6787), .ZN(n5035) );
  INV_X1 U5262 ( .A(n7598), .ZN(n6716) );
  INV_X1 U5263 ( .A(n6990), .ZN(n6714) );
  BUF_X1 U5264 ( .A(n6754), .Z(n6829) );
  NOR2_X1 U5265 ( .A1(n6409), .A2(n8749), .ZN(n4527) );
  AND2_X1 U5266 ( .A1(n9027), .A2(n6583), .ZN(n5079) );
  AND2_X1 U5267 ( .A1(n4401), .A2(n8919), .ZN(n4830) );
  OR2_X1 U5268 ( .A1(n9327), .A2(n9206), .ZN(n9142) );
  AND2_X1 U5269 ( .A1(n6305), .A2(n6551), .ZN(n6306) );
  OR2_X1 U5270 ( .A1(n8911), .A2(n9204), .ZN(n6548) );
  NOR2_X1 U5271 ( .A1(n4985), .A2(n9347), .ZN(n4984) );
  NAND2_X1 U5272 ( .A1(n6248), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n6261) );
  NAND2_X1 U5273 ( .A1(n7816), .A2(n5078), .ZN(n6927) );
  AND2_X1 U5274 ( .A1(n6229), .A2(n6527), .ZN(n5078) );
  INV_X1 U5275 ( .A(n6637), .ZN(n4662) );
  NAND2_X1 U5276 ( .A1(n10575), .A2(n8841), .ZN(n6636) );
  AND2_X1 U5277 ( .A1(n6637), .A2(n6636), .ZN(n7711) );
  NAND2_X1 U5278 ( .A1(n6625), .A2(n6624), .ZN(n6929) );
  NOR2_X1 U5279 ( .A1(n9028), .A2(n9275), .ZN(n8633) );
  AOI21_X1 U5280 ( .B1(n10531), .B2(n6837), .A(n6836), .ZN(n7533) );
  INV_X1 U5281 ( .A(n8417), .ZN(n6832) );
  AND2_X1 U5282 ( .A1(n6099), .A2(n6677), .ZN(n5081) );
  BUF_X1 U5283 ( .A(n6097), .Z(n4541) );
  OR2_X1 U5284 ( .A1(n6271), .A2(n6170), .ZN(n6242) );
  OR2_X1 U5285 ( .A1(n6224), .A2(n6223), .ZN(n6230) );
  INV_X2 U5286 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n6222) );
  INV_X1 U5287 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n6089) );
  AND2_X1 U5288 ( .A1(n6949), .A2(n7806), .ZN(n6953) );
  NAND2_X1 U5289 ( .A1(n8513), .A2(n4448), .ZN(n4951) );
  NOR2_X1 U5290 ( .A1(n8514), .A2(n4959), .ZN(n4953) );
  AND2_X1 U5291 ( .A1(n9605), .A2(n10334), .ZN(n9607) );
  OR2_X1 U5292 ( .A1(n10329), .A2(n9607), .ZN(n9609) );
  NOR2_X1 U5293 ( .A1(n9623), .A2(n10234), .ZN(n4569) );
  INV_X1 U5294 ( .A(SI_20_), .ZN(n9816) );
  NAND2_X1 U5295 ( .A1(n10114), .A2(n10133), .ZN(n5776) );
  OR2_X1 U5296 ( .A1(n10226), .A2(n10156), .ZN(n5987) );
  INV_X1 U5297 ( .A(n5848), .ZN(n5983) );
  OR2_X1 U5298 ( .A1(n8066), .A2(n8207), .ZN(n8033) );
  INV_X1 U5299 ( .A(n7889), .ZN(n4807) );
  INV_X1 U5300 ( .A(n7921), .ZN(n4906) );
  INV_X1 U5301 ( .A(n6043), .ZN(n5014) );
  INV_X1 U5302 ( .A(n5005), .ZN(n5004) );
  INV_X1 U5303 ( .A(n5260), .ZN(n4618) );
  AND2_X1 U5304 ( .A1(n5229), .A2(n5228), .ZN(n5301) );
  OAI21_X1 U5305 ( .B1(n5328), .B2(n5220), .A(n5219), .ZN(n5314) );
  NOR2_X1 U5306 ( .A1(n5336), .A2(n4722), .ZN(n4721) );
  INV_X1 U5307 ( .A(n5204), .ZN(n4722) );
  NAND2_X1 U5308 ( .A1(n4607), .A2(n5360), .ZN(n4723) );
  AND2_X1 U5309 ( .A1(n5725), .A2(n5832), .ZN(n4912) );
  AOI21_X1 U5310 ( .B1(n4428), .B2(n4601), .A(n4598), .ZN(n4597) );
  INV_X1 U5311 ( .A(n5195), .ZN(n4598) );
  INV_X1 U5312 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n5723) );
  NAND2_X1 U5313 ( .A1(n5174), .A2(n5173), .ZN(n5438) );
  AOI21_X1 U5314 ( .B1(n4894), .B2(n4891), .A(n4890), .ZN(n4889) );
  INV_X1 U5315 ( .A(n5166), .ZN(n4890) );
  INV_X1 U5316 ( .A(n5161), .ZN(n4891) );
  INV_X1 U5317 ( .A(n4894), .ZN(n4892) );
  INV_X1 U5318 ( .A(n5516), .ZN(n4728) );
  AND2_X1 U5319 ( .A1(n5152), .A2(n5148), .ZN(n5097) );
  OR2_X1 U5320 ( .A1(n5641), .A2(P1_IR_REG_7__SCAN_IN), .ZN(n5535) );
  NAND2_X1 U5321 ( .A1(n4872), .A2(n5133), .ZN(n5639) );
  NAND2_X1 U5322 ( .A1(n5111), .A2(n5110), .ZN(n5565) );
  OR2_X1 U5323 ( .A1(n6430), .A2(n6896), .ZN(n6442) );
  NAND2_X1 U5324 ( .A1(n8681), .A2(n6800), .ZN(n5042) );
  OR2_X1 U5325 ( .A1(n6802), .A2(n6801), .ZN(n5041) );
  INV_X1 U5326 ( .A(n8769), .ZN(n5043) );
  NAND2_X1 U5327 ( .A1(n6324), .A2(n6323), .ZN(n6342) );
  INV_X1 U5328 ( .A(n6340), .ZN(n6324) );
  INV_X1 U5329 ( .A(n4526), .ZN(n6372) );
  NAND2_X1 U5330 ( .A1(n4526), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n6388) );
  OR2_X1 U5331 ( .A1(n7932), .A2(n5019), .ZN(n5018) );
  INV_X1 U5332 ( .A(n6759), .ZN(n5019) );
  NAND2_X1 U5333 ( .A1(n6276), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n6299) );
  INV_X1 U5334 ( .A(n6297), .ZN(n6276) );
  NAND2_X1 U5335 ( .A1(n4525), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n6287) );
  INV_X1 U5336 ( .A(n6299), .ZN(n4525) );
  AND2_X1 U5337 ( .A1(n6752), .A2(n6747), .ZN(n5002) );
  AOI22_X1 U5338 ( .A1(n5055), .A2(n5059), .B1(n4437), .B2(n5057), .ZN(n5053)
         );
  OR2_X2 U5339 ( .A1(n8743), .A2(n5054), .ZN(n5052) );
  NOR2_X1 U5340 ( .A1(n5055), .A2(n5057), .ZN(n5054) );
  NAND2_X1 U5341 ( .A1(n4878), .A2(n4420), .ZN(n4876) );
  NAND2_X1 U5342 ( .A1(n6626), .A2(n4397), .ZN(n6620) );
  NAND2_X1 U5343 ( .A1(n4876), .A2(n4874), .ZN(n4877) );
  NOR2_X1 U5344 ( .A1(n4875), .A2(n6658), .ZN(n4874) );
  INV_X1 U5345 ( .A(n6623), .ZN(n4875) );
  OAI21_X1 U5346 ( .B1(n7272), .B2(n7575), .A(n4646), .ZN(n4645) );
  NAND2_X1 U5347 ( .A1(n7272), .A2(n7575), .ZN(n4646) );
  NOR2_X1 U5348 ( .A1(n4645), .A2(n4644), .ZN(n7263) );
  NAND2_X1 U5349 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), 
        .ZN(n4644) );
  AOI21_X1 U5350 ( .B1(n7239), .B2(n7143), .A(n7142), .ZN(n7145) );
  AND2_X1 U5351 ( .A1(n7315), .A2(n7316), .ZN(n7313) );
  AOI21_X1 U5352 ( .B1(n4654), .B2(n4417), .A(n4408), .ZN(n4653) );
  NOR2_X1 U5353 ( .A1(n8857), .A2(n4638), .ZN(n8878) );
  NOR2_X1 U5354 ( .A1(n8869), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n4638) );
  NAND2_X1 U5355 ( .A1(n8878), .A2(n8877), .ZN(n8876) );
  NAND2_X1 U5356 ( .A1(n8850), .A2(n8849), .ZN(n8848) );
  NOR2_X1 U5357 ( .A1(n8873), .A2(n4516), .ZN(n8544) );
  AND2_X1 U5358 ( .A1(n8543), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n4516) );
  INV_X1 U5359 ( .A(n8946), .ZN(n8899) );
  NOR2_X1 U5360 ( .A1(n8946), .A2(n8634), .ZN(n8900) );
  NAND2_X1 U5361 ( .A1(n8945), .A2(n6451), .ZN(n8970) );
  OR2_X1 U5362 ( .A1(n8932), .A2(n8931), .ZN(n8956) );
  NAND2_X1 U5363 ( .A1(n6463), .A2(n6462), .ZN(n8964) );
  INV_X1 U5364 ( .A(n8953), .ZN(n9016) );
  NAND2_X1 U5365 ( .A1(n9046), .A2(n5079), .ZN(n9038) );
  NAND2_X1 U5366 ( .A1(n5105), .A2(n4447), .ZN(n4858) );
  AND2_X1 U5367 ( .A1(n8632), .A2(n4548), .ZN(n9057) );
  AND2_X1 U5368 ( .A1(n6405), .A2(n6404), .ZN(n9077) );
  NOR2_X1 U5369 ( .A1(n4989), .A2(n9296), .ZN(n4987) );
  NOR2_X1 U5370 ( .A1(n9068), .A2(n9291), .ZN(n8632) );
  AND2_X1 U5371 ( .A1(n9301), .A2(n8921), .ZN(n4507) );
  AND2_X1 U5372 ( .A1(n6574), .A2(n6571), .ZN(n9120) );
  NAND2_X1 U5373 ( .A1(n4400), .A2(n4434), .ZN(n4834) );
  NOR2_X1 U5375 ( .A1(n9191), .A2(n9321), .ZN(n9165) );
  INV_X1 U5376 ( .A(n9230), .ZN(n4845) );
  AND2_X1 U5377 ( .A1(n4982), .A2(n8097), .ZN(n9209) );
  AND2_X1 U5378 ( .A1(n9337), .A2(n4407), .ZN(n4982) );
  INV_X1 U5379 ( .A(n6640), .ZN(n5067) );
  AND2_X1 U5380 ( .A1(n7102), .A2(n7121), .ZN(n9220) );
  NOR2_X1 U5381 ( .A1(n6919), .A2(n4851), .ZN(n4850) );
  NAND2_X1 U5382 ( .A1(n6198), .A2(n6197), .ZN(n7783) );
  INV_X1 U5383 ( .A(n6507), .ZN(n4542) );
  CLKBUF_X1 U5384 ( .A(n7554), .Z(n7713) );
  INV_X1 U5385 ( .A(n9225), .ZN(n9200) );
  INV_X1 U5386 ( .A(n9222), .ZN(n9205) );
  NAND2_X1 U5387 ( .A1(n6929), .A2(n6928), .ZN(n9225) );
  INV_X1 U5388 ( .A(n9287), .ZN(n10588) );
  OR3_X1 U5389 ( .A1(n7534), .A2(n7533), .A3(n7532), .ZN(n7562) );
  AND2_X1 U5390 ( .A1(n6903), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6680) );
  XNOR2_X1 U5391 ( .A(n6120), .B(P2_IR_REG_21__SCAN_IN), .ZN(n6697) );
  OAI21_X1 U5392 ( .B1(n6488), .B2(n6119), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n6120) );
  NAND2_X1 U5393 ( .A1(n7858), .A2(n7870), .ZN(n4933) );
  OR2_X1 U5394 ( .A1(n8591), .A2(n8590), .ZN(n5089) );
  OAI21_X1 U5395 ( .B1(n8318), .B2(n4967), .A(n4966), .ZN(n9413) );
  AND2_X1 U5396 ( .A1(n4970), .A2(n4968), .ZN(n4966) );
  AOI21_X1 U5397 ( .B1(n4969), .B2(n4971), .A(n8448), .ZN(n4968) );
  INV_X1 U5398 ( .A(n5089), .ZN(n4928) );
  NOR2_X1 U5399 ( .A1(n4928), .A2(n4925), .ZN(n4924) );
  INV_X1 U5400 ( .A(n9458), .ZN(n4925) );
  OR3_X1 U5401 ( .A1(n5407), .A2(n9824), .A3(n9505), .ZN(n5375) );
  NAND2_X1 U5402 ( .A1(n5430), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n5433) );
  AND2_X1 U5403 ( .A1(n9490), .A2(n8571), .ZN(n8572) );
  NAND2_X1 U5404 ( .A1(n7735), .A2(n7734), .ZN(n7859) );
  NAND2_X1 U5405 ( .A1(n8584), .A2(n8583), .ZN(n4930) );
  AND2_X1 U5406 ( .A1(n4970), .A2(n4964), .ZN(n4963) );
  NAND2_X1 U5407 ( .A1(n4969), .A2(n4971), .ZN(n4964) );
  NAND2_X1 U5408 ( .A1(n7414), .A2(n4451), .ZN(n9591) );
  NAND2_X1 U5409 ( .A1(n7193), .A2(n7081), .ZN(n7220) );
  NOR2_X1 U5410 ( .A1(n7395), .A2(n4704), .ZN(n4703) );
  INV_X1 U5411 ( .A(n7391), .ZN(n4704) );
  NOR2_X1 U5412 ( .A1(n7464), .A2(n4559), .ZN(n4558) );
  INV_X1 U5413 ( .A(n7461), .ZN(n4559) );
  INV_X1 U5414 ( .A(n4556), .ZN(n4555) );
  OAI21_X1 U5415 ( .B1(n7464), .B2(n4557), .A(n7616), .ZN(n4556) );
  NAND2_X1 U5416 ( .A1(n4562), .A2(n7461), .ZN(n4557) );
  NOR2_X1 U5417 ( .A1(n10343), .A2(n10344), .ZN(n10342) );
  NOR2_X1 U5418 ( .A1(n10338), .A2(n4584), .ZN(n9620) );
  AND2_X1 U5419 ( .A1(n9619), .A2(n9864), .ZN(n4584) );
  AND2_X1 U5420 ( .A1(n5570), .A2(n4920), .ZN(n4919) );
  INV_X1 U5421 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n4920) );
  XNOR2_X1 U5422 ( .A(n9615), .B(n9614), .ZN(n9630) );
  INV_X1 U5423 ( .A(n5695), .ZN(n9669) );
  NAND2_X1 U5424 ( .A1(n9715), .A2(n4610), .ZN(n9701) );
  NOR2_X1 U5425 ( .A1(n9697), .A2(n4611), .ZN(n4610) );
  NAND2_X1 U5426 ( .A1(n8423), .A2(n6041), .ZN(n10012) );
  NAND2_X1 U5427 ( .A1(n6040), .A2(n6039), .ZN(n8425) );
  NAND2_X1 U5428 ( .A1(n5391), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n5407) );
  NOR2_X1 U5429 ( .A1(n4908), .A2(n10226), .ZN(n4907) );
  INV_X1 U5430 ( .A(n4909), .ZN(n4908) );
  AND2_X1 U5431 ( .A1(n8033), .A2(n5968), .ZN(n8068) );
  INV_X1 U5432 ( .A(n8068), .ZN(n8059) );
  AND4_X1 U5433 ( .A1(n5559), .A2(n5558), .A3(n5557), .A4(n5556), .ZN(n8008)
         );
  NAND2_X1 U5434 ( .A1(n5007), .A2(n6016), .ZN(n7836) );
  INV_X1 U5435 ( .A(n7834), .ZN(n5007) );
  INV_X1 U5436 ( .A(n10415), .ZN(n6014) );
  NAND2_X1 U5437 ( .A1(n7345), .A2(n7349), .ZN(n6004) );
  OR2_X1 U5438 ( .A1(n5737), .A2(n6054), .ZN(n5738) );
  AND2_X1 U5439 ( .A1(n10428), .A2(n7496), .ZN(n7363) );
  NAND2_X1 U5440 ( .A1(n5713), .A2(n5712), .ZN(n9646) );
  AND2_X1 U5441 ( .A1(n10084), .A2(n5989), .ZN(n5103) );
  NAND2_X1 U5442 ( .A1(n5465), .A2(n5464), .ZN(n8450) );
  AND2_X1 U5443 ( .A1(n7234), .A2(n6951), .ZN(n10240) );
  AND2_X1 U5444 ( .A1(n6070), .A2(n6069), .ZN(n10427) );
  AND2_X1 U5445 ( .A1(n5257), .A2(n5256), .ZN(n4615) );
  XNOR2_X1 U5446 ( .A(n5248), .B(n5247), .ZN(n9384) );
  NAND2_X1 U5447 ( .A1(n5268), .A2(n5267), .ZN(n5272) );
  NOR2_X1 U5448 ( .A1(P1_IR_REG_29__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), .ZN(
        n5270) );
  XNOR2_X1 U5449 ( .A(n5699), .B(n5698), .ZN(n8640) );
  NAND2_X1 U5450 ( .A1(n5943), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5947) );
  NAND2_X1 U5451 ( .A1(n5947), .A2(n5946), .ZN(n5949) );
  XNOR2_X1 U5452 ( .A(n5314), .B(n5313), .ZN(n8402) );
  NAND2_X1 U5453 ( .A1(n4886), .A2(n4884), .ZN(n5400) );
  INV_X1 U5454 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n5460) );
  AND2_X1 U5455 ( .A1(n5507), .A2(n5506), .ZN(n7390) );
  NAND2_X1 U5456 ( .A1(n6127), .A2(n5582), .ZN(n4873) );
  NAND2_X1 U5457 ( .A1(n7631), .A2(n6351), .ZN(n6321) );
  NAND2_X1 U5458 ( .A1(n6408), .A2(n6407), .ZN(n9278) );
  AND2_X1 U5459 ( .A1(n6475), .A2(n6474), .ZN(n8969) );
  AND2_X1 U5460 ( .A1(n6427), .A2(n6426), .ZN(n9036) );
  OR2_X1 U5461 ( .A1(n9021), .A2(n6467), .ZN(n6427) );
  OR2_X1 U5462 ( .A1(n9031), .A2(n6467), .ZN(n6416) );
  OR2_X1 U5463 ( .A1(n6328), .A2(n6327), .ZN(n9175) );
  NAND2_X1 U5464 ( .A1(n6175), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n6190) );
  NAND2_X1 U5465 ( .A1(n4738), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n4737) );
  NAND2_X1 U5466 ( .A1(n7124), .A2(n7125), .ZN(n7136) );
  NAND2_X1 U5467 ( .A1(n7210), .A2(n7211), .ZN(n7297) );
  NAND2_X1 U5468 ( .A1(n4518), .A2(n4517), .ZN(n4635) );
  OR2_X1 U5469 ( .A1(n8558), .A2(n10510), .ZN(n4517) );
  NAND2_X1 U5470 ( .A1(n8557), .A2(n10506), .ZN(n4518) );
  OAI211_X1 U5471 ( .C1(n8557), .C2(n10511), .A(n4749), .B(n10509), .ZN(n4748)
         );
  NAND2_X1 U5472 ( .A1(n8558), .A2(n10505), .ZN(n4749) );
  NAND2_X1 U5473 ( .A1(n6940), .A2(n9188), .ZN(n9060) );
  NOR2_X1 U5474 ( .A1(n9258), .A2(n4684), .ZN(n4683) );
  OR2_X1 U5475 ( .A1(n10598), .A2(n9878), .ZN(n4871) );
  NAND2_X1 U5476 ( .A1(n8978), .A2(n8980), .ZN(n4867) );
  OAI21_X1 U5477 ( .B1(n8989), .B2(n8978), .A(n4866), .ZN(n4865) );
  NAND2_X1 U5478 ( .A1(n9413), .A2(n9411), .ZN(n9416) );
  OR2_X1 U5479 ( .A1(n9680), .A2(n5434), .ZN(n5312) );
  INV_X1 U5480 ( .A(n9520), .ZN(n9547) );
  NAND2_X1 U5481 ( .A1(n7502), .A2(n7501), .ZN(n9560) );
  AND2_X1 U5482 ( .A1(n5828), .A2(n5829), .ZN(n4755) );
  OR2_X1 U5483 ( .A1(n5955), .A2(n5954), .ZN(n4717) );
  INV_X1 U5484 ( .A(n8026), .ZN(n9583) );
  INV_X1 U5485 ( .A(n8008), .ZN(n9584) );
  INV_X1 U5486 ( .A(n7088), .ZN(n4694) );
  INV_X1 U5487 ( .A(n7183), .ZN(n4695) );
  NOR2_X1 U5488 ( .A1(n7250), .A2(n4590), .ZN(n7386) );
  NOR2_X1 U5489 ( .A1(n7254), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n4590) );
  AOI21_X1 U5490 ( .B1(n4534), .B2(n4496), .A(n4532), .ZN(n4588) );
  NAND2_X1 U5491 ( .A1(n4533), .A2(n4589), .ZN(n4532) );
  INV_X1 U5492 ( .A(n9630), .ZN(n4534) );
  NOR2_X1 U5493 ( .A1(n10363), .A2(n9733), .ZN(n4589) );
  AOI21_X1 U5494 ( .B1(n9630), .B2(n10383), .A(n9632), .ZN(n4586) );
  AOI21_X1 U5495 ( .B1(n4568), .B2(n10364), .A(n4566), .ZN(n4565) );
  NAND2_X1 U5496 ( .A1(n9624), .A2(n4568), .ZN(n4564) );
  NAND3_X1 U5497 ( .A1(n10465), .A2(n10428), .A3(n7930), .ZN(n10145) );
  NOR3_X2 U5498 ( .A1(n9651), .A2(n6066), .A3(n6065), .ZN(n6695) );
  NOR3_X1 U5499 ( .A1(n9653), .A2(n10243), .A3(n6051), .ZN(n6066) );
  NOR3_X1 U5500 ( .A1(n6516), .A2(n6510), .A3(n6509), .ZN(n6525) );
  NAND2_X1 U5501 ( .A1(n5742), .A2(n5741), .ZN(n4510) );
  NOR2_X1 U5502 ( .A1(n4811), .A2(n6950), .ZN(n4509) );
  INV_X1 U5503 ( .A(n4773), .ZN(n4772) );
  NAND2_X1 U5504 ( .A1(n5761), .A2(n4551), .ZN(n4768) );
  NOR3_X1 U5505 ( .A1(n4779), .A2(n6950), .A3(n5854), .ZN(n4551) );
  INV_X1 U5506 ( .A(n5758), .ZN(n4779) );
  AOI21_X1 U5507 ( .B1(n4773), .B2(n4770), .A(n4458), .ZN(n4769) );
  INV_X1 U5508 ( .A(n4775), .ZN(n4770) );
  NOR2_X1 U5509 ( .A1(n4778), .A2(n6950), .ZN(n4774) );
  INV_X1 U5510 ( .A(n6571), .ZN(n4819) );
  NAND2_X1 U5511 ( .A1(n6577), .A2(n4397), .ZN(n4818) );
  MUX2_X1 U5512 ( .A(n6565), .B(n6564), .S(n4394), .Z(n6566) );
  NAND2_X1 U5513 ( .A1(n4750), .A2(n6950), .ZN(n4631) );
  NAND2_X1 U5514 ( .A1(n5775), .A2(n4751), .ZN(n4632) );
  INV_X1 U5515 ( .A(n5841), .ZN(n4750) );
  NOR2_X1 U5516 ( .A1(n4814), .A2(n4813), .ZN(n4812) );
  INV_X1 U5517 ( .A(n4816), .ZN(n4815) );
  AOI21_X1 U5518 ( .B1(n4796), .B2(n6601), .A(n4431), .ZN(n4794) );
  AOI21_X1 U5519 ( .B1(n4794), .B2(n4792), .A(n8963), .ZN(n4791) );
  INV_X1 U5520 ( .A(n4796), .ZN(n4792) );
  INV_X1 U5521 ( .A(n5776), .ZN(n5842) );
  INV_X1 U5522 ( .A(n7349), .ZN(n5739) );
  INV_X1 U5523 ( .A(n5100), .ZN(n4600) );
  NAND2_X1 U5524 ( .A1(n4791), .A2(n4793), .ZN(n4790) );
  INV_X1 U5525 ( .A(n4794), .ZN(n4793) );
  NOR2_X1 U5526 ( .A1(n6610), .A2(n6628), .ZN(n4795) );
  AOI21_X1 U5527 ( .B1(n5074), .B2(n5076), .A(n5075), .ZN(n5072) );
  NOR2_X1 U5528 ( .A1(n6476), .A2(n6608), .ZN(n5074) );
  INV_X1 U5529 ( .A(n8101), .ZN(n4985) );
  INV_X1 U5530 ( .A(n6587), .ZN(n4674) );
  INV_X1 U5531 ( .A(n4673), .ZN(n4672) );
  OAI21_X1 U5532 ( .B1(n5079), .B2(n4674), .A(n9016), .ZN(n4673) );
  NAND2_X1 U5533 ( .A1(n7696), .A2(n6907), .ZN(n6501) );
  AND2_X1 U5534 ( .A1(n5339), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n5317) );
  NOR2_X1 U5535 ( .A1(n5365), .A2(n8527), .ZN(n5339) );
  NOR2_X1 U5536 ( .A1(n5346), .A2(n10042), .ZN(n5960) );
  INV_X1 U5537 ( .A(n6031), .ZN(n5021) );
  AND2_X1 U5538 ( .A1(n6035), .A2(n5023), .ZN(n5020) );
  NAND2_X1 U5539 ( .A1(n5024), .A2(n6034), .ZN(n5023) );
  NOR2_X1 U5540 ( .A1(n10086), .A2(n10111), .ZN(n6035) );
  INV_X1 U5541 ( .A(n6033), .ZN(n5024) );
  OAI21_X1 U5542 ( .B1(n6016), .B2(n5006), .A(n7889), .ZN(n5005) );
  INV_X1 U5543 ( .A(n5280), .ZN(n4734) );
  AOI21_X1 U5544 ( .B1(n4733), .B2(n5280), .A(n4491), .ZN(n4732) );
  INV_X1 U5545 ( .A(n5235), .ZN(n4733) );
  INV_X1 U5546 ( .A(n5313), .ZN(n4714) );
  INV_X1 U5547 ( .A(n5224), .ZN(n4712) );
  INV_X1 U5548 ( .A(n5209), .ZN(n4726) );
  INV_X1 U5549 ( .A(n5216), .ZN(n4725) );
  NAND2_X1 U5550 ( .A1(n5190), .A2(n5189), .ZN(n5195) );
  INV_X1 U5551 ( .A(SI_19_), .ZN(n5189) );
  NAND2_X1 U5552 ( .A1(n5171), .A2(n5170), .ZN(n5174) );
  INV_X1 U5553 ( .A(SI_13_), .ZN(n5162) );
  AND2_X1 U5554 ( .A1(n5501), .A2(n5498), .ZN(n5144) );
  OAI21_X1 U5555 ( .B1(n7001), .B2(n5130), .A(n5129), .ZN(n5132) );
  NOR2_X1 U5556 ( .A1(n6614), .A2(n6617), .ZN(n4879) );
  NAND2_X1 U5557 ( .A1(n6627), .A2(n4394), .ZN(n6619) );
  OR2_X1 U5558 ( .A1(n6161), .A2(n6147), .ZN(n6148) );
  OR2_X1 U5559 ( .A1(n6161), .A2(n6140), .ZN(n6141) );
  NAND2_X1 U5560 ( .A1(n8538), .A2(n4519), .ZN(n8540) );
  OR2_X1 U5561 ( .A1(n8539), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n4519) );
  NOR2_X1 U5562 ( .A1(n9259), .A2(n9261), .ZN(n4986) );
  NAND2_X1 U5563 ( .A1(n10288), .A2(n6351), .ZN(n6604) );
  OR2_X1 U5564 ( .A1(n9268), .A2(n8991), .ZN(n8960) );
  OR2_X1 U5565 ( .A1(n9291), .A2(n9092), .ZN(n6406) );
  AND2_X1 U5566 ( .A1(n6559), .A2(n9142), .ZN(n6347) );
  NAND2_X1 U5567 ( .A1(n5063), .A2(n9184), .ZN(n5062) );
  INV_X1 U5568 ( .A(n6537), .ZN(n5071) );
  NAND2_X1 U5569 ( .A1(n4524), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n6297) );
  INV_X1 U5570 ( .A(n6261), .ZN(n4524) );
  NAND2_X1 U5571 ( .A1(n8048), .A2(n6241), .ZN(n8090) );
  AND2_X1 U5572 ( .A1(n6233), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n6248) );
  NOR2_X1 U5573 ( .A1(n7671), .A2(n10569), .ZN(n7569) );
  NOR2_X1 U5574 ( .A1(n7556), .A2(n8759), .ZN(n7719) );
  NAND2_X1 U5575 ( .A1(n6501), .A2(n6908), .ZN(n7579) );
  OR2_X1 U5576 ( .A1(P2_IR_REG_27__SCAN_IN), .A2(P2_IR_REG_28__SCAN_IN), .ZN(
        n6109) );
  INV_X1 U5577 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n6107) );
  NAND2_X1 U5578 ( .A1(n6661), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6662) );
  NOR2_X1 U5579 ( .A1(P2_IR_REG_18__SCAN_IN), .A2(P2_IR_REG_17__SCAN_IN), .ZN(
        n5031) );
  INV_X1 U5580 ( .A(n7865), .ZN(n7425) );
  OR2_X1 U5581 ( .A1(n4951), .A2(n4950), .ZN(n4946) );
  NAND2_X1 U5582 ( .A1(n4954), .A2(n4955), .ZN(n4949) );
  NAND2_X1 U5583 ( .A1(n8566), .A2(n8520), .ZN(n4955) );
  NOR2_X1 U5584 ( .A1(n5668), .A2(n5632), .ZN(n5552) );
  AOI22_X1 U5585 ( .A1(n8459), .A2(n4439), .B1(n4941), .B2(n4404), .ZN(n4938)
         );
  INV_X1 U5586 ( .A(n8486), .ZN(n4943) );
  NAND2_X1 U5587 ( .A1(n8520), .A2(n4959), .ZN(n4958) );
  INV_X1 U5588 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n5510) );
  NOR2_X1 U5589 ( .A1(n5523), .A2(n5522), .ZN(n5491) );
  NAND2_X1 U5590 ( .A1(n4939), .A2(n8472), .ZN(n9436) );
  INV_X1 U5591 ( .A(n8473), .ZN(n4940) );
  AND2_X1 U5592 ( .A1(n8440), .A2(n8439), .ZN(n4974) );
  INV_X1 U5593 ( .A(n4975), .ZN(n4972) );
  AND2_X1 U5594 ( .A1(n5445), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n5430) );
  NOR2_X1 U5595 ( .A1(n5478), .A2(n9766), .ZN(n5445) );
  AND2_X1 U5596 ( .A1(n6875), .A2(n4764), .ZN(n4763) );
  NAND2_X1 U5597 ( .A1(n9646), .A2(n6002), .ZN(n5897) );
  NAND2_X1 U5598 ( .A1(n6049), .A2(n6050), .ZN(n5028) );
  NOR2_X1 U5599 ( .A1(n9690), .A2(n10190), .ZN(n4904) );
  NAND2_X1 U5600 ( .A1(n5013), .A2(n6043), .ZN(n5012) );
  INV_X1 U5601 ( .A(n6042), .ZN(n5013) );
  NOR2_X1 U5602 ( .A1(n5014), .A2(n5010), .ZN(n5009) );
  INV_X1 U5603 ( .A(n6041), .ZN(n5010) );
  INV_X1 U5604 ( .A(n5960), .ZN(n5795) );
  INV_X1 U5605 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n9824) );
  NOR2_X1 U5606 ( .A1(n5433), .A2(n9791), .ZN(n5391) );
  INV_X1 U5607 ( .A(n6034), .ZN(n5025) );
  NAND2_X1 U5608 ( .A1(n4403), .A2(n5049), .ZN(n5045) );
  NAND2_X1 U5609 ( .A1(n5762), .A2(n5856), .ZN(n6024) );
  NAND2_X1 U5610 ( .A1(n5048), .A2(n6019), .ZN(n5047) );
  INV_X1 U5611 ( .A(n7905), .ZN(n5048) );
  NOR2_X1 U5612 ( .A1(n8163), .A2(n10475), .ZN(n4901) );
  AND3_X1 U5613 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .A3(P1_REG3_REG_5__SCAN_IN), .ZN(n5655) );
  INV_X1 U5614 ( .A(n5991), .ZN(n4550) );
  NAND2_X1 U5615 ( .A1(n10084), .A2(n4822), .ZN(n10069) );
  NOR2_X2 U5616 ( .A1(n8180), .A2(n8287), .ZN(n8220) );
  INV_X1 U5617 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n5261) );
  NOR2_X1 U5618 ( .A1(n5266), .A2(n4918), .ZN(n5267) );
  INV_X1 U5619 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n5266) );
  OAI21_X1 U5620 ( .B1(n5314), .B2(n4713), .A(n4710), .ZN(n5293) );
  AOI21_X1 U5621 ( .B1(n5301), .B2(n4712), .A(n4711), .ZN(n4710) );
  NAND2_X1 U5622 ( .A1(n4714), .A2(n5301), .ZN(n4713) );
  INV_X1 U5623 ( .A(n5229), .ZN(n4711) );
  AND2_X1 U5624 ( .A1(n5235), .A2(n5234), .ZN(n5294) );
  NAND2_X1 U5625 ( .A1(n5200), .A2(n5199), .ZN(n5359) );
  INV_X1 U5626 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n5724) );
  INV_X1 U5627 ( .A(n5180), .ZN(n4885) );
  OR2_X1 U5628 ( .A1(n5188), .A2(n5187), .ZN(n5399) );
  NAND2_X1 U5629 ( .A1(n5158), .A2(n5157), .ZN(n5161) );
  INV_X1 U5630 ( .A(SI_12_), .ZN(n5157) );
  OR2_X1 U5631 ( .A1(n5532), .A2(n5459), .ZN(n5503) );
  INV_X1 U5632 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n5536) );
  NAND2_X1 U5633 ( .A1(n5639), .A2(n5134), .ZN(n5137) );
  AOI21_X1 U5634 ( .B1(n5126), .B2(n4418), .A(n5104), .ZN(n5127) );
  INV_X1 U5635 ( .A(n5128), .ZN(n7002) );
  INV_X1 U5636 ( .A(n6705), .ZN(n6754) );
  NAND2_X1 U5637 ( .A1(n6325), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n6365) );
  INV_X1 U5638 ( .A(n6342), .ZN(n6325) );
  INV_X1 U5639 ( .A(n8717), .ZN(n5037) );
  NAND2_X1 U5640 ( .A1(n5001), .A2(n6714), .ZN(n8756) );
  INV_X1 U5641 ( .A(n6989), .ZN(n5001) );
  OR2_X1 U5642 ( .A1(n8678), .A2(n8681), .ZN(n8679) );
  OR2_X1 U5643 ( .A1(n6789), .A2(n6788), .ZN(n5033) );
  NAND2_X1 U5644 ( .A1(n6176), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n6204) );
  OAI21_X1 U5645 ( .B1(n5000), .B2(n6989), .A(n6726), .ZN(n7606) );
  NAND2_X1 U5646 ( .A1(n6714), .A2(n4441), .ZN(n5000) );
  AND3_X1 U5647 ( .A1(n6369), .A2(n6368), .A3(n6367), .ZN(n8918) );
  AND4_X1 U5648 ( .A1(n6346), .A2(n6345), .A3(n6344), .A4(n6343), .ZN(n8833)
         );
  AND2_X1 U5649 ( .A1(n6167), .A2(n6165), .ZN(n4543) );
  NAND2_X1 U5650 ( .A1(n6468), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n6166) );
  NAND2_X1 U5651 ( .A1(n6175), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n4836) );
  OAI21_X1 U5652 ( .B1(n7145), .B2(n7113), .A(n7112), .ZN(n7131) );
  AND2_X1 U5653 ( .A1(n4637), .A2(n4636), .ZN(n7157) );
  INV_X1 U5654 ( .A(n7129), .ZN(n4636) );
  NAND2_X1 U5655 ( .A1(n7131), .A2(n7130), .ZN(n4637) );
  OAI21_X1 U5656 ( .B1(n7157), .B2(n7156), .A(n7155), .ZN(n7170) );
  NOR2_X1 U5657 ( .A1(n7313), .A2(n4736), .ZN(n7301) );
  AND2_X1 U5658 ( .A1(n7299), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n4736) );
  NAND2_X1 U5659 ( .A1(n7336), .A2(n7337), .ZN(n7477) );
  AND2_X1 U5660 ( .A1(n6271), .A2(n6270), .ZN(n6292) );
  NAND2_X1 U5661 ( .A1(n7645), .A2(n4740), .ZN(n7647) );
  OR2_X1 U5662 ( .A1(n7646), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n4740) );
  NAND2_X1 U5663 ( .A1(n7647), .A2(n7648), .ZN(n7766) );
  AOI21_X1 U5664 ( .B1(n4650), .B2(n4652), .A(n4426), .ZN(n4648) );
  NAND2_X1 U5665 ( .A1(n7766), .A2(n4739), .ZN(n7768) );
  OR2_X1 U5666 ( .A1(n7767), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n4739) );
  NAND2_X1 U5667 ( .A1(n7768), .A2(n7769), .ZN(n8538) );
  OR2_X1 U5668 ( .A1(n7640), .A2(n7639), .ZN(n4642) );
  OR2_X1 U5669 ( .A1(n7763), .A2(n7762), .ZN(n4640) );
  AND2_X1 U5670 ( .A1(n4640), .A2(n4639), .ZN(n8552) );
  NAND2_X1 U5671 ( .A1(n8550), .A2(n9747), .ZN(n4639) );
  NAND2_X1 U5672 ( .A1(n8876), .A2(n4497), .ZN(n8887) );
  NOR2_X1 U5673 ( .A1(n8887), .A2(n8886), .ZN(n8885) );
  NAND2_X1 U5674 ( .A1(n6612), .A2(n6611), .ZN(n6628) );
  NAND2_X1 U5675 ( .A1(n6604), .A2(n6603), .ZN(n9259) );
  NAND2_X1 U5676 ( .A1(n9007), .A2(n8987), .ZN(n8981) );
  AND2_X1 U5677 ( .A1(n6458), .A2(n6457), .ZN(n8992) );
  OR2_X1 U5678 ( .A1(n8970), .A2(n6467), .ZN(n6458) );
  AND2_X1 U5679 ( .A1(n6442), .A2(n6431), .ZN(n9008) );
  NAND2_X1 U5680 ( .A1(n4527), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n6430) );
  INV_X1 U5681 ( .A(n4527), .ZN(n6420) );
  OR2_X1 U5682 ( .A1(n6388), .A2(n6387), .ZN(n6399) );
  NAND2_X1 U5683 ( .A1(n6398), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n6409) );
  INV_X1 U5684 ( .A(n6399), .ZN(n6398) );
  INV_X1 U5685 ( .A(n9044), .ZN(n9054) );
  NAND2_X1 U5686 ( .A1(n8923), .A2(n8922), .ZN(n9066) );
  AND3_X1 U5687 ( .A1(n6376), .A2(n6375), .A3(n6374), .ZN(n9091) );
  NAND2_X1 U5688 ( .A1(n9103), .A2(n6577), .ZN(n9088) );
  AND2_X1 U5689 ( .A1(n6580), .A2(n9072), .ZN(n9087) );
  INV_X1 U5690 ( .A(n4989), .ZN(n4988) );
  NAND2_X1 U5691 ( .A1(n4829), .A2(n4831), .ZN(n9099) );
  INV_X1 U5692 ( .A(n4832), .ZN(n4831) );
  OAI21_X1 U5693 ( .B1(n4834), .B2(n4833), .A(n8920), .ZN(n4832) );
  NAND2_X1 U5694 ( .A1(n9127), .A2(n4991), .ZN(n9113) );
  NAND2_X1 U5695 ( .A1(n9127), .A2(n9133), .ZN(n9128) );
  NAND2_X1 U5696 ( .A1(n9180), .A2(n9184), .ZN(n9143) );
  NAND2_X1 U5697 ( .A1(n9209), .A2(n8631), .ZN(n9191) );
  NAND2_X1 U5698 ( .A1(n6307), .A2(n6306), .ZN(n9180) );
  AND4_X1 U5699 ( .A1(n6291), .A2(n6290), .A3(n6289), .A4(n6288), .ZN(n9204)
         );
  AND4_X1 U5700 ( .A1(n6316), .A2(n6315), .A3(n6314), .A4(n6313), .ZN(n9206)
         );
  INV_X1 U5701 ( .A(n8295), .ZN(n4863) );
  AND2_X1 U5702 ( .A1(n8298), .A2(n6632), .ZN(n9230) );
  NAND2_X1 U5703 ( .A1(n8097), .A2(n4984), .ZN(n9226) );
  AND4_X1 U5704 ( .A1(n6303), .A2(n6302), .A3(n6301), .A4(n6300), .ZN(n8304)
         );
  NAND2_X1 U5705 ( .A1(n6256), .A2(n8090), .ZN(n8093) );
  NAND2_X1 U5706 ( .A1(n8097), .A2(n8101), .ZN(n8119) );
  NAND2_X1 U5707 ( .A1(n6927), .A2(n6530), .ZN(n8048) );
  NOR2_X1 U5708 ( .A1(n7556), .A2(n7824), .ZN(n4992) );
  NAND2_X1 U5709 ( .A1(n7816), .A2(n6527), .ZN(n6925) );
  NAND2_X1 U5710 ( .A1(n4661), .A2(n4660), .ZN(n4659) );
  NAND2_X1 U5711 ( .A1(n7779), .A2(n4662), .ZN(n4661) );
  AND2_X1 U5712 ( .A1(n7102), .A2(n7105), .ZN(n9222) );
  NAND2_X1 U5713 ( .A1(n4429), .A2(n4993), .ZN(n7810) );
  INV_X1 U5714 ( .A(n7556), .ZN(n4993) );
  NOR2_X1 U5715 ( .A1(n7556), .A2(n4994), .ZN(n7782) );
  NAND2_X1 U5716 ( .A1(n7680), .A2(n10575), .ZN(n4994) );
  INV_X1 U5717 ( .A(n7711), .ZN(n7776) );
  NAND2_X1 U5718 ( .A1(n6192), .A2(n6146), .ZN(n4979) );
  INV_X1 U5719 ( .A(n4981), .ZN(n4980) );
  NAND2_X1 U5720 ( .A1(n7521), .A2(n10569), .ZN(n7696) );
  AND2_X1 U5721 ( .A1(n8940), .A2(n8939), .ZN(n9253) );
  OR2_X1 U5722 ( .A1(n8938), .A2(n8955), .ZN(n8939) );
  OR2_X1 U5723 ( .A1(n9259), .A2(n8941), .ZN(n9243) );
  NAND2_X1 U5724 ( .A1(n9259), .A2(n9356), .ZN(n4685) );
  OAI21_X1 U5725 ( .B1(n8989), .B2(n8979), .A(n8978), .ZN(n4866) );
  NAND2_X1 U5726 ( .A1(n6232), .A2(n6231), .ZN(n9355) );
  INV_X1 U5727 ( .A(n10590), .ZN(n9357) );
  INV_X1 U5728 ( .A(n6717), .ZN(n10575) );
  AND2_X1 U5729 ( .A1(n6833), .A2(n6832), .ZN(n10531) );
  OAI21_X1 U5730 ( .B1(n6662), .B2(n6665), .A(n6676), .ZN(n6903) );
  INV_X1 U5731 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n5083) );
  INV_X1 U5732 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n6665) );
  AND3_X1 U5733 ( .A1(n5092), .A2(n5081), .A3(n6490), .ZN(n5082) );
  NAND2_X1 U5734 ( .A1(n6662), .A2(n6665), .ZN(n6676) );
  XNOR2_X1 U5735 ( .A(n6242), .B(P2_IR_REG_9__SCAN_IN), .ZN(n7299) );
  AND2_X1 U5736 ( .A1(n6210), .A2(n6195), .ZN(n7167) );
  NOR2_X1 U5737 ( .A1(n9427), .A2(n9426), .ZN(n9486) );
  INV_X1 U5738 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n9915) );
  NAND2_X1 U5739 ( .A1(n9500), .A2(n9502), .ZN(n9448) );
  NAND2_X1 U5740 ( .A1(n4952), .A2(n4951), .ZN(n8524) );
  INV_X1 U5741 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n5522) );
  AND2_X1 U5742 ( .A1(n7859), .A2(n7858), .ZN(n9523) );
  AND2_X1 U5743 ( .A1(n5425), .A2(n5424), .ZN(n10156) );
  NAND2_X1 U5744 ( .A1(n5664), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n4757) );
  NAND2_X1 U5745 ( .A1(n6979), .A2(n4696), .ZN(n7277) );
  NAND2_X1 U5746 ( .A1(n7280), .A2(n7062), .ZN(n7412) );
  NOR2_X1 U5747 ( .A1(n7063), .A2(n4701), .ZN(n4700) );
  INV_X1 U5748 ( .A(n7062), .ZN(n4701) );
  NAND2_X1 U5749 ( .A1(n4583), .A2(n4582), .ZN(n7407) );
  NAND2_X1 U5750 ( .A1(n4579), .A2(n4578), .ZN(n7053) );
  NAND2_X1 U5751 ( .A1(n4583), .A2(n4443), .ZN(n4579) );
  NAND2_X1 U5752 ( .A1(n4581), .A2(n7051), .ZN(n4578) );
  NAND2_X1 U5753 ( .A1(n7182), .A2(n4692), .ZN(n7215) );
  AND2_X1 U5754 ( .A1(n7090), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n4692) );
  NAND2_X1 U5755 ( .A1(n4561), .A2(n4415), .ZN(n4560) );
  INV_X1 U5756 ( .A(n7462), .ZN(n4561) );
  OR2_X1 U5757 ( .A1(n9607), .A2(n9606), .ZN(n10330) );
  INV_X1 U5758 ( .A(n9609), .ZN(n9608) );
  OR2_X1 U5759 ( .A1(n10359), .A2(n10358), .ZN(n10355) );
  NAND2_X1 U5760 ( .A1(n4570), .A2(n4567), .ZN(n10377) );
  INV_X1 U5761 ( .A(n4569), .ZN(n4567) );
  AND2_X1 U5762 ( .A1(n10393), .A2(n4577), .ZN(n4574) );
  NAND2_X1 U5763 ( .A1(n10377), .A2(n10378), .ZN(n4575) );
  NAND2_X1 U5764 ( .A1(n9631), .A2(n10395), .ZN(n4533) );
  NOR2_X1 U5765 ( .A1(n4573), .A2(n4569), .ZN(n4568) );
  INV_X1 U5766 ( .A(n4574), .ZN(n4573) );
  INV_X1 U5767 ( .A(n4572), .ZN(n4566) );
  AOI21_X1 U5768 ( .B1(n10393), .B2(n4414), .A(n9628), .ZN(n4572) );
  XNOR2_X1 U5769 ( .A(n4595), .B(n6051), .ZN(n4594) );
  NAND2_X1 U5770 ( .A1(n6878), .A2(n5999), .ZN(n4595) );
  AND2_X1 U5771 ( .A1(n5287), .A2(n9656), .ZN(n8620) );
  NAND2_X1 U5772 ( .A1(n9732), .A2(n4904), .ZN(n9691) );
  NAND2_X1 U5773 ( .A1(n9732), .A2(n9708), .ZN(n9703) );
  AND2_X1 U5774 ( .A1(n5358), .A2(n5357), .ZN(n9721) );
  OR2_X1 U5775 ( .A1(n10017), .A2(n5434), .ZN(n5358) );
  AND2_X1 U5776 ( .A1(n5795), .A2(n5991), .ZN(n8430) );
  AND2_X1 U5777 ( .A1(n8426), .A2(n5778), .ZN(n10070) );
  NAND2_X1 U5778 ( .A1(n10085), .A2(n5988), .ZN(n10084) );
  AND2_X1 U5779 ( .A1(n5843), .A2(n5989), .ZN(n10086) );
  AND2_X1 U5780 ( .A1(n5412), .A2(n5411), .ZN(n10107) );
  NAND2_X1 U5781 ( .A1(n10102), .A2(n10111), .ZN(n10085) );
  AND2_X1 U5782 ( .A1(n5398), .A2(n5397), .ZN(n10133) );
  NAND2_X1 U5783 ( .A1(n8215), .A2(n5979), .ZN(n4502) );
  NAND2_X1 U5784 ( .A1(n10144), .A2(n10153), .ZN(n6032) );
  AND2_X1 U5785 ( .A1(n5767), .A2(n5983), .ZN(n10143) );
  NAND2_X1 U5786 ( .A1(n8221), .A2(n4909), .ZN(n10160) );
  NAND2_X1 U5787 ( .A1(n8221), .A2(n9557), .ZN(n10159) );
  AND3_X1 U5788 ( .A1(n5437), .A2(n5436), .A3(n5435), .ZN(n10132) );
  INV_X1 U5789 ( .A(n6024), .ZN(n8174) );
  NAND2_X1 U5790 ( .A1(n5046), .A2(n4399), .ZN(n8169) );
  OR2_X1 U5791 ( .A1(n7906), .A2(n5049), .ZN(n5046) );
  AND4_X1 U5792 ( .A1(n5529), .A2(n5528), .A3(n5527), .A4(n5526), .ZN(n8202)
         );
  AND4_X1 U5793 ( .A1(n5497), .A2(n5496), .A3(n5495), .A4(n5494), .ZN(n8264)
         );
  AND2_X1 U5794 ( .A1(n8138), .A2(n5971), .ZN(n8035) );
  NAND2_X1 U5795 ( .A1(n4899), .A2(n4901), .ZN(n8061) );
  NAND2_X1 U5796 ( .A1(n4628), .A2(n5743), .ZN(n4753) );
  AOI21_X1 U5797 ( .B1(n5744), .B2(n4628), .A(n4811), .ZN(n4627) );
  AOI21_X1 U5798 ( .B1(n5592), .B2(P2_DATAO_REG_7__SCAN_IN), .A(n4433), .ZN(
        n4759) );
  NAND2_X1 U5799 ( .A1(n6999), .A2(n5675), .ZN(n4760) );
  NOR2_X1 U5800 ( .A1(n6055), .A2(n9531), .ZN(n4905) );
  AND2_X1 U5801 ( .A1(n5867), .A2(n5911), .ZN(n7842) );
  AND3_X1 U5802 ( .A1(n4906), .A2(n6010), .A3(n10421), .ZN(n10417) );
  OR2_X1 U5803 ( .A1(n7921), .A2(n7924), .ZN(n10416) );
  INV_X1 U5804 ( .A(n5011), .ZN(n9728) );
  AOI21_X1 U5805 ( .B1(n10012), .B2(n6042), .A(n5014), .ZN(n5011) );
  NAND2_X1 U5806 ( .A1(n5406), .A2(n5405), .ZN(n10217) );
  NAND2_X1 U5807 ( .A1(n5444), .A2(n5443), .ZN(n8454) );
  OR2_X1 U5808 ( .A1(n7791), .A2(n6950), .ZN(n10473) );
  OAI21_X1 U5809 ( .B1(n4784), .B2(n7796), .A(n7795), .ZN(n7797) );
  INV_X1 U5810 ( .A(n10473), .ZN(n10465) );
  NAND2_X1 U5811 ( .A1(n6073), .A2(n6072), .ZN(n7358) );
  XNOR2_X1 U5812 ( .A(n5711), .B(n5710), .ZN(n8627) );
  NAND2_X2 U5813 ( .A1(n5265), .A2(n5269), .ZN(n10306) );
  MUX2_X1 U5814 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5264), .S(
        P1_IR_REG_27__SCAN_IN), .Z(n5265) );
  OAI21_X1 U5815 ( .B1(n5314), .B2(n5313), .A(n5224), .ZN(n5302) );
  OAI21_X2 U5816 ( .B1(n5942), .B2(P1_IR_REG_23__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5951) );
  NAND2_X1 U5817 ( .A1(n4727), .A2(n5209), .ZN(n5348) );
  NAND2_X1 U5818 ( .A1(n4723), .A2(n4721), .ZN(n4727) );
  NAND2_X1 U5819 ( .A1(n5731), .A2(n4453), .ZN(n5736) );
  NAND2_X1 U5820 ( .A1(n4723), .A2(n5204), .ZN(n4606) );
  NAND2_X1 U5821 ( .A1(n5731), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5727) );
  XNOR2_X1 U5822 ( .A(n5359), .B(n5360), .ZN(n7929) );
  INV_X1 U5823 ( .A(n4917), .ZN(n4916) );
  OAI21_X1 U5824 ( .B1(n5723), .B2(n4918), .A(n5724), .ZN(n4917) );
  NAND2_X1 U5825 ( .A1(n4915), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5403) );
  NAND2_X1 U5826 ( .A1(n5415), .A2(n5723), .ZN(n4915) );
  XNOR2_X1 U5827 ( .A(n5386), .B(n5385), .ZN(n7655) );
  NAND2_X1 U5828 ( .A1(n4528), .A2(n5413), .ZN(n5384) );
  INV_X1 U5829 ( .A(n5414), .ZN(n4528) );
  OAI21_X1 U5830 ( .B1(n5484), .B2(n4892), .A(n4889), .ZN(n5455) );
  XNOR2_X1 U5831 ( .A(n4544), .B(n5097), .ZN(n7030) );
  NAND2_X1 U5832 ( .A1(n5502), .A2(n5501), .ZN(n4544) );
  XNOR2_X1 U5833 ( .A(n5531), .B(n5530), .ZN(n7024) );
  NOR2_X1 U5834 ( .A1(n5570), .A2(n4918), .ZN(n5593) );
  NOR2_X1 U5836 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n10636), .ZN(n8380) );
  NAND2_X1 U5837 ( .A1(n7750), .A2(n6747), .ZN(n7986) );
  AND4_X1 U5838 ( .A1(n6266), .A2(n6265), .A3(n6264), .A4(n6263), .ZN(n8088)
         );
  NAND2_X1 U5839 ( .A1(n8816), .A2(n9220), .ZN(n8786) );
  OR2_X1 U5840 ( .A1(n6860), .A2(n6863), .ZN(n8712) );
  INV_X1 U5841 ( .A(n5040), .ZN(n5039) );
  OAI21_X1 U5842 ( .B1(n8769), .B2(n5042), .A(n5041), .ZN(n5040) );
  AND2_X1 U5843 ( .A1(n5056), .A2(n5061), .ZN(n8711) );
  NAND2_X1 U5844 ( .A1(n8743), .A2(n6817), .ZN(n5056) );
  NAND2_X1 U5845 ( .A1(n8718), .A2(n6787), .ZN(n8736) );
  NAND2_X1 U5846 ( .A1(n8679), .A2(n6800), .ZN(n8770) );
  AOI21_X1 U5847 ( .B1(n4427), .B2(n5019), .A(n5017), .ZN(n5016) );
  INV_X1 U5848 ( .A(n8074), .ZN(n5017) );
  NAND2_X1 U5849 ( .A1(n6755), .A2(n7932), .ZN(n7935) );
  NAND2_X1 U5850 ( .A1(n7033), .A2(n6351), .ZN(n4546) );
  INV_X1 U5851 ( .A(n8712), .ZN(n8816) );
  OR2_X1 U5852 ( .A1(n6860), .A2(n6852), .ZN(n8821) );
  INV_X1 U5853 ( .A(n8818), .ZN(n8761) );
  AND2_X1 U5854 ( .A1(n5053), .A2(n5051), .ZN(n5050) );
  INV_X1 U5855 ( .A(n6892), .ZN(n5051) );
  NAND2_X1 U5856 ( .A1(n5052), .A2(n5053), .ZN(n6893) );
  NAND2_X1 U5857 ( .A1(n7522), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8818) );
  AOI21_X1 U5858 ( .B1(n4876), .B2(n6623), .A(n4820), .ZN(n6659) );
  OAI21_X1 U5859 ( .B1(n6657), .B2(n6658), .A(n4396), .ZN(n4820) );
  NAND2_X1 U5860 ( .A1(n4877), .A2(n4396), .ZN(n6656) );
  INV_X1 U5861 ( .A(n8992), .ZN(n8941) );
  OR2_X1 U5862 ( .A1(n7099), .A2(n10565), .ZN(n8832) );
  INV_X1 U5863 ( .A(n9092), .ZN(n9048) );
  AND4_X1 U5864 ( .A1(n6281), .A2(n6280), .A3(n6279), .A4(n6278), .ZN(n8914)
         );
  AND2_X1 U5865 ( .A1(n4677), .A2(n4676), .ZN(n4675) );
  NAND2_X1 U5866 ( .A1(n7269), .A2(n7268), .ZN(n7267) );
  NOR3_X1 U5867 ( .A1(n10510), .A2(n7263), .A3(n4643), .ZN(n7265) );
  AND2_X1 U5868 ( .A1(n4645), .A2(n7264), .ZN(n4643) );
  NAND2_X1 U5869 ( .A1(n7245), .A2(n4514), .ZN(n7149) );
  NAND2_X1 U5870 ( .A1(n4515), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n4514) );
  NAND2_X1 U5871 ( .A1(n7149), .A2(n7150), .ZN(n7148) );
  NAND2_X1 U5872 ( .A1(n7136), .A2(n4450), .ZN(n7138) );
  NAND2_X1 U5873 ( .A1(n7138), .A2(n7139), .ZN(n7161) );
  NAND2_X1 U5874 ( .A1(n7163), .A2(n7164), .ZN(n7175) );
  NAND2_X1 U5875 ( .A1(n7297), .A2(n4444), .ZN(n7315) );
  AOI21_X1 U5876 ( .B1(n7309), .B2(n7308), .A(n4417), .ZN(n7332) );
  NAND2_X1 U5877 ( .A1(n4649), .A2(n4653), .ZN(n7475) );
  NAND2_X1 U5878 ( .A1(n7309), .A2(n4654), .ZN(n4649) );
  INV_X1 U5879 ( .A(n4642), .ZN(n7759) );
  AND2_X1 U5880 ( .A1(n4642), .A2(n4641), .ZN(n7763) );
  NAND2_X1 U5881 ( .A1(n7761), .A2(n7760), .ZN(n4641) );
  INV_X1 U5882 ( .A(n4640), .ZN(n8549) );
  NAND2_X1 U5883 ( .A1(n8848), .A2(n4421), .ZN(n4743) );
  OAI21_X1 U5884 ( .B1(n4742), .B2(n4741), .A(n4413), .ZN(n8873) );
  NAND2_X1 U5885 ( .A1(n4421), .A2(n4745), .ZN(n4742) );
  INV_X1 U5886 ( .A(n8848), .ZN(n4741) );
  INV_X1 U5887 ( .A(n10511), .ZN(n10506) );
  NAND2_X1 U5888 ( .A1(n6484), .A2(n6483), .ZN(n8630) );
  INV_X1 U5889 ( .A(n8901), .ZN(n9241) );
  OR2_X1 U5890 ( .A1(n6450), .A2(n6868), .ZN(n8945) );
  NAND2_X1 U5891 ( .A1(n6466), .A2(n6465), .ZN(n9245) );
  NAND2_X1 U5892 ( .A1(n8968), .A2(n4490), .ZN(n9258) );
  NAND2_X1 U5893 ( .A1(n8402), .A2(n6351), .ZN(n6419) );
  NAND2_X1 U5894 ( .A1(n9038), .A2(n6587), .ZN(n9017) );
  NAND2_X1 U5895 ( .A1(n9046), .A2(n6583), .ZN(n9035) );
  NAND2_X1 U5896 ( .A1(n4857), .A2(n4858), .ZN(n9026) );
  NAND2_X1 U5897 ( .A1(n8923), .A2(n4859), .ZN(n4857) );
  INV_X1 U5898 ( .A(n8632), .ZN(n9067) );
  AND2_X1 U5899 ( .A1(n6362), .A2(n6361), .ZN(n9117) );
  NAND2_X1 U5900 ( .A1(n4835), .A2(n4834), .ZN(n9112) );
  NAND2_X1 U5901 ( .A1(n4547), .A2(n4401), .ZN(n4835) );
  NAND2_X1 U5902 ( .A1(n4547), .A2(n8916), .ZN(n9126) );
  OR2_X1 U5903 ( .A1(n9209), .A2(n8308), .ZN(n9338) );
  AND2_X1 U5904 ( .A1(n4844), .A2(n4841), .ZN(n8291) );
  INV_X1 U5905 ( .A(n8110), .ZN(n4841) );
  NAND2_X1 U5906 ( .A1(n8112), .A2(n8111), .ZN(n4844) );
  NAND2_X1 U5907 ( .A1(n4849), .A2(n6918), .ZN(n7809) );
  NAND2_X1 U5908 ( .A1(n7550), .A2(n4850), .ZN(n4849) );
  NAND2_X1 U5909 ( .A1(n7554), .A2(n6518), .ZN(n4658) );
  NAND2_X1 U5910 ( .A1(n5077), .A2(n6507), .ZN(n7553) );
  NAND2_X1 U5911 ( .A1(n6849), .A2(n7532), .ZN(n9188) );
  INV_X1 U5912 ( .A(n8974), .ZN(n9234) );
  INV_X1 U5913 ( .A(n10523), .ZN(n9190) );
  INV_X2 U5914 ( .A(n10603), .ZN(n10605) );
  CLKBUF_X1 U5915 ( .A(n10546), .Z(n10567) );
  INV_X1 U5916 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n8404) );
  INV_X1 U5917 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n8255) );
  XNOR2_X1 U5918 ( .A(n6678), .B(n6677), .ZN(n8256) );
  NAND2_X1 U5919 ( .A1(n6676), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6678) );
  INV_X1 U5920 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n9862) );
  INV_X1 U5921 ( .A(n6624), .ZN(n8535) );
  INV_X1 U5922 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n8532) );
  INV_X1 U5923 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n7707) );
  INV_X1 U5924 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n7632) );
  INV_X1 U5925 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n9860) );
  INV_X1 U5926 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n7307) );
  INV_X1 U5927 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n9873) );
  INV_X1 U5928 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n7034) );
  INV_X1 U5929 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n7031) );
  INV_X1 U5930 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n7025) );
  INV_X1 U5931 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n9741) );
  INV_X1 U5932 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n5118) );
  NAND2_X1 U5933 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_31__SCAN_IN), .ZN(
        n4735) );
  OAI21_X1 U5934 ( .B1(n7859), .B2(n4935), .A(n4424), .ZN(n8000) );
  NAND2_X1 U5935 ( .A1(n7859), .A2(n4936), .ZN(n4934) );
  INV_X1 U5936 ( .A(n4933), .ZN(n4936) );
  NAND2_X1 U5937 ( .A1(n9539), .A2(n5089), .ZN(n9404) );
  AND3_X1 U5938 ( .A1(n5453), .A2(n5452), .A3(n5451), .ZN(n10155) );
  AND4_X1 U5939 ( .A1(n5546), .A2(n5545), .A3(n5544), .A4(n5543), .ZN(n8026)
         );
  AND2_X1 U5940 ( .A1(n5381), .A2(n5380), .ZN(n10091) );
  NAND2_X1 U5941 ( .A1(n4923), .A2(n4926), .ZN(n8618) );
  INV_X1 U5942 ( .A(n4927), .ZN(n4926) );
  OAI21_X1 U5943 ( .B1(n4929), .B2(n4928), .A(n8598), .ZN(n4927) );
  AND4_X1 U5944 ( .A1(n5482), .A2(n5481), .A3(n5480), .A4(n5479), .ZN(n8327)
         );
  NAND2_X1 U5945 ( .A1(n9548), .A2(n9552), .ZN(n9472) );
  AND4_X1 U5946 ( .A1(n5471), .A2(n5470), .A3(n5469), .A4(n5468), .ZN(n8441)
         );
  NAND2_X1 U5947 ( .A1(n8318), .A2(n8275), .ZN(n4978) );
  AND2_X1 U5948 ( .A1(n5370), .A2(n5369), .ZN(n10074) );
  AND4_X1 U5949 ( .A1(n5515), .A2(n5514), .A3(n5513), .A4(n5512), .ZN(n8207)
         );
  OR2_X1 U5950 ( .A1(n7439), .A2(n10290), .ZN(n9494) );
  OR2_X1 U5951 ( .A1(n7439), .A2(n7366), .ZN(n9555) );
  AND2_X1 U5952 ( .A1(n7501), .A2(n7363), .ZN(n9532) );
  INV_X1 U5953 ( .A(n9555), .ZN(n9534) );
  INV_X1 U5954 ( .A(n9494), .ZN(n9553) );
  NAND2_X1 U5955 ( .A1(n8453), .A2(n9416), .ZN(n9551) );
  NAND2_X1 U5956 ( .A1(n8459), .A2(n8458), .ZN(n9552) );
  INV_X1 U5957 ( .A(n5720), .ZN(n9641) );
  INV_X1 U5958 ( .A(n10025), .ZN(n9570) );
  INV_X1 U5959 ( .A(n9721), .ZN(n9571) );
  INV_X1 U5960 ( .A(n10156), .ZN(n10104) );
  INV_X1 U5961 ( .A(n8202), .ZN(n9581) );
  NAND4_X1 U5962 ( .A1(n5589), .A2(n5588), .A3(n5587), .A4(n5586), .ZN(n9588)
         );
  INV_X1 U5963 ( .A(n7495), .ZN(n9589) );
  NAND2_X1 U5964 ( .A1(n5715), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n5613) );
  NAND4_X1 U5965 ( .A1(n5579), .A2(n5578), .A3(n5577), .A4(n5576), .ZN(n9590)
         );
  NAND2_X1 U5966 ( .A1(n7407), .A2(n4580), .ZN(n9596) );
  INV_X1 U5967 ( .A(n4581), .ZN(n4580) );
  AND2_X1 U5968 ( .A1(n7089), .A2(n7088), .ZN(n7184) );
  NAND2_X1 U5969 ( .A1(n7182), .A2(n7090), .ZN(n7091) );
  OR2_X1 U5970 ( .A1(n7226), .A2(n7093), .ZN(n7256) );
  AOI21_X1 U5971 ( .B1(n7220), .B2(n7084), .A(n7083), .ZN(n7219) );
  NOR2_X1 U5972 ( .A1(n7219), .A2(n7085), .ZN(n7250) );
  NAND2_X1 U5973 ( .A1(n7392), .A2(n7391), .ZN(n7394) );
  NAND2_X1 U5974 ( .A1(n4560), .A2(n7461), .ZN(n7463) );
  AND2_X1 U5975 ( .A1(n4560), .A2(n4558), .ZN(n7617) );
  AND2_X1 U5976 ( .A1(n7468), .A2(n7466), .ZN(n4702) );
  AND2_X1 U5977 ( .A1(n7467), .A2(n7466), .ZN(n7469) );
  OR2_X1 U5978 ( .A1(n4555), .A2(n7618), .ZN(n4554) );
  NAND2_X1 U5979 ( .A1(n7462), .A2(n4558), .ZN(n4553) );
  XNOR2_X1 U5980 ( .A(n9620), .B(n9621), .ZN(n10351) );
  NAND2_X1 U5981 ( .A1(n10351), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n10350) );
  AND2_X1 U5982 ( .A1(n4575), .A2(n4577), .ZN(n10394) );
  NAND2_X1 U5983 ( .A1(n4575), .A2(n4574), .ZN(n10392) );
  INV_X1 U5984 ( .A(n10248), .ZN(n9642) );
  NAND2_X1 U5985 ( .A1(n9647), .A2(n9646), .ZN(n4523) );
  NAND2_X1 U5986 ( .A1(n4690), .A2(n6875), .ZN(n6874) );
  INV_X1 U5987 ( .A(n6873), .ZN(n4690) );
  XNOR2_X1 U5988 ( .A(n9665), .B(n9669), .ZN(n10181) );
  NAND2_X1 U5989 ( .A1(n5026), .A2(n6050), .ZN(n9665) );
  OR2_X1 U5990 ( .A1(n9689), .A2(n9688), .ZN(n10184) );
  NAND2_X1 U5991 ( .A1(n9715), .A2(n5993), .ZN(n9698) );
  INV_X1 U5992 ( .A(n6057), .ZN(n10013) );
  AND2_X1 U5993 ( .A1(n10077), .A2(n10076), .ZN(n10211) );
  INV_X1 U5994 ( .A(n10217), .ZN(n10098) );
  NAND2_X1 U5995 ( .A1(n7904), .A2(n6019), .ZN(n8060) );
  OAI21_X1 U5996 ( .B1(n5744), .B2(n5743), .A(n5908), .ZN(n7887) );
  NAND2_X1 U5997 ( .A1(n7836), .A2(n6017), .ZN(n7890) );
  NAND2_X1 U5998 ( .A1(n4999), .A2(n6011), .ZN(n10414) );
  NAND2_X1 U5999 ( .A1(n7892), .A2(n7891), .ZN(n10424) );
  INV_X1 U6000 ( .A(n10424), .ZN(n10142) );
  XNOR2_X1 U6001 ( .A(n7790), .B(n4784), .ZN(n10442) );
  INV_X1 U6002 ( .A(n7979), .ZN(n7529) );
  INV_X1 U6003 ( .A(n10114), .ZN(n10270) );
  INV_X1 U6004 ( .A(n8450), .ZN(n9423) );
  INV_X1 U6005 ( .A(n10434), .ZN(n10435) );
  AND2_X1 U6006 ( .A1(n4520), .A2(n5952), .ZN(n10428) );
  AND2_X1 U6007 ( .A1(n5253), .A2(n5258), .ZN(n4616) );
  INV_X1 U6008 ( .A(n5289), .ZN(n10285) );
  OR2_X1 U6009 ( .A1(n5947), .A2(n5946), .ZN(n5948) );
  INV_X1 U6010 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n8332) );
  INV_X1 U6011 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n7995) );
  INV_X1 U6012 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n9929) );
  INV_X1 U6013 ( .A(n6949), .ZN(n7930) );
  INV_X1 U6014 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n7808) );
  INV_X1 U6015 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n7709) );
  INV_X1 U6016 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n7653) );
  INV_X1 U6017 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n7507) );
  INV_X1 U6018 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n7456) );
  OR3_X1 U6019 ( .A1(n5473), .A2(P1_IR_REG_13__SCAN_IN), .A3(
        P1_IR_REG_12__SCAN_IN), .ZN(n5461) );
  INV_X1 U6020 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n7274) );
  INV_X1 U6021 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n7079) );
  INV_X1 U6022 ( .A(n7622), .ZN(n7460) );
  INV_X1 U6023 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n7035) );
  INV_X1 U6024 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n7026) );
  INV_X1 U6025 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n7014) );
  XNOR2_X1 U6026 ( .A(n5641), .B(n5640), .ZN(n7185) );
  XNOR2_X1 U6027 ( .A(n5677), .B(P1_IR_REG_6__SCAN_IN), .ZN(n7087) );
  AND2_X1 U6028 ( .A1(n5676), .A2(n5652), .ZN(n9595) );
  AND3_X1 U6029 ( .A1(n4699), .A2(n4698), .A3(n4697), .ZN(n7059) );
  NAND2_X1 U6030 ( .A1(n4918), .A2(n5249), .ZN(n4697) );
  INV_X1 U6031 ( .A(n5570), .ZN(n4699) );
  NAND2_X1 U6032 ( .A1(n5569), .A2(P1_IR_REG_2__SCAN_IN), .ZN(n4698) );
  OAI21_X1 U6033 ( .B1(n7001), .B2(n5620), .A(n5619), .ZN(n5621) );
  AOI21_X1 U6034 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(P1_ADDR_REG_10__SCAN_IN), 
        .A(n10632), .ZN(n10631) );
  NOR2_X1 U6035 ( .A1(n10631), .A2(n10630), .ZN(n10629) );
  AOI21_X1 U6036 ( .B1(P2_ADDR_REG_11__SCAN_IN), .B2(P1_ADDR_REG_11__SCAN_IN), 
        .A(n10629), .ZN(n10628) );
  OAI21_X1 U6037 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(P2_ADDR_REG_12__SCAN_IN), 
        .A(n10626), .ZN(n10624) );
  INV_X1 U6038 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n8560) );
  AOI21_X1 U6039 ( .B1(n4748), .B2(n6625), .A(n4747), .ZN(n4746) );
  NAND2_X1 U6040 ( .A1(n4635), .A2(n7706), .ZN(n4634) );
  OAI21_X1 U6041 ( .B1(n8863), .B2(n8560), .A(n8559), .ZN(n4747) );
  OR2_X1 U6042 ( .A1(n10605), .A2(n4681), .ZN(n4680) );
  NAND2_X1 U6043 ( .A1(n9365), .A2(n10605), .ZN(n4682) );
  INV_X1 U6044 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n4681) );
  NAND2_X1 U6045 ( .A1(n10598), .A2(n10583), .ZN(n4870) );
  INV_X1 U6046 ( .A(n4869), .ZN(n4868) );
  OAI21_X1 U6047 ( .B1(n4425), .B2(n10596), .A(n4871), .ZN(n4869) );
  NAND2_X1 U6048 ( .A1(n9498), .A2(n4521), .ZN(P1_U3227) );
  AND2_X1 U6049 ( .A1(n9497), .A2(n4492), .ZN(n4521) );
  NOR2_X1 U6050 ( .A1(n5957), .A2(n4716), .ZN(n4715) );
  NAND2_X1 U6051 ( .A1(n4587), .A2(n4585), .ZN(n9634) );
  OAI21_X1 U6052 ( .B1(n9631), .B2(n7629), .A(n4586), .ZN(n4585) );
  INV_X1 U6053 ( .A(n4588), .ZN(n4587) );
  OAI22_X1 U6054 ( .A1(n6691), .A2(n10275), .B1(n10492), .B2(n6085), .ZN(n6086) );
  NAND2_X1 U6055 ( .A1(n8619), .A2(n6889), .ZN(n6890) );
  OR2_X1 U6056 ( .A1(n6624), .A2(n6499), .ZN(n4397) );
  INV_X1 U6057 ( .A(n8844), .ZN(n6911) );
  INV_X1 U6058 ( .A(n7894), .ZN(n4758) );
  AND2_X1 U6059 ( .A1(n4901), .A2(n4900), .ZN(n4398) );
  XNOR2_X2 U6060 ( .A(n5727), .B(P1_IR_REG_21__SCAN_IN), .ZN(n6949) );
  INV_X1 U6061 ( .A(n6817), .ZN(n5059) );
  AND2_X1 U6062 ( .A1(n8059), .A2(n5047), .ZN(n4399) );
  OR2_X1 U6063 ( .A1(n9312), .A2(n9147), .ZN(n4400) );
  AND2_X1 U6064 ( .A1(n4400), .A2(n8916), .ZN(n4401) );
  AND2_X1 U6065 ( .A1(n6138), .A2(n6137), .ZN(n4402) );
  INV_X1 U6066 ( .A(n9502), .ZN(n4959) );
  AND2_X1 U6067 ( .A1(n4399), .A2(n4438), .ZN(n4403) );
  INV_X1 U6068 ( .A(n6051), .ZN(n4709) );
  OR2_X1 U6069 ( .A1(n8473), .A2(n4943), .ZN(n4404) );
  NAND2_X1 U6070 ( .A1(n5908), .A2(n4807), .ZN(n4809) );
  INV_X1 U6071 ( .A(n4809), .ZN(n4628) );
  AND2_X1 U6072 ( .A1(n5250), .A2(n5261), .ZN(n4405) );
  AND2_X1 U6073 ( .A1(n4462), .A2(n4757), .ZN(n7850) );
  AND2_X1 U6074 ( .A1(n6378), .A2(n6377), .ZN(n9086) );
  INV_X1 U6075 ( .A(n9086), .ZN(n9296) );
  NAND2_X1 U6076 ( .A1(n5836), .A2(n7994), .ZN(n4406) );
  NAND2_X1 U6077 ( .A1(n5037), .A2(n6786), .ZN(n8718) );
  AND2_X1 U6078 ( .A1(n4984), .A2(n4983), .ZN(n4407) );
  AND2_X1 U6079 ( .A1(n7335), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n4408) );
  INV_X1 U6080 ( .A(n6010), .ZN(n7924) );
  AND2_X1 U6081 ( .A1(n5610), .A2(n5609), .ZN(n6010) );
  NAND2_X1 U6082 ( .A1(n7894), .A2(n7850), .ZN(n5855) );
  INV_X1 U6083 ( .A(n5855), .ZN(n4811) );
  AND2_X1 U6084 ( .A1(n9197), .A2(n8912), .ZN(n4409) );
  AND2_X1 U6085 ( .A1(n5347), .A2(n4721), .ZN(n4410) );
  AND2_X1 U6086 ( .A1(n4904), .A2(n4903), .ZN(n4411) );
  NOR2_X1 U6087 ( .A1(n6109), .A2(P2_IR_REG_29__SCAN_IN), .ZN(n4412) );
  INV_X1 U6088 ( .A(n9197), .ZN(n4798) );
  INV_X1 U6089 ( .A(n9027), .ZN(n4856) );
  OR2_X1 U6090 ( .A1(n8537), .A2(n8874), .ZN(n4413) );
  NOR2_X1 U6091 ( .A1(n10378), .A2(n4576), .ZN(n4414) );
  OR2_X1 U6092 ( .A1(n7393), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n4415) );
  INV_X1 U6093 ( .A(n5346), .ZN(n6053) );
  INV_X2 U6094 ( .A(n8593), .ZN(n6956) );
  NAND2_X1 U6095 ( .A1(n8690), .A2(n6920), .ZN(n4416) );
  NAND2_X1 U6096 ( .A1(n8962), .A2(n6607), .ZN(n8989) );
  NAND2_X1 U6097 ( .A1(n6275), .A2(n6274), .ZN(n9331) );
  NAND2_X1 U6098 ( .A1(n9551), .A2(n9550), .ZN(n9548) );
  AND2_X1 U6099 ( .A1(n7299), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n4417) );
  INV_X1 U6100 ( .A(n6510), .ZN(n4660) );
  NAND2_X1 U6101 ( .A1(n5646), .A2(n5606), .ZN(n4418) );
  NAND2_X1 U6102 ( .A1(n8195), .A2(n8196), .ZN(n4419) );
  AND2_X1 U6103 ( .A1(n6620), .A2(n6619), .ZN(n4420) );
  INV_X1 U6104 ( .A(n8520), .ZN(n4960) );
  NAND2_X1 U6105 ( .A1(n5701), .A2(n5700), .ZN(n6058) );
  AND2_X1 U6106 ( .A1(n8541), .A2(n4744), .ZN(n4421) );
  OR4_X1 U6107 ( .A1(n5941), .A2(n9632), .A3(n5940), .A4(n5953), .ZN(n4422) );
  NAND3_X1 U6108 ( .A1(n6604), .A2(n8941), .A3(n6603), .ZN(n6605) );
  OR2_X1 U6109 ( .A1(n10178), .A2(n9567), .ZN(n4423) );
  AND2_X1 U6110 ( .A1(n7877), .A2(n4932), .ZN(n4424) );
  INV_X1 U6111 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n6170) );
  INV_X1 U6112 ( .A(n8521), .ZN(n4962) );
  AND2_X1 U6113 ( .A1(n5570), .A2(n5250), .ZN(n5456) );
  NAND2_X2 U6114 ( .A1(n6174), .A2(n6173), .ZN(n8759) );
  XNOR2_X1 U6115 ( .A(n5167), .B(SI_14_), .ZN(n5454) );
  NAND2_X1 U6116 ( .A1(n6032), .A2(n6031), .ZN(n10124) );
  AND2_X1 U6117 ( .A1(n9264), .A2(n9263), .ZN(n4425) );
  INV_X1 U6118 ( .A(n6951), .ZN(n4911) );
  AND2_X1 U6119 ( .A1(n7478), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n4426) );
  AND2_X1 U6120 ( .A1(n8075), .A2(n5018), .ZN(n4427) );
  AND2_X1 U6121 ( .A1(n4599), .A2(n5194), .ZN(n4428) );
  AND3_X1 U6122 ( .A1(n7680), .A2(n10575), .A3(n10579), .ZN(n4429) );
  AND2_X1 U6123 ( .A1(n6139), .A2(n4836), .ZN(n4430) );
  AND2_X1 U6124 ( .A1(n6602), .A2(n4394), .ZN(n4431) );
  INV_X1 U6125 ( .A(n8275), .ZN(n4971) );
  INV_X1 U6126 ( .A(n8066), .ZN(n4900) );
  NAND2_X1 U6127 ( .A1(n5895), .A2(n5896), .ZN(n6051) );
  AND2_X1 U6128 ( .A1(n6518), .A2(n7779), .ZN(n4432) );
  INV_X1 U6129 ( .A(n9198), .ZN(n4667) );
  AND2_X1 U6130 ( .A1(n5678), .A2(n7185), .ZN(n4433) );
  NOR2_X1 U6131 ( .A1(n4625), .A2(n4622), .ZN(n5273) );
  AND2_X1 U6132 ( .A1(n9312), .A2(n9147), .ZN(n4434) );
  AND2_X1 U6133 ( .A1(n5999), .A2(n5837), .ZN(n6875) );
  AND3_X1 U6134 ( .A1(n5504), .A2(n5249), .A3(n5640), .ZN(n4435) );
  AND3_X1 U6135 ( .A1(n6023), .A2(n5045), .A3(n6024), .ZN(n4436) );
  OR2_X1 U6136 ( .A1(n5059), .A2(n6818), .ZN(n4437) );
  AND2_X1 U6137 ( .A1(n8170), .A2(n8167), .ZN(n4438) );
  AND2_X1 U6138 ( .A1(n4941), .A2(n8458), .ZN(n4439) );
  OR2_X1 U6139 ( .A1(n5382), .A2(n5188), .ZN(n4440) );
  NAND3_X1 U6140 ( .A1(n6883), .A2(n10418), .A3(n6882), .ZN(n4442) );
  INV_X1 U6141 ( .A(n10111), .ZN(n4604) );
  AND2_X1 U6142 ( .A1(n4582), .A2(n7051), .ZN(n4443) );
  INV_X1 U6143 ( .A(n5022), .ZN(n10108) );
  AOI21_X1 U6144 ( .B1(n10124), .B2(n6033), .A(n5025), .ZN(n5022) );
  OR2_X1 U6145 ( .A1(n7298), .A2(n9796), .ZN(n4444) );
  NAND2_X1 U6146 ( .A1(n5890), .A2(n5993), .ZN(n4445) );
  INV_X1 U6147 ( .A(n10190), .ZN(n9708) );
  AND2_X1 U6148 ( .A1(n4743), .A2(n8537), .ZN(n4446) );
  INV_X1 U6149 ( .A(n5085), .ZN(n4977) );
  INV_X1 U6150 ( .A(n4860), .ZN(n4859) );
  NAND2_X1 U6151 ( .A1(n5105), .A2(n8922), .ZN(n4860) );
  NAND2_X1 U6152 ( .A1(n9075), .A2(n8925), .ZN(n4447) );
  NAND2_X1 U6153 ( .A1(n8520), .A2(n4962), .ZN(n4448) );
  INV_X1 U6154 ( .A(n9261), .ZN(n8987) );
  NAND2_X1 U6155 ( .A1(n6439), .A2(n6438), .ZN(n9261) );
  INV_X1 U6156 ( .A(n8989), .ZN(n8980) );
  OR2_X1 U6157 ( .A1(n5025), .A2(n5021), .ZN(n4449) );
  AND2_X1 U6158 ( .A1(n5680), .A2(n5679), .ZN(n7867) );
  AND2_X1 U6159 ( .A1(n5980), .A2(n10151), .ZN(n8337) );
  INV_X1 U6160 ( .A(n8337), .ZN(n4782) );
  OR2_X1 U6161 ( .A1(n7137), .A2(n7679), .ZN(n4450) );
  AND2_X1 U6162 ( .A1(n7066), .A2(n7064), .ZN(n4451) );
  INV_X1 U6163 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n5249) );
  INV_X1 U6164 ( .A(n10042), .ZN(n10022) );
  AND2_X1 U6165 ( .A1(n5345), .A2(n5344), .ZN(n10042) );
  AND2_X1 U6166 ( .A1(n5928), .A2(n5997), .ZN(n5995) );
  INV_X1 U6167 ( .A(n5995), .ZN(n9683) );
  INV_X1 U6168 ( .A(n4823), .ZN(n4822) );
  NAND2_X1 U6169 ( .A1(n10070), .A2(n5989), .ZN(n4823) );
  AND2_X1 U6170 ( .A1(n4857), .A2(n4855), .ZN(n4452) );
  AND2_X1 U6171 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), .ZN(
        n4453) );
  AND2_X1 U6172 ( .A1(n9065), .A2(n6581), .ZN(n4454) );
  OR2_X1 U6173 ( .A1(n9636), .A2(n10236), .ZN(n4455) );
  AND2_X1 U6174 ( .A1(n9347), .A2(n9221), .ZN(n4456) );
  NAND2_X1 U6175 ( .A1(n10350), .A2(n9622), .ZN(n10365) );
  AND2_X1 U6176 ( .A1(n5877), .A2(n5850), .ZN(n4457) );
  NAND2_X1 U6177 ( .A1(n6815), .A2(n6816), .ZN(n5061) );
  INV_X1 U6178 ( .A(n4655), .ZN(n4654) );
  NAND2_X1 U6179 ( .A1(n4657), .A2(n4656), .ZN(n4655) );
  OAI21_X1 U6180 ( .B1(n5695), .B2(n5028), .A(n4423), .ZN(n5027) );
  OR2_X1 U6181 ( .A1(n4774), .A2(n4782), .ZN(n4458) );
  INV_X1 U6182 ( .A(n4957), .ZN(n4956) );
  NAND2_X1 U6183 ( .A1(n4961), .A2(n4958), .ZN(n4957) );
  AND3_X1 U6184 ( .A1(n5695), .A2(n5694), .A3(n5995), .ZN(n4459) );
  OR2_X1 U6185 ( .A1(n9257), .A2(n10590), .ZN(n4460) );
  AND2_X1 U6186 ( .A1(n4889), .A2(n5454), .ZN(n4461) );
  AND3_X1 U6187 ( .A1(n5636), .A2(n5635), .A3(n5637), .ZN(n4462) );
  AND2_X1 U6188 ( .A1(n4850), .A2(n4416), .ZN(n4463) );
  NOR2_X1 U6189 ( .A1(n5962), .A2(n10048), .ZN(n4464) );
  AND2_X1 U6190 ( .A1(n6548), .A2(n9198), .ZN(n8299) );
  OR2_X1 U6191 ( .A1(n4660), .A2(n4397), .ZN(n4465) );
  NOR2_X1 U6192 ( .A1(n8735), .A2(n5036), .ZN(n4466) );
  AND2_X1 U6193 ( .A1(n8338), .A2(n5850), .ZN(n8216) );
  AND2_X1 U6194 ( .A1(n5043), .A2(n6800), .ZN(n4467) );
  NOR2_X1 U6195 ( .A1(P1_IR_REG_28__SCAN_IN), .A2(P1_IR_REG_29__SCAN_IN), .ZN(
        n4468) );
  INV_X1 U6196 ( .A(n7325), .ZN(n4996) );
  AND2_X1 U6197 ( .A1(n8989), .A2(n8979), .ZN(n4469) );
  AND2_X1 U6198 ( .A1(n5904), .A2(n8130), .ZN(n4470) );
  NAND2_X1 U6199 ( .A1(n8927), .A2(n6417), .ZN(n9027) );
  INV_X1 U6200 ( .A(n6017), .ZN(n5006) );
  AND2_X1 U6201 ( .A1(n4941), .A2(n9550), .ZN(n4471) );
  NAND2_X1 U6202 ( .A1(n10475), .A2(n9584), .ZN(n4472) );
  AND2_X1 U6203 ( .A1(n10143), .A2(n5982), .ZN(n4473) );
  AND2_X1 U6204 ( .A1(n7233), .A2(n4784), .ZN(n4474) );
  AND2_X1 U6205 ( .A1(n6774), .A2(n6767), .ZN(n4475) );
  AND2_X1 U6206 ( .A1(n6529), .A2(n6229), .ZN(n4476) );
  INV_X1 U6207 ( .A(n8919), .ZN(n4833) );
  AND2_X1 U6208 ( .A1(n9054), .A2(n6591), .ZN(n4477) );
  AND2_X1 U6209 ( .A1(n4790), .A2(n4795), .ZN(n4478) );
  AND2_X1 U6210 ( .A1(n4825), .A2(n4442), .ZN(n4479) );
  AND2_X1 U6211 ( .A1(n6044), .A2(n5012), .ZN(n4480) );
  INV_X1 U6212 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n5832) );
  AND2_X1 U6213 ( .A1(n5034), .A2(n5033), .ZN(n4481) );
  AND2_X1 U6214 ( .A1(n4946), .A2(n4949), .ZN(n4482) );
  NAND2_X1 U6215 ( .A1(n4861), .A2(n4862), .ZN(n4483) );
  AND2_X1 U6216 ( .A1(n4965), .A2(n4972), .ZN(n4967) );
  NAND2_X1 U6217 ( .A1(n4822), .A2(n4821), .ZN(n4484) );
  INV_X1 U6218 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n6118) );
  INV_X2 U6219 ( .A(n10148), .ZN(n10123) );
  NAND2_X1 U6220 ( .A1(n5330), .A2(n5329), .ZN(n9729) );
  INV_X1 U6221 ( .A(n9729), .ZN(n4503) );
  AND2_X1 U6222 ( .A1(n9127), .A2(n4988), .ZN(n4485) );
  NAND2_X1 U6223 ( .A1(n7837), .A2(n4758), .ZN(n7965) );
  NAND2_X1 U6224 ( .A1(n7935), .A2(n6759), .ZN(n8076) );
  INV_X2 U6225 ( .A(n10596), .ZN(n10598) );
  NAND2_X1 U6226 ( .A1(n4689), .A2(n6018), .ZN(n7961) );
  NAND2_X1 U6227 ( .A1(n8093), .A2(n6537), .ZN(n8113) );
  NAND2_X1 U6228 ( .A1(n4658), .A2(n6637), .ZN(n7778) );
  NAND2_X1 U6229 ( .A1(n4837), .A2(n4838), .ZN(n9229) );
  INV_X1 U6230 ( .A(n5993), .ZN(n4611) );
  AND2_X1 U6231 ( .A1(n8913), .A2(n8912), .ZN(n4486) );
  INV_X1 U6232 ( .A(n9286), .ZN(n4548) );
  NAND2_X1 U6233 ( .A1(n5296), .A2(n5295), .ZN(n10178) );
  INV_X1 U6234 ( .A(n10178), .ZN(n4903) );
  NAND2_X1 U6235 ( .A1(n6371), .A2(n6370), .ZN(n9301) );
  INV_X1 U6236 ( .A(n9301), .ZN(n4990) );
  NAND2_X1 U6237 ( .A1(n6922), .A2(n6924), .ZN(n8112) );
  NAND2_X1 U6238 ( .A1(n6768), .A2(n6767), .ZN(n8654) );
  NAND2_X1 U6239 ( .A1(n4541), .A2(n6171), .ZN(n4487) );
  OR2_X1 U6240 ( .A1(n8969), .A2(n9205), .ZN(n4488) );
  NAND2_X1 U6241 ( .A1(n4863), .A2(n8294), .ZN(n8913) );
  XNOR2_X1 U6242 ( .A(n5202), .B(SI_21_), .ZN(n5360) );
  NAND2_X1 U6243 ( .A1(n4398), .A2(n4899), .ZN(n4902) );
  AND2_X1 U6244 ( .A1(n8097), .A2(n4407), .ZN(n4489) );
  INV_X1 U6245 ( .A(n6950), .ZN(n7994) );
  AND2_X1 U6246 ( .A1(n8967), .A2(n4488), .ZN(n4490) );
  INV_X1 U6247 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n6285) );
  NOR2_X1 U6248 ( .A1(n7965), .A2(n10475), .ZN(n7907) );
  AND2_X1 U6249 ( .A1(n5238), .A2(n9775), .ZN(n4491) );
  OR2_X1 U6250 ( .A1(n4503), .A2(n9556), .ZN(n4492) );
  INV_X1 U6251 ( .A(n7618), .ZN(n4563) );
  AND2_X1 U6252 ( .A1(n4978), .A2(n4977), .ZN(n4493) );
  AND2_X1 U6253 ( .A1(n7335), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n4494) );
  AND2_X1 U6254 ( .A1(n4558), .A2(n4563), .ZN(n4495) );
  NAND2_X1 U6255 ( .A1(n5374), .A2(n5373), .ZN(n10075) );
  INV_X1 U6256 ( .A(n10075), .ZN(n4897) );
  INV_X1 U6257 ( .A(n10243), .ZN(n10489) );
  AND3_X1 U6258 ( .A1(n4906), .A2(n4905), .A3(n6010), .ZN(n7837) );
  AND2_X1 U6259 ( .A1(n6001), .A2(n6000), .ZN(n10406) );
  INV_X1 U6260 ( .A(n10406), .ZN(n10101) );
  INV_X1 U6261 ( .A(n10418), .ZN(n10158) );
  OAI22_X1 U6262 ( .A1(n7790), .A2(n4784), .B1(n7802), .B2(n5737), .ZN(n7345)
         );
  INV_X1 U6263 ( .A(n9342), .ZN(n4983) );
  INV_X1 U6264 ( .A(n4577), .ZN(n4576) );
  NAND2_X1 U6265 ( .A1(n9626), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n4577) );
  INV_X1 U6266 ( .A(n10364), .ZN(n4571) );
  AND2_X1 U6267 ( .A1(n6975), .A2(n8421), .ZN(n4496) );
  INV_X1 U6268 ( .A(n8874), .ZN(n4745) );
  OR2_X1 U6269 ( .A1(n8881), .A2(n9918), .ZN(n4497) );
  AND2_X1 U6270 ( .A1(n4553), .A2(n4555), .ZN(n4498) );
  OR2_X1 U6271 ( .A1(n6478), .A2(n8908), .ZN(n4499) );
  INV_X1 U6272 ( .A(n10421), .ZN(n6055) );
  AND2_X1 U6273 ( .A1(n5654), .A2(n5653), .ZN(n10421) );
  NAND2_X1 U6274 ( .A1(n7414), .A2(n7064), .ZN(n4500) );
  INV_X1 U6275 ( .A(n4415), .ZN(n4562) );
  INV_X1 U6276 ( .A(n9733), .ZN(n9632) );
  AND2_X1 U6277 ( .A1(n7407), .A2(n7049), .ZN(n4501) );
  NAND2_X1 U6278 ( .A1(n4502), .A2(n4473), .ZN(n5984) );
  OAI21_X1 U6279 ( .B1(n5871), .B2(n7899), .A(n5851), .ZN(n5965) );
  NAND2_X2 U6280 ( .A1(n10020), .A2(n10021), .ZN(n9716) );
  AND2_X2 U6281 ( .A1(n4602), .A2(n4549), .ZN(n10020) );
  NAND2_X1 U6282 ( .A1(n5137), .A2(n5136), .ZN(n5548) );
  NAND2_X1 U6283 ( .A1(n9673), .A2(n5998), .ZN(n6876) );
  AND2_X2 U6284 ( .A1(n6057), .A2(n4503), .ZN(n9732) );
  NOR2_X2 U6285 ( .A1(n10014), .A2(n10201), .ZN(n6057) );
  OAI21_X1 U6286 ( .B1(n5730), .B2(n4504), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n5264) );
  NAND2_X1 U6287 ( .A1(n10492), .A2(n10240), .ZN(n10275) );
  NAND2_X1 U6288 ( .A1(n6030), .A2(n6029), .ZN(n10144) );
  NOR2_X1 U6289 ( .A1(n5729), .A2(n5260), .ZN(n4505) );
  NAND2_X1 U6290 ( .A1(n7919), .A2(n7920), .ZN(n4999) );
  NAND2_X1 U6291 ( .A1(n6026), .A2(n6025), .ZN(n8214) );
  NAND2_X1 U6292 ( .A1(n6046), .A2(n6045), .ZN(n9711) );
  NAND2_X1 U6293 ( .A1(n4530), .A2(n6028), .ZN(n8335) );
  NAND2_X1 U6294 ( .A1(n5003), .A2(n5004), .ZN(n4689) );
  NAND2_X1 U6295 ( .A1(n4824), .A2(n10489), .ZN(n4691) );
  OAI21_X1 U6296 ( .B1(n7961), .B2(n7962), .A(n4472), .ZN(n4688) );
  INV_X1 U6297 ( .A(n4505), .ZN(n4504) );
  NAND2_X2 U6298 ( .A1(n5863), .A2(n5862), .ZN(n7349) );
  AND2_X2 U6299 ( .A1(n6966), .A2(n7001), .ZN(n5591) );
  INV_X1 U6300 ( .A(n4688), .ZN(n7906) );
  INV_X1 U6301 ( .A(n8626), .ZN(n4824) );
  INV_X1 U6302 ( .A(n5575), .ZN(n7946) );
  NAND2_X1 U6303 ( .A1(n4998), .A2(n4999), .ZN(n10412) );
  NAND2_X1 U6304 ( .A1(n8214), .A2(n6027), .ZN(n4530) );
  NAND2_X1 U6305 ( .A1(n4691), .A2(n4479), .ZN(n6887) );
  NAND2_X1 U6306 ( .A1(n4506), .A2(n5068), .ZN(n9219) );
  NAND2_X2 U6307 ( .A1(n6537), .A2(n6540), .ZN(n8109) );
  INV_X1 U6308 ( .A(n8111), .ZN(n4839) );
  NOR2_X2 U6309 ( .A1(n9185), .A2(n9184), .ZN(n9183) );
  NAND3_X1 U6310 ( .A1(n5830), .A2(n4755), .A3(n4508), .ZN(n4614) );
  NAND4_X1 U6311 ( .A1(n5825), .A2(n5939), .A3(n5824), .A4(n5895), .ZN(n4508)
         );
  OR2_X1 U6312 ( .A1(n5750), .A2(n6950), .ZN(n4630) );
  AOI21_X1 U6313 ( .B1(n5761), .B2(n5760), .A(n5759), .ZN(n5764) );
  AOI21_X2 U6314 ( .B1(n7914), .B2(n5909), .A(n5740), .ZN(n10401) );
  BUF_X4 U6315 ( .A(n5567), .Z(n5592) );
  XNOR2_X2 U6316 ( .A(n5472), .B(n5099), .ZN(n7273) );
  NAND2_X1 U6317 ( .A1(n4896), .A2(n5137), .ZN(n5499) );
  NAND2_X1 U6318 ( .A1(n4513), .A2(n4511), .ZN(n4789) );
  OR2_X1 U6319 ( .A1(n6598), .A2(n4394), .ZN(n4512) );
  INV_X1 U6320 ( .A(n7120), .ZN(n4515) );
  NOR2_X1 U6321 ( .A1(n7334), .A2(n4494), .ZN(n7336) );
  AND2_X1 U6322 ( .A1(n6255), .A2(n8089), .ZN(n6256) );
  NAND2_X1 U6323 ( .A1(n4529), .A2(n4476), .ZN(n6533) );
  NAND2_X1 U6324 ( .A1(n4746), .A2(n4634), .ZN(P2_U3264) );
  OAI211_X1 U6325 ( .C1(n6557), .C2(n6556), .A(n9173), .B(n6555), .ZN(n6568)
         );
  OAI21_X1 U6326 ( .B1(n4806), .B2(n6547), .A(n4804), .ZN(n4803) );
  NAND3_X1 U6327 ( .A1(n6348), .A2(n5062), .A3(n5064), .ZN(n4664) );
  OAI21_X2 U6328 ( .B1(n5439), .B2(n5438), .A(n5174), .ZN(n5426) );
  AND2_X1 U6329 ( .A1(n6955), .A2(n6954), .ZN(n6960) );
  NAND2_X1 U6330 ( .A1(n7492), .A2(n7491), .ZN(n7728) );
  NAND2_X1 U6331 ( .A1(n8000), .A2(n7999), .ZN(n8152) );
  AND3_X2 U6332 ( .A1(n4623), .A2(n4624), .A3(n5250), .ZN(n4921) );
  NAND2_X1 U6333 ( .A1(n5114), .A2(n5565), .ZN(n4609) );
  NAND2_X1 U6334 ( .A1(n4522), .A2(n5127), .ZN(n5674) );
  NOR2_X1 U6335 ( .A1(n4464), .A2(n4550), .ZN(n4549) );
  AND2_X1 U6336 ( .A1(n5126), .A2(n5604), .ZN(n4608) );
  NAND2_X1 U6337 ( .A1(n6888), .A2(n9666), .ZN(n6883) );
  NAND2_X1 U6338 ( .A1(n4898), .A2(n4897), .ZN(n10076) );
  NAND2_X1 U6339 ( .A1(n10057), .A2(n6053), .ZN(n10014) );
  NAND2_X1 U6340 ( .A1(n9637), .A2(n9636), .ZN(n9645) );
  NAND2_X1 U6341 ( .A1(n4608), .A2(n5605), .ZN(n4522) );
  NAND2_X1 U6342 ( .A1(n10176), .A2(n4455), .ZN(P1_U3553) );
  INV_X1 U6343 ( .A(n10092), .ZN(n4898) );
  NOR2_X2 U6344 ( .A1(n10076), .A2(n10061), .ZN(n10057) );
  INV_X1 U6345 ( .A(n6462), .ZN(n5076) );
  INV_X1 U6346 ( .A(n6306), .ZN(n5063) );
  NAND2_X1 U6347 ( .A1(n6592), .A2(n4477), .ZN(n6594) );
  AND2_X1 U6348 ( .A1(n6594), .A2(n6593), .ZN(n6596) );
  NAND2_X1 U6349 ( .A1(n4609), .A2(n5116), .ZN(n5605) );
  OAI21_X1 U6350 ( .B1(n4815), .B2(n4812), .A(n4454), .ZN(n6592) );
  AOI21_X1 U6351 ( .B1(n6545), .B2(n6544), .A(n6543), .ZN(n4806) );
  INV_X1 U6352 ( .A(n6519), .ZN(n4827) );
  NAND3_X1 U6353 ( .A1(n6526), .A2(n7817), .A3(n4465), .ZN(n4529) );
  INV_X1 U6354 ( .A(n6575), .ZN(n4814) );
  AND2_X2 U6355 ( .A1(n10087), .A2(n5776), .ZN(n10111) );
  NAND3_X1 U6356 ( .A1(n4531), .A2(n4484), .A3(n5990), .ZN(n4602) );
  NAND2_X1 U6357 ( .A1(n10102), .A2(n4603), .ZN(n4531) );
  NAND2_X1 U6358 ( .A1(n7541), .A2(n6160), .ZN(n5077) );
  NAND2_X1 U6359 ( .A1(n5977), .A2(n5976), .ZN(n8175) );
  NAND2_X1 U6360 ( .A1(n5969), .A2(n5968), .ZN(n4783) );
  NAND2_X1 U6361 ( .A1(n7467), .A2(n4702), .ZN(n7624) );
  NAND2_X1 U6362 ( .A1(n7092), .A2(n7225), .ZN(n7226) );
  NOR2_X1 U6363 ( .A1(n4695), .A2(n4694), .ZN(n4693) );
  NAND2_X1 U6364 ( .A1(n8018), .A2(n8017), .ZN(n8193) );
  NAND2_X1 U6365 ( .A1(n7431), .A2(n7430), .ZN(n7447) );
  OAI21_X2 U6366 ( .B1(n9500), .B2(n4960), .A(n4956), .ZN(n9424) );
  INV_X1 U6367 ( .A(n5254), .ZN(n4922) );
  NAND2_X1 U6369 ( .A1(n9500), .A2(n4953), .ZN(n4952) );
  NAND2_X1 U6370 ( .A1(n8524), .A2(n8523), .ZN(n9425) );
  NAND2_X1 U6371 ( .A1(n4938), .A2(n4937), .ZN(n8492) );
  AND2_X4 U6372 ( .A1(n5289), .A2(n5288), .ZN(n5705) );
  NAND2_X1 U6373 ( .A1(n4754), .A2(n4626), .ZN(n5745) );
  NAND2_X1 U6374 ( .A1(n4633), .A2(n4761), .ZN(n5825) );
  INV_X1 U6375 ( .A(n5825), .ZN(n5823) );
  NAND2_X1 U6376 ( .A1(n9219), .A2(n4666), .ZN(n6307) );
  NOR2_X1 U6377 ( .A1(n7552), .A2(n4542), .ZN(n4663) );
  NAND2_X1 U6378 ( .A1(n7712), .A2(n6503), .ZN(n7552) );
  NAND2_X1 U6379 ( .A1(n9118), .A2(n6571), .ZN(n9104) );
  NAND2_X1 U6380 ( .A1(n9002), .A2(n6629), .ZN(n8961) );
  INV_X1 U6381 ( .A(n5070), .ZN(n5069) );
  NAND2_X2 U6382 ( .A1(n6247), .A2(n6246), .ZN(n8243) );
  NAND2_X2 U6383 ( .A1(n9090), .A2(n6395), .ZN(n9043) );
  XNOR2_X2 U6384 ( .A(n5414), .B(n5413), .ZN(n7631) );
  AOI21_X2 U6385 ( .B1(n8910), .B2(n9225), .A(n8909), .ZN(n9250) );
  INV_X1 U6386 ( .A(n8290), .ZN(n4843) );
  NAND2_X1 U6387 ( .A1(n4682), .A2(n4680), .ZN(P2_U3548) );
  INV_X1 U6388 ( .A(n4842), .ZN(n4840) );
  NAND2_X1 U6389 ( .A1(n4460), .A2(n4685), .ZN(n4684) );
  NAND2_X1 U6390 ( .A1(n4788), .A2(n5695), .ZN(n9673) );
  AOI21_X2 U6391 ( .B1(n8175), .B2(n8174), .A(n5978), .ZN(n8215) );
  INV_X1 U6392 ( .A(n6876), .ZN(n4787) );
  OAI21_X1 U6393 ( .B1(n6887), .B2(n10168), .A(n5088), .ZN(n6886) );
  OAI21_X1 U6394 ( .B1(n6887), .B2(n10490), .A(n5094), .ZN(n6891) );
  NAND2_X1 U6395 ( .A1(n9260), .A2(n4683), .ZN(n9365) );
  INV_X1 U6396 ( .A(n8623), .ZN(n4825) );
  NAND2_X1 U6397 ( .A1(n4893), .A2(n5161), .ZN(n5472) );
  NOR2_X2 U6398 ( .A1(n5840), .A2(n5839), .ZN(n5845) );
  INV_X1 U6399 ( .A(n5359), .ZN(n4607) );
  OAI21_X1 U6400 ( .B1(n4422), .B2(n5956), .A(n4717), .ZN(n4716) );
  NAND2_X1 U6401 ( .A1(n4614), .A2(n5903), .ZN(n4613) );
  NAND2_X1 U6402 ( .A1(n4613), .A2(n4470), .ZN(n4612) );
  INV_X1 U6403 ( .A(n4969), .ZN(n4965) );
  NAND2_X1 U6404 ( .A1(n7462), .A2(n4495), .ZN(n4552) );
  NAND2_X1 U6405 ( .A1(n4552), .A2(n4554), .ZN(n9616) );
  NAND2_X1 U6406 ( .A1(n4564), .A2(n4565), .ZN(n9629) );
  NAND2_X1 U6407 ( .A1(n10365), .A2(n4571), .ZN(n4570) );
  INV_X1 U6408 ( .A(n7048), .ZN(n4582) );
  NAND2_X1 U6409 ( .A1(n9597), .A2(n7049), .ZN(n4581) );
  INV_X1 U6410 ( .A(n7405), .ZN(n4583) );
  NAND2_X1 U6411 ( .A1(n5426), .A2(n4428), .ZN(n4596) );
  NAND2_X1 U6412 ( .A1(n4596), .A2(n4597), .ZN(n5371) );
  NAND2_X1 U6413 ( .A1(n5484), .A2(n4461), .ZN(n4605) );
  OAI21_X2 U6414 ( .B1(n5517), .B2(n4728), .A(n5156), .ZN(n5484) );
  NAND2_X1 U6415 ( .A1(n9701), .A2(n5996), .ZN(n9685) );
  NAND3_X1 U6416 ( .A1(n4785), .A2(n6005), .A3(n5862), .ZN(n7914) );
  NAND2_X1 U6417 ( .A1(n4612), .A2(n4715), .ZN(P1_U3240) );
  NAND4_X1 U6418 ( .A1(n5258), .A2(n5257), .A3(n5256), .A4(n5255), .ZN(n5729)
         );
  NAND4_X1 U6419 ( .A1(n5253), .A2(n5458), .A3(n5251), .A4(n5252), .ZN(n5254)
         );
  NAND4_X1 U6420 ( .A1(n4617), .A2(n4616), .A3(n4615), .A4(n4468), .ZN(n4622)
         );
  NAND3_X1 U6422 ( .A1(n4765), .A2(n5751), .A3(n4630), .ZN(n4629) );
  NAND3_X1 U6423 ( .A1(n5786), .A2(n4632), .A3(n4631), .ZN(n5781) );
  NAND4_X1 U6424 ( .A1(n5819), .A2(n5818), .A3(n5998), .A4(n6875), .ZN(n4633)
         );
  NAND2_X1 U6425 ( .A1(n7309), .A2(n4650), .ZN(n4647) );
  NAND2_X1 U6426 ( .A1(n4647), .A2(n4648), .ZN(n7636) );
  INV_X1 U6427 ( .A(n7636), .ZN(n7634) );
  AOI21_X2 U6428 ( .B1(n7554), .B2(n4432), .A(n4659), .ZN(n7818) );
  NAND2_X1 U6429 ( .A1(n5077), .A2(n4663), .ZN(n7554) );
  NAND3_X1 U6430 ( .A1(n4665), .A2(n6350), .A3(n4664), .ZN(n9134) );
  NAND3_X1 U6431 ( .A1(n6307), .A2(n6348), .A3(n5062), .ZN(n4665) );
  NAND2_X1 U6432 ( .A1(n9046), .A2(n4672), .ZN(n4669) );
  NAND2_X1 U6433 ( .A1(n4669), .A2(n4670), .ZN(n9002) );
  INV_X1 U6434 ( .A(n6122), .ZN(n4679) );
  NAND3_X1 U6435 ( .A1(n6124), .A2(n6123), .A3(n4675), .ZN(n6700) );
  NAND3_X1 U6436 ( .A1(n6122), .A2(n6136), .A3(P2_REG3_REG_0__SCAN_IN), .ZN(
        n4676) );
  NAND3_X1 U6437 ( .A1(n4679), .A2(n4678), .A3(P2_REG0_REG_0__SCAN_IN), .ZN(
        n4677) );
  NOR2_X4 U6438 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n5568) );
  NAND3_X1 U6439 ( .A1(n10144), .A2(n10153), .A3(n5020), .ZN(n4686) );
  NAND2_X1 U6440 ( .A1(n4687), .A2(n4686), .ZN(n10046) );
  NAND2_X1 U6441 ( .A1(n7089), .A2(n4693), .ZN(n7182) );
  MUX2_X1 U6442 ( .A(P1_REG2_REG_2__SCAN_IN), .B(n6976), .S(n7059), .Z(n4696)
         );
  NAND2_X1 U6443 ( .A1(n4700), .A2(n7280), .ZN(n7414) );
  NAND2_X1 U6444 ( .A1(n7392), .A2(n4703), .ZN(n7467) );
  INV_X2 U6445 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n9635) );
  NAND3_X1 U6446 ( .A1(n4709), .A2(n5897), .A3(n4708), .ZN(n4707) );
  AND2_X2 U6447 ( .A1(n5998), .A2(n5836), .ZN(n5695) );
  NAND2_X1 U6448 ( .A1(n5359), .A2(n4410), .ZN(n4720) );
  NAND3_X1 U6449 ( .A1(n5347), .A2(n4721), .A3(n5201), .ZN(n4719) );
  INV_X1 U6450 ( .A(n5236), .ZN(n4729) );
  OAI21_X1 U6451 ( .B1(n5236), .B2(n4734), .A(n4732), .ZN(n5699) );
  OAI21_X1 U6452 ( .B1(n4729), .B2(n4731), .A(n4730), .ZN(n5239) );
  NAND2_X1 U6453 ( .A1(n5236), .A2(n5235), .ZN(n5281) );
  MUX2_X1 U6454 ( .A(n7672), .B(P2_REG2_REG_1__SCAN_IN), .S(n7272), .Z(n7269)
         );
  XNOR2_X1 U6455 ( .A(n4735), .B(n6129), .ZN(n7272) );
  NAND2_X1 U6456 ( .A1(n7148), .A2(n4737), .ZN(n7124) );
  INV_X1 U6457 ( .A(n7153), .ZN(n4738) );
  NAND2_X1 U6458 ( .A1(n8848), .A2(n8541), .ZN(n8866) );
  INV_X1 U6459 ( .A(n4743), .ZN(n8864) );
  INV_X1 U6460 ( .A(n8865), .ZN(n4744) );
  NAND3_X1 U6461 ( .A1(n4709), .A2(n5813), .A3(n5814), .ZN(n4762) );
  OR2_X1 U6462 ( .A1(n5764), .A2(n4772), .ZN(n4771) );
  NAND3_X1 U6463 ( .A1(n4771), .A2(n4769), .A3(n4768), .ZN(n5771) );
  NAND2_X1 U6464 ( .A1(n4783), .A2(n5970), .ZN(n5977) );
  NAND2_X1 U6465 ( .A1(n4783), .A2(n8033), .ZN(n8034) );
  NAND3_X1 U6466 ( .A1(n5909), .A2(n5739), .A3(n4474), .ZN(n5642) );
  XNOR2_X2 U6467 ( .A(n5737), .B(n7802), .ZN(n4784) );
  NAND2_X2 U6468 ( .A1(n9716), .A2(n5992), .ZN(n9715) );
  NAND2_X1 U6469 ( .A1(n4785), .A2(n5862), .ZN(n5907) );
  NAND2_X1 U6470 ( .A1(n4787), .A2(n4786), .ZN(n6877) );
  INV_X1 U6471 ( .A(n6875), .ZN(n4786) );
  INV_X1 U6472 ( .A(n9670), .ZN(n4788) );
  NAND2_X1 U6473 ( .A1(n4789), .A2(n4478), .ZN(n6616) );
  NAND2_X1 U6474 ( .A1(n5867), .A2(n5855), .ZN(n4810) );
  NAND3_X1 U6475 ( .A1(n6574), .A2(n6576), .A3(n4394), .ZN(n4813) );
  AND2_X1 U6476 ( .A1(n7712), .A2(n6636), .ZN(n6518) );
  NOR2_X2 U6477 ( .A1(P1_IR_REG_18__SCAN_IN), .A2(P1_IR_REG_16__SCAN_IN), .ZN(
        n5257) );
  NOR2_X2 U6478 ( .A1(P1_IR_REG_17__SCAN_IN), .A2(P1_IR_REG_20__SCAN_IN), .ZN(
        n5255) );
  NOR2_X2 U6479 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P1_IR_REG_15__SCAN_IN), .ZN(
        n5256) );
  NAND2_X1 U6480 ( .A1(n8842), .A2(n7680), .ZN(n7712) );
  XNOR2_X1 U6481 ( .A(n5648), .B(n5649), .ZN(n6998) );
  XNOR2_X1 U6482 ( .A(n4873), .B(n5618), .ZN(n5622) );
  NOR2_X1 U6483 ( .A1(n10330), .A2(n10331), .ZN(n10329) );
  NAND2_X1 U6484 ( .A1(n5986), .A2(n5985), .ZN(n10135) );
  INV_X1 U6485 ( .A(n10131), .ZN(n5986) );
  NAND2_X1 U6486 ( .A1(n9149), .A2(n4830), .ZN(n4829) );
  NAND3_X1 U6487 ( .A1(n4430), .A2(n4402), .A3(n7671), .ZN(n6907) );
  NOR2_X1 U6488 ( .A1(n8110), .A2(n4843), .ZN(n4842) );
  NAND3_X1 U6489 ( .A1(n4837), .A2(n4838), .A3(n4845), .ZN(n8293) );
  AOI21_X2 U6490 ( .B1(n4842), .B2(n4839), .A(n4456), .ZN(n4838) );
  NAND2_X1 U6491 ( .A1(n6921), .A2(n6918), .ZN(n4848) );
  NAND2_X1 U6492 ( .A1(n7550), .A2(n4463), .ZN(n4846) );
  NAND2_X1 U6493 ( .A1(n4847), .A2(n4846), .ZN(n6922) );
  NAND2_X1 U6494 ( .A1(n7550), .A2(n6915), .ZN(n7710) );
  INV_X1 U6495 ( .A(n6915), .ZN(n4851) );
  AOI21_X1 U6496 ( .B1(n4409), .B2(n8295), .A(n4483), .ZN(n9185) );
  NAND3_X1 U6497 ( .A1(n8299), .A2(n8912), .A3(n9197), .ZN(n4861) );
  NAND2_X1 U6498 ( .A1(n9215), .A2(n8914), .ZN(n4862) );
  NAND2_X1 U6499 ( .A1(n9000), .A2(n4469), .ZN(n4864) );
  OAI211_X1 U6500 ( .C1(n9000), .C2(n4867), .A(n4865), .B(n4864), .ZN(n9265)
         );
  OAI21_X1 U6501 ( .B1(n9265), .B2(n4870), .A(n4868), .ZN(P2_U3515) );
  OAI21_X1 U6502 ( .B1(n9265), .B2(n9350), .A(n4425), .ZN(n9366) );
  NAND2_X1 U6503 ( .A1(n5674), .A2(n5131), .ZN(n4872) );
  NAND2_X1 U6504 ( .A1(n4873), .A2(n5108), .ZN(n5111) );
  NAND2_X1 U6505 ( .A1(n4880), .A2(n4879), .ZN(n4878) );
  NAND2_X1 U6506 ( .A1(n6616), .A2(n6615), .ZN(n4880) );
  NAND2_X4 U6507 ( .A1(n4883), .A2(n4881), .ZN(n5128) );
  NAND3_X1 U6508 ( .A1(n4889), .A2(n4892), .A3(n5454), .ZN(n4888) );
  NAND2_X1 U6509 ( .A1(n5499), .A2(n5144), .ZN(n5151) );
  INV_X1 U6510 ( .A(n7965), .ZN(n4899) );
  NAND3_X1 U6511 ( .A1(n4899), .A2(n4398), .A3(n8208), .ZN(n8146) );
  AND2_X2 U6512 ( .A1(n9732), .A2(n4411), .ZN(n9666) );
  AND2_X2 U6513 ( .A1(n8221), .A2(n4907), .ZN(n10127) );
  NAND2_X1 U6514 ( .A1(n5726), .A2(n5725), .ZN(n5831) );
  NAND2_X1 U6515 ( .A1(n5726), .A2(n4912), .ZN(n5731) );
  NAND2_X1 U6516 ( .A1(n5415), .A2(n4916), .ZN(n4914) );
  NAND3_X1 U6517 ( .A1(n4922), .A2(n4921), .A3(n4919), .ZN(n5441) );
  NAND2_X1 U6518 ( .A1(n9457), .A2(n9458), .ZN(n4931) );
  NAND2_X1 U6519 ( .A1(n9457), .A2(n4924), .ZN(n4923) );
  NAND2_X1 U6520 ( .A1(n4931), .A2(n4929), .ZN(n9539) );
  AND2_X1 U6521 ( .A1(n4931), .A2(n4930), .ZN(n9541) );
  INV_X1 U6522 ( .A(n7875), .ZN(n4935) );
  NAND2_X1 U6523 ( .A1(n4933), .A2(n7875), .ZN(n4932) );
  NAND2_X1 U6524 ( .A1(n4934), .A2(n7875), .ZN(n7876) );
  NAND2_X1 U6525 ( .A1(n9551), .A2(n4471), .ZN(n4937) );
  NAND3_X1 U6526 ( .A1(n9548), .A2(n9552), .A3(n4940), .ZN(n4939) );
  NAND2_X1 U6527 ( .A1(n4944), .A2(n4482), .ZN(n8573) );
  NOR2_X1 U6528 ( .A1(n8519), .A2(n4962), .ZN(n4961) );
  OAI21_X1 U6529 ( .B1(n8318), .B2(n4967), .A(n4963), .ZN(n8449) );
  NAND2_X1 U6530 ( .A1(n7569), .A2(n6941), .ZN(n7582) );
  OAI22_X1 U6531 ( .A1(n6157), .A2(n5113), .B1(n7103), .B2(n7120), .ZN(n4981)
         );
  NAND2_X1 U6532 ( .A1(n9007), .A2(n4986), .ZN(n8946) );
  NAND2_X1 U6533 ( .A1(n9127), .A2(n4987), .ZN(n9068) );
  NAND2_X1 U6534 ( .A1(n4429), .A2(n4992), .ZN(n7812) );
  INV_X2 U6535 ( .A(n6812), .ZN(n7520) );
  INV_X1 U6536 ( .A(n6863), .ZN(n4995) );
  INV_X2 U6537 ( .A(n6696), .ZN(n6657) );
  NAND2_X1 U6538 ( .A1(n4996), .A2(n6812), .ZN(n6709) );
  NAND2_X1 U6539 ( .A1(n4997), .A2(n6666), .ZN(n6661) );
  AND2_X1 U6540 ( .A1(n6014), .A2(n6011), .ZN(n4998) );
  NAND2_X1 U6541 ( .A1(n7606), .A2(n6729), .ZN(n7660) );
  NAND2_X2 U6542 ( .A1(n8655), .A2(n6775), .ZN(n8820) );
  NAND2_X1 U6543 ( .A1(n6768), .A2(n4475), .ZN(n8655) );
  NAND2_X1 U6544 ( .A1(n7834), .A2(n6017), .ZN(n5003) );
  NAND2_X1 U6545 ( .A1(n5008), .A2(n4480), .ZN(n6046) );
  NAND2_X1 U6546 ( .A1(n8423), .A2(n5009), .ZN(n5008) );
  NAND2_X1 U6547 ( .A1(n5015), .A2(n5016), .ZN(n8186) );
  NAND2_X1 U6548 ( .A1(n6755), .A2(n4427), .ZN(n5015) );
  OR2_X2 U6549 ( .A1(n9678), .A2(n6049), .ZN(n5026) );
  NAND3_X1 U6550 ( .A1(n4541), .A2(n6171), .A3(n6098), .ZN(n6317) );
  NAND2_X1 U6551 ( .A1(n8717), .A2(n4466), .ZN(n5032) );
  NAND2_X1 U6552 ( .A1(n5032), .A2(n4481), .ZN(n8805) );
  NAND2_X1 U6553 ( .A1(n8678), .A2(n4467), .ZN(n5038) );
  NAND2_X1 U6554 ( .A1(n5038), .A2(n5039), .ZN(n8701) );
  NAND2_X1 U6555 ( .A1(n5044), .A2(n4436), .ZN(n6026) );
  NAND2_X1 U6556 ( .A1(n7906), .A2(n4403), .ZN(n5044) );
  INV_X1 U6557 ( .A(n6019), .ZN(n5049) );
  NAND2_X1 U6558 ( .A1(n7906), .A2(n7905), .ZN(n7904) );
  INV_X1 U6559 ( .A(n8708), .ZN(n5060) );
  NAND2_X1 U6560 ( .A1(n8844), .A2(n6812), .ZN(n6702) );
  XNOR2_X2 U6561 ( .A(n5065), .B(P2_IR_REG_30__SCAN_IN), .ZN(n6122) );
  AND2_X2 U6562 ( .A1(n9385), .A2(n5066), .ZN(n6136) );
  NAND2_X1 U6563 ( .A1(n8090), .A2(n5069), .ZN(n5068) );
  OAI21_X1 U6564 ( .B1(n6256), .B2(n5071), .A(n6639), .ZN(n5070) );
  INV_X1 U6565 ( .A(n5074), .ZN(n5073) );
  NAND2_X1 U6566 ( .A1(n8964), .A2(n6605), .ZN(n8905) );
  NAND2_X1 U6567 ( .A1(n6477), .A2(n4499), .ZN(n6481) );
  NAND2_X1 U6568 ( .A1(n7818), .A2(n7817), .ZN(n7816) );
  NAND2_X2 U6569 ( .A1(n9043), .A2(n6585), .ZN(n9046) );
  NAND3_X2 U6570 ( .A1(n5080), .A2(n6171), .A3(n6097), .ZN(n6673) );
  AND4_X2 U6571 ( .A1(n5092), .A2(n6490), .A3(n5081), .A4(n5083), .ZN(n5080)
         );
  NAND3_X1 U6572 ( .A1(n5082), .A2(n6171), .A3(n4541), .ZN(n6670) );
  OR2_X1 U6573 ( .A1(n7582), .A2(n7546), .ZN(n7556) );
  NAND2_X1 U6574 ( .A1(n9266), .A2(n10583), .ZN(n9272) );
  XNOR2_X1 U6575 ( .A(n5115), .B(SI_2_), .ZN(n5566) );
  OAI21_X1 U6576 ( .B1(n5128), .B2(n5123), .A(n5122), .ZN(n5124) );
  NAND2_X1 U6577 ( .A1(n5128), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n5122) );
  OAI21_X1 U6578 ( .B1(n5128), .B2(n5118), .A(n5117), .ZN(n5125) );
  NAND2_X1 U6579 ( .A1(n5128), .A2(P2_DATAO_REG_5__SCAN_IN), .ZN(n5117) );
  OAI21_X1 U6580 ( .B1(n5128), .B2(n5113), .A(n5112), .ZN(n5115) );
  NAND2_X1 U6581 ( .A1(n5128), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n5112) );
  OR2_X2 U6582 ( .A1(n9638), .A2(n10158), .ZN(n10166) );
  OR2_X1 U6583 ( .A1(n9253), .A2(n9252), .ZN(n9254) );
  AND2_X1 U6584 ( .A1(n10314), .A2(n10306), .ZN(n10395) );
  NAND2_X2 U6585 ( .A1(n8492), .A2(n8491), .ZN(n9500) );
  INV_X1 U6586 ( .A(n9637), .ZN(n9647) );
  XNOR2_X1 U6587 ( .A(n6709), .B(n6707), .ZN(n8794) );
  NOR2_X1 U6588 ( .A1(n8644), .A2(n8643), .ZN(n8647) );
  NAND2_X1 U6589 ( .A1(n8840), .A2(n6812), .ZN(n6727) );
  NAND2_X2 U6590 ( .A1(n8665), .A2(n6811), .ZN(n8743) );
  OR2_X1 U6591 ( .A1(n6131), .A2(n7029), .ZN(n6132) );
  NAND2_X2 U6592 ( .A1(n6186), .A2(n6185), .ZN(n6717) );
  AOI211_X2 U6593 ( .C1(n6725), .C2(n7603), .A(n7602), .B(n7605), .ZN(n6726)
         );
  AND2_X1 U6594 ( .A1(n6724), .A2(n6723), .ZN(n7602) );
  CLKBUF_X1 U6595 ( .A(n8805), .Z(n8807) );
  INV_X1 U6596 ( .A(n7907), .ZN(n7966) );
  OR2_X1 U6597 ( .A1(n6966), .A2(n5571), .ZN(n5572) );
  NAND2_X1 U6598 ( .A1(n7563), .A2(n6910), .ZN(n7564) );
  NAND2_X1 U6599 ( .A1(n6908), .A2(n6907), .ZN(n7563) );
  NAND2_X1 U6600 ( .A1(n8899), .A2(n8898), .ZN(n8948) );
  AND2_X1 U6601 ( .A1(n6700), .A2(n10569), .ZN(n6909) );
  NAND3_X2 U6602 ( .A1(n5631), .A2(n5630), .A3(n5629), .ZN(n7802) );
  CLKBUF_X1 U6603 ( .A(n8335), .Z(n8336) );
  AOI211_X1 U6604 ( .C1(n8800), .C2(n7584), .A(n10590), .B(n7583), .ZN(n7692)
         );
  XNOR2_X1 U6605 ( .A(n6705), .B(n8800), .ZN(n6707) );
  NAND4_X2 U6606 ( .A1(n5616), .A2(n5613), .A3(n5614), .A4(n5615), .ZN(n5737)
         );
  OAI21_X1 U6607 ( .B1(n6673), .B2(n6109), .A(n6108), .ZN(n6111) );
  AOI21_X1 U6608 ( .B1(n8915), .B2(n9206), .A(n9183), .ZN(n9164) );
  NOR2_X1 U6609 ( .A1(n6870), .A2(n6869), .ZN(n5084) );
  INV_X1 U6610 ( .A(n8821), .ZN(n6894) );
  NOR2_X1 U6611 ( .A1(n8274), .A2(n8273), .ZN(n5085) );
  AND2_X1 U6612 ( .A1(n9652), .A2(n10489), .ZN(n5086) );
  INV_X1 U6613 ( .A(n8619), .ZN(n6888) );
  INV_X1 U6614 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n5113) );
  NOR2_X1 U6615 ( .A1(n6691), .A2(n10236), .ZN(n5087) );
  OR2_X1 U6616 ( .A1(n10504), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n5088) );
  AND2_X1 U6617 ( .A1(n9251), .A2(n9250), .ZN(n5090) );
  AND2_X1 U6618 ( .A1(n5097), .A2(n5500), .ZN(n5091) );
  AND2_X1 U6619 ( .A1(n6490), .A2(n6489), .ZN(n5093) );
  OR2_X1 U6620 ( .A1(n10492), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n5094) );
  OR2_X1 U6621 ( .A1(P1_REG0_REG_31__SCAN_IN), .A2(n10492), .ZN(n5095) );
  INV_X1 U6622 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n5632) );
  AND2_X1 U6623 ( .A1(n5592), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(n5096) );
  OR2_X1 U6624 ( .A1(P2_IR_REG_29__SCAN_IN), .A2(P2_IR_REG_31__SCAN_IN), .ZN(
        n5098) );
  AND2_X1 U6625 ( .A1(n5166), .A2(n5165), .ZN(n5099) );
  AND2_X1 U6626 ( .A1(n5180), .A2(n5179), .ZN(n5100) );
  INV_X1 U6627 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n6260) );
  INV_X1 U6628 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n5130) );
  INV_X1 U6629 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n5123) );
  INV_X1 U6630 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n5120) );
  AND2_X2 U6631 ( .A1(n6690), .A2(n6689), .ZN(n10504) );
  INV_X1 U6632 ( .A(n10504), .ZN(n10168) );
  NAND2_X2 U6633 ( .A1(n7839), .A2(n10145), .ZN(n10148) );
  INV_X1 U6634 ( .A(n5611), .ZN(n5585) );
  OR2_X1 U6635 ( .A1(n8840), .A2(n7783), .ZN(n5101) );
  AND3_X1 U6636 ( .A1(n9271), .A2(n9270), .A3(n9269), .ZN(n5102) );
  INV_X1 U6637 ( .A(n5279), .ZN(n5937) );
  NAND2_X1 U6638 ( .A1(n10248), .A2(n9641), .ZN(n5279) );
  INV_X1 U6639 ( .A(n8633), .ZN(n9020) );
  AND2_X1 U6640 ( .A1(n5125), .A2(SI_5_), .ZN(n5104) );
  AND2_X1 U6641 ( .A1(n6384), .A2(n6383), .ZN(n9076) );
  INV_X1 U6642 ( .A(n8299), .ZN(n8294) );
  INV_X1 U6643 ( .A(n8163), .ZN(n6056) );
  INV_X1 U6644 ( .A(n6924), .ZN(n6229) );
  NAND2_X1 U6645 ( .A1(n6812), .A2(n6928), .ZN(n6497) );
  INV_X1 U6646 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n6489) );
  INV_X1 U6647 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n6094) );
  NAND2_X1 U6648 ( .A1(n6618), .A2(n6621), .ZN(n6626) );
  INV_X1 U6649 ( .A(n7659), .ZN(n6734) );
  INV_X1 U6650 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n6193) );
  AND2_X1 U6651 ( .A1(n6037), .A2(n10050), .ZN(n6038) );
  INV_X1 U6652 ( .A(n8069), .ZN(n5969) );
  INV_X1 U6653 ( .A(SI_16_), .ZN(n5176) );
  AND2_X1 U6654 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_REG3_REG_7__SCAN_IN), 
        .ZN(n6200) );
  NOR2_X1 U6655 ( .A1(n7715), .A2(n7520), .ZN(n6715) );
  OR2_X1 U6656 ( .A1(n9426), .A2(n9485), .ZN(n8571) );
  INV_X1 U6657 ( .A(n6953), .ZN(n7423) );
  AND2_X1 U6658 ( .A1(n5317), .A2(n5284), .ZN(n5305) );
  INV_X1 U6659 ( .A(SI_25_), .ZN(n9887) );
  INV_X1 U6660 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n5722) );
  NOR2_X1 U6661 ( .A1(n5183), .A2(n5182), .ZN(n5188) );
  INV_X1 U6662 ( .A(SI_15_), .ZN(n5170) );
  NAND2_X1 U6663 ( .A1(n7001), .A2(P2_DATAO_REG_6__SCAN_IN), .ZN(n5129) );
  NAND2_X1 U6664 ( .A1(n5128), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n5119) );
  INV_X1 U6665 ( .A(n8657), .ZN(n6774) );
  INV_X1 U6666 ( .A(n8720), .ZN(n6786) );
  NAND2_X1 U6667 ( .A1(n6716), .A2(n7599), .ZN(n7601) );
  INV_X1 U6668 ( .A(n9245), .ZN(n8898) );
  INV_X1 U6669 ( .A(n7817), .ZN(n6921) );
  INV_X1 U6670 ( .A(n6909), .ZN(n6910) );
  INV_X1 U6671 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n9791) );
  INV_X1 U6672 ( .A(n7738), .ZN(n7734) );
  INV_X1 U6673 ( .A(n9646), .ZN(n9636) );
  AND2_X1 U6674 ( .A1(n5320), .A2(n5319), .ZN(n9706) );
  INV_X1 U6675 ( .A(n8430), .ZN(n8424) );
  INV_X1 U6676 ( .A(n10130), .ZN(n5985) );
  INV_X1 U6677 ( .A(n7842), .ZN(n6016) );
  OR2_X1 U6678 ( .A1(n6949), .A2(n6950), .ZN(n7359) );
  OR2_X1 U6679 ( .A1(n5699), .A2(n5696), .ZN(n5708) );
  AND3_X1 U6680 ( .A1(n5724), .A2(n5723), .A3(n5722), .ZN(n5725) );
  NAND2_X1 U6681 ( .A1(n5163), .A2(n5162), .ZN(n5166) );
  AND2_X1 U6682 ( .A1(n6828), .A2(n6826), .ZN(n8643) );
  NAND2_X1 U6683 ( .A1(n7706), .A2(n6698), .ZN(n6863) );
  BUF_X4 U6684 ( .A(n6175), .Z(n6468) );
  INV_X1 U6685 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n9890) );
  OR2_X1 U6686 ( .A1(n8901), .A2(n9245), .ZN(n8634) );
  NAND2_X1 U6687 ( .A1(n8960), .A2(n6629), .ZN(n9003) );
  NAND2_X1 U6688 ( .A1(n9086), .A2(n9076), .ZN(n8922) );
  AND2_X1 U6689 ( .A1(n6624), .A2(n6697), .ZN(n7102) );
  OR2_X1 U6690 ( .A1(n7812), .A2(n6944), .ZN(n8052) );
  OR2_X1 U6691 ( .A1(n6938), .A2(n7534), .ZN(n6940) );
  OR2_X1 U6692 ( .A1(n6940), .A2(n6625), .ZN(n7718) );
  INV_X1 U6693 ( .A(n9220), .ZN(n9203) );
  NOR2_X1 U6694 ( .A1(n10590), .A2(n7706), .ZN(n7532) );
  OR2_X1 U6695 ( .A1(n8576), .A2(n8575), .ZN(n8577) );
  OR2_X1 U6696 ( .A1(n7357), .A2(n7356), .ZN(n7509) );
  INV_X1 U6697 ( .A(n5904), .ZN(n5956) );
  INV_X1 U6698 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n7619) );
  INV_X1 U6699 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n9766) );
  INV_X1 U6700 ( .A(n10363), .ZN(n10390) );
  INV_X1 U6701 ( .A(n9697), .ZN(n5994) );
  NAND2_X1 U6702 ( .A1(n7512), .A2(n7511), .ZN(n7839) );
  INV_X1 U6703 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n10167) );
  AND2_X1 U6704 ( .A1(n9660), .A2(n6062), .ZN(n6063) );
  AND2_X1 U6705 ( .A1(n9717), .A2(n5923), .ZN(n10021) );
  AND2_X1 U6706 ( .A1(n7900), .A2(n7899), .ZN(n7962) );
  AND2_X1 U6707 ( .A1(n5216), .A2(n5215), .ZN(n5347) );
  AND2_X1 U6708 ( .A1(n5199), .A2(n5198), .ZN(n5372) );
  INV_X1 U6709 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n5620) );
  NAND2_X1 U6710 ( .A1(n8816), .A2(n9222), .ZN(n8785) );
  NAND2_X1 U6711 ( .A1(n6850), .A2(n9188), .ZN(n8825) );
  OR2_X1 U6712 ( .A1(n8945), .A2(n6467), .ZN(n6475) );
  AND2_X1 U6713 ( .A1(n6394), .A2(n6393), .ZN(n9092) );
  AND2_X1 U6714 ( .A1(n7108), .A2(n7107), .ZN(n10505) );
  AND2_X1 U6715 ( .A1(n7123), .A2(n7105), .ZN(n8870) );
  AND2_X1 U6716 ( .A1(n6631), .A2(n6630), .ZN(n9136) );
  INV_X1 U6717 ( .A(n9188), .ZN(n10517) );
  NAND2_X1 U6718 ( .A1(n6835), .A2(n10563), .ZN(n7561) );
  INV_X1 U6719 ( .A(n10583), .ZN(n9350) );
  NAND2_X1 U6720 ( .A1(n7666), .A2(n10586), .ZN(n10583) );
  INV_X1 U6721 ( .A(n7561), .ZN(n7535) );
  NAND2_X1 U6722 ( .A1(n7099), .A2(n6680), .ZN(n10530) );
  INV_X1 U6723 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n6677) );
  AND2_X1 U6724 ( .A1(n6245), .A2(n6257), .ZN(n7335) );
  XNOR2_X1 U6725 ( .A(n5902), .B(P1_IR_REG_23__SCAN_IN), .ZN(n6902) );
  OR2_X1 U6726 ( .A1(n9402), .A2(n8607), .ZN(n8598) );
  INV_X1 U6727 ( .A(n9560), .ZN(n9542) );
  NOR2_X1 U6728 ( .A1(n7509), .A2(n7358), .ZN(n7371) );
  AND2_X1 U6729 ( .A1(n9532), .A2(n10240), .ZN(n9518) );
  INV_X1 U6730 ( .A(n10399), .ZN(n10319) );
  AND2_X1 U6731 ( .A1(n4496), .A2(n7366), .ZN(n10383) );
  AND2_X1 U6732 ( .A1(n4496), .A2(n10290), .ZN(n10363) );
  INV_X1 U6733 ( .A(n9659), .ZN(n10422) );
  AND2_X1 U6734 ( .A1(n10148), .A2(n7801), .ZN(n10150) );
  INV_X1 U6735 ( .A(n10236), .ZN(n6884) );
  AND2_X1 U6736 ( .A1(n10278), .A2(n7363), .ZN(n6689) );
  AND2_X1 U6737 ( .A1(n7424), .A2(n10473), .ZN(n10243) );
  AND2_X1 U6738 ( .A1(n7497), .A2(P1_STATE_REG_SCAN_IN), .ZN(n5952) );
  AND2_X1 U6739 ( .A1(n5488), .A2(n5487), .ZN(n7622) );
  INV_X1 U6740 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n9917) );
  NOR2_X1 U6741 ( .A1(n10637), .A2(n8380), .ZN(n8381) );
  OAI21_X1 U6742 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(P1_ADDR_REG_17__SCAN_IN), 
        .A(n10611), .ZN(n10640) );
  INV_X1 U6743 ( .A(n8863), .ZN(n10508) );
  INV_X1 U6744 ( .A(n8825), .ZN(n8695) );
  AND3_X1 U6745 ( .A1(n6114), .A2(n6113), .A3(n6112), .ZN(n8908) );
  NAND2_X1 U6746 ( .A1(n6416), .A2(n6415), .ZN(n9049) );
  INV_X1 U6747 ( .A(n10505), .ZN(n10510) );
  OR2_X1 U6748 ( .A1(n10529), .A2(n6943), .ZN(n10523) );
  INV_X1 U6749 ( .A(n9060), .ZN(n10529) );
  OR2_X1 U6750 ( .A1(n10529), .A2(n7667), .ZN(n9231) );
  OR2_X1 U6751 ( .A1(n7562), .A2(n7561), .ZN(n10603) );
  NAND2_X1 U6752 ( .A1(n9272), .A2(n5102), .ZN(n9367) );
  OR3_X1 U6753 ( .A1(n9341), .A2(n9340), .A3(n9339), .ZN(n9380) );
  OR2_X1 U6754 ( .A1(n7562), .A2(n7535), .ZN(n10596) );
  NOR2_X1 U6755 ( .A1(n10531), .A2(n10530), .ZN(n10546) );
  INV_X1 U6756 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n9836) );
  INV_X1 U6757 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n9948) );
  INV_X1 U6758 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n7077) );
  NAND2_X1 U6759 ( .A1(n7371), .A2(n7370), .ZN(n9520) );
  INV_X1 U6760 ( .A(n9518), .ZN(n9556) );
  INV_X1 U6761 ( .A(n9699), .ZN(n9568) );
  INV_X1 U6762 ( .A(n10133), .ZN(n9574) );
  INV_X1 U6763 ( .A(n10395), .ZN(n7629) );
  OR2_X1 U6764 ( .A1(P1_U3083), .A2(n6965), .ZN(n10399) );
  INV_X1 U6765 ( .A(n10150), .ZN(n10400) );
  AND2_X1 U6766 ( .A1(n10045), .A2(n10044), .ZN(n10208) );
  NAND2_X1 U6767 ( .A1(n10504), .A2(n10240), .ZN(n10236) );
  INV_X1 U6768 ( .A(n8454), .ZN(n9557) );
  OR2_X1 U6769 ( .A1(n7510), .A2(n6688), .ZN(n10490) );
  INV_X2 U6770 ( .A(n10490), .ZN(n10492) );
  AND2_X1 U6771 ( .A1(n10429), .A2(n10428), .ZN(n10434) );
  INV_X1 U6772 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n8407) );
  INV_X1 U6773 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n9886) );
  INV_X1 U6774 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n9936) );
  OAI21_X1 U6775 ( .B1(n7292), .B2(n8376), .A(n8375), .ZN(n10658) );
  NOR2_X1 U6776 ( .A1(n10634), .A2(n10633), .ZN(n10632) );
  OAI21_X1 U6777 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(P1_ADDR_REG_13__SCAN_IN), 
        .A(n10623), .ZN(n10621) );
  INV_X2 U6778 ( .A(n8832), .ZN(P2_U3966) );
  AND2_X1 U6779 ( .A1(SI_0_), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n5106) );
  NAND2_X1 U6780 ( .A1(n5128), .A2(n5106), .ZN(n5582) );
  AND2_X1 U6781 ( .A1(SI_0_), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n5107) );
  NAND2_X1 U6782 ( .A1(n7002), .A2(n5107), .ZN(n6127) );
  NAND2_X1 U6783 ( .A1(n5128), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n5619) );
  INV_X1 U6784 ( .A(SI_1_), .ZN(n5618) );
  OAI211_X1 U6785 ( .C1(n5128), .C2(n5620), .A(n5619), .B(n5618), .ZN(n5108)
         );
  INV_X1 U6786 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n7028) );
  NAND2_X1 U6787 ( .A1(n5128), .A2(n7028), .ZN(n5109) );
  OAI211_X1 U6788 ( .C1(n5128), .C2(P1_DATAO_REG_1__SCAN_IN), .A(n5109), .B(
        SI_1_), .ZN(n5110) );
  INV_X1 U6789 ( .A(n5566), .ZN(n5114) );
  NAND2_X1 U6790 ( .A1(n5115), .A2(SI_2_), .ZN(n5116) );
  XNOR2_X1 U6791 ( .A(n5125), .B(SI_5_), .ZN(n5648) );
  OAI21_X1 U6792 ( .B1(n5128), .B2(n5120), .A(n5119), .ZN(n5608) );
  NOR2_X1 U6793 ( .A1(n5608), .A2(SI_4_), .ZN(n5121) );
  XNOR2_X1 U6794 ( .A(n5124), .B(SI_3_), .ZN(n5590) );
  INV_X1 U6795 ( .A(n5590), .ZN(n5604) );
  NAND2_X1 U6796 ( .A1(n5608), .A2(SI_4_), .ZN(n5646) );
  NAND2_X1 U6797 ( .A1(n5124), .A2(SI_3_), .ZN(n5606) );
  BUF_X8 U6798 ( .A(n5128), .Z(n7001) );
  XNOR2_X1 U6799 ( .A(n5132), .B(SI_6_), .ZN(n5673) );
  INV_X1 U6800 ( .A(n5673), .ZN(n5131) );
  NAND2_X1 U6801 ( .A1(n5132), .A2(SI_6_), .ZN(n5133) );
  MUX2_X1 U6802 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .S(n7001), .Z(n5135) );
  XNOR2_X1 U6803 ( .A(n5135), .B(SI_7_), .ZN(n5638) );
  INV_X1 U6804 ( .A(n5638), .ZN(n5134) );
  NAND2_X1 U6805 ( .A1(n5135), .A2(SI_7_), .ZN(n5136) );
  MUX2_X1 U6806 ( .A(n9741), .B(n7014), .S(n7001), .Z(n5139) );
  INV_X1 U6807 ( .A(SI_8_), .ZN(n5138) );
  NAND2_X1 U6808 ( .A1(n5139), .A2(n5138), .ZN(n5498) );
  INV_X1 U6809 ( .A(n5139), .ZN(n5140) );
  NAND2_X1 U6810 ( .A1(n5140), .A2(SI_8_), .ZN(n5141) );
  NAND2_X1 U6811 ( .A1(n5498), .A2(n5141), .ZN(n5547) );
  INV_X1 U6812 ( .A(n5547), .ZN(n5142) );
  MUX2_X1 U6813 ( .A(n7025), .B(n7026), .S(n7001), .Z(n5149) );
  INV_X1 U6814 ( .A(SI_9_), .ZN(n5143) );
  NAND2_X1 U6815 ( .A1(n5149), .A2(n5143), .ZN(n5501) );
  MUX2_X1 U6816 ( .A(n7031), .B(n9936), .S(n7001), .Z(n5146) );
  NAND2_X1 U6817 ( .A1(n5146), .A2(n5145), .ZN(n5152) );
  INV_X1 U6818 ( .A(n5146), .ZN(n5147) );
  NAND2_X1 U6819 ( .A1(n5147), .A2(SI_10_), .ZN(n5148) );
  INV_X1 U6820 ( .A(n5149), .ZN(n5150) );
  NAND2_X1 U6821 ( .A1(n5150), .A2(SI_9_), .ZN(n5500) );
  NAND2_X1 U6822 ( .A1(n5151), .A2(n5091), .ZN(n5153) );
  MUX2_X1 U6823 ( .A(n7034), .B(n7035), .S(n7001), .Z(n5154) );
  XNOR2_X1 U6824 ( .A(n5154), .B(SI_11_), .ZN(n5516) );
  INV_X1 U6825 ( .A(n5154), .ZN(n5155) );
  NAND2_X1 U6826 ( .A1(n5155), .A2(SI_11_), .ZN(n5156) );
  MUX2_X1 U6827 ( .A(n7077), .B(n7079), .S(n7001), .Z(n5158) );
  INV_X1 U6828 ( .A(n5158), .ZN(n5159) );
  NAND2_X1 U6829 ( .A1(n5159), .A2(SI_12_), .ZN(n5160) );
  NAND2_X1 U6830 ( .A1(n5161), .A2(n5160), .ZN(n5483) );
  MUX2_X1 U6831 ( .A(n9873), .B(n7274), .S(n7001), .Z(n5163) );
  INV_X1 U6832 ( .A(n5163), .ZN(n5164) );
  NAND2_X1 U6833 ( .A1(n5164), .A2(SI_13_), .ZN(n5165) );
  MUX2_X1 U6834 ( .A(n7307), .B(n9886), .S(n7001), .Z(n5167) );
  INV_X1 U6835 ( .A(n5167), .ZN(n5168) );
  NAND2_X1 U6836 ( .A1(n5168), .A2(SI_14_), .ZN(n5169) );
  MUX2_X1 U6837 ( .A(n9860), .B(n7456), .S(n7001), .Z(n5171) );
  INV_X1 U6838 ( .A(n5171), .ZN(n5172) );
  NAND2_X1 U6839 ( .A1(n5172), .A2(SI_15_), .ZN(n5173) );
  MUX2_X1 U6840 ( .A(n5175), .B(n7507), .S(n7001), .Z(n5177) );
  INV_X1 U6841 ( .A(n5177), .ZN(n5178) );
  NAND2_X1 U6842 ( .A1(n5178), .A2(SI_16_), .ZN(n5179) );
  MUX2_X1 U6843 ( .A(n7632), .B(n7653), .S(n7001), .Z(n5184) );
  XNOR2_X1 U6844 ( .A(n5184), .B(SI_17_), .ZN(n5413) );
  INV_X1 U6845 ( .A(n5413), .ZN(n5382) );
  MUX2_X1 U6846 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .S(n7001), .Z(n5181) );
  NAND2_X1 U6847 ( .A1(n5181), .A2(SI_18_), .ZN(n5186) );
  INV_X1 U6848 ( .A(n5186), .ZN(n5183) );
  XNOR2_X1 U6849 ( .A(n5181), .B(SI_18_), .ZN(n5385) );
  INV_X1 U6850 ( .A(n5184), .ZN(n5185) );
  NAND2_X1 U6851 ( .A1(n5185), .A2(SI_17_), .ZN(n5383) );
  AND2_X1 U6852 ( .A1(n5383), .A2(n5186), .ZN(n5187) );
  MUX2_X1 U6853 ( .A(n7707), .B(n7709), .S(n7001), .Z(n5190) );
  INV_X1 U6854 ( .A(n5190), .ZN(n5191) );
  NAND2_X1 U6855 ( .A1(n5191), .A2(SI_19_), .ZN(n5192) );
  NAND2_X1 U6856 ( .A1(n5195), .A2(n5192), .ZN(n5401) );
  INV_X1 U6857 ( .A(n5401), .ZN(n5193) );
  MUX2_X1 U6858 ( .A(n9948), .B(n7808), .S(n7001), .Z(n5196) );
  INV_X1 U6859 ( .A(n5196), .ZN(n5197) );
  NAND2_X1 U6860 ( .A1(n5197), .A2(SI_20_), .ZN(n5198) );
  NAND2_X1 U6861 ( .A1(n5371), .A2(n5372), .ZN(n5200) );
  MUX2_X1 U6862 ( .A(n8532), .B(n9929), .S(n7001), .Z(n5202) );
  INV_X1 U6863 ( .A(n5360), .ZN(n5201) );
  INV_X1 U6864 ( .A(n5202), .ZN(n5203) );
  NAND2_X1 U6865 ( .A1(n5203), .A2(SI_21_), .ZN(n5204) );
  MUX2_X1 U6866 ( .A(n9862), .B(n7995), .S(n7001), .Z(n5206) );
  INV_X1 U6867 ( .A(SI_22_), .ZN(n5205) );
  NAND2_X1 U6868 ( .A1(n5206), .A2(n5205), .ZN(n5209) );
  INV_X1 U6869 ( .A(n5206), .ZN(n5207) );
  NAND2_X1 U6870 ( .A1(n5207), .A2(SI_22_), .ZN(n5208) );
  NAND2_X1 U6871 ( .A1(n5209), .A2(n5208), .ZN(n5336) );
  INV_X1 U6872 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n5211) );
  INV_X1 U6873 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n5210) );
  MUX2_X1 U6874 ( .A(n5211), .B(n5210), .S(n7001), .Z(n5213) );
  INV_X1 U6875 ( .A(SI_23_), .ZN(n5212) );
  NAND2_X1 U6876 ( .A1(n5213), .A2(n5212), .ZN(n5216) );
  INV_X1 U6877 ( .A(n5213), .ZN(n5214) );
  NAND2_X1 U6878 ( .A1(n5214), .A2(SI_23_), .ZN(n5215) );
  MUX2_X1 U6879 ( .A(n8255), .B(n8332), .S(n7001), .Z(n5217) );
  XNOR2_X1 U6880 ( .A(n5217), .B(SI_24_), .ZN(n5327) );
  INV_X1 U6881 ( .A(n5327), .ZN(n5220) );
  INV_X1 U6882 ( .A(n5217), .ZN(n5218) );
  NAND2_X1 U6883 ( .A1(n5218), .A2(SI_24_), .ZN(n5219) );
  MUX2_X1 U6884 ( .A(n8404), .B(n8407), .S(n7001), .Z(n5221) );
  NAND2_X1 U6885 ( .A1(n5221), .A2(n9887), .ZN(n5224) );
  INV_X1 U6886 ( .A(n5221), .ZN(n5222) );
  NAND2_X1 U6887 ( .A1(n5222), .A2(SI_25_), .ZN(n5223) );
  NAND2_X1 U6888 ( .A1(n5224), .A2(n5223), .ZN(n5313) );
  INV_X1 U6889 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n8418) );
  MUX2_X1 U6890 ( .A(n9836), .B(n8418), .S(n7001), .Z(n5226) );
  INV_X1 U6891 ( .A(SI_26_), .ZN(n5225) );
  NAND2_X1 U6892 ( .A1(n5226), .A2(n5225), .ZN(n5229) );
  INV_X1 U6893 ( .A(n5226), .ZN(n5227) );
  NAND2_X1 U6894 ( .A1(n5227), .A2(SI_26_), .ZN(n5228) );
  INV_X1 U6895 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n9396) );
  INV_X1 U6896 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n5230) );
  MUX2_X1 U6897 ( .A(n9396), .B(n5230), .S(n7001), .Z(n5232) );
  INV_X1 U6898 ( .A(SI_27_), .ZN(n5231) );
  NAND2_X1 U6899 ( .A1(n5232), .A2(n5231), .ZN(n5235) );
  INV_X1 U6900 ( .A(n5232), .ZN(n5233) );
  NAND2_X1 U6901 ( .A1(n5233), .A2(SI_27_), .ZN(n5234) );
  NAND2_X1 U6902 ( .A1(n5293), .A2(n5294), .ZN(n5236) );
  MUX2_X1 U6903 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(P2_DATAO_REG_28__SCAN_IN), 
        .S(n7001), .Z(n5237) );
  INV_X1 U6904 ( .A(SI_28_), .ZN(n9775) );
  XNOR2_X1 U6905 ( .A(n5237), .B(n9775), .ZN(n5280) );
  INV_X1 U6906 ( .A(n5237), .ZN(n5238) );
  INV_X1 U6907 ( .A(SI_29_), .ZN(n5696) );
  MUX2_X1 U6908 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(P2_DATAO_REG_29__SCAN_IN), 
        .S(n7001), .Z(n5697) );
  NAND2_X1 U6909 ( .A1(n5239), .A2(n5697), .ZN(n5707) );
  MUX2_X1 U6910 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(P1_DATAO_REG_30__SCAN_IN), 
        .S(n4545), .Z(n5709) );
  NAND2_X1 U6911 ( .A1(n5709), .A2(SI_30_), .ZN(n5240) );
  NAND3_X1 U6912 ( .A1(n5707), .A2(n5708), .A3(n5240), .ZN(n5244) );
  INV_X1 U6913 ( .A(n5709), .ZN(n5242) );
  INV_X1 U6914 ( .A(SI_30_), .ZN(n5241) );
  NAND2_X1 U6915 ( .A1(n5242), .A2(n5241), .ZN(n5243) );
  NAND2_X1 U6916 ( .A1(n5244), .A2(n5243), .ZN(n5248) );
  INV_X1 U6917 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n5245) );
  INV_X1 U6918 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n6482) );
  MUX2_X1 U6919 ( .A(n5245), .B(n6482), .S(n4545), .Z(n5246) );
  XNOR2_X1 U6920 ( .A(n5246), .B(SI_31_), .ZN(n5247) );
  NOR2_X2 U6921 ( .A1(P1_IR_REG_14__SCAN_IN), .A2(P1_IR_REG_8__SCAN_IN), .ZN(
        n5252) );
  NOR2_X2 U6922 ( .A1(P1_IR_REG_5__SCAN_IN), .A2(P1_IR_REG_4__SCAN_IN), .ZN(
        n5251) );
  INV_X2 U6923 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n5950) );
  NAND4_X1 U6925 ( .A1(n5946), .A2(n5950), .A3(n5259), .A4(n5944), .ZN(n5260)
         );
  NAND2_X1 U6926 ( .A1(n5269), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5262) );
  NAND2_X1 U6927 ( .A1(n5263), .A2(n5268), .ZN(n5617) );
  NAND2_X2 U6928 ( .A1(n5617), .A2(n10306), .ZN(n6966) );
  INV_X1 U6929 ( .A(n5273), .ZN(n10279) );
  NOR2_X1 U6930 ( .A1(n5273), .A2(n5270), .ZN(n5271) );
  XNOR2_X2 U6931 ( .A(n5275), .B(n5274), .ZN(n8629) );
  INV_X2 U6932 ( .A(n5585), .ZN(n5664) );
  NAND2_X1 U6933 ( .A1(n5664), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n5278) );
  AND2_X2 U6934 ( .A1(n8629), .A2(n10285), .ZN(n5612) );
  NAND2_X1 U6935 ( .A1(n5716), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n5277) );
  AND2_X4 U6936 ( .A1(n10285), .A2(n5288), .ZN(n5715) );
  NAND2_X1 U6937 ( .A1(n5715), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n5276) );
  AND3_X1 U6938 ( .A1(n5278), .A2(n5277), .A3(n5276), .ZN(n5720) );
  NAND2_X1 U6939 ( .A1(n10288), .A2(n5591), .ZN(n5283) );
  NAND2_X1 U6940 ( .A1(n5592), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n5282) );
  NAND2_X1 U6941 ( .A1(n5655), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n5668) );
  NAND2_X1 U6942 ( .A1(n5552), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n5555) );
  OR2_X2 U6943 ( .A1(n5555), .A2(n9915), .ZN(n5542) );
  OR2_X2 U6944 ( .A1(n5542), .A2(n5510), .ZN(n5523) );
  NAND2_X1 U6945 ( .A1(n5491), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n5493) );
  OR2_X2 U6946 ( .A1(n5493), .A2(n7619), .ZN(n5478) );
  INV_X1 U6947 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n9505) );
  INV_X1 U6948 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n5363) );
  OR2_X2 U6949 ( .A1(n5375), .A2(n5363), .ZN(n5365) );
  INV_X1 U6950 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n8527) );
  AND2_X1 U6951 ( .A1(P1_REG3_REG_24__SCAN_IN), .A2(P1_REG3_REG_25__SCAN_IN), 
        .ZN(n5284) );
  INV_X1 U6952 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n9405) );
  INV_X1 U6953 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n5285) );
  OAI21_X1 U6954 ( .B1(n5307), .B2(n9405), .A(n5285), .ZN(n5287) );
  NAND2_X1 U6955 ( .A1(P1_REG3_REG_27__SCAN_IN), .A2(P1_REG3_REG_28__SCAN_IN), 
        .ZN(n5286) );
  OR2_X2 U6956 ( .A1(n5307), .A2(n5286), .ZN(n9656) );
  INV_X1 U6957 ( .A(P1_REG2_REG_28__SCAN_IN), .ZN(n9900) );
  INV_X2 U6958 ( .A(n5585), .ZN(n5714) );
  NAND2_X1 U6959 ( .A1(n5714), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n5291) );
  NAND2_X1 U6960 ( .A1(n5716), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n5290) );
  OAI211_X1 U6961 ( .C1(n9900), .C2(n5422), .A(n5291), .B(n5290), .ZN(n5292)
         );
  AOI21_X2 U6962 ( .B1(n8620), .B2(n5705), .A(n5292), .ZN(n9671) );
  OR2_X2 U6963 ( .A1(n8619), .A2(n9671), .ZN(n5999) );
  NAND2_X1 U6964 ( .A1(n8619), .A2(n9671), .ZN(n5837) );
  NAND2_X1 U6965 ( .A1(n8420), .A2(n5591), .ZN(n5296) );
  NAND2_X1 U6966 ( .A1(n5592), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n5295) );
  XNOR2_X1 U6967 ( .A(n5307), .B(P1_REG3_REG_27__SCAN_IN), .ZN(n9667) );
  INV_X1 U6968 ( .A(P1_REG2_REG_27__SCAN_IN), .ZN(n5299) );
  NAND2_X1 U6969 ( .A1(n5714), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n5298) );
  NAND2_X1 U6970 ( .A1(n5716), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n5297) );
  OAI211_X1 U6971 ( .C1(n5299), .C2(n5422), .A(n5298), .B(n5297), .ZN(n5300)
         );
  AOI21_X2 U6972 ( .B1(n9667), .B2(n5705), .A(n5300), .ZN(n9687) );
  OR2_X2 U6973 ( .A1(n10178), .A2(n9687), .ZN(n5998) );
  NAND2_X1 U6974 ( .A1(n10178), .A2(n9687), .ZN(n5836) );
  XNOR2_X1 U6975 ( .A(n5302), .B(n5301), .ZN(n8416) );
  INV_X2 U6976 ( .A(n5574), .ZN(n5675) );
  NAND2_X1 U6977 ( .A1(n8416), .A2(n5675), .ZN(n5304) );
  NAND2_X1 U6978 ( .A1(n5592), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n5303) );
  INV_X1 U6979 ( .A(n5305), .ZN(n5319) );
  INV_X1 U6980 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n9802) );
  NAND2_X1 U6981 ( .A1(n5319), .A2(n9802), .ZN(n5306) );
  NAND2_X1 U6982 ( .A1(n5307), .A2(n5306), .ZN(n9680) );
  INV_X1 U6983 ( .A(P1_REG2_REG_26__SCAN_IN), .ZN(n9679) );
  NAND2_X1 U6984 ( .A1(n5714), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n5309) );
  NAND2_X1 U6985 ( .A1(n5716), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n5308) );
  OAI211_X1 U6986 ( .C1(n9679), .C2(n5422), .A(n5309), .B(n5308), .ZN(n5310)
         );
  INV_X1 U6987 ( .A(n5310), .ZN(n5311) );
  OR2_X1 U6988 ( .A1(n9690), .A2(n9699), .ZN(n5928) );
  AND2_X1 U6989 ( .A1(n9690), .A2(n9699), .ZN(n5834) );
  INV_X1 U6990 ( .A(n5834), .ZN(n5997) );
  NAND2_X1 U6991 ( .A1(n8402), .A2(n5591), .ZN(n5316) );
  NAND2_X1 U6992 ( .A1(n5592), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n5315) );
  INV_X1 U6993 ( .A(n5317), .ZN(n5353) );
  INV_X1 U6994 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n9493) );
  INV_X1 U6995 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n5318) );
  OAI21_X1 U6996 ( .B1(n5353), .B2(n9493), .A(n5318), .ZN(n5320) );
  NAND2_X1 U6997 ( .A1(n9706), .A2(n5705), .ZN(n5326) );
  INV_X1 U6998 ( .A(P1_REG2_REG_25__SCAN_IN), .ZN(n5323) );
  NAND2_X1 U6999 ( .A1(n5714), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n5322) );
  NAND2_X1 U7000 ( .A1(n5716), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n5321) );
  OAI211_X1 U7001 ( .C1(n5323), .C2(n5422), .A(n5322), .B(n5321), .ZN(n5324)
         );
  INV_X1 U7002 ( .A(n5324), .ZN(n5325) );
  OR2_X2 U7003 ( .A1(n10190), .A2(n9722), .ZN(n9682) );
  NAND2_X1 U7004 ( .A1(n10190), .A2(n9722), .ZN(n5890) );
  XNOR2_X1 U7005 ( .A(n5328), .B(n5327), .ZN(n8254) );
  NAND2_X1 U7006 ( .A1(n8254), .A2(n5675), .ZN(n5330) );
  NAND2_X1 U7007 ( .A1(n5592), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n5329) );
  XNOR2_X1 U7008 ( .A(n5353), .B(P1_REG3_REG_24__SCAN_IN), .ZN(n9723) );
  NAND2_X1 U7009 ( .A1(n9723), .A2(n5705), .ZN(n5335) );
  INV_X1 U7010 ( .A(P1_REG2_REG_24__SCAN_IN), .ZN(n9725) );
  NAND2_X1 U7011 ( .A1(n5664), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n5332) );
  NAND2_X1 U7012 ( .A1(n5716), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n5331) );
  OAI211_X1 U7013 ( .C1(n9725), .C2(n5422), .A(n5332), .B(n5331), .ZN(n5333)
         );
  INV_X1 U7014 ( .A(n5333), .ZN(n5334) );
  OR2_X1 U7015 ( .A1(n9729), .A2(n10025), .ZN(n5888) );
  NAND2_X1 U7016 ( .A1(n9729), .A2(n10025), .ZN(n5993) );
  AND2_X2 U7017 ( .A1(n5888), .A2(n5993), .ZN(n9727) );
  NAND2_X1 U7018 ( .A1(n7993), .A2(n5591), .ZN(n5338) );
  NAND2_X1 U7019 ( .A1(n5592), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n5337) );
  INV_X1 U7020 ( .A(n5339), .ZN(n5351) );
  NAND2_X1 U7021 ( .A1(n5365), .A2(n8527), .ZN(n5340) );
  NAND2_X1 U7022 ( .A1(n5351), .A2(n5340), .ZN(n10031) );
  OR2_X1 U7023 ( .A1(n10031), .A2(n5434), .ZN(n5345) );
  INV_X1 U7024 ( .A(P1_REG2_REG_22__SCAN_IN), .ZN(n10030) );
  NAND2_X1 U7025 ( .A1(n5664), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n5342) );
  NAND2_X1 U7026 ( .A1(n5716), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n5341) );
  OAI211_X1 U7027 ( .C1(n10030), .C2(n5422), .A(n5342), .B(n5341), .ZN(n5343)
         );
  INV_X1 U7028 ( .A(n5343), .ZN(n5344) );
  XNOR2_X1 U7029 ( .A(n5348), .B(n5347), .ZN(n8127) );
  NAND2_X1 U7030 ( .A1(n8127), .A2(n5675), .ZN(n5350) );
  NAND2_X1 U7031 ( .A1(n5592), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n5349) );
  INV_X1 U7032 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n9430) );
  NAND2_X1 U7033 ( .A1(n5351), .A2(n9430), .ZN(n5352) );
  NAND2_X1 U7034 ( .A1(n5353), .A2(n5352), .ZN(n10017) );
  INV_X1 U7035 ( .A(P1_REG2_REG_23__SCAN_IN), .ZN(n10016) );
  NAND2_X1 U7036 ( .A1(n5714), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n5355) );
  NAND2_X1 U7037 ( .A1(n5716), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n5354) );
  OAI211_X1 U7038 ( .C1(n10016), .C2(n5422), .A(n5355), .B(n5354), .ZN(n5356)
         );
  INV_X1 U7039 ( .A(n5356), .ZN(n5357) );
  OR2_X2 U7040 ( .A1(n10201), .A2(n9721), .ZN(n9717) );
  NAND2_X1 U7041 ( .A1(n10201), .A2(n9721), .ZN(n5923) );
  NAND2_X1 U7042 ( .A1(n7929), .A2(n5591), .ZN(n5362) );
  NAND2_X1 U7043 ( .A1(n5592), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n5361) );
  NAND2_X1 U7044 ( .A1(n5375), .A2(n5363), .ZN(n5364) );
  AND2_X1 U7045 ( .A1(n5365), .A2(n5364), .ZN(n10052) );
  NAND2_X1 U7046 ( .A1(n10052), .A2(n5705), .ZN(n5370) );
  INV_X1 U7047 ( .A(P1_REG2_REG_21__SCAN_IN), .ZN(n10053) );
  NAND2_X1 U7048 ( .A1(n5714), .A2(P1_REG1_REG_21__SCAN_IN), .ZN(n5367) );
  NAND2_X1 U7049 ( .A1(n5716), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n5366) );
  OAI211_X1 U7050 ( .C1(n5422), .C2(n10053), .A(n5367), .B(n5366), .ZN(n5368)
         );
  INV_X1 U7051 ( .A(n5368), .ZN(n5369) );
  NAND2_X1 U7052 ( .A1(n10061), .A2(n10074), .ZN(n5783) );
  XNOR2_X1 U7053 ( .A(n5371), .B(n5372), .ZN(n7774) );
  NAND2_X1 U7054 ( .A1(n7774), .A2(n5591), .ZN(n5374) );
  NAND2_X1 U7055 ( .A1(n5592), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n5373) );
  OAI21_X1 U7056 ( .B1(n5407), .B2(n9824), .A(n9505), .ZN(n5376) );
  NAND2_X1 U7057 ( .A1(n5376), .A2(n5375), .ZN(n10066) );
  OR2_X1 U7058 ( .A1(n10066), .A2(n5434), .ZN(n5381) );
  INV_X1 U7059 ( .A(P1_REG2_REG_20__SCAN_IN), .ZN(n10067) );
  NAND2_X1 U7060 ( .A1(n5664), .A2(P1_REG1_REG_20__SCAN_IN), .ZN(n5378) );
  NAND2_X1 U7061 ( .A1(n5716), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n5377) );
  OAI211_X1 U7062 ( .C1(n10067), .C2(n5422), .A(n5378), .B(n5377), .ZN(n5379)
         );
  INV_X1 U7063 ( .A(n5379), .ZN(n5380) );
  AND2_X1 U7064 ( .A1(n10075), .A2(n10091), .ZN(n5838) );
  INV_X1 U7065 ( .A(n5838), .ZN(n5778) );
  NAND2_X1 U7066 ( .A1(n5384), .A2(n5383), .ZN(n5386) );
  NAND2_X1 U7067 ( .A1(n7655), .A2(n5591), .ZN(n5390) );
  NAND2_X1 U7068 ( .A1(n5388), .A2(n5387), .ZN(n5721) );
  XNOR2_X1 U7069 ( .A(n5403), .B(P1_IR_REG_18__SCAN_IN), .ZN(n9627) );
  AOI22_X1 U7070 ( .A1(n5592), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n9627), .B2(
        n5678), .ZN(n5389) );
  INV_X1 U7071 ( .A(n5391), .ZN(n5419) );
  INV_X1 U7072 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n5392) );
  NAND2_X1 U7073 ( .A1(n5419), .A2(n5392), .ZN(n5393) );
  NAND2_X1 U7074 ( .A1(n5407), .A2(n5393), .ZN(n10115) );
  OR2_X1 U7075 ( .A1(n10115), .A2(n5434), .ZN(n5398) );
  INV_X1 U7076 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n10116) );
  NAND2_X1 U7077 ( .A1(n5714), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n5395) );
  NAND2_X1 U7078 ( .A1(n5716), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n5394) );
  OAI211_X1 U7079 ( .C1(n10116), .C2(n5422), .A(n5395), .B(n5394), .ZN(n5396)
         );
  INV_X1 U7080 ( .A(n5396), .ZN(n5397) );
  NAND2_X1 U7081 ( .A1(n5400), .A2(n5399), .ZN(n5402) );
  XNOR2_X1 U7082 ( .A(n5402), .B(n5401), .ZN(n7705) );
  NAND2_X1 U7083 ( .A1(n7705), .A2(n5675), .ZN(n5406) );
  AOI22_X1 U7085 ( .A1(n9632), .A2(n5678), .B1(n5592), .B2(
        P2_DATAO_REG_19__SCAN_IN), .ZN(n5405) );
  XNOR2_X1 U7086 ( .A(n5407), .B(P1_REG3_REG_19__SCAN_IN), .ZN(n10095) );
  NAND2_X1 U7087 ( .A1(n10095), .A2(n5705), .ZN(n5412) );
  INV_X1 U7088 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n9614) );
  NAND2_X1 U7089 ( .A1(n5664), .A2(P1_REG1_REG_19__SCAN_IN), .ZN(n5409) );
  NAND2_X1 U7090 ( .A1(n5716), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n5408) );
  OAI211_X1 U7091 ( .C1(n5422), .C2(n9614), .A(n5409), .B(n5408), .ZN(n5410)
         );
  INV_X1 U7092 ( .A(n5410), .ZN(n5411) );
  OR2_X1 U7093 ( .A1(n10217), .A2(n10107), .ZN(n5843) );
  NAND2_X1 U7094 ( .A1(n10217), .A2(n10107), .ZN(n5989) );
  NAND2_X1 U7095 ( .A1(n7631), .A2(n5675), .ZN(n5417) );
  XNOR2_X1 U7096 ( .A(n5415), .B(P1_IR_REG_17__SCAN_IN), .ZN(n9626) );
  AOI22_X1 U7097 ( .A1(n5592), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n5678), .B2(
        n9626), .ZN(n5416) );
  NAND2_X1 U7098 ( .A1(n5433), .A2(n9791), .ZN(n5418) );
  AND2_X1 U7099 ( .A1(n5419), .A2(n5418), .ZN(n10137) );
  NAND2_X1 U7100 ( .A1(n10137), .A2(n5705), .ZN(n5425) );
  INV_X1 U7101 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n10128) );
  NAND2_X1 U7102 ( .A1(n5664), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n5421) );
  NAND2_X1 U7103 ( .A1(n5716), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n5420) );
  OAI211_X1 U7104 ( .C1(n10128), .C2(n5422), .A(n5421), .B(n5420), .ZN(n5423)
         );
  INV_X1 U7105 ( .A(n5423), .ZN(n5424) );
  NAND2_X1 U7106 ( .A1(n10226), .A2(n10156), .ZN(n5772) );
  NAND2_X1 U7107 ( .A1(n5987), .A2(n5772), .ZN(n10130) );
  XNOR2_X1 U7108 ( .A(n5426), .B(n5100), .ZN(n7458) );
  NAND2_X1 U7109 ( .A1(n7458), .A2(n5675), .ZN(n5429) );
  NAND2_X1 U7110 ( .A1(n5441), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5427) );
  XNOR2_X1 U7111 ( .A(n5427), .B(P1_IR_REG_16__SCAN_IN), .ZN(n10362) );
  AOI22_X1 U7112 ( .A1(n5592), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n5678), .B2(
        n10362), .ZN(n5428) );
  INV_X1 U7113 ( .A(n5430), .ZN(n5448) );
  INV_X1 U7114 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n5431) );
  NAND2_X1 U7115 ( .A1(n5448), .A2(n5431), .ZN(n5432) );
  NAND2_X1 U7116 ( .A1(n5433), .A2(n5432), .ZN(n10146) );
  OR2_X1 U7117 ( .A1(n10146), .A2(n5434), .ZN(n5437) );
  AOI22_X1 U7118 ( .A1(n5664), .A2(P1_REG1_REG_16__SCAN_IN), .B1(n5612), .B2(
        P1_REG0_REG_16__SCAN_IN), .ZN(n5436) );
  NAND2_X1 U7119 ( .A1(n5715), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n5435) );
  OR2_X1 U7120 ( .A1(n10230), .A2(n10132), .ZN(n5767) );
  XNOR2_X1 U7121 ( .A(n5439), .B(n5438), .ZN(n7455) );
  NAND2_X1 U7122 ( .A1(n7455), .A2(n5675), .ZN(n5444) );
  NAND2_X1 U7123 ( .A1(n5730), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5440) );
  MUX2_X1 U7124 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5440), .S(
        P1_IR_REG_15__SCAN_IN), .Z(n5442) );
  AND2_X1 U7125 ( .A1(n5442), .A2(n5441), .ZN(n10346) );
  AOI22_X1 U7126 ( .A1(n5592), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n5678), .B2(
        n10346), .ZN(n5443) );
  INV_X1 U7127 ( .A(n5445), .ZN(n5467) );
  INV_X1 U7128 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n5446) );
  NAND2_X1 U7129 ( .A1(n5467), .A2(n5446), .ZN(n5447) );
  AND2_X1 U7130 ( .A1(n5448), .A2(n5447), .ZN(n9561) );
  NAND2_X1 U7131 ( .A1(n9561), .A2(n5705), .ZN(n5453) );
  NAND2_X1 U7132 ( .A1(n5664), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n5450) );
  NAND2_X1 U7133 ( .A1(n5716), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n5449) );
  AND2_X1 U7134 ( .A1(n5450), .A2(n5449), .ZN(n5452) );
  NAND2_X1 U7135 ( .A1(n5715), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n5451) );
  OR2_X1 U7136 ( .A1(n8454), .A2(n10155), .ZN(n5980) );
  NAND2_X1 U7137 ( .A1(n8454), .A2(n10155), .ZN(n10151) );
  XNOR2_X1 U7138 ( .A(n5455), .B(n5454), .ZN(n7306) );
  NAND2_X1 U7139 ( .A1(n7306), .A2(n5675), .ZN(n5465) );
  NAND2_X1 U7140 ( .A1(n5456), .A2(n5457), .ZN(n5532) );
  NOR2_X1 U7141 ( .A1(P1_IR_REG_6__SCAN_IN), .A2(P1_IR_REG_5__SCAN_IN), .ZN(
        n5533) );
  NAND4_X1 U7142 ( .A1(n5533), .A2(n5640), .A3(n5458), .A4(n5536), .ZN(n5459)
         );
  NAND2_X1 U7143 ( .A1(n5518), .A2(n5460), .ZN(n5473) );
  NAND2_X1 U7144 ( .A1(n5461), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5463) );
  INV_X1 U7145 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n5462) );
  XNOR2_X1 U7146 ( .A(n5463), .B(n5462), .ZN(n9619) );
  INV_X1 U7147 ( .A(n9619), .ZN(n10334) );
  AOI22_X1 U7148 ( .A1(n10334), .A2(n5678), .B1(n5592), .B2(
        P2_DATAO_REG_14__SCAN_IN), .ZN(n5464) );
  NAND2_X1 U7149 ( .A1(n5478), .A2(n9766), .ZN(n5466) );
  AND2_X1 U7150 ( .A1(n5467), .A2(n5466), .ZN(n9420) );
  NAND2_X1 U7151 ( .A1(n9420), .A2(n5705), .ZN(n5471) );
  NAND2_X1 U7152 ( .A1(n5714), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n5470) );
  NAND2_X1 U7153 ( .A1(n5716), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n5469) );
  NAND2_X1 U7154 ( .A1(n5715), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n5468) );
  NAND2_X1 U7155 ( .A1(n8450), .A2(n8441), .ZN(n5850) );
  NAND2_X1 U7156 ( .A1(n7273), .A2(n5675), .ZN(n5476) );
  NAND2_X1 U7157 ( .A1(n5473), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5486) );
  INV_X1 U7158 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n5485) );
  NAND2_X1 U7159 ( .A1(n5486), .A2(n5485), .ZN(n5488) );
  NAND2_X1 U7160 ( .A1(n5488), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5474) );
  XNOR2_X1 U7161 ( .A(n5474), .B(P1_IR_REG_13__SCAN_IN), .ZN(n9602) );
  AOI22_X1 U7162 ( .A1(n9602), .A2(n5678), .B1(n5592), .B2(
        P2_DATAO_REG_13__SCAN_IN), .ZN(n5475) );
  NAND2_X1 U7163 ( .A1(n5714), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n5482) );
  NAND2_X1 U7164 ( .A1(n5493), .A2(n7619), .ZN(n5477) );
  AND2_X1 U7165 ( .A1(n5478), .A2(n5477), .ZN(n8283) );
  NAND2_X1 U7166 ( .A1(n5705), .A2(n8283), .ZN(n5481) );
  NAND2_X1 U7167 ( .A1(n5716), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n5480) );
  NAND2_X1 U7168 ( .A1(n5715), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n5479) );
  OR2_X1 U7169 ( .A1(n8287), .A2(n8327), .ZN(n5762) );
  NAND2_X1 U7170 ( .A1(n8287), .A2(n8327), .ZN(n5856) );
  XNOR2_X1 U7171 ( .A(n5484), .B(n5483), .ZN(n7076) );
  NAND2_X1 U7172 ( .A1(n7076), .A2(n5675), .ZN(n5490) );
  OR2_X1 U7173 ( .A1(n5486), .A2(n5485), .ZN(n5487) );
  AOI22_X1 U7174 ( .A1(n5592), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n5678), .B2(
        n7622), .ZN(n5489) );
  NAND2_X1 U7175 ( .A1(n5664), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n5497) );
  INV_X1 U7176 ( .A(n5491), .ZN(n5525) );
  INV_X1 U7177 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n9805) );
  NAND2_X1 U7178 ( .A1(n5525), .A2(n9805), .ZN(n5492) );
  AND2_X1 U7179 ( .A1(n5493), .A2(n5492), .ZN(n8324) );
  NAND2_X1 U7180 ( .A1(n5705), .A2(n8324), .ZN(n5496) );
  NAND2_X1 U7181 ( .A1(n5716), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n5495) );
  NAND2_X1 U7182 ( .A1(n5715), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n5494) );
  OR2_X1 U7183 ( .A1(n8329), .A2(n8264), .ZN(n5973) );
  NAND2_X1 U7184 ( .A1(n8329), .A2(n8264), .ZN(n5974) );
  NAND2_X1 U7185 ( .A1(n5499), .A2(n5498), .ZN(n5531) );
  AND2_X1 U7186 ( .A1(n5501), .A2(n5500), .ZN(n5530) );
  NAND2_X1 U7187 ( .A1(n5531), .A2(n5530), .ZN(n5502) );
  NAND2_X1 U7188 ( .A1(n7030), .A2(n5675), .ZN(n5509) );
  NAND2_X1 U7189 ( .A1(n5503), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5505) );
  MUX2_X1 U7190 ( .A(n5505), .B(P1_IR_REG_31__SCAN_IN), .S(n5504), .Z(n5507)
         );
  INV_X1 U7191 ( .A(n5518), .ZN(n5506) );
  AOI22_X1 U7192 ( .A1(n5592), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n5678), .B2(
        n7390), .ZN(n5508) );
  NAND2_X1 U7193 ( .A1(n5542), .A2(n5510), .ZN(n5511) );
  AND2_X1 U7194 ( .A1(n5523), .A2(n5511), .ZN(n8027) );
  NAND2_X1 U7195 ( .A1(n5705), .A2(n8027), .ZN(n5515) );
  NAND2_X1 U7196 ( .A1(n5714), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n5514) );
  NAND2_X1 U7197 ( .A1(n5716), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n5513) );
  NAND2_X1 U7198 ( .A1(n5715), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n5512) );
  NAND2_X1 U7199 ( .A1(n8066), .A2(n8207), .ZN(n5968) );
  XNOR2_X1 U7200 ( .A(n5517), .B(n5516), .ZN(n7033) );
  NAND2_X1 U7201 ( .A1(n7033), .A2(n5675), .ZN(n5521) );
  OR2_X1 U7202 ( .A1(n5518), .A2(n4918), .ZN(n5519) );
  XNOR2_X1 U7203 ( .A(n5519), .B(P1_IR_REG_11__SCAN_IN), .ZN(n7393) );
  AOI22_X1 U7204 ( .A1(n5592), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n5678), .B2(
        n7393), .ZN(n5520) );
  NAND2_X1 U7205 ( .A1(n5716), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n5529) );
  NAND2_X1 U7206 ( .A1(n5523), .A2(n5522), .ZN(n5524) );
  AND2_X1 U7207 ( .A1(n5525), .A2(n5524), .ZN(n8211) );
  NAND2_X1 U7208 ( .A1(n5705), .A2(n8211), .ZN(n5528) );
  NAND2_X1 U7209 ( .A1(n5664), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n5527) );
  NAND2_X1 U7210 ( .A1(n5715), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n5526) );
  OR2_X1 U7211 ( .A1(n10239), .A2(n8202), .ZN(n8138) );
  NAND2_X1 U7212 ( .A1(n10239), .A2(n8202), .ZN(n5971) );
  NAND2_X1 U7213 ( .A1(n7024), .A2(n5675), .ZN(n5540) );
  NAND2_X1 U7214 ( .A1(n5532), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5651) );
  OR2_X1 U7215 ( .A1(n5533), .A2(n4918), .ZN(n5534) );
  NAND2_X1 U7216 ( .A1(n5651), .A2(n5534), .ZN(n5641) );
  NAND2_X1 U7217 ( .A1(n5535), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5549) );
  NAND2_X1 U7218 ( .A1(n5549), .A2(n5536), .ZN(n5537) );
  NAND2_X1 U7219 ( .A1(n5537), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5538) );
  XNOR2_X1 U7220 ( .A(n5538), .B(P1_IR_REG_9__SCAN_IN), .ZN(n7254) );
  AOI22_X1 U7221 ( .A1(n5592), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n5678), .B2(
        n7254), .ZN(n5539) );
  NAND2_X1 U7222 ( .A1(n5540), .A2(n5539), .ZN(n8163) );
  NAND2_X1 U7223 ( .A1(n5555), .A2(n9915), .ZN(n5541) );
  AND2_X1 U7224 ( .A1(n5542), .A2(n5541), .ZN(n8162) );
  NAND2_X1 U7225 ( .A1(n5705), .A2(n8162), .ZN(n5546) );
  NAND2_X1 U7226 ( .A1(n5714), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n5545) );
  NAND2_X1 U7227 ( .A1(n5716), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n5544) );
  NAND2_X1 U7228 ( .A1(n5715), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n5543) );
  OR2_X1 U7229 ( .A1(n8163), .A2(n8026), .ZN(n5748) );
  NAND2_X1 U7230 ( .A1(n8163), .A2(n8026), .ZN(n5851) );
  NAND2_X1 U7231 ( .A1(n5748), .A2(n5851), .ZN(n7905) );
  XNOR2_X1 U7232 ( .A(n5548), .B(n5547), .ZN(n7012) );
  NAND2_X1 U7233 ( .A1(n7012), .A2(n5675), .ZN(n5551) );
  XNOR2_X1 U7234 ( .A(n5549), .B(P1_IR_REG_8__SCAN_IN), .ZN(n7082) );
  AOI22_X1 U7235 ( .A1(n5592), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n5678), .B2(
        n7082), .ZN(n5550) );
  NAND2_X1 U7236 ( .A1(n5551), .A2(n5550), .ZN(n10475) );
  NAND2_X1 U7237 ( .A1(n5664), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n5559) );
  INV_X1 U7238 ( .A(n5552), .ZN(n5634) );
  INV_X1 U7239 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n5553) );
  NAND2_X1 U7240 ( .A1(n5634), .A2(n5553), .ZN(n5554) );
  AND2_X1 U7241 ( .A1(n5555), .A2(n5554), .ZN(n8235) );
  NAND2_X1 U7242 ( .A1(n5705), .A2(n8235), .ZN(n5558) );
  NAND2_X1 U7243 ( .A1(n5716), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n5557) );
  NAND2_X1 U7244 ( .A1(n5715), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n5556) );
  NAND2_X1 U7245 ( .A1(n10475), .A2(n8008), .ZN(n7899) );
  NAND2_X1 U7246 ( .A1(n5705), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n5564) );
  NAND2_X1 U7247 ( .A1(n5611), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n5561) );
  NAND2_X1 U7248 ( .A1(n5612), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n5560) );
  AND2_X1 U7249 ( .A1(n5561), .A2(n5560), .ZN(n5563) );
  NAND2_X1 U7250 ( .A1(n5715), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n5562) );
  AND3_X2 U7251 ( .A1(n5564), .A2(n5563), .A3(n5562), .ZN(n7495) );
  INV_X1 U7252 ( .A(n5591), .ZN(n5574) );
  XNOR2_X1 U7253 ( .A(n5566), .B(n5565), .ZN(n6146) );
  INV_X1 U7254 ( .A(n6146), .ZN(n7004) );
  NAND2_X1 U7255 ( .A1(n5567), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n5573) );
  NOR2_X1 U7256 ( .A1(n5568), .A2(n4918), .ZN(n5569) );
  INV_X1 U7257 ( .A(n7059), .ZN(n5571) );
  OAI211_X1 U7258 ( .C1(n5574), .C2(n7004), .A(n5573), .B(n5572), .ZN(n5575)
         );
  NAND2_X1 U7259 ( .A1(n7495), .A2(n5575), .ZN(n5862) );
  NAND2_X1 U7260 ( .A1(n5705), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n5579) );
  NAND2_X1 U7261 ( .A1(n5611), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n5578) );
  NAND2_X1 U7262 ( .A1(n5612), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n5577) );
  NAND2_X1 U7263 ( .A1(n5715), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n5576) );
  INV_X1 U7264 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n10307) );
  INV_X1 U7265 ( .A(SI_0_), .ZN(n5581) );
  INV_X1 U7266 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n5580) );
  OAI21_X1 U7267 ( .B1(n4545), .B2(n5581), .A(n5580), .ZN(n5583) );
  NAND2_X1 U7268 ( .A1(n5583), .A2(n5582), .ZN(n10295) );
  MUX2_X1 U7269 ( .A(n10307), .B(n10295), .S(n6966), .Z(n7794) );
  INV_X1 U7270 ( .A(n7796), .ZN(n5584) );
  NAND2_X1 U7271 ( .A1(n9590), .A2(n7794), .ZN(n5860) );
  AND2_X1 U7272 ( .A1(n5584), .A2(n5860), .ZN(n7233) );
  NAND2_X1 U7273 ( .A1(n5611), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n5589) );
  INV_X1 U7274 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n5598) );
  NAND2_X1 U7275 ( .A1(n5705), .A2(n5598), .ZN(n5588) );
  NAND2_X1 U7276 ( .A1(n5612), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n5587) );
  NAND2_X1 U7277 ( .A1(n5715), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n5586) );
  XNOR2_X1 U7278 ( .A(n5605), .B(n5590), .ZN(n6995) );
  NAND2_X1 U7279 ( .A1(n5591), .A2(n6995), .ZN(n5597) );
  NAND2_X1 U7280 ( .A1(n5592), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n5596) );
  MUX2_X1 U7281 ( .A(n4918), .B(n5593), .S(P1_IR_REG_3__SCAN_IN), .Z(n5594) );
  NAND2_X1 U7282 ( .A1(n5678), .A2(n7284), .ZN(n5595) );
  NAND2_X1 U7283 ( .A1(n9588), .A2(n7979), .ZN(n7913) );
  NAND2_X1 U7284 ( .A1(n5714), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n5602) );
  XNOR2_X1 U7285 ( .A(n5598), .B(P1_REG3_REG_4__SCAN_IN), .ZN(n7923) );
  NAND2_X1 U7286 ( .A1(n5705), .A2(n7923), .ZN(n5601) );
  NAND2_X1 U7287 ( .A1(n5612), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n5600) );
  NAND2_X1 U7288 ( .A1(n5715), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n5599) );
  NAND4_X1 U7289 ( .A1(n5602), .A2(n5601), .A3(n5600), .A4(n5599), .ZN(n9587)
         );
  OR2_X1 U7290 ( .A1(n5456), .A2(n4918), .ZN(n5603) );
  XNOR2_X1 U7291 ( .A(n5603), .B(P1_IR_REG_4__SCAN_IN), .ZN(n7421) );
  AOI22_X1 U7292 ( .A1(n5592), .A2(P2_DATAO_REG_4__SCAN_IN), .B1(n5678), .B2(
        n7421), .ZN(n5610) );
  NAND2_X1 U7293 ( .A1(n5605), .A2(n5604), .ZN(n5607) );
  NAND2_X1 U7294 ( .A1(n5607), .A2(n5606), .ZN(n5645) );
  XNOR2_X1 U7295 ( .A(n5608), .B(SI_4_), .ZN(n5643) );
  XNOR2_X1 U7296 ( .A(n5645), .B(n5643), .ZN(n6996) );
  NAND2_X1 U7297 ( .A1(n6996), .A2(n5675), .ZN(n5609) );
  NAND2_X1 U7298 ( .A1(n9587), .A2(n6010), .ZN(n6008) );
  NAND2_X1 U7299 ( .A1(n7913), .A2(n6008), .ZN(n5865) );
  INV_X1 U7300 ( .A(n5865), .ZN(n5909) );
  NAND2_X1 U7301 ( .A1(n5611), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n5616) );
  NAND2_X1 U7302 ( .A1(n5705), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n5615) );
  NAND2_X1 U7303 ( .A1(n5612), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n5614) );
  INV_X1 U7304 ( .A(n10290), .ZN(n7366) );
  XNOR2_X2 U7305 ( .A(n5622), .B(n5621), .ZN(n7029) );
  NAND2_X1 U7306 ( .A1(n4545), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n5623) );
  OAI21_X1 U7307 ( .B1(n7029), .B2(n4545), .A(n5623), .ZN(n5624) );
  NAND2_X1 U7308 ( .A1(n7366), .A2(n5624), .ZN(n5631) );
  INV_X1 U7309 ( .A(n10306), .ZN(n6962) );
  NAND2_X1 U7310 ( .A1(n7029), .A2(n7001), .ZN(n5625) );
  OAI211_X1 U7311 ( .C1(n7001), .C2(P2_DATAO_REG_1__SCAN_IN), .A(n6962), .B(
        n5625), .ZN(n5630) );
  NAND2_X1 U7312 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5626) );
  MUX2_X1 U7313 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5626), .S(
        P1_IR_REG_1__SCAN_IN), .Z(n5628) );
  INV_X1 U7314 ( .A(n5568), .ZN(n5627) );
  NAND2_X1 U7315 ( .A1(n5628), .A2(n5627), .ZN(n10317) );
  INV_X1 U7316 ( .A(n10317), .ZN(n6978) );
  NAND3_X1 U7317 ( .A1(n10290), .A2(n6978), .A3(n10306), .ZN(n5629) );
  NAND2_X1 U7318 ( .A1(n5668), .A2(n5632), .ZN(n5633) );
  AND2_X1 U7319 ( .A1(n5634), .A2(n5633), .ZN(n7893) );
  NAND2_X1 U7320 ( .A1(n5705), .A2(n7893), .ZN(n5637) );
  NAND2_X1 U7321 ( .A1(n5612), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n5636) );
  NAND2_X1 U7322 ( .A1(n5715), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n5635) );
  XNOR2_X1 U7323 ( .A(n5639), .B(n5638), .ZN(n6999) );
  NOR2_X1 U7324 ( .A1(n5642), .A2(n7889), .ZN(n5684) );
  INV_X1 U7325 ( .A(n9587), .ZN(n10402) );
  NAND2_X1 U7326 ( .A1(n10402), .A2(n7924), .ZN(n6009) );
  INV_X1 U7327 ( .A(n9588), .ZN(n7440) );
  NAND2_X1 U7328 ( .A1(n7440), .A2(n7529), .ZN(n6005) );
  NAND2_X1 U7329 ( .A1(n6009), .A2(n6005), .ZN(n5663) );
  INV_X1 U7330 ( .A(n5643), .ZN(n5644) );
  NAND2_X1 U7331 ( .A1(n5645), .A2(n5644), .ZN(n5647) );
  NAND2_X1 U7332 ( .A1(n5647), .A2(n5646), .ZN(n5649) );
  NAND2_X1 U7333 ( .A1(n6998), .A2(n5675), .ZN(n5654) );
  INV_X1 U7334 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n5650) );
  NAND2_X1 U7335 ( .A1(n5651), .A2(n5650), .ZN(n5676) );
  OR2_X1 U7336 ( .A1(n5651), .A2(n5650), .ZN(n5652) );
  AOI22_X1 U7337 ( .A1(n5592), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n5678), .B2(
        n9595), .ZN(n5653) );
  NAND2_X1 U7338 ( .A1(n5714), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n5662) );
  INV_X1 U7339 ( .A(n5655), .ZN(n5666) );
  INV_X1 U7340 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n5657) );
  NAND2_X1 U7341 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .ZN(n5656) );
  NAND2_X1 U7342 ( .A1(n5657), .A2(n5656), .ZN(n5658) );
  AND2_X1 U7343 ( .A1(n5666), .A2(n5658), .ZN(n10410) );
  NAND2_X1 U7344 ( .A1(n5705), .A2(n10410), .ZN(n5661) );
  NAND2_X1 U7345 ( .A1(n5612), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n5660) );
  NAND2_X1 U7346 ( .A1(n5715), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n5659) );
  NAND4_X1 U7347 ( .A1(n5662), .A2(n5661), .A3(n5660), .A4(n5659), .ZN(n9586)
         );
  NAND2_X1 U7348 ( .A1(n10421), .A2(n9586), .ZN(n6012) );
  NAND3_X1 U7349 ( .A1(n5663), .A2(n6008), .A3(n6012), .ZN(n5682) );
  NAND2_X1 U7350 ( .A1(n5664), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n5672) );
  INV_X1 U7351 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n5665) );
  NAND2_X1 U7352 ( .A1(n5666), .A2(n5665), .ZN(n5667) );
  AND2_X1 U7353 ( .A1(n5668), .A2(n5667), .ZN(n9533) );
  NAND2_X1 U7354 ( .A1(n5705), .A2(n9533), .ZN(n5671) );
  NAND2_X1 U7355 ( .A1(n5612), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n5670) );
  NAND2_X1 U7356 ( .A1(n5715), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n5669) );
  NAND4_X1 U7357 ( .A1(n5672), .A2(n5671), .A3(n5670), .A4(n5669), .ZN(n9585)
         );
  INV_X1 U7358 ( .A(n9585), .ZN(n10404) );
  XNOR2_X1 U7359 ( .A(n5674), .B(n5673), .ZN(n6997) );
  NAND2_X1 U7360 ( .A1(n6997), .A2(n5675), .ZN(n5680) );
  NAND2_X1 U7361 ( .A1(n5676), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5677) );
  AOI22_X1 U7362 ( .A1(n5592), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n5678), .B2(
        n7087), .ZN(n5679) );
  INV_X1 U7363 ( .A(n7867), .ZN(n9531) );
  NAND2_X1 U7364 ( .A1(n10404), .A2(n9531), .ZN(n5867) );
  INV_X1 U7365 ( .A(n9586), .ZN(n7741) );
  NAND2_X1 U7366 ( .A1(n7741), .A2(n6055), .ZN(n6013) );
  AND2_X1 U7367 ( .A1(n5867), .A2(n6013), .ZN(n5681) );
  AND2_X1 U7368 ( .A1(n5682), .A2(n5681), .ZN(n5910) );
  NAND2_X1 U7369 ( .A1(n7867), .A2(n9585), .ZN(n5911) );
  NAND2_X1 U7370 ( .A1(n6012), .A2(n5911), .ZN(n5683) );
  NAND2_X1 U7371 ( .A1(n5683), .A2(n5867), .ZN(n5908) );
  NAND4_X1 U7372 ( .A1(n7962), .A2(n5684), .A3(n5910), .A4(n5908), .ZN(n5685)
         );
  NOR2_X1 U7373 ( .A1(n7905), .A2(n5685), .ZN(n5686) );
  NAND4_X1 U7374 ( .A1(n8139), .A2(n8068), .A3(n8035), .A4(n5686), .ZN(n5687)
         );
  NOR2_X1 U7375 ( .A1(n6024), .A2(n5687), .ZN(n5688) );
  NAND4_X1 U7376 ( .A1(n10143), .A2(n8337), .A3(n8216), .A4(n5688), .ZN(n5689)
         );
  NOR2_X1 U7377 ( .A1(n10130), .A2(n5689), .ZN(n5690) );
  NAND4_X1 U7378 ( .A1(n10070), .A2(n10111), .A3(n10086), .A4(n5690), .ZN(
        n5691) );
  NOR2_X1 U7379 ( .A1(n10050), .A2(n5691), .ZN(n5692) );
  NAND4_X1 U7380 ( .A1(n9727), .A2(n8430), .A3(n10021), .A4(n5692), .ZN(n5693)
         );
  NOR2_X1 U7381 ( .A1(n9697), .A2(n5693), .ZN(n5694) );
  XNOR2_X1 U7382 ( .A(n5697), .B(n5696), .ZN(n5698) );
  NAND2_X1 U7383 ( .A1(n8640), .A2(n5591), .ZN(n5701) );
  NAND2_X1 U7384 ( .A1(n5592), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n5700) );
  INV_X1 U7385 ( .A(n9656), .ZN(n5706) );
  INV_X1 U7386 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n6692) );
  NAND2_X1 U7387 ( .A1(n5715), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n5703) );
  NAND2_X1 U7388 ( .A1(n5716), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n5702) );
  OAI211_X1 U7389 ( .C1(n6692), .C2(n5585), .A(n5703), .B(n5702), .ZN(n5704)
         );
  AOI21_X1 U7390 ( .B1(n5706), .B2(n5705), .A(n5704), .ZN(n8610) );
  OR2_X1 U7391 ( .A1(n6058), .A2(n8610), .ZN(n5895) );
  NAND2_X1 U7392 ( .A1(n6058), .A2(n8610), .ZN(n5896) );
  NAND2_X1 U7393 ( .A1(n5708), .A2(n5707), .ZN(n5711) );
  XNOR2_X1 U7394 ( .A(n5709), .B(SI_30_), .ZN(n5710) );
  NAND2_X1 U7395 ( .A1(n8627), .A2(n5591), .ZN(n5713) );
  NAND2_X1 U7396 ( .A1(n5592), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n5712) );
  NAND2_X1 U7397 ( .A1(n5714), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n5719) );
  NAND2_X1 U7398 ( .A1(n5715), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n5718) );
  NAND2_X1 U7399 ( .A1(n5716), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n5717) );
  AND3_X1 U7400 ( .A1(n5719), .A2(n5718), .A3(n5717), .ZN(n6002) );
  NOR2_X1 U7401 ( .A1(n9646), .A2(n6002), .ZN(n5820) );
  AOI21_X1 U7402 ( .B1(n5720), .B2(n9642), .A(n5820), .ZN(n5900) );
  INV_X1 U7403 ( .A(n5721), .ZN(n5726) );
  AOI21_X1 U7404 ( .B1(n5728), .B2(n5900), .A(n6949), .ZN(n5941) );
  NAND2_X1 U7405 ( .A1(n5941), .A2(n9632), .ZN(n5903) );
  INV_X1 U7406 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n5734) );
  NAND2_X1 U7407 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(P1_IR_REG_21__SCAN_IN), 
        .ZN(n5732) );
  NAND2_X1 U7408 ( .A1(n5732), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5733) );
  OAI21_X1 U7409 ( .B1(n5734), .B2(P1_IR_REG_31__SCAN_IN), .A(n5733), .ZN(
        n5735) );
  MUX2_X1 U7410 ( .A(n5837), .B(n5999), .S(n7994), .Z(n5814) );
  INV_X1 U7411 ( .A(n5888), .ZN(n5805) );
  INV_X1 U7412 ( .A(n6009), .ZN(n5740) );
  NAND2_X1 U7413 ( .A1(n5744), .A2(n6012), .ZN(n7843) );
  NAND2_X1 U7414 ( .A1(n7843), .A2(n7842), .ZN(n5742) );
  AND2_X1 U7415 ( .A1(n5913), .A2(n5911), .ZN(n5741) );
  INV_X1 U7416 ( .A(n5867), .ZN(n5743) );
  NAND2_X1 U7417 ( .A1(n5745), .A2(n7900), .ZN(n5749) );
  NAND2_X1 U7418 ( .A1(n5749), .A2(n7899), .ZN(n5746) );
  NAND2_X1 U7419 ( .A1(n5746), .A2(n5748), .ZN(n5747) );
  NAND2_X1 U7420 ( .A1(n5748), .A2(n7900), .ZN(n5871) );
  INV_X1 U7421 ( .A(n5871), .ZN(n5964) );
  AOI21_X1 U7422 ( .B1(n5749), .B2(n5964), .A(n5965), .ZN(n5750) );
  MUX2_X1 U7423 ( .A(n8207), .B(n4900), .S(n6950), .Z(n5752) );
  INV_X1 U7424 ( .A(n8207), .ZN(n9582) );
  OR2_X1 U7425 ( .A1(n8066), .A2(n9582), .ZN(n8032) );
  NAND2_X1 U7426 ( .A1(n5752), .A2(n8032), .ZN(n5751) );
  INV_X1 U7427 ( .A(n5752), .ZN(n5753) );
  OAI21_X1 U7428 ( .B1(n4900), .B2(n8207), .A(n5753), .ZN(n5754) );
  AND2_X1 U7429 ( .A1(n8035), .A2(n5754), .ZN(n5755) );
  NAND2_X1 U7430 ( .A1(n5974), .A2(n5971), .ZN(n5854) );
  INV_X1 U7431 ( .A(n5974), .ZN(n5757) );
  INV_X1 U7432 ( .A(n5973), .ZN(n5756) );
  MUX2_X1 U7433 ( .A(n5757), .B(n5756), .S(n7994), .Z(n5759) );
  INV_X1 U7434 ( .A(n8216), .ZN(n6027) );
  INV_X1 U7435 ( .A(n5856), .ZN(n5978) );
  NOR2_X1 U7436 ( .A1(n6027), .A2(n5978), .ZN(n5758) );
  NAND2_X1 U7437 ( .A1(n8338), .A2(n5762), .ZN(n5877) );
  NAND2_X1 U7438 ( .A1(n5973), .A2(n8138), .ZN(n5873) );
  INV_X1 U7439 ( .A(n5873), .ZN(n5760) );
  INV_X1 U7440 ( .A(n5762), .ZN(n5763) );
  NAND2_X1 U7441 ( .A1(n5983), .A2(n10151), .ZN(n5765) );
  NAND2_X1 U7442 ( .A1(n5767), .A2(n5980), .ZN(n5881) );
  MUX2_X1 U7443 ( .A(n5765), .B(n5881), .S(n6950), .Z(n5766) );
  INV_X1 U7444 ( .A(n5766), .ZN(n5770) );
  INV_X1 U7445 ( .A(n5767), .ZN(n5768) );
  MUX2_X1 U7446 ( .A(n5848), .B(n5768), .S(n7994), .Z(n5769) );
  NAND2_X1 U7447 ( .A1(n10226), .A2(n10104), .ZN(n6034) );
  OAI21_X1 U7448 ( .B1(n6950), .B2(n10104), .A(n6034), .ZN(n5774) );
  NAND2_X1 U7449 ( .A1(n5776), .A2(n5772), .ZN(n5849) );
  AND2_X1 U7450 ( .A1(n5849), .A2(n7994), .ZN(n5773) );
  AND2_X1 U7451 ( .A1(n10087), .A2(n5987), .ZN(n5841) );
  NAND3_X1 U7452 ( .A1(n5781), .A2(n5989), .A3(n5776), .ZN(n5777) );
  NAND2_X1 U7453 ( .A1(n5777), .A2(n5843), .ZN(n5780) );
  NAND2_X1 U7454 ( .A1(n5991), .A2(n5783), .ZN(n5840) );
  INV_X1 U7455 ( .A(n5840), .ZN(n5779) );
  NAND4_X1 U7456 ( .A1(n5780), .A2(n6950), .A3(n5779), .A4(n5778), .ZN(n5801)
         );
  NAND2_X1 U7457 ( .A1(n5782), .A2(n10098), .ZN(n5790) );
  INV_X1 U7458 ( .A(n8426), .ZN(n5784) );
  OAI21_X1 U7459 ( .B1(n10050), .B2(n5784), .A(n5783), .ZN(n5785) );
  AND2_X1 U7460 ( .A1(n5785), .A2(n5795), .ZN(n5793) );
  INV_X1 U7461 ( .A(n5786), .ZN(n5787) );
  NAND2_X1 U7462 ( .A1(n5787), .A2(n10087), .ZN(n5788) );
  INV_X1 U7463 ( .A(n10107), .ZN(n10071) );
  NAND2_X1 U7464 ( .A1(n5788), .A2(n10071), .ZN(n5789) );
  NAND4_X1 U7465 ( .A1(n5790), .A2(n5793), .A3(n7994), .A4(n5789), .ZN(n5800)
         );
  INV_X1 U7466 ( .A(n10070), .ZN(n6037) );
  NAND2_X1 U7467 ( .A1(n8426), .A2(n6950), .ZN(n5791) );
  NAND2_X1 U7468 ( .A1(n6037), .A2(n5791), .ZN(n5792) );
  NAND2_X1 U7469 ( .A1(n10048), .A2(n5792), .ZN(n5798) );
  INV_X1 U7470 ( .A(n5793), .ZN(n5794) );
  NAND3_X1 U7471 ( .A1(n5794), .A2(n7994), .A3(n5991), .ZN(n5797) );
  NAND3_X1 U7472 ( .A1(n5840), .A2(n6950), .A3(n5795), .ZN(n5796) );
  OAI211_X1 U7473 ( .C1(n8424), .C2(n5798), .A(n5797), .B(n5796), .ZN(n5799)
         );
  NAND3_X1 U7474 ( .A1(n5801), .A2(n5800), .A3(n5799), .ZN(n5804) );
  NAND2_X1 U7475 ( .A1(n5888), .A2(n9717), .ZN(n5815) );
  AND2_X1 U7476 ( .A1(n5993), .A2(n5923), .ZN(n5886) );
  INV_X1 U7477 ( .A(n5886), .ZN(n5802) );
  NOR2_X1 U7478 ( .A1(n5815), .A2(n5802), .ZN(n5803) );
  NAND2_X1 U7479 ( .A1(n5804), .A2(n5803), .ZN(n5816) );
  NAND3_X1 U7480 ( .A1(n9690), .A2(n9699), .A3(n6950), .ZN(n5807) );
  OAI21_X1 U7481 ( .B1(n5836), .B2(n7994), .A(n5807), .ZN(n5808) );
  NAND2_X1 U7482 ( .A1(n5808), .A2(n5998), .ZN(n5811) );
  INV_X1 U7483 ( .A(n5928), .ZN(n5809) );
  NAND3_X1 U7484 ( .A1(n5836), .A2(n5809), .A3(n7994), .ZN(n5810) );
  OAI211_X1 U7485 ( .C1(n4406), .C2(n5998), .A(n5811), .B(n5810), .ZN(n5812)
         );
  NAND2_X1 U7486 ( .A1(n5812), .A2(n6875), .ZN(n5813) );
  INV_X1 U7487 ( .A(n5815), .ZN(n5926) );
  OAI211_X1 U7488 ( .C1(n4611), .C2(n5926), .A(n5816), .B(n9682), .ZN(n5817)
         );
  NAND2_X1 U7489 ( .A1(n5817), .A2(n5890), .ZN(n5819) );
  NOR2_X1 U7490 ( .A1(n9683), .A2(n7994), .ZN(n5818) );
  INV_X1 U7491 ( .A(n5820), .ZN(n5821) );
  NAND2_X1 U7492 ( .A1(n5821), .A2(n9641), .ZN(n5822) );
  NAND2_X1 U7493 ( .A1(n5822), .A2(n9642), .ZN(n5939) );
  NAND3_X1 U7494 ( .A1(n5823), .A2(n6904), .A3(n5939), .ZN(n5830) );
  AND2_X1 U7495 ( .A1(n5279), .A2(n9632), .ZN(n5829) );
  NAND2_X1 U7496 ( .A1(n6949), .A2(n7994), .ZN(n5824) );
  INV_X1 U7497 ( .A(n6002), .ZN(n9565) );
  NAND2_X1 U7498 ( .A1(n9565), .A2(n9641), .ZN(n5826) );
  NAND2_X1 U7499 ( .A1(n9646), .A2(n5826), .ZN(n5827) );
  NAND2_X1 U7500 ( .A1(n5827), .A2(n5896), .ZN(n5933) );
  NAND2_X1 U7501 ( .A1(n5939), .A2(n5933), .ZN(n5828) );
  NAND2_X1 U7502 ( .A1(n5831), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5833) );
  NAND2_X1 U7503 ( .A1(n9632), .A2(n7806), .ZN(n7791) );
  NAND2_X1 U7504 ( .A1(n5998), .A2(n5834), .ZN(n5835) );
  NAND3_X1 U7505 ( .A1(n5837), .A2(n5836), .A3(n5835), .ZN(n5931) );
  AND2_X1 U7506 ( .A1(n8427), .A2(n5838), .ZN(n5839) );
  NAND2_X1 U7507 ( .A1(n5845), .A2(n5989), .ZN(n5905) );
  OR3_X1 U7508 ( .A1(n5905), .A2(n5842), .A3(n5841), .ZN(n5847) );
  NAND3_X1 U7509 ( .A1(n8427), .A2(n8426), .A3(n5843), .ZN(n5844) );
  AOI21_X1 U7510 ( .B1(n5845), .B2(n5844), .A(n5960), .ZN(n5846) );
  NAND2_X1 U7511 ( .A1(n5847), .A2(n5846), .ZN(n5925) );
  OR2_X1 U7512 ( .A1(n5849), .A2(n5848), .ZN(n5883) );
  NAND2_X1 U7513 ( .A1(n10151), .A2(n5850), .ZN(n5876) );
  NAND2_X1 U7514 ( .A1(n5968), .A2(n5851), .ZN(n5852) );
  AND2_X1 U7515 ( .A1(n5852), .A2(n8033), .ZN(n5853) );
  NOR2_X1 U7516 ( .A1(n5854), .A2(n5853), .ZN(n5870) );
  NAND4_X1 U7517 ( .A1(n5870), .A2(n5856), .A3(n5855), .A4(n7899), .ZN(n5857)
         );
  OR2_X1 U7518 ( .A1(n5876), .A2(n5857), .ZN(n5858) );
  NOR2_X1 U7519 ( .A1(n5883), .A2(n5858), .ZN(n5906) );
  NAND2_X1 U7520 ( .A1(n5737), .A2(n6054), .ZN(n5859) );
  NAND3_X1 U7521 ( .A1(n5860), .A2(n6949), .A3(n5859), .ZN(n5861) );
  NAND2_X1 U7522 ( .A1(n5862), .A2(n5861), .ZN(n5864) );
  OAI21_X1 U7523 ( .B1(n7348), .B2(n5864), .A(n5863), .ZN(n5866) );
  AOI21_X1 U7524 ( .B1(n5866), .B2(n6005), .A(n5865), .ZN(n5869) );
  NAND3_X1 U7525 ( .A1(n5867), .A2(n6013), .A3(n6009), .ZN(n5868) );
  OAI211_X1 U7526 ( .C1(n5869), .C2(n5868), .A(n5913), .B(n5908), .ZN(n5884)
         );
  INV_X1 U7527 ( .A(n8033), .ZN(n5872) );
  OAI21_X1 U7528 ( .B1(n5872), .B2(n5871), .A(n5870), .ZN(n5875) );
  NAND2_X1 U7529 ( .A1(n5873), .A2(n5974), .ZN(n5874) );
  AOI21_X1 U7530 ( .B1(n5875), .B2(n5874), .A(n5978), .ZN(n5878) );
  INV_X1 U7531 ( .A(n5876), .ZN(n5979) );
  OAI21_X1 U7532 ( .B1(n5878), .B2(n5877), .A(n5979), .ZN(n5879) );
  INV_X1 U7533 ( .A(n5879), .ZN(n5880) );
  NOR2_X1 U7534 ( .A1(n5881), .A2(n5880), .ZN(n5882) );
  NOR2_X1 U7535 ( .A1(n5883), .A2(n5882), .ZN(n5917) );
  AOI21_X1 U7536 ( .B1(n5906), .B2(n5884), .A(n5917), .ZN(n5885) );
  OAI21_X1 U7537 ( .B1(n5905), .B2(n5885), .A(n9717), .ZN(n5887) );
  OAI21_X1 U7538 ( .B1(n5925), .B2(n5887), .A(n5886), .ZN(n5889) );
  NAND3_X1 U7539 ( .A1(n5889), .A2(n9682), .A3(n5888), .ZN(n5891) );
  NAND2_X1 U7540 ( .A1(n5891), .A2(n5890), .ZN(n5892) );
  NAND2_X1 U7541 ( .A1(n5892), .A2(n5928), .ZN(n5893) );
  NOR2_X1 U7542 ( .A1(n9669), .A2(n5893), .ZN(n5894) );
  NOR2_X1 U7543 ( .A1(n5931), .A2(n5894), .ZN(n5898) );
  NAND2_X1 U7544 ( .A1(n5895), .A2(n5999), .ZN(n5935) );
  OAI211_X1 U7545 ( .C1(n5898), .C2(n5935), .A(n5897), .B(n5896), .ZN(n5899)
         );
  MUX2_X1 U7546 ( .A(n7791), .B(n6951), .S(n5901), .Z(n5904) );
  NAND2_X1 U7547 ( .A1(n5942), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5902) );
  AND2_X1 U7548 ( .A1(n6902), .A2(P1_STATE_REG_SCAN_IN), .ZN(n8130) );
  INV_X1 U7549 ( .A(n7806), .ZN(n6059) );
  INV_X1 U7550 ( .A(n8130), .ZN(n5953) );
  NOR3_X1 U7551 ( .A1(n5956), .A2(n6059), .A3(n5953), .ZN(n5957) );
  INV_X1 U7552 ( .A(n5905), .ZN(n5922) );
  INV_X1 U7553 ( .A(n5906), .ZN(n5920) );
  NAND3_X1 U7554 ( .A1(n5907), .A2(n5909), .A3(n5908), .ZN(n5916) );
  INV_X1 U7555 ( .A(n5910), .ZN(n5912) );
  NAND2_X1 U7556 ( .A1(n5912), .A2(n5911), .ZN(n5915) );
  INV_X1 U7557 ( .A(n5913), .ZN(n5914) );
  AOI21_X1 U7558 ( .B1(n5916), .B2(n5915), .A(n5914), .ZN(n5919) );
  INV_X1 U7559 ( .A(n5917), .ZN(n5918) );
  OAI21_X1 U7560 ( .B1(n5920), .B2(n5919), .A(n5918), .ZN(n5921) );
  AND2_X1 U7561 ( .A1(n5922), .A2(n5921), .ZN(n5924) );
  OAI21_X1 U7562 ( .B1(n5925), .B2(n5924), .A(n5923), .ZN(n5927) );
  AOI21_X1 U7563 ( .B1(n5927), .B2(n5926), .A(n4445), .ZN(n5930) );
  NAND2_X1 U7564 ( .A1(n5928), .A2(n9682), .ZN(n5929) );
  NOR2_X1 U7565 ( .A1(n5930), .A2(n5929), .ZN(n5932) );
  AOI21_X1 U7566 ( .B1(n5932), .B2(n5998), .A(n5931), .ZN(n5936) );
  INV_X1 U7567 ( .A(n5933), .ZN(n5934) );
  OAI21_X1 U7568 ( .B1(n5936), .B2(n5935), .A(n5934), .ZN(n5938) );
  AOI211_X1 U7569 ( .C1(n5939), .C2(n5938), .A(n7930), .B(n5937), .ZN(n5940)
         );
  NAND2_X1 U7570 ( .A1(n5951), .A2(n5950), .ZN(n5943) );
  XNOR2_X1 U7571 ( .A(n5950), .B(n5951), .ZN(n8334) );
  NAND2_X1 U7572 ( .A1(n7360), .A2(n10428), .ZN(n7364) );
  NOR3_X1 U7573 ( .A1(n7364), .A2(n10290), .A3(n10306), .ZN(n5955) );
  OAI21_X1 U7574 ( .B1(n6950), .B2(n5953), .A(P1_B_REG_SCAN_IN), .ZN(n5954) );
  INV_X1 U7575 ( .A(P1_B_REG_SCAN_IN), .ZN(n5958) );
  NOR2_X1 U7576 ( .A1(n10306), .A2(n5958), .ZN(n5959) );
  OR2_X1 U7577 ( .A1(n10405), .A2(n5959), .ZN(n9639) );
  INV_X1 U7578 ( .A(n8427), .ZN(n5961) );
  INV_X1 U7579 ( .A(n5963), .ZN(n5962) );
  AND2_X1 U7580 ( .A1(n8426), .A2(n5963), .ZN(n5990) );
  INV_X1 U7581 ( .A(n5965), .ZN(n5966) );
  NAND2_X1 U7582 ( .A1(n5967), .A2(n5966), .ZN(n8069) );
  AND3_X1 U7583 ( .A1(n5973), .A2(n8033), .A3(n8138), .ZN(n5970) );
  INV_X1 U7584 ( .A(n5971), .ZN(n5972) );
  NAND2_X1 U7585 ( .A1(n5973), .A2(n5972), .ZN(n5975) );
  AND2_X1 U7586 ( .A1(n5975), .A2(n5974), .ZN(n5976) );
  NAND2_X1 U7587 ( .A1(n5980), .A2(n8338), .ZN(n5981) );
  NAND2_X1 U7588 ( .A1(n5981), .A2(n10151), .ZN(n5982) );
  NAND2_X1 U7589 ( .A1(n5984), .A2(n5983), .ZN(n10131) );
  NAND2_X2 U7590 ( .A1(n10135), .A2(n5987), .ZN(n10102) );
  AND2_X1 U7591 ( .A1(n10086), .A2(n10087), .ZN(n5988) );
  AND2_X1 U7592 ( .A1(n9727), .A2(n9717), .ZN(n5992) );
  AND2_X1 U7593 ( .A1(n5995), .A2(n9682), .ZN(n5996) );
  NAND2_X1 U7594 ( .A1(n9685), .A2(n5997), .ZN(n9670) );
  NAND2_X1 U7595 ( .A1(n6876), .A2(n6875), .ZN(n6878) );
  NAND2_X1 U7596 ( .A1(n9632), .A2(n6950), .ZN(n6001) );
  NAND2_X1 U7597 ( .A1(n6949), .A2(n6059), .ZN(n6000) );
  INV_X1 U7598 ( .A(n7794), .ZN(n7235) );
  AND2_X1 U7599 ( .A1(n9590), .A2(n7235), .ZN(n7790) );
  NAND2_X1 U7600 ( .A1(n7495), .A2(n4391), .ZN(n6003) );
  NAND2_X1 U7601 ( .A1(n6004), .A2(n6003), .ZN(n7377) );
  NAND2_X1 U7602 ( .A1(n6005), .A2(n7913), .ZN(n7380) );
  NAND2_X1 U7603 ( .A1(n7377), .A2(n7380), .ZN(n6007) );
  NAND2_X1 U7604 ( .A1(n7440), .A2(n7979), .ZN(n6006) );
  NAND2_X1 U7605 ( .A1(n6007), .A2(n6006), .ZN(n7919) );
  NAND2_X1 U7606 ( .A1(n6009), .A2(n6008), .ZN(n7920) );
  NAND2_X1 U7607 ( .A1(n10402), .A2(n6010), .ZN(n6011) );
  NAND2_X1 U7608 ( .A1(n6055), .A2(n9586), .ZN(n6015) );
  NAND2_X1 U7609 ( .A1(n10412), .A2(n6015), .ZN(n7834) );
  NAND2_X1 U7610 ( .A1(n10404), .A2(n7867), .ZN(n6017) );
  OR2_X1 U7611 ( .A1(n4756), .A2(n7894), .ZN(n6018) );
  OR2_X1 U7612 ( .A1(n8163), .A2(n9583), .ZN(n6019) );
  INV_X1 U7613 ( .A(n8264), .ZN(n9580) );
  NAND2_X1 U7614 ( .A1(n8329), .A2(n9580), .ZN(n8170) );
  NAND2_X1 U7615 ( .A1(n10239), .A2(n9581), .ZN(n8167) );
  NAND2_X1 U7616 ( .A1(n8032), .A2(n9581), .ZN(n6020) );
  INV_X1 U7617 ( .A(n10239), .ZN(n8208) );
  NAND2_X1 U7618 ( .A1(n6020), .A2(n8208), .ZN(n6021) );
  OAI21_X1 U7619 ( .B1(n8032), .B2(n9581), .A(n6021), .ZN(n6022) );
  OR2_X1 U7620 ( .A1(n8139), .A2(n6022), .ZN(n8171) );
  NAND2_X1 U7621 ( .A1(n8171), .A2(n8170), .ZN(n6023) );
  INV_X1 U7622 ( .A(n8327), .ZN(n9579) );
  NAND2_X1 U7623 ( .A1(n8287), .A2(n9579), .ZN(n6025) );
  INV_X1 U7624 ( .A(n8441), .ZN(n9578) );
  NAND2_X1 U7625 ( .A1(n8450), .A2(n9578), .ZN(n6028) );
  NAND2_X1 U7626 ( .A1(n8335), .A2(n4782), .ZN(n6030) );
  INV_X1 U7627 ( .A(n10155), .ZN(n9577) );
  NAND2_X1 U7628 ( .A1(n8454), .A2(n9577), .ZN(n6029) );
  INV_X1 U7629 ( .A(n10143), .ZN(n10153) );
  INV_X1 U7630 ( .A(n10132), .ZN(n9575) );
  NAND2_X1 U7631 ( .A1(n10230), .A2(n9575), .ZN(n6031) );
  OR2_X1 U7632 ( .A1(n10226), .A2(n10104), .ZN(n6033) );
  NAND2_X1 U7633 ( .A1(n10114), .A2(n9574), .ZN(n10082) );
  OAI22_X1 U7634 ( .A1(n10086), .A2(n10082), .B1(n10107), .B2(n10098), .ZN(
        n6036) );
  NAND2_X1 U7635 ( .A1(n10046), .A2(n6038), .ZN(n6040) );
  INV_X1 U7636 ( .A(n10091), .ZN(n9573) );
  AND2_X1 U7637 ( .A1(n10075), .A2(n9573), .ZN(n10047) );
  INV_X1 U7638 ( .A(n10074), .ZN(n9572) );
  AOI22_X1 U7639 ( .A1(n10050), .A2(n10047), .B1(n9572), .B2(n10061), .ZN(
        n6039) );
  NAND2_X1 U7640 ( .A1(n8425), .A2(n8424), .ZN(n8423) );
  NAND2_X1 U7641 ( .A1(n5346), .A2(n10022), .ZN(n6041) );
  OR2_X1 U7642 ( .A1(n10201), .A2(n9571), .ZN(n6042) );
  NAND2_X1 U7643 ( .A1(n10201), .A2(n9571), .ZN(n6043) );
  INV_X1 U7644 ( .A(n9727), .ZN(n6044) );
  NAND2_X1 U7645 ( .A1(n9729), .A2(n9570), .ZN(n6045) );
  INV_X1 U7646 ( .A(n9711), .ZN(n6047) );
  INV_X1 U7647 ( .A(n9722), .ZN(n9569) );
  OR2_X1 U7648 ( .A1(n10190), .A2(n9569), .ZN(n6048) );
  NOR2_X1 U7649 ( .A1(n9690), .A2(n9568), .ZN(n6049) );
  NAND2_X1 U7650 ( .A1(n9690), .A2(n9568), .ZN(n6050) );
  INV_X1 U7651 ( .A(n9687), .ZN(n9567) );
  INV_X1 U7652 ( .A(n9671), .ZN(n9566) );
  NAND2_X1 U7653 ( .A1(n8619), .A2(n9566), .ZN(n9652) );
  AND2_X1 U7654 ( .A1(n6051), .A2(n5086), .ZN(n6052) );
  NAND2_X1 U7655 ( .A1(n9653), .A2(n6052), .ZN(n6064) );
  NAND2_X1 U7656 ( .A1(n7794), .A2(n6054), .ZN(n7793) );
  INV_X1 U7657 ( .A(n4391), .ZN(n7435) );
  NOR2_X2 U7658 ( .A1(n7793), .A2(n5575), .ZN(n7378) );
  NAND2_X1 U7659 ( .A1(n7378), .A2(n7979), .ZN(n7921) );
  OR2_X2 U7660 ( .A1(n8146), .A2(n8329), .ZN(n8180) );
  AND2_X2 U7661 ( .A1(n10127), .A2(n10270), .ZN(n10112) );
  NAND2_X1 U7662 ( .A1(n10112), .A2(n10098), .ZN(n10092) );
  NOR2_X2 U7663 ( .A1(n6883), .A2(n6058), .ZN(n9637) );
  NOR2_X2 U7664 ( .A1(n7359), .A2(n6059), .ZN(n10418) );
  NAND2_X1 U7665 ( .A1(n6883), .A2(n6058), .ZN(n6060) );
  NAND3_X1 U7666 ( .A1(n9647), .A2(n10418), .A3(n6060), .ZN(n9660) );
  INV_X1 U7667 ( .A(n9652), .ZN(n6061) );
  NAND3_X1 U7668 ( .A1(n4709), .A2(n6061), .A3(n10489), .ZN(n6062) );
  NAND2_X1 U7669 ( .A1(n6064), .A2(n6063), .ZN(n6065) );
  INV_X1 U7670 ( .A(n6067), .ZN(n6070) );
  NAND2_X1 U7671 ( .A1(n8405), .A2(P1_B_REG_SCAN_IN), .ZN(n6068) );
  MUX2_X1 U7672 ( .A(P1_B_REG_SCAN_IN), .B(n6068), .S(n8334), .Z(n6069) );
  INV_X1 U7673 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n6071) );
  NAND2_X1 U7674 ( .A1(n10427), .A2(n6071), .ZN(n6073) );
  NAND2_X1 U7675 ( .A1(n6067), .A2(n8334), .ZN(n6072) );
  NAND2_X1 U7676 ( .A1(n7367), .A2(n6951), .ZN(n7496) );
  NAND2_X1 U7677 ( .A1(n7358), .A2(n7363), .ZN(n7510) );
  INV_X1 U7678 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n7009) );
  NAND2_X1 U7679 ( .A1(n10427), .A2(n7009), .ZN(n6075) );
  NAND2_X1 U7680 ( .A1(n6067), .A2(n8405), .ZN(n6074) );
  NAND2_X1 U7681 ( .A1(n6075), .A2(n6074), .ZN(n7356) );
  NOR4_X1 U7682 ( .A1(P1_D_REG_15__SCAN_IN), .A2(P1_D_REG_17__SCAN_IN), .A3(
        P1_D_REG_18__SCAN_IN), .A4(P1_D_REG_19__SCAN_IN), .ZN(n6079) );
  NOR4_X1 U7683 ( .A1(P1_D_REG_10__SCAN_IN), .A2(P1_D_REG_12__SCAN_IN), .A3(
        P1_D_REG_16__SCAN_IN), .A4(P1_D_REG_14__SCAN_IN), .ZN(n6078) );
  NOR4_X1 U7684 ( .A1(P1_D_REG_25__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_29__SCAN_IN), .ZN(n6077) );
  NOR4_X1 U7685 ( .A1(P1_D_REG_20__SCAN_IN), .A2(P1_D_REG_24__SCAN_IN), .A3(
        P1_D_REG_22__SCAN_IN), .A4(P1_D_REG_23__SCAN_IN), .ZN(n6076) );
  NAND4_X1 U7686 ( .A1(n6079), .A2(n6078), .A3(n6077), .A4(n6076), .ZN(n6084)
         );
  NOR2_X1 U7687 ( .A1(P1_D_REG_11__SCAN_IN), .A2(P1_D_REG_21__SCAN_IN), .ZN(
        n9763) );
  NOR4_X1 U7688 ( .A1(P1_D_REG_30__SCAN_IN), .A2(P1_D_REG_31__SCAN_IN), .A3(
        P1_D_REG_7__SCAN_IN), .A4(P1_D_REG_26__SCAN_IN), .ZN(n6082) );
  NOR4_X1 U7689 ( .A1(P1_D_REG_5__SCAN_IN), .A2(P1_D_REG_6__SCAN_IN), .A3(
        P1_D_REG_8__SCAN_IN), .A4(P1_D_REG_9__SCAN_IN), .ZN(n6081) );
  NOR4_X1 U7690 ( .A1(P1_D_REG_13__SCAN_IN), .A2(P1_D_REG_2__SCAN_IN), .A3(
        P1_D_REG_3__SCAN_IN), .A4(P1_D_REG_4__SCAN_IN), .ZN(n6080) );
  NAND4_X1 U7691 ( .A1(n9763), .A2(n6082), .A3(n6081), .A4(n6080), .ZN(n6083)
         );
  OAI21_X1 U7692 ( .B1(n6084), .B2(n6083), .A(n10427), .ZN(n7355) );
  OAI211_X1 U7693 ( .C1(n6949), .C2(n10473), .A(n7356), .B(n7355), .ZN(n6688)
         );
  INV_X1 U7694 ( .A(n6058), .ZN(n6691) );
  INV_X1 U7695 ( .A(n7359), .ZN(n7234) );
  INV_X1 U7696 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n6085) );
  INV_X1 U7697 ( .A(n6086), .ZN(n6087) );
  OAI21_X1 U7698 ( .B1(n6695), .B2(n10490), .A(n6087), .ZN(P1_U3520) );
  NOR2_X2 U7699 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n6145) );
  NOR2_X1 U7700 ( .A1(P2_IR_REG_3__SCAN_IN), .A2(P2_IR_REG_2__SCAN_IN), .ZN(
        n6088) );
  NOR2_X1 U7701 ( .A1(P2_IR_REG_9__SCAN_IN), .A2(P2_IR_REG_5__SCAN_IN), .ZN(
        n6093) );
  NAND4_X1 U7702 ( .A1(n6093), .A2(n6092), .A3(n6091), .A4(n6090), .ZN(n6096)
         );
  NAND4_X1 U7703 ( .A1(n6094), .A2(n6269), .A3(n6222), .A4(n6329), .ZN(n6095)
         );
  NOR2_X2 U7704 ( .A1(n6096), .A2(n6095), .ZN(n6097) );
  INV_X2 U7705 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n6492) );
  NOR2_X1 U7706 ( .A1(P2_IR_REG_23__SCAN_IN), .A2(P2_IR_REG_25__SCAN_IN), .ZN(
        n6099) );
  INV_X1 U7707 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n6100) );
  AOI21_X1 U7708 ( .B1(n6683), .B2(P2_IR_REG_28__SCAN_IN), .A(n6101), .ZN(
        n6103) );
  OR2_X2 U7709 ( .A1(n6683), .A2(P2_IR_REG_27__SCAN_IN), .ZN(n6102) );
  NAND2_X4 U7710 ( .A1(n6103), .A2(n6102), .ZN(n7103) );
  NAND2_X1 U7711 ( .A1(n7103), .A2(n4545), .ZN(n6131) );
  NAND2_X1 U7712 ( .A1(n8627), .A2(n6351), .ZN(n6105) );
  NAND2_X2 U7713 ( .A1(n7103), .A2(n7001), .ZN(n6157) );
  INV_X1 U7714 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n9391) );
  OR2_X1 U7715 ( .A1(n6157), .A2(n9391), .ZN(n6104) );
  INV_X1 U7716 ( .A(n6673), .ZN(n6106) );
  NAND2_X1 U7717 ( .A1(n6106), .A2(n4412), .ZN(n6110) );
  NOR2_X1 U7718 ( .A1(n6107), .A2(n6170), .ZN(n6108) );
  NAND2_X1 U7719 ( .A1(n6468), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n6114) );
  NAND2_X1 U7720 ( .A1(n6452), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n6113) );
  NAND2_X1 U7721 ( .A1(n6469), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n6112) );
  NAND2_X1 U7722 ( .A1(n6468), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n6117) );
  NAND2_X1 U7723 ( .A1(n6452), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n6116) );
  NAND2_X1 U7724 ( .A1(n6469), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n6115) );
  NAND3_X1 U7725 ( .A1(n6117), .A2(n6116), .A3(n6115), .ZN(n8830) );
  NOR2_X1 U7726 ( .A1(n8830), .A2(n8533), .ZN(n6478) );
  NAND2_X1 U7727 ( .A1(n6175), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n6124) );
  NAND2_X1 U7728 ( .A1(n6187), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n6123) );
  INV_X1 U7729 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n6121) );
  INV_X1 U7730 ( .A(n6700), .ZN(n7521) );
  NAND2_X1 U7731 ( .A1(n4545), .A2(SI_0_), .ZN(n6126) );
  INV_X1 U7732 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n6125) );
  NAND2_X1 U7733 ( .A1(n6126), .A2(n6125), .ZN(n6128) );
  AND2_X1 U7734 ( .A1(n6128), .A2(n6127), .ZN(n9400) );
  MUX2_X1 U7735 ( .A(P2_IR_REG_0__SCAN_IN), .B(n9400), .S(n7103), .Z(n10569)
         );
  INV_X1 U7736 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n6129) );
  OAI22_X1 U7737 ( .A1(n6157), .A2(n5620), .B1(n7103), .B2(n7272), .ZN(n6130)
         );
  INV_X1 U7738 ( .A(n6130), .ZN(n6133) );
  NAND2_X1 U7739 ( .A1(n4679), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n6135) );
  OR2_X1 U7740 ( .A1(n6136), .A2(n6135), .ZN(n6139) );
  NAND2_X1 U7741 ( .A1(n6199), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n6138) );
  NAND2_X1 U7742 ( .A1(n6187), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n6137) );
  INV_X1 U7743 ( .A(n7671), .ZN(n7571) );
  NAND2_X1 U7744 ( .A1(n8844), .A2(n7571), .ZN(n6908) );
  NAND2_X1 U7745 ( .A1(n6199), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n6144) );
  NAND2_X1 U7746 ( .A1(n6175), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n6143) );
  NAND2_X1 U7747 ( .A1(n6187), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n6142) );
  INV_X1 U7748 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n6140) );
  OR2_X1 U7749 ( .A1(n6145), .A2(n6170), .ZN(n6153) );
  INV_X1 U7750 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n6152) );
  XNOR2_X1 U7751 ( .A(n6153), .B(n6152), .ZN(n7120) );
  NAND2_X1 U7752 ( .A1(n7325), .A2(n8800), .ZN(n6511) );
  NAND2_X1 U7753 ( .A1(n4996), .A2(n6941), .ZN(n6513) );
  OAI21_X2 U7754 ( .B1(n7579), .B2(n7578), .A(n6511), .ZN(n7541) );
  INV_X1 U7755 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n6991) );
  NAND2_X1 U7756 ( .A1(n6199), .A2(n6991), .ZN(n6151) );
  NAND2_X1 U7757 ( .A1(n6175), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n6150) );
  NAND2_X1 U7758 ( .A1(n6187), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n6149) );
  INV_X1 U7759 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n6147) );
  NAND2_X1 U7760 ( .A1(n6153), .A2(n6152), .ZN(n6154) );
  NAND2_X1 U7761 ( .A1(n6154), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6156) );
  INV_X1 U7762 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n6155) );
  XNOR2_X1 U7763 ( .A(n6156), .B(n6155), .ZN(n7153) );
  NAND2_X1 U7764 ( .A1(n6995), .A2(n6192), .ZN(n6159) );
  INV_X2 U7765 ( .A(n6157), .ZN(n6196) );
  NAND2_X1 U7766 ( .A1(n6196), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n6158) );
  OAI211_X1 U7767 ( .C1(n7103), .C2(n7153), .A(n6159), .B(n6158), .ZN(n7546)
         );
  NAND2_X1 U7768 ( .A1(n7580), .A2(n7546), .ZN(n6507) );
  INV_X1 U7769 ( .A(n7580), .ZN(n8843) );
  INV_X1 U7770 ( .A(n7546), .ZN(n10524) );
  INV_X1 U7771 ( .A(n7540), .ZN(n6160) );
  NAND2_X1 U7772 ( .A1(n6411), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n6167) );
  INV_X1 U7773 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n6162) );
  NAND2_X1 U7774 ( .A1(n6991), .A2(n6162), .ZN(n6163) );
  NAND2_X1 U7775 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n6178) );
  AND2_X1 U7776 ( .A1(n6163), .A2(n6178), .ZN(n8760) );
  NAND2_X1 U7777 ( .A1(n6199), .A2(n8760), .ZN(n6165) );
  NAND2_X1 U7778 ( .A1(n6452), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n6164) );
  NAND2_X1 U7779 ( .A1(n6996), .A2(n6351), .ZN(n6174) );
  INV_X2 U7780 ( .A(n7103), .ZN(n7106) );
  NOR2_X1 U7781 ( .A1(n6168), .A2(n6170), .ZN(n6169) );
  MUX2_X1 U7782 ( .A(n6170), .B(n6169), .S(P2_IR_REG_4__SCAN_IN), .Z(n6172) );
  NOR2_X1 U7783 ( .A1(n6172), .A2(n6171), .ZN(n7128) );
  AOI22_X1 U7784 ( .A1(n6196), .A2(P1_DATAO_REG_4__SCAN_IN), .B1(n7106), .B2(
        n7128), .ZN(n6173) );
  NAND2_X1 U7785 ( .A1(n7715), .A2(n8759), .ZN(n6503) );
  INV_X1 U7786 ( .A(n7715), .ZN(n8842) );
  INV_X1 U7787 ( .A(n8759), .ZN(n7680) );
  NAND2_X1 U7788 ( .A1(n6411), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n6183) );
  NAND2_X1 U7789 ( .A1(n6175), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n6182) );
  INV_X1 U7790 ( .A(n6178), .ZN(n6176) );
  INV_X1 U7791 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n6177) );
  NAND2_X1 U7792 ( .A1(n6178), .A2(n6177), .ZN(n6179) );
  AND2_X1 U7793 ( .A1(n6204), .A2(n6179), .ZN(n8731) );
  NAND2_X1 U7794 ( .A1(n6199), .A2(n8731), .ZN(n6181) );
  NAND2_X1 U7795 ( .A1(n6187), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n6180) );
  NAND4_X1 U7796 ( .A1(n6183), .A2(n6182), .A3(n6181), .A4(n6180), .ZN(n8841)
         );
  NAND2_X1 U7797 ( .A1(n6998), .A2(n6351), .ZN(n6186) );
  OR2_X1 U7798 ( .A1(n6171), .A2(n6170), .ZN(n6184) );
  XNOR2_X1 U7799 ( .A(n6184), .B(P2_IR_REG_5__SCAN_IN), .ZN(n7135) );
  AOI22_X1 U7800 ( .A1(n6196), .A2(P1_DATAO_REG_5__SCAN_IN), .B1(n7106), .B2(
        n7135), .ZN(n6185) );
  INV_X1 U7801 ( .A(n8841), .ZN(n7781) );
  NAND2_X1 U7802 ( .A1(n7781), .A2(n6717), .ZN(n6637) );
  NAND2_X1 U7803 ( .A1(n6411), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n6191) );
  XNOR2_X1 U7804 ( .A(n6204), .B(P2_REG3_REG_6__SCAN_IN), .ZN(n7784) );
  NAND2_X1 U7805 ( .A1(n6199), .A2(n7784), .ZN(n6189) );
  NAND2_X1 U7806 ( .A1(n6187), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n6188) );
  NAND2_X1 U7807 ( .A1(n6997), .A2(n6192), .ZN(n6198) );
  NAND2_X1 U7808 ( .A1(n6171), .A2(n6193), .ZN(n6224) );
  NAND2_X1 U7809 ( .A1(n6224), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6194) );
  NAND2_X1 U7810 ( .A1(n6194), .A2(n6222), .ZN(n6210) );
  OR2_X1 U7811 ( .A1(n6194), .A2(n6222), .ZN(n6195) );
  AOI22_X1 U7812 ( .A1(n6196), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n7106), .B2(
        n7167), .ZN(n6197) );
  XNOR2_X1 U7813 ( .A(n8840), .B(n7783), .ZN(n7779) );
  INV_X1 U7814 ( .A(n7783), .ZN(n10579) );
  NOR2_X1 U7815 ( .A1(n8840), .A2(n10579), .ZN(n6510) );
  NAND2_X1 U7816 ( .A1(n6469), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n6209) );
  NAND2_X1 U7817 ( .A1(n6468), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n6208) );
  INV_X1 U7818 ( .A(n6204), .ZN(n6201) );
  NAND2_X1 U7819 ( .A1(n6201), .A2(n6200), .ZN(n6215) );
  INV_X1 U7820 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n6203) );
  INV_X1 U7821 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n6202) );
  OAI21_X1 U7822 ( .B1(n6204), .B2(n6203), .A(n6202), .ZN(n6205) );
  AND2_X1 U7823 ( .A1(n6215), .A2(n6205), .ZN(n7813) );
  NAND2_X1 U7824 ( .A1(n6437), .A2(n7813), .ZN(n6207) );
  NAND2_X1 U7825 ( .A1(n6452), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n6206) );
  AND4_X2 U7826 ( .A1(n6209), .A2(n6208), .A3(n6207), .A4(n6206), .ZN(n8690)
         );
  NAND2_X1 U7827 ( .A1(n6999), .A2(n6351), .ZN(n6213) );
  NAND2_X1 U7828 ( .A1(n6210), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6211) );
  XNOR2_X1 U7829 ( .A(n6211), .B(P2_IR_REG_7__SCAN_IN), .ZN(n7174) );
  AOI22_X1 U7830 ( .A1(n6196), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n7106), .B2(
        n7174), .ZN(n6212) );
  NAND2_X1 U7831 ( .A1(n6213), .A2(n6212), .ZN(n7824) );
  NAND2_X1 U7832 ( .A1(n8690), .A2(n7824), .ZN(n6528) );
  INV_X1 U7833 ( .A(n7824), .ZN(n6920) );
  INV_X1 U7834 ( .A(n8690), .ZN(n8839) );
  NAND2_X1 U7835 ( .A1(n6920), .A2(n8839), .ZN(n6527) );
  NAND2_X1 U7836 ( .A1(n6469), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n6220) );
  NAND2_X1 U7837 ( .A1(n6468), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n6219) );
  INV_X1 U7838 ( .A(n6215), .ZN(n6214) );
  NAND2_X1 U7839 ( .A1(n6214), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n6235) );
  INV_X1 U7840 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n9876) );
  NAND2_X1 U7841 ( .A1(n6215), .A2(n9876), .ZN(n6216) );
  AND2_X1 U7842 ( .A1(n6235), .A2(n6216), .ZN(n8693) );
  NAND2_X1 U7843 ( .A1(n6437), .A2(n8693), .ZN(n6218) );
  NAND2_X1 U7844 ( .A1(n6452), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n6217) );
  NAND4_X1 U7845 ( .A1(n6220), .A2(n6219), .A3(n6218), .A4(n6217), .ZN(n8838)
         );
  NAND2_X1 U7846 ( .A1(n7012), .A2(n6351), .ZN(n6227) );
  INV_X1 U7847 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n6221) );
  NAND2_X1 U7848 ( .A1(n6222), .A2(n6221), .ZN(n6223) );
  NAND2_X1 U7849 ( .A1(n6230), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6225) );
  XNOR2_X1 U7850 ( .A(n6225), .B(P2_IR_REG_8__SCAN_IN), .ZN(n7206) );
  AOI22_X1 U7851 ( .A1(n6196), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n7106), .B2(
        n7206), .ZN(n6226) );
  NAND2_X1 U7852 ( .A1(n6227), .A2(n6226), .ZN(n6944) );
  OR2_X1 U7853 ( .A1(n8838), .A2(n6944), .ZN(n6228) );
  NAND2_X1 U7854 ( .A1(n6944), .A2(n8838), .ZN(n8043) );
  INV_X1 U7855 ( .A(n8838), .ZN(n8046) );
  NAND2_X1 U7856 ( .A1(n6944), .A2(n8046), .ZN(n6530) );
  NAND2_X1 U7857 ( .A1(n7024), .A2(n6351), .ZN(n6232) );
  AOI22_X1 U7858 ( .A1(n6196), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n7106), .B2(
        n7299), .ZN(n6231) );
  NAND2_X1 U7859 ( .A1(n6411), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n6240) );
  NAND2_X1 U7860 ( .A1(n6468), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n6239) );
  INV_X1 U7861 ( .A(n6235), .ZN(n6233) );
  INV_X1 U7862 ( .A(n6248), .ZN(n6249) );
  INV_X1 U7863 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n6234) );
  NAND2_X1 U7864 ( .A1(n6235), .A2(n6234), .ZN(n6236) );
  AND2_X1 U7865 ( .A1(n6249), .A2(n6236), .ZN(n8053) );
  NAND2_X1 U7866 ( .A1(n6437), .A2(n8053), .ZN(n6238) );
  NAND2_X1 U7867 ( .A1(n6452), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n6237) );
  NAND4_X1 U7868 ( .A1(n6240), .A2(n6239), .A3(n6238), .A4(n6237), .ZN(n8837)
         );
  OR2_X1 U7869 ( .A1(n9355), .A2(n7988), .ZN(n6538) );
  NAND2_X1 U7870 ( .A1(n9355), .A2(n7988), .ZN(n8089) );
  INV_X1 U7871 ( .A(n8047), .ZN(n6241) );
  NAND2_X1 U7872 ( .A1(n7030), .A2(n6351), .ZN(n6247) );
  INV_X1 U7873 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n6268) );
  AOI21_X1 U7874 ( .B1(n6242), .B2(n6268), .A(n6170), .ZN(n6243) );
  NAND2_X1 U7875 ( .A1(n6243), .A2(P2_IR_REG_10__SCAN_IN), .ZN(n6245) );
  INV_X1 U7876 ( .A(n6243), .ZN(n6244) );
  NAND2_X1 U7877 ( .A1(n6244), .A2(n6269), .ZN(n6257) );
  AOI22_X1 U7878 ( .A1(n7335), .A2(n7106), .B1(n6196), .B2(
        P1_DATAO_REG_10__SCAN_IN), .ZN(n6246) );
  NAND2_X1 U7879 ( .A1(n6469), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n6254) );
  NAND2_X1 U7880 ( .A1(n6468), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n6253) );
  INV_X1 U7881 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n7294) );
  NAND2_X1 U7882 ( .A1(n6249), .A2(n7294), .ZN(n6250) );
  AND2_X1 U7883 ( .A1(n6261), .A2(n6250), .ZN(n8099) );
  NAND2_X1 U7884 ( .A1(n6437), .A2(n8099), .ZN(n6252) );
  NAND2_X1 U7885 ( .A1(n6452), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n6251) );
  OR2_X2 U7886 ( .A1(n8243), .A2(n8115), .ZN(n6537) );
  NAND2_X1 U7887 ( .A1(n8243), .A2(n8115), .ZN(n6540) );
  INV_X1 U7888 ( .A(n8109), .ZN(n6255) );
  NAND2_X1 U7889 ( .A1(n6257), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6258) );
  XNOR2_X1 U7890 ( .A(n6258), .B(P2_IR_REG_11__SCAN_IN), .ZN(n7478) );
  AOI22_X1 U7891 ( .A1(n7478), .A2(n7106), .B1(n6196), .B2(
        P1_DATAO_REG_11__SCAN_IN), .ZN(n6259) );
  NAND2_X1 U7892 ( .A1(n6411), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n6266) );
  NAND2_X1 U7893 ( .A1(n6468), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n6265) );
  NAND2_X1 U7894 ( .A1(n6261), .A2(n6260), .ZN(n6262) );
  AND2_X1 U7895 ( .A1(n6297), .A2(n6262), .ZN(n8121) );
  NAND2_X1 U7896 ( .A1(n6437), .A2(n8121), .ZN(n6264) );
  NAND2_X1 U7897 ( .A1(n6452), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n6263) );
  NAND2_X1 U7898 ( .A1(n9347), .A2(n8088), .ZN(n6639) );
  NAND2_X1 U7899 ( .A1(n7306), .A2(n6351), .ZN(n6275) );
  INV_X1 U7900 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n6267) );
  AND3_X1 U7901 ( .A1(n6269), .A2(n6268), .A3(n6267), .ZN(n6270) );
  INV_X1 U7902 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n6272) );
  NAND2_X1 U7903 ( .A1(n6292), .A2(n6272), .ZN(n6333) );
  NAND2_X1 U7904 ( .A1(n6333), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6282) );
  INV_X1 U7905 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n6330) );
  NAND2_X1 U7906 ( .A1(n6282), .A2(n6330), .ZN(n6273) );
  NAND2_X1 U7907 ( .A1(n6273), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6308) );
  XNOR2_X1 U7908 ( .A(n6308), .B(P2_IR_REG_14__SCAN_IN), .ZN(n8539) );
  AOI22_X1 U7909 ( .A1(n8539), .A2(n7106), .B1(n6464), .B2(
        P1_DATAO_REG_14__SCAN_IN), .ZN(n6274) );
  NAND2_X1 U7910 ( .A1(n6468), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n6281) );
  NAND2_X1 U7911 ( .A1(n6411), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n6280) );
  NAND2_X1 U7912 ( .A1(n6287), .A2(n9890), .ZN(n6277) );
  AND2_X1 U7913 ( .A1(n6340), .A2(n6277), .ZN(n9213) );
  NAND2_X1 U7914 ( .A1(n6437), .A2(n9213), .ZN(n6279) );
  NAND2_X1 U7915 ( .A1(n6452), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n6278) );
  NAND2_X1 U7916 ( .A1(n9331), .A2(n8914), .ZN(n6552) );
  NAND2_X1 U7917 ( .A1(n7273), .A2(n6351), .ZN(n6284) );
  XNOR2_X1 U7918 ( .A(n6282), .B(P2_IR_REG_13__SCAN_IN), .ZN(n7767) );
  AOI22_X1 U7919 ( .A1(n7767), .A2(n7106), .B1(n6464), .B2(
        P1_DATAO_REG_13__SCAN_IN), .ZN(n6283) );
  NAND2_X2 U7920 ( .A1(n6284), .A2(n6283), .ZN(n8911) );
  NAND2_X1 U7921 ( .A1(n6468), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n6291) );
  NAND2_X1 U7922 ( .A1(n6469), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n6290) );
  NAND2_X1 U7923 ( .A1(n6299), .A2(n6285), .ZN(n6286) );
  AND2_X1 U7924 ( .A1(n6287), .A2(n6286), .ZN(n8309) );
  NAND2_X1 U7925 ( .A1(n6437), .A2(n8309), .ZN(n6289) );
  NAND2_X1 U7926 ( .A1(n6452), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n6288) );
  NAND2_X1 U7927 ( .A1(n8911), .A2(n9204), .ZN(n9198) );
  NAND2_X1 U7928 ( .A1(n7076), .A2(n6351), .ZN(n6295) );
  OR2_X1 U7929 ( .A1(n6292), .A2(n6170), .ZN(n6293) );
  XNOR2_X1 U7930 ( .A(n6293), .B(P2_IR_REG_12__SCAN_IN), .ZN(n7646) );
  AOI22_X1 U7931 ( .A1(n7646), .A2(n7106), .B1(n6196), .B2(
        P1_DATAO_REG_12__SCAN_IN), .ZN(n6294) );
  NAND2_X1 U7932 ( .A1(n6469), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n6303) );
  NAND2_X1 U7933 ( .A1(n6468), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n6302) );
  INV_X1 U7934 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n6296) );
  NAND2_X1 U7935 ( .A1(n6297), .A2(n6296), .ZN(n6298) );
  AND2_X1 U7936 ( .A1(n6299), .A2(n6298), .ZN(n9227) );
  NAND2_X1 U7937 ( .A1(n6437), .A2(n9227), .ZN(n6301) );
  NAND2_X1 U7938 ( .A1(n6452), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n6300) );
  NAND2_X1 U7939 ( .A1(n9342), .A2(n8304), .ZN(n6632) );
  INV_X1 U7940 ( .A(n6548), .ZN(n6549) );
  OR2_X2 U7941 ( .A1(n9342), .A2(n8304), .ZN(n8298) );
  INV_X1 U7942 ( .A(n8298), .ZN(n6304) );
  OAI211_X1 U7943 ( .C1(n6549), .C2(n6304), .A(n6552), .B(n9198), .ZN(n6305)
         );
  OR2_X1 U7944 ( .A1(n9331), .A2(n8914), .ZN(n6551) );
  NAND2_X1 U7945 ( .A1(n7455), .A2(n6351), .ZN(n6312) );
  INV_X1 U7946 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n6331) );
  NAND2_X1 U7947 ( .A1(n6308), .A2(n6331), .ZN(n6309) );
  NAND2_X1 U7948 ( .A1(n6309), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6310) );
  XNOR2_X1 U7949 ( .A(n6310), .B(P2_IR_REG_15__SCAN_IN), .ZN(n8852) );
  AOI22_X1 U7950 ( .A1(n8852), .A2(n7106), .B1(n6464), .B2(
        P1_DATAO_REG_15__SCAN_IN), .ZN(n6311) );
  NAND2_X1 U7951 ( .A1(n6469), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n6316) );
  NAND2_X1 U7952 ( .A1(n6468), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n6315) );
  XNOR2_X1 U7953 ( .A(n6340), .B(P2_REG3_REG_15__SCAN_IN), .ZN(n8815) );
  NAND2_X1 U7954 ( .A1(n6437), .A2(n8815), .ZN(n6314) );
  NAND2_X1 U7955 ( .A1(n6452), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n6313) );
  NAND2_X1 U7956 ( .A1(n9327), .A2(n9206), .ZN(n6554) );
  NAND2_X1 U7957 ( .A1(n4487), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6318) );
  MUX2_X1 U7958 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6318), .S(
        P2_IR_REG_17__SCAN_IN), .Z(n6319) );
  AND2_X1 U7959 ( .A1(n6317), .A2(n6319), .ZN(n8543) );
  AOI22_X1 U7960 ( .A1(n6196), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n7106), .B2(
        n8543), .ZN(n6320) );
  NAND2_X2 U7961 ( .A1(n6321), .A2(n6320), .ZN(n9317) );
  INV_X1 U7962 ( .A(n6468), .ZN(n6435) );
  INV_X1 U7963 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n9918) );
  INV_X1 U7964 ( .A(n6452), .ZN(n6472) );
  INV_X1 U7965 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n6322) );
  OAI22_X1 U7966 ( .A1(n6435), .A2(n9918), .B1(n6472), .B2(n6322), .ZN(n6328)
         );
  AND2_X1 U7967 ( .A1(P2_REG3_REG_16__SCAN_IN), .A2(P2_REG3_REG_15__SCAN_IN), 
        .ZN(n6323) );
  INV_X1 U7968 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n9937) );
  NAND2_X1 U7969 ( .A1(n6342), .A2(n9937), .ZN(n6326) );
  NAND2_X1 U7970 ( .A1(n6365), .A2(n6326), .ZN(n9154) );
  INV_X1 U7971 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n9927) );
  OAI22_X1 U7972 ( .A1(n9154), .A2(n6467), .B1(n6455), .B2(n9927), .ZN(n6327)
         );
  INV_X1 U7973 ( .A(n9175), .ZN(n8721) );
  OR2_X2 U7974 ( .A1(n9317), .A2(n8721), .ZN(n6562) );
  NAND2_X1 U7975 ( .A1(n7458), .A2(n6351), .ZN(n6337) );
  NAND3_X1 U7976 ( .A1(n6331), .A2(n6330), .A3(n6329), .ZN(n6332) );
  OAI21_X1 U7977 ( .B1(n6333), .B2(n6332), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n6334) );
  MUX2_X1 U7978 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6334), .S(
        P2_IR_REG_16__SCAN_IN), .Z(n6335) );
  AND2_X1 U7979 ( .A1(n4487), .A2(n6335), .ZN(n8869) );
  AOI22_X1 U7980 ( .A1(n8869), .A2(n7106), .B1(n6464), .B2(
        P1_DATAO_REG_16__SCAN_IN), .ZN(n6336) );
  NAND2_X2 U7981 ( .A1(n6337), .A2(n6336), .ZN(n9321) );
  NAND2_X1 U7982 ( .A1(n6469), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n6346) );
  NAND2_X1 U7983 ( .A1(n6468), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n6345) );
  INV_X1 U7984 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n6339) );
  INV_X1 U7985 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n6338) );
  OAI21_X1 U7986 ( .B1(n6340), .B2(n6339), .A(n6338), .ZN(n6341) );
  AND2_X1 U7987 ( .A1(n6342), .A2(n6341), .ZN(n9166) );
  NAND2_X1 U7988 ( .A1(n6437), .A2(n9166), .ZN(n6344) );
  NAND2_X1 U7989 ( .A1(n6452), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n6343) );
  OR2_X1 U7990 ( .A1(n9321), .A2(n8833), .ZN(n6559) );
  NAND2_X1 U7991 ( .A1(n9317), .A2(n8721), .ZN(n6563) );
  NAND2_X1 U7992 ( .A1(n9321), .A2(n8833), .ZN(n6558) );
  NAND2_X1 U7993 ( .A1(n6563), .A2(n6558), .ZN(n6349) );
  NAND2_X1 U7994 ( .A1(n6349), .A2(n6562), .ZN(n6350) );
  NAND2_X1 U7995 ( .A1(n7655), .A2(n6351), .ZN(n6354) );
  NAND2_X1 U7996 ( .A1(n6317), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6352) );
  XNOR2_X1 U7997 ( .A(n6352), .B(P2_IR_REG_18__SCAN_IN), .ZN(n8547) );
  AOI22_X1 U7998 ( .A1(n6196), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n7106), .B2(
        n8547), .ZN(n6353) );
  NAND2_X2 U7999 ( .A1(n6354), .A2(n6353), .ZN(n9312) );
  INV_X1 U8000 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n9913) );
  NAND2_X1 U8001 ( .A1(n6468), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n6356) );
  NAND2_X1 U8002 ( .A1(n6452), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n6355) );
  OAI211_X1 U8003 ( .C1(n6455), .C2(n9913), .A(n6356), .B(n6355), .ZN(n6357)
         );
  INV_X1 U8004 ( .A(n6357), .ZN(n6359) );
  XNOR2_X1 U8005 ( .A(n6365), .B(P2_REG3_REG_18__SCAN_IN), .ZN(n9131) );
  NAND2_X1 U8006 ( .A1(n9131), .A2(n6437), .ZN(n6358) );
  NAND2_X1 U8007 ( .A1(n6359), .A2(n6358), .ZN(n9147) );
  INV_X1 U8008 ( .A(n9147), .ZN(n8917) );
  OR2_X1 U8009 ( .A1(n9312), .A2(n8917), .ZN(n6631) );
  NAND2_X1 U8010 ( .A1(n9134), .A2(n6631), .ZN(n6360) );
  NAND2_X1 U8011 ( .A1(n9312), .A2(n8917), .ZN(n6630) );
  NAND2_X1 U8012 ( .A1(n6360), .A2(n6630), .ZN(n9119) );
  NAND2_X1 U8013 ( .A1(n7705), .A2(n6351), .ZN(n6362) );
  XNOR2_X2 U8014 ( .A(n6493), .B(n6492), .ZN(n7706) );
  AOI22_X1 U8015 ( .A1(n6196), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n7106), .B2(
        n6625), .ZN(n6361) );
  INV_X1 U8016 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n6363) );
  OAI21_X1 U8017 ( .B1(n6365), .B2(n6363), .A(n9884), .ZN(n6366) );
  NAND2_X1 U8018 ( .A1(P2_REG3_REG_19__SCAN_IN), .A2(P2_REG3_REG_18__SCAN_IN), 
        .ZN(n6364) );
  AND2_X1 U8019 ( .A1(n6366), .A2(n6372), .ZN(n9115) );
  NAND2_X1 U8020 ( .A1(n9115), .A2(n6437), .ZN(n6369) );
  AOI22_X1 U8021 ( .A1(n6468), .A2(P2_REG1_REG_19__SCAN_IN), .B1(n6452), .B2(
        P2_REG2_REG_19__SCAN_IN), .ZN(n6368) );
  NAND2_X1 U8022 ( .A1(n6411), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n6367) );
  OR2_X1 U8023 ( .A1(n9307), .A2(n8918), .ZN(n6574) );
  NAND2_X1 U8024 ( .A1(n9307), .A2(n8918), .ZN(n6571) );
  NAND2_X1 U8025 ( .A1(n9119), .A2(n9120), .ZN(n9118) );
  NAND2_X1 U8026 ( .A1(n7774), .A2(n6351), .ZN(n6371) );
  OR2_X1 U8027 ( .A1(n6157), .A2(n9948), .ZN(n6370) );
  INV_X1 U8028 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n8771) );
  NAND2_X1 U8029 ( .A1(n6372), .A2(n8771), .ZN(n6373) );
  NAND2_X1 U8030 ( .A1(n6388), .A2(n6373), .ZN(n9100) );
  OR2_X1 U8031 ( .A1(n9100), .A2(n6467), .ZN(n6376) );
  AOI22_X1 U8032 ( .A1(n6468), .A2(P2_REG1_REG_20__SCAN_IN), .B1(n6469), .B2(
        P2_REG0_REG_20__SCAN_IN), .ZN(n6375) );
  NAND2_X1 U8033 ( .A1(n6452), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n6374) );
  OR2_X1 U8034 ( .A1(n9301), .A2(n9091), .ZN(n6576) );
  NAND2_X1 U8035 ( .A1(n9301), .A2(n9091), .ZN(n6577) );
  NAND2_X1 U8036 ( .A1(n6576), .A2(n6577), .ZN(n9098) );
  INV_X1 U8037 ( .A(n9098), .ZN(n9105) );
  NAND2_X1 U8038 ( .A1(n9104), .A2(n9105), .ZN(n9103) );
  NAND2_X1 U8039 ( .A1(n7929), .A2(n6351), .ZN(n6378) );
  NAND2_X1 U8040 ( .A1(n6464), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n6377) );
  XNOR2_X1 U8041 ( .A(n6388), .B(P2_REG3_REG_21__SCAN_IN), .ZN(n9084) );
  NAND2_X1 U8042 ( .A1(n9084), .A2(n6437), .ZN(n6384) );
  INV_X1 U8043 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n6381) );
  NAND2_X1 U8044 ( .A1(n6468), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n6380) );
  NAND2_X1 U8045 ( .A1(n6469), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n6379) );
  OAI211_X1 U8046 ( .C1(n6381), .C2(n6472), .A(n6380), .B(n6379), .ZN(n6382)
         );
  INV_X1 U8047 ( .A(n6382), .ZN(n6383) );
  OR2_X1 U8048 ( .A1(n9296), .A2(n9076), .ZN(n6580) );
  NAND2_X1 U8049 ( .A1(n9296), .A2(n9076), .ZN(n9072) );
  NAND2_X1 U8050 ( .A1(n7993), .A2(n6351), .ZN(n6386) );
  OR2_X1 U8051 ( .A1(n6157), .A2(n9862), .ZN(n6385) );
  INV_X1 U8052 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n9925) );
  INV_X1 U8053 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n8783) );
  OAI21_X1 U8054 ( .B1(n6388), .B2(n9925), .A(n8783), .ZN(n6389) );
  NAND2_X1 U8055 ( .A1(P2_REG3_REG_21__SCAN_IN), .A2(P2_REG3_REG_22__SCAN_IN), 
        .ZN(n6387) );
  AND2_X1 U8056 ( .A1(n6389), .A2(n6399), .ZN(n9069) );
  NAND2_X1 U8057 ( .A1(n9069), .A2(n6437), .ZN(n6394) );
  INV_X1 U8058 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n9794) );
  NAND2_X1 U8059 ( .A1(n6468), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n6391) );
  NAND2_X1 U8060 ( .A1(n6452), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n6390) );
  OAI211_X1 U8061 ( .C1(n6455), .C2(n9794), .A(n6391), .B(n6390), .ZN(n6392)
         );
  INV_X1 U8062 ( .A(n6392), .ZN(n6393) );
  NAND2_X1 U8063 ( .A1(n9291), .A2(n9092), .ZN(n6591) );
  NAND2_X1 U8064 ( .A1(n6406), .A2(n6591), .ZN(n9075) );
  INV_X1 U8065 ( .A(n9075), .ZN(n9065) );
  AND2_X1 U8066 ( .A1(n9065), .A2(n9072), .ZN(n6395) );
  NAND2_X1 U8067 ( .A1(n8127), .A2(n6351), .ZN(n6397) );
  NAND2_X1 U8068 ( .A1(n6464), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n6396) );
  INV_X1 U8069 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n8671) );
  NAND2_X1 U8070 ( .A1(n6399), .A2(n8671), .ZN(n6400) );
  NAND2_X1 U8071 ( .A1(n6409), .A2(n6400), .ZN(n9058) );
  OR2_X1 U8072 ( .A1(n9058), .A2(n6467), .ZN(n6405) );
  INV_X1 U8073 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n9059) );
  NAND2_X1 U8074 ( .A1(n6468), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n6402) );
  NAND2_X1 U8075 ( .A1(n6469), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n6401) );
  OAI211_X1 U8076 ( .C1(n9059), .C2(n6472), .A(n6402), .B(n6401), .ZN(n6403)
         );
  INV_X1 U8077 ( .A(n6403), .ZN(n6404) );
  OR2_X1 U8078 ( .A1(n9286), .A2(n9077), .ZN(n6593) );
  NAND2_X1 U8079 ( .A1(n9286), .A2(n9077), .ZN(n6583) );
  INV_X1 U8080 ( .A(n6406), .ZN(n9045) );
  NOR2_X1 U8081 ( .A1(n9044), .A2(n9045), .ZN(n6585) );
  NAND2_X1 U8082 ( .A1(n8254), .A2(n6351), .ZN(n6408) );
  NAND2_X1 U8083 ( .A1(n6464), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n6407) );
  INV_X1 U8084 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n8749) );
  NAND2_X1 U8085 ( .A1(n6409), .A2(n8749), .ZN(n6410) );
  NAND2_X1 U8086 ( .A1(n6420), .A2(n6410), .ZN(n9031) );
  INV_X1 U8087 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n9875) );
  NAND2_X1 U8088 ( .A1(n6452), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n6413) );
  NAND2_X1 U8089 ( .A1(n6411), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n6412) );
  OAI211_X1 U8090 ( .C1(n6435), .C2(n9875), .A(n6413), .B(n6412), .ZN(n6414)
         );
  INV_X1 U8091 ( .A(n6414), .ZN(n6415) );
  NAND2_X1 U8092 ( .A1(n9278), .A2(n9049), .ZN(n6417) );
  INV_X1 U8093 ( .A(n9049), .ZN(n8672) );
  OR2_X1 U8094 ( .A1(n9278), .A2(n8672), .ZN(n6587) );
  NAND2_X1 U8095 ( .A1(n6464), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n6418) );
  INV_X1 U8096 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n9966) );
  NAND2_X1 U8097 ( .A1(n6420), .A2(n9966), .ZN(n6421) );
  NAND2_X1 U8098 ( .A1(n6430), .A2(n6421), .ZN(n9021) );
  INV_X1 U8099 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n6424) );
  NAND2_X1 U8100 ( .A1(n6469), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n6423) );
  NAND2_X1 U8101 ( .A1(n6452), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n6422) );
  OAI211_X1 U8102 ( .C1(n6435), .C2(n6424), .A(n6423), .B(n6422), .ZN(n6425)
         );
  INV_X1 U8103 ( .A(n6425), .ZN(n6426) );
  NAND2_X1 U8104 ( .A1(n9275), .A2(n9036), .ZN(n6589) );
  NAND2_X1 U8105 ( .A1(n8416), .A2(n6351), .ZN(n6429) );
  NAND2_X1 U8106 ( .A1(n6464), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n6428) );
  INV_X1 U8107 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n6896) );
  NAND2_X1 U8108 ( .A1(n6430), .A2(n6896), .ZN(n6431) );
  INV_X1 U8109 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n6434) );
  NAND2_X1 U8110 ( .A1(n6469), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n6433) );
  NAND2_X1 U8111 ( .A1(n6452), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n6432) );
  OAI211_X1 U8112 ( .C1(n6435), .C2(n6434), .A(n6433), .B(n6432), .ZN(n6436)
         );
  AOI21_X1 U8113 ( .B1(n9008), .B2(n6437), .A(n6436), .ZN(n8991) );
  NAND2_X1 U8114 ( .A1(n9268), .A2(n8991), .ZN(n6629) );
  NAND2_X1 U8115 ( .A1(n8420), .A2(n6351), .ZN(n6439) );
  NAND2_X1 U8116 ( .A1(n6464), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n6438) );
  INV_X1 U8117 ( .A(n6442), .ZN(n6440) );
  NAND2_X1 U8118 ( .A1(n6440), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n6450) );
  INV_X1 U8119 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n6441) );
  NAND2_X1 U8120 ( .A1(n6442), .A2(n6441), .ZN(n6443) );
  NAND2_X1 U8121 ( .A1(n6450), .A2(n6443), .ZN(n8984) );
  INV_X1 U8122 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n9878) );
  NAND2_X1 U8123 ( .A1(n6468), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n6445) );
  NAND2_X1 U8124 ( .A1(n6452), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n6444) );
  OAI211_X1 U8125 ( .C1(n6455), .C2(n9878), .A(n6445), .B(n6444), .ZN(n6446)
         );
  INV_X1 U8126 ( .A(n6446), .ZN(n6447) );
  AND2_X1 U8127 ( .A1(n8962), .A2(n8960), .ZN(n6449) );
  INV_X1 U8128 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n6868) );
  NAND2_X1 U8129 ( .A1(n6450), .A2(n6868), .ZN(n6451) );
  INV_X1 U8130 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n9889) );
  NAND2_X1 U8131 ( .A1(n6468), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n6454) );
  NAND2_X1 U8132 ( .A1(n6452), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n6453) );
  OAI211_X1 U8133 ( .C1(n6455), .C2(n9889), .A(n6454), .B(n6453), .ZN(n6456)
         );
  INV_X1 U8134 ( .A(n6456), .ZN(n6457) );
  OR2_X1 U8135 ( .A1(n6604), .A2(n8941), .ZN(n6461) );
  INV_X1 U8136 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n9806) );
  OR2_X1 U8137 ( .A1(n6157), .A2(n9806), .ZN(n6603) );
  NAND2_X1 U8138 ( .A1(n9261), .A2(n8928), .ZN(n6607) );
  INV_X1 U8139 ( .A(n6603), .ZN(n6459) );
  NAND2_X1 U8140 ( .A1(n8992), .A2(n6459), .ZN(n6460) );
  AND4_X1 U8141 ( .A1(n6461), .A2(n6605), .A3(n6607), .A4(n6460), .ZN(n6462)
         );
  NAND2_X1 U8142 ( .A1(n8640), .A2(n6351), .ZN(n6466) );
  NAND2_X1 U8143 ( .A1(n6464), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n6465) );
  INV_X1 U8144 ( .A(P2_REG2_REG_29__SCAN_IN), .ZN(n8944) );
  NAND2_X1 U8145 ( .A1(n6468), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n6471) );
  NAND2_X1 U8146 ( .A1(n6469), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n6470) );
  OAI211_X1 U8147 ( .C1(n8944), .C2(n6472), .A(n6471), .B(n6470), .ZN(n6473)
         );
  INV_X1 U8148 ( .A(n6473), .ZN(n6474) );
  INV_X1 U8149 ( .A(n6612), .ZN(n6476) );
  NAND2_X1 U8150 ( .A1(n9245), .A2(n8969), .ZN(n6611) );
  INV_X1 U8151 ( .A(n6477), .ZN(n6480) );
  INV_X1 U8152 ( .A(n6478), .ZN(n6479) );
  AOI22_X1 U8153 ( .A1(n9241), .A2(n6481), .B1(n6480), .B2(n6479), .ZN(n6486)
         );
  NAND2_X1 U8154 ( .A1(n9384), .A2(n6351), .ZN(n6484) );
  OR2_X1 U8155 ( .A1(n6157), .A2(n6482), .ZN(n6483) );
  INV_X1 U8156 ( .A(n8830), .ZN(n6485) );
  OR2_X1 U8157 ( .A1(n8630), .A2(n6485), .ZN(n6622) );
  NAND2_X1 U8158 ( .A1(n8901), .A2(n8908), .ZN(n6613) );
  NAND2_X1 U8159 ( .A1(n6622), .A2(n6613), .ZN(n6627) );
  NAND2_X1 U8160 ( .A1(n8630), .A2(n6485), .ZN(n6621) );
  OAI21_X1 U8161 ( .B1(n6486), .B2(n6627), .A(n6621), .ZN(n6487) );
  XNOR2_X1 U8162 ( .A(n6487), .B(n6625), .ZN(n6498) );
  INV_X1 U8163 ( .A(n6488), .ZN(n6491) );
  NAND2_X1 U8164 ( .A1(n6491), .A2(n5093), .ZN(n6668) );
  NAND2_X1 U8165 ( .A1(n6493), .A2(n6492), .ZN(n6494) );
  INV_X1 U8166 ( .A(n4396), .ZN(n6848) );
  NAND2_X1 U8167 ( .A1(n6848), .A2(n6697), .ZN(n6928) );
  NAND2_X1 U8168 ( .A1(n6498), .A2(n6497), .ZN(n6660) );
  NAND2_X1 U8169 ( .A1(n6625), .A2(n6697), .ZN(n6499) );
  INV_X1 U8170 ( .A(n6511), .ZN(n6500) );
  NOR2_X1 U8171 ( .A1(n6500), .A2(n4394), .ZN(n6505) );
  INV_X1 U8172 ( .A(n10569), .ZN(n7570) );
  AND2_X1 U8173 ( .A1(n6700), .A2(n7570), .ZN(n6633) );
  NOR2_X1 U8174 ( .A1(n6633), .A2(n8533), .ZN(n6502) );
  OAI211_X1 U8175 ( .C1(n6501), .C2(n6502), .A(n6513), .B(n6908), .ZN(n6504)
         );
  NAND2_X1 U8176 ( .A1(n6637), .A2(n6503), .ZN(n6506) );
  INV_X1 U8177 ( .A(n6506), .ZN(n6508) );
  AOI22_X1 U8178 ( .A1(n6519), .A2(n6637), .B1(n6508), .B2(n6507), .ZN(n6509)
         );
  NAND2_X1 U8179 ( .A1(n8840), .A2(n10579), .ZN(n6520) );
  INV_X1 U8180 ( .A(n6908), .ZN(n6512) );
  OAI211_X1 U8181 ( .C1(n6512), .C2(n6633), .A(n6511), .B(n6907), .ZN(n6514)
         );
  NAND3_X1 U8182 ( .A1(n6514), .A2(n4394), .A3(n6513), .ZN(n6515) );
  OAI211_X1 U8183 ( .C1(n6516), .C2(n4397), .A(n6520), .B(n6515), .ZN(n6524)
         );
  AOI22_X1 U8184 ( .A1(n6519), .A2(n6636), .B1(n6518), .B2(n6517), .ZN(n6522)
         );
  INV_X1 U8185 ( .A(n6520), .ZN(n6521) );
  OAI21_X1 U8186 ( .B1(n6522), .B2(n6521), .A(n4394), .ZN(n6523) );
  OAI21_X1 U8187 ( .B1(n6525), .B2(n6524), .A(n6523), .ZN(n6526) );
  MUX2_X1 U8188 ( .A(n6528), .B(n6527), .S(n4394), .Z(n6529) );
  INV_X1 U8189 ( .A(n6944), .ZN(n10589) );
  NAND2_X1 U8190 ( .A1(n10589), .A2(n8838), .ZN(n6531) );
  MUX2_X1 U8191 ( .A(n6531), .B(n6530), .S(n4394), .Z(n6532) );
  NAND3_X1 U8192 ( .A1(n6533), .A2(n8089), .A3(n6532), .ZN(n6545) );
  AND2_X1 U8193 ( .A1(n8837), .A2(n4394), .ZN(n6535) );
  OAI21_X1 U8194 ( .B1(n4394), .B2(n8837), .A(n9355), .ZN(n6534) );
  OAI21_X1 U8195 ( .B1(n6535), .B2(n9355), .A(n6534), .ZN(n6536) );
  NAND3_X1 U8196 ( .A1(n6537), .A2(n6540), .A3(n6536), .ZN(n6539) );
  INV_X1 U8197 ( .A(n6539), .ZN(n6544) );
  OAI211_X1 U8198 ( .C1(n6539), .C2(n6538), .A(n6537), .B(n6640), .ZN(n6542)
         );
  NAND2_X1 U8199 ( .A1(n6639), .A2(n6540), .ZN(n6541) );
  MUX2_X1 U8200 ( .A(n6542), .B(n6541), .S(n4394), .Z(n6543) );
  NAND2_X1 U8201 ( .A1(n6632), .A2(n6639), .ZN(n6546) );
  NAND2_X1 U8202 ( .A1(n8298), .A2(n6640), .ZN(n6547) );
  MUX2_X1 U8203 ( .A(n6549), .B(n4667), .S(n4394), .Z(n6550) );
  NAND2_X1 U8204 ( .A1(n6551), .A2(n6552), .ZN(n9197) );
  MUX2_X1 U8205 ( .A(n6552), .B(n6551), .S(n4394), .Z(n6553) );
  NAND2_X1 U8206 ( .A1(n9184), .A2(n6553), .ZN(n6556) );
  NAND2_X1 U8207 ( .A1(n6559), .A2(n6558), .ZN(n9163) );
  INV_X1 U8208 ( .A(n9163), .ZN(n9173) );
  MUX2_X1 U8209 ( .A(n9142), .B(n6554), .S(n4394), .Z(n6555) );
  INV_X1 U8210 ( .A(n6558), .ZN(n9144) );
  INV_X1 U8211 ( .A(n6559), .ZN(n6560) );
  MUX2_X1 U8212 ( .A(n9144), .B(n6560), .S(n4394), .Z(n6561) );
  NAND2_X1 U8213 ( .A1(n6562), .A2(n6563), .ZN(n9150) );
  NOR2_X1 U8214 ( .A1(n6561), .A2(n9150), .ZN(n6567) );
  NAND2_X1 U8215 ( .A1(n6631), .A2(n6562), .ZN(n6565) );
  NAND2_X1 U8216 ( .A1(n6630), .A2(n6563), .ZN(n6564) );
  AOI21_X1 U8217 ( .B1(n6568), .B2(n6567), .A(n6566), .ZN(n6573) );
  INV_X1 U8218 ( .A(n6630), .ZN(n6569) );
  OAI21_X1 U8219 ( .B1(n6573), .B2(n6569), .A(n6574), .ZN(n6570) );
  INV_X1 U8220 ( .A(n6631), .ZN(n6572) );
  OAI21_X1 U8221 ( .B1(n6573), .B2(n6572), .A(n6571), .ZN(n6575) );
  NAND2_X1 U8222 ( .A1(n6580), .A2(n6576), .ZN(n6579) );
  NAND2_X1 U8223 ( .A1(n9072), .A2(n6577), .ZN(n6578) );
  MUX2_X1 U8224 ( .A(n6579), .B(n6578), .S(n4394), .Z(n6582) );
  MUX2_X1 U8225 ( .A(n9072), .B(n6580), .S(n4394), .Z(n6581) );
  INV_X1 U8226 ( .A(n6583), .ZN(n6584) );
  AOI21_X1 U8227 ( .B1(n6592), .B2(n6585), .A(n6584), .ZN(n6590) );
  NAND2_X1 U8228 ( .A1(n9278), .A2(n8672), .ZN(n6586) );
  MUX2_X1 U8229 ( .A(n6587), .B(n6586), .S(n4394), .Z(n6588) );
  NAND2_X1 U8230 ( .A1(n9016), .A2(n6588), .ZN(n6599) );
  OAI211_X1 U8231 ( .C1(n6590), .C2(n6599), .A(n6629), .B(n6589), .ZN(n6598)
         );
  OAI21_X1 U8232 ( .B1(n6596), .B2(n6599), .A(n6595), .ZN(n6597) );
  OAI21_X1 U8233 ( .B1(n6599), .B2(n9027), .A(n8960), .ZN(n6601) );
  MUX2_X1 U8234 ( .A(n8960), .B(n6629), .S(n4394), .Z(n6600) );
  INV_X1 U8235 ( .A(n8962), .ZN(n6602) );
  NAND2_X1 U8236 ( .A1(n9259), .A2(n8992), .ZN(n6606) );
  NAND2_X1 U8237 ( .A1(n6605), .A2(n6606), .ZN(n8963) );
  INV_X1 U8238 ( .A(n8963), .ZN(n8958) );
  INV_X1 U8239 ( .A(n6605), .ZN(n6608) );
  OAI21_X1 U8240 ( .B1(n6608), .B2(n6607), .A(n6606), .ZN(n6609) );
  MUX2_X1 U8241 ( .A(n6609), .B(n6608), .S(n4394), .Z(n6610) );
  MUX2_X1 U8242 ( .A(n6612), .B(n6611), .S(n4394), .Z(n6615) );
  INV_X1 U8243 ( .A(n6613), .ZN(n6614) );
  NOR2_X1 U8244 ( .A1(n8901), .A2(n8908), .ZN(n6617) );
  INV_X1 U8245 ( .A(n6617), .ZN(n6618) );
  MUX2_X1 U8246 ( .A(n6622), .B(n6621), .S(n4394), .Z(n6623) );
  INV_X2 U8247 ( .A(n7706), .ZN(n6625) );
  INV_X1 U8248 ( .A(n6929), .ZN(n6658) );
  INV_X1 U8249 ( .A(n6626), .ZN(n6652) );
  INV_X1 U8250 ( .A(n6627), .ZN(n6651) );
  INV_X1 U8251 ( .A(n6628), .ZN(n9242) );
  INV_X1 U8252 ( .A(n9087), .ZN(n6647) );
  INV_X1 U8253 ( .A(n9150), .ZN(n6645) );
  INV_X1 U8254 ( .A(n6501), .ZN(n6634) );
  INV_X1 U8255 ( .A(n6633), .ZN(n7697) );
  NAND4_X1 U8256 ( .A1(n6908), .A2(n6848), .A3(n6634), .A4(n7697), .ZN(n6635)
         );
  NOR4_X1 U8257 ( .A1(n6635), .A2(n7540), .A3(n7578), .A4(n7552), .ZN(n6638)
         );
  NAND4_X1 U8258 ( .A1(n6638), .A2(n7711), .A3(n7817), .A4(n7779), .ZN(n6641)
         );
  NOR4_X1 U8259 ( .A1(n6641), .A2(n8290), .A3(n6924), .A4(n8047), .ZN(n6642)
         );
  NAND4_X1 U8260 ( .A1(n8299), .A2(n9230), .A3(n6255), .A4(n6642), .ZN(n6643)
         );
  NOR4_X1 U8261 ( .A1(n9163), .A2(n5064), .A3(n9197), .A4(n6643), .ZN(n6644)
         );
  NAND4_X1 U8262 ( .A1(n9120), .A2(n9136), .A3(n6645), .A4(n6644), .ZN(n6646)
         );
  NOR4_X1 U8263 ( .A1(n9075), .A2(n6647), .A3(n9098), .A4(n6646), .ZN(n6648)
         );
  NAND4_X1 U8264 ( .A1(n9016), .A2(n9054), .A3(n6648), .A4(n9027), .ZN(n6649)
         );
  NOR4_X1 U8265 ( .A1(n8963), .A2(n8989), .A3(n9003), .A4(n6649), .ZN(n6650)
         );
  NAND4_X1 U8266 ( .A1(n6652), .A2(n6651), .A3(n9242), .A4(n6650), .ZN(n6653)
         );
  XNOR2_X1 U8267 ( .A(n6653), .B(n6625), .ZN(n6654) );
  NAND2_X1 U8268 ( .A1(n6654), .A2(n8533), .ZN(n6655) );
  NAND3_X1 U8269 ( .A1(n6660), .A2(n6656), .A3(n6655), .ZN(n6664) );
  NAND2_X1 U8270 ( .A1(n6660), .A2(n6659), .ZN(n6663) );
  OR2_X1 U8271 ( .A1(n6903), .A2(P2_U3152), .ZN(n7098) );
  INV_X1 U8272 ( .A(n7098), .ZN(n8128) );
  NAND3_X1 U8273 ( .A1(n6664), .A2(n6663), .A3(n8128), .ZN(n6687) );
  NAND3_X1 U8274 ( .A1(n6666), .A2(n6665), .A3(n6677), .ZN(n6667) );
  OAI21_X1 U8275 ( .B1(n6668), .B2(n6667), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n6669) );
  MUX2_X1 U8276 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6669), .S(
        P2_IR_REG_25__SCAN_IN), .Z(n6671) );
  NAND2_X1 U8277 ( .A1(n6671), .A2(n6670), .ZN(n8403) );
  INV_X1 U8278 ( .A(n8403), .ZN(n6675) );
  NAND2_X1 U8279 ( .A1(n6670), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6672) );
  MUX2_X1 U8280 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6672), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n6674) );
  NAND2_X1 U8281 ( .A1(n6674), .A2(n6673), .ZN(n8417) );
  NAND2_X1 U8282 ( .A1(n6675), .A2(n6832), .ZN(n6679) );
  OR2_X1 U8283 ( .A1(n6673), .A2(P2_IR_REG_27__SCAN_IN), .ZN(n6681) );
  NAND2_X1 U8284 ( .A1(n6681), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6682) );
  XNOR2_X1 U8285 ( .A(n6682), .B(P2_IR_REG_28__SCAN_IN), .ZN(n7121) );
  XNOR2_X1 U8286 ( .A(n6683), .B(P2_IR_REG_27__SCAN_IN), .ZN(n8635) );
  INV_X1 U8287 ( .A(n8635), .ZN(n9397) );
  NOR4_X1 U8288 ( .A1(n10530), .A2(n9203), .A3(n9397), .A4(n6863), .ZN(n6685)
         );
  OAI21_X1 U8289 ( .B1(n7098), .B2(n6624), .A(P2_B_REG_SCAN_IN), .ZN(n6684) );
  OR2_X1 U8290 ( .A1(n6685), .A2(n6684), .ZN(n6686) );
  NAND2_X1 U8291 ( .A1(n6687), .A2(n6686), .ZN(P2_U3244) );
  INV_X1 U8292 ( .A(n6688), .ZN(n6690) );
  INV_X1 U8293 ( .A(n7358), .ZN(n10278) );
  NOR2_X1 U8294 ( .A1(n10504), .A2(n6692), .ZN(n6693) );
  NOR2_X1 U8295 ( .A1(n5087), .A2(n6693), .ZN(n6694) );
  OAI21_X1 U8296 ( .B1(n6695), .B2(n10168), .A(n6694), .ZN(P1_U3552) );
  NAND3_X1 U8297 ( .A1(n6696), .A2(n8533), .A3(n6929), .ZN(n6699) );
  NAND2_X1 U8298 ( .A1(n4396), .A2(n6697), .ZN(n6939) );
  NAND2_X2 U8299 ( .A1(n6699), .A2(n6939), .ZN(n6705) );
  XNOR2_X1 U8300 ( .A(n6703), .B(n6702), .ZN(n7323) );
  NAND2_X1 U8301 ( .A1(n6909), .A2(n6812), .ZN(n7526) );
  NAND2_X1 U8302 ( .A1(n6754), .A2(n7570), .ZN(n6701) );
  AND2_X1 U8303 ( .A1(n7526), .A2(n6701), .ZN(n7324) );
  NAND2_X1 U8304 ( .A1(n7323), .A2(n7324), .ZN(n7322) );
  INV_X1 U8305 ( .A(n6703), .ZN(n8792) );
  NAND2_X1 U8306 ( .A1(n6702), .A2(n8792), .ZN(n6704) );
  NAND2_X1 U8307 ( .A1(n7322), .A2(n6704), .ZN(n6706) );
  NAND2_X1 U8308 ( .A1(n6706), .A2(n8794), .ZN(n8797) );
  INV_X1 U8309 ( .A(n6707), .ZN(n6708) );
  NAND2_X1 U8310 ( .A1(n6709), .A2(n6708), .ZN(n6710) );
  NAND2_X1 U8311 ( .A1(n8797), .A2(n6710), .ZN(n6989) );
  NOR2_X1 U8312 ( .A1(n7580), .A2(n4395), .ZN(n6720) );
  XNOR2_X1 U8313 ( .A(n6705), .B(n7546), .ZN(n8763) );
  INV_X1 U8314 ( .A(n6720), .ZN(n6712) );
  INV_X1 U8315 ( .A(n8763), .ZN(n6711) );
  NAND2_X1 U8316 ( .A1(n6712), .A2(n6711), .ZN(n6713) );
  NAND2_X1 U8317 ( .A1(n7600), .A2(n6713), .ZN(n6990) );
  XNOR2_X1 U8318 ( .A(n8759), .B(n6705), .ZN(n7598) );
  INV_X1 U8319 ( .A(n6715), .ZN(n7599) );
  XNOR2_X1 U8320 ( .A(n6717), .B(n6705), .ZN(n6724) );
  INV_X1 U8321 ( .A(n6724), .ZN(n7611) );
  AND2_X1 U8322 ( .A1(n8841), .A2(n6812), .ZN(n6723) );
  INV_X1 U8323 ( .A(n6723), .ZN(n6718) );
  NAND2_X1 U8324 ( .A1(n7600), .A2(n7599), .ZN(n6719) );
  NAND2_X1 U8325 ( .A1(n6719), .A2(n7598), .ZN(n6722) );
  NAND3_X1 U8326 ( .A1(n6715), .A2(n6720), .A3(n8763), .ZN(n6721) );
  NAND2_X1 U8327 ( .A1(n6722), .A2(n6721), .ZN(n6725) );
  XNOR2_X1 U8328 ( .A(n6754), .B(n7783), .ZN(n6728) );
  XNOR2_X1 U8329 ( .A(n6728), .B(n6727), .ZN(n7605) );
  NAND2_X1 U8330 ( .A1(n6728), .A2(n6727), .ZN(n6729) );
  INV_X1 U8331 ( .A(n7660), .ZN(n6735) );
  NOR2_X1 U8332 ( .A1(n8690), .A2(n7520), .ZN(n6730) );
  XNOR2_X1 U8333 ( .A(n7824), .B(n6821), .ZN(n6731) );
  NAND2_X1 U8334 ( .A1(n6730), .A2(n6731), .ZN(n6736) );
  INV_X1 U8335 ( .A(n6730), .ZN(n6732) );
  INV_X1 U8336 ( .A(n6731), .ZN(n8689) );
  NAND2_X1 U8337 ( .A1(n6732), .A2(n8689), .ZN(n6733) );
  NAND2_X1 U8338 ( .A1(n6736), .A2(n6733), .ZN(n7659) );
  NAND2_X1 U8339 ( .A1(n6735), .A2(n6734), .ZN(n7657) );
  NAND2_X1 U8340 ( .A1(n7657), .A2(n6736), .ZN(n6741) );
  XNOR2_X1 U8341 ( .A(n6944), .B(n6821), .ZN(n6737) );
  AND2_X1 U8342 ( .A1(n8838), .A2(n6812), .ZN(n6738) );
  NAND2_X1 U8343 ( .A1(n6737), .A2(n6738), .ZN(n6742) );
  INV_X1 U8344 ( .A(n6737), .ZN(n7747) );
  INV_X1 U8345 ( .A(n6738), .ZN(n6739) );
  NAND2_X1 U8346 ( .A1(n7747), .A2(n6739), .ZN(n6740) );
  AND2_X1 U8347 ( .A1(n6742), .A2(n6740), .ZN(n8687) );
  NAND2_X1 U8348 ( .A1(n6741), .A2(n8687), .ZN(n7746) );
  XNOR2_X1 U8349 ( .A(n9355), .B(n6821), .ZN(n6744) );
  NAND2_X1 U8350 ( .A1(n8837), .A2(n6812), .ZN(n6745) );
  XNOR2_X1 U8351 ( .A(n6744), .B(n6745), .ZN(n7757) );
  AND2_X1 U8352 ( .A1(n7757), .A2(n6742), .ZN(n6743) );
  INV_X1 U8353 ( .A(n6744), .ZN(n6746) );
  NAND2_X1 U8354 ( .A1(n6746), .A2(n6745), .ZN(n6747) );
  XNOR2_X1 U8355 ( .A(n4985), .B(n6821), .ZN(n6748) );
  NOR2_X1 U8356 ( .A1(n8115), .A2(n7520), .ZN(n6749) );
  NAND2_X1 U8357 ( .A1(n6748), .A2(n6749), .ZN(n6753) );
  INV_X1 U8358 ( .A(n6748), .ZN(n7934) );
  INV_X1 U8359 ( .A(n6749), .ZN(n6750) );
  NAND2_X1 U8360 ( .A1(n7934), .A2(n6750), .ZN(n6751) );
  NAND2_X1 U8361 ( .A1(n6753), .A2(n6751), .ZN(n7987) );
  INV_X1 U8362 ( .A(n7987), .ZN(n6752) );
  NAND2_X1 U8363 ( .A1(n7931), .A2(n6753), .ZN(n6755) );
  XNOR2_X1 U8364 ( .A(n9347), .B(n6829), .ZN(n6756) );
  NOR2_X1 U8365 ( .A1(n8088), .A2(n7520), .ZN(n6757) );
  XNOR2_X1 U8366 ( .A(n6756), .B(n6757), .ZN(n7932) );
  INV_X1 U8367 ( .A(n6756), .ZN(n6758) );
  NAND2_X1 U8368 ( .A1(n6758), .A2(n6757), .ZN(n6759) );
  XNOR2_X1 U8369 ( .A(n9342), .B(n6829), .ZN(n6760) );
  OR2_X1 U8370 ( .A1(n8304), .A2(n7520), .ZN(n6761) );
  NAND2_X1 U8371 ( .A1(n6760), .A2(n6761), .ZN(n8075) );
  INV_X1 U8372 ( .A(n6760), .ZN(n6763) );
  INV_X1 U8373 ( .A(n6761), .ZN(n6762) );
  NAND2_X1 U8374 ( .A1(n6763), .A2(n6762), .ZN(n8074) );
  XNOR2_X1 U8375 ( .A(n8911), .B(n6829), .ZN(n6764) );
  NOR2_X1 U8376 ( .A1(n9204), .A2(n7520), .ZN(n6765) );
  XNOR2_X1 U8377 ( .A(n6764), .B(n6765), .ZN(n8187) );
  NAND2_X1 U8378 ( .A1(n8186), .A2(n8187), .ZN(n6768) );
  INV_X1 U8379 ( .A(n6764), .ZN(n6766) );
  NAND2_X1 U8380 ( .A1(n6766), .A2(n6765), .ZN(n6767) );
  XNOR2_X1 U8381 ( .A(n9331), .B(n6829), .ZN(n6769) );
  OR2_X1 U8382 ( .A1(n8914), .A2(n4395), .ZN(n6770) );
  NAND2_X1 U8383 ( .A1(n6769), .A2(n6770), .ZN(n6775) );
  INV_X1 U8384 ( .A(n6769), .ZN(n6772) );
  INV_X1 U8385 ( .A(n6770), .ZN(n6771) );
  NAND2_X1 U8386 ( .A1(n6772), .A2(n6771), .ZN(n6773) );
  NAND2_X1 U8387 ( .A1(n6775), .A2(n6773), .ZN(n8657) );
  XNOR2_X1 U8388 ( .A(n9327), .B(n6829), .ZN(n8819) );
  NAND2_X1 U8389 ( .A1(n8820), .A2(n8819), .ZN(n6776) );
  NOR2_X1 U8390 ( .A1(n9206), .A2(n7520), .ZN(n8822) );
  NAND2_X1 U8391 ( .A1(n6776), .A2(n8822), .ZN(n6780) );
  INV_X1 U8392 ( .A(n8820), .ZN(n6778) );
  INV_X1 U8393 ( .A(n8819), .ZN(n6777) );
  NAND2_X1 U8394 ( .A1(n6778), .A2(n6777), .ZN(n6779) );
  XNOR2_X1 U8395 ( .A(n9321), .B(n6829), .ZN(n6781) );
  OR2_X1 U8396 ( .A1(n8833), .A2(n4395), .ZN(n6782) );
  NAND2_X1 U8397 ( .A1(n6781), .A2(n6782), .ZN(n6787) );
  INV_X1 U8398 ( .A(n6781), .ZN(n6784) );
  INV_X1 U8399 ( .A(n6782), .ZN(n6783) );
  NAND2_X1 U8400 ( .A1(n6784), .A2(n6783), .ZN(n6785) );
  NAND2_X1 U8401 ( .A1(n6787), .A2(n6785), .ZN(n8720) );
  XNOR2_X1 U8402 ( .A(n9317), .B(n6829), .ZN(n6789) );
  NAND2_X1 U8403 ( .A1(n9175), .A2(n6812), .ZN(n6788) );
  XNOR2_X1 U8404 ( .A(n6789), .B(n6788), .ZN(n8735) );
  XNOR2_X1 U8405 ( .A(n9312), .B(n6821), .ZN(n6792) );
  NAND2_X1 U8406 ( .A1(n9147), .A2(n6812), .ZN(n6790) );
  XNOR2_X1 U8407 ( .A(n6792), .B(n6790), .ZN(n8806) );
  NAND2_X1 U8408 ( .A1(n8805), .A2(n8806), .ZN(n6794) );
  INV_X1 U8409 ( .A(n6790), .ZN(n6791) );
  NAND2_X1 U8410 ( .A1(n6792), .A2(n6791), .ZN(n6793) );
  NAND2_X1 U8411 ( .A1(n6794), .A2(n6793), .ZN(n8678) );
  XNOR2_X1 U8412 ( .A(n9117), .B(n6821), .ZN(n6795) );
  OR2_X1 U8413 ( .A1(n8918), .A2(n7520), .ZN(n6796) );
  NAND2_X1 U8414 ( .A1(n6795), .A2(n6796), .ZN(n6800) );
  INV_X1 U8415 ( .A(n6795), .ZN(n6798) );
  INV_X1 U8416 ( .A(n6796), .ZN(n6797) );
  NAND2_X1 U8417 ( .A1(n6798), .A2(n6797), .ZN(n6799) );
  NAND2_X1 U8418 ( .A1(n6800), .A2(n6799), .ZN(n8681) );
  XNOR2_X1 U8419 ( .A(n9301), .B(n6829), .ZN(n6802) );
  INV_X1 U8420 ( .A(n9091), .ZN(n8921) );
  NAND2_X1 U8421 ( .A1(n8921), .A2(n6812), .ZN(n6801) );
  XNOR2_X1 U8422 ( .A(n6802), .B(n6801), .ZN(n8769) );
  XNOR2_X1 U8423 ( .A(n9086), .B(n6821), .ZN(n6805) );
  NOR2_X1 U8424 ( .A1(n9076), .A2(n7520), .ZN(n6807) );
  XNOR2_X1 U8425 ( .A(n6805), .B(n6807), .ZN(n8702) );
  NAND2_X1 U8426 ( .A1(n8701), .A2(n8702), .ZN(n8777) );
  XNOR2_X1 U8427 ( .A(n9291), .B(n6829), .ZN(n6804) );
  NAND2_X1 U8428 ( .A1(n9048), .A2(n6812), .ZN(n8781) );
  AND2_X1 U8429 ( .A1(n6804), .A2(n8781), .ZN(n6803) );
  OR2_X2 U8430 ( .A1(n8777), .A2(n6803), .ZN(n8665) );
  NOR2_X1 U8431 ( .A1(n9077), .A2(n4395), .ZN(n6814) );
  XNOR2_X1 U8432 ( .A(n9286), .B(n6821), .ZN(n6813) );
  INV_X1 U8433 ( .A(n6804), .ZN(n8778) );
  INV_X1 U8434 ( .A(n6805), .ZN(n6808) );
  NAND2_X1 U8435 ( .A1(n6808), .A2(n6807), .ZN(n8776) );
  NAND2_X1 U8436 ( .A1(n8776), .A2(n8781), .ZN(n6806) );
  NAND2_X1 U8437 ( .A1(n8778), .A2(n6806), .ZN(n6810) );
  NAND3_X1 U8438 ( .A1(n6808), .A2(n6807), .A3(n9048), .ZN(n6809) );
  NAND2_X1 U8439 ( .A1(n6810), .A2(n6809), .ZN(n8663) );
  AOI21_X1 U8440 ( .B1(n6814), .B2(n6813), .A(n8663), .ZN(n6811) );
  XNOR2_X1 U8441 ( .A(n9278), .B(n6829), .ZN(n8744) );
  NAND2_X1 U8442 ( .A1(n9049), .A2(n6812), .ZN(n8747) );
  INV_X1 U8443 ( .A(n6813), .ZN(n8666) );
  INV_X1 U8444 ( .A(n6814), .ZN(n8668) );
  AND2_X1 U8445 ( .A1(n8666), .A2(n8668), .ZN(n8741) );
  AOI21_X1 U8446 ( .B1(n8744), .B2(n8747), .A(n8741), .ZN(n6817) );
  INV_X1 U8447 ( .A(n8747), .ZN(n6816) );
  INV_X1 U8448 ( .A(n8744), .ZN(n6815) );
  INV_X1 U8449 ( .A(n9275), .ZN(n8935) );
  XNOR2_X1 U8450 ( .A(n8935), .B(n6821), .ZN(n6818) );
  NOR2_X1 U8451 ( .A1(n9036), .A2(n7520), .ZN(n8708) );
  INV_X1 U8452 ( .A(n6818), .ZN(n8709) );
  XNOR2_X1 U8453 ( .A(n9268), .B(n6821), .ZN(n8645) );
  NOR2_X1 U8454 ( .A1(n8991), .A2(n4395), .ZN(n6819) );
  NAND2_X1 U8455 ( .A1(n8645), .A2(n6819), .ZN(n6820) );
  OAI21_X1 U8456 ( .B1(n8645), .B2(n6819), .A(n6820), .ZN(n6892) );
  INV_X1 U8457 ( .A(n6820), .ZN(n6827) );
  XNOR2_X1 U8458 ( .A(n9261), .B(n6821), .ZN(n6822) );
  NOR2_X1 U8459 ( .A1(n8928), .A2(n7520), .ZN(n6823) );
  NAND2_X1 U8460 ( .A1(n6822), .A2(n6823), .ZN(n6828) );
  INV_X1 U8461 ( .A(n6822), .ZN(n6825) );
  INV_X1 U8462 ( .A(n6823), .ZN(n6824) );
  NAND2_X1 U8463 ( .A1(n6825), .A2(n6824), .ZN(n6826) );
  NAND2_X1 U8464 ( .A1(n8648), .A2(n6828), .ZN(n6859) );
  INV_X1 U8465 ( .A(n9259), .ZN(n6853) );
  NOR2_X1 U8466 ( .A1(n8992), .A2(n4395), .ZN(n6830) );
  XNOR2_X1 U8467 ( .A(n6830), .B(n6829), .ZN(n6857) );
  XNOR2_X1 U8468 ( .A(n8256), .B(P2_B_REG_SCAN_IN), .ZN(n6831) );
  NAND2_X1 U8469 ( .A1(n6831), .A2(n8403), .ZN(n6833) );
  INV_X1 U8470 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n6834) );
  NAND2_X1 U8471 ( .A1(n10531), .A2(n6834), .ZN(n6835) );
  NAND2_X1 U8472 ( .A1(n8256), .A2(n8417), .ZN(n10563) );
  INV_X1 U8473 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n6837) );
  NAND2_X1 U8474 ( .A1(n8403), .A2(n8417), .ZN(n10566) );
  INV_X1 U8475 ( .A(n10566), .ZN(n6836) );
  NOR4_X1 U8476 ( .A1(P2_D_REG_5__SCAN_IN), .A2(P2_D_REG_6__SCAN_IN), .A3(
        P2_D_REG_8__SCAN_IN), .A4(P2_D_REG_9__SCAN_IN), .ZN(n6846) );
  INV_X1 U8477 ( .A(P2_D_REG_10__SCAN_IN), .ZN(n10554) );
  INV_X1 U8478 ( .A(P2_D_REG_3__SCAN_IN), .ZN(n10561) );
  INV_X1 U8479 ( .A(P2_D_REG_4__SCAN_IN), .ZN(n10560) );
  INV_X1 U8480 ( .A(P2_D_REG_11__SCAN_IN), .ZN(n10553) );
  NAND4_X1 U8481 ( .A1(n10554), .A2(n10561), .A3(n10560), .A4(n10553), .ZN(
        n6843) );
  NOR4_X1 U8482 ( .A1(P2_D_REG_17__SCAN_IN), .A2(P2_D_REG_18__SCAN_IN), .A3(
        P2_D_REG_19__SCAN_IN), .A4(P2_D_REG_20__SCAN_IN), .ZN(n6841) );
  NOR4_X1 U8483 ( .A1(P2_D_REG_15__SCAN_IN), .A2(P2_D_REG_12__SCAN_IN), .A3(
        P2_D_REG_13__SCAN_IN), .A4(P2_D_REG_16__SCAN_IN), .ZN(n6840) );
  NOR4_X1 U8484 ( .A1(P2_D_REG_26__SCAN_IN), .A2(P2_D_REG_27__SCAN_IN), .A3(
        P2_D_REG_28__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n6839) );
  NOR4_X1 U8485 ( .A1(P2_D_REG_21__SCAN_IN), .A2(P2_D_REG_23__SCAN_IN), .A3(
        P2_D_REG_24__SCAN_IN), .A4(P2_D_REG_25__SCAN_IN), .ZN(n6838) );
  NAND4_X1 U8486 ( .A1(n6841), .A2(n6840), .A3(n6839), .A4(n6838), .ZN(n6842)
         );
  NOR4_X1 U8487 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        n6843), .A4(n6842), .ZN(n6845) );
  NOR4_X1 U8488 ( .A1(P2_D_REG_7__SCAN_IN), .A2(P2_D_REG_14__SCAN_IN), .A3(
        P2_D_REG_22__SCAN_IN), .A4(P2_D_REG_2__SCAN_IN), .ZN(n6844) );
  NAND3_X1 U8489 ( .A1(n6846), .A2(n6845), .A3(n6844), .ZN(n6847) );
  NAND2_X1 U8490 ( .A1(n10531), .A2(n6847), .ZN(n6937) );
  NAND3_X1 U8491 ( .A1(n7535), .A2(n7533), .A3(n6937), .ZN(n6862) );
  NAND2_X1 U8492 ( .A1(n6657), .A2(n6848), .ZN(n6943) );
  OR2_X1 U8493 ( .A1(n6860), .A2(n6943), .ZN(n6850) );
  INV_X1 U8494 ( .A(n10530), .ZN(n6849) );
  NOR3_X1 U8495 ( .A1(n6853), .A2(n6857), .A3(n8825), .ZN(n6851) );
  AOI21_X1 U8496 ( .B1(n6853), .B2(n6857), .A(n6851), .ZN(n6855) );
  AND2_X1 U8497 ( .A1(n6657), .A2(n6863), .ZN(n9287) );
  INV_X1 U8498 ( .A(n7102), .ZN(n7037) );
  NAND2_X1 U8499 ( .A1(n10588), .A2(n7037), .ZN(n6852) );
  OAI21_X1 U8500 ( .B1(n6853), .B2(n8695), .A(n8821), .ZN(n6854) );
  OAI21_X1 U8501 ( .B1(n6859), .B2(n6855), .A(n6854), .ZN(n6872) );
  NAND3_X1 U8502 ( .A1(n9259), .A2(n8695), .A3(n6857), .ZN(n6856) );
  OAI21_X1 U8503 ( .B1(n9259), .B2(n6857), .A(n6856), .ZN(n6858) );
  INV_X1 U8504 ( .A(n7121), .ZN(n7105) );
  OAI22_X1 U8505 ( .A1(n8969), .A2(n8785), .B1(n8928), .B2(n8786), .ZN(n6870)
         );
  INV_X1 U8506 ( .A(n7532), .ZN(n6861) );
  NAND2_X1 U8507 ( .A1(n6862), .A2(n6861), .ZN(n6867) );
  AND2_X1 U8508 ( .A1(n7102), .A2(n6863), .ZN(n6935) );
  INV_X1 U8509 ( .A(n6903), .ZN(n6864) );
  NOR2_X1 U8510 ( .A1(n6935), .A2(n6864), .ZN(n6865) );
  AND2_X1 U8511 ( .A1(n7099), .A2(n6865), .ZN(n6866) );
  NAND2_X1 U8512 ( .A1(n6867), .A2(n6866), .ZN(n7522) );
  OAI22_X1 U8513 ( .A1(n8970), .A2(n8818), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n6868), .ZN(n6869) );
  OAI21_X1 U8514 ( .B1(n6872), .B2(n6871), .A(n5084), .ZN(P2_U3222) );
  NAND2_X1 U8515 ( .A1(n9653), .A2(n6874), .ZN(n8626) );
  NAND3_X1 U8516 ( .A1(n6878), .A2(n10101), .A3(n6877), .ZN(n6881) );
  OAI22_X1 U8517 ( .A1(n9687), .A2(n10403), .B1(n8610), .B2(n10405), .ZN(n6879) );
  INV_X1 U8518 ( .A(n6879), .ZN(n6880) );
  NAND2_X1 U8519 ( .A1(n6881), .A2(n6880), .ZN(n8623) );
  OR2_X1 U8520 ( .A1(n6888), .A2(n9666), .ZN(n6882) );
  NAND2_X1 U8521 ( .A1(n8619), .A2(n6884), .ZN(n6885) );
  NAND2_X1 U8522 ( .A1(n6886), .A2(n6885), .ZN(P1_U3551) );
  INV_X1 U8523 ( .A(n10275), .ZN(n6889) );
  NAND2_X1 U8524 ( .A1(n6891), .A2(n6890), .ZN(P1_U3519) );
  NAND2_X1 U8525 ( .A1(n6893), .A2(n6892), .ZN(n6895) );
  NAND2_X1 U8526 ( .A1(n6895), .A2(n6894), .ZN(n6901) );
  INV_X1 U8527 ( .A(n9268), .ZN(n8929) );
  OAI22_X1 U8528 ( .A1(n8928), .A2(n9205), .B1(n9036), .B2(n9203), .ZN(n9267)
         );
  INV_X1 U8529 ( .A(n9267), .ZN(n9010) );
  OAI22_X1 U8530 ( .A1(n9010), .A2(n8712), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n6896), .ZN(n6897) );
  AOI21_X1 U8531 ( .B1(n9008), .B2(n8761), .A(n6897), .ZN(n6898) );
  OAI21_X1 U8532 ( .B1(n8929), .B2(n8695), .A(n6898), .ZN(n6899) );
  INV_X1 U8533 ( .A(n6899), .ZN(n6900) );
  OAI21_X1 U8534 ( .B1(n8644), .B2(n6901), .A(n6900), .ZN(P2_U3242) );
  NOR2_X1 U8535 ( .A1(n4520), .A2(n6902), .ZN(n6965) );
  NAND2_X1 U8536 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6903), .ZN(n10565) );
  NAND2_X1 U8537 ( .A1(n4520), .A2(n6904), .ZN(n6905) );
  NAND2_X1 U8538 ( .A1(n6905), .A2(n7497), .ZN(n6975) );
  NAND2_X1 U8539 ( .A1(n6975), .A2(n6966), .ZN(n6906) );
  NAND2_X1 U8540 ( .A1(n6906), .A2(P1_STATE_REG_SCAN_IN), .ZN(P1_U3083) );
  NAND2_X1 U8541 ( .A1(n6911), .A2(n7571), .ZN(n6912) );
  NAND2_X1 U8542 ( .A1(n7564), .A2(n6912), .ZN(n7577) );
  NAND2_X1 U8543 ( .A1(n7577), .A2(n7578), .ZN(n7576) );
  NAND2_X1 U8544 ( .A1(n7325), .A2(n6941), .ZN(n6913) );
  NAND2_X1 U8545 ( .A1(n7576), .A2(n6913), .ZN(n7536) );
  NAND2_X1 U8546 ( .A1(n7536), .A2(n7540), .ZN(n7538) );
  NAND2_X1 U8547 ( .A1(n7580), .A2(n10524), .ZN(n6914) );
  NAND2_X1 U8548 ( .A1(n7538), .A2(n6914), .ZN(n7551) );
  NAND2_X1 U8549 ( .A1(n7551), .A2(n7552), .ZN(n7550) );
  NAND2_X1 U8550 ( .A1(n7715), .A2(n7680), .ZN(n6915) );
  NOR2_X1 U8551 ( .A1(n8841), .A2(n6717), .ZN(n7775) );
  INV_X1 U8552 ( .A(n7775), .ZN(n6916) );
  NAND2_X1 U8553 ( .A1(n5101), .A2(n6916), .ZN(n6919) );
  AND2_X1 U8554 ( .A1(n5101), .A2(n6717), .ZN(n6917) );
  AOI22_X1 U8555 ( .A1(n7711), .A2(n6917), .B1(n8840), .B2(n7783), .ZN(n6918)
         );
  OAI21_X1 U8556 ( .B1(n6922), .B2(n6924), .A(n8112), .ZN(n10587) );
  XNOR2_X1 U8557 ( .A(n6624), .B(n6939), .ZN(n6923) );
  NAND2_X1 U8558 ( .A1(n6923), .A2(n7706), .ZN(n7666) );
  OR2_X1 U8559 ( .A1(n10587), .A2(n7666), .ZN(n6934) );
  NAND2_X1 U8560 ( .A1(n6925), .A2(n6924), .ZN(n6926) );
  NAND2_X1 U8561 ( .A1(n6927), .A2(n6926), .ZN(n6932) );
  NAND2_X1 U8562 ( .A1(n8837), .A2(n9222), .ZN(n6930) );
  OAI21_X1 U8563 ( .B1(n8690), .B2(n9203), .A(n6930), .ZN(n6931) );
  AOI21_X1 U8564 ( .B1(n6932), .B2(n9225), .A(n6931), .ZN(n6933) );
  NAND2_X1 U8565 ( .A1(n6934), .A2(n6933), .ZN(n10592) );
  NAND2_X1 U8566 ( .A1(n7533), .A2(n7561), .ZN(n6938) );
  NOR2_X1 U8567 ( .A1(n10530), .A2(n6935), .ZN(n6936) );
  NAND2_X1 U8568 ( .A1(n6937), .A2(n6936), .ZN(n7534) );
  MUX2_X1 U8569 ( .A(n10592), .B(P2_REG2_REG_8__SCAN_IN), .S(n4392), .Z(n6948)
         );
  OR2_X1 U8570 ( .A1(n6939), .A2(n7706), .ZN(n7665) );
  NOR2_X1 U8571 ( .A1(n4392), .A2(n7665), .ZN(n10519) );
  INV_X1 U8572 ( .A(n10519), .ZN(n8105) );
  NOR2_X1 U8573 ( .A1(n10587), .A2(n8105), .ZN(n6947) );
  NAND2_X1 U8574 ( .A1(n9158), .A2(n9357), .ZN(n8974) );
  NAND2_X1 U8575 ( .A1(n7812), .A2(n6944), .ZN(n6942) );
  NAND2_X1 U8576 ( .A1(n8052), .A2(n6942), .ZN(n10591) );
  AOI22_X1 U8577 ( .A1(n9190), .A2(n6944), .B1(n8693), .B2(n10517), .ZN(n6945)
         );
  OAI21_X1 U8578 ( .B1(n8974), .B2(n10591), .A(n6945), .ZN(n6946) );
  OR3_X1 U8579 ( .A1(n6948), .A2(n6947), .A3(n6946), .ZN(P2_U3288) );
  INV_X2 U8580 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3084) );
  OR2_X1 U8581 ( .A1(n6951), .A2(n6950), .ZN(n6952) );
  OR2_X1 U8582 ( .A1(n8599), .A2(n7798), .ZN(n6955) );
  INV_X1 U8583 ( .A(n4520), .ZN(n6957) );
  AOI22_X1 U8584 ( .A1(n6956), .A2(n7235), .B1(n6957), .B2(
        P1_IR_REG_0__SCAN_IN), .ZN(n6954) );
  NAND2_X1 U8585 ( .A1(n9590), .A2(n6956), .ZN(n6959) );
  NAND2_X1 U8586 ( .A1(n6957), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n6958) );
  OAI211_X1 U8587 ( .C1(n7865), .C2(n7794), .A(n6959), .B(n6958), .ZN(n7428)
         );
  NAND2_X1 U8588 ( .A1(n6960), .A2(n7428), .ZN(n7431) );
  OAI21_X1 U8589 ( .B1(n6960), .B2(n7428), .A(n7431), .ZN(n7372) );
  NOR2_X1 U8590 ( .A1(n10306), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n6961) );
  NOR2_X1 U8591 ( .A1(n10290), .A2(n6961), .ZN(n10308) );
  NAND3_X1 U8592 ( .A1(n7372), .A2(n10308), .A3(n10306), .ZN(n6964) );
  NAND2_X1 U8593 ( .A1(n10308), .A2(n6962), .ZN(n6963) );
  MUX2_X1 U8594 ( .A(n10308), .B(n6963), .S(n10307), .Z(n10312) );
  INV_X1 U8595 ( .A(P1_U4006), .ZN(n9576) );
  AOI21_X1 U8596 ( .B1(n6964), .B2(n10312), .A(n9576), .ZN(n7418) );
  NOR2_X1 U8597 ( .A1(n10399), .A2(n9917), .ZN(n6987) );
  INV_X1 U8598 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n6974) );
  AND2_X1 U8599 ( .A1(n6966), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6967) );
  AND2_X1 U8600 ( .A1(n6975), .A2(n6967), .ZN(n10314) );
  NAND2_X1 U8601 ( .A1(n6978), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n6969) );
  INV_X1 U8602 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n10493) );
  NAND2_X1 U8603 ( .A1(n10317), .A2(n10493), .ZN(n6968) );
  AND2_X1 U8604 ( .A1(n6969), .A2(n6968), .ZN(n10321) );
  AND2_X1 U8605 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(
        n10322) );
  NAND2_X1 U8606 ( .A1(n10321), .A2(n10322), .ZN(n10320) );
  NAND2_X1 U8607 ( .A1(n10320), .A2(n6969), .ZN(n7041) );
  INV_X1 U8608 ( .A(n7041), .ZN(n6971) );
  INV_X1 U8609 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n6970) );
  XNOR2_X1 U8610 ( .A(n7059), .B(n6970), .ZN(n7042) );
  XNOR2_X1 U8611 ( .A(n6971), .B(n7042), .ZN(n6972) );
  NAND2_X1 U8612 ( .A1(n10395), .A2(n6972), .ZN(n6973) );
  OAI21_X1 U8613 ( .B1(P1_STATE_REG_SCAN_IN), .B2(n6974), .A(n6973), .ZN(n6986) );
  NOR2_X1 U8614 ( .A1(n10306), .A2(P1_U3084), .ZN(n8421) );
  INV_X1 U8615 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n6976) );
  INV_X1 U8616 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n6977) );
  MUX2_X1 U8617 ( .A(n6977), .B(P1_REG2_REG_1__SCAN_IN), .S(n10317), .Z(n10324) );
  AND2_X1 U8618 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(
        n10325) );
  NAND2_X1 U8619 ( .A1(n10324), .A2(n10325), .ZN(n10323) );
  NAND2_X1 U8620 ( .A1(n6978), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n6980) );
  NAND2_X1 U8621 ( .A1(n10323), .A2(n6980), .ZN(n6979) );
  MUX2_X1 U8622 ( .A(n6976), .B(P1_REG2_REG_2__SCAN_IN), .S(n7059), .Z(n6981)
         );
  NAND3_X1 U8623 ( .A1(n6981), .A2(n10323), .A3(n6980), .ZN(n6982) );
  NAND3_X1 U8624 ( .A1(n10383), .A2(n7277), .A3(n6982), .ZN(n6984) );
  NAND2_X1 U8625 ( .A1(n10363), .A2(n7059), .ZN(n6983) );
  NAND2_X1 U8626 ( .A1(n6984), .A2(n6983), .ZN(n6985) );
  OR4_X1 U8627 ( .A1(n7418), .A2(n6987), .A3(n6986), .A4(n6985), .ZN(P1_U3243)
         );
  INV_X1 U8628 ( .A(n8756), .ZN(n6988) );
  AOI211_X1 U8629 ( .C1(n6990), .C2(n6989), .A(n8821), .B(n6988), .ZN(n6994)
         );
  MUX2_X1 U8630 ( .A(P2_U3152), .B(n8761), .S(n6991), .Z(n6993) );
  AOI22_X1 U8631 ( .A1(n9220), .A2(n4996), .B1(n8842), .B2(n9222), .ZN(n7542)
         );
  OAI22_X1 U8632 ( .A1(n8695), .A2(n10524), .B1(n7542), .B2(n8712), .ZN(n6992)
         );
  OR3_X1 U8633 ( .A1(n6994), .A2(n6993), .A3(n6992), .ZN(P2_U3220) );
  NOR2_X1 U8634 ( .A1(n4545), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9388) );
  INV_X2 U8635 ( .A(n9388), .ZN(n9395) );
  AND2_X1 U8636 ( .A1(n4545), .A2(P2_U3152), .ZN(n9392) );
  INV_X2 U8637 ( .A(n9392), .ZN(n9399) );
  OAI222_X1 U8638 ( .A1(n9395), .A2(n5113), .B1(n9399), .B2(n7004), .C1(
        P2_U3152), .C2(n7120), .ZN(P2_U3356) );
  INV_X1 U8639 ( .A(n6995), .ZN(n7010) );
  OAI222_X1 U8640 ( .A1(n9395), .A2(n5123), .B1(n9399), .B2(n7010), .C1(
        P2_U3152), .C2(n7153), .ZN(P2_U3355) );
  INV_X1 U8641 ( .A(n6996), .ZN(n7021) );
  INV_X1 U8642 ( .A(n7128), .ZN(n7137) );
  OAI222_X1 U8643 ( .A1(n9395), .A2(n5120), .B1(n9399), .B2(n7021), .C1(
        P2_U3152), .C2(n7137), .ZN(P2_U3354) );
  INV_X1 U8644 ( .A(n6997), .ZN(n7019) );
  INV_X1 U8645 ( .A(n7167), .ZN(n7177) );
  OAI222_X1 U8646 ( .A1(n9395), .A2(n5130), .B1(n9399), .B2(n7019), .C1(
        P2_U3152), .C2(n7177), .ZN(P2_U3352) );
  INV_X1 U8647 ( .A(n6998), .ZN(n7006) );
  INV_X1 U8648 ( .A(n7135), .ZN(n7162) );
  OAI222_X1 U8649 ( .A1(n9395), .A2(n5118), .B1(n9399), .B2(n7006), .C1(
        P2_U3152), .C2(n7162), .ZN(P2_U3353) );
  INV_X1 U8650 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n7000) );
  INV_X1 U8651 ( .A(n6999), .ZN(n7015) );
  INV_X1 U8652 ( .A(n7174), .ZN(n7209) );
  OAI222_X1 U8653 ( .A1(n9395), .A2(n7000), .B1(n9399), .B2(n7015), .C1(
        P2_U3152), .C2(n7209), .ZN(P2_U3351) );
  NAND2_X1 U8654 ( .A1(n7001), .A2(P1_U3084), .ZN(n10292) );
  CLKBUF_X1 U8655 ( .A(n10292), .Z(n10283) );
  INV_X1 U8656 ( .A(n10294), .ZN(n10281) );
  AOI22_X1 U8657 ( .A1(n7059), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_2__SCAN_IN), .B2(n10281), .ZN(n7003) );
  OAI21_X1 U8658 ( .B1(n7004), .B2(n10283), .A(n7003), .ZN(P1_U3351) );
  AOI22_X1 U8659 ( .A1(n9595), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_5__SCAN_IN), .B2(n10281), .ZN(n7005) );
  OAI21_X1 U8660 ( .B1(n7006), .B2(n10283), .A(n7005), .ZN(P1_U3348) );
  INV_X1 U8661 ( .A(n7356), .ZN(n7007) );
  NAND2_X1 U8662 ( .A1(n7007), .A2(n10428), .ZN(n7008) );
  OAI21_X1 U8663 ( .B1(n7009), .B2(n10428), .A(n7008), .ZN(P1_U3441) );
  INV_X1 U8664 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n7011) );
  INV_X1 U8665 ( .A(n7284), .ZN(n7282) );
  OAI222_X1 U8666 ( .A1(n10294), .A2(n7011), .B1(n10283), .B2(n7010), .C1(
        P1_U3084), .C2(n7282), .ZN(P1_U3350) );
  INV_X1 U8667 ( .A(n7012), .ZN(n7013) );
  INV_X1 U8668 ( .A(n7206), .ZN(n7298) );
  OAI222_X1 U8669 ( .A1(n9395), .A2(n9741), .B1(n9399), .B2(n7013), .C1(
        P2_U3152), .C2(n7298), .ZN(P2_U3350) );
  INV_X1 U8670 ( .A(n7082), .ZN(n7229) );
  OAI222_X1 U8671 ( .A1(n10294), .A2(n7014), .B1(n10283), .B2(n7013), .C1(
        P1_U3084), .C2(n7229), .ZN(P1_U3345) );
  INV_X1 U8672 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n7017) );
  INV_X1 U8673 ( .A(n7185), .ZN(n7016) );
  OAI222_X1 U8674 ( .A1(n7017), .A2(n10294), .B1(P1_U3084), .B2(n7016), .C1(
        n10283), .C2(n7015), .ZN(P1_U3346) );
  INV_X1 U8675 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n7020) );
  INV_X1 U8676 ( .A(n7087), .ZN(n7018) );
  OAI222_X1 U8677 ( .A1(n10294), .A2(n7020), .B1(n10283), .B2(n7019), .C1(
        P1_U3084), .C2(n7018), .ZN(P1_U3347) );
  INV_X1 U8678 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n7022) );
  INV_X1 U8679 ( .A(n7421), .ZN(n7410) );
  OAI222_X1 U8680 ( .A1(n10294), .A2(n7022), .B1(n10283), .B2(n7021), .C1(
        P1_U3084), .C2(n7410), .ZN(P1_U3349) );
  NAND2_X1 U8681 ( .A1(n8832), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n7023) );
  OAI21_X1 U8682 ( .B1(n8832), .B2(n8908), .A(n7023), .ZN(P2_U3582) );
  INV_X1 U8683 ( .A(n7024), .ZN(n7027) );
  INV_X1 U8684 ( .A(n7299), .ZN(n7310) );
  OAI222_X1 U8685 ( .A1(n9399), .A2(n7027), .B1(n7310), .B2(P2_U3152), .C1(
        n7025), .C2(n9395), .ZN(P2_U3349) );
  INV_X1 U8686 ( .A(n7254), .ZN(n7251) );
  OAI222_X1 U8687 ( .A1(P1_U3084), .A2(n7251), .B1(n10283), .B2(n7027), .C1(
        n7026), .C2(n10294), .ZN(P1_U3344) );
  INV_X1 U8688 ( .A(n7030), .ZN(n7032) );
  INV_X1 U8689 ( .A(n7335), .ZN(n7330) );
  OAI222_X1 U8690 ( .A1(n9399), .A2(n7032), .B1(n7330), .B2(P2_U3152), .C1(
        n7031), .C2(n9395), .ZN(P2_U3348) );
  INV_X1 U8691 ( .A(n7390), .ZN(n7252) );
  OAI222_X1 U8692 ( .A1(n10294), .A2(n9936), .B1(n10283), .B2(n7032), .C1(
        n7252), .C2(P1_U3084), .ZN(P1_U3343) );
  INV_X1 U8693 ( .A(n7033), .ZN(n7036) );
  INV_X1 U8694 ( .A(n7478), .ZN(n7339) );
  OAI222_X1 U8695 ( .A1(n9399), .A2(n7036), .B1(n7339), .B2(P2_U3152), .C1(
        n7034), .C2(n9395), .ZN(P2_U3347) );
  INV_X1 U8696 ( .A(n7393), .ZN(n7388) );
  OAI222_X1 U8697 ( .A1(P1_U3084), .A2(n7388), .B1(n10292), .B2(n7036), .C1(
        n7035), .C2(n10294), .ZN(P1_U3342) );
  OAI21_X1 U8698 ( .B1(n10530), .B2(n7037), .A(n7103), .ZN(n7039) );
  NAND2_X1 U8699 ( .A1(n10530), .A2(n7098), .ZN(n7038) );
  NAND2_X1 U8700 ( .A1(n7039), .A2(n7038), .ZN(n8863) );
  NOR2_X1 U8701 ( .A1(n10508), .A2(P2_U3966), .ZN(P2_U3151) );
  NAND2_X1 U8702 ( .A1(P1_U4006), .A2(n9641), .ZN(n7040) );
  OAI21_X1 U8703 ( .B1(P1_U4006), .B2(n6482), .A(n7040), .ZN(P1_U3586) );
  NAND2_X1 U8704 ( .A1(n7042), .A2(n7041), .ZN(n7044) );
  NAND2_X1 U8705 ( .A1(n7059), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n7043) );
  NAND2_X1 U8706 ( .A1(n7044), .A2(n7043), .ZN(n7283) );
  INV_X1 U8707 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n7045) );
  MUX2_X1 U8708 ( .A(P1_REG1_REG_3__SCAN_IN), .B(n7045), .S(n7284), .Z(n7046)
         );
  NAND2_X1 U8709 ( .A1(n7283), .A2(n7046), .ZN(n7285) );
  NAND2_X1 U8710 ( .A1(n7284), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n7047) );
  NAND2_X1 U8711 ( .A1(n7285), .A2(n7047), .ZN(n7405) );
  INV_X1 U8712 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n7404) );
  MUX2_X1 U8713 ( .A(n7404), .B(P1_REG1_REG_4__SCAN_IN), .S(n7421), .Z(n7048)
         );
  NAND2_X1 U8714 ( .A1(n7410), .A2(n7404), .ZN(n7049) );
  INV_X1 U8715 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n7050) );
  MUX2_X1 U8716 ( .A(P1_REG1_REG_5__SCAN_IN), .B(n7050), .S(n9595), .Z(n9597)
         );
  NAND2_X1 U8717 ( .A1(n9595), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n7051) );
  INV_X1 U8718 ( .A(n7053), .ZN(n7056) );
  INV_X1 U8719 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n10497) );
  MUX2_X1 U8720 ( .A(P1_REG1_REG_6__SCAN_IN), .B(n10497), .S(n7087), .Z(n7052)
         );
  INV_X1 U8721 ( .A(n7052), .ZN(n7055) );
  NAND2_X1 U8722 ( .A1(n7053), .A2(n7052), .ZN(n7191) );
  INV_X1 U8723 ( .A(n7191), .ZN(n7054) );
  AOI21_X1 U8724 ( .B1(n7056), .B2(n7055), .A(n7054), .ZN(n7075) );
  AND2_X1 U8725 ( .A1(P1_U3084), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n9530) );
  INV_X1 U8726 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n7057) );
  NOR2_X1 U8727 ( .A1(n10399), .A2(n7057), .ZN(n7058) );
  AOI211_X1 U8728 ( .C1(n10363), .C2(n7087), .A(n9530), .B(n7058), .ZN(n7074)
         );
  NAND2_X1 U8729 ( .A1(n7059), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n7276) );
  NAND2_X1 U8730 ( .A1(n7277), .A2(n7276), .ZN(n7061) );
  INV_X1 U8731 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n7978) );
  MUX2_X1 U8732 ( .A(P1_REG2_REG_3__SCAN_IN), .B(n7978), .S(n7284), .Z(n7060)
         );
  NAND2_X1 U8733 ( .A1(n7061), .A2(n7060), .ZN(n7280) );
  NAND2_X1 U8734 ( .A1(n7284), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n7062) );
  INV_X1 U8735 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n7411) );
  MUX2_X1 U8736 ( .A(n7411), .B(P1_REG2_REG_4__SCAN_IN), .S(n7421), .Z(n7063)
         );
  NAND2_X1 U8737 ( .A1(n7410), .A2(n7411), .ZN(n7064) );
  INV_X1 U8738 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n7065) );
  MUX2_X1 U8739 ( .A(P1_REG2_REG_5__SCAN_IN), .B(n7065), .S(n9595), .Z(n7066)
         );
  NAND2_X1 U8740 ( .A1(n9595), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n7071) );
  NAND2_X1 U8741 ( .A1(n9591), .A2(n7071), .ZN(n7069) );
  INV_X1 U8742 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n7067) );
  MUX2_X1 U8743 ( .A(P1_REG2_REG_6__SCAN_IN), .B(n7067), .S(n7087), .Z(n7068)
         );
  NAND2_X1 U8744 ( .A1(n7069), .A2(n7068), .ZN(n7089) );
  MUX2_X1 U8745 ( .A(n7067), .B(P1_REG2_REG_6__SCAN_IN), .S(n7087), .Z(n7070)
         );
  NAND3_X1 U8746 ( .A1(n9591), .A2(n7071), .A3(n7070), .ZN(n7072) );
  NAND3_X1 U8747 ( .A1(n10383), .A2(n7089), .A3(n7072), .ZN(n7073) );
  OAI211_X1 U8748 ( .C1(n7075), .C2(n7629), .A(n7074), .B(n7073), .ZN(P1_U3247) );
  INV_X1 U8749 ( .A(n7076), .ZN(n7078) );
  INV_X1 U8750 ( .A(n7646), .ZN(n7638) );
  OAI222_X1 U8751 ( .A1(n9395), .A2(n7077), .B1(n9399), .B2(n7078), .C1(
        P2_U3152), .C2(n7638), .ZN(P2_U3346) );
  OAI222_X1 U8752 ( .A1(n10294), .A2(n7079), .B1(n10283), .B2(n7078), .C1(
        P1_U3084), .C2(n7460), .ZN(P1_U3341) );
  INV_X1 U8753 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n10502) );
  MUX2_X1 U8754 ( .A(n10502), .B(P1_REG1_REG_9__SCAN_IN), .S(n7254), .Z(n7085)
         );
  OR2_X1 U8755 ( .A1(n7087), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n7189) );
  NAND2_X1 U8756 ( .A1(n7191), .A2(n7189), .ZN(n7080) );
  INV_X1 U8757 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n10499) );
  MUX2_X1 U8758 ( .A(P1_REG1_REG_7__SCAN_IN), .B(n10499), .S(n7185), .Z(n7188)
         );
  NAND2_X1 U8759 ( .A1(n7080), .A2(n7188), .ZN(n7193) );
  OR2_X1 U8760 ( .A1(n7185), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n7081) );
  NAND2_X1 U8761 ( .A1(n7082), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n7084) );
  NOR2_X1 U8762 ( .A1(n7082), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n7083) );
  AOI21_X1 U8763 ( .B1(n7085), .B2(n7219), .A(n7250), .ZN(n7097) );
  NAND2_X1 U8764 ( .A1(P1_U3084), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n8159) );
  OAI21_X1 U8765 ( .B1(n10390), .B2(n7251), .A(n8159), .ZN(n7086) );
  AOI21_X1 U8766 ( .B1(n10319), .B2(P1_ADDR_REG_9__SCAN_IN), .A(n7086), .ZN(
        n7096) );
  NAND2_X1 U8767 ( .A1(n7087), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n7088) );
  INV_X1 U8768 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n9859) );
  MUX2_X1 U8769 ( .A(P1_REG2_REG_7__SCAN_IN), .B(n9859), .S(n7185), .Z(n7183)
         );
  OR2_X1 U8770 ( .A1(n7185), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n7090) );
  NAND2_X1 U8771 ( .A1(n7215), .A2(n7229), .ZN(n7092) );
  INV_X1 U8772 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n7969) );
  NAND2_X1 U8773 ( .A1(n7091), .A2(n7969), .ZN(n7225) );
  INV_X1 U8774 ( .A(n7226), .ZN(n7216) );
  XNOR2_X1 U8775 ( .A(n7254), .B(P1_REG2_REG_9__SCAN_IN), .ZN(n7093) );
  INV_X1 U8776 ( .A(n7093), .ZN(n7094) );
  OAI211_X1 U8777 ( .C1(n7216), .C2(n7094), .A(n10383), .B(n7256), .ZN(n7095)
         );
  OAI211_X1 U8778 ( .C1(n7097), .C2(n7629), .A(n7096), .B(n7095), .ZN(P1_U3250) );
  NAND2_X1 U8779 ( .A1(n7121), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9393) );
  OAI21_X1 U8780 ( .B1(n7099), .B2(n9393), .A(n7098), .ZN(n7100) );
  INV_X1 U8781 ( .A(n7100), .ZN(n7101) );
  OAI21_X1 U8782 ( .B1(n10530), .B2(n7102), .A(n7101), .ZN(n7108) );
  NAND2_X1 U8783 ( .A1(n7108), .A2(n7103), .ZN(n7104) );
  NAND2_X1 U8784 ( .A1(n7104), .A2(n8832), .ZN(n7123) );
  INV_X1 U8785 ( .A(n8870), .ZN(n10509) );
  AND2_X1 U8786 ( .A1(P2_U3152), .A2(P2_REG3_REG_4__SCAN_IN), .ZN(n7119) );
  NOR2_X1 U8787 ( .A1(n7106), .A2(n8635), .ZN(n7107) );
  INV_X1 U8788 ( .A(n7272), .ZN(n7110) );
  INV_X1 U8789 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n7575) );
  INV_X1 U8790 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n7262) );
  INV_X1 U8791 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n7109) );
  AOI21_X1 U8792 ( .B1(n7110), .B2(P2_REG1_REG_1__SCAN_IN), .A(n7263), .ZN(
        n7242) );
  INV_X1 U8793 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n7588) );
  MUX2_X1 U8794 ( .A(P2_REG1_REG_2__SCAN_IN), .B(n7588), .S(n7120), .Z(n7241)
         );
  OR2_X1 U8795 ( .A1(n7242), .A2(n7241), .ZN(n7239) );
  NAND2_X1 U8796 ( .A1(n4515), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n7143) );
  INV_X1 U8797 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n7591) );
  MUX2_X1 U8798 ( .A(P2_REG1_REG_3__SCAN_IN), .B(n7591), .S(n7153), .Z(n7142)
         );
  NOR2_X1 U8799 ( .A1(n7153), .A2(n7591), .ZN(n7113) );
  INV_X1 U8800 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n7111) );
  MUX2_X1 U8801 ( .A(P2_REG1_REG_4__SCAN_IN), .B(n7111), .S(n7128), .Z(n7112)
         );
  INV_X1 U8802 ( .A(n7145), .ZN(n7116) );
  INV_X1 U8803 ( .A(n7113), .ZN(n7115) );
  MUX2_X1 U8804 ( .A(n7111), .B(P2_REG1_REG_4__SCAN_IN), .S(n7128), .Z(n7114)
         );
  NAND3_X1 U8805 ( .A1(n7116), .A2(n7115), .A3(n7114), .ZN(n7117) );
  AND3_X1 U8806 ( .A1(n10505), .A2(n7131), .A3(n7117), .ZN(n7118) );
  AOI211_X1 U8807 ( .C1(n10508), .C2(P2_ADDR_REG_4__SCAN_IN), .A(n7119), .B(
        n7118), .ZN(n7127) );
  INV_X1 U8808 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n7679) );
  MUX2_X1 U8809 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n7679), .S(n7128), .Z(n7125)
         );
  INV_X1 U8810 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n7672) );
  AND2_X1 U8811 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(
        n7268) );
  OAI21_X1 U8812 ( .B1(n7272), .B2(n7672), .A(n7267), .ZN(n7246) );
  XNOR2_X1 U8813 ( .A(n7120), .B(P2_REG2_REG_2__SCAN_IN), .ZN(n7247) );
  NAND2_X1 U8814 ( .A1(n7246), .A2(n7247), .ZN(n7245) );
  XNOR2_X1 U8815 ( .A(n7153), .B(P2_REG2_REG_3__SCAN_IN), .ZN(n7150) );
  AND2_X1 U8816 ( .A1(n7121), .A2(n8635), .ZN(n7122) );
  NAND2_X1 U8817 ( .A1(n7123), .A2(n7122), .ZN(n10511) );
  OAI211_X1 U8818 ( .C1(n7125), .C2(n7124), .A(n10506), .B(n7136), .ZN(n7126)
         );
  OAI211_X1 U8819 ( .C1(n10509), .C2(n7137), .A(n7127), .B(n7126), .ZN(
        P2_U3249) );
  AND2_X1 U8820 ( .A1(P2_U3152), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n7134) );
  NAND2_X1 U8821 ( .A1(n7128), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n7130) );
  INV_X1 U8822 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n10600) );
  MUX2_X1 U8823 ( .A(n10600), .B(P2_REG1_REG_5__SCAN_IN), .S(n7135), .Z(n7129)
         );
  AND3_X1 U8824 ( .A1(n7131), .A2(n7130), .A3(n7129), .ZN(n7132) );
  NOR3_X1 U8825 ( .A1(n10510), .A2(n7157), .A3(n7132), .ZN(n7133) );
  AOI211_X1 U8826 ( .C1(n10508), .C2(P2_ADDR_REG_5__SCAN_IN), .A(n7134), .B(
        n7133), .ZN(n7141) );
  INV_X1 U8827 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n9825) );
  MUX2_X1 U8828 ( .A(P2_REG2_REG_5__SCAN_IN), .B(n9825), .S(n7135), .Z(n7139)
         );
  OAI211_X1 U8829 ( .C1(n7139), .C2(n7138), .A(n10506), .B(n7161), .ZN(n7140)
         );
  OAI211_X1 U8830 ( .C1(n10509), .C2(n7162), .A(n7141), .B(n7140), .ZN(
        P2_U3250) );
  NOR2_X1 U8831 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6991), .ZN(n7147) );
  AND3_X1 U8832 ( .A1(n7239), .A2(n7143), .A3(n7142), .ZN(n7144) );
  NOR3_X1 U8833 ( .A1(n10510), .A2(n7145), .A3(n7144), .ZN(n7146) );
  AOI211_X1 U8834 ( .C1(n10508), .C2(P2_ADDR_REG_3__SCAN_IN), .A(n7147), .B(
        n7146), .ZN(n7152) );
  OAI211_X1 U8835 ( .C1(n7150), .C2(n7149), .A(n10506), .B(n7148), .ZN(n7151)
         );
  OAI211_X1 U8836 ( .C1(n10509), .C2(n7153), .A(n7152), .B(n7151), .ZN(
        P2_U3248) );
  AND2_X1 U8837 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_U3152), .ZN(n7609) );
  NOR2_X1 U8838 ( .A1(n7162), .A2(n10600), .ZN(n7156) );
  INV_X1 U8839 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n7154) );
  MUX2_X1 U8840 ( .A(P2_REG1_REG_6__SCAN_IN), .B(n7154), .S(n7167), .Z(n7155)
         );
  INV_X1 U8841 ( .A(n7170), .ZN(n7159) );
  NOR3_X1 U8842 ( .A1(n7157), .A2(n7156), .A3(n7155), .ZN(n7158) );
  NOR3_X1 U8843 ( .A1(n10510), .A2(n7159), .A3(n7158), .ZN(n7160) );
  AOI211_X1 U8844 ( .C1(n10508), .C2(P2_ADDR_REG_6__SCAN_IN), .A(n7609), .B(
        n7160), .ZN(n7166) );
  XOR2_X1 U8845 ( .A(P2_REG2_REG_6__SCAN_IN), .B(n7167), .Z(n7164) );
  OAI21_X1 U8846 ( .B1(n9825), .B2(n7162), .A(n7161), .ZN(n7163) );
  OAI211_X1 U8847 ( .C1(n7164), .C2(n7163), .A(n10506), .B(n7175), .ZN(n7165)
         );
  OAI211_X1 U8848 ( .C1(n10509), .C2(n7177), .A(n7166), .B(n7165), .ZN(
        P2_U3251) );
  AND2_X1 U8849 ( .A1(P2_U3152), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n7173) );
  NAND2_X1 U8850 ( .A1(n7167), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n7169) );
  INV_X1 U8851 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n7830) );
  MUX2_X1 U8852 ( .A(n7830), .B(P2_REG1_REG_7__SCAN_IN), .S(n7174), .Z(n7168)
         );
  AOI21_X1 U8853 ( .B1(n7170), .B2(n7169), .A(n7168), .ZN(n7201) );
  AND3_X1 U8854 ( .A1(n7170), .A2(n7169), .A3(n7168), .ZN(n7171) );
  NOR3_X1 U8855 ( .A1(n10510), .A2(n7201), .A3(n7171), .ZN(n7172) );
  AOI211_X1 U8856 ( .C1(n10508), .C2(P2_ADDR_REG_7__SCAN_IN), .A(n7173), .B(
        n7172), .ZN(n7181) );
  XOR2_X1 U8857 ( .A(P2_REG2_REG_7__SCAN_IN), .B(n7174), .Z(n7179) );
  INV_X1 U8858 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n7176) );
  OAI21_X1 U8859 ( .B1(n7177), .B2(n7176), .A(n7175), .ZN(n7178) );
  NAND2_X1 U8860 ( .A1(n7178), .A2(n7179), .ZN(n7207) );
  OAI211_X1 U8861 ( .C1(n7179), .C2(n7178), .A(n10506), .B(n7207), .ZN(n7180)
         );
  OAI211_X1 U8862 ( .C1(n10509), .C2(n7209), .A(n7181), .B(n7180), .ZN(
        P2_U3252) );
  OAI21_X1 U8863 ( .B1(n7184), .B2(n7183), .A(n7182), .ZN(n7196) );
  INV_X1 U8864 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n7187) );
  NOR2_X1 U8865 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n5632), .ZN(n7878) );
  AOI21_X1 U8866 ( .B1(n10363), .B2(n7185), .A(n7878), .ZN(n7186) );
  OAI21_X1 U8867 ( .B1(n10399), .B2(n7187), .A(n7186), .ZN(n7195) );
  INV_X1 U8868 ( .A(n7188), .ZN(n7190) );
  NAND3_X1 U8869 ( .A1(n7191), .A2(n7190), .A3(n7189), .ZN(n7192) );
  AOI21_X1 U8870 ( .B1(n7193), .B2(n7192), .A(n7629), .ZN(n7194) );
  AOI211_X1 U8871 ( .C1(n10383), .C2(n7196), .A(n7195), .B(n7194), .ZN(n7197)
         );
  INV_X1 U8872 ( .A(n7197), .ZN(P1_U3248) );
  NOR2_X1 U8873 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9876), .ZN(n7205) );
  NOR2_X1 U8874 ( .A1(n7209), .A2(n7830), .ZN(n7200) );
  INV_X1 U8875 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n7198) );
  MUX2_X1 U8876 ( .A(P2_REG1_REG_8__SCAN_IN), .B(n7198), .S(n7206), .Z(n7199)
         );
  OAI21_X1 U8877 ( .B1(n7201), .B2(n7200), .A(n7199), .ZN(n7293) );
  INV_X1 U8878 ( .A(n7293), .ZN(n7203) );
  NOR3_X1 U8879 ( .A1(n7201), .A2(n7200), .A3(n7199), .ZN(n7202) );
  NOR3_X1 U8880 ( .A1(n7203), .A2(n7202), .A3(n10510), .ZN(n7204) );
  AOI211_X1 U8881 ( .C1(n10508), .C2(P2_ADDR_REG_8__SCAN_IN), .A(n7205), .B(
        n7204), .ZN(n7213) );
  INV_X1 U8882 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n9796) );
  MUX2_X1 U8883 ( .A(P2_REG2_REG_8__SCAN_IN), .B(n9796), .S(n7206), .Z(n7211)
         );
  INV_X1 U8884 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n7208) );
  OAI21_X1 U8885 ( .B1(n7209), .B2(n7208), .A(n7207), .ZN(n7210) );
  OAI211_X1 U8886 ( .C1(n7211), .C2(n7210), .A(n10506), .B(n7297), .ZN(n7212)
         );
  OAI211_X1 U8887 ( .C1(n10509), .C2(n7298), .A(n7213), .B(n7212), .ZN(
        P2_U3253) );
  INV_X1 U8888 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n7214) );
  OAI21_X1 U8889 ( .B1(n7214), .B2(n7220), .A(n7219), .ZN(n7218) );
  INV_X1 U8890 ( .A(n10383), .ZN(n10357) );
  AOI21_X1 U8891 ( .B1(n7216), .B2(n7215), .A(n10357), .ZN(n7217) );
  AOI211_X1 U8892 ( .C1(n10395), .C2(n7218), .A(n10363), .B(n7217), .ZN(n7230)
         );
  INV_X1 U8893 ( .A(n7219), .ZN(n7224) );
  AOI21_X1 U8894 ( .B1(n7214), .B2(n7220), .A(n7629), .ZN(n7223) );
  INV_X1 U8895 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n7221) );
  NAND2_X1 U8896 ( .A1(P1_U3084), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n8233) );
  OAI21_X1 U8897 ( .B1(n10399), .B2(n7221), .A(n8233), .ZN(n7222) );
  AOI21_X1 U8898 ( .B1(n7224), .B2(n7223), .A(n7222), .ZN(n7228) );
  NAND3_X1 U8899 ( .A1(n7226), .A2(n10383), .A3(n7225), .ZN(n7227) );
  OAI211_X1 U8900 ( .C1(n7230), .C2(n7229), .A(n7228), .B(n7227), .ZN(P1_U3249) );
  INV_X1 U8901 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n7238) );
  INV_X1 U8902 ( .A(n7360), .ZN(n7231) );
  NAND2_X1 U8903 ( .A1(n7231), .A2(n7359), .ZN(n7232) );
  INV_X1 U8904 ( .A(n5737), .ZN(n7441) );
  OAI22_X1 U8905 ( .A1(n7233), .A2(n7232), .B1(n7441), .B2(n10405), .ZN(n7517)
         );
  INV_X1 U8906 ( .A(n7517), .ZN(n7236) );
  NAND2_X1 U8907 ( .A1(n7235), .A2(n7234), .ZN(n7513) );
  NAND2_X1 U8908 ( .A1(n7236), .A2(n7513), .ZN(n10244) );
  NAND2_X1 U8909 ( .A1(n10244), .A2(n10492), .ZN(n7237) );
  OAI21_X1 U8910 ( .B1(n10492), .B2(n7238), .A(n7237), .ZN(P1_U3454) );
  INV_X1 U8911 ( .A(P2_ADDR_REG_2__SCAN_IN), .ZN(n8372) );
  INV_X1 U8912 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n7687) );
  OAI22_X1 U8913 ( .A1(n8863), .A2(n8372), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7687), .ZN(n7244) );
  INV_X1 U8914 ( .A(n7239), .ZN(n7240) );
  AOI211_X1 U8915 ( .C1(n7242), .C2(n7241), .A(n7240), .B(n10510), .ZN(n7243)
         );
  AOI211_X1 U8916 ( .C1(n8870), .C2(n4515), .A(n7244), .B(n7243), .ZN(n7249)
         );
  OAI211_X1 U8917 ( .C1(n7247), .C2(n7246), .A(n10506), .B(n7245), .ZN(n7248)
         );
  NAND2_X1 U8918 ( .A1(n7249), .A2(n7248), .ZN(P2_U3247) );
  XNOR2_X1 U8919 ( .A(n7390), .B(P1_REG1_REG_10__SCAN_IN), .ZN(n7385) );
  XOR2_X1 U8920 ( .A(n7385), .B(n7386), .Z(n7261) );
  NAND2_X1 U8921 ( .A1(P1_U3084), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n8024) );
  OAI21_X1 U8922 ( .B1(n10390), .B2(n7252), .A(n8024), .ZN(n7253) );
  AOI21_X1 U8923 ( .B1(n10319), .B2(P1_ADDR_REG_10__SCAN_IN), .A(n7253), .ZN(
        n7260) );
  NAND2_X1 U8924 ( .A1(n7254), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n7255) );
  NAND2_X1 U8925 ( .A1(n7256), .A2(n7255), .ZN(n7258) );
  INV_X1 U8926 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n8064) );
  XNOR2_X1 U8927 ( .A(n7390), .B(n8064), .ZN(n7257) );
  NAND2_X1 U8928 ( .A1(n7258), .A2(n7257), .ZN(n7392) );
  OAI211_X1 U8929 ( .C1(n7258), .C2(n7257), .A(n7392), .B(n10383), .ZN(n7259)
         );
  OAI211_X1 U8930 ( .C1(n7261), .C2(n7629), .A(n7260), .B(n7259), .ZN(P1_U3251) );
  INV_X1 U8931 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n7668) );
  NOR2_X1 U8932 ( .A1(n7668), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7266) );
  OR2_X1 U8933 ( .A1(n7262), .A2(n7109), .ZN(n7264) );
  AOI211_X1 U8934 ( .C1(n10508), .C2(P2_ADDR_REG_1__SCAN_IN), .A(n7266), .B(
        n7265), .ZN(n7271) );
  OAI211_X1 U8935 ( .C1(n7269), .C2(n7268), .A(n10506), .B(n7267), .ZN(n7270)
         );
  OAI211_X1 U8936 ( .C1(n10509), .C2(n7272), .A(n7271), .B(n7270), .ZN(
        P2_U3246) );
  INV_X1 U8937 ( .A(n7273), .ZN(n7275) );
  INV_X1 U8938 ( .A(n7767), .ZN(n7761) );
  OAI222_X1 U8939 ( .A1(n9399), .A2(n7275), .B1(n7761), .B2(P2_U3152), .C1(
        n9873), .C2(n9395), .ZN(P2_U3345) );
  INV_X1 U8940 ( .A(n9602), .ZN(n9618) );
  OAI222_X1 U8941 ( .A1(P1_U3084), .A2(n9618), .B1(n10283), .B2(n7275), .C1(
        n7274), .C2(n10294), .ZN(P1_U3340) );
  INV_X1 U8942 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n7292) );
  MUX2_X1 U8943 ( .A(n7978), .B(P1_REG2_REG_3__SCAN_IN), .S(n7284), .Z(n7278)
         );
  NAND3_X1 U8944 ( .A1(n7278), .A2(n7277), .A3(n7276), .ZN(n7279) );
  NAND3_X1 U8945 ( .A1(n10383), .A2(n7280), .A3(n7279), .ZN(n7281) );
  OAI21_X1 U8946 ( .B1(n10390), .B2(n7282), .A(n7281), .ZN(n7290) );
  INV_X1 U8947 ( .A(n7283), .ZN(n7288) );
  MUX2_X1 U8948 ( .A(n7045), .B(P1_REG1_REG_3__SCAN_IN), .S(n7284), .Z(n7287)
         );
  INV_X1 U8949 ( .A(n7285), .ZN(n7286) );
  AOI211_X1 U8950 ( .C1(n7288), .C2(n7287), .A(n7286), .B(n7629), .ZN(n7289)
         );
  AOI211_X1 U8951 ( .C1(P1_REG3_REG_3__SCAN_IN), .C2(P1_U3084), .A(n7290), .B(
        n7289), .ZN(n7291) );
  OAI21_X1 U8952 ( .B1(n10399), .B2(n7292), .A(n7291), .ZN(P1_U3244) );
  XNOR2_X1 U8953 ( .A(n7335), .B(P2_REG1_REG_10__SCAN_IN), .ZN(n7331) );
  OAI21_X1 U8954 ( .B1(n7198), .B2(n7298), .A(n7293), .ZN(n7309) );
  XOR2_X1 U8955 ( .A(P2_REG1_REG_9__SCAN_IN), .B(n7299), .Z(n7308) );
  XOR2_X1 U8956 ( .A(n7331), .B(n7332), .Z(n7304) );
  NOR2_X1 U8957 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7294), .ZN(n7295) );
  AOI21_X1 U8958 ( .B1(n10508), .B2(P2_ADDR_REG_10__SCAN_IN), .A(n7295), .ZN(
        n7296) );
  OAI21_X1 U8959 ( .B1(n10509), .B2(n7330), .A(n7296), .ZN(n7303) );
  XOR2_X1 U8960 ( .A(P2_REG2_REG_9__SCAN_IN), .B(n7299), .Z(n7316) );
  XNOR2_X1 U8961 ( .A(n7335), .B(P2_REG2_REG_10__SCAN_IN), .ZN(n7300) );
  NOR2_X1 U8962 ( .A1(n7301), .A2(n7300), .ZN(n7334) );
  AOI211_X1 U8963 ( .C1(n7301), .C2(n7300), .A(n10511), .B(n7334), .ZN(n7302)
         );
  AOI211_X1 U8964 ( .C1(n10505), .C2(n7304), .A(n7303), .B(n7302), .ZN(n7305)
         );
  INV_X1 U8965 ( .A(n7305), .ZN(P2_U3255) );
  INV_X1 U8966 ( .A(n7306), .ZN(n7320) );
  INV_X1 U8967 ( .A(n8539), .ZN(n8550) );
  OAI222_X1 U8968 ( .A1(n9399), .A2(n7320), .B1(n8550), .B2(P2_U3152), .C1(
        n7307), .C2(n9395), .ZN(P2_U3344) );
  XNOR2_X1 U8969 ( .A(n7309), .B(n7308), .ZN(n7319) );
  NAND2_X1 U8970 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(P2_U3152), .ZN(n7752) );
  INV_X1 U8971 ( .A(n7752), .ZN(n7312) );
  NOR2_X1 U8972 ( .A1(n10509), .A2(n7310), .ZN(n7311) );
  AOI211_X1 U8973 ( .C1(n10508), .C2(P2_ADDR_REG_9__SCAN_IN), .A(n7312), .B(
        n7311), .ZN(n7318) );
  INV_X1 U8974 ( .A(n7313), .ZN(n7314) );
  OAI211_X1 U8975 ( .C1(n7316), .C2(n7315), .A(n7314), .B(n10506), .ZN(n7317)
         );
  OAI211_X1 U8976 ( .C1(n7319), .C2(n10510), .A(n7318), .B(n7317), .ZN(
        P2_U3254) );
  OAI222_X1 U8977 ( .A1(P1_U3084), .A2(n9619), .B1(n10292), .B2(n7320), .C1(
        n9886), .C2(n10294), .ZN(P1_U3339) );
  NAND2_X1 U8978 ( .A1(n8832), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n7321) );
  OAI21_X1 U8979 ( .B1(n9036), .B2(n8832), .A(n7321), .ZN(P2_U3577) );
  OAI21_X1 U8980 ( .B1(n7324), .B2(n7323), .A(n7322), .ZN(n7326) );
  OAI22_X1 U8981 ( .A1(n7521), .A2(n9203), .B1(n7325), .B2(n9205), .ZN(n7567)
         );
  AOI22_X1 U8982 ( .A1(n6894), .A2(n7326), .B1(n8816), .B2(n7567), .ZN(n7329)
         );
  INV_X1 U8983 ( .A(n7522), .ZN(n7327) );
  NAND2_X1 U8984 ( .A1(n7327), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8801) );
  AOI22_X1 U8985 ( .A1(n8801), .A2(P2_REG3_REG_1__SCAN_IN), .B1(n8825), .B2(
        n7671), .ZN(n7328) );
  NAND2_X1 U8986 ( .A1(n7329), .A2(n7328), .ZN(P2_U3224) );
  INV_X1 U8987 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n8249) );
  INV_X1 U8988 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n7333) );
  XNOR2_X1 U8989 ( .A(n7478), .B(n7333), .ZN(n7474) );
  XNOR2_X1 U8990 ( .A(n7475), .B(n7474), .ZN(n7344) );
  XOR2_X1 U8991 ( .A(P2_REG2_REG_11__SCAN_IN), .B(n7478), .Z(n7337) );
  OAI21_X1 U8992 ( .B1(n7337), .B2(n7336), .A(n7477), .ZN(n7338) );
  NAND2_X1 U8993 ( .A1(n7338), .A2(n10506), .ZN(n7343) );
  NOR2_X1 U8994 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6260), .ZN(n7341) );
  NOR2_X1 U8995 ( .A1(n10509), .A2(n7339), .ZN(n7340) );
  AOI211_X1 U8996 ( .C1(n10508), .C2(P2_ADDR_REG_11__SCAN_IN), .A(n7341), .B(
        n7340), .ZN(n7342) );
  OAI211_X1 U8997 ( .C1(n7344), .C2(n10510), .A(n7343), .B(n7342), .ZN(
        P2_U3256) );
  XNOR2_X1 U8998 ( .A(n7349), .B(n7345), .ZN(n7950) );
  INV_X1 U8999 ( .A(n10240), .ZN(n10485) );
  INV_X1 U9000 ( .A(n7793), .ZN(n7347) );
  INV_X1 U9001 ( .A(n7378), .ZN(n7346) );
  OAI211_X1 U9002 ( .C1(n4391), .C2(n7347), .A(n7346), .B(n10418), .ZN(n7943)
         );
  OAI21_X1 U9003 ( .B1(n4391), .B2(n10485), .A(n7943), .ZN(n7353) );
  XNOR2_X1 U9004 ( .A(n7348), .B(n7349), .ZN(n7352) );
  INV_X1 U9005 ( .A(n7424), .ZN(n10482) );
  NAND2_X1 U9006 ( .A1(n7950), .A2(n10482), .ZN(n7351) );
  INV_X1 U9007 ( .A(n10405), .ZN(n8217) );
  AOI22_X1 U9008 ( .A1(n10103), .A2(n5737), .B1(n9588), .B2(n8217), .ZN(n7350)
         );
  OAI211_X1 U9009 ( .C1(n10406), .C2(n7352), .A(n7351), .B(n7350), .ZN(n7947)
         );
  AOI211_X1 U9010 ( .C1(n10465), .C2(n7950), .A(n7353), .B(n7947), .ZN(n10445)
         );
  NAND2_X1 U9011 ( .A1(n10168), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n7354) );
  OAI21_X1 U9012 ( .B1(n10445), .B2(n10168), .A(n7354), .ZN(P1_U3525) );
  INV_X1 U9013 ( .A(n7355), .ZN(n7357) );
  INV_X1 U9014 ( .A(n7371), .ZN(n7374) );
  NOR2_X1 U9015 ( .A1(n7359), .A2(n7806), .ZN(n7801) );
  OAI21_X1 U9016 ( .B1(n7360), .B2(n7801), .A(n10428), .ZN(n7361) );
  INV_X1 U9017 ( .A(n7361), .ZN(n7362) );
  NAND2_X1 U9018 ( .A1(n7374), .A2(n7362), .ZN(n7501) );
  INV_X1 U9019 ( .A(n7364), .ZN(n7365) );
  NAND2_X1 U9020 ( .A1(n7371), .A2(n7365), .ZN(n7439) );
  NOR2_X1 U9021 ( .A1(n10240), .A2(n7367), .ZN(n7373) );
  INV_X1 U9022 ( .A(n7373), .ZN(n7369) );
  INV_X1 U9023 ( .A(n10428), .ZN(n7368) );
  NOR2_X1 U9024 ( .A1(n7369), .A2(n7368), .ZN(n7370) );
  AOI22_X1 U9025 ( .A1(n9534), .A2(n5737), .B1(n9547), .B2(n7372), .ZN(n7376)
         );
  NAND2_X1 U9026 ( .A1(n7374), .A2(n7373), .ZN(n7499) );
  NAND2_X1 U9027 ( .A1(n9532), .A2(n7499), .ZN(n7452) );
  NAND2_X1 U9028 ( .A1(n7452), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n7375) );
  OAI211_X1 U9029 ( .C1(n9556), .C2(n7794), .A(n7376), .B(n7375), .ZN(P1_U3230) );
  XNOR2_X1 U9030 ( .A(n7377), .B(n7380), .ZN(n7975) );
  OR2_X1 U9031 ( .A1(n7378), .A2(n7979), .ZN(n7379) );
  AND3_X1 U9032 ( .A1(n7921), .A2(n10418), .A3(n7379), .ZN(n7981) );
  XNOR2_X1 U9033 ( .A(n7380), .B(n5907), .ZN(n7381) );
  OAI222_X1 U9034 ( .A1(n7381), .A2(n10406), .B1(n10405), .B2(n10402), .C1(
        n10403), .C2(n7495), .ZN(n7976) );
  AOI211_X1 U9035 ( .C1(n10489), .C2(n7975), .A(n7981), .B(n7976), .ZN(n7531)
         );
  INV_X1 U9036 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n7382) );
  OAI22_X1 U9037 ( .A1(n10275), .A2(n7979), .B1(n10492), .B2(n7382), .ZN(n7383) );
  INV_X1 U9038 ( .A(n7383), .ZN(n7384) );
  OAI21_X1 U9039 ( .B1(n7531), .B2(n10490), .A(n7384), .ZN(P1_U3463) );
  OAI22_X1 U9040 ( .A1(n7386), .A2(n7385), .B1(n7390), .B2(
        P1_REG1_REG_10__SCAN_IN), .ZN(n7462) );
  NAND2_X1 U9041 ( .A1(n7393), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n7461) );
  NAND2_X1 U9042 ( .A1(n4415), .A2(n7461), .ZN(n7387) );
  XNOR2_X1 U9043 ( .A(n7462), .B(n7387), .ZN(n7401) );
  NAND2_X1 U9044 ( .A1(P1_U3084), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n8205) );
  OAI21_X1 U9045 ( .B1(n10390), .B2(n7388), .A(n8205), .ZN(n7389) );
  AOI21_X1 U9046 ( .B1(n10319), .B2(P1_ADDR_REG_11__SCAN_IN), .A(n7389), .ZN(
        n7400) );
  NAND2_X1 U9047 ( .A1(n7390), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n7391) );
  AND2_X1 U9048 ( .A1(n7393), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n7395) );
  OR2_X1 U9049 ( .A1(n7393), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n7466) );
  INV_X1 U9050 ( .A(n7466), .ZN(n7397) );
  OAI21_X1 U9051 ( .B1(n7397), .B2(n7395), .A(n7394), .ZN(n7396) );
  OAI21_X1 U9052 ( .B1(n7467), .B2(n7397), .A(n7396), .ZN(n7398) );
  NAND2_X1 U9053 ( .A1(n7398), .A2(n10383), .ZN(n7399) );
  OAI211_X1 U9054 ( .C1(n7401), .C2(n7629), .A(n7400), .B(n7399), .ZN(P1_U3252) );
  NAND3_X1 U9055 ( .A1(n10383), .A2(P1_REG2_REG_4__SCAN_IN), .A3(n7412), .ZN(
        n7403) );
  NAND3_X1 U9056 ( .A1(n10395), .A2(P1_REG1_REG_4__SCAN_IN), .A3(n7405), .ZN(
        n7402) );
  NAND3_X1 U9057 ( .A1(n10390), .A2(n7403), .A3(n7402), .ZN(n7420) );
  INV_X1 U9058 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n9855) );
  NAND3_X1 U9059 ( .A1(n7405), .A2(n7404), .A3(n7410), .ZN(n7406) );
  NAND2_X1 U9060 ( .A1(n7407), .A2(n7406), .ZN(n7409) );
  NAND2_X1 U9061 ( .A1(P1_U3084), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n7739) );
  INV_X1 U9062 ( .A(n7739), .ZN(n7408) );
  AOI21_X1 U9063 ( .B1(n10395), .B2(n7409), .A(n7408), .ZN(n7417) );
  NAND3_X1 U9064 ( .A1(n7412), .A2(n7411), .A3(n7410), .ZN(n7413) );
  NAND2_X1 U9065 ( .A1(n7414), .A2(n7413), .ZN(n7415) );
  NAND2_X1 U9066 ( .A1(n10383), .A2(n7415), .ZN(n7416) );
  OAI211_X1 U9067 ( .C1(n9855), .C2(n10399), .A(n7417), .B(n7416), .ZN(n7419)
         );
  AOI211_X1 U9068 ( .C1(n7421), .C2(n7420), .A(n7419), .B(n7418), .ZN(n7422)
         );
  INV_X1 U9069 ( .A(n7422), .ZN(P1_U3245) );
  AOI22_X1 U9070 ( .A1(n5737), .A2(n6956), .B1(n8592), .B2(n7802), .ZN(n7426)
         );
  XNOR2_X1 U9071 ( .A(n8476), .B(n7426), .ZN(n7448) );
  NOR2_X1 U9072 ( .A1(n8593), .A2(n6054), .ZN(n7427) );
  AOI21_X1 U9073 ( .B1(n8496), .B2(n5737), .A(n7427), .ZN(n7446) );
  INV_X1 U9074 ( .A(n7428), .ZN(n7429) );
  NAND2_X1 U9075 ( .A1(n7429), .A2(n8476), .ZN(n7430) );
  OAI21_X1 U9076 ( .B1(n7448), .B2(n7446), .A(n7447), .ZN(n7433) );
  NAND2_X1 U9077 ( .A1(n7448), .A2(n7446), .ZN(n7432) );
  NAND2_X1 U9078 ( .A1(n7433), .A2(n7432), .ZN(n7487) );
  OAI22_X1 U9079 ( .A1(n7495), .A2(n8593), .B1(n4391), .B2(n7865), .ZN(n7434)
         );
  XNOR2_X1 U9080 ( .A(n7434), .B(n8476), .ZN(n7490) );
  OR2_X1 U9081 ( .A1(n7495), .A2(n8599), .ZN(n7437) );
  NAND2_X1 U9082 ( .A1(n6956), .A2(n7435), .ZN(n7436) );
  NAND2_X1 U9083 ( .A1(n7437), .A2(n7436), .ZN(n7489) );
  INV_X1 U9084 ( .A(n7489), .ZN(n7438) );
  XNOR2_X1 U9085 ( .A(n7490), .B(n7438), .ZN(n7488) );
  XOR2_X1 U9086 ( .A(n7487), .B(n7488), .Z(n7445) );
  OAI22_X1 U9087 ( .A1(n7441), .A2(n9494), .B1(n9555), .B2(n7440), .ZN(n7443)
         );
  NOR2_X1 U9088 ( .A1(n9556), .A2(n4391), .ZN(n7442) );
  AOI211_X1 U9089 ( .C1(P1_REG3_REG_2__SCAN_IN), .C2(n7452), .A(n7443), .B(
        n7442), .ZN(n7444) );
  OAI21_X1 U9090 ( .B1(n9520), .B2(n7445), .A(n7444), .ZN(P1_U3235) );
  XNOR2_X1 U9091 ( .A(n7447), .B(n7446), .ZN(n7449) );
  XNOR2_X1 U9092 ( .A(n7448), .B(n7449), .ZN(n7454) );
  INV_X1 U9093 ( .A(n9590), .ZN(n7798) );
  OAI22_X1 U9094 ( .A1(n7798), .A2(n9494), .B1(n9555), .B2(n7495), .ZN(n7451)
         );
  NOR2_X1 U9095 ( .A1(n9556), .A2(n6054), .ZN(n7450) );
  AOI211_X1 U9096 ( .C1(P1_REG3_REG_1__SCAN_IN), .C2(n7452), .A(n7451), .B(
        n7450), .ZN(n7453) );
  OAI21_X1 U9097 ( .B1(n9520), .B2(n7454), .A(n7453), .ZN(P1_U3220) );
  INV_X1 U9098 ( .A(n7455), .ZN(n7457) );
  INV_X1 U9099 ( .A(n10346), .ZN(n9621) );
  OAI222_X1 U9100 ( .A1(n10294), .A2(n7456), .B1(n10283), .B2(n7457), .C1(
        P1_U3084), .C2(n9621), .ZN(P1_U3338) );
  INV_X1 U9101 ( .A(n8852), .ZN(n8551) );
  OAI222_X1 U9102 ( .A1(n9395), .A2(n9860), .B1(n9399), .B2(n7457), .C1(
        P2_U3152), .C2(n8551), .ZN(P2_U3343) );
  INV_X1 U9103 ( .A(n7458), .ZN(n7508) );
  AOI22_X1 U9104 ( .A1(n8869), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_16__SCAN_IN), .B2(n9388), .ZN(n7459) );
  OAI21_X1 U9105 ( .B1(n7508), .B2(n9399), .A(n7459), .ZN(P2_U3342) );
  INV_X1 U9106 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n8355) );
  NAND2_X1 U9107 ( .A1(n7460), .A2(n8355), .ZN(n7616) );
  OAI21_X1 U9108 ( .B1(n7460), .B2(n8355), .A(n7616), .ZN(n7464) );
  AOI21_X1 U9109 ( .B1(n7464), .B2(n7463), .A(n7617), .ZN(n7472) );
  NOR2_X1 U9110 ( .A1(n9805), .A2(P1_STATE_REG_SCAN_IN), .ZN(n8323) );
  INV_X1 U9111 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n9939) );
  NOR2_X1 U9112 ( .A1(n10399), .A2(n9939), .ZN(n7465) );
  AOI211_X1 U9113 ( .C1(n10363), .C2(n7622), .A(n8323), .B(n7465), .ZN(n7471)
         );
  INV_X1 U9114 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n9819) );
  XNOR2_X1 U9115 ( .A(n7622), .B(n9819), .ZN(n7468) );
  OAI211_X1 U9116 ( .C1(n7469), .C2(n7468), .A(n7624), .B(n10383), .ZN(n7470)
         );
  OAI211_X1 U9117 ( .C1(n7472), .C2(n7629), .A(n7471), .B(n7470), .ZN(P1_U3253) );
  NAND2_X1 U9118 ( .A1(n9576), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n7473) );
  OAI21_X1 U9119 ( .B1(n8610), .B2(n9576), .A(n7473), .ZN(P1_U3584) );
  XNOR2_X1 U9120 ( .A(n7646), .B(P2_REG1_REG_12__SCAN_IN), .ZN(n7635) );
  XNOR2_X1 U9121 ( .A(n7634), .B(n7635), .ZN(n7486) );
  INV_X1 U9122 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n7476) );
  MUX2_X1 U9123 ( .A(P2_REG2_REG_12__SCAN_IN), .B(n7476), .S(n7646), .Z(n7480)
         );
  OAI21_X1 U9124 ( .B1(P2_REG2_REG_11__SCAN_IN), .B2(n7478), .A(n7477), .ZN(
        n7479) );
  NAND2_X1 U9125 ( .A1(n7479), .A2(n7480), .ZN(n7645) );
  OAI21_X1 U9126 ( .B1(n7480), .B2(n7479), .A(n7645), .ZN(n7481) );
  NAND2_X1 U9127 ( .A1(n7481), .A2(n10506), .ZN(n7485) );
  INV_X1 U9128 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n7482) );
  NAND2_X1 U9129 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(P2_U3152), .ZN(n8078) );
  OAI21_X1 U9130 ( .B1(n8863), .B2(n7482), .A(n8078), .ZN(n7483) );
  AOI21_X1 U9131 ( .B1(n8870), .B2(n7646), .A(n7483), .ZN(n7484) );
  OAI211_X1 U9132 ( .C1(n7486), .C2(n10510), .A(n7485), .B(n7484), .ZN(
        P2_U3257) );
  NAND2_X1 U9133 ( .A1(n7488), .A2(n7487), .ZN(n7492) );
  OR2_X1 U9134 ( .A1(n7490), .A2(n7489), .ZN(n7491) );
  NAND2_X1 U9135 ( .A1(n9588), .A2(n6956), .ZN(n7493) );
  OAI21_X1 U9136 ( .B1(n7979), .B2(n7865), .A(n7493), .ZN(n7494) );
  XNOR2_X1 U9137 ( .A(n8476), .B(n7494), .ZN(n7729) );
  AOI22_X1 U9138 ( .A1(n8496), .A2(n9588), .B1(n7529), .B2(n6956), .ZN(n7730)
         );
  XNOR2_X1 U9139 ( .A(n7729), .B(n7730), .ZN(n7727) );
  XOR2_X1 U9140 ( .A(n7728), .B(n7727), .Z(n7506) );
  OAI22_X1 U9141 ( .A1(n7495), .A2(n9494), .B1(n9555), .B2(n10402), .ZN(n7504)
         );
  NAND4_X1 U9142 ( .A1(n7499), .A2(n4520), .A3(n7497), .A4(n7496), .ZN(n7500)
         );
  NAND2_X1 U9143 ( .A1(n7500), .A2(P1_STATE_REG_SCAN_IN), .ZN(n7502) );
  MUX2_X1 U9144 ( .A(n9560), .B(P1_U3084), .S(P1_REG3_REG_3__SCAN_IN), .Z(
        n7503) );
  AOI211_X1 U9145 ( .C1(n9518), .C2(n7529), .A(n7504), .B(n7503), .ZN(n7505)
         );
  OAI21_X1 U9146 ( .B1(n9520), .B2(n7506), .A(n7505), .ZN(P1_U3216) );
  INV_X1 U9147 ( .A(n10362), .ZN(n9623) );
  OAI222_X1 U9148 ( .A1(P1_U3084), .A2(n9623), .B1(n10292), .B2(n7508), .C1(
        n7507), .C2(n10294), .ZN(P1_U3337) );
  INV_X1 U9149 ( .A(n7509), .ZN(n7512) );
  INV_X1 U9150 ( .A(n7510), .ZN(n7511) );
  INV_X1 U9151 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n7519) );
  INV_X1 U9152 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n7515) );
  INV_X1 U9153 ( .A(n7791), .ZN(n7514) );
  OAI22_X1 U9154 ( .A1(n10145), .A2(n7515), .B1(n7514), .B2(n7513), .ZN(n7516)
         );
  OAI21_X1 U9155 ( .B1(n7517), .B2(n7516), .A(n10148), .ZN(n7518) );
  OAI21_X1 U9156 ( .B1(n10148), .B2(n7519), .A(n7518), .ZN(P1_U3291) );
  NOR2_X1 U9157 ( .A1(n8821), .A2(n7520), .ZN(n8826) );
  INV_X1 U9158 ( .A(n8826), .ZN(n8793) );
  OAI22_X1 U9159 ( .A1(n8793), .A2(n7521), .B1(n8821), .B2(n7570), .ZN(n7527)
         );
  AND2_X1 U9160 ( .A1(P2_U3152), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n10507) );
  AOI21_X1 U9161 ( .B1(n7522), .B2(P2_REG3_REG_0__SCAN_IN), .A(n10507), .ZN(
        n7524) );
  NAND2_X1 U9162 ( .A1(n8825), .A2(n10569), .ZN(n7523) );
  OAI211_X1 U9163 ( .C1(n8785), .C2(n6911), .A(n7524), .B(n7523), .ZN(n7525)
         );
  AOI21_X1 U9164 ( .B1(n7527), .B2(n7526), .A(n7525), .ZN(n7528) );
  INV_X1 U9165 ( .A(n7528), .ZN(P2_U3234) );
  AOI22_X1 U9166 ( .A1(n6884), .A2(n7529), .B1(n10168), .B2(
        P1_REG1_REG_3__SCAN_IN), .ZN(n7530) );
  OAI21_X1 U9167 ( .B1(n7531), .B2(n10168), .A(n7530), .ZN(P1_U3526) );
  OR2_X1 U9168 ( .A1(n7536), .A2(n7540), .ZN(n7537) );
  NAND2_X1 U9169 ( .A1(n7538), .A2(n7537), .ZN(n10518) );
  INV_X1 U9170 ( .A(n10518), .ZN(n7548) );
  AND2_X1 U9171 ( .A1(n4396), .A2(n6625), .ZN(n7539) );
  NAND2_X1 U9172 ( .A1(n7539), .A2(n8535), .ZN(n10586) );
  INV_X1 U9173 ( .A(n7666), .ZN(n8086) );
  XNOR2_X1 U9174 ( .A(n7541), .B(n7540), .ZN(n7543) );
  OAI21_X1 U9175 ( .B1(n7543), .B2(n9200), .A(n7542), .ZN(n7544) );
  AOI21_X1 U9176 ( .B1(n8086), .B2(n10518), .A(n7544), .ZN(n10528) );
  INV_X2 U9177 ( .A(n10588), .ZN(n9356) );
  AOI21_X1 U9178 ( .B1(n7582), .B2(n7546), .A(n10590), .ZN(n7545) );
  AND2_X1 U9179 ( .A1(n7545), .A2(n7556), .ZN(n10520) );
  AOI21_X1 U9180 ( .B1(n9356), .B2(n7546), .A(n10520), .ZN(n7547) );
  OAI211_X1 U9181 ( .C1(n7548), .C2(n10586), .A(n10528), .B(n7547), .ZN(n7589)
         );
  NAND2_X1 U9182 ( .A1(n7589), .A2(n10598), .ZN(n7549) );
  OAI21_X1 U9183 ( .B1(n10598), .B2(n6147), .A(n7549), .ZN(P2_U3460) );
  INV_X1 U9184 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n7560) );
  OAI21_X1 U9185 ( .B1(n7551), .B2(n7552), .A(n7550), .ZN(n7684) );
  INV_X1 U9186 ( .A(n7684), .ZN(n7558) );
  AOI21_X1 U9187 ( .B1(n7553), .B2(n7552), .A(n9200), .ZN(n7555) );
  OAI22_X1 U9188 ( .A1(n7781), .A2(n9205), .B1(n7580), .B2(n9203), .ZN(n8758)
         );
  AOI21_X1 U9189 ( .B1(n7555), .B2(n7713), .A(n8758), .ZN(n7681) );
  AOI211_X1 U9190 ( .C1(n8759), .C2(n7556), .A(n10590), .B(n7719), .ZN(n7677)
         );
  AOI21_X1 U9191 ( .B1(n9356), .B2(n8759), .A(n7677), .ZN(n7557) );
  OAI211_X1 U9192 ( .C1(n7558), .C2(n9350), .A(n7681), .B(n7557), .ZN(n7594)
         );
  NAND2_X1 U9193 ( .A1(n7594), .A2(n10598), .ZN(n7559) );
  OAI21_X1 U9194 ( .B1(n10598), .B2(n7560), .A(n7559), .ZN(P2_U3463) );
  INV_X1 U9195 ( .A(n7563), .ZN(n7566) );
  INV_X1 U9196 ( .A(n7564), .ZN(n7565) );
  AOI21_X1 U9197 ( .B1(n7566), .B2(n6909), .A(n7565), .ZN(n7676) );
  XNOR2_X1 U9198 ( .A(n7563), .B(n7696), .ZN(n7568) );
  AOI21_X1 U9199 ( .B1(n7568), .B2(n9225), .A(n7567), .ZN(n7673) );
  INV_X1 U9200 ( .A(n7569), .ZN(n7584) );
  OAI211_X1 U9201 ( .C1(n7571), .C2(n7570), .A(n7584), .B(n9357), .ZN(n7669)
         );
  INV_X1 U9202 ( .A(n7669), .ZN(n7572) );
  AOI21_X1 U9203 ( .B1(n9356), .B2(n7671), .A(n7572), .ZN(n7573) );
  OAI211_X1 U9204 ( .C1(n7676), .C2(n9350), .A(n7673), .B(n7573), .ZN(n7596)
         );
  NAND2_X1 U9205 ( .A1(n7596), .A2(n10605), .ZN(n7574) );
  OAI21_X1 U9206 ( .B1(n10605), .B2(n7575), .A(n7574), .ZN(P2_U3521) );
  OAI21_X1 U9207 ( .B1(n7577), .B2(n7578), .A(n7576), .ZN(n7693) );
  INV_X1 U9208 ( .A(n7693), .ZN(n7586) );
  XNOR2_X1 U9209 ( .A(n7579), .B(n7578), .ZN(n7581) );
  OAI22_X1 U9210 ( .A1(n7580), .A2(n9205), .B1(n6911), .B2(n9203), .ZN(n8798)
         );
  AOI21_X1 U9211 ( .B1(n7581), .B2(n9225), .A(n8798), .ZN(n7689) );
  INV_X1 U9212 ( .A(n7582), .ZN(n7583) );
  AOI21_X1 U9213 ( .B1(n9356), .B2(n8800), .A(n7692), .ZN(n7585) );
  OAI211_X1 U9214 ( .C1(n7586), .C2(n9350), .A(n7689), .B(n7585), .ZN(n7592)
         );
  NAND2_X1 U9215 ( .A1(n7592), .A2(n10605), .ZN(n7587) );
  OAI21_X1 U9216 ( .B1(n10605), .B2(n7588), .A(n7587), .ZN(P2_U3522) );
  NAND2_X1 U9217 ( .A1(n7589), .A2(n10605), .ZN(n7590) );
  OAI21_X1 U9218 ( .B1(n10605), .B2(n7591), .A(n7590), .ZN(P2_U3523) );
  NAND2_X1 U9219 ( .A1(n7592), .A2(n10598), .ZN(n7593) );
  OAI21_X1 U9220 ( .B1(n10598), .B2(n6140), .A(n7593), .ZN(P2_U3457) );
  NAND2_X1 U9221 ( .A1(n7594), .A2(n10605), .ZN(n7595) );
  OAI21_X1 U9222 ( .B1(n10605), .B2(n7111), .A(n7595), .ZN(P2_U3524) );
  INV_X1 U9223 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n9950) );
  NAND2_X1 U9224 ( .A1(n7596), .A2(n10598), .ZN(n7597) );
  OAI21_X1 U9225 ( .B1(n10598), .B2(n9950), .A(n7597), .ZN(P2_U3454) );
  XNOR2_X1 U9226 ( .A(n7599), .B(n7598), .ZN(n8762) );
  NAND3_X1 U9227 ( .A1(n8756), .A2(n7600), .A3(n8762), .ZN(n8755) );
  NAND2_X1 U9228 ( .A1(n8755), .A2(n7601), .ZN(n8727) );
  INV_X1 U9229 ( .A(n7602), .ZN(n7604) );
  NAND2_X1 U9230 ( .A1(n7604), .A2(n7603), .ZN(n8728) );
  NOR2_X1 U9231 ( .A1(n8727), .A2(n8728), .ZN(n8726) );
  INV_X1 U9232 ( .A(n7606), .ZN(n7607) );
  AOI21_X1 U9233 ( .B1(n8726), .B2(n7605), .A(n7607), .ZN(n7615) );
  OAI22_X1 U9234 ( .A1(n8785), .A2(n8690), .B1(n8695), .B2(n10579), .ZN(n7608)
         );
  AOI211_X1 U9235 ( .C1(n7784), .C2(n8761), .A(n7609), .B(n7608), .ZN(n7614)
         );
  INV_X1 U9236 ( .A(n7605), .ZN(n7610) );
  NOR3_X1 U9237 ( .A1(n8793), .A2(n7611), .A3(n7610), .ZN(n7612) );
  INV_X1 U9238 ( .A(n8786), .ZN(n8697) );
  OAI21_X1 U9239 ( .B1(n7612), .B2(n8697), .A(n8841), .ZN(n7613) );
  OAI211_X1 U9240 ( .C1(n7615), .C2(n8821), .A(n7614), .B(n7613), .ZN(P2_U3241) );
  XNOR2_X1 U9241 ( .A(n9602), .B(P1_REG1_REG_13__SCAN_IN), .ZN(n7618) );
  AOI21_X1 U9242 ( .B1(n4498), .B2(n7618), .A(n9616), .ZN(n7630) );
  NOR2_X1 U9243 ( .A1(n7619), .A2(P1_STATE_REG_SCAN_IN), .ZN(n8282) );
  INV_X1 U9244 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n7620) );
  NOR2_X1 U9245 ( .A1(n10399), .A2(n7620), .ZN(n7621) );
  AOI211_X1 U9246 ( .C1(n10363), .C2(n9602), .A(n8282), .B(n7621), .ZN(n7628)
         );
  NAND2_X1 U9247 ( .A1(n7622), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n7623) );
  NAND2_X1 U9248 ( .A1(n7624), .A2(n7623), .ZN(n7626) );
  INV_X1 U9249 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n9803) );
  MUX2_X1 U9250 ( .A(P1_REG2_REG_13__SCAN_IN), .B(n9803), .S(n9602), .Z(n7625)
         );
  NAND2_X1 U9251 ( .A1(n7626), .A2(n7625), .ZN(n9604) );
  OAI211_X1 U9252 ( .C1(n7626), .C2(n7625), .A(n9604), .B(n10383), .ZN(n7627)
         );
  OAI211_X1 U9253 ( .C1(n7630), .C2(n7629), .A(n7628), .B(n7627), .ZN(P1_U3254) );
  INV_X1 U9254 ( .A(n7631), .ZN(n7654) );
  INV_X1 U9255 ( .A(n8543), .ZN(n8881) );
  OAI222_X1 U9256 ( .A1(n9399), .A2(n7654), .B1(n8881), .B2(P2_U3152), .C1(
        n7632), .C2(n9395), .ZN(P2_U3341) );
  NAND2_X1 U9257 ( .A1(n8832), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n7633) );
  OAI21_X1 U9258 ( .B1(n8969), .B2(n8832), .A(n7633), .ZN(P2_U3581) );
  INV_X1 U9259 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n9964) );
  NOR2_X1 U9260 ( .A1(n7636), .A2(n7635), .ZN(n7637) );
  AOI21_X1 U9261 ( .B1(n7638), .B2(n9964), .A(n7637), .ZN(n7640) );
  INV_X1 U9262 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n7760) );
  AOI22_X1 U9263 ( .A1(n7767), .A2(n7760), .B1(P2_REG1_REG_13__SCAN_IN), .B2(
        n7761), .ZN(n7639) );
  AOI21_X1 U9264 ( .B1(n7640), .B2(n7639), .A(n7759), .ZN(n7652) );
  INV_X1 U9265 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n7642) );
  AND2_X1 U9266 ( .A1(P2_U3152), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n8189) );
  INV_X1 U9267 ( .A(n8189), .ZN(n7641) );
  OAI21_X1 U9268 ( .B1(n8863), .B2(n7642), .A(n7641), .ZN(n7643) );
  AOI21_X1 U9269 ( .B1(n8870), .B2(n7767), .A(n7643), .ZN(n7651) );
  NOR2_X1 U9270 ( .A1(n7767), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n7644) );
  AOI21_X1 U9271 ( .B1(P2_REG2_REG_13__SCAN_IN), .B2(n7767), .A(n7644), .ZN(
        n7648) );
  OAI21_X1 U9272 ( .B1(n7648), .B2(n7647), .A(n7766), .ZN(n7649) );
  NAND2_X1 U9273 ( .A1(n7649), .A2(n10506), .ZN(n7650) );
  OAI211_X1 U9274 ( .C1(n7652), .C2(n10510), .A(n7651), .B(n7650), .ZN(
        P2_U3258) );
  INV_X1 U9275 ( .A(n9626), .ZN(n10375) );
  OAI222_X1 U9276 ( .A1(P1_U3084), .A2(n10375), .B1(n10292), .B2(n7654), .C1(
        n7653), .C2(n10294), .ZN(P1_U3336) );
  INV_X1 U9277 ( .A(n7655), .ZN(n7686) );
  AOI22_X1 U9278 ( .A1(n8547), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_18__SCAN_IN), .B2(n9388), .ZN(n7656) );
  OAI21_X1 U9279 ( .B1(n7686), .B2(n9399), .A(n7656), .ZN(P2_U3340) );
  INV_X1 U9280 ( .A(n7657), .ZN(n7658) );
  AOI211_X1 U9281 ( .C1(n7660), .C2(n7659), .A(n8821), .B(n7658), .ZN(n7664)
         );
  INV_X1 U9282 ( .A(n8840), .ZN(n7716) );
  INV_X1 U9283 ( .A(n8785), .ZN(n8694) );
  AOI22_X1 U9284 ( .A1(n8694), .A2(n8838), .B1(n8761), .B2(n7813), .ZN(n7662)
         );
  AOI22_X1 U9285 ( .A1(n8825), .A2(n7824), .B1(P2_REG3_REG_7__SCAN_IN), .B2(
        P2_U3152), .ZN(n7661) );
  OAI211_X1 U9286 ( .C1(n7716), .C2(n8786), .A(n7662), .B(n7661), .ZN(n7663)
         );
  OR2_X1 U9287 ( .A1(n7664), .A2(n7663), .ZN(P2_U3215) );
  AND2_X1 U9288 ( .A1(n7666), .A2(n7665), .ZN(n7667) );
  OAI22_X1 U9289 ( .A1(n7718), .A2(n7669), .B1(n7668), .B2(n9188), .ZN(n7670)
         );
  AOI21_X1 U9290 ( .B1(n9190), .B2(n7671), .A(n7670), .ZN(n7675) );
  MUX2_X1 U9291 ( .A(n7673), .B(n7672), .S(n4392), .Z(n7674) );
  OAI211_X1 U9292 ( .C1(n7676), .C2(n9231), .A(n7675), .B(n7674), .ZN(P2_U3295) );
  INV_X1 U9293 ( .A(n9231), .ZN(n9056) );
  AOI22_X1 U9294 ( .A1(n9158), .A2(n7677), .B1(n8760), .B2(n10517), .ZN(n7678)
         );
  OAI21_X1 U9295 ( .B1(n7679), .B2(n9060), .A(n7678), .ZN(n7683) );
  OAI22_X1 U9296 ( .A1(n7681), .A2(n4392), .B1(n7680), .B2(n10523), .ZN(n7682)
         );
  AOI211_X1 U9297 ( .C1(n9056), .C2(n7684), .A(n7683), .B(n7682), .ZN(n7685)
         );
  INV_X1 U9298 ( .A(n7685), .ZN(P2_U3292) );
  INV_X1 U9299 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n9827) );
  INV_X1 U9300 ( .A(n9627), .ZN(n10389) );
  OAI222_X1 U9301 ( .A1(n10294), .A2(n9827), .B1(n10292), .B2(n7686), .C1(
        P1_U3084), .C2(n10389), .ZN(P1_U3335) );
  NOR2_X1 U9302 ( .A1(n9188), .A2(n7687), .ZN(n7691) );
  NAND2_X1 U9303 ( .A1(n4392), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n7688) );
  OAI21_X1 U9304 ( .B1(n7689), .B2(n4392), .A(n7688), .ZN(n7690) );
  AOI211_X1 U9305 ( .C1(n9158), .C2(n7692), .A(n7691), .B(n7690), .ZN(n7695)
         );
  AOI22_X1 U9306 ( .A1(n9056), .A2(n7693), .B1(n9190), .B2(n8800), .ZN(n7694)
         );
  NAND2_X1 U9307 ( .A1(n7695), .A2(n7694), .ZN(P2_U3294) );
  AND2_X1 U9308 ( .A1(n7697), .A2(n7696), .ZN(n7700) );
  INV_X1 U9309 ( .A(n7700), .ZN(n10570) );
  NOR2_X1 U9310 ( .A1(n6911), .A2(n9205), .ZN(n7698) );
  AOI21_X1 U9311 ( .B1(n10570), .B2(n9225), .A(n7698), .ZN(n10571) );
  INV_X1 U9312 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n7699) );
  OAI22_X1 U9313 ( .A1(n4392), .A2(n10571), .B1(n7699), .B2(n9188), .ZN(n7702)
         );
  NOR2_X1 U9314 ( .A1(n9231), .A2(n7700), .ZN(n7701) );
  AOI211_X1 U9315 ( .C1(n4392), .C2(P2_REG2_REG_0__SCAN_IN), .A(n7702), .B(
        n7701), .ZN(n7704) );
  OAI21_X1 U9316 ( .B1(n9234), .B2(n9190), .A(n10569), .ZN(n7703) );
  NAND2_X1 U9317 ( .A1(n7704), .A2(n7703), .ZN(P2_U3296) );
  INV_X1 U9318 ( .A(n7705), .ZN(n7708) );
  OAI222_X1 U9319 ( .A1(n9395), .A2(n7707), .B1(n9399), .B2(n7708), .C1(
        P2_U3152), .C2(n7706), .ZN(P2_U3339) );
  OAI222_X1 U9320 ( .A1(n10294), .A2(n7709), .B1(n10292), .B2(n7708), .C1(
        P1_U3084), .C2(n9733), .ZN(P1_U3334) );
  XNOR2_X1 U9321 ( .A(n7710), .B(n7776), .ZN(n10577) );
  INV_X1 U9322 ( .A(n10577), .ZN(n7725) );
  NAND2_X1 U9323 ( .A1(n7713), .A2(n7712), .ZN(n7714) );
  XNOR2_X1 U9324 ( .A(n7714), .B(n7776), .ZN(n7717) );
  OAI22_X1 U9325 ( .A1(n7716), .A2(n9205), .B1(n7715), .B2(n9203), .ZN(n8730)
         );
  AOI21_X1 U9326 ( .B1(n7717), .B2(n9225), .A(n8730), .ZN(n10574) );
  MUX2_X1 U9327 ( .A(n10574), .B(n9825), .S(n4392), .Z(n7724) );
  INV_X1 U9328 ( .A(n7718), .ZN(n9158) );
  OAI21_X1 U9329 ( .B1(n7719), .B2(n10575), .A(n9357), .ZN(n7720) );
  OR2_X1 U9330 ( .A1(n7720), .A2(n7782), .ZN(n10573) );
  INV_X1 U9331 ( .A(n8731), .ZN(n7721) );
  OAI22_X1 U9332 ( .A1(n7718), .A2(n10573), .B1(n7721), .B2(n9188), .ZN(n7722)
         );
  AOI21_X1 U9333 ( .B1(n9190), .B2(n6717), .A(n7722), .ZN(n7723) );
  OAI211_X1 U9334 ( .C1(n7725), .C2(n9231), .A(n7724), .B(n7723), .ZN(P2_U3291) );
  AOI22_X1 U9335 ( .A1(n7924), .A2(n8592), .B1(n9587), .B2(n6956), .ZN(n7726)
         );
  XNOR2_X1 U9336 ( .A(n7726), .B(n8476), .ZN(n7857) );
  AOI22_X1 U9337 ( .A1(n8496), .A2(n9587), .B1(n7924), .B2(n6956), .ZN(n7856)
         );
  XNOR2_X1 U9338 ( .A(n7857), .B(n7856), .ZN(n7738) );
  NAND2_X1 U9339 ( .A1(n7728), .A2(n7727), .ZN(n7733) );
  INV_X1 U9340 ( .A(n7729), .ZN(n7731) );
  NAND2_X1 U9341 ( .A1(n7731), .A2(n7730), .ZN(n7732) );
  NAND2_X1 U9342 ( .A1(n7733), .A2(n7732), .ZN(n7737) );
  INV_X1 U9343 ( .A(n7737), .ZN(n7735) );
  INV_X1 U9344 ( .A(n7859), .ZN(n7736) );
  AOI211_X1 U9345 ( .C1(n7738), .C2(n7737), .A(n9520), .B(n7736), .ZN(n7745)
         );
  NAND2_X1 U9346 ( .A1(n9553), .A2(n9588), .ZN(n7740) );
  OAI211_X1 U9347 ( .C1(n7741), .C2(n9555), .A(n7740), .B(n7739), .ZN(n7744)
         );
  INV_X1 U9348 ( .A(n7923), .ZN(n7742) );
  INV_X1 U9349 ( .A(n9532), .ZN(n9452) );
  NAND2_X1 U9350 ( .A1(n7924), .A2(n10240), .ZN(n10446) );
  OAI22_X1 U9351 ( .A1(n9542), .A2(n7742), .B1(n9452), .B2(n10446), .ZN(n7743)
         );
  OR3_X1 U9352 ( .A1(n7745), .A2(n7744), .A3(n7743), .ZN(P1_U3228) );
  INV_X1 U9353 ( .A(n7746), .ZN(n7749) );
  NOR3_X1 U9354 ( .A1(n8793), .A2(n8046), .A3(n7747), .ZN(n7748) );
  AOI21_X1 U9355 ( .B1(n7749), .B2(n6894), .A(n7748), .ZN(n7758) );
  INV_X1 U9356 ( .A(n7750), .ZN(n7755) );
  INV_X1 U9357 ( .A(n9355), .ZN(n8056) );
  OAI22_X1 U9358 ( .A1(n8786), .A2(n8046), .B1(n8695), .B2(n8056), .ZN(n7754)
         );
  NAND2_X1 U9359 ( .A1(n8761), .A2(n8053), .ZN(n7751) );
  OAI211_X1 U9360 ( .C1(n8785), .C2(n8115), .A(n7752), .B(n7751), .ZN(n7753)
         );
  AOI211_X1 U9361 ( .C1(n7755), .C2(n6894), .A(n7754), .B(n7753), .ZN(n7756)
         );
  OAI21_X1 U9362 ( .B1(n7758), .B2(n7757), .A(n7756), .ZN(P2_U3233) );
  INV_X1 U9363 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n9747) );
  AOI22_X1 U9364 ( .A1(n8539), .A2(n9747), .B1(P2_REG1_REG_14__SCAN_IN), .B2(
        n8550), .ZN(n7762) );
  AOI21_X1 U9365 ( .B1(n7763), .B2(n7762), .A(n8549), .ZN(n7773) );
  NOR2_X1 U9366 ( .A1(n9890), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8659) );
  INV_X1 U9367 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n7764) );
  NOR2_X1 U9368 ( .A1(n8863), .A2(n7764), .ZN(n7765) );
  AOI211_X1 U9369 ( .C1(n8870), .C2(n8539), .A(n8659), .B(n7765), .ZN(n7772)
         );
  INV_X1 U9370 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n9817) );
  AOI22_X1 U9371 ( .A1(n8539), .A2(P2_REG2_REG_14__SCAN_IN), .B1(n9817), .B2(
        n8550), .ZN(n7769) );
  OAI21_X1 U9372 ( .B1(n7769), .B2(n7768), .A(n8538), .ZN(n7770) );
  NAND2_X1 U9373 ( .A1(n7770), .A2(n10506), .ZN(n7771) );
  OAI211_X1 U9374 ( .C1(n7773), .C2(n10510), .A(n7772), .B(n7771), .ZN(
        P2_U3259) );
  INV_X1 U9375 ( .A(n7774), .ZN(n7807) );
  OAI222_X1 U9376 ( .A1(n9399), .A2(n7807), .B1(n4396), .B2(P2_U3152), .C1(
        n9948), .C2(n9395), .ZN(P2_U3338) );
  AOI21_X1 U9377 ( .B1(n7710), .B2(n7776), .A(n7775), .ZN(n7777) );
  XNOR2_X1 U9378 ( .A(n7777), .B(n7779), .ZN(n10584) );
  INV_X1 U9379 ( .A(n10584), .ZN(n7789) );
  XOR2_X1 U9380 ( .A(n7778), .B(n7779), .Z(n7780) );
  OAI222_X1 U9381 ( .A1(n9205), .A2(n8690), .B1(n9203), .B2(n7781), .C1(n9200), 
        .C2(n7780), .ZN(n10581) );
  OAI21_X1 U9382 ( .B1(n7782), .B2(n10579), .A(n7810), .ZN(n10580) );
  NAND2_X1 U9383 ( .A1(n9190), .A2(n7783), .ZN(n7786) );
  AOI22_X1 U9384 ( .A1(n4392), .A2(P2_REG2_REG_6__SCAN_IN), .B1(n7784), .B2(
        n10517), .ZN(n7785) );
  OAI211_X1 U9385 ( .C1(n10580), .C2(n8974), .A(n7786), .B(n7785), .ZN(n7787)
         );
  AOI21_X1 U9386 ( .B1(n10581), .B2(n9060), .A(n7787), .ZN(n7788) );
  OAI21_X1 U9387 ( .B1(n9231), .B2(n7789), .A(n7788), .ZN(P2_U3290) );
  INV_X1 U9388 ( .A(n10442), .ZN(n7805) );
  NOR2_X1 U9389 ( .A1(n7791), .A2(n7930), .ZN(n7792) );
  NAND2_X1 U9390 ( .A1(n10148), .A2(n7792), .ZN(n7892) );
  OAI211_X1 U9391 ( .C1(n6054), .C2(n7794), .A(n10418), .B(n7793), .ZN(n10437)
         );
  AOI222_X1 U9392 ( .A1(n7797), .A2(n10101), .B1(n10482), .B2(n10442), .C1(
        n9589), .C2(n8217), .ZN(n10439) );
  INV_X1 U9393 ( .A(n10145), .ZN(n10411) );
  NOR2_X1 U9394 ( .A1(n7798), .A2(n10403), .ZN(n10436) );
  AOI21_X1 U9395 ( .B1(n10411), .B2(P1_REG3_REG_1__SCAN_IN), .A(n10436), .ZN(
        n7799) );
  OAI211_X1 U9396 ( .C1(n9632), .C2(n10437), .A(n10439), .B(n7799), .ZN(n7800)
         );
  NAND2_X1 U9397 ( .A1(n7800), .A2(n10148), .ZN(n7804) );
  AOI22_X1 U9398 ( .A1(n10150), .A2(n7802), .B1(n10123), .B2(
        P1_REG2_REG_1__SCAN_IN), .ZN(n7803) );
  OAI211_X1 U9399 ( .C1(n7805), .C2(n7892), .A(n7804), .B(n7803), .ZN(P1_U3290) );
  OAI222_X1 U9400 ( .A1(n10294), .A2(n7808), .B1(n10292), .B2(n7807), .C1(
        n7806), .C2(P1_U3084), .ZN(P1_U3333) );
  XOR2_X1 U9401 ( .A(n7809), .B(n7817), .Z(n7828) );
  NAND2_X1 U9402 ( .A1(n7810), .A2(n7824), .ZN(n7811) );
  AND2_X1 U9403 ( .A1(n7812), .A2(n7811), .ZN(n7825) );
  INV_X1 U9404 ( .A(n7825), .ZN(n7815) );
  AOI22_X1 U9405 ( .A1(n4392), .A2(P2_REG2_REG_7__SCAN_IN), .B1(n7813), .B2(
        n10517), .ZN(n7814) );
  OAI21_X1 U9406 ( .B1(n8974), .B2(n7815), .A(n7814), .ZN(n7822) );
  OAI211_X1 U9407 ( .C1(n7818), .C2(n7817), .A(n7816), .B(n9225), .ZN(n7820)
         );
  AOI22_X1 U9408 ( .A1(n9220), .A2(n8840), .B1(n8838), .B2(n9222), .ZN(n7819)
         );
  AND2_X1 U9409 ( .A1(n7820), .A2(n7819), .ZN(n7827) );
  NOR2_X1 U9410 ( .A1(n7827), .A2(n4392), .ZN(n7821) );
  AOI211_X1 U9411 ( .C1(n9190), .C2(n7824), .A(n7822), .B(n7821), .ZN(n7823)
         );
  OAI21_X1 U9412 ( .B1(n9231), .B2(n7828), .A(n7823), .ZN(P2_U3289) );
  AOI22_X1 U9413 ( .A1(n7825), .A2(n9357), .B1(n9356), .B2(n7824), .ZN(n7826)
         );
  OAI211_X1 U9414 ( .C1(n7828), .C2(n9350), .A(n7827), .B(n7826), .ZN(n7831)
         );
  NAND2_X1 U9415 ( .A1(n7831), .A2(n10605), .ZN(n7829) );
  OAI21_X1 U9416 ( .B1(n10605), .B2(n7830), .A(n7829), .ZN(P2_U3527) );
  INV_X1 U9417 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n7833) );
  NAND2_X1 U9418 ( .A1(n7831), .A2(n10598), .ZN(n7832) );
  OAI21_X1 U9419 ( .B1(n10598), .B2(n7833), .A(n7832), .ZN(P2_U3472) );
  INV_X1 U9420 ( .A(n7892), .ZN(n7951) );
  NAND2_X1 U9421 ( .A1(n7834), .A2(n7842), .ZN(n7835) );
  NAND2_X1 U9422 ( .A1(n7836), .A2(n7835), .ZN(n10464) );
  INV_X1 U9423 ( .A(n7837), .ZN(n7838) );
  OAI211_X1 U9424 ( .C1(n7867), .C2(n10417), .A(n7838), .B(n10418), .ZN(n10461) );
  INV_X1 U9425 ( .A(n7839), .ZN(n7840) );
  NAND2_X1 U9426 ( .A1(n7840), .A2(n9733), .ZN(n9659) );
  AOI22_X1 U9427 ( .A1(n10150), .A2(n9531), .B1(n10411), .B2(n9533), .ZN(n7841) );
  OAI21_X1 U9428 ( .B1(n10461), .B2(n9659), .A(n7841), .ZN(n7848) );
  XNOR2_X1 U9429 ( .A(n7843), .B(n7842), .ZN(n7846) );
  NAND2_X1 U9430 ( .A1(n10464), .A2(n10482), .ZN(n7845) );
  AOI22_X1 U9431 ( .A1(n4756), .A2(n8217), .B1(n10103), .B2(n9586), .ZN(n7844)
         );
  OAI211_X1 U9432 ( .C1(n10406), .C2(n7846), .A(n7845), .B(n7844), .ZN(n10462)
         );
  MUX2_X1 U9433 ( .A(n10462), .B(P1_REG2_REG_6__SCAN_IN), .S(n10123), .Z(n7847) );
  AOI211_X1 U9434 ( .C1(n7951), .C2(n10464), .A(n7848), .B(n7847), .ZN(n7849)
         );
  INV_X1 U9435 ( .A(n7849), .ZN(P1_U3285) );
  NAND2_X1 U9436 ( .A1(n7894), .A2(n8592), .ZN(n7852) );
  OR2_X1 U9437 ( .A1(n7850), .A2(n8593), .ZN(n7851) );
  NAND2_X1 U9438 ( .A1(n7852), .A2(n7851), .ZN(n7853) );
  XNOR2_X1 U9439 ( .A(n7853), .B(n8476), .ZN(n7996) );
  NAND2_X1 U9440 ( .A1(n4756), .A2(n8496), .ZN(n7855) );
  NAND2_X1 U9441 ( .A1(n7894), .A2(n6956), .ZN(n7854) );
  AND2_X1 U9442 ( .A1(n7855), .A2(n7854), .ZN(n7997) );
  XNOR2_X1 U9443 ( .A(n7996), .B(n7997), .ZN(n7877) );
  OR2_X1 U9444 ( .A1(n7857), .A2(n7856), .ZN(n7858) );
  NAND2_X1 U9445 ( .A1(n8496), .A2(n9586), .ZN(n7861) );
  OR2_X1 U9446 ( .A1(n10421), .A2(n8593), .ZN(n7860) );
  NAND2_X1 U9447 ( .A1(n7861), .A2(n7860), .ZN(n7954) );
  NAND2_X1 U9448 ( .A1(n9586), .A2(n6956), .ZN(n7862) );
  OAI21_X1 U9449 ( .B1(n10421), .B2(n7865), .A(n7862), .ZN(n7863) );
  XNOR2_X1 U9450 ( .A(n7863), .B(n8476), .ZN(n7871) );
  NAND2_X1 U9451 ( .A1(n9585), .A2(n6956), .ZN(n7864) );
  OAI21_X1 U9452 ( .B1(n7867), .B2(n7865), .A(n7864), .ZN(n7866) );
  XNOR2_X1 U9453 ( .A(n8476), .B(n7866), .ZN(n9526) );
  NAND2_X1 U9454 ( .A1(n8496), .A2(n9585), .ZN(n7869) );
  OR2_X1 U9455 ( .A1(n7867), .A2(n8593), .ZN(n7868) );
  NAND2_X1 U9456 ( .A1(n7869), .A2(n7868), .ZN(n9525) );
  AOI22_X1 U9457 ( .A1(n7954), .A2(n7871), .B1(n9526), .B2(n9525), .ZN(n7870)
         );
  OAI21_X1 U9458 ( .B1(n7871), .B2(n7954), .A(n9525), .ZN(n7874) );
  INV_X1 U9459 ( .A(n9526), .ZN(n7873) );
  INV_X1 U9460 ( .A(n7871), .ZN(n9524) );
  NOR2_X1 U9461 ( .A1(n7954), .A2(n9525), .ZN(n7872) );
  AOI22_X1 U9462 ( .A1(n7874), .A2(n7873), .B1(n9524), .B2(n7872), .ZN(n7875)
         );
  OAI21_X1 U9463 ( .B1(n7877), .B2(n7876), .A(n8000), .ZN(n7885) );
  AOI21_X1 U9464 ( .B1(n9553), .B2(n9585), .A(n7878), .ZN(n7883) );
  NAND2_X1 U9465 ( .A1(n7894), .A2(n10240), .ZN(n10467) );
  INV_X1 U9466 ( .A(n10467), .ZN(n7879) );
  NAND2_X1 U9467 ( .A1(n9532), .A2(n7879), .ZN(n7882) );
  NAND2_X1 U9468 ( .A1(n9560), .A2(n7893), .ZN(n7881) );
  NAND2_X1 U9469 ( .A1(n9534), .A2(n9584), .ZN(n7880) );
  NAND4_X1 U9470 ( .A1(n7883), .A2(n7882), .A3(n7881), .A4(n7880), .ZN(n7884)
         );
  AOI21_X1 U9471 ( .B1(n7885), .B2(n9547), .A(n7884), .ZN(n7886) );
  INV_X1 U9472 ( .A(n7886), .ZN(P1_U3211) );
  XNOR2_X1 U9473 ( .A(n7887), .B(n7889), .ZN(n7888) );
  AOI222_X1 U9474 ( .A1(n7888), .A2(n10101), .B1(n9585), .B2(n10103), .C1(
        n9584), .C2(n8217), .ZN(n10469) );
  MUX2_X1 U9475 ( .A(n9859), .B(n10469), .S(n10148), .Z(n7898) );
  XNOR2_X1 U9476 ( .A(n7890), .B(n7889), .ZN(n10471) );
  NAND2_X1 U9477 ( .A1(n10148), .A2(n10482), .ZN(n7891) );
  OAI211_X1 U9478 ( .C1(n7837), .C2(n4758), .A(n10418), .B(n7965), .ZN(n10468)
         );
  AOI22_X1 U9479 ( .A1(n10150), .A2(n7894), .B1(n7893), .B2(n10411), .ZN(n7895) );
  OAI21_X1 U9480 ( .B1(n10468), .B2(n9659), .A(n7895), .ZN(n7896) );
  AOI21_X1 U9481 ( .B1(n10471), .B2(n10424), .A(n7896), .ZN(n7897) );
  NAND2_X1 U9482 ( .A1(n7898), .A2(n7897), .ZN(P1_U3284) );
  INV_X1 U9483 ( .A(n7899), .ZN(n7901) );
  OAI21_X1 U9484 ( .B1(n7963), .B2(n7901), .A(n7900), .ZN(n7902) );
  XOR2_X1 U9485 ( .A(n7905), .B(n7902), .Z(n7903) );
  OAI222_X1 U9486 ( .A1(n10405), .A2(n8207), .B1(n10403), .B2(n8008), .C1(
        n7903), .C2(n10406), .ZN(n10486) );
  INV_X1 U9487 ( .A(n10486), .ZN(n7912) );
  OAI21_X1 U9488 ( .B1(n7906), .B2(n7905), .A(n7904), .ZN(n10488) );
  OAI211_X1 U9489 ( .C1(n7907), .C2(n6056), .A(n10418), .B(n8061), .ZN(n10484)
         );
  AOI22_X1 U9490 ( .A1(n10123), .A2(P1_REG2_REG_9__SCAN_IN), .B1(n8162), .B2(
        n10411), .ZN(n7909) );
  NAND2_X1 U9491 ( .A1(n10150), .A2(n8163), .ZN(n7908) );
  OAI211_X1 U9492 ( .C1(n10484), .C2(n9659), .A(n7909), .B(n7908), .ZN(n7910)
         );
  AOI21_X1 U9493 ( .B1(n10488), .B2(n10424), .A(n7910), .ZN(n7911) );
  OAI21_X1 U9494 ( .B1(n7912), .B2(n10123), .A(n7911), .ZN(P1_U3282) );
  NAND2_X1 U9495 ( .A1(n7914), .A2(n7913), .ZN(n7915) );
  XNOR2_X1 U9496 ( .A(n7920), .B(n7915), .ZN(n7916) );
  NAND2_X1 U9497 ( .A1(n7916), .A2(n10101), .ZN(n7918) );
  AOI22_X1 U9498 ( .A1(n10103), .A2(n9588), .B1(n9586), .B2(n8217), .ZN(n7917)
         );
  AND2_X1 U9499 ( .A1(n7918), .A2(n7917), .ZN(n10451) );
  XNOR2_X1 U9500 ( .A(n7919), .B(n7920), .ZN(n10449) );
  AOI21_X1 U9501 ( .B1(n7921), .B2(n7924), .A(n10158), .ZN(n7922) );
  NAND2_X1 U9502 ( .A1(n7922), .A2(n10416), .ZN(n10447) );
  AOI22_X1 U9503 ( .A1(n10123), .A2(P1_REG2_REG_4__SCAN_IN), .B1(n7923), .B2(
        n10411), .ZN(n7926) );
  NAND2_X1 U9504 ( .A1(n10150), .A2(n7924), .ZN(n7925) );
  OAI211_X1 U9505 ( .C1(n10447), .C2(n9659), .A(n7926), .B(n7925), .ZN(n7927)
         );
  AOI21_X1 U9506 ( .B1(n10449), .B2(n10424), .A(n7927), .ZN(n7928) );
  OAI21_X1 U9507 ( .B1(n10451), .B2(n10123), .A(n7928), .ZN(P1_U3287) );
  INV_X1 U9508 ( .A(n7929), .ZN(n8534) );
  OAI222_X1 U9509 ( .A1(n10294), .A2(n9929), .B1(n10283), .B2(n8534), .C1(
        n7930), .C2(P1_U3084), .ZN(P1_U3332) );
  INV_X1 U9510 ( .A(n7932), .ZN(n7933) );
  AOI21_X1 U9511 ( .B1(n7931), .B2(n7933), .A(n8821), .ZN(n7937) );
  NOR3_X1 U9512 ( .A1(n8793), .A2(n8115), .A3(n7934), .ZN(n7936) );
  OAI21_X1 U9513 ( .B1(n7937), .B2(n7936), .A(n7935), .ZN(n7942) );
  INV_X1 U9514 ( .A(n8121), .ZN(n7938) );
  OAI22_X1 U9515 ( .A1(n8818), .A2(n7938), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n6260), .ZN(n7940) );
  OAI22_X1 U9516 ( .A1(n8115), .A2(n8786), .B1(n8785), .B2(n8304), .ZN(n7939)
         );
  AOI211_X1 U9517 ( .C1(n9347), .C2(n8825), .A(n7940), .B(n7939), .ZN(n7941)
         );
  NAND2_X1 U9518 ( .A1(n7942), .A2(n7941), .ZN(P2_U3238) );
  INV_X1 U9519 ( .A(n7943), .ZN(n7944) );
  AOI22_X1 U9520 ( .A1(n10422), .A2(n7944), .B1(P1_REG3_REG_2__SCAN_IN), .B2(
        n10411), .ZN(n7945) );
  OAI21_X1 U9521 ( .B1(n10400), .B2(n4391), .A(n7945), .ZN(n7949) );
  MUX2_X1 U9522 ( .A(P1_REG2_REG_2__SCAN_IN), .B(n7947), .S(n10148), .Z(n7948)
         );
  AOI211_X1 U9523 ( .C1(n7951), .C2(n7950), .A(n7949), .B(n7948), .ZN(n7952)
         );
  INV_X1 U9524 ( .A(n7952), .ZN(P1_U3289) );
  XNOR2_X1 U9525 ( .A(n9523), .B(n9524), .ZN(n7953) );
  NOR2_X1 U9526 ( .A1(n7953), .A2(n7954), .ZN(n9522) );
  AOI21_X1 U9527 ( .B1(n7954), .B2(n7953), .A(n9522), .ZN(n7960) );
  OR2_X1 U9528 ( .A1(n10485), .A2(n10421), .ZN(n10453) );
  NOR2_X1 U9529 ( .A1(n9452), .A2(n10453), .ZN(n7958) );
  NAND2_X1 U9530 ( .A1(P1_U3084), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n9600) );
  INV_X1 U9531 ( .A(n9600), .ZN(n7955) );
  AOI21_X1 U9532 ( .B1(n9553), .B2(n9587), .A(n7955), .ZN(n7956) );
  OAI21_X1 U9533 ( .B1(n10404), .B2(n9555), .A(n7956), .ZN(n7957) );
  AOI211_X1 U9534 ( .C1(n10410), .C2(n9560), .A(n7958), .B(n7957), .ZN(n7959)
         );
  OAI21_X1 U9535 ( .B1(n7960), .B2(n9520), .A(n7959), .ZN(P1_U3225) );
  XOR2_X1 U9536 ( .A(n7961), .B(n7962), .Z(n10481) );
  INV_X1 U9537 ( .A(n10481), .ZN(n10474) );
  XNOR2_X1 U9538 ( .A(n7963), .B(n7962), .ZN(n7964) );
  AOI222_X1 U9539 ( .A1(n9583), .A2(n8217), .B1(n10101), .B2(n7964), .C1(n4756), .C2(n10103), .ZN(n10477) );
  INV_X1 U9540 ( .A(n10477), .ZN(n7973) );
  AOI21_X1 U9541 ( .B1(n7965), .B2(n10475), .A(n10158), .ZN(n7967) );
  NAND2_X1 U9542 ( .A1(n7967), .A2(n7966), .ZN(n10476) );
  INV_X1 U9543 ( .A(n8235), .ZN(n7968) );
  OAI22_X1 U9544 ( .A1(n10148), .A2(n7969), .B1(n7968), .B2(n10145), .ZN(n7970) );
  AOI21_X1 U9545 ( .B1(n10150), .B2(n10475), .A(n7970), .ZN(n7971) );
  OAI21_X1 U9546 ( .B1(n10476), .B2(n9659), .A(n7971), .ZN(n7972) );
  AOI21_X1 U9547 ( .B1(n7973), .B2(n10148), .A(n7972), .ZN(n7974) );
  OAI21_X1 U9548 ( .B1(n10142), .B2(n10474), .A(n7974), .ZN(P1_U3283) );
  INV_X1 U9549 ( .A(n7975), .ZN(n7984) );
  INV_X1 U9550 ( .A(n7976), .ZN(n7977) );
  MUX2_X1 U9551 ( .A(n7978), .B(n7977), .S(n10148), .Z(n7983) );
  OAI22_X1 U9552 ( .A1(n10400), .A2(n7979), .B1(P1_REG3_REG_3__SCAN_IN), .B2(
        n10145), .ZN(n7980) );
  AOI21_X1 U9553 ( .B1(n10422), .B2(n7981), .A(n7980), .ZN(n7982) );
  OAI211_X1 U9554 ( .C1(n10142), .C2(n7984), .A(n7983), .B(n7982), .ZN(
        P1_U3288) );
  INV_X1 U9555 ( .A(n7931), .ZN(n7985) );
  AOI211_X1 U9556 ( .C1(n7987), .C2(n7986), .A(n8821), .B(n7985), .ZN(n7992)
         );
  OAI22_X1 U9557 ( .A1(n7988), .A2(n8786), .B1(n8785), .B2(n8088), .ZN(n7991)
         );
  INV_X1 U9558 ( .A(n8243), .ZN(n8101) );
  AOI22_X1 U9559 ( .A1(n8761), .A2(n8099), .B1(P2_REG3_REG_10__SCAN_IN), .B2(
        P2_U3152), .ZN(n7989) );
  OAI21_X1 U9560 ( .B1(n8101), .B2(n8695), .A(n7989), .ZN(n7990) );
  OR3_X1 U9561 ( .A1(n7992), .A2(n7991), .A3(n7990), .ZN(P2_U3219) );
  INV_X1 U9562 ( .A(n7993), .ZN(n8536) );
  OAI222_X1 U9563 ( .A1(n10294), .A2(n7995), .B1(n10292), .B2(n8536), .C1(
        P1_U3084), .C2(n7994), .ZN(P1_U3331) );
  INV_X1 U9564 ( .A(n7996), .ZN(n7998) );
  NAND2_X1 U9565 ( .A1(n7998), .A2(n7997), .ZN(n7999) );
  NAND2_X1 U9566 ( .A1(n8163), .A2(n8592), .ZN(n8002) );
  OR2_X1 U9567 ( .A1(n8026), .A2(n8593), .ZN(n8001) );
  NAND2_X1 U9568 ( .A1(n8002), .A2(n8001), .ZN(n8003) );
  XNOR2_X1 U9569 ( .A(n8003), .B(n8476), .ZN(n8156) );
  NAND2_X1 U9570 ( .A1(n8163), .A2(n4535), .ZN(n8005) );
  NAND2_X1 U9571 ( .A1(n9583), .A2(n8496), .ZN(n8004) );
  NAND2_X1 U9572 ( .A1(n8005), .A2(n8004), .ZN(n8155) );
  NAND2_X1 U9573 ( .A1(n10475), .A2(n4535), .ZN(n8007) );
  NAND2_X1 U9574 ( .A1(n9584), .A2(n8496), .ZN(n8006) );
  NAND2_X1 U9575 ( .A1(n8007), .A2(n8006), .ZN(n8153) );
  NAND2_X1 U9576 ( .A1(n10475), .A2(n8592), .ZN(n8010) );
  OR2_X1 U9577 ( .A1(n8008), .A2(n8593), .ZN(n8009) );
  NAND2_X1 U9578 ( .A1(n8010), .A2(n8009), .ZN(n8011) );
  XNOR2_X1 U9579 ( .A(n8011), .B(n8476), .ZN(n8231) );
  AOI22_X1 U9580 ( .A1(n8156), .A2(n8155), .B1(n8153), .B2(n8231), .ZN(n8012)
         );
  NAND2_X1 U9581 ( .A1(n8152), .A2(n8012), .ZN(n8018) );
  INV_X1 U9582 ( .A(n8156), .ZN(n8016) );
  OAI21_X1 U9583 ( .B1(n8231), .B2(n8153), .A(n8155), .ZN(n8015) );
  NOR2_X1 U9584 ( .A1(n8155), .A2(n8153), .ZN(n8014) );
  INV_X1 U9585 ( .A(n8231), .ZN(n8013) );
  AOI22_X1 U9586 ( .A1(n8016), .A2(n8015), .B1(n8014), .B2(n8013), .ZN(n8017)
         );
  NAND2_X1 U9587 ( .A1(n8066), .A2(n8592), .ZN(n8020) );
  OR2_X1 U9588 ( .A1(n8207), .A2(n8593), .ZN(n8019) );
  NAND2_X1 U9589 ( .A1(n8020), .A2(n8019), .ZN(n8021) );
  XNOR2_X1 U9590 ( .A(n8021), .B(n8563), .ZN(n8195) );
  NOR2_X1 U9591 ( .A1(n8207), .A2(n8599), .ZN(n8022) );
  AOI21_X1 U9592 ( .B1(n8066), .B2(n6956), .A(n8022), .ZN(n8196) );
  XNOR2_X1 U9593 ( .A(n8195), .B(n8196), .ZN(n8023) );
  XNOR2_X1 U9594 ( .A(n8193), .B(n8023), .ZN(n8031) );
  NAND2_X1 U9595 ( .A1(n9534), .A2(n9581), .ZN(n8025) );
  OAI211_X1 U9596 ( .C1(n8026), .C2(n9494), .A(n8025), .B(n8024), .ZN(n8029)
         );
  INV_X1 U9597 ( .A(n8027), .ZN(n8063) );
  NOR2_X1 U9598 ( .A1(n9542), .A2(n8063), .ZN(n8028) );
  AOI211_X1 U9599 ( .C1(n9518), .C2(n8066), .A(n8029), .B(n8028), .ZN(n8030)
         );
  OAI21_X1 U9600 ( .B1(n8031), .B2(n9520), .A(n8030), .ZN(P1_U3215) );
  NAND2_X1 U9601 ( .A1(n8169), .A2(n8032), .ZN(n8134) );
  XNOR2_X1 U9602 ( .A(n8134), .B(n8035), .ZN(n10242) );
  NAND2_X1 U9603 ( .A1(n8034), .A2(n8035), .ZN(n8140) );
  OAI211_X1 U9604 ( .C1(n8035), .C2(n8034), .A(n8140), .B(n10101), .ZN(n8037)
         );
  OR2_X1 U9605 ( .A1(n8264), .A2(n10405), .ZN(n8036) );
  OAI211_X1 U9606 ( .C1(n8207), .C2(n10403), .A(n8037), .B(n8036), .ZN(n10237)
         );
  INV_X1 U9607 ( .A(n8146), .ZN(n8038) );
  AOI211_X1 U9608 ( .C1(n10239), .C2(n4902), .A(n10158), .B(n8038), .ZN(n10238) );
  NAND2_X1 U9609 ( .A1(n10238), .A2(n10422), .ZN(n8040) );
  AOI22_X1 U9610 ( .A1(n10123), .A2(P1_REG2_REG_11__SCAN_IN), .B1(n8211), .B2(
        n10411), .ZN(n8039) );
  OAI211_X1 U9611 ( .C1(n8208), .C2(n10400), .A(n8040), .B(n8039), .ZN(n8041)
         );
  AOI21_X1 U9612 ( .B1(n10237), .B2(n10148), .A(n8041), .ZN(n8042) );
  OAI21_X1 U9613 ( .B1(n10242), .B2(n10142), .A(n8042), .ZN(P1_U3280) );
  AND2_X1 U9614 ( .A1(n8112), .A2(n8043), .ZN(n8045) );
  NAND2_X1 U9615 ( .A1(n8047), .A2(n8043), .ZN(n8106) );
  INV_X1 U9616 ( .A(n8106), .ZN(n8044) );
  NAND2_X1 U9617 ( .A1(n8112), .A2(n8044), .ZN(n8084) );
  OAI21_X1 U9618 ( .B1(n8045), .B2(n8047), .A(n8084), .ZN(n9354) );
  OAI22_X1 U9619 ( .A1(n8046), .A2(n9203), .B1(n8115), .B2(n9205), .ZN(n8051)
         );
  XNOR2_X1 U9620 ( .A(n8048), .B(n8047), .ZN(n8049) );
  NOR2_X1 U9621 ( .A1(n8049), .A2(n9200), .ZN(n8050) );
  AOI211_X1 U9622 ( .C1(n8086), .C2(n9354), .A(n8051), .B(n8050), .ZN(n9360)
         );
  NOR2_X2 U9623 ( .A1(n8052), .A2(n9355), .ZN(n8097) );
  AOI21_X1 U9624 ( .B1(n9355), .B2(n8052), .A(n8097), .ZN(n9358) );
  NAND2_X1 U9625 ( .A1(n9358), .A2(n9234), .ZN(n8055) );
  AOI22_X1 U9626 ( .A1(n4392), .A2(P2_REG2_REG_9__SCAN_IN), .B1(n8053), .B2(
        n10517), .ZN(n8054) );
  OAI211_X1 U9627 ( .C1(n8056), .C2(n10523), .A(n8055), .B(n8054), .ZN(n8057)
         );
  AOI21_X1 U9628 ( .B1(n9354), .B2(n10519), .A(n8057), .ZN(n8058) );
  OAI21_X1 U9629 ( .B1(n9360), .B2(n4392), .A(n8058), .ZN(P2_U3287) );
  XNOR2_X1 U9630 ( .A(n8060), .B(n8059), .ZN(n10300) );
  AOI21_X1 U9631 ( .B1(n8061), .B2(n8066), .A(n10158), .ZN(n8062) );
  NAND2_X1 U9632 ( .A1(n4902), .A2(n8062), .ZN(n10297) );
  OAI22_X1 U9633 ( .A1(n10148), .A2(n8064), .B1(n8063), .B2(n10145), .ZN(n8065) );
  AOI21_X1 U9634 ( .B1(n10150), .B2(n8066), .A(n8065), .ZN(n8067) );
  OAI21_X1 U9635 ( .B1(n10297), .B2(n9659), .A(n8067), .ZN(n8072) );
  XNOR2_X1 U9636 ( .A(n8069), .B(n8068), .ZN(n8070) );
  AOI222_X1 U9637 ( .A1(n9581), .A2(n8217), .B1(n10101), .B2(n8070), .C1(n9583), .C2(n10103), .ZN(n10298) );
  NOR2_X1 U9638 ( .A1(n10298), .A2(n10123), .ZN(n8071) );
  AOI211_X1 U9639 ( .C1(n10424), .C2(n10300), .A(n8072), .B(n8071), .ZN(n8073)
         );
  INV_X1 U9640 ( .A(n8073), .ZN(P1_U3281) );
  NAND2_X1 U9641 ( .A1(n8075), .A2(n8074), .ZN(n8077) );
  XOR2_X1 U9642 ( .A(n8077), .B(n8076), .Z(n8083) );
  INV_X1 U9643 ( .A(n9227), .ZN(n8079) );
  OAI21_X1 U9644 ( .B1(n8818), .B2(n8079), .A(n8078), .ZN(n8081) );
  OAI22_X1 U9645 ( .A1(n8088), .A2(n8786), .B1(n8785), .B2(n9204), .ZN(n8080)
         );
  AOI211_X1 U9646 ( .C1(n9342), .C2(n8825), .A(n8081), .B(n8080), .ZN(n8082)
         );
  OAI21_X1 U9647 ( .B1(n8083), .B2(n8821), .A(n8082), .ZN(P2_U3226) );
  OR2_X1 U9648 ( .A1(n9355), .A2(n8837), .ZN(n8108) );
  NAND2_X1 U9649 ( .A1(n8084), .A2(n8108), .ZN(n8085) );
  XNOR2_X1 U9650 ( .A(n8109), .B(n8085), .ZN(n8087) );
  INV_X1 U9651 ( .A(n8087), .ZN(n8246) );
  NAND2_X1 U9652 ( .A1(n8087), .A2(n8086), .ZN(n8096) );
  INV_X1 U9653 ( .A(n8088), .ZN(n9221) );
  AOI22_X1 U9654 ( .A1(n9221), .A2(n9222), .B1(n9220), .B2(n8837), .ZN(n8095)
         );
  NAND2_X1 U9655 ( .A1(n8090), .A2(n8089), .ZN(n8091) );
  NAND2_X1 U9656 ( .A1(n8091), .A2(n8109), .ZN(n8092) );
  NAND3_X1 U9657 ( .A1(n8093), .A2(n9225), .A3(n8092), .ZN(n8094) );
  NAND3_X1 U9658 ( .A1(n8096), .A2(n8095), .A3(n8094), .ZN(n8248) );
  NAND2_X1 U9659 ( .A1(n8248), .A2(n9060), .ZN(n8104) );
  OR2_X1 U9660 ( .A1(n8097), .A2(n8101), .ZN(n8098) );
  AND2_X1 U9661 ( .A1(n8098), .A2(n8119), .ZN(n8244) );
  AOI22_X1 U9662 ( .A1(n4392), .A2(P2_REG2_REG_10__SCAN_IN), .B1(n8099), .B2(
        n10517), .ZN(n8100) );
  OAI21_X1 U9663 ( .B1(n10523), .B2(n8101), .A(n8100), .ZN(n8102) );
  AOI21_X1 U9664 ( .B1(n8244), .B2(n9234), .A(n8102), .ZN(n8103) );
  OAI211_X1 U9665 ( .C1(n8246), .C2(n8105), .A(n8104), .B(n8103), .ZN(P2_U3286) );
  INV_X1 U9666 ( .A(n8115), .ZN(n8836) );
  AND2_X1 U9667 ( .A1(n8243), .A2(n8836), .ZN(n8107) );
  NOR2_X1 U9668 ( .A1(n8106), .A2(n8107), .ZN(n8111) );
  AOI21_X1 U9669 ( .B1(n8109), .B2(n8108), .A(n8107), .ZN(n8110) );
  XNOR2_X1 U9670 ( .A(n8291), .B(n8290), .ZN(n9351) );
  XNOR2_X1 U9671 ( .A(n8113), .B(n8290), .ZN(n8114) );
  NAND2_X1 U9672 ( .A1(n8114), .A2(n9225), .ZN(n8118) );
  OAI22_X1 U9673 ( .A1(n8304), .A2(n9205), .B1(n8115), .B2(n9203), .ZN(n8116)
         );
  INV_X1 U9674 ( .A(n8116), .ZN(n8117) );
  NAND2_X1 U9675 ( .A1(n8118), .A2(n8117), .ZN(n9353) );
  NAND2_X1 U9676 ( .A1(n9353), .A2(n9060), .ZN(n8126) );
  NAND2_X1 U9677 ( .A1(n8119), .A2(n9347), .ZN(n8120) );
  AND2_X1 U9678 ( .A1(n9226), .A2(n8120), .ZN(n9348) );
  INV_X1 U9679 ( .A(n9347), .ZN(n8123) );
  AOI22_X1 U9680 ( .A1(n4392), .A2(P2_REG2_REG_11__SCAN_IN), .B1(n8121), .B2(
        n10517), .ZN(n8122) );
  OAI21_X1 U9681 ( .B1(n10523), .B2(n8123), .A(n8122), .ZN(n8124) );
  AOI21_X1 U9682 ( .B1(n9348), .B2(n9234), .A(n8124), .ZN(n8125) );
  OAI211_X1 U9683 ( .C1(n9351), .C2(n9231), .A(n8126), .B(n8125), .ZN(P2_U3285) );
  INV_X1 U9684 ( .A(n8127), .ZN(n8132) );
  AOI21_X1 U9685 ( .B1(P1_DATAO_REG_23__SCAN_IN), .B2(n9388), .A(n8128), .ZN(
        n8129) );
  OAI21_X1 U9686 ( .B1(n8132), .B2(n9399), .A(n8129), .ZN(P2_U3335) );
  AOI21_X1 U9687 ( .B1(P2_DATAO_REG_23__SCAN_IN), .B2(n10281), .A(n8130), .ZN(
        n8131) );
  OAI21_X1 U9688 ( .B1(n8132), .B2(n10283), .A(n8131), .ZN(P1_U3330) );
  NOR2_X1 U9689 ( .A1(n10239), .A2(n9581), .ZN(n8133) );
  OAI21_X1 U9690 ( .B1(n8134), .B2(n8133), .A(n8167), .ZN(n8135) );
  XNOR2_X1 U9691 ( .A(n8135), .B(n8139), .ZN(n8351) );
  INV_X1 U9692 ( .A(n8351), .ZN(n8151) );
  NAND2_X1 U9693 ( .A1(n8140), .A2(n8138), .ZN(n8137) );
  INV_X1 U9694 ( .A(n8139), .ZN(n8136) );
  NAND2_X1 U9695 ( .A1(n8137), .A2(n8136), .ZN(n8142) );
  NAND3_X1 U9696 ( .A1(n8140), .A2(n8139), .A3(n8138), .ZN(n8141) );
  AOI21_X1 U9697 ( .B1(n8142), .B2(n8141), .A(n10406), .ZN(n8144) );
  OAI22_X1 U9698 ( .A1(n8202), .A2(n10403), .B1(n8327), .B2(n10405), .ZN(n8143) );
  OR2_X1 U9699 ( .A1(n8144), .A2(n8143), .ZN(n8349) );
  INV_X1 U9700 ( .A(n8329), .ZN(n8357) );
  INV_X1 U9701 ( .A(n8180), .ZN(n8145) );
  AOI211_X1 U9702 ( .C1(n8329), .C2(n8146), .A(n10158), .B(n8145), .ZN(n8350)
         );
  NAND2_X1 U9703 ( .A1(n8350), .A2(n10422), .ZN(n8148) );
  AOI22_X1 U9704 ( .A1(n10123), .A2(P1_REG2_REG_12__SCAN_IN), .B1(n8324), .B2(
        n10411), .ZN(n8147) );
  OAI211_X1 U9705 ( .C1(n8357), .C2(n10400), .A(n8148), .B(n8147), .ZN(n8149)
         );
  AOI21_X1 U9706 ( .B1(n8349), .B2(n10148), .A(n8149), .ZN(n8150) );
  OAI21_X1 U9707 ( .B1(n8151), .B2(n10142), .A(n8150), .ZN(P1_U3279) );
  INV_X1 U9708 ( .A(n8153), .ZN(n8154) );
  NAND2_X1 U9709 ( .A1(n8152), .A2(n8154), .ZN(n8229) );
  NOR2_X1 U9710 ( .A1(n8152), .A2(n8154), .ZN(n8228) );
  AOI21_X1 U9711 ( .B1(n8231), .B2(n8229), .A(n8228), .ZN(n8158) );
  XNOR2_X1 U9712 ( .A(n8156), .B(n8155), .ZN(n8157) );
  XNOR2_X1 U9713 ( .A(n8158), .B(n8157), .ZN(n8166) );
  NAND2_X1 U9714 ( .A1(n9553), .A2(n9584), .ZN(n8160) );
  OAI211_X1 U9715 ( .C1(n8207), .C2(n9555), .A(n8160), .B(n8159), .ZN(n8161)
         );
  AOI21_X1 U9716 ( .B1(n8162), .B2(n9560), .A(n8161), .ZN(n8165) );
  NAND2_X1 U9717 ( .A1(n9518), .A2(n8163), .ZN(n8164) );
  OAI211_X1 U9718 ( .C1(n8166), .C2(n9520), .A(n8165), .B(n8164), .ZN(P1_U3229) );
  INV_X1 U9719 ( .A(n8167), .ZN(n8168) );
  NOR2_X1 U9720 ( .A1(n8169), .A2(n8168), .ZN(n8172) );
  OAI21_X1 U9721 ( .B1(n8172), .B2(n8171), .A(n8170), .ZN(n8173) );
  XNOR2_X1 U9722 ( .A(n8173), .B(n8174), .ZN(n8360) );
  INV_X1 U9723 ( .A(n8360), .ZN(n8185) );
  XNOR2_X1 U9724 ( .A(n8175), .B(n8174), .ZN(n8176) );
  NAND2_X1 U9725 ( .A1(n8176), .A2(n10101), .ZN(n8179) );
  OAI22_X1 U9726 ( .A1(n8264), .A2(n10403), .B1(n8441), .B2(n10405), .ZN(n8177) );
  INV_X1 U9727 ( .A(n8177), .ZN(n8178) );
  NAND2_X1 U9728 ( .A1(n8179), .A2(n8178), .ZN(n8358) );
  INV_X1 U9729 ( .A(n8287), .ZN(n8365) );
  AOI211_X1 U9730 ( .C1(n8287), .C2(n8180), .A(n10158), .B(n8220), .ZN(n8359)
         );
  NAND2_X1 U9731 ( .A1(n8359), .A2(n10422), .ZN(n8182) );
  AOI22_X1 U9732 ( .A1(n10123), .A2(P1_REG2_REG_13__SCAN_IN), .B1(n8283), .B2(
        n10411), .ZN(n8181) );
  OAI211_X1 U9733 ( .C1(n8365), .C2(n10400), .A(n8182), .B(n8181), .ZN(n8183)
         );
  AOI21_X1 U9734 ( .B1(n10148), .B2(n8358), .A(n8183), .ZN(n8184) );
  OAI21_X1 U9735 ( .B1(n8185), .B2(n10142), .A(n8184), .ZN(P1_U3278) );
  XNOR2_X1 U9736 ( .A(n8186), .B(n8187), .ZN(n8192) );
  OAI22_X1 U9737 ( .A1(n8304), .A2(n8786), .B1(n8785), .B2(n8914), .ZN(n8188)
         );
  AOI211_X1 U9738 ( .C1(n8761), .C2(n8309), .A(n8189), .B(n8188), .ZN(n8191)
         );
  NAND2_X1 U9739 ( .A1(n8911), .A2(n8825), .ZN(n8190) );
  OAI211_X1 U9740 ( .C1(n8192), .C2(n8821), .A(n8191), .B(n8190), .ZN(P2_U3236) );
  INV_X1 U9741 ( .A(n8193), .ZN(n8194) );
  INV_X1 U9742 ( .A(n8195), .ZN(n8198) );
  INV_X1 U9743 ( .A(n8196), .ZN(n8197) );
  NAND2_X1 U9744 ( .A1(n8198), .A2(n8197), .ZN(n8260) );
  NAND2_X1 U9745 ( .A1(n8318), .A2(n8260), .ZN(n8204) );
  NAND2_X1 U9746 ( .A1(n10239), .A2(n8592), .ZN(n8200) );
  OR2_X1 U9747 ( .A1(n8202), .A2(n8593), .ZN(n8199) );
  NAND2_X1 U9748 ( .A1(n8200), .A2(n8199), .ZN(n8201) );
  XNOR2_X1 U9749 ( .A(n8201), .B(n8476), .ZN(n8259) );
  NOR2_X1 U9750 ( .A1(n8202), .A2(n8599), .ZN(n8203) );
  AOI21_X1 U9751 ( .B1(n10239), .B2(n6956), .A(n8203), .ZN(n8257) );
  XNOR2_X1 U9752 ( .A(n8259), .B(n8257), .ZN(n8271) );
  XNOR2_X1 U9753 ( .A(n8271), .B(n8204), .ZN(n8213) );
  NAND2_X1 U9754 ( .A1(n9534), .A2(n9580), .ZN(n8206) );
  OAI211_X1 U9755 ( .C1(n8207), .C2(n9494), .A(n8206), .B(n8205), .ZN(n8210)
         );
  NOR2_X1 U9756 ( .A1(n9556), .A2(n8208), .ZN(n8209) );
  AOI211_X1 U9757 ( .C1(n8211), .C2(n9560), .A(n8210), .B(n8209), .ZN(n8212)
         );
  OAI21_X1 U9758 ( .B1(n8213), .B2(n9520), .A(n8212), .ZN(P1_U3234) );
  XNOR2_X1 U9759 ( .A(n8214), .B(n8216), .ZN(n8397) );
  INV_X1 U9760 ( .A(n8397), .ZN(n8227) );
  NAND2_X1 U9761 ( .A1(n8215), .A2(n8216), .ZN(n8339) );
  OAI211_X1 U9762 ( .C1(n8215), .C2(n8216), .A(n8339), .B(n10101), .ZN(n8219)
         );
  NAND2_X1 U9763 ( .A1(n9577), .A2(n8217), .ZN(n8218) );
  OAI211_X1 U9764 ( .C1(n8327), .C2(n10403), .A(n8219), .B(n8218), .ZN(n8395)
         );
  INV_X1 U9765 ( .A(n8220), .ZN(n8222) );
  AOI211_X1 U9766 ( .C1(n8450), .C2(n8222), .A(n10158), .B(n8221), .ZN(n8396)
         );
  NAND2_X1 U9767 ( .A1(n8396), .A2(n10422), .ZN(n8224) );
  AOI22_X1 U9768 ( .A1(n10123), .A2(P1_REG2_REG_14__SCAN_IN), .B1(n9420), .B2(
        n10411), .ZN(n8223) );
  OAI211_X1 U9769 ( .C1(n9423), .C2(n10400), .A(n8224), .B(n8223), .ZN(n8225)
         );
  AOI21_X1 U9770 ( .B1(n10148), .B2(n8395), .A(n8225), .ZN(n8226) );
  OAI21_X1 U9771 ( .B1(n8227), .B2(n10142), .A(n8226), .ZN(P1_U3277) );
  INV_X1 U9772 ( .A(n8228), .ZN(n8230) );
  NAND2_X1 U9773 ( .A1(n8230), .A2(n8229), .ZN(n8232) );
  XNOR2_X1 U9774 ( .A(n8232), .B(n8231), .ZN(n8241) );
  INV_X1 U9775 ( .A(n8233), .ZN(n8234) );
  AOI21_X1 U9776 ( .B1(n9553), .B2(n4756), .A(n8234), .ZN(n8239) );
  NAND2_X1 U9777 ( .A1(n9518), .A2(n10475), .ZN(n8238) );
  NAND2_X1 U9778 ( .A1(n9560), .A2(n8235), .ZN(n8237) );
  NAND2_X1 U9779 ( .A1(n9534), .A2(n9583), .ZN(n8236) );
  NAND4_X1 U9780 ( .A1(n8239), .A2(n8238), .A3(n8237), .A4(n8236), .ZN(n8240)
         );
  AOI21_X1 U9781 ( .B1(n8241), .B2(n9547), .A(n8240), .ZN(n8242) );
  INV_X1 U9782 ( .A(n8242), .ZN(P1_U3219) );
  AOI22_X1 U9783 ( .A1(n8244), .A2(n9357), .B1(n9356), .B2(n8243), .ZN(n8245)
         );
  OAI21_X1 U9784 ( .B1(n8246), .B2(n10586), .A(n8245), .ZN(n8247) );
  NOR2_X1 U9785 ( .A1(n8248), .A2(n8247), .ZN(n8251) );
  MUX2_X1 U9786 ( .A(n8249), .B(n8251), .S(n10605), .Z(n8250) );
  INV_X1 U9787 ( .A(n8250), .ZN(P2_U3530) );
  INV_X1 U9788 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n8252) );
  MUX2_X1 U9789 ( .A(n8252), .B(n8251), .S(n10598), .Z(n8253) );
  INV_X1 U9790 ( .A(n8253), .ZN(P2_U3481) );
  INV_X1 U9791 ( .A(n8254), .ZN(n8333) );
  OAI222_X1 U9792 ( .A1(n9399), .A2(n8333), .B1(P2_U3152), .B2(n8256), .C1(
        n8255), .C2(n9395), .ZN(P2_U3334) );
  INV_X1 U9793 ( .A(n8257), .ZN(n8258) );
  NAND2_X1 U9794 ( .A1(n8259), .A2(n8258), .ZN(n8270) );
  AND2_X1 U9795 ( .A1(n8260), .A2(n8270), .ZN(n8317) );
  NAND2_X1 U9796 ( .A1(n8329), .A2(n8592), .ZN(n8262) );
  OR2_X1 U9797 ( .A1(n8264), .A2(n8593), .ZN(n8261) );
  NAND2_X1 U9798 ( .A1(n8262), .A2(n8261), .ZN(n8263) );
  XNOR2_X1 U9799 ( .A(n8263), .B(n8563), .ZN(n8269) );
  INV_X1 U9800 ( .A(n8269), .ZN(n8267) );
  NOR2_X1 U9801 ( .A1(n8264), .A2(n8599), .ZN(n8265) );
  AOI21_X1 U9802 ( .B1(n8329), .B2(n6956), .A(n8265), .ZN(n8268) );
  INV_X1 U9803 ( .A(n8268), .ZN(n8266) );
  NAND2_X1 U9804 ( .A1(n8267), .A2(n8266), .ZN(n8316) );
  AND2_X1 U9805 ( .A1(n8317), .A2(n8316), .ZN(n8275) );
  INV_X1 U9806 ( .A(n8316), .ZN(n8274) );
  NAND2_X1 U9807 ( .A1(n8269), .A2(n8268), .ZN(n8315) );
  INV_X1 U9808 ( .A(n8270), .ZN(n8272) );
  OR2_X1 U9809 ( .A1(n8272), .A2(n8271), .ZN(n8319) );
  AND2_X1 U9810 ( .A1(n8315), .A2(n8319), .ZN(n8273) );
  NAND2_X1 U9811 ( .A1(n8287), .A2(n4535), .ZN(n8277) );
  NAND2_X1 U9812 ( .A1(n9579), .A2(n8496), .ZN(n8276) );
  NAND2_X1 U9813 ( .A1(n8277), .A2(n8276), .ZN(n8439) );
  NAND2_X1 U9814 ( .A1(n8287), .A2(n8592), .ZN(n8279) );
  OR2_X1 U9815 ( .A1(n8327), .A2(n8593), .ZN(n8278) );
  NAND2_X1 U9816 ( .A1(n8279), .A2(n8278), .ZN(n8280) );
  XNOR2_X1 U9817 ( .A(n8280), .B(n8476), .ZN(n8440) );
  XOR2_X1 U9818 ( .A(n8439), .B(n8440), .Z(n8281) );
  XNOR2_X1 U9819 ( .A(n4493), .B(n8281), .ZN(n8289) );
  AOI21_X1 U9820 ( .B1(n9553), .B2(n9580), .A(n8282), .ZN(n8285) );
  NAND2_X1 U9821 ( .A1(n9560), .A2(n8283), .ZN(n8284) );
  OAI211_X1 U9822 ( .C1(n8441), .C2(n9555), .A(n8285), .B(n8284), .ZN(n8286)
         );
  AOI21_X1 U9823 ( .B1(n9518), .B2(n8287), .A(n8286), .ZN(n8288) );
  OAI21_X1 U9824 ( .B1(n8289), .B2(n9520), .A(n8288), .ZN(P1_U3232) );
  INV_X1 U9825 ( .A(n8304), .ZN(n8835) );
  OR2_X1 U9826 ( .A1(n9342), .A2(n8835), .ZN(n8292) );
  NAND2_X1 U9827 ( .A1(n8295), .A2(n8299), .ZN(n8296) );
  NAND2_X1 U9828 ( .A1(n8913), .A2(n8296), .ZN(n9336) );
  NAND2_X1 U9829 ( .A1(n9219), .A2(n9230), .ZN(n8301) );
  NAND2_X1 U9830 ( .A1(n8301), .A2(n8298), .ZN(n8297) );
  NAND2_X1 U9831 ( .A1(n8297), .A2(n8294), .ZN(n8302) );
  AND2_X1 U9832 ( .A1(n8299), .A2(n8298), .ZN(n8300) );
  NAND2_X1 U9833 ( .A1(n8301), .A2(n8300), .ZN(n9201) );
  NAND2_X1 U9834 ( .A1(n8302), .A2(n9201), .ZN(n8303) );
  NAND2_X1 U9835 ( .A1(n8303), .A2(n9225), .ZN(n8307) );
  OAI22_X1 U9836 ( .A1(n8914), .A2(n9205), .B1(n8304), .B2(n9203), .ZN(n8305)
         );
  INV_X1 U9837 ( .A(n8305), .ZN(n8306) );
  NAND2_X1 U9838 ( .A1(n8307), .A2(n8306), .ZN(n9340) );
  NAND2_X1 U9839 ( .A1(n9340), .A2(n9060), .ZN(n8314) );
  INV_X1 U9840 ( .A(n8911), .ZN(n9337) );
  NOR2_X1 U9841 ( .A1(n4489), .A2(n9337), .ZN(n8308) );
  INV_X1 U9842 ( .A(n9338), .ZN(n8312) );
  AOI22_X1 U9843 ( .A1(n4392), .A2(P2_REG2_REG_13__SCAN_IN), .B1(n8309), .B2(
        n10517), .ZN(n8310) );
  OAI21_X1 U9844 ( .B1(n9337), .B2(n10523), .A(n8310), .ZN(n8311) );
  AOI21_X1 U9845 ( .B1(n8312), .B2(n9234), .A(n8311), .ZN(n8313) );
  OAI211_X1 U9846 ( .C1(n9336), .C2(n9231), .A(n8314), .B(n8313), .ZN(P2_U3283) );
  NAND2_X1 U9847 ( .A1(n8316), .A2(n8315), .ZN(n8322) );
  NAND2_X1 U9848 ( .A1(n8318), .A2(n8317), .ZN(n8320) );
  AND2_X1 U9849 ( .A1(n8319), .A2(n8320), .ZN(n8321) );
  XOR2_X1 U9850 ( .A(n8322), .B(n8321), .Z(n8331) );
  AOI21_X1 U9851 ( .B1(n9553), .B2(n9581), .A(n8323), .ZN(n8326) );
  NAND2_X1 U9852 ( .A1(n9560), .A2(n8324), .ZN(n8325) );
  OAI211_X1 U9853 ( .C1(n8327), .C2(n9555), .A(n8326), .B(n8325), .ZN(n8328)
         );
  AOI21_X1 U9854 ( .B1(n9518), .B2(n8329), .A(n8328), .ZN(n8330) );
  OAI21_X1 U9855 ( .B1(n8331), .B2(n9520), .A(n8330), .ZN(P1_U3222) );
  OAI222_X1 U9856 ( .A1(P1_U3084), .A2(n8334), .B1(n10292), .B2(n8333), .C1(
        n8332), .C2(n10294), .ZN(P1_U3329) );
  XNOR2_X1 U9857 ( .A(n8336), .B(n8337), .ZN(n8410) );
  INV_X1 U9858 ( .A(n8410), .ZN(n8348) );
  NAND3_X1 U9859 ( .A1(n8339), .A2(n8337), .A3(n8338), .ZN(n10152) );
  INV_X1 U9860 ( .A(n10152), .ZN(n8341) );
  AOI21_X1 U9861 ( .B1(n8339), .B2(n8338), .A(n8337), .ZN(n8340) );
  NOR2_X1 U9862 ( .A1(n8341), .A2(n8340), .ZN(n8342) );
  OAI222_X1 U9863 ( .A1(n10405), .A2(n10132), .B1(n10403), .B2(n8441), .C1(
        n8342), .C2(n10406), .ZN(n8408) );
  OR2_X1 U9864 ( .A1(n8221), .A2(n9557), .ZN(n8343) );
  AND3_X1 U9865 ( .A1(n10159), .A2(n8343), .A3(n10418), .ZN(n8409) );
  NAND2_X1 U9866 ( .A1(n8409), .A2(n10422), .ZN(n8345) );
  AOI22_X1 U9867 ( .A1(n10123), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n9561), .B2(
        n10411), .ZN(n8344) );
  OAI211_X1 U9868 ( .C1(n9557), .C2(n10400), .A(n8345), .B(n8344), .ZN(n8346)
         );
  AOI21_X1 U9869 ( .B1(n8408), .B2(n10148), .A(n8346), .ZN(n8347) );
  OAI21_X1 U9870 ( .B1(n10142), .B2(n8348), .A(n8347), .ZN(P1_U3276) );
  INV_X1 U9871 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n8352) );
  AOI211_X1 U9872 ( .C1(n8351), .C2(n10489), .A(n8350), .B(n8349), .ZN(n8354)
         );
  MUX2_X1 U9873 ( .A(n8352), .B(n8354), .S(n10492), .Z(n8353) );
  OAI21_X1 U9874 ( .B1(n8357), .B2(n10275), .A(n8353), .ZN(P1_U3490) );
  MUX2_X1 U9875 ( .A(n8355), .B(n8354), .S(n10504), .Z(n8356) );
  OAI21_X1 U9876 ( .B1(n8357), .B2(n10236), .A(n8356), .ZN(P1_U3535) );
  INV_X1 U9877 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n8361) );
  AOI211_X1 U9878 ( .C1(n8360), .C2(n10489), .A(n8359), .B(n8358), .ZN(n8363)
         );
  MUX2_X1 U9879 ( .A(n8361), .B(n8363), .S(n10492), .Z(n8362) );
  OAI21_X1 U9880 ( .B1(n8365), .B2(n10275), .A(n8362), .ZN(P1_U3493) );
  INV_X1 U9881 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n9617) );
  MUX2_X1 U9882 ( .A(n9617), .B(n8363), .S(n10504), .Z(n8364) );
  OAI21_X1 U9883 ( .B1(n8365), .B2(n10236), .A(n8364), .ZN(P1_U3536) );
  INV_X1 U9884 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n10641) );
  NOR2_X1 U9885 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n8366) );
  AOI21_X1 U9886 ( .B1(P1_ADDR_REG_17__SCAN_IN), .B2(P2_ADDR_REG_17__SCAN_IN), 
        .A(n8366), .ZN(n10613) );
  NOR2_X1 U9887 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n8367) );
  AOI21_X1 U9888 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(P2_ADDR_REG_16__SCAN_IN), 
        .A(n8367), .ZN(n10616) );
  NOR2_X1 U9889 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n8368) );
  AOI21_X1 U9890 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(P2_ADDR_REG_15__SCAN_IN), 
        .A(n8368), .ZN(n10619) );
  NOR2_X1 U9891 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n8369) );
  AOI21_X1 U9892 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(P2_ADDR_REG_14__SCAN_IN), 
        .A(n8369), .ZN(n10622) );
  NOR2_X1 U9893 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n8370) );
  AOI21_X1 U9894 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(P2_ADDR_REG_13__SCAN_IN), 
        .A(n8370), .ZN(n10625) );
  INV_X1 U9895 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n10650) );
  NAND2_X1 U9896 ( .A1(n7221), .A2(n10650), .ZN(n10649) );
  NOR2_X1 U9897 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n8378) );
  INV_X1 U9898 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n8371) );
  AOI22_X1 U9899 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(n8371), .B1(
        P2_ADDR_REG_4__SCAN_IN), .B2(n9855), .ZN(n10659) );
  INV_X1 U9900 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n8376) );
  AOI22_X1 U9901 ( .A1(P2_ADDR_REG_3__SCAN_IN), .A2(P1_ADDR_REG_3__SCAN_IN), 
        .B1(n7292), .B2(n8376), .ZN(n10657) );
  NAND2_X1 U9902 ( .A1(P1_ADDR_REG_2__SCAN_IN), .A2(P2_ADDR_REG_2__SCAN_IN), 
        .ZN(n8374) );
  AOI22_X1 U9903 ( .A1(P1_ADDR_REG_2__SCAN_IN), .A2(P2_ADDR_REG_2__SCAN_IN), 
        .B1(n8372), .B2(n9917), .ZN(n10655) );
  AOI21_X1 U9904 ( .B1(P1_ADDR_REG_0__SCAN_IN), .B2(P2_ADDR_REG_0__SCAN_IN), 
        .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n10606) );
  INV_X1 U9905 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n10610) );
  NAND3_X1 U9906 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(P1_ADDR_REG_0__SCAN_IN), 
        .A3(P2_ADDR_REG_0__SCAN_IN), .ZN(n10608) );
  OAI21_X1 U9907 ( .B1(n10606), .B2(n10610), .A(n10608), .ZN(n10654) );
  NAND2_X1 U9908 ( .A1(n10655), .A2(n10654), .ZN(n8373) );
  NAND2_X1 U9909 ( .A1(n8374), .A2(n8373), .ZN(n10656) );
  NAND2_X1 U9910 ( .A1(n10657), .A2(n10656), .ZN(n8375) );
  NOR2_X1 U9911 ( .A1(n10659), .A2(n10658), .ZN(n8377) );
  NOR2_X1 U9912 ( .A1(n8378), .A2(n8377), .ZN(n8379) );
  NOR2_X1 U9913 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n8379), .ZN(n10637) );
  AND2_X1 U9914 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n8379), .ZN(n10636) );
  NAND2_X1 U9915 ( .A1(n8381), .A2(P1_ADDR_REG_6__SCAN_IN), .ZN(n8383) );
  XOR2_X1 U9916 ( .A(n8381), .B(P1_ADDR_REG_6__SCAN_IN), .Z(n10635) );
  NAND2_X1 U9917 ( .A1(n10635), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n8382) );
  NAND2_X1 U9918 ( .A1(n8383), .A2(n8382), .ZN(n8384) );
  NAND2_X1 U9919 ( .A1(P1_ADDR_REG_7__SCAN_IN), .A2(n8384), .ZN(n8386) );
  XOR2_X1 U9920 ( .A(P1_ADDR_REG_7__SCAN_IN), .B(n8384), .Z(n10653) );
  NAND2_X1 U9921 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(n10653), .ZN(n8385) );
  NAND2_X1 U9922 ( .A1(n8386), .A2(n8385), .ZN(n10651) );
  AOI22_X1 U9923 ( .A1(P1_ADDR_REG_8__SCAN_IN), .A2(P2_ADDR_REG_8__SCAN_IN), 
        .B1(n10649), .B2(n10651), .ZN(n8387) );
  INV_X1 U9924 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n8388) );
  NAND2_X1 U9925 ( .A1(n8387), .A2(n8388), .ZN(n10646) );
  OR2_X1 U9926 ( .A1(n8388), .A2(n8387), .ZN(n10647) );
  INV_X1 U9927 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n10648) );
  NAND2_X1 U9928 ( .A1(n10647), .A2(n10648), .ZN(n10644) );
  NAND2_X1 U9929 ( .A1(n10646), .A2(n10644), .ZN(n10634) );
  NAND2_X1 U9930 ( .A1(P1_ADDR_REG_10__SCAN_IN), .A2(P2_ADDR_REG_10__SCAN_IN), 
        .ZN(n8389) );
  OAI21_X1 U9931 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(P2_ADDR_REG_10__SCAN_IN), 
        .A(n8389), .ZN(n10633) );
  NAND2_X1 U9932 ( .A1(P1_ADDR_REG_11__SCAN_IN), .A2(P2_ADDR_REG_11__SCAN_IN), 
        .ZN(n8390) );
  OAI21_X1 U9933 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(P2_ADDR_REG_11__SCAN_IN), 
        .A(n8390), .ZN(n10630) );
  NOR2_X1 U9934 ( .A1(P1_ADDR_REG_12__SCAN_IN), .A2(P2_ADDR_REG_12__SCAN_IN), 
        .ZN(n8391) );
  AOI21_X1 U9935 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(P1_ADDR_REG_12__SCAN_IN), 
        .A(n8391), .ZN(n10627) );
  NAND2_X1 U9936 ( .A1(n10628), .A2(n10627), .ZN(n10626) );
  NAND2_X1 U9937 ( .A1(n10625), .A2(n10624), .ZN(n10623) );
  NAND2_X1 U9938 ( .A1(n10622), .A2(n10621), .ZN(n10620) );
  OAI21_X1 U9939 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(P1_ADDR_REG_14__SCAN_IN), 
        .A(n10620), .ZN(n10618) );
  NAND2_X1 U9940 ( .A1(n10619), .A2(n10618), .ZN(n10617) );
  OAI21_X1 U9941 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(P1_ADDR_REG_15__SCAN_IN), 
        .A(n10617), .ZN(n10615) );
  NAND2_X1 U9942 ( .A1(n10616), .A2(n10615), .ZN(n10614) );
  OAI21_X1 U9943 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(P1_ADDR_REG_16__SCAN_IN), 
        .A(n10614), .ZN(n10612) );
  NAND2_X1 U9944 ( .A1(n10613), .A2(n10612), .ZN(n10611) );
  NOR2_X1 U9945 ( .A1(n10641), .A2(n10640), .ZN(n8392) );
  NAND2_X1 U9946 ( .A1(n10641), .A2(n10640), .ZN(n10639) );
  OAI21_X1 U9947 ( .B1(P1_ADDR_REG_18__SCAN_IN), .B2(n8392), .A(n10639), .ZN(
        n8394) );
  XNOR2_X1 U9948 ( .A(n8560), .B(P1_ADDR_REG_19__SCAN_IN), .ZN(n8393) );
  XNOR2_X1 U9949 ( .A(n8394), .B(n8393), .ZN(ADD_1071_U4) );
  INV_X1 U9950 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n8398) );
  AOI211_X1 U9951 ( .C1(n8397), .C2(n10489), .A(n8396), .B(n8395), .ZN(n8400)
         );
  MUX2_X1 U9952 ( .A(n8398), .B(n8400), .S(n10492), .Z(n8399) );
  OAI21_X1 U9953 ( .B1(n9423), .B2(n10275), .A(n8399), .ZN(P1_U3496) );
  INV_X1 U9954 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n9864) );
  MUX2_X1 U9955 ( .A(n9864), .B(n8400), .S(n10504), .Z(n8401) );
  OAI21_X1 U9956 ( .B1(n9423), .B2(n10236), .A(n8401), .ZN(P1_U3537) );
  INV_X1 U9957 ( .A(n8402), .ZN(n8406) );
  OAI222_X1 U9958 ( .A1(n9395), .A2(n8404), .B1(n9399), .B2(n8406), .C1(n8403), 
        .C2(P2_U3152), .ZN(P2_U3333) );
  OAI222_X1 U9959 ( .A1(n10294), .A2(n8407), .B1(n10292), .B2(n8406), .C1(
        P1_U3084), .C2(n8405), .ZN(P1_U3328) );
  INV_X1 U9960 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n8411) );
  AOI211_X1 U9961 ( .C1(n8410), .C2(n10489), .A(n8409), .B(n8408), .ZN(n8413)
         );
  MUX2_X1 U9962 ( .A(n8411), .B(n8413), .S(n10504), .Z(n8412) );
  OAI21_X1 U9963 ( .B1(n9557), .B2(n10236), .A(n8412), .ZN(P1_U3538) );
  INV_X1 U9964 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n8414) );
  MUX2_X1 U9965 ( .A(n8414), .B(n8413), .S(n10492), .Z(n8415) );
  OAI21_X1 U9966 ( .B1(n9557), .B2(n10275), .A(n8415), .ZN(P1_U3499) );
  INV_X1 U9967 ( .A(n8416), .ZN(n8419) );
  OAI222_X1 U9968 ( .A1(n9399), .A2(n8419), .B1(P2_U3152), .B2(n8417), .C1(
        n9836), .C2(n9395), .ZN(P2_U3332) );
  OAI222_X1 U9969 ( .A1(P1_U3084), .A2(n6067), .B1(n10292), .B2(n8419), .C1(
        n8418), .C2(n10294), .ZN(P1_U3327) );
  INV_X1 U9970 ( .A(n8420), .ZN(n9398) );
  AOI21_X1 U9971 ( .B1(n10281), .B2(P2_DATAO_REG_27__SCAN_IN), .A(n8421), .ZN(
        n8422) );
  OAI21_X1 U9972 ( .B1(n9398), .B2(n10283), .A(n8422), .ZN(P1_U3326) );
  INV_X1 U9973 ( .A(P1_REG0_REG_22__SCAN_IN), .ZN(n8434) );
  OAI21_X1 U9974 ( .B1(n8425), .B2(n8424), .A(n8423), .ZN(n10035) );
  OAI211_X1 U9975 ( .C1(n6053), .C2(n10057), .A(n10418), .B(n10014), .ZN(
        n10034) );
  OAI21_X1 U9976 ( .B1(n10035), .B2(n10243), .A(n10034), .ZN(n8433) );
  NAND2_X1 U9977 ( .A1(n10069), .A2(n8426), .ZN(n10041) );
  NAND2_X1 U9978 ( .A1(n10041), .A2(n10048), .ZN(n10040) );
  NAND2_X1 U9979 ( .A1(n10040), .A2(n8427), .ZN(n8429) );
  NAND2_X1 U9980 ( .A1(n8429), .A2(n8430), .ZN(n8428) );
  OAI211_X1 U9981 ( .C1(n8430), .C2(n8429), .A(n8428), .B(n10101), .ZN(n8432)
         );
  NAND2_X1 U9982 ( .A1(n9572), .A2(n10103), .ZN(n8431) );
  OAI211_X1 U9983 ( .C1(n9721), .C2(n10405), .A(n8432), .B(n8431), .ZN(n10038)
         );
  NOR2_X1 U9984 ( .A1(n8433), .A2(n10038), .ZN(n8436) );
  MUX2_X1 U9985 ( .A(n8434), .B(n8436), .S(n10492), .Z(n8435) );
  OAI21_X1 U9986 ( .B1(n6053), .B2(n10275), .A(n8435), .ZN(P1_U3513) );
  INV_X1 U9987 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n8437) );
  MUX2_X1 U9988 ( .A(n8437), .B(n8436), .S(n10504), .Z(n8438) );
  OAI21_X1 U9989 ( .B1(n6053), .B2(n10236), .A(n8438), .ZN(P1_U3545) );
  NAND2_X1 U9990 ( .A1(n8450), .A2(n8592), .ZN(n8443) );
  OR2_X1 U9991 ( .A1(n8441), .A2(n8593), .ZN(n8442) );
  NAND2_X1 U9992 ( .A1(n8443), .A2(n8442), .ZN(n8444) );
  XNOR2_X1 U9993 ( .A(n8444), .B(n8476), .ZN(n8448) );
  NAND2_X1 U9994 ( .A1(n8449), .A2(n8448), .ZN(n9412) );
  NAND2_X1 U9995 ( .A1(n8454), .A2(n8592), .ZN(n8446) );
  NAND2_X1 U9996 ( .A1(n9577), .A2(n4535), .ZN(n8445) );
  NAND2_X1 U9997 ( .A1(n8446), .A2(n8445), .ZN(n8447) );
  XNOR2_X1 U9998 ( .A(n8447), .B(n8563), .ZN(n8457) );
  AND2_X1 U9999 ( .A1(n9412), .A2(n8457), .ZN(n8453) );
  NAND2_X1 U10000 ( .A1(n8450), .A2(n4535), .ZN(n8452) );
  NAND2_X1 U10001 ( .A1(n9578), .A2(n8496), .ZN(n8451) );
  NAND2_X1 U10002 ( .A1(n8452), .A2(n8451), .ZN(n9411) );
  NAND2_X1 U10003 ( .A1(n8454), .A2(n4535), .ZN(n8456) );
  NAND2_X1 U10004 ( .A1(n9577), .A2(n8496), .ZN(n8455) );
  NAND2_X1 U10005 ( .A1(n8456), .A2(n8455), .ZN(n9550) );
  NAND2_X1 U10006 ( .A1(n9416), .A2(n9412), .ZN(n8459) );
  INV_X1 U10007 ( .A(n8457), .ZN(n8458) );
  NAND2_X1 U10008 ( .A1(n10226), .A2(n8592), .ZN(n8461) );
  NAND2_X1 U10009 ( .A1(n10104), .A2(n4535), .ZN(n8460) );
  NAND2_X1 U10010 ( .A1(n8461), .A2(n8460), .ZN(n8462) );
  XNOR2_X1 U10011 ( .A(n8462), .B(n8563), .ZN(n9477) );
  NOR2_X1 U10012 ( .A1(n10156), .A2(n8599), .ZN(n8463) );
  AOI21_X1 U10013 ( .B1(n10226), .B2(n4535), .A(n8463), .ZN(n8469) );
  NOR2_X1 U10014 ( .A1(n10132), .A2(n8599), .ZN(n8464) );
  AOI21_X1 U10015 ( .B1(n10230), .B2(n4535), .A(n8464), .ZN(n8468) );
  NAND2_X1 U10016 ( .A1(n10230), .A2(n8592), .ZN(n8466) );
  NAND2_X1 U10017 ( .A1(n9575), .A2(n4535), .ZN(n8465) );
  NAND2_X1 U10018 ( .A1(n8466), .A2(n8465), .ZN(n8467) );
  XNOR2_X1 U10019 ( .A(n8467), .B(n8563), .ZN(n9474) );
  OAI22_X1 U10020 ( .A1(n9477), .A2(n8469), .B1(n8468), .B2(n9474), .ZN(n8473)
         );
  INV_X1 U10021 ( .A(n9474), .ZN(n9471) );
  INV_X1 U10022 ( .A(n8468), .ZN(n9470) );
  INV_X1 U10023 ( .A(n8469), .ZN(n9476) );
  OAI21_X1 U10024 ( .B1(n9471), .B2(n9470), .A(n9476), .ZN(n8471) );
  NOR2_X1 U10025 ( .A1(n9476), .A2(n9470), .ZN(n8470) );
  AOI22_X1 U10026 ( .A1(n8471), .A2(n9477), .B1(n9474), .B2(n8470), .ZN(n8472)
         );
  NAND2_X1 U10027 ( .A1(n10217), .A2(n8592), .ZN(n8475) );
  OR2_X1 U10028 ( .A1(n10107), .A2(n8593), .ZN(n8474) );
  NAND2_X1 U10029 ( .A1(n8475), .A2(n8474), .ZN(n8477) );
  XNOR2_X1 U10030 ( .A(n8477), .B(n8476), .ZN(n9440) );
  NAND2_X1 U10031 ( .A1(n10217), .A2(n4535), .ZN(n8479) );
  OR2_X1 U10032 ( .A1(n10107), .A2(n8599), .ZN(n8478) );
  NAND2_X1 U10033 ( .A1(n8479), .A2(n8478), .ZN(n9439) );
  NAND2_X1 U10034 ( .A1(n9440), .A2(n9439), .ZN(n9438) );
  NAND2_X1 U10035 ( .A1(n10114), .A2(n8592), .ZN(n8481) );
  NAND2_X1 U10036 ( .A1(n9574), .A2(n4535), .ZN(n8480) );
  NAND2_X1 U10037 ( .A1(n8481), .A2(n8480), .ZN(n8482) );
  XNOR2_X1 U10038 ( .A(n8482), .B(n8476), .ZN(n8487) );
  NAND2_X1 U10039 ( .A1(n10114), .A2(n4535), .ZN(n8484) );
  NAND2_X1 U10040 ( .A1(n9574), .A2(n8496), .ZN(n8483) );
  NAND2_X1 U10041 ( .A1(n8484), .A2(n8483), .ZN(n9513) );
  NAND2_X1 U10042 ( .A1(n8487), .A2(n9513), .ZN(n8485) );
  AND2_X1 U10043 ( .A1(n9438), .A2(n8485), .ZN(n8486) );
  OAI21_X1 U10044 ( .B1(n8487), .B2(n9513), .A(n9439), .ZN(n8490) );
  INV_X1 U10045 ( .A(n9440), .ZN(n8489) );
  INV_X1 U10046 ( .A(n8487), .ZN(n9437) );
  NOR2_X1 U10047 ( .A1(n9439), .A2(n9513), .ZN(n8488) );
  AOI22_X1 U10048 ( .A1(n8490), .A2(n8489), .B1(n9437), .B2(n8488), .ZN(n8491)
         );
  NAND2_X1 U10049 ( .A1(n10075), .A2(n8592), .ZN(n8494) );
  NAND2_X1 U10050 ( .A1(n9573), .A2(n4535), .ZN(n8493) );
  NAND2_X1 U10051 ( .A1(n8494), .A2(n8493), .ZN(n8495) );
  XNOR2_X1 U10052 ( .A(n8495), .B(n8476), .ZN(n8499) );
  NAND2_X1 U10053 ( .A1(n10075), .A2(n6956), .ZN(n8498) );
  NAND2_X1 U10054 ( .A1(n9573), .A2(n8496), .ZN(n8497) );
  NAND2_X1 U10055 ( .A1(n8498), .A2(n8497), .ZN(n8500) );
  NAND2_X1 U10056 ( .A1(n8499), .A2(n8500), .ZN(n9502) );
  INV_X1 U10057 ( .A(n8499), .ZN(n8502) );
  INV_X1 U10058 ( .A(n8500), .ZN(n8501) );
  NAND2_X1 U10059 ( .A1(n8502), .A2(n8501), .ZN(n9501) );
  NAND2_X1 U10060 ( .A1(n10061), .A2(n8592), .ZN(n8504) );
  NAND2_X1 U10061 ( .A1(n9572), .A2(n4535), .ZN(n8503) );
  NAND2_X1 U10062 ( .A1(n8504), .A2(n8503), .ZN(n8505) );
  XNOR2_X1 U10063 ( .A(n8505), .B(n8476), .ZN(n8511) );
  INV_X1 U10064 ( .A(n8511), .ZN(n8507) );
  NOR2_X1 U10065 ( .A1(n10074), .A2(n8599), .ZN(n8506) );
  AOI21_X1 U10066 ( .B1(n10061), .B2(n4535), .A(n8506), .ZN(n8510) );
  NAND2_X1 U10067 ( .A1(n8507), .A2(n8510), .ZN(n8509) );
  AND2_X1 U10068 ( .A1(n9501), .A2(n8509), .ZN(n8520) );
  NOR2_X1 U10069 ( .A1(n10042), .A2(n8599), .ZN(n8508) );
  AOI21_X1 U10070 ( .B1(n5346), .B2(n4535), .A(n8508), .ZN(n8521) );
  INV_X1 U10071 ( .A(n8509), .ZN(n8512) );
  XNOR2_X1 U10072 ( .A(n8511), .B(n8510), .ZN(n9450) );
  OR2_X1 U10073 ( .A1(n8512), .A2(n9450), .ZN(n8518) );
  OR2_X1 U10074 ( .A1(n8521), .A2(n8518), .ZN(n8513) );
  INV_X1 U10075 ( .A(n8513), .ZN(n8514) );
  NAND2_X1 U10076 ( .A1(n5346), .A2(n8592), .ZN(n8516) );
  NAND2_X1 U10077 ( .A1(n10022), .A2(n6956), .ZN(n8515) );
  NAND2_X1 U10078 ( .A1(n8516), .A2(n8515), .ZN(n8517) );
  XNOR2_X1 U10079 ( .A(n8517), .B(n8563), .ZN(n8523) );
  INV_X1 U10080 ( .A(n8518), .ZN(n8519) );
  INV_X1 U10081 ( .A(n9424), .ZN(n8522) );
  NOR2_X1 U10082 ( .A1(n9425), .A2(n8522), .ZN(n8526) );
  AOI21_X1 U10083 ( .B1(n8524), .B2(n9424), .A(n8523), .ZN(n8525) );
  OAI21_X1 U10084 ( .B1(n8526), .B2(n8525), .A(n9547), .ZN(n8531) );
  OAI22_X1 U10085 ( .A1(n10074), .A2(n9494), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8527), .ZN(n8529) );
  NOR2_X1 U10086 ( .A1(n9542), .A2(n10031), .ZN(n8528) );
  AOI211_X1 U10087 ( .C1(n9571), .C2(n9534), .A(n8529), .B(n8528), .ZN(n8530)
         );
  OAI211_X1 U10088 ( .C1(n6053), .C2(n9556), .A(n8531), .B(n8530), .ZN(
        P1_U3233) );
  OAI222_X1 U10089 ( .A1(n9399), .A2(n8534), .B1(n8533), .B2(P2_U3152), .C1(
        n8532), .C2(n9395), .ZN(P2_U3337) );
  OAI222_X1 U10090 ( .A1(n9395), .A2(n9862), .B1(n9399), .B2(n8536), .C1(
        P2_U3152), .C2(n8535), .ZN(P2_U3336) );
  NAND2_X1 U10091 ( .A1(n8869), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n8537) );
  OAI21_X1 U10092 ( .B1(n8869), .B2(P2_REG2_REG_16__SCAN_IN), .A(n8537), .ZN(
        n8865) );
  NAND2_X1 U10093 ( .A1(n8551), .A2(n8540), .ZN(n8541) );
  XNOR2_X1 U10094 ( .A(n8540), .B(n8852), .ZN(n8850) );
  INV_X1 U10095 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n8849) );
  NAND2_X1 U10096 ( .A1(n8543), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n8542) );
  OAI21_X1 U10097 ( .B1(n8543), .B2(P2_REG2_REG_17__SCAN_IN), .A(n8542), .ZN(
        n8874) );
  XNOR2_X1 U10098 ( .A(n8544), .B(n8547), .ZN(n8893) );
  INV_X1 U10099 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n8892) );
  NAND2_X1 U10100 ( .A1(n8893), .A2(n8892), .ZN(n8891) );
  INV_X1 U10101 ( .A(n8547), .ZN(n8897) );
  NAND2_X1 U10102 ( .A1(n8544), .A2(n8897), .ZN(n8545) );
  NAND2_X1 U10103 ( .A1(n8891), .A2(n8545), .ZN(n8546) );
  XNOR2_X1 U10104 ( .A(P2_REG2_REG_19__SCAN_IN), .B(n8546), .ZN(n8557) );
  OR2_X1 U10105 ( .A1(n8547), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n8554) );
  NAND2_X1 U10106 ( .A1(n8547), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n8548) );
  NAND2_X1 U10107 ( .A1(n8554), .A2(n8548), .ZN(n8886) );
  XNOR2_X1 U10108 ( .A(n8881), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n8877) );
  INV_X1 U10109 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n9924) );
  XNOR2_X1 U10110 ( .A(n8869), .B(P2_REG1_REG_16__SCAN_IN), .ZN(n8858) );
  NAND2_X1 U10111 ( .A1(n8852), .A2(n8552), .ZN(n8553) );
  XNOR2_X1 U10112 ( .A(n8552), .B(n8551), .ZN(n8846) );
  NAND2_X1 U10113 ( .A1(P2_REG1_REG_15__SCAN_IN), .A2(n8846), .ZN(n8845) );
  NAND2_X1 U10114 ( .A1(n8553), .A2(n8845), .ZN(n8859) );
  NOR2_X1 U10115 ( .A1(n8858), .A2(n8859), .ZN(n8857) );
  INV_X1 U10116 ( .A(n8554), .ZN(n8555) );
  NOR2_X1 U10117 ( .A1(n8885), .A2(n8555), .ZN(n8556) );
  XNOR2_X1 U10118 ( .A(n8556), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n8558) );
  NAND2_X1 U10119 ( .A1(P2_REG3_REG_19__SCAN_IN), .A2(P2_U3152), .ZN(n8559) );
  NAND2_X1 U10120 ( .A1(n10201), .A2(n8592), .ZN(n8562) );
  NAND2_X1 U10121 ( .A1(n9571), .A2(n4535), .ZN(n8561) );
  NAND2_X1 U10122 ( .A1(n8562), .A2(n8561), .ZN(n8564) );
  XNOR2_X1 U10123 ( .A(n8564), .B(n8563), .ZN(n9426) );
  NOR2_X1 U10124 ( .A1(n9721), .A2(n8599), .ZN(n8565) );
  AOI21_X1 U10125 ( .B1(n10201), .B2(n4535), .A(n8565), .ZN(n9485) );
  NAND2_X1 U10126 ( .A1(n9426), .A2(n9485), .ZN(n8566) );
  NAND2_X1 U10127 ( .A1(n9729), .A2(n8592), .ZN(n8568) );
  OR2_X1 U10128 ( .A1(n10025), .A2(n8593), .ZN(n8567) );
  NAND2_X1 U10129 ( .A1(n8568), .A2(n8567), .ZN(n8569) );
  XNOR2_X1 U10130 ( .A(n8569), .B(n8476), .ZN(n8576) );
  NOR2_X1 U10131 ( .A1(n10025), .A2(n8599), .ZN(n8570) );
  AOI21_X1 U10132 ( .B1(n9729), .B2(n4535), .A(n8570), .ZN(n8574) );
  XNOR2_X1 U10133 ( .A(n8576), .B(n8574), .ZN(n9490) );
  NAND2_X1 U10134 ( .A1(n8573), .A2(n8572), .ZN(n9489) );
  INV_X1 U10135 ( .A(n8574), .ZN(n8575) );
  OAI22_X1 U10136 ( .A1(n9708), .A2(n8593), .B1(n9722), .B2(n8599), .ZN(n8582)
         );
  NAND2_X1 U10137 ( .A1(n10190), .A2(n8592), .ZN(n8579) );
  OR2_X1 U10138 ( .A1(n9722), .A2(n8593), .ZN(n8578) );
  NAND2_X1 U10139 ( .A1(n8579), .A2(n8578), .ZN(n8580) );
  XNOR2_X1 U10140 ( .A(n8580), .B(n8476), .ZN(n8581) );
  XOR2_X1 U10141 ( .A(n8582), .B(n8581), .Z(n9458) );
  INV_X1 U10142 ( .A(n8581), .ZN(n8584) );
  INV_X1 U10143 ( .A(n8582), .ZN(n8583) );
  NAND2_X1 U10144 ( .A1(n9690), .A2(n8592), .ZN(n8586) );
  NAND2_X1 U10145 ( .A1(n9568), .A2(n6956), .ZN(n8585) );
  NAND2_X1 U10146 ( .A1(n8586), .A2(n8585), .ZN(n8587) );
  XNOR2_X1 U10147 ( .A(n8587), .B(n8476), .ZN(n8589) );
  NOR2_X1 U10148 ( .A1(n9699), .A2(n8599), .ZN(n8588) );
  AOI21_X1 U10149 ( .B1(n9690), .B2(n4535), .A(n8588), .ZN(n8590) );
  XNOR2_X1 U10150 ( .A(n8589), .B(n8590), .ZN(n9540) );
  INV_X1 U10151 ( .A(n8589), .ZN(n8591) );
  NAND2_X1 U10152 ( .A1(n10178), .A2(n8592), .ZN(n8595) );
  OR2_X1 U10153 ( .A1(n9687), .A2(n8593), .ZN(n8594) );
  NAND2_X1 U10154 ( .A1(n8595), .A2(n8594), .ZN(n8596) );
  XNOR2_X1 U10155 ( .A(n8596), .B(n8476), .ZN(n9402) );
  NOR2_X1 U10156 ( .A1(n9687), .A2(n8599), .ZN(n8597) );
  AOI21_X1 U10157 ( .B1(n10178), .B2(n4535), .A(n8597), .ZN(n9401) );
  INV_X1 U10158 ( .A(n9401), .ZN(n8607) );
  NAND2_X1 U10159 ( .A1(n8619), .A2(n6956), .ZN(n8601) );
  OR2_X1 U10160 ( .A1(n9671), .A2(n8599), .ZN(n8600) );
  NAND2_X1 U10161 ( .A1(n8601), .A2(n8600), .ZN(n8602) );
  XNOR2_X1 U10162 ( .A(n8602), .B(n8476), .ZN(n8605) );
  AOI22_X1 U10163 ( .A1(n8619), .A2(n8592), .B1(n4535), .B2(n9566), .ZN(n8604)
         );
  XNOR2_X1 U10164 ( .A(n8605), .B(n8604), .ZN(n8612) );
  INV_X1 U10165 ( .A(n8612), .ZN(n8606) );
  NAND2_X1 U10166 ( .A1(n8606), .A2(n9547), .ZN(n8617) );
  NAND2_X1 U10167 ( .A1(n9402), .A2(n8607), .ZN(n8611) );
  NAND4_X1 U10168 ( .A1(n8618), .A2(n9547), .A3(n8612), .A4(n8611), .ZN(n8616)
         );
  NAND2_X1 U10169 ( .A1(n9567), .A2(n9553), .ZN(n8609) );
  AOI22_X1 U10170 ( .A1(n8620), .A2(n9560), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3084), .ZN(n8608) );
  OAI211_X1 U10171 ( .C1(n8610), .C2(n9555), .A(n8609), .B(n8608), .ZN(n8614)
         );
  NOR3_X1 U10172 ( .A1(n8612), .A2(n9520), .A3(n8611), .ZN(n8613) );
  AOI211_X1 U10173 ( .C1(n9518), .C2(n8619), .A(n8614), .B(n8613), .ZN(n8615)
         );
  OAI211_X1 U10174 ( .C1(n8618), .C2(n8617), .A(n8616), .B(n8615), .ZN(
        P1_U3218) );
  AOI22_X1 U10175 ( .A1(n8619), .A2(n10150), .B1(n10123), .B2(
        P1_REG2_REG_28__SCAN_IN), .ZN(n8625) );
  INV_X1 U10176 ( .A(n8620), .ZN(n8621) );
  OAI22_X1 U10177 ( .A1(n4442), .A2(n9632), .B1(n10145), .B2(n8621), .ZN(n8622) );
  OAI21_X1 U10178 ( .B1(n8623), .B2(n8622), .A(n10148), .ZN(n8624) );
  OAI211_X1 U10179 ( .C1(n8626), .C2(n10142), .A(n8625), .B(n8624), .ZN(
        P1_U3263) );
  INV_X1 U10180 ( .A(n8627), .ZN(n9390) );
  INV_X1 U10181 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n8628) );
  OAI222_X1 U10182 ( .A1(P1_U3084), .A2(n8629), .B1(n10283), .B2(n9390), .C1(
        n8628), .C2(n10294), .ZN(P1_U3323) );
  INV_X1 U10183 ( .A(n9278), .ZN(n9034) );
  INV_X1 U10184 ( .A(n9327), .ZN(n8915) );
  INV_X1 U10185 ( .A(n9331), .ZN(n9215) );
  AND2_X1 U10186 ( .A1(n8915), .A2(n9215), .ZN(n8631) );
  INV_X1 U10187 ( .A(n9317), .ZN(n9156) );
  AND2_X2 U10188 ( .A1(n9165), .A2(n9156), .ZN(n9127) );
  INV_X1 U10189 ( .A(n9312), .ZN(n9133) );
  NAND2_X1 U10190 ( .A1(n9034), .A2(n9057), .ZN(n9028) );
  XOR2_X1 U10191 ( .A(n8630), .B(n8900), .Z(n9237) );
  NAND2_X1 U10192 ( .A1(n8635), .A2(P2_B_REG_SCAN_IN), .ZN(n8636) );
  NAND2_X1 U10193 ( .A1(n9222), .A2(n8636), .ZN(n8907) );
  INV_X1 U10194 ( .A(n8907), .ZN(n8637) );
  NAND2_X1 U10195 ( .A1(n8830), .A2(n8637), .ZN(n9239) );
  NOR2_X1 U10196 ( .A1(n4392), .A2(n9239), .ZN(n8902) );
  AOI21_X1 U10197 ( .B1(n4392), .B2(P2_REG2_REG_31__SCAN_IN), .A(n8902), .ZN(
        n8639) );
  NAND2_X1 U10198 ( .A1(n8630), .A2(n9190), .ZN(n8638) );
  OAI211_X1 U10199 ( .C1(n9237), .C2(n8974), .A(n8639), .B(n8638), .ZN(
        P2_U3265) );
  INV_X1 U10200 ( .A(n8640), .ZN(n10286) );
  INV_X1 U10201 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n8641) );
  OAI222_X1 U10202 ( .A1(n9399), .A2(n10286), .B1(n8642), .B2(P2_U3152), .C1(
        n8641), .C2(n9395), .ZN(P2_U3329) );
  INV_X1 U10203 ( .A(n8991), .ZN(n8831) );
  NAND3_X1 U10204 ( .A1(n8645), .A2(n8826), .A3(n8831), .ZN(n8646) );
  OAI21_X1 U10205 ( .B1(n8647), .B2(n8821), .A(n8646), .ZN(n8649) );
  NAND2_X1 U10206 ( .A1(n8649), .A2(n8648), .ZN(n8653) );
  NOR2_X1 U10207 ( .A1(n8984), .A2(n8818), .ZN(n8651) );
  OAI22_X1 U10208 ( .A1(n8992), .A2(n8785), .B1(n8991), .B2(n8786), .ZN(n8650)
         );
  AOI211_X1 U10209 ( .C1(P2_REG3_REG_27__SCAN_IN), .C2(P2_U3152), .A(n8651), 
        .B(n8650), .ZN(n8652) );
  OAI211_X1 U10210 ( .C1(n8987), .C2(n8695), .A(n8653), .B(n8652), .ZN(
        P2_U3216) );
  INV_X1 U10211 ( .A(n8655), .ZN(n8656) );
  AOI21_X1 U10212 ( .B1(n8657), .B2(n8654), .A(n8656), .ZN(n8662) );
  OAI22_X1 U10213 ( .A1(n9204), .A2(n8786), .B1(n8785), .B2(n9206), .ZN(n8658)
         );
  AOI211_X1 U10214 ( .C1(n8761), .C2(n9213), .A(n8659), .B(n8658), .ZN(n8661)
         );
  NAND2_X1 U10215 ( .A1(n9331), .A2(n8825), .ZN(n8660) );
  OAI211_X1 U10216 ( .C1(n8662), .C2(n8821), .A(n8661), .B(n8660), .ZN(
        P2_U3217) );
  INV_X1 U10217 ( .A(n8663), .ZN(n8664) );
  NAND2_X1 U10218 ( .A1(n8665), .A2(n8664), .ZN(n8667) );
  XNOR2_X1 U10219 ( .A(n8667), .B(n8666), .ZN(n8669) );
  NAND3_X1 U10220 ( .A1(n8669), .A2(n6894), .A3(n8668), .ZN(n8677) );
  INV_X1 U10221 ( .A(n8669), .ZN(n8670) );
  INV_X1 U10222 ( .A(n9077), .ZN(n8924) );
  NAND3_X1 U10223 ( .A1(n8670), .A2(n8826), .A3(n8924), .ZN(n8676) );
  OAI22_X1 U10224 ( .A1(n8818), .A2(n9058), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8671), .ZN(n8674) );
  OAI22_X1 U10225 ( .A1(n9092), .A2(n8786), .B1(n8785), .B2(n8672), .ZN(n8673)
         );
  AOI211_X1 U10226 ( .C1(n9286), .C2(n8825), .A(n8674), .B(n8673), .ZN(n8675)
         );
  NAND3_X1 U10227 ( .A1(n8677), .A2(n8676), .A3(n8675), .ZN(P2_U3218) );
  INV_X1 U10228 ( .A(n8679), .ZN(n8680) );
  AOI21_X1 U10229 ( .B1(n8678), .B2(n8681), .A(n8680), .ZN(n8686) );
  INV_X1 U10230 ( .A(n9115), .ZN(n8683) );
  OAI22_X1 U10231 ( .A1(n9091), .A2(n9205), .B1(n8917), .B2(n9203), .ZN(n9121)
         );
  AOI22_X1 U10232 ( .A1(n8816), .A2(n9121), .B1(P2_REG3_REG_19__SCAN_IN), .B2(
        P2_U3152), .ZN(n8682) );
  OAI21_X1 U10233 ( .B1(n8683), .B2(n8818), .A(n8682), .ZN(n8684) );
  AOI21_X1 U10234 ( .B1(n9307), .B2(n8825), .A(n8684), .ZN(n8685) );
  OAI21_X1 U10235 ( .B1(n8686), .B2(n8821), .A(n8685), .ZN(P2_U3221) );
  INV_X1 U10236 ( .A(n8687), .ZN(n8688) );
  AOI21_X1 U10237 ( .B1(n7657), .B2(n8688), .A(n8821), .ZN(n8692) );
  NOR3_X1 U10238 ( .A1(n8793), .A2(n8690), .A3(n8689), .ZN(n8691) );
  OAI21_X1 U10239 ( .B1(n8692), .B2(n8691), .A(n7746), .ZN(n8700) );
  AOI22_X1 U10240 ( .A1(n8694), .A2(n8837), .B1(n8761), .B2(n8693), .ZN(n8699)
         );
  OAI22_X1 U10241 ( .A1(n8695), .A2(n10589), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9876), .ZN(n8696) );
  AOI21_X1 U10242 ( .B1(n8697), .B2(n8839), .A(n8696), .ZN(n8698) );
  NAND3_X1 U10243 ( .A1(n8700), .A2(n8699), .A3(n8698), .ZN(P2_U3223) );
  XNOR2_X1 U10244 ( .A(n8701), .B(n8702), .ZN(n8707) );
  INV_X1 U10245 ( .A(n9084), .ZN(n8703) );
  OAI22_X1 U10246 ( .A1(n8818), .A2(n8703), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9925), .ZN(n8705) );
  OAI22_X1 U10247 ( .A1(n9091), .A2(n8786), .B1(n8785), .B2(n9092), .ZN(n8704)
         );
  AOI211_X1 U10248 ( .C1(n9296), .C2(n8825), .A(n8705), .B(n8704), .ZN(n8706)
         );
  OAI21_X1 U10249 ( .B1(n8707), .B2(n8821), .A(n8706), .ZN(P2_U3225) );
  XNOR2_X1 U10250 ( .A(n8709), .B(n8708), .ZN(n8710) );
  XNOR2_X1 U10251 ( .A(n8711), .B(n8710), .ZN(n8716) );
  NOR2_X1 U10252 ( .A1(n8818), .A2(n9021), .ZN(n8714) );
  AOI22_X1 U10253 ( .A1(n8831), .A2(n9222), .B1(n9220), .B2(n9049), .ZN(n9018)
         );
  OAI22_X1 U10254 ( .A1(n9018), .A2(n8712), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9966), .ZN(n8713) );
  AOI211_X1 U10255 ( .C1(n9275), .C2(n8825), .A(n8714), .B(n8713), .ZN(n8715)
         );
  OAI21_X1 U10256 ( .B1(n8716), .B2(n8821), .A(n8715), .ZN(P2_U3227) );
  INV_X1 U10257 ( .A(n8718), .ZN(n8719) );
  AOI21_X1 U10258 ( .B1(n8720), .B2(n8717), .A(n8719), .ZN(n8725) );
  AND2_X1 U10259 ( .A1(P2_U3152), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n8860) );
  OAI22_X1 U10260 ( .A1(n9206), .A2(n8786), .B1(n8785), .B2(n8721), .ZN(n8722)
         );
  AOI211_X1 U10261 ( .C1(n8761), .C2(n9166), .A(n8860), .B(n8722), .ZN(n8724)
         );
  NAND2_X1 U10262 ( .A1(n9321), .A2(n8825), .ZN(n8723) );
  OAI211_X1 U10263 ( .C1(n8725), .C2(n8821), .A(n8724), .B(n8723), .ZN(
        P2_U3228) );
  AOI211_X1 U10264 ( .C1(n8728), .C2(n8727), .A(n8821), .B(n8726), .ZN(n8729)
         );
  INV_X1 U10265 ( .A(n8729), .ZN(n8734) );
  AOI22_X1 U10266 ( .A1(n8816), .A2(n8730), .B1(P2_REG3_REG_5__SCAN_IN), .B2(
        P2_U3152), .ZN(n8733) );
  AOI22_X1 U10267 ( .A1(n8761), .A2(n8731), .B1(n8825), .B2(n6717), .ZN(n8732)
         );
  NAND3_X1 U10268 ( .A1(n8734), .A2(n8733), .A3(n8732), .ZN(P2_U3229) );
  XNOR2_X1 U10269 ( .A(n8736), .B(n8735), .ZN(n8740) );
  OAI22_X1 U10270 ( .A1(n8818), .A2(n9154), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9937), .ZN(n8738) );
  OAI22_X1 U10271 ( .A1(n8833), .A2(n8786), .B1(n8785), .B2(n8917), .ZN(n8737)
         );
  AOI211_X1 U10272 ( .C1(n9317), .C2(n8825), .A(n8738), .B(n8737), .ZN(n8739)
         );
  OAI21_X1 U10273 ( .B1(n8740), .B2(n8821), .A(n8739), .ZN(P2_U3230) );
  INV_X1 U10274 ( .A(n8741), .ZN(n8742) );
  NAND2_X1 U10275 ( .A1(n8743), .A2(n8742), .ZN(n8745) );
  XNOR2_X1 U10276 ( .A(n8745), .B(n8744), .ZN(n8746) );
  NAND3_X1 U10277 ( .A1(n8746), .A2(n8826), .A3(n9049), .ZN(n8754) );
  INV_X1 U10278 ( .A(n8746), .ZN(n8748) );
  NAND3_X1 U10279 ( .A1(n8748), .A2(n6894), .A3(n8747), .ZN(n8753) );
  OAI22_X1 U10280 ( .A1(n8818), .A2(n9031), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8749), .ZN(n8751) );
  OAI22_X1 U10281 ( .A1(n9077), .A2(n8786), .B1(n8785), .B2(n9036), .ZN(n8750)
         );
  AOI211_X1 U10282 ( .C1(n9278), .C2(n8825), .A(n8751), .B(n8750), .ZN(n8752)
         );
  NAND3_X1 U10283 ( .A1(n8754), .A2(n8753), .A3(n8752), .ZN(P2_U3231) );
  OAI21_X1 U10284 ( .B1(n8762), .B2(n8756), .A(n8755), .ZN(n8757) );
  NAND2_X1 U10285 ( .A1(n8757), .A2(n6894), .ZN(n8768) );
  AOI22_X1 U10286 ( .A1(n8816), .A2(n8758), .B1(P2_REG3_REG_4__SCAN_IN), .B2(
        P2_U3152), .ZN(n8767) );
  AOI22_X1 U10287 ( .A1(n8761), .A2(n8760), .B1(n8825), .B2(n8759), .ZN(n8766)
         );
  INV_X1 U10288 ( .A(n8762), .ZN(n8764) );
  NAND4_X1 U10289 ( .A1(n8826), .A2(n8764), .A3(n8843), .A4(n8763), .ZN(n8765)
         );
  NAND4_X1 U10290 ( .A1(n8768), .A2(n8767), .A3(n8766), .A4(n8765), .ZN(
        P2_U3232) );
  XNOR2_X1 U10291 ( .A(n8770), .B(n8769), .ZN(n8775) );
  OAI22_X1 U10292 ( .A1(n8818), .A2(n9100), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8771), .ZN(n8773) );
  OAI22_X1 U10293 ( .A1(n8918), .A2(n8786), .B1(n8785), .B2(n9076), .ZN(n8772)
         );
  AOI211_X1 U10294 ( .C1(n9301), .C2(n8825), .A(n8773), .B(n8772), .ZN(n8774)
         );
  OAI21_X1 U10295 ( .B1(n8775), .B2(n8821), .A(n8774), .ZN(P2_U3235) );
  NAND2_X1 U10296 ( .A1(n8777), .A2(n8776), .ZN(n8779) );
  XNOR2_X1 U10297 ( .A(n8779), .B(n8778), .ZN(n8780) );
  NAND3_X1 U10298 ( .A1(n8780), .A2(n8826), .A3(n9048), .ZN(n8791) );
  INV_X1 U10299 ( .A(n8780), .ZN(n8782) );
  NAND3_X1 U10300 ( .A1(n8782), .A2(n6894), .A3(n8781), .ZN(n8790) );
  INV_X1 U10301 ( .A(n9069), .ZN(n8784) );
  OAI22_X1 U10302 ( .A1(n8818), .A2(n8784), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8783), .ZN(n8788) );
  OAI22_X1 U10303 ( .A1(n9076), .A2(n8786), .B1(n8785), .B2(n9077), .ZN(n8787)
         );
  AOI211_X1 U10304 ( .C1(n9291), .C2(n8825), .A(n8788), .B(n8787), .ZN(n8789)
         );
  NAND3_X1 U10305 ( .A1(n8791), .A2(n8790), .A3(n8789), .ZN(P2_U3237) );
  OAI22_X1 U10306 ( .A1(n8793), .A2(n6911), .B1(n8792), .B2(n8821), .ZN(n8796)
         );
  INV_X1 U10307 ( .A(n8794), .ZN(n8795) );
  NAND3_X1 U10308 ( .A1(n8796), .A2(n8795), .A3(n7322), .ZN(n8804) );
  INV_X1 U10309 ( .A(n8797), .ZN(n8799) );
  AOI22_X1 U10310 ( .A1(n8799), .A2(n6894), .B1(n8816), .B2(n8798), .ZN(n8803)
         );
  AOI22_X1 U10311 ( .A1(n8801), .A2(P2_REG3_REG_2__SCAN_IN), .B1(n8825), .B2(
        n8800), .ZN(n8802) );
  NAND3_X1 U10312 ( .A1(n8804), .A2(n8803), .A3(n8802), .ZN(P2_U3239) );
  XNOR2_X1 U10313 ( .A(n8807), .B(n8806), .ZN(n8814) );
  INV_X1 U10314 ( .A(n9131), .ZN(n8811) );
  OR2_X1 U10315 ( .A1(n8918), .A2(n9205), .ZN(n8809) );
  NAND2_X1 U10316 ( .A1(n9175), .A2(n9220), .ZN(n8808) );
  NAND2_X1 U10317 ( .A1(n8809), .A2(n8808), .ZN(n9137) );
  NAND2_X1 U10318 ( .A1(n8816), .A2(n9137), .ZN(n8810) );
  NAND2_X1 U10319 ( .A1(P2_U3152), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n8884) );
  OAI211_X1 U10320 ( .C1(n8818), .C2(n8811), .A(n8810), .B(n8884), .ZN(n8812)
         );
  AOI21_X1 U10321 ( .B1(n9312), .B2(n8825), .A(n8812), .ZN(n8813) );
  OAI21_X1 U10322 ( .B1(n8814), .B2(n8821), .A(n8813), .ZN(P2_U3240) );
  INV_X1 U10323 ( .A(n8815), .ZN(n9187) );
  OAI22_X1 U10324 ( .A1(n8833), .A2(n9205), .B1(n8914), .B2(n9203), .ZN(n9181)
         );
  AOI22_X1 U10325 ( .A1(n8816), .A2(n9181), .B1(P2_REG3_REG_15__SCAN_IN), .B2(
        P2_U3152), .ZN(n8817) );
  OAI21_X1 U10326 ( .B1(n9187), .B2(n8818), .A(n8817), .ZN(n8824) );
  XNOR2_X1 U10327 ( .A(n8820), .B(n8819), .ZN(n8827) );
  NOR3_X1 U10328 ( .A1(n8827), .A2(n8822), .A3(n8821), .ZN(n8823) );
  AOI211_X1 U10329 ( .C1(n9327), .C2(n8825), .A(n8824), .B(n8823), .ZN(n8829)
         );
  INV_X1 U10330 ( .A(n9206), .ZN(n9174) );
  NAND3_X1 U10331 ( .A1(n8827), .A2(n8826), .A3(n9174), .ZN(n8828) );
  NAND2_X1 U10332 ( .A1(n8829), .A2(n8828), .ZN(P2_U3243) );
  MUX2_X1 U10333 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(n8830), .S(P2_U3966), .Z(
        P2_U3583) );
  MUX2_X1 U10334 ( .A(n8941), .B(P2_DATAO_REG_28__SCAN_IN), .S(n8832), .Z(
        P2_U3580) );
  INV_X1 U10335 ( .A(n8928), .ZN(n8966) );
  MUX2_X1 U10336 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n8966), .S(P2_U3966), .Z(
        P2_U3579) );
  MUX2_X1 U10337 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(n8831), .S(P2_U3966), .Z(
        P2_U3578) );
  MUX2_X1 U10338 ( .A(n9049), .B(P2_DATAO_REG_24__SCAN_IN), .S(n8832), .Z(
        P2_U3576) );
  MUX2_X1 U10339 ( .A(n8924), .B(P2_DATAO_REG_23__SCAN_IN), .S(n8832), .Z(
        P2_U3575) );
  MUX2_X1 U10340 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n9048), .S(P2_U3966), .Z(
        P2_U3574) );
  INV_X1 U10341 ( .A(n9076), .ZN(n9107) );
  MUX2_X1 U10342 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n9107), .S(P2_U3966), .Z(
        P2_U3573) );
  MUX2_X1 U10343 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n8921), .S(P2_U3966), .Z(
        P2_U3572) );
  INV_X1 U10344 ( .A(n8918), .ZN(n9106) );
  MUX2_X1 U10345 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n9106), .S(P2_U3966), .Z(
        P2_U3571) );
  MUX2_X1 U10346 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(n9147), .S(P2_U3966), .Z(
        P2_U3570) );
  MUX2_X1 U10347 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n9175), .S(P2_U3966), .Z(
        P2_U3569) );
  INV_X1 U10348 ( .A(n8833), .ZN(n9148) );
  MUX2_X1 U10349 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n9148), .S(P2_U3966), .Z(
        P2_U3568) );
  MUX2_X1 U10350 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(n9174), .S(P2_U3966), .Z(
        P2_U3567) );
  INV_X1 U10351 ( .A(n8914), .ZN(n8834) );
  MUX2_X1 U10352 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(n8834), .S(P2_U3966), .Z(
        P2_U3566) );
  INV_X1 U10353 ( .A(n9204), .ZN(n9223) );
  MUX2_X1 U10354 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(n9223), .S(P2_U3966), .Z(
        P2_U3565) );
  MUX2_X1 U10355 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(n8835), .S(P2_U3966), .Z(
        P2_U3564) );
  MUX2_X1 U10356 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(n9221), .S(P2_U3966), .Z(
        P2_U3563) );
  MUX2_X1 U10357 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(n8836), .S(P2_U3966), .Z(
        P2_U3562) );
  MUX2_X1 U10358 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(n8837), .S(P2_U3966), .Z(
        P2_U3561) );
  MUX2_X1 U10359 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(n8838), .S(P2_U3966), .Z(
        P2_U3560) );
  MUX2_X1 U10360 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(n8839), .S(P2_U3966), .Z(
        P2_U3559) );
  MUX2_X1 U10361 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(n8840), .S(P2_U3966), .Z(
        P2_U3558) );
  MUX2_X1 U10362 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(n8841), .S(P2_U3966), .Z(
        P2_U3557) );
  MUX2_X1 U10363 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(n8842), .S(P2_U3966), .Z(
        P2_U3556) );
  MUX2_X1 U10364 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(n8843), .S(P2_U3966), .Z(
        P2_U3555) );
  MUX2_X1 U10365 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(n4996), .S(P2_U3966), .Z(
        P2_U3554) );
  MUX2_X1 U10366 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(n8844), .S(P2_U3966), .Z(
        P2_U3553) );
  MUX2_X1 U10367 ( .A(P2_DATAO_REG_0__SCAN_IN), .B(n6700), .S(P2_U3966), .Z(
        P2_U3552) );
  OAI211_X1 U10368 ( .C1(n8846), .C2(P2_REG1_REG_15__SCAN_IN), .A(n10505), .B(
        n8845), .ZN(n8856) );
  AND2_X1 U10369 ( .A1(P2_U3152), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n8847) );
  AOI21_X1 U10370 ( .B1(n10508), .B2(P2_ADDR_REG_15__SCAN_IN), .A(n8847), .ZN(
        n8855) );
  OAI21_X1 U10371 ( .B1(n8850), .B2(n8849), .A(n8848), .ZN(n8851) );
  NAND2_X1 U10372 ( .A1(n8851), .A2(n10506), .ZN(n8854) );
  NAND2_X1 U10373 ( .A1(n8870), .A2(n8852), .ZN(n8853) );
  NAND4_X1 U10374 ( .A1(n8856), .A2(n8855), .A3(n8854), .A4(n8853), .ZN(
        P2_U3260) );
  AOI21_X1 U10375 ( .B1(n8859), .B2(n8858), .A(n8857), .ZN(n8872) );
  INV_X1 U10376 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n8862) );
  INV_X1 U10377 ( .A(n8860), .ZN(n8861) );
  OAI21_X1 U10378 ( .B1(n8863), .B2(n8862), .A(n8861), .ZN(n8868) );
  AOI211_X1 U10379 ( .C1(n8866), .C2(n8865), .A(n8864), .B(n10511), .ZN(n8867)
         );
  AOI211_X1 U10380 ( .C1(n8870), .C2(n8869), .A(n8868), .B(n8867), .ZN(n8871)
         );
  OAI21_X1 U10381 ( .B1(n8872), .B2(n10510), .A(n8871), .ZN(P2_U3261) );
  AOI211_X1 U10382 ( .C1(n4446), .C2(n8874), .A(n8873), .B(n10511), .ZN(n8883)
         );
  NOR2_X1 U10383 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9937), .ZN(n8875) );
  AOI21_X1 U10384 ( .B1(n10508), .B2(P2_ADDR_REG_17__SCAN_IN), .A(n8875), .ZN(
        n8880) );
  OAI211_X1 U10385 ( .C1(n8878), .C2(n8877), .A(n10505), .B(n8876), .ZN(n8879)
         );
  OAI211_X1 U10386 ( .C1(n10509), .C2(n8881), .A(n8880), .B(n8879), .ZN(n8882)
         );
  OR2_X1 U10387 ( .A1(n8883), .A2(n8882), .ZN(P2_U3262) );
  INV_X1 U10388 ( .A(n8884), .ZN(n8890) );
  AOI21_X1 U10389 ( .B1(n8887), .B2(n8886), .A(n8885), .ZN(n8888) );
  NOR2_X1 U10390 ( .A1(n10510), .A2(n8888), .ZN(n8889) );
  AOI211_X1 U10391 ( .C1(n10508), .C2(P2_ADDR_REG_18__SCAN_IN), .A(n8890), .B(
        n8889), .ZN(n8896) );
  OAI21_X1 U10392 ( .B1(n8893), .B2(n8892), .A(n8891), .ZN(n8894) );
  NAND2_X1 U10393 ( .A1(n10506), .A2(n8894), .ZN(n8895) );
  OAI211_X1 U10394 ( .C1(n10509), .C2(n8897), .A(n8896), .B(n8895), .ZN(
        P2_U3263) );
  AOI21_X1 U10395 ( .B1(n8901), .B2(n8948), .A(n8900), .ZN(n9238) );
  NAND2_X1 U10396 ( .A1(n9238), .A2(n9234), .ZN(n8904) );
  AOI21_X1 U10397 ( .B1(n4392), .B2(P2_REG2_REG_30__SCAN_IN), .A(n8902), .ZN(
        n8903) );
  OAI211_X1 U10398 ( .C1(n9241), .C2(n10523), .A(n8904), .B(n8903), .ZN(
        P2_U3266) );
  XNOR2_X1 U10399 ( .A(n8905), .B(n6628), .ZN(n8910) );
  NAND2_X1 U10400 ( .A1(n8941), .A2(n9220), .ZN(n8906) );
  OAI21_X1 U10401 ( .B1(n8908), .B2(n8907), .A(n8906), .ZN(n8909) );
  NAND2_X1 U10402 ( .A1(n8911), .A2(n9223), .ZN(n8912) );
  AOI22_X1 U10403 ( .A1(n9164), .A2(n9163), .B1(n9321), .B2(n9148), .ZN(n9151)
         );
  NAND2_X1 U10404 ( .A1(n9151), .A2(n9150), .ZN(n9149) );
  NAND2_X1 U10405 ( .A1(n9117), .A2(n8918), .ZN(n8919) );
  NAND2_X1 U10406 ( .A1(n9307), .A2(n9106), .ZN(n8920) );
  NAND2_X1 U10407 ( .A1(n9286), .A2(n8924), .ZN(n8925) );
  INV_X1 U10408 ( .A(n8925), .ZN(n8926) );
  INV_X1 U10409 ( .A(n9291), .ZN(n9071) );
  NAND2_X1 U10410 ( .A1(n9071), .A2(n9092), .ZN(n9052) );
  NAND2_X1 U10411 ( .A1(n8987), .A2(n8928), .ZN(n8937) );
  INV_X1 U10412 ( .A(n8937), .ZN(n8932) );
  NAND2_X1 U10413 ( .A1(n8929), .A2(n8991), .ZN(n8936) );
  INV_X1 U10414 ( .A(n8936), .ZN(n8930) );
  AND2_X1 U10415 ( .A1(n8989), .A2(n8978), .ZN(n8931) );
  AND2_X1 U10416 ( .A1(n8956), .A2(n8963), .ZN(n8934) );
  AND2_X1 U10417 ( .A1(n8953), .A2(n8934), .ZN(n8933) );
  NAND2_X1 U10418 ( .A1(n8954), .A2(n8933), .ZN(n8940) );
  INV_X1 U10419 ( .A(n8934), .ZN(n8938) );
  NAND2_X1 U10420 ( .A1(n8935), .A2(n9036), .ZN(n8999) );
  AND2_X1 U10421 ( .A1(n8999), .A2(n8936), .ZN(n8979) );
  AND2_X1 U10422 ( .A1(n8979), .A2(n8937), .ZN(n8955) );
  NAND2_X1 U10423 ( .A1(n9253), .A2(n9243), .ZN(n8942) );
  XNOR2_X1 U10424 ( .A(n8942), .B(n6628), .ZN(n8943) );
  NAND2_X1 U10425 ( .A1(n8943), .A2(n9056), .ZN(n8952) );
  OAI22_X1 U10426 ( .A1(n8945), .A2(n9188), .B1(n9060), .B2(n8944), .ZN(n8950)
         );
  NAND2_X1 U10427 ( .A1(n9245), .A2(n8946), .ZN(n8947) );
  NAND2_X1 U10428 ( .A1(n8948), .A2(n8947), .ZN(n9248) );
  NOR2_X1 U10429 ( .A1(n9248), .A2(n8974), .ZN(n8949) );
  AOI211_X1 U10430 ( .C1(n9190), .C2(n9245), .A(n8950), .B(n8949), .ZN(n8951)
         );
  OAI211_X1 U10431 ( .C1(n9250), .C2(n10529), .A(n8952), .B(n8951), .ZN(
        P2_U3267) );
  NAND2_X1 U10432 ( .A1(n9000), .A2(n8955), .ZN(n8957) );
  NAND2_X1 U10433 ( .A1(n8957), .A2(n8956), .ZN(n8959) );
  XNOR2_X1 U10434 ( .A(n8959), .B(n8958), .ZN(n9256) );
  INV_X1 U10435 ( .A(n9256), .ZN(n8977) );
  NAND2_X1 U10436 ( .A1(n8961), .A2(n8960), .ZN(n8988) );
  NAND2_X1 U10437 ( .A1(n8988), .A2(n8980), .ZN(n8994) );
  NAND3_X1 U10438 ( .A1(n8994), .A2(n8963), .A3(n8962), .ZN(n8965) );
  NAND3_X1 U10439 ( .A1(n8965), .A2(n8964), .A3(n9225), .ZN(n8968) );
  NAND2_X1 U10440 ( .A1(n8966), .A2(n9220), .ZN(n8967) );
  XNOR2_X1 U10441 ( .A(n9259), .B(n8981), .ZN(n9257) );
  INV_X1 U10442 ( .A(n8970), .ZN(n8971) );
  AOI22_X1 U10443 ( .A1(n8971), .A2(n10517), .B1(P2_REG2_REG_28__SCAN_IN), 
        .B2(n4392), .ZN(n8973) );
  NAND2_X1 U10444 ( .A1(n9259), .A2(n9190), .ZN(n8972) );
  OAI211_X1 U10445 ( .C1(n9257), .C2(n8974), .A(n8973), .B(n8972), .ZN(n8975)
         );
  AOI21_X1 U10446 ( .B1(n9258), .B2(n9060), .A(n8975), .ZN(n8976) );
  OAI21_X1 U10447 ( .B1(n8977), .B2(n9231), .A(n8976), .ZN(P2_U3268) );
  INV_X1 U10448 ( .A(n9007), .ZN(n8983) );
  INV_X1 U10449 ( .A(n8981), .ZN(n8982) );
  AOI21_X1 U10450 ( .B1(n9261), .B2(n8983), .A(n8982), .ZN(n9262) );
  INV_X1 U10451 ( .A(n8984), .ZN(n8985) );
  AOI22_X1 U10452 ( .A1(n8985), .A2(n10517), .B1(P2_REG2_REG_27__SCAN_IN), 
        .B2(n4392), .ZN(n8986) );
  OAI21_X1 U10453 ( .B1(n8987), .B2(n10523), .A(n8986), .ZN(n8997) );
  INV_X1 U10454 ( .A(n8988), .ZN(n8990) );
  AOI21_X1 U10455 ( .B1(n8990), .B2(n8989), .A(n9200), .ZN(n8995) );
  OAI22_X1 U10456 ( .A1(n8992), .A2(n9205), .B1(n8991), .B2(n9203), .ZN(n8993)
         );
  AOI21_X1 U10457 ( .B1(n8995), .B2(n8994), .A(n8993), .ZN(n9264) );
  NOR2_X1 U10458 ( .A1(n9264), .A2(n4392), .ZN(n8996) );
  AOI211_X1 U10459 ( .C1(n9234), .C2(n9262), .A(n8997), .B(n8996), .ZN(n8998)
         );
  OAI21_X1 U10460 ( .B1(n9265), .B2(n9231), .A(n8998), .ZN(P2_U3269) );
  NAND2_X1 U10461 ( .A1(n9000), .A2(n8999), .ZN(n9001) );
  XNOR2_X1 U10462 ( .A(n9001), .B(n9003), .ZN(n9266) );
  INV_X1 U10463 ( .A(n9266), .ZN(n9015) );
  AOI22_X1 U10464 ( .A1(n9268), .A2(n9190), .B1(n4392), .B2(
        P2_REG2_REG_26__SCAN_IN), .ZN(n9014) );
  XNOR2_X1 U10465 ( .A(n9002), .B(n9003), .ZN(n9004) );
  NAND2_X1 U10466 ( .A1(n9004), .A2(n9225), .ZN(n9270) );
  INV_X1 U10467 ( .A(n9270), .ZN(n9012) );
  NAND2_X1 U10468 ( .A1(n9268), .A2(n9020), .ZN(n9005) );
  NAND2_X1 U10469 ( .A1(n9005), .A2(n9357), .ZN(n9006) );
  OR2_X1 U10470 ( .A1(n9007), .A2(n9006), .ZN(n9271) );
  NAND2_X1 U10471 ( .A1(n9008), .A2(n10517), .ZN(n9009) );
  OAI211_X1 U10472 ( .C1(n9271), .C2(n6625), .A(n9010), .B(n9009), .ZN(n9011)
         );
  OAI21_X1 U10473 ( .B1(n9012), .B2(n9011), .A(n9060), .ZN(n9013) );
  OAI211_X1 U10474 ( .C1(n9015), .C2(n9231), .A(n9014), .B(n9013), .ZN(
        P2_U3270) );
  XNOR2_X1 U10475 ( .A(n8954), .B(n9016), .ZN(n9277) );
  AOI22_X1 U10476 ( .A1(n9275), .A2(n9190), .B1(n10529), .B2(
        P2_REG2_REG_25__SCAN_IN), .ZN(n9025) );
  XNOR2_X1 U10477 ( .A(n9017), .B(n9016), .ZN(n9019) );
  OAI21_X1 U10478 ( .B1(n9019), .B2(n9200), .A(n9018), .ZN(n9273) );
  AOI211_X1 U10479 ( .C1(n9275), .C2(n9028), .A(n10590), .B(n8633), .ZN(n9274)
         );
  INV_X1 U10480 ( .A(n9274), .ZN(n9022) );
  OAI22_X1 U10481 ( .A1(n9022), .A2(n6625), .B1(n9188), .B2(n9021), .ZN(n9023)
         );
  OAI21_X1 U10482 ( .B1(n9273), .B2(n9023), .A(n9060), .ZN(n9024) );
  OAI211_X1 U10483 ( .C1(n9277), .C2(n9231), .A(n9025), .B(n9024), .ZN(
        P2_U3271) );
  AOI21_X1 U10484 ( .B1(n9027), .B2(n9026), .A(n4452), .ZN(n9282) );
  INV_X1 U10485 ( .A(n9057), .ZN(n9030) );
  INV_X1 U10486 ( .A(n9028), .ZN(n9029) );
  AOI21_X1 U10487 ( .B1(n9278), .B2(n9030), .A(n9029), .ZN(n9279) );
  INV_X1 U10488 ( .A(n9031), .ZN(n9032) );
  AOI22_X1 U10489 ( .A1(n4392), .A2(P2_REG2_REG_24__SCAN_IN), .B1(n9032), .B2(
        n10517), .ZN(n9033) );
  OAI21_X1 U10490 ( .B1(n9034), .B2(n10523), .A(n9033), .ZN(n9041) );
  AOI21_X1 U10491 ( .B1(n9035), .B2(n4856), .A(n9200), .ZN(n9039) );
  OAI22_X1 U10492 ( .A1(n9036), .A2(n9205), .B1(n9077), .B2(n9203), .ZN(n9037)
         );
  AOI21_X1 U10493 ( .B1(n9039), .B2(n9038), .A(n9037), .ZN(n9281) );
  NOR2_X1 U10494 ( .A1(n9281), .A2(n4392), .ZN(n9040) );
  AOI211_X1 U10495 ( .C1(n9279), .C2(n9234), .A(n9041), .B(n9040), .ZN(n9042)
         );
  OAI21_X1 U10496 ( .B1(n9282), .B2(n9231), .A(n9042), .ZN(P2_U3272) );
  INV_X1 U10497 ( .A(n9043), .ZN(n9073) );
  OAI21_X1 U10498 ( .B1(n9073), .B2(n9045), .A(n9044), .ZN(n9047) );
  NAND2_X1 U10499 ( .A1(n9047), .A2(n9046), .ZN(n9050) );
  AOI222_X1 U10500 ( .A1(n9225), .A2(n9050), .B1(n9049), .B2(n9222), .C1(n9048), .C2(n9220), .ZN(n9289) );
  NAND2_X1 U10501 ( .A1(n9066), .A2(n9075), .ZN(n9053) );
  NAND2_X1 U10502 ( .A1(n9053), .A2(n9051), .ZN(n9284) );
  NAND2_X1 U10503 ( .A1(n9053), .A2(n9052), .ZN(n9055) );
  NAND2_X1 U10504 ( .A1(n9055), .A2(n9054), .ZN(n9283) );
  NAND3_X1 U10505 ( .A1(n9284), .A2(n9283), .A3(n9056), .ZN(n9064) );
  AOI211_X1 U10506 ( .C1(n9286), .C2(n9067), .A(n10590), .B(n9057), .ZN(n9285)
         );
  NOR2_X1 U10507 ( .A1(n4548), .A2(n10523), .ZN(n9062) );
  OAI22_X1 U10508 ( .A1(n9060), .A2(n9059), .B1(n9058), .B2(n9188), .ZN(n9061)
         );
  AOI211_X1 U10509 ( .C1(n9285), .C2(n9158), .A(n9062), .B(n9061), .ZN(n9063)
         );
  OAI211_X1 U10510 ( .C1(n4392), .C2(n9289), .A(n9064), .B(n9063), .ZN(
        P2_U3273) );
  XNOR2_X1 U10511 ( .A(n9066), .B(n9065), .ZN(n9295) );
  AOI21_X1 U10512 ( .B1(n9291), .B2(n9068), .A(n8632), .ZN(n9292) );
  AOI22_X1 U10513 ( .A1(n4392), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n9069), .B2(
        n10517), .ZN(n9070) );
  OAI21_X1 U10514 ( .B1(n9071), .B2(n10523), .A(n9070), .ZN(n9081) );
  NAND2_X1 U10515 ( .A1(n9090), .A2(n9072), .ZN(n9074) );
  AOI211_X1 U10516 ( .C1(n9075), .C2(n9074), .A(n9200), .B(n9073), .ZN(n9079)
         );
  OAI22_X1 U10517 ( .A1(n9077), .A2(n9205), .B1(n9076), .B2(n9203), .ZN(n9078)
         );
  NOR2_X1 U10518 ( .A1(n9079), .A2(n9078), .ZN(n9294) );
  NOR2_X1 U10519 ( .A1(n9294), .A2(n4392), .ZN(n9080) );
  AOI211_X1 U10520 ( .C1(n9292), .C2(n9234), .A(n9081), .B(n9080), .ZN(n9082)
         );
  OAI21_X1 U10521 ( .B1(n9295), .B2(n9231), .A(n9082), .ZN(P2_U3274) );
  XNOR2_X1 U10522 ( .A(n9083), .B(n9087), .ZN(n9300) );
  XNOR2_X1 U10523 ( .A(n9296), .B(n4485), .ZN(n9297) );
  AOI22_X1 U10524 ( .A1(n4392), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n9084), .B2(
        n10517), .ZN(n9085) );
  OAI21_X1 U10525 ( .B1(n9086), .B2(n10523), .A(n9085), .ZN(n9096) );
  OR2_X1 U10526 ( .A1(n9088), .A2(n9087), .ZN(n9089) );
  NAND2_X1 U10527 ( .A1(n9090), .A2(n9089), .ZN(n9094) );
  OAI22_X1 U10528 ( .A1(n9092), .A2(n9205), .B1(n9091), .B2(n9203), .ZN(n9093)
         );
  AOI21_X1 U10529 ( .B1(n9094), .B2(n9225), .A(n9093), .ZN(n9299) );
  NOR2_X1 U10530 ( .A1(n9299), .A2(n4392), .ZN(n9095) );
  AOI211_X1 U10531 ( .C1(n9297), .C2(n9234), .A(n9096), .B(n9095), .ZN(n9097)
         );
  OAI21_X1 U10532 ( .B1(n9300), .B2(n9231), .A(n9097), .ZN(P2_U3275) );
  XNOR2_X1 U10533 ( .A(n9099), .B(n9098), .ZN(n9305) );
  AOI21_X1 U10534 ( .B1(n9301), .B2(n9113), .A(n4485), .ZN(n9302) );
  INV_X1 U10535 ( .A(n9100), .ZN(n9101) );
  AOI22_X1 U10536 ( .A1(n4392), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n9101), .B2(
        n10517), .ZN(n9102) );
  OAI21_X1 U10537 ( .B1(n4990), .B2(n10523), .A(n9102), .ZN(n9110) );
  OAI21_X1 U10538 ( .B1(n9105), .B2(n9104), .A(n9103), .ZN(n9108) );
  AOI222_X1 U10539 ( .A1(n9225), .A2(n9108), .B1(n9107), .B2(n9222), .C1(n9106), .C2(n9220), .ZN(n9304) );
  NOR2_X1 U10540 ( .A1(n9304), .A2(n4392), .ZN(n9109) );
  AOI211_X1 U10541 ( .C1(n9302), .C2(n9234), .A(n9110), .B(n9109), .ZN(n9111)
         );
  OAI21_X1 U10542 ( .B1(n9305), .B2(n9231), .A(n9111), .ZN(P2_U3276) );
  XOR2_X1 U10543 ( .A(n9112), .B(n9120), .Z(n9310) );
  INV_X1 U10544 ( .A(n9113), .ZN(n9114) );
  AOI211_X1 U10545 ( .C1(n9307), .C2(n9128), .A(n10590), .B(n9114), .ZN(n9306)
         );
  AOI22_X1 U10546 ( .A1(n4392), .A2(P2_REG2_REG_19__SCAN_IN), .B1(n9115), .B2(
        n10517), .ZN(n9116) );
  OAI21_X1 U10547 ( .B1(n9117), .B2(n10523), .A(n9116), .ZN(n9124) );
  OAI21_X1 U10548 ( .B1(n9120), .B2(n9119), .A(n9118), .ZN(n9122) );
  AOI21_X1 U10549 ( .B1(n9122), .B2(n9225), .A(n9121), .ZN(n9309) );
  NOR2_X1 U10550 ( .A1(n9309), .A2(n10529), .ZN(n9123) );
  AOI211_X1 U10551 ( .C1(n9306), .C2(n9158), .A(n9124), .B(n9123), .ZN(n9125)
         );
  OAI21_X1 U10552 ( .B1(n9310), .B2(n9231), .A(n9125), .ZN(P2_U3277) );
  XNOR2_X1 U10553 ( .A(n9126), .B(n9136), .ZN(n9315) );
  INV_X1 U10554 ( .A(n9127), .ZN(n9130) );
  INV_X1 U10555 ( .A(n9128), .ZN(n9129) );
  AOI211_X1 U10556 ( .C1(n9312), .C2(n9130), .A(n10590), .B(n9129), .ZN(n9311)
         );
  AOI22_X1 U10557 ( .A1(n4392), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n9131), .B2(
        n10517), .ZN(n9132) );
  OAI21_X1 U10558 ( .B1(n9133), .B2(n10523), .A(n9132), .ZN(n9140) );
  INV_X1 U10559 ( .A(n9134), .ZN(n9135) );
  XOR2_X1 U10560 ( .A(n9136), .B(n9135), .Z(n9138) );
  AOI21_X1 U10561 ( .B1(n9138), .B2(n9225), .A(n9137), .ZN(n9314) );
  NOR2_X1 U10562 ( .A1(n9314), .A2(n4392), .ZN(n9139) );
  AOI211_X1 U10563 ( .C1(n9311), .C2(n9158), .A(n9140), .B(n9139), .ZN(n9141)
         );
  OAI21_X1 U10564 ( .B1(n9315), .B2(n9231), .A(n9141), .ZN(P2_U3278) );
  NAND2_X1 U10565 ( .A1(n9143), .A2(n9142), .ZN(n9169) );
  NOR2_X1 U10566 ( .A1(n9169), .A2(n9163), .ZN(n9170) );
  NOR2_X1 U10567 ( .A1(n9170), .A2(n9144), .ZN(n9145) );
  XNOR2_X1 U10568 ( .A(n9145), .B(n9150), .ZN(n9146) );
  AOI222_X1 U10569 ( .A1(n9148), .A2(n9220), .B1(n9147), .B2(n9222), .C1(n9225), .C2(n9146), .ZN(n9319) );
  OAI21_X1 U10570 ( .B1(n9151), .B2(n9150), .A(n4547), .ZN(n9152) );
  INV_X1 U10571 ( .A(n9152), .ZN(n9320) );
  NAND2_X1 U10572 ( .A1(n4392), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n9153) );
  OAI21_X1 U10573 ( .B1(n9188), .B2(n9154), .A(n9153), .ZN(n9155) );
  AOI21_X1 U10574 ( .B1(n9317), .B2(n9190), .A(n9155), .ZN(n9160) );
  OAI21_X1 U10575 ( .B1(n9165), .B2(n9156), .A(n9357), .ZN(n9157) );
  NOR2_X1 U10576 ( .A1(n9157), .A2(n9127), .ZN(n9316) );
  NAND2_X1 U10577 ( .A1(n9316), .A2(n9158), .ZN(n9159) );
  OAI211_X1 U10578 ( .C1(n9320), .C2(n9231), .A(n9160), .B(n9159), .ZN(n9161)
         );
  INV_X1 U10579 ( .A(n9161), .ZN(n9162) );
  OAI21_X1 U10580 ( .B1(n4392), .B2(n9319), .A(n9162), .ZN(P2_U3279) );
  XNOR2_X1 U10581 ( .A(n9164), .B(n9163), .ZN(n9325) );
  AOI21_X1 U10582 ( .B1(n9321), .B2(n9191), .A(n9165), .ZN(n9322) );
  INV_X1 U10583 ( .A(n9321), .ZN(n9168) );
  AOI22_X1 U10584 ( .A1(n4392), .A2(P2_REG2_REG_16__SCAN_IN), .B1(n9166), .B2(
        n10517), .ZN(n9167) );
  OAI21_X1 U10585 ( .B1(n9168), .B2(n10523), .A(n9167), .ZN(n9178) );
  INV_X1 U10586 ( .A(n9169), .ZN(n9172) );
  INV_X1 U10587 ( .A(n9170), .ZN(n9171) );
  OAI21_X1 U10588 ( .B1(n9173), .B2(n9172), .A(n9171), .ZN(n9176) );
  AOI222_X1 U10589 ( .A1(n9225), .A2(n9176), .B1(n9175), .B2(n9222), .C1(n9174), .C2(n9220), .ZN(n9324) );
  NOR2_X1 U10590 ( .A1(n9324), .A2(n4392), .ZN(n9177) );
  AOI211_X1 U10591 ( .C1(n9322), .C2(n9234), .A(n9178), .B(n9177), .ZN(n9179)
         );
  OAI21_X1 U10592 ( .B1(n9231), .B2(n9325), .A(n9179), .ZN(P2_U3280) );
  XNOR2_X1 U10593 ( .A(n9180), .B(n5064), .ZN(n9182) );
  AOI21_X1 U10594 ( .B1(n9182), .B2(n9225), .A(n9181), .ZN(n9329) );
  AOI21_X1 U10595 ( .B1(n9185), .B2(n9184), .A(n9183), .ZN(n9330) );
  NAND2_X1 U10596 ( .A1(n4392), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n9186) );
  OAI21_X1 U10597 ( .B1(n9188), .B2(n9187), .A(n9186), .ZN(n9189) );
  AOI21_X1 U10598 ( .B1(n9327), .B2(n9190), .A(n9189), .ZN(n9194) );
  NAND2_X1 U10599 ( .A1(n9209), .A2(n9215), .ZN(n9210) );
  AOI21_X1 U10600 ( .B1(n9210), .B2(n9327), .A(n10590), .ZN(n9192) );
  AND2_X1 U10601 ( .A1(n9192), .A2(n9191), .ZN(n9326) );
  NAND2_X1 U10602 ( .A1(n9326), .A2(n9158), .ZN(n9193) );
  OAI211_X1 U10603 ( .C1(n9330), .C2(n9231), .A(n9194), .B(n9193), .ZN(n9195)
         );
  INV_X1 U10604 ( .A(n9195), .ZN(n9196) );
  OAI21_X1 U10605 ( .B1(n10529), .B2(n9329), .A(n9196), .ZN(P2_U3281) );
  NOR2_X1 U10606 ( .A1(n9197), .A2(n4667), .ZN(n9202) );
  AOI21_X1 U10607 ( .B1(n9201), .B2(n9198), .A(n4798), .ZN(n9199) );
  AOI211_X1 U10608 ( .C1(n9202), .C2(n9201), .A(n9200), .B(n9199), .ZN(n9208)
         );
  OAI22_X1 U10609 ( .A1(n9206), .A2(n9205), .B1(n9204), .B2(n9203), .ZN(n9207)
         );
  NOR2_X1 U10610 ( .A1(n9208), .A2(n9207), .ZN(n9334) );
  INV_X1 U10611 ( .A(n9209), .ZN(n9212) );
  INV_X1 U10612 ( .A(n9210), .ZN(n9211) );
  AOI21_X1 U10613 ( .B1(n9331), .B2(n9212), .A(n9211), .ZN(n9332) );
  AOI22_X1 U10614 ( .A1(n4392), .A2(P2_REG2_REG_14__SCAN_IN), .B1(n9213), .B2(
        n10517), .ZN(n9214) );
  OAI21_X1 U10615 ( .B1(n9215), .B2(n10523), .A(n9214), .ZN(n9217) );
  XNOR2_X1 U10616 ( .A(n4486), .B(n4798), .ZN(n9335) );
  NOR2_X1 U10617 ( .A1(n9335), .A2(n9231), .ZN(n9216) );
  AOI211_X1 U10618 ( .C1(n9332), .C2(n9234), .A(n9217), .B(n9216), .ZN(n9218)
         );
  OAI21_X1 U10619 ( .B1(n9334), .B2(n4392), .A(n9218), .ZN(P2_U3282) );
  XOR2_X1 U10620 ( .A(n9219), .B(n9230), .Z(n9224) );
  AOI222_X1 U10621 ( .A1(n9225), .A2(n9224), .B1(n9223), .B2(n9222), .C1(n9221), .C2(n9220), .ZN(n9345) );
  AOI21_X1 U10622 ( .B1(n9342), .B2(n9226), .A(n4489), .ZN(n9343) );
  AOI22_X1 U10623 ( .A1(n4392), .A2(P2_REG2_REG_12__SCAN_IN), .B1(n9227), .B2(
        n10517), .ZN(n9228) );
  OAI21_X1 U10624 ( .B1(n10523), .B2(n4983), .A(n9228), .ZN(n9233) );
  XOR2_X1 U10625 ( .A(n9229), .B(n9230), .Z(n9346) );
  NOR2_X1 U10626 ( .A1(n9346), .A2(n9231), .ZN(n9232) );
  AOI211_X1 U10627 ( .C1(n9343), .C2(n9234), .A(n9233), .B(n9232), .ZN(n9235)
         );
  OAI21_X1 U10628 ( .B1(n9345), .B2(n4392), .A(n9235), .ZN(P2_U3284) );
  NAND2_X1 U10629 ( .A1(n8630), .A2(n9356), .ZN(n9236) );
  OAI211_X1 U10630 ( .C1(n9237), .C2(n10590), .A(n9239), .B(n9236), .ZN(n9362)
         );
  MUX2_X1 U10631 ( .A(P2_REG1_REG_31__SCAN_IN), .B(n9362), .S(n10605), .Z(
        P2_U3551) );
  NAND2_X1 U10632 ( .A1(n9238), .A2(n9357), .ZN(n9240) );
  OAI211_X1 U10633 ( .C1(n9241), .C2(n10588), .A(n9240), .B(n9239), .ZN(n9363)
         );
  MUX2_X1 U10634 ( .A(P2_REG1_REG_30__SCAN_IN), .B(n9363), .S(n10605), .Z(
        P2_U3550) );
  NAND4_X1 U10635 ( .A1(n9253), .A2(n9242), .A3(n10583), .A4(n9243), .ZN(n9255) );
  INV_X1 U10636 ( .A(n9243), .ZN(n9244) );
  NAND3_X1 U10637 ( .A1(n6628), .A2(n9244), .A3(n10583), .ZN(n9247) );
  NAND2_X1 U10638 ( .A1(n9245), .A2(n9356), .ZN(n9246) );
  OAI211_X1 U10639 ( .C1(n10590), .C2(n9248), .A(n9247), .B(n9246), .ZN(n9249)
         );
  INV_X1 U10640 ( .A(n9249), .ZN(n9251) );
  NAND2_X1 U10641 ( .A1(n6628), .A2(n10583), .ZN(n9252) );
  NAND3_X1 U10642 ( .A1(n9255), .A2(n5090), .A3(n9254), .ZN(n9364) );
  MUX2_X1 U10643 ( .A(P2_REG1_REG_29__SCAN_IN), .B(n9364), .S(n10605), .Z(
        P2_U3549) );
  NAND2_X1 U10644 ( .A1(n9256), .A2(n10583), .ZN(n9260) );
  AOI22_X1 U10645 ( .A1(n9262), .A2(n9357), .B1(n9356), .B2(n9261), .ZN(n9263)
         );
  MUX2_X1 U10646 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n9366), .S(n10605), .Z(
        P2_U3547) );
  AOI21_X1 U10647 ( .B1(n9268), .B2(n9356), .A(n9267), .ZN(n9269) );
  MUX2_X1 U10648 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n9367), .S(n10605), .Z(
        P2_U3546) );
  AOI211_X1 U10649 ( .C1(n9356), .C2(n9275), .A(n9274), .B(n9273), .ZN(n9276)
         );
  OAI21_X1 U10650 ( .B1(n9277), .B2(n9350), .A(n9276), .ZN(n9368) );
  MUX2_X1 U10651 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n9368), .S(n10605), .Z(
        P2_U3545) );
  AOI22_X1 U10652 ( .A1(n9279), .A2(n9357), .B1(n9356), .B2(n9278), .ZN(n9280)
         );
  OAI211_X1 U10653 ( .C1(n9282), .C2(n9350), .A(n9281), .B(n9280), .ZN(n9369)
         );
  MUX2_X1 U10654 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n9369), .S(n10605), .Z(
        P2_U3544) );
  NAND3_X1 U10655 ( .A1(n9284), .A2(n9283), .A3(n10583), .ZN(n9290) );
  AOI21_X1 U10656 ( .B1(n9287), .B2(n9286), .A(n9285), .ZN(n9288) );
  NAND3_X1 U10657 ( .A1(n9290), .A2(n9289), .A3(n9288), .ZN(n9370) );
  MUX2_X1 U10658 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n9370), .S(n10605), .Z(
        P2_U3543) );
  AOI22_X1 U10659 ( .A1(n9292), .A2(n9357), .B1(n9356), .B2(n9291), .ZN(n9293)
         );
  OAI211_X1 U10660 ( .C1(n9295), .C2(n9350), .A(n9294), .B(n9293), .ZN(n9371)
         );
  MUX2_X1 U10661 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n9371), .S(n10605), .Z(
        P2_U3542) );
  AOI22_X1 U10662 ( .A1(n9297), .A2(n9357), .B1(n9356), .B2(n9296), .ZN(n9298)
         );
  OAI211_X1 U10663 ( .C1(n9300), .C2(n9350), .A(n9299), .B(n9298), .ZN(n9372)
         );
  MUX2_X1 U10664 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n9372), .S(n10605), .Z(
        P2_U3541) );
  AOI22_X1 U10665 ( .A1(n9302), .A2(n9357), .B1(n9356), .B2(n9301), .ZN(n9303)
         );
  OAI211_X1 U10666 ( .C1(n9305), .C2(n9350), .A(n9304), .B(n9303), .ZN(n9373)
         );
  MUX2_X1 U10667 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n9373), .S(n10605), .Z(
        P2_U3540) );
  AOI21_X1 U10668 ( .B1(n9356), .B2(n9307), .A(n9306), .ZN(n9308) );
  OAI211_X1 U10669 ( .C1(n9310), .C2(n9350), .A(n9309), .B(n9308), .ZN(n9374)
         );
  MUX2_X1 U10670 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n9374), .S(n10605), .Z(
        P2_U3539) );
  AOI21_X1 U10671 ( .B1(n9356), .B2(n9312), .A(n9311), .ZN(n9313) );
  OAI211_X1 U10672 ( .C1(n9315), .C2(n9350), .A(n9314), .B(n9313), .ZN(n9375)
         );
  MUX2_X1 U10673 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n9375), .S(n10605), .Z(
        P2_U3538) );
  AOI21_X1 U10674 ( .B1(n9356), .B2(n9317), .A(n9316), .ZN(n9318) );
  OAI211_X1 U10675 ( .C1(n9320), .C2(n9350), .A(n9319), .B(n9318), .ZN(n9376)
         );
  MUX2_X1 U10676 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n9376), .S(n10605), .Z(
        P2_U3537) );
  AOI22_X1 U10677 ( .A1(n9322), .A2(n9357), .B1(n9356), .B2(n9321), .ZN(n9323)
         );
  OAI211_X1 U10678 ( .C1(n9325), .C2(n9350), .A(n9324), .B(n9323), .ZN(n9377)
         );
  MUX2_X1 U10679 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n9377), .S(n10605), .Z(
        P2_U3536) );
  AOI21_X1 U10680 ( .B1(n9356), .B2(n9327), .A(n9326), .ZN(n9328) );
  OAI211_X1 U10681 ( .C1(n9330), .C2(n9350), .A(n9329), .B(n9328), .ZN(n9378)
         );
  MUX2_X1 U10682 ( .A(P2_REG1_REG_15__SCAN_IN), .B(n9378), .S(n10605), .Z(
        P2_U3535) );
  AOI22_X1 U10683 ( .A1(n9332), .A2(n9357), .B1(n9356), .B2(n9331), .ZN(n9333)
         );
  OAI211_X1 U10684 ( .C1(n9350), .C2(n9335), .A(n9334), .B(n9333), .ZN(n9379)
         );
  MUX2_X1 U10685 ( .A(P2_REG1_REG_14__SCAN_IN), .B(n9379), .S(n10605), .Z(
        P2_U3534) );
  NOR2_X1 U10686 ( .A1(n9336), .A2(n9350), .ZN(n9341) );
  OAI22_X1 U10687 ( .A1(n9338), .A2(n10590), .B1(n9337), .B2(n10588), .ZN(
        n9339) );
  MUX2_X1 U10688 ( .A(n9380), .B(P2_REG1_REG_13__SCAN_IN), .S(n10603), .Z(
        P2_U3533) );
  AOI22_X1 U10689 ( .A1(n9343), .A2(n9357), .B1(n9356), .B2(n9342), .ZN(n9344)
         );
  OAI211_X1 U10690 ( .C1(n9350), .C2(n9346), .A(n9345), .B(n9344), .ZN(n9381)
         );
  MUX2_X1 U10691 ( .A(P2_REG1_REG_12__SCAN_IN), .B(n9381), .S(n10605), .Z(
        P2_U3532) );
  AOI22_X1 U10692 ( .A1(n9348), .A2(n9357), .B1(n9356), .B2(n9347), .ZN(n9349)
         );
  OAI21_X1 U10693 ( .B1(n9351), .B2(n9350), .A(n9349), .ZN(n9352) );
  OR2_X1 U10694 ( .A1(n9353), .A2(n9352), .ZN(n9382) );
  MUX2_X1 U10695 ( .A(n9382), .B(P2_REG1_REG_11__SCAN_IN), .S(n10603), .Z(
        P2_U3531) );
  INV_X1 U10696 ( .A(n9354), .ZN(n9361) );
  AOI22_X1 U10697 ( .A1(n9358), .A2(n9357), .B1(n9356), .B2(n9355), .ZN(n9359)
         );
  OAI211_X1 U10698 ( .C1(n9361), .C2(n10586), .A(n9360), .B(n9359), .ZN(n9383)
         );
  MUX2_X1 U10699 ( .A(P2_REG1_REG_9__SCAN_IN), .B(n9383), .S(n10605), .Z(
        P2_U3529) );
  MUX2_X1 U10700 ( .A(P2_REG0_REG_31__SCAN_IN), .B(n9362), .S(n10598), .Z(
        P2_U3519) );
  MUX2_X1 U10701 ( .A(P2_REG0_REG_30__SCAN_IN), .B(n9363), .S(n10598), .Z(
        P2_U3518) );
  MUX2_X1 U10702 ( .A(P2_REG0_REG_29__SCAN_IN), .B(n9364), .S(n10598), .Z(
        P2_U3517) );
  MUX2_X1 U10703 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n9365), .S(n10598), .Z(
        P2_U3516) );
  MUX2_X1 U10704 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n9367), .S(n10598), .Z(
        P2_U3514) );
  MUX2_X1 U10705 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n9368), .S(n10598), .Z(
        P2_U3513) );
  MUX2_X1 U10706 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n9369), .S(n10598), .Z(
        P2_U3512) );
  MUX2_X1 U10707 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n9370), .S(n10598), .Z(
        P2_U3511) );
  MUX2_X1 U10708 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n9371), .S(n10598), .Z(
        P2_U3510) );
  MUX2_X1 U10709 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n9372), .S(n10598), .Z(
        P2_U3509) );
  MUX2_X1 U10710 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n9373), .S(n10598), .Z(
        P2_U3508) );
  MUX2_X1 U10711 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n9374), .S(n10598), .Z(
        P2_U3507) );
  MUX2_X1 U10712 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n9375), .S(n10598), .Z(
        P2_U3505) );
  MUX2_X1 U10713 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n9376), .S(n10598), .Z(
        P2_U3502) );
  MUX2_X1 U10714 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n9377), .S(n10598), .Z(
        P2_U3499) );
  MUX2_X1 U10715 ( .A(P2_REG0_REG_15__SCAN_IN), .B(n9378), .S(n10598), .Z(
        P2_U3496) );
  MUX2_X1 U10716 ( .A(P2_REG0_REG_14__SCAN_IN), .B(n9379), .S(n10598), .Z(
        P2_U3493) );
  MUX2_X1 U10717 ( .A(n9380), .B(P2_REG0_REG_13__SCAN_IN), .S(n10596), .Z(
        P2_U3490) );
  MUX2_X1 U10718 ( .A(P2_REG0_REG_12__SCAN_IN), .B(n9381), .S(n10598), .Z(
        P2_U3487) );
  MUX2_X1 U10719 ( .A(n9382), .B(P2_REG0_REG_11__SCAN_IN), .S(n10596), .Z(
        P2_U3484) );
  MUX2_X1 U10720 ( .A(P2_REG0_REG_9__SCAN_IN), .B(n9383), .S(n10598), .Z(
        P2_U3478) );
  INV_X1 U10721 ( .A(n9384), .ZN(n10284) );
  NOR4_X1 U10722 ( .A1(n9385), .A2(P2_IR_REG_30__SCAN_IN), .A3(P2_U3152), .A4(
        n6170), .ZN(n9387) );
  AOI21_X1 U10723 ( .B1(n9388), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n9387), .ZN(
        n9389) );
  OAI21_X1 U10724 ( .B1(n10284), .B2(n9399), .A(n9389), .ZN(P2_U3327) );
  OAI222_X1 U10725 ( .A1(n9395), .A2(n9391), .B1(n9399), .B2(n9390), .C1(
        P2_U3152), .C2(n4679), .ZN(P2_U3328) );
  NAND2_X1 U10726 ( .A1(n10288), .A2(n9392), .ZN(n9394) );
  OAI211_X1 U10727 ( .C1(n9395), .C2(n9806), .A(n9394), .B(n9393), .ZN(
        P2_U3330) );
  OAI222_X1 U10728 ( .A1(n9399), .A2(n9398), .B1(n9397), .B2(P2_U3152), .C1(
        n9396), .C2(n9395), .ZN(P2_U3331) );
  MUX2_X1 U10729 ( .A(n9400), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3358) );
  XNOR2_X1 U10730 ( .A(n9402), .B(n9401), .ZN(n9403) );
  XNOR2_X1 U10731 ( .A(n9404), .B(n9403), .ZN(n9410) );
  OAI22_X1 U10732 ( .A1(n9699), .A2(n9494), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9405), .ZN(n9406) );
  AOI21_X1 U10733 ( .B1(n9667), .B2(n9560), .A(n9406), .ZN(n9407) );
  OAI21_X1 U10734 ( .B1(n9671), .B2(n9555), .A(n9407), .ZN(n9408) );
  AOI21_X1 U10735 ( .B1(n10178), .B2(n9518), .A(n9408), .ZN(n9409) );
  OAI21_X1 U10736 ( .B1(n9410), .B2(n9520), .A(n9409), .ZN(P1_U3212) );
  INV_X1 U10737 ( .A(n9412), .ZN(n9417) );
  AOI21_X1 U10738 ( .B1(n9413), .B2(n9412), .A(n9411), .ZN(n9414) );
  NOR2_X1 U10739 ( .A1(n9414), .A2(n9520), .ZN(n9415) );
  OAI21_X1 U10740 ( .B1(n9417), .B2(n9416), .A(n9415), .ZN(n9422) );
  NOR2_X1 U10741 ( .A1(n9766), .A2(P1_STATE_REG_SCAN_IN), .ZN(n10333) );
  AOI21_X1 U10742 ( .B1(n9553), .B2(n9579), .A(n10333), .ZN(n9418) );
  OAI21_X1 U10743 ( .B1(n10155), .B2(n9555), .A(n9418), .ZN(n9419) );
  AOI21_X1 U10744 ( .B1(n9420), .B2(n9560), .A(n9419), .ZN(n9421) );
  OAI211_X1 U10745 ( .C1(n9423), .C2(n9556), .A(n9422), .B(n9421), .ZN(
        P1_U3213) );
  NAND2_X1 U10746 ( .A1(n9425), .A2(n9424), .ZN(n9427) );
  INV_X1 U10747 ( .A(n9486), .ZN(n9428) );
  NAND2_X1 U10748 ( .A1(n9427), .A2(n9426), .ZN(n9487) );
  NAND2_X1 U10749 ( .A1(n9428), .A2(n9487), .ZN(n9429) );
  XNOR2_X1 U10750 ( .A(n9429), .B(n9485), .ZN(n9435) );
  NOR2_X1 U10751 ( .A1(n9542), .A2(n10017), .ZN(n9432) );
  OAI22_X1 U10752 ( .A1(n10042), .A2(n9494), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9430), .ZN(n9431) );
  AOI211_X1 U10753 ( .C1(n9570), .C2(n9534), .A(n9432), .B(n9431), .ZN(n9434)
         );
  NAND2_X1 U10754 ( .A1(n10201), .A2(n9518), .ZN(n9433) );
  OAI211_X1 U10755 ( .C1(n9435), .C2(n9520), .A(n9434), .B(n9433), .ZN(
        P1_U3214) );
  NAND2_X1 U10756 ( .A1(n9436), .A2(n9437), .ZN(n9510) );
  NOR2_X1 U10757 ( .A1(n9436), .A2(n9437), .ZN(n9512) );
  AOI21_X1 U10758 ( .B1(n9513), .B2(n9510), .A(n9512), .ZN(n9442) );
  OAI21_X1 U10759 ( .B1(n9440), .B2(n9439), .A(n9438), .ZN(n9441) );
  XNOR2_X1 U10760 ( .A(n9442), .B(n9441), .ZN(n9447) );
  NAND2_X1 U10761 ( .A1(n9553), .A2(n9574), .ZN(n9443) );
  NAND2_X1 U10762 ( .A1(P1_U3084), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n9633) );
  OAI211_X1 U10763 ( .C1(n10091), .C2(n9555), .A(n9443), .B(n9633), .ZN(n9445)
         );
  NOR2_X1 U10764 ( .A1(n10098), .A2(n9556), .ZN(n9444) );
  AOI211_X1 U10765 ( .C1(n10095), .C2(n9560), .A(n9445), .B(n9444), .ZN(n9446)
         );
  OAI21_X1 U10766 ( .B1(n9447), .B2(n9520), .A(n9446), .ZN(P1_U3217) );
  NAND2_X1 U10767 ( .A1(n9448), .A2(n9501), .ZN(n9449) );
  XOR2_X1 U10768 ( .A(n9450), .B(n9449), .Z(n9456) );
  AOI22_X1 U10769 ( .A1(n10022), .A2(n9534), .B1(P1_REG3_REG_21__SCAN_IN), 
        .B2(P1_U3084), .ZN(n9451) );
  OAI21_X1 U10770 ( .B1(n10091), .B2(n9494), .A(n9451), .ZN(n9454) );
  NAND2_X1 U10771 ( .A1(n10061), .A2(n10240), .ZN(n10207) );
  NOR2_X1 U10772 ( .A1(n10207), .A2(n9452), .ZN(n9453) );
  AOI211_X1 U10773 ( .C1(n10052), .C2(n9560), .A(n9454), .B(n9453), .ZN(n9455)
         );
  OAI21_X1 U10774 ( .B1(n9456), .B2(n9520), .A(n9455), .ZN(P1_U3221) );
  XOR2_X1 U10775 ( .A(n9458), .B(n9457), .Z(n9463) );
  AOI22_X1 U10776 ( .A1(n9706), .A2(n9560), .B1(P1_REG3_REG_25__SCAN_IN), .B2(
        P1_U3084), .ZN(n9460) );
  NAND2_X1 U10777 ( .A1(n9570), .A2(n9553), .ZN(n9459) );
  OAI211_X1 U10778 ( .C1(n9699), .C2(n9555), .A(n9460), .B(n9459), .ZN(n9461)
         );
  AOI21_X1 U10779 ( .B1(n10190), .B2(n9518), .A(n9461), .ZN(n9462) );
  OAI21_X1 U10780 ( .B1(n9463), .B2(n9520), .A(n9462), .ZN(P1_U3223) );
  XNOR2_X1 U10781 ( .A(n9474), .B(n9470), .ZN(n9464) );
  XNOR2_X1 U10782 ( .A(n9472), .B(n9464), .ZN(n9469) );
  AND2_X1 U10783 ( .A1(P1_U3084), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n10361) );
  NOR2_X1 U10784 ( .A1(n9494), .A2(n10155), .ZN(n9465) );
  AOI211_X1 U10785 ( .C1(n9534), .C2(n10104), .A(n10361), .B(n9465), .ZN(n9466) );
  OAI21_X1 U10786 ( .B1(n9542), .B2(n10146), .A(n9466), .ZN(n9467) );
  AOI21_X1 U10787 ( .B1(n10230), .B2(n9518), .A(n9467), .ZN(n9468) );
  OAI21_X1 U10788 ( .B1(n9469), .B2(n9520), .A(n9468), .ZN(P1_U3224) );
  INV_X1 U10789 ( .A(n9472), .ZN(n9475) );
  OAI21_X1 U10790 ( .B1(n9472), .B2(n9471), .A(n9470), .ZN(n9473) );
  OAI21_X1 U10791 ( .B1(n9475), .B2(n9474), .A(n9473), .ZN(n9479) );
  XNOR2_X1 U10792 ( .A(n9477), .B(n9476), .ZN(n9478) );
  XNOR2_X1 U10793 ( .A(n9479), .B(n9478), .ZN(n9484) );
  NAND2_X1 U10794 ( .A1(n9553), .A2(n9575), .ZN(n9480) );
  NAND2_X1 U10795 ( .A1(P1_U3084), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n10373)
         );
  OAI211_X1 U10796 ( .C1(n10133), .C2(n9555), .A(n9480), .B(n10373), .ZN(n9481) );
  AOI21_X1 U10797 ( .B1(n10137), .B2(n9560), .A(n9481), .ZN(n9483) );
  NAND2_X1 U10798 ( .A1(n10226), .A2(n9518), .ZN(n9482) );
  OAI211_X1 U10799 ( .C1(n9484), .C2(n9520), .A(n9483), .B(n9482), .ZN(
        P1_U3226) );
  INV_X1 U10800 ( .A(n9485), .ZN(n9488) );
  AOI21_X1 U10801 ( .B1(n9488), .B2(n9487), .A(n9486), .ZN(n9491) );
  OAI21_X1 U10802 ( .B1(n9491), .B2(n9490), .A(n9489), .ZN(n9492) );
  NAND2_X1 U10803 ( .A1(n9492), .A2(n9547), .ZN(n9498) );
  OAI22_X1 U10804 ( .A1(n9721), .A2(n9494), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9493), .ZN(n9496) );
  NOR2_X1 U10805 ( .A1(n9722), .A2(n9555), .ZN(n9495) );
  AOI211_X1 U10806 ( .C1(n9723), .C2(n9560), .A(n9496), .B(n9495), .ZN(n9497)
         );
  INV_X1 U10807 ( .A(n9501), .ZN(n9499) );
  NOR2_X1 U10808 ( .A1(n9448), .A2(n9499), .ZN(n9504) );
  AOI21_X1 U10809 ( .B1(n9502), .B2(n9501), .A(n9500), .ZN(n9503) );
  OAI21_X1 U10810 ( .B1(n9504), .B2(n9503), .A(n9547), .ZN(n9509) );
  OAI22_X1 U10811 ( .A1(n10074), .A2(n9555), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9505), .ZN(n9507) );
  NOR2_X1 U10812 ( .A1(n9542), .A2(n10066), .ZN(n9506) );
  AOI211_X1 U10813 ( .C1(n9553), .C2(n10071), .A(n9507), .B(n9506), .ZN(n9508)
         );
  OAI211_X1 U10814 ( .C1(n4897), .C2(n9556), .A(n9509), .B(n9508), .ZN(
        P1_U3231) );
  INV_X1 U10815 ( .A(n9510), .ZN(n9511) );
  NOR2_X1 U10816 ( .A1(n9512), .A2(n9511), .ZN(n9514) );
  XNOR2_X1 U10817 ( .A(n9514), .B(n9513), .ZN(n9521) );
  NAND2_X1 U10818 ( .A1(P1_U3084), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n10387)
         );
  OAI21_X1 U10819 ( .B1(n9555), .B2(n10107), .A(n10387), .ZN(n9515) );
  AOI21_X1 U10820 ( .B1(n9553), .B2(n10104), .A(n9515), .ZN(n9516) );
  OAI21_X1 U10821 ( .B1(n9542), .B2(n10115), .A(n9516), .ZN(n9517) );
  AOI21_X1 U10822 ( .B1(n10114), .B2(n9518), .A(n9517), .ZN(n9519) );
  OAI21_X1 U10823 ( .B1(n9521), .B2(n9520), .A(n9519), .ZN(P1_U3236) );
  AOI21_X1 U10824 ( .B1(n9524), .B2(n9523), .A(n9522), .ZN(n9528) );
  XNOR2_X1 U10825 ( .A(n9526), .B(n9525), .ZN(n9527) );
  XNOR2_X1 U10826 ( .A(n9528), .B(n9527), .ZN(n9529) );
  NAND2_X1 U10827 ( .A1(n9529), .A2(n9547), .ZN(n9538) );
  AOI21_X1 U10828 ( .B1(n9553), .B2(n9586), .A(n9530), .ZN(n9537) );
  AND2_X1 U10829 ( .A1(n9531), .A2(n10240), .ZN(n10459) );
  AOI22_X1 U10830 ( .A1(n9560), .A2(n9533), .B1(n9532), .B2(n10459), .ZN(n9536) );
  NAND2_X1 U10831 ( .A1(n9534), .A2(n4756), .ZN(n9535) );
  NAND4_X1 U10832 ( .A1(n9538), .A2(n9537), .A3(n9536), .A4(n9535), .ZN(
        P1_U3237) );
  INV_X1 U10833 ( .A(n9690), .ZN(n10256) );
  OAI211_X1 U10834 ( .C1(n9541), .C2(n9540), .A(n9539), .B(n9547), .ZN(n9546)
         );
  OAI22_X1 U10835 ( .A1(n9680), .A2(n9542), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9802), .ZN(n9544) );
  NOR2_X1 U10836 ( .A1(n9687), .A2(n9555), .ZN(n9543) );
  AOI211_X1 U10837 ( .C1(n9553), .C2(n9569), .A(n9544), .B(n9543), .ZN(n9545)
         );
  OAI211_X1 U10838 ( .C1(n10256), .C2(n9556), .A(n9546), .B(n9545), .ZN(
        P1_U3238) );
  INV_X1 U10839 ( .A(n9552), .ZN(n9549) );
  OAI21_X1 U10840 ( .B1(n9549), .B2(n9548), .A(n9547), .ZN(n9564) );
  AOI21_X1 U10841 ( .B1(n9552), .B2(n9551), .A(n9550), .ZN(n9563) );
  NAND2_X1 U10842 ( .A1(n9553), .A2(n9578), .ZN(n9554) );
  NAND2_X1 U10843 ( .A1(P1_U3084), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n10347)
         );
  OAI211_X1 U10844 ( .C1(n10132), .C2(n9555), .A(n9554), .B(n10347), .ZN(n9559) );
  NOR2_X1 U10845 ( .A1(n9557), .A2(n9556), .ZN(n9558) );
  AOI211_X1 U10846 ( .C1(n9561), .C2(n9560), .A(n9559), .B(n9558), .ZN(n9562)
         );
  OAI21_X1 U10847 ( .B1(n9564), .B2(n9563), .A(n9562), .ZN(P1_U3239) );
  MUX2_X1 U10848 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n9565), .S(P1_U4006), .Z(
        P1_U3585) );
  MUX2_X1 U10849 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n9566), .S(P1_U4006), .Z(
        P1_U3583) );
  MUX2_X1 U10850 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n9567), .S(P1_U4006), .Z(
        P1_U3582) );
  MUX2_X1 U10851 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n9568), .S(P1_U4006), .Z(
        P1_U3581) );
  MUX2_X1 U10852 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n9569), .S(P1_U4006), .Z(
        P1_U3580) );
  MUX2_X1 U10853 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n9570), .S(P1_U4006), .Z(
        P1_U3579) );
  MUX2_X1 U10854 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n9571), .S(P1_U4006), .Z(
        P1_U3578) );
  MUX2_X1 U10855 ( .A(n10022), .B(P1_DATAO_REG_22__SCAN_IN), .S(n9576), .Z(
        P1_U3577) );
  MUX2_X1 U10856 ( .A(n9572), .B(P1_DATAO_REG_21__SCAN_IN), .S(n9576), .Z(
        P1_U3576) );
  MUX2_X1 U10857 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n9573), .S(P1_U4006), .Z(
        P1_U3575) );
  MUX2_X1 U10858 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n10071), .S(P1_U4006), .Z(
        P1_U3574) );
  MUX2_X1 U10859 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n9574), .S(P1_U4006), .Z(
        P1_U3573) );
  MUX2_X1 U10860 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n10104), .S(P1_U4006), .Z(
        P1_U3572) );
  MUX2_X1 U10861 ( .A(n9575), .B(P1_DATAO_REG_16__SCAN_IN), .S(n9576), .Z(
        P1_U3571) );
  MUX2_X1 U10862 ( .A(n9577), .B(P1_DATAO_REG_15__SCAN_IN), .S(n9576), .Z(
        P1_U3570) );
  MUX2_X1 U10863 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n9578), .S(P1_U4006), .Z(
        P1_U3569) );
  MUX2_X1 U10864 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n9579), .S(P1_U4006), .Z(
        P1_U3568) );
  MUX2_X1 U10865 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n9580), .S(P1_U4006), .Z(
        P1_U3567) );
  MUX2_X1 U10866 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n9581), .S(P1_U4006), .Z(
        P1_U3566) );
  MUX2_X1 U10867 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n9582), .S(P1_U4006), .Z(
        P1_U3565) );
  MUX2_X1 U10868 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n9583), .S(P1_U4006), .Z(
        P1_U3564) );
  MUX2_X1 U10869 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n9584), .S(P1_U4006), .Z(
        P1_U3563) );
  MUX2_X1 U10870 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n4756), .S(P1_U4006), .Z(
        P1_U3562) );
  MUX2_X1 U10871 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n9585), .S(P1_U4006), .Z(
        P1_U3561) );
  MUX2_X1 U10872 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n9586), .S(P1_U4006), .Z(
        P1_U3560) );
  MUX2_X1 U10873 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n9587), .S(P1_U4006), .Z(
        P1_U3559) );
  MUX2_X1 U10874 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n9588), .S(P1_U4006), .Z(
        P1_U3558) );
  MUX2_X1 U10875 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n9589), .S(P1_U4006), .Z(
        P1_U3557) );
  MUX2_X1 U10876 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n5737), .S(P1_U4006), .Z(
        P1_U3556) );
  MUX2_X1 U10877 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(n9590), .S(P1_U4006), .Z(
        P1_U3555) );
  MUX2_X1 U10878 ( .A(n7065), .B(P1_REG2_REG_5__SCAN_IN), .S(n9595), .Z(n9593)
         );
  INV_X1 U10879 ( .A(n9591), .ZN(n9592) );
  AOI211_X1 U10880 ( .C1(n4500), .C2(n9593), .A(n9592), .B(n10357), .ZN(n9594)
         );
  AOI21_X1 U10881 ( .B1(n10363), .B2(n9595), .A(n9594), .ZN(n9601) );
  NAND2_X1 U10882 ( .A1(n10319), .A2(P1_ADDR_REG_5__SCAN_IN), .ZN(n9599) );
  OAI211_X1 U10883 ( .C1(n4501), .C2(n9597), .A(n10395), .B(n9596), .ZN(n9598)
         );
  NAND4_X1 U10884 ( .A1(n9601), .A2(n9600), .A3(n9599), .A4(n9598), .ZN(
        P1_U3246) );
  NAND2_X1 U10885 ( .A1(n9602), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n9603) );
  NAND2_X1 U10886 ( .A1(n9604), .A2(n9603), .ZN(n9605) );
  NOR2_X1 U10887 ( .A1(n9605), .A2(n10334), .ZN(n9606) );
  INV_X1 U10888 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n10331) );
  NOR2_X1 U10889 ( .A1(n9608), .A2(n9621), .ZN(n9610) );
  INV_X1 U10890 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n10343) );
  XNOR2_X1 U10891 ( .A(n10346), .B(n9609), .ZN(n10344) );
  NOR2_X1 U10892 ( .A1(n9610), .A2(n10342), .ZN(n10359) );
  XNOR2_X1 U10893 ( .A(n10362), .B(P1_REG2_REG_16__SCAN_IN), .ZN(n10358) );
  NAND2_X1 U10894 ( .A1(n10362), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n9611) );
  NAND2_X1 U10895 ( .A1(n10355), .A2(n9611), .ZN(n10372) );
  XNOR2_X1 U10896 ( .A(n9626), .B(n10128), .ZN(n10371) );
  NAND2_X1 U10897 ( .A1(n10372), .A2(n10371), .ZN(n10370) );
  NAND2_X1 U10898 ( .A1(n9626), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n9612) );
  NAND2_X1 U10899 ( .A1(n10370), .A2(n9612), .ZN(n10386) );
  MUX2_X1 U10900 ( .A(P1_REG2_REG_18__SCAN_IN), .B(n10116), .S(n9627), .Z(
        n10385) );
  NAND2_X1 U10901 ( .A1(n10386), .A2(n10385), .ZN(n10384) );
  NAND2_X1 U10902 ( .A1(n9627), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n9613) );
  NAND2_X1 U10903 ( .A1(n10384), .A2(n9613), .ZN(n9615) );
  AOI21_X1 U10904 ( .B1(n9618), .B2(n9617), .A(n9616), .ZN(n10336) );
  XNOR2_X1 U10905 ( .A(n9619), .B(n9864), .ZN(n10335) );
  NOR2_X1 U10906 ( .A1(n10336), .A2(n10335), .ZN(n10338) );
  NAND2_X1 U10907 ( .A1(n10346), .A2(n9620), .ZN(n9622) );
  INV_X1 U10908 ( .A(n10365), .ZN(n9624) );
  XNOR2_X1 U10909 ( .A(n10362), .B(P1_REG1_REG_16__SCAN_IN), .ZN(n10364) );
  INV_X1 U10910 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n10234) );
  INV_X1 U10911 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n9625) );
  XNOR2_X1 U10912 ( .A(n9626), .B(n9625), .ZN(n10378) );
  NOR2_X1 U10913 ( .A1(n9627), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n9628) );
  AOI21_X1 U10914 ( .B1(n9627), .B2(P1_REG1_REG_18__SCAN_IN), .A(n9628), .ZN(
        n10393) );
  XOR2_X1 U10915 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n9629), .Z(n9631) );
  OAI211_X1 U10916 ( .C1(n9635), .C2(n10399), .A(n9634), .B(n9633), .ZN(
        P1_U3260) );
  XNOR2_X1 U10917 ( .A(n9645), .B(n9642), .ZN(n9638) );
  INV_X1 U10918 ( .A(n9639), .ZN(n9640) );
  NAND2_X1 U10919 ( .A1(n9641), .A2(n9640), .ZN(n10172) );
  NOR2_X1 U10920 ( .A1(n10123), .A2(n10172), .ZN(n9648) );
  AOI21_X1 U10921 ( .B1(n10123), .B2(P1_REG2_REG_31__SCAN_IN), .A(n9648), .ZN(
        n9644) );
  NAND2_X1 U10922 ( .A1(n9642), .A2(n10150), .ZN(n9643) );
  OAI211_X1 U10923 ( .C1(n10166), .C2(n9659), .A(n9644), .B(n9643), .ZN(
        P1_U3261) );
  NAND2_X1 U10924 ( .A1(n10174), .A2(n10422), .ZN(n9650) );
  AOI21_X1 U10925 ( .B1(n10123), .B2(P1_REG2_REG_30__SCAN_IN), .A(n9648), .ZN(
        n9649) );
  OAI211_X1 U10926 ( .C1(n9636), .C2(n10400), .A(n9650), .B(n9649), .ZN(
        P1_U3262) );
  INV_X1 U10927 ( .A(n9651), .ZN(n9664) );
  NAND2_X1 U10928 ( .A1(n9653), .A2(n9652), .ZN(n9654) );
  XNOR2_X1 U10929 ( .A(n9654), .B(n4709), .ZN(n9662) );
  INV_X1 U10930 ( .A(P1_REG2_REG_29__SCAN_IN), .ZN(n9655) );
  OAI22_X1 U10931 ( .A1(n9656), .A2(n10145), .B1(n9655), .B2(n10148), .ZN(
        n9657) );
  AOI21_X1 U10932 ( .B1(n6058), .B2(n10150), .A(n9657), .ZN(n9658) );
  OAI21_X1 U10933 ( .B1(n9660), .B2(n9659), .A(n9658), .ZN(n9661) );
  AOI21_X1 U10934 ( .B1(n9662), .B2(n10424), .A(n9661), .ZN(n9663) );
  OAI21_X1 U10935 ( .B1(n9664), .B2(n10123), .A(n9663), .ZN(P1_U3355) );
  AOI211_X1 U10936 ( .C1(n10178), .C2(n9691), .A(n10158), .B(n9666), .ZN(
        n10177) );
  AOI22_X1 U10937 ( .A1(n9667), .A2(n10411), .B1(P1_REG2_REG_27__SCAN_IN), 
        .B2(n10123), .ZN(n9668) );
  OAI21_X1 U10938 ( .B1(n4903), .B2(n10400), .A(n9668), .ZN(n9676) );
  AOI21_X1 U10939 ( .B1(n9670), .B2(n9669), .A(n10406), .ZN(n9674) );
  OAI22_X1 U10940 ( .A1(n9671), .A2(n10405), .B1(n9699), .B2(n10403), .ZN(
        n9672) );
  AOI21_X1 U10941 ( .B1(n9674), .B2(n9673), .A(n9672), .ZN(n10180) );
  NOR2_X1 U10942 ( .A1(n10180), .A2(n10123), .ZN(n9675) );
  AOI211_X1 U10943 ( .C1(n10422), .C2(n10177), .A(n9676), .B(n9675), .ZN(n9677) );
  OAI21_X1 U10944 ( .B1(n10142), .B2(n10181), .A(n9677), .ZN(P1_U3264) );
  XNOR2_X1 U10945 ( .A(n9678), .B(n9683), .ZN(n10182) );
  NAND2_X1 U10946 ( .A1(n10182), .A2(n10424), .ZN(n9696) );
  OAI22_X1 U10947 ( .A1(n9680), .A2(n10145), .B1(n9679), .B2(n10148), .ZN(
        n9681) );
  AOI21_X1 U10948 ( .B1(n9690), .B2(n10150), .A(n9681), .ZN(n9695) );
  NAND2_X1 U10949 ( .A1(n9701), .A2(n9682), .ZN(n9684) );
  NAND2_X1 U10950 ( .A1(n9684), .A2(n9683), .ZN(n9686) );
  AOI21_X1 U10951 ( .B1(n9686), .B2(n9685), .A(n10406), .ZN(n9689) );
  OAI22_X1 U10952 ( .A1(n9687), .A2(n10405), .B1(n9722), .B2(n10403), .ZN(
        n9688) );
  NAND2_X1 U10953 ( .A1(n10184), .A2(n10148), .ZN(n9694) );
  AOI21_X1 U10954 ( .B1(n9690), .B2(n9703), .A(n10158), .ZN(n9692) );
  AND2_X1 U10955 ( .A1(n9692), .A2(n9691), .ZN(n10183) );
  NAND2_X1 U10956 ( .A1(n10183), .A2(n10422), .ZN(n9693) );
  NAND4_X1 U10957 ( .A1(n9696), .A2(n9695), .A3(n9694), .A4(n9693), .ZN(
        P1_U3265) );
  AOI21_X1 U10958 ( .B1(n9698), .B2(n9697), .A(n10406), .ZN(n9702) );
  OAI22_X1 U10959 ( .A1(n9699), .A2(n10405), .B1(n10025), .B2(n10403), .ZN(
        n9700) );
  AOI21_X1 U10960 ( .B1(n9702), .B2(n9701), .A(n9700), .ZN(n10192) );
  INV_X1 U10961 ( .A(n9732), .ZN(n9705) );
  INV_X1 U10962 ( .A(n9703), .ZN(n9704) );
  AOI211_X1 U10963 ( .C1(n10190), .C2(n9705), .A(n10158), .B(n9704), .ZN(
        n10189) );
  AOI22_X1 U10964 ( .A1(n9706), .A2(n10411), .B1(P1_REG2_REG_25__SCAN_IN), 
        .B2(n10123), .ZN(n9707) );
  OAI21_X1 U10965 ( .B1(n9708), .B2(n10400), .A(n9707), .ZN(n9713) );
  INV_X1 U10966 ( .A(n9709), .ZN(n9710) );
  AOI21_X1 U10967 ( .B1(n5994), .B2(n9711), .A(n9710), .ZN(n10193) );
  NOR2_X1 U10968 ( .A1(n10193), .A2(n10142), .ZN(n9712) );
  AOI211_X1 U10969 ( .C1(n10189), .C2(n10422), .A(n9713), .B(n9712), .ZN(n9714) );
  OAI21_X1 U10970 ( .B1(n10123), .B2(n10192), .A(n9714), .ZN(P1_U3266) );
  INV_X1 U10971 ( .A(n9715), .ZN(n9719) );
  AOI21_X1 U10972 ( .B1(n9716), .B2(n9717), .A(n9727), .ZN(n9718) );
  NOR2_X1 U10973 ( .A1(n9719), .A2(n9718), .ZN(n9720) );
  OAI222_X1 U10974 ( .A1(n10405), .A2(n9722), .B1(n10403), .B2(n9721), .C1(
        n9720), .C2(n10406), .ZN(n10194) );
  NAND2_X1 U10975 ( .A1(n10194), .A2(n10148), .ZN(n9737) );
  NAND2_X1 U10976 ( .A1(n9723), .A2(n10411), .ZN(n9724) );
  OAI21_X1 U10977 ( .B1(n10148), .B2(n9725), .A(n9724), .ZN(n9726) );
  AOI21_X1 U10978 ( .B1(n9729), .B2(n10150), .A(n9726), .ZN(n9736) );
  XNOR2_X1 U10979 ( .A(n9728), .B(n9727), .ZN(n10196) );
  NAND2_X1 U10980 ( .A1(n10196), .A2(n10424), .ZN(n9735) );
  NAND2_X1 U10981 ( .A1(n9729), .A2(n10013), .ZN(n9730) );
  NAND2_X1 U10982 ( .A1(n9730), .A2(n10418), .ZN(n9731) );
  NOR2_X1 U10983 ( .A1(n9732), .A2(n9731), .ZN(n10195) );
  AND2_X1 U10984 ( .A1(n10148), .A2(n9733), .ZN(n10119) );
  NAND2_X1 U10985 ( .A1(n10195), .A2(n10119), .ZN(n9734) );
  NAND4_X1 U10986 ( .A1(n9737), .A2(n9736), .A3(n9735), .A4(n9734), .ZN(
        P1_U3267) );
  NOR4_X1 U10987 ( .A1(P2_DATAO_REG_18__SCAN_IN), .A2(P2_DATAO_REG_20__SCAN_IN), .A3(P1_DATAO_REG_17__SCAN_IN), .A4(n9948), .ZN(n9761) );
  NOR4_X1 U10988 ( .A1(P1_DATAO_REG_22__SCAN_IN), .A2(P1_DATAO_REG_21__SCAN_IN), .A3(P2_DATAO_REG_21__SCAN_IN), .A4(n9816), .ZN(n9760) );
  NOR4_X1 U10989 ( .A1(n10234), .A2(n9864), .A3(P2_DATAO_REG_2__SCAN_IN), .A4(
        P1_REG2_REG_13__SCAN_IN), .ZN(n9738) );
  NAND3_X1 U10990 ( .A1(n9738), .A2(P1_DATAO_REG_3__SCAN_IN), .A3(
        P1_REG0_REG_18__SCAN_IN), .ZN(n9746) );
  INV_X1 U10991 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n10301) );
  NOR4_X1 U10992 ( .A1(P1_REG2_REG_12__SCAN_IN), .A2(P1_REG1_REG_7__SCAN_IN), 
        .A3(n10301), .A4(n10502), .ZN(n9744) );
  NOR4_X1 U10993 ( .A1(P1_DATAO_REG_15__SCAN_IN), .A2(P2_DATAO_REG_14__SCAN_IN), .A3(SI_12_), .A4(n9873), .ZN(n9740) );
  NOR4_X1 U10994 ( .A1(P1_REG2_REG_7__SCAN_IN), .A2(P1_REG2_REG_6__SCAN_IN), 
        .A3(P1_REG1_REG_2__SCAN_IN), .A4(n7050), .ZN(n9739) );
  NAND4_X1 U10995 ( .A1(n9741), .A2(P2_DATAO_REG_7__SCAN_IN), .A3(n9740), .A4(
        n9739), .ZN(n9742) );
  NOR3_X1 U10996 ( .A1(n9742), .A2(n9936), .A3(P1_DATAO_REG_6__SCAN_IN), .ZN(
        n9743) );
  NAND2_X1 U10997 ( .A1(n9744), .A2(n9743), .ZN(n9745) );
  NOR4_X1 U10998 ( .A1(SI_5_), .A2(SI_4_), .A3(n9746), .A4(n9745), .ZN(n9759)
         );
  NOR4_X1 U10999 ( .A1(P2_REG0_REG_3__SCAN_IN), .A2(P2_REG2_REG_8__SCAN_IN), 
        .A3(P2_REG0_REG_22__SCAN_IN), .A4(n9876), .ZN(n9748) );
  NAND3_X1 U11000 ( .A1(SI_29_), .A2(n9748), .A3(n9747), .ZN(n9757) );
  INV_X1 U11001 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n9911) );
  NAND4_X1 U11002 ( .A1(P2_D_REG_7__SCAN_IN), .A2(P2_REG0_REG_18__SCAN_IN), 
        .A3(P2_REG1_REG_24__SCAN_IN), .A4(n9911), .ZN(n9749) );
  NOR3_X1 U11003 ( .A1(P2_D_REG_22__SCAN_IN), .A2(P2_REG1_REG_17__SCAN_IN), 
        .A3(n9749), .ZN(n9755) );
  INV_X1 U11004 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n9879) );
  NAND4_X1 U11005 ( .A1(P1_REG2_REG_28__SCAN_IN), .A2(P2_IR_REG_26__SCAN_IN), 
        .A3(P2_D_REG_11__SCAN_IN), .A4(n9879), .ZN(n9753) );
  NAND4_X1 U11006 ( .A1(P2_REG3_REG_21__SCAN_IN), .A2(P1_REG2_REG_26__SCAN_IN), 
        .A3(P2_REG3_REG_3__SCAN_IN), .A4(n9924), .ZN(n9752) );
  NAND4_X1 U11007 ( .A1(P2_REG3_REG_25__SCAN_IN), .A2(P2_IR_REG_27__SCAN_IN), 
        .A3(P2_REG3_REG_17__SCAN_IN), .A4(n10167), .ZN(n9751) );
  NAND4_X1 U11008 ( .A1(P2_REG0_REG_27__SCAN_IN), .A2(P2_REG3_REG_19__SCAN_IN), 
        .A3(P2_REG2_REG_14__SCAN_IN), .A4(n7672), .ZN(n9750) );
  NOR4_X1 U11009 ( .A1(n9753), .A2(n9752), .A3(n9751), .A4(n9750), .ZN(n9754)
         );
  NAND4_X1 U11010 ( .A1(P2_IR_REG_18__SCAN_IN), .A2(P2_D_REG_14__SCAN_IN), 
        .A3(n9755), .A4(n9754), .ZN(n9756) );
  NOR4_X1 U11011 ( .A1(P2_IR_REG_20__SCAN_IN), .A2(n9950), .A3(n9757), .A4(
        n9756), .ZN(n9758) );
  NAND4_X1 U11012 ( .A1(n9761), .A2(n9760), .A3(n9759), .A4(n9758), .ZN(n9789)
         );
  INV_X1 U11013 ( .A(n10649), .ZN(n9762) );
  NAND4_X1 U11014 ( .A1(n9763), .A2(P2_REG1_REG_12__SCAN_IN), .A3(n9762), .A4(
        n10361), .ZN(n9770) );
  NOR2_X1 U11015 ( .A1(P1_WR_REG_SCAN_IN), .A2(P2_WR_REG_SCAN_IN), .ZN(n9765)
         );
  INV_X1 U11016 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n9895) );
  NOR4_X1 U11017 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P1_ADDR_REG_2__SCAN_IN), 
        .A3(P2_ADDR_REG_18__SCAN_IN), .A4(n9895), .ZN(n9764) );
  NAND4_X1 U11018 ( .A1(n9765), .A2(P1_ADDR_REG_4__SCAN_IN), .A3(
        P2_ADDR_REG_3__SCAN_IN), .A4(n9764), .ZN(n9769) );
  NAND4_X1 U11019 ( .A1(P1_REG3_REG_12__SCAN_IN), .A2(P1_REG3_REG_17__SCAN_IN), 
        .A3(n9766), .A4(n9824), .ZN(n9768) );
  NAND4_X1 U11020 ( .A1(P1_IR_REG_24__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .A3(P1_REG3_REG_7__SCAN_IN), .A4(P1_REG3_REG_9__SCAN_IN), .ZN(n9767)
         );
  NOR4_X1 U11021 ( .A1(n9770), .A2(n9769), .A3(n9768), .A4(n9767), .ZN(n9787)
         );
  NAND4_X1 U11022 ( .A1(P1_REG3_REG_25__SCAN_IN), .A2(P1_REG3_REG_28__SCAN_IN), 
        .A3(P2_D_REG_4__SCAN_IN), .A4(n8944), .ZN(n9771) );
  NOR3_X1 U11023 ( .A1(P2_REG0_REG_17__SCAN_IN), .A2(P2_REG2_REG_12__SCAN_IN), 
        .A3(n9771), .ZN(n9786) );
  NOR4_X1 U11024 ( .A1(P2_IR_REG_4__SCAN_IN), .A2(P2_IR_REG_25__SCAN_IN), .A3(
        P2_IR_REG_29__SCAN_IN), .A4(P1_REG2_REG_0__SCAN_IN), .ZN(n9773) );
  NOR2_X1 U11025 ( .A1(n9889), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n9772) );
  NAND4_X1 U11026 ( .A1(n9773), .A2(P2_REG3_REG_14__SCAN_IN), .A3(
        P2_REG1_REG_11__SCAN_IN), .A4(n9772), .ZN(n9784) );
  NOR4_X1 U11027 ( .A1(P1_REG3_REG_26__SCAN_IN), .A2(P1_REG3_REG_27__SCAN_IN), 
        .A3(P2_D_REG_3__SCAN_IN), .A4(n9806), .ZN(n9774) );
  NAND3_X1 U11028 ( .A1(P1_REG2_REG_30__SCAN_IN), .A2(n9774), .A3(n9059), .ZN(
        n9783) );
  NAND4_X1 U11029 ( .A1(P2_REG0_REG_14__SCAN_IN), .A2(P2_REG1_REG_10__SCAN_IN), 
        .A3(P2_REG2_REG_5__SCAN_IN), .A4(n6381), .ZN(n9782) );
  NAND4_X1 U11030 ( .A1(n9939), .A2(P2_D_REG_10__SCAN_IN), .A3(
        P1_D_REG_7__SCAN_IN), .A4(P1_D_REG_13__SCAN_IN), .ZN(n9780) );
  NAND4_X1 U11031 ( .A1(n9775), .A2(SI_25_), .A3(P1_IR_REG_16__SCAN_IN), .A4(
        P1_REG3_REG_0__SCAN_IN), .ZN(n9779) );
  NOR4_X1 U11032 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .A3(
        P1_IR_REG_10__SCAN_IN), .A4(P1_IR_REG_25__SCAN_IN), .ZN(n9776) );
  NAND4_X1 U11033 ( .A1(P1_IR_REG_28__SCAN_IN), .A2(n9776), .A3(n7045), .A4(
        P2_ADDR_REG_15__SCAN_IN), .ZN(n9778) );
  INV_X1 U11034 ( .A(P1_D_REG_26__SCAN_IN), .ZN(n9777) );
  OR4_X1 U11035 ( .A1(n9780), .A2(n9779), .A3(n9778), .A4(n9777), .ZN(n9781)
         );
  NOR4_X1 U11036 ( .A1(n9784), .A2(n9783), .A3(n9782), .A4(n9781), .ZN(n9785)
         );
  NAND3_X1 U11037 ( .A1(n9787), .A2(n9786), .A3(n9785), .ZN(n9788) );
  OAI21_X1 U11038 ( .B1(n9789), .B2(n9788), .A(P1_DATAO_REG_26__SCAN_IN), .ZN(
        n10011) );
  AOI22_X1 U11039 ( .A1(n10502), .A2(keyinput79), .B1(n9791), .B2(keyinput102), 
        .ZN(n9790) );
  OAI221_X1 U11040 ( .B1(n10502), .B2(keyinput79), .C1(n9791), .C2(keyinput102), .A(n9790), .ZN(n9800) );
  INV_X1 U11041 ( .A(P1_D_REG_21__SCAN_IN), .ZN(n10430) );
  INV_X1 U11042 ( .A(P1_D_REG_13__SCAN_IN), .ZN(n10431) );
  AOI22_X1 U11043 ( .A1(n10430), .A2(keyinput120), .B1(keyinput66), .B2(n10431), .ZN(n9792) );
  OAI221_X1 U11044 ( .B1(n10430), .B2(keyinput120), .C1(n10431), .C2(
        keyinput66), .A(n9792), .ZN(n9799) );
  AOI22_X1 U11045 ( .A1(n10167), .A2(keyinput41), .B1(n9794), .B2(keyinput26), 
        .ZN(n9793) );
  OAI221_X1 U11046 ( .B1(n10167), .B2(keyinput41), .C1(n9794), .C2(keyinput26), 
        .A(n9793), .ZN(n9798) );
  INV_X1 U11047 ( .A(P1_D_REG_11__SCAN_IN), .ZN(n10432) );
  AOI22_X1 U11048 ( .A1(n10432), .A2(keyinput40), .B1(keyinput24), .B2(n9796), 
        .ZN(n9795) );
  OAI221_X1 U11049 ( .B1(n10432), .B2(keyinput40), .C1(n9796), .C2(keyinput24), 
        .A(n9795), .ZN(n9797) );
  NOR4_X1 U11050 ( .A1(n9800), .A2(n9799), .A3(n9798), .A4(n9797), .ZN(n9814)
         );
  AOI22_X1 U11051 ( .A1(n9803), .A2(keyinput17), .B1(n9802), .B2(keyinput20), 
        .ZN(n9801) );
  OAI221_X1 U11052 ( .B1(n9803), .B2(keyinput17), .C1(n9802), .C2(keyinput20), 
        .A(n9801), .ZN(n9812) );
  AOI22_X1 U11053 ( .A1(n9806), .A2(keyinput9), .B1(keyinput77), .B2(n9805), 
        .ZN(n9804) );
  OAI221_X1 U11054 ( .B1(n9806), .B2(keyinput9), .C1(n9805), .C2(keyinput77), 
        .A(n9804), .ZN(n9811) );
  AOI22_X1 U11055 ( .A1(n9777), .A2(keyinput42), .B1(keyinput54), .B2(n5285), 
        .ZN(n9807) );
  OAI221_X1 U11056 ( .B1(n9777), .B2(keyinput42), .C1(n5285), .C2(keyinput54), 
        .A(n9807), .ZN(n9810) );
  AOI22_X1 U11057 ( .A1(n10561), .A2(keyinput56), .B1(n9405), .B2(keyinput28), 
        .ZN(n9808) );
  OAI221_X1 U11058 ( .B1(n10561), .B2(keyinput56), .C1(n9405), .C2(keyinput28), 
        .A(n9808), .ZN(n9809) );
  NOR4_X1 U11059 ( .A1(n9812), .A2(n9811), .A3(n9810), .A4(n9809), .ZN(n9813)
         );
  NAND2_X1 U11060 ( .A1(n9814), .A2(n9813), .ZN(n10010) );
  AOI22_X1 U11061 ( .A1(n9817), .A2(keyinput43), .B1(n9816), .B2(keyinput38), 
        .ZN(n9815) );
  OAI221_X1 U11062 ( .B1(n9817), .B2(keyinput43), .C1(n9816), .C2(keyinput38), 
        .A(n9815), .ZN(n9822) );
  INV_X1 U11063 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n9820) );
  AOI22_X1 U11064 ( .A1(n9820), .A2(keyinput108), .B1(n9819), .B2(keyinput10), 
        .ZN(n9818) );
  OAI221_X1 U11065 ( .B1(n9820), .B2(keyinput108), .C1(n9819), .C2(keyinput10), 
        .A(n9818), .ZN(n9821) );
  NOR2_X1 U11066 ( .A1(n9822), .A2(n9821), .ZN(n9852) );
  AOI22_X1 U11067 ( .A1(n9825), .A2(keyinput97), .B1(n9824), .B2(keyinput92), 
        .ZN(n9823) );
  OAI221_X1 U11068 ( .B1(n9825), .B2(keyinput97), .C1(n9824), .C2(keyinput92), 
        .A(n9823), .ZN(n9829) );
  INV_X1 U11069 ( .A(P1_WR_REG_SCAN_IN), .ZN(n10304) );
  AOI22_X1 U11070 ( .A1(n10304), .A2(keyinput116), .B1(n9827), .B2(keyinput93), 
        .ZN(n9826) );
  OAI221_X1 U11071 ( .B1(n10304), .B2(keyinput116), .C1(n9827), .C2(keyinput93), .A(n9826), .ZN(n9828) );
  NOR2_X1 U11072 ( .A1(n9829), .A2(n9828), .ZN(n9851) );
  XNOR2_X1 U11073 ( .A(SI_12_), .B(keyinput121), .ZN(n9833) );
  XNOR2_X1 U11074 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(keyinput21), .ZN(n9832)
         );
  XNOR2_X1 U11075 ( .A(SI_4_), .B(keyinput119), .ZN(n9831) );
  XNOR2_X1 U11076 ( .A(P1_IR_REG_0__SCAN_IN), .B(keyinput88), .ZN(n9830) );
  NAND4_X1 U11077 ( .A1(n9833), .A2(n9832), .A3(n9831), .A4(n9830), .ZN(n9838)
         );
  XNOR2_X1 U11078 ( .A(SI_5_), .B(keyinput46), .ZN(n9835) );
  XNOR2_X1 U11079 ( .A(keyinput0), .B(P2_REG2_REG_29__SCAN_IN), .ZN(n9834) );
  OAI211_X1 U11080 ( .C1(keyinput35), .C2(n9836), .A(n9835), .B(n9834), .ZN(
        n9837) );
  NOR2_X1 U11081 ( .A1(n9838), .A2(n9837), .ZN(n9850) );
  XNOR2_X1 U11082 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(keyinput3), .ZN(n9842) );
  XNOR2_X1 U11083 ( .A(P1_IR_REG_3__SCAN_IN), .B(keyinput125), .ZN(n9841) );
  XNOR2_X1 U11084 ( .A(P1_IR_REG_25__SCAN_IN), .B(keyinput78), .ZN(n9840) );
  XNOR2_X1 U11085 ( .A(P1_IR_REG_10__SCAN_IN), .B(keyinput122), .ZN(n9839) );
  NAND4_X1 U11086 ( .A1(n9842), .A2(n9841), .A3(n9840), .A4(n9839), .ZN(n9848)
         );
  XNOR2_X1 U11087 ( .A(P1_REG1_REG_2__SCAN_IN), .B(keyinput11), .ZN(n9846) );
  XNOR2_X1 U11088 ( .A(P1_REG0_REG_18__SCAN_IN), .B(keyinput114), .ZN(n9845)
         );
  XNOR2_X1 U11089 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(keyinput29), .ZN(n9844) );
  XNOR2_X1 U11090 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(keyinput32), .ZN(n9843) );
  NAND4_X1 U11091 ( .A1(n9846), .A2(n9845), .A3(n9844), .A4(n9843), .ZN(n9847)
         );
  NOR2_X1 U11092 ( .A1(n9848), .A2(n9847), .ZN(n9849) );
  AND4_X1 U11093 ( .A1(n9852), .A2(n9851), .A3(n9850), .A4(n9849), .ZN(n9871)
         );
  AOI22_X1 U11094 ( .A1(n6147), .A2(keyinput31), .B1(n7045), .B2(keyinput12), 
        .ZN(n9853) );
  OAI221_X1 U11095 ( .B1(n6147), .B2(keyinput31), .C1(n7045), .C2(keyinput12), 
        .A(n9853), .ZN(n9857) );
  AOI22_X1 U11096 ( .A1(n9775), .A2(keyinput65), .B1(keyinput126), .B2(n9855), 
        .ZN(n9854) );
  OAI221_X1 U11097 ( .B1(n9775), .B2(keyinput65), .C1(n9855), .C2(keyinput126), 
        .A(n9854), .ZN(n9856) );
  NOR2_X1 U11098 ( .A1(n9857), .A2(n9856), .ZN(n9870) );
  AOI22_X1 U11099 ( .A1(n9860), .A2(keyinput25), .B1(keyinput117), .B2(n9859), 
        .ZN(n9858) );
  OAI221_X1 U11100 ( .B1(n9860), .B2(keyinput25), .C1(n9859), .C2(keyinput117), 
        .A(n9858), .ZN(n9868) );
  AOI22_X1 U11101 ( .A1(n9059), .A2(keyinput124), .B1(n9862), .B2(keyinput105), 
        .ZN(n9861) );
  OAI221_X1 U11102 ( .B1(n9059), .B2(keyinput124), .C1(n9862), .C2(keyinput105), .A(n9861), .ZN(n9867) );
  INV_X1 U11103 ( .A(P1_REG2_REG_30__SCAN_IN), .ZN(n9865) );
  AOI22_X1 U11104 ( .A1(n9865), .A2(keyinput1), .B1(n9864), .B2(keyinput94), 
        .ZN(n9863) );
  OAI221_X1 U11105 ( .B1(n9865), .B2(keyinput1), .C1(n9864), .C2(keyinput94), 
        .A(n9863), .ZN(n9866) );
  NOR3_X1 U11106 ( .A1(n9868), .A2(n9867), .A3(n9866), .ZN(n9869) );
  NAND3_X1 U11107 ( .A1(n9871), .A2(n9870), .A3(n9869), .ZN(n9909) );
  AOI22_X1 U11108 ( .A1(n9873), .A2(keyinput86), .B1(keyinput47), .B2(n5632), 
        .ZN(n9872) );
  OAI221_X1 U11109 ( .B1(n9873), .B2(keyinput86), .C1(n5632), .C2(keyinput47), 
        .A(n9872), .ZN(n9882) );
  AOI22_X1 U11110 ( .A1(n9876), .A2(keyinput30), .B1(keyinput5), .B2(n9875), 
        .ZN(n9874) );
  OAI221_X1 U11111 ( .B1(n9876), .B2(keyinput30), .C1(n9875), .C2(keyinput5), 
        .A(n9874), .ZN(n9881) );
  AOI22_X1 U11112 ( .A1(n9879), .A2(keyinput100), .B1(keyinput103), .B2(n9878), 
        .ZN(n9877) );
  OAI221_X1 U11113 ( .B1(n9879), .B2(keyinput100), .C1(n9878), .C2(keyinput103), .A(n9877), .ZN(n9880) );
  NOR3_X1 U11114 ( .A1(n9882), .A2(n9881), .A3(n9880), .ZN(n9907) );
  INV_X1 U11115 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n9884) );
  AOI22_X1 U11116 ( .A1(n9884), .A2(keyinput81), .B1(n7067), .B2(keyinput96), 
        .ZN(n9883) );
  OAI221_X1 U11117 ( .B1(n9884), .B2(keyinput81), .C1(n7067), .C2(keyinput96), 
        .A(n9883), .ZN(n9893) );
  AOI22_X1 U11118 ( .A1(n9887), .A2(keyinput39), .B1(keyinput68), .B2(n9886), 
        .ZN(n9885) );
  OAI221_X1 U11119 ( .B1(n9887), .B2(keyinput39), .C1(n9886), .C2(keyinput68), 
        .A(n9885), .ZN(n9892) );
  AOI22_X1 U11120 ( .A1(n9890), .A2(keyinput52), .B1(keyinput127), .B2(n9889), 
        .ZN(n9888) );
  OAI221_X1 U11121 ( .B1(n9890), .B2(keyinput52), .C1(n9889), .C2(keyinput127), 
        .A(n9888), .ZN(n9891) );
  NOR3_X1 U11122 ( .A1(n9893), .A2(n9892), .A3(n9891), .ZN(n9906) );
  AOI22_X1 U11123 ( .A1(n10650), .A2(keyinput64), .B1(keyinput4), .B2(n9895), 
        .ZN(n9894) );
  OAI221_X1 U11124 ( .B1(n10650), .B2(keyinput64), .C1(n9895), .C2(keyinput4), 
        .A(n9894), .ZN(n9898) );
  INV_X1 U11125 ( .A(P2_D_REG_7__SCAN_IN), .ZN(n10557) );
  INV_X1 U11126 ( .A(P2_D_REG_14__SCAN_IN), .ZN(n10550) );
  AOI22_X1 U11127 ( .A1(n10557), .A2(keyinput51), .B1(keyinput18), .B2(n10550), 
        .ZN(n9896) );
  OAI221_X1 U11128 ( .B1(n10557), .B2(keyinput51), .C1(n10550), .C2(keyinput18), .A(n9896), .ZN(n9897) );
  NOR2_X1 U11129 ( .A1(n9898), .A2(n9897), .ZN(n9905) );
  AOI22_X1 U11130 ( .A1(n9900), .A2(keyinput107), .B1(keyinput111), .B2(n10553), .ZN(n9899) );
  OAI221_X1 U11131 ( .B1(n9900), .B2(keyinput107), .C1(n10553), .C2(
        keyinput111), .A(n9899), .ZN(n9903) );
  AOI22_X1 U11132 ( .A1(n5318), .A2(keyinput36), .B1(keyinput95), .B2(n10560), 
        .ZN(n9901) );
  OAI221_X1 U11133 ( .B1(n5318), .B2(keyinput36), .C1(n10560), .C2(keyinput95), 
        .A(n9901), .ZN(n9902) );
  NOR2_X1 U11134 ( .A1(n9903), .A2(n9902), .ZN(n9904) );
  NAND4_X1 U11135 ( .A1(n9907), .A2(n9906), .A3(n9905), .A4(n9904), .ZN(n9908)
         );
  NOR2_X1 U11136 ( .A1(n9909), .A2(n9908), .ZN(n10008) );
  AOI22_X1 U11137 ( .A1(n9911), .A2(keyinput101), .B1(keyinput76), .B2(n7221), 
        .ZN(n9910) );
  OAI221_X1 U11138 ( .B1(n9911), .B2(keyinput101), .C1(n7221), .C2(keyinput76), 
        .A(n9910), .ZN(n9922) );
  AOI22_X1 U11139 ( .A1(n9913), .A2(keyinput23), .B1(keyinput44), .B2(n10641), 
        .ZN(n9912) );
  OAI221_X1 U11140 ( .B1(n9913), .B2(keyinput23), .C1(n10641), .C2(keyinput44), 
        .A(n9912), .ZN(n9921) );
  INV_X1 U11141 ( .A(P2_D_REG_22__SCAN_IN), .ZN(n10541) );
  AOI22_X1 U11142 ( .A1(n9915), .A2(keyinput60), .B1(keyinput87), .B2(n10541), 
        .ZN(n9914) );
  OAI221_X1 U11143 ( .B1(n9915), .B2(keyinput60), .C1(n10541), .C2(keyinput87), 
        .A(n9914), .ZN(n9920) );
  AOI22_X1 U11144 ( .A1(n9918), .A2(keyinput57), .B1(keyinput70), .B2(n9917), 
        .ZN(n9916) );
  OAI221_X1 U11145 ( .B1(n9918), .B2(keyinput57), .C1(n9917), .C2(keyinput70), 
        .A(n9916), .ZN(n9919) );
  NOR4_X1 U11146 ( .A1(n9922), .A2(n9921), .A3(n9920), .A4(n9919), .ZN(n10007)
         );
  AOI22_X1 U11147 ( .A1(n9925), .A2(keyinput113), .B1(keyinput104), .B2(n9924), 
        .ZN(n9923) );
  OAI221_X1 U11148 ( .B1(n9925), .B2(keyinput113), .C1(n9924), .C2(keyinput104), .A(n9923), .ZN(n9934) );
  AOI22_X1 U11149 ( .A1(n7050), .A2(keyinput91), .B1(keyinput61), .B2(n9927), 
        .ZN(n9926) );
  OAI221_X1 U11150 ( .B1(n7050), .B2(keyinput91), .C1(n9927), .C2(keyinput61), 
        .A(n9926), .ZN(n9933) );
  AOI22_X1 U11151 ( .A1(n9679), .A2(keyinput33), .B1(n9929), .B2(keyinput71), 
        .ZN(n9928) );
  OAI221_X1 U11152 ( .B1(n9679), .B2(keyinput33), .C1(n9929), .C2(keyinput71), 
        .A(n9928), .ZN(n9932) );
  AOI22_X1 U11153 ( .A1(n6991), .A2(keyinput2), .B1(n5950), .B2(keyinput50), 
        .ZN(n9930) );
  OAI221_X1 U11154 ( .B1(n6991), .B2(keyinput2), .C1(n5950), .C2(keyinput50), 
        .A(n9930), .ZN(n9931) );
  NOR4_X1 U11155 ( .A1(n9934), .A2(n9933), .A3(n9932), .A4(n9931), .ZN(n10006)
         );
  AOI22_X1 U11156 ( .A1(n9937), .A2(keyinput73), .B1(n9936), .B2(keyinput15), 
        .ZN(n9935) );
  OAI221_X1 U11157 ( .B1(n9937), .B2(keyinput73), .C1(n9936), .C2(keyinput15), 
        .A(n9935), .ZN(n9938) );
  INV_X1 U11158 ( .A(n9938), .ZN(n9943) );
  XNOR2_X1 U11159 ( .A(keyinput27), .B(n9939), .ZN(n9941) );
  XNOR2_X1 U11160 ( .A(keyinput72), .B(n7515), .ZN(n9940) );
  NOR2_X1 U11161 ( .A1(n9941), .A2(n9940), .ZN(n9942) );
  NAND2_X1 U11162 ( .A1(n9943), .A2(n9942), .ZN(n9946) );
  AOI22_X1 U11163 ( .A1(n7476), .A2(keyinput75), .B1(n10301), .B2(keyinput6), 
        .ZN(n9944) );
  OAI221_X1 U11164 ( .B1(n7476), .B2(keyinput75), .C1(n10301), .C2(keyinput6), 
        .A(n9944), .ZN(n9945) );
  NOR2_X1 U11165 ( .A1(n9946), .A2(n9945), .ZN(n9962) );
  AOI22_X1 U11166 ( .A1(n9948), .A2(keyinput69), .B1(keyinput8), .B2(n5696), 
        .ZN(n9947) );
  OAI221_X1 U11167 ( .B1(n9948), .B2(keyinput69), .C1(n5696), .C2(keyinput8), 
        .A(n9947), .ZN(n9952) );
  INV_X1 U11168 ( .A(P1_D_REG_7__SCAN_IN), .ZN(n10433) );
  AOI22_X1 U11169 ( .A1(n9950), .A2(keyinput19), .B1(n10433), .B2(keyinput106), 
        .ZN(n9949) );
  OAI221_X1 U11170 ( .B1(n9950), .B2(keyinput19), .C1(n10433), .C2(keyinput106), .A(n9949), .ZN(n9951) );
  NOR2_X1 U11171 ( .A1(n9952), .A2(n9951), .ZN(n9961) );
  INV_X1 U11172 ( .A(P2_WR_REG_SCAN_IN), .ZN(n10305) );
  INV_X1 U11173 ( .A(keyinput110), .ZN(n9953) );
  XNOR2_X1 U11174 ( .A(n10305), .B(n9953), .ZN(n9960) );
  INV_X1 U11175 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n9955) );
  AOI22_X1 U11176 ( .A1(n9955), .A2(keyinput85), .B1(n6381), .B2(keyinput118), 
        .ZN(n9954) );
  OAI221_X1 U11177 ( .B1(n9955), .B2(keyinput85), .C1(n6381), .C2(keyinput118), 
        .A(n9954), .ZN(n9958) );
  AOI22_X1 U11178 ( .A1(n10499), .A2(keyinput49), .B1(n10234), .B2(keyinput55), 
        .ZN(n9956) );
  OAI221_X1 U11179 ( .B1(n10499), .B2(keyinput49), .C1(n10234), .C2(keyinput55), .A(n9956), .ZN(n9957) );
  NOR2_X1 U11180 ( .A1(n9958), .A2(n9957), .ZN(n9959) );
  NAND4_X1 U11181 ( .A1(n9962), .A2(n9961), .A3(n9960), .A4(n9959), .ZN(n10004) );
  AOI22_X1 U11182 ( .A1(n7292), .A2(keyinput13), .B1(n9964), .B2(keyinput62), 
        .ZN(n9963) );
  OAI221_X1 U11183 ( .B1(n7292), .B2(keyinput13), .C1(n9964), .C2(keyinput62), 
        .A(n9963), .ZN(n9968) );
  AOI22_X1 U11184 ( .A1(n7672), .A2(keyinput14), .B1(n9966), .B2(keyinput74), 
        .ZN(n9965) );
  OAI221_X1 U11185 ( .B1(n7672), .B2(keyinput14), .C1(n9966), .C2(keyinput74), 
        .A(n9965), .ZN(n9967) );
  NOR2_X1 U11186 ( .A1(n9968), .A2(n9967), .ZN(n10002) );
  XNOR2_X1 U11187 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(keyinput82), .ZN(n9972)
         );
  XNOR2_X1 U11188 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(keyinput109), .ZN(n9971)
         );
  XNOR2_X1 U11189 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(keyinput83), .ZN(n9970)
         );
  XNOR2_X1 U11190 ( .A(P1_REG3_REG_16__SCAN_IN), .B(keyinput80), .ZN(n9969) );
  NAND4_X1 U11191 ( .A1(n9972), .A2(n9971), .A3(n9970), .A4(n9969), .ZN(n9978)
         );
  XNOR2_X1 U11192 ( .A(P1_REG3_REG_4__SCAN_IN), .B(keyinput63), .ZN(n9976) );
  XNOR2_X1 U11193 ( .A(P1_STATE_REG_SCAN_IN), .B(keyinput98), .ZN(n9975) );
  XNOR2_X1 U11194 ( .A(P1_REG3_REG_14__SCAN_IN), .B(keyinput67), .ZN(n9974) );
  XNOR2_X1 U11195 ( .A(P2_IR_REG_20__SCAN_IN), .B(keyinput58), .ZN(n9973) );
  NAND4_X1 U11196 ( .A1(n9976), .A2(n9975), .A3(n9974), .A4(n9973), .ZN(n9977)
         );
  NOR2_X1 U11197 ( .A1(n9978), .A2(n9977), .ZN(n10001) );
  XNOR2_X1 U11198 ( .A(P2_IR_REG_18__SCAN_IN), .B(keyinput59), .ZN(n9982) );
  XNOR2_X1 U11199 ( .A(P2_IR_REG_27__SCAN_IN), .B(keyinput48), .ZN(n9981) );
  XNOR2_X1 U11200 ( .A(P2_IR_REG_26__SCAN_IN), .B(keyinput22), .ZN(n9980) );
  XNOR2_X1 U11201 ( .A(P2_REG1_REG_10__SCAN_IN), .B(keyinput99), .ZN(n9979) );
  NAND4_X1 U11202 ( .A1(n9982), .A2(n9981), .A3(n9980), .A4(n9979), .ZN(n9988)
         );
  XNOR2_X1 U11203 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(keyinput123), .ZN(n9986)
         );
  XNOR2_X1 U11204 ( .A(P2_REG1_REG_14__SCAN_IN), .B(keyinput7), .ZN(n9985) );
  XNOR2_X1 U11205 ( .A(P2_IR_REG_25__SCAN_IN), .B(keyinput90), .ZN(n9984) );
  XNOR2_X1 U11206 ( .A(P2_IR_REG_4__SCAN_IN), .B(keyinput112), .ZN(n9983) );
  NAND4_X1 U11207 ( .A1(n9986), .A2(n9985), .A3(n9984), .A4(n9983), .ZN(n9987)
         );
  NOR2_X1 U11208 ( .A1(n9988), .A2(n9987), .ZN(n10000) );
  XNOR2_X1 U11209 ( .A(P1_REG2_REG_0__SCAN_IN), .B(keyinput53), .ZN(n9992) );
  XNOR2_X1 U11210 ( .A(P2_REG1_REG_11__SCAN_IN), .B(keyinput89), .ZN(n9991) );
  XNOR2_X1 U11211 ( .A(P1_IR_REG_28__SCAN_IN), .B(keyinput37), .ZN(n9990) );
  XNOR2_X1 U11212 ( .A(P2_REG0_REG_12__SCAN_IN), .B(keyinput45), .ZN(n9989) );
  NAND4_X1 U11213 ( .A1(n9992), .A2(n9991), .A3(n9990), .A4(n9989), .ZN(n9998)
         );
  XNOR2_X1 U11214 ( .A(P1_IR_REG_16__SCAN_IN), .B(keyinput34), .ZN(n9996) );
  XNOR2_X1 U11215 ( .A(P2_IR_REG_29__SCAN_IN), .B(keyinput16), .ZN(n9995) );
  XNOR2_X1 U11216 ( .A(keyinput115), .B(P2_D_REG_10__SCAN_IN), .ZN(n9994) );
  XNOR2_X1 U11217 ( .A(keyinput84), .B(P2_ADDR_REG_3__SCAN_IN), .ZN(n9993) );
  NAND4_X1 U11218 ( .A1(n9996), .A2(n9995), .A3(n9994), .A4(n9993), .ZN(n9997)
         );
  NOR2_X1 U11219 ( .A1(n9998), .A2(n9997), .ZN(n9999) );
  NAND4_X1 U11220 ( .A1(n10002), .A2(n10001), .A3(n10000), .A4(n9999), .ZN(
        n10003) );
  NOR2_X1 U11221 ( .A1(n10004), .A2(n10003), .ZN(n10005) );
  NAND4_X1 U11222 ( .A1(n10008), .A2(n10007), .A3(n10006), .A4(n10005), .ZN(
        n10009) );
  AOI211_X1 U11223 ( .C1(n10011), .C2(keyinput35), .A(n10010), .B(n10009), 
        .ZN(n10029) );
  XOR2_X1 U11224 ( .A(n10012), .B(n10021), .Z(n10203) );
  AOI211_X1 U11225 ( .C1(n10201), .C2(n10014), .A(n6057), .B(n10158), .ZN(
        n10199) );
  INV_X1 U11226 ( .A(n10201), .ZN(n10015) );
  NOR2_X1 U11227 ( .A1(n10015), .A2(n10400), .ZN(n10019) );
  OAI22_X1 U11228 ( .A1(n10017), .A2(n10145), .B1(n10016), .B2(n10148), .ZN(
        n10018) );
  AOI211_X1 U11229 ( .C1(n10199), .C2(n10119), .A(n10019), .B(n10018), .ZN(
        n10027) );
  OAI211_X1 U11230 ( .C1(n10021), .C2(n10020), .A(n9716), .B(n10101), .ZN(
        n10024) );
  NAND2_X1 U11231 ( .A1(n10022), .A2(n10103), .ZN(n10023) );
  OAI211_X1 U11232 ( .C1(n10025), .C2(n10405), .A(n10024), .B(n10023), .ZN(
        n10200) );
  NAND2_X1 U11233 ( .A1(n10200), .A2(n10148), .ZN(n10026) );
  OAI211_X1 U11234 ( .C1(n10203), .C2(n10142), .A(n10027), .B(n10026), .ZN(
        n10028) );
  XOR2_X1 U11235 ( .A(n10029), .B(n10028), .Z(P1_U3268) );
  INV_X1 U11236 ( .A(n10119), .ZN(n10058) );
  OAI22_X1 U11237 ( .A1(n10031), .A2(n10145), .B1(n10030), .B2(n10148), .ZN(
        n10032) );
  AOI21_X1 U11238 ( .B1(n5346), .B2(n10150), .A(n10032), .ZN(n10033) );
  OAI21_X1 U11239 ( .B1(n10034), .B2(n10058), .A(n10033), .ZN(n10037) );
  NOR2_X1 U11240 ( .A1(n10035), .A2(n10142), .ZN(n10036) );
  AOI211_X1 U11241 ( .C1(n10148), .C2(n10038), .A(n10037), .B(n10036), .ZN(
        n10039) );
  INV_X1 U11242 ( .A(n10039), .ZN(P1_U3269) );
  OAI211_X1 U11243 ( .C1(n10041), .C2(n10048), .A(n10040), .B(n10101), .ZN(
        n10045) );
  OAI22_X1 U11244 ( .A1(n10042), .A2(n10405), .B1(n10091), .B2(n10403), .ZN(
        n10043) );
  INV_X1 U11245 ( .A(n10043), .ZN(n10044) );
  INV_X1 U11246 ( .A(n10046), .ZN(n10065) );
  NOR2_X1 U11247 ( .A1(n10065), .A2(n10070), .ZN(n10064) );
  NOR2_X1 U11248 ( .A1(n10064), .A2(n10047), .ZN(n10049) );
  NAND2_X1 U11249 ( .A1(n10049), .A2(n10048), .ZN(n10205) );
  INV_X1 U11250 ( .A(n10049), .ZN(n10051) );
  NAND2_X1 U11251 ( .A1(n10051), .A2(n10050), .ZN(n10204) );
  NAND3_X1 U11252 ( .A1(n10205), .A2(n10424), .A3(n10204), .ZN(n10063) );
  INV_X1 U11253 ( .A(n10052), .ZN(n10054) );
  OAI22_X1 U11254 ( .A1(n10054), .A2(n10145), .B1(n10053), .B2(n10148), .ZN(
        n10060) );
  NAND2_X1 U11255 ( .A1(n10076), .A2(n10061), .ZN(n10055) );
  NAND2_X1 U11256 ( .A1(n10055), .A2(n10418), .ZN(n10056) );
  OR2_X1 U11257 ( .A1(n10057), .A2(n10056), .ZN(n10206) );
  NOR2_X1 U11258 ( .A1(n10206), .A2(n10058), .ZN(n10059) );
  AOI211_X1 U11259 ( .C1(n10150), .C2(n10061), .A(n10060), .B(n10059), .ZN(
        n10062) );
  OAI211_X1 U11260 ( .C1(n10123), .C2(n10208), .A(n10063), .B(n10062), .ZN(
        P1_U3270) );
  AOI21_X1 U11261 ( .B1(n10065), .B2(n10070), .A(n10064), .ZN(n10212) );
  NAND2_X1 U11262 ( .A1(n10212), .A2(n10424), .ZN(n10081) );
  OAI22_X1 U11263 ( .A1(n10148), .A2(n10067), .B1(n10066), .B2(n10145), .ZN(
        n10068) );
  AOI21_X1 U11264 ( .B1(n10075), .B2(n10150), .A(n10068), .ZN(n10080) );
  OAI211_X1 U11265 ( .C1(n5103), .C2(n10070), .A(n10069), .B(n10101), .ZN(
        n10073) );
  NAND2_X1 U11266 ( .A1(n10071), .A2(n10103), .ZN(n10072) );
  OAI211_X1 U11267 ( .C1(n10074), .C2(n10405), .A(n10073), .B(n10072), .ZN(
        n10210) );
  NAND2_X1 U11268 ( .A1(n10210), .A2(n10148), .ZN(n10079) );
  AOI21_X1 U11269 ( .B1(n10092), .B2(n10075), .A(n10158), .ZN(n10077) );
  NAND2_X1 U11270 ( .A1(n10211), .A2(n10119), .ZN(n10078) );
  NAND4_X1 U11271 ( .A1(n10081), .A2(n10080), .A3(n10079), .A4(n10078), .ZN(
        P1_U3271) );
  NAND2_X1 U11272 ( .A1(n10108), .A2(n4604), .ZN(n10109) );
  NAND2_X1 U11273 ( .A1(n10109), .A2(n10082), .ZN(n10083) );
  XOR2_X1 U11274 ( .A(n10086), .B(n10083), .Z(n10219) );
  INV_X1 U11275 ( .A(n10084), .ZN(n10089) );
  AOI21_X1 U11276 ( .B1(n10085), .B2(n10087), .A(n10086), .ZN(n10088) );
  NOR2_X1 U11277 ( .A1(n10089), .A2(n10088), .ZN(n10090) );
  OAI222_X1 U11278 ( .A1(n10405), .A2(n10091), .B1(n10403), .B2(n10133), .C1(
        n10090), .C2(n10406), .ZN(n10215) );
  INV_X1 U11279 ( .A(n10112), .ZN(n10094) );
  INV_X1 U11280 ( .A(n10092), .ZN(n10093) );
  AOI211_X1 U11281 ( .C1(n10217), .C2(n10094), .A(n10158), .B(n10093), .ZN(
        n10216) );
  NAND2_X1 U11282 ( .A1(n10216), .A2(n10422), .ZN(n10097) );
  AOI22_X1 U11283 ( .A1(n10123), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n10095), 
        .B2(n10411), .ZN(n10096) );
  OAI211_X1 U11284 ( .C1(n10098), .C2(n10400), .A(n10097), .B(n10096), .ZN(
        n10099) );
  AOI21_X1 U11285 ( .B1(n10215), .B2(n10148), .A(n10099), .ZN(n10100) );
  OAI21_X1 U11286 ( .B1(n10219), .B2(n10142), .A(n10100), .ZN(P1_U3272) );
  OAI211_X1 U11287 ( .C1(n10111), .C2(n10102), .A(n10085), .B(n10101), .ZN(
        n10106) );
  NAND2_X1 U11288 ( .A1(n10104), .A2(n10103), .ZN(n10105) );
  OAI211_X1 U11289 ( .C1(n10107), .C2(n10405), .A(n10106), .B(n10105), .ZN(
        n10220) );
  INV_X1 U11290 ( .A(n10220), .ZN(n10122) );
  INV_X1 U11291 ( .A(n10109), .ZN(n10110) );
  AOI21_X1 U11292 ( .B1(n5022), .B2(n10111), .A(n10110), .ZN(n10222) );
  NAND2_X1 U11293 ( .A1(n10222), .A2(n10424), .ZN(n10121) );
  INV_X1 U11294 ( .A(n10127), .ZN(n10113) );
  AOI211_X1 U11295 ( .C1(n10114), .C2(n10113), .A(n10158), .B(n10112), .ZN(
        n10221) );
  NOR2_X1 U11296 ( .A1(n10270), .A2(n10400), .ZN(n10118) );
  OAI22_X1 U11297 ( .A1(n10148), .A2(n10116), .B1(n10115), .B2(n10145), .ZN(
        n10117) );
  AOI211_X1 U11298 ( .C1(n10221), .C2(n10119), .A(n10118), .B(n10117), .ZN(
        n10120) );
  OAI211_X1 U11299 ( .C1(n10123), .C2(n10122), .A(n10121), .B(n10120), .ZN(
        P1_U3273) );
  XNOR2_X1 U11300 ( .A(n10124), .B(n10130), .ZN(n10229) );
  NAND2_X1 U11301 ( .A1(n10160), .A2(n10226), .ZN(n10125) );
  NAND2_X1 U11302 ( .A1(n10125), .A2(n10418), .ZN(n10126) );
  NOR2_X1 U11303 ( .A1(n10127), .A2(n10126), .ZN(n10225) );
  INV_X1 U11304 ( .A(n10226), .ZN(n10129) );
  OAI22_X1 U11305 ( .A1(n10129), .A2(n10400), .B1(n10128), .B2(n10148), .ZN(
        n10140) );
  AOI21_X1 U11306 ( .B1(n10131), .B2(n10130), .A(n10406), .ZN(n10136) );
  OAI22_X1 U11307 ( .A1(n10133), .A2(n10405), .B1(n10132), .B2(n10403), .ZN(
        n10134) );
  AOI21_X1 U11308 ( .B1(n10136), .B2(n10135), .A(n10134), .ZN(n10228) );
  NAND2_X1 U11309 ( .A1(n10411), .A2(n10137), .ZN(n10138) );
  AOI21_X1 U11310 ( .B1(n10228), .B2(n10138), .A(n10123), .ZN(n10139) );
  AOI211_X1 U11311 ( .C1(n10225), .C2(n10422), .A(n10140), .B(n10139), .ZN(
        n10141) );
  OAI21_X1 U11312 ( .B1(n10142), .B2(n10229), .A(n10141), .ZN(P1_U3274) );
  XNOR2_X1 U11313 ( .A(n10144), .B(n10143), .ZN(n10233) );
  NAND2_X1 U11314 ( .A1(n10233), .A2(n10424), .ZN(n10165) );
  INV_X1 U11315 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n10147) );
  OAI22_X1 U11316 ( .A1(n10148), .A2(n10147), .B1(n10146), .B2(n10145), .ZN(
        n10149) );
  AOI21_X1 U11317 ( .B1(n10230), .B2(n10150), .A(n10149), .ZN(n10164) );
  NAND2_X1 U11318 ( .A1(n10152), .A2(n10151), .ZN(n10154) );
  XNOR2_X1 U11319 ( .A(n10154), .B(n10153), .ZN(n10157) );
  OAI222_X1 U11320 ( .A1(n10157), .A2(n10406), .B1(n10405), .B2(n10156), .C1(
        n10403), .C2(n10155), .ZN(n10231) );
  NAND2_X1 U11321 ( .A1(n10231), .A2(n10148), .ZN(n10163) );
  AOI21_X1 U11322 ( .B1(n10159), .B2(n10230), .A(n10158), .ZN(n10161) );
  AND2_X1 U11323 ( .A1(n10161), .A2(n10160), .ZN(n10232) );
  NAND2_X1 U11324 ( .A1(n10232), .A2(n10422), .ZN(n10162) );
  NAND4_X1 U11325 ( .A1(n10165), .A2(n10164), .A3(n10163), .A4(n10162), .ZN(
        P1_U3275) );
  NAND2_X1 U11326 ( .A1(n10166), .A2(n10172), .ZN(n10245) );
  OR2_X1 U11327 ( .A1(n10245), .A2(n10168), .ZN(n10170) );
  NAND2_X1 U11328 ( .A1(n10168), .A2(n10167), .ZN(n10169) );
  NAND2_X1 U11329 ( .A1(n10170), .A2(n10169), .ZN(n10171) );
  OAI21_X1 U11330 ( .B1(n10248), .B2(n10236), .A(n10171), .ZN(P1_U3554) );
  INV_X1 U11331 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n10175) );
  INV_X1 U11332 ( .A(n10172), .ZN(n10173) );
  NOR2_X1 U11333 ( .A1(n10174), .A2(n10173), .ZN(n10249) );
  MUX2_X1 U11334 ( .A(n10175), .B(n10249), .S(n10504), .Z(n10176) );
  AOI21_X1 U11335 ( .B1(n10240), .B2(n10178), .A(n10177), .ZN(n10179) );
  OAI211_X1 U11336 ( .C1(n10181), .C2(n10243), .A(n10180), .B(n10179), .ZN(
        n10252) );
  MUX2_X1 U11337 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n10252), .S(n10504), .Z(
        P1_U3550) );
  INV_X1 U11338 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n10187) );
  NAND2_X1 U11339 ( .A1(n10182), .A2(n10489), .ZN(n10186) );
  NOR2_X1 U11340 ( .A1(n10184), .A2(n10183), .ZN(n10185) );
  AND2_X1 U11341 ( .A1(n10186), .A2(n10185), .ZN(n10253) );
  MUX2_X1 U11342 ( .A(n10187), .B(n10253), .S(n10504), .Z(n10188) );
  OAI21_X1 U11343 ( .B1(n10256), .B2(n10236), .A(n10188), .ZN(P1_U3549) );
  AOI21_X1 U11344 ( .B1(n10240), .B2(n10190), .A(n10189), .ZN(n10191) );
  OAI211_X1 U11345 ( .C1(n10193), .C2(n10243), .A(n10192), .B(n10191), .ZN(
        n10257) );
  MUX2_X1 U11346 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n10257), .S(n10504), .Z(
        P1_U3548) );
  INV_X1 U11347 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n10197) );
  AOI211_X1 U11348 ( .C1(n10196), .C2(n10489), .A(n10195), .B(n10194), .ZN(
        n10258) );
  MUX2_X1 U11349 ( .A(n10197), .B(n10258), .S(n10504), .Z(n10198) );
  OAI21_X1 U11350 ( .B1(n4503), .B2(n10236), .A(n10198), .ZN(P1_U3547) );
  AOI211_X1 U11351 ( .C1(n10240), .C2(n10201), .A(n10200), .B(n10199), .ZN(
        n10202) );
  OAI21_X1 U11352 ( .B1(n10243), .B2(n10203), .A(n10202), .ZN(n10261) );
  MUX2_X1 U11353 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n10261), .S(n10504), .Z(
        P1_U3546) );
  NAND3_X1 U11354 ( .A1(n10205), .A2(n10489), .A3(n10204), .ZN(n10209) );
  NAND4_X1 U11355 ( .A1(n10209), .A2(n10208), .A3(n10207), .A4(n10206), .ZN(
        n10262) );
  MUX2_X1 U11356 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n10262), .S(n10504), .Z(
        P1_U3544) );
  INV_X1 U11357 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n10213) );
  AOI211_X1 U11358 ( .C1(n10212), .C2(n10489), .A(n10211), .B(n10210), .ZN(
        n10263) );
  MUX2_X1 U11359 ( .A(n10213), .B(n10263), .S(n10504), .Z(n10214) );
  OAI21_X1 U11360 ( .B1(n4897), .B2(n10236), .A(n10214), .ZN(P1_U3543) );
  AOI211_X1 U11361 ( .C1(n10240), .C2(n10217), .A(n10216), .B(n10215), .ZN(
        n10218) );
  OAI21_X1 U11362 ( .B1(n10243), .B2(n10219), .A(n10218), .ZN(n10266) );
  MUX2_X1 U11363 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n10266), .S(n10504), .Z(
        P1_U3542) );
  INV_X1 U11364 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n10223) );
  AOI211_X1 U11365 ( .C1(n10222), .C2(n10489), .A(n10221), .B(n10220), .ZN(
        n10267) );
  MUX2_X1 U11366 ( .A(n10223), .B(n10267), .S(n10504), .Z(n10224) );
  OAI21_X1 U11367 ( .B1(n10270), .B2(n10236), .A(n10224), .ZN(P1_U3541) );
  AOI21_X1 U11368 ( .B1(n10240), .B2(n10226), .A(n10225), .ZN(n10227) );
  OAI211_X1 U11369 ( .C1(n10229), .C2(n10243), .A(n10228), .B(n10227), .ZN(
        n10271) );
  MUX2_X1 U11370 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n10271), .S(n10504), .Z(
        P1_U3540) );
  INV_X1 U11371 ( .A(n10230), .ZN(n10276) );
  AOI211_X1 U11372 ( .C1(n10233), .C2(n10489), .A(n10232), .B(n10231), .ZN(
        n10272) );
  MUX2_X1 U11373 ( .A(n10234), .B(n10272), .S(n10504), .Z(n10235) );
  OAI21_X1 U11374 ( .B1(n10276), .B2(n10236), .A(n10235), .ZN(P1_U3539) );
  AOI211_X1 U11375 ( .C1(n10240), .C2(n10239), .A(n10238), .B(n10237), .ZN(
        n10241) );
  OAI21_X1 U11376 ( .B1(n10243), .B2(n10242), .A(n10241), .ZN(n10277) );
  MUX2_X1 U11377 ( .A(P1_REG1_REG_11__SCAN_IN), .B(n10277), .S(n10504), .Z(
        P1_U3534) );
  MUX2_X1 U11378 ( .A(P1_REG1_REG_0__SCAN_IN), .B(n10244), .S(n10504), .Z(
        P1_U3523) );
  OR2_X1 U11379 ( .A1(n10245), .A2(n10490), .ZN(n10246) );
  NAND2_X1 U11380 ( .A1(n10246), .A2(n5095), .ZN(n10247) );
  OAI21_X1 U11381 ( .B1(n10248), .B2(n10275), .A(n10247), .ZN(P1_U3522) );
  INV_X1 U11382 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n10250) );
  MUX2_X1 U11383 ( .A(n10250), .B(n10249), .S(n10492), .Z(n10251) );
  OAI21_X1 U11384 ( .B1(n9636), .B2(n10275), .A(n10251), .ZN(P1_U3521) );
  MUX2_X1 U11385 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n10252), .S(n10492), .Z(
        P1_U3518) );
  INV_X1 U11386 ( .A(P1_REG0_REG_26__SCAN_IN), .ZN(n10254) );
  MUX2_X1 U11387 ( .A(n10254), .B(n10253), .S(n10492), .Z(n10255) );
  OAI21_X1 U11388 ( .B1(n10256), .B2(n10275), .A(n10255), .ZN(P1_U3517) );
  MUX2_X1 U11389 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n10257), .S(n10492), .Z(
        P1_U3516) );
  INV_X1 U11390 ( .A(P1_REG0_REG_24__SCAN_IN), .ZN(n10259) );
  MUX2_X1 U11391 ( .A(n10259), .B(n10258), .S(n10492), .Z(n10260) );
  OAI21_X1 U11392 ( .B1(n4503), .B2(n10275), .A(n10260), .ZN(P1_U3515) );
  MUX2_X1 U11393 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n10261), .S(n10492), .Z(
        P1_U3514) );
  MUX2_X1 U11394 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n10262), .S(n10492), .Z(
        P1_U3512) );
  INV_X1 U11395 ( .A(P1_REG0_REG_20__SCAN_IN), .ZN(n10264) );
  MUX2_X1 U11396 ( .A(n10264), .B(n10263), .S(n10492), .Z(n10265) );
  OAI21_X1 U11397 ( .B1(n4897), .B2(n10275), .A(n10265), .ZN(P1_U3511) );
  MUX2_X1 U11398 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n10266), .S(n10492), .Z(
        P1_U3510) );
  INV_X1 U11399 ( .A(P1_REG0_REG_18__SCAN_IN), .ZN(n10268) );
  MUX2_X1 U11400 ( .A(n10268), .B(n10267), .S(n10492), .Z(n10269) );
  OAI21_X1 U11401 ( .B1(n10270), .B2(n10275), .A(n10269), .ZN(P1_U3508) );
  MUX2_X1 U11402 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n10271), .S(n10492), .Z(
        P1_U3505) );
  INV_X1 U11403 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n10273) );
  MUX2_X1 U11404 ( .A(n10273), .B(n10272), .S(n10492), .Z(n10274) );
  OAI21_X1 U11405 ( .B1(n10276), .B2(n10275), .A(n10274), .ZN(P1_U3502) );
  MUX2_X1 U11406 ( .A(P1_REG0_REG_11__SCAN_IN), .B(n10277), .S(n10492), .Z(
        P1_U3487) );
  MUX2_X1 U11407 ( .A(P1_D_REG_0__SCAN_IN), .B(n10278), .S(n10428), .Z(
        P1_U3440) );
  NOR4_X1 U11408 ( .A1(n10279), .A2(P1_IR_REG_30__SCAN_IN), .A3(n4918), .A4(
        P1_U3084), .ZN(n10280) );
  AOI21_X1 U11409 ( .B1(n10281), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n10280), 
        .ZN(n10282) );
  OAI21_X1 U11410 ( .B1(n10284), .B2(n10283), .A(n10282), .ZN(P1_U3322) );
  INV_X1 U11411 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n10287) );
  OAI222_X1 U11412 ( .A1(n10294), .A2(n10287), .B1(n10292), .B2(n10286), .C1(
        n10285), .C2(P1_U3084), .ZN(P1_U3324) );
  INV_X1 U11413 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n10293) );
  INV_X1 U11414 ( .A(n10288), .ZN(n10291) );
  OAI222_X1 U11415 ( .A1(n10294), .A2(n10293), .B1(n10292), .B2(n10291), .C1(
        n10290), .C2(P1_U3084), .ZN(P1_U3325) );
  INV_X1 U11416 ( .A(n10295), .ZN(n10296) );
  MUX2_X1 U11417 ( .A(n10296), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3353) );
  OAI211_X1 U11418 ( .C1(n4900), .C2(n10485), .A(n10298), .B(n10297), .ZN(
        n10299) );
  AOI21_X1 U11419 ( .B1(n10489), .B2(n10300), .A(n10299), .ZN(n10303) );
  AOI22_X1 U11420 ( .A1(n10492), .A2(n10303), .B1(n10301), .B2(n10490), .ZN(
        P1_U3484) );
  INV_X1 U11421 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n10302) );
  AOI22_X1 U11422 ( .A1(n10504), .A2(n10303), .B1(n10302), .B2(n10168), .ZN(
        P1_U3533) );
  AOI22_X1 U11423 ( .A1(P1_WR_REG_SCAN_IN), .A2(n10305), .B1(P2_WR_REG_SCAN_IN), .B2(n10304), .ZN(U123) );
  XNOR2_X1 U11424 ( .A(P2_RD_REG_SCAN_IN), .B(P1_RD_REG_SCAN_IN), .ZN(U126) );
  NAND2_X1 U11425 ( .A1(n10306), .A2(P1_IR_REG_0__SCAN_IN), .ZN(n10310) );
  NAND2_X1 U11426 ( .A1(n10308), .A2(n10307), .ZN(n10309) );
  MUX2_X1 U11427 ( .A(n10310), .B(n10309), .S(P1_REG1_REG_0__SCAN_IN), .Z(
        n10311) );
  NAND2_X1 U11428 ( .A1(n10312), .A2(n10311), .ZN(n10313) );
  AOI22_X1 U11429 ( .A1(n10319), .A2(P1_ADDR_REG_0__SCAN_IN), .B1(n10314), 
        .B2(n10313), .ZN(n10315) );
  OAI21_X1 U11430 ( .B1(P1_STATE_REG_SCAN_IN), .B2(n7515), .A(n10315), .ZN(
        P1_U3241) );
  INV_X1 U11431 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n10316) );
  OAI22_X1 U11432 ( .A1(n10390), .A2(n10317), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n10316), .ZN(n10318) );
  AOI21_X1 U11433 ( .B1(n10319), .B2(P1_ADDR_REG_1__SCAN_IN), .A(n10318), .ZN(
        n10328) );
  OAI211_X1 U11434 ( .C1(n10322), .C2(n10321), .A(n10395), .B(n10320), .ZN(
        n10327) );
  OAI211_X1 U11435 ( .C1(n10325), .C2(n10324), .A(n10383), .B(n10323), .ZN(
        n10326) );
  NAND3_X1 U11436 ( .A1(n10328), .A2(n10327), .A3(n10326), .ZN(P1_U3242) );
  INV_X1 U11437 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n10341) );
  AOI211_X1 U11438 ( .C1(n10331), .C2(n10330), .A(n10357), .B(n10329), .ZN(
        n10332) );
  AOI211_X1 U11439 ( .C1(n10363), .C2(n10334), .A(n10333), .B(n10332), .ZN(
        n10340) );
  AND2_X1 U11440 ( .A1(n10336), .A2(n10335), .ZN(n10337) );
  OAI21_X1 U11441 ( .B1(n10338), .B2(n10337), .A(n10395), .ZN(n10339) );
  OAI211_X1 U11442 ( .C1(n10341), .C2(n10399), .A(n10340), .B(n10339), .ZN(
        P1_U3255) );
  INV_X1 U11443 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n10354) );
  AOI21_X1 U11444 ( .B1(n10344), .B2(n10343), .A(n10342), .ZN(n10345) );
  NAND2_X1 U11445 ( .A1(n10383), .A2(n10345), .ZN(n10349) );
  NAND2_X1 U11446 ( .A1(n10363), .A2(n10346), .ZN(n10348) );
  AND3_X1 U11447 ( .A1(n10349), .A2(n10348), .A3(n10347), .ZN(n10353) );
  OAI211_X1 U11448 ( .C1(P1_REG1_REG_15__SCAN_IN), .C2(n10351), .A(n10395), 
        .B(n10350), .ZN(n10352) );
  OAI211_X1 U11449 ( .C1(n10354), .C2(n10399), .A(n10353), .B(n10352), .ZN(
        P1_U3256) );
  INV_X1 U11450 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n10369) );
  INV_X1 U11451 ( .A(n10355), .ZN(n10356) );
  AOI211_X1 U11452 ( .C1(n10359), .C2(n10358), .A(n10357), .B(n10356), .ZN(
        n10360) );
  AOI211_X1 U11453 ( .C1(n10363), .C2(n10362), .A(n10361), .B(n10360), .ZN(
        n10368) );
  XNOR2_X1 U11454 ( .A(n10365), .B(n10364), .ZN(n10366) );
  NAND2_X1 U11455 ( .A1(n10366), .A2(n10395), .ZN(n10367) );
  OAI211_X1 U11456 ( .C1(n10369), .C2(n10399), .A(n10368), .B(n10367), .ZN(
        P1_U3257) );
  INV_X1 U11457 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n10382) );
  OAI211_X1 U11458 ( .C1(n10372), .C2(n10371), .A(n10370), .B(n10383), .ZN(
        n10374) );
  OAI211_X1 U11459 ( .C1(n10390), .C2(n10375), .A(n10374), .B(n10373), .ZN(
        n10376) );
  INV_X1 U11460 ( .A(n10376), .ZN(n10381) );
  XOR2_X1 U11461 ( .A(n10378), .B(n10377), .Z(n10379) );
  NAND2_X1 U11462 ( .A1(n10379), .A2(n10395), .ZN(n10380) );
  OAI211_X1 U11463 ( .C1(n10382), .C2(n10399), .A(n10381), .B(n10380), .ZN(
        P1_U3258) );
  INV_X1 U11464 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n10642) );
  OAI211_X1 U11465 ( .C1(n10386), .C2(n10385), .A(n10384), .B(n10383), .ZN(
        n10388) );
  OAI211_X1 U11466 ( .C1(n10390), .C2(n10389), .A(n10388), .B(n10387), .ZN(
        n10391) );
  INV_X1 U11467 ( .A(n10391), .ZN(n10398) );
  OAI21_X1 U11468 ( .B1(n10394), .B2(n10393), .A(n10392), .ZN(n10396) );
  NAND2_X1 U11469 ( .A1(n10396), .A2(n10395), .ZN(n10397) );
  OAI211_X1 U11470 ( .C1(n10642), .C2(n10399), .A(n10398), .B(n10397), .ZN(
        P1_U3259) );
  NOR2_X1 U11471 ( .A1(n10400), .A2(n10421), .ZN(n10409) );
  XNOR2_X1 U11472 ( .A(n10401), .B(n10415), .ZN(n10407) );
  OAI222_X1 U11473 ( .A1(n10407), .A2(n10406), .B1(n10405), .B2(n10404), .C1(
        n10403), .C2(n10402), .ZN(n10455) );
  MUX2_X1 U11474 ( .A(n10455), .B(P1_REG2_REG_5__SCAN_IN), .S(n10123), .Z(
        n10408) );
  AOI211_X1 U11475 ( .C1(n10411), .C2(n10410), .A(n10409), .B(n10408), .ZN(
        n10426) );
  INV_X1 U11476 ( .A(n10412), .ZN(n10413) );
  AOI21_X1 U11477 ( .B1(n10415), .B2(n10414), .A(n10413), .ZN(n10457) );
  INV_X1 U11478 ( .A(n10416), .ZN(n10420) );
  INV_X1 U11479 ( .A(n10417), .ZN(n10419) );
  OAI211_X1 U11480 ( .C1(n10421), .C2(n10420), .A(n10419), .B(n10418), .ZN(
        n10454) );
  INV_X1 U11481 ( .A(n10454), .ZN(n10423) );
  AOI22_X1 U11482 ( .A1(n10457), .A2(n10424), .B1(n10423), .B2(n10422), .ZN(
        n10425) );
  NAND2_X1 U11483 ( .A1(n10426), .A2(n10425), .ZN(P1_U3286) );
  INV_X1 U11484 ( .A(n10427), .ZN(n10429) );
  AND2_X1 U11485 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n10435), .ZN(P1_U3292) );
  AND2_X1 U11486 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n10435), .ZN(P1_U3293) );
  AND2_X1 U11487 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n10435), .ZN(P1_U3294) );
  AND2_X1 U11488 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n10435), .ZN(P1_U3295) );
  AND2_X1 U11489 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n10435), .ZN(P1_U3296) );
  NOR2_X1 U11490 ( .A1(n10434), .A2(n9777), .ZN(P1_U3297) );
  AND2_X1 U11491 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n10435), .ZN(P1_U3298) );
  AND2_X1 U11492 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n10435), .ZN(P1_U3299) );
  AND2_X1 U11493 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n10435), .ZN(P1_U3300) );
  AND2_X1 U11494 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n10435), .ZN(P1_U3301) );
  NOR2_X1 U11495 ( .A1(n10434), .A2(n10430), .ZN(P1_U3302) );
  AND2_X1 U11496 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n10435), .ZN(P1_U3303) );
  AND2_X1 U11497 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n10435), .ZN(P1_U3304) );
  AND2_X1 U11498 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n10435), .ZN(P1_U3305) );
  AND2_X1 U11499 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n10435), .ZN(P1_U3306) );
  AND2_X1 U11500 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n10435), .ZN(P1_U3307) );
  AND2_X1 U11501 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n10435), .ZN(P1_U3308) );
  AND2_X1 U11502 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n10435), .ZN(P1_U3309) );
  NOR2_X1 U11503 ( .A1(n10434), .A2(n10431), .ZN(P1_U3310) );
  AND2_X1 U11504 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n10435), .ZN(P1_U3311) );
  NOR2_X1 U11505 ( .A1(n10434), .A2(n10432), .ZN(P1_U3312) );
  AND2_X1 U11506 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n10435), .ZN(P1_U3313) );
  AND2_X1 U11507 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n10435), .ZN(P1_U3314) );
  AND2_X1 U11508 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n10435), .ZN(P1_U3315) );
  NOR2_X1 U11509 ( .A1(n10434), .A2(n10433), .ZN(P1_U3316) );
  AND2_X1 U11510 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n10435), .ZN(P1_U3317) );
  AND2_X1 U11511 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n10435), .ZN(P1_U3318) );
  AND2_X1 U11512 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n10435), .ZN(P1_U3319) );
  AND2_X1 U11513 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n10435), .ZN(P1_U3320) );
  AND2_X1 U11514 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n10435), .ZN(P1_U3321) );
  INV_X1 U11515 ( .A(n10436), .ZN(n10438) );
  OAI211_X1 U11516 ( .C1(n6054), .C2(n10485), .A(n10438), .B(n10437), .ZN(
        n10441) );
  INV_X1 U11517 ( .A(n10439), .ZN(n10440) );
  AOI211_X1 U11518 ( .C1(n10465), .C2(n10442), .A(n10441), .B(n10440), .ZN(
        n10494) );
  INV_X1 U11519 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n10443) );
  AOI22_X1 U11520 ( .A1(n10492), .A2(n10494), .B1(n10443), .B2(n10490), .ZN(
        P1_U3457) );
  INV_X1 U11521 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n10444) );
  AOI22_X1 U11522 ( .A1(n10492), .A2(n10445), .B1(n10444), .B2(n10490), .ZN(
        P1_U3460) );
  NAND2_X1 U11523 ( .A1(n10447), .A2(n10446), .ZN(n10448) );
  AOI21_X1 U11524 ( .B1(n10449), .B2(n10489), .A(n10448), .ZN(n10450) );
  AND2_X1 U11525 ( .A1(n10451), .A2(n10450), .ZN(n10495) );
  INV_X1 U11526 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n10452) );
  AOI22_X1 U11527 ( .A1(n10492), .A2(n10495), .B1(n10452), .B2(n10490), .ZN(
        P1_U3466) );
  NAND2_X1 U11528 ( .A1(n10454), .A2(n10453), .ZN(n10456) );
  AOI211_X1 U11529 ( .C1(n10457), .C2(n10489), .A(n10456), .B(n10455), .ZN(
        n10496) );
  INV_X1 U11530 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n10458) );
  AOI22_X1 U11531 ( .A1(n10492), .A2(n10496), .B1(n10458), .B2(n10490), .ZN(
        P1_U3469) );
  INV_X1 U11532 ( .A(n10459), .ZN(n10460) );
  NAND2_X1 U11533 ( .A1(n10461), .A2(n10460), .ZN(n10463) );
  AOI211_X1 U11534 ( .C1(n10465), .C2(n10464), .A(n10463), .B(n10462), .ZN(
        n10498) );
  INV_X1 U11535 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n10466) );
  AOI22_X1 U11536 ( .A1(n10492), .A2(n10498), .B1(n10466), .B2(n10490), .ZN(
        P1_U3472) );
  NAND3_X1 U11537 ( .A1(n10469), .A2(n10468), .A3(n10467), .ZN(n10470) );
  AOI21_X1 U11538 ( .B1(n10489), .B2(n10471), .A(n10470), .ZN(n10500) );
  INV_X1 U11539 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n10472) );
  AOI22_X1 U11540 ( .A1(n10492), .A2(n10500), .B1(n10472), .B2(n10490), .ZN(
        P1_U3475) );
  NOR2_X1 U11541 ( .A1(n10474), .A2(n10473), .ZN(n10480) );
  INV_X1 U11542 ( .A(n10475), .ZN(n10478) );
  OAI211_X1 U11543 ( .C1(n10478), .C2(n10485), .A(n10477), .B(n10476), .ZN(
        n10479) );
  AOI211_X1 U11544 ( .C1(n10482), .C2(n10481), .A(n10480), .B(n10479), .ZN(
        n10501) );
  INV_X1 U11545 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n10483) );
  AOI22_X1 U11546 ( .A1(n10492), .A2(n10501), .B1(n10483), .B2(n10490), .ZN(
        P1_U3478) );
  OAI21_X1 U11547 ( .B1(n6056), .B2(n10485), .A(n10484), .ZN(n10487) );
  AOI211_X1 U11548 ( .C1(n10489), .C2(n10488), .A(n10487), .B(n10486), .ZN(
        n10503) );
  INV_X1 U11549 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n10491) );
  AOI22_X1 U11550 ( .A1(n10492), .A2(n10503), .B1(n10491), .B2(n10490), .ZN(
        P1_U3481) );
  AOI22_X1 U11551 ( .A1(n10504), .A2(n10494), .B1(n10493), .B2(n10168), .ZN(
        P1_U3524) );
  AOI22_X1 U11552 ( .A1(n10504), .A2(n10495), .B1(n7404), .B2(n10168), .ZN(
        P1_U3527) );
  AOI22_X1 U11553 ( .A1(n10504), .A2(n10496), .B1(n7050), .B2(n10168), .ZN(
        P1_U3528) );
  AOI22_X1 U11554 ( .A1(n10504), .A2(n10498), .B1(n10497), .B2(n10168), .ZN(
        P1_U3529) );
  AOI22_X1 U11555 ( .A1(n10504), .A2(n10500), .B1(n10499), .B2(n10168), .ZN(
        P1_U3530) );
  AOI22_X1 U11556 ( .A1(n10504), .A2(n10501), .B1(n7214), .B2(n10168), .ZN(
        P1_U3531) );
  AOI22_X1 U11557 ( .A1(n10504), .A2(n10503), .B1(n10502), .B2(n10168), .ZN(
        P1_U3532) );
  AOI22_X1 U11558 ( .A1(n10506), .A2(P2_REG2_REG_0__SCAN_IN), .B1(
        P2_REG1_REG_0__SCAN_IN), .B2(n10505), .ZN(n10516) );
  AOI21_X1 U11559 ( .B1(n10508), .B2(P2_ADDR_REG_0__SCAN_IN), .A(n10507), .ZN(
        n10515) );
  OAI21_X1 U11560 ( .B1(P2_REG1_REG_0__SCAN_IN), .B2(n10510), .A(n10509), .ZN(
        n10513) );
  NOR2_X1 U11561 ( .A1(n10511), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n10512) );
  OAI21_X1 U11562 ( .B1(n10513), .B2(n10512), .A(P2_IR_REG_0__SCAN_IN), .ZN(
        n10514) );
  OAI211_X1 U11563 ( .C1(P2_IR_REG_0__SCAN_IN), .C2(n10516), .A(n10515), .B(
        n10514), .ZN(P2_U3245) );
  AOI22_X1 U11564 ( .A1(n10517), .A2(n6991), .B1(P2_REG2_REG_3__SCAN_IN), .B2(
        n10529), .ZN(n10527) );
  NAND2_X1 U11565 ( .A1(n10519), .A2(n10518), .ZN(n10522) );
  NAND2_X1 U11566 ( .A1(n9158), .A2(n10520), .ZN(n10521) );
  OAI211_X1 U11567 ( .C1(n10524), .C2(n10523), .A(n10522), .B(n10521), .ZN(
        n10525) );
  INV_X1 U11568 ( .A(n10525), .ZN(n10526) );
  OAI211_X1 U11569 ( .C1(n10529), .C2(n10528), .A(n10527), .B(n10526), .ZN(
        P2_U3293) );
  INV_X1 U11570 ( .A(P2_D_REG_31__SCAN_IN), .ZN(n10532) );
  NOR2_X1 U11571 ( .A1(n10567), .A2(n10532), .ZN(P2_U3297) );
  INV_X1 U11572 ( .A(P2_D_REG_30__SCAN_IN), .ZN(n10533) );
  NOR2_X1 U11573 ( .A1(n10567), .A2(n10533), .ZN(P2_U3298) );
  INV_X1 U11574 ( .A(P2_D_REG_29__SCAN_IN), .ZN(n10534) );
  NOR2_X1 U11575 ( .A1(n10567), .A2(n10534), .ZN(P2_U3299) );
  INV_X1 U11576 ( .A(P2_D_REG_28__SCAN_IN), .ZN(n10535) );
  NOR2_X1 U11577 ( .A1(n10567), .A2(n10535), .ZN(P2_U3300) );
  INV_X1 U11578 ( .A(P2_D_REG_27__SCAN_IN), .ZN(n10536) );
  NOR2_X1 U11579 ( .A1(n10546), .A2(n10536), .ZN(P2_U3301) );
  INV_X1 U11580 ( .A(P2_D_REG_26__SCAN_IN), .ZN(n10537) );
  NOR2_X1 U11581 ( .A1(n10546), .A2(n10537), .ZN(P2_U3302) );
  INV_X1 U11582 ( .A(P2_D_REG_25__SCAN_IN), .ZN(n10538) );
  NOR2_X1 U11583 ( .A1(n10546), .A2(n10538), .ZN(P2_U3303) );
  INV_X1 U11584 ( .A(P2_D_REG_24__SCAN_IN), .ZN(n10539) );
  NOR2_X1 U11585 ( .A1(n10546), .A2(n10539), .ZN(P2_U3304) );
  INV_X1 U11586 ( .A(P2_D_REG_23__SCAN_IN), .ZN(n10540) );
  NOR2_X1 U11587 ( .A1(n10546), .A2(n10540), .ZN(P2_U3305) );
  NOR2_X1 U11588 ( .A1(n10546), .A2(n10541), .ZN(P2_U3306) );
  INV_X1 U11589 ( .A(P2_D_REG_21__SCAN_IN), .ZN(n10542) );
  NOR2_X1 U11590 ( .A1(n10546), .A2(n10542), .ZN(P2_U3307) );
  INV_X1 U11591 ( .A(P2_D_REG_20__SCAN_IN), .ZN(n10543) );
  NOR2_X1 U11592 ( .A1(n10546), .A2(n10543), .ZN(P2_U3308) );
  INV_X1 U11593 ( .A(P2_D_REG_19__SCAN_IN), .ZN(n10544) );
  NOR2_X1 U11594 ( .A1(n10546), .A2(n10544), .ZN(P2_U3309) );
  INV_X1 U11595 ( .A(P2_D_REG_18__SCAN_IN), .ZN(n10545) );
  NOR2_X1 U11596 ( .A1(n10546), .A2(n10545), .ZN(P2_U3310) );
  INV_X1 U11597 ( .A(P2_D_REG_17__SCAN_IN), .ZN(n10547) );
  NOR2_X1 U11598 ( .A1(n10567), .A2(n10547), .ZN(P2_U3311) );
  INV_X1 U11599 ( .A(P2_D_REG_16__SCAN_IN), .ZN(n10548) );
  NOR2_X1 U11600 ( .A1(n10567), .A2(n10548), .ZN(P2_U3312) );
  INV_X1 U11601 ( .A(P2_D_REG_15__SCAN_IN), .ZN(n10549) );
  NOR2_X1 U11602 ( .A1(n10567), .A2(n10549), .ZN(P2_U3313) );
  NOR2_X1 U11603 ( .A1(n10567), .A2(n10550), .ZN(P2_U3314) );
  INV_X1 U11604 ( .A(P2_D_REG_13__SCAN_IN), .ZN(n10551) );
  NOR2_X1 U11605 ( .A1(n10567), .A2(n10551), .ZN(P2_U3315) );
  INV_X1 U11606 ( .A(P2_D_REG_12__SCAN_IN), .ZN(n10552) );
  NOR2_X1 U11607 ( .A1(n10567), .A2(n10552), .ZN(P2_U3316) );
  NOR2_X1 U11608 ( .A1(n10567), .A2(n10553), .ZN(P2_U3317) );
  NOR2_X1 U11609 ( .A1(n10567), .A2(n10554), .ZN(P2_U3318) );
  INV_X1 U11610 ( .A(P2_D_REG_9__SCAN_IN), .ZN(n10555) );
  NOR2_X1 U11611 ( .A1(n10567), .A2(n10555), .ZN(P2_U3319) );
  INV_X1 U11612 ( .A(P2_D_REG_8__SCAN_IN), .ZN(n10556) );
  NOR2_X1 U11613 ( .A1(n10567), .A2(n10556), .ZN(P2_U3320) );
  NOR2_X1 U11614 ( .A1(n10567), .A2(n10557), .ZN(P2_U3321) );
  INV_X1 U11615 ( .A(P2_D_REG_6__SCAN_IN), .ZN(n10558) );
  NOR2_X1 U11616 ( .A1(n10567), .A2(n10558), .ZN(P2_U3322) );
  INV_X1 U11617 ( .A(P2_D_REG_5__SCAN_IN), .ZN(n10559) );
  NOR2_X1 U11618 ( .A1(n10567), .A2(n10559), .ZN(P2_U3323) );
  NOR2_X1 U11619 ( .A1(n10567), .A2(n10560), .ZN(P2_U3324) );
  NOR2_X1 U11620 ( .A1(n10567), .A2(n10561), .ZN(P2_U3325) );
  INV_X1 U11621 ( .A(P2_D_REG_2__SCAN_IN), .ZN(n10562) );
  NOR2_X1 U11622 ( .A1(n10567), .A2(n10562), .ZN(P2_U3326) );
  OAI22_X1 U11623 ( .A1(P2_D_REG_0__SCAN_IN), .A2(n10567), .B1(n10563), .B2(
        n10565), .ZN(n10564) );
  INV_X1 U11624 ( .A(n10564), .ZN(P2_U3437) );
  OAI22_X1 U11625 ( .A1(P2_D_REG_1__SCAN_IN), .A2(n10567), .B1(n10566), .B2(
        n10565), .ZN(n10568) );
  INV_X1 U11626 ( .A(n10568), .ZN(P2_U3438) );
  AOI22_X1 U11627 ( .A1(n10570), .A2(n10583), .B1(n10569), .B2(n6657), .ZN(
        n10572) );
  AND2_X1 U11628 ( .A1(n10572), .A2(n10571), .ZN(n10599) );
  AOI22_X1 U11629 ( .A1(n10598), .A2(n10599), .B1(n6121), .B2(n10596), .ZN(
        P2_U3451) );
  OAI211_X1 U11630 ( .C1(n10575), .C2(n10588), .A(n10574), .B(n10573), .ZN(
        n10576) );
  AOI21_X1 U11631 ( .B1(n10583), .B2(n10577), .A(n10576), .ZN(n10601) );
  INV_X1 U11632 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n10578) );
  AOI22_X1 U11633 ( .A1(n10598), .A2(n10601), .B1(n10578), .B2(n10596), .ZN(
        P2_U3466) );
  OAI22_X1 U11634 ( .A1(n10580), .A2(n10590), .B1(n10579), .B2(n10588), .ZN(
        n10582) );
  AOI211_X1 U11635 ( .C1(n10584), .C2(n10583), .A(n10582), .B(n10581), .ZN(
        n10602) );
  INV_X1 U11636 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n10585) );
  AOI22_X1 U11637 ( .A1(n10598), .A2(n10602), .B1(n10585), .B2(n10596), .ZN(
        P2_U3469) );
  INV_X1 U11638 ( .A(n10586), .ZN(n10595) );
  INV_X1 U11639 ( .A(n10587), .ZN(n10594) );
  OAI22_X1 U11640 ( .A1(n10591), .A2(n10590), .B1(n10589), .B2(n10588), .ZN(
        n10593) );
  AOI211_X1 U11641 ( .C1(n10595), .C2(n10594), .A(n10593), .B(n10592), .ZN(
        n10604) );
  INV_X1 U11642 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n10597) );
  AOI22_X1 U11643 ( .A1(n10598), .A2(n10604), .B1(n10597), .B2(n10596), .ZN(
        P2_U3475) );
  AOI22_X1 U11644 ( .A1(n10605), .A2(n10599), .B1(n7109), .B2(n10603), .ZN(
        P2_U3520) );
  AOI22_X1 U11645 ( .A1(n10605), .A2(n10601), .B1(n10600), .B2(n10603), .ZN(
        P2_U3525) );
  AOI22_X1 U11646 ( .A1(n10605), .A2(n10602), .B1(n7154), .B2(n10603), .ZN(
        P2_U3526) );
  AOI22_X1 U11647 ( .A1(n10605), .A2(n10604), .B1(n7198), .B2(n10603), .ZN(
        P2_U3528) );
  INV_X1 U11648 ( .A(n10606), .ZN(n10607) );
  NAND2_X1 U11649 ( .A1(n10608), .A2(n10607), .ZN(n10609) );
  XOR2_X1 U11650 ( .A(n10610), .B(n10609), .Z(ADD_1071_U5) );
  XOR2_X1 U11651 ( .A(P1_ADDR_REG_0__SCAN_IN), .B(P2_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1071_U46) );
  OAI21_X1 U11652 ( .B1(n10613), .B2(n10612), .A(n10611), .ZN(ADD_1071_U56) );
  OAI21_X1 U11653 ( .B1(n10616), .B2(n10615), .A(n10614), .ZN(ADD_1071_U57) );
  OAI21_X1 U11654 ( .B1(n10619), .B2(n10618), .A(n10617), .ZN(ADD_1071_U58) );
  OAI21_X1 U11655 ( .B1(n10622), .B2(n10621), .A(n10620), .ZN(ADD_1071_U59) );
  OAI21_X1 U11656 ( .B1(n10625), .B2(n10624), .A(n10623), .ZN(ADD_1071_U60) );
  OAI21_X1 U11657 ( .B1(n10628), .B2(n10627), .A(n10626), .ZN(ADD_1071_U61) );
  AOI21_X1 U11658 ( .B1(n10631), .B2(n10630), .A(n10629), .ZN(ADD_1071_U62) );
  AOI21_X1 U11659 ( .B1(n10634), .B2(n10633), .A(n10632), .ZN(ADD_1071_U63) );
  XOR2_X1 U11660 ( .A(n10635), .B(P2_ADDR_REG_6__SCAN_IN), .Z(ADD_1071_U50) );
  NOR2_X1 U11661 ( .A1(n10637), .A2(n10636), .ZN(n10638) );
  XOR2_X1 U11662 ( .A(P1_ADDR_REG_5__SCAN_IN), .B(n10638), .Z(ADD_1071_U51) );
  OAI21_X1 U11663 ( .B1(n10641), .B2(n10640), .A(n10639), .ZN(n10643) );
  XOR2_X1 U11664 ( .A(n10643), .B(n10642), .Z(ADD_1071_U55) );
  INV_X1 U11665 ( .A(n10646), .ZN(n10645) );
  OAI222_X1 U11666 ( .A1(n10648), .A2(n10647), .B1(n10648), .B2(n10646), .C1(
        n10645), .C2(n10644), .ZN(ADD_1071_U47) );
  OAI21_X1 U11667 ( .B1(n10650), .B2(n7221), .A(n10649), .ZN(n10652) );
  XNOR2_X1 U11668 ( .A(n10652), .B(n10651), .ZN(ADD_1071_U48) );
  XOR2_X1 U11669 ( .A(P2_ADDR_REG_7__SCAN_IN), .B(n10653), .Z(ADD_1071_U49) );
  XOR2_X1 U11670 ( .A(n10655), .B(n10654), .Z(ADD_1071_U54) );
  XOR2_X1 U11671 ( .A(n10657), .B(n10656), .Z(ADD_1071_U53) );
  XNOR2_X1 U11672 ( .A(n10659), .B(n10658), .ZN(ADD_1071_U52) );
  AND2_X1 U4917 ( .A1(n5568), .A2(n5249), .ZN(n5570) );
  CLKBUF_X1 U5374 ( .A(n6161), .Z(n6455) );
  CLKBUF_X1 U5835 ( .A(n9149), .Z(n4547) );
  CLKBUF_X1 U6368 ( .A(n6956), .Z(n4535) );
  INV_X1 U6421 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n5944) );
  CLKBUF_X1 U6924 ( .A(n7002), .Z(n4545) );
  XNOR2_X1 U7084 ( .A(n5404), .B(n5722), .ZN(n9733) );
endmodule

