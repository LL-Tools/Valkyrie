

module b20_C_gen_AntiSAT_k_256_6 ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, 
        P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, 
        P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, 
        P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, 
        P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, 
        P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, 
        P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, 
        P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, 
        P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, 
        P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, 
        P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, 
        P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, 
        P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, 
        P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, 
        P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, 
        P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, 
        P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, 
        P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, 
        P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, 
        P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, 
        P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, 
        P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, 
        P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, 
        P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, 
        P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, 
        P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN, 
        P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN, 
        P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN, 
        P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN, 
        P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN, 
        P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN, 
        P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN, 
        P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN, 
        P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN, 
        P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN, 
        P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN, 
        P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN, 
        P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN, 
        P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN, 
        P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN, 
        P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN, 
        P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN, 
        P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN, 
        P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN, 
        P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN, 
        P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN, 
        P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN, 
        P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN, 
        P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN, 
        P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN, 
        P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN, 
        P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, 
        P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, 
        P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, 
        P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN, 
        P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN, 
        P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN, 
        P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN, 
        P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN, 
        P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN, 
        P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN, 
        P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN, 
        P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN, 
        P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN, 
        P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN, 
        P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN, 
        P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN, 
        P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN, 
        P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN, 
        P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN, 
        P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN, 
        P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN, 
        P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN, 
        P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, 
        P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN, 
        P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN, 
        P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN, 
        P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN, 
        P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN, 
        P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, keyinput_f0, 
        keyinput_f1, keyinput_f2, keyinput_f3, keyinput_f4, keyinput_f5, 
        keyinput_f6, keyinput_f7, keyinput_f8, keyinput_f9, keyinput_f10, 
        keyinput_f11, keyinput_f12, keyinput_f13, keyinput_f14, keyinput_f15, 
        keyinput_f16, keyinput_f17, keyinput_f18, keyinput_f19, keyinput_f20, 
        keyinput_f21, keyinput_f22, keyinput_f23, keyinput_f24, keyinput_f25, 
        keyinput_f26, keyinput_f27, keyinput_f28, keyinput_f29, keyinput_f30, 
        keyinput_f31, keyinput_f32, keyinput_f33, keyinput_f34, keyinput_f35, 
        keyinput_f36, keyinput_f37, keyinput_f38, keyinput_f39, keyinput_f40, 
        keyinput_f41, keyinput_f42, keyinput_f43, keyinput_f44, keyinput_f45, 
        keyinput_f46, keyinput_f47, keyinput_f48, keyinput_f49, keyinput_f50, 
        keyinput_f51, keyinput_f52, keyinput_f53, keyinput_f54, keyinput_f55, 
        keyinput_f56, keyinput_f57, keyinput_f58, keyinput_f59, keyinput_f60, 
        keyinput_f61, keyinput_f62, keyinput_f63, keyinput_f64, keyinput_f65, 
        keyinput_f66, keyinput_f67, keyinput_f68, keyinput_f69, keyinput_f70, 
        keyinput_f71, keyinput_f72, keyinput_f73, keyinput_f74, keyinput_f75, 
        keyinput_f76, keyinput_f77, keyinput_f78, keyinput_f79, keyinput_f80, 
        keyinput_f81, keyinput_f82, keyinput_f83, keyinput_f84, keyinput_f85, 
        keyinput_f86, keyinput_f87, keyinput_f88, keyinput_f89, keyinput_f90, 
        keyinput_f91, keyinput_f92, keyinput_f93, keyinput_f94, keyinput_f95, 
        keyinput_f96, keyinput_f97, keyinput_f98, keyinput_f99, keyinput_f100, 
        keyinput_f101, keyinput_f102, keyinput_f103, keyinput_f104, 
        keyinput_f105, keyinput_f106, keyinput_f107, keyinput_f108, 
        keyinput_f109, keyinput_f110, keyinput_f111, keyinput_f112, 
        keyinput_f113, keyinput_f114, keyinput_f115, keyinput_f116, 
        keyinput_f117, keyinput_f118, keyinput_f119, keyinput_f120, 
        keyinput_f121, keyinput_f122, keyinput_f123, keyinput_f124, 
        keyinput_f125, keyinput_f126, keyinput_f127, keyinput_g0, keyinput_g1, 
        keyinput_g2, keyinput_g3, keyinput_g4, keyinput_g5, keyinput_g6, 
        keyinput_g7, keyinput_g8, keyinput_g9, keyinput_g10, keyinput_g11, 
        keyinput_g12, keyinput_g13, keyinput_g14, keyinput_g15, keyinput_g16, 
        keyinput_g17, keyinput_g18, keyinput_g19, keyinput_g20, keyinput_g21, 
        keyinput_g22, keyinput_g23, keyinput_g24, keyinput_g25, keyinput_g26, 
        keyinput_g27, keyinput_g28, keyinput_g29, keyinput_g30, keyinput_g31, 
        keyinput_g32, keyinput_g33, keyinput_g34, keyinput_g35, keyinput_g36, 
        keyinput_g37, keyinput_g38, keyinput_g39, keyinput_g40, keyinput_g41, 
        keyinput_g42, keyinput_g43, keyinput_g44, keyinput_g45, keyinput_g46, 
        keyinput_g47, keyinput_g48, keyinput_g49, keyinput_g50, keyinput_g51, 
        keyinput_g52, keyinput_g53, keyinput_g54, keyinput_g55, keyinput_g56, 
        keyinput_g57, keyinput_g58, keyinput_g59, keyinput_g60, keyinput_g61, 
        keyinput_g62, keyinput_g63, keyinput_g64, keyinput_g65, keyinput_g66, 
        keyinput_g67, keyinput_g68, keyinput_g69, keyinput_g70, keyinput_g71, 
        keyinput_g72, keyinput_g73, keyinput_g74, keyinput_g75, keyinput_g76, 
        keyinput_g77, keyinput_g78, keyinput_g79, keyinput_g80, keyinput_g81, 
        keyinput_g82, keyinput_g83, keyinput_g84, keyinput_g85, keyinput_g86, 
        keyinput_g87, keyinput_g88, keyinput_g89, keyinput_g90, keyinput_g91, 
        keyinput_g92, keyinput_g93, keyinput_g94, keyinput_g95, keyinput_g96, 
        keyinput_g97, keyinput_g98, keyinput_g99, keyinput_g100, keyinput_g101, 
        keyinput_g102, keyinput_g103, keyinput_g104, keyinput_g105, 
        keyinput_g106, keyinput_g107, keyinput_g108, keyinput_g109, 
        keyinput_g110, keyinput_g111, keyinput_g112, keyinput_g113, 
        keyinput_g114, keyinput_g115, keyinput_g116, keyinput_g117, 
        keyinput_g118, keyinput_g119, keyinput_g120, keyinput_g121, 
        keyinput_g122, keyinput_g123, keyinput_g124, keyinput_g125, 
        keyinput_g126, keyinput_g127, ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, 
        ADD_1068_U57, ADD_1068_U58, ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, 
        ADD_1068_U62, ADD_1068_U63, ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, 
        ADD_1068_U50, ADD_1068_U51, ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, 
        ADD_1068_U5, ADD_1068_U46, U126, U123, P1_U3355, P1_U3354, P1_U3353, 
        P1_U3352, P1_U3351, P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, 
        P1_U3345, P1_U3344, P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, 
        P1_U3338, P1_U3337, P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, 
        P1_U3331, P1_U3330, P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, 
        P1_U3324, P1_U3439, P1_U3440, P1_U3323, P1_U3322, P1_U3321, P1_U3320, 
        P1_U3319, P1_U3318, P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, 
        P1_U3312, P1_U3311, P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, 
        P1_U3305, P1_U3304, P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, 
        P1_U3298, P1_U3297, P1_U3296, P1_U3295, P1_U3294, P1_U3453, P1_U3456, 
        P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, 
        P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, 
        P1_U3501, P1_U3504, P1_U3507, P1_U3509, P1_U3510, P1_U3511, P1_U3512, 
        P1_U3513, P1_U3514, P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, 
        P1_U3520, P1_U3521, P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, 
        P1_U3527, P1_U3528, P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, 
        P1_U3534, P1_U3535, P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, 
        P1_U3541, P1_U3542, P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, 
        P1_U3548, P1_U3549, P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3293, 
        P1_U3292, P1_U3291, P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, 
        P1_U3285, P1_U3284, P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, 
        P1_U3278, P1_U3277, P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, 
        P1_U3271, P1_U3270, P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, 
        P1_U3356, P1_U3264, P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, 
        P1_U3258, P1_U3257, P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, 
        P1_U3251, P1_U3250, P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, 
        P1_U3244, P1_U3243, P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, 
        P1_U3559, P1_U3560, P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, 
        P1_U3566, P1_U3567, P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, 
        P1_U3573, P1_U3574, P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, 
        P1_U3580, P1_U3581, P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3242, 
        P1_U3241, P1_U3240, P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, 
        P1_U3234, P1_U3233, P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, 
        P1_U3227, P1_U3226, P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, 
        P1_U3220, P1_U3219, P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, 
        P1_U3213, P1_U3086, P1_U3085, P1_U3973, P2_U3295, P2_U3294, P2_U3293, 
        P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, 
        P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, 
        P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, 
        P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, 
        P2_U3264, P2_U3376, P2_U3377, P2_U3263, P2_U3262, P2_U3261, P2_U3260, 
        P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, 
        P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, 
        P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, 
        P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3390, P2_U3393, 
        P2_U3396, P2_U3399, P2_U3402, P2_U3405, P2_U3408, P2_U3411, P2_U3414, 
        P2_U3417, P2_U3420, P2_U3423, P2_U3426, P2_U3429, P2_U3432, P2_U3435, 
        P2_U3438, P2_U3441, P2_U3444, P2_U3446, P2_U3447, P2_U3448, P2_U3449, 
        P2_U3450, P2_U3451, P2_U3452, P2_U3453, P2_U3454, P2_U3455, P2_U3456, 
        P2_U3457, P2_U3458, P2_U3459, P2_U3460, P2_U3461, P2_U3462, P2_U3463, 
        P2_U3464, P2_U3465, P2_U3466, P2_U3467, P2_U3468, P2_U3469, P2_U3470, 
        P2_U3471, P2_U3472, P2_U3473, P2_U3474, P2_U3475, P2_U3476, P2_U3477, 
        P2_U3478, P2_U3479, P2_U3480, P2_U3481, P2_U3482, P2_U3483, P2_U3484, 
        P2_U3485, P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3233, 
        P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, 
        P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, 
        P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, 
        P2_U3211, P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, 
        P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, 
        P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, 
        P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3184, 
        P2_U3183, P2_U3182, P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, 
        P2_U3496, P2_U3497, P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, 
        P2_U3503, P2_U3504, P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, 
        P2_U3510, P2_U3511, P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, 
        P2_U3517, P2_U3518, P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3296, 
        P2_U3181, P2_U3180, P2_U3179, P2_U3178, P2_U3177, P2_U3176, P2_U3175, 
        P2_U3174, P2_U3173, P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, 
        P2_U3167, P2_U3166, P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, 
        P2_U3160, P2_U3159, P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, 
        P2_U3153, P2_U3151, P2_U3150, P2_U3893 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN,
         P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN,
         P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN,
         P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN,
         P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN,
         P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN,
         P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN,
         P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN,
         P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN,
         P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN,
         P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN,
         P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN,
         P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN,
         P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN,
         P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN,
         P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN,
         P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN,
         P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN,
         P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN,
         P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN,
         P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN,
         P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN,
         P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN,
         P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN,
         P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN,
         P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN,
         P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN,
         P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN,
         P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN,
         P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN,
         P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN,
         P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN,
         P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN,
         P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN,
         P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN,
         P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN,
         P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN,
         P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN,
         P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN,
         P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN,
         P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN,
         P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN,
         P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN,
         P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN,
         P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN,
         P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN,
         P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN,
         P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN,
         P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN,
         P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN,
         P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN,
         P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN,
         P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN,
         P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN,
         P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN,
         P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN,
         P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN,
         P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN,
         P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN,
         P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN,
         P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN,
         P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN,
         P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN,
         P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN,
         P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN,
         P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN,
         P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN,
         P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN,
         P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN,
         P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN,
         P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN,
         P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN,
         P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN,
         P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN,
         P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN,
         P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN,
         P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN,
         P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN,
         P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN,
         P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN,
         P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN,
         P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN,
         P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN,
         P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN,
         P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN,
         P1_REG3_REG_4__SCAN_IN, P1_REG3_REG_24__SCAN_IN,
         P1_REG3_REG_17__SCAN_IN, P1_REG3_REG_5__SCAN_IN,
         P1_REG3_REG_16__SCAN_IN, P1_REG3_REG_25__SCAN_IN,
         P1_REG3_REG_12__SCAN_IN, P1_REG3_REG_21__SCAN_IN,
         P1_REG3_REG_1__SCAN_IN, P1_REG3_REG_8__SCAN_IN,
         P1_REG3_REG_28__SCAN_IN, P1_REG3_REG_19__SCAN_IN,
         P1_REG3_REG_3__SCAN_IN, P1_REG3_REG_10__SCAN_IN,
         P1_REG3_REG_23__SCAN_IN, P1_REG3_REG_14__SCAN_IN,
         P1_REG3_REG_27__SCAN_IN, P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN,
         P1_RD_REG_SCAN_IN, P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN,
         P2_IR_REG_1__SCAN_IN, P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN,
         P2_IR_REG_4__SCAN_IN, P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN,
         P2_IR_REG_7__SCAN_IN, P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN,
         P2_IR_REG_10__SCAN_IN, P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN,
         P2_IR_REG_13__SCAN_IN, P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN,
         P2_IR_REG_16__SCAN_IN, P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN,
         P2_IR_REG_19__SCAN_IN, P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN,
         P2_IR_REG_22__SCAN_IN, P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN,
         P2_IR_REG_25__SCAN_IN, P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN,
         P2_IR_REG_28__SCAN_IN, P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN,
         P2_IR_REG_31__SCAN_IN, P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN,
         P2_D_REG_2__SCAN_IN, P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN,
         P2_D_REG_5__SCAN_IN, P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN,
         P2_D_REG_8__SCAN_IN, P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN,
         P2_D_REG_11__SCAN_IN, P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN,
         P2_D_REG_14__SCAN_IN, P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN,
         P2_D_REG_17__SCAN_IN, P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN,
         P2_D_REG_20__SCAN_IN, P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN,
         P2_D_REG_23__SCAN_IN, P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN,
         P2_D_REG_26__SCAN_IN, P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN,
         P2_D_REG_29__SCAN_IN, P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN,
         P2_REG0_REG_0__SCAN_IN, P2_REG0_REG_1__SCAN_IN,
         P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN,
         P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN,
         P2_REG0_REG_6__SCAN_IN, P2_REG0_REG_7__SCAN_IN,
         P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN,
         P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN,
         P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN,
         P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN,
         P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN,
         P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN,
         P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN,
         P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN,
         P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN,
         P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN,
         P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN,
         P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN,
         P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN,
         P2_REG1_REG_2__SCAN_IN, P2_REG1_REG_3__SCAN_IN,
         P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN,
         P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN,
         P2_REG1_REG_8__SCAN_IN, P2_REG1_REG_9__SCAN_IN,
         P2_REG1_REG_10__SCAN_IN, P2_REG1_REG_11__SCAN_IN,
         P2_REG1_REG_12__SCAN_IN, P2_REG1_REG_13__SCAN_IN,
         P2_REG1_REG_14__SCAN_IN, P2_REG1_REG_15__SCAN_IN,
         P2_REG1_REG_16__SCAN_IN, P2_REG1_REG_17__SCAN_IN,
         P2_REG1_REG_18__SCAN_IN, P2_REG1_REG_19__SCAN_IN,
         P2_REG1_REG_20__SCAN_IN, P2_REG1_REG_21__SCAN_IN,
         P2_REG1_REG_22__SCAN_IN, P2_REG1_REG_23__SCAN_IN,
         P2_REG1_REG_24__SCAN_IN, P2_REG1_REG_25__SCAN_IN,
         P2_REG1_REG_26__SCAN_IN, P2_REG1_REG_27__SCAN_IN,
         P2_REG1_REG_28__SCAN_IN, P2_REG1_REG_29__SCAN_IN,
         P2_REG1_REG_30__SCAN_IN, P2_REG1_REG_31__SCAN_IN,
         P2_REG2_REG_0__SCAN_IN, P2_REG2_REG_1__SCAN_IN,
         P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN,
         P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN,
         P2_REG2_REG_6__SCAN_IN, P2_REG2_REG_7__SCAN_IN,
         P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN,
         P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN,
         P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN,
         P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN,
         P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN,
         P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN,
         P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN,
         P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN,
         P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN,
         P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN,
         P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN,
         P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN,
         P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN,
         P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN,
         P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN,
         P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN,
         P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN,
         P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN,
         P2_ADDR_REG_7__SCAN_IN, P2_ADDR_REG_6__SCAN_IN,
         P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN,
         P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN,
         P2_ADDR_REG_1__SCAN_IN, P2_ADDR_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, keyinput_f0, keyinput_f1, keyinput_f2,
         keyinput_f3, keyinput_f4, keyinput_f5, keyinput_f6, keyinput_f7,
         keyinput_f8, keyinput_f9, keyinput_f10, keyinput_f11, keyinput_f12,
         keyinput_f13, keyinput_f14, keyinput_f15, keyinput_f16, keyinput_f17,
         keyinput_f18, keyinput_f19, keyinput_f20, keyinput_f21, keyinput_f22,
         keyinput_f23, keyinput_f24, keyinput_f25, keyinput_f26, keyinput_f27,
         keyinput_f28, keyinput_f29, keyinput_f30, keyinput_f31, keyinput_f32,
         keyinput_f33, keyinput_f34, keyinput_f35, keyinput_f36, keyinput_f37,
         keyinput_f38, keyinput_f39, keyinput_f40, keyinput_f41, keyinput_f42,
         keyinput_f43, keyinput_f44, keyinput_f45, keyinput_f46, keyinput_f47,
         keyinput_f48, keyinput_f49, keyinput_f50, keyinput_f51, keyinput_f52,
         keyinput_f53, keyinput_f54, keyinput_f55, keyinput_f56, keyinput_f57,
         keyinput_f58, keyinput_f59, keyinput_f60, keyinput_f61, keyinput_f62,
         keyinput_f63, keyinput_f64, keyinput_f65, keyinput_f66, keyinput_f67,
         keyinput_f68, keyinput_f69, keyinput_f70, keyinput_f71, keyinput_f72,
         keyinput_f73, keyinput_f74, keyinput_f75, keyinput_f76, keyinput_f77,
         keyinput_f78, keyinput_f79, keyinput_f80, keyinput_f81, keyinput_f82,
         keyinput_f83, keyinput_f84, keyinput_f85, keyinput_f86, keyinput_f87,
         keyinput_f88, keyinput_f89, keyinput_f90, keyinput_f91, keyinput_f92,
         keyinput_f93, keyinput_f94, keyinput_f95, keyinput_f96, keyinput_f97,
         keyinput_f98, keyinput_f99, keyinput_f100, keyinput_f101,
         keyinput_f102, keyinput_f103, keyinput_f104, keyinput_f105,
         keyinput_f106, keyinput_f107, keyinput_f108, keyinput_f109,
         keyinput_f110, keyinput_f111, keyinput_f112, keyinput_f113,
         keyinput_f114, keyinput_f115, keyinput_f116, keyinput_f117,
         keyinput_f118, keyinput_f119, keyinput_f120, keyinput_f121,
         keyinput_f122, keyinput_f123, keyinput_f124, keyinput_f125,
         keyinput_f126, keyinput_f127, keyinput_g0, keyinput_g1, keyinput_g2,
         keyinput_g3, keyinput_g4, keyinput_g5, keyinput_g6, keyinput_g7,
         keyinput_g8, keyinput_g9, keyinput_g10, keyinput_g11, keyinput_g12,
         keyinput_g13, keyinput_g14, keyinput_g15, keyinput_g16, keyinput_g17,
         keyinput_g18, keyinput_g19, keyinput_g20, keyinput_g21, keyinput_g22,
         keyinput_g23, keyinput_g24, keyinput_g25, keyinput_g26, keyinput_g27,
         keyinput_g28, keyinput_g29, keyinput_g30, keyinput_g31, keyinput_g32,
         keyinput_g33, keyinput_g34, keyinput_g35, keyinput_g36, keyinput_g37,
         keyinput_g38, keyinput_g39, keyinput_g40, keyinput_g41, keyinput_g42,
         keyinput_g43, keyinput_g44, keyinput_g45, keyinput_g46, keyinput_g47,
         keyinput_g48, keyinput_g49, keyinput_g50, keyinput_g51, keyinput_g52,
         keyinput_g53, keyinput_g54, keyinput_g55, keyinput_g56, keyinput_g57,
         keyinput_g58, keyinput_g59, keyinput_g60, keyinput_g61, keyinput_g62,
         keyinput_g63, keyinput_g64, keyinput_g65, keyinput_g66, keyinput_g67,
         keyinput_g68, keyinput_g69, keyinput_g70, keyinput_g71, keyinput_g72,
         keyinput_g73, keyinput_g74, keyinput_g75, keyinput_g76, keyinput_g77,
         keyinput_g78, keyinput_g79, keyinput_g80, keyinput_g81, keyinput_g82,
         keyinput_g83, keyinput_g84, keyinput_g85, keyinput_g86, keyinput_g87,
         keyinput_g88, keyinput_g89, keyinput_g90, keyinput_g91, keyinput_g92,
         keyinput_g93, keyinput_g94, keyinput_g95, keyinput_g96, keyinput_g97,
         keyinput_g98, keyinput_g99, keyinput_g100, keyinput_g101,
         keyinput_g102, keyinput_g103, keyinput_g104, keyinput_g105,
         keyinput_g106, keyinput_g107, keyinput_g108, keyinput_g109,
         keyinput_g110, keyinput_g111, keyinput_g112, keyinput_g113,
         keyinput_g114, keyinput_g115, keyinput_g116, keyinput_g117,
         keyinput_g118, keyinput_g119, keyinput_g120, keyinput_g121,
         keyinput_g122, keyinput_g123, keyinput_g124, keyinput_g125,
         keyinput_g126, keyinput_g127;
  output ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58,
         ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63,
         ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51,
         ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46,
         U126, U123, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351,
         P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344,
         P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337,
         P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330,
         P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439,
         P1_U3440, P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318,
         P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311,
         P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304,
         P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297,
         P1_U3296, P1_U3295, P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462,
         P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483,
         P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504,
         P1_U3507, P1_U3509, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291,
         P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284,
         P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277,
         P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270,
         P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264,
         P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257,
         P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250,
         P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243,
         P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240,
         P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233,
         P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226,
         P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219,
         P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086,
         P1_U3085, P1_U3973, P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291,
         P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284,
         P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277,
         P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270,
         P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376,
         P2_U3377, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258,
         P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251,
         P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244,
         P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237,
         P2_U3236, P2_U3235, P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399,
         P2_U3402, P2_U3405, P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420,
         P2_U3423, P2_U3426, P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441,
         P2_U3444, P2_U3446, P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451,
         P2_U3452, P2_U3453, P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458,
         P2_U3459, P2_U3460, P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465,
         P2_U3466, P2_U3467, P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472,
         P2_U3473, P2_U3474, P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479,
         P2_U3480, P2_U3481, P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486,
         P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231,
         P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224,
         P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217,
         P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210,
         P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203,
         P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196,
         P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189,
         P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182,
         P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497,
         P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504,
         P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511,
         P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518,
         P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180,
         P2_U3179, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173,
         P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166,
         P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159,
         P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151,
         P2_U3150, P2_U3893;
  wire   n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516,
         n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526,
         n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536,
         n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546,
         n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556,
         n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566,
         n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576,
         n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586,
         n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596,
         n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606,
         n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616,
         n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626,
         n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636,
         n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646,
         n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656,
         n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666,
         n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676,
         n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686,
         n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696,
         n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706,
         n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716,
         n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726,
         n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736,
         n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746,
         n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756,
         n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766,
         n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776,
         n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786,
         n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796,
         n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806,
         n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816,
         n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826,
         n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836,
         n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846,
         n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856,
         n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866,
         n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876,
         n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886,
         n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896,
         n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906,
         n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916,
         n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926,
         n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936,
         n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946,
         n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956,
         n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966,
         n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976,
         n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986,
         n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996,
         n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006,
         n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016,
         n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026,
         n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036,
         n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046,
         n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056,
         n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066,
         n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076,
         n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086,
         n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096,
         n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106,
         n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116,
         n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126,
         n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136,
         n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146,
         n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156,
         n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166,
         n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176,
         n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186,
         n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196,
         n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206,
         n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216,
         n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226,
         n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236,
         n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246,
         n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256,
         n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266,
         n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276,
         n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286,
         n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296,
         n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306,
         n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316,
         n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326,
         n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336,
         n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346,
         n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356,
         n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366,
         n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376,
         n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386,
         n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396,
         n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406,
         n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416,
         n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426,
         n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436,
         n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446,
         n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456,
         n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466,
         n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476,
         n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486,
         n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496,
         n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506,
         n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516,
         n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526,
         n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536,
         n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546,
         n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556,
         n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566,
         n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576,
         n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586,
         n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596,
         n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606,
         n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616,
         n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626,
         n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636,
         n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646,
         n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656,
         n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666,
         n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676,
         n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686,
         n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696,
         n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706,
         n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716,
         n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726,
         n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736,
         n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746,
         n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756,
         n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766,
         n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776,
         n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786,
         n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796,
         n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806,
         n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816,
         n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826,
         n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836,
         n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846,
         n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856,
         n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866,
         n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876,
         n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886,
         n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896,
         n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906,
         n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916,
         n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926,
         n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936,
         n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946,
         n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956,
         n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966,
         n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976,
         n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986,
         n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996,
         n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006,
         n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016,
         n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026,
         n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036,
         n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046,
         n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056,
         n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066,
         n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076,
         n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086,
         n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096,
         n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106,
         n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116,
         n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126,
         n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136,
         n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146,
         n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156,
         n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166,
         n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176,
         n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186,
         n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196,
         n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206,
         n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216,
         n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226,
         n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236,
         n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246,
         n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256,
         n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266,
         n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276,
         n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286,
         n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296,
         n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306,
         n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316,
         n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326,
         n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336,
         n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346,
         n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356,
         n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366,
         n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376,
         n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386,
         n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396,
         n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406,
         n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416,
         n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426,
         n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436,
         n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446,
         n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456,
         n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466,
         n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476,
         n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486,
         n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496,
         n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506,
         n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516,
         n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526,
         n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536,
         n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546,
         n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556,
         n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566,
         n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576,
         n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586,
         n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596,
         n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606,
         n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616,
         n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626,
         n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636,
         n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646,
         n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656,
         n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666,
         n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676,
         n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686,
         n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696,
         n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706,
         n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716,
         n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726,
         n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736,
         n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746,
         n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756,
         n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766,
         n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776,
         n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786,
         n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796,
         n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806,
         n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816,
         n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826,
         n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836,
         n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846,
         n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856,
         n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866,
         n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876,
         n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886,
         n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896,
         n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906,
         n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916,
         n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926,
         n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936,
         n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946,
         n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956,
         n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966,
         n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976,
         n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986,
         n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996,
         n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006,
         n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016,
         n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026,
         n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036,
         n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046,
         n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056,
         n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066,
         n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076,
         n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086,
         n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096,
         n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106,
         n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116,
         n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126,
         n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136,
         n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146,
         n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156,
         n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166,
         n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176,
         n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186,
         n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196,
         n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206,
         n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216,
         n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226,
         n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236,
         n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246,
         n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256,
         n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266,
         n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276,
         n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286,
         n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296,
         n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306,
         n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316,
         n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326,
         n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336,
         n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346,
         n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356,
         n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366,
         n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376,
         n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386,
         n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396,
         n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406,
         n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416,
         n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426,
         n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436,
         n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446,
         n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456,
         n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466,
         n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476,
         n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486,
         n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496,
         n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506,
         n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516,
         n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526,
         n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536,
         n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546,
         n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556,
         n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566,
         n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576,
         n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586,
         n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596,
         n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606,
         n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616,
         n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626,
         n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636,
         n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646,
         n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656,
         n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666,
         n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676,
         n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686,
         n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696,
         n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706,
         n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716,
         n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726,
         n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736,
         n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746,
         n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756,
         n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766,
         n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776,
         n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786,
         n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796,
         n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806,
         n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816,
         n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826,
         n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836,
         n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846,
         n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856,
         n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866,
         n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876,
         n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886,
         n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896,
         n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906,
         n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916,
         n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926,
         n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936,
         n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946,
         n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956,
         n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966,
         n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976,
         n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986,
         n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996,
         n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006,
         n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016,
         n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026,
         n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036,
         n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046,
         n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056,
         n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066,
         n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076,
         n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086,
         n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096,
         n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106,
         n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116,
         n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126,
         n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136,
         n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146,
         n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156,
         n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166,
         n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176,
         n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186,
         n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196,
         n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206,
         n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216,
         n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226,
         n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236,
         n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246,
         n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256,
         n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266,
         n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276,
         n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286,
         n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296,
         n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306,
         n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316,
         n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326,
         n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336,
         n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346,
         n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356,
         n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366,
         n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376,
         n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386,
         n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396,
         n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406,
         n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416,
         n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426,
         n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436,
         n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446,
         n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456,
         n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466,
         n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476,
         n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486,
         n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496,
         n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506,
         n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516,
         n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526,
         n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536,
         n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546,
         n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556,
         n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566,
         n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576,
         n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586,
         n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596,
         n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606,
         n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616,
         n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626,
         n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636,
         n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646,
         n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656,
         n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666,
         n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676,
         n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686,
         n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696,
         n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706,
         n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716,
         n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726,
         n8727, n8728, n8729, n8730, n8731, n8733, n8734, n8735, n8736, n8737,
         n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747,
         n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757,
         n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767,
         n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777,
         n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787,
         n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797,
         n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807,
         n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817,
         n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827,
         n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837,
         n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847,
         n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857,
         n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867,
         n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877,
         n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887,
         n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897,
         n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907,
         n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917,
         n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927,
         n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937,
         n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947,
         n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957,
         n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967,
         n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977,
         n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987,
         n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997,
         n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007,
         n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017,
         n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027,
         n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037,
         n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047,
         n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057,
         n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067,
         n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077,
         n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087,
         n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097,
         n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107,
         n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117,
         n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127,
         n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137,
         n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147,
         n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157,
         n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167,
         n9168, n9169, n9170, n9171, n9173, n9174, n9175, n9176, n9177, n9178,
         n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188,
         n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198,
         n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208,
         n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218,
         n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228,
         n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238,
         n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248,
         n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258,
         n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268,
         n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278,
         n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288,
         n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298,
         n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308,
         n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318,
         n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328,
         n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338,
         n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348,
         n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358,
         n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368,
         n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378,
         n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388,
         n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398,
         n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408,
         n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418,
         n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428,
         n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438,
         n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448,
         n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458,
         n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468,
         n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478,
         n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488,
         n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498,
         n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508,
         n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518,
         n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528,
         n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538,
         n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548,
         n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558,
         n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568,
         n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578,
         n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588,
         n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598,
         n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608,
         n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618,
         n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628,
         n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638,
         n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648,
         n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658,
         n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668,
         n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678,
         n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688,
         n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698,
         n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708,
         n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718,
         n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728,
         n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738,
         n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748,
         n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758,
         n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768,
         n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778,
         n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788,
         n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798,
         n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808,
         n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818,
         n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828,
         n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838,
         n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848,
         n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858,
         n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868,
         n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878,
         n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888,
         n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898,
         n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908,
         n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918,
         n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928,
         n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938,
         n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948,
         n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958,
         n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968,
         n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978,
         n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988,
         n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998,
         n9999, n10000, n10001, n10002, n10003, n10004, n10005, n10006, n10007,
         n10008, n10009, n10010, n10011, n10012, n10013, n10014, n10015,
         n10016, n10017, n10018, n10019, n10020, n10021, n10022, n10023,
         n10024, n10025, n10026, n10027, n10028, n10029, n10030, n10031,
         n10032, n10033, n10034, n10035, n10036, n10037, n10038, n10039,
         n10040, n10041, n10042, n10043, n10044, n10045, n10046, n10047,
         n10048, n10049, n10050, n10051, n10052, n10053, n10054, n10055,
         n10056, n10057, n10058, n10059, n10060, n10061, n10062, n10063,
         n10064, n10065, n10066, n10067, n10068, n10069, n10070, n10071,
         n10072, n10073, n10074, n10075, n10076, n10077, n10078, n10079,
         n10080, n10081, n10082, n10083, n10084, n10085, n10086, n10087,
         n10088, n10089, n10090, n10091, n10092, n10093, n10094, n10095,
         n10096, n10097, n10098, n10099, n10100, n10101, n10102, n10103,
         n10104, n10105, n10106, n10107, n10108, n10109, n10110, n10111,
         n10112, n10113, n10114, n10115, n10116, n10117, n10118, n10119,
         n10120, n10121, n10122, n10123, n10124, n10125, n10126, n10127,
         n10128, n10129, n10130, n10131, n10132, n10133, n10134, n10135,
         n10136, n10137, n10138, n10139, n10140, n10141, n10142, n10143,
         n10144, n10145, n10146, n10147, n10148, n10149, n10150, n10151,
         n10152, n10153, n10154, n10155, n10156, n10157, n10158, n10159,
         n10160, n10161, n10162, n10163, n10164, n10165, n10166, n10167,
         n10168, n10169, n10170, n10171, n10172, n10173, n10174, n10175,
         n10176, n10177, n10178, n10179, n10180, n10181, n10182, n10183,
         n10184, n10185, n10186, n10187, n10188, n10189, n10190, n10191,
         n10192, n10193, n10194, n10195, n10196, n10197, n10198, n10199,
         n10200, n10201, n10202, n10203, n10204, n10205, n10206, n10207,
         n10208, n10209, n10210, n10211, n10212, n10213, n10214, n10215,
         n10216, n10217, n10218, n10219, n10220, n10221, n10222, n10223,
         n10224, n10225, n10226, n10227, n10228, n10229, n10230, n10231,
         n10232, n10233, n10234, n10235, n10236, n10237, n10238, n10239,
         n10240, n10241, n10242, n10243, n10244, n10245, n10246, n10247,
         n10248, n10249, n10250, n10251, n10252, n10253, n10254, n10255,
         n10256, n10257, n10258, n10259, n10260, n10261, n10262, n10263,
         n10264, n10265, n10266, n10267, n10268, n10269, n10270, n10271,
         n10272, n10273, n10274, n10275, n10276, n10277, n10278, n10279,
         n10280, n10281, n10282, n10283, n10284, n10285, n10286, n10287,
         n10288, n10289, n10290, n10291, n10292, n10293, n10294, n10295,
         n10296, n10297, n10298, n10299, n10300, n10301, n10302, n10303,
         n10304, n10305, n10306, n10307, n10308, n10309, n10310, n10311,
         n10312, n10313, n10314, n10315, n10316, n10317, n10318, n10319,
         n10320, n10321, n10322, n10323, n10324, n10325, n10326, n10327,
         n10328, n10329, n10330, n10331, n10332, n10333, n10334, n10335,
         n10336, n10337, n10338, n10339, n10340, n10341, n10342, n10343,
         n10344, n10345, n10346, n10347, n10348, n10349, n10350, n10351,
         n10352, n10353, n10354, n10355, n10356, n10357, n10358, n10359,
         n10360, n10361, n10362, n10363, n10364, n10365, n10366, n10367,
         n10368, n10369, n10370, n10371, n10372, n10373, n10374, n10375,
         n10376, n10377, n10378, n10379, n10380, n10381, n10382, n10383,
         n10384, n10385, n10386, n10387, n10388, n10389, n10390, n10391,
         n10392, n10393, n10394, n10395, n10396, n10397, n10398, n10399,
         n10400, n10401, n10402, n10403, n10404, n10405, n10406, n10407,
         n10408, n10409, n10410, n10411, n10412, n10413, n10414, n10415,
         n10416, n10417, n10418, n10419, n10420, n10421, n10422, n10423,
         n10424, n10425, n10426, n10427, n10428, n10429, n10430, n10431,
         n10432, n10433, n10434, n10435, n10436, n10437, n10438, n10439,
         n10440, n10441, n10442, n10443, n10444, n10445, n10446, n10447,
         n10448, n10449, n10450, n10451, n10452, n10453, n10454, n10455,
         n10456, n10457, n10458, n10459, n10460, n10461, n10462, n10463,
         n10464, n10465, n10466, n10467, n10468, n10469, n10470, n10471,
         n10472, n10473, n10474, n10475, n10476, n10477, n10478, n10479,
         n10480, n10481, n10482, n10483, n10484, n10485, n10486, n10487,
         n10488, n10489, n10490, n10491, n10492, n10493, n10494, n10495,
         n10496, n10497, n10498, n10499, n10500, n10501, n10502, n10503,
         n10504, n10505, n10506, n10507, n10508, n10509, n10510, n10511,
         n10512, n10513, n10514, n10515, n10516, n10517, n10518, n10519,
         n10520, n10521, n10522, n10523, n10524, n10525, n10526, n10527,
         n10528, n10529, n10530, n10531, n10532, n10533, n10534, n10535,
         n10536, n10537, n10538, n10539, n10540, n10541, n10542, n10543,
         n10544, n10545, n10546, n10547, n10548, n10549, n10550, n10551,
         n10552, n10553, n10554, n10555, n10556, n10557, n10558, n10559,
         n10560, n10561, n10562, n10563, n10564, n10565, n10566, n10567,
         n10568, n10569, n10570, n10571, n10572, n10573, n10574, n10575,
         n10576, n10577, n10578, n10579, n10580, n10581, n10582, n10583,
         n10584, n10585, n10586, n10587, n10588, n10589, n10590, n10591,
         n10592, n10593, n10594, n10595, n10596, n10597, n10598, n10599,
         n10600, n10601, n10602, n10603, n10604, n10605, n10606, n10607,
         n10608, n10609, n10610, n10611, n10612, n10613, n10614, n10615,
         n10616, n10617, n10618, n10619, n10620, n10621, n10622, n10623,
         n10624, n10625, n10626, n10627, n10628, n10629, n10630, n10631,
         n10632, n10633, n10634, n10635, n10636, n10637, n10638, n10639,
         n10640, n10641, n10642, n10643, n10644, n10645, n10646, n10647,
         n10648, n10649, n10650, n10651, n10652, n10653, n10654, n10655,
         n10656, n10657, n10658, n10659, n10660, n10661, n10662, n10663,
         n10664, n10665, n10666;

  NOR2_X1 U5013 ( .A1(n7406), .A2(n7396), .ZN(n7397) );
  NAND2_X1 U5014 ( .A1(n5494), .A2(n5493), .ZN(n10197) );
  INV_X1 U5015 ( .A(n5339), .ZN(n8198) );
  CLKBUF_X2 U5016 ( .A(n5358), .Z(n4507) );
  NAND3_X1 U5017 ( .A1(n5950), .A2(n5949), .A3(n5948), .ZN(n7257) );
  OR3_X2 U5018 ( .A1(n6411), .A2(n7899), .A3(n7919), .ZN(n5925) );
  INV_X1 U5019 ( .A(n6619), .ZN(n9206) );
  OR2_X1 U5020 ( .A1(n5824), .A2(n8584), .ZN(n8212) );
  INV_X1 U5021 ( .A(n8203), .ZN(n8174) );
  CLKBUF_X3 U5022 ( .A(n9736), .Z(n4515) );
  INV_X1 U5023 ( .A(n5635), .ZN(n7535) );
  AND2_X1 U5024 ( .A1(n5784), .A2(n5783), .ZN(n4694) );
  INV_X1 U5025 ( .A(n7431), .ZN(n7011) );
  AND2_X1 U5026 ( .A1(n7652), .A2(n4761), .ZN(n9754) );
  AOI21_X1 U5027 ( .B1(n6691), .B2(n6501), .A(n4633), .ZN(n10060) );
  NAND2_X1 U5028 ( .A1(n6536), .A2(n6535), .ZN(n9961) );
  INV_X1 U5029 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n5848) );
  XNOR2_X1 U5030 ( .A(n10197), .B(n7940), .ZN(n8236) );
  CLKBUF_X3 U5031 ( .A(n9642), .Z(n4509) );
  XNOR2_X1 U5032 ( .A(n5850), .B(n5849), .ZN(n6411) );
  XNOR2_X1 U5033 ( .A(n4813), .B(P1_IR_REG_19__SCAN_IN), .ZN(n9642) );
  OAI21_X1 U5034 ( .B1(n7729), .B2(n4977), .A(n4975), .ZN(n7941) );
  NAND2_X4 U5035 ( .A1(n5925), .A2(n5867), .ZN(n9214) );
  OAI21_X2 U5036 ( .B1(n7832), .B2(n5010), .A(n5008), .ZN(n7920) );
  NAND2_X2 U5037 ( .A1(n6546), .A2(n6545), .ZN(n7832) );
  INV_X4 U5038 ( .A(n5382), .ZN(n5346) );
  AOI21_X2 U5039 ( .B1(n8846), .B2(n8845), .A(n8844), .ZN(n8854) );
  NAND2_X1 U5040 ( .A1(n5341), .A2(n6671), .ZN(n5358) );
  OAI222_X1 U5041 ( .A1(n9905), .A2(n7966), .B1(P1_U3086), .B2(n6411), .C1(
        n10530), .C2(n9903), .ZN(P1_U3329) );
  INV_X2 U5042 ( .A(n5875), .ZN(n9901) );
  NAND2_X4 U5043 ( .A1(n4747), .A2(n4746), .ZN(n5217) );
  INV_X2 U5044 ( .A(n10147), .ZN(n6841) );
  NAND2_X2 U5045 ( .A1(n5323), .A2(n5324), .ZN(n10147) );
  CLKBUF_X1 U5046 ( .A(n6506), .Z(n4508) );
  XNOR2_X1 U5047 ( .A(n5844), .B(n5843), .ZN(n6506) );
  AOI21_X2 U5048 ( .B1(n9275), .B2(n5131), .A(n5128), .ZN(n9231) );
  OAI21_X2 U5049 ( .B1(n7982), .B2(n7981), .A(n7980), .ZN(n8005) );
  CLKBUF_X1 U5050 ( .A(n8596), .Z(n8597) );
  NAND2_X1 U5051 ( .A1(n7546), .A2(n7547), .ZN(n7729) );
  OAI21_X1 U5052 ( .B1(n5469), .B2(n4786), .A(n4783), .ZN(n5520) );
  NAND4_X1 U5053 ( .A1(n5352), .A2(n5351), .A3(n5350), .A4(n5349), .ZN(n10149)
         );
  NOR2_X2 U5054 ( .A1(n7096), .A2(n10011), .ZN(n6586) );
  CLKBUF_X2 U5055 ( .A(P1_U3973), .Z(n4511) );
  NAND2_X2 U5056 ( .A1(n6768), .A2(n5225), .ZN(n5908) );
  NAND2_X2 U5058 ( .A1(n6442), .A2(n6506), .ZN(n6768) );
  INV_X1 U5059 ( .A(n5217), .ZN(n5225) );
  OR2_X1 U5060 ( .A1(n9848), .A2(n10100), .ZN(n9768) );
  NOR2_X1 U5061 ( .A1(n8512), .A2(n4740), .ZN(n8519) );
  AOI21_X1 U5062 ( .B1(n9253), .B2(n6408), .A(n6409), .ZN(n6454) );
  OR2_X1 U5063 ( .A1(n9554), .A2(n10034), .ZN(n4611) );
  MUX2_X1 U5064 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n9088), .S(n10199), .Z(n9092) );
  OAI21_X1 U5065 ( .B1(n9285), .B2(n5126), .A(n5123), .ZN(n6631) );
  AOI21_X1 U5066 ( .B1(n8505), .B2(n8504), .A(n4742), .ZN(n4741) );
  OR2_X1 U5067 ( .A1(n4541), .A2(n9195), .ZN(n9365) );
  AND2_X1 U5068 ( .A1(n4612), .A2(n4522), .ZN(n4608) );
  NAND2_X1 U5069 ( .A1(n6568), .A2(n6567), .ZN(n9565) );
  NOR2_X1 U5070 ( .A1(n4614), .A2(n6612), .ZN(n4613) );
  NAND2_X1 U5071 ( .A1(n8686), .A2(n8690), .ZN(n8563) );
  AOI211_X1 U5072 ( .C1(n9993), .C2(n9936), .A(n9935), .B(n9934), .ZN(n9938)
         );
  NAND2_X1 U5073 ( .A1(n5590), .A2(n5589), .ZN(n9153) );
  NAND2_X1 U5074 ( .A1(n5510), .A2(n5509), .ZN(n7947) );
  NAND2_X1 U5075 ( .A1(n5062), .A2(n5060), .ZN(n4745) );
  INV_X2 U5076 ( .A(n10159), .ZN(n9029) );
  INV_X1 U5077 ( .A(n10060), .ZN(n9306) );
  NAND2_X1 U5078 ( .A1(n8293), .A2(n8298), .ZN(n8459) );
  INV_X1 U5079 ( .A(n10024), .ZN(n7396) );
  NOR2_X1 U5080 ( .A1(n7257), .A2(n9992), .ZN(n7407) );
  AND3_X1 U5081 ( .A1(n5989), .A2(n5988), .A3(n5987), .ZN(n10024) );
  INV_X2 U5082 ( .A(n7074), .ZN(n8580) );
  INV_X2 U5083 ( .A(n9221), .ZN(n4510) );
  NAND2_X1 U5084 ( .A1(n5364), .A2(n5363), .ZN(n10165) );
  NAND4_X1 U5085 ( .A1(n5966), .A2(n5965), .A3(n5964), .A4(n5963), .ZN(n9421)
         );
  OAI21_X1 U5086 ( .B1(n5401), .B2(n5232), .A(n5231), .ZN(n5434) );
  AND2_X2 U5087 ( .A1(n6837), .A2(n4963), .ZN(n7074) );
  CLKBUF_X3 U5088 ( .A(n6620), .Z(n4512) );
  NAND4_X1 U5089 ( .A1(n5985), .A2(n5984), .A3(n5983), .A4(n5982), .ZN(n7416)
         );
  INV_X2 U5090 ( .A(n5319), .ZN(n5776) );
  BUF_X2 U5091 ( .A(n5319), .Z(n7532) );
  INV_X2 U5092 ( .A(n6697), .ZN(n6747) );
  NAND2_X1 U5093 ( .A1(n5157), .A2(n7700), .ZN(n5529) );
  NAND2_X1 U5094 ( .A1(n5819), .A2(n8260), .ZN(n10151) );
  OAI21_X1 U5095 ( .B1(n5356), .B2(n4700), .A(n4697), .ZN(n5393) );
  INV_X1 U5096 ( .A(n5511), .ZN(n5157) );
  INV_X1 U5097 ( .A(n9214), .ZN(n6339) );
  OR2_X1 U5098 ( .A1(n6313), .A2(n5937), .ZN(n5941) );
  NAND2_X1 U5099 ( .A1(n5341), .A2(n5225), .ZN(n5339) );
  INV_X2 U5100 ( .A(n5939), .ZN(n6872) );
  INV_X4 U5101 ( .A(n5961), .ZN(n6313) );
  INV_X2 U5102 ( .A(n5908), .ZN(n4673) );
  INV_X1 U5103 ( .A(n9168), .ZN(n5193) );
  INV_X2 U5104 ( .A(n5890), .ZN(n5900) );
  INV_X1 U5105 ( .A(n6434), .ZN(n7103) );
  NAND2_X1 U5106 ( .A1(n5771), .A2(n5772), .ZN(n5341) );
  AND2_X1 U5107 ( .A1(n7759), .A2(n7601), .ZN(n6434) );
  XNOR2_X1 U5108 ( .A(n5618), .B(n5617), .ZN(n8859) );
  XNOR2_X1 U5109 ( .A(n5870), .B(n5869), .ZN(n5874) );
  XNOR2_X1 U5110 ( .A(n6430), .B(n6429), .ZN(n7759) );
  NAND2_X1 U5111 ( .A1(n7601), .A2(n4509), .ZN(n5866) );
  AND2_X1 U5112 ( .A1(n5789), .A2(n4529), .ZN(n5803) );
  INV_X1 U5113 ( .A(n8456), .ZN(n7601) );
  NAND2_X1 U5114 ( .A1(n5859), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6430) );
  OR2_X1 U5115 ( .A1(n5871), .A2(n5848), .ZN(n5873) );
  NAND2_X1 U5116 ( .A1(n9896), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5870) );
  INV_X2 U5117 ( .A(n9166), .ZN(n9171) );
  XNOR2_X1 U5118 ( .A(n5860), .B(P1_IR_REG_21__SCAN_IN), .ZN(n8456) );
  INV_X1 U5119 ( .A(n5136), .ZN(n5847) );
  OAI21_X1 U5120 ( .B1(n5136), .B2(n4771), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n5844) );
  NAND2_X2 U5121 ( .A1(n5217), .A2(P2_U3151), .ZN(n8539) );
  NAND3_X1 U5122 ( .A1(n4814), .A2(n4815), .A3(n5135), .ZN(n5136) );
  XNOR2_X1 U5123 ( .A(n5340), .B(n5359), .ZN(n6947) );
  AND2_X1 U5124 ( .A1(n4521), .A2(n5834), .ZN(n4814) );
  AND2_X1 U5125 ( .A1(n5185), .A2(n4576), .ZN(n5082) );
  AND2_X2 U5126 ( .A1(n5832), .A2(n6155), .ZN(n5834) );
  AND2_X1 U5127 ( .A1(n5142), .A2(n10441), .ZN(n5135) );
  AND2_X1 U5128 ( .A1(n4542), .A2(n5000), .ZN(n4815) );
  AND2_X1 U5129 ( .A1(n5833), .A2(n5836), .ZN(n5000) );
  AND3_X1 U5130 ( .A1(n5831), .A2(n6201), .A3(n6158), .ZN(n5832) );
  INV_X4 U5131 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3151) );
  NOR2_X1 U5132 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(P1_IR_REG_2__SCAN_IN), .ZN(
        n5833) );
  INV_X4 U5133 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  NOR2_X2 U5134 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5906) );
  INV_X1 U5135 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n5484) );
  INV_X1 U5136 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n5390) );
  NOR2_X1 U5137 ( .A1(P2_IR_REG_3__SCAN_IN), .A2(P2_IR_REG_2__SCAN_IN), .ZN(
        n5179) );
  NOR2_X2 U5138 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n6944) );
  NOR2_X1 U5139 ( .A1(P2_IR_REG_4__SCAN_IN), .A2(P2_IR_REG_9__SCAN_IN), .ZN(
        n5174) );
  NOR2_X1 U5140 ( .A1(P2_IR_REG_13__SCAN_IN), .A2(P2_IR_REG_12__SCAN_IN), .ZN(
        n5173) );
  NOR2_X1 U5141 ( .A1(P2_IR_REG_6__SCAN_IN), .A2(P2_IR_REG_10__SCAN_IN), .ZN(
        n5172) );
  INV_X1 U5142 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n5489) );
  NOR2_X1 U5143 ( .A1(P1_IR_REG_11__SCAN_IN), .A2(P1_IR_REG_10__SCAN_IN), .ZN(
        n6155) );
  INV_X1 U5144 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n5862) );
  NOR2_X1 U5145 ( .A1(P1_IR_REG_16__SCAN_IN), .A2(P1_IR_REG_9__SCAN_IN), .ZN(
        n5830) );
  INV_X1 U5146 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n6432) );
  NOR2_X1 U5147 ( .A1(P1_IR_REG_4__SCAN_IN), .A2(P1_IR_REG_6__SCAN_IN), .ZN(
        n5828) );
  NOR2_X1 U5148 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(P1_IR_REG_7__SCAN_IN), .ZN(
        n5829) );
  NOR2_X1 U5149 ( .A1(P1_IR_REG_26__SCAN_IN), .A2(P1_IR_REG_25__SCAN_IN), .ZN(
        n5840) );
  INV_X1 U5150 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n6201) );
  OAI21_X2 U5151 ( .B1(n9663), .B2(n5025), .A(n5023), .ZN(n9632) );
  OAI21_X4 U5152 ( .B1(n9679), .B2(n6558), .A(n6557), .ZN(n9663) );
  AOI21_X2 U5153 ( .B1(n5518), .B2(n4548), .A(n5141), .ZN(n7900) );
  INV_X4 U5154 ( .A(n6768), .ZN(n4823) );
  NAND2_X1 U5155 ( .A1(n5925), .A2(n5865), .ZN(n6620) );
  NAND2_X2 U5156 ( .A1(n9276), .A2(n9277), .ZN(n9275) );
  NAND2_X1 U5157 ( .A1(n5874), .A2(n5875), .ZN(n5890) );
  OAI21_X2 U5158 ( .B1(n7306), .B2(n5398), .A(n5397), .ZN(n7457) );
  OAI21_X2 U5159 ( .B1(n7266), .B2(n5755), .A(n5756), .ZN(n7306) );
  OAI22_X2 U5160 ( .A1(n7500), .A2(n5433), .B1(n8740), .B2(n7507), .ZN(n7632)
         );
  NAND2_X2 U5161 ( .A1(n5414), .A2(n5413), .ZN(n7500) );
  OAI21_X2 U5162 ( .B1(n9711), .B2(n5029), .A(n5027), .ZN(n9679) );
  OAI21_X2 U5163 ( .B1(n9735), .B2(n6554), .A(n6553), .ZN(n9711) );
  INV_X1 U5164 ( .A(n5908), .ZN(n4514) );
  NAND2_X1 U5165 ( .A1(n4705), .A2(n4701), .ZN(n8166) );
  INV_X1 U5166 ( .A(n8162), .ZN(n4705) );
  NAND2_X1 U5167 ( .A1(n4703), .A2(n4702), .ZN(n4701) );
  NOR2_X1 U5168 ( .A1(n4912), .A2(n5566), .ZN(n4911) );
  NOR2_X1 U5169 ( .A1(n4516), .A2(n5550), .ZN(n4912) );
  NAND2_X1 U5170 ( .A1(n4867), .A2(n4534), .ZN(n4862) );
  INV_X1 U5171 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n5309) );
  INV_X1 U5172 ( .A(n5874), .ZN(n5876) );
  INV_X1 U5173 ( .A(n6027), .ZN(n6577) );
  XNOR2_X1 U5174 ( .A(n10165), .B(n7074), .ZN(n7114) );
  AND2_X1 U5175 ( .A1(n8331), .A2(n8330), .ZN(n9543) );
  INV_X1 U5176 ( .A(n6154), .ZN(n6501) );
  XNOR2_X1 U5177 ( .A(n6480), .B(SI_29_), .ZN(n9170) );
  INV_X1 U5178 ( .A(n8379), .ZN(n8386) );
  INV_X1 U5179 ( .A(n8420), .ZN(n4821) );
  NAND2_X1 U5180 ( .A1(n8146), .A2(n4719), .ZN(n8140) );
  AND2_X1 U5181 ( .A1(n8150), .A2(n8245), .ZN(n4719) );
  NAND2_X1 U5182 ( .A1(n4819), .A2(n4818), .ZN(n4817) );
  INV_X1 U5183 ( .A(n8426), .ZN(n4818) );
  NAND2_X1 U5184 ( .A1(n4820), .A2(n9655), .ZN(n4819) );
  AOI21_X1 U5185 ( .B1(n4834), .B2(n4831), .A(n4654), .ZN(n4653) );
  AND2_X1 U5186 ( .A1(n8433), .A2(n4832), .ZN(n4831) );
  NAND2_X1 U5187 ( .A1(n4835), .A2(n8440), .ZN(n4654) );
  OAI21_X1 U5188 ( .B1(n8436), .B2(n8431), .A(n8438), .ZN(n4834) );
  INV_X1 U5189 ( .A(n5039), .ZN(n5037) );
  INV_X1 U5190 ( .A(n4716), .ZN(n4715) );
  AOI21_X1 U5191 ( .B1(n8170), .B2(n8203), .A(n8178), .ZN(n4716) );
  NOR2_X1 U5192 ( .A1(n4956), .A2(n5383), .ZN(n4951) );
  NAND2_X1 U5193 ( .A1(n5522), .A2(n5064), .ZN(n5062) );
  AND2_X1 U5194 ( .A1(n5248), .A2(n5065), .ZN(n5064) );
  NAND2_X1 U5195 ( .A1(n5536), .A2(SI_14_), .ZN(n5065) );
  NAND2_X1 U5196 ( .A1(n8674), .A2(n4549), .ZN(n4968) );
  NOR2_X1 U5197 ( .A1(n9081), .A2(n5095), .ZN(n5094) );
  NOR2_X1 U5198 ( .A1(n9084), .A2(n8882), .ZN(n5095) );
  NOR2_X1 U5199 ( .A1(n5093), .A2(n8215), .ZN(n5091) );
  INV_X1 U5200 ( .A(n9081), .ZN(n5093) );
  NOR2_X1 U5201 ( .A1(n4533), .A2(n7061), .ZN(n4865) );
  OR2_X1 U5202 ( .A1(n6937), .A2(n4533), .ZN(n4860) );
  INV_X1 U5203 ( .A(n4868), .ZN(n4867) );
  OR2_X1 U5204 ( .A1(n7172), .A2(n4854), .ZN(n4853) );
  INV_X1 U5205 ( .A(n7148), .ZN(n4854) );
  AND2_X1 U5206 ( .A1(n4567), .A2(n4888), .ZN(n4518) );
  NAND2_X1 U5207 ( .A1(n4889), .A2(n4890), .ZN(n4888) );
  AND2_X1 U5208 ( .A1(n9095), .A2(n8914), .ZN(n4890) );
  OR2_X1 U5209 ( .A1(n8628), .A2(n8667), .ZN(n8175) );
  OR2_X1 U5210 ( .A1(n8699), .A2(n8994), .ZN(n8245) );
  AOI21_X1 U5211 ( .B1(n4911), .B2(n4516), .A(n4559), .ZN(n4910) );
  OR2_X1 U5212 ( .A1(n8647), .A2(n8653), .ZN(n8144) );
  OR2_X1 U5213 ( .A1(n7953), .A2(n7985), .ZN(n8055) );
  NAND2_X1 U5214 ( .A1(n9158), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5308) );
  INV_X1 U5215 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n5085) );
  AND2_X1 U5216 ( .A1(n9526), .A2(n8493), .ZN(n8484) );
  AOI21_X1 U5217 ( .B1(n8452), .B2(n8451), .A(n4647), .ZN(n4841) );
  NAND2_X1 U5218 ( .A1(n4649), .A2(n4648), .ZN(n4647) );
  INV_X1 U5219 ( .A(n4842), .ZN(n4649) );
  OAI21_X1 U5220 ( .B1(n8451), .B2(n8444), .A(n8445), .ZN(n4842) );
  INV_X1 U5221 ( .A(n8484), .ZN(n8510) );
  INV_X1 U5222 ( .A(n4772), .ZN(n4631) );
  AOI21_X1 U5223 ( .B1(n4772), .B2(n4630), .A(n4629), .ZN(n4628) );
  INV_X1 U5224 ( .A(n8430), .ZN(n4629) );
  INV_X1 U5225 ( .A(n4773), .ZN(n4630) );
  INV_X1 U5226 ( .A(n8431), .ZN(n8435) );
  NAND2_X1 U5227 ( .A1(n4750), .A2(n4748), .ZN(n9600) );
  AND2_X1 U5228 ( .A1(n4749), .A2(n6363), .ZN(n4748) );
  OR2_X1 U5229 ( .A1(n9688), .A2(n9232), .ZN(n8335) );
  OR2_X1 U5230 ( .A1(n6548), .A2(n5011), .ZN(n5010) );
  INV_X1 U5231 ( .A(n6547), .ZN(n5011) );
  NOR2_X1 U5232 ( .A1(n7842), .A2(n7765), .ZN(n4763) );
  OAI21_X1 U5233 ( .B1(n6480), .B2(n10358), .A(n6479), .ZN(n6498) );
  NAND2_X1 U5234 ( .A1(n5294), .A2(n5293), .ZN(n5705) );
  AND2_X1 U5235 ( .A1(n5289), .A2(n5288), .ZN(n5678) );
  NAND2_X1 U5236 ( .A1(n5244), .A2(SI_13_), .ZN(n5248) );
  NAND2_X1 U5237 ( .A1(n5520), .A2(n5519), .ZN(n5522) );
  OR2_X1 U5238 ( .A1(n6018), .A2(P1_IR_REG_5__SCAN_IN), .ZN(n6070) );
  AND2_X1 U5239 ( .A1(n8205), .A2(n6668), .ZN(n4964) );
  AND2_X1 U5240 ( .A1(n7117), .A2(n7115), .ZN(n4966) );
  INV_X1 U5241 ( .A(n7120), .ZN(n7117) );
  AOI21_X1 U5242 ( .B1(n4983), .B2(n4979), .A(n4540), .ZN(n4978) );
  INV_X1 U5243 ( .A(n7728), .ZN(n4979) );
  INV_X1 U5244 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n5743) );
  OR2_X1 U5246 ( .A1(n4926), .A2(n7239), .ZN(n6993) );
  NAND2_X1 U5247 ( .A1(n7056), .A2(n4932), .ZN(n7058) );
  NAND2_X1 U5248 ( .A1(n4929), .A2(n4928), .ZN(n4932) );
  NAND2_X1 U5249 ( .A1(n4927), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n4928) );
  NAND2_X1 U5250 ( .A1(n6964), .A2(n4930), .ZN(n4929) );
  AND2_X1 U5251 ( .A1(n7156), .A2(n7148), .ZN(n4855) );
  NOR2_X1 U5252 ( .A1(n7578), .A2(n7795), .ZN(n7693) );
  OR2_X1 U5253 ( .A1(n4944), .A2(n4946), .ZN(n4940) );
  NAND2_X1 U5254 ( .A1(n4944), .A2(n4942), .ZN(n4941) );
  NAND2_X1 U5255 ( .A1(n8823), .A2(n8862), .ZN(n4942) );
  NAND2_X1 U5256 ( .A1(n5168), .A2(n5167), .ZN(n5708) );
  INV_X1 U5257 ( .A(n5696), .ZN(n5168) );
  OR2_X1 U5258 ( .A1(n8737), .A2(n7777), .ZN(n4598) );
  AOI21_X1 U5260 ( .B1(n4919), .B2(n4918), .A(n4556), .ZN(n4917) );
  INV_X1 U5261 ( .A(n4922), .ZN(n4918) );
  INV_X1 U5262 ( .A(n10151), .ZN(n9003) );
  OR2_X1 U5263 ( .A1(n9067), .A2(n9007), .ZN(n8150) );
  INV_X1 U5264 ( .A(n4507), .ZN(n5619) );
  OAI21_X1 U5265 ( .B1(n5792), .B2(n4915), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n4914) );
  NAND2_X1 U5266 ( .A1(n4569), .A2(n4527), .ZN(n4915) );
  NAND2_X1 U5267 ( .A1(n6219), .A2(n6222), .ZN(n4811) );
  INV_X1 U5268 ( .A(n9176), .ZN(n6222) );
  AOI21_X1 U5269 ( .B1(n4801), .B2(n4803), .A(n4799), .ZN(n4798) );
  NAND2_X1 U5270 ( .A1(n9336), .A2(n4801), .ZN(n4800) );
  INV_X1 U5271 ( .A(n9286), .ZN(n4799) );
  AND2_X1 U5272 ( .A1(n6410), .A2(n5124), .ZN(n5123) );
  NAND2_X1 U5273 ( .A1(n9254), .A2(n5125), .ZN(n5124) );
  INV_X1 U5274 ( .A(n6376), .ZN(n5125) );
  AOI21_X1 U5275 ( .B1(n8507), .B2(n8455), .A(n8454), .ZN(n8503) );
  INV_X1 U5276 ( .A(n5866), .ZN(n8454) );
  AND4_X1 U5277 ( .A1(n6211), .A2(n6210), .A3(n6209), .A4(n6208), .ZN(n7927)
         );
  OR2_X1 U5278 ( .A1(n6571), .A2(n6570), .ZN(n9548) );
  OR2_X1 U5279 ( .A1(n9770), .A2(n7235), .ZN(n5015) );
  NAND2_X1 U5280 ( .A1(n5018), .A2(n5017), .ZN(n6568) );
  AND2_X1 U5281 ( .A1(n5019), .A2(n4586), .ZN(n5017) );
  AOI21_X1 U5282 ( .B1(n5026), .B2(n5024), .A(n4584), .ZN(n5023) );
  INV_X1 U5283 ( .A(n5026), .ZN(n5025) );
  NAND2_X1 U5284 ( .A1(n7812), .A2(n8468), .ZN(n6546) );
  OR2_X1 U5285 ( .A1(n9831), .A2(n8509), .ZN(n6510) );
  OR2_X1 U5286 ( .A1(n6498), .A2(n6497), .ZN(n6500) );
  NAND2_X1 U5287 ( .A1(n5038), .A2(n5039), .ZN(n5642) );
  NAND2_X1 U5288 ( .A1(n5630), .A2(n5040), .ZN(n5038) );
  AND2_X1 U5289 ( .A1(n5239), .A2(n5236), .ZN(n5059) );
  INV_X1 U5290 ( .A(n5781), .ZN(n6655) );
  NAND2_X1 U5291 ( .A1(n5721), .A2(n5720), .ZN(n8590) );
  INV_X1 U5292 ( .A(n5772), .ZN(n8266) );
  AOI21_X1 U5293 ( .B1(n9540), .B2(n9837), .A(n9539), .ZN(n9763) );
  OR2_X1 U5294 ( .A1(n9893), .A2(n6510), .ZN(n9970) );
  AOI21_X1 U5295 ( .B1(n9170), .B2(n6501), .A(n5144), .ZN(n9852) );
  INV_X1 U5296 ( .A(n4845), .ZN(n4844) );
  OAI21_X1 U5297 ( .B1(n8348), .B2(n8453), .A(n8349), .ZN(n4845) );
  AND2_X1 U5298 ( .A1(n8370), .A2(n8369), .ZN(n4662) );
  INV_X1 U5299 ( .A(n4661), .ZN(n4660) );
  NAND2_X1 U5300 ( .A1(n4720), .A2(n8137), .ZN(n8146) );
  NAND2_X1 U5301 ( .A1(n4722), .A2(n4721), .ZN(n4720) );
  OAI21_X1 U5302 ( .B1(n4704), .B2(n8154), .A(n8161), .ZN(n4703) );
  NOR2_X1 U5303 ( .A1(n8156), .A2(n8155), .ZN(n4704) );
  OAI21_X1 U5304 ( .B1(n8166), .B2(n8163), .A(n8219), .ZN(n8165) );
  NOR2_X1 U5305 ( .A1(n8439), .A2(n8453), .ZN(n4837) );
  AOI21_X1 U5306 ( .B1(n8436), .B2(n8435), .A(n4839), .ZN(n4838) );
  INV_X1 U5307 ( .A(n8438), .ZN(n4839) );
  INV_X1 U5308 ( .A(n5718), .ZN(n5058) );
  INV_X1 U5309 ( .A(n5057), .ZN(n5056) );
  OAI21_X1 U5310 ( .B1(n5305), .B2(n5058), .A(n5730), .ZN(n5057) );
  INV_X1 U5311 ( .A(n5640), .ZN(n5271) );
  AND2_X1 U5312 ( .A1(n6381), .A2(n6380), .ZN(n6395) );
  NOR2_X1 U5313 ( .A1(n6349), .A2(n9189), .ZN(n6381) );
  NOR2_X1 U5314 ( .A1(n5536), .A2(SI_14_), .ZN(n5063) );
  INV_X1 U5315 ( .A(n4787), .ZN(n4785) );
  NAND2_X1 U5316 ( .A1(n4634), .A2(SI_7_), .ZN(n5228) );
  INV_X1 U5317 ( .A(n8701), .ZN(n4987) );
  AOI21_X1 U5318 ( .B1(n4992), .B2(n4990), .A(n8702), .ZN(n4989) );
  INV_X1 U5319 ( .A(n8546), .ZN(n4990) );
  AOI21_X1 U5320 ( .B1(n4713), .B2(n8183), .A(n4711), .ZN(n8194) );
  NAND2_X1 U5321 ( .A1(n4712), .A2(n8184), .ZN(n4711) );
  OAI21_X1 U5322 ( .B1(n4717), .B2(n4715), .A(n4714), .ZN(n4713) );
  NOR2_X1 U5323 ( .A1(n5091), .A2(n5090), .ZN(n5089) );
  INV_X1 U5324 ( .A(n8212), .ZN(n5090) );
  OR2_X1 U5325 ( .A1(n4539), .A2(n6976), .ZN(n4927) );
  OAI21_X1 U5326 ( .B1(n7060), .B2(n4952), .A(n4948), .ZN(n7126) );
  NOR2_X1 U5327 ( .A1(n4951), .A2(n4949), .ZN(n4948) );
  NOR2_X1 U5328 ( .A1(n6949), .A2(n4950), .ZN(n4949) );
  AND3_X1 U5329 ( .A1(n4871), .A2(n4872), .A3(n4590), .ZN(n8761) );
  OAI21_X1 U5330 ( .B1(n8184), .B2(n4561), .A(n4886), .ZN(n4885) );
  NAND2_X1 U5331 ( .A1(n8184), .A2(n4518), .ZN(n4886) );
  INV_X1 U5332 ( .A(n8106), .ZN(n5759) );
  INV_X1 U5333 ( .A(n8176), .ZN(n4691) );
  NOR2_X1 U5334 ( .A1(n5691), .A2(n4923), .ZN(n4922) );
  INV_X1 U5335 ( .A(n5676), .ZN(n4923) );
  OR2_X1 U5336 ( .A1(n9119), .A2(n8694), .ZN(n8219) );
  OR2_X1 U5337 ( .A1(n9125), .A2(n8684), .ZN(n8046) );
  AOI21_X1 U5338 ( .B1(n4897), .B2(n8989), .A(n4895), .ZN(n4894) );
  INV_X1 U5339 ( .A(n8969), .ZN(n4895) );
  OR2_X1 U5340 ( .A1(n9131), .A2(n8678), .ZN(n8049) );
  AND2_X1 U5341 ( .A1(n5639), .A2(n4546), .ZN(n4897) );
  NAND2_X1 U5342 ( .A1(n7969), .A2(n4911), .ZN(n4909) );
  OR2_X1 U5343 ( .A1(n7970), .A2(n8129), .ZN(n8133) );
  NAND2_X1 U5344 ( .A1(n4683), .A2(n8232), .ZN(n4682) );
  AND2_X1 U5345 ( .A1(n5185), .A2(n5181), .ZN(n5086) );
  NOR2_X1 U5346 ( .A1(n5423), .A2(P2_IR_REG_6__SCAN_IN), .ZN(n5486) );
  OR2_X1 U5347 ( .A1(n5399), .A2(P2_IR_REG_5__SCAN_IN), .ZN(n5423) );
  NAND2_X1 U5348 ( .A1(n4514), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n4672) );
  NAND2_X1 U5349 ( .A1(n4823), .A2(n9425), .ZN(n4822) );
  NAND2_X1 U5350 ( .A1(n9933), .A2(n8445), .ZN(n8494) );
  AOI21_X1 U5351 ( .B1(n7887), .B2(P1_REG2_REG_14__SCAN_IN), .A(n7886), .ZN(
        n7888) );
  INV_X1 U5352 ( .A(n8442), .ZN(n8330) );
  INV_X1 U5353 ( .A(n8441), .ZN(n8331) );
  NOR2_X1 U5354 ( .A1(n6566), .A2(n5022), .ZN(n5021) );
  INV_X1 U5355 ( .A(n6565), .ZN(n5022) );
  AND2_X1 U5356 ( .A1(n9617), .A2(n9618), .ZN(n4773) );
  AOI21_X1 U5357 ( .B1(n6560), .B2(n6559), .A(n4557), .ZN(n5026) );
  NOR2_X1 U5358 ( .A1(n9719), .A2(n9739), .ZN(n4768) );
  NAND2_X1 U5359 ( .A1(n9835), .A2(n9834), .ZN(n6602) );
  NAND2_X1 U5360 ( .A1(n7873), .A2(n9177), .ZN(n8379) );
  INV_X1 U5361 ( .A(n5005), .ZN(n5004) );
  OAI21_X1 U5362 ( .B1(n9962), .B2(n5006), .A(n7663), .ZN(n5005) );
  INV_X1 U5363 ( .A(n6537), .ZN(n5006) );
  AND2_X1 U5364 ( .A1(n7665), .A2(n6593), .ZN(n8349) );
  INV_X1 U5365 ( .A(n8293), .ZN(n4658) );
  NAND2_X1 U5366 ( .A1(n4619), .A2(n4617), .ZN(n9636) );
  AOI21_X1 U5367 ( .B1(n4532), .B2(n4622), .A(n4618), .ZN(n4617) );
  NAND2_X1 U5368 ( .A1(n9680), .A2(n4532), .ZN(n4619) );
  INV_X1 U5369 ( .A(n8281), .ZN(n4618) );
  AND2_X1 U5370 ( .A1(n6417), .A2(n6715), .ZN(n7100) );
  AND2_X1 U5371 ( .A1(n6514), .A2(n6513), .ZN(n7101) );
  AOI21_X1 U5372 ( .B1(n5051), .B2(n5053), .A(n5050), .ZN(n5049) );
  INV_X1 U5373 ( .A(n5289), .ZN(n5050) );
  INV_X1 U5374 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n5838) );
  NAND2_X1 U5375 ( .A1(n4754), .A2(n4752), .ZN(n5651) );
  AOI21_X1 U5376 ( .B1(n4755), .B2(n4760), .A(n4753), .ZN(n4752) );
  INV_X1 U5377 ( .A(n5034), .ZN(n4753) );
  NAND2_X1 U5378 ( .A1(n4756), .A2(n4757), .ZN(n5630) );
  OR2_X1 U5379 ( .A1(n5586), .A2(n4760), .ZN(n4756) );
  NOR2_X1 U5380 ( .A1(n5264), .A2(n5047), .ZN(n5046) );
  INV_X1 U5381 ( .A(n5260), .ZN(n5047) );
  OAI21_X1 U5382 ( .B1(n5264), .B2(n5045), .A(n5263), .ZN(n5044) );
  NAND2_X1 U5383 ( .A1(n5585), .A2(n5260), .ZN(n5045) );
  NAND2_X1 U5384 ( .A1(n5252), .A2(n5251), .ZN(n5569) );
  NAND2_X1 U5385 ( .A1(n4745), .A2(n5061), .ZN(n5251) );
  NOR2_X1 U5386 ( .A1(n5479), .A2(n4788), .ZN(n4787) );
  INV_X1 U5387 ( .A(n5240), .ZN(n4788) );
  NAND2_X1 U5388 ( .A1(n5238), .A2(SI_10_), .ZN(n5240) );
  OAI22_X1 U5389 ( .A1(n5434), .A2(n5435), .B1(SI_8_), .B2(n5233), .ZN(n5452)
         );
  OAI21_X1 U5390 ( .B1(SI_7_), .B2(n4634), .A(n5228), .ZN(n5417) );
  OAI22_X1 U5391 ( .A1(n5393), .A2(n5224), .B1(SI_5_), .B2(n5223), .ZN(n5401)
         );
  INV_X1 U5392 ( .A(n5216), .ZN(n4699) );
  INV_X1 U5393 ( .A(P1_RD_REG_SCAN_IN), .ZN(n4696) );
  NOR2_X1 U5394 ( .A1(n8651), .A2(n4993), .ZN(n4992) );
  INV_X1 U5395 ( .A(n5139), .ZN(n4993) );
  INV_X1 U5396 ( .A(n8563), .ZN(n8565) );
  NAND2_X1 U5397 ( .A1(n4968), .A2(n4553), .ZN(n8686) );
  OR2_X1 U5398 ( .A1(n8685), .A2(n8971), .ZN(n4973) );
  INV_X1 U5399 ( .A(n4978), .ZN(n4976) );
  INV_X1 U5400 ( .A(n7850), .ZN(n4984) );
  AND2_X2 U5401 ( .A1(n8268), .A2(n6834), .ZN(n8203) );
  AND2_X1 U5402 ( .A1(n5584), .A2(n5583), .ZN(n8653) );
  NAND2_X1 U5403 ( .A1(n4936), .A2(n4934), .ZN(n7056) );
  OR2_X1 U5404 ( .A1(n6964), .A2(n4539), .ZN(n4936) );
  NAND2_X1 U5405 ( .A1(n6936), .A2(n6976), .ZN(n7062) );
  OR2_X1 U5406 ( .A1(n6981), .A2(n5347), .ZN(n7064) );
  AND2_X1 U5407 ( .A1(n4860), .A2(n4596), .ZN(n4858) );
  NAND2_X1 U5408 ( .A1(n7126), .A2(n7163), .ZN(n7168) );
  OAI21_X1 U5409 ( .B1(n7145), .B2(n4854), .A(n4530), .ZN(n7209) );
  INV_X1 U5410 ( .A(n4855), .ZN(n4852) );
  AOI21_X1 U5411 ( .B1(n4530), .B2(n4854), .A(n4848), .ZN(n4847) );
  OR2_X1 U5412 ( .A1(n7335), .A2(n7339), .ZN(n4879) );
  NOR2_X1 U5413 ( .A1(n7693), .A2(n7694), .ZN(n7697) );
  INV_X1 U5414 ( .A(n4635), .ZN(n7691) );
  OR2_X1 U5415 ( .A1(n7697), .A2(n7696), .ZN(n4960) );
  OR2_X1 U5416 ( .A1(n7569), .A2(n4874), .ZN(n4871) );
  OR2_X1 U5417 ( .A1(n7683), .A2(n5497), .ZN(n4874) );
  NAND2_X1 U5418 ( .A1(n7682), .A2(n4873), .ZN(n4872) );
  INV_X1 U5419 ( .A(n7683), .ZN(n4873) );
  NOR2_X1 U5420 ( .A1(n10125), .A2(n10124), .ZN(n10123) );
  NAND2_X1 U5421 ( .A1(n4645), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n4644) );
  NOR2_X1 U5422 ( .A1(n10119), .A2(n4958), .ZN(n8788) );
  NOR2_X1 U5423 ( .A1(n8764), .A2(n8747), .ZN(n4958) );
  XNOR2_X1 U5424 ( .A(n4869), .B(n8765), .ZN(n8766) );
  OR2_X1 U5425 ( .A1(n10123), .A2(n4870), .ZN(n4869) );
  NOR2_X1 U5426 ( .A1(n8764), .A2(n8763), .ZN(n4870) );
  NOR2_X1 U5427 ( .A1(n8766), .A2(n8767), .ZN(n8775) );
  NOR2_X1 U5428 ( .A1(n8801), .A2(n4880), .ZN(n8842) );
  AND2_X1 U5429 ( .A1(n8810), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n4880) );
  OR2_X1 U5430 ( .A1(n8803), .A2(n9077), .ZN(n8846) );
  AOI21_X1 U5431 ( .B1(n8821), .B2(n4945), .A(n8858), .ZN(n4944) );
  NOR2_X1 U5432 ( .A1(n8808), .A2(n8807), .ZN(n8820) );
  NAND2_X1 U5433 ( .A1(n5164), .A2(n5163), .ZN(n5668) );
  INV_X1 U5434 ( .A(n5645), .ZN(n5164) );
  OR2_X1 U5435 ( .A1(n5633), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n5645) );
  NAND2_X1 U5436 ( .A1(n9019), .A2(n4721), .ZN(n5081) );
  AND2_X1 U5437 ( .A1(n5594), .A2(n5593), .ZN(n9005) );
  OR2_X1 U5438 ( .A1(n5578), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n5591) );
  AND2_X1 U5439 ( .A1(n5759), .A2(n8115), .ZN(n4683) );
  OR2_X1 U5440 ( .A1(n7645), .A2(n7730), .ZN(n8115) );
  OR2_X1 U5441 ( .A1(n7618), .A2(n8232), .ZN(n4684) );
  INV_X1 U5442 ( .A(n4901), .ZN(n4900) );
  OAI21_X1 U5443 ( .B1(n7456), .B2(n5099), .A(n5096), .ZN(n7618) );
  INV_X1 U5444 ( .A(n5100), .ZN(n5099) );
  AOI21_X1 U5445 ( .B1(n5100), .B2(n5098), .A(n5097), .ZN(n5096) );
  AND2_X1 U5446 ( .A1(n4693), .A2(n4692), .ZN(n5100) );
  NAND2_X1 U5447 ( .A1(n4903), .A2(n5449), .ZN(n7634) );
  NOR2_X1 U5448 ( .A1(n8090), .A2(n8096), .ZN(n5105) );
  OR2_X1 U5449 ( .A1(n8096), .A2(n5104), .ZN(n4693) );
  NAND2_X1 U5450 ( .A1(n8081), .A2(n8091), .ZN(n5104) );
  OR2_X1 U5451 ( .A1(n5406), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5428) );
  NAND2_X1 U5452 ( .A1(n5150), .A2(n7282), .ZN(n5380) );
  INV_X1 U5453 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n5150) );
  NAND2_X1 U5454 ( .A1(n5757), .A2(n5756), .ZN(n8220) );
  NOR2_X1 U5455 ( .A1(n8897), .A2(n8172), .ZN(n5074) );
  NAND2_X1 U5456 ( .A1(n4687), .A2(n4685), .ZN(n5075) );
  NOR2_X1 U5457 ( .A1(n4686), .A2(n8173), .ZN(n4685) );
  INV_X1 U5458 ( .A(n4688), .ZN(n4686) );
  OR2_X1 U5459 ( .A1(n8173), .A2(n8172), .ZN(n8912) );
  NOR2_X1 U5460 ( .A1(n4690), .A2(n4689), .ZN(n4688) );
  INV_X1 U5461 ( .A(n8175), .ZN(n4689) );
  NOR2_X1 U5462 ( .A1(n8218), .A2(n4691), .ZN(n4690) );
  OR2_X1 U5463 ( .A1(n5765), .A2(n4691), .ZN(n4687) );
  INV_X1 U5464 ( .A(n8945), .ZN(n8925) );
  NAND2_X1 U5465 ( .A1(n5677), .A2(n4922), .ZN(n4921) );
  NAND2_X1 U5466 ( .A1(n6842), .A2(n8203), .ZN(n9008) );
  OR2_X1 U5467 ( .A1(n9113), .A2(n8925), .ZN(n8218) );
  NAND2_X1 U5468 ( .A1(n8992), .A2(n8991), .ZN(n4898) );
  NAND2_X1 U5469 ( .A1(n4898), .A2(n4897), .ZN(n8967) );
  AND2_X1 U5470 ( .A1(n5762), .A2(n8965), .ZN(n8979) );
  AOI21_X1 U5471 ( .B1(n9018), .B2(n5079), .A(n5077), .ZN(n5076) );
  INV_X1 U5472 ( .A(n5079), .ZN(n5078) );
  INV_X1 U5473 ( .A(n8245), .ZN(n5077) );
  AOI21_X1 U5474 ( .B1(n4907), .B2(n4906), .A(n4905), .ZN(n4904) );
  INV_X1 U5475 ( .A(n9020), .ZN(n4905) );
  NAND2_X1 U5476 ( .A1(n4909), .A2(n4910), .ZN(n8025) );
  NAND2_X1 U5477 ( .A1(n4909), .A2(n4907), .ZN(n9021) );
  NAND2_X1 U5478 ( .A1(n4679), .A2(n8057), .ZN(n4675) );
  NOR2_X1 U5479 ( .A1(n5110), .A2(n5109), .ZN(n5108) );
  AND2_X1 U5480 ( .A1(n8144), .A2(n8141), .ZN(n8242) );
  NAND2_X1 U5481 ( .A1(n4526), .A2(n5116), .ZN(n5113) );
  NAND2_X1 U5482 ( .A1(n5761), .A2(n8054), .ZN(n5115) );
  NOR2_X1 U5483 ( .A1(n8129), .A2(n5112), .ZN(n5111) );
  INV_X1 U5484 ( .A(n8054), .ZN(n5112) );
  AND2_X1 U5485 ( .A1(n8135), .A2(n8143), .ZN(n8240) );
  NAND2_X1 U5486 ( .A1(n4676), .A2(n8057), .ZN(n7905) );
  NAND2_X1 U5487 ( .A1(n7856), .A2(n8235), .ZN(n4676) );
  INV_X1 U5488 ( .A(n9008), .ZN(n10148) );
  AND2_X1 U5489 ( .A1(n5405), .A2(n5404), .ZN(n10177) );
  XNOR2_X1 U5490 ( .A(n5803), .B(n5790), .ZN(n5794) );
  INV_X1 U5491 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n4916) );
  AND2_X1 U5492 ( .A1(n5085), .A2(n5186), .ZN(n5083) );
  AND2_X1 U5493 ( .A1(n5572), .A2(n4573), .ZN(n5748) );
  INV_X1 U5494 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n4995) );
  INV_X1 U5495 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n5359) );
  INV_X1 U5496 ( .A(n5133), .ZN(n5132) );
  OR2_X1 U5497 ( .A1(n6141), .A2(n6140), .ZN(n6167) );
  INV_X1 U5498 ( .A(n5931), .ZN(n5926) );
  NOR2_X1 U5499 ( .A1(n4809), .A2(n6128), .ZN(n4808) );
  INV_X1 U5500 ( .A(n6113), .ZN(n4809) );
  XNOR2_X1 U5501 ( .A(n5953), .B(n9210), .ZN(n5958) );
  NOR2_X1 U5502 ( .A1(n6442), .A2(n8498), .ZN(n9199) );
  NAND2_X1 U5503 ( .A1(n6442), .A2(n6766), .ZN(n9338) );
  NAND2_X1 U5504 ( .A1(n6247), .A2(n6246), .ZN(n9388) );
  NAND2_X1 U5505 ( .A1(n8506), .A2(n7528), .ZN(n4744) );
  NAND2_X1 U5506 ( .A1(n8329), .A2(n8328), .ZN(n4743) );
  INV_X1 U5507 ( .A(n8508), .ZN(n4751) );
  INV_X1 U5508 ( .A(n4841), .ZN(n4840) );
  AND2_X1 U5509 ( .A1(n6402), .A2(n6401), .ZN(n9257) );
  AND2_X1 U5510 ( .A1(n6355), .A2(n6354), .ZN(n9339) );
  AND2_X1 U5511 ( .A1(n5882), .A2(n5881), .ZN(n9233) );
  AND3_X1 U5512 ( .A1(n5893), .A2(n5892), .A3(n5891), .ZN(n9232) );
  AND4_X1 U5513 ( .A1(n6284), .A2(n6283), .A3(n6282), .A4(n6281), .ZN(n9367)
         );
  AND4_X1 U5514 ( .A1(n6263), .A2(n6262), .A3(n6261), .A4(n6260), .ZN(n9279)
         );
  AND4_X1 U5515 ( .A1(n6124), .A2(n6123), .A3(n6122), .A4(n6121), .ZN(n7740)
         );
  AND4_X1 U5516 ( .A1(n6104), .A2(n6103), .A3(n6102), .A4(n6101), .ZN(n7669)
         );
  AND4_X1 U5517 ( .A1(n6086), .A2(n6085), .A3(n6084), .A4(n6083), .ZN(n7717)
         );
  AND4_X1 U5518 ( .A1(n6051), .A2(n6050), .A3(n6049), .A4(n6048), .ZN(n7668)
         );
  NAND2_X1 U5519 ( .A1(n9469), .A2(n4736), .ZN(n4735) );
  NAND2_X1 U5520 ( .A1(n9464), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n4736) );
  NAND2_X1 U5521 ( .A1(n4735), .A2(n4734), .ZN(n4733) );
  INV_X1 U5522 ( .A(n6808), .ZN(n4734) );
  AND2_X1 U5523 ( .A1(n5833), .A2(n5906), .ZN(n6008) );
  INV_X1 U5524 ( .A(n9933), .ZN(n8451) );
  AOI21_X1 U5525 ( .B1(n9555), .B2(n6577), .A(n6576), .ZN(n9538) );
  AOI21_X1 U5526 ( .B1(n5021), .B2(n6564), .A(n5020), .ZN(n5019) );
  NOR2_X1 U5527 ( .A1(n9609), .A2(n9401), .ZN(n5020) );
  AND2_X1 U5528 ( .A1(n6603), .A2(n9600), .ZN(n4772) );
  NAND2_X1 U5529 ( .A1(n9635), .A2(n4773), .ZN(n9619) );
  NAND2_X1 U5530 ( .A1(n9636), .A2(n9637), .ZN(n9635) );
  NOR2_X1 U5531 ( .A1(n9662), .A2(n4624), .ZN(n4623) );
  INV_X1 U5532 ( .A(n8335), .ZN(n4624) );
  NAND2_X1 U5533 ( .A1(n9680), .A2(n8335), .ZN(n9665) );
  AOI21_X1 U5534 ( .B1(n5030), .B2(n5028), .A(n4543), .ZN(n5027) );
  INV_X1 U5535 ( .A(n5030), .ZN(n5029) );
  INV_X1 U5536 ( .A(n6556), .ZN(n5028) );
  NAND2_X1 U5537 ( .A1(n9705), .A2(n8334), .ZN(n9682) );
  INV_X1 U5538 ( .A(n8478), .ZN(n9681) );
  NAND2_X1 U5539 ( .A1(n9730), .A2(n8408), .ZN(n9713) );
  AND2_X1 U5540 ( .A1(n8408), .A2(n8289), .ZN(n9734) );
  INV_X1 U5541 ( .A(n9734), .ZN(n9728) );
  OAI21_X1 U5542 ( .B1(n7920), .B2(n6549), .A(n6550), .ZN(n9829) );
  OAI21_X1 U5543 ( .B1(n7820), .B2(n8383), .A(n4562), .ZN(n7924) );
  NAND2_X1 U5544 ( .A1(n4776), .A2(n8380), .ZN(n4774) );
  AND2_X1 U5545 ( .A1(n8381), .A2(n8380), .ZN(n9752) );
  OR2_X1 U5546 ( .A1(n7873), .A2(n9177), .ZN(n8385) );
  NAND2_X1 U5547 ( .A1(n7820), .A2(n4775), .ZN(n9748) );
  INV_X1 U5548 ( .A(n4776), .ZN(n4775) );
  NAND2_X1 U5549 ( .A1(n8385), .A2(n8379), .ZN(n7822) );
  OR2_X1 U5550 ( .A1(n7823), .A2(n7822), .ZN(n7820) );
  INV_X1 U5551 ( .A(n8471), .ZN(n7751) );
  OR2_X1 U5552 ( .A1(n9419), .A2(n10039), .ZN(n9963) );
  INV_X1 U5553 ( .A(n8349), .ZN(n9962) );
  NAND2_X1 U5554 ( .A1(n6588), .A2(n8340), .ZN(n7465) );
  INV_X1 U5555 ( .A(n9837), .ZN(n9982) );
  OR2_X1 U5556 ( .A1(n7103), .A2(n8504), .ZN(n9831) );
  INV_X1 U5557 ( .A(n9559), .ZN(n4614) );
  NAND2_X1 U5558 ( .A1(n6394), .A2(n6393), .ZN(n9591) );
  NAND2_X1 U5559 ( .A1(n4750), .A2(n6363), .ZN(n9625) );
  INV_X1 U5560 ( .A(n7565), .ZN(n10043) );
  AND3_X1 U5561 ( .A1(n5971), .A2(n5970), .A3(n5969), .ZN(n10017) );
  NAND2_X1 U5562 ( .A1(n6500), .A2(n6499), .ZN(n8537) );
  AND2_X1 U5563 ( .A1(n4828), .A2(P1_IR_REG_28__SCAN_IN), .ZN(n4827) );
  OR2_X1 U5564 ( .A1(n4830), .A2(n4829), .ZN(n4828) );
  AND2_X1 U5565 ( .A1(n5840), .A2(n5843), .ZN(n4830) );
  INV_X1 U5566 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n4829) );
  INV_X1 U5567 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n5843) );
  XNOR2_X1 U5568 ( .A(n5705), .B(n5704), .ZN(n7949) );
  NAND2_X1 U5569 ( .A1(n5136), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5854) );
  NAND2_X1 U5570 ( .A1(n5854), .A2(n5853), .ZN(n5856) );
  NAND2_X1 U5571 ( .A1(n4815), .A2(n4814), .ZN(n5857) );
  NAND2_X1 U5572 ( .A1(n5664), .A2(n5285), .ZN(n5679) );
  OAI21_X1 U5573 ( .B1(n5586), .B2(n5585), .A(n5260), .ZN(n5598) );
  INV_X1 U5574 ( .A(n4745), .ZN(n5553) );
  NAND2_X1 U5575 ( .A1(n5522), .A2(n5248), .ZN(n5535) );
  OAI21_X1 U5576 ( .B1(n5242), .B2(SI_12_), .A(n5243), .ZN(n5504) );
  AND2_X1 U5577 ( .A1(n4790), .A2(n4538), .ZN(n4789) );
  INV_X1 U5578 ( .A(n5504), .ZN(n4790) );
  NAND2_X1 U5579 ( .A1(n5452), .A2(n5451), .ZN(n5237) );
  NOR2_X1 U5580 ( .A1(n6070), .A2(n6069), .ZN(n6073) );
  NAND2_X1 U5581 ( .A1(n5338), .A2(n5213), .ZN(n5353) );
  AND2_X1 U5582 ( .A1(n5448), .A2(n5447), .ZN(n7621) );
  AND2_X1 U5583 ( .A1(n5534), .A2(n5533), .ZN(n7985) );
  OR2_X1 U5584 ( .A1(n8578), .A2(n8587), .ZN(n8579) );
  NAND2_X1 U5585 ( .A1(n8545), .A2(n8544), .ZN(n8642) );
  OR2_X1 U5586 ( .A1(n8543), .A2(n8542), .ZN(n8544) );
  AND2_X1 U5587 ( .A1(n5703), .A2(n5702), .ZN(n8667) );
  NAND2_X1 U5588 ( .A1(n7082), .A2(n7081), .ZN(n7116) );
  INV_X1 U5589 ( .A(n7085), .ZN(n7081) );
  AND3_X1 U5590 ( .A1(n5626), .A2(n5625), .A3(n5624), .ZN(n9007) );
  INV_X1 U5591 ( .A(n8667), .ZN(n8935) );
  INV_X1 U5592 ( .A(n8678), .ZN(n8982) );
  OR2_X1 U5593 ( .A1(n5432), .A2(n5431), .ZN(n8740) );
  OR2_X1 U5594 ( .A1(n5387), .A2(n5386), .ZN(n7458) );
  OR2_X1 U5595 ( .A1(n7532), .A2(n5347), .ZN(n5350) );
  OAI21_X1 U5596 ( .B1(n7530), .B2(n5321), .A(n5067), .ZN(n5322) );
  NAND2_X1 U5597 ( .A1(n5635), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n5315) );
  NAND2_X1 U5598 ( .A1(n6915), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n6989) );
  NAND2_X1 U5599 ( .A1(n7145), .A2(n7172), .ZN(n7176) );
  XNOR2_X1 U5600 ( .A(n8842), .B(n8841), .ZN(n8803) );
  INV_X1 U5601 ( .A(n8846), .ZN(n8840) );
  OR2_X1 U5602 ( .A1(n4642), .A2(n8820), .ZN(n4641) );
  AND2_X1 U5603 ( .A1(n8808), .A2(n8807), .ZN(n4642) );
  OR2_X1 U5604 ( .A1(n6932), .A2(n8266), .ZN(n10127) );
  NAND2_X1 U5605 ( .A1(n5621), .A2(n5620), .ZN(n9067) );
  OAI21_X1 U5606 ( .B1(n6696), .B2(n5339), .A(n5472), .ZN(n7777) );
  INV_X1 U5607 ( .A(n10141), .ZN(n9031) );
  NAND2_X1 U5608 ( .A1(n5735), .A2(n5734), .ZN(n5824) );
  NAND2_X1 U5609 ( .A1(n8200), .A2(n8199), .ZN(n9081) );
  AND2_X1 U5610 ( .A1(n5785), .A2(n6829), .ZN(n5786) );
  NOR2_X1 U5611 ( .A1(n6456), .A2(n6455), .ZN(n6457) );
  XNOR2_X1 U5612 ( .A(n4597), .B(n8581), .ZN(n6458) );
  NOR2_X1 U5613 ( .A1(n8587), .A2(n9006), .ZN(n6455) );
  NAND2_X1 U5614 ( .A1(n6628), .A2(n5122), .ZN(n5121) );
  NAND2_X1 U5615 ( .A1(n5123), .A2(n5126), .ZN(n5122) );
  NAND2_X1 U5616 ( .A1(n6493), .A2(n6492), .ZN(n9556) );
  NAND2_X1 U5617 ( .A1(n6331), .A2(n6330), .ZN(n9671) );
  AND2_X1 U5618 ( .A1(n6437), .A2(n9970), .ZN(n9946) );
  AND2_X1 U5619 ( .A1(n6445), .A2(n6435), .ZN(n9948) );
  INV_X1 U5620 ( .A(n9337), .ZN(n9404) );
  NOR2_X1 U5621 ( .A1(n7355), .A2(n4723), .ZN(n7357) );
  AND2_X1 U5622 ( .A1(n7360), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n4723) );
  NAND2_X1 U5623 ( .A1(n7357), .A2(n7356), .ZN(n7490) );
  NOR2_X1 U5624 ( .A1(n7491), .A2(n7492), .ZN(n7606) );
  NAND2_X1 U5625 ( .A1(n5863), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4813) );
  OAI21_X1 U5626 ( .B1(n9507), .B2(n4695), .A(n8536), .ZN(n4727) );
  NAND2_X1 U5627 ( .A1(n6613), .A2(n9837), .ZN(n4612) );
  NAND2_X1 U5628 ( .A1(n9573), .A2(n8286), .ZN(n9532) );
  NAND2_X1 U5629 ( .A1(n5016), .A2(n4517), .ZN(n9542) );
  NAND2_X1 U5630 ( .A1(n5016), .A2(n5015), .ZN(n6579) );
  NAND2_X1 U5631 ( .A1(n9974), .A2(n7262), .ZN(n9929) );
  NAND2_X1 U5632 ( .A1(n6164), .A2(n6163), .ZN(n7842) );
  NAND2_X1 U5633 ( .A1(n9763), .A2(n4796), .ZN(n9848) );
  AND2_X1 U5634 ( .A1(n9764), .A2(n9765), .ZN(n4796) );
  AND2_X1 U5635 ( .A1(n6416), .A2(n6415), .ZN(n9894) );
  NAND2_X1 U5636 ( .A1(n4846), .A2(n4844), .ZN(n4843) );
  NAND2_X1 U5637 ( .A1(n4664), .A2(n8423), .ZN(n4820) );
  NOR2_X1 U5638 ( .A1(n8160), .A2(n8953), .ZN(n4702) );
  NAND2_X1 U5639 ( .A1(n4817), .A2(n4816), .ZN(n8429) );
  AND2_X1 U5640 ( .A1(n9617), .A2(n8425), .ZN(n4816) );
  NOR2_X1 U5641 ( .A1(n4536), .A2(n4836), .ZN(n4835) );
  NOR2_X1 U5642 ( .A1(n8433), .A2(n8453), .ZN(n4836) );
  AND2_X1 U5643 ( .A1(n8434), .A2(n4833), .ZN(n4832) );
  AND2_X1 U5644 ( .A1(n8432), .A2(n8453), .ZN(n4833) );
  NOR2_X1 U5645 ( .A1(n5044), .A2(n5614), .ZN(n5042) );
  NOR2_X1 U5646 ( .A1(n4718), .A2(n8203), .ZN(n4717) );
  INV_X1 U5647 ( .A(n8171), .ZN(n4718) );
  AND2_X1 U5648 ( .A1(n8910), .A2(n8177), .ZN(n4714) );
  INV_X1 U5649 ( .A(n8182), .ZN(n4712) );
  AOI21_X1 U5650 ( .B1(n4653), .B2(n4652), .A(n4651), .ZN(n4650) );
  INV_X1 U5651 ( .A(n9543), .ZN(n4651) );
  OR2_X1 U5652 ( .A1(n4623), .A2(n4622), .ZN(n4621) );
  INV_X1 U5653 ( .A(n8422), .ZN(n4622) );
  NAND2_X1 U5654 ( .A1(n5055), .A2(n5054), .ZN(n6478) );
  AOI21_X1 U5655 ( .B1(n5056), .B2(n5058), .A(n4591), .ZN(n5054) );
  INV_X1 U5656 ( .A(n5052), .ZN(n5051) );
  OAI21_X1 U5657 ( .B1(n5284), .B2(n5053), .A(n5678), .ZN(n5052) );
  INV_X1 U5658 ( .A(n5285), .ZN(n5053) );
  AOI21_X1 U5659 ( .B1(n5035), .B2(n5036), .A(n4585), .ZN(n5034) );
  INV_X1 U5660 ( .A(n5040), .ZN(n5035) );
  AND2_X1 U5661 ( .A1(n4757), .A2(n5036), .ZN(n4755) );
  AOI21_X1 U5662 ( .B1(n5042), .B2(n4759), .A(n4758), .ZN(n4757) );
  INV_X1 U5663 ( .A(n5269), .ZN(n4758) );
  INV_X1 U5664 ( .A(n5046), .ZN(n4759) );
  INV_X1 U5665 ( .A(n5042), .ZN(n4760) );
  INV_X1 U5666 ( .A(SI_17_), .ZN(n10511) );
  OR2_X1 U5667 ( .A1(n6667), .A2(P2_D_REG_0__SCAN_IN), .ZN(n4965) );
  INV_X1 U5668 ( .A(n8620), .ZN(n4974) );
  OR2_X1 U5669 ( .A1(n8640), .A2(n9026), .ZN(n8546) );
  NOR2_X1 U5670 ( .A1(n4710), .A2(n8254), .ZN(n4709) );
  NOR2_X1 U5671 ( .A1(n4931), .A2(n7284), .ZN(n4930) );
  INV_X1 U5672 ( .A(n6965), .ZN(n4931) );
  INV_X1 U5673 ( .A(n6949), .ZN(n4957) );
  INV_X1 U5674 ( .A(n4865), .ZN(n4859) );
  NAND2_X1 U5675 ( .A1(n4849), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n4848) );
  NAND2_X1 U5676 ( .A1(n4855), .A2(n4850), .ZN(n4849) );
  OR2_X1 U5677 ( .A1(n7576), .A2(n4636), .ZN(n4635) );
  NOR2_X1 U5678 ( .A1(n7382), .A2(n7774), .ZN(n4636) );
  AND2_X1 U5679 ( .A1(n4960), .A2(n4959), .ZN(n8745) );
  NAND2_X1 U5680 ( .A1(n8759), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n4959) );
  INV_X1 U5681 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n10602) );
  INV_X1 U5682 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n10556) );
  INV_X1 U5683 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n7700) );
  OAI21_X1 U5684 ( .B1(n5449), .B2(n4902), .A(n5463), .ZN(n4901) );
  AND2_X1 U5685 ( .A1(n8114), .A2(n8113), .ZN(n4692) );
  INV_X1 U5686 ( .A(n5105), .ZN(n5098) );
  INV_X1 U5687 ( .A(n8101), .ZN(n5097) );
  AND2_X1 U5688 ( .A1(n8729), .A2(n8901), .ZN(n8173) );
  NOR2_X1 U5689 ( .A1(n9009), .A2(n5080), .ZN(n5079) );
  INV_X1 U5690 ( .A(n8053), .ZN(n5080) );
  INV_X1 U5691 ( .A(n8242), .ZN(n4913) );
  INV_X1 U5692 ( .A(n4911), .ZN(n4906) );
  OR2_X1 U5693 ( .A1(n9153), .A2(n9005), .ZN(n8243) );
  INV_X1 U5694 ( .A(n8143), .ZN(n5109) );
  INV_X1 U5695 ( .A(n5111), .ZN(n5110) );
  NAND2_X1 U5696 ( .A1(n4678), .A2(n8057), .ZN(n4677) );
  INV_X1 U5697 ( .A(n8235), .ZN(n4678) );
  INV_X1 U5698 ( .A(P2_B_REG_SCAN_IN), .ZN(n5790) );
  INV_X1 U5699 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n5186) );
  NOR2_X1 U5700 ( .A1(n4523), .A2(P2_IR_REG_17__SCAN_IN), .ZN(n4996) );
  NOR2_X1 U5701 ( .A1(n6297), .A2(n5888), .ZN(n5887) );
  AND2_X1 U5702 ( .A1(n6231), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n6255) );
  NOR2_X1 U5703 ( .A1(n4802), .A2(n9287), .ZN(n4801) );
  NOR2_X1 U5704 ( .A1(n4803), .A2(n4528), .ZN(n4802) );
  INV_X1 U5705 ( .A(n4804), .ZN(n4803) );
  NOR2_X1 U5706 ( .A1(n8484), .A2(n8448), .ZN(n8449) );
  AND2_X1 U5707 ( .A1(n9531), .A2(n4781), .ZN(n4780) );
  NAND2_X1 U5708 ( .A1(n9564), .A2(n8286), .ZN(n4781) );
  INV_X1 U5709 ( .A(n6560), .ZN(n5024) );
  AND2_X1 U5710 ( .A1(n9702), .A2(n5031), .ZN(n5030) );
  NAND2_X1 U5711 ( .A1(n6555), .A2(n6556), .ZN(n5031) );
  NOR2_X1 U5712 ( .A1(n9815), .A2(n4767), .ZN(n4766) );
  INV_X1 U5713 ( .A(n4768), .ZN(n4767) );
  OR2_X1 U5714 ( .A1(n9815), .A2(n9316), .ZN(n8334) );
  NOR2_X1 U5715 ( .A1(n6167), .A2(n6166), .ZN(n6165) );
  NAND2_X1 U5716 ( .A1(n9752), .A2(n8385), .ZN(n4776) );
  INV_X1 U5717 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n6140) );
  INV_X1 U5718 ( .A(n8344), .ZN(n8340) );
  NAND2_X1 U5719 ( .A1(n7397), .A2(n7420), .ZN(n7418) );
  NAND2_X1 U5720 ( .A1(n7898), .A2(n6501), .ZN(n4750) );
  XNOR2_X1 U5721 ( .A(n6478), .B(n6477), .ZN(n6480) );
  AND2_X1 U5722 ( .A1(n5718), .A2(n5304), .ZN(n5305) );
  AND2_X1 U5723 ( .A1(n5299), .A2(n5298), .ZN(n5704) );
  AND2_X1 U5724 ( .A1(n5293), .A2(n5292), .ZN(n5693) );
  NAND2_X1 U5725 ( .A1(n5270), .A2(n5627), .ZN(n5039) );
  OR2_X1 U5726 ( .A1(n5270), .A2(n5627), .ZN(n5040) );
  INV_X1 U5727 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n5837) );
  AND3_X1 U5728 ( .A1(n5830), .A2(n5828), .A3(n5829), .ZN(n4999) );
  INV_X1 U5729 ( .A(SI_20_), .ZN(n5627) );
  NAND2_X1 U5730 ( .A1(n5257), .A2(n10511), .ZN(n5260) );
  INV_X1 U5731 ( .A(SI_16_), .ZN(n10554) );
  INV_X1 U5732 ( .A(n5063), .ZN(n5060) );
  AOI21_X1 U5733 ( .B1(n4785), .B2(n4789), .A(n4784), .ZN(n4783) );
  INV_X1 U5734 ( .A(n4789), .ZN(n4786) );
  INV_X1 U5735 ( .A(n5243), .ZN(n4784) );
  AND2_X1 U5736 ( .A1(n5248), .A2(n5247), .ZN(n5519) );
  OR2_X1 U5737 ( .A1(n6157), .A2(n6156), .ZN(n6161) );
  XNOR2_X1 U5738 ( .A(n5241), .B(SI_11_), .ZN(n5479) );
  OR2_X1 U5739 ( .A1(n6114), .A2(P1_IR_REG_9__SCAN_IN), .ZN(n6157) );
  INV_X1 U5740 ( .A(SI_5_), .ZN(n10574) );
  NAND2_X1 U5741 ( .A1(n4970), .A2(n4974), .ZN(n4969) );
  INV_X1 U5742 ( .A(n4971), .ZN(n4970) );
  AOI21_X1 U5743 ( .B1(n8672), .B2(n8673), .A(n4972), .ZN(n4971) );
  INV_X1 U5744 ( .A(n8619), .ZN(n4972) );
  AND2_X1 U5745 ( .A1(n8712), .A2(n8572), .ZN(n8631) );
  OR2_X1 U5746 ( .A1(n8547), .A2(n8653), .ZN(n5139) );
  NAND2_X1 U5747 ( .A1(n8642), .A2(n8546), .ZN(n4994) );
  AND2_X1 U5748 ( .A1(n8630), .A2(n8568), .ZN(n8661) );
  OAI21_X1 U5749 ( .B1(n8674), .B2(n8673), .A(n8672), .ZN(n8671) );
  NOR2_X1 U5750 ( .A1(n7952), .A2(n5140), .ZN(n7955) );
  AND2_X1 U5751 ( .A1(n4967), .A2(n4525), .ZN(n8688) );
  XNOR2_X1 U5752 ( .A(n7074), .B(n7431), .ZN(n6880) );
  XNOR2_X1 U5753 ( .A(n10143), .B(n7074), .ZN(n7077) );
  AOI21_X1 U5754 ( .B1(n4989), .B2(n4991), .A(n4987), .ZN(n4986) );
  INV_X1 U5755 ( .A(n4992), .ZN(n4991) );
  OR2_X1 U5756 ( .A1(n5092), .A2(n5091), .ZN(n5088) );
  NOR2_X1 U5757 ( .A1(n5094), .A2(n8214), .ZN(n5092) );
  NAND2_X1 U5758 ( .A1(n5818), .A2(n8205), .ZN(n8258) );
  XNOR2_X1 U5759 ( .A(n5310), .B(n5309), .ZN(n5772) );
  NAND2_X1 U5760 ( .A1(n4537), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5310) );
  INV_X1 U5762 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n6943) );
  NAND2_X1 U5763 ( .A1(n6964), .A2(n6965), .ZN(n6963) );
  NAND2_X1 U5764 ( .A1(n6962), .A2(n6961), .ZN(n6960) );
  NAND2_X1 U5765 ( .A1(n6963), .A2(n4937), .ZN(n4933) );
  INV_X1 U5766 ( .A(n4927), .ZN(n4937) );
  NAND2_X1 U5767 ( .A1(n7060), .A2(n4956), .ZN(n4955) );
  AND2_X1 U5768 ( .A1(n4863), .A2(n4862), .ZN(n4861) );
  NOR2_X1 U5769 ( .A1(n4865), .A2(n5385), .ZN(n4863) );
  NAND2_X1 U5770 ( .A1(n4864), .A2(n4867), .ZN(n7173) );
  NAND2_X1 U5771 ( .A1(n7060), .A2(n6949), .ZN(n4947) );
  OR2_X1 U5772 ( .A1(n5486), .A2(n5488), .ZN(n5454) );
  AND2_X1 U5773 ( .A1(n7156), .A2(n7127), .ZN(n4639) );
  OAI21_X1 U5774 ( .B1(n7126), .B2(n4638), .A(n4560), .ZN(n7193) );
  OR2_X1 U5775 ( .A1(n7163), .A2(n4638), .ZN(n4637) );
  INV_X1 U5776 ( .A(n7127), .ZN(n4638) );
  NOR2_X1 U5777 ( .A1(n7378), .A2(n4961), .ZN(n7381) );
  INV_X1 U5778 ( .A(n7318), .ZN(n4961) );
  NOR2_X1 U5779 ( .A1(n7381), .A2(n7380), .ZN(n7576) );
  XNOR2_X1 U5780 ( .A(n4635), .B(n7581), .ZN(n7578) );
  AOI21_X1 U5781 ( .B1(P2_REG1_REG_10__SCAN_IN), .B2(n7577), .A(n7568), .ZN(
        n7680) );
  XNOR2_X1 U5782 ( .A(n8745), .B(n8760), .ZN(n10104) );
  NOR2_X1 U5783 ( .A1(n8762), .A2(n10108), .ZN(n10125) );
  NOR2_X1 U5784 ( .A1(n10104), .A2(n10105), .ZN(n10103) );
  NOR2_X1 U5785 ( .A1(n8790), .A2(n8791), .ZN(n8794) );
  INV_X1 U5786 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n8869) );
  NAND2_X1 U5787 ( .A1(n4885), .A2(n4887), .ZN(n4884) );
  NAND2_X1 U5788 ( .A1(n8254), .A2(n4518), .ZN(n4887) );
  NAND2_X1 U5789 ( .A1(n8899), .A2(n4882), .ZN(n4881) );
  AND2_X1 U5790 ( .A1(n4885), .A2(n4579), .ZN(n4882) );
  NAND2_X1 U5791 ( .A1(n5170), .A2(n5169), .ZN(n5722) );
  INV_X1 U5792 ( .A(n5710), .ZN(n5170) );
  NAND2_X1 U5793 ( .A1(n5166), .A2(n5165), .ZN(n5696) );
  AND3_X1 U5794 ( .A1(n5638), .A2(n5637), .A3(n5636), .ZN(n8995) );
  NAND2_X1 U5795 ( .A1(n5161), .A2(n10556), .ZN(n5605) );
  INV_X1 U5796 ( .A(n5591), .ZN(n5161) );
  NAND2_X1 U5797 ( .A1(n5160), .A2(n5159), .ZN(n5578) );
  INV_X1 U5798 ( .A(n5560), .ZN(n5160) );
  NAND2_X1 U5799 ( .A1(n5158), .A2(n10513), .ZN(n5543) );
  INV_X1 U5800 ( .A(n5529), .ZN(n5158) );
  AND2_X1 U5801 ( .A1(n8206), .A2(n8873), .ZN(n6467) );
  INV_X1 U5802 ( .A(n8735), .ZN(n7959) );
  NAND2_X1 U5803 ( .A1(n5156), .A2(n5155), .ZN(n5473) );
  INV_X1 U5804 ( .A(n5457), .ZN(n5156) );
  OR2_X1 U5805 ( .A1(n5442), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n5457) );
  NAND2_X1 U5806 ( .A1(n5154), .A2(n5153), .ZN(n5442) );
  INV_X1 U5807 ( .A(n5428), .ZN(n5154) );
  NAND2_X1 U5808 ( .A1(n5152), .A2(n5151), .ZN(n5406) );
  INV_X1 U5809 ( .A(n8058), .ZN(n5751) );
  AND2_X1 U5810 ( .A1(n8882), .A2(n8881), .ZN(n9082) );
  NAND2_X1 U5811 ( .A1(n5695), .A2(n5694), .ZN(n8628) );
  AOI21_X1 U5812 ( .B1(n4894), .B2(n4896), .A(n4892), .ZN(n4891) );
  INV_X1 U5813 ( .A(n4897), .ZN(n4896) );
  NOR2_X1 U5814 ( .A1(n8050), .A2(n5069), .ZN(n5068) );
  INV_X1 U5815 ( .A(n8150), .ZN(n5069) );
  NAND2_X1 U5816 ( .A1(n5081), .A2(n5079), .ZN(n9072) );
  NAND2_X1 U5817 ( .A1(n5604), .A2(n5603), .ZN(n8699) );
  AND2_X1 U5818 ( .A1(n4682), .A2(n8119), .ZN(n4681) );
  OR2_X1 U5819 ( .A1(n8174), .A2(n6835), .ZN(n6899) );
  XNOR2_X1 U5820 ( .A(n5795), .B(P2_IR_REG_26__SCAN_IN), .ZN(n5804) );
  NAND2_X1 U5821 ( .A1(n5084), .A2(n5086), .ZN(n5787) );
  XNOR2_X1 U5822 ( .A(n5745), .B(P2_IR_REG_21__SCAN_IN), .ZN(n6834) );
  OR2_X1 U5823 ( .A1(n5748), .A2(n5488), .ZN(n5745) );
  AND2_X1 U5824 ( .A1(n5486), .A2(n5485), .ZN(n5490) );
  XNOR2_X1 U5825 ( .A(n5400), .B(P2_IR_REG_6__SCAN_IN), .ZN(n7147) );
  INV_X1 U5826 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n5388) );
  INV_X1 U5827 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n6044) );
  NOR2_X1 U5828 ( .A1(n9186), .A2(n4805), .ZN(n4804) );
  INV_X1 U5829 ( .A(n4807), .ZN(n4805) );
  NAND2_X1 U5830 ( .A1(n6346), .A2(n9333), .ZN(n4807) );
  NAND2_X1 U5831 ( .A1(n9336), .A2(n4528), .ZN(n4806) );
  CLKBUF_X1 U5832 ( .A(n9908), .Z(n9909) );
  OR2_X1 U5833 ( .A1(n6311), .A2(n6295), .ZN(n6297) );
  OR2_X1 U5834 ( .A1(n6045), .A2(n6044), .ZN(n6079) );
  INV_X1 U5835 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n6078) );
  NAND2_X1 U5836 ( .A1(n7557), .A2(n6066), .ZN(n6094) );
  NAND2_X1 U5837 ( .A1(n5910), .A2(n5909), .ZN(n4824) );
  INV_X1 U5838 ( .A(n5134), .ZN(n5130) );
  AND2_X1 U5839 ( .A1(n9313), .A2(n9312), .ZN(n5134) );
  INV_X1 U5840 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n6166) );
  AND2_X1 U5841 ( .A1(n6376), .A2(n6375), .ZN(n9286) );
  AND2_X1 U5842 ( .A1(n6327), .A2(n6292), .ZN(n5133) );
  NAND2_X1 U5843 ( .A1(n9322), .A2(n9324), .ZN(n9323) );
  INV_X1 U5844 ( .A(n9347), .ZN(n5119) );
  NAND2_X1 U5845 ( .A1(n6255), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n6309) );
  INV_X1 U5846 ( .A(n9254), .ZN(n5126) );
  NOR2_X1 U5847 ( .A1(n6446), .A2(n9893), .ZN(n6445) );
  XNOR2_X1 U5848 ( .A(n6433), .B(n6432), .ZN(n6769) );
  AND4_X1 U5849 ( .A1(n6317), .A2(n6316), .A3(n6315), .A4(n6314), .ZN(n9281)
         );
  AND4_X1 U5850 ( .A1(n6238), .A2(n6237), .A3(n6236), .A4(n6235), .ZN(n9269)
         );
  AND4_X1 U5851 ( .A1(n6192), .A2(n6191), .A3(n6190), .A4(n6189), .ZN(n9177)
         );
  AND4_X1 U5852 ( .A1(n6172), .A2(n6171), .A3(n6170), .A4(n6169), .ZN(n7824)
         );
  AND4_X1 U5853 ( .A1(n6146), .A2(n6145), .A3(n6144), .A4(n6143), .ZN(n7807)
         );
  AOI21_X1 U5854 ( .B1(n6860), .B2(P1_REG2_REG_8__SCAN_IN), .A(n6859), .ZN(
        n6863) );
  AOI21_X1 U5855 ( .B1(P1_REG2_REG_11__SCAN_IN), .B2(n7360), .A(n7359), .ZN(
        n7481) );
  XNOR2_X1 U5856 ( .A(n7879), .B(n4737), .ZN(n9484) );
  NOR2_X1 U5857 ( .A1(n7878), .A2(n4738), .ZN(n7879) );
  AND2_X1 U5858 ( .A1(n7887), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n4738) );
  NOR2_X1 U5859 ( .A1(n9484), .A2(n6230), .ZN(n9485) );
  NOR2_X1 U5860 ( .A1(n7889), .A2(n9475), .ZN(n7893) );
  AND2_X1 U5861 ( .A1(n4999), .A2(n6248), .ZN(n5835) );
  AOI21_X1 U5862 ( .B1(P1_REG2_REG_16__SCAN_IN), .B2(n8528), .A(n8521), .ZN(
        n9492) );
  AOI21_X1 U5863 ( .B1(n4780), .B2(n4782), .A(n4779), .ZN(n4778) );
  INV_X1 U5864 ( .A(n8286), .ZN(n4782) );
  INV_X1 U5865 ( .A(n9533), .ZN(n4779) );
  NOR2_X1 U5866 ( .A1(n9566), .A2(n9556), .ZN(n9546) );
  NAND2_X1 U5867 ( .A1(n9546), .A2(n9852), .ZN(n9545) );
  AOI21_X1 U5868 ( .B1(n9568), .B2(n6577), .A(n6441), .ZN(n6622) );
  INV_X1 U5869 ( .A(n9199), .ZN(n9537) );
  AND2_X1 U5870 ( .A1(n8433), .A2(n9533), .ZN(n9531) );
  AND2_X1 U5871 ( .A1(n6572), .A2(n9548), .ZN(n9555) );
  NAND2_X1 U5872 ( .A1(n4627), .A2(n9584), .ZN(n4626) );
  NAND2_X1 U5873 ( .A1(n4628), .A2(n4631), .ZN(n4627) );
  NAND2_X1 U5874 ( .A1(n4770), .A2(n9570), .ZN(n9566) );
  OAI21_X1 U5875 ( .B1(n9635), .B2(n4631), .A(n4628), .ZN(n9585) );
  AND2_X1 U5876 ( .A1(n6382), .A2(n6396), .ZN(n9608) );
  AND2_X1 U5877 ( .A1(n8427), .A2(n9600), .ZN(n9617) );
  OAI21_X1 U5878 ( .B1(n9713), .B2(n9712), .A(n8410), .ZN(n9703) );
  OR2_X1 U5879 ( .A1(n9703), .A2(n9702), .ZN(n9705) );
  NAND2_X1 U5880 ( .A1(n4515), .A2(n4766), .ZN(n9696) );
  INV_X1 U5881 ( .A(n8475), .ZN(n9712) );
  NAND2_X1 U5882 ( .A1(n4515), .A2(n6494), .ZN(n9737) );
  NAND2_X1 U5883 ( .A1(n6602), .A2(n8398), .ZN(n4794) );
  NOR2_X1 U5884 ( .A1(n9728), .A2(n4793), .ZN(n4792) );
  INV_X1 U5885 ( .A(n8398), .ZN(n4793) );
  NAND2_X1 U5886 ( .A1(n7924), .A2(n8394), .ZN(n9835) );
  INV_X1 U5887 ( .A(n5009), .ZN(n5008) );
  OAI21_X1 U5888 ( .B1(n7822), .B2(n5010), .A(n5012), .ZN(n5009) );
  AND2_X1 U5889 ( .A1(n9755), .A2(n4520), .ZN(n4761) );
  INV_X1 U5890 ( .A(n7822), .ZN(n8470) );
  NAND2_X1 U5891 ( .A1(n7652), .A2(n4763), .ZN(n7828) );
  NAND2_X1 U5892 ( .A1(n6542), .A2(n6541), .ZN(n7752) );
  NAND2_X1 U5893 ( .A1(n6598), .A2(n7739), .ZN(n7805) );
  AND2_X1 U5894 ( .A1(n8369), .A2(n8371), .ZN(n8471) );
  NAND3_X1 U5895 ( .A1(n8308), .A2(n8464), .A3(n6597), .ZN(n7739) );
  OR2_X1 U5896 ( .A1(n6079), .A2(n6078), .ZN(n6099) );
  INV_X1 U5897 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n6866) );
  NAND2_X1 U5898 ( .A1(n5002), .A2(n5001), .ZN(n7720) );
  AOI21_X1 U5899 ( .B1(n5004), .B2(n5006), .A(n4555), .ZN(n5001) );
  OR2_X1 U5900 ( .A1(n8358), .A2(n6538), .ZN(n7719) );
  OR2_X1 U5901 ( .A1(n9975), .A2(n9941), .ZN(n7709) );
  NAND2_X1 U5902 ( .A1(n9976), .A2(n10043), .ZN(n9975) );
  NOR2_X1 U5903 ( .A1(n6000), .A2(n7520), .ZN(n6023) );
  NAND2_X1 U5904 ( .A1(n4657), .A2(n8459), .ZN(n4655) );
  NAND2_X1 U5905 ( .A1(n8294), .A2(n4657), .ZN(n4656) );
  NOR2_X1 U5906 ( .A1(n6587), .A2(n4658), .ZN(n4657) );
  NAND2_X1 U5907 ( .A1(n4998), .A2(n9994), .ZN(n9992) );
  XNOR2_X1 U5908 ( .A(n5914), .B(n6524), .ZN(n4997) );
  AND2_X1 U5909 ( .A1(n8493), .A2(n6509), .ZN(n9935) );
  NAND2_X1 U5910 ( .A1(n6378), .A2(n6377), .ZN(n9609) );
  NAND2_X1 U5911 ( .A1(n5846), .A2(n5845), .ZN(n9800) );
  NAND2_X1 U5912 ( .A1(n5007), .A2(n6547), .ZN(n9751) );
  NAND2_X1 U5913 ( .A1(n7832), .A2(n7822), .ZN(n5007) );
  INV_X1 U5914 ( .A(n7655), .ZN(n10068) );
  INV_X1 U5915 ( .A(n6096), .ZN(n4633) );
  AND2_X1 U5916 ( .A1(n6434), .A2(n6581), .ZN(n10074) );
  INV_X1 U5917 ( .A(n10074), .ZN(n10067) );
  AND2_X1 U5918 ( .A1(n6515), .A2(n7101), .ZN(n6518) );
  XNOR2_X1 U5919 ( .A(n5731), .B(n5730), .ZN(n8274) );
  NAND2_X1 U5920 ( .A1(n5719), .A2(n5718), .ZN(n5731) );
  NAND2_X1 U5921 ( .A1(n5279), .A2(n5278), .ZN(n5661) );
  NAND2_X1 U5922 ( .A1(n5043), .A2(n5041), .ZN(n5615) );
  INV_X1 U5923 ( .A(n5044), .ZN(n5041) );
  NOR2_X1 U5924 ( .A1(n6161), .A2(P1_IR_REG_12__SCAN_IN), .ZN(n6202) );
  AND2_X1 U5925 ( .A1(n5422), .A2(n5421), .ZN(n6678) );
  AOI21_X1 U5926 ( .B1(n4699), .B2(n5373), .A(n4698), .ZN(n4697) );
  INV_X1 U5927 ( .A(n5373), .ZN(n4700) );
  INV_X1 U5928 ( .A(n5222), .ZN(n4698) );
  INV_X1 U5929 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n6007) );
  NAND2_X1 U5930 ( .A1(n5216), .A2(n4706), .ZN(n5354) );
  NAND2_X1 U5931 ( .A1(n4708), .A2(n4707), .ZN(n4706) );
  INV_X1 U5932 ( .A(SI_3_), .ZN(n4707) );
  INV_X1 U5933 ( .A(n5214), .ZN(n4708) );
  NAND2_X1 U5934 ( .A1(n5202), .A2(n5326), .ZN(n4739) );
  NAND2_X1 U5935 ( .A1(n5204), .A2(n5203), .ZN(n5205) );
  INV_X1 U5936 ( .A(n5325), .ZN(n5204) );
  NAND2_X1 U5937 ( .A1(n7443), .A2(n7442), .ZN(n7446) );
  AND2_X1 U5938 ( .A1(n5658), .A2(n5657), .ZN(n8684) );
  NAND2_X1 U5939 ( .A1(n7729), .A2(n7728), .ZN(n4985) );
  NAND2_X1 U5940 ( .A1(n4967), .A2(n4969), .ZN(n8622) );
  INV_X1 U5941 ( .A(n8736), .ZN(n7940) );
  AND2_X1 U5942 ( .A1(n4994), .A2(n4992), .ZN(n8703) );
  NAND2_X1 U5943 ( .A1(n4994), .A2(n5139), .ZN(n8650) );
  NAND2_X1 U5944 ( .A1(n4981), .A2(n4983), .ZN(n4977) );
  NAND2_X1 U5945 ( .A1(n4976), .A2(n4981), .ZN(n4975) );
  INV_X1 U5946 ( .A(n7942), .ZN(n4981) );
  INV_X1 U5947 ( .A(n4982), .ZN(n7852) );
  OAI21_X1 U5948 ( .B1(n7729), .B2(n4980), .A(n4978), .ZN(n4982) );
  NAND2_X1 U5949 ( .A1(n7300), .A2(n7299), .ZN(n7443) );
  NAND2_X1 U5950 ( .A1(n8008), .A2(n8007), .ZN(n8545) );
  INV_X1 U5951 ( .A(n8658), .ZN(n8717) );
  INV_X1 U5952 ( .A(n8859), .ZN(n8873) );
  XNOR2_X1 U5953 ( .A(n5744), .B(P2_IR_REG_22__SCAN_IN), .ZN(n8268) );
  INV_X1 U5954 ( .A(n8216), .ZN(n8882) );
  INV_X1 U5955 ( .A(n8684), .ZN(n8971) );
  INV_X1 U5956 ( .A(n7985), .ZN(n7981) );
  NAND2_X1 U5957 ( .A1(n5776), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n5334) );
  NOR2_X1 U5958 ( .A1(n6994), .A2(n4925), .ZN(n6999) );
  NAND2_X1 U5959 ( .A1(n7056), .A2(n4933), .ZN(n6979) );
  OR2_X1 U5960 ( .A1(n4954), .A2(n4953), .ZN(n7166) );
  NAND2_X1 U5961 ( .A1(n4955), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n4954) );
  INV_X1 U5962 ( .A(n7164), .ZN(n4953) );
  NAND2_X1 U5963 ( .A1(n4856), .A2(n7209), .ZN(n7150) );
  NAND2_X1 U5964 ( .A1(n7176), .A2(n4855), .ZN(n4856) );
  NAND2_X1 U5965 ( .A1(n4640), .A2(n7193), .ZN(n7129) );
  NAND2_X1 U5966 ( .A1(n4877), .A2(n4879), .ZN(n7336) );
  NOR2_X1 U5967 ( .A1(n4878), .A2(n7366), .ZN(n7365) );
  AND2_X1 U5968 ( .A1(n4877), .A2(n4878), .ZN(n7369) );
  OR2_X1 U5969 ( .A1(n7569), .A2(n5497), .ZN(n4876) );
  INV_X1 U5970 ( .A(n4960), .ZN(n8744) );
  NAND2_X1 U5971 ( .A1(n4872), .A2(n4871), .ZN(n8758) );
  XNOR2_X1 U5972 ( .A(n8788), .B(n8789), .ZN(n8748) );
  NOR2_X1 U5973 ( .A1(n8748), .A2(n7998), .ZN(n8790) );
  NOR2_X1 U5974 ( .A1(n8776), .A2(n8775), .ZN(n8779) );
  INV_X1 U5975 ( .A(n4869), .ZN(n8774) );
  NOR2_X1 U5976 ( .A1(n8779), .A2(n8778), .ZN(n8801) );
  NAND2_X1 U5977 ( .A1(n4944), .A2(n8862), .ZN(n4943) );
  NAND2_X1 U5978 ( .A1(n4941), .A2(n4940), .ZN(n4939) );
  XNOR2_X1 U5979 ( .A(n8211), .B(n8184), .ZN(n8895) );
  AND2_X1 U5980 ( .A1(n6472), .A2(n5137), .ZN(n6473) );
  NAND2_X1 U5981 ( .A1(n5081), .A2(n8053), .ZN(n9010) );
  OR2_X1 U5982 ( .A1(n6467), .A2(n10187), .ZN(n10142) );
  NAND2_X1 U5983 ( .A1(n4684), .A2(n8115), .ZN(n7771) );
  NAND2_X1 U5984 ( .A1(n7634), .A2(n5450), .ZN(n7619) );
  NAND2_X1 U5985 ( .A1(n5101), .A2(n5103), .ZN(n7629) );
  AND2_X1 U5986 ( .A1(n4693), .A2(n8113), .ZN(n5103) );
  NAND2_X1 U5987 ( .A1(n7456), .A2(n5105), .ZN(n5101) );
  NAND2_X1 U5988 ( .A1(n5102), .A2(n8081), .ZN(n7498) );
  OR2_X1 U5989 ( .A1(n7456), .A2(n8091), .ZN(n5102) );
  INV_X1 U5990 ( .A(n8225), .ZN(n5072) );
  NAND2_X1 U5991 ( .A1(n7270), .A2(n8077), .ZN(n5073) );
  AND2_X1 U5992 ( .A1(n5362), .A2(n4535), .ZN(n5363) );
  NAND2_X1 U5993 ( .A1(n6730), .A2(n6465), .ZN(n10141) );
  NAND2_X1 U5994 ( .A1(n8187), .A2(n8186), .ZN(n9084) );
  NAND2_X1 U5995 ( .A1(n5312), .A2(n5311), .ZN(n9095) );
  NAND2_X1 U5996 ( .A1(n5075), .A2(n8043), .ZN(n8896) );
  NAND2_X1 U5997 ( .A1(n5707), .A2(n5706), .ZN(n9102) );
  NAND2_X1 U5998 ( .A1(n4687), .A2(n4688), .ZN(n8911) );
  NAND2_X1 U5999 ( .A1(n4921), .A2(n5690), .ZN(n8921) );
  NAND2_X1 U6000 ( .A1(n5765), .A2(n8218), .ZN(n8920) );
  NAND2_X1 U6001 ( .A1(n5681), .A2(n5680), .ZN(n9113) );
  NAND2_X1 U6002 ( .A1(n5677), .A2(n5676), .ZN(n8933) );
  NAND2_X1 U6003 ( .A1(n5667), .A2(n5666), .ZN(n9119) );
  NAND2_X1 U6004 ( .A1(n5653), .A2(n5652), .ZN(n9125) );
  NAND2_X1 U6005 ( .A1(n5644), .A2(n5643), .ZN(n9131) );
  NAND2_X1 U6006 ( .A1(n5632), .A2(n5631), .ZN(n9137) );
  AND2_X1 U6007 ( .A1(n4898), .A2(n4546), .ZN(n8980) );
  NAND2_X1 U6008 ( .A1(n8988), .A2(n8150), .ZN(n8978) );
  AND2_X1 U6009 ( .A1(n9028), .A2(n9027), .ZN(n9150) );
  NAND2_X1 U6010 ( .A1(n5575), .A2(n5574), .ZN(n8647) );
  AND2_X1 U6011 ( .A1(n8028), .A2(n8027), .ZN(n8038) );
  NAND2_X1 U6012 ( .A1(n5559), .A2(n5558), .ZN(n8006) );
  NAND2_X1 U6013 ( .A1(n5106), .A2(n5113), .ZN(n7989) );
  NAND2_X1 U6014 ( .A1(n7905), .A2(n5111), .ZN(n5106) );
  NAND2_X1 U6015 ( .A1(n5542), .A2(n5541), .ZN(n8015) );
  NAND2_X1 U6016 ( .A1(n5114), .A2(n8054), .ZN(n7974) );
  OR2_X1 U6017 ( .A1(n7905), .A2(n5761), .ZN(n5114) );
  NAND2_X1 U6018 ( .A1(n5526), .A2(n5525), .ZN(n7953) );
  INV_X1 U6019 ( .A(n9148), .ZN(n9152) );
  INV_X1 U6020 ( .A(n7428), .ZN(n7435) );
  AND2_X1 U6021 ( .A1(n6734), .A2(n6726), .ZN(n6730) );
  INV_X1 U6022 ( .A(n5792), .ZN(n4674) );
  NAND2_X1 U6023 ( .A1(n5189), .A2(n5188), .ZN(n8538) );
  CLKBUF_X1 U6024 ( .A(n5771), .Z(n8276) );
  NAND2_X1 U6025 ( .A1(n5792), .A2(n5793), .ZN(n7935) );
  NAND2_X1 U6026 ( .A1(n4529), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5791) );
  INV_X1 U6027 ( .A(n5803), .ZN(n7910) );
  INV_X1 U6028 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n7757) );
  INV_X1 U6029 ( .A(n8268), .ZN(n7758) );
  INV_X1 U6030 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n7616) );
  INV_X1 U6031 ( .A(n6834), .ZN(n5818) );
  INV_X1 U6032 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n7512) );
  INV_X1 U6033 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n7427) );
  INV_X1 U6034 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n7313) );
  INV_X1 U6035 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n5360) );
  NAND2_X1 U6036 ( .A1(n4646), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5361) );
  NAND2_X1 U6037 ( .A1(n4857), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5340) );
  INV_X1 U6038 ( .A(n6944), .ZN(n4857) );
  XNOR2_X1 U6039 ( .A(n5329), .B(n5328), .ZN(n6991) );
  NAND2_X1 U6040 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_31__SCAN_IN), .ZN(
        n5328) );
  AND2_X1 U6041 ( .A1(n6769), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6650) );
  INV_X1 U6042 ( .A(n4811), .ZN(n4810) );
  NAND2_X1 U6043 ( .A1(n6219), .A2(n6223), .ZN(n9175) );
  NAND2_X1 U6044 ( .A1(n4806), .A2(n4807), .ZN(n9185) );
  AND2_X1 U6045 ( .A1(n9225), .A2(n9948), .ZN(n9217) );
  CLKBUF_X1 U6046 ( .A(n9296), .Z(n9297) );
  INV_X1 U6047 ( .A(n5129), .ZN(n5128) );
  NOR2_X1 U6048 ( .A1(n5134), .A2(n5132), .ZN(n5131) );
  AOI21_X1 U6049 ( .B1(n5130), .B2(n4519), .A(n4565), .ZN(n5129) );
  AND2_X1 U6050 ( .A1(n5127), .A2(n9388), .ZN(n9264) );
  NAND2_X1 U6051 ( .A1(n6253), .A2(n6252), .ZN(n9833) );
  AOI21_X1 U6052 ( .B1(n9275), .B2(n5133), .A(n4519), .ZN(n9315) );
  NAND2_X1 U6053 ( .A1(n6307), .A2(n6306), .ZN(n9719) );
  AND3_X1 U6054 ( .A1(n6021), .A2(n6020), .A3(n6019), .ZN(n10039) );
  NAND2_X1 U6055 ( .A1(n9252), .A2(n9254), .ZN(n9253) );
  OAI21_X1 U6056 ( .B1(n9857), .B2(n9946), .A(n6450), .ZN(n6451) );
  INV_X1 U6057 ( .A(n9946), .ZN(n9395) );
  INV_X1 U6058 ( .A(n9948), .ZN(n9916) );
  INV_X1 U6059 ( .A(n4741), .ZN(n4740) );
  NAND2_X1 U6060 ( .A1(n4744), .A2(n4743), .ZN(n4742) );
  NAND2_X1 U6061 ( .A1(n4568), .A2(n4669), .ZN(n4668) );
  NAND2_X1 U6062 ( .A1(n8508), .A2(n4509), .ZN(n4670) );
  NOR2_X1 U6063 ( .A1(n8515), .A2(n8511), .ZN(n4669) );
  INV_X1 U6064 ( .A(n9281), .ZN(n9407) );
  INV_X1 U6065 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n5207) );
  OR2_X1 U6066 ( .A1(n5939), .A2(n5938), .ZN(n5940) );
  OR2_X1 U6067 ( .A1(n6027), .A2(n7106), .ZN(n5920) );
  OAI21_X1 U6068 ( .B1(n9436), .B2(n5937), .A(n4603), .ZN(n9443) );
  NAND2_X1 U6069 ( .A1(n9436), .A2(n5937), .ZN(n4603) );
  NAND2_X1 U6070 ( .A1(n9442), .A2(n9443), .ZN(n9441) );
  AOI21_X1 U6071 ( .B1(n9464), .B2(P1_REG2_REG_5__SCAN_IN), .A(n9465), .ZN(
        n6806) );
  INV_X1 U6072 ( .A(n4733), .ZN(n6807) );
  INV_X1 U6073 ( .A(n4735), .ZN(n6809) );
  NAND2_X1 U6074 ( .A1(n6810), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n4732) );
  NOR2_X1 U6075 ( .A1(n6855), .A2(n4725), .ZN(n6858) );
  AND2_X1 U6076 ( .A1(n6860), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n4725) );
  NAND2_X1 U6077 ( .A1(n6858), .A2(n6857), .ZN(n7039) );
  NOR2_X1 U6078 ( .A1(n7043), .A2(n7042), .ZN(n7225) );
  NAND2_X1 U6079 ( .A1(n7039), .A2(n4724), .ZN(n7043) );
  OR2_X1 U6080 ( .A1(n7040), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n4724) );
  NAND2_X1 U6081 ( .A1(n7490), .A2(n7489), .ZN(n7491) );
  AOI21_X1 U6082 ( .B1(P1_REG2_REG_13__SCAN_IN), .B2(n7607), .A(n7602), .ZN(
        n7605) );
  AND2_X1 U6083 ( .A1(n5066), .A2(n6502), .ZN(n9933) );
  NAND2_X1 U6084 ( .A1(n8537), .A2(n6501), .ZN(n5066) );
  NAND2_X1 U6085 ( .A1(n5014), .A2(n5013), .ZN(n9544) );
  AOI21_X1 U6086 ( .B1(n4517), .B2(n9574), .A(n4551), .ZN(n5013) );
  NAND2_X1 U6087 ( .A1(n5018), .A2(n5019), .ZN(n9583) );
  OAI21_X1 U6088 ( .B1(n9616), .B2(n6564), .A(n6565), .ZN(n9599) );
  NAND2_X1 U6089 ( .A1(n9619), .A2(n4772), .ZN(n9604) );
  NAND2_X1 U6090 ( .A1(n6348), .A2(n6347), .ZN(n9791) );
  NAND2_X1 U6091 ( .A1(n4620), .A2(n8422), .ZN(n9656) );
  NAND2_X1 U6092 ( .A1(n9680), .A2(n4623), .ZN(n4620) );
  INV_X1 U6093 ( .A(n9800), .ZN(n9654) );
  OR2_X1 U6094 ( .A1(n9666), .A2(n9982), .ZN(n9669) );
  NAND2_X1 U6095 ( .A1(n9748), .A2(n8380), .ZN(n7925) );
  NAND2_X1 U6096 ( .A1(n6229), .A2(n6228), .ZN(n9396) );
  NAND2_X1 U6097 ( .A1(n5003), .A2(n6537), .ZN(n7660) );
  NAND2_X1 U6098 ( .A1(n9961), .A2(n9962), .ZN(n5003) );
  OR2_X1 U6099 ( .A1(n10000), .A2(n7108), .ZN(n9990) );
  OAI21_X1 U6100 ( .B1(n8294), .B2(n8459), .A(n8293), .ZN(n7392) );
  OR2_X1 U6101 ( .A1(n7109), .A2(n4509), .ZN(n9612) );
  INV_X1 U6102 ( .A(n9612), .ZN(n9996) );
  INV_X1 U6103 ( .A(n9990), .ZN(n9633) );
  NAND2_X1 U6104 ( .A1(n10100), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n4606) );
  NAND2_X1 U6105 ( .A1(n4611), .A2(n4609), .ZN(n6617) );
  INV_X1 U6106 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n4616) );
  INV_X1 U6107 ( .A(n9609), .ZN(n9861) );
  INV_X1 U6108 ( .A(n9396), .ZN(n9892) );
  AND2_X1 U6109 ( .A1(n4572), .A2(n4524), .ZN(n5032) );
  XNOR2_X1 U6110 ( .A(n6489), .B(n6488), .ZN(n9895) );
  AOI21_X1 U6111 ( .B1(n4827), .B2(n4829), .A(n4570), .ZN(n4826) );
  INV_X1 U6112 ( .A(n5840), .ZN(n4771) );
  INV_X1 U6113 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n10526) );
  OR2_X1 U6114 ( .A1(n5854), .A2(n5853), .ZN(n5855) );
  INV_X1 U6115 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n10588) );
  XNOR2_X1 U6116 ( .A(n5852), .B(n10441), .ZN(n7899) );
  INV_X1 U6117 ( .A(n5857), .ZN(n5839) );
  INV_X1 U6118 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n10389) );
  INV_X1 U6119 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n10406) );
  INV_X1 U6120 ( .A(n4509), .ZN(n8509) );
  INV_X1 U6121 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n10347) );
  NAND2_X1 U6122 ( .A1(n4791), .A2(n4789), .ZN(n5507) );
  NAND2_X1 U6123 ( .A1(n4791), .A2(n4538), .ZN(n5505) );
  NAND2_X1 U6124 ( .A1(n5468), .A2(n5469), .ZN(n6696) );
  NAND2_X1 U6125 ( .A1(n5237), .A2(n5236), .ZN(n5467) );
  OR2_X1 U6126 ( .A1(n6075), .A2(n6074), .ZN(n6688) );
  NAND2_X1 U6127 ( .A1(n5374), .A2(n5373), .ZN(n5376) );
  NAND2_X1 U6128 ( .A1(n5356), .A2(n5216), .ZN(n5374) );
  AOI22_X1 U6129 ( .A1(n4566), .A2(P1_IR_REG_0__SCAN_IN), .B1(n4731), .B2(
        n5848), .ZN(n4730) );
  NAND2_X1 U6130 ( .A1(n7116), .A2(n7115), .ZN(n7119) );
  NAND2_X1 U6131 ( .A1(n8872), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n6922) );
  AOI21_X1 U6132 ( .B1(n4641), .B2(n8878), .A(n4595), .ZN(n8817) );
  NAND2_X1 U6133 ( .A1(n4602), .A2(n4601), .ZN(P2_U3487) );
  INV_X1 U6134 ( .A(n9040), .ZN(n4601) );
  OAI22_X1 U6135 ( .A1(n8890), .A2(n9148), .B1(n10199), .B2(n5825), .ZN(n5826)
         );
  OAI21_X1 U6136 ( .B1(n9570), .B2(n9946), .A(n6638), .ZN(n6639) );
  AOI21_X1 U6137 ( .B1(n4728), .B2(n4509), .A(n4727), .ZN(n4726) );
  AND2_X1 U6138 ( .A1(n4612), .A2(n9222), .ZN(n9563) );
  NAND2_X1 U6139 ( .A1(n4607), .A2(n4604), .ZN(P1_U3550) );
  INV_X1 U6140 ( .A(n4605), .ZN(n4604) );
  NAND2_X1 U6141 ( .A1(n6617), .A2(n10102), .ZN(n4607) );
  OAI21_X1 U6142 ( .B1(n6616), .B2(n9846), .A(n4606), .ZN(n4605) );
  OAI21_X1 U6143 ( .B1(n9848), .B2(n10082), .A(n9850), .ZN(n9851) );
  NAND2_X1 U6144 ( .A1(n10082), .A2(n9849), .ZN(n9850) );
  NAND4_X2 U6145 ( .A1(n5904), .A2(n5903), .A3(n5902), .A4(n5901), .ZN(n5914)
         );
  NOR2_X1 U6146 ( .A1(n8015), .A2(n8734), .ZN(n4516) );
  AND2_X1 U6147 ( .A1(n6578), .A2(n5015), .ZN(n4517) );
  NAND2_X1 U6148 ( .A1(n9416), .A2(n10060), .ZN(n4632) );
  OR2_X1 U6149 ( .A1(n6326), .A2(n6325), .ZN(n4519) );
  AND2_X1 U6150 ( .A1(n4763), .A2(n4762), .ZN(n4520) );
  AND3_X1 U6151 ( .A1(n4564), .A2(n5906), .A3(n6248), .ZN(n4521) );
  AND2_X1 U6152 ( .A1(n4613), .A2(n10084), .ZN(n4522) );
  NAND2_X1 U6153 ( .A1(n8212), .A2(n8190), .ZN(n8254) );
  NAND2_X1 U6154 ( .A1(n5600), .A2(n5617), .ZN(n4523) );
  AND2_X1 U6155 ( .A1(n5843), .A2(n5033), .ZN(n4524) );
  AND2_X1 U6156 ( .A1(n4969), .A2(n4552), .ZN(n4525) );
  NAND2_X1 U6157 ( .A1(n5115), .A2(n8130), .ZN(n4526) );
  AND2_X1 U6158 ( .A1(n4916), .A2(n5309), .ZN(n4527) );
  OAI21_X1 U6159 ( .B1(n5113), .B2(n5109), .A(n8135), .ZN(n5107) );
  OR2_X1 U6160 ( .A1(n6346), .A2(n9333), .ZN(n4528) );
  INV_X1 U6161 ( .A(n8862), .ZN(n4946) );
  INV_X1 U6162 ( .A(n5910), .ZN(n6154) );
  INV_X2 U6163 ( .A(n7530), .ZN(n5348) );
  NAND2_X1 U6164 ( .A1(n4671), .A2(n4824), .ZN(n6524) );
  INV_X1 U6165 ( .A(n6524), .ZN(n4998) );
  NAND4_X1 U6166 ( .A1(n5920), .A2(n5919), .A3(n5918), .A4(n5917), .ZN(n5927)
         );
  NAND3_X1 U6167 ( .A1(n5084), .A2(n5086), .A3(n5085), .ZN(n4529) );
  AND2_X1 U6168 ( .A1(n4853), .A2(n7149), .ZN(n4530) );
  OR2_X1 U6169 ( .A1(n9649), .A2(n9791), .ZN(n4531) );
  INV_X1 U6170 ( .A(n7420), .ZN(n10031) );
  AND3_X1 U6171 ( .A1(n6012), .A2(n6011), .A3(n6010), .ZN(n7420) );
  AND2_X1 U6172 ( .A1(n4621), .A2(n9655), .ZN(n4532) );
  AOI21_X1 U6173 ( .B1(n8507), .B2(n4670), .A(n4668), .ZN(n8512) );
  OR2_X1 U6174 ( .A1(n4534), .A2(n6950), .ZN(n4533) );
  AND2_X1 U6175 ( .A1(n7073), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n4534) );
  OR2_X1 U6176 ( .A1(n5781), .A2(n6976), .ZN(n4535) );
  AND3_X1 U6177 ( .A1(n8439), .A2(n8453), .A3(n8433), .ZN(n4536) );
  OR2_X1 U6178 ( .A1(n5792), .A2(P2_IR_REG_26__SCAN_IN), .ZN(n4537) );
  OR2_X1 U6179 ( .A1(n5241), .A2(SI_11_), .ZN(n4538) );
  INV_X1 U6180 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n5181) );
  XNOR2_X1 U6181 ( .A(n8590), .B(n8902), .ZN(n8581) );
  INV_X1 U6182 ( .A(n9018), .ZN(n4721) );
  INV_X1 U6183 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n9159) );
  NAND2_X1 U6184 ( .A1(n6139), .A2(n6138), .ZN(n7765) );
  AND2_X1 U6185 ( .A1(n6947), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n4539) );
  AND2_X1 U6186 ( .A1(n7850), .A2(n8737), .ZN(n4540) );
  OR2_X1 U6187 ( .A1(n5477), .A2(n5476), .ZN(n8737) );
  NAND2_X1 U6188 ( .A1(n8660), .A2(n4962), .ZN(n8604) );
  AND2_X1 U6189 ( .A1(n9275), .A2(n6292), .ZN(n4541) );
  AND4_X1 U6190 ( .A1(n5829), .A2(n5830), .A3(n5828), .A4(n5838), .ZN(n4542)
         );
  AND2_X1 U6191 ( .A1(n9815), .A2(n9406), .ZN(n4543) );
  AND2_X1 U6192 ( .A1(n5635), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n4544) );
  AND2_X1 U6193 ( .A1(n4806), .A2(n4804), .ZN(n4545) );
  NAND2_X1 U6194 ( .A1(n9067), .A2(n8981), .ZN(n4546) );
  AND2_X1 U6195 ( .A1(n4733), .A2(n4732), .ZN(n4547) );
  INV_X1 U6196 ( .A(n8193), .ZN(n4710) );
  INV_X1 U6197 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n5617) );
  NAND2_X1 U6198 ( .A1(n5907), .A2(n4730), .ZN(n6785) );
  NAND2_X1 U6199 ( .A1(n9214), .A2(n6620), .ZN(n4797) );
  XNOR2_X1 U6200 ( .A(n9095), .B(n8587), .ZN(n8897) );
  NAND2_X1 U6201 ( .A1(n5839), .A2(n5142), .ZN(n5851) );
  AOI21_X1 U6202 ( .B1(n9635), .B2(n4628), .A(n4626), .ZN(n4625) );
  INV_X1 U6203 ( .A(n5729), .ZN(n4889) );
  NAND2_X1 U6204 ( .A1(n7947), .A2(n8735), .ZN(n4548) );
  NAND2_X1 U6205 ( .A1(n6294), .A2(n6293), .ZN(n9815) );
  INV_X1 U6206 ( .A(n4770), .ZN(n9590) );
  NOR2_X1 U6207 ( .A1(n9607), .A2(n9591), .ZN(n4770) );
  AND2_X1 U6208 ( .A1(n6491), .A2(n6490), .ZN(n9526) );
  INV_X1 U6209 ( .A(n9526), .ZN(n4648) );
  AND2_X1 U6210 ( .A1(n4974), .A2(n8672), .ZN(n4549) );
  INV_X1 U6211 ( .A(n9739), .ZN(n6494) );
  AND2_X1 U6212 ( .A1(n7444), .A2(n7442), .ZN(n4550) );
  AND2_X1 U6213 ( .A1(n9556), .A2(n9541), .ZN(n4551) );
  OR2_X1 U6214 ( .A1(n8561), .A2(n8982), .ZN(n4552) );
  OR2_X1 U6215 ( .A1(n7947), .A2(n7959), .ZN(n8057) );
  INV_X1 U6216 ( .A(n4632), .ZN(n8358) );
  INV_X1 U6217 ( .A(n4983), .ZN(n4980) );
  NAND2_X1 U6218 ( .A1(n4984), .A2(n7845), .ZN(n4983) );
  AND2_X1 U6219 ( .A1(n4525), .A2(n4973), .ZN(n4553) );
  AND2_X1 U6220 ( .A1(n4921), .A2(n4919), .ZN(n4554) );
  NOR2_X1 U6221 ( .A1(n9941), .A2(n9417), .ZN(n4555) );
  NOR2_X1 U6222 ( .A1(n8628), .A2(n8935), .ZN(n4556) );
  NOR2_X1 U6223 ( .A1(n9800), .A2(n9403), .ZN(n4557) );
  OR2_X1 U6224 ( .A1(n9137), .A2(n8995), .ZN(n5762) );
  INV_X1 U6225 ( .A(n6586), .ZN(n4659) );
  AND2_X1 U6226 ( .A1(n5108), .A2(n4677), .ZN(n4558) );
  NOR2_X1 U6227 ( .A1(n8006), .A2(n8733), .ZN(n4559) );
  AND2_X1 U6228 ( .A1(n4637), .A2(n7149), .ZN(n4560) );
  AND2_X1 U6229 ( .A1(n4518), .A2(n5729), .ZN(n4561) );
  XNOR2_X1 U6230 ( .A(n5913), .B(n4512), .ZN(n5933) );
  AND2_X1 U6231 ( .A1(n4774), .A2(n7926), .ZN(n4562) );
  NAND2_X1 U6232 ( .A1(n4739), .A2(n5205), .ZN(n4563) );
  INV_X1 U6233 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n5599) );
  INV_X1 U6234 ( .A(n4920), .ZN(n4919) );
  NAND2_X1 U6235 ( .A1(n8178), .A2(n5690), .ZN(n4920) );
  NAND2_X1 U6236 ( .A1(n8574), .A2(n8713), .ZN(n8716) );
  INV_X1 U6237 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n5488) );
  AND2_X1 U6238 ( .A1(n5837), .A2(n5862), .ZN(n4564) );
  AND2_X1 U6239 ( .A1(n6329), .A2(n6328), .ZN(n4565) );
  INV_X1 U6240 ( .A(n8464), .ZN(n7657) );
  AND2_X1 U6241 ( .A1(n8370), .A2(n8368), .ZN(n8464) );
  AND2_X1 U6242 ( .A1(n8175), .A2(n8176), .ZN(n8922) );
  AND2_X1 U6243 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n4566) );
  OR2_X1 U6244 ( .A1(n9089), .A2(n8191), .ZN(n4567) );
  OR2_X1 U6245 ( .A1(n8510), .A2(n8509), .ZN(n4568) );
  NOR2_X1 U6246 ( .A1(P2_IR_REG_28__SCAN_IN), .A2(P2_IR_REG_29__SCAN_IN), .ZN(
        n4569) );
  AND2_X1 U6247 ( .A1(n5033), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4570) );
  NAND4_X1 U6248 ( .A1(n4521), .A2(n5000), .A3(n5834), .A4(n4999), .ZN(n4571)
         );
  INV_X1 U6249 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n5033) );
  AND2_X1 U6250 ( .A1(n5840), .A2(n5872), .ZN(n4572) );
  INV_X1 U6251 ( .A(n8129), .ZN(n5116) );
  INV_X1 U6252 ( .A(n7156), .ZN(n7149) );
  AND2_X1 U6253 ( .A1(n5425), .A2(n5436), .ZN(n7156) );
  AND2_X1 U6254 ( .A1(n4996), .A2(n4995), .ZN(n4573) );
  NOR2_X1 U6255 ( .A1(n8824), .A2(n8823), .ZN(n4574) );
  AND2_X1 U6256 ( .A1(n8078), .A2(n8077), .ZN(n4575) );
  INV_X1 U6257 ( .A(n5450), .ZN(n4902) );
  AND2_X1 U6258 ( .A1(n5181), .A2(n5083), .ZN(n4576) );
  AND2_X1 U6259 ( .A1(n8577), .A2(n8576), .ZN(n4577) );
  NAND2_X1 U6260 ( .A1(n6204), .A2(n6203), .ZN(n10073) );
  OR2_X1 U6261 ( .A1(n7630), .A2(n7621), .ZN(n8114) );
  INV_X1 U6262 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n10441) );
  AND2_X1 U6263 ( .A1(n4524), .A2(n5840), .ZN(n4578) );
  NAND2_X1 U6264 ( .A1(n8184), .A2(n4889), .ZN(n4579) );
  INV_X1 U6265 ( .A(n4908), .ZN(n4907) );
  NAND2_X1 U6266 ( .A1(n4913), .A2(n4910), .ZN(n4908) );
  AND2_X1 U6267 ( .A1(n4648), .A2(n8495), .ZN(n8508) );
  XNOR2_X1 U6268 ( .A(n5391), .B(n5390), .ZN(n6950) );
  NAND2_X1 U6269 ( .A1(n7900), .A2(n8238), .ZN(n7969) );
  AND2_X1 U6270 ( .A1(n6368), .A2(n6367), .ZN(n9256) );
  INV_X1 U6271 ( .A(n9256), .ZN(n4749) );
  INV_X1 U6272 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n4795) );
  AOI21_X1 U6273 ( .B1(n7969), .B2(n5550), .A(n4516), .ZN(n7990) );
  INV_X1 U6274 ( .A(n7382), .ZN(n7577) );
  INV_X1 U6275 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n6158) );
  INV_X1 U6276 ( .A(n8968), .ZN(n4892) );
  NAND2_X1 U6277 ( .A1(n5715), .A2(n5714), .ZN(n8901) );
  NAND2_X1 U6278 ( .A1(n6496), .A2(n6495), .ZN(n9770) );
  INV_X1 U6279 ( .A(n9770), .ZN(n9570) );
  NOR2_X1 U6280 ( .A1(n9832), .A2(n9833), .ZN(n9736) );
  AND2_X1 U6281 ( .A1(n5120), .A2(n6133), .ZN(n4580) );
  NAND2_X1 U6282 ( .A1(n4684), .A2(n4683), .ZN(n7789) );
  NOR2_X1 U6283 ( .A1(n10103), .A2(n8746), .ZN(n4581) );
  NAND2_X1 U6284 ( .A1(n4515), .A2(n4768), .ZN(n4769) );
  NAND2_X1 U6285 ( .A1(n9791), .A2(n9402), .ZN(n4582) );
  AND2_X1 U6286 ( .A1(n4810), .A2(n6223), .ZN(n4583) );
  AND2_X1 U6287 ( .A1(n9800), .A2(n9403), .ZN(n4584) );
  NOR2_X1 U6288 ( .A1(P1_IR_REG_14__SCAN_IN), .A2(P1_IR_REG_15__SCAN_IN), .ZN(
        n6248) );
  AND2_X1 U6289 ( .A1(n5271), .A2(SI_21_), .ZN(n4585) );
  OR2_X1 U6290 ( .A1(n9591), .A2(n9400), .ZN(n4586) );
  NOR2_X1 U6291 ( .A1(n5063), .A2(n5061), .ZN(n4587) );
  NOR2_X1 U6292 ( .A1(n5272), .A2(n5037), .ZN(n5036) );
  AND2_X1 U6293 ( .A1(n7820), .A2(n8385), .ZN(n4588) );
  INV_X1 U6294 ( .A(SI_15_), .ZN(n5061) );
  NAND2_X1 U6295 ( .A1(n6184), .A2(n6183), .ZN(n7873) );
  INV_X1 U6296 ( .A(n7873), .ZN(n4762) );
  NAND2_X1 U6297 ( .A1(n5886), .A2(n5885), .ZN(n9688) );
  INV_X1 U6298 ( .A(n9688), .ZN(n4765) );
  INV_X1 U6299 ( .A(n9483), .ZN(n4737) );
  NAND2_X1 U6300 ( .A1(n7652), .A2(n9358), .ZN(n7745) );
  OAI21_X1 U6301 ( .B1(n7254), .B2(n6586), .A(n8297), .ZN(n8294) );
  NAND2_X1 U6302 ( .A1(n4965), .A2(n6668), .ZN(n6833) );
  XNOR2_X1 U6303 ( .A(n4985), .B(n8737), .ZN(n7851) );
  INV_X1 U6304 ( .A(n8764), .ZN(n10135) );
  OAI22_X1 U6305 ( .A1(n7856), .A2(n4675), .B1(n4558), .B2(n5107), .ZN(n8030)
         );
  NAND2_X1 U6306 ( .A1(n7443), .A2(n4550), .ZN(n7543) );
  NAND2_X1 U6307 ( .A1(n5981), .A2(n5980), .ZN(n7345) );
  XNOR2_X1 U6308 ( .A(n6094), .B(n6092), .ZN(n9939) );
  OAI21_X1 U6309 ( .B1(n7515), .B2(n6042), .A(n6041), .ZN(n7556) );
  AND2_X1 U6310 ( .A1(n8308), .A2(n6597), .ZN(n4589) );
  NAND2_X1 U6311 ( .A1(n7652), .A2(n4520), .ZN(n4764) );
  OR2_X1 U6312 ( .A1(n7699), .A2(n7687), .ZN(n4590) );
  AND2_X1 U6313 ( .A1(n5733), .A2(n10359), .ZN(n4591) );
  AND2_X1 U6314 ( .A1(n7335), .A2(n7339), .ZN(n7366) );
  AND2_X1 U6315 ( .A1(n4876), .A2(n4875), .ZN(n4592) );
  NAND2_X1 U6316 ( .A1(n4947), .A2(n6950), .ZN(n7164) );
  INV_X1 U6317 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n6429) );
  AND2_X1 U6318 ( .A1(n8872), .A2(n8841), .ZN(n4593) );
  NAND2_X1 U6319 ( .A1(n5981), .A2(n4812), .ZN(n7347) );
  INV_X1 U6320 ( .A(n8823), .ZN(n4945) );
  AND2_X1 U6321 ( .A1(n4858), .A2(n4866), .ZN(n4594) );
  NAND2_X1 U6322 ( .A1(n7116), .A2(n4966), .ZN(n7246) );
  OR2_X1 U6323 ( .A1(n8809), .A2(n4593), .ZN(n4595) );
  AND2_X1 U6324 ( .A1(n4859), .A2(n4862), .ZN(n4596) );
  INV_X1 U6325 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n4731) );
  INV_X1 U6326 ( .A(n7172), .ZN(n4850) );
  XNOR2_X1 U6327 ( .A(n5864), .B(P1_IR_REG_20__SCAN_IN), .ZN(n8504) );
  INV_X1 U6328 ( .A(n8504), .ZN(n7528) );
  INV_X1 U6329 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n4695) );
  OAI21_X1 U6330 ( .B1(n7061), .B2(n4534), .A(n6950), .ZN(n4868) );
  NOR2_X1 U6331 ( .A1(n4957), .A2(n6950), .ZN(n4956) );
  INV_X1 U6332 ( .A(n6950), .ZN(n4950) );
  NOR2_X1 U6333 ( .A1(n6950), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n4952) );
  NAND2_X1 U6334 ( .A1(n5613), .A2(n5612), .ZN(n8992) );
  OAI21_X2 U6336 ( .B1(n5677), .B2(n4920), .A(n4917), .ZN(n8913) );
  NAND2_X1 U6337 ( .A1(n4893), .A2(n4891), .ZN(n8952) );
  NAND2_X1 U6338 ( .A1(n9023), .A2(n5596), .ZN(n9002) );
  INV_X1 U6339 ( .A(n9041), .ZN(n4602) );
  OAI21_X1 U6340 ( .B1(n7792), .B2(n5502), .A(n5503), .ZN(n7857) );
  NAND2_X1 U6341 ( .A1(n5595), .A2(n9018), .ZN(n9023) );
  NAND2_X1 U6342 ( .A1(n4674), .A2(n4527), .ZN(n9158) );
  NAND2_X1 U6343 ( .A1(n8957), .A2(n5660), .ZN(n8944) );
  NAND2_X1 U6344 ( .A1(n5180), .A2(n5389), .ZN(n5570) );
  NAND2_X1 U6345 ( .A1(n10144), .A2(n5345), .ZN(n7279) );
  OAI21_X1 U6346 ( .B1(n7772), .B2(n5478), .A(n4598), .ZN(n7792) );
  NAND2_X1 U6347 ( .A1(n9168), .A2(n8538), .ZN(n7530) );
  XNOR2_X2 U6348 ( .A(n5191), .B(P2_IR_REG_29__SCAN_IN), .ZN(n9168) );
  NAND2_X1 U6349 ( .A1(n10145), .A2(n10146), .ZN(n10144) );
  NOR2_X1 U6350 ( .A1(n4600), .A2(n4544), .ZN(n4599) );
  AOI21_X1 U6351 ( .B1(n8913), .B2(n5717), .A(n5716), .ZN(n8898) );
  AOI21_X2 U6352 ( .B1(n7942), .B2(n8736), .A(n7941), .ZN(n7944) );
  XNOR2_X1 U6353 ( .A(n6880), .B(n6841), .ZN(n6878) );
  XNOR2_X2 U6354 ( .A(n8743), .B(n10143), .ZN(n10146) );
  NAND2_X2 U6355 ( .A1(n4599), .A2(n5334), .ZN(n8743) );
  NAND2_X1 U6356 ( .A1(n5070), .A2(n6839), .ZN(n8058) );
  INV_X1 U6357 ( .A(n7857), .ZN(n5518) );
  AND2_X2 U6358 ( .A1(n5192), .A2(n9168), .ZN(n5635) );
  NAND2_X1 U6359 ( .A1(n5333), .A2(n5335), .ZN(n4600) );
  NAND2_X1 U6360 ( .A1(n5465), .A2(n5464), .ZN(n7772) );
  NAND2_X1 U6361 ( .A1(n9263), .A2(n9267), .ZN(n9276) );
  NAND2_X1 U6362 ( .A1(n4988), .A2(n4986), .ZN(n8700) );
  NAND3_X1 U6363 ( .A1(n4965), .A2(n5818), .A3(n4964), .ZN(n4963) );
  AOI21_X1 U6364 ( .B1(n7298), .B2(n7297), .A(n7296), .ZN(n7300) );
  AND2_X1 U6365 ( .A1(n5995), .A2(n5980), .ZN(n4812) );
  NAND2_X2 U6366 ( .A1(n6841), .A2(n7431), .ZN(n8066) );
  NAND2_X1 U6367 ( .A1(n4924), .A2(n5366), .ZN(n7266) );
  OAI21_X1 U6368 ( .B1(n8535), .B2(n4509), .A(n4726), .ZN(P1_U3262) );
  NAND2_X1 U6369 ( .A1(n8534), .A2(n9517), .ZN(n4729) );
  OAI211_X1 U6370 ( .C1(n8533), .C2(n9510), .A(n4729), .B(n7885), .ZN(n4728)
         );
  NAND2_X2 U6371 ( .A1(n8944), .A2(n5675), .ZN(n5677) );
  NAND2_X1 U6372 ( .A1(n7279), .A2(n5365), .ZN(n4924) );
  OAI21_X1 U6373 ( .B1(n7969), .B2(n4908), .A(n4904), .ZN(n5595) );
  AND2_X1 U6374 ( .A1(n4612), .A2(n4613), .ZN(n4609) );
  NAND2_X1 U6375 ( .A1(n4611), .A2(n4608), .ZN(n4610) );
  NAND2_X1 U6376 ( .A1(n4610), .A2(n4615), .ZN(n6618) );
  NAND2_X1 U6377 ( .A1(n10082), .A2(n4616), .ZN(n4615) );
  INV_X1 U6378 ( .A(n4625), .ZN(n9571) );
  NAND2_X1 U6379 ( .A1(n7805), .A2(n6600), .ZN(n6601) );
  INV_X2 U6380 ( .A(n5225), .ZN(n6672) );
  MUX2_X1 U6381 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(P1_DATAO_REG_7__SCAN_IN), 
        .S(n5225), .Z(n4634) );
  NAND2_X1 U6382 ( .A1(n7168), .A2(n4639), .ZN(n4640) );
  NAND3_X1 U6383 ( .A1(n4640), .A2(n7193), .A3(P2_REG2_REG_7__SCAN_IN), .ZN(
        n7197) );
  OAI21_X1 U6384 ( .B1(n4644), .B2(n10104), .A(n4643), .ZN(n10119) );
  NAND2_X1 U6385 ( .A1(n8746), .A2(n4645), .ZN(n4643) );
  INV_X1 U6386 ( .A(n10120), .ZN(n4645) );
  NAND2_X1 U6387 ( .A1(n6944), .A2(n5359), .ZN(n4646) );
  NOR2_X2 U6388 ( .A1(n4650), .A2(n8443), .ZN(n8452) );
  OAI21_X1 U6389 ( .B1(n4838), .B2(n8437), .A(n4837), .ZN(n4652) );
  NAND3_X1 U6390 ( .A1(n4656), .A2(n8299), .A3(n4655), .ZN(n8345) );
  NAND2_X1 U6391 ( .A1(n8361), .A2(n8360), .ZN(n8367) );
  OAI21_X1 U6392 ( .B1(n8361), .B2(n8358), .A(n4660), .ZN(n4663) );
  OAI21_X1 U6393 ( .B1(n8360), .B2(n8358), .A(n8368), .ZN(n4661) );
  NAND2_X1 U6394 ( .A1(n4663), .A2(n4662), .ZN(n8375) );
  NAND2_X1 U6395 ( .A1(n4665), .A2(n8419), .ZN(n4664) );
  NAND3_X1 U6396 ( .A1(n4667), .A2(n4821), .A3(n4666), .ZN(n4665) );
  NAND2_X1 U6397 ( .A1(n8415), .A2(n8453), .ZN(n4666) );
  NAND2_X1 U6398 ( .A1(n8416), .A2(n8444), .ZN(n4667) );
  NAND3_X1 U6399 ( .A1(n4840), .A2(n4751), .A3(n5145), .ZN(n8507) );
  AND2_X1 U6400 ( .A1(n4672), .A2(n4822), .ZN(n4671) );
  NAND2_X2 U6401 ( .A1(n5084), .A2(n5082), .ZN(n5792) );
  NAND2_X1 U6402 ( .A1(n8030), .A2(n8242), .ZN(n8031) );
  INV_X1 U6403 ( .A(n5107), .ZN(n4679) );
  NAND2_X1 U6404 ( .A1(n4680), .A2(n4681), .ZN(n5760) );
  NAND2_X1 U6405 ( .A1(n7618), .A2(n4683), .ZN(n4680) );
  OAI21_X2 U6406 ( .B1(n8895), .B2(n10137), .A(n4694), .ZN(n8889) );
  NAND3_X1 U6407 ( .A1(n8869), .A2(n4696), .A3(n4695), .ZN(n4747) );
  MUX2_X1 U6408 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(P2_DATAO_REG_3__SCAN_IN), 
        .S(n5217), .Z(n5214) );
  NAND2_X2 U6409 ( .A1(n5237), .A2(n5059), .ZN(n5469) );
  NOR2_X2 U6410 ( .A1(n8194), .A2(n4709), .ZN(n8188) );
  NAND3_X1 U6411 ( .A1(n8136), .A2(n8141), .A3(n8203), .ZN(n4722) );
  MUX2_X1 U6412 ( .A(n10085), .B(P1_REG1_REG_1__SCAN_IN), .S(n6785), .Z(n9424)
         );
  NAND3_X1 U6413 ( .A1(n4739), .A2(n5205), .A3(n5212), .ZN(n5338) );
  MUX2_X1 U6414 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .S(n5217), .Z(n5325) );
  NAND3_X1 U6415 ( .A1(n5200), .A2(P1_ADDR_REG_19__SCAN_IN), .A3(
        P2_ADDR_REG_19__SCAN_IN), .ZN(n4746) );
  NAND2_X1 U6416 ( .A1(n5586), .A2(n4755), .ZN(n4754) );
  NAND2_X1 U6417 ( .A1(n5586), .A2(n5046), .ZN(n5043) );
  NOR2_X2 U6418 ( .A1(n7418), .A2(n7475), .ZN(n9976) );
  INV_X1 U6419 ( .A(n4764), .ZN(n9753) );
  NAND3_X2 U6420 ( .A1(n4515), .A2(n4765), .A3(n4766), .ZN(n9686) );
  INV_X1 U6421 ( .A(n4769), .ZN(n9718) );
  NAND2_X1 U6422 ( .A1(n6604), .A2(n4780), .ZN(n4777) );
  NAND2_X1 U6423 ( .A1(n4777), .A2(n4778), .ZN(n9534) );
  NAND2_X1 U6424 ( .A1(n6604), .A2(n9574), .ZN(n9573) );
  NAND2_X1 U6425 ( .A1(n5469), .A2(n4787), .ZN(n4791) );
  NAND2_X1 U6426 ( .A1(n5469), .A2(n5240), .ZN(n5480) );
  NAND2_X1 U6427 ( .A1(n6602), .A2(n4792), .ZN(n9730) );
  NAND2_X1 U6428 ( .A1(n4794), .A2(n9728), .ZN(n9729) );
  NAND2_X1 U6429 ( .A1(n4797), .A2(n6524), .ZN(n5911) );
  INV_X1 U6430 ( .A(n4797), .ZN(n6619) );
  NAND2_X1 U6431 ( .A1(n4797), .A2(n7110), .ZN(n5923) );
  NAND2_X1 U6432 ( .A1(n4797), .A2(n7257), .ZN(n5951) );
  NAND2_X2 U6433 ( .A1(n4800), .A2(n4798), .ZN(n9285) );
  NAND3_X1 U6434 ( .A1(n5127), .A2(n9265), .A3(n9388), .ZN(n9263) );
  NAND2_X1 U6435 ( .A1(n6130), .A2(n9346), .ZN(n9908) );
  NAND2_X1 U6436 ( .A1(n9299), .A2(n4808), .ZN(n9346) );
  NAND2_X1 U6437 ( .A1(n9299), .A2(n6113), .ZN(n6129) );
  NAND2_X1 U6438 ( .A1(n4811), .A2(n6223), .ZN(n6244) );
  NAND2_X1 U6439 ( .A1(n7347), .A2(n5998), .ZN(n7515) );
  NAND4_X1 U6440 ( .A1(n5835), .A2(n5834), .A3(n5836), .A4(n6008), .ZN(n5861)
         );
  AND2_X2 U6441 ( .A1(n6768), .A2(n6671), .ZN(n5910) );
  NAND2_X1 U6442 ( .A1(n4825), .A2(n4826), .ZN(n5842) );
  NAND2_X1 U6443 ( .A1(n5847), .A2(n4827), .ZN(n4825) );
  NAND2_X1 U6444 ( .A1(n4843), .A2(n8353), .ZN(n8361) );
  NAND3_X1 U6445 ( .A1(n8347), .A2(n8453), .A3(n8346), .ZN(n4846) );
  NAND2_X1 U6446 ( .A1(n6585), .A2(n6584), .ZN(n7254) );
  NAND2_X1 U6447 ( .A1(n7145), .A2(n4530), .ZN(n4851) );
  OAI211_X1 U6448 ( .C1(n7145), .C2(n4852), .A(n4851), .B(n4847), .ZN(n7211)
         );
  NAND3_X1 U6449 ( .A1(n4866), .A2(n4861), .A3(n4860), .ZN(n7174) );
  NAND2_X1 U6450 ( .A1(n6937), .A2(n7061), .ZN(n7066) );
  OR2_X1 U6451 ( .A1(n6937), .A2(n4534), .ZN(n4864) );
  NAND2_X1 U6452 ( .A1(n6937), .A2(n4867), .ZN(n4866) );
  INV_X1 U6453 ( .A(n4876), .ZN(n7681) );
  INV_X1 U6454 ( .A(n7682), .ZN(n4875) );
  NAND2_X1 U6455 ( .A1(n4879), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n4878) );
  INV_X1 U6456 ( .A(n7366), .ZN(n4877) );
  NAND2_X1 U6457 ( .A1(n6908), .A2(n4997), .ZN(n6585) );
  NOR2_X1 U6458 ( .A1(n10110), .A2(n10109), .ZN(n10108) );
  NOR2_X1 U6459 ( .A1(n8854), .A2(n8853), .ZN(n8856) );
  NAND2_X1 U6460 ( .A1(n6960), .A2(n6935), .ZN(n6936) );
  NAND3_X1 U6461 ( .A1(n4883), .A2(n4881), .A3(n10151), .ZN(n5784) );
  NAND2_X1 U6463 ( .A1(n8992), .A2(n4894), .ZN(n4893) );
  INV_X1 U6464 ( .A(n7632), .ZN(n4903) );
  NAND2_X1 U6465 ( .A1(n4899), .A2(n4900), .ZN(n5465) );
  NAND2_X1 U6466 ( .A1(n7632), .A2(n5450), .ZN(n4899) );
  INV_X1 U6467 ( .A(n4914), .ZN(n5187) );
  AND2_X1 U6468 ( .A1(n4926), .A2(n7239), .ZN(n4925) );
  OAI21_X1 U6469 ( .B1(n6991), .B2(n6945), .A(n6946), .ZN(n4926) );
  INV_X1 U6470 ( .A(n4935), .ZN(n4934) );
  OAI21_X1 U6471 ( .B1(n6965), .B2(n4539), .A(n6976), .ZN(n4935) );
  NOR2_X1 U6472 ( .A1(n8820), .A2(n8821), .ZN(n8824) );
  OAI211_X1 U6473 ( .C1(n4943), .C2(n8820), .A(n4939), .B(n4938), .ZN(n8877)
         );
  NAND3_X1 U6474 ( .A1(n8820), .A2(n4945), .A3(n4946), .ZN(n4938) );
  NAND2_X1 U6475 ( .A1(n7164), .A2(n4955), .ZN(n6951) );
  MUX2_X1 U6476 ( .A(n9174), .B(P2_IR_REG_0__SCAN_IN), .S(P2_STATE_REG_SCAN_IN), .Z(P2_U3295) );
  MUX2_X1 U6477 ( .A(P2_IR_REG_0__SCAN_IN), .B(n9174), .S(n5781), .Z(n6839) );
  NAND2_X1 U6478 ( .A1(n7319), .A2(n7339), .ZN(n7318) );
  NAND3_X1 U6479 ( .A1(n4962), .A2(n8660), .A3(n8694), .ZN(n8605) );
  NAND2_X2 U6480 ( .A1(n8565), .A2(n8564), .ZN(n8660) );
  NAND2_X1 U6481 ( .A1(n8563), .A2(n8562), .ZN(n4962) );
  CLKBUF_X1 U6482 ( .A(n4968), .Z(n4967) );
  NAND2_X1 U6483 ( .A1(n8716), .A2(n8576), .ZN(n8594) );
  NAND2_X1 U6484 ( .A1(n8716), .A2(n4577), .ZN(n8596) );
  NAND2_X1 U6485 ( .A1(n8642), .A2(n4989), .ZN(n4988) );
  NAND2_X1 U6486 ( .A1(n5572), .A2(n4996), .ZN(n5746) );
  NAND2_X1 U6487 ( .A1(n5572), .A2(n5599), .ZN(n5742) );
  INV_X1 U6488 ( .A(n4997), .ZN(n6523) );
  XNOR2_X1 U6489 ( .A(n9981), .B(n4997), .ZN(n9983) );
  XNOR2_X1 U6490 ( .A(n9980), .B(n4997), .ZN(n10007) );
  NAND4_X1 U6491 ( .A1(n8462), .A2(n8463), .A3(n8464), .A4(n4997), .ZN(n8467)
         );
  NAND2_X1 U6492 ( .A1(n9961), .A2(n5004), .ZN(n5002) );
  OAI21_X2 U6493 ( .B1(n7752), .B2(n6543), .A(n6544), .ZN(n7812) );
  OR2_X1 U6494 ( .A1(n10073), .A2(n9411), .ZN(n5012) );
  NAND2_X1 U6495 ( .A1(n9565), .A2(n4517), .ZN(n5014) );
  OR2_X1 U6496 ( .A1(n9565), .A2(n9574), .ZN(n5016) );
  NAND2_X1 U6497 ( .A1(n9616), .A2(n5021), .ZN(n5018) );
  OAI21_X1 U6498 ( .B1(n9663), .B2(n6559), .A(n6560), .ZN(n9648) );
  OAI21_X1 U6499 ( .B1(n9711), .B2(n6555), .A(n6556), .ZN(n9695) );
  AND2_X1 U6500 ( .A1(n5847), .A2(n4578), .ZN(n5871) );
  NAND2_X1 U6501 ( .A1(n5847), .A2(n5032), .ZN(n9896) );
  INV_X1 U6502 ( .A(n5651), .ZN(n5277) );
  NAND2_X1 U6503 ( .A1(n5661), .A2(n5051), .ZN(n5048) );
  NAND2_X1 U6504 ( .A1(n5048), .A2(n5049), .ZN(n5692) );
  NAND2_X1 U6505 ( .A1(n5661), .A2(n5284), .ZN(n5664) );
  NAND2_X1 U6506 ( .A1(n5306), .A2(n5056), .ZN(n5055) );
  NAND2_X1 U6507 ( .A1(n5306), .A2(n5305), .ZN(n5719) );
  NAND2_X1 U6508 ( .A1(n5062), .A2(n4587), .ZN(n5250) );
  NAND3_X1 U6509 ( .A1(n5192), .A2(n9169), .A3(P2_REG2_REG_1__SCAN_IN), .ZN(
        n5067) );
  NAND2_X1 U6510 ( .A1(n8988), .A2(n5068), .ZN(n8964) );
  NAND2_X1 U6511 ( .A1(n8964), .A2(n8052), .ZN(n5763) );
  NAND2_X1 U6512 ( .A1(n7011), .A2(n10147), .ZN(n8061) );
  NAND2_X1 U6513 ( .A1(n8066), .A2(n8061), .ZN(n7005) );
  NAND3_X1 U6514 ( .A1(n5751), .A2(n8066), .A3(n8061), .ZN(n7006) );
  INV_X1 U6515 ( .A(n5317), .ZN(n5070) );
  INV_X1 U6516 ( .A(n6839), .ZN(n5071) );
  NAND2_X1 U6517 ( .A1(n7270), .A2(n4575), .ZN(n5758) );
  XNOR2_X1 U6518 ( .A(n5073), .B(n5072), .ZN(n7439) );
  NAND2_X1 U6519 ( .A1(n5075), .A2(n5074), .ZN(n5767) );
  OAI21_X1 U6520 ( .B1(n9019), .B2(n5078), .A(n5076), .ZN(n8990) );
  INV_X1 U6521 ( .A(n5570), .ZN(n5084) );
  NOR2_X1 U6522 ( .A1(n5570), .A2(P2_IR_REG_16__SCAN_IN), .ZN(n5572) );
  NAND2_X1 U6523 ( .A1(n8213), .A2(n5089), .ZN(n5087) );
  NAND2_X1 U6524 ( .A1(n5087), .A2(n5088), .ZN(n8261) );
  NAND2_X1 U6525 ( .A1(n9908), .A2(n9346), .ZN(n5118) );
  INV_X1 U6526 ( .A(n9909), .ZN(n5120) );
  NAND2_X1 U6527 ( .A1(n5118), .A2(n5117), .ZN(n9238) );
  AOI21_X1 U6528 ( .B1(n9346), .B2(n9910), .A(n5119), .ZN(n5117) );
  AOI21_X1 U6529 ( .B1(n9285), .B2(n5123), .A(n5121), .ZN(n9218) );
  NAND2_X1 U6530 ( .A1(n9285), .A2(n6376), .ZN(n9252) );
  NAND2_X1 U6531 ( .A1(n9387), .A2(n9390), .ZN(n5127) );
  NAND3_X1 U6532 ( .A1(n5835), .A2(n5834), .A3(n6008), .ZN(n6273) );
  NAND2_X1 U6533 ( .A1(n6500), .A2(n6485), .ZN(n6489) );
  INV_X1 U6534 ( .A(n5661), .ZN(n5663) );
  OAI21_X1 U6535 ( .B1(n6458), .B2(n9003), .A(n6457), .ZN(n9088) );
  INV_X4 U6536 ( .A(n5225), .ZN(n6671) );
  MUX2_X1 U6537 ( .A(n8442), .B(n8441), .S(n8444), .Z(n8443) );
  NOR2_X1 U6538 ( .A1(n7944), .A2(n7943), .ZN(n7952) );
  AND2_X1 U6539 ( .A1(n9852), .A2(n9399), .ZN(n8441) );
  NAND2_X1 U6540 ( .A1(n8451), .A2(n8444), .ZN(n8447) );
  NOR2_X1 U6541 ( .A1(n9545), .A2(n8451), .ZN(n6503) );
  OAI21_X1 U6542 ( .B1(n5217), .B2(n5207), .A(n5206), .ZN(n5208) );
  NAND2_X1 U6543 ( .A1(n5217), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n5206) );
  MUX2_X2 U6544 ( .A(n6646), .B(n6645), .S(n10213), .Z(n6649) );
  NOR2_X2 U6545 ( .A1(n8889), .A2(n5786), .ZN(n6645) );
  NAND2_X1 U6546 ( .A1(n9542), .A2(n6580), .ZN(n9554) );
  OAI21_X1 U6547 ( .B1(n9218), .B2(n6632), .A(n9948), .ZN(n6641) );
  NAND2_X1 U6548 ( .A1(n5187), .A2(P2_IR_REG_30__SCAN_IN), .ZN(n5189) );
  NAND2_X1 U6549 ( .A1(n5856), .A2(n5855), .ZN(n7919) );
  NAND2_X1 U6550 ( .A1(n5856), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5850) );
  NOR2_X1 U6551 ( .A1(n5931), .A2(n4512), .ZN(n5932) );
  NAND2_X1 U6552 ( .A1(n5926), .A2(n5138), .ZN(n6894) );
  NAND2_X1 U6553 ( .A1(n5925), .A2(n5883), .ZN(n5905) );
  AOI21_X2 U6554 ( .B1(n8700), .B2(n8612), .A(n8611), .ZN(n8674) );
  OR2_X1 U6555 ( .A1(n10159), .A2(n6469), .ZN(n9035) );
  INV_X2 U6556 ( .A(n10201), .ZN(n10199) );
  OAI21_X1 U6557 ( .B1(n7591), .B2(n7592), .A(n7593), .ZN(n7546) );
  INV_X1 U6558 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n5153) );
  OR2_X1 U6559 ( .A1(n9029), .A2(n6471), .ZN(n5137) );
  OR2_X1 U6560 ( .A1(n5925), .A2(n9954), .ZN(n5138) );
  AND2_X1 U6561 ( .A1(n7951), .A2(n8735), .ZN(n5140) );
  AND2_X1 U6562 ( .A1(n5517), .A2(n7959), .ZN(n5141) );
  AND3_X1 U6563 ( .A1(n5858), .A2(n6432), .A3(n6429), .ZN(n5142) );
  INV_X1 U6564 ( .A(n9025), .ZN(n9006) );
  NAND2_X1 U6565 ( .A1(n9377), .A2(n6035), .ZN(n5143) );
  NAND2_X1 U6566 ( .A1(n5674), .A2(n5673), .ZN(n8958) );
  INV_X1 U6567 ( .A(n9076), .ZN(n6647) );
  INV_X1 U6568 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n5849) );
  INV_X1 U6569 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n5872) );
  INV_X1 U6570 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n5155) );
  INV_X1 U6571 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n6067) );
  AND2_X1 U6572 ( .A1(n4673), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n5144) );
  NAND2_X1 U6573 ( .A1(n8450), .A2(n8449), .ZN(n5145) );
  OR2_X1 U6574 ( .A1(n9526), .A2(n9891), .ZN(n5146) );
  OR2_X1 U6575 ( .A1(n9526), .A2(n9846), .ZN(n5147) );
  AND2_X1 U6576 ( .A1(n7109), .A2(n9970), .ZN(n10000) );
  AND2_X2 U6577 ( .A1(n6518), .A2(n7102), .ZN(n10084) );
  INV_X1 U6578 ( .A(n10102), .ZN(n10100) );
  INV_X1 U6579 ( .A(n5824), .ZN(n8890) );
  NAND2_X1 U6580 ( .A1(n6036), .A2(n6037), .ZN(n5148) );
  OR2_X1 U6581 ( .A1(n5341), .A2(n6991), .ZN(n5149) );
  NAND2_X1 U6582 ( .A1(n8493), .A2(n8445), .ZN(n8446) );
  INV_X1 U6583 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n5176) );
  INV_X1 U6584 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n5831) );
  INV_X1 U6585 ( .A(n9910), .ZN(n6133) );
  INV_X1 U6586 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n5836) );
  INV_X1 U6587 ( .A(n8979), .ZN(n5639) );
  AND4_X1 U6588 ( .A1(n5184), .A2(n5183), .A3(n5182), .A4(n5617), .ZN(n5185)
         );
  NAND2_X1 U6589 ( .A1(n5143), .A2(n5148), .ZN(n6042) );
  NOR4_X1 U6590 ( .A1(n8484), .A2(n8508), .A3(n8491), .A4(n8483), .ZN(n8502)
         );
  NAND2_X1 U6591 ( .A1(n8575), .A2(n8924), .ZN(n8576) );
  INV_X1 U6592 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n5151) );
  INV_X1 U6593 ( .A(n8228), .ZN(n5449) );
  INV_X1 U6594 ( .A(n5905), .ZN(n9212) );
  NAND2_X1 U6595 ( .A1(n6180), .A2(n9240), .ZN(n9242) );
  OR2_X1 U6596 ( .A1(n6335), .A2(n9340), .ZN(n6349) );
  NOR2_X1 U6597 ( .A1(n6233), .A2(n6232), .ZN(n6231) );
  OR2_X1 U6598 ( .A1(n6478), .A2(n6477), .ZN(n6479) );
  INV_X1 U6599 ( .A(SI_22_), .ZN(n10600) );
  INV_X1 U6600 ( .A(SI_19_), .ZN(n5265) );
  OR2_X1 U6601 ( .A1(n5402), .A2(n5230), .ZN(n5232) );
  INV_X1 U6602 ( .A(n5208), .ZN(n5210) );
  INV_X1 U6603 ( .A(n5622), .ZN(n5162) );
  INV_X2 U6604 ( .A(n8266), .ZN(n8860) );
  OR2_X1 U6605 ( .A1(n6913), .A2(P2_U3151), .ZN(n6919) );
  INV_X1 U6606 ( .A(n5682), .ZN(n5166) );
  INV_X1 U6607 ( .A(n7581), .ZN(n7692) );
  INV_X1 U6608 ( .A(n6217), .ZN(n6215) );
  INV_X1 U6609 ( .A(n6407), .ZN(n9207) );
  OR2_X1 U6610 ( .A1(n6309), .A2(n6308), .ZN(n6311) );
  NAND2_X1 U6611 ( .A1(n6561), .A2(n4582), .ZN(n6563) );
  AND2_X1 U6612 ( .A1(n8409), .A2(n8410), .ZN(n8475) );
  OR2_X1 U6613 ( .A1(n6206), .A2(n6205), .ZN(n6233) );
  INV_X1 U6614 ( .A(n9564), .ZN(n9574) );
  AND2_X1 U6615 ( .A1(n7528), .A2(n8509), .ZN(n8328) );
  OR2_X1 U6616 ( .A1(n6714), .A2(n6428), .ZN(n6513) );
  INV_X1 U6617 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n5858) );
  NAND2_X1 U6618 ( .A1(n5242), .A2(SI_12_), .ZN(n5243) );
  INV_X1 U6619 ( .A(SI_9_), .ZN(n10614) );
  NAND2_X1 U6620 ( .A1(n5162), .A2(n10602), .ZN(n5633) );
  OR2_X1 U6621 ( .A1(n5605), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n5622) );
  AND2_X1 U6622 ( .A1(n7538), .A2(n7537), .ZN(n8216) );
  AND2_X1 U6623 ( .A1(n5199), .A2(n5198), .ZN(n8587) );
  OR2_X1 U6624 ( .A1(n5722), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n8883) );
  OR3_X1 U6625 ( .A1(n5668), .A2(P2_REG3_REG_22__SCAN_IN), .A3(
        P2_REG3_REG_23__SCAN_IN), .ZN(n5682) );
  INV_X1 U6626 ( .A(n9024), .ZN(n8994) );
  OR2_X1 U6627 ( .A1(n5543), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n5560) );
  INV_X1 U6628 ( .A(n8133), .ZN(n8241) );
  AND2_X1 U6629 ( .A1(n5774), .A2(n8203), .ZN(n9025) );
  INV_X1 U6630 ( .A(n8737), .ZN(n7845) );
  AND2_X1 U6631 ( .A1(n8114), .A2(n8101), .ZN(n8228) );
  INV_X1 U6632 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n9160) );
  NOR2_X1 U6633 ( .A1(n6099), .A2(n6866), .ZN(n6098) );
  AND2_X1 U6634 ( .A1(n6629), .A2(n6630), .ZN(n6628) );
  INV_X1 U6635 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n7520) );
  AND2_X1 U6636 ( .A1(n6409), .A2(n6408), .ZN(n6410) );
  NAND2_X1 U6637 ( .A1(n6395), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n6571) );
  NAND2_X1 U6638 ( .A1(n6872), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n5985) );
  INV_X1 U6639 ( .A(n6688), .ZN(n6860) );
  INV_X1 U6640 ( .A(n6442), .ZN(n7016) );
  INV_X1 U6641 ( .A(n8479), .ZN(n9637) );
  INV_X1 U6642 ( .A(n8473), .ZN(n9834) );
  OR2_X1 U6643 ( .A1(n7465), .A2(n7477), .ZN(n9964) );
  OR2_X1 U6644 ( .A1(n10000), .A2(n7261), .ZN(n9974) );
  INV_X1 U6645 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n9766) );
  INV_X1 U6646 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n9849) );
  INV_X1 U6647 ( .A(n8328), .ZN(n6581) );
  INV_X1 U6648 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n5853) );
  INV_X1 U6649 ( .A(n5466), .ZN(n5239) );
  INV_X1 U6650 ( .A(n5353), .ZN(n5355) );
  NAND2_X1 U6651 ( .A1(n7087), .A2(n8271), .ZN(n8709) );
  INV_X1 U6652 ( .A(n8587), .ZN(n8914) );
  AND2_X1 U6653 ( .A1(n7086), .A2(n6652), .ZN(n6912) );
  INV_X1 U6654 ( .A(n8870), .ZN(n10118) );
  INV_X1 U6655 ( .A(n10129), .ZN(n8814) );
  INV_X1 U6656 ( .A(n8254), .ZN(n8184) );
  INV_X1 U6657 ( .A(n9014), .ZN(n9032) );
  AND2_X1 U6658 ( .A1(n8218), .A2(n8217), .ZN(n8934) );
  NAND2_X1 U6659 ( .A1(n7758), .A2(n5818), .ZN(n10187) );
  NAND2_X1 U6660 ( .A1(n10137), .A2(n10182), .ZN(n10192) );
  AND2_X1 U6661 ( .A1(n5799), .A2(n5798), .ZN(n6664) );
  NAND2_X1 U6662 ( .A1(n5796), .A2(n5804), .ZN(n6667) );
  XNOR2_X1 U6663 ( .A(n5437), .B(P2_IR_REG_8__SCAN_IN), .ZN(n7332) );
  AND3_X1 U6664 ( .A1(n6338), .A2(n6337), .A3(n6336), .ZN(n9337) );
  INV_X1 U6665 ( .A(n9517), .ZN(n7891) );
  INV_X1 U6666 ( .A(n9510), .ZN(n9499) );
  INV_X1 U6667 ( .A(n8474), .ZN(n7926) );
  OR2_X1 U6668 ( .A1(n8455), .A2(n6605), .ZN(n9837) );
  INV_X1 U6669 ( .A(n9831), .ZN(n9993) );
  INV_X1 U6670 ( .A(n10070), .ZN(n10034) );
  NAND2_X1 U6671 ( .A1(n9960), .A2(n10077), .ZN(n10070) );
  NAND2_X1 U6672 ( .A1(n6414), .A2(n6413), .ZN(n6714) );
  AND2_X1 U6673 ( .A1(n6740), .A2(n6739), .ZN(n8658) );
  AND2_X1 U6674 ( .A1(n7538), .A2(n5741), .ZN(n8584) );
  NAND2_X1 U6675 ( .A1(n5689), .A2(n5688), .ZN(n8945) );
  INV_X1 U6676 ( .A(n8653), .ZN(n9026) );
  INV_X1 U6677 ( .A(n8872), .ZN(n10136) );
  INV_X1 U6678 ( .A(n8878), .ZN(n10131) );
  AND2_X1 U6679 ( .A1(n6470), .A2(n10141), .ZN(n10159) );
  NAND2_X1 U6680 ( .A1(n5824), .A2(n6647), .ZN(n6648) );
  INV_X1 U6681 ( .A(n5826), .ZN(n5827) );
  OR2_X1 U6682 ( .A1(n10201), .A2(n10187), .ZN(n9148) );
  OR2_X1 U6683 ( .A1(n10201), .A2(n10193), .ZN(n9156) );
  AND2_X1 U6684 ( .A1(n5823), .A2(n5822), .ZN(n10201) );
  OR2_X1 U6685 ( .A1(n5492), .A2(n5491), .ZN(n7581) );
  NAND2_X1 U6686 ( .A1(n9218), .A2(n9217), .ZN(n9228) );
  NAND2_X1 U6687 ( .A1(n6447), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9920) );
  INV_X1 U6688 ( .A(n7765), .ZN(n9358) );
  INV_X1 U6689 ( .A(n6451), .ZN(n6452) );
  INV_X1 U6690 ( .A(n9257), .ZN(n9400) );
  INV_X1 U6691 ( .A(n9339), .ZN(n9402) );
  OR2_X1 U6692 ( .A1(n6770), .A2(n6781), .ZN(n9507) );
  INV_X1 U6693 ( .A(n9929), .ZN(n9726) );
  INV_X1 U6694 ( .A(n9742), .ZN(n9988) );
  NAND2_X1 U6695 ( .A1(n10102), .A2(n10074), .ZN(n9846) );
  AND2_X2 U6696 ( .A1(n6518), .A2(n9894), .ZN(n10102) );
  NAND2_X1 U6697 ( .A1(n10084), .A2(n10074), .ZN(n9891) );
  INV_X1 U6698 ( .A(n10084), .ZN(n10082) );
  NAND2_X1 U6699 ( .A1(n6895), .A2(n6714), .ZN(n10001) );
  NAND2_X1 U6700 ( .A1(n5925), .A2(n6650), .ZN(n9893) );
  INV_X1 U6701 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n7761) );
  INV_X1 U6702 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n10395) );
  OAI21_X1 U6703 ( .B1(n6476), .B2(n10159), .A(n6475), .ZN(P2_U3205) );
  NOR2_X1 U6704 ( .A1(n5925), .A2(n6651), .ZN(P1_U3973) );
  OAI21_X1 U6705 ( .B1(n9891), .B2(n6616), .A(n6618), .ZN(P1_U3518) );
  INV_X2 U6706 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n7282) );
  INV_X1 U6707 ( .A(n5380), .ZN(n5152) );
  OR2_X2 U6708 ( .A1(n5473), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n5495) );
  OR2_X2 U6709 ( .A1(n5495), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n5511) );
  INV_X1 U6710 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n5159) );
  INV_X1 U6711 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n5163) );
  INV_X1 U6712 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n5165) );
  INV_X1 U6713 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n5167) );
  OR2_X2 U6714 ( .A1(n5708), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n5710) );
  INV_X1 U6715 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n5169) );
  NAND2_X1 U6716 ( .A1(n5710), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n5171) );
  NAND2_X1 U6717 ( .A1(n5722), .A2(n5171), .ZN(n8906) );
  NOR2_X1 U6718 ( .A1(P2_IR_REG_8__SCAN_IN), .A2(P2_IR_REG_14__SCAN_IN), .ZN(
        n5175) );
  NAND4_X1 U6719 ( .A1(n5175), .A2(n5174), .A3(n5173), .A4(n5172), .ZN(n5178)
         );
  NAND4_X1 U6720 ( .A1(n5484), .A2(n5390), .A3(n5489), .A4(n5176), .ZN(n5177)
         );
  NOR2_X1 U6721 ( .A1(n5178), .A2(n5177), .ZN(n5180) );
  AND2_X2 U6722 ( .A1(n6944), .A2(n5179), .ZN(n5389) );
  NOR2_X1 U6723 ( .A1(P2_IR_REG_22__SCAN_IN), .A2(P2_IR_REG_18__SCAN_IN), .ZN(
        n5184) );
  NOR2_X1 U6724 ( .A1(P2_IR_REG_17__SCAN_IN), .A2(P2_IR_REG_21__SCAN_IN), .ZN(
        n5183) );
  NOR2_X1 U6725 ( .A1(P2_IR_REG_23__SCAN_IN), .A2(P2_IR_REG_20__SCAN_IN), .ZN(
        n5182) );
  INV_X1 U6726 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n9161) );
  NAND2_X1 U6727 ( .A1(n4914), .A2(n9161), .ZN(n5188) );
  INV_X1 U6728 ( .A(n8538), .ZN(n5192) );
  NAND2_X1 U6729 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_28__SCAN_IN), 
        .ZN(n5190) );
  NAND2_X1 U6730 ( .A1(n5308), .A2(n5190), .ZN(n5191) );
  NAND2_X1 U6731 ( .A1(n5192), .A2(n5193), .ZN(n5382) );
  NAND2_X1 U6732 ( .A1(n8906), .A2(n5346), .ZN(n5199) );
  INV_X1 U6733 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n5196) );
  NAND2_X1 U6734 ( .A1(n5775), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n5195) );
  NAND2_X1 U6735 ( .A1(n8538), .A2(n5193), .ZN(n5319) );
  NAND2_X1 U6736 ( .A1(n5776), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n5194) );
  OAI211_X1 U6737 ( .C1(n7535), .C2(n5196), .A(n5195), .B(n5194), .ZN(n5197)
         );
  INV_X1 U6738 ( .A(n5197), .ZN(n5198) );
  INV_X1 U6739 ( .A(P2_RD_REG_SCAN_IN), .ZN(n5200) );
  NAND2_X1 U6740 ( .A1(n5325), .A2(SI_1_), .ZN(n5202) );
  MUX2_X1 U6741 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(P2_DATAO_REG_0__SCAN_IN), 
        .S(n5217), .Z(n5201) );
  NAND2_X1 U6742 ( .A1(n5201), .A2(SI_0_), .ZN(n5326) );
  INV_X1 U6743 ( .A(SI_1_), .ZN(n5203) );
  NAND2_X1 U6744 ( .A1(n5208), .A2(SI_2_), .ZN(n5213) );
  INV_X1 U6745 ( .A(SI_2_), .ZN(n5209) );
  NAND2_X1 U6746 ( .A1(n5210), .A2(n5209), .ZN(n5211) );
  NAND2_X1 U6747 ( .A1(n5213), .A2(n5211), .ZN(n5336) );
  INV_X1 U6748 ( .A(n5336), .ZN(n5212) );
  NAND2_X1 U6749 ( .A1(n5214), .A2(SI_3_), .ZN(n5216) );
  INV_X1 U6750 ( .A(n5354), .ZN(n5215) );
  NAND2_X1 U6751 ( .A1(n5353), .A2(n5215), .ZN(n5356) );
  MUX2_X1 U6752 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(P2_DATAO_REG_4__SCAN_IN), 
        .S(n5217), .Z(n5218) );
  NAND2_X1 U6753 ( .A1(n5218), .A2(SI_4_), .ZN(n5222) );
  INV_X1 U6754 ( .A(n5218), .ZN(n5220) );
  INV_X1 U6755 ( .A(SI_4_), .ZN(n5219) );
  NAND2_X1 U6756 ( .A1(n5220), .A2(n5219), .ZN(n5221) );
  AND2_X1 U6757 ( .A1(n5222), .A2(n5221), .ZN(n5373) );
  MUX2_X1 U6758 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(P2_DATAO_REG_5__SCAN_IN), 
        .S(n6672), .Z(n5223) );
  XNOR2_X1 U6759 ( .A(n5223), .B(n10574), .ZN(n5392) );
  INV_X1 U6760 ( .A(n5392), .ZN(n5224) );
  MUX2_X1 U6761 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .S(n6671), .Z(n5226) );
  NAND2_X1 U6762 ( .A1(n5226), .A2(SI_6_), .ZN(n5415) );
  OAI21_X1 U6763 ( .B1(n5226), .B2(SI_6_), .A(n5415), .ZN(n5402) );
  INV_X1 U6764 ( .A(n5228), .ZN(n5227) );
  INV_X1 U6765 ( .A(n5417), .ZN(n5419) );
  NOR2_X1 U6766 ( .A1(n5227), .A2(n5419), .ZN(n5230) );
  AND2_X1 U6767 ( .A1(n5415), .A2(n5228), .ZN(n5229) );
  OR2_X1 U6768 ( .A1(n5230), .A2(n5229), .ZN(n5231) );
  MUX2_X1 U6769 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(P2_DATAO_REG_8__SCAN_IN), 
        .S(n6671), .Z(n5233) );
  XNOR2_X1 U6770 ( .A(n5233), .B(SI_8_), .ZN(n5435) );
  MUX2_X1 U6771 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(P2_DATAO_REG_9__SCAN_IN), 
        .S(n6672), .Z(n5234) );
  XNOR2_X1 U6772 ( .A(n5234), .B(n10614), .ZN(n5451) );
  INV_X1 U6773 ( .A(n5234), .ZN(n5235) );
  NAND2_X1 U6774 ( .A1(n5235), .A2(n10614), .ZN(n5236) );
  MUX2_X1 U6775 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(P2_DATAO_REG_10__SCAN_IN), 
        .S(n6671), .Z(n5238) );
  OAI21_X1 U6776 ( .B1(n5238), .B2(SI_10_), .A(n5240), .ZN(n5466) );
  MUX2_X1 U6777 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(P2_DATAO_REG_11__SCAN_IN), 
        .S(n6671), .Z(n5241) );
  MUX2_X1 U6778 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(P2_DATAO_REG_12__SCAN_IN), 
        .S(n6671), .Z(n5242) );
  MUX2_X1 U6779 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(P2_DATAO_REG_13__SCAN_IN), 
        .S(n6671), .Z(n5244) );
  INV_X1 U6780 ( .A(n5244), .ZN(n5246) );
  INV_X1 U6781 ( .A(SI_13_), .ZN(n5245) );
  NAND2_X1 U6782 ( .A1(n5246), .A2(n5245), .ZN(n5247) );
  MUX2_X1 U6783 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(P2_DATAO_REG_14__SCAN_IN), 
        .S(n6671), .Z(n5536) );
  MUX2_X1 U6784 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(P2_DATAO_REG_15__SCAN_IN), 
        .S(n6672), .Z(n5551) );
  INV_X1 U6785 ( .A(n5551), .ZN(n5249) );
  NAND2_X1 U6786 ( .A1(n5250), .A2(n5249), .ZN(n5252) );
  NAND2_X1 U6787 ( .A1(n5569), .A2(n10554), .ZN(n5253) );
  MUX2_X1 U6788 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(P2_DATAO_REG_16__SCAN_IN), 
        .S(n6672), .Z(n5567) );
  NAND2_X1 U6789 ( .A1(n5253), .A2(n5567), .ZN(n5256) );
  INV_X1 U6790 ( .A(n5569), .ZN(n5254) );
  NAND2_X1 U6791 ( .A1(n5254), .A2(SI_16_), .ZN(n5255) );
  NAND2_X1 U6792 ( .A1(n5256), .A2(n5255), .ZN(n5586) );
  MUX2_X1 U6793 ( .A(n7313), .B(n10347), .S(n6671), .Z(n5257) );
  INV_X1 U6794 ( .A(n5257), .ZN(n5258) );
  NAND2_X1 U6795 ( .A1(n5258), .A2(SI_17_), .ZN(n5259) );
  NAND2_X1 U6796 ( .A1(n5260), .A2(n5259), .ZN(n5585) );
  MUX2_X1 U6797 ( .A(n7427), .B(n10395), .S(n6672), .Z(n5261) );
  XNOR2_X1 U6798 ( .A(n5261), .B(SI_18_), .ZN(n5597) );
  INV_X1 U6799 ( .A(n5597), .ZN(n5264) );
  INV_X1 U6800 ( .A(n5261), .ZN(n5262) );
  NAND2_X1 U6801 ( .A1(n5262), .A2(SI_18_), .ZN(n5263) );
  MUX2_X1 U6802 ( .A(n7512), .B(n10406), .S(n6671), .Z(n5266) );
  NAND2_X1 U6803 ( .A1(n5266), .A2(n5265), .ZN(n5269) );
  INV_X1 U6804 ( .A(n5266), .ZN(n5267) );
  NAND2_X1 U6805 ( .A1(n5267), .A2(SI_19_), .ZN(n5268) );
  NAND2_X1 U6806 ( .A1(n5269), .A2(n5268), .ZN(n5614) );
  MUX2_X1 U6807 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(P2_DATAO_REG_20__SCAN_IN), 
        .S(n6671), .Z(n5628) );
  INV_X1 U6808 ( .A(n5628), .ZN(n5270) );
  MUX2_X1 U6809 ( .A(n7616), .B(n10389), .S(n6671), .Z(n5640) );
  NOR2_X1 U6810 ( .A1(n5271), .A2(SI_21_), .ZN(n5272) );
  MUX2_X1 U6811 ( .A(n7757), .B(n7761), .S(n6671), .Z(n5273) );
  NAND2_X1 U6812 ( .A1(n5273), .A2(n10600), .ZN(n5278) );
  INV_X1 U6813 ( .A(n5273), .ZN(n5274) );
  NAND2_X1 U6814 ( .A1(n5274), .A2(SI_22_), .ZN(n5275) );
  NAND2_X1 U6815 ( .A1(n5278), .A2(n5275), .ZN(n5650) );
  INV_X1 U6816 ( .A(n5650), .ZN(n5276) );
  NAND2_X1 U6817 ( .A1(n5277), .A2(n5276), .ZN(n5279) );
  INV_X1 U6818 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n7800) );
  INV_X1 U6819 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n5280) );
  MUX2_X1 U6820 ( .A(n7800), .B(n5280), .S(n6671), .Z(n5281) );
  INV_X1 U6821 ( .A(SI_23_), .ZN(n10557) );
  NAND2_X1 U6822 ( .A1(n5281), .A2(n10557), .ZN(n5285) );
  INV_X1 U6823 ( .A(n5281), .ZN(n5282) );
  NAND2_X1 U6824 ( .A1(n5282), .A2(SI_23_), .ZN(n5283) );
  NAND2_X1 U6825 ( .A1(n5285), .A2(n5283), .ZN(n5662) );
  INV_X1 U6826 ( .A(n5662), .ZN(n5284) );
  INV_X1 U6827 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n7908) );
  MUX2_X1 U6828 ( .A(n7908), .B(n10588), .S(n6672), .Z(n5286) );
  INV_X1 U6829 ( .A(SI_24_), .ZN(n10524) );
  NAND2_X1 U6830 ( .A1(n5286), .A2(n10524), .ZN(n5289) );
  INV_X1 U6831 ( .A(n5286), .ZN(n5287) );
  NAND2_X1 U6832 ( .A1(n5287), .A2(SI_24_), .ZN(n5288) );
  INV_X1 U6833 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n7933) );
  MUX2_X1 U6834 ( .A(n7933), .B(n10526), .S(n5217), .Z(n5290) );
  INV_X1 U6835 ( .A(SI_25_), .ZN(n10584) );
  NAND2_X1 U6836 ( .A1(n5290), .A2(n10584), .ZN(n5293) );
  INV_X1 U6837 ( .A(n5290), .ZN(n5291) );
  NAND2_X1 U6838 ( .A1(n5291), .A2(SI_25_), .ZN(n5292) );
  NAND2_X1 U6839 ( .A1(n5692), .A2(n5693), .ZN(n5294) );
  INV_X1 U6840 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n7965) );
  INV_X1 U6841 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n10530) );
  MUX2_X1 U6842 ( .A(n7965), .B(n10530), .S(n5217), .Z(n5296) );
  INV_X1 U6843 ( .A(SI_26_), .ZN(n5295) );
  NAND2_X1 U6844 ( .A1(n5296), .A2(n5295), .ZN(n5299) );
  INV_X1 U6845 ( .A(n5296), .ZN(n5297) );
  NAND2_X1 U6846 ( .A1(n5297), .A2(SI_26_), .ZN(n5298) );
  NAND2_X1 U6847 ( .A1(n5705), .A2(n5704), .ZN(n5300) );
  NAND2_X1 U6848 ( .A1(n5300), .A2(n5299), .ZN(n5306) );
  INV_X1 U6849 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n8540) );
  INV_X1 U6850 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n5301) );
  MUX2_X1 U6851 ( .A(n8540), .B(n5301), .S(n5217), .Z(n5302) );
  INV_X1 U6852 ( .A(SI_27_), .ZN(n10572) );
  NAND2_X1 U6853 ( .A1(n5302), .A2(n10572), .ZN(n5718) );
  INV_X1 U6854 ( .A(n5302), .ZN(n5303) );
  NAND2_X1 U6855 ( .A1(n5303), .A2(SI_27_), .ZN(n5304) );
  OR2_X1 U6856 ( .A1(n5306), .A2(n5305), .ZN(n5307) );
  NAND2_X1 U6857 ( .A1(n5719), .A2(n5307), .ZN(n8273) );
  XNOR2_X1 U6858 ( .A(n5308), .B(n9160), .ZN(n5771) );
  NAND2_X1 U6859 ( .A1(n8273), .A2(n8198), .ZN(n5312) );
  OR2_X1 U6860 ( .A1(n4507), .A2(n8540), .ZN(n5311) );
  NAND2_X1 U6861 ( .A1(n5346), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n5316) );
  NAND2_X1 U6862 ( .A1(n5348), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n5314) );
  INV_X1 U6863 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n6914) );
  OR2_X1 U6864 ( .A1(n5319), .A2(n6914), .ZN(n5313) );
  NAND4_X1 U6865 ( .A1(n5316), .A2(n5315), .A3(n5314), .A4(n5313), .ZN(n5317)
         );
  NAND2_X1 U6866 ( .A1(n5225), .A2(SI_0_), .ZN(n5318) );
  XNOR2_X1 U6867 ( .A(n5318), .B(P1_DATAO_REG_0__SCAN_IN), .ZN(n9174) );
  NAND2_X1 U6868 ( .A1(n5317), .A2(n6839), .ZN(n7008) );
  INV_X1 U6869 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n6992) );
  INV_X1 U6870 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n6925) );
  OAI22_X1 U6871 ( .A1(n5382), .A2(n6992), .B1(n6925), .B2(n5319), .ZN(n5320)
         );
  INV_X1 U6872 ( .A(n5320), .ZN(n5324) );
  INV_X1 U6873 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n5321) );
  INV_X1 U6874 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n7239) );
  INV_X1 U6875 ( .A(n5322), .ZN(n5323) );
  OR2_X1 U6876 ( .A1(n5358), .A2(n4795), .ZN(n5331) );
  XNOR2_X1 U6877 ( .A(n5325), .B(SI_1_), .ZN(n5327) );
  XNOR2_X1 U6878 ( .A(n5327), .B(n5326), .ZN(n6675) );
  OR2_X1 U6879 ( .A1(n5339), .A2(n6675), .ZN(n5330) );
  INV_X1 U6880 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n5329) );
  NAND3_X2 U6881 ( .A1(n5331), .A2(n5330), .A3(n5149), .ZN(n7431) );
  NAND2_X1 U6882 ( .A1(n7008), .A2(n7005), .ZN(n7007) );
  NAND2_X1 U6883 ( .A1(n6841), .A2(n7011), .ZN(n5332) );
  NAND2_X1 U6884 ( .A1(n7007), .A2(n5332), .ZN(n10145) );
  NAND2_X1 U6885 ( .A1(n5346), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n5335) );
  NAND2_X1 U6886 ( .A1(n5348), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n5333) );
  OR2_X1 U6887 ( .A1(n4507), .A2(n5207), .ZN(n5344) );
  NAND2_X1 U6888 ( .A1(n4563), .A2(n5336), .ZN(n5337) );
  NAND2_X1 U6889 ( .A1(n5338), .A2(n5337), .ZN(n6677) );
  OR2_X1 U6890 ( .A1(n5339), .A2(n6677), .ZN(n5343) );
  OR2_X1 U6891 ( .A1(n5341), .A2(n6947), .ZN(n5342) );
  AND3_X2 U6892 ( .A1(n5344), .A2(n5343), .A3(n5342), .ZN(n10143) );
  INV_X1 U6893 ( .A(n8743), .ZN(n7078) );
  NAND2_X1 U6894 ( .A1(n7078), .A2(n10143), .ZN(n5345) );
  NAND2_X1 U6895 ( .A1(n5346), .A2(n7282), .ZN(n5352) );
  NAND2_X1 U6896 ( .A1(n5635), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n5351) );
  INV_X1 U6897 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n5347) );
  NAND2_X1 U6898 ( .A1(n5348), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n5349) );
  NAND2_X1 U6899 ( .A1(n5355), .A2(n5354), .ZN(n5357) );
  NAND2_X1 U6900 ( .A1(n5357), .A2(n5356), .ZN(n6673) );
  OR2_X1 U6901 ( .A1(n5339), .A2(n6673), .ZN(n5364) );
  INV_X1 U6902 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n6674) );
  OR2_X1 U6903 ( .A1(n4507), .A2(n6674), .ZN(n5362) );
  XNOR2_X1 U6904 ( .A(n5361), .B(n5360), .ZN(n6976) );
  NAND2_X1 U6905 ( .A1(n10149), .A2(n10165), .ZN(n5365) );
  INV_X1 U6906 ( .A(n10149), .ZN(n5752) );
  INV_X1 U6907 ( .A(n10165), .ZN(n5753) );
  NAND2_X1 U6908 ( .A1(n5752), .A2(n5753), .ZN(n5366) );
  NAND2_X1 U6909 ( .A1(n5635), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n5371) );
  NAND2_X1 U6910 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n5367) );
  NAND2_X1 U6911 ( .A1(n5380), .A2(n5367), .ZN(n7272) );
  NAND2_X1 U6912 ( .A1(n5346), .A2(n7272), .ZN(n5370) );
  NAND2_X1 U6913 ( .A1(n5776), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n5369) );
  NAND2_X1 U6914 ( .A1(n5348), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n5368) );
  NAND4_X1 U6915 ( .A1(n5371), .A2(n5370), .A3(n5369), .A4(n5368), .ZN(n8742)
         );
  OR2_X1 U6916 ( .A1(n5389), .A2(n5488), .ZN(n5372) );
  XNOR2_X1 U6917 ( .A(n5372), .B(n5388), .ZN(n7073) );
  OR2_X1 U6918 ( .A1(n5374), .A2(n5373), .ZN(n5375) );
  NAND2_X1 U6919 ( .A1(n5376), .A2(n5375), .ZN(n6676) );
  OR2_X1 U6920 ( .A1(n5339), .A2(n6676), .ZN(n5379) );
  INV_X1 U6921 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n5377) );
  OR2_X1 U6922 ( .A1(n4507), .A2(n5377), .ZN(n5378) );
  OAI211_X1 U6923 ( .C1(n5781), .C2(n7073), .A(n5379), .B(n5378), .ZN(n7273)
         );
  NOR2_X1 U6924 ( .A1(n8742), .A2(n7273), .ZN(n5755) );
  NAND2_X1 U6925 ( .A1(n8742), .A2(n7273), .ZN(n5756) );
  NAND2_X1 U6926 ( .A1(n5380), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n5381) );
  AND2_X1 U6927 ( .A1(n5406), .A2(n5381), .ZN(n7434) );
  INV_X1 U6928 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n5383) );
  OAI22_X1 U6929 ( .A1(n7434), .A2(n5581), .B1(n7535), .B2(n5383), .ZN(n5387)
         );
  INV_X1 U6930 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n5385) );
  NAND2_X1 U6931 ( .A1(n5348), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n5384) );
  OAI21_X1 U6932 ( .B1(n5385), .B2(n7532), .A(n5384), .ZN(n5386) );
  NAND2_X1 U6933 ( .A1(n5389), .A2(n5388), .ZN(n5399) );
  NAND2_X1 U6934 ( .A1(n5399), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5391) );
  XNOR2_X1 U6935 ( .A(n5393), .B(n5392), .ZN(n6681) );
  OR2_X1 U6936 ( .A1(n5339), .A2(n6681), .ZN(n5395) );
  INV_X1 U6937 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n6680) );
  OR2_X1 U6938 ( .A1(n4507), .A2(n6680), .ZN(n5394) );
  OAI211_X1 U6939 ( .C1(n5781), .C2(n6950), .A(n5395), .B(n5394), .ZN(n7428)
         );
  AND2_X1 U6940 ( .A1(n7458), .A2(n7428), .ZN(n5398) );
  INV_X1 U6941 ( .A(n7458), .ZN(n5396) );
  NAND2_X1 U6942 ( .A1(n5396), .A2(n7435), .ZN(n5397) );
  NAND2_X1 U6943 ( .A1(n5423), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5400) );
  AOI22_X1 U6944 ( .A1(n5619), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n6655), .B2(
        n7147), .ZN(n5405) );
  OR2_X1 U6945 ( .A1(n5401), .A2(n5402), .ZN(n5416) );
  NAND2_X1 U6946 ( .A1(n5401), .A2(n5402), .ZN(n5403) );
  AND2_X1 U6947 ( .A1(n5416), .A2(n5403), .ZN(n6662) );
  NAND2_X1 U6948 ( .A1(n6662), .A2(n8198), .ZN(n5404) );
  NAND2_X1 U6949 ( .A1(n7457), .A2(n10177), .ZN(n5412) );
  NAND2_X1 U6950 ( .A1(n5635), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n5411) );
  NAND2_X1 U6951 ( .A1(n5406), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5407) );
  NAND2_X1 U6952 ( .A1(n5428), .A2(n5407), .ZN(n7461) );
  NAND2_X1 U6953 ( .A1(n5346), .A2(n7461), .ZN(n5410) );
  NAND2_X1 U6954 ( .A1(n5776), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n5409) );
  NAND2_X1 U6955 ( .A1(n5348), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n5408) );
  NAND4_X1 U6956 ( .A1(n5411), .A2(n5410), .A3(n5409), .A4(n5408), .ZN(n8741)
         );
  NAND2_X1 U6957 ( .A1(n5412), .A2(n8741), .ZN(n5414) );
  OR2_X2 U6958 ( .A1(n7457), .A2(n10177), .ZN(n5413) );
  AND2_X1 U6959 ( .A1(n5416), .A2(n5415), .ZN(n5418) );
  NAND2_X1 U6960 ( .A1(n5418), .A2(n5417), .ZN(n5422) );
  INV_X1 U6961 ( .A(n5418), .ZN(n5420) );
  NAND2_X1 U6962 ( .A1(n5420), .A2(n5419), .ZN(n5421) );
  NAND2_X1 U6963 ( .A1(n6678), .A2(n8198), .ZN(n5427) );
  INV_X1 U6964 ( .A(n5454), .ZN(n5424) );
  NAND2_X1 U6965 ( .A1(n5424), .A2(P2_IR_REG_7__SCAN_IN), .ZN(n5425) );
  NAND2_X1 U6966 ( .A1(n5454), .A2(n5484), .ZN(n5436) );
  AOI22_X1 U6967 ( .A1(n5619), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n6655), .B2(
        n7156), .ZN(n5426) );
  NAND2_X1 U6968 ( .A1(n5427), .A2(n5426), .ZN(n7507) );
  NAND2_X1 U6969 ( .A1(n5428), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n5429) );
  AND2_X1 U6970 ( .A1(n5442), .A2(n5429), .ZN(n7505) );
  INV_X1 U6971 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n7137) );
  OAI22_X1 U6972 ( .A1(n7505), .A2(n5581), .B1(n7535), .B2(n7137), .ZN(n5432)
         );
  INV_X1 U6973 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n7136) );
  NAND2_X1 U6974 ( .A1(n5348), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n5430) );
  OAI21_X1 U6975 ( .B1(n7136), .B2(n7532), .A(n5430), .ZN(n5431) );
  AND2_X1 U6976 ( .A1(n7507), .A2(n8740), .ZN(n5433) );
  XNOR2_X1 U6977 ( .A(n5434), .B(n5435), .ZN(n6686) );
  NAND2_X1 U6978 ( .A1(n6686), .A2(n8198), .ZN(n5439) );
  NAND2_X1 U6979 ( .A1(n5436), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5437) );
  AOI22_X1 U6980 ( .A1(n5619), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n6655), .B2(
        n7332), .ZN(n5438) );
  NAND2_X1 U6981 ( .A1(n5439), .A2(n5438), .ZN(n7630) );
  INV_X1 U6982 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n7315) );
  INV_X1 U6983 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n10209) );
  OR2_X1 U6984 ( .A1(n7532), .A2(n10209), .ZN(n5440) );
  OAI21_X1 U6985 ( .B1(n7535), .B2(n7315), .A(n5440), .ZN(n5441) );
  INV_X1 U6986 ( .A(n5441), .ZN(n5448) );
  NAND2_X1 U6987 ( .A1(n5442), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n5443) );
  AND2_X1 U6988 ( .A1(n5457), .A2(n5443), .ZN(n7631) );
  INV_X1 U6989 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n5444) );
  OR2_X1 U6990 ( .A1(n7530), .A2(n5444), .ZN(n5445) );
  OAI21_X1 U6991 ( .B1(n5581), .B2(n7631), .A(n5445), .ZN(n5446) );
  INV_X1 U6992 ( .A(n5446), .ZN(n5447) );
  NAND2_X1 U6993 ( .A1(n7630), .A2(n7621), .ZN(n8101) );
  INV_X1 U6994 ( .A(n7621), .ZN(n8739) );
  NAND2_X1 U6995 ( .A1(n7630), .A2(n8739), .ZN(n5450) );
  XNOR2_X1 U6996 ( .A(n5452), .B(n5451), .ZN(n6691) );
  NAND2_X1 U6997 ( .A1(n6691), .A2(n8198), .ZN(n5456) );
  OAI21_X1 U6998 ( .B1(P2_IR_REG_7__SCAN_IN), .B2(P2_IR_REG_8__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5453) );
  NAND2_X1 U6999 ( .A1(n5454), .A2(n5453), .ZN(n5470) );
  XNOR2_X1 U7000 ( .A(n5470), .B(P2_IR_REG_9__SCAN_IN), .ZN(n7339) );
  INV_X1 U7001 ( .A(n7339), .ZN(n7323) );
  AOI22_X1 U7002 ( .A1(n5619), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n6655), .B2(
        n7323), .ZN(n5455) );
  NAND2_X1 U7003 ( .A1(n5456), .A2(n5455), .ZN(n7645) );
  NAND2_X1 U7004 ( .A1(n5635), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n5462) );
  NAND2_X1 U7005 ( .A1(n5457), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n5458) );
  NAND2_X1 U7006 ( .A1(n5473), .A2(n5458), .ZN(n7622) );
  NAND2_X1 U7007 ( .A1(n5346), .A2(n7622), .ZN(n5461) );
  INV_X1 U7008 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n7322) );
  OR2_X1 U7009 ( .A1(n7532), .A2(n7322), .ZN(n5460) );
  NAND2_X1 U7010 ( .A1(n5775), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n5459) );
  NAND4_X1 U7011 ( .A1(n5462), .A2(n5461), .A3(n5460), .A4(n5459), .ZN(n8738)
         );
  OR2_X1 U7012 ( .A1(n7645), .A2(n8738), .ZN(n5463) );
  NAND2_X1 U7013 ( .A1(n7645), .A2(n8738), .ZN(n5464) );
  NAND2_X1 U7014 ( .A1(n5467), .A2(n5466), .ZN(n5468) );
  OAI21_X1 U7015 ( .B1(n5470), .B2(P2_IR_REG_9__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5471) );
  XNOR2_X1 U7016 ( .A(n5471), .B(P2_IR_REG_10__SCAN_IN), .ZN(n7382) );
  AOI22_X1 U7017 ( .A1(n5619), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n6655), .B2(
        n7382), .ZN(n5472) );
  NAND2_X1 U7018 ( .A1(n5473), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n5474) );
  AND2_X1 U7019 ( .A1(n5495), .A2(n5474), .ZN(n7775) );
  INV_X1 U7020 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n7774) );
  OAI22_X1 U7021 ( .A1(n7775), .A2(n5581), .B1(n7535), .B2(n7774), .ZN(n5477)
         );
  INV_X1 U7022 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n7370) );
  NAND2_X1 U7023 ( .A1(n5775), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n5475) );
  OAI21_X1 U7024 ( .B1(n7370), .B2(n7532), .A(n5475), .ZN(n5476) );
  AND2_X1 U7025 ( .A1(n7777), .A2(n8737), .ZN(n5478) );
  XNOR2_X1 U7026 ( .A(n5480), .B(n5479), .ZN(n6712) );
  NAND2_X1 U7027 ( .A1(n6712), .A2(n8198), .ZN(n5494) );
  INV_X1 U7028 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n5483) );
  INV_X1 U7029 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n5482) );
  INV_X1 U7030 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n5481) );
  AND4_X1 U7031 ( .A1(n5484), .A2(n5483), .A3(n5482), .A4(n5481), .ZN(n5485)
         );
  NOR2_X1 U7032 ( .A1(n5490), .A2(n5488), .ZN(n5487) );
  MUX2_X1 U7033 ( .A(n5488), .B(n5487), .S(P2_IR_REG_11__SCAN_IN), .Z(n5492)
         );
  NAND2_X1 U7034 ( .A1(n5490), .A2(n5489), .ZN(n5523) );
  INV_X1 U7035 ( .A(n5523), .ZN(n5491) );
  AOI22_X1 U7036 ( .A1(n5619), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n6655), .B2(
        n7692), .ZN(n5493) );
  NAND2_X1 U7037 ( .A1(n5635), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n5501) );
  NAND2_X1 U7038 ( .A1(n5495), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n5496) );
  NAND2_X1 U7039 ( .A1(n5511), .A2(n5496), .ZN(n7794) );
  NAND2_X1 U7040 ( .A1(n5346), .A2(n7794), .ZN(n5500) );
  INV_X1 U7041 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n5497) );
  OR2_X1 U7042 ( .A1(n7532), .A2(n5497), .ZN(n5499) );
  NAND2_X1 U7043 ( .A1(n5775), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n5498) );
  NAND4_X1 U7044 ( .A1(n5501), .A2(n5500), .A3(n5499), .A4(n5498), .ZN(n8736)
         );
  NOR2_X1 U7045 ( .A1(n10197), .A2(n8736), .ZN(n5502) );
  NAND2_X1 U7046 ( .A1(n10197), .A2(n8736), .ZN(n5503) );
  NAND2_X1 U7047 ( .A1(n5505), .A2(n5504), .ZN(n5506) );
  NAND2_X1 U7048 ( .A1(n5507), .A2(n5506), .ZN(n6720) );
  OR2_X1 U7049 ( .A1(n6720), .A2(n5339), .ZN(n5510) );
  NAND2_X1 U7050 ( .A1(n5523), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5508) );
  XNOR2_X1 U7051 ( .A(n5508), .B(P2_IR_REG_12__SCAN_IN), .ZN(n7699) );
  AOI22_X1 U7052 ( .A1(n5619), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n6655), .B2(
        n7699), .ZN(n5509) );
  NAND2_X1 U7053 ( .A1(n5635), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n5516) );
  NAND2_X1 U7054 ( .A1(n5511), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n5512) );
  NAND2_X1 U7055 ( .A1(n5529), .A2(n5512), .ZN(n7937) );
  NAND2_X1 U7056 ( .A1(n5346), .A2(n7937), .ZN(n5515) );
  INV_X1 U7057 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n7687) );
  OR2_X1 U7058 ( .A1(n7532), .A2(n7687), .ZN(n5514) );
  NAND2_X1 U7059 ( .A1(n5775), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n5513) );
  NAND4_X1 U7060 ( .A1(n5516), .A2(n5515), .A3(n5514), .A4(n5513), .ZN(n8735)
         );
  INV_X1 U7061 ( .A(n7947), .ZN(n5517) );
  OR2_X1 U7062 ( .A1(n5520), .A2(n5519), .ZN(n5521) );
  AND2_X1 U7063 ( .A1(n5522), .A2(n5521), .ZN(n6849) );
  NAND2_X1 U7064 ( .A1(n6849), .A2(n8198), .ZN(n5526) );
  OR2_X1 U7065 ( .A1(n5523), .A2(P2_IR_REG_12__SCAN_IN), .ZN(n5524) );
  NAND2_X1 U7066 ( .A1(n5524), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5539) );
  XNOR2_X1 U7067 ( .A(n5539), .B(P2_IR_REG_13__SCAN_IN), .ZN(n8760) );
  AOI22_X1 U7068 ( .A1(n5619), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n6655), .B2(
        n8760), .ZN(n5525) );
  INV_X1 U7069 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n10105) );
  INV_X1 U7070 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n10110) );
  OR2_X1 U7071 ( .A1(n7532), .A2(n10110), .ZN(n5527) );
  OAI21_X1 U7072 ( .B1(n7535), .B2(n10105), .A(n5527), .ZN(n5528) );
  INV_X1 U7073 ( .A(n5528), .ZN(n5534) );
  NAND2_X1 U7074 ( .A1(n5529), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n5530) );
  AND2_X1 U7075 ( .A1(n5543), .A2(n5530), .ZN(n7957) );
  INV_X1 U7076 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n7911) );
  OR2_X1 U7077 ( .A1(n7530), .A2(n7911), .ZN(n5531) );
  OAI21_X1 U7078 ( .B1(n5581), .B2(n7957), .A(n5531), .ZN(n5532) );
  INV_X1 U7079 ( .A(n5532), .ZN(n5533) );
  NAND2_X1 U7080 ( .A1(n7953), .A2(n7985), .ZN(n8054) );
  NAND2_X1 U7081 ( .A1(n8055), .A2(n8054), .ZN(n8238) );
  NAND2_X1 U7082 ( .A1(n7953), .A2(n7981), .ZN(n7968) );
  XNOR2_X1 U7083 ( .A(n5536), .B(SI_14_), .ZN(n5537) );
  XNOR2_X1 U7084 ( .A(n5535), .B(n5537), .ZN(n6889) );
  NAND2_X1 U7085 ( .A1(n6889), .A2(n8198), .ZN(n5542) );
  INV_X1 U7086 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n5538) );
  NAND2_X1 U7087 ( .A1(n5539), .A2(n5538), .ZN(n5540) );
  NAND2_X1 U7088 ( .A1(n5540), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5555) );
  XNOR2_X1 U7089 ( .A(n5555), .B(P2_IR_REG_14__SCAN_IN), .ZN(n8764) );
  AOI22_X1 U7090 ( .A1(n5619), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n6655), .B2(
        n8764), .ZN(n5541) );
  NAND2_X1 U7091 ( .A1(n5635), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n5548) );
  NAND2_X1 U7092 ( .A1(n5543), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n5544) );
  NAND2_X1 U7093 ( .A1(n5560), .A2(n5544), .ZN(n8020) );
  NAND2_X1 U7094 ( .A1(n5346), .A2(n8020), .ZN(n5547) );
  INV_X1 U7095 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n8763) );
  OR2_X1 U7096 ( .A1(n7532), .A2(n8763), .ZN(n5546) );
  NAND2_X1 U7097 ( .A1(n5348), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n5545) );
  NAND4_X1 U7098 ( .A1(n5548), .A2(n5547), .A3(n5546), .A4(n5545), .ZN(n8734)
         );
  NAND2_X1 U7099 ( .A1(n8015), .A2(n8734), .ZN(n5549) );
  AND2_X1 U7100 ( .A1(n7968), .A2(n5549), .ZN(n5550) );
  XNOR2_X1 U7101 ( .A(n5551), .B(SI_15_), .ZN(n5552) );
  XNOR2_X1 U7102 ( .A(n5553), .B(n5552), .ZN(n7032) );
  NAND2_X1 U7103 ( .A1(n7032), .A2(n8198), .ZN(n5559) );
  INV_X1 U7104 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n5554) );
  NAND2_X1 U7105 ( .A1(n5555), .A2(n5554), .ZN(n5556) );
  NAND2_X1 U7106 ( .A1(n5556), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5557) );
  XNOR2_X1 U7107 ( .A(n5557), .B(P2_IR_REG_15__SCAN_IN), .ZN(n8789) );
  AOI22_X1 U7108 ( .A1(n5619), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n6655), .B2(
        n8789), .ZN(n5558) );
  NAND2_X1 U7109 ( .A1(n5635), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n5565) );
  NAND2_X1 U7110 ( .A1(n5560), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n5561) );
  NAND2_X1 U7111 ( .A1(n5578), .A2(n5561), .ZN(n8011) );
  NAND2_X1 U7112 ( .A1(n5346), .A2(n8011), .ZN(n5564) );
  INV_X1 U7113 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n8767) );
  OR2_X1 U7114 ( .A1(n7532), .A2(n8767), .ZN(n5563) );
  NAND2_X1 U7115 ( .A1(n5775), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n5562) );
  NAND4_X1 U7116 ( .A1(n5565), .A2(n5564), .A3(n5563), .A4(n5562), .ZN(n8733)
         );
  AND2_X1 U7117 ( .A1(n8006), .A2(n8733), .ZN(n5566) );
  XNOR2_X1 U7118 ( .A(n5567), .B(n10554), .ZN(n5568) );
  XNOR2_X1 U7119 ( .A(n5569), .B(n5568), .ZN(n7183) );
  NAND2_X1 U7120 ( .A1(n7183), .A2(n8198), .ZN(n5575) );
  NAND2_X1 U7121 ( .A1(n5570), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5571) );
  MUX2_X1 U7122 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5571), .S(
        P2_IR_REG_16__SCAN_IN), .Z(n5573) );
  INV_X1 U7123 ( .A(n5572), .ZN(n5587) );
  AND2_X1 U7124 ( .A1(n5573), .A2(n5587), .ZN(n8784) );
  AOI22_X1 U7125 ( .A1(n5619), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n6655), .B2(
        n8784), .ZN(n5574) );
  INV_X1 U7126 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n8037) );
  INV_X1 U7127 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n8777) );
  OR2_X1 U7128 ( .A1(n7532), .A2(n8777), .ZN(n5576) );
  OAI21_X1 U7129 ( .B1(n7535), .B2(n8037), .A(n5576), .ZN(n5577) );
  INV_X1 U7130 ( .A(n5577), .ZN(n5584) );
  NAND2_X1 U7131 ( .A1(n5578), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n5579) );
  AND2_X1 U7132 ( .A1(n5591), .A2(n5579), .ZN(n8645) );
  INV_X1 U7133 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n8029) );
  OR2_X1 U7134 ( .A1(n7530), .A2(n8029), .ZN(n5580) );
  OAI21_X1 U7135 ( .B1(n5581), .B2(n8645), .A(n5580), .ZN(n5582) );
  INV_X1 U7136 ( .A(n5582), .ZN(n5583) );
  NAND2_X1 U7137 ( .A1(n8647), .A2(n8653), .ZN(n8141) );
  NAND2_X1 U7138 ( .A1(n8647), .A2(n9026), .ZN(n9020) );
  XNOR2_X1 U7139 ( .A(n5586), .B(n5585), .ZN(n7312) );
  NAND2_X1 U7140 ( .A1(n7312), .A2(n8198), .ZN(n5590) );
  NAND2_X1 U7141 ( .A1(n5587), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5588) );
  XNOR2_X1 U7142 ( .A(n5588), .B(P2_IR_REG_17__SCAN_IN), .ZN(n8841) );
  AOI22_X1 U7143 ( .A1(n5619), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n6655), .B2(
        n8841), .ZN(n5589) );
  AOI22_X1 U7144 ( .A1(n5635), .A2(P2_REG2_REG_17__SCAN_IN), .B1(n5776), .B2(
        P2_REG1_REG_17__SCAN_IN), .ZN(n5594) );
  NAND2_X1 U7145 ( .A1(n5591), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n5592) );
  NAND2_X1 U7146 ( .A1(n5605), .A2(n5592), .ZN(n9030) );
  AOI22_X1 U7147 ( .A1(n5346), .A2(n9030), .B1(n5775), .B2(
        P2_REG0_REG_17__SCAN_IN), .ZN(n5593) );
  NAND2_X1 U7148 ( .A1(n9153), .A2(n9005), .ZN(n8053) );
  NAND2_X1 U7149 ( .A1(n8243), .A2(n8053), .ZN(n9018) );
  INV_X1 U7150 ( .A(n9005), .ZN(n8731) );
  NAND2_X1 U7151 ( .A1(n9153), .A2(n8731), .ZN(n5596) );
  XNOR2_X1 U7152 ( .A(n5598), .B(n5597), .ZN(n7426) );
  NAND2_X1 U7153 ( .A1(n7426), .A2(n8198), .ZN(n5604) );
  NAND2_X1 U7154 ( .A1(n5742), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5601) );
  INV_X1 U7155 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n5600) );
  NAND2_X1 U7156 ( .A1(n5601), .A2(n5600), .ZN(n5616) );
  OR2_X1 U7157 ( .A1(n5601), .A2(n5600), .ZN(n5602) );
  AND2_X1 U7158 ( .A1(n5616), .A2(n5602), .ZN(n8865) );
  AOI22_X1 U7159 ( .A1(n5619), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n6655), .B2(
        n8865), .ZN(n5603) );
  NAND2_X1 U7160 ( .A1(n5605), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n5606) );
  NAND2_X1 U7161 ( .A1(n5622), .A2(n5606), .ZN(n9012) );
  NAND2_X1 U7162 ( .A1(n9012), .A2(n5346), .ZN(n5610) );
  NAND2_X1 U7163 ( .A1(n5635), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n5609) );
  NAND2_X1 U7164 ( .A1(n5776), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n5608) );
  NAND2_X1 U7165 ( .A1(n5348), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n5607) );
  NAND4_X1 U7166 ( .A1(n5610), .A2(n5609), .A3(n5608), .A4(n5607), .ZN(n9024)
         );
  OR2_X1 U7167 ( .A1(n8699), .A2(n9024), .ZN(n5611) );
  NAND2_X1 U7168 ( .A1(n9002), .A2(n5611), .ZN(n5613) );
  NAND2_X1 U7169 ( .A1(n8699), .A2(n9024), .ZN(n5612) );
  XNOR2_X1 U7170 ( .A(n5615), .B(n5614), .ZN(n7511) );
  NAND2_X1 U7171 ( .A1(n7511), .A2(n8198), .ZN(n5621) );
  NAND2_X1 U7172 ( .A1(n5616), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5618) );
  AOI22_X1 U7173 ( .A1(n5619), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n8873), .B2(
        n6655), .ZN(n5620) );
  NAND2_X1 U7174 ( .A1(n5622), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n5623) );
  NAND2_X1 U7175 ( .A1(n5633), .A2(n5623), .ZN(n8996) );
  NAND2_X1 U7176 ( .A1(n8996), .A2(n5346), .ZN(n5626) );
  AOI22_X1 U7177 ( .A1(n5635), .A2(P2_REG2_REG_19__SCAN_IN), .B1(n5776), .B2(
        P2_REG1_REG_19__SCAN_IN), .ZN(n5625) );
  NAND2_X1 U7178 ( .A1(n5348), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n5624) );
  NAND2_X1 U7179 ( .A1(n9067), .A2(n9007), .ZN(n8151) );
  NAND2_X1 U7180 ( .A1(n8150), .A2(n8151), .ZN(n8991) );
  INV_X1 U7181 ( .A(n9007), .ZN(n8981) );
  XNOR2_X1 U7182 ( .A(n5628), .B(n5627), .ZN(n5629) );
  XNOR2_X1 U7183 ( .A(n5630), .B(n5629), .ZN(n7526) );
  NAND2_X1 U7184 ( .A1(n7526), .A2(n8198), .ZN(n5632) );
  INV_X1 U7185 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n7554) );
  OR2_X1 U7186 ( .A1(n4507), .A2(n7554), .ZN(n5631) );
  NAND2_X1 U7187 ( .A1(n5633), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n5634) );
  NAND2_X1 U7188 ( .A1(n5645), .A2(n5634), .ZN(n8985) );
  NAND2_X1 U7189 ( .A1(n8985), .A2(n5346), .ZN(n5638) );
  AOI22_X1 U7190 ( .A1(n5635), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n5776), .B2(
        P2_REG1_REG_20__SCAN_IN), .ZN(n5637) );
  NAND2_X1 U7191 ( .A1(n5775), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n5636) );
  NAND2_X1 U7192 ( .A1(n9137), .A2(n8995), .ZN(n8965) );
  INV_X1 U7193 ( .A(n8995), .ZN(n8972) );
  OR2_X1 U7194 ( .A1(n9137), .A2(n8972), .ZN(n8969) );
  XNOR2_X1 U7195 ( .A(n5640), .B(SI_21_), .ZN(n5641) );
  XNOR2_X1 U7196 ( .A(n5642), .B(n5641), .ZN(n7600) );
  NAND2_X1 U7197 ( .A1(n7600), .A2(n8198), .ZN(n5644) );
  OR2_X1 U7198 ( .A1(n4507), .A2(n7616), .ZN(n5643) );
  NAND2_X1 U7199 ( .A1(n5645), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n5646) );
  NAND2_X1 U7200 ( .A1(n5668), .A2(n5646), .ZN(n8975) );
  INV_X1 U7201 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n8974) );
  NAND2_X1 U7202 ( .A1(n5775), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n5648) );
  NAND2_X1 U7203 ( .A1(n5776), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n5647) );
  OAI211_X1 U7204 ( .C1(n7535), .C2(n8974), .A(n5648), .B(n5647), .ZN(n5649)
         );
  AOI21_X1 U7205 ( .B1(n8975), .B2(n5346), .A(n5649), .ZN(n8678) );
  NAND2_X1 U7206 ( .A1(n9131), .A2(n8678), .ZN(n8157) );
  NAND2_X1 U7207 ( .A1(n8049), .A2(n8157), .ZN(n8968) );
  OR2_X1 U7208 ( .A1(n9131), .A2(n8982), .ZN(n8954) );
  NAND2_X1 U7209 ( .A1(n8952), .A2(n8954), .ZN(n5659) );
  XNOR2_X1 U7210 ( .A(n5651), .B(n5650), .ZN(n7756) );
  NAND2_X1 U7211 ( .A1(n7756), .A2(n8198), .ZN(n5653) );
  OR2_X1 U7212 ( .A1(n4507), .A2(n7757), .ZN(n5652) );
  XNOR2_X1 U7213 ( .A(n5668), .B(P2_REG3_REG_22__SCAN_IN), .ZN(n8961) );
  NAND2_X1 U7214 ( .A1(n8961), .A2(n5346), .ZN(n5658) );
  INV_X1 U7215 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n8960) );
  NAND2_X1 U7216 ( .A1(n5775), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n5655) );
  NAND2_X1 U7217 ( .A1(n5776), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n5654) );
  OAI211_X1 U7218 ( .C1(n7535), .C2(n8960), .A(n5655), .B(n5654), .ZN(n5656)
         );
  INV_X1 U7219 ( .A(n5656), .ZN(n5657) );
  NAND2_X1 U7220 ( .A1(n9125), .A2(n8684), .ZN(n8045) );
  NAND2_X1 U7221 ( .A1(n8046), .A2(n8045), .ZN(n8953) );
  NAND2_X1 U7222 ( .A1(n5659), .A2(n8953), .ZN(n8957) );
  OR2_X1 U7223 ( .A1(n9125), .A2(n8971), .ZN(n5660) );
  NAND2_X1 U7224 ( .A1(n5663), .A2(n5662), .ZN(n5665) );
  NAND2_X1 U7225 ( .A1(n5665), .A2(n5664), .ZN(n7802) );
  NAND2_X1 U7226 ( .A1(n7802), .A2(n8198), .ZN(n5667) );
  OR2_X1 U7227 ( .A1(n4507), .A2(n7800), .ZN(n5666) );
  OAI21_X1 U7228 ( .B1(n5668), .B2(P2_REG3_REG_22__SCAN_IN), .A(
        P2_REG3_REG_23__SCAN_IN), .ZN(n5669) );
  NAND2_X1 U7229 ( .A1(n5669), .A2(n5682), .ZN(n8948) );
  NAND2_X1 U7230 ( .A1(n8948), .A2(n5346), .ZN(n5674) );
  INV_X1 U7231 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n8947) );
  NAND2_X1 U7232 ( .A1(n5348), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n5671) );
  NAND2_X1 U7233 ( .A1(n5776), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n5670) );
  OAI211_X1 U7234 ( .C1(n7535), .C2(n8947), .A(n5671), .B(n5670), .ZN(n5672)
         );
  INV_X1 U7235 ( .A(n5672), .ZN(n5673) );
  NAND2_X1 U7236 ( .A1(n9119), .A2(n8958), .ZN(n5675) );
  OR2_X1 U7237 ( .A1(n9119), .A2(n8958), .ZN(n5676) );
  XNOR2_X1 U7238 ( .A(n5679), .B(n5678), .ZN(n7898) );
  NAND2_X1 U7239 ( .A1(n7898), .A2(n8198), .ZN(n5681) );
  OR2_X1 U7240 ( .A1(n4507), .A2(n7908), .ZN(n5680) );
  NAND2_X1 U7241 ( .A1(n5682), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n5683) );
  NAND2_X1 U7242 ( .A1(n5696), .A2(n5683), .ZN(n8939) );
  NAND2_X1 U7243 ( .A1(n8939), .A2(n5346), .ZN(n5689) );
  INV_X1 U7244 ( .A(P2_REG2_REG_24__SCAN_IN), .ZN(n5686) );
  NAND2_X1 U7245 ( .A1(n5776), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n5685) );
  NAND2_X1 U7246 ( .A1(n5348), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n5684) );
  OAI211_X1 U7247 ( .C1(n5686), .C2(n7535), .A(n5685), .B(n5684), .ZN(n5687)
         );
  INV_X1 U7248 ( .A(n5687), .ZN(n5688) );
  NOR2_X1 U7249 ( .A1(n9113), .A2(n8945), .ZN(n5691) );
  NAND2_X1 U7250 ( .A1(n9113), .A2(n8945), .ZN(n5690) );
  XNOR2_X1 U7251 ( .A(n5692), .B(n5693), .ZN(n7918) );
  NAND2_X1 U7252 ( .A1(n7918), .A2(n8198), .ZN(n5695) );
  OR2_X1 U7253 ( .A1(n4507), .A2(n7933), .ZN(n5694) );
  NAND2_X1 U7254 ( .A1(n5696), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n5697) );
  NAND2_X1 U7255 ( .A1(n5708), .A2(n5697), .ZN(n8635) );
  NAND2_X1 U7256 ( .A1(n8635), .A2(n5346), .ZN(n5703) );
  INV_X1 U7257 ( .A(P2_REG2_REG_25__SCAN_IN), .ZN(n5700) );
  NAND2_X1 U7258 ( .A1(n5776), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n5699) );
  NAND2_X1 U7259 ( .A1(n5775), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n5698) );
  OAI211_X1 U7260 ( .C1(n7535), .C2(n5700), .A(n5699), .B(n5698), .ZN(n5701)
         );
  INV_X1 U7261 ( .A(n5701), .ZN(n5702) );
  NAND2_X1 U7262 ( .A1(n8628), .A2(n8667), .ZN(n8176) );
  NAND2_X1 U7263 ( .A1(n7949), .A2(n8198), .ZN(n5707) );
  OR2_X1 U7264 ( .A1(n4507), .A2(n7965), .ZN(n5706) );
  NAND2_X1 U7265 ( .A1(n5708), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n5709) );
  NAND2_X1 U7266 ( .A1(n5710), .A2(n5709), .ZN(n8917) );
  NAND2_X1 U7267 ( .A1(n8917), .A2(n5346), .ZN(n5715) );
  INV_X1 U7268 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n8916) );
  NAND2_X1 U7269 ( .A1(n5348), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n5712) );
  NAND2_X1 U7270 ( .A1(n5776), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n5711) );
  OAI211_X1 U7271 ( .C1(n7535), .C2(n8916), .A(n5712), .B(n5711), .ZN(n5713)
         );
  INV_X1 U7272 ( .A(n5713), .ZN(n5714) );
  NAND2_X1 U7273 ( .A1(n9102), .A2(n8901), .ZN(n5717) );
  NOR2_X1 U7274 ( .A1(n9102), .A2(n8901), .ZN(n5716) );
  AND2_X2 U7275 ( .A1(n8898), .A2(n8897), .ZN(n8899) );
  MUX2_X1 U7276 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(P2_DATAO_REG_28__SCAN_IN), 
        .S(n5217), .Z(n5732) );
  INV_X1 U7277 ( .A(SI_28_), .ZN(n10359) );
  XNOR2_X1 U7278 ( .A(n5732), .B(n10359), .ZN(n5730) );
  NAND2_X1 U7279 ( .A1(n8274), .A2(n8198), .ZN(n5721) );
  INV_X1 U7280 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n8275) );
  OR2_X1 U7281 ( .A1(n4507), .A2(n8275), .ZN(n5720) );
  NAND2_X1 U7282 ( .A1(n5722), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n5723) );
  NAND2_X1 U7283 ( .A1(n8883), .A2(n5723), .ZN(n8585) );
  NAND2_X1 U7284 ( .A1(n8585), .A2(n5346), .ZN(n5728) );
  INV_X1 U7285 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n6471) );
  NAND2_X1 U7286 ( .A1(n5775), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n5725) );
  NAND2_X1 U7287 ( .A1(n5776), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n5724) );
  OAI211_X1 U7288 ( .C1(n7535), .C2(n6471), .A(n5725), .B(n5724), .ZN(n5726)
         );
  INV_X1 U7289 ( .A(n5726), .ZN(n5727) );
  NAND2_X2 U7290 ( .A1(n5728), .A2(n5727), .ZN(n8902) );
  NOR2_X1 U7291 ( .A1(n8590), .A2(n8902), .ZN(n5729) );
  INV_X1 U7292 ( .A(n8902), .ZN(n8191) );
  INV_X1 U7293 ( .A(n8590), .ZN(n9089) );
  INV_X1 U7294 ( .A(n5732), .ZN(n5733) );
  INV_X1 U7295 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n9173) );
  INV_X1 U7296 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n10338) );
  MUX2_X1 U7297 ( .A(n9173), .B(n10338), .S(n5217), .Z(n6477) );
  NAND2_X1 U7298 ( .A1(n9170), .A2(n8198), .ZN(n5735) );
  OR2_X1 U7299 ( .A1(n4507), .A2(n9173), .ZN(n5734) );
  INV_X1 U7300 ( .A(n8883), .ZN(n5736) );
  NAND2_X1 U7301 ( .A1(n5736), .A2(n5346), .ZN(n7538) );
  INV_X1 U7302 ( .A(P2_REG2_REG_29__SCAN_IN), .ZN(n5739) );
  NAND2_X1 U7303 ( .A1(n5348), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n5738) );
  NAND2_X1 U7304 ( .A1(n5776), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n5737) );
  OAI211_X1 U7305 ( .C1(n7535), .C2(n5739), .A(n5738), .B(n5737), .ZN(n5740)
         );
  INV_X1 U7306 ( .A(n5740), .ZN(n5741) );
  NAND2_X1 U7307 ( .A1(n5824), .A2(n8584), .ZN(n8190) );
  NAND2_X1 U7308 ( .A1(n5748), .A2(n5743), .ZN(n5800) );
  NAND2_X1 U7309 ( .A1(n5800), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5744) );
  NAND2_X1 U7310 ( .A1(n8268), .A2(n8873), .ZN(n5819) );
  NAND2_X1 U7311 ( .A1(n5746), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5747) );
  MUX2_X1 U7312 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5747), .S(
        P2_IR_REG_20__SCAN_IN), .Z(n5750) );
  INV_X1 U7313 ( .A(n5748), .ZN(n5749) );
  NAND2_X1 U7314 ( .A1(n5750), .A2(n5749), .ZN(n8206) );
  INV_X1 U7315 ( .A(n8206), .ZN(n8205) );
  NAND2_X1 U7316 ( .A1(n6834), .A2(n8205), .ZN(n8260) );
  NAND2_X1 U7317 ( .A1(n7006), .A2(n8066), .ZN(n10140) );
  INV_X1 U7318 ( .A(n10146), .ZN(n10139) );
  NAND2_X1 U7319 ( .A1(n10140), .A2(n10139), .ZN(n10138) );
  INV_X1 U7320 ( .A(n10143), .ZN(n10160) );
  NAND2_X1 U7321 ( .A1(n7078), .A2(n10160), .ZN(n8068) );
  NAND2_X1 U7322 ( .A1(n10138), .A2(n8068), .ZN(n7281) );
  NAND2_X1 U7323 ( .A1(n5752), .A2(n10165), .ZN(n8084) );
  NAND2_X1 U7324 ( .A1(n10149), .A2(n5753), .ZN(n8076) );
  AND2_X1 U7325 ( .A1(n8084), .A2(n8076), .ZN(n8222) );
  NAND2_X1 U7326 ( .A1(n7281), .A2(n8222), .ZN(n5754) );
  NAND2_X1 U7327 ( .A1(n5754), .A2(n8084), .ZN(n7271) );
  INV_X1 U7328 ( .A(n5755), .ZN(n5757) );
  NAND2_X1 U7329 ( .A1(n7271), .A2(n8220), .ZN(n7270) );
  INV_X1 U7330 ( .A(n8742), .ZN(n7308) );
  NAND2_X1 U7331 ( .A1(n7308), .A2(n7273), .ZN(n8077) );
  NOR2_X1 U7332 ( .A1(n7458), .A2(n7435), .ZN(n8089) );
  NAND2_X1 U7333 ( .A1(n7458), .A2(n7435), .ZN(n8085) );
  NAND2_X1 U7334 ( .A1(n5758), .A2(n8085), .ZN(n7456) );
  AND2_X1 U7335 ( .A1(n8741), .A2(n10177), .ZN(n8091) );
  INV_X1 U7336 ( .A(n8741), .ZN(n7501) );
  INV_X1 U7337 ( .A(n10177), .ZN(n7462) );
  NAND2_X1 U7338 ( .A1(n7501), .A2(n7462), .ZN(n8081) );
  INV_X1 U7339 ( .A(n7507), .ZN(n10181) );
  NAND2_X1 U7340 ( .A1(n10181), .A2(n8740), .ZN(n8113) );
  INV_X1 U7341 ( .A(n8740), .ZN(n7540) );
  NAND2_X1 U7342 ( .A1(n7507), .A2(n7540), .ZN(n8100) );
  NAND2_X1 U7343 ( .A1(n8113), .A2(n8100), .ZN(n8096) );
  INV_X1 U7344 ( .A(n8738), .ZN(n7730) );
  NAND2_X1 U7345 ( .A1(n7645), .A2(n7730), .ZN(n8102) );
  NAND2_X1 U7346 ( .A1(n8115), .A2(n8102), .ZN(n8232) );
  INV_X1 U7347 ( .A(n7777), .ZN(n7785) );
  AND2_X1 U7348 ( .A1(n7785), .A2(n8737), .ZN(n8106) );
  AND2_X1 U7349 ( .A1(n7777), .A2(n7845), .ZN(n7790) );
  AOI21_X1 U7350 ( .B1(n10197), .B2(n7940), .A(n7790), .ZN(n8119) );
  OR2_X1 U7351 ( .A1(n10197), .A2(n7940), .ZN(n8108) );
  NAND2_X1 U7352 ( .A1(n5760), .A2(n8108), .ZN(n7856) );
  NAND2_X1 U7353 ( .A1(n7947), .A2(n7959), .ZN(n8056) );
  AND2_X2 U7354 ( .A1(n8057), .A2(n8056), .ZN(n8235) );
  INV_X1 U7355 ( .A(n8055), .ZN(n5761) );
  INV_X1 U7356 ( .A(n8734), .ZN(n8003) );
  OR2_X1 U7357 ( .A1(n8015), .A2(n8003), .ZN(n8130) );
  AND2_X1 U7358 ( .A1(n8015), .A2(n8003), .ZN(n8129) );
  INV_X1 U7359 ( .A(n8733), .ZN(n8542) );
  NAND2_X1 U7360 ( .A1(n8006), .A2(n8542), .ZN(n8143) );
  OR2_X1 U7361 ( .A1(n8006), .A2(n8542), .ZN(n8135) );
  NAND2_X1 U7362 ( .A1(n8031), .A2(n8141), .ZN(n9019) );
  NAND2_X1 U7363 ( .A1(n8699), .A2(n8994), .ZN(n8138) );
  NAND2_X1 U7364 ( .A1(n8245), .A2(n8138), .ZN(n9009) );
  INV_X1 U7365 ( .A(n8991), .ZN(n8989) );
  NAND2_X1 U7366 ( .A1(n8990), .A2(n8989), .ZN(n8988) );
  INV_X1 U7367 ( .A(n5762), .ZN(n8050) );
  AND2_X1 U7368 ( .A1(n8157), .A2(n8965), .ZN(n8052) );
  NAND2_X1 U7369 ( .A1(n5763), .A2(n8049), .ZN(n8951) );
  INV_X1 U7370 ( .A(n8046), .ZN(n5764) );
  AOI21_X1 U7371 ( .B1(n8951), .B2(n8045), .A(n5764), .ZN(n8942) );
  INV_X1 U7372 ( .A(n8958), .ZN(n8694) );
  NAND2_X1 U7373 ( .A1(n8942), .A2(n8219), .ZN(n8931) );
  NAND2_X1 U7374 ( .A1(n9113), .A2(n8925), .ZN(n8217) );
  NAND2_X1 U7375 ( .A1(n9119), .A2(n8694), .ZN(n8930) );
  AND2_X1 U7376 ( .A1(n8217), .A2(n8930), .ZN(n8167) );
  NAND2_X1 U7377 ( .A1(n8931), .A2(n8167), .ZN(n5765) );
  INV_X1 U7378 ( .A(n9102), .ZN(n8729) );
  INV_X1 U7379 ( .A(n8901), .ZN(n8924) );
  NAND2_X1 U7380 ( .A1(n9102), .A2(n8924), .ZN(n8043) );
  INV_X1 U7381 ( .A(n8897), .ZN(n5766) );
  OR2_X1 U7382 ( .A1(n9095), .A2(n8587), .ZN(n8179) );
  NAND2_X1 U7383 ( .A1(n5767), .A2(n8179), .ZN(n6466) );
  NAND2_X1 U7384 ( .A1(n6466), .A2(n8581), .ZN(n5769) );
  OR2_X1 U7385 ( .A1(n8590), .A2(n8191), .ZN(n5768) );
  NAND2_X1 U7386 ( .A1(n5769), .A2(n5768), .ZN(n8211) );
  NAND2_X1 U7387 ( .A1(n8206), .A2(n8859), .ZN(n6835) );
  NAND2_X1 U7388 ( .A1(n8268), .A2(n8859), .ZN(n6459) );
  NAND2_X1 U7389 ( .A1(n6459), .A2(n6835), .ZN(n5770) );
  NAND3_X1 U7390 ( .A1(n6899), .A2(n10187), .A3(n5770), .ZN(n10137) );
  INV_X1 U7391 ( .A(n8276), .ZN(n6920) );
  NAND2_X1 U7392 ( .A1(n6920), .A2(n8266), .ZN(n5773) );
  NAND2_X1 U7393 ( .A1(n5781), .A2(n5773), .ZN(n6842) );
  INV_X1 U7394 ( .A(n6842), .ZN(n5774) );
  INV_X1 U7395 ( .A(P2_REG2_REG_30__SCAN_IN), .ZN(n8888) );
  NAND2_X1 U7396 ( .A1(n5775), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n5778) );
  NAND2_X1 U7397 ( .A1(n5776), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n5777) );
  OAI211_X1 U7398 ( .C1(n7535), .C2(n8888), .A(n5778), .B(n5777), .ZN(n5779)
         );
  INV_X1 U7399 ( .A(n5779), .ZN(n5780) );
  NAND2_X1 U7400 ( .A1(n7538), .A2(n5780), .ZN(n8730) );
  AND2_X1 U7401 ( .A1(n5781), .A2(P2_B_REG_SCAN_IN), .ZN(n5782) );
  NOR2_X1 U7402 ( .A1(n9008), .A2(n5782), .ZN(n8881) );
  AOI22_X1 U7403 ( .A1(n9025), .A2(n8902), .B1(n8730), .B2(n8881), .ZN(n5783)
         );
  INV_X1 U7404 ( .A(n8895), .ZN(n5785) );
  AND2_X1 U7405 ( .A1(n6467), .A2(n7758), .ZN(n6829) );
  NAND2_X1 U7406 ( .A1(n5787), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5788) );
  MUX2_X1 U7407 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5788), .S(
        P2_IR_REG_24__SCAN_IN), .Z(n5789) );
  MUX2_X1 U7408 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5791), .S(
        P2_IR_REG_25__SCAN_IN), .Z(n5793) );
  NAND2_X1 U7409 ( .A1(n5794), .A2(n7935), .ZN(n5796) );
  NAND2_X1 U7410 ( .A1(n5792), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5795) );
  INV_X1 U7411 ( .A(n6667), .ZN(n5797) );
  INV_X1 U7412 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n6666) );
  NAND2_X1 U7413 ( .A1(n5797), .A2(n6666), .ZN(n5799) );
  INV_X1 U7414 ( .A(n5804), .ZN(n7967) );
  NAND2_X1 U7415 ( .A1(n7967), .A2(n7935), .ZN(n5798) );
  NAND2_X1 U7416 ( .A1(n7967), .A2(n7910), .ZN(n6668) );
  INV_X1 U7417 ( .A(n6833), .ZN(n6464) );
  NAND2_X1 U7418 ( .A1(n6664), .A2(n6464), .ZN(n6723) );
  INV_X1 U7419 ( .A(n6723), .ZN(n5817) );
  OAI21_X1 U7420 ( .B1(n5800), .B2(P2_IR_REG_22__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5802) );
  INV_X1 U7421 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n5801) );
  XNOR2_X1 U7422 ( .A(n5802), .B(n5801), .ZN(n7086) );
  AND2_X1 U7423 ( .A1(n7086), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6734) );
  INV_X1 U7424 ( .A(n7935), .ZN(n5805) );
  NAND3_X1 U7425 ( .A1(n5805), .A2(n5804), .A3(n5803), .ZN(n6726) );
  NOR2_X1 U7426 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .ZN(
        n5809) );
  NOR4_X1 U7427 ( .A1(P2_D_REG_4__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .A3(
        P2_D_REG_22__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n5808) );
  NOR4_X1 U7428 ( .A1(P2_D_REG_12__SCAN_IN), .A2(P2_D_REG_25__SCAN_IN), .A3(
        P2_D_REG_24__SCAN_IN), .A4(P2_D_REG_23__SCAN_IN), .ZN(n5807) );
  NOR4_X1 U7429 ( .A1(P2_D_REG_16__SCAN_IN), .A2(P2_D_REG_28__SCAN_IN), .A3(
        P2_D_REG_27__SCAN_IN), .A4(P2_D_REG_26__SCAN_IN), .ZN(n5806) );
  NAND4_X1 U7430 ( .A1(n5809), .A2(n5808), .A3(n5807), .A4(n5806), .ZN(n5815)
         );
  NOR4_X1 U7431 ( .A1(P2_D_REG_14__SCAN_IN), .A2(P2_D_REG_13__SCAN_IN), .A3(
        P2_D_REG_21__SCAN_IN), .A4(P2_D_REG_8__SCAN_IN), .ZN(n5813) );
  NOR4_X1 U7432 ( .A1(P2_D_REG_18__SCAN_IN), .A2(P2_D_REG_9__SCAN_IN), .A3(
        P2_D_REG_17__SCAN_IN), .A4(P2_D_REG_15__SCAN_IN), .ZN(n5812) );
  NOR4_X1 U7433 ( .A1(P2_D_REG_7__SCAN_IN), .A2(P2_D_REG_6__SCAN_IN), .A3(
        P2_D_REG_5__SCAN_IN), .A4(P2_D_REG_2__SCAN_IN), .ZN(n5811) );
  NOR4_X1 U7434 ( .A1(P2_D_REG_11__SCAN_IN), .A2(P2_D_REG_10__SCAN_IN), .A3(
        P2_D_REG_20__SCAN_IN), .A4(P2_D_REG_19__SCAN_IN), .ZN(n5810) );
  NAND4_X1 U7435 ( .A1(n5813), .A2(n5812), .A3(n5811), .A4(n5810), .ZN(n5814)
         );
  NOR2_X1 U7436 ( .A1(n5815), .A2(n5814), .ZN(n5816) );
  OR2_X1 U7437 ( .A1(n6667), .A2(n5816), .ZN(n6721) );
  AND3_X1 U7438 ( .A1(n5817), .A2(n6730), .A3(n6721), .ZN(n6741) );
  OR2_X1 U7439 ( .A1(n8258), .A2(n5819), .ZN(n6737) );
  NAND2_X1 U7440 ( .A1(n6899), .A2(n6737), .ZN(n5820) );
  NAND2_X1 U7441 ( .A1(n6741), .A2(n5820), .ZN(n5823) );
  NAND2_X1 U7442 ( .A1(n6833), .A2(n6721), .ZN(n5821) );
  NOR2_X1 U7443 ( .A1(n5821), .A2(n6664), .ZN(n6731) );
  AND2_X1 U7444 ( .A1(n6731), .A2(n6730), .ZN(n6844) );
  NAND3_X1 U7445 ( .A1(n8174), .A2(n6737), .A3(n10187), .ZN(n6735) );
  NAND2_X1 U7446 ( .A1(n6735), .A2(n10142), .ZN(n6722) );
  NAND2_X1 U7447 ( .A1(n6844), .A2(n6722), .ZN(n5822) );
  INV_X1 U7448 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n5825) );
  OAI21_X1 U7449 ( .B1(n6645), .B2(n10201), .A(n5827), .ZN(P2_U3456) );
  INV_X1 U7450 ( .A(n5871), .ZN(n5841) );
  NAND2_X1 U7451 ( .A1(n5842), .A2(n5841), .ZN(n6442) );
  NAND2_X1 U7452 ( .A1(n7756), .A2(n6501), .ZN(n5846) );
  NAND2_X1 U7453 ( .A1(n4673), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n5845) );
  NAND2_X1 U7454 ( .A1(n5851), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5852) );
  NAND2_X1 U7455 ( .A1(n5857), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5860) );
  NAND2_X1 U7456 ( .A1(n5860), .A2(n5858), .ZN(n5859) );
  NAND2_X1 U7457 ( .A1(n5861), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6305) );
  NAND2_X1 U7458 ( .A1(n6305), .A2(n5862), .ZN(n5863) );
  NAND2_X1 U7459 ( .A1(n4571), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5864) );
  NAND2_X1 U7460 ( .A1(n8456), .A2(n8504), .ZN(n8511) );
  NAND3_X1 U7461 ( .A1(n7103), .A2(n5866), .A3(n8511), .ZN(n5865) );
  OR2_X1 U7462 ( .A1(n7759), .A2(n4509), .ZN(n6582) );
  NAND3_X1 U7463 ( .A1(n6582), .A2(n7528), .A3(n5866), .ZN(n5867) );
  NAND2_X1 U7464 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n6000) );
  NAND2_X1 U7465 ( .A1(n6023), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n6045) );
  NAND2_X1 U7466 ( .A1(n6098), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n6141) );
  NAND2_X1 U7467 ( .A1(n6165), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n6206) );
  INV_X1 U7468 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n6205) );
  INV_X1 U7469 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n6232) );
  INV_X1 U7470 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n6308) );
  INV_X1 U7471 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n6295) );
  INV_X1 U7472 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n5888) );
  NAND2_X1 U7473 ( .A1(n5887), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n6335) );
  INV_X1 U7474 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n9340) );
  NAND2_X1 U7475 ( .A1(n6335), .A2(n9340), .ZN(n5868) );
  AND2_X1 U7476 ( .A1(n6349), .A2(n5868), .ZN(n9652) );
  INV_X1 U7477 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n5869) );
  XNOR2_X2 U7478 ( .A(n5873), .B(P1_IR_REG_29__SCAN_IN), .ZN(n5875) );
  NAND2_X4 U7479 ( .A1(n5876), .A2(n5875), .ZN(n6027) );
  NAND2_X1 U7480 ( .A1(n9652), .A2(n6577), .ZN(n5882) );
  INV_X1 U7481 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n5879) );
  NAND2_X2 U7482 ( .A1(n5874), .A2(n9901), .ZN(n5939) );
  NAND2_X1 U7483 ( .A1(n6872), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n5878) );
  AND2_X4 U7484 ( .A1(n5876), .A2(n9901), .ZN(n5961) );
  NAND2_X1 U7485 ( .A1(n5961), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n5877) );
  OAI211_X1 U7486 ( .C1(n4513), .C2(n5879), .A(n5878), .B(n5877), .ZN(n5880)
         );
  INV_X1 U7487 ( .A(n5880), .ZN(n5881) );
  AND2_X1 U7488 ( .A1(n8456), .A2(n7528), .ZN(n5883) );
  INV_X2 U7489 ( .A(n5905), .ZN(n6407) );
  OAI22_X1 U7490 ( .A1(n9654), .A2(n6619), .B1(n9233), .B2(n9207), .ZN(n5884)
         );
  XNOR2_X1 U7491 ( .A(n5884), .B(n4512), .ZN(n6346) );
  INV_X1 U7492 ( .A(n6346), .ZN(n9334) );
  NAND2_X1 U7493 ( .A1(n7526), .A2(n5910), .ZN(n5886) );
  NAND2_X1 U7494 ( .A1(n4673), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n5885) );
  NAND2_X1 U7495 ( .A1(n9688), .A2(n9206), .ZN(n5895) );
  INV_X1 U7496 ( .A(n5887), .ZN(n6333) );
  NAND2_X1 U7497 ( .A1(n6297), .A2(n5888), .ZN(n5889) );
  AND2_X1 U7498 ( .A1(n6333), .A2(n5889), .ZN(n9689) );
  NAND2_X1 U7499 ( .A1(n9689), .A2(n6577), .ZN(n5893) );
  AOI22_X1 U7500 ( .A1(n5900), .A2(P1_REG1_REG_20__SCAN_IN), .B1(n6872), .B2(
        P1_REG0_REG_20__SCAN_IN), .ZN(n5892) );
  NAND2_X1 U7501 ( .A1(n5961), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n5891) );
  OR2_X1 U7502 ( .A1(n9232), .A2(n9207), .ZN(n5894) );
  NAND2_X1 U7503 ( .A1(n5895), .A2(n5894), .ZN(n5896) );
  INV_X2 U7504 ( .A(n4512), .ZN(n9210) );
  XNOR2_X1 U7505 ( .A(n5896), .B(n9210), .ZN(n9313) );
  INV_X1 U7506 ( .A(n9313), .ZN(n6329) );
  NOR2_X1 U7507 ( .A1(n9232), .A2(n9214), .ZN(n5897) );
  AOI21_X1 U7508 ( .B1(n9688), .B2(n6407), .A(n5897), .ZN(n9312) );
  INV_X1 U7509 ( .A(n9312), .ZN(n6328) );
  INV_X1 U7510 ( .A(n5939), .ZN(n5898) );
  NAND2_X1 U7511 ( .A1(n5898), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n5904) );
  INV_X1 U7512 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n5899) );
  OR2_X1 U7513 ( .A1(n6027), .A2(n5899), .ZN(n5903) );
  NAND2_X1 U7514 ( .A1(n5900), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n5902) );
  NAND2_X1 U7515 ( .A1(n5961), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n5901) );
  NAND2_X1 U7516 ( .A1(n5914), .A2(n9212), .ZN(n5912) );
  INV_X1 U7517 ( .A(n5906), .ZN(n5907) );
  INV_X1 U7518 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n6658) );
  INV_X1 U7519 ( .A(n6675), .ZN(n5909) );
  NAND2_X1 U7520 ( .A1(n5912), .A2(n5911), .ZN(n5913) );
  AND2_X1 U7521 ( .A1(n6524), .A2(n6407), .ZN(n5915) );
  AOI21_X1 U7522 ( .B1(n5914), .B2(n6339), .A(n5915), .ZN(n5934) );
  XNOR2_X1 U7523 ( .A(n5933), .B(n5934), .ZN(n7092) );
  INV_X1 U7524 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n7106) );
  NAND2_X1 U7525 ( .A1(n5961), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n5919) );
  NAND2_X1 U7526 ( .A1(n5900), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n5918) );
  INV_X1 U7527 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n5916) );
  OR2_X1 U7528 ( .A1(n5939), .A2(n5916), .ZN(n5917) );
  NAND2_X1 U7529 ( .A1(n5927), .A2(n6407), .ZN(n5924) );
  INV_X1 U7530 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n10397) );
  NAND2_X1 U7531 ( .A1(n6671), .A2(SI_0_), .ZN(n5922) );
  INV_X1 U7532 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n5921) );
  XNOR2_X1 U7533 ( .A(n5922), .B(n5921), .ZN(n9906) );
  MUX2_X1 U7534 ( .A(n10397), .B(n9906), .S(n6768), .Z(n9994) );
  INV_X1 U7535 ( .A(n9994), .ZN(n7110) );
  NAND2_X1 U7536 ( .A1(n5924), .A2(n5923), .ZN(n5931) );
  INV_X1 U7537 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n9954) );
  NAND2_X1 U7538 ( .A1(n5927), .A2(n6339), .ZN(n5930) );
  OAI22_X1 U7539 ( .A1(n9994), .A2(n5905), .B1(n5925), .B2(n10397), .ZN(n5928)
         );
  INV_X1 U7540 ( .A(n5928), .ZN(n5929) );
  NAND2_X1 U7541 ( .A1(n5930), .A2(n5929), .ZN(n6893) );
  AOI21_X1 U7542 ( .B1(n6894), .B2(n6893), .A(n5932), .ZN(n7094) );
  NAND2_X1 U7543 ( .A1(n7092), .A2(n7094), .ZN(n7093) );
  INV_X1 U7544 ( .A(n5933), .ZN(n5935) );
  NAND2_X1 U7545 ( .A1(n5935), .A2(n5934), .ZN(n5936) );
  NAND2_X1 U7546 ( .A1(n7093), .A2(n5936), .ZN(n7185) );
  NAND2_X1 U7547 ( .A1(n5900), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n5943) );
  INV_X1 U7548 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n9433) );
  OR2_X1 U7549 ( .A1(n6027), .A2(n9433), .ZN(n5942) );
  INV_X1 U7550 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n5937) );
  INV_X1 U7551 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n5938) );
  NAND4_X2 U7552 ( .A1(n5943), .A2(n5942), .A3(n5941), .A4(n5940), .ZN(n7096)
         );
  NAND2_X1 U7553 ( .A1(n7096), .A2(n6407), .ZN(n5952) );
  OR2_X1 U7554 ( .A1(n6154), .A2(n6677), .ZN(n5950) );
  NOR2_X1 U7555 ( .A1(n5906), .A2(n5848), .ZN(n5944) );
  NAND2_X1 U7556 ( .A1(n5944), .A2(P1_IR_REG_2__SCAN_IN), .ZN(n5947) );
  INV_X1 U7557 ( .A(n5944), .ZN(n5946) );
  INV_X1 U7558 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n5945) );
  NAND2_X1 U7559 ( .A1(n5946), .A2(n5945), .ZN(n5967) );
  AND2_X1 U7560 ( .A1(n5947), .A2(n5967), .ZN(n9436) );
  NAND2_X1 U7561 ( .A1(n4823), .A2(n9436), .ZN(n5949) );
  INV_X1 U7562 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n6659) );
  OR2_X1 U7563 ( .A1(n5908), .A2(n6659), .ZN(n5948) );
  NAND2_X1 U7564 ( .A1(n5952), .A2(n5951), .ZN(n5953) );
  NAND2_X1 U7565 ( .A1(n7096), .A2(n6339), .ZN(n5955) );
  NAND2_X1 U7566 ( .A1(n7257), .A2(n9212), .ZN(n5954) );
  NAND2_X1 U7567 ( .A1(n5955), .A2(n5954), .ZN(n5956) );
  XNOR2_X1 U7568 ( .A(n5958), .B(n5956), .ZN(n7186) );
  NAND2_X1 U7569 ( .A1(n7185), .A2(n7186), .ZN(n5960) );
  INV_X1 U7570 ( .A(n5956), .ZN(n5957) );
  NAND2_X1 U7571 ( .A1(n5958), .A2(n5957), .ZN(n5959) );
  NAND2_X1 U7572 ( .A1(n5960), .A2(n5959), .ZN(n7287) );
  NAND2_X1 U7573 ( .A1(n5900), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n5966) );
  OR2_X1 U7574 ( .A1(n6027), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n5965) );
  INV_X1 U7575 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n6773) );
  OR2_X1 U7576 ( .A1(n6313), .A2(n6773), .ZN(n5964) );
  INV_X1 U7577 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n5962) );
  OR2_X1 U7578 ( .A1(n5939), .A2(n5962), .ZN(n5963) );
  NAND2_X1 U7579 ( .A1(n9421), .A2(n6407), .ZN(n5973) );
  INV_X1 U7580 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n6661) );
  OR2_X1 U7581 ( .A1(n5908), .A2(n6661), .ZN(n5971) );
  OR2_X1 U7582 ( .A1(n6154), .A2(n6673), .ZN(n5970) );
  NAND2_X1 U7583 ( .A1(n5967), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5968) );
  XNOR2_X1 U7584 ( .A(n5968), .B(P1_IR_REG_3__SCAN_IN), .ZN(n9451) );
  NAND2_X1 U7585 ( .A1(n4823), .A2(n9451), .ZN(n5969) );
  INV_X1 U7586 ( .A(n10017), .ZN(n7409) );
  NAND2_X1 U7587 ( .A1(n7409), .A2(n4797), .ZN(n5972) );
  NAND2_X1 U7588 ( .A1(n5973), .A2(n5972), .ZN(n5974) );
  XNOR2_X1 U7589 ( .A(n5974), .B(n9210), .ZN(n5979) );
  NAND2_X1 U7590 ( .A1(n9421), .A2(n6339), .ZN(n5976) );
  NAND2_X1 U7591 ( .A1(n7409), .A2(n6407), .ZN(n5975) );
  NAND2_X1 U7592 ( .A1(n5976), .A2(n5975), .ZN(n5977) );
  XNOR2_X1 U7593 ( .A(n5979), .B(n5977), .ZN(n7288) );
  NAND2_X1 U7594 ( .A1(n7287), .A2(n7288), .ZN(n5981) );
  INV_X1 U7595 ( .A(n5977), .ZN(n5978) );
  NAND2_X1 U7596 ( .A1(n5979), .A2(n5978), .ZN(n5980) );
  INV_X1 U7597 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n6792) );
  OR2_X1 U7598 ( .A1(n4513), .A2(n6792), .ZN(n5984) );
  OAI21_X1 U7599 ( .B1(P1_REG3_REG_4__SCAN_IN), .B2(P1_REG3_REG_3__SCAN_IN), 
        .A(n6000), .ZN(n7399) );
  OR2_X1 U7600 ( .A1(n6027), .A2(n7399), .ZN(n5983) );
  INV_X1 U7601 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n7395) );
  OR2_X1 U7602 ( .A1(n6313), .A2(n7395), .ZN(n5982) );
  NAND2_X1 U7603 ( .A1(n7416), .A2(n6407), .ZN(n5991) );
  INV_X1 U7604 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n6660) );
  OR2_X1 U7605 ( .A1(n5908), .A2(n6660), .ZN(n5989) );
  OR2_X1 U7606 ( .A1(n6154), .A2(n6676), .ZN(n5988) );
  OR2_X1 U7607 ( .A1(n6008), .A2(n5848), .ZN(n5986) );
  XNOR2_X1 U7608 ( .A(n5986), .B(P1_IR_REG_4__SCAN_IN), .ZN(n7023) );
  NAND2_X1 U7609 ( .A1(n4823), .A2(n7023), .ZN(n5987) );
  NAND2_X1 U7610 ( .A1(n7396), .A2(n4797), .ZN(n5990) );
  NAND2_X1 U7611 ( .A1(n5991), .A2(n5990), .ZN(n5992) );
  XNOR2_X1 U7612 ( .A(n5992), .B(n4512), .ZN(n5997) );
  NAND2_X1 U7613 ( .A1(n7416), .A2(n6339), .ZN(n5994) );
  NAND2_X1 U7614 ( .A1(n7396), .A2(n9212), .ZN(n5993) );
  NAND2_X1 U7615 ( .A1(n5994), .A2(n5993), .ZN(n5996) );
  XNOR2_X1 U7616 ( .A(n5997), .B(n5996), .ZN(n7346) );
  INV_X1 U7617 ( .A(n7346), .ZN(n5995) );
  NAND2_X1 U7618 ( .A1(n5997), .A2(n5996), .ZN(n5998) );
  NAND2_X1 U7619 ( .A1(n5900), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n6005) );
  INV_X1 U7620 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n5999) );
  OR2_X1 U7621 ( .A1(n5939), .A2(n5999), .ZN(n6004) );
  AND2_X1 U7622 ( .A1(n6000), .A2(n7520), .ZN(n6001) );
  OR2_X1 U7623 ( .A1(n6001), .A2(n6023), .ZN(n7525) );
  OR2_X1 U7624 ( .A1(n6027), .A2(n7525), .ZN(n6003) );
  INV_X1 U7625 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n7421) );
  OR2_X1 U7626 ( .A1(n6313), .A2(n7421), .ZN(n6002) );
  NAND4_X1 U7627 ( .A1(n6005), .A2(n6004), .A3(n6003), .A4(n6002), .ZN(n9420)
         );
  NAND2_X1 U7628 ( .A1(n9420), .A2(n9212), .ZN(n6014) );
  OR2_X1 U7629 ( .A1(n6154), .A2(n6681), .ZN(n6012) );
  INV_X1 U7630 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n6006) );
  OR2_X1 U7631 ( .A1(n5908), .A2(n6006), .ZN(n6011) );
  NAND2_X1 U7632 ( .A1(n6008), .A2(n6007), .ZN(n6018) );
  NAND2_X1 U7633 ( .A1(n6018), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6009) );
  XNOR2_X1 U7634 ( .A(n6009), .B(P1_IR_REG_5__SCAN_IN), .ZN(n9464) );
  NAND2_X1 U7635 ( .A1(n4823), .A2(n9464), .ZN(n6010) );
  NAND2_X1 U7636 ( .A1(n10031), .A2(n9206), .ZN(n6013) );
  NAND2_X1 U7637 ( .A1(n6014), .A2(n6013), .ZN(n6015) );
  XNOR2_X1 U7638 ( .A(n6015), .B(n4512), .ZN(n9377) );
  NAND2_X1 U7639 ( .A1(n9420), .A2(n6339), .ZN(n6017) );
  NAND2_X1 U7640 ( .A1(n10031), .A2(n9212), .ZN(n6016) );
  NAND2_X1 U7641 ( .A1(n6017), .A2(n6016), .ZN(n6035) );
  NAND2_X1 U7642 ( .A1(n6662), .A2(n6501), .ZN(n6021) );
  NAND2_X1 U7643 ( .A1(n6070), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6052) );
  XNOR2_X1 U7644 ( .A(n6052), .B(P1_IR_REG_6__SCAN_IN), .ZN(n6810) );
  NAND2_X1 U7645 ( .A1(n4823), .A2(n6810), .ZN(n6020) );
  NAND2_X1 U7646 ( .A1(n4673), .A2(P2_DATAO_REG_6__SCAN_IN), .ZN(n6019) );
  NAND2_X1 U7647 ( .A1(n5900), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n6031) );
  INV_X1 U7648 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n6022) );
  OR2_X1 U7649 ( .A1(n5939), .A2(n6022), .ZN(n6030) );
  INV_X1 U7650 ( .A(n6023), .ZN(n6025) );
  INV_X1 U7651 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n6024) );
  NAND2_X1 U7652 ( .A1(n6025), .A2(n6024), .ZN(n6026) );
  NAND2_X1 U7653 ( .A1(n6045), .A2(n6026), .ZN(n9382) );
  OR2_X1 U7654 ( .A1(n6027), .A2(n9382), .ZN(n6029) );
  INV_X1 U7655 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n7470) );
  OR2_X1 U7656 ( .A1(n6313), .A2(n7470), .ZN(n6028) );
  NAND4_X1 U7657 ( .A1(n6031), .A2(n6030), .A3(n6029), .A4(n6028), .ZN(n9419)
         );
  NAND2_X1 U7658 ( .A1(n9419), .A2(n9212), .ZN(n6032) );
  OAI21_X1 U7659 ( .B1(n10039), .B2(n6619), .A(n6032), .ZN(n6033) );
  XNOR2_X1 U7660 ( .A(n6033), .B(n4512), .ZN(n6036) );
  NAND2_X1 U7661 ( .A1(n9419), .A2(n6339), .ZN(n6034) );
  OAI21_X1 U7662 ( .B1(n10039), .B2(n9207), .A(n6034), .ZN(n6037) );
  INV_X1 U7663 ( .A(n6035), .ZN(n7518) );
  INV_X1 U7664 ( .A(n9377), .ZN(n7516) );
  NAND3_X1 U7665 ( .A1(n5148), .A2(n7518), .A3(n7516), .ZN(n6040) );
  INV_X1 U7666 ( .A(n6036), .ZN(n6039) );
  INV_X1 U7667 ( .A(n6037), .ZN(n6038) );
  NAND2_X1 U7668 ( .A1(n6039), .A2(n6038), .ZN(n9375) );
  AND2_X1 U7669 ( .A1(n6040), .A2(n9375), .ZN(n6041) );
  NAND2_X1 U7670 ( .A1(n6872), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n6051) );
  INV_X1 U7671 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n6043) );
  OR2_X1 U7672 ( .A1(n4513), .A2(n6043), .ZN(n6050) );
  NAND2_X1 U7673 ( .A1(n6045), .A2(n6044), .ZN(n6046) );
  NAND2_X1 U7674 ( .A1(n6079), .A2(n6046), .ZN(n9969) );
  OR2_X1 U7675 ( .A1(n6027), .A2(n9969), .ZN(n6049) );
  INV_X1 U7676 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n6047) );
  OR2_X1 U7677 ( .A1(n6313), .A2(n6047), .ZN(n6048) );
  NAND2_X1 U7678 ( .A1(n6678), .A2(n6501), .ZN(n6056) );
  NAND2_X1 U7679 ( .A1(n6052), .A2(n6067), .ZN(n6053) );
  NAND2_X1 U7680 ( .A1(n6053), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6054) );
  XNOR2_X1 U7681 ( .A(n6054), .B(P1_IR_REG_7__SCAN_IN), .ZN(n6821) );
  AOI22_X1 U7682 ( .A1(n4673), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n4823), .B2(
        n6821), .ZN(n6055) );
  NAND2_X1 U7683 ( .A1(n6056), .A2(n6055), .ZN(n7565) );
  NAND2_X1 U7684 ( .A1(n7565), .A2(n9206), .ZN(n6057) );
  OAI21_X1 U7685 ( .B1(n7668), .B2(n9207), .A(n6057), .ZN(n6058) );
  XNOR2_X1 U7686 ( .A(n6058), .B(n9210), .ZN(n6061) );
  OR2_X1 U7687 ( .A1(n7668), .A2(n9214), .ZN(n6060) );
  NAND2_X1 U7688 ( .A1(n7565), .A2(n9212), .ZN(n6059) );
  AND2_X1 U7689 ( .A1(n6060), .A2(n6059), .ZN(n6062) );
  NAND2_X1 U7690 ( .A1(n6061), .A2(n6062), .ZN(n6066) );
  INV_X1 U7691 ( .A(n6061), .ZN(n6064) );
  INV_X1 U7692 ( .A(n6062), .ZN(n6063) );
  NAND2_X1 U7693 ( .A1(n6064), .A2(n6063), .ZN(n6065) );
  AND2_X1 U7694 ( .A1(n6066), .A2(n6065), .ZN(n7558) );
  NAND2_X1 U7695 ( .A1(n7556), .A2(n7558), .ZN(n7557) );
  NAND2_X1 U7696 ( .A1(n6686), .A2(n6501), .ZN(n6077) );
  INV_X1 U7697 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n6068) );
  NAND2_X1 U7698 ( .A1(n6068), .A2(n6067), .ZN(n6069) );
  NOR2_X1 U7699 ( .A1(n6073), .A2(n5848), .ZN(n6071) );
  MUX2_X1 U7700 ( .A(n5848), .B(n6071), .S(P1_IR_REG_8__SCAN_IN), .Z(n6075) );
  INV_X1 U7701 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n6072) );
  NAND2_X1 U7702 ( .A1(n6073), .A2(n6072), .ZN(n6114) );
  INV_X1 U7703 ( .A(n6114), .ZN(n6074) );
  AOI22_X1 U7704 ( .A1(n4673), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n4823), .B2(
        n6860), .ZN(n6076) );
  NAND2_X1 U7705 ( .A1(n6077), .A2(n6076), .ZN(n9941) );
  NAND2_X1 U7706 ( .A1(n9941), .A2(n9206), .ZN(n6088) );
  NAND2_X1 U7707 ( .A1(n5900), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n6086) );
  NAND2_X1 U7708 ( .A1(n6079), .A2(n6078), .ZN(n6080) );
  NAND2_X1 U7709 ( .A1(n6099), .A2(n6080), .ZN(n9952) );
  OR2_X1 U7710 ( .A1(n6027), .A2(n9952), .ZN(n6085) );
  INV_X1 U7711 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n6081) );
  OR2_X1 U7712 ( .A1(n6313), .A2(n6081), .ZN(n6084) );
  INV_X1 U7713 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n6082) );
  OR2_X1 U7714 ( .A1(n5939), .A2(n6082), .ZN(n6083) );
  OR2_X1 U7715 ( .A1(n7717), .A2(n9207), .ZN(n6087) );
  NAND2_X1 U7716 ( .A1(n6088), .A2(n6087), .ZN(n6089) );
  XNOR2_X1 U7717 ( .A(n6089), .B(n4512), .ZN(n6092) );
  NAND2_X1 U7718 ( .A1(n9941), .A2(n9212), .ZN(n6091) );
  OR2_X1 U7719 ( .A1(n7717), .A2(n9214), .ZN(n6090) );
  AND2_X1 U7720 ( .A1(n6091), .A2(n6090), .ZN(n9940) );
  NAND2_X1 U7721 ( .A1(n9939), .A2(n9940), .ZN(n9296) );
  INV_X1 U7722 ( .A(n6092), .ZN(n6093) );
  NAND2_X1 U7723 ( .A1(n6094), .A2(n6093), .ZN(n9298) );
  NAND2_X1 U7724 ( .A1(n6114), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6095) );
  XNOR2_X1 U7725 ( .A(n6095), .B(P1_IR_REG_9__SCAN_IN), .ZN(n7040) );
  AOI22_X1 U7726 ( .A1(n4673), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n4823), .B2(
        n7040), .ZN(n6096) );
  NAND2_X1 U7727 ( .A1(n9306), .A2(n9206), .ZN(n6106) );
  NAND2_X1 U7728 ( .A1(n6872), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n6104) );
  INV_X1 U7729 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n6097) );
  OR2_X1 U7730 ( .A1(n4513), .A2(n6097), .ZN(n6103) );
  INV_X1 U7731 ( .A(n6098), .ZN(n6119) );
  NAND2_X1 U7732 ( .A1(n6099), .A2(n6866), .ZN(n6100) );
  NAND2_X1 U7733 ( .A1(n6119), .A2(n6100), .ZN(n9307) );
  OR2_X1 U7734 ( .A1(n6027), .A2(n9307), .ZN(n6102) );
  INV_X1 U7735 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n7721) );
  OR2_X1 U7736 ( .A1(n6313), .A2(n7721), .ZN(n6101) );
  OR2_X1 U7737 ( .A1(n7669), .A2(n9207), .ZN(n6105) );
  NAND2_X1 U7738 ( .A1(n6106), .A2(n6105), .ZN(n6107) );
  XNOR2_X1 U7739 ( .A(n6107), .B(n4512), .ZN(n6110) );
  NOR2_X1 U7740 ( .A1(n7669), .A2(n9214), .ZN(n6108) );
  AOI21_X1 U7741 ( .B1(n9306), .B2(n6407), .A(n6108), .ZN(n6111) );
  XNOR2_X1 U7742 ( .A(n6110), .B(n6111), .ZN(n9300) );
  AND2_X1 U7743 ( .A1(n9298), .A2(n9300), .ZN(n6109) );
  NAND2_X1 U7744 ( .A1(n9296), .A2(n6109), .ZN(n9299) );
  INV_X1 U7745 ( .A(n6110), .ZN(n6112) );
  OR2_X1 U7746 ( .A1(n6112), .A2(n6111), .ZN(n6113) );
  OR2_X1 U7747 ( .A1(n6696), .A2(n6154), .ZN(n6116) );
  NAND2_X1 U7748 ( .A1(n6157), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6135) );
  XNOR2_X1 U7749 ( .A(n6135), .B(P1_IR_REG_10__SCAN_IN), .ZN(n7226) );
  AOI22_X1 U7750 ( .A1(n4673), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n4823), .B2(
        n7226), .ZN(n6115) );
  NAND2_X1 U7751 ( .A1(n6116), .A2(n6115), .ZN(n7655) );
  NAND2_X1 U7752 ( .A1(n7655), .A2(n9206), .ZN(n6126) );
  NAND2_X1 U7753 ( .A1(n5900), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n6124) );
  INV_X1 U7754 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n7651) );
  OR2_X1 U7755 ( .A1(n6313), .A2(n7651), .ZN(n6123) );
  INV_X1 U7756 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n6117) );
  OR2_X1 U7757 ( .A1(n5939), .A2(n6117), .ZN(n6122) );
  INV_X1 U7758 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n6118) );
  NAND2_X1 U7759 ( .A1(n6119), .A2(n6118), .ZN(n6120) );
  NAND2_X1 U7760 ( .A1(n6141), .A2(n6120), .ZN(n9921) );
  OR2_X1 U7761 ( .A1(n6027), .A2(n9921), .ZN(n6121) );
  OR2_X1 U7762 ( .A1(n7740), .A2(n9207), .ZN(n6125) );
  NAND2_X1 U7763 ( .A1(n6126), .A2(n6125), .ZN(n6127) );
  XNOR2_X1 U7764 ( .A(n6127), .B(n4512), .ZN(n6128) );
  NAND2_X1 U7765 ( .A1(n6129), .A2(n6128), .ZN(n6130) );
  NAND2_X1 U7766 ( .A1(n7655), .A2(n9212), .ZN(n6132) );
  OR2_X1 U7767 ( .A1(n7740), .A2(n9214), .ZN(n6131) );
  NAND2_X1 U7768 ( .A1(n6132), .A2(n6131), .ZN(n9910) );
  NAND2_X1 U7769 ( .A1(n6712), .A2(n5910), .ZN(n6139) );
  INV_X1 U7770 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n6134) );
  NAND2_X1 U7771 ( .A1(n6135), .A2(n6134), .ZN(n6136) );
  NAND2_X1 U7772 ( .A1(n6136), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6137) );
  XNOR2_X1 U7773 ( .A(n6137), .B(P1_IR_REG_11__SCAN_IN), .ZN(n7360) );
  AOI22_X1 U7774 ( .A1(n4673), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n4823), .B2(
        n7360), .ZN(n6138) );
  NAND2_X1 U7775 ( .A1(n7765), .A2(n9206), .ZN(n6148) );
  NAND2_X1 U7776 ( .A1(n6872), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n6146) );
  NAND2_X1 U7777 ( .A1(n6141), .A2(n6140), .ZN(n6142) );
  NAND2_X1 U7778 ( .A1(n6167), .A2(n6142), .ZN(n9352) );
  OR2_X1 U7779 ( .A1(n6027), .A2(n9352), .ZN(n6145) );
  INV_X1 U7780 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n7227) );
  OR2_X1 U7781 ( .A1(n4513), .A2(n7227), .ZN(n6144) );
  INV_X1 U7782 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n7748) );
  OR2_X1 U7783 ( .A1(n6313), .A2(n7748), .ZN(n6143) );
  OR2_X1 U7784 ( .A1(n7807), .A2(n9207), .ZN(n6147) );
  NAND2_X1 U7785 ( .A1(n6148), .A2(n6147), .ZN(n6149) );
  XNOR2_X1 U7786 ( .A(n6149), .B(n9210), .ZN(n6152) );
  NOR2_X1 U7787 ( .A1(n7807), .A2(n9214), .ZN(n6150) );
  AOI21_X1 U7788 ( .B1(n7765), .B2(n6407), .A(n6150), .ZN(n6151) );
  NAND2_X1 U7789 ( .A1(n6152), .A2(n6151), .ZN(n9239) );
  OR2_X1 U7790 ( .A1(n6152), .A2(n6151), .ZN(n6153) );
  AND2_X1 U7791 ( .A1(n9239), .A2(n6153), .ZN(n9347) );
  NAND2_X1 U7792 ( .A1(n9238), .A2(n9239), .ZN(n6180) );
  OR2_X1 U7793 ( .A1(n6720), .A2(n6154), .ZN(n6164) );
  INV_X1 U7794 ( .A(n6155), .ZN(n6156) );
  NAND2_X1 U7795 ( .A1(n6161), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6159) );
  MUX2_X1 U7796 ( .A(n6159), .B(P1_IR_REG_31__SCAN_IN), .S(n6158), .Z(n6160)
         );
  INV_X1 U7797 ( .A(n6160), .ZN(n6162) );
  NOR2_X1 U7798 ( .A1(n6162), .A2(n6202), .ZN(n7358) );
  AOI22_X1 U7799 ( .A1(n4673), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n4823), .B2(
        n7358), .ZN(n6163) );
  NAND2_X1 U7800 ( .A1(n7842), .A2(n9206), .ZN(n6174) );
  NAND2_X1 U7801 ( .A1(n6872), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n6172) );
  INV_X1 U7802 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n7487) );
  OR2_X1 U7803 ( .A1(n4513), .A2(n7487), .ZN(n6171) );
  INV_X1 U7804 ( .A(n6165), .ZN(n6186) );
  NAND2_X1 U7805 ( .A1(n6167), .A2(n6166), .ZN(n6168) );
  NAND2_X1 U7806 ( .A1(n6186), .A2(n6168), .ZN(n9245) );
  OR2_X1 U7807 ( .A1(n6027), .A2(n9245), .ZN(n6170) );
  INV_X1 U7808 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n7814) );
  OR2_X1 U7809 ( .A1(n6313), .A2(n7814), .ZN(n6169) );
  OR2_X1 U7810 ( .A1(n7824), .A2(n9207), .ZN(n6173) );
  NAND2_X1 U7811 ( .A1(n6174), .A2(n6173), .ZN(n6175) );
  XNOR2_X1 U7812 ( .A(n6175), .B(n9210), .ZN(n6178) );
  NOR2_X1 U7813 ( .A1(n7824), .A2(n9214), .ZN(n6176) );
  AOI21_X1 U7814 ( .B1(n7842), .B2(n6407), .A(n6176), .ZN(n6177) );
  NAND2_X1 U7815 ( .A1(n6178), .A2(n6177), .ZN(n6181) );
  OR2_X1 U7816 ( .A1(n6178), .A2(n6177), .ZN(n6179) );
  AND2_X1 U7817 ( .A1(n6181), .A2(n6179), .ZN(n9240) );
  NAND2_X1 U7818 ( .A1(n9242), .A2(n6181), .ZN(n9322) );
  NAND2_X1 U7819 ( .A1(n6849), .A2(n5910), .ZN(n6184) );
  OR2_X1 U7820 ( .A1(n6202), .A2(n5848), .ZN(n6182) );
  XNOR2_X1 U7821 ( .A(n6182), .B(P1_IR_REG_13__SCAN_IN), .ZN(n7607) );
  AOI22_X1 U7822 ( .A1(n4673), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n4823), .B2(
        n7607), .ZN(n6183) );
  NAND2_X1 U7823 ( .A1(n7873), .A2(n9206), .ZN(n6194) );
  NAND2_X1 U7824 ( .A1(n5900), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n6192) );
  INV_X1 U7825 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n7829) );
  OR2_X1 U7826 ( .A1(n6313), .A2(n7829), .ZN(n6191) );
  INV_X1 U7827 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n6185) );
  NAND2_X1 U7828 ( .A1(n6186), .A2(n6185), .ZN(n6187) );
  NAND2_X1 U7829 ( .A1(n6206), .A2(n6187), .ZN(n9327) );
  OR2_X1 U7830 ( .A1(n6027), .A2(n9327), .ZN(n6190) );
  INV_X1 U7831 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n6188) );
  OR2_X1 U7832 ( .A1(n5939), .A2(n6188), .ZN(n6189) );
  OR2_X1 U7833 ( .A1(n9177), .A2(n9207), .ZN(n6193) );
  NAND2_X1 U7834 ( .A1(n6194), .A2(n6193), .ZN(n6195) );
  XNOR2_X1 U7835 ( .A(n6195), .B(n4512), .ZN(n6197) );
  NOR2_X1 U7836 ( .A1(n9177), .A2(n9214), .ZN(n6196) );
  AOI21_X1 U7837 ( .B1(n7873), .B2(n6407), .A(n6196), .ZN(n6198) );
  XNOR2_X1 U7838 ( .A(n6197), .B(n6198), .ZN(n9324) );
  INV_X1 U7839 ( .A(n6197), .ZN(n6199) );
  NAND2_X1 U7840 ( .A1(n6199), .A2(n6198), .ZN(n6200) );
  NAND2_X1 U7841 ( .A1(n9323), .A2(n6200), .ZN(n6218) );
  INV_X1 U7842 ( .A(n6218), .ZN(n6216) );
  NAND2_X1 U7843 ( .A1(n6889), .A2(n5910), .ZN(n6204) );
  NAND2_X1 U7844 ( .A1(n6202), .A2(n6201), .ZN(n6250) );
  NAND2_X1 U7845 ( .A1(n6250), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6225) );
  XNOR2_X1 U7846 ( .A(n6225), .B(P1_IR_REG_14__SCAN_IN), .ZN(n7887) );
  AOI22_X1 U7847 ( .A1(n4673), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n4823), .B2(
        n7887), .ZN(n6203) );
  NAND2_X1 U7848 ( .A1(n10073), .A2(n9206), .ZN(n6213) );
  NAND2_X1 U7849 ( .A1(n6872), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n6211) );
  INV_X1 U7850 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n7608) );
  OR2_X1 U7851 ( .A1(n4513), .A2(n7608), .ZN(n6210) );
  INV_X1 U7852 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n9757) );
  OR2_X1 U7853 ( .A1(n6313), .A2(n9757), .ZN(n6209) );
  NAND2_X1 U7854 ( .A1(n6206), .A2(n6205), .ZN(n6207) );
  NAND2_X1 U7855 ( .A1(n6233), .A2(n6207), .ZN(n9756) );
  OR2_X1 U7856 ( .A1(n6027), .A2(n9756), .ZN(n6208) );
  OR2_X1 U7857 ( .A1(n7927), .A2(n9207), .ZN(n6212) );
  NAND2_X1 U7858 ( .A1(n6213), .A2(n6212), .ZN(n6214) );
  XNOR2_X1 U7859 ( .A(n6214), .B(n9210), .ZN(n6217) );
  NAND2_X1 U7860 ( .A1(n6216), .A2(n6215), .ZN(n6219) );
  NAND2_X1 U7861 ( .A1(n6218), .A2(n6217), .ZN(n6223) );
  NAND2_X1 U7862 ( .A1(n10073), .A2(n6407), .ZN(n6221) );
  OR2_X1 U7863 ( .A1(n7927), .A2(n9214), .ZN(n6220) );
  NAND2_X1 U7864 ( .A1(n6221), .A2(n6220), .ZN(n9176) );
  NAND2_X1 U7865 ( .A1(n7032), .A2(n6501), .ZN(n6229) );
  INV_X1 U7866 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n6224) );
  NAND2_X1 U7867 ( .A1(n6225), .A2(n6224), .ZN(n6226) );
  NAND2_X1 U7868 ( .A1(n6226), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6227) );
  XNOR2_X1 U7869 ( .A(n6227), .B(P1_IR_REG_15__SCAN_IN), .ZN(n9483) );
  AOI22_X1 U7870 ( .A1(n4673), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n4823), .B2(
        n9483), .ZN(n6228) );
  NAND2_X1 U7871 ( .A1(n9396), .A2(n9206), .ZN(n6240) );
  NAND2_X1 U7872 ( .A1(n6872), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n6238) );
  INV_X1 U7873 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n6230) );
  OR2_X1 U7874 ( .A1(n4513), .A2(n6230), .ZN(n6237) );
  INV_X1 U7875 ( .A(n6231), .ZN(n6257) );
  NAND2_X1 U7876 ( .A1(n6233), .A2(n6232), .ZN(n6234) );
  NAND2_X1 U7877 ( .A1(n6257), .A2(n6234), .ZN(n9393) );
  OR2_X1 U7878 ( .A1(n6027), .A2(n9393), .ZN(n6236) );
  INV_X1 U7879 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n7921) );
  OR2_X1 U7880 ( .A1(n6313), .A2(n7921), .ZN(n6235) );
  OR2_X1 U7881 ( .A1(n9269), .A2(n9207), .ZN(n6239) );
  NAND2_X1 U7882 ( .A1(n6240), .A2(n6239), .ZN(n6241) );
  XNOR2_X1 U7883 ( .A(n6241), .B(n9210), .ZN(n6245) );
  NAND2_X1 U7884 ( .A1(n6244), .A2(n6245), .ZN(n9387) );
  NAND2_X1 U7885 ( .A1(n9396), .A2(n6407), .ZN(n6243) );
  OR2_X1 U7886 ( .A1(n9269), .A2(n9214), .ZN(n6242) );
  NAND2_X1 U7887 ( .A1(n6243), .A2(n6242), .ZN(n9390) );
  INV_X1 U7888 ( .A(n6244), .ZN(n6247) );
  INV_X1 U7889 ( .A(n6245), .ZN(n6246) );
  NAND2_X1 U7890 ( .A1(n7183), .A2(n6501), .ZN(n6253) );
  INV_X1 U7891 ( .A(n6248), .ZN(n6249) );
  OAI21_X1 U7892 ( .B1(n6250), .B2(n6249), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n6251) );
  XNOR2_X1 U7893 ( .A(n6251), .B(P1_IR_REG_16__SCAN_IN), .ZN(n8528) );
  AOI22_X1 U7894 ( .A1(n4673), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n4823), .B2(
        n8528), .ZN(n6252) );
  NAND2_X1 U7895 ( .A1(n9833), .A2(n9206), .ZN(n6265) );
  NAND2_X1 U7896 ( .A1(n5961), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n6263) );
  INV_X1 U7897 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n6254) );
  OR2_X1 U7898 ( .A1(n4513), .A2(n6254), .ZN(n6262) );
  INV_X1 U7899 ( .A(n6255), .ZN(n6279) );
  INV_X1 U7900 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n6256) );
  NAND2_X1 U7901 ( .A1(n6257), .A2(n6256), .ZN(n6258) );
  NAND2_X1 U7902 ( .A1(n6279), .A2(n6258), .ZN(n9923) );
  OR2_X1 U7903 ( .A1(n6027), .A2(n9923), .ZN(n6261) );
  INV_X1 U7904 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n6259) );
  OR2_X1 U7905 ( .A1(n5939), .A2(n6259), .ZN(n6260) );
  OR2_X1 U7906 ( .A1(n9279), .A2(n9207), .ZN(n6264) );
  NAND2_X1 U7907 ( .A1(n6265), .A2(n6264), .ZN(n6266) );
  XNOR2_X1 U7908 ( .A(n6266), .B(n4512), .ZN(n6269) );
  NAND2_X1 U7909 ( .A1(n9833), .A2(n6407), .ZN(n6268) );
  OR2_X1 U7910 ( .A1(n9279), .A2(n9214), .ZN(n6267) );
  NAND2_X1 U7911 ( .A1(n6268), .A2(n6267), .ZN(n6270) );
  NAND2_X1 U7912 ( .A1(n6269), .A2(n6270), .ZN(n9265) );
  INV_X1 U7913 ( .A(n6269), .ZN(n6272) );
  INV_X1 U7914 ( .A(n6270), .ZN(n6271) );
  NAND2_X1 U7915 ( .A1(n6272), .A2(n6271), .ZN(n9267) );
  NAND2_X1 U7916 ( .A1(n7312), .A2(n6501), .ZN(n6276) );
  NAND2_X1 U7917 ( .A1(n6273), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6274) );
  XNOR2_X1 U7918 ( .A(n6274), .B(P1_IR_REG_17__SCAN_IN), .ZN(n9501) );
  AOI22_X1 U7919 ( .A1(n4673), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n4823), .B2(
        n9501), .ZN(n6275) );
  NAND2_X2 U7920 ( .A1(n6276), .A2(n6275), .ZN(n9739) );
  NAND2_X1 U7921 ( .A1(n9739), .A2(n9206), .ZN(n6286) );
  NAND2_X1 U7922 ( .A1(n6872), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n6284) );
  INV_X1 U7923 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n6277) );
  OR2_X1 U7924 ( .A1(n4513), .A2(n6277), .ZN(n6283) );
  INV_X1 U7925 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n6278) );
  NAND2_X1 U7926 ( .A1(n6279), .A2(n6278), .ZN(n6280) );
  NAND2_X1 U7927 ( .A1(n6309), .A2(n6280), .ZN(n9740) );
  OR2_X1 U7928 ( .A1(n6027), .A2(n9740), .ZN(n6282) );
  INV_X1 U7929 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n9741) );
  OR2_X1 U7930 ( .A1(n6313), .A2(n9741), .ZN(n6281) );
  OR2_X1 U7931 ( .A1(n9367), .A2(n9207), .ZN(n6285) );
  NAND2_X1 U7932 ( .A1(n6286), .A2(n6285), .ZN(n6287) );
  XNOR2_X1 U7933 ( .A(n6287), .B(n4512), .ZN(n6289) );
  NOR2_X1 U7934 ( .A1(n9367), .A2(n9214), .ZN(n6288) );
  AOI21_X1 U7935 ( .B1(n9739), .B2(n6407), .A(n6288), .ZN(n6290) );
  XNOR2_X1 U7936 ( .A(n6289), .B(n6290), .ZN(n9277) );
  INV_X1 U7937 ( .A(n6289), .ZN(n6291) );
  NAND2_X1 U7938 ( .A1(n6291), .A2(n6290), .ZN(n6292) );
  NAND2_X1 U7939 ( .A1(n7511), .A2(n5910), .ZN(n6294) );
  AOI22_X1 U7940 ( .A1(n4673), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n4509), .B2(
        n4823), .ZN(n6293) );
  NAND2_X1 U7941 ( .A1(n6311), .A2(n6295), .ZN(n6296) );
  NAND2_X1 U7942 ( .A1(n6297), .A2(n6296), .ZN(n9698) );
  INV_X1 U7943 ( .A(P1_REG0_REG_19__SCAN_IN), .ZN(n6298) );
  OR2_X1 U7944 ( .A1(n5939), .A2(n6298), .ZN(n6300) );
  INV_X1 U7945 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n8530) );
  OR2_X1 U7946 ( .A1(n4513), .A2(n8530), .ZN(n6299) );
  AND2_X1 U7947 ( .A1(n6300), .A2(n6299), .ZN(n6302) );
  NAND2_X1 U7948 ( .A1(n5961), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n6301) );
  OAI211_X1 U7949 ( .C1(n9698), .C2(n6027), .A(n6302), .B(n6301), .ZN(n9406)
         );
  AOI22_X1 U7950 ( .A1(n9815), .A2(n9206), .B1(n6407), .B2(n9406), .ZN(n6303)
         );
  XNOR2_X1 U7951 ( .A(n6303), .B(n4512), .ZN(n9196) );
  AND2_X1 U7952 ( .A1(n9406), .A2(n6339), .ZN(n6304) );
  AOI21_X1 U7953 ( .B1(n9815), .B2(n6407), .A(n6304), .ZN(n9197) );
  NAND2_X1 U7954 ( .A1(n7426), .A2(n6501), .ZN(n6307) );
  XNOR2_X1 U7955 ( .A(n6305), .B(P1_IR_REG_18__SCAN_IN), .ZN(n9515) );
  AOI22_X1 U7956 ( .A1(n4673), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n4823), .B2(
        n9515), .ZN(n6306) );
  NAND2_X1 U7957 ( .A1(n9719), .A2(n9206), .ZN(n6319) );
  NAND2_X1 U7958 ( .A1(n6872), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n6317) );
  INV_X1 U7959 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n9823) );
  OR2_X1 U7960 ( .A1(n4513), .A2(n9823), .ZN(n6316) );
  NAND2_X1 U7961 ( .A1(n6309), .A2(n6308), .ZN(n6310) );
  NAND2_X1 U7962 ( .A1(n6311), .A2(n6310), .ZN(n9720) );
  OR2_X1 U7963 ( .A1(n9720), .A2(n6027), .ZN(n6315) );
  INV_X1 U7964 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n6312) );
  OR2_X1 U7965 ( .A1(n6313), .A2(n6312), .ZN(n6314) );
  NAND2_X1 U7966 ( .A1(n9407), .A2(n6407), .ZN(n6318) );
  NAND2_X1 U7967 ( .A1(n6319), .A2(n6318), .ZN(n6320) );
  XNOR2_X1 U7968 ( .A(n6320), .B(n4512), .ZN(n9195) );
  INV_X1 U7969 ( .A(n9195), .ZN(n6323) );
  NAND2_X1 U7970 ( .A1(n9719), .A2(n9212), .ZN(n6322) );
  NAND2_X1 U7971 ( .A1(n9407), .A2(n6339), .ZN(n6321) );
  NAND2_X1 U7972 ( .A1(n6322), .A2(n6321), .ZN(n9194) );
  INV_X1 U7973 ( .A(n9194), .ZN(n9361) );
  AOI22_X1 U7974 ( .A1(n9196), .A2(n9197), .B1(n6323), .B2(n9361), .ZN(n6327)
         );
  NAND2_X1 U7975 ( .A1(n9195), .A2(n9194), .ZN(n6324) );
  AOI21_X1 U7976 ( .B1(n9197), .B2(n6324), .A(n9196), .ZN(n6326) );
  NOR2_X1 U7977 ( .A1(n6324), .A2(n9197), .ZN(n6325) );
  NAND2_X1 U7978 ( .A1(n7600), .A2(n6501), .ZN(n6331) );
  NAND2_X1 U7979 ( .A1(n4673), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n6330) );
  INV_X1 U7980 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n6332) );
  NAND2_X1 U7981 ( .A1(n6333), .A2(n6332), .ZN(n6334) );
  NAND2_X1 U7982 ( .A1(n6335), .A2(n6334), .ZN(n9672) );
  OR2_X1 U7983 ( .A1(n9672), .A2(n6027), .ZN(n6338) );
  AOI22_X1 U7984 ( .A1(n5900), .A2(P1_REG1_REG_21__SCAN_IN), .B1(n6872), .B2(
        P1_REG0_REG_21__SCAN_IN), .ZN(n6337) );
  NAND2_X1 U7985 ( .A1(n5961), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n6336) );
  AOI22_X1 U7986 ( .A1(n9671), .A2(n6407), .B1(n6339), .B2(n9404), .ZN(n6345)
         );
  NAND2_X1 U7987 ( .A1(n9671), .A2(n9206), .ZN(n6341) );
  NAND2_X1 U7988 ( .A1(n9404), .A2(n6407), .ZN(n6340) );
  NAND2_X1 U7989 ( .A1(n6341), .A2(n6340), .ZN(n6342) );
  XNOR2_X1 U7990 ( .A(n6342), .B(n4512), .ZN(n6343) );
  XOR2_X1 U7991 ( .A(n6345), .B(n6343), .Z(n9230) );
  INV_X1 U7992 ( .A(n6343), .ZN(n6344) );
  OAI22_X2 U7993 ( .A1(n9231), .A2(n9230), .B1(n6345), .B2(n6344), .ZN(n9336)
         );
  OAI22_X1 U7994 ( .A1(n9654), .A2(n9207), .B1(n9233), .B2(n9214), .ZN(n9333)
         );
  NAND2_X1 U7995 ( .A1(n7802), .A2(n6501), .ZN(n6348) );
  NAND2_X1 U7996 ( .A1(n4673), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n6347) );
  NAND2_X1 U7997 ( .A1(n9791), .A2(n9206), .ZN(n6357) );
  INV_X1 U7998 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n9189) );
  INV_X1 U7999 ( .A(n6381), .ZN(n6379) );
  NAND2_X1 U8000 ( .A1(n6349), .A2(n9189), .ZN(n6350) );
  NAND2_X1 U8001 ( .A1(n6379), .A2(n6350), .ZN(n9639) );
  OR2_X1 U8002 ( .A1(n9639), .A2(n6027), .ZN(n6355) );
  INV_X1 U8003 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n9798) );
  NAND2_X1 U8004 ( .A1(n6872), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n6352) );
  NAND2_X1 U8005 ( .A1(n5961), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n6351) );
  OAI211_X1 U8006 ( .C1(n4513), .C2(n9798), .A(n6352), .B(n6351), .ZN(n6353)
         );
  INV_X1 U8007 ( .A(n6353), .ZN(n6354) );
  NAND2_X1 U8008 ( .A1(n9402), .A2(n6407), .ZN(n6356) );
  NAND2_X1 U8009 ( .A1(n6357), .A2(n6356), .ZN(n6358) );
  XNOR2_X1 U8010 ( .A(n6358), .B(n9210), .ZN(n6361) );
  NOR2_X1 U8011 ( .A1(n9339), .A2(n9214), .ZN(n6359) );
  AOI21_X1 U8012 ( .B1(n9791), .B2(n6407), .A(n6359), .ZN(n6360) );
  NAND2_X1 U8013 ( .A1(n6361), .A2(n6360), .ZN(n6362) );
  OAI21_X1 U8014 ( .B1(n6361), .B2(n6360), .A(n6362), .ZN(n9186) );
  INV_X1 U8015 ( .A(n6362), .ZN(n9287) );
  NAND2_X1 U8016 ( .A1(n4673), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n6363) );
  NAND2_X1 U8017 ( .A1(n9625), .A2(n9206), .ZN(n6370) );
  XNOR2_X1 U8018 ( .A(n6379), .B(P1_REG3_REG_24__SCAN_IN), .ZN(n9626) );
  NAND2_X1 U8019 ( .A1(n9626), .A2(n6577), .ZN(n6368) );
  INV_X1 U8020 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n9789) );
  NAND2_X1 U8021 ( .A1(n5961), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n6365) );
  NAND2_X1 U8022 ( .A1(n6872), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n6364) );
  OAI211_X1 U8023 ( .C1(n4513), .C2(n9789), .A(n6365), .B(n6364), .ZN(n6366)
         );
  INV_X1 U8024 ( .A(n6366), .ZN(n6367) );
  OR2_X1 U8025 ( .A1(n9256), .A2(n9207), .ZN(n6369) );
  NAND2_X1 U8026 ( .A1(n6370), .A2(n6369), .ZN(n6371) );
  XNOR2_X1 U8027 ( .A(n6371), .B(n9210), .ZN(n6374) );
  NOR2_X1 U8028 ( .A1(n9256), .A2(n9214), .ZN(n6372) );
  AOI21_X1 U8029 ( .B1(n9625), .B2(n6407), .A(n6372), .ZN(n6373) );
  NAND2_X1 U8030 ( .A1(n6374), .A2(n6373), .ZN(n6376) );
  OR2_X1 U8031 ( .A1(n6374), .A2(n6373), .ZN(n6375) );
  NAND2_X1 U8032 ( .A1(n7918), .A2(n6501), .ZN(n6378) );
  NAND2_X1 U8033 ( .A1(n4673), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n6377) );
  INV_X1 U8034 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n9291) );
  INV_X1 U8035 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n9258) );
  OAI21_X1 U8036 ( .B1(n6379), .B2(n9291), .A(n9258), .ZN(n6382) );
  AND2_X1 U8037 ( .A1(P1_REG3_REG_24__SCAN_IN), .A2(P1_REG3_REG_25__SCAN_IN), 
        .ZN(n6380) );
  INV_X1 U8038 ( .A(n6395), .ZN(n6396) );
  INV_X1 U8039 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n9784) );
  NAND2_X1 U8040 ( .A1(n5961), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n6384) );
  NAND2_X1 U8041 ( .A1(n6872), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n6383) );
  OAI211_X1 U8042 ( .C1(n4513), .C2(n9784), .A(n6384), .B(n6383), .ZN(n6385)
         );
  AOI21_X1 U8043 ( .B1(n9608), .B2(n6577), .A(n6385), .ZN(n9290) );
  OAI22_X1 U8044 ( .A1(n9861), .A2(n9207), .B1(n9290), .B2(n9214), .ZN(n6390)
         );
  NAND2_X1 U8045 ( .A1(n9609), .A2(n9206), .ZN(n6387) );
  OR2_X1 U8046 ( .A1(n9290), .A2(n9207), .ZN(n6386) );
  NAND2_X1 U8047 ( .A1(n6387), .A2(n6386), .ZN(n6388) );
  XNOR2_X1 U8048 ( .A(n6388), .B(n4512), .ZN(n6389) );
  XOR2_X1 U8049 ( .A(n6390), .B(n6389), .Z(n9254) );
  INV_X1 U8050 ( .A(n6389), .ZN(n6392) );
  INV_X1 U8051 ( .A(n6390), .ZN(n6391) );
  NAND2_X1 U8052 ( .A1(n6392), .A2(n6391), .ZN(n6408) );
  NAND2_X1 U8053 ( .A1(n7949), .A2(n5910), .ZN(n6394) );
  NAND2_X1 U8054 ( .A1(n4673), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n6393) );
  NAND2_X1 U8055 ( .A1(n9591), .A2(n9206), .ZN(n6404) );
  INV_X1 U8056 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n6448) );
  NAND2_X1 U8057 ( .A1(n6396), .A2(n6448), .ZN(n6397) );
  NAND2_X1 U8058 ( .A1(n6571), .A2(n6397), .ZN(n9592) );
  OR2_X1 U8059 ( .A1(n9592), .A2(n6027), .ZN(n6402) );
  INV_X1 U8060 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n9778) );
  NAND2_X1 U8061 ( .A1(n5961), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n6399) );
  NAND2_X1 U8062 ( .A1(n6872), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n6398) );
  OAI211_X1 U8063 ( .C1(n4513), .C2(n9778), .A(n6399), .B(n6398), .ZN(n6400)
         );
  INV_X1 U8064 ( .A(n6400), .ZN(n6401) );
  NAND2_X1 U8065 ( .A1(n9400), .A2(n9212), .ZN(n6403) );
  NAND2_X1 U8066 ( .A1(n6404), .A2(n6403), .ZN(n6405) );
  XNOR2_X1 U8067 ( .A(n6405), .B(n4512), .ZN(n6625) );
  NOR2_X1 U8068 ( .A1(n9257), .A2(n9214), .ZN(n6406) );
  AOI21_X1 U8069 ( .B1(n9591), .B2(n6407), .A(n6406), .ZN(n6626) );
  XNOR2_X1 U8070 ( .A(n6625), .B(n6626), .ZN(n6409) );
  INV_X1 U8071 ( .A(n6411), .ZN(n6414) );
  NAND2_X1 U8072 ( .A1(n7919), .A2(P1_B_REG_SCAN_IN), .ZN(n6412) );
  MUX2_X1 U8073 ( .A(P1_B_REG_SCAN_IN), .B(n6412), .S(n7899), .Z(n6413) );
  OR2_X1 U8074 ( .A1(n6714), .A2(P1_D_REG_0__SCAN_IN), .ZN(n6416) );
  NAND2_X1 U8075 ( .A1(n6411), .A2(n7899), .ZN(n6415) );
  OR2_X1 U8076 ( .A1(n6714), .A2(P1_D_REG_1__SCAN_IN), .ZN(n6417) );
  NAND2_X1 U8077 ( .A1(n6411), .A2(n7919), .ZN(n6715) );
  NOR4_X1 U8078 ( .A1(P1_D_REG_18__SCAN_IN), .A2(P1_D_REG_19__SCAN_IN), .A3(
        P1_D_REG_20__SCAN_IN), .A4(P1_D_REG_21__SCAN_IN), .ZN(n6421) );
  NOR4_X1 U8079 ( .A1(P1_D_REG_16__SCAN_IN), .A2(P1_D_REG_14__SCAN_IN), .A3(
        P1_D_REG_15__SCAN_IN), .A4(P1_D_REG_17__SCAN_IN), .ZN(n6420) );
  NOR4_X1 U8080 ( .A1(P1_D_REG_26__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n6419) );
  NOR4_X1 U8081 ( .A1(P1_D_REG_22__SCAN_IN), .A2(P1_D_REG_23__SCAN_IN), .A3(
        P1_D_REG_24__SCAN_IN), .A4(P1_D_REG_25__SCAN_IN), .ZN(n6418) );
  NAND4_X1 U8082 ( .A1(n6421), .A2(n6420), .A3(n6419), .A4(n6418), .ZN(n6427)
         );
  NOR2_X1 U8083 ( .A1(P1_D_REG_5__SCAN_IN), .A2(P1_D_REG_4__SCAN_IN), .ZN(
        n6425) );
  NOR4_X1 U8084 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        P1_D_REG_2__SCAN_IN), .A4(P1_D_REG_3__SCAN_IN), .ZN(n6424) );
  NOR4_X1 U8085 ( .A1(P1_D_REG_10__SCAN_IN), .A2(P1_D_REG_11__SCAN_IN), .A3(
        P1_D_REG_12__SCAN_IN), .A4(P1_D_REG_13__SCAN_IN), .ZN(n6423) );
  NOR4_X1 U8086 ( .A1(P1_D_REG_6__SCAN_IN), .A2(P1_D_REG_7__SCAN_IN), .A3(
        P1_D_REG_8__SCAN_IN), .A4(P1_D_REG_9__SCAN_IN), .ZN(n6422) );
  NAND4_X1 U8087 ( .A1(n6425), .A2(n6424), .A3(n6423), .A4(n6422), .ZN(n6426)
         );
  NOR2_X1 U8088 ( .A1(n6427), .A2(n6426), .ZN(n6428) );
  NAND3_X1 U8089 ( .A1(n9894), .A2(n7100), .A3(n6513), .ZN(n6446) );
  NAND2_X1 U8090 ( .A1(n6430), .A2(n6429), .ZN(n6431) );
  NAND2_X1 U8091 ( .A1(n6431), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6433) );
  INV_X1 U8092 ( .A(n7759), .ZN(n8515) );
  NAND2_X1 U8093 ( .A1(n8515), .A2(n8456), .ZN(n8498) );
  AND2_X1 U8094 ( .A1(n10067), .A2(n8498), .ZN(n6435) );
  NAND2_X1 U8095 ( .A1(n6631), .A2(n9948), .ZN(n6453) );
  INV_X1 U8096 ( .A(n9591), .ZN(n9857) );
  OR2_X1 U8097 ( .A1(n7103), .A2(n7528), .ZN(n7108) );
  INV_X1 U8098 ( .A(n7108), .ZN(n6436) );
  NAND2_X1 U8099 ( .A1(n6445), .A2(n6436), .ZN(n6437) );
  XNOR2_X1 U8100 ( .A(n6571), .B(P1_REG3_REG_27__SCAN_IN), .ZN(n9568) );
  INV_X1 U8101 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n6440) );
  NAND2_X1 U8102 ( .A1(n5961), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n6439) );
  NAND2_X1 U8103 ( .A1(n6872), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n6438) );
  OAI211_X1 U8104 ( .C1(n4513), .C2(n6440), .A(n6439), .B(n6438), .ZN(n6441)
         );
  INV_X1 U8105 ( .A(n8498), .ZN(n6766) );
  OR2_X1 U8106 ( .A1(n6622), .A2(n9338), .ZN(n6444) );
  OR2_X1 U8107 ( .A1(n9290), .A2(n9537), .ZN(n6443) );
  NAND2_X1 U8108 ( .A1(n6444), .A2(n6443), .ZN(n9587) );
  NAND2_X1 U8109 ( .A1(n6445), .A2(n8328), .ZN(n9221) );
  NOR2_X1 U8110 ( .A1(n8498), .A2(n8328), .ZN(n6512) );
  AOI21_X1 U8111 ( .B1(n6446), .B2(n6510), .A(n6512), .ZN(n6896) );
  NAND3_X1 U8112 ( .A1(n6896), .A2(n5925), .A3(n6769), .ZN(n6447) );
  OAI22_X1 U8113 ( .A1(n9592), .A2(n9920), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n6448), .ZN(n6449) );
  AOI21_X1 U8114 ( .B1(n9587), .B2(n4510), .A(n6449), .ZN(n6450) );
  OAI21_X1 U8115 ( .B1(n6454), .B2(n6453), .A(n6452), .ZN(P1_U3240) );
  NOR2_X1 U8116 ( .A1(n9008), .A2(n8584), .ZN(n6456) );
  INV_X1 U8117 ( .A(n9088), .ZN(n6476) );
  NAND2_X1 U8118 ( .A1(n8203), .A2(n6835), .ZN(n6725) );
  AND3_X1 U8119 ( .A1(n6730), .A2(n6721), .A3(n6725), .ZN(n6644) );
  OR2_X1 U8120 ( .A1(n6459), .A2(n8206), .ZN(n6460) );
  NAND2_X1 U8121 ( .A1(n6460), .A2(n8174), .ZN(n6462) );
  NAND2_X1 U8122 ( .A1(n6462), .A2(n6664), .ZN(n6461) );
  OAI21_X1 U8123 ( .B1(n6462), .B2(n6833), .A(n6461), .ZN(n6642) );
  INV_X1 U8124 ( .A(n6642), .ZN(n6463) );
  OAI211_X1 U8125 ( .C1(n6664), .C2(n6464), .A(n6644), .B(n6463), .ZN(n6470)
         );
  NAND2_X1 U8126 ( .A1(n6829), .A2(n5818), .ZN(n6643) );
  INV_X1 U8127 ( .A(n6643), .ZN(n6465) );
  XNOR2_X1 U8128 ( .A(n6466), .B(n8581), .ZN(n9090) );
  AND2_X1 U8129 ( .A1(n6467), .A2(n6834), .ZN(n7499) );
  INV_X1 U8130 ( .A(n7499), .ZN(n6468) );
  AND2_X1 U8131 ( .A1(n10137), .A2(n6468), .ZN(n6469) );
  OR2_X1 U8132 ( .A1(n6470), .A2(n10142), .ZN(n9014) );
  AOI22_X1 U8133 ( .A1(n8590), .A2(n9032), .B1(n9031), .B2(n8585), .ZN(n6472)
         );
  OAI21_X1 U8134 ( .B1(n9090), .B2(n9035), .A(n6473), .ZN(n6474) );
  INV_X1 U8135 ( .A(n6474), .ZN(n6475) );
  INV_X1 U8136 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n6516) );
  INV_X1 U8137 ( .A(SI_29_), .ZN(n10358) );
  INV_X1 U8138 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n8185) );
  INV_X1 U8139 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n10372) );
  MUX2_X1 U8140 ( .A(n8185), .B(n10372), .S(n5217), .Z(n6482) );
  INV_X1 U8141 ( .A(SI_30_), .ZN(n6481) );
  NAND2_X1 U8142 ( .A1(n6482), .A2(n6481), .ZN(n6485) );
  INV_X1 U8143 ( .A(n6482), .ZN(n6483) );
  NAND2_X1 U8144 ( .A1(n6483), .A2(SI_30_), .ZN(n6484) );
  NAND2_X1 U8145 ( .A1(n6485), .A2(n6484), .ZN(n6497) );
  INV_X1 U8146 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n9163) );
  INV_X1 U8147 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n6486) );
  MUX2_X1 U8148 ( .A(n9163), .B(n6486), .S(n5217), .Z(n6487) );
  XNOR2_X1 U8149 ( .A(n6487), .B(SI_31_), .ZN(n6488) );
  NAND2_X1 U8150 ( .A1(n9895), .A2(n5910), .ZN(n6491) );
  NAND2_X1 U8151 ( .A1(n4673), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(n6490) );
  NAND2_X1 U8152 ( .A1(n8274), .A2(n5910), .ZN(n6493) );
  NAND2_X1 U8153 ( .A1(n4673), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n6492) );
  INV_X1 U8154 ( .A(n9815), .ZN(n9701) );
  NAND2_X1 U8155 ( .A1(n7407), .A2(n10017), .ZN(n7406) );
  INV_X1 U8156 ( .A(n10039), .ZN(n7475) );
  NOR2_X2 U8157 ( .A1(n7709), .A2(n9306), .ZN(n7711) );
  AND2_X2 U8158 ( .A1(n7711), .A2(n10068), .ZN(n7652) );
  INV_X1 U8159 ( .A(n10073), .ZN(n9755) );
  NAND2_X1 U8160 ( .A1(n9754), .A2(n9892), .ZN(n9832) );
  NOR2_X2 U8161 ( .A1(n9671), .A2(n9686), .ZN(n9670) );
  NAND2_X1 U8162 ( .A1(n9654), .A2(n9670), .ZN(n9649) );
  NOR2_X2 U8163 ( .A1(n4531), .A2(n9625), .ZN(n9624) );
  NAND2_X1 U8164 ( .A1(n9861), .A2(n9624), .ZN(n9607) );
  NAND2_X1 U8165 ( .A1(n8273), .A2(n5910), .ZN(n6496) );
  NAND2_X1 U8166 ( .A1(n4673), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n6495) );
  NAND2_X1 U8167 ( .A1(n6498), .A2(n6497), .ZN(n6499) );
  NAND2_X1 U8168 ( .A1(n4673), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n6502) );
  XNOR2_X1 U8169 ( .A(n4648), .B(n6503), .ZN(n9523) );
  NAND2_X1 U8170 ( .A1(n5961), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n6505) );
  NAND2_X1 U8171 ( .A1(n6872), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n6504) );
  OAI211_X1 U8172 ( .C1(n4513), .C2(n6516), .A(n6505), .B(n6504), .ZN(n8493)
         );
  INV_X1 U8173 ( .A(P1_B_REG_SCAN_IN), .ZN(n6507) );
  NOR2_X1 U8174 ( .A1(n4508), .A2(n6507), .ZN(n6508) );
  OR2_X1 U8175 ( .A1(n9338), .A2(n6508), .ZN(n9535) );
  INV_X1 U8176 ( .A(n9535), .ZN(n6509) );
  AOI21_X1 U8177 ( .B1(n9523), .B2(n9993), .A(n9935), .ZN(n6519) );
  INV_X1 U8178 ( .A(n6510), .ZN(n6511) );
  NOR2_X1 U8179 ( .A1(n7100), .A2(n6511), .ZN(n6515) );
  NOR2_X1 U8180 ( .A1(n9893), .A2(n6512), .ZN(n6514) );
  MUX2_X1 U8181 ( .A(n6516), .B(n6519), .S(n10102), .Z(n6517) );
  NAND2_X1 U8182 ( .A1(n6517), .A2(n5147), .ZN(P1_U3553) );
  INV_X1 U8183 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n6520) );
  INV_X1 U8184 ( .A(n9894), .ZN(n7102) );
  MUX2_X1 U8185 ( .A(n6520), .B(n6519), .S(n10084), .Z(n6521) );
  NAND2_X1 U8186 ( .A1(n6521), .A2(n5146), .ZN(P1_U3521) );
  INV_X1 U8187 ( .A(n9556), .ZN(n6616) );
  AND2_X1 U8188 ( .A1(n5927), .A2(n7110), .ZN(n9980) );
  INV_X1 U8189 ( .A(n9980), .ZN(n6522) );
  NAND2_X1 U8190 ( .A1(n6523), .A2(n6522), .ZN(n6526) );
  OR2_X1 U8191 ( .A1(n5914), .A2(n6524), .ZN(n6525) );
  NAND2_X1 U8192 ( .A1(n6526), .A2(n6525), .ZN(n7260) );
  INV_X1 U8193 ( .A(n7257), .ZN(n10011) );
  NAND2_X1 U8194 ( .A1(n7096), .A2(n10011), .ZN(n8297) );
  NAND2_X1 U8195 ( .A1(n4659), .A2(n8297), .ZN(n8460) );
  NAND2_X1 U8196 ( .A1(n7260), .A2(n8460), .ZN(n6528) );
  OR2_X1 U8197 ( .A1(n7257), .A2(n7096), .ZN(n6527) );
  NAND2_X1 U8198 ( .A1(n6528), .A2(n6527), .ZN(n7405) );
  OR2_X1 U8199 ( .A1(n9421), .A2(n10017), .ZN(n8293) );
  NAND2_X1 U8200 ( .A1(n9421), .A2(n10017), .ZN(n8298) );
  NAND2_X1 U8201 ( .A1(n7405), .A2(n8459), .ZN(n6530) );
  OR2_X1 U8202 ( .A1(n7409), .A2(n9421), .ZN(n6529) );
  NAND2_X1 U8203 ( .A1(n6530), .A2(n6529), .ZN(n7390) );
  NOR2_X1 U8204 ( .A1(n7416), .A2(n10024), .ZN(n6587) );
  INV_X1 U8205 ( .A(n6587), .ZN(n8303) );
  NAND2_X1 U8206 ( .A1(n7416), .A2(n10024), .ZN(n8299) );
  NAND2_X1 U8207 ( .A1(n8303), .A2(n8299), .ZN(n8458) );
  NAND2_X1 U8208 ( .A1(n7390), .A2(n8458), .ZN(n6532) );
  OR2_X1 U8209 ( .A1(n7396), .A2(n7416), .ZN(n6531) );
  NAND2_X1 U8210 ( .A1(n6532), .A2(n6531), .ZN(n7414) );
  OR2_X1 U8211 ( .A1(n9420), .A2(n7420), .ZN(n8343) );
  AND2_X1 U8212 ( .A1(n9420), .A2(n7420), .ZN(n8344) );
  NAND2_X1 U8213 ( .A1(n8343), .A2(n8340), .ZN(n8461) );
  NAND2_X1 U8214 ( .A1(n7414), .A2(n8461), .ZN(n6534) );
  OR2_X1 U8215 ( .A1(n10031), .A2(n9420), .ZN(n6533) );
  NAND2_X1 U8216 ( .A1(n6534), .A2(n6533), .ZN(n7476) );
  NAND2_X1 U8217 ( .A1(n9419), .A2(n10039), .ZN(n8346) );
  NAND2_X1 U8218 ( .A1(n9963), .A2(n8346), .ZN(n7477) );
  NAND2_X1 U8219 ( .A1(n7476), .A2(n7477), .ZN(n6536) );
  OR2_X1 U8220 ( .A1(n7475), .A2(n9419), .ZN(n6535) );
  NAND2_X1 U8221 ( .A1(n7668), .A2(n7565), .ZN(n7665) );
  INV_X1 U8222 ( .A(n7668), .ZN(n9418) );
  NAND2_X1 U8223 ( .A1(n10043), .A2(n9418), .ZN(n6593) );
  NAND2_X1 U8224 ( .A1(n10043), .A2(n7668), .ZN(n6537) );
  OR2_X1 U8225 ( .A1(n9941), .A2(n7717), .ZN(n8354) );
  NAND2_X1 U8226 ( .A1(n9941), .A2(n7717), .ZN(n8355) );
  NAND2_X1 U8227 ( .A1(n8354), .A2(n8355), .ZN(n7663) );
  INV_X1 U8228 ( .A(n7717), .ZN(n9417) );
  INV_X1 U8229 ( .A(n7669), .ZN(n9416) );
  NAND2_X1 U8230 ( .A1(n9306), .A2(n7669), .ZN(n8362) );
  INV_X1 U8231 ( .A(n8362), .ZN(n6538) );
  NAND2_X1 U8232 ( .A1(n7720), .A2(n7719), .ZN(n6540) );
  OR2_X1 U8233 ( .A1(n9306), .A2(n9416), .ZN(n6539) );
  NAND2_X1 U8234 ( .A1(n6540), .A2(n6539), .ZN(n7656) );
  INV_X1 U8235 ( .A(n7740), .ZN(n9415) );
  NAND2_X1 U8236 ( .A1(n10068), .A2(n9415), .ZN(n8370) );
  NAND2_X1 U8237 ( .A1(n7655), .A2(n7740), .ZN(n8368) );
  NAND2_X1 U8238 ( .A1(n7656), .A2(n7657), .ZN(n6542) );
  NAND2_X1 U8239 ( .A1(n10068), .A2(n7740), .ZN(n6541) );
  INV_X1 U8240 ( .A(n7807), .ZN(n9414) );
  NOR2_X1 U8241 ( .A1(n7765), .A2(n9414), .ZN(n6543) );
  NAND2_X1 U8242 ( .A1(n7765), .A2(n9414), .ZN(n6544) );
  NOR2_X1 U8243 ( .A1(n7842), .A2(n7824), .ZN(n8373) );
  INV_X1 U8244 ( .A(n8373), .ZN(n8312) );
  NAND2_X1 U8245 ( .A1(n7842), .A2(n7824), .ZN(n8372) );
  NAND2_X1 U8246 ( .A1(n8312), .A2(n8372), .ZN(n8468) );
  INV_X1 U8247 ( .A(n7824), .ZN(n9413) );
  NAND2_X1 U8248 ( .A1(n7842), .A2(n9413), .ZN(n6545) );
  INV_X1 U8249 ( .A(n9177), .ZN(n9412) );
  NAND2_X1 U8250 ( .A1(n7873), .A2(n9412), .ZN(n6547) );
  INV_X1 U8251 ( .A(n7927), .ZN(n9411) );
  AND2_X1 U8252 ( .A1(n10073), .A2(n9411), .ZN(n6548) );
  INV_X1 U8253 ( .A(n9269), .ZN(n9410) );
  NOR2_X1 U8254 ( .A1(n9396), .A2(n9410), .ZN(n6549) );
  NAND2_X1 U8255 ( .A1(n9396), .A2(n9410), .ZN(n6550) );
  INV_X1 U8256 ( .A(n9833), .ZN(n9927) );
  INV_X1 U8257 ( .A(n9279), .ZN(n9409) );
  AND2_X1 U8258 ( .A1(n9927), .A2(n9409), .ZN(n8389) );
  INV_X1 U8259 ( .A(n8389), .ZN(n8396) );
  NAND2_X1 U8260 ( .A1(n9833), .A2(n9279), .ZN(n8398) );
  NAND2_X1 U8261 ( .A1(n8396), .A2(n8398), .ZN(n8473) );
  NAND2_X1 U8262 ( .A1(n9829), .A2(n8473), .ZN(n6552) );
  NAND2_X1 U8263 ( .A1(n9833), .A2(n9409), .ZN(n6551) );
  NAND2_X1 U8264 ( .A1(n6552), .A2(n6551), .ZN(n9735) );
  INV_X1 U8265 ( .A(n9367), .ZN(n9408) );
  AND2_X1 U8266 ( .A1(n9739), .A2(n9408), .ZN(n6554) );
  OR2_X1 U8267 ( .A1(n9739), .A2(n9408), .ZN(n6553) );
  NOR2_X1 U8268 ( .A1(n9719), .A2(n9407), .ZN(n6555) );
  NAND2_X1 U8269 ( .A1(n9719), .A2(n9407), .ZN(n6556) );
  INV_X1 U8270 ( .A(n9406), .ZN(n9316) );
  AND2_X1 U8271 ( .A1(n9815), .A2(n9316), .ZN(n8290) );
  INV_X1 U8272 ( .A(n8290), .ZN(n8411) );
  NAND2_X1 U8273 ( .A1(n8334), .A2(n8411), .ZN(n9702) );
  INV_X1 U8274 ( .A(n9232), .ZN(n9405) );
  AND2_X1 U8275 ( .A1(n9688), .A2(n9405), .ZN(n6558) );
  OR2_X1 U8276 ( .A1(n9688), .A2(n9405), .ZN(n6557) );
  NOR2_X1 U8277 ( .A1(n9671), .A2(n9404), .ZN(n6559) );
  NAND2_X1 U8278 ( .A1(n9671), .A2(n9404), .ZN(n6560) );
  INV_X1 U8279 ( .A(n9233), .ZN(n9403) );
  INV_X1 U8280 ( .A(n9632), .ZN(n6561) );
  OR2_X1 U8281 ( .A1(n9791), .A2(n9402), .ZN(n6562) );
  NAND2_X1 U8282 ( .A1(n6563), .A2(n6562), .ZN(n9616) );
  NOR2_X1 U8283 ( .A1(n9625), .A2(n4749), .ZN(n6564) );
  NAND2_X1 U8284 ( .A1(n9625), .A2(n4749), .ZN(n6565) );
  INV_X1 U8285 ( .A(n9290), .ZN(n9401) );
  AND2_X1 U8286 ( .A1(n9609), .A2(n9401), .ZN(n6566) );
  NAND2_X1 U8287 ( .A1(n9591), .A2(n9400), .ZN(n6567) );
  OR2_X1 U8288 ( .A1(n9770), .A2(n6622), .ZN(n8434) );
  NAND2_X1 U8289 ( .A1(n9770), .A2(n6622), .ZN(n8286) );
  NAND2_X1 U8290 ( .A1(n8434), .A2(n8286), .ZN(n9564) );
  INV_X1 U8291 ( .A(n6622), .ZN(n7235) );
  INV_X1 U8292 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n6635) );
  INV_X1 U8293 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n6569) );
  OAI21_X1 U8294 ( .B1(n6571), .B2(n6635), .A(n6569), .ZN(n6572) );
  NAND2_X1 U8295 ( .A1(P1_REG3_REG_28__SCAN_IN), .A2(P1_REG3_REG_27__SCAN_IN), 
        .ZN(n6570) );
  INV_X1 U8296 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n6575) );
  NAND2_X1 U8297 ( .A1(n6872), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n6574) );
  NAND2_X1 U8298 ( .A1(n5961), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n6573) );
  OAI211_X1 U8299 ( .C1(n4513), .C2(n6575), .A(n6574), .B(n6573), .ZN(n6576)
         );
  OR2_X1 U8300 ( .A1(n9556), .A2(n9538), .ZN(n8433) );
  NAND2_X1 U8301 ( .A1(n9556), .A2(n9538), .ZN(n9533) );
  INV_X1 U8302 ( .A(n9531), .ZN(n6578) );
  NAND2_X1 U8303 ( .A1(n6579), .A2(n9531), .ZN(n6580) );
  OR2_X1 U8304 ( .A1(n8498), .A2(n6581), .ZN(n8513) );
  NAND2_X1 U8305 ( .A1(n6582), .A2(n6581), .ZN(n6583) );
  NAND3_X1 U8306 ( .A1(n7103), .A2(n8513), .A3(n6583), .ZN(n9960) );
  NAND2_X1 U8307 ( .A1(n7759), .A2(n4509), .ZN(n8444) );
  OR2_X1 U8308 ( .A1(n8444), .A2(n8504), .ZN(n10077) );
  AND2_X1 U8309 ( .A1(n9861), .A2(n9401), .ZN(n8431) );
  NAND2_X1 U8310 ( .A1(n9609), .A2(n9290), .ZN(n8430) );
  NAND2_X1 U8311 ( .A1(n8435), .A2(n8430), .ZN(n9601) );
  INV_X1 U8312 ( .A(n9601), .ZN(n6603) );
  NAND2_X1 U8313 ( .A1(n9625), .A2(n9256), .ZN(n8427) );
  NAND2_X1 U8314 ( .A1(n9791), .A2(n9339), .ZN(n9618) );
  NOR2_X1 U8315 ( .A1(n5927), .A2(n9994), .ZN(n6908) );
  OR2_X1 U8316 ( .A1(n5914), .A2(n4998), .ZN(n6584) );
  INV_X1 U8317 ( .A(n8461), .ZN(n7415) );
  NAND2_X1 U8318 ( .A1(n8345), .A2(n7415), .ZN(n6588) );
  NAND2_X1 U8319 ( .A1(n8355), .A2(n7665), .ZN(n8350) );
  INV_X1 U8320 ( .A(n9963), .ZN(n6589) );
  NOR2_X1 U8321 ( .A1(n8350), .A2(n6589), .ZN(n6590) );
  NAND2_X1 U8322 ( .A1(n6590), .A2(n8362), .ZN(n8465) );
  INV_X1 U8323 ( .A(n8465), .ZN(n6591) );
  NAND2_X1 U8324 ( .A1(n7465), .A2(n6591), .ZN(n6597) );
  NAND3_X1 U8325 ( .A1(n4632), .A2(n8354), .A3(n8350), .ZN(n6592) );
  NAND2_X1 U8326 ( .A1(n6592), .A2(n8362), .ZN(n8305) );
  NAND2_X1 U8327 ( .A1(n8354), .A2(n6593), .ZN(n8351) );
  INV_X1 U8328 ( .A(n8346), .ZN(n6594) );
  NOR2_X1 U8329 ( .A1(n8351), .A2(n6594), .ZN(n6595) );
  NAND2_X1 U8330 ( .A1(n4632), .A2(n6595), .ZN(n8466) );
  INV_X1 U8331 ( .A(n8466), .ZN(n6596) );
  OR2_X1 U8332 ( .A1(n8305), .A2(n6596), .ZN(n8308) );
  OR2_X1 U8333 ( .A1(n7765), .A2(n7807), .ZN(n8369) );
  NAND2_X1 U8334 ( .A1(n7765), .A2(n7807), .ZN(n8371) );
  INV_X1 U8335 ( .A(n8368), .ZN(n7737) );
  NOR2_X1 U8336 ( .A1(n7751), .A2(n7737), .ZN(n6598) );
  INV_X1 U8337 ( .A(n8369), .ZN(n6599) );
  NOR2_X1 U8338 ( .A1(n8468), .A2(n6599), .ZN(n6600) );
  NAND2_X1 U8339 ( .A1(n6601), .A2(n8372), .ZN(n7823) );
  OR2_X1 U8340 ( .A1(n10073), .A2(n7927), .ZN(n8381) );
  NAND2_X1 U8341 ( .A1(n10073), .A2(n7927), .ZN(n8380) );
  OR2_X1 U8342 ( .A1(n9396), .A2(n9269), .ZN(n8292) );
  NAND2_X1 U8343 ( .A1(n9396), .A2(n9269), .ZN(n8394) );
  NAND2_X1 U8344 ( .A1(n8292), .A2(n8394), .ZN(n8474) );
  OR2_X1 U8345 ( .A1(n9739), .A2(n9367), .ZN(n8408) );
  NAND2_X1 U8346 ( .A1(n9739), .A2(n9367), .ZN(n8289) );
  OR2_X1 U8347 ( .A1(n9719), .A2(n9281), .ZN(n8409) );
  NAND2_X1 U8348 ( .A1(n9719), .A2(n9281), .ZN(n8410) );
  NAND2_X1 U8349 ( .A1(n9688), .A2(n9232), .ZN(n8405) );
  NAND2_X1 U8350 ( .A1(n8335), .A2(n8405), .ZN(n8478) );
  NAND2_X1 U8351 ( .A1(n9682), .A2(n9681), .ZN(n9680) );
  XNOR2_X1 U8352 ( .A(n9671), .B(n9404), .ZN(n9664) );
  INV_X1 U8353 ( .A(n9664), .ZN(n9662) );
  NAND2_X1 U8354 ( .A1(n9671), .A2(n9337), .ZN(n8422) );
  XNOR2_X1 U8355 ( .A(n9800), .B(n9233), .ZN(n9647) );
  INV_X1 U8356 ( .A(n9647), .ZN(n9655) );
  NAND2_X1 U8357 ( .A1(n9800), .A2(n9233), .ZN(n8281) );
  OR2_X1 U8358 ( .A1(n9791), .A2(n9339), .ZN(n8424) );
  NAND2_X1 U8359 ( .A1(n8424), .A2(n9618), .ZN(n8479) );
  XNOR2_X1 U8360 ( .A(n9591), .B(n9257), .ZN(n9582) );
  INV_X1 U8361 ( .A(n9582), .ZN(n9584) );
  NAND2_X1 U8362 ( .A1(n9591), .A2(n9257), .ZN(n9572) );
  NAND2_X1 U8363 ( .A1(n9571), .A2(n9572), .ZN(n6604) );
  XNOR2_X1 U8364 ( .A(n9532), .B(n9531), .ZN(n6613) );
  AND2_X1 U8365 ( .A1(n8515), .A2(n4509), .ZN(n8455) );
  INV_X1 U8366 ( .A(n8511), .ZN(n6605) );
  OR2_X1 U8367 ( .A1(n6622), .A2(n9537), .ZN(n6611) );
  NAND2_X1 U8368 ( .A1(n6872), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n6607) );
  NAND2_X1 U8369 ( .A1(n5961), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n6606) );
  OAI211_X1 U8370 ( .C1(n4513), .C2(n9766), .A(n6607), .B(n6606), .ZN(n6608)
         );
  INV_X1 U8371 ( .A(n6608), .ZN(n6609) );
  OAI21_X1 U8372 ( .B1(n9548), .B2(n6027), .A(n6609), .ZN(n9399) );
  INV_X1 U8373 ( .A(n9338), .ZN(n9368) );
  NAND2_X1 U8374 ( .A1(n9399), .A2(n9368), .ZN(n6610) );
  AND2_X1 U8375 ( .A1(n6611), .A2(n6610), .ZN(n9222) );
  INV_X1 U8376 ( .A(n9222), .ZN(n6612) );
  NAND2_X1 U8377 ( .A1(n9556), .A2(n9566), .ZN(n6614) );
  NAND2_X1 U8378 ( .A1(n6614), .A2(n9993), .ZN(n6615) );
  OR2_X1 U8379 ( .A1(n9546), .A2(n6615), .ZN(n9559) );
  OAI22_X1 U8380 ( .A1(n9570), .A2(n6619), .B1(n6622), .B2(n9207), .ZN(n6621)
         );
  XNOR2_X1 U8381 ( .A(n6621), .B(n4512), .ZN(n6624) );
  OAI22_X1 U8382 ( .A1(n9570), .A2(n9207), .B1(n6622), .B2(n9214), .ZN(n6623)
         );
  NOR2_X1 U8383 ( .A1(n6624), .A2(n6623), .ZN(n9224) );
  AOI21_X1 U8384 ( .B1(n6624), .B2(n6623), .A(n9224), .ZN(n6629) );
  INV_X1 U8385 ( .A(n6625), .ZN(n6627) );
  OR2_X1 U8386 ( .A1(n6627), .A2(n6626), .ZN(n6630) );
  AOI21_X1 U8387 ( .B1(n6631), .B2(n6630), .A(n6629), .ZN(n6632) );
  OR2_X1 U8388 ( .A1(n9538), .A2(n9338), .ZN(n6634) );
  NAND2_X1 U8389 ( .A1(n9400), .A2(n9199), .ZN(n6633) );
  NAND2_X1 U8390 ( .A1(n6634), .A2(n6633), .ZN(n9576) );
  INV_X1 U8391 ( .A(n9568), .ZN(n6636) );
  OAI22_X1 U8392 ( .A1(n6636), .A2(n9920), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n6635), .ZN(n6637) );
  AOI21_X1 U8393 ( .B1(n9576), .B2(n4510), .A(n6637), .ZN(n6638) );
  INV_X1 U8394 ( .A(n6639), .ZN(n6640) );
  NAND2_X1 U8395 ( .A1(n6641), .A2(n6640), .ZN(P1_U3214) );
  INV_X1 U8396 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n6646) );
  AND4_X2 U8397 ( .A1(n6644), .A2(n6723), .A3(n6643), .A4(n6642), .ZN(n10213)
         );
  INV_X1 U8398 ( .A(n10187), .ZN(n10198) );
  NAND2_X1 U8399 ( .A1(n10213), .A2(n10198), .ZN(n9076) );
  NAND2_X1 U8400 ( .A1(n6649), .A2(n6648), .ZN(P2_U3488) );
  INV_X1 U8401 ( .A(n6650), .ZN(n6651) );
  NAND2_X1 U8402 ( .A1(n8203), .A2(n7086), .ZN(n6654) );
  INV_X1 U8403 ( .A(n6726), .ZN(n6652) );
  INV_X1 U8404 ( .A(n6912), .ZN(n6653) );
  NAND2_X1 U8405 ( .A1(n6654), .A2(n6653), .ZN(n6913) );
  OR2_X1 U8406 ( .A1(n6655), .A2(n6913), .ZN(n6656) );
  NAND2_X1 U8407 ( .A1(n6656), .A2(P2_STATE_REG_SCAN_IN), .ZN(P2_U3150) );
  AND2_X2 U8408 ( .A1(n6912), .A2(P2_STATE_REG_SCAN_IN), .ZN(P2_U3893) );
  INV_X1 U8409 ( .A(n9464), .ZN(n6657) );
  AND2_X1 U8410 ( .A1(n5217), .A2(P1_U3086), .ZN(n7801) );
  INV_X2 U8411 ( .A(n7801), .ZN(n9905) );
  NOR2_X1 U8412 ( .A1(n5217), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9898) );
  INV_X2 U8413 ( .A(n9898), .ZN(n9903) );
  OAI222_X1 U8414 ( .A1(n6657), .A2(P1_U3086), .B1(n9905), .B2(n6681), .C1(
        n9903), .C2(n6006), .ZN(P1_U3350) );
  OAI222_X1 U8415 ( .A1(n9903), .A2(n6658), .B1(n6785), .B2(P1_U3086), .C1(
        n9905), .C2(n6675), .ZN(P1_U3354) );
  INV_X1 U8416 ( .A(n9436), .ZN(n6787) );
  OAI222_X1 U8417 ( .A1(n9903), .A2(n6659), .B1(n6787), .B2(P1_U3086), .C1(
        n9905), .C2(n6677), .ZN(P1_U3353) );
  INV_X1 U8418 ( .A(n7023), .ZN(n6791) );
  OAI222_X1 U8419 ( .A1(n9903), .A2(n6660), .B1(n6791), .B2(P1_U3086), .C1(
        n9905), .C2(n6676), .ZN(P1_U3351) );
  INV_X1 U8420 ( .A(n9451), .ZN(n6789) );
  OAI222_X1 U8421 ( .A1(n9903), .A2(n6661), .B1(n6789), .B2(P1_U3086), .C1(
        n9905), .C2(n6673), .ZN(P1_U3352) );
  INV_X1 U8422 ( .A(n6662), .ZN(n6683) );
  AOI22_X1 U8423 ( .A1(n6810), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_6__SCAN_IN), .B2(n9898), .ZN(n6663) );
  OAI21_X1 U8424 ( .B1(n6683), .B2(n9905), .A(n6663), .ZN(P1_U3349) );
  NAND2_X1 U8425 ( .A1(n6730), .A2(n6664), .ZN(n6665) );
  OAI21_X1 U8426 ( .B1(n6730), .B2(n6666), .A(n6665), .ZN(P2_U3377) );
  NAND2_X1 U8427 ( .A1(n6730), .A2(n6667), .ZN(n6697) );
  INV_X1 U8428 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n6670) );
  INV_X1 U8429 ( .A(n6668), .ZN(n6669) );
  AOI22_X1 U8430 ( .A1(n6697), .A2(n6670), .B1(n6734), .B2(n6669), .ZN(
        P2_U3376) );
  NOR2_X1 U8431 ( .A1(n5217), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9166) );
  OAI222_X1 U8432 ( .A1(n8539), .A2(n6674), .B1(n9171), .B2(n6673), .C1(
        P2_U3151), .C2(n6976), .ZN(P2_U3292) );
  OAI222_X1 U8433 ( .A1(n8539), .A2(n4795), .B1(n9171), .B2(n6675), .C1(
        P2_U3151), .C2(n6991), .ZN(P2_U3294) );
  OAI222_X1 U8434 ( .A1(n7073), .A2(P2_U3151), .B1(n8539), .B2(n5377), .C1(
        n6676), .C2(n9171), .ZN(P2_U3291) );
  OAI222_X1 U8435 ( .A1(n6947), .A2(P2_U3151), .B1(n8539), .B2(n5207), .C1(
        n6677), .C2(n9171), .ZN(P2_U3293) );
  INV_X1 U8436 ( .A(n6678), .ZN(n6685) );
  AOI22_X1 U8437 ( .A1(n6821), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_7__SCAN_IN), .B2(n9898), .ZN(n6679) );
  OAI21_X1 U8438 ( .B1(n6685), .B2(n9905), .A(n6679), .ZN(P1_U3348) );
  OAI222_X1 U8439 ( .A1(n6950), .A2(P2_U3151), .B1(n9171), .B2(n6681), .C1(
        n6680), .C2(n8539), .ZN(P2_U3290) );
  INV_X1 U8440 ( .A(n7147), .ZN(n7171) );
  INV_X1 U8441 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n6682) );
  OAI222_X1 U8442 ( .A1(P2_U3151), .A2(n7171), .B1(n9171), .B2(n6683), .C1(
        n6682), .C2(n8539), .ZN(P2_U3289) );
  INV_X1 U8443 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n6684) );
  OAI222_X1 U8444 ( .A1(P2_U3151), .A2(n7149), .B1(n9171), .B2(n6685), .C1(
        n6684), .C2(n8539), .ZN(P2_U3288) );
  INV_X1 U8445 ( .A(n7332), .ZN(n7200) );
  INV_X1 U8446 ( .A(n6686), .ZN(n6689) );
  INV_X1 U8447 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n6687) );
  OAI222_X1 U8448 ( .A1(n7200), .A2(P2_U3151), .B1(n9171), .B2(n6689), .C1(
        n6687), .C2(n8539), .ZN(P2_U3287) );
  INV_X1 U8449 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n6690) );
  OAI222_X1 U8450 ( .A1(n9903), .A2(n6690), .B1(n9905), .B2(n6689), .C1(
        P1_U3086), .C2(n6688), .ZN(P1_U3347) );
  INV_X1 U8451 ( .A(n6691), .ZN(n6692) );
  INV_X1 U8452 ( .A(n7040), .ZN(n6869) );
  INV_X1 U8453 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n10369) );
  OAI222_X1 U8454 ( .A1(n9905), .A2(n6692), .B1(n6869), .B2(P1_U3086), .C1(
        n10369), .C2(n9903), .ZN(P1_U3346) );
  INV_X1 U8455 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n6693) );
  OAI222_X1 U8456 ( .A1(n8539), .A2(n6693), .B1(P2_U3151), .B2(n7339), .C1(
        n6692), .C2(n9171), .ZN(P2_U3286) );
  INV_X1 U8457 ( .A(n7226), .ZN(n6694) );
  INV_X1 U8458 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n10371) );
  OAI222_X1 U8459 ( .A1(n9905), .A2(n6696), .B1(n6694), .B2(P1_U3086), .C1(
        n10371), .C2(n9903), .ZN(P1_U3345) );
  INV_X1 U8460 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n6695) );
  OAI222_X1 U8461 ( .A1(P2_U3151), .A2(n7577), .B1(n9171), .B2(n6696), .C1(
        n6695), .C2(n8539), .ZN(P2_U3285) );
  INV_X1 U8462 ( .A(P2_D_REG_19__SCAN_IN), .ZN(n6698) );
  NOR2_X1 U8463 ( .A1(n6747), .A2(n6698), .ZN(P2_U3246) );
  INV_X1 U8464 ( .A(P2_D_REG_12__SCAN_IN), .ZN(n6699) );
  NOR2_X1 U8465 ( .A1(n6747), .A2(n6699), .ZN(P2_U3253) );
  INV_X1 U8466 ( .A(P2_D_REG_11__SCAN_IN), .ZN(n6700) );
  NOR2_X1 U8467 ( .A1(n6747), .A2(n6700), .ZN(P2_U3254) );
  INV_X1 U8468 ( .A(P2_D_REG_13__SCAN_IN), .ZN(n6701) );
  NOR2_X1 U8469 ( .A1(n6747), .A2(n6701), .ZN(P2_U3252) );
  INV_X1 U8470 ( .A(P2_D_REG_14__SCAN_IN), .ZN(n6702) );
  NOR2_X1 U8471 ( .A1(n6747), .A2(n6702), .ZN(P2_U3251) );
  INV_X1 U8472 ( .A(P2_D_REG_15__SCAN_IN), .ZN(n6703) );
  NOR2_X1 U8473 ( .A1(n6747), .A2(n6703), .ZN(P2_U3250) );
  INV_X1 U8474 ( .A(P2_D_REG_18__SCAN_IN), .ZN(n6704) );
  NOR2_X1 U8475 ( .A1(n6747), .A2(n6704), .ZN(P2_U3247) );
  INV_X1 U8476 ( .A(P2_D_REG_8__SCAN_IN), .ZN(n6705) );
  NOR2_X1 U8477 ( .A1(n6747), .A2(n6705), .ZN(P2_U3257) );
  INV_X1 U8478 ( .A(P2_D_REG_17__SCAN_IN), .ZN(n6706) );
  NOR2_X1 U8479 ( .A1(n6747), .A2(n6706), .ZN(P2_U3248) );
  INV_X1 U8480 ( .A(P2_D_REG_10__SCAN_IN), .ZN(n6707) );
  NOR2_X1 U8481 ( .A1(n6747), .A2(n6707), .ZN(P2_U3255) );
  INV_X1 U8482 ( .A(P2_D_REG_9__SCAN_IN), .ZN(n6708) );
  NOR2_X1 U8483 ( .A1(n6747), .A2(n6708), .ZN(P2_U3256) );
  INV_X1 U8484 ( .A(P2_D_REG_16__SCAN_IN), .ZN(n6709) );
  NOR2_X1 U8485 ( .A1(n6747), .A2(n6709), .ZN(P2_U3249) );
  INV_X1 U8486 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n10412) );
  NAND2_X1 U8487 ( .A1(n7981), .A2(P2_U3893), .ZN(n6710) );
  OAI21_X1 U8488 ( .B1(P2_U3893), .B2(n10412), .A(n6710), .ZN(P2_U3504) );
  NAND2_X1 U8489 ( .A1(n7458), .A2(P2_U3893), .ZN(n6711) );
  OAI21_X1 U8490 ( .B1(P2_U3893), .B2(n6006), .A(n6711), .ZN(P2_U3496) );
  INV_X1 U8491 ( .A(n6712), .ZN(n6718) );
  AOI22_X1 U8492 ( .A1(n7360), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_11__SCAN_IN), .B2(n9898), .ZN(n6713) );
  OAI21_X1 U8493 ( .B1(n6718), .B2(n9905), .A(n6713), .ZN(P1_U3344) );
  INV_X1 U8494 ( .A(n9893), .ZN(n6895) );
  INV_X1 U8495 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n10420) );
  INV_X1 U8496 ( .A(n10001), .ZN(n10002) );
  OAI21_X1 U8497 ( .B1(n10002), .B2(P1_D_REG_1__SCAN_IN), .A(n6715), .ZN(n6716) );
  OAI21_X1 U8498 ( .B1(n6895), .B2(n10420), .A(n6716), .ZN(P1_U3440) );
  INV_X1 U8499 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n6717) );
  OAI222_X1 U8500 ( .A1(n7581), .A2(P2_U3151), .B1(n9171), .B2(n6718), .C1(
        n6717), .C2(n8539), .ZN(P2_U3284) );
  INV_X1 U8501 ( .A(n7699), .ZN(n8759) );
  INV_X1 U8502 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n6719) );
  OAI222_X1 U8503 ( .A1(P2_U3151), .A2(n8759), .B1(n9171), .B2(n6720), .C1(
        n6719), .C2(n8539), .ZN(P2_U3283) );
  INV_X1 U8504 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n10410) );
  INV_X1 U8505 ( .A(n7358), .ZN(n7488) );
  OAI222_X1 U8506 ( .A1(n9903), .A2(n10410), .B1(n7488), .B2(P1_U3086), .C1(
        n9905), .C2(n6720), .ZN(P1_U3343) );
  INV_X1 U8507 ( .A(n6721), .ZN(n6724) );
  OAI21_X1 U8508 ( .B1(n6724), .B2(n6723), .A(n6722), .ZN(n6728) );
  OR2_X1 U8509 ( .A1(n6731), .A2(n6737), .ZN(n6727) );
  NAND4_X1 U8510 ( .A1(n6728), .A2(n6727), .A3(n6726), .A4(n6725), .ZN(n6729)
         );
  NAND2_X1 U8511 ( .A1(n6729), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6733) );
  INV_X1 U8512 ( .A(n6899), .ZN(n6743) );
  NAND2_X1 U8513 ( .A1(n6730), .A2(n6743), .ZN(n8267) );
  OR2_X1 U8514 ( .A1(n8267), .A2(n6731), .ZN(n6732) );
  AND2_X1 U8515 ( .A1(n6733), .A2(n6732), .ZN(n7087) );
  AND2_X1 U8516 ( .A1(n7087), .A2(n6734), .ZN(n6884) );
  INV_X1 U8517 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n6904) );
  NAND2_X1 U8518 ( .A1(n5317), .A2(n5071), .ZN(n8062) );
  AND2_X1 U8519 ( .A1(n8058), .A2(n8062), .ZN(n8221) );
  INV_X1 U8520 ( .A(n8221), .ZN(n6900) );
  INV_X1 U8521 ( .A(n6735), .ZN(n6736) );
  NAND2_X1 U8522 ( .A1(n6741), .A2(n6736), .ZN(n6740) );
  INV_X1 U8523 ( .A(n6737), .ZN(n6738) );
  NAND2_X1 U8524 ( .A1(n6844), .A2(n6738), .ZN(n6739) );
  NAND2_X1 U8525 ( .A1(n6741), .A2(n10198), .ZN(n6742) );
  NAND2_X1 U8526 ( .A1(n6742), .A2(n10141), .ZN(n8655) );
  INV_X1 U8527 ( .A(n8655), .ZN(n8728) );
  AND2_X1 U8528 ( .A1(n6842), .A2(n6743), .ZN(n6744) );
  NAND2_X1 U8529 ( .A1(n6844), .A2(n6744), .ZN(n8707) );
  OAI22_X1 U8530 ( .A1(n8728), .A2(n5071), .B1(n6841), .B2(n8707), .ZN(n6745)
         );
  AOI21_X1 U8531 ( .B1(n6900), .B2(n8717), .A(n6745), .ZN(n6746) );
  OAI21_X1 U8532 ( .B1(n6884), .B2(n6904), .A(n6746), .ZN(P2_U3172) );
  INV_X1 U8533 ( .A(P2_D_REG_4__SCAN_IN), .ZN(n6748) );
  NOR2_X1 U8534 ( .A1(n6747), .A2(n6748), .ZN(P2_U3261) );
  INV_X1 U8535 ( .A(P2_D_REG_6__SCAN_IN), .ZN(n6749) );
  NOR2_X1 U8536 ( .A1(n6747), .A2(n6749), .ZN(P2_U3259) );
  INV_X1 U8537 ( .A(P2_D_REG_27__SCAN_IN), .ZN(n6750) );
  NOR2_X1 U8538 ( .A1(n6747), .A2(n6750), .ZN(P2_U3238) );
  INV_X1 U8539 ( .A(P2_D_REG_5__SCAN_IN), .ZN(n6751) );
  NOR2_X1 U8540 ( .A1(n6747), .A2(n6751), .ZN(P2_U3260) );
  INV_X1 U8541 ( .A(P2_D_REG_7__SCAN_IN), .ZN(n6752) );
  NOR2_X1 U8542 ( .A1(n6747), .A2(n6752), .ZN(P2_U3258) );
  INV_X1 U8543 ( .A(P2_D_REG_20__SCAN_IN), .ZN(n6753) );
  NOR2_X1 U8544 ( .A1(n6747), .A2(n6753), .ZN(P2_U3245) );
  INV_X1 U8545 ( .A(P2_D_REG_31__SCAN_IN), .ZN(n6754) );
  NOR2_X1 U8546 ( .A1(n6747), .A2(n6754), .ZN(P2_U3234) );
  INV_X1 U8547 ( .A(P2_D_REG_22__SCAN_IN), .ZN(n6755) );
  NOR2_X1 U8548 ( .A1(n6747), .A2(n6755), .ZN(P2_U3243) );
  INV_X1 U8549 ( .A(P2_D_REG_24__SCAN_IN), .ZN(n6756) );
  NOR2_X1 U8550 ( .A1(n6747), .A2(n6756), .ZN(P2_U3241) );
  INV_X1 U8551 ( .A(P2_D_REG_21__SCAN_IN), .ZN(n6757) );
  NOR2_X1 U8552 ( .A1(n6747), .A2(n6757), .ZN(P2_U3244) );
  INV_X1 U8553 ( .A(P2_D_REG_2__SCAN_IN), .ZN(n6758) );
  NOR2_X1 U8554 ( .A1(n6747), .A2(n6758), .ZN(P2_U3263) );
  INV_X1 U8555 ( .A(P2_D_REG_3__SCAN_IN), .ZN(n6759) );
  NOR2_X1 U8556 ( .A1(n6747), .A2(n6759), .ZN(P2_U3262) );
  INV_X1 U8557 ( .A(P2_D_REG_28__SCAN_IN), .ZN(n6760) );
  NOR2_X1 U8558 ( .A1(n6747), .A2(n6760), .ZN(P2_U3237) );
  INV_X1 U8559 ( .A(P2_D_REG_25__SCAN_IN), .ZN(n6761) );
  NOR2_X1 U8560 ( .A1(n6747), .A2(n6761), .ZN(P2_U3240) );
  INV_X1 U8561 ( .A(P2_D_REG_29__SCAN_IN), .ZN(n6762) );
  NOR2_X1 U8562 ( .A1(n6747), .A2(n6762), .ZN(P2_U3236) );
  INV_X1 U8563 ( .A(P2_D_REG_30__SCAN_IN), .ZN(n6763) );
  NOR2_X1 U8564 ( .A1(n6747), .A2(n6763), .ZN(P2_U3235) );
  INV_X1 U8565 ( .A(P2_D_REG_26__SCAN_IN), .ZN(n6764) );
  NOR2_X1 U8566 ( .A1(n6747), .A2(n6764), .ZN(P2_U3239) );
  INV_X1 U8567 ( .A(P2_D_REG_23__SCAN_IN), .ZN(n6765) );
  NOR2_X1 U8568 ( .A1(n6747), .A2(n6765), .ZN(P2_U3242) );
  NAND2_X1 U8569 ( .A1(n6766), .A2(n6769), .ZN(n6767) );
  NAND2_X1 U8570 ( .A1(n6768), .A2(n6767), .ZN(n6780) );
  INV_X1 U8571 ( .A(n6780), .ZN(n6770) );
  INV_X1 U8572 ( .A(n6769), .ZN(n7803) );
  OAI21_X1 U8573 ( .B1(n5925), .B2(n7803), .A(P1_STATE_REG_SCAN_IN), .ZN(n6781) );
  INV_X1 U8574 ( .A(n9507), .ZN(n9956) );
  NOR2_X1 U8575 ( .A1(n9956), .A2(n4511), .ZN(P1_U3085) );
  INV_X1 U8576 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n9986) );
  MUX2_X1 U8577 ( .A(n9986), .B(P1_REG2_REG_1__SCAN_IN), .S(n6785), .Z(n9428)
         );
  AND2_X1 U8578 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(
        n9427) );
  NAND2_X1 U8579 ( .A1(n9428), .A2(n9427), .ZN(n9426) );
  INV_X1 U8580 ( .A(n6785), .ZN(n9425) );
  NAND2_X1 U8581 ( .A1(n9425), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n6771) );
  NAND2_X1 U8582 ( .A1(n9426), .A2(n6771), .ZN(n9442) );
  NAND2_X1 U8583 ( .A1(n9436), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n6772) );
  NAND2_X1 U8584 ( .A1(n9441), .A2(n6772), .ZN(n9456) );
  XNOR2_X1 U8585 ( .A(n9451), .B(n6773), .ZN(n9457) );
  NAND2_X1 U8586 ( .A1(n9456), .A2(n9457), .ZN(n9455) );
  NAND2_X1 U8587 ( .A1(n9451), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n6774) );
  NAND2_X1 U8588 ( .A1(n9455), .A2(n6774), .ZN(n7025) );
  MUX2_X1 U8589 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n7395), .S(n7023), .Z(n7026)
         );
  NAND2_X1 U8590 ( .A1(n7025), .A2(n7026), .ZN(n7024) );
  NAND2_X1 U8591 ( .A1(n7023), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n6775) );
  NAND2_X1 U8592 ( .A1(n7024), .A2(n6775), .ZN(n9467) );
  OR2_X1 U8593 ( .A1(n9464), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n6777) );
  NAND2_X1 U8594 ( .A1(P1_REG2_REG_5__SCAN_IN), .A2(n9464), .ZN(n6776) );
  AND2_X1 U8595 ( .A1(n6777), .A2(n6776), .ZN(n9468) );
  AND2_X1 U8596 ( .A1(n9467), .A2(n9468), .ZN(n9465) );
  NAND2_X1 U8597 ( .A1(P1_REG2_REG_6__SCAN_IN), .A2(n6810), .ZN(n6778) );
  OAI21_X1 U8598 ( .B1(P1_REG2_REG_6__SCAN_IN), .B2(n6810), .A(n6778), .ZN(
        n6805) );
  NOR2_X1 U8599 ( .A1(n6806), .A2(n6805), .ZN(n6804) );
  AOI21_X1 U8600 ( .B1(n6810), .B2(P1_REG2_REG_6__SCAN_IN), .A(n6804), .ZN(
        n6784) );
  NAND2_X1 U8601 ( .A1(n6821), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n6779) );
  OAI21_X1 U8602 ( .B1(n6821), .B2(P1_REG2_REG_7__SCAN_IN), .A(n6779), .ZN(
        n6783) );
  NOR2_X1 U8603 ( .A1(n6784), .A2(n6783), .ZN(n6817) );
  OR2_X1 U8604 ( .A1(n6781), .A2(n6780), .ZN(n9958) );
  INV_X1 U8605 ( .A(n4508), .ZN(n6782) );
  NAND2_X1 U8606 ( .A1(n7016), .A2(n6782), .ZN(n8514) );
  NOR2_X2 U8607 ( .A1(n9958), .A2(n8514), .ZN(n9517) );
  AOI211_X1 U8608 ( .C1(n6784), .C2(n6783), .A(n6817), .B(n7891), .ZN(n6803)
         );
  INV_X1 U8609 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n6790) );
  INV_X1 U8610 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n6788) );
  MUX2_X1 U8611 ( .A(P1_REG1_REG_2__SCAN_IN), .B(n6788), .S(n9436), .Z(n9439)
         );
  INV_X1 U8612 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n10085) );
  AND2_X1 U8613 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(
        n9423) );
  NAND2_X1 U8614 ( .A1(n9424), .A2(n9423), .ZN(n9422) );
  NAND2_X1 U8615 ( .A1(n9425), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n6786) );
  NAND2_X1 U8616 ( .A1(n9422), .A2(n6786), .ZN(n9438) );
  NAND2_X1 U8617 ( .A1(n9439), .A2(n9438), .ZN(n9437) );
  OAI21_X1 U8618 ( .B1(n6788), .B2(n6787), .A(n9437), .ZN(n9453) );
  XOR2_X1 U8619 ( .A(P1_REG1_REG_3__SCAN_IN), .B(n9451), .Z(n9454) );
  NAND2_X1 U8620 ( .A1(n9453), .A2(n9454), .ZN(n9452) );
  OAI21_X1 U8621 ( .B1(n6790), .B2(n6789), .A(n9452), .ZN(n7021) );
  MUX2_X1 U8622 ( .A(P1_REG1_REG_4__SCAN_IN), .B(n6792), .S(n7023), .Z(n7022)
         );
  NAND2_X1 U8623 ( .A1(n7021), .A2(n7022), .ZN(n7020) );
  OAI21_X1 U8624 ( .B1(n6792), .B2(n6791), .A(n7020), .ZN(n9470) );
  NAND2_X1 U8625 ( .A1(P1_REG1_REG_5__SCAN_IN), .A2(n9464), .ZN(n6793) );
  OAI21_X1 U8626 ( .B1(n9464), .B2(P1_REG1_REG_5__SCAN_IN), .A(n6793), .ZN(
        n6794) );
  INV_X1 U8627 ( .A(n6794), .ZN(n9471) );
  NAND2_X1 U8628 ( .A1(n9470), .A2(n9471), .ZN(n9469) );
  NAND2_X1 U8629 ( .A1(P1_REG1_REG_6__SCAN_IN), .A2(n6810), .ZN(n6795) );
  OAI21_X1 U8630 ( .B1(n6810), .B2(P1_REG1_REG_6__SCAN_IN), .A(n6795), .ZN(
        n6808) );
  NAND2_X1 U8631 ( .A1(n6821), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n6796) );
  OAI21_X1 U8632 ( .B1(n6821), .B2(P1_REG1_REG_7__SCAN_IN), .A(n6796), .ZN(
        n6798) );
  NOR2_X1 U8633 ( .A1(n4547), .A2(n6798), .ZN(n6820) );
  INV_X1 U8634 ( .A(n9958), .ZN(n6797) );
  NAND2_X1 U8635 ( .A1(n6797), .A2(n4508), .ZN(n9510) );
  AOI211_X1 U8636 ( .C1(n4547), .C2(n6798), .A(n6820), .B(n9510), .ZN(n6802)
         );
  INV_X1 U8637 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n6800) );
  NOR2_X2 U8638 ( .A1(n9958), .A2(n7016), .ZN(n9516) );
  NAND2_X1 U8639 ( .A1(n9516), .A2(n6821), .ZN(n6799) );
  NAND2_X1 U8640 ( .A1(P1_REG3_REG_7__SCAN_IN), .A2(P1_U3086), .ZN(n7562) );
  OAI211_X1 U8641 ( .C1(n6800), .C2(n9507), .A(n6799), .B(n7562), .ZN(n6801)
         );
  OR3_X1 U8642 ( .A1(n6803), .A2(n6802), .A3(n6801), .ZN(P1_U3250) );
  AOI211_X1 U8643 ( .C1(n6806), .C2(n6805), .A(n6804), .B(n7891), .ZN(n6816)
         );
  AOI211_X1 U8644 ( .C1(n6809), .C2(n6808), .A(n6807), .B(n9510), .ZN(n6815)
         );
  INV_X1 U8645 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n6813) );
  NAND2_X1 U8646 ( .A1(n9516), .A2(n6810), .ZN(n6812) );
  NAND2_X1 U8647 ( .A1(P1_REG3_REG_6__SCAN_IN), .A2(P1_U3086), .ZN(n6811) );
  OAI211_X1 U8648 ( .C1(n6813), .C2(n9507), .A(n6812), .B(n6811), .ZN(n6814)
         );
  OR3_X1 U8649 ( .A1(n6816), .A2(n6815), .A3(n6814), .ZN(P1_U3249) );
  AOI21_X1 U8650 ( .B1(P1_REG2_REG_7__SCAN_IN), .B2(n6821), .A(n6817), .ZN(
        n6819) );
  XNOR2_X1 U8651 ( .A(n6860), .B(P1_REG2_REG_8__SCAN_IN), .ZN(n6818) );
  NOR2_X1 U8652 ( .A1(n6818), .A2(n6819), .ZN(n6859) );
  AOI211_X1 U8653 ( .C1(n6819), .C2(n6818), .A(n6859), .B(n7891), .ZN(n6828)
         );
  AOI21_X1 U8654 ( .B1(n6821), .B2(P1_REG1_REG_7__SCAN_IN), .A(n6820), .ZN(
        n6823) );
  XNOR2_X1 U8655 ( .A(n6860), .B(P1_REG1_REG_8__SCAN_IN), .ZN(n6822) );
  NOR2_X1 U8656 ( .A1(n6822), .A2(n6823), .ZN(n6855) );
  AOI211_X1 U8657 ( .C1(n6823), .C2(n6822), .A(n6855), .B(n9510), .ZN(n6827)
         );
  INV_X1 U8658 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n6825) );
  NAND2_X1 U8659 ( .A1(n9516), .A2(n6860), .ZN(n6824) );
  NAND2_X1 U8660 ( .A1(P1_U3086), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n9942) );
  OAI211_X1 U8661 ( .C1(n6825), .C2(n9507), .A(n6824), .B(n9942), .ZN(n6826)
         );
  OR3_X1 U8662 ( .A1(n6828), .A2(n6827), .A3(n6826), .ZN(P1_U3251) );
  INV_X1 U8663 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n6832) );
  INV_X1 U8664 ( .A(n6829), .ZN(n10182) );
  OAI21_X1 U8665 ( .B1(n10151), .B2(n10192), .A(n6900), .ZN(n6830) );
  OR2_X1 U8666 ( .A1(n6841), .A2(n9008), .ZN(n6901) );
  OAI211_X1 U8667 ( .C1(n10187), .C2(n5071), .A(n6830), .B(n6901), .ZN(n6853)
         );
  NAND2_X1 U8668 ( .A1(n6853), .A2(n10199), .ZN(n6831) );
  OAI21_X1 U8669 ( .B1(n6832), .B2(n10199), .A(n6831), .ZN(P2_U3390) );
  NAND2_X1 U8670 ( .A1(n6834), .A2(n8206), .ZN(n6836) );
  AND2_X1 U8671 ( .A1(n6836), .A2(n6835), .ZN(n6837) );
  INV_X1 U8672 ( .A(n7074), .ZN(n6838) );
  OR2_X1 U8673 ( .A1(n6839), .A2(n6838), .ZN(n6840) );
  NAND2_X1 U8674 ( .A1(n8058), .A2(n6840), .ZN(n6879) );
  XOR2_X1 U8675 ( .A(n6878), .B(n6879), .Z(n6848) );
  INV_X1 U8676 ( .A(n8707), .ZN(n8725) );
  NOR2_X1 U8677 ( .A1(n6842), .A2(n6899), .ZN(n6843) );
  NAND2_X1 U8678 ( .A1(n6844), .A2(n6843), .ZN(n8677) );
  OAI22_X1 U8679 ( .A1(n7011), .A2(n8728), .B1(n5070), .B2(n8677), .ZN(n6846)
         );
  NOR2_X1 U8680 ( .A1(n6884), .A2(n6992), .ZN(n6845) );
  AOI211_X1 U8681 ( .C1(n8725), .C2(n8743), .A(n6846), .B(n6845), .ZN(n6847)
         );
  OAI21_X1 U8682 ( .B1(n8658), .B2(n6848), .A(n6847), .ZN(P2_U3162) );
  INV_X1 U8683 ( .A(n6849), .ZN(n6852) );
  INV_X1 U8684 ( .A(n7607), .ZN(n6850) );
  OAI222_X1 U8685 ( .A1(n9905), .A2(n6852), .B1(n9903), .B2(n10412), .C1(
        P1_U3086), .C2(n6850), .ZN(P1_U3342) );
  INV_X1 U8686 ( .A(n8760), .ZN(n10117) );
  INV_X1 U8687 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n6851) );
  OAI222_X1 U8688 ( .A1(P2_U3151), .A2(n10117), .B1(n9171), .B2(n6852), .C1(
        n6851), .C2(n8539), .ZN(P2_U3282) );
  NAND2_X1 U8689 ( .A1(n6853), .A2(n10213), .ZN(n6854) );
  OAI21_X1 U8690 ( .B1(n10213), .B2(n6914), .A(n6854), .ZN(P2_U3459) );
  INV_X1 U8691 ( .A(n9516), .ZN(n7885) );
  NOR2_X1 U8692 ( .A1(P1_REG1_REG_9__SCAN_IN), .A2(n7040), .ZN(n6856) );
  AOI21_X1 U8693 ( .B1(n7040), .B2(P1_REG1_REG_9__SCAN_IN), .A(n6856), .ZN(
        n6857) );
  OAI21_X1 U8694 ( .B1(n6858), .B2(n6857), .A(n7039), .ZN(n6865) );
  NOR2_X1 U8695 ( .A1(P1_REG2_REG_9__SCAN_IN), .A2(n7040), .ZN(n6861) );
  AOI21_X1 U8696 ( .B1(n7040), .B2(P1_REG2_REG_9__SCAN_IN), .A(n6861), .ZN(
        n6862) );
  NAND2_X1 U8697 ( .A1(n6862), .A2(n6863), .ZN(n7035) );
  OAI21_X1 U8698 ( .B1(n6863), .B2(n6862), .A(n7035), .ZN(n6864) );
  AOI22_X1 U8699 ( .A1(n9499), .A2(n6865), .B1(n9517), .B2(n6864), .ZN(n6868)
         );
  NOR2_X1 U8700 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6866), .ZN(n9304) );
  AOI21_X1 U8701 ( .B1(n9956), .B2(P1_ADDR_REG_9__SCAN_IN), .A(n9304), .ZN(
        n6867) );
  OAI211_X1 U8702 ( .C1(n6869), .C2(n7885), .A(n6868), .B(n6867), .ZN(P1_U3252) );
  NAND2_X1 U8703 ( .A1(n8493), .A2(n4511), .ZN(n6870) );
  OAI21_X1 U8704 ( .B1(n4511), .B2(n9163), .A(n6870), .ZN(P1_U3585) );
  NAND2_X1 U8705 ( .A1(n7416), .A2(n4511), .ZN(n6871) );
  OAI21_X1 U8706 ( .B1(n4511), .B2(n5377), .A(n6871), .ZN(P1_U3558) );
  INV_X1 U8707 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n6875) );
  NAND2_X1 U8708 ( .A1(n5961), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n6874) );
  NAND2_X1 U8709 ( .A1(n6872), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n6873) );
  OAI211_X1 U8710 ( .C1(n4513), .C2(n6875), .A(n6874), .B(n6873), .ZN(n8445)
         );
  NAND2_X1 U8711 ( .A1(n8445), .A2(n4511), .ZN(n6876) );
  OAI21_X1 U8712 ( .B1(n8185), .B2(n4511), .A(n6876), .ZN(P1_U3584) );
  NAND2_X1 U8713 ( .A1(n7096), .A2(n4511), .ZN(n6877) );
  OAI21_X1 U8714 ( .B1(n4511), .B2(n5207), .A(n6877), .ZN(P1_U3556) );
  XNOR2_X1 U8715 ( .A(n7077), .B(n8743), .ZN(n7075) );
  NAND2_X1 U8716 ( .A1(n6879), .A2(n6878), .ZN(n6883) );
  INV_X1 U8717 ( .A(n6880), .ZN(n6881) );
  NAND2_X1 U8718 ( .A1(n6841), .A2(n6881), .ZN(n6882) );
  NAND2_X1 U8719 ( .A1(n6883), .A2(n6882), .ZN(n7076) );
  XOR2_X1 U8720 ( .A(n7075), .B(n7076), .Z(n6888) );
  OAI22_X1 U8721 ( .A1(n8728), .A2(n10143), .B1(n6841), .B2(n8677), .ZN(n6886)
         );
  INV_X1 U8722 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n10583) );
  NOR2_X1 U8723 ( .A1(n6884), .A2(n10583), .ZN(n6885) );
  AOI211_X1 U8724 ( .C1(n8725), .C2(n10149), .A(n6886), .B(n6885), .ZN(n6887)
         );
  OAI21_X1 U8725 ( .B1(n6888), .B2(n8658), .A(n6887), .ZN(P2_U3177) );
  INV_X1 U8726 ( .A(n6889), .ZN(n6892) );
  INV_X1 U8727 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n6890) );
  OAI222_X1 U8728 ( .A1(n10135), .A2(P2_U3151), .B1(n9171), .B2(n6892), .C1(
        n6890), .C2(n8539), .ZN(P2_U3281) );
  INV_X1 U8729 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n10293) );
  INV_X1 U8730 ( .A(n7887), .ZN(n6891) );
  OAI222_X1 U8731 ( .A1(n9903), .A2(n10293), .B1(n9905), .B2(n6892), .C1(
        P1_U3086), .C2(n6891), .ZN(P1_U3341) );
  XNOR2_X1 U8732 ( .A(n6894), .B(n6893), .ZN(n7014) );
  AND2_X1 U8733 ( .A1(n5914), .A2(n9368), .ZN(n6909) );
  NAND2_X1 U8734 ( .A1(n6896), .A2(n6895), .ZN(n7189) );
  AOI22_X1 U8735 ( .A1(n4510), .A2(n6909), .B1(n7189), .B2(
        P1_REG3_REG_0__SCAN_IN), .ZN(n6898) );
  NAND2_X1 U8736 ( .A1(n9395), .A2(n7110), .ZN(n6897) );
  OAI211_X1 U8737 ( .C1(n7014), .C2(n9916), .A(n6898), .B(n6897), .ZN(P1_U3232) );
  NAND3_X1 U8738 ( .A1(n6900), .A2(n6899), .A3(n10187), .ZN(n6902) );
  AOI21_X1 U8739 ( .B1(n6902), .B2(n6901), .A(n10159), .ZN(n6907) );
  INV_X1 U8740 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n6903) );
  NOR2_X1 U8741 ( .A1(n9029), .A2(n6903), .ZN(n6906) );
  OAI22_X1 U8742 ( .A1(n9014), .A2(n5071), .B1(n6904), .B2(n10141), .ZN(n6905)
         );
  OR3_X1 U8743 ( .A1(n6907), .A2(n6906), .A3(n6905), .ZN(P2_U3233) );
  INV_X1 U8744 ( .A(n6908), .ZN(n9981) );
  NAND2_X1 U8745 ( .A1(n5927), .A2(n9994), .ZN(n8296) );
  NAND2_X1 U8746 ( .A1(n9981), .A2(n8296), .ZN(n8457) );
  OAI21_X1 U8747 ( .B1(n9837), .B2(n10070), .A(n8457), .ZN(n6910) );
  INV_X1 U8748 ( .A(n6909), .ZN(n7104) );
  OAI211_X1 U8749 ( .C1(n7103), .C2(n9994), .A(n6910), .B(n7104), .ZN(n9847)
         );
  NAND2_X1 U8750 ( .A1(n9847), .A2(n10084), .ZN(n6911) );
  OAI21_X1 U8751 ( .B1(n10084), .B2(n5916), .A(n6911), .ZN(P1_U3453) );
  OR2_X1 U8752 ( .A1(P2_U3150), .A2(n6912), .ZN(n8870) );
  INV_X1 U8753 ( .A(P2_ADDR_REG_0__SCAN_IN), .ZN(n6924) );
  NOR2_X1 U8754 ( .A1(n6919), .A2(n8276), .ZN(n6952) );
  INV_X1 U8755 ( .A(n6952), .ZN(n6932) );
  NAND2_X1 U8756 ( .A1(P2_U3893), .A2(n8276), .ZN(n10129) );
  MUX2_X1 U8757 ( .A(n6903), .B(n6914), .S(n8860), .Z(n6915) );
  MUX2_X1 U8758 ( .A(P2_REG2_REG_0__SCAN_IN), .B(P2_REG1_REG_0__SCAN_IN), .S(
        n8860), .Z(n6916) );
  NAND2_X1 U8759 ( .A1(n6916), .A2(n6943), .ZN(n6917) );
  AOI22_X1 U8760 ( .A1(n6932), .A2(n10129), .B1(n6989), .B2(n6917), .ZN(n6918)
         );
  AOI21_X1 U8761 ( .B1(P2_REG3_REG_0__SCAN_IN), .B2(P2_U3151), .A(n6918), .ZN(
        n6923) );
  NOR2_X1 U8762 ( .A1(n6919), .A2(n8860), .ZN(n6921) );
  MUX2_X1 U8763 ( .A(n6921), .B(P2_U3893), .S(n6920), .Z(n8872) );
  OAI211_X1 U8764 ( .C1(n8870), .C2(n6924), .A(n6923), .B(n6922), .ZN(P2_U3182) );
  MUX2_X1 U8765 ( .A(P2_REG2_REG_4__SCAN_IN), .B(P2_REG1_REG_4__SCAN_IN), .S(
        n8860), .Z(n6931) );
  MUX2_X1 U8766 ( .A(n7239), .B(n6925), .S(n8860), .Z(n6926) );
  XNOR2_X1 U8767 ( .A(n6926), .B(n6991), .ZN(n6990) );
  INV_X1 U8768 ( .A(n6926), .ZN(n6927) );
  AOI22_X1 U8769 ( .A1(n6990), .A2(n6989), .B1(n6927), .B2(n6991), .ZN(n6959)
         );
  MUX2_X1 U8770 ( .A(P2_REG2_REG_2__SCAN_IN), .B(P2_REG1_REG_2__SCAN_IN), .S(
        n8860), .Z(n6928) );
  XNOR2_X1 U8771 ( .A(n6928), .B(n6947), .ZN(n6958) );
  INV_X1 U8772 ( .A(n6947), .ZN(n6971) );
  INV_X1 U8773 ( .A(n6928), .ZN(n6929) );
  OAI22_X1 U8774 ( .A1(n6959), .A2(n6958), .B1(n6971), .B2(n6929), .ZN(n6974)
         );
  MUX2_X1 U8775 ( .A(P2_REG2_REG_3__SCAN_IN), .B(P2_REG1_REG_3__SCAN_IN), .S(
        n8860), .Z(n6930) );
  XNOR2_X1 U8776 ( .A(n6930), .B(n6976), .ZN(n6975) );
  NOR2_X1 U8777 ( .A1(n6974), .A2(n6975), .ZN(n7052) );
  NOR2_X1 U8778 ( .A1(n6930), .A2(n6976), .ZN(n7051) );
  XNOR2_X1 U8779 ( .A(n6931), .B(n7073), .ZN(n7050) );
  NOR3_X1 U8780 ( .A1(n7052), .A2(n7051), .A3(n7050), .ZN(n7049) );
  AOI21_X1 U8781 ( .B1(n6931), .B2(n7073), .A(n7049), .ZN(n7133) );
  MUX2_X1 U8782 ( .A(P2_REG2_REG_5__SCAN_IN), .B(P2_REG1_REG_5__SCAN_IN), .S(
        n8860), .Z(n7130) );
  XNOR2_X1 U8783 ( .A(n7130), .B(n6950), .ZN(n7132) );
  XNOR2_X1 U8784 ( .A(n7133), .B(n7132), .ZN(n6957) );
  INV_X1 U8785 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n6941) );
  INV_X1 U8786 ( .A(n10127), .ZN(n8847) );
  INV_X1 U8787 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n10202) );
  MUX2_X1 U8788 ( .A(P2_REG1_REG_2__SCAN_IN), .B(n10202), .S(n6947), .Z(n6962)
         );
  AND2_X1 U8789 ( .A1(n6943), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n6933) );
  NAND2_X1 U8790 ( .A1(n6944), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n6934) );
  OAI21_X1 U8791 ( .B1(n6991), .B2(n6933), .A(n6934), .ZN(n6997) );
  OR2_X1 U8792 ( .A1(n6997), .A2(n6925), .ZN(n6995) );
  NAND2_X1 U8793 ( .A1(n6995), .A2(n6934), .ZN(n6961) );
  NAND2_X1 U8794 ( .A1(n6947), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n6935) );
  OAI21_X1 U8795 ( .B1(n6936), .B2(n6976), .A(n7062), .ZN(n6981) );
  NAND2_X1 U8796 ( .A1(n7064), .A2(n7062), .ZN(n6937) );
  INV_X1 U8797 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n10205) );
  MUX2_X1 U8798 ( .A(P2_REG1_REG_4__SCAN_IN), .B(n10205), .S(n7073), .Z(n7061)
         );
  OAI21_X1 U8799 ( .B1(n4594), .B2(P2_REG1_REG_5__SCAN_IN), .A(n7174), .ZN(
        n6938) );
  NAND2_X1 U8800 ( .A1(n8847), .A2(n6938), .ZN(n6940) );
  NOR2_X1 U8801 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n5151), .ZN(n7247) );
  INV_X1 U8802 ( .A(n7247), .ZN(n6939) );
  OAI211_X1 U8803 ( .C1(n6941), .C2(n8870), .A(n6940), .B(n6939), .ZN(n6955)
         );
  INV_X1 U8804 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n6942) );
  MUX2_X1 U8805 ( .A(P2_REG2_REG_2__SCAN_IN), .B(n6942), .S(n6947), .Z(n6965)
         );
  AND2_X1 U8806 ( .A1(n6943), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n6945) );
  NAND2_X1 U8807 ( .A1(n6944), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n6946) );
  NAND2_X1 U8808 ( .A1(n6993), .A2(n6946), .ZN(n6964) );
  INV_X1 U8809 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n7284) );
  NAND2_X1 U8810 ( .A1(n7058), .A2(n7056), .ZN(n6948) );
  INV_X1 U8811 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n7275) );
  MUX2_X1 U8812 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n7275), .S(n7073), .Z(n7055)
         );
  NAND2_X1 U8813 ( .A1(n6948), .A2(n7055), .ZN(n7060) );
  NAND2_X1 U8814 ( .A1(n7073), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n6949) );
  NAND2_X1 U8815 ( .A1(n6951), .A2(n5383), .ZN(n6953) );
  AND2_X1 U8816 ( .A1(n6952), .A2(n8266), .ZN(n8878) );
  AOI21_X1 U8817 ( .B1(n7166), .B2(n6953), .A(n10131), .ZN(n6954) );
  AOI211_X1 U8818 ( .C1(n8872), .C2(n4950), .A(n6955), .B(n6954), .ZN(n6956)
         );
  OAI21_X1 U8819 ( .B1(n6957), .B2(n10129), .A(n6956), .ZN(P2_U3187) );
  XNOR2_X1 U8820 ( .A(n6959), .B(n6958), .ZN(n6973) );
  OAI21_X1 U8821 ( .B1(n6962), .B2(n6961), .A(n6960), .ZN(n6967) );
  OAI21_X1 U8822 ( .B1(n6965), .B2(n6964), .A(n6963), .ZN(n6966) );
  AOI22_X1 U8823 ( .A1(n8847), .A2(n6967), .B1(n8878), .B2(n6966), .ZN(n6969)
         );
  NAND2_X1 U8824 ( .A1(n10118), .A2(P2_ADDR_REG_2__SCAN_IN), .ZN(n6968) );
  OAI211_X1 U8825 ( .C1(P2_STATE_REG_SCAN_IN), .C2(n10583), .A(n6969), .B(
        n6968), .ZN(n6970) );
  AOI21_X1 U8826 ( .B1(n6971), .B2(n8872), .A(n6970), .ZN(n6972) );
  OAI21_X1 U8827 ( .B1(n10129), .B2(n6973), .A(n6972), .ZN(P2_U3184) );
  AOI21_X1 U8828 ( .B1(n6975), .B2(n6974), .A(n7052), .ZN(n6988) );
  INV_X1 U8829 ( .A(n6976), .ZN(n6986) );
  INV_X1 U8830 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n6977) );
  OAI22_X1 U8831 ( .A1(n8870), .A2(n6977), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7282), .ZN(n6985) );
  INV_X1 U8832 ( .A(n7058), .ZN(n6978) );
  AOI21_X1 U8833 ( .B1(n7284), .B2(n6979), .A(n6978), .ZN(n6983) );
  INV_X1 U8834 ( .A(n7064), .ZN(n6980) );
  AOI21_X1 U8835 ( .B1(n5347), .B2(n6981), .A(n6980), .ZN(n6982) );
  OAI22_X1 U8836 ( .A1(n10131), .A2(n6983), .B1(n6982), .B2(n10127), .ZN(n6984) );
  AOI211_X1 U8837 ( .C1(n6986), .C2(n8872), .A(n6985), .B(n6984), .ZN(n6987)
         );
  OAI21_X1 U8838 ( .B1(n6988), .B2(n10129), .A(n6987), .ZN(P2_U3185) );
  XNOR2_X1 U8839 ( .A(n6990), .B(n6989), .ZN(n7004) );
  INV_X1 U8840 ( .A(n6991), .ZN(n7002) );
  INV_X1 U8841 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n10217) );
  OAI22_X1 U8842 ( .A1(n8870), .A2(n10217), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n6992), .ZN(n7001) );
  INV_X1 U8843 ( .A(n6993), .ZN(n6994) );
  INV_X1 U8844 ( .A(n6995), .ZN(n6996) );
  AOI21_X1 U8845 ( .B1(n6925), .B2(n6997), .A(n6996), .ZN(n6998) );
  OAI22_X1 U8846 ( .A1(n10131), .A2(n6999), .B1(n6998), .B2(n10127), .ZN(n7000) );
  AOI211_X1 U8847 ( .C1(n7002), .C2(n8872), .A(n7001), .B(n7000), .ZN(n7003)
         );
  OAI21_X1 U8848 ( .B1(n10129), .B2(n7004), .A(n7003), .ZN(P2_U3183) );
  INV_X1 U8849 ( .A(n7005), .ZN(n8223) );
  OAI21_X1 U8850 ( .B1(n8223), .B2(n5751), .A(n7006), .ZN(n7237) );
  OAI21_X1 U8851 ( .B1(n7008), .B2(n7005), .A(n7007), .ZN(n7009) );
  AOI222_X1 U8852 ( .A1(n10151), .A2(n7009), .B1(n8743), .B2(n10148), .C1(
        n5317), .C2(n9025), .ZN(n7238) );
  INV_X1 U8853 ( .A(n7238), .ZN(n7010) );
  AOI21_X1 U8854 ( .B1(n10192), .B2(n7237), .A(n7010), .ZN(n7433) );
  OAI22_X1 U8855 ( .A1(n7011), .A2(n9148), .B1(n10199), .B2(n5321), .ZN(n7012)
         );
  INV_X1 U8856 ( .A(n7012), .ZN(n7013) );
  OAI21_X1 U8857 ( .B1(n7433), .B2(n10201), .A(n7013), .ZN(P2_U3393) );
  NAND3_X1 U8858 ( .A1(n7014), .A2(n7016), .A3(n4508), .ZN(n7019) );
  INV_X1 U8859 ( .A(n8514), .ZN(n7017) );
  OR2_X1 U8860 ( .A1(n4508), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n7015) );
  NAND2_X1 U8861 ( .A1(n7016), .A2(n7015), .ZN(n9953) );
  AOI22_X1 U8862 ( .A1(n7017), .A2(n9427), .B1(n9953), .B2(n10397), .ZN(n7018)
         );
  NAND3_X1 U8863 ( .A1(n7019), .A2(P1_U3973), .A3(n7018), .ZN(n9447) );
  OAI211_X1 U8864 ( .C1(n7022), .C2(n7021), .A(n9499), .B(n7020), .ZN(n7030)
         );
  AND2_X1 U8865 ( .A1(P1_U3086), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n7352) );
  AOI21_X1 U8866 ( .B1(n9956), .B2(P1_ADDR_REG_4__SCAN_IN), .A(n7352), .ZN(
        n7029) );
  NAND2_X1 U8867 ( .A1(n9516), .A2(n7023), .ZN(n7028) );
  OAI211_X1 U8868 ( .C1(n7026), .C2(n7025), .A(n9517), .B(n7024), .ZN(n7027)
         );
  AND4_X1 U8869 ( .A1(n7030), .A2(n7029), .A3(n7028), .A4(n7027), .ZN(n7031)
         );
  NAND2_X1 U8870 ( .A1(n9447), .A2(n7031), .ZN(P1_U3247) );
  INV_X1 U8871 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n10586) );
  INV_X1 U8872 ( .A(n7032), .ZN(n7034) );
  OAI222_X1 U8873 ( .A1(n9903), .A2(n10586), .B1(n9905), .B2(n7034), .C1(
        P1_U3086), .C2(n4737), .ZN(P1_U3340) );
  INV_X1 U8874 ( .A(n8789), .ZN(n8765) );
  INV_X1 U8875 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n7033) );
  OAI222_X1 U8876 ( .A1(n8765), .A2(P2_U3151), .B1(n9171), .B2(n7034), .C1(
        n7033), .C2(n8539), .ZN(P2_U3280) );
  OAI21_X1 U8877 ( .B1(P1_REG2_REG_9__SCAN_IN), .B2(n7040), .A(n7035), .ZN(
        n7038) );
  NAND2_X1 U8878 ( .A1(n7226), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n7036) );
  OAI21_X1 U8879 ( .B1(n7226), .B2(P1_REG2_REG_10__SCAN_IN), .A(n7036), .ZN(
        n7037) );
  NOR2_X1 U8880 ( .A1(n7037), .A2(n7038), .ZN(n7221) );
  AOI211_X1 U8881 ( .C1(n7038), .C2(n7037), .A(n7221), .B(n7891), .ZN(n7048)
         );
  NAND2_X1 U8882 ( .A1(n7226), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n7041) );
  OAI21_X1 U8883 ( .B1(n7226), .B2(P1_REG1_REG_10__SCAN_IN), .A(n7041), .ZN(
        n7042) );
  AOI211_X1 U8884 ( .C1(n7043), .C2(n7042), .A(n7225), .B(n9510), .ZN(n7047)
         );
  INV_X1 U8885 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n7045) );
  NAND2_X1 U8886 ( .A1(n9516), .A2(n7226), .ZN(n7044) );
  NAND2_X1 U8887 ( .A1(P1_U3086), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n9911) );
  OAI211_X1 U8888 ( .C1(n7045), .C2(n9507), .A(n7044), .B(n9911), .ZN(n7046)
         );
  OR3_X1 U8889 ( .A1(n7048), .A2(n7047), .A3(n7046), .ZN(P1_U3253) );
  INV_X1 U8890 ( .A(n7049), .ZN(n7054) );
  OAI21_X1 U8891 ( .B1(n7052), .B2(n7051), .A(n7050), .ZN(n7053) );
  NAND3_X1 U8892 ( .A1(n7054), .A2(n8814), .A3(n7053), .ZN(n7072) );
  INV_X1 U8893 ( .A(n7055), .ZN(n7057) );
  NAND3_X1 U8894 ( .A1(n7058), .A2(n7057), .A3(n7056), .ZN(n7059) );
  AOI21_X1 U8895 ( .B1(n7060), .B2(n7059), .A(n10131), .ZN(n7070) );
  INV_X1 U8896 ( .A(n7061), .ZN(n7063) );
  NAND3_X1 U8897 ( .A1(n7064), .A2(n7063), .A3(n7062), .ZN(n7065) );
  AOI21_X1 U8898 ( .B1(n7066), .B2(n7065), .A(n10127), .ZN(n7069) );
  INV_X1 U8899 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n7067) );
  NAND2_X1 U8900 ( .A1(P2_U3151), .A2(P2_REG3_REG_4__SCAN_IN), .ZN(n7121) );
  OAI21_X1 U8901 ( .B1(n8870), .B2(n7067), .A(n7121), .ZN(n7068) );
  NOR3_X1 U8902 ( .A1(n7070), .A2(n7069), .A3(n7068), .ZN(n7071) );
  OAI211_X1 U8903 ( .C1(n10136), .C2(n7073), .A(n7072), .B(n7071), .ZN(
        P2_U3186) );
  XNOR2_X1 U8904 ( .A(n7114), .B(n10149), .ZN(n7085) );
  NAND2_X1 U8905 ( .A1(n7076), .A2(n7075), .ZN(n7080) );
  NAND2_X1 U8906 ( .A1(n7078), .A2(n7077), .ZN(n7079) );
  NAND2_X1 U8907 ( .A1(n7080), .A2(n7079), .ZN(n7084) );
  INV_X1 U8908 ( .A(n7084), .ZN(n7082) );
  INV_X1 U8909 ( .A(n7116), .ZN(n7083) );
  AOI211_X1 U8910 ( .C1(n7085), .C2(n7084), .A(n8658), .B(n7083), .ZN(n7091)
         );
  OR2_X1 U8911 ( .A1(n7086), .A2(P2_U3151), .ZN(n8271) );
  INV_X1 U8912 ( .A(n8709), .ZN(n8722) );
  MUX2_X1 U8913 ( .A(n8722), .B(P2_STATE_REG_SCAN_IN), .S(
        P2_REG3_REG_3__SCAN_IN), .Z(n7089) );
  INV_X1 U8914 ( .A(n8677), .ZN(n8720) );
  AOI22_X1 U8915 ( .A1(n8720), .A2(n8743), .B1(n8655), .B2(n10165), .ZN(n7088)
         );
  OAI211_X1 U8916 ( .C1(n7308), .C2(n8707), .A(n7089), .B(n7088), .ZN(n7090)
         );
  OR2_X1 U8917 ( .A1(n7091), .A2(n7090), .ZN(P2_U3158) );
  OAI21_X1 U8918 ( .B1(n7092), .B2(n7094), .A(n7093), .ZN(n7095) );
  NAND2_X1 U8919 ( .A1(n7095), .A2(n9948), .ZN(n7099) );
  INV_X1 U8920 ( .A(n5927), .ZN(n7097) );
  INV_X1 U8921 ( .A(n7096), .ZN(n7289) );
  OAI22_X1 U8922 ( .A1(n7097), .A2(n9537), .B1(n7289), .B2(n9338), .ZN(n9985)
         );
  AOI22_X1 U8923 ( .A1(n9985), .A2(n4510), .B1(P1_REG3_REG_1__SCAN_IN), .B2(
        n7189), .ZN(n7098) );
  OAI211_X1 U8924 ( .C1(n4998), .C2(n9946), .A(n7099), .B(n7098), .ZN(P1_U3222) );
  INV_X1 U8925 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n7113) );
  NAND3_X1 U8926 ( .A1(n7102), .A2(n7101), .A3(n7100), .ZN(n7109) );
  INV_X2 U8927 ( .A(n10000), .ZN(n9742) );
  NAND3_X1 U8928 ( .A1(n8457), .A2(n8513), .A3(n7103), .ZN(n7105) );
  OAI211_X1 U8929 ( .C1(n9970), .C2(n7106), .A(n7105), .B(n7104), .ZN(n7107)
         );
  NAND2_X1 U8930 ( .A1(n7107), .A2(n9742), .ZN(n7112) );
  NOR2_X1 U8931 ( .A1(n9612), .A2(n9831), .ZN(n9709) );
  OAI21_X1 U8932 ( .B1(n9633), .B2(n9709), .A(n7110), .ZN(n7111) );
  OAI211_X1 U8933 ( .C1(n7113), .C2(n9742), .A(n7112), .B(n7111), .ZN(P1_U3293) );
  XNOR2_X1 U8934 ( .A(n7273), .B(n7074), .ZN(n7243) );
  XNOR2_X1 U8935 ( .A(n7243), .B(n8742), .ZN(n7120) );
  NAND2_X1 U8936 ( .A1(n7114), .A2(n10149), .ZN(n7115) );
  INV_X1 U8937 ( .A(n7246), .ZN(n7118) );
  AOI21_X1 U8938 ( .B1(n7120), .B2(n7119), .A(n7118), .ZN(n7125) );
  INV_X1 U8939 ( .A(n7273), .ZN(n10170) );
  AOI22_X1 U8940 ( .A1(n8720), .A2(n10149), .B1(n8725), .B2(n7458), .ZN(n7122)
         );
  OAI211_X1 U8941 ( .C1(n10170), .C2(n8728), .A(n7122), .B(n7121), .ZN(n7123)
         );
  AOI21_X1 U8942 ( .B1(n7272), .B2(n8709), .A(n7123), .ZN(n7124) );
  OAI21_X1 U8943 ( .B1(n7125), .B2(n8658), .A(n7124), .ZN(P2_U3170) );
  XNOR2_X1 U8944 ( .A(n7147), .B(P2_REG2_REG_6__SCAN_IN), .ZN(n7163) );
  INV_X1 U8945 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n7460) );
  OR2_X1 U8946 ( .A1(n7147), .A2(n7460), .ZN(n7127) );
  INV_X1 U8947 ( .A(n7197), .ZN(n7128) );
  AOI21_X1 U8948 ( .B1(n7137), .B2(n7129), .A(n7128), .ZN(n7159) );
  INV_X1 U8949 ( .A(n7130), .ZN(n7131) );
  OAI22_X1 U8950 ( .A1(n7133), .A2(n7132), .B1(n4950), .B2(n7131), .ZN(n7162)
         );
  INV_X1 U8951 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n7146) );
  MUX2_X1 U8952 ( .A(n7460), .B(n7146), .S(n8860), .Z(n7134) );
  NAND2_X1 U8953 ( .A1(n7134), .A2(n7147), .ZN(n7135) );
  OAI21_X1 U8954 ( .B1(n7134), .B2(n7147), .A(n7135), .ZN(n7161) );
  NOR2_X1 U8955 ( .A1(n7162), .A2(n7161), .ZN(n7160) );
  INV_X1 U8956 ( .A(n7135), .ZN(n7142) );
  MUX2_X1 U8957 ( .A(n7137), .B(n7136), .S(n8860), .Z(n7138) );
  NAND2_X1 U8958 ( .A1(n7138), .A2(n7156), .ZN(n7204) );
  INV_X1 U8959 ( .A(n7138), .ZN(n7139) );
  NAND2_X1 U8960 ( .A1(n7139), .A2(n7149), .ZN(n7140) );
  AND2_X1 U8961 ( .A1(n7204), .A2(n7140), .ZN(n7141) );
  OAI21_X1 U8962 ( .B1(n7160), .B2(n7142), .A(n7141), .ZN(n7205) );
  INV_X1 U8963 ( .A(n7205), .ZN(n7144) );
  NOR3_X1 U8964 ( .A1(n7160), .A2(n7142), .A3(n7141), .ZN(n7143) );
  OAI21_X1 U8965 ( .B1(n7144), .B2(n7143), .A(n8814), .ZN(n7158) );
  NAND2_X1 U8966 ( .A1(n7174), .A2(n7173), .ZN(n7145) );
  XNOR2_X1 U8967 ( .A(n7147), .B(P2_REG1_REG_6__SCAN_IN), .ZN(n7172) );
  OR2_X1 U8968 ( .A1(n7147), .A2(n7146), .ZN(n7148) );
  NAND2_X1 U8969 ( .A1(n7150), .A2(n7136), .ZN(n7151) );
  AOI21_X1 U8970 ( .B1(n7211), .B2(n7151), .A(n10127), .ZN(n7155) );
  INV_X1 U8971 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n7153) );
  NOR2_X1 U8972 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n5153), .ZN(n7448) );
  INV_X1 U8973 ( .A(n7448), .ZN(n7152) );
  OAI21_X1 U8974 ( .B1(n8870), .B2(n7153), .A(n7152), .ZN(n7154) );
  AOI211_X1 U8975 ( .C1(n8872), .C2(n7156), .A(n7155), .B(n7154), .ZN(n7157)
         );
  OAI211_X1 U8976 ( .C1(n7159), .C2(n10131), .A(n7158), .B(n7157), .ZN(
        P2_U3189) );
  AOI21_X1 U8977 ( .B1(n7162), .B2(n7161), .A(n7160), .ZN(n7181) );
  INV_X1 U8978 ( .A(n7163), .ZN(n7165) );
  NAND3_X1 U8979 ( .A1(n7166), .A2(n7165), .A3(n7164), .ZN(n7167) );
  AOI21_X1 U8980 ( .B1(n7168), .B2(n7167), .A(n10131), .ZN(n7179) );
  INV_X1 U8981 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n10529) );
  NOR2_X1 U8982 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10529), .ZN(n7302) );
  INV_X1 U8983 ( .A(n7302), .ZN(n7170) );
  NAND2_X1 U8984 ( .A1(n10118), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n7169) );
  OAI211_X1 U8985 ( .C1(n10136), .C2(n7171), .A(n7170), .B(n7169), .ZN(n7178)
         );
  NAND3_X1 U8986 ( .A1(n7174), .A2(n4850), .A3(n7173), .ZN(n7175) );
  AOI21_X1 U8987 ( .B1(n7176), .B2(n7175), .A(n10127), .ZN(n7177) );
  NOR3_X1 U8988 ( .A1(n7179), .A2(n7178), .A3(n7177), .ZN(n7180) );
  OAI21_X1 U8989 ( .B1(n7181), .B2(n10129), .A(n7180), .ZN(P2_U3188) );
  NAND2_X1 U8990 ( .A1(n8958), .A2(P2_U3893), .ZN(n7182) );
  OAI21_X1 U8991 ( .B1(P2_U3893), .B2(n5280), .A(n7182), .ZN(P2_U3514) );
  INV_X1 U8992 ( .A(n8784), .ZN(n8810) );
  INV_X1 U8993 ( .A(n7183), .ZN(n7220) );
  INV_X1 U8994 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n7184) );
  OAI222_X1 U8995 ( .A1(P2_U3151), .A2(n8810), .B1(n9171), .B2(n7220), .C1(
        n7184), .C2(n8539), .ZN(P2_U3279) );
  XNOR2_X1 U8996 ( .A(n7186), .B(n7185), .ZN(n7187) );
  NAND2_X1 U8997 ( .A1(n7187), .A2(n9948), .ZN(n7191) );
  INV_X1 U8998 ( .A(n9421), .ZN(n7350) );
  INV_X1 U8999 ( .A(n5914), .ZN(n7188) );
  OAI22_X1 U9000 ( .A1(n7350), .A2(n9338), .B1(n7188), .B2(n9537), .ZN(n7255)
         );
  AOI22_X1 U9001 ( .A1(n7255), .A2(n4510), .B1(P1_REG3_REG_2__SCAN_IN), .B2(
        n7189), .ZN(n7190) );
  OAI211_X1 U9002 ( .C1(n10011), .C2(n9946), .A(n7191), .B(n7190), .ZN(
        P1_U3237) );
  INV_X1 U9003 ( .A(n7193), .ZN(n7192) );
  XNOR2_X1 U9004 ( .A(n7332), .B(P2_REG2_REG_8__SCAN_IN), .ZN(n7194) );
  NOR2_X1 U9005 ( .A1(n7192), .A2(n7194), .ZN(n7198) );
  NAND2_X1 U9006 ( .A1(n7197), .A2(n7193), .ZN(n7195) );
  NAND2_X1 U9007 ( .A1(n7195), .A2(n7194), .ZN(n7317) );
  INV_X1 U9008 ( .A(n7317), .ZN(n7196) );
  AOI21_X1 U9009 ( .B1(n7198), .B2(n7197), .A(n7196), .ZN(n7219) );
  MUX2_X1 U9010 ( .A(n7315), .B(n10209), .S(n8860), .Z(n7199) );
  NAND2_X1 U9011 ( .A1(n7199), .A2(n7332), .ZN(n7321) );
  INV_X1 U9012 ( .A(n7199), .ZN(n7201) );
  NAND2_X1 U9013 ( .A1(n7201), .A2(n7200), .ZN(n7202) );
  NAND2_X1 U9014 ( .A1(n7321), .A2(n7202), .ZN(n7203) );
  AOI21_X1 U9015 ( .B1(n7205), .B2(n7204), .A(n7203), .ZN(n7329) );
  AND3_X1 U9016 ( .A1(n7205), .A2(n7204), .A3(n7203), .ZN(n7206) );
  OAI21_X1 U9017 ( .B1(n7329), .B2(n7206), .A(n8814), .ZN(n7218) );
  NAND2_X1 U9018 ( .A1(n7211), .A2(n7209), .ZN(n7207) );
  XNOR2_X1 U9019 ( .A(n7332), .B(P2_REG1_REG_8__SCAN_IN), .ZN(n7208) );
  NAND2_X1 U9020 ( .A1(n7207), .A2(n7208), .ZN(n7334) );
  INV_X1 U9021 ( .A(n7208), .ZN(n7210) );
  NAND3_X1 U9022 ( .A1(n7211), .A2(n7210), .A3(n7209), .ZN(n7212) );
  AOI21_X1 U9023 ( .B1(n7334), .B2(n7212), .A(n10127), .ZN(n7216) );
  INV_X1 U9024 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n7214) );
  INV_X1 U9025 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n10533) );
  NOR2_X1 U9026 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10533), .ZN(n7588) );
  INV_X1 U9027 ( .A(n7588), .ZN(n7213) );
  OAI21_X1 U9028 ( .B1(n8870), .B2(n7214), .A(n7213), .ZN(n7215) );
  AOI211_X1 U9029 ( .C1(n8872), .C2(n7332), .A(n7216), .B(n7215), .ZN(n7217)
         );
  OAI211_X1 U9030 ( .C1(n7219), .C2(n10131), .A(n7218), .B(n7217), .ZN(
        P2_U3190) );
  INV_X1 U9031 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n10387) );
  INV_X1 U9032 ( .A(n8528), .ZN(n7884) );
  OAI222_X1 U9033 ( .A1(n9903), .A2(n10387), .B1(n7884), .B2(P1_U3086), .C1(
        n9905), .C2(n7220), .ZN(P1_U3339) );
  AOI21_X1 U9034 ( .B1(P1_REG2_REG_10__SCAN_IN), .B2(n7226), .A(n7221), .ZN(
        n7224) );
  NAND2_X1 U9035 ( .A1(n7360), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n7222) );
  OAI21_X1 U9036 ( .B1(n7360), .B2(P1_REG2_REG_11__SCAN_IN), .A(n7222), .ZN(
        n7223) );
  NOR2_X1 U9037 ( .A1(n7224), .A2(n7223), .ZN(n7359) );
  AOI211_X1 U9038 ( .C1(n7224), .C2(n7223), .A(n7359), .B(n7891), .ZN(n7234)
         );
  AOI21_X1 U9039 ( .B1(n7226), .B2(P1_REG1_REG_10__SCAN_IN), .A(n7225), .ZN(
        n7229) );
  MUX2_X1 U9040 ( .A(n7227), .B(P1_REG1_REG_11__SCAN_IN), .S(n7360), .Z(n7228)
         );
  NOR2_X1 U9041 ( .A1(n7229), .A2(n7228), .ZN(n7355) );
  AOI211_X1 U9042 ( .C1(n7229), .C2(n7228), .A(n7355), .B(n9510), .ZN(n7233)
         );
  INV_X1 U9043 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n7231) );
  NAND2_X1 U9044 ( .A1(n9516), .A2(n7360), .ZN(n7230) );
  NAND2_X1 U9045 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_U3086), .ZN(n9351) );
  OAI211_X1 U9046 ( .C1(n7231), .C2(n9507), .A(n7230), .B(n9351), .ZN(n7232)
         );
  OR3_X1 U9047 ( .A1(n7234), .A2(n7233), .A3(n7232), .ZN(P1_U3254) );
  NAND2_X1 U9048 ( .A1(n7235), .A2(n4511), .ZN(n7236) );
  OAI21_X1 U9049 ( .B1(n4511), .B2(n8540), .A(n7236), .ZN(P1_U3581) );
  INV_X1 U9050 ( .A(n7237), .ZN(n7242) );
  MUX2_X1 U9051 ( .A(n7239), .B(n7238), .S(n9029), .Z(n7241) );
  AOI22_X1 U9052 ( .A1(n9032), .A2(n7431), .B1(n9031), .B2(
        P2_REG3_REG_1__SCAN_IN), .ZN(n7240) );
  OAI211_X1 U9053 ( .C1(n9035), .C2(n7242), .A(n7241), .B(n7240), .ZN(P2_U3232) );
  INV_X1 U9054 ( .A(n7243), .ZN(n7244) );
  NAND2_X1 U9055 ( .A1(n7308), .A2(n7244), .ZN(n7245) );
  NAND2_X1 U9056 ( .A1(n7246), .A2(n7245), .ZN(n7298) );
  XNOR2_X1 U9057 ( .A(n7428), .B(n8580), .ZN(n7294) );
  XNOR2_X1 U9058 ( .A(n7294), .B(n7458), .ZN(n7297) );
  XOR2_X1 U9059 ( .A(n7298), .B(n7297), .Z(n7253) );
  INV_X1 U9060 ( .A(n7434), .ZN(n7251) );
  AOI21_X1 U9061 ( .B1(n8720), .B2(n8742), .A(n7247), .ZN(n7249) );
  NAND2_X1 U9062 ( .A1(n8655), .A2(n7428), .ZN(n7248) );
  OAI211_X1 U9063 ( .C1(n7501), .C2(n8707), .A(n7249), .B(n7248), .ZN(n7250)
         );
  AOI21_X1 U9064 ( .B1(n7251), .B2(n8709), .A(n7250), .ZN(n7252) );
  OAI21_X1 U9065 ( .B1(n7253), .B2(n8658), .A(n7252), .ZN(P2_U3167) );
  XOR2_X1 U9066 ( .A(n8460), .B(n7254), .Z(n7256) );
  AOI21_X1 U9067 ( .B1(n7256), .B2(n9837), .A(n7255), .ZN(n10012) );
  AOI211_X1 U9068 ( .C1(n7257), .C2(n9992), .A(n9831), .B(n7407), .ZN(n10009)
         );
  NOR2_X1 U9069 ( .A1(n9990), .A2(n10011), .ZN(n7259) );
  OAI22_X1 U9070 ( .A1(n9742), .A2(n5937), .B1(n9433), .B2(n9970), .ZN(n7258)
         );
  AOI211_X1 U9071 ( .C1(n10009), .C2(n9996), .A(n7259), .B(n7258), .ZN(n7264)
         );
  XNOR2_X1 U9072 ( .A(n7260), .B(n8460), .ZN(n10015) );
  NAND3_X1 U9073 ( .A1(n8456), .A2(n7528), .A3(n4509), .ZN(n7261) );
  OR2_X1 U9074 ( .A1(n10000), .A2(n9960), .ZN(n7262) );
  NAND2_X1 U9075 ( .A1(n10015), .A2(n9929), .ZN(n7263) );
  OAI211_X1 U9076 ( .C1(n10012), .C2(n9988), .A(n7264), .B(n7263), .ZN(
        P1_U3291) );
  INV_X1 U9077 ( .A(n8220), .ZN(n7265) );
  XNOR2_X1 U9078 ( .A(n7266), .B(n7265), .ZN(n7267) );
  NAND2_X1 U9079 ( .A1(n7267), .A2(n10151), .ZN(n7269) );
  AOI22_X1 U9080 ( .A1(n9025), .A2(n10149), .B1(n7458), .B2(n10148), .ZN(n7268) );
  NAND2_X1 U9081 ( .A1(n7269), .A2(n7268), .ZN(n10171) );
  INV_X1 U9082 ( .A(n10171), .ZN(n7278) );
  OAI21_X1 U9083 ( .B1(n7271), .B2(n8220), .A(n7270), .ZN(n10173) );
  INV_X1 U9084 ( .A(n9035), .ZN(n8021) );
  AOI22_X1 U9085 ( .A1(n9032), .A2(n7273), .B1(n9031), .B2(n7272), .ZN(n7274)
         );
  OAI21_X1 U9086 ( .B1(n7275), .B2(n9029), .A(n7274), .ZN(n7276) );
  AOI21_X1 U9087 ( .B1(n10173), .B2(n8021), .A(n7276), .ZN(n7277) );
  OAI21_X1 U9088 ( .B1(n7278), .B2(n10159), .A(n7277), .ZN(P2_U3229) );
  XOR2_X1 U9089 ( .A(n7279), .B(n8222), .Z(n7280) );
  AOI222_X1 U9090 ( .A1(n10151), .A2(n7280), .B1(n8742), .B2(n10148), .C1(
        n8743), .C2(n9025), .ZN(n10168) );
  XNOR2_X1 U9091 ( .A(n7281), .B(n8222), .ZN(n10166) );
  AOI22_X1 U9092 ( .A1(n9032), .A2(n10165), .B1(n9031), .B2(n7282), .ZN(n7283)
         );
  OAI21_X1 U9093 ( .B1(n7284), .B2(n9029), .A(n7283), .ZN(n7285) );
  AOI21_X1 U9094 ( .B1(n10166), .B2(n8021), .A(n7285), .ZN(n7286) );
  OAI21_X1 U9095 ( .B1(n10168), .B2(n10159), .A(n7286), .ZN(P2_U3230) );
  XOR2_X1 U9096 ( .A(n7288), .B(n7287), .Z(n7293) );
  INV_X1 U9097 ( .A(n7416), .ZN(n7290) );
  OAI22_X1 U9098 ( .A1(n7290), .A2(n9338), .B1(n7289), .B2(n9537), .ZN(n7403)
         );
  AOI22_X1 U9099 ( .A1(n7409), .A2(n9395), .B1(n7403), .B2(n4510), .ZN(n7292)
         );
  MUX2_X1 U9100 ( .A(n9920), .B(P1_STATE_REG_SCAN_IN), .S(
        P1_REG3_REG_3__SCAN_IN), .Z(n7291) );
  OAI211_X1 U9101 ( .C1(n7293), .C2(n9916), .A(n7292), .B(n7291), .ZN(P1_U3218) );
  INV_X1 U9102 ( .A(n7461), .ZN(n7305) );
  INV_X1 U9103 ( .A(n7294), .ZN(n7295) );
  NOR2_X1 U9104 ( .A1(n7295), .A2(n7458), .ZN(n7296) );
  XNOR2_X1 U9105 ( .A(n10177), .B(n8580), .ZN(n7441) );
  XNOR2_X1 U9106 ( .A(n7441), .B(n7501), .ZN(n7299) );
  OAI211_X1 U9107 ( .C1(n7300), .C2(n7299), .A(n7443), .B(n8717), .ZN(n7304)
         );
  OAI22_X1 U9108 ( .A1(n10177), .A2(n8728), .B1(n7540), .B2(n8707), .ZN(n7301)
         );
  AOI211_X1 U9109 ( .C1(n8720), .C2(n7458), .A(n7302), .B(n7301), .ZN(n7303)
         );
  OAI211_X1 U9110 ( .C1(n7305), .C2(n8722), .A(n7304), .B(n7303), .ZN(P2_U3179) );
  XNOR2_X1 U9111 ( .A(n7458), .B(n7435), .ZN(n8225) );
  XNOR2_X1 U9112 ( .A(n7306), .B(n8225), .ZN(n7307) );
  OAI222_X1 U9113 ( .A1(n9008), .A2(n7501), .B1(n9006), .B2(n7308), .C1(n9003), 
        .C2(n7307), .ZN(n7436) );
  AOI21_X1 U9114 ( .B1(n10192), .B2(n7439), .A(n7436), .ZN(n7430) );
  INV_X1 U9115 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n7309) );
  OAI22_X1 U9116 ( .A1(n7435), .A2(n9148), .B1(n10199), .B2(n7309), .ZN(n7310)
         );
  INV_X1 U9117 ( .A(n7310), .ZN(n7311) );
  OAI21_X1 U9118 ( .B1(n7430), .B2(n10201), .A(n7311), .ZN(P2_U3405) );
  INV_X1 U9119 ( .A(n7312), .ZN(n7314) );
  INV_X1 U9120 ( .A(n9501), .ZN(n8526) );
  OAI222_X1 U9121 ( .A1(n9903), .A2(n10347), .B1(n9905), .B2(n7314), .C1(
        P1_U3086), .C2(n8526), .ZN(P1_U3338) );
  INV_X1 U9122 ( .A(n8841), .ZN(n8802) );
  OAI222_X1 U9123 ( .A1(n8802), .A2(P2_U3151), .B1(n9171), .B2(n7314), .C1(
        n7313), .C2(n8539), .ZN(P2_U3278) );
  OR2_X1 U9124 ( .A1(n7332), .A2(n7315), .ZN(n7316) );
  NAND2_X1 U9125 ( .A1(n7317), .A2(n7316), .ZN(n7319) );
  OAI21_X1 U9126 ( .B1(n7339), .B2(n7319), .A(n7318), .ZN(n7320) );
  INV_X1 U9127 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n7624) );
  NOR2_X1 U9128 ( .A1(n7624), .A2(n7320), .ZN(n7378) );
  AOI21_X1 U9129 ( .B1(n7320), .B2(n7624), .A(n7378), .ZN(n7344) );
  INV_X1 U9130 ( .A(n7321), .ZN(n7328) );
  MUX2_X1 U9131 ( .A(n7624), .B(n7322), .S(n8860), .Z(n7324) );
  NAND2_X1 U9132 ( .A1(n7324), .A2(n7323), .ZN(n7375) );
  INV_X1 U9133 ( .A(n7324), .ZN(n7325) );
  NAND2_X1 U9134 ( .A1(n7325), .A2(n7339), .ZN(n7326) );
  AND2_X1 U9135 ( .A1(n7375), .A2(n7326), .ZN(n7327) );
  OAI21_X1 U9136 ( .B1(n7329), .B2(n7328), .A(n7327), .ZN(n7376) );
  INV_X1 U9137 ( .A(n7376), .ZN(n7331) );
  NOR3_X1 U9138 ( .A1(n7329), .A2(n7328), .A3(n7327), .ZN(n7330) );
  OAI21_X1 U9139 ( .B1(n7331), .B2(n7330), .A(n8814), .ZN(n7343) );
  OR2_X1 U9140 ( .A1(n7332), .A2(n10209), .ZN(n7333) );
  NAND2_X1 U9141 ( .A1(n7334), .A2(n7333), .ZN(n7335) );
  AOI21_X1 U9142 ( .B1(n7336), .B2(n7322), .A(n7365), .ZN(n7337) );
  NOR2_X1 U9143 ( .A1(n7337), .A2(n10127), .ZN(n7341) );
  NOR2_X1 U9144 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n5155), .ZN(n7548) );
  INV_X1 U9145 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n7338) );
  OAI22_X1 U9146 ( .A1(n10136), .A2(n7339), .B1(n8870), .B2(n7338), .ZN(n7340)
         );
  NOR3_X1 U9147 ( .A1(n7341), .A2(n7548), .A3(n7340), .ZN(n7342) );
  OAI211_X1 U9148 ( .C1(n7344), .C2(n10131), .A(n7343), .B(n7342), .ZN(
        P2_U3191) );
  AOI21_X1 U9149 ( .B1(n7345), .B2(n7346), .A(n9916), .ZN(n7348) );
  NAND2_X1 U9150 ( .A1(n7348), .A2(n7347), .ZN(n7354) );
  INV_X1 U9151 ( .A(n9420), .ZN(n7349) );
  OAI22_X1 U9152 ( .A1(n7350), .A2(n9537), .B1(n7349), .B2(n9338), .ZN(n7393)
         );
  NOR2_X1 U9153 ( .A1(n9946), .A2(n10024), .ZN(n7351) );
  AOI211_X1 U9154 ( .C1(n4510), .C2(n7393), .A(n7352), .B(n7351), .ZN(n7353)
         );
  OAI211_X1 U9155 ( .C1(n9920), .C2(n7399), .A(n7354), .B(n7353), .ZN(P1_U3230) );
  MUX2_X1 U9156 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n7487), .S(n7358), .Z(n7356)
         );
  OAI21_X1 U9157 ( .B1(n7357), .B2(n7356), .A(n7490), .ZN(n7362) );
  XNOR2_X1 U9158 ( .A(n7358), .B(n7814), .ZN(n7482) );
  XNOR2_X1 U9159 ( .A(n7482), .B(n7481), .ZN(n7361) );
  AOI22_X1 U9160 ( .A1(n9499), .A2(n7362), .B1(n9517), .B2(n7361), .ZN(n7364)
         );
  AND2_X1 U9161 ( .A1(P1_U3086), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n9247) );
  AOI21_X1 U9162 ( .B1(n9956), .B2(P1_ADDR_REG_12__SCAN_IN), .A(n9247), .ZN(
        n7363) );
  OAI211_X1 U9163 ( .C1(n7488), .C2(n7885), .A(n7364), .B(n7363), .ZN(P1_U3255) );
  NAND2_X1 U9164 ( .A1(P2_REG1_REG_10__SCAN_IN), .A2(n7577), .ZN(n7367) );
  OAI21_X1 U9165 ( .B1(P2_REG1_REG_10__SCAN_IN), .B2(n7577), .A(n7367), .ZN(
        n7368) );
  NOR2_X1 U9166 ( .A1(n7369), .A2(n7368), .ZN(n7568) );
  AOI21_X1 U9167 ( .B1(n7369), .B2(n7368), .A(n7568), .ZN(n7389) );
  MUX2_X1 U9168 ( .A(n7774), .B(n7370), .S(n8860), .Z(n7371) );
  NAND2_X1 U9169 ( .A1(n7371), .A2(n7382), .ZN(n7570) );
  INV_X1 U9170 ( .A(n7371), .ZN(n7372) );
  NAND2_X1 U9171 ( .A1(n7372), .A2(n7577), .ZN(n7373) );
  NAND2_X1 U9172 ( .A1(n7570), .A2(n7373), .ZN(n7374) );
  AOI21_X1 U9173 ( .B1(n7376), .B2(n7375), .A(n7374), .ZN(n7572) );
  AND3_X1 U9174 ( .A1(n7376), .A2(n7375), .A3(n7374), .ZN(n7377) );
  OAI21_X1 U9175 ( .B1(n7572), .B2(n7377), .A(n8814), .ZN(n7388) );
  NAND2_X1 U9176 ( .A1(P2_REG2_REG_10__SCAN_IN), .A2(n7577), .ZN(n7379) );
  OAI21_X1 U9177 ( .B1(P2_REG2_REG_10__SCAN_IN), .B2(n7577), .A(n7379), .ZN(
        n7380) );
  AOI21_X1 U9178 ( .B1(n7381), .B2(n7380), .A(n7576), .ZN(n7385) );
  AOI22_X1 U9179 ( .A1(n8872), .A2(n7382), .B1(n10118), .B2(
        P2_ADDR_REG_10__SCAN_IN), .ZN(n7384) );
  INV_X1 U9180 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n10385) );
  NOR2_X1 U9181 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10385), .ZN(n7732) );
  INV_X1 U9182 ( .A(n7732), .ZN(n7383) );
  OAI211_X1 U9183 ( .C1(n7385), .C2(n10131), .A(n7384), .B(n7383), .ZN(n7386)
         );
  INV_X1 U9184 ( .A(n7386), .ZN(n7387) );
  OAI211_X1 U9185 ( .C1(n7389), .C2(n10127), .A(n7388), .B(n7387), .ZN(
        P2_U3192) );
  INV_X1 U9186 ( .A(n8458), .ZN(n7391) );
  XNOR2_X1 U9187 ( .A(n7390), .B(n7391), .ZN(n10023) );
  XOR2_X1 U9188 ( .A(n8458), .B(n7392), .Z(n7394) );
  AOI21_X1 U9189 ( .B1(n7394), .B2(n9837), .A(n7393), .ZN(n10022) );
  MUX2_X1 U9190 ( .A(n7395), .B(n10022), .S(n9742), .Z(n7402) );
  AOI21_X1 U9191 ( .B1(n7406), .B2(n7396), .A(n9831), .ZN(n7398) );
  INV_X1 U9192 ( .A(n7397), .ZN(n7419) );
  AND2_X1 U9193 ( .A1(n7398), .A2(n7419), .ZN(n10026) );
  OAI22_X1 U9194 ( .A1(n9990), .A2(n10024), .B1(n9970), .B2(n7399), .ZN(n7400)
         );
  AOI21_X1 U9195 ( .B1(n10026), .B2(n9996), .A(n7400), .ZN(n7401) );
  OAI211_X1 U9196 ( .C1(n9726), .C2(n10023), .A(n7402), .B(n7401), .ZN(
        P1_U3289) );
  XNOR2_X1 U9197 ( .A(n8294), .B(n8459), .ZN(n7404) );
  AOI21_X1 U9198 ( .B1(n7404), .B2(n9837), .A(n7403), .ZN(n10018) );
  XNOR2_X1 U9199 ( .A(n7405), .B(n8459), .ZN(n10021) );
  OAI211_X1 U9200 ( .C1(n7407), .C2(n10017), .A(n7406), .B(n9993), .ZN(n10016)
         );
  INV_X1 U9201 ( .A(n9970), .ZN(n9987) );
  INV_X1 U9202 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n7408) );
  AOI22_X1 U9203 ( .A1(n9988), .A2(P1_REG2_REG_3__SCAN_IN), .B1(n9987), .B2(
        n7408), .ZN(n7411) );
  NAND2_X1 U9204 ( .A1(n9633), .A2(n7409), .ZN(n7410) );
  OAI211_X1 U9205 ( .C1(n10016), .C2(n9612), .A(n7411), .B(n7410), .ZN(n7412)
         );
  AOI21_X1 U9206 ( .B1(n10021), .B2(n9929), .A(n7412), .ZN(n7413) );
  OAI21_X1 U9207 ( .B1(n10018), .B2(n9988), .A(n7413), .ZN(P1_U3290) );
  XNOR2_X1 U9208 ( .A(n7414), .B(n7415), .ZN(n10033) );
  XNOR2_X1 U9209 ( .A(n8345), .B(n7415), .ZN(n7417) );
  AOI22_X1 U9210 ( .A1(n9199), .A2(n7416), .B1(n9419), .B2(n9368), .ZN(n7521)
         );
  OAI21_X1 U9211 ( .B1(n7417), .B2(n9982), .A(n7521), .ZN(n10035) );
  NAND2_X1 U9212 ( .A1(n10035), .A2(n9742), .ZN(n7425) );
  INV_X1 U9213 ( .A(n7418), .ZN(n7472) );
  AOI211_X1 U9214 ( .C1(n10031), .C2(n7419), .A(n9831), .B(n7472), .ZN(n10030)
         );
  NOR2_X1 U9215 ( .A1(n9990), .A2(n7420), .ZN(n7423) );
  OAI22_X1 U9216 ( .A1(n9742), .A2(n7421), .B1(n7525), .B2(n9970), .ZN(n7422)
         );
  AOI211_X1 U9217 ( .C1(n10030), .C2(n9996), .A(n7423), .B(n7422), .ZN(n7424)
         );
  OAI211_X1 U9218 ( .C1(n9726), .C2(n10033), .A(n7425), .B(n7424), .ZN(
        P1_U3288) );
  INV_X1 U9219 ( .A(n7426), .ZN(n7454) );
  INV_X1 U9220 ( .A(n8865), .ZN(n8822) );
  OAI222_X1 U9221 ( .A1(n8539), .A2(n7427), .B1(n9171), .B2(n7454), .C1(
        P2_U3151), .C2(n8822), .ZN(P2_U3277) );
  INV_X1 U9222 ( .A(n10213), .ZN(n10211) );
  AOI22_X1 U9223 ( .A1(n6647), .A2(n7428), .B1(n10211), .B2(
        P2_REG1_REG_5__SCAN_IN), .ZN(n7429) );
  OAI21_X1 U9224 ( .B1(n7430), .B2(n10211), .A(n7429), .ZN(P2_U3464) );
  AOI22_X1 U9225 ( .A1(n6647), .A2(n7431), .B1(n10211), .B2(
        P2_REG1_REG_1__SCAN_IN), .ZN(n7432) );
  OAI21_X1 U9226 ( .B1(n7433), .B2(n10211), .A(n7432), .ZN(P2_U3460) );
  OAI22_X1 U9227 ( .A1(n9014), .A2(n7435), .B1(n7434), .B2(n10141), .ZN(n7438)
         );
  MUX2_X1 U9228 ( .A(P2_REG2_REG_5__SCAN_IN), .B(n7436), .S(n9029), .Z(n7437)
         );
  AOI211_X1 U9229 ( .C1(n8021), .C2(n7439), .A(n7438), .B(n7437), .ZN(n7440)
         );
  INV_X1 U9230 ( .A(n7440), .ZN(P2_U3228) );
  XNOR2_X1 U9231 ( .A(n7507), .B(n8580), .ZN(n7541) );
  XNOR2_X1 U9232 ( .A(n7541), .B(n7540), .ZN(n7447) );
  NAND2_X1 U9233 ( .A1(n7441), .A2(n8741), .ZN(n7442) );
  INV_X1 U9234 ( .A(n7447), .ZN(n7444) );
  INV_X1 U9235 ( .A(n7543), .ZN(n7445) );
  AOI21_X1 U9236 ( .B1(n7447), .B2(n7446), .A(n7445), .ZN(n7453) );
  AOI21_X1 U9237 ( .B1(n8741), .B2(n8720), .A(n7448), .ZN(n7449) );
  OAI21_X1 U9238 ( .B1(n7621), .B2(n8707), .A(n7449), .ZN(n7451) );
  NOR2_X1 U9239 ( .A1(n8722), .A2(n7505), .ZN(n7450) );
  AOI211_X1 U9240 ( .C1(n7507), .C2(n8655), .A(n7451), .B(n7450), .ZN(n7452)
         );
  OAI21_X1 U9241 ( .B1(n7453), .B2(n8658), .A(n7452), .ZN(P2_U3153) );
  INV_X1 U9242 ( .A(n9515), .ZN(n7455) );
  OAI222_X1 U9243 ( .A1(n9903), .A2(n10395), .B1(n7455), .B2(P1_U3086), .C1(
        n9905), .C2(n7454), .ZN(P1_U3337) );
  XNOR2_X1 U9244 ( .A(n8741), .B(n10177), .ZN(n8226) );
  XOR2_X1 U9245 ( .A(n7456), .B(n8226), .Z(n10175) );
  XNOR2_X1 U9246 ( .A(n7457), .B(n8226), .ZN(n7459) );
  AOI222_X1 U9247 ( .A1(n10151), .A2(n7459), .B1(n8740), .B2(n10148), .C1(
        n7458), .C2(n9025), .ZN(n10176) );
  MUX2_X1 U9248 ( .A(n7460), .B(n10176), .S(n9029), .Z(n7464) );
  AOI22_X1 U9249 ( .A1(n9032), .A2(n7462), .B1(n9031), .B2(n7461), .ZN(n7463)
         );
  OAI211_X1 U9250 ( .C1(n9035), .C2(n10175), .A(n7464), .B(n7463), .ZN(
        P2_U3227) );
  NAND2_X1 U9251 ( .A1(n7465), .A2(n7477), .ZN(n7466) );
  NAND2_X1 U9252 ( .A1(n9964), .A2(n7466), .ZN(n7469) );
  OR2_X1 U9253 ( .A1(n7668), .A2(n9338), .ZN(n7468) );
  NAND2_X1 U9254 ( .A1(n9420), .A2(n9199), .ZN(n7467) );
  NAND2_X1 U9255 ( .A1(n7468), .A2(n7467), .ZN(n9381) );
  AOI21_X1 U9256 ( .B1(n7469), .B2(n9837), .A(n9381), .ZN(n10038) );
  OAI22_X1 U9257 ( .A1(n9742), .A2(n7470), .B1(n9382), .B2(n9970), .ZN(n7474)
         );
  INV_X1 U9258 ( .A(n9976), .ZN(n7471) );
  OAI211_X1 U9259 ( .C1(n10039), .C2(n7472), .A(n7471), .B(n9993), .ZN(n10037)
         );
  NOR2_X1 U9260 ( .A1(n10037), .A2(n9612), .ZN(n7473) );
  AOI211_X1 U9261 ( .C1(n9633), .C2(n7475), .A(n7474), .B(n7473), .ZN(n7479)
         );
  XNOR2_X1 U9262 ( .A(n7476), .B(n7477), .ZN(n10041) );
  NAND2_X1 U9263 ( .A1(n10041), .A2(n9929), .ZN(n7478) );
  OAI211_X1 U9264 ( .C1(n10038), .C2(n10000), .A(n7479), .B(n7478), .ZN(
        P1_U3287) );
  NAND2_X1 U9265 ( .A1(n7607), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n7480) );
  OAI21_X1 U9266 ( .B1(n7607), .B2(P1_REG2_REG_13__SCAN_IN), .A(n7480), .ZN(
        n7485) );
  AOI22_X1 U9267 ( .A1(n7482), .A2(n7481), .B1(n7488), .B2(n7814), .ZN(n7483)
         );
  INV_X1 U9268 ( .A(n7483), .ZN(n7484) );
  NOR2_X1 U9269 ( .A1(n7485), .A2(n7484), .ZN(n7602) );
  AOI211_X1 U9270 ( .C1(n7485), .C2(n7484), .A(n7602), .B(n7891), .ZN(n7497)
         );
  INV_X1 U9271 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n7486) );
  MUX2_X1 U9272 ( .A(n7486), .B(P1_REG1_REG_13__SCAN_IN), .S(n7607), .Z(n7492)
         );
  NAND2_X1 U9273 ( .A1(n7488), .A2(n7487), .ZN(n7489) );
  AOI211_X1 U9274 ( .C1(n7492), .C2(n7491), .A(n7606), .B(n9510), .ZN(n7496)
         );
  INV_X1 U9275 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n7494) );
  NAND2_X1 U9276 ( .A1(n9516), .A2(n7607), .ZN(n7493) );
  NAND2_X1 U9277 ( .A1(P1_REG3_REG_13__SCAN_IN), .A2(P1_U3086), .ZN(n9326) );
  OAI211_X1 U9278 ( .C1(n7494), .C2(n9507), .A(n7493), .B(n9326), .ZN(n7495)
         );
  OR3_X1 U9279 ( .A1(n7497), .A2(n7496), .A3(n7495), .ZN(P1_U3256) );
  XNOR2_X1 U9280 ( .A(n7498), .B(n8096), .ZN(n10183) );
  NAND2_X1 U9281 ( .A1(n9029), .A2(n7499), .ZN(n10155) );
  INV_X1 U9282 ( .A(n8096), .ZN(n8229) );
  XNOR2_X1 U9283 ( .A(n7500), .B(n8229), .ZN(n7503) );
  OAI22_X1 U9284 ( .A1(n7501), .A2(n9006), .B1(n7621), .B2(n9008), .ZN(n7502)
         );
  AOI21_X1 U9285 ( .B1(n7503), .B2(n10151), .A(n7502), .ZN(n7504) );
  OAI21_X1 U9286 ( .B1(n10183), .B2(n10137), .A(n7504), .ZN(n10185) );
  NAND2_X1 U9287 ( .A1(n10185), .A2(n9029), .ZN(n7509) );
  OAI22_X1 U9288 ( .A1(n9029), .A2(n7137), .B1(n7505), .B2(n10141), .ZN(n7506)
         );
  AOI21_X1 U9289 ( .B1(n9032), .B2(n7507), .A(n7506), .ZN(n7508) );
  OAI211_X1 U9290 ( .C1(n10183), .C2(n10155), .A(n7509), .B(n7508), .ZN(
        P2_U3226) );
  INV_X1 U9291 ( .A(P2_U3893), .ZN(n8832) );
  NAND2_X1 U9292 ( .A1(n8832), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n7510) );
  OAI21_X1 U9293 ( .B1(n8584), .B2(n8832), .A(n7510), .ZN(P2_U3520) );
  INV_X1 U9294 ( .A(n7511), .ZN(n7513) );
  OAI222_X1 U9295 ( .A1(n8859), .A2(P2_U3151), .B1(n9171), .B2(n7513), .C1(
        n7512), .C2(n8539), .ZN(P2_U3276) );
  OAI222_X1 U9296 ( .A1(n9903), .A2(n10406), .B1(n9905), .B2(n7513), .C1(
        P1_U3086), .C2(n8509), .ZN(P1_U3336) );
  NAND2_X1 U9297 ( .A1(n8914), .A2(P2_U3893), .ZN(n7514) );
  OAI21_X1 U9298 ( .B1(P2_U3893), .B2(n5301), .A(n7514), .ZN(P2_U3518) );
  XNOR2_X1 U9299 ( .A(n7515), .B(n7516), .ZN(n7517) );
  NAND2_X1 U9300 ( .A1(n7517), .A2(n7518), .ZN(n9376) );
  OAI21_X1 U9301 ( .B1(n7518), .B2(n7517), .A(n9376), .ZN(n7519) );
  NAND2_X1 U9302 ( .A1(n7519), .A2(n9948), .ZN(n7524) );
  OAI22_X1 U9303 ( .A1(n7521), .A2(n9221), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n7520), .ZN(n7522) );
  AOI21_X1 U9304 ( .B1(n10031), .B2(n9395), .A(n7522), .ZN(n7523) );
  OAI211_X1 U9305 ( .C1(n9920), .C2(n7525), .A(n7524), .B(n7523), .ZN(P1_U3227) );
  INV_X1 U9306 ( .A(n7526), .ZN(n7555) );
  INV_X1 U9307 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n7527) );
  OAI222_X1 U9308 ( .A1(n9905), .A2(n7555), .B1(n7528), .B2(P1_U3086), .C1(
        n7527), .C2(n9903), .ZN(P1_U3335) );
  INV_X1 U9309 ( .A(P2_REG2_REG_31__SCAN_IN), .ZN(n8885) );
  INV_X1 U9310 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n7529) );
  OR2_X1 U9311 ( .A1(n7530), .A2(n7529), .ZN(n7534) );
  INV_X1 U9312 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n7531) );
  OR2_X1 U9313 ( .A1(n7532), .A2(n7531), .ZN(n7533) );
  OAI211_X1 U9314 ( .C1(n7535), .C2(n8885), .A(n7534), .B(n7533), .ZN(n7536)
         );
  INV_X1 U9315 ( .A(n7536), .ZN(n7537) );
  NAND2_X1 U9316 ( .A1(n8882), .A2(P2_U3893), .ZN(n7539) );
  OAI21_X1 U9317 ( .B1(P2_U3893), .B2(n6486), .A(n7539), .ZN(P2_U3522) );
  INV_X1 U9318 ( .A(n7645), .ZN(n7553) );
  NAND2_X1 U9319 ( .A1(n7541), .A2(n7540), .ZN(n7542) );
  NAND2_X1 U9320 ( .A1(n7543), .A2(n7542), .ZN(n7591) );
  XNOR2_X1 U9321 ( .A(n7630), .B(n8580), .ZN(n7544) );
  AND2_X1 U9322 ( .A1(n7544), .A2(n7621), .ZN(n7592) );
  INV_X1 U9323 ( .A(n7544), .ZN(n7545) );
  NAND2_X1 U9324 ( .A1(n7545), .A2(n8739), .ZN(n7593) );
  XNOR2_X1 U9325 ( .A(n7645), .B(n8580), .ZN(n7726) );
  XNOR2_X1 U9326 ( .A(n7726), .B(n8738), .ZN(n7547) );
  OAI211_X1 U9327 ( .C1(n7546), .C2(n7547), .A(n7729), .B(n8717), .ZN(n7552)
         );
  AOI21_X1 U9328 ( .B1(n8739), .B2(n8720), .A(n7548), .ZN(n7549) );
  OAI21_X1 U9329 ( .B1(n7845), .B2(n8707), .A(n7549), .ZN(n7550) );
  AOI21_X1 U9330 ( .B1(n7622), .B2(n8709), .A(n7550), .ZN(n7551) );
  OAI211_X1 U9331 ( .C1(n7553), .C2(n8728), .A(n7552), .B(n7551), .ZN(P2_U3171) );
  OAI222_X1 U9332 ( .A1(P2_U3151), .A2(n8206), .B1(n9171), .B2(n7555), .C1(
        n7554), .C2(n8539), .ZN(P2_U3275) );
  OAI21_X1 U9333 ( .B1(n7558), .B2(n7556), .A(n7557), .ZN(n7559) );
  NAND2_X1 U9334 ( .A1(n7559), .A2(n9948), .ZN(n7567) );
  OR2_X1 U9335 ( .A1(n7717), .A2(n9338), .ZN(n7561) );
  NAND2_X1 U9336 ( .A1(n9419), .A2(n9199), .ZN(n7560) );
  NAND2_X1 U9337 ( .A1(n7561), .A2(n7560), .ZN(n9968) );
  INV_X1 U9338 ( .A(n9968), .ZN(n7563) );
  OAI21_X1 U9339 ( .B1(n7563), .B2(n9221), .A(n7562), .ZN(n7564) );
  AOI21_X1 U9340 ( .B1(n7565), .B2(n9395), .A(n7564), .ZN(n7566) );
  OAI211_X1 U9341 ( .C1(n9920), .C2(n9969), .A(n7567), .B(n7566), .ZN(P1_U3213) );
  XOR2_X1 U9342 ( .A(n7680), .B(n7581), .Z(n7569) );
  AOI21_X1 U9343 ( .B1(n5497), .B2(n7569), .A(n7681), .ZN(n7586) );
  INV_X1 U9344 ( .A(n7570), .ZN(n7571) );
  NOR2_X1 U9345 ( .A1(n7572), .A2(n7571), .ZN(n7574) );
  MUX2_X1 U9346 ( .A(P2_REG2_REG_11__SCAN_IN), .B(P2_REG1_REG_11__SCAN_IN), 
        .S(n8860), .Z(n7684) );
  XNOR2_X1 U9347 ( .A(n7684), .B(n7581), .ZN(n7573) );
  NOR2_X1 U9348 ( .A1(n7574), .A2(n7573), .ZN(n7685) );
  AOI21_X1 U9349 ( .B1(n7574), .B2(n7573), .A(n7685), .ZN(n7575) );
  NOR2_X1 U9350 ( .A1(n7575), .A2(n10129), .ZN(n7584) );
  INV_X1 U9351 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n10411) );
  NOR2_X1 U9352 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10411), .ZN(n7847) );
  INV_X1 U9353 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n7795) );
  AOI21_X1 U9354 ( .B1(n7795), .B2(n7578), .A(n7693), .ZN(n7579) );
  NOR2_X1 U9355 ( .A1(n7579), .A2(n10131), .ZN(n7583) );
  INV_X1 U9356 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n7580) );
  OAI22_X1 U9357 ( .A1(n10136), .A2(n7581), .B1(n8870), .B2(n7580), .ZN(n7582)
         );
  NOR4_X1 U9358 ( .A1(n7584), .A2(n7847), .A3(n7583), .A4(n7582), .ZN(n7585)
         );
  OAI21_X1 U9359 ( .B1(n7586), .B2(n10127), .A(n7585), .ZN(P2_U3193) );
  INV_X1 U9360 ( .A(n7631), .ZN(n7587) );
  NAND2_X1 U9361 ( .A1(n8709), .A2(n7587), .ZN(n7590) );
  AOI21_X1 U9362 ( .B1(n8720), .B2(n8740), .A(n7588), .ZN(n7589) );
  OAI211_X1 U9363 ( .C1(n7730), .C2(n8707), .A(n7590), .B(n7589), .ZN(n7598)
         );
  INV_X1 U9364 ( .A(n7592), .ZN(n7594) );
  NAND2_X1 U9365 ( .A1(n7594), .A2(n7593), .ZN(n7595) );
  XNOR2_X1 U9366 ( .A(n7591), .B(n7595), .ZN(n7596) );
  NOR2_X1 U9367 ( .A1(n7596), .A2(n8658), .ZN(n7597) );
  AOI211_X1 U9368 ( .C1(n7630), .C2(n8655), .A(n7598), .B(n7597), .ZN(n7599)
         );
  INV_X1 U9369 ( .A(n7599), .ZN(P2_U3161) );
  INV_X1 U9370 ( .A(n7600), .ZN(n7617) );
  OAI222_X1 U9371 ( .A1(n9905), .A2(n7617), .B1(n7601), .B2(P1_U3086), .C1(
        n10389), .C2(n9903), .ZN(P1_U3334) );
  NAND2_X1 U9372 ( .A1(P1_REG2_REG_14__SCAN_IN), .A2(n7887), .ZN(n7603) );
  OAI21_X1 U9373 ( .B1(P1_REG2_REG_14__SCAN_IN), .B2(n7887), .A(n7603), .ZN(
        n7604) );
  NOR2_X1 U9374 ( .A1(n7605), .A2(n7604), .ZN(n7886) );
  AOI211_X1 U9375 ( .C1(n7605), .C2(n7604), .A(n7886), .B(n7891), .ZN(n7615)
         );
  AOI21_X1 U9376 ( .B1(n7607), .B2(P1_REG1_REG_13__SCAN_IN), .A(n7606), .ZN(
        n7610) );
  MUX2_X1 U9377 ( .A(n7608), .B(P1_REG1_REG_14__SCAN_IN), .S(n7887), .Z(n7609)
         );
  NOR2_X1 U9378 ( .A1(n7610), .A2(n7609), .ZN(n7878) );
  AOI211_X1 U9379 ( .C1(n7610), .C2(n7609), .A(n7878), .B(n9510), .ZN(n7614)
         );
  INV_X1 U9380 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n7612) );
  NAND2_X1 U9381 ( .A1(n9516), .A2(n7887), .ZN(n7611) );
  NAND2_X1 U9382 ( .A1(P1_U3086), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n9180) );
  OAI211_X1 U9383 ( .C1(n7612), .C2(n9507), .A(n7611), .B(n9180), .ZN(n7613)
         );
  OR3_X1 U9384 ( .A1(n7615), .A2(n7614), .A3(n7613), .ZN(P1_U3257) );
  OAI222_X1 U9385 ( .A1(P2_U3151), .A2(n5818), .B1(n9171), .B2(n7617), .C1(
        n7616), .C2(n8539), .ZN(P2_U3274) );
  XOR2_X1 U9386 ( .A(n8232), .B(n7618), .Z(n7641) );
  INV_X1 U9387 ( .A(n7641), .ZN(n7628) );
  XNOR2_X1 U9388 ( .A(n7619), .B(n8232), .ZN(n7620) );
  OAI222_X1 U9389 ( .A1(n9006), .A2(n7621), .B1(n9008), .B2(n7845), .C1(n7620), 
        .C2(n9003), .ZN(n7640) );
  NAND2_X1 U9390 ( .A1(n7640), .A2(n9029), .ZN(n7627) );
  INV_X1 U9391 ( .A(n7622), .ZN(n7623) );
  OAI22_X1 U9392 ( .A1(n9029), .A2(n7624), .B1(n7623), .B2(n10141), .ZN(n7625)
         );
  AOI21_X1 U9393 ( .B1(n7645), .B2(n9032), .A(n7625), .ZN(n7626) );
  OAI211_X1 U9394 ( .C1(n9035), .C2(n7628), .A(n7627), .B(n7626), .ZN(P2_U3224) );
  XOR2_X1 U9395 ( .A(n8228), .B(n7629), .Z(n10191) );
  INV_X1 U9396 ( .A(n7630), .ZN(n10188) );
  OAI22_X1 U9397 ( .A1(n10188), .A2(n9014), .B1(n7631), .B2(n10141), .ZN(n7638) );
  NAND2_X1 U9398 ( .A1(n7632), .A2(n8228), .ZN(n7633) );
  NAND3_X1 U9399 ( .A1(n7634), .A2(n10151), .A3(n7633), .ZN(n7636) );
  AOI22_X1 U9400 ( .A1(n10148), .A2(n8738), .B1(n8740), .B2(n9025), .ZN(n7635)
         );
  NAND2_X1 U9401 ( .A1(n7636), .A2(n7635), .ZN(n10189) );
  MUX2_X1 U9402 ( .A(n10189), .B(P2_REG2_REG_8__SCAN_IN), .S(n10159), .Z(n7637) );
  AOI211_X1 U9403 ( .C1(n8021), .C2(n10191), .A(n7638), .B(n7637), .ZN(n7639)
         );
  INV_X1 U9404 ( .A(n7639), .ZN(P2_U3225) );
  AOI21_X1 U9405 ( .B1(n7641), .B2(n10192), .A(n7640), .ZN(n7647) );
  INV_X1 U9406 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n7642) );
  NOR2_X1 U9407 ( .A1(n10199), .A2(n7642), .ZN(n7643) );
  AOI21_X1 U9408 ( .B1(n7645), .B2(n9152), .A(n7643), .ZN(n7644) );
  OAI21_X1 U9409 ( .B1(n7647), .B2(n10201), .A(n7644), .ZN(P2_U3417) );
  AOI22_X1 U9410 ( .A1(n7645), .A2(n6647), .B1(n10211), .B2(
        P2_REG1_REG_9__SCAN_IN), .ZN(n7646) );
  OAI21_X1 U9411 ( .B1(n7647), .B2(n10211), .A(n7646), .ZN(P2_U3468) );
  OAI21_X1 U9412 ( .B1(n4589), .B2(n8464), .A(n7739), .ZN(n7650) );
  OR2_X1 U9413 ( .A1(n7669), .A2(n9537), .ZN(n7649) );
  OR2_X1 U9414 ( .A1(n7807), .A2(n9338), .ZN(n7648) );
  NAND2_X1 U9415 ( .A1(n7649), .A2(n7648), .ZN(n9914) );
  AOI21_X1 U9416 ( .B1(n7650), .B2(n9837), .A(n9914), .ZN(n10066) );
  OAI22_X1 U9417 ( .A1(n9742), .A2(n7651), .B1(n9921), .B2(n9970), .ZN(n7654)
         );
  INV_X1 U9418 ( .A(n7652), .ZN(n7747) );
  OAI211_X1 U9419 ( .C1(n10068), .C2(n7711), .A(n7747), .B(n9993), .ZN(n10065)
         );
  NOR2_X1 U9420 ( .A1(n10065), .A2(n9612), .ZN(n7653) );
  AOI211_X1 U9421 ( .C1(n9633), .C2(n7655), .A(n7654), .B(n7653), .ZN(n7659)
         );
  XNOR2_X1 U9422 ( .A(n7656), .B(n7657), .ZN(n10071) );
  NAND2_X1 U9423 ( .A1(n10071), .A2(n9929), .ZN(n7658) );
  OAI211_X1 U9424 ( .C1(n10000), .C2(n10066), .A(n7659), .B(n7658), .ZN(
        P1_U3283) );
  XOR2_X1 U9425 ( .A(n7663), .B(n7660), .Z(n10050) );
  NAND2_X1 U9426 ( .A1(n9964), .A2(n9963), .ZN(n7661) );
  NAND2_X1 U9427 ( .A1(n7661), .A2(n8349), .ZN(n9966) );
  INV_X1 U9428 ( .A(n8350), .ZN(n7662) );
  NAND2_X1 U9429 ( .A1(n9966), .A2(n7662), .ZN(n7714) );
  INV_X1 U9430 ( .A(n7714), .ZN(n7667) );
  INV_X1 U9431 ( .A(n7663), .ZN(n7664) );
  AOI21_X1 U9432 ( .B1(n9966), .B2(n7665), .A(n7664), .ZN(n7666) );
  AOI211_X1 U9433 ( .C1(n7667), .C2(n8354), .A(n9982), .B(n7666), .ZN(n7672)
         );
  OR2_X1 U9434 ( .A1(n7668), .A2(n9537), .ZN(n7671) );
  OR2_X1 U9435 ( .A1(n7669), .A2(n9338), .ZN(n7670) );
  NAND2_X1 U9436 ( .A1(n7671), .A2(n7670), .ZN(n9944) );
  NOR2_X1 U9437 ( .A1(n7672), .A2(n9944), .ZN(n10052) );
  INV_X1 U9438 ( .A(n10052), .ZN(n7678) );
  AOI21_X1 U9439 ( .B1(n9975), .B2(n9941), .A(n9831), .ZN(n7673) );
  NAND2_X1 U9440 ( .A1(n7673), .A2(n7709), .ZN(n10051) );
  NAND2_X1 U9441 ( .A1(n9988), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n7674) );
  OAI21_X1 U9442 ( .B1(n9970), .B2(n9952), .A(n7674), .ZN(n7675) );
  AOI21_X1 U9443 ( .B1(n9633), .B2(n9941), .A(n7675), .ZN(n7676) );
  OAI21_X1 U9444 ( .B1(n10051), .B2(n9612), .A(n7676), .ZN(n7677) );
  AOI21_X1 U9445 ( .B1(n7678), .B2(n9742), .A(n7677), .ZN(n7679) );
  OAI21_X1 U9446 ( .B1(n9726), .B2(n10050), .A(n7679), .ZN(P1_U3285) );
  NOR2_X1 U9447 ( .A1(n7692), .A2(n7680), .ZN(n7682) );
  AOI22_X1 U9448 ( .A1(P2_REG1_REG_12__SCAN_IN), .A2(n7699), .B1(n8759), .B2(
        n7687), .ZN(n7683) );
  AOI21_X1 U9449 ( .B1(n4592), .B2(n7683), .A(n8758), .ZN(n7708) );
  INV_X1 U9450 ( .A(n7684), .ZN(n7686) );
  AOI21_X1 U9451 ( .B1(n7692), .B2(n7686), .A(n7685), .ZN(n8751) );
  INV_X1 U9452 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n7862) );
  MUX2_X1 U9453 ( .A(n7862), .B(n7687), .S(n8860), .Z(n7688) );
  NOR2_X1 U9454 ( .A1(n7688), .A2(n7699), .ZN(n8750) );
  INV_X1 U9455 ( .A(n8750), .ZN(n7689) );
  NAND2_X1 U9456 ( .A1(n7688), .A2(n7699), .ZN(n8749) );
  NAND2_X1 U9457 ( .A1(n7689), .A2(n8749), .ZN(n7690) );
  XNOR2_X1 U9458 ( .A(n8751), .B(n7690), .ZN(n7706) );
  NOR2_X1 U9459 ( .A1(n7692), .A2(n7691), .ZN(n7694) );
  MUX2_X1 U9460 ( .A(n7862), .B(P2_REG2_REG_12__SCAN_IN), .S(n7699), .Z(n7695)
         );
  INV_X1 U9461 ( .A(n7695), .ZN(n7696) );
  AOI21_X1 U9462 ( .B1(n7697), .B2(n7696), .A(n8744), .ZN(n7698) );
  NOR2_X1 U9463 ( .A1(n7698), .A2(n10131), .ZN(n7705) );
  INV_X1 U9464 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n7703) );
  NAND2_X1 U9465 ( .A1(n8872), .A2(n7699), .ZN(n7702) );
  NOR2_X1 U9466 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7700), .ZN(n7936) );
  INV_X1 U9467 ( .A(n7936), .ZN(n7701) );
  OAI211_X1 U9468 ( .C1(n7703), .C2(n8870), .A(n7702), .B(n7701), .ZN(n7704)
         );
  AOI211_X1 U9469 ( .C1(n7706), .C2(n8814), .A(n7705), .B(n7704), .ZN(n7707)
         );
  OAI21_X1 U9470 ( .B1(n7708), .B2(n10127), .A(n7707), .ZN(P2_U3194) );
  NAND2_X1 U9471 ( .A1(n7709), .A2(n9306), .ZN(n7710) );
  NAND2_X1 U9472 ( .A1(n7710), .A2(n9993), .ZN(n7712) );
  OR2_X1 U9473 ( .A1(n7712), .A2(n7711), .ZN(n7713) );
  OR2_X1 U9474 ( .A1(n7740), .A2(n9338), .ZN(n9302) );
  NAND2_X1 U9475 ( .A1(n7713), .A2(n9302), .ZN(n10058) );
  NAND2_X1 U9476 ( .A1(n7714), .A2(n8354), .ZN(n7715) );
  XNOR2_X1 U9477 ( .A(n7715), .B(n7719), .ZN(n7716) );
  NAND2_X1 U9478 ( .A1(n7716), .A2(n9837), .ZN(n7718) );
  OR2_X1 U9479 ( .A1(n7717), .A2(n9537), .ZN(n9303) );
  NAND2_X1 U9480 ( .A1(n7718), .A2(n9303), .ZN(n10063) );
  AOI21_X1 U9481 ( .B1(n8509), .B2(n10058), .A(n10063), .ZN(n7725) );
  XNOR2_X1 U9482 ( .A(n7720), .B(n7719), .ZN(n10057) );
  NOR2_X1 U9483 ( .A1(n10060), .A2(n9990), .ZN(n7723) );
  OAI22_X1 U9484 ( .A1(n9742), .A2(n7721), .B1(n9307), .B2(n9970), .ZN(n7722)
         );
  AOI211_X1 U9485 ( .C1(n10057), .C2(n9929), .A(n7723), .B(n7722), .ZN(n7724)
         );
  OAI21_X1 U9486 ( .B1(n7725), .B2(n9988), .A(n7724), .ZN(P1_U3284) );
  INV_X1 U9487 ( .A(n7726), .ZN(n7727) );
  NAND2_X1 U9488 ( .A1(n7727), .A2(n8738), .ZN(n7728) );
  XNOR2_X1 U9489 ( .A(n7785), .B(n8580), .ZN(n7850) );
  XOR2_X1 U9490 ( .A(n7851), .B(n7850), .Z(n7736) );
  NOR2_X1 U9491 ( .A1(n7730), .A2(n8677), .ZN(n7731) );
  AOI211_X1 U9492 ( .C1(n8725), .C2(n8736), .A(n7732), .B(n7731), .ZN(n7733)
         );
  OAI21_X1 U9493 ( .B1(n7775), .B2(n8722), .A(n7733), .ZN(n7734) );
  AOI21_X1 U9494 ( .B1(n7777), .B2(n8655), .A(n7734), .ZN(n7735) );
  OAI21_X1 U9495 ( .B1(n7736), .B2(n8658), .A(n7735), .ZN(P2_U3157) );
  AOI21_X1 U9496 ( .B1(n7751), .B2(n7737), .A(n9982), .ZN(n7738) );
  OAI211_X1 U9497 ( .C1(n8471), .C2(n7739), .A(n7805), .B(n7738), .ZN(n7744)
         );
  OR2_X1 U9498 ( .A1(n7824), .A2(n9338), .ZN(n7742) );
  OR2_X1 U9499 ( .A1(n7740), .A2(n9537), .ZN(n7741) );
  NAND2_X1 U9500 ( .A1(n7742), .A2(n7741), .ZN(n9355) );
  INV_X1 U9501 ( .A(n9355), .ZN(n7743) );
  NAND2_X1 U9502 ( .A1(n7744), .A2(n7743), .ZN(n7763) );
  INV_X1 U9503 ( .A(n7763), .ZN(n7755) );
  INV_X1 U9504 ( .A(n7745), .ZN(n7746) );
  AOI211_X1 U9505 ( .C1(n7765), .C2(n7747), .A(n9831), .B(n7746), .ZN(n7762)
         );
  NOR2_X1 U9506 ( .A1(n9358), .A2(n9990), .ZN(n7750) );
  OAI22_X1 U9507 ( .A1(n9742), .A2(n7748), .B1(n9352), .B2(n9970), .ZN(n7749)
         );
  AOI211_X1 U9508 ( .C1(n7762), .C2(n9996), .A(n7750), .B(n7749), .ZN(n7754)
         );
  XNOR2_X1 U9509 ( .A(n7752), .B(n7751), .ZN(n7764) );
  NAND2_X1 U9510 ( .A1(n7764), .A2(n9929), .ZN(n7753) );
  OAI211_X1 U9511 ( .C1(n10000), .C2(n7755), .A(n7754), .B(n7753), .ZN(
        P1_U3282) );
  INV_X1 U9512 ( .A(n7756), .ZN(n7760) );
  OAI222_X1 U9513 ( .A1(n7758), .A2(P2_U3151), .B1(n9171), .B2(n7760), .C1(
        n7757), .C2(n8539), .ZN(P2_U3273) );
  OAI222_X1 U9514 ( .A1(n9903), .A2(n7761), .B1(n9905), .B2(n7760), .C1(
        P1_U3086), .C2(n7759), .ZN(P1_U3333) );
  AOI211_X1 U9515 ( .C1(n7764), .C2(n10070), .A(n7763), .B(n7762), .ZN(n7770)
         );
  INV_X1 U9516 ( .A(n9846), .ZN(n7872) );
  AOI22_X1 U9517 ( .A1(n7765), .A2(n7872), .B1(n10100), .B2(
        P1_REG1_REG_11__SCAN_IN), .ZN(n7766) );
  OAI21_X1 U9518 ( .B1(n7770), .B2(n10100), .A(n7766), .ZN(P1_U3533) );
  INV_X1 U9519 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n7767) );
  OAI22_X1 U9520 ( .A1(n9358), .A2(n9891), .B1(n10084), .B2(n7767), .ZN(n7768)
         );
  INV_X1 U9521 ( .A(n7768), .ZN(n7769) );
  OAI21_X1 U9522 ( .B1(n7770), .B2(n10082), .A(n7769), .ZN(P1_U3486) );
  XNOR2_X1 U9523 ( .A(n7777), .B(n8737), .ZN(n8233) );
  XNOR2_X1 U9524 ( .A(n7771), .B(n8233), .ZN(n7781) );
  XNOR2_X1 U9525 ( .A(n7772), .B(n8233), .ZN(n7773) );
  AOI222_X1 U9526 ( .A1(n10151), .A2(n7773), .B1(n8736), .B2(n10148), .C1(
        n8738), .C2(n9025), .ZN(n7780) );
  MUX2_X1 U9527 ( .A(n7774), .B(n7780), .S(n9029), .Z(n7779) );
  INV_X1 U9528 ( .A(n7775), .ZN(n7776) );
  AOI22_X1 U9529 ( .A1(n7777), .A2(n9032), .B1(n9031), .B2(n7776), .ZN(n7778)
         );
  OAI211_X1 U9530 ( .C1(n9035), .C2(n7781), .A(n7779), .B(n7778), .ZN(P2_U3223) );
  INV_X1 U9531 ( .A(n10192), .ZN(n10193) );
  OAI21_X1 U9532 ( .B1(n10193), .B2(n7781), .A(n7780), .ZN(n7787) );
  INV_X1 U9533 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n7782) );
  OAI22_X1 U9534 ( .A1(n7785), .A2(n9148), .B1(n7782), .B2(n10199), .ZN(n7783)
         );
  AOI21_X1 U9535 ( .B1(n7787), .B2(n10199), .A(n7783), .ZN(n7784) );
  INV_X1 U9536 ( .A(n7784), .ZN(P2_U3420) );
  OAI22_X1 U9537 ( .A1(n7785), .A2(n9076), .B1(n10213), .B2(n7370), .ZN(n7786)
         );
  AOI21_X1 U9538 ( .B1(n7787), .B2(n10213), .A(n7786), .ZN(n7788) );
  INV_X1 U9539 ( .A(n7788), .ZN(P2_U3469) );
  INV_X1 U9540 ( .A(n7790), .ZN(n8103) );
  NAND2_X1 U9541 ( .A1(n7789), .A2(n8103), .ZN(n7791) );
  XNOR2_X1 U9542 ( .A(n7791), .B(n8236), .ZN(n10194) );
  XOR2_X1 U9543 ( .A(n8236), .B(n7792), .Z(n7793) );
  OAI222_X1 U9544 ( .A1(n9008), .A2(n7959), .B1(n9006), .B2(n7845), .C1(n7793), 
        .C2(n9003), .ZN(n10195) );
  NAND2_X1 U9545 ( .A1(n10195), .A2(n9029), .ZN(n7798) );
  INV_X1 U9546 ( .A(n7794), .ZN(n7849) );
  OAI22_X1 U9547 ( .A1(n9029), .A2(n7795), .B1(n7849), .B2(n10141), .ZN(n7796)
         );
  AOI21_X1 U9548 ( .B1(n10197), .B2(n9032), .A(n7796), .ZN(n7797) );
  OAI211_X1 U9549 ( .C1(n10194), .C2(n9035), .A(n7798), .B(n7797), .ZN(
        P2_U3222) );
  NAND2_X1 U9550 ( .A1(n7802), .A2(n9166), .ZN(n7799) );
  OAI211_X1 U9551 ( .C1(n7800), .C2(n8539), .A(n7799), .B(n8271), .ZN(P2_U3272) );
  NAND2_X1 U9552 ( .A1(n7802), .A2(n7801), .ZN(n7804) );
  NAND2_X1 U9553 ( .A1(n7803), .A2(P1_STATE_REG_SCAN_IN), .ZN(n8518) );
  OAI211_X1 U9554 ( .C1(n5280), .C2(n9903), .A(n7804), .B(n8518), .ZN(P1_U3332) );
  NAND2_X1 U9555 ( .A1(n7805), .A2(n8369), .ZN(n7806) );
  XOR2_X1 U9556 ( .A(n8468), .B(n7806), .Z(n7811) );
  OR2_X1 U9557 ( .A1(n9177), .A2(n9338), .ZN(n7809) );
  OR2_X1 U9558 ( .A1(n7807), .A2(n9537), .ZN(n7808) );
  NAND2_X1 U9559 ( .A1(n7809), .A2(n7808), .ZN(n9248) );
  INV_X1 U9560 ( .A(n9248), .ZN(n7810) );
  OAI21_X1 U9561 ( .B1(n7811), .B2(n9982), .A(n7810), .ZN(n7836) );
  INV_X1 U9562 ( .A(n7836), .ZN(n7819) );
  XOR2_X1 U9563 ( .A(n8468), .B(n7812), .Z(n7838) );
  NAND2_X1 U9564 ( .A1(n7838), .A2(n9929), .ZN(n7818) );
  INV_X1 U9565 ( .A(n7828), .ZN(n7813) );
  AOI211_X1 U9566 ( .C1(n7842), .C2(n7745), .A(n9831), .B(n7813), .ZN(n7837)
         );
  INV_X1 U9567 ( .A(n7842), .ZN(n9251) );
  NOR2_X1 U9568 ( .A1(n9251), .A2(n9990), .ZN(n7816) );
  OAI22_X1 U9569 ( .A1(n9742), .A2(n7814), .B1(n9245), .B2(n9970), .ZN(n7815)
         );
  AOI211_X1 U9570 ( .C1(n7837), .C2(n9996), .A(n7816), .B(n7815), .ZN(n7817)
         );
  OAI211_X1 U9571 ( .C1(n10000), .C2(n7819), .A(n7818), .B(n7817), .ZN(
        P1_U3281) );
  INV_X1 U9572 ( .A(n7820), .ZN(n7821) );
  AOI211_X1 U9573 ( .C1(n7823), .C2(n7822), .A(n9982), .B(n7821), .ZN(n7827)
         );
  OR2_X1 U9574 ( .A1(n7824), .A2(n9537), .ZN(n7826) );
  OR2_X1 U9575 ( .A1(n7927), .A2(n9338), .ZN(n7825) );
  NAND2_X1 U9576 ( .A1(n7826), .A2(n7825), .ZN(n9330) );
  OR2_X1 U9577 ( .A1(n7827), .A2(n9330), .ZN(n7869) );
  INV_X1 U9578 ( .A(n7869), .ZN(n7835) );
  AOI211_X1 U9579 ( .C1(n7873), .C2(n7828), .A(n9831), .B(n9753), .ZN(n7870)
         );
  NOR2_X1 U9580 ( .A1(n4762), .A2(n9990), .ZN(n7831) );
  OAI22_X1 U9581 ( .A1(n9742), .A2(n7829), .B1(n9327), .B2(n9970), .ZN(n7830)
         );
  AOI211_X1 U9582 ( .C1(n7870), .C2(n9996), .A(n7831), .B(n7830), .ZN(n7834)
         );
  XNOR2_X1 U9583 ( .A(n7832), .B(n8470), .ZN(n7871) );
  NAND2_X1 U9584 ( .A1(n7871), .A2(n9929), .ZN(n7833) );
  OAI211_X1 U9585 ( .C1(n7835), .C2(n10000), .A(n7834), .B(n7833), .ZN(
        P1_U3280) );
  AOI211_X1 U9586 ( .C1(n7838), .C2(n10070), .A(n7837), .B(n7836), .ZN(n7844)
         );
  INV_X1 U9587 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n7839) );
  OAI22_X1 U9588 ( .A1(n9251), .A2(n9891), .B1(n10084), .B2(n7839), .ZN(n7840)
         );
  INV_X1 U9589 ( .A(n7840), .ZN(n7841) );
  OAI21_X1 U9590 ( .B1(n7844), .B2(n10082), .A(n7841), .ZN(P1_U3489) );
  AOI22_X1 U9591 ( .A1(n7842), .A2(n7872), .B1(n10100), .B2(
        P1_REG1_REG_12__SCAN_IN), .ZN(n7843) );
  OAI21_X1 U9592 ( .B1(n7844), .B2(n10100), .A(n7843), .ZN(P1_U3534) );
  NOR2_X1 U9593 ( .A1(n7845), .A2(n8677), .ZN(n7846) );
  AOI211_X1 U9594 ( .C1(n8725), .C2(n8735), .A(n7847), .B(n7846), .ZN(n7848)
         );
  OAI21_X1 U9595 ( .B1(n7849), .B2(n8722), .A(n7848), .ZN(n7854) );
  XNOR2_X1 U9596 ( .A(n8236), .B(n8580), .ZN(n7942) );
  AOI211_X1 U9597 ( .C1(n7942), .C2(n7852), .A(n8658), .B(n7941), .ZN(n7853)
         );
  AOI211_X1 U9598 ( .C1(n10197), .C2(n8655), .A(n7854), .B(n7853), .ZN(n7855)
         );
  INV_X1 U9599 ( .A(n7855), .ZN(P2_U3176) );
  XNOR2_X1 U9600 ( .A(n7856), .B(n8235), .ZN(n7868) );
  INV_X1 U9601 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n7859) );
  XNOR2_X1 U9602 ( .A(n7857), .B(n8235), .ZN(n7858) );
  AOI222_X1 U9603 ( .A1(n10151), .A2(n7858), .B1(n7981), .B2(n10148), .C1(
        n8736), .C2(n9025), .ZN(n7865) );
  MUX2_X1 U9604 ( .A(n7859), .B(n7865), .S(n10199), .Z(n7861) );
  NAND2_X1 U9605 ( .A1(n7947), .A2(n9152), .ZN(n7860) );
  OAI211_X1 U9606 ( .C1(n7868), .C2(n9156), .A(n7861), .B(n7860), .ZN(P2_U3426) );
  MUX2_X1 U9607 ( .A(n7862), .B(n7865), .S(n9029), .Z(n7864) );
  AOI22_X1 U9608 ( .A1(n7947), .A2(n9032), .B1(n9031), .B2(n7937), .ZN(n7863)
         );
  OAI211_X1 U9609 ( .C1(n7868), .C2(n9035), .A(n7864), .B(n7863), .ZN(P2_U3221) );
  NAND2_X1 U9610 ( .A1(n10213), .A2(n10192), .ZN(n9080) );
  MUX2_X1 U9611 ( .A(n7687), .B(n7865), .S(n10213), .Z(n7867) );
  NAND2_X1 U9612 ( .A1(n7947), .A2(n6647), .ZN(n7866) );
  OAI211_X1 U9613 ( .C1(n7868), .C2(n9080), .A(n7867), .B(n7866), .ZN(P2_U3471) );
  AOI211_X1 U9614 ( .C1(n7871), .C2(n10070), .A(n7870), .B(n7869), .ZN(n7877)
         );
  AOI22_X1 U9615 ( .A1(n7873), .A2(n7872), .B1(n10100), .B2(
        P1_REG1_REG_13__SCAN_IN), .ZN(n7874) );
  OAI21_X1 U9616 ( .B1(n7877), .B2(n10100), .A(n7874), .ZN(P1_U3535) );
  OAI22_X1 U9617 ( .A1(n4762), .A2(n9891), .B1(n10084), .B2(n6188), .ZN(n7875)
         );
  INV_X1 U9618 ( .A(n7875), .ZN(n7876) );
  OAI21_X1 U9619 ( .B1(n7877), .B2(n10082), .A(n7876), .ZN(P1_U3492) );
  AOI22_X1 U9620 ( .A1(n8528), .A2(P1_REG1_REG_16__SCAN_IN), .B1(n6254), .B2(
        n7884), .ZN(n7882) );
  NOR2_X1 U9621 ( .A1(n7879), .A2(n4737), .ZN(n7880) );
  NOR2_X1 U9622 ( .A1(n7880), .A2(n9485), .ZN(n7881) );
  NAND2_X1 U9623 ( .A1(n7882), .A2(n7881), .ZN(n8527) );
  OAI21_X1 U9624 ( .B1(n7882), .B2(n7881), .A(n8527), .ZN(n7896) );
  NAND2_X1 U9625 ( .A1(P1_U3086), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n9270) );
  NAND2_X1 U9626 ( .A1(n9956), .A2(P1_ADDR_REG_16__SCAN_IN), .ZN(n7883) );
  OAI211_X1 U9627 ( .C1(n7885), .C2(n7884), .A(n9270), .B(n7883), .ZN(n7895)
         );
  NOR2_X1 U9628 ( .A1(n7888), .A2(n4737), .ZN(n7889) );
  XOR2_X1 U9629 ( .A(n9483), .B(n7888), .Z(n9478) );
  NOR2_X1 U9630 ( .A1(n7921), .A2(n9478), .ZN(n9475) );
  NAND2_X1 U9631 ( .A1(n8528), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n7890) );
  OAI21_X1 U9632 ( .B1(n8528), .B2(P1_REG2_REG_16__SCAN_IN), .A(n7890), .ZN(
        n7892) );
  NOR2_X1 U9633 ( .A1(n7893), .A2(n7892), .ZN(n8521) );
  AOI211_X1 U9634 ( .C1(n7893), .C2(n7892), .A(n8521), .B(n7891), .ZN(n7894)
         );
  AOI211_X1 U9635 ( .C1(n9499), .C2(n7896), .A(n7895), .B(n7894), .ZN(n7897)
         );
  INV_X1 U9636 ( .A(n7897), .ZN(P1_U3259) );
  INV_X1 U9637 ( .A(n7898), .ZN(n7909) );
  OAI222_X1 U9638 ( .A1(n9905), .A2(n7909), .B1(P1_U3086), .B2(n7899), .C1(
        n10588), .C2(n9903), .ZN(P1_U3331) );
  OAI211_X1 U9639 ( .C1(n7900), .C2(n8238), .A(n7969), .B(n10151), .ZN(n7902)
         );
  AOI22_X1 U9640 ( .A1(n9025), .A2(n8735), .B1(n8734), .B2(n10148), .ZN(n7901)
         );
  AND2_X1 U9641 ( .A1(n7902), .A2(n7901), .ZN(n7914) );
  INV_X1 U9642 ( .A(n7914), .ZN(n7904) );
  INV_X1 U9643 ( .A(n7953), .ZN(n7964) );
  OAI22_X1 U9644 ( .A1(n7964), .A2(n10142), .B1(n7957), .B2(n10141), .ZN(n7903) );
  OAI21_X1 U9645 ( .B1(n7904), .B2(n7903), .A(n9029), .ZN(n7907) );
  XNOR2_X1 U9646 ( .A(n7905), .B(n8238), .ZN(n7915) );
  AOI22_X1 U9647 ( .A1(n7915), .A2(n8021), .B1(P2_REG2_REG_13__SCAN_IN), .B2(
        n10159), .ZN(n7906) );
  NAND2_X1 U9648 ( .A1(n7907), .A2(n7906), .ZN(P2_U3220) );
  OAI222_X1 U9649 ( .A1(n7910), .A2(P2_U3151), .B1(n9171), .B2(n7909), .C1(
        n7908), .C2(n8539), .ZN(P2_U3271) );
  MUX2_X1 U9650 ( .A(n7914), .B(n7911), .S(n10201), .Z(n7913) );
  INV_X1 U9651 ( .A(n9156), .ZN(n9096) );
  AOI22_X1 U9652 ( .A1(n7915), .A2(n9096), .B1(n9152), .B2(n7953), .ZN(n7912)
         );
  NAND2_X1 U9653 ( .A1(n7913), .A2(n7912), .ZN(P2_U3429) );
  MUX2_X1 U9654 ( .A(n7914), .B(n10110), .S(n10211), .Z(n7917) );
  INV_X1 U9655 ( .A(n9080), .ZN(n9043) );
  AOI22_X1 U9656 ( .A1(n7915), .A2(n9043), .B1(n6647), .B2(n7953), .ZN(n7916)
         );
  NAND2_X1 U9657 ( .A1(n7917), .A2(n7916), .ZN(P2_U3472) );
  INV_X1 U9658 ( .A(n7918), .ZN(n7934) );
  OAI222_X1 U9659 ( .A1(n9905), .A2(n7934), .B1(P1_U3086), .B2(n7919), .C1(
        n10526), .C2(n9903), .ZN(P1_U3330) );
  XNOR2_X1 U9660 ( .A(n7920), .B(n7926), .ZN(n9843) );
  OAI22_X1 U9661 ( .A1(n9742), .A2(n7921), .B1(n9393), .B2(n9970), .ZN(n7923)
         );
  OAI211_X1 U9662 ( .C1(n9754), .C2(n9892), .A(n9993), .B(n9832), .ZN(n9841)
         );
  NOR2_X1 U9663 ( .A1(n9841), .A2(n9612), .ZN(n7922) );
  AOI211_X1 U9664 ( .C1(n9633), .C2(n9396), .A(n7923), .B(n7922), .ZN(n7932)
         );
  OAI21_X1 U9665 ( .B1(n7926), .B2(n7925), .A(n7924), .ZN(n7930) );
  OR2_X1 U9666 ( .A1(n7927), .A2(n9537), .ZN(n7929) );
  OR2_X1 U9667 ( .A1(n9279), .A2(n9338), .ZN(n7928) );
  NAND2_X1 U9668 ( .A1(n7929), .A2(n7928), .ZN(n9391) );
  AOI21_X1 U9669 ( .B1(n7930), .B2(n9837), .A(n9391), .ZN(n9842) );
  OR2_X1 U9670 ( .A1(n9842), .A2(n10000), .ZN(n7931) );
  OAI211_X1 U9671 ( .C1(n9843), .C2(n9726), .A(n7932), .B(n7931), .ZN(P1_U3278) );
  OAI222_X1 U9672 ( .A1(n7935), .A2(P2_U3151), .B1(n9171), .B2(n7934), .C1(
        n7933), .C2(n8539), .ZN(P2_U3270) );
  AOI21_X1 U9673 ( .B1(n7981), .B2(n8725), .A(n7936), .ZN(n7939) );
  NAND2_X1 U9674 ( .A1(n8709), .A2(n7937), .ZN(n7938) );
  OAI211_X1 U9675 ( .C1(n7940), .C2(n8677), .A(n7939), .B(n7938), .ZN(n7946)
         );
  XNOR2_X1 U9676 ( .A(n7947), .B(n8580), .ZN(n7950) );
  XNOR2_X1 U9677 ( .A(n7950), .B(n7959), .ZN(n7943) );
  AOI211_X1 U9678 ( .C1(n7944), .C2(n7943), .A(n8658), .B(n7952), .ZN(n7945)
         );
  AOI211_X1 U9679 ( .C1(n7947), .C2(n8655), .A(n7946), .B(n7945), .ZN(n7948)
         );
  INV_X1 U9680 ( .A(n7948), .ZN(P2_U3164) );
  INV_X1 U9681 ( .A(n7949), .ZN(n7966) );
  INV_X1 U9682 ( .A(n7950), .ZN(n7951) );
  XNOR2_X1 U9683 ( .A(n7953), .B(n8580), .ZN(n7979) );
  XNOR2_X1 U9684 ( .A(n7979), .B(n7981), .ZN(n7954) );
  NAND2_X1 U9685 ( .A1(n7955), .A2(n7954), .ZN(n7980) );
  OAI21_X1 U9686 ( .B1(n7955), .B2(n7954), .A(n7980), .ZN(n7956) );
  NAND2_X1 U9687 ( .A1(n7956), .A2(n8717), .ZN(n7963) );
  INV_X1 U9688 ( .A(n7957), .ZN(n7961) );
  AOI22_X1 U9689 ( .A1(n8725), .A2(n8734), .B1(P2_REG3_REG_13__SCAN_IN), .B2(
        P2_U3151), .ZN(n7958) );
  OAI21_X1 U9690 ( .B1(n7959), .B2(n8677), .A(n7958), .ZN(n7960) );
  AOI21_X1 U9691 ( .B1(n7961), .B2(n8709), .A(n7960), .ZN(n7962) );
  OAI211_X1 U9692 ( .C1(n7964), .C2(n8728), .A(n7963), .B(n7962), .ZN(P2_U3174) );
  OAI222_X1 U9693 ( .A1(n7967), .A2(P2_U3151), .B1(n9171), .B2(n7966), .C1(
        n7965), .C2(n8539), .ZN(P2_U3269) );
  INV_X1 U9694 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n7973) );
  NAND2_X1 U9695 ( .A1(n7969), .A2(n7968), .ZN(n7971) );
  INV_X1 U9696 ( .A(n8130), .ZN(n7970) );
  XNOR2_X1 U9697 ( .A(n7971), .B(n8241), .ZN(n7972) );
  AOI222_X1 U9698 ( .A1(n10151), .A2(n7972), .B1(n7981), .B2(n9025), .C1(n8733), .C2(n10148), .ZN(n8017) );
  MUX2_X1 U9699 ( .A(n7973), .B(n8017), .S(n10199), .Z(n7976) );
  XNOR2_X1 U9700 ( .A(n7974), .B(n8241), .ZN(n8022) );
  AOI22_X1 U9701 ( .A1(n8022), .A2(n9096), .B1(n9152), .B2(n8015), .ZN(n7975)
         );
  NAND2_X1 U9702 ( .A1(n7976), .A2(n7975), .ZN(P2_U3432) );
  MUX2_X1 U9703 ( .A(n8763), .B(n8017), .S(n10213), .Z(n7978) );
  AOI22_X1 U9704 ( .A1(n8022), .A2(n9043), .B1(n6647), .B2(n8015), .ZN(n7977)
         );
  NAND2_X1 U9705 ( .A1(n7978), .A2(n7977), .ZN(P2_U3473) );
  INV_X1 U9706 ( .A(n7979), .ZN(n7982) );
  XNOR2_X1 U9707 ( .A(n8015), .B(n8580), .ZN(n8002) );
  XNOR2_X1 U9708 ( .A(n8002), .B(n8734), .ZN(n8004) );
  XOR2_X1 U9709 ( .A(n8005), .B(n8004), .Z(n7988) );
  NAND2_X1 U9710 ( .A1(n8709), .A2(n8020), .ZN(n7984) );
  AOI22_X1 U9711 ( .A1(n8725), .A2(n8733), .B1(P2_REG3_REG_14__SCAN_IN), .B2(
        P2_U3151), .ZN(n7983) );
  OAI211_X1 U9712 ( .C1(n7985), .C2(n8677), .A(n7984), .B(n7983), .ZN(n7986)
         );
  AOI21_X1 U9713 ( .B1(n8015), .B2(n8655), .A(n7986), .ZN(n7987) );
  OAI21_X1 U9714 ( .B1(n7988), .B2(n8658), .A(n7987), .ZN(P2_U3155) );
  XNOR2_X1 U9715 ( .A(n7989), .B(n8240), .ZN(n8001) );
  INV_X1 U9716 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n7992) );
  XNOR2_X1 U9717 ( .A(n7990), .B(n8240), .ZN(n7991) );
  AOI222_X1 U9718 ( .A1(n10151), .A2(n7991), .B1(n8734), .B2(n9025), .C1(n9026), .C2(n10148), .ZN(n7997) );
  MUX2_X1 U9719 ( .A(n7992), .B(n7997), .S(n10199), .Z(n7994) );
  NAND2_X1 U9720 ( .A1(n8006), .A2(n9152), .ZN(n7993) );
  OAI211_X1 U9721 ( .C1(n8001), .C2(n9156), .A(n7994), .B(n7993), .ZN(P2_U3435) );
  MUX2_X1 U9722 ( .A(n8767), .B(n7997), .S(n10213), .Z(n7996) );
  NAND2_X1 U9723 ( .A1(n8006), .A2(n6647), .ZN(n7995) );
  OAI211_X1 U9724 ( .C1(n9080), .C2(n8001), .A(n7996), .B(n7995), .ZN(P2_U3474) );
  INV_X1 U9725 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n7998) );
  MUX2_X1 U9726 ( .A(n7998), .B(n7997), .S(n9029), .Z(n8000) );
  AOI22_X1 U9727 ( .A1(n8006), .A2(n9032), .B1(n9031), .B2(n8011), .ZN(n7999)
         );
  OAI211_X1 U9728 ( .C1(n8001), .C2(n9035), .A(n8000), .B(n7999), .ZN(P2_U3218) );
  INV_X1 U9729 ( .A(n8006), .ZN(n8014) );
  AOI22_X2 U9730 ( .A1(n8005), .A2(n8004), .B1(n8003), .B2(n8002), .ZN(n8008)
         );
  XNOR2_X1 U9731 ( .A(n8006), .B(n8580), .ZN(n8543) );
  XNOR2_X1 U9732 ( .A(n8543), .B(n8733), .ZN(n8007) );
  OAI211_X1 U9733 ( .C1(n8008), .C2(n8007), .A(n8545), .B(n8717), .ZN(n8013)
         );
  NAND2_X1 U9734 ( .A1(n8720), .A2(n8734), .ZN(n8009) );
  NAND2_X1 U9735 ( .A1(P2_U3151), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n8755) );
  OAI211_X1 U9736 ( .C1(n8653), .C2(n8707), .A(n8009), .B(n8755), .ZN(n8010)
         );
  AOI21_X1 U9737 ( .B1(n8011), .B2(n8709), .A(n8010), .ZN(n8012) );
  OAI211_X1 U9738 ( .C1(n8014), .C2(n8728), .A(n8013), .B(n8012), .ZN(P2_U3181) );
  INV_X1 U9739 ( .A(n8015), .ZN(n8016) );
  NOR2_X1 U9740 ( .A1(n8016), .A2(n10142), .ZN(n8019) );
  INV_X1 U9741 ( .A(n8017), .ZN(n8018) );
  AOI211_X1 U9742 ( .C1(n9031), .C2(n8020), .A(n8019), .B(n8018), .ZN(n8024)
         );
  AOI22_X1 U9743 ( .A1(n8022), .A2(n8021), .B1(P2_REG2_REG_14__SCAN_IN), .B2(
        n10159), .ZN(n8023) );
  OAI21_X1 U9744 ( .B1(n8024), .B2(n10159), .A(n8023), .ZN(P2_U3219) );
  NAND2_X1 U9745 ( .A1(n8025), .A2(n8242), .ZN(n8026) );
  NAND3_X1 U9746 ( .A1(n9021), .A2(n10151), .A3(n8026), .ZN(n8028) );
  AOI22_X1 U9747 ( .A1(n8731), .A2(n10148), .B1(n9025), .B2(n8733), .ZN(n8027)
         );
  MUX2_X1 U9748 ( .A(n8038), .B(n8029), .S(n10201), .Z(n8033) );
  OAI21_X1 U9749 ( .B1(n8030), .B2(n8242), .A(n8031), .ZN(n8036) );
  AOI22_X1 U9750 ( .A1(n8036), .A2(n9096), .B1(n9152), .B2(n8647), .ZN(n8032)
         );
  NAND2_X1 U9751 ( .A1(n8033), .A2(n8032), .ZN(P2_U3438) );
  MUX2_X1 U9752 ( .A(n8777), .B(n8038), .S(n10213), .Z(n8035) );
  AOI22_X1 U9753 ( .A1(n8036), .A2(n9043), .B1(n6647), .B2(n8647), .ZN(n8034)
         );
  NAND2_X1 U9754 ( .A1(n8035), .A2(n8034), .ZN(P2_U3475) );
  INV_X1 U9755 ( .A(n8036), .ZN(n8042) );
  MUX2_X1 U9756 ( .A(n8038), .B(n8037), .S(n10159), .Z(n8041) );
  INV_X1 U9757 ( .A(n8645), .ZN(n8039) );
  AOI22_X1 U9758 ( .A1(n8647), .A2(n9032), .B1(n9031), .B2(n8039), .ZN(n8040)
         );
  OAI211_X1 U9759 ( .C1(n8042), .C2(n9035), .A(n8041), .B(n8040), .ZN(P2_U3217) );
  MUX2_X1 U9760 ( .A(n8902), .B(n8590), .S(n8174), .Z(n8193) );
  INV_X1 U9761 ( .A(n8043), .ZN(n8172) );
  MUX2_X1 U9762 ( .A(n8172), .B(n8173), .S(n8203), .Z(n8044) );
  NOR2_X1 U9763 ( .A1(n8044), .A2(n8897), .ZN(n8183) );
  INV_X1 U9764 ( .A(n8045), .ZN(n8048) );
  NAND2_X1 U9765 ( .A1(n8219), .A2(n8046), .ZN(n8047) );
  MUX2_X1 U9766 ( .A(n8048), .B(n8047), .S(n8203), .Z(n8162) );
  INV_X1 U9767 ( .A(n8049), .ZN(n8158) );
  NOR2_X1 U9768 ( .A1(n8158), .A2(n8050), .ZN(n8051) );
  MUX2_X1 U9769 ( .A(n8052), .B(n8051), .S(n8203), .Z(n8161) );
  NAND2_X1 U9770 ( .A1(n8138), .A2(n8053), .ZN(n8246) );
  NAND2_X1 U9771 ( .A1(n8246), .A2(n8203), .ZN(n8137) );
  MUX2_X1 U9772 ( .A(n8055), .B(n8054), .S(n8203), .Z(n8128) );
  INV_X1 U9773 ( .A(n8238), .ZN(n8126) );
  MUX2_X1 U9774 ( .A(n8057), .B(n8056), .S(n8174), .Z(n8125) );
  INV_X1 U9775 ( .A(n8119), .ZN(n8123) );
  NAND2_X1 U9776 ( .A1(n8058), .A2(n5818), .ZN(n8059) );
  NAND2_X1 U9777 ( .A1(n8059), .A2(n8062), .ZN(n8060) );
  NAND2_X1 U9778 ( .A1(n8060), .A2(n8066), .ZN(n8065) );
  AND2_X1 U9779 ( .A1(n8061), .A2(n8174), .ZN(n8064) );
  AOI21_X1 U9780 ( .B1(n8062), .B2(n8061), .A(n8174), .ZN(n8063) );
  AOI21_X1 U9781 ( .B1(n8065), .B2(n8064), .A(n8063), .ZN(n8074) );
  OAI21_X1 U9782 ( .B1(n8066), .B2(n8174), .A(n10139), .ZN(n8073) );
  NAND2_X1 U9783 ( .A1(n8743), .A2(n10143), .ZN(n8067) );
  NAND2_X1 U9784 ( .A1(n8076), .A2(n8067), .ZN(n8070) );
  NAND2_X1 U9785 ( .A1(n8084), .A2(n8068), .ZN(n8069) );
  MUX2_X1 U9786 ( .A(n8070), .B(n8069), .S(n8174), .Z(n8071) );
  INV_X1 U9787 ( .A(n8071), .ZN(n8072) );
  OAI21_X1 U9788 ( .B1(n8074), .B2(n8073), .A(n8072), .ZN(n8075) );
  NAND2_X1 U9789 ( .A1(n8075), .A2(n8220), .ZN(n8088) );
  INV_X1 U9790 ( .A(n8076), .ZN(n8079) );
  INV_X1 U9791 ( .A(n8089), .ZN(n8078) );
  OAI211_X1 U9792 ( .C1(n8088), .C2(n8079), .A(n8078), .B(n8077), .ZN(n8083)
         );
  INV_X1 U9793 ( .A(n8085), .ZN(n8080) );
  NOR2_X1 U9794 ( .A1(n8080), .A2(n8091), .ZN(n8082) );
  INV_X1 U9795 ( .A(n8081), .ZN(n8090) );
  AOI21_X1 U9796 ( .B1(n8083), .B2(n8082), .A(n8090), .ZN(n8095) );
  INV_X1 U9797 ( .A(n8084), .ZN(n8087) );
  NAND2_X1 U9798 ( .A1(n8742), .A2(n10170), .ZN(n8086) );
  OAI211_X1 U9799 ( .C1(n8088), .C2(n8087), .A(n8086), .B(n8085), .ZN(n8093)
         );
  NOR2_X1 U9800 ( .A1(n8090), .A2(n8089), .ZN(n8092) );
  AOI21_X1 U9801 ( .B1(n8093), .B2(n8092), .A(n8091), .ZN(n8094) );
  MUX2_X1 U9802 ( .A(n8095), .B(n8094), .S(n8203), .Z(n8099) );
  NAND2_X1 U9803 ( .A1(n8115), .A2(n8114), .ZN(n8104) );
  INV_X1 U9804 ( .A(n8104), .ZN(n8098) );
  NAND2_X1 U9805 ( .A1(n8102), .A2(n8101), .ZN(n8116) );
  NOR3_X1 U9806 ( .A1(n8106), .A2(n8116), .A3(n8096), .ZN(n8097) );
  NAND4_X1 U9807 ( .A1(n8099), .A2(n8098), .A3(n8097), .A4(n8108), .ZN(n8122)
         );
  AND2_X1 U9808 ( .A1(n8101), .A2(n8100), .ZN(n8105) );
  OAI211_X1 U9809 ( .C1(n8105), .C2(n8104), .A(n8103), .B(n8102), .ZN(n8107)
         );
  NAND4_X1 U9810 ( .A1(n8108), .A2(n8107), .A3(n8203), .A4(n5759), .ZN(n8112)
         );
  AND2_X1 U9811 ( .A1(n8736), .A2(n8174), .ZN(n8110) );
  OAI21_X1 U9812 ( .B1(n8174), .B2(n8736), .A(n10197), .ZN(n8109) );
  OAI21_X1 U9813 ( .B1(n8110), .B2(n10197), .A(n8109), .ZN(n8111) );
  AND3_X1 U9814 ( .A1(n8235), .A2(n8112), .A3(n8111), .ZN(n8121) );
  AND2_X1 U9815 ( .A1(n8114), .A2(n8113), .ZN(n8117) );
  OAI211_X1 U9816 ( .C1(n8117), .C2(n8116), .A(n5759), .B(n8115), .ZN(n8118)
         );
  NAND3_X1 U9817 ( .A1(n8119), .A2(n8174), .A3(n8118), .ZN(n8120) );
  OAI211_X1 U9818 ( .C1(n8123), .C2(n8122), .A(n8121), .B(n8120), .ZN(n8124)
         );
  NAND3_X1 U9819 ( .A1(n8126), .A2(n8125), .A3(n8124), .ZN(n8127) );
  NAND2_X1 U9820 ( .A1(n8128), .A2(n8127), .ZN(n8132) );
  MUX2_X1 U9821 ( .A(n8130), .B(n5116), .S(n8174), .Z(n8131) );
  OAI21_X1 U9822 ( .B1(n8133), .B2(n8132), .A(n8131), .ZN(n8134) );
  NAND2_X1 U9823 ( .A1(n8240), .A2(n8134), .ZN(n8142) );
  NAND3_X1 U9824 ( .A1(n8142), .A2(n8144), .A3(n8135), .ZN(n8136) );
  INV_X1 U9825 ( .A(n8138), .ZN(n8139) );
  MUX2_X1 U9826 ( .A(n8140), .B(n8139), .S(n8174), .Z(n8156) );
  NAND4_X1 U9827 ( .A1(n8146), .A2(n8143), .A3(n8142), .A4(n8141), .ZN(n8148)
         );
  NAND2_X1 U9828 ( .A1(n8144), .A2(n8174), .ZN(n8145) );
  NAND2_X1 U9829 ( .A1(n8146), .A2(n8145), .ZN(n8147) );
  NAND4_X1 U9830 ( .A1(n8148), .A2(n8147), .A3(n8243), .A4(n8245), .ZN(n8149)
         );
  NAND2_X1 U9831 ( .A1(n8149), .A2(n8151), .ZN(n8155) );
  NAND2_X1 U9832 ( .A1(n8979), .A2(n8150), .ZN(n8153) );
  NAND2_X1 U9833 ( .A1(n8965), .A2(n8151), .ZN(n8152) );
  MUX2_X1 U9834 ( .A(n8153), .B(n8152), .S(n8203), .Z(n8154) );
  INV_X1 U9835 ( .A(n8157), .ZN(n8159) );
  MUX2_X1 U9836 ( .A(n8159), .B(n8158), .S(n8174), .Z(n8160) );
  INV_X1 U9837 ( .A(n8930), .ZN(n8163) );
  INV_X1 U9838 ( .A(n8218), .ZN(n8164) );
  AOI21_X1 U9839 ( .B1(n8165), .B2(n8217), .A(n8164), .ZN(n8171) );
  INV_X1 U9840 ( .A(n8166), .ZN(n8169) );
  INV_X1 U9841 ( .A(n8167), .ZN(n8168) );
  OAI21_X1 U9842 ( .B1(n8169), .B2(n8168), .A(n8218), .ZN(n8170) );
  INV_X1 U9843 ( .A(n8922), .ZN(n8178) );
  INV_X1 U9844 ( .A(n8912), .ZN(n8910) );
  MUX2_X1 U9845 ( .A(n8176), .B(n8175), .S(n8174), .Z(n8177) );
  INV_X1 U9846 ( .A(n8179), .ZN(n8181) );
  INV_X1 U9847 ( .A(n9095), .ZN(n8603) );
  NOR2_X1 U9848 ( .A1(n8603), .A2(n8914), .ZN(n8180) );
  MUX2_X1 U9849 ( .A(n8181), .B(n8180), .S(n8203), .Z(n8182) );
  NAND2_X1 U9850 ( .A1(n8537), .A2(n8198), .ZN(n8187) );
  OR2_X1 U9851 ( .A1(n4507), .A2(n8185), .ZN(n8186) );
  INV_X1 U9852 ( .A(n8730), .ZN(n8189) );
  OR2_X1 U9853 ( .A1(n9084), .A2(n8189), .ZN(n8215) );
  OAI211_X1 U9854 ( .C1(n8188), .C2(n8590), .A(n8212), .B(n8215), .ZN(n8197)
         );
  INV_X1 U9855 ( .A(n8188), .ZN(n8192) );
  NAND2_X1 U9856 ( .A1(n9084), .A2(n8189), .ZN(n8253) );
  NAND2_X1 U9857 ( .A1(n8253), .A2(n8190), .ZN(n8214) );
  AOI21_X1 U9858 ( .B1(n8192), .B2(n8191), .A(n8214), .ZN(n8196) );
  INV_X1 U9859 ( .A(n8194), .ZN(n8195) );
  OAI22_X1 U9860 ( .A1(n8196), .A2(n8203), .B1(n4710), .B2(n8195), .ZN(n8210)
         );
  OAI21_X1 U9861 ( .B1(n8197), .B2(n8210), .A(n8253), .ZN(n8201) );
  NAND2_X1 U9862 ( .A1(n9895), .A2(n8198), .ZN(n8200) );
  OR2_X1 U9863 ( .A1(n4507), .A2(n9163), .ZN(n8199) );
  NAND2_X1 U9864 ( .A1(n9081), .A2(n8216), .ZN(n8202) );
  NAND3_X1 U9865 ( .A1(n8201), .A2(n8203), .A3(n8202), .ZN(n8264) );
  INV_X1 U9866 ( .A(n8202), .ZN(n8204) );
  INV_X1 U9867 ( .A(n8215), .ZN(n8255) );
  NOR3_X1 U9868 ( .A1(n8204), .A2(n8203), .A3(n8255), .ZN(n8209) );
  NOR2_X1 U9869 ( .A1(n8882), .A2(n8205), .ZN(n8207) );
  OAI22_X1 U9870 ( .A1(n9081), .A2(n8207), .B1(n8216), .B2(n8206), .ZN(n8208)
         );
  AOI21_X1 U9871 ( .B1(n8210), .B2(n8209), .A(n8208), .ZN(n8263) );
  INV_X1 U9872 ( .A(n8211), .ZN(n8213) );
  NOR2_X1 U9873 ( .A1(n9081), .A2(n8216), .ZN(n8257) );
  NAND2_X1 U9874 ( .A1(n8219), .A2(n8930), .ZN(n8943) );
  NAND4_X1 U9875 ( .A1(n8223), .A2(n8222), .A3(n8221), .A4(n8220), .ZN(n8224)
         );
  NOR2_X1 U9876 ( .A1(n8224), .A2(n10146), .ZN(n8230) );
  NOR2_X1 U9877 ( .A1(n8226), .A2(n8225), .ZN(n8227) );
  NAND4_X1 U9878 ( .A1(n8230), .A2(n8229), .A3(n8228), .A4(n8227), .ZN(n8231)
         );
  NOR2_X1 U9879 ( .A1(n8232), .A2(n8231), .ZN(n8234) );
  NAND3_X1 U9880 ( .A1(n8235), .A2(n8234), .A3(n8233), .ZN(n8237) );
  NOR3_X1 U9881 ( .A1(n8238), .A2(n8237), .A3(n8236), .ZN(n8239) );
  AND4_X1 U9882 ( .A1(n8242), .A2(n8241), .A3(n8240), .A4(n8239), .ZN(n8244)
         );
  NAND3_X1 U9883 ( .A1(n8245), .A2(n8244), .A3(n8243), .ZN(n8247) );
  NOR2_X1 U9884 ( .A1(n8247), .A2(n8246), .ZN(n8248) );
  NAND3_X1 U9885 ( .A1(n8979), .A2(n8989), .A3(n8248), .ZN(n8249) );
  NOR4_X1 U9886 ( .A1(n8943), .A2(n8953), .A3(n8968), .A4(n8249), .ZN(n8250)
         );
  NAND3_X1 U9887 ( .A1(n8922), .A2(n8934), .A3(n8250), .ZN(n8251) );
  NOR2_X1 U9888 ( .A1(n8912), .A2(n8251), .ZN(n8252) );
  NAND4_X1 U9889 ( .A1(n8253), .A2(n8252), .A3(n5766), .A4(n8581), .ZN(n8256)
         );
  NOR4_X1 U9890 ( .A1(n8257), .A2(n8256), .A3(n8255), .A4(n8254), .ZN(n8259)
         );
  OAI22_X1 U9891 ( .A1(n8261), .A2(n8260), .B1(n8259), .B2(n8258), .ZN(n8262)
         );
  AOI21_X1 U9892 ( .B1(n8264), .B2(n8263), .A(n8262), .ZN(n8265) );
  XNOR2_X1 U9893 ( .A(n8265), .B(n8873), .ZN(n8272) );
  NOR3_X1 U9894 ( .A1(n8267), .A2(n8266), .A3(n8276), .ZN(n8270) );
  OAI21_X1 U9895 ( .B1(n8271), .B2(n8268), .A(P2_B_REG_SCAN_IN), .ZN(n8269) );
  OAI22_X1 U9896 ( .A1(n8272), .A2(n8271), .B1(n8270), .B2(n8269), .ZN(
        P2_U3296) );
  INV_X1 U9897 ( .A(n8273), .ZN(n8541) );
  OAI222_X1 U9898 ( .A1(n4508), .A2(P1_U3086), .B1(n9905), .B2(n8541), .C1(
        n9903), .C2(n5301), .ZN(P1_U3328) );
  INV_X1 U9899 ( .A(n8274), .ZN(n9904) );
  OAI222_X1 U9900 ( .A1(P2_U3151), .A2(n8276), .B1(n9171), .B2(n9904), .C1(
        n8275), .C2(n8539), .ZN(P2_U3267) );
  INV_X1 U9901 ( .A(n8434), .ZN(n8277) );
  OR2_X1 U9902 ( .A1(n9591), .A2(n9257), .ZN(n8432) );
  INV_X1 U9903 ( .A(n8432), .ZN(n8437) );
  NOR2_X1 U9904 ( .A1(n8277), .A2(n8437), .ZN(n8487) );
  OR2_X1 U9905 ( .A1(n9800), .A2(n9233), .ZN(n8278) );
  NAND2_X1 U9906 ( .A1(n8424), .A2(n8278), .ZN(n8333) );
  NAND2_X1 U9907 ( .A1(n8333), .A2(n9618), .ZN(n8279) );
  NAND2_X1 U9908 ( .A1(n9600), .A2(n8279), .ZN(n8280) );
  NAND2_X1 U9909 ( .A1(n8280), .A2(n8427), .ZN(n8288) );
  OR2_X1 U9910 ( .A1(n9671), .A2(n9337), .ZN(n8421) );
  INV_X1 U9911 ( .A(n8421), .ZN(n8283) );
  AND2_X1 U9912 ( .A1(n8422), .A2(n8405), .ZN(n8418) );
  NAND2_X1 U9913 ( .A1(n9618), .A2(n8281), .ZN(n8332) );
  INV_X1 U9914 ( .A(n8332), .ZN(n8282) );
  OAI211_X1 U9915 ( .C1(n8283), .C2(n8418), .A(n8427), .B(n8282), .ZN(n8284)
         );
  NAND3_X1 U9916 ( .A1(n8435), .A2(n8288), .A3(n8284), .ZN(n8285) );
  NAND2_X1 U9917 ( .A1(n8285), .A2(n8430), .ZN(n8287) );
  NAND2_X1 U9918 ( .A1(n9533), .A2(n8286), .ZN(n8439) );
  AOI21_X1 U9919 ( .B1(n8487), .B2(n8287), .A(n8439), .ZN(n8490) );
  AND2_X1 U9920 ( .A1(n8421), .A2(n8335), .ZN(n8417) );
  NAND3_X1 U9921 ( .A1(n8288), .A2(n8435), .A3(n8417), .ZN(n8485) );
  AND2_X1 U9922 ( .A1(n8334), .A2(n8409), .ZN(n8336) );
  NAND2_X1 U9923 ( .A1(n8410), .A2(n8289), .ZN(n8291) );
  AOI21_X1 U9924 ( .B1(n8336), .B2(n8291), .A(n8290), .ZN(n8406) );
  AND2_X1 U9925 ( .A1(n8396), .A2(n8292), .ZN(n8382) );
  INV_X1 U9926 ( .A(n8382), .ZN(n8319) );
  AND2_X1 U9927 ( .A1(n8394), .A2(n8380), .ZN(n8388) );
  INV_X1 U9928 ( .A(n8388), .ZN(n8317) );
  NAND2_X1 U9929 ( .A1(n8294), .A2(n8293), .ZN(n8339) );
  INV_X1 U9930 ( .A(n8339), .ZN(n8302) );
  NAND2_X1 U9931 ( .A1(n5914), .A2(n4998), .ZN(n8295) );
  NAND4_X1 U9932 ( .A1(n8297), .A2(n8296), .A3(n8456), .A4(n8295), .ZN(n8301)
         );
  AND2_X1 U9933 ( .A1(n8299), .A2(n8298), .ZN(n8338) );
  INV_X1 U9934 ( .A(n8338), .ZN(n8300) );
  AOI21_X1 U9935 ( .B1(n8302), .B2(n8301), .A(n8300), .ZN(n8304) );
  NAND2_X1 U9936 ( .A1(n8303), .A2(n8343), .ZN(n8337) );
  OAI21_X1 U9937 ( .B1(n8304), .B2(n8337), .A(n8340), .ZN(n8307) );
  INV_X1 U9938 ( .A(n8305), .ZN(n8306) );
  NAND3_X1 U9939 ( .A1(n8307), .A2(n8306), .A3(n9963), .ZN(n8309) );
  AND2_X1 U9940 ( .A1(n8371), .A2(n8368), .ZN(n8363) );
  INV_X1 U9941 ( .A(n8363), .ZN(n8310) );
  AOI21_X1 U9942 ( .B1(n8309), .B2(n8308), .A(n8310), .ZN(n8314) );
  OR2_X1 U9943 ( .A1(n8310), .A2(n8370), .ZN(n8311) );
  AND3_X1 U9944 ( .A1(n8312), .A2(n8311), .A3(n8369), .ZN(n8365) );
  INV_X1 U9945 ( .A(n8365), .ZN(n8313) );
  OAI211_X1 U9946 ( .C1(n8314), .C2(n8313), .A(n8379), .B(n8372), .ZN(n8315)
         );
  AND3_X1 U9947 ( .A1(n8381), .A2(n8385), .A3(n8315), .ZN(n8316) );
  NOR2_X1 U9948 ( .A1(n8317), .A2(n8316), .ZN(n8318) );
  OAI21_X1 U9949 ( .B1(n8319), .B2(n8318), .A(n8398), .ZN(n8320) );
  NAND3_X1 U9950 ( .A1(n8336), .A2(n8408), .A3(n8320), .ZN(n8321) );
  AND2_X1 U9951 ( .A1(n8406), .A2(n8321), .ZN(n8322) );
  OAI21_X1 U9952 ( .B1(n8485), .B2(n8322), .A(n9572), .ZN(n8323) );
  NAND2_X1 U9953 ( .A1(n8487), .A2(n8323), .ZN(n8324) );
  NAND2_X1 U9954 ( .A1(n8331), .A2(n8433), .ZN(n8488) );
  AOI21_X1 U9955 ( .B1(n8490), .B2(n8324), .A(n8488), .ZN(n8326) );
  INV_X1 U9956 ( .A(n8445), .ZN(n9536) );
  NAND2_X1 U9957 ( .A1(n8451), .A2(n9536), .ZN(n8325) );
  NOR2_X1 U9958 ( .A1(n9852), .A2(n9399), .ZN(n8442) );
  NAND2_X1 U9959 ( .A1(n8325), .A2(n8330), .ZN(n8491) );
  OAI21_X1 U9960 ( .B1(n8326), .B2(n8491), .A(n8494), .ZN(n8327) );
  INV_X1 U9961 ( .A(n8493), .ZN(n8495) );
  AOI21_X1 U9962 ( .B1(n8327), .B2(n8510), .A(n8508), .ZN(n8329) );
  NOR2_X1 U9963 ( .A1(n8329), .A2(n8509), .ZN(n8506) );
  INV_X1 U9964 ( .A(n8444), .ZN(n8453) );
  MUX2_X1 U9965 ( .A(n8333), .B(n8332), .S(n8444), .Z(n8426) );
  AOI21_X1 U9966 ( .B1(n8335), .B2(n8334), .A(n8444), .ZN(n8420) );
  INV_X1 U9967 ( .A(n8336), .ZN(n8407) );
  AOI21_X1 U9968 ( .B1(n8339), .B2(n8338), .A(n8337), .ZN(n8342) );
  NAND2_X1 U9969 ( .A1(n8346), .A2(n8340), .ZN(n8341) );
  OAI21_X1 U9970 ( .B1(n8342), .B2(n8341), .A(n9963), .ZN(n8348) );
  OAI211_X1 U9971 ( .C1(n8345), .C2(n8344), .A(n9963), .B(n8343), .ZN(n8347)
         );
  MUX2_X1 U9972 ( .A(n8351), .B(n8350), .S(n8444), .Z(n8352) );
  INV_X1 U9973 ( .A(n8352), .ZN(n8353) );
  INV_X1 U9974 ( .A(n8354), .ZN(n8357) );
  NAND2_X1 U9975 ( .A1(n8362), .A2(n8355), .ZN(n8356) );
  MUX2_X1 U9976 ( .A(n8357), .B(n8356), .S(n8453), .Z(n8359) );
  NOR2_X1 U9977 ( .A1(n8359), .A2(n8358), .ZN(n8360) );
  NAND3_X1 U9978 ( .A1(n8367), .A2(n8363), .A3(n8362), .ZN(n8366) );
  INV_X1 U9979 ( .A(n8372), .ZN(n8364) );
  AOI21_X1 U9980 ( .B1(n8366), .B2(n8365), .A(n8364), .ZN(n8377) );
  AND2_X1 U9981 ( .A1(n8372), .A2(n8371), .ZN(n8374) );
  AOI21_X1 U9982 ( .B1(n8375), .B2(n8374), .A(n8373), .ZN(n8376) );
  MUX2_X1 U9983 ( .A(n8377), .B(n8376), .S(n8453), .Z(n8387) );
  INV_X1 U9984 ( .A(n8385), .ZN(n8378) );
  AOI21_X1 U9985 ( .B1(n8387), .B2(n8379), .A(n8378), .ZN(n8384) );
  INV_X1 U9986 ( .A(n8380), .ZN(n8383) );
  OAI211_X1 U9987 ( .C1(n8384), .C2(n8383), .A(n8382), .B(n8381), .ZN(n8393)
         );
  OAI211_X1 U9988 ( .C1(n8387), .C2(n8386), .A(n9752), .B(n8385), .ZN(n8391)
         );
  AND2_X1 U9989 ( .A1(n8398), .A2(n8388), .ZN(n8390) );
  AOI21_X1 U9990 ( .B1(n8391), .B2(n8390), .A(n8389), .ZN(n8392) );
  MUX2_X1 U9991 ( .A(n8393), .B(n8392), .S(n8453), .Z(n8403) );
  INV_X1 U9992 ( .A(n8394), .ZN(n8395) );
  NAND2_X1 U9993 ( .A1(n8396), .A2(n8395), .ZN(n8397) );
  OAI211_X1 U9994 ( .C1(n9396), .C2(n8444), .A(n8397), .B(n8398), .ZN(n8401)
         );
  NAND2_X1 U9995 ( .A1(n8398), .A2(n9410), .ZN(n8399) );
  NAND2_X1 U9996 ( .A1(n8399), .A2(n8453), .ZN(n8400) );
  NAND2_X1 U9997 ( .A1(n8401), .A2(n8400), .ZN(n8402) );
  NAND2_X1 U9998 ( .A1(n8403), .A2(n8402), .ZN(n8404) );
  NAND2_X1 U9999 ( .A1(n8404), .A2(n9734), .ZN(n8414) );
  OAI211_X1 U10000 ( .C1(n8407), .C2(n8414), .A(n8406), .B(n8405), .ZN(n8416)
         );
  AND2_X1 U10001 ( .A1(n8409), .A2(n8408), .ZN(n8413) );
  NAND2_X1 U10002 ( .A1(n8411), .A2(n8410), .ZN(n8412) );
  AOI21_X1 U10003 ( .B1(n8414), .B2(n8413), .A(n8412), .ZN(n8415) );
  MUX2_X1 U10004 ( .A(n8418), .B(n8417), .S(n8444), .Z(n8419) );
  MUX2_X1 U10005 ( .A(n8422), .B(n8421), .S(n8453), .Z(n8423) );
  MUX2_X1 U10006 ( .A(n9618), .B(n8424), .S(n8444), .Z(n8425) );
  MUX2_X1 U10007 ( .A(n9600), .B(n8427), .S(n8444), .Z(n8428) );
  NAND2_X1 U10008 ( .A1(n8429), .A2(n8428), .ZN(n8436) );
  AND2_X1 U10009 ( .A1(n9572), .A2(n8430), .ZN(n8438) );
  OR3_X1 U10010 ( .A1(n8439), .A2(n8453), .A3(n8434), .ZN(n8440) );
  NAND2_X1 U10011 ( .A1(n8452), .A2(n9933), .ZN(n8450) );
  NAND2_X1 U10012 ( .A1(n8447), .A2(n8446), .ZN(n8448) );
  NOR3_X1 U10013 ( .A1(n8458), .A2(n8457), .A3(n8456), .ZN(n8463) );
  NOR3_X1 U10014 ( .A1(n8461), .A2(n8460), .A3(n8459), .ZN(n8462) );
  NOR4_X1 U10015 ( .A1(n8468), .A2(n8467), .A3(n8466), .A4(n8465), .ZN(n8469)
         );
  NAND4_X1 U10016 ( .A1(n9752), .A2(n8471), .A3(n8470), .A4(n8469), .ZN(n8472)
         );
  NOR4_X1 U10017 ( .A1(n9728), .A2(n8474), .A3(n8473), .A4(n8472), .ZN(n8476)
         );
  NAND2_X1 U10018 ( .A1(n8476), .A2(n8475), .ZN(n8477) );
  NOR4_X1 U10019 ( .A1(n8479), .A2(n9702), .A3(n8478), .A4(n8477), .ZN(n8480)
         );
  NAND4_X1 U10020 ( .A1(n9617), .A2(n8480), .A3(n9664), .A4(n9655), .ZN(n8481)
         );
  NOR4_X1 U10021 ( .A1(n9564), .A2(n9582), .A3(n9601), .A4(n8481), .ZN(n8482)
         );
  NAND4_X1 U10022 ( .A1(n8494), .A2(n9531), .A3(n8482), .A4(n8331), .ZN(n8483)
         );
  OAI21_X1 U10023 ( .B1(n8485), .B2(n9682), .A(n9572), .ZN(n8486) );
  NAND2_X1 U10024 ( .A1(n8487), .A2(n8486), .ZN(n8489) );
  AOI21_X1 U10025 ( .B1(n8490), .B2(n8489), .A(n8488), .ZN(n8497) );
  INV_X1 U10026 ( .A(n8491), .ZN(n8492) );
  OAI21_X1 U10027 ( .B1(n9933), .B2(n8493), .A(n8492), .ZN(n8496) );
  OAI22_X1 U10028 ( .A1(n8497), .A2(n8496), .B1(n8495), .B2(n8494), .ZN(n8499)
         );
  AOI211_X1 U10029 ( .C1(n8499), .C2(n8510), .A(n8498), .B(n8508), .ZN(n8500)
         );
  NOR2_X1 U10030 ( .A1(n8502), .A2(n8500), .ZN(n8501) );
  OAI22_X1 U10031 ( .A1(n8503), .A2(n8502), .B1(n4509), .B2(n8501), .ZN(n8505)
         );
  NOR3_X1 U10032 ( .A1(n8514), .A2(n9893), .A3(n8513), .ZN(n8517) );
  OAI21_X1 U10033 ( .B1(n8518), .B2(n8515), .A(P1_B_REG_SCAN_IN), .ZN(n8516)
         );
  OAI22_X1 U10034 ( .A1(n8519), .A2(n8518), .B1(n8517), .B2(n8516), .ZN(
        P1_U3242) );
  NOR2_X1 U10035 ( .A1(P1_REG2_REG_17__SCAN_IN), .A2(n9501), .ZN(n8520) );
  AOI21_X1 U10036 ( .B1(n9501), .B2(P1_REG2_REG_17__SCAN_IN), .A(n8520), .ZN(
        n9493) );
  NAND2_X1 U10037 ( .A1(n9493), .A2(n9492), .ZN(n9491) );
  OAI21_X1 U10038 ( .B1(P1_REG2_REG_17__SCAN_IN), .B2(n9501), .A(n9491), .ZN(
        n8522) );
  INV_X1 U10039 ( .A(n8522), .ZN(n9520) );
  NAND2_X1 U10040 ( .A1(n9515), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n8524) );
  OAI21_X1 U10041 ( .B1(n9515), .B2(P1_REG2_REG_18__SCAN_IN), .A(n8524), .ZN(
        n8523) );
  INV_X1 U10042 ( .A(n8523), .ZN(n9519) );
  NAND2_X1 U10043 ( .A1(n9520), .A2(n9519), .ZN(n9518) );
  NAND2_X1 U10044 ( .A1(n9518), .A2(n8524), .ZN(n8525) );
  XNOR2_X1 U10045 ( .A(n8525), .B(P1_REG2_REG_19__SCAN_IN), .ZN(n8534) );
  INV_X1 U10046 ( .A(n8534), .ZN(n8532) );
  AOI22_X1 U10047 ( .A1(P1_REG1_REG_17__SCAN_IN), .A2(n9501), .B1(n8526), .B2(
        n6277), .ZN(n9498) );
  OAI21_X1 U10048 ( .B1(n8528), .B2(P1_REG1_REG_16__SCAN_IN), .A(n8527), .ZN(
        n9497) );
  NAND2_X1 U10049 ( .A1(n9498), .A2(n9497), .ZN(n9496) );
  OAI21_X1 U10050 ( .B1(n9501), .B2(P1_REG1_REG_17__SCAN_IN), .A(n9496), .ZN(
        n9512) );
  NAND2_X1 U10051 ( .A1(n9515), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n8529) );
  OAI21_X1 U10052 ( .B1(n9515), .B2(P1_REG1_REG_18__SCAN_IN), .A(n8529), .ZN(
        n9511) );
  OR2_X1 U10053 ( .A1(n9512), .A2(n9511), .ZN(n9508) );
  NAND2_X1 U10054 ( .A1(n9508), .A2(n8529), .ZN(n8531) );
  XNOR2_X1 U10055 ( .A(n8531), .B(n8530), .ZN(n8533) );
  AOI22_X1 U10056 ( .A1(n8532), .A2(n9517), .B1(n9499), .B2(n8533), .ZN(n8535)
         );
  NAND2_X1 U10057 ( .A1(P1_REG3_REG_19__SCAN_IN), .A2(P1_U3086), .ZN(n8536) );
  INV_X1 U10058 ( .A(n8537), .ZN(n8593) );
  OAI222_X1 U10059 ( .A1(P2_U3151), .A2(n8538), .B1(n9171), .B2(n8593), .C1(
        n8539), .C2(n8185), .ZN(P2_U3265) );
  OAI222_X1 U10060 ( .A1(n8860), .A2(P2_U3151), .B1(n9171), .B2(n8541), .C1(
        n8540), .C2(n8539), .ZN(P2_U3268) );
  XNOR2_X1 U10061 ( .A(n9125), .B(n7074), .ZN(n8685) );
  XNOR2_X1 U10062 ( .A(n8647), .B(n7074), .ZN(n8640) );
  INV_X1 U10063 ( .A(n8640), .ZN(n8547) );
  XNOR2_X1 U10064 ( .A(n9153), .B(n8580), .ZN(n8548) );
  NAND2_X1 U10065 ( .A1(n8548), .A2(n9005), .ZN(n8549) );
  OAI21_X1 U10066 ( .B1(n8548), .B2(n9005), .A(n8549), .ZN(n8651) );
  INV_X1 U10067 ( .A(n8549), .ZN(n8702) );
  XNOR2_X1 U10068 ( .A(n8699), .B(n8580), .ZN(n8550) );
  NAND2_X1 U10069 ( .A1(n8550), .A2(n8994), .ZN(n8612) );
  INV_X1 U10070 ( .A(n8550), .ZN(n8551) );
  NAND2_X1 U10071 ( .A1(n8551), .A2(n9024), .ZN(n8552) );
  AND2_X1 U10072 ( .A1(n8612), .A2(n8552), .ZN(n8701) );
  XNOR2_X1 U10073 ( .A(n9067), .B(n8580), .ZN(n8553) );
  NAND2_X1 U10074 ( .A1(n8553), .A2(n9007), .ZN(n8556) );
  INV_X1 U10075 ( .A(n8553), .ZN(n8554) );
  NAND2_X1 U10076 ( .A1(n8554), .A2(n8981), .ZN(n8555) );
  NAND2_X1 U10077 ( .A1(n8556), .A2(n8555), .ZN(n8611) );
  INV_X1 U10078 ( .A(n8556), .ZN(n8673) );
  XNOR2_X1 U10079 ( .A(n9137), .B(n8580), .ZN(n8557) );
  NAND2_X1 U10080 ( .A1(n8557), .A2(n8995), .ZN(n8619) );
  INV_X1 U10081 ( .A(n8557), .ZN(n8558) );
  NAND2_X1 U10082 ( .A1(n8558), .A2(n8972), .ZN(n8559) );
  AND2_X1 U10083 ( .A1(n8619), .A2(n8559), .ZN(n8672) );
  XNOR2_X1 U10084 ( .A(n9131), .B(n8580), .ZN(n8560) );
  XNOR2_X1 U10085 ( .A(n8560), .B(n8678), .ZN(n8620) );
  INV_X1 U10086 ( .A(n8560), .ZN(n8561) );
  NAND2_X1 U10087 ( .A1(n8685), .A2(n8971), .ZN(n8690) );
  XNOR2_X1 U10088 ( .A(n9119), .B(n8580), .ZN(n8564) );
  INV_X1 U10089 ( .A(n8564), .ZN(n8562) );
  NAND2_X1 U10090 ( .A1(n8605), .A2(n8660), .ZN(n8569) );
  XNOR2_X1 U10091 ( .A(n9113), .B(n8580), .ZN(n8566) );
  NAND2_X1 U10092 ( .A1(n8566), .A2(n8925), .ZN(n8630) );
  INV_X1 U10093 ( .A(n8566), .ZN(n8567) );
  NAND2_X1 U10094 ( .A1(n8567), .A2(n8945), .ZN(n8568) );
  NAND2_X1 U10095 ( .A1(n8569), .A2(n8661), .ZN(n8629) );
  NAND2_X1 U10096 ( .A1(n8629), .A2(n8630), .ZN(n8573) );
  XNOR2_X1 U10097 ( .A(n8628), .B(n8580), .ZN(n8570) );
  NAND2_X1 U10098 ( .A1(n8570), .A2(n8667), .ZN(n8712) );
  INV_X1 U10099 ( .A(n8570), .ZN(n8571) );
  NAND2_X1 U10100 ( .A1(n8571), .A2(n8935), .ZN(n8572) );
  NAND2_X1 U10101 ( .A1(n8573), .A2(n8631), .ZN(n8633) );
  NAND2_X1 U10102 ( .A1(n8633), .A2(n8712), .ZN(n8574) );
  XNOR2_X1 U10103 ( .A(n9102), .B(n8580), .ZN(n8575) );
  XNOR2_X1 U10104 ( .A(n8575), .B(n8901), .ZN(n8713) );
  XNOR2_X1 U10105 ( .A(n9095), .B(n8580), .ZN(n8578) );
  XNOR2_X1 U10106 ( .A(n8578), .B(n8587), .ZN(n8595) );
  INV_X1 U10107 ( .A(n8595), .ZN(n8577) );
  NAND2_X1 U10108 ( .A1(n8596), .A2(n8579), .ZN(n8583) );
  XNOR2_X1 U10109 ( .A(n8581), .B(n8580), .ZN(n8582) );
  XNOR2_X1 U10110 ( .A(n8583), .B(n8582), .ZN(n8592) );
  NOR2_X1 U10111 ( .A1(n8584), .A2(n8707), .ZN(n8589) );
  AOI22_X1 U10112 ( .A1(n8585), .A2(n8709), .B1(P2_REG3_REG_28__SCAN_IN), .B2(
        P2_U3151), .ZN(n8586) );
  OAI21_X1 U10113 ( .B1(n8587), .B2(n8677), .A(n8586), .ZN(n8588) );
  AOI211_X1 U10114 ( .C1(n8590), .C2(n8655), .A(n8589), .B(n8588), .ZN(n8591)
         );
  OAI21_X1 U10115 ( .B1(n8592), .B2(n8658), .A(n8591), .ZN(P2_U3160) );
  OAI222_X1 U10116 ( .A1(n9903), .A2(n10372), .B1(n9905), .B2(n8593), .C1(
        P1_U3086), .C2(n5874), .ZN(P1_U3325) );
  AOI21_X1 U10117 ( .B1(n8594), .B2(n8595), .A(n8658), .ZN(n8598) );
  NAND2_X1 U10118 ( .A1(n8598), .A2(n8597), .ZN(n8602) );
  AOI22_X1 U10119 ( .A1(n8906), .A2(n8709), .B1(P2_REG3_REG_27__SCAN_IN), .B2(
        P2_U3151), .ZN(n8599) );
  OAI21_X1 U10120 ( .B1(n8924), .B2(n8677), .A(n8599), .ZN(n8600) );
  AOI21_X1 U10121 ( .B1(n8725), .B2(n8902), .A(n8600), .ZN(n8601) );
  OAI211_X1 U10122 ( .C1(n8603), .C2(n8728), .A(n8602), .B(n8601), .ZN(
        P2_U3154) );
  INV_X1 U10123 ( .A(n8605), .ZN(n8663) );
  AOI21_X1 U10124 ( .B1(n8958), .B2(n8604), .A(n8663), .ZN(n8610) );
  AOI22_X1 U10125 ( .A1(n8945), .A2(n8725), .B1(P2_REG3_REG_23__SCAN_IN), .B2(
        P2_U3151), .ZN(n8607) );
  NAND2_X1 U10126 ( .A1(n8948), .A2(n8709), .ZN(n8606) );
  OAI211_X1 U10127 ( .C1(n8684), .C2(n8677), .A(n8607), .B(n8606), .ZN(n8608)
         );
  AOI21_X1 U10128 ( .B1(n9119), .B2(n8655), .A(n8608), .ZN(n8609) );
  OAI21_X1 U10129 ( .B1(n8610), .B2(n8658), .A(n8609), .ZN(P2_U3156) );
  INV_X1 U10130 ( .A(n9067), .ZN(n8618) );
  AND3_X1 U10131 ( .A1(n8700), .A2(n8612), .A3(n8611), .ZN(n8613) );
  OAI21_X1 U10132 ( .B1(n8674), .B2(n8613), .A(n8717), .ZN(n8617) );
  NAND2_X1 U10133 ( .A1(n9024), .A2(n8720), .ZN(n8614) );
  NAND2_X1 U10134 ( .A1(P2_U3151), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n8868) );
  OAI211_X1 U10135 ( .C1(n8995), .C2(n8707), .A(n8614), .B(n8868), .ZN(n8615)
         );
  AOI21_X1 U10136 ( .B1(n8996), .B2(n8709), .A(n8615), .ZN(n8616) );
  OAI211_X1 U10137 ( .C1(n8618), .C2(n8728), .A(n8617), .B(n8616), .ZN(
        P2_U3159) );
  INV_X1 U10138 ( .A(n9131), .ZN(n8627) );
  AND3_X1 U10139 ( .A1(n8671), .A2(n8620), .A3(n8619), .ZN(n8621) );
  OAI21_X1 U10140 ( .B1(n8622), .B2(n8621), .A(n8717), .ZN(n8626) );
  AOI22_X1 U10141 ( .A1(n8972), .A2(n8720), .B1(P2_REG3_REG_21__SCAN_IN), .B2(
        P2_U3151), .ZN(n8623) );
  OAI21_X1 U10142 ( .B1(n8684), .B2(n8707), .A(n8623), .ZN(n8624) );
  AOI21_X1 U10143 ( .B1(n8975), .B2(n8709), .A(n8624), .ZN(n8625) );
  OAI211_X1 U10144 ( .C1(n8627), .C2(n8728), .A(n8626), .B(n8625), .ZN(
        P2_U3163) );
  INV_X1 U10145 ( .A(n8628), .ZN(n9107) );
  INV_X1 U10146 ( .A(n8629), .ZN(n8664) );
  INV_X1 U10147 ( .A(n8630), .ZN(n8632) );
  NOR3_X1 U10148 ( .A1(n8664), .A2(n8632), .A3(n8631), .ZN(n8634) );
  INV_X1 U10149 ( .A(n8633), .ZN(n8715) );
  OAI21_X1 U10150 ( .B1(n8634), .B2(n8715), .A(n8717), .ZN(n8639) );
  INV_X1 U10151 ( .A(n8635), .ZN(n8926) );
  AOI22_X1 U10152 ( .A1(n8945), .A2(n8720), .B1(P2_REG3_REG_25__SCAN_IN), .B2(
        P2_U3151), .ZN(n8636) );
  OAI21_X1 U10153 ( .B1(n8926), .B2(n8722), .A(n8636), .ZN(n8637) );
  AOI21_X1 U10154 ( .B1(n8725), .B2(n8901), .A(n8637), .ZN(n8638) );
  OAI211_X1 U10155 ( .C1(n9107), .C2(n8728), .A(n8639), .B(n8638), .ZN(
        P2_U3165) );
  XNOR2_X1 U10156 ( .A(n8640), .B(n8653), .ZN(n8641) );
  XNOR2_X1 U10157 ( .A(n8642), .B(n8641), .ZN(n8649) );
  NAND2_X1 U10158 ( .A1(P2_U3151), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n8785) );
  OAI21_X1 U10159 ( .B1(n9005), .B2(n8707), .A(n8785), .ZN(n8643) );
  AOI21_X1 U10160 ( .B1(n8720), .B2(n8733), .A(n8643), .ZN(n8644) );
  OAI21_X1 U10161 ( .B1(n8645), .B2(n8722), .A(n8644), .ZN(n8646) );
  AOI21_X1 U10162 ( .B1(n8647), .B2(n8655), .A(n8646), .ZN(n8648) );
  OAI21_X1 U10163 ( .B1(n8649), .B2(n8658), .A(n8648), .ZN(P2_U3166) );
  AOI21_X1 U10164 ( .B1(n8651), .B2(n8650), .A(n8703), .ZN(n8659) );
  NAND2_X1 U10165 ( .A1(n9024), .A2(n8725), .ZN(n8652) );
  NAND2_X1 U10166 ( .A1(P2_U3151), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n8804) );
  OAI211_X1 U10167 ( .C1(n8653), .C2(n8677), .A(n8652), .B(n8804), .ZN(n8654)
         );
  AOI21_X1 U10168 ( .B1(n9030), .B2(n8709), .A(n8654), .ZN(n8657) );
  NAND2_X1 U10169 ( .A1(n9153), .A2(n8655), .ZN(n8656) );
  OAI211_X1 U10170 ( .C1(n8659), .C2(n8658), .A(n8657), .B(n8656), .ZN(
        P2_U3168) );
  INV_X1 U10171 ( .A(n9113), .ZN(n8937) );
  INV_X1 U10172 ( .A(n8660), .ZN(n8662) );
  NOR3_X1 U10173 ( .A1(n8663), .A2(n8662), .A3(n8661), .ZN(n8665) );
  OAI21_X1 U10174 ( .B1(n8665), .B2(n8664), .A(n8717), .ZN(n8670) );
  AOI22_X1 U10175 ( .A1(n8958), .A2(n8720), .B1(P2_REG3_REG_24__SCAN_IN), .B2(
        P2_U3151), .ZN(n8666) );
  OAI21_X1 U10176 ( .B1(n8667), .B2(n8707), .A(n8666), .ZN(n8668) );
  AOI21_X1 U10177 ( .B1(n8939), .B2(n8709), .A(n8668), .ZN(n8669) );
  OAI211_X1 U10178 ( .C1(n8937), .C2(n8728), .A(n8670), .B(n8669), .ZN(
        P2_U3169) );
  INV_X1 U10179 ( .A(n9137), .ZN(n8683) );
  INV_X1 U10180 ( .A(n8671), .ZN(n8676) );
  NOR3_X1 U10181 ( .A1(n8674), .A2(n8673), .A3(n8672), .ZN(n8675) );
  OAI21_X1 U10182 ( .B1(n8676), .B2(n8675), .A(n8717), .ZN(n8682) );
  NOR2_X1 U10183 ( .A1(n9007), .A2(n8677), .ZN(n8680) );
  INV_X1 U10184 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n10613) );
  OAI22_X1 U10185 ( .A1(n8678), .A2(n8707), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10613), .ZN(n8679) );
  AOI211_X1 U10186 ( .C1(n8985), .C2(n8709), .A(n8680), .B(n8679), .ZN(n8681)
         );
  OAI211_X1 U10187 ( .C1(n8683), .C2(n8728), .A(n8682), .B(n8681), .ZN(
        P2_U3173) );
  INV_X1 U10188 ( .A(n9125), .ZN(n8698) );
  INV_X1 U10189 ( .A(n8688), .ZN(n8691) );
  XNOR2_X1 U10190 ( .A(n8685), .B(n8684), .ZN(n8687) );
  OAI21_X1 U10191 ( .B1(n8688), .B2(n8687), .A(n8686), .ZN(n8689) );
  OAI21_X1 U10192 ( .B1(n8691), .B2(n8690), .A(n8689), .ZN(n8692) );
  NAND2_X1 U10193 ( .A1(n8692), .A2(n8717), .ZN(n8697) );
  AOI22_X1 U10194 ( .A1(n8982), .A2(n8720), .B1(P2_REG3_REG_22__SCAN_IN), .B2(
        P2_U3151), .ZN(n8693) );
  OAI21_X1 U10195 ( .B1(n8694), .B2(n8707), .A(n8693), .ZN(n8695) );
  AOI21_X1 U10196 ( .B1(n8961), .B2(n8709), .A(n8695), .ZN(n8696) );
  OAI211_X1 U10197 ( .C1(n8698), .C2(n8728), .A(n8697), .B(n8696), .ZN(
        P2_U3175) );
  INV_X1 U10198 ( .A(n8699), .ZN(n9149) );
  INV_X1 U10199 ( .A(n8700), .ZN(n8705) );
  NOR3_X1 U10200 ( .A1(n8703), .A2(n8702), .A3(n8701), .ZN(n8704) );
  OAI21_X1 U10201 ( .B1(n8705), .B2(n8704), .A(n8717), .ZN(n8711) );
  NAND2_X1 U10202 ( .A1(n8731), .A2(n8720), .ZN(n8706) );
  NAND2_X1 U10203 ( .A1(P2_U3151), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n8834) );
  OAI211_X1 U10204 ( .C1(n9007), .C2(n8707), .A(n8706), .B(n8834), .ZN(n8708)
         );
  AOI21_X1 U10205 ( .B1(n9012), .B2(n8709), .A(n8708), .ZN(n8710) );
  OAI211_X1 U10206 ( .C1(n9149), .C2(n8728), .A(n8711), .B(n8710), .ZN(
        P2_U3178) );
  INV_X1 U10207 ( .A(n8712), .ZN(n8714) );
  NOR3_X1 U10208 ( .A1(n8715), .A2(n8714), .A3(n8713), .ZN(n8719) );
  INV_X1 U10209 ( .A(n8716), .ZN(n8718) );
  OAI21_X1 U10210 ( .B1(n8719), .B2(n8718), .A(n8717), .ZN(n8727) );
  INV_X1 U10211 ( .A(n8917), .ZN(n8723) );
  AOI22_X1 U10212 ( .A1(n8935), .A2(n8720), .B1(P2_REG3_REG_26__SCAN_IN), .B2(
        P2_U3151), .ZN(n8721) );
  OAI21_X1 U10213 ( .B1(n8723), .B2(n8722), .A(n8721), .ZN(n8724) );
  AOI21_X1 U10214 ( .B1(n8725), .B2(n8914), .A(n8724), .ZN(n8726) );
  OAI211_X1 U10215 ( .C1(n8729), .C2(n8728), .A(n8727), .B(n8726), .ZN(
        P2_U3180) );
  MUX2_X1 U10216 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(n8730), .S(P2_U3893), .Z(
        P2_U3521) );
  MUX2_X1 U10217 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(n8902), .S(P2_U3893), .Z(
        P2_U3519) );
  MUX2_X1 U10218 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(n8901), .S(P2_U3893), .Z(
        P2_U3517) );
  MUX2_X1 U10219 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n8935), .S(P2_U3893), .Z(
        P2_U3516) );
  MUX2_X1 U10220 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(n8945), .S(P2_U3893), .Z(
        P2_U3515) );
  MUX2_X1 U10221 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n8971), .S(P2_U3893), .Z(
        P2_U3513) );
  MUX2_X1 U10222 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n8982), .S(P2_U3893), .Z(
        P2_U3512) );
  MUX2_X1 U10223 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n8972), .S(P2_U3893), .Z(
        P2_U3511) );
  MUX2_X1 U10224 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n8981), .S(P2_U3893), .Z(
        P2_U3510) );
  MUX2_X1 U10225 ( .A(n9024), .B(P2_DATAO_REG_18__SCAN_IN), .S(n8832), .Z(
        P2_U3509) );
  MUX2_X1 U10226 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n8731), .S(P2_U3893), .Z(
        P2_U3508) );
  MUX2_X1 U10227 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n9026), .S(P2_U3893), .Z(
        P2_U3507) );
  MUX2_X1 U10228 ( .A(n8733), .B(P2_DATAO_REG_15__SCAN_IN), .S(n8832), .Z(
        P2_U3506) );
  MUX2_X1 U10229 ( .A(n8734), .B(P2_DATAO_REG_14__SCAN_IN), .S(n8832), .Z(
        P2_U3505) );
  MUX2_X1 U10230 ( .A(n8735), .B(P2_DATAO_REG_12__SCAN_IN), .S(n8832), .Z(
        P2_U3503) );
  MUX2_X1 U10231 ( .A(n8736), .B(P2_DATAO_REG_11__SCAN_IN), .S(n8832), .Z(
        P2_U3502) );
  MUX2_X1 U10232 ( .A(n8737), .B(P2_DATAO_REG_10__SCAN_IN), .S(n8832), .Z(
        P2_U3501) );
  MUX2_X1 U10233 ( .A(n8738), .B(P2_DATAO_REG_9__SCAN_IN), .S(n8832), .Z(
        P2_U3500) );
  MUX2_X1 U10234 ( .A(n8739), .B(P2_DATAO_REG_8__SCAN_IN), .S(n8832), .Z(
        P2_U3499) );
  MUX2_X1 U10235 ( .A(n8740), .B(P2_DATAO_REG_7__SCAN_IN), .S(n8832), .Z(
        P2_U3498) );
  MUX2_X1 U10236 ( .A(n8741), .B(P2_DATAO_REG_6__SCAN_IN), .S(n8832), .Z(
        P2_U3497) );
  MUX2_X1 U10237 ( .A(n8742), .B(P2_DATAO_REG_4__SCAN_IN), .S(n8832), .Z(
        P2_U3495) );
  MUX2_X1 U10238 ( .A(n10149), .B(P2_DATAO_REG_3__SCAN_IN), .S(n8832), .Z(
        P2_U3494) );
  MUX2_X1 U10239 ( .A(n8743), .B(P2_DATAO_REG_2__SCAN_IN), .S(n8832), .Z(
        P2_U3493) );
  MUX2_X1 U10240 ( .A(n10147), .B(P2_DATAO_REG_1__SCAN_IN), .S(n8832), .Z(
        P2_U3492) );
  MUX2_X1 U10241 ( .A(n5317), .B(P2_DATAO_REG_0__SCAN_IN), .S(n8832), .Z(
        P2_U3491) );
  NOR2_X1 U10242 ( .A1(n8760), .A2(n8745), .ZN(n8746) );
  INV_X1 U10243 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n8747) );
  AOI22_X1 U10244 ( .A1(P2_REG2_REG_14__SCAN_IN), .A2(n8764), .B1(n10135), 
        .B2(n8747), .ZN(n10120) );
  AOI21_X1 U10245 ( .B1(n8748), .B2(n7998), .A(n8790), .ZN(n8773) );
  OAI21_X1 U10246 ( .B1(n8751), .B2(n8750), .A(n8749), .ZN(n10106) );
  MUX2_X1 U10247 ( .A(P2_REG2_REG_13__SCAN_IN), .B(P2_REG1_REG_13__SCAN_IN), 
        .S(n8860), .Z(n8752) );
  XNOR2_X1 U10248 ( .A(n8752), .B(n8760), .ZN(n10107) );
  INV_X1 U10249 ( .A(n8752), .ZN(n8753) );
  AOI22_X1 U10250 ( .A1(n10106), .A2(n10107), .B1(n8760), .B2(n8753), .ZN(
        n10121) );
  MUX2_X1 U10251 ( .A(P2_REG2_REG_14__SCAN_IN), .B(P2_REG1_REG_14__SCAN_IN), 
        .S(n8860), .Z(n8754) );
  XNOR2_X1 U10252 ( .A(n8754), .B(n10135), .ZN(n10122) );
  OAI22_X1 U10253 ( .A1(n10121), .A2(n10122), .B1(n8754), .B2(n10135), .ZN(
        n8783) );
  MUX2_X1 U10254 ( .A(P2_REG2_REG_15__SCAN_IN), .B(P2_REG1_REG_15__SCAN_IN), 
        .S(n8860), .Z(n8780) );
  XNOR2_X1 U10255 ( .A(n8780), .B(n8789), .ZN(n8782) );
  XNOR2_X1 U10256 ( .A(n8783), .B(n8782), .ZN(n8771) );
  INV_X1 U10257 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n8757) );
  NAND2_X1 U10258 ( .A1(n8872), .A2(n8789), .ZN(n8756) );
  OAI211_X1 U10259 ( .C1(n8757), .C2(n8870), .A(n8756), .B(n8755), .ZN(n8770)
         );
  NOR2_X1 U10260 ( .A1(n8760), .A2(n8761), .ZN(n8762) );
  XOR2_X1 U10261 ( .A(n8761), .B(n10117), .Z(n10109) );
  AOI22_X1 U10262 ( .A1(P2_REG1_REG_14__SCAN_IN), .A2(n8764), .B1(n10135), 
        .B2(n8763), .ZN(n10124) );
  AOI21_X1 U10263 ( .B1(n8767), .B2(n8766), .A(n8775), .ZN(n8768) );
  NOR2_X1 U10264 ( .A1(n8768), .A2(n10127), .ZN(n8769) );
  AOI211_X1 U10265 ( .C1(n8814), .C2(n8771), .A(n8770), .B(n8769), .ZN(n8772)
         );
  OAI21_X1 U10266 ( .B1(n8773), .B2(n10131), .A(n8772), .ZN(P2_U3197) );
  NOR2_X1 U10267 ( .A1(n8789), .A2(n8774), .ZN(n8776) );
  AOI22_X1 U10268 ( .A1(P2_REG1_REG_16__SCAN_IN), .A2(n8784), .B1(n8810), .B2(
        n8777), .ZN(n8778) );
  AOI21_X1 U10269 ( .B1(n8779), .B2(n8778), .A(n8801), .ZN(n8800) );
  INV_X1 U10270 ( .A(n8780), .ZN(n8781) );
  AOI22_X1 U10271 ( .A1(n8783), .A2(n8782), .B1(n8789), .B2(n8781), .ZN(n8813)
         );
  MUX2_X1 U10272 ( .A(P2_REG2_REG_16__SCAN_IN), .B(P2_REG1_REG_16__SCAN_IN), 
        .S(n8860), .Z(n8811) );
  XNOR2_X1 U10273 ( .A(n8811), .B(n8810), .ZN(n8812) );
  XNOR2_X1 U10274 ( .A(n8813), .B(n8812), .ZN(n8798) );
  INV_X1 U10275 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n8787) );
  NAND2_X1 U10276 ( .A1(n8872), .A2(n8784), .ZN(n8786) );
  OAI211_X1 U10277 ( .C1(n8787), .C2(n8870), .A(n8786), .B(n8785), .ZN(n8797)
         );
  NOR2_X1 U10278 ( .A1(n8789), .A2(n8788), .ZN(n8791) );
  NAND2_X1 U10279 ( .A1(P2_REG2_REG_16__SCAN_IN), .A2(n8810), .ZN(n8792) );
  OAI21_X1 U10280 ( .B1(n8810), .B2(P2_REG2_REG_16__SCAN_IN), .A(n8792), .ZN(
        n8793) );
  NOR2_X1 U10281 ( .A1(n8794), .A2(n8793), .ZN(n8806) );
  AOI21_X1 U10282 ( .B1(n8794), .B2(n8793), .A(n8806), .ZN(n8795) );
  NOR2_X1 U10283 ( .A1(n8795), .A2(n10131), .ZN(n8796) );
  AOI211_X1 U10284 ( .C1(n8814), .C2(n8798), .A(n8797), .B(n8796), .ZN(n8799)
         );
  OAI21_X1 U10285 ( .B1(n8800), .B2(n10127), .A(n8799), .ZN(P2_U3198) );
  INV_X1 U10286 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n9077) );
  AOI21_X1 U10287 ( .B1(n9077), .B2(n8803), .A(n8840), .ZN(n8818) );
  INV_X1 U10288 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n8805) );
  OAI21_X1 U10289 ( .B1(n8870), .B2(n8805), .A(n8804), .ZN(n8809) );
  AOI21_X1 U10290 ( .B1(P2_REG2_REG_16__SCAN_IN), .B2(n8810), .A(n8806), .ZN(
        n8819) );
  XNOR2_X1 U10291 ( .A(n8841), .B(n8819), .ZN(n8808) );
  INV_X1 U10292 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n8807) );
  OAI22_X1 U10293 ( .A1(n8813), .A2(n8812), .B1(n8811), .B2(n8810), .ZN(n8828)
         );
  MUX2_X1 U10294 ( .A(P2_REG2_REG_17__SCAN_IN), .B(P2_REG1_REG_17__SCAN_IN), 
        .S(n8860), .Z(n8825) );
  XNOR2_X1 U10295 ( .A(n8825), .B(n8841), .ZN(n8827) );
  XNOR2_X1 U10296 ( .A(n8828), .B(n8827), .ZN(n8815) );
  NAND2_X1 U10297 ( .A1(n8815), .A2(n8814), .ZN(n8816) );
  OAI211_X1 U10298 ( .C1(n8818), .C2(n10127), .A(n8817), .B(n8816), .ZN(
        P2_U3199) );
  NOR2_X1 U10299 ( .A1(n8841), .A2(n8819), .ZN(n8821) );
  NAND2_X1 U10300 ( .A1(n8822), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n8857) );
  OAI21_X1 U10301 ( .B1(n8822), .B2(P2_REG2_REG_18__SCAN_IN), .A(n8857), .ZN(
        n8823) );
  AOI21_X1 U10302 ( .B1(n8824), .B2(n8823), .A(n4574), .ZN(n8851) );
  INV_X1 U10303 ( .A(n8825), .ZN(n8826) );
  AOI22_X1 U10304 ( .A1(n8828), .A2(n8827), .B1(n8841), .B2(n8826), .ZN(n8830)
         );
  MUX2_X1 U10305 ( .A(P2_REG2_REG_18__SCAN_IN), .B(P2_REG1_REG_18__SCAN_IN), 
        .S(n8860), .Z(n8829) );
  NOR2_X1 U10306 ( .A1(n8830), .A2(n8829), .ZN(n8863) );
  NAND2_X1 U10307 ( .A1(n8830), .A2(n8829), .ZN(n8864) );
  INV_X1 U10308 ( .A(n8864), .ZN(n8831) );
  NOR2_X1 U10309 ( .A1(n8863), .A2(n8831), .ZN(n8836) );
  INV_X1 U10310 ( .A(n8836), .ZN(n8833) );
  OAI21_X1 U10311 ( .B1(n8833), .B2(n8832), .A(n10136), .ZN(n8839) );
  INV_X1 U10312 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n8835) );
  OAI21_X1 U10313 ( .B1(n8870), .B2(n8835), .A(n8834), .ZN(n8838) );
  NOR3_X1 U10314 ( .A1(n8836), .A2(n8865), .A3(n10129), .ZN(n8837) );
  AOI211_X1 U10315 ( .C1(n8865), .C2(n8839), .A(n8838), .B(n8837), .ZN(n8850)
         );
  OR2_X1 U10316 ( .A1(n8842), .A2(n8841), .ZN(n8845) );
  INV_X1 U10317 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n9074) );
  OR2_X1 U10318 ( .A1(n8865), .A2(n9074), .ZN(n8852) );
  NAND2_X1 U10319 ( .A1(n8865), .A2(n9074), .ZN(n8843) );
  NAND2_X1 U10320 ( .A1(n8852), .A2(n8843), .ZN(n8844) );
  AND3_X1 U10321 ( .A1(n8846), .A2(n8845), .A3(n8844), .ZN(n8848) );
  OAI21_X1 U10322 ( .B1(n8854), .B2(n8848), .A(n8847), .ZN(n8849) );
  OAI211_X1 U10323 ( .C1(n8851), .C2(n10131), .A(n8850), .B(n8849), .ZN(
        P2_U3200) );
  INV_X1 U10324 ( .A(n8852), .ZN(n8853) );
  XNOR2_X1 U10325 ( .A(n8859), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n8861) );
  INV_X1 U10326 ( .A(n8861), .ZN(n8855) );
  XNOR2_X1 U10327 ( .A(n8856), .B(n8855), .ZN(n8880) );
  INV_X1 U10328 ( .A(n8857), .ZN(n8858) );
  XNOR2_X1 U10329 ( .A(n8859), .B(P2_REG2_REG_19__SCAN_IN), .ZN(n8862) );
  MUX2_X1 U10330 ( .A(n8862), .B(n8861), .S(n8860), .Z(n8867) );
  AOI21_X1 U10331 ( .B1(n8865), .B2(n8864), .A(n8863), .ZN(n8866) );
  XOR2_X1 U10332 ( .A(n8867), .B(n8866), .Z(n8875) );
  OAI21_X1 U10333 ( .B1(n8870), .B2(n8869), .A(n8868), .ZN(n8871) );
  AOI21_X1 U10334 ( .B1(n8873), .B2(n8872), .A(n8871), .ZN(n8874) );
  OAI21_X1 U10335 ( .B1(n8875), .B2(n10129), .A(n8874), .ZN(n8876) );
  AOI21_X1 U10336 ( .B1(n8878), .B2(n8877), .A(n8876), .ZN(n8879) );
  OAI21_X1 U10337 ( .B1(n8880), .B2(n10127), .A(n8879), .ZN(P2_U3201) );
  NAND2_X1 U10338 ( .A1(n9081), .A2(n9032), .ZN(n8884) );
  NOR2_X1 U10339 ( .A1(n8883), .A2(n10141), .ZN(n8892) );
  AOI21_X1 U10340 ( .B1(n9082), .B2(n9029), .A(n8892), .ZN(n8886) );
  OAI211_X1 U10341 ( .C1(n9029), .C2(n8885), .A(n8884), .B(n8886), .ZN(
        P2_U3202) );
  NAND2_X1 U10342 ( .A1(n9084), .A2(n9032), .ZN(n8887) );
  OAI211_X1 U10343 ( .C1(n9029), .C2(n8888), .A(n8887), .B(n8886), .ZN(
        P2_U3203) );
  NAND2_X1 U10344 ( .A1(n8889), .A2(n9029), .ZN(n8894) );
  NOR2_X1 U10345 ( .A1(n8890), .A2(n9014), .ZN(n8891) );
  AOI211_X1 U10346 ( .C1(n10159), .C2(P2_REG2_REG_29__SCAN_IN), .A(n8892), .B(
        n8891), .ZN(n8893) );
  OAI211_X1 U10347 ( .C1(n8895), .C2(n10155), .A(n8894), .B(n8893), .ZN(
        P2_U3204) );
  XNOR2_X1 U10348 ( .A(n8896), .B(n5766), .ZN(n9097) );
  INV_X1 U10349 ( .A(n9097), .ZN(n8909) );
  OAI21_X1 U10350 ( .B1(n8898), .B2(n8897), .A(n10151), .ZN(n8900) );
  OR2_X1 U10351 ( .A1(n8900), .A2(n8899), .ZN(n8904) );
  AOI22_X1 U10352 ( .A1(n8902), .A2(n10148), .B1(n9025), .B2(n8901), .ZN(n8903) );
  NAND2_X1 U10353 ( .A1(n8904), .A2(n8903), .ZN(n9093) );
  MUX2_X1 U10354 ( .A(n9093), .B(P2_REG2_REG_27__SCAN_IN), .S(n10159), .Z(
        n8905) );
  INV_X1 U10355 ( .A(n8905), .ZN(n8908) );
  AOI22_X1 U10356 ( .A1(n9095), .A2(n9032), .B1(n9031), .B2(n8906), .ZN(n8907)
         );
  OAI211_X1 U10357 ( .C1(n8909), .C2(n9035), .A(n8908), .B(n8907), .ZN(
        P2_U3206) );
  XNOR2_X1 U10358 ( .A(n8911), .B(n8910), .ZN(n9105) );
  XNOR2_X1 U10359 ( .A(n8913), .B(n8912), .ZN(n8915) );
  AOI222_X1 U10360 ( .A1(n10151), .A2(n8915), .B1(n8914), .B2(n10148), .C1(
        n8935), .C2(n9025), .ZN(n9100) );
  MUX2_X1 U10361 ( .A(n8916), .B(n9100), .S(n9029), .Z(n8919) );
  AOI22_X1 U10362 ( .A1(n9102), .A2(n9032), .B1(n9031), .B2(n8917), .ZN(n8918)
         );
  OAI211_X1 U10363 ( .C1(n9105), .C2(n9035), .A(n8919), .B(n8918), .ZN(
        P2_U3207) );
  XNOR2_X1 U10364 ( .A(n8920), .B(n8922), .ZN(n9108) );
  AOI21_X1 U10365 ( .B1(n8922), .B2(n8921), .A(n4554), .ZN(n8923) );
  OAI222_X1 U10366 ( .A1(n9006), .A2(n8925), .B1(n9008), .B2(n8924), .C1(n9003), .C2(n8923), .ZN(n9106) );
  OAI22_X1 U10367 ( .A1(n9107), .A2(n10142), .B1(n8926), .B2(n10141), .ZN(
        n8927) );
  OAI21_X1 U10368 ( .B1(n9106), .B2(n8927), .A(n9029), .ZN(n8929) );
  NAND2_X1 U10369 ( .A1(n10159), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n8928) );
  OAI211_X1 U10370 ( .C1(n9108), .C2(n9035), .A(n8929), .B(n8928), .ZN(
        P2_U3208) );
  NAND2_X1 U10371 ( .A1(n8931), .A2(n8930), .ZN(n8932) );
  XOR2_X1 U10372 ( .A(n8934), .B(n8932), .Z(n9116) );
  XOR2_X1 U10373 ( .A(n8934), .B(n8933), .Z(n8936) );
  AOI222_X1 U10374 ( .A1(n10151), .A2(n8936), .B1(n8958), .B2(n9025), .C1(
        n8935), .C2(n10148), .ZN(n9111) );
  OAI21_X1 U10375 ( .B1(n8937), .B2(n10142), .A(n9111), .ZN(n8938) );
  NAND2_X1 U10376 ( .A1(n8938), .A2(n9029), .ZN(n8941) );
  AOI22_X1 U10377 ( .A1(n8939), .A2(n9031), .B1(n10159), .B2(
        P2_REG2_REG_24__SCAN_IN), .ZN(n8940) );
  OAI211_X1 U10378 ( .C1(n9116), .C2(n9035), .A(n8941), .B(n8940), .ZN(
        P2_U3209) );
  XNOR2_X1 U10379 ( .A(n8942), .B(n8943), .ZN(n9122) );
  XNOR2_X1 U10380 ( .A(n8944), .B(n8943), .ZN(n8946) );
  AOI222_X1 U10381 ( .A1(n10151), .A2(n8946), .B1(n8945), .B2(n10148), .C1(
        n8971), .C2(n9025), .ZN(n9117) );
  MUX2_X1 U10382 ( .A(n8947), .B(n9117), .S(n9029), .Z(n8950) );
  AOI22_X1 U10383 ( .A1(n9119), .A2(n9032), .B1(n9031), .B2(n8948), .ZN(n8949)
         );
  OAI211_X1 U10384 ( .C1(n9122), .C2(n9035), .A(n8950), .B(n8949), .ZN(
        P2_U3210) );
  XOR2_X1 U10385 ( .A(n8953), .B(n8951), .Z(n9128) );
  INV_X1 U10386 ( .A(n8953), .ZN(n8955) );
  NAND3_X1 U10387 ( .A1(n8952), .A2(n8955), .A3(n8954), .ZN(n8956) );
  NAND2_X1 U10388 ( .A1(n8957), .A2(n8956), .ZN(n8959) );
  AOI222_X1 U10389 ( .A1(n10151), .A2(n8959), .B1(n8958), .B2(n10148), .C1(
        n8982), .C2(n9025), .ZN(n9123) );
  MUX2_X1 U10390 ( .A(n8960), .B(n9123), .S(n9029), .Z(n8963) );
  AOI22_X1 U10391 ( .A1(n9125), .A2(n9032), .B1(n9031), .B2(n8961), .ZN(n8962)
         );
  OAI211_X1 U10392 ( .C1(n9128), .C2(n9035), .A(n8963), .B(n8962), .ZN(
        P2_U3211) );
  NAND2_X1 U10393 ( .A1(n8964), .A2(n8965), .ZN(n8966) );
  XNOR2_X1 U10394 ( .A(n8966), .B(n8968), .ZN(n9134) );
  NAND3_X1 U10395 ( .A1(n8967), .A2(n4892), .A3(n8969), .ZN(n8970) );
  NAND2_X1 U10396 ( .A1(n8952), .A2(n8970), .ZN(n8973) );
  AOI222_X1 U10397 ( .A1(n10151), .A2(n8973), .B1(n8972), .B2(n9025), .C1(
        n8971), .C2(n10148), .ZN(n9129) );
  MUX2_X1 U10398 ( .A(n8974), .B(n9129), .S(n9029), .Z(n8977) );
  AOI22_X1 U10399 ( .A1(n9131), .A2(n9032), .B1(n9031), .B2(n8975), .ZN(n8976)
         );
  OAI211_X1 U10400 ( .C1(n9134), .C2(n9035), .A(n8977), .B(n8976), .ZN(
        P2_U3212) );
  XNOR2_X1 U10401 ( .A(n8978), .B(n8979), .ZN(n9140) );
  INV_X1 U10402 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n8984) );
  OAI21_X1 U10403 ( .B1(n8980), .B2(n5639), .A(n8967), .ZN(n8983) );
  AOI222_X1 U10404 ( .A1(n10151), .A2(n8983), .B1(n8982), .B2(n10148), .C1(
        n8981), .C2(n9025), .ZN(n9135) );
  MUX2_X1 U10405 ( .A(n8984), .B(n9135), .S(n9029), .Z(n8987) );
  AOI22_X1 U10406 ( .A1(n9137), .A2(n9032), .B1(n9031), .B2(n8985), .ZN(n8986)
         );
  OAI211_X1 U10407 ( .C1(n9140), .C2(n9035), .A(n8987), .B(n8986), .ZN(
        P2_U3213) );
  OAI21_X1 U10408 ( .B1(n8990), .B2(n8989), .A(n8988), .ZN(n9144) );
  XNOR2_X1 U10409 ( .A(n8992), .B(n8991), .ZN(n8993) );
  OAI222_X1 U10410 ( .A1(n9008), .A2(n8995), .B1(n9006), .B2(n8994), .C1(n8993), .C2(n9003), .ZN(n9066) );
  NAND2_X1 U10411 ( .A1(n9066), .A2(n9029), .ZN(n9001) );
  INV_X1 U10412 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n8998) );
  INV_X1 U10413 ( .A(n8996), .ZN(n8997) );
  OAI22_X1 U10414 ( .A1(n9029), .A2(n8998), .B1(n8997), .B2(n10141), .ZN(n8999) );
  AOI21_X1 U10415 ( .B1(n9067), .B2(n9032), .A(n8999), .ZN(n9000) );
  OAI211_X1 U10416 ( .C1(n9144), .C2(n9035), .A(n9001), .B(n9000), .ZN(
        P2_U3214) );
  XNOR2_X1 U10417 ( .A(n9002), .B(n9009), .ZN(n9004) );
  OAI222_X1 U10418 ( .A1(n9008), .A2(n9007), .B1(n9006), .B2(n9005), .C1(n9004), .C2(n9003), .ZN(n9071) );
  INV_X1 U10419 ( .A(n9072), .ZN(n9011) );
  AND2_X1 U10420 ( .A1(n9010), .A2(n9009), .ZN(n9070) );
  NOR3_X1 U10421 ( .A1(n9011), .A2(n9070), .A3(n9035), .ZN(n9016) );
  AOI22_X1 U10422 ( .A1(n10159), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n9031), 
        .B2(n9012), .ZN(n9013) );
  OAI21_X1 U10423 ( .B1(n9149), .B2(n9014), .A(n9013), .ZN(n9015) );
  AOI211_X1 U10424 ( .C1(n9071), .C2(n9029), .A(n9016), .B(n9015), .ZN(n9017)
         );
  INV_X1 U10425 ( .A(n9017), .ZN(P2_U3215) );
  XNOR2_X1 U10426 ( .A(n9019), .B(n9018), .ZN(n9157) );
  NAND3_X1 U10427 ( .A1(n9021), .A2(n4721), .A3(n9020), .ZN(n9022) );
  NAND3_X1 U10428 ( .A1(n9023), .A2(n10151), .A3(n9022), .ZN(n9028) );
  AOI22_X1 U10429 ( .A1(n9026), .A2(n9025), .B1(n10148), .B2(n9024), .ZN(n9027) );
  MUX2_X1 U10430 ( .A(n8807), .B(n9150), .S(n9029), .Z(n9034) );
  AOI22_X1 U10431 ( .A1(n9153), .A2(n9032), .B1(n9031), .B2(n9030), .ZN(n9033)
         );
  OAI211_X1 U10432 ( .C1(n9157), .C2(n9035), .A(n9034), .B(n9033), .ZN(
        P2_U3216) );
  NAND2_X1 U10433 ( .A1(n9081), .A2(n6647), .ZN(n9036) );
  NAND2_X1 U10434 ( .A1(n9082), .A2(n10213), .ZN(n9037) );
  OAI211_X1 U10435 ( .C1(n10213), .C2(n7531), .A(n9036), .B(n9037), .ZN(
        P2_U3490) );
  INV_X1 U10436 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n9039) );
  NAND2_X1 U10437 ( .A1(n9084), .A2(n6647), .ZN(n9038) );
  OAI211_X1 U10438 ( .C1(n10213), .C2(n9039), .A(n9038), .B(n9037), .ZN(
        P2_U3489) );
  MUX2_X1 U10439 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n9088), .S(n10213), .Z(
        n9041) );
  OAI22_X1 U10440 ( .A1(n9090), .A2(n9080), .B1(n9089), .B2(n9076), .ZN(n9040)
         );
  MUX2_X1 U10441 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n9093), .S(n10213), .Z(
        n9042) );
  INV_X1 U10442 ( .A(n9042), .ZN(n9045) );
  AOI22_X1 U10443 ( .A1(n9097), .A2(n9043), .B1(n6647), .B2(n9095), .ZN(n9044)
         );
  NAND2_X1 U10444 ( .A1(n9045), .A2(n9044), .ZN(P2_U3486) );
  INV_X1 U10445 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n9046) );
  MUX2_X1 U10446 ( .A(n9046), .B(n9100), .S(n10213), .Z(n9048) );
  NAND2_X1 U10447 ( .A1(n9102), .A2(n6647), .ZN(n9047) );
  OAI211_X1 U10448 ( .C1(n9105), .C2(n9080), .A(n9048), .B(n9047), .ZN(
        P2_U3485) );
  MUX2_X1 U10449 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n9106), .S(n10213), .Z(
        n9050) );
  OAI22_X1 U10450 ( .A1(n9108), .A2(n9080), .B1(n9107), .B2(n9076), .ZN(n9049)
         );
  OR2_X1 U10451 ( .A1(n9050), .A2(n9049), .ZN(P2_U3484) );
  INV_X1 U10452 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n9051) );
  MUX2_X1 U10453 ( .A(n9051), .B(n9111), .S(n10213), .Z(n9053) );
  NAND2_X1 U10454 ( .A1(n9113), .A2(n6647), .ZN(n9052) );
  OAI211_X1 U10455 ( .C1(n9080), .C2(n9116), .A(n9053), .B(n9052), .ZN(
        P2_U3483) );
  INV_X1 U10456 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n9054) );
  MUX2_X1 U10457 ( .A(n9054), .B(n9117), .S(n10213), .Z(n9056) );
  NAND2_X1 U10458 ( .A1(n9119), .A2(n6647), .ZN(n9055) );
  OAI211_X1 U10459 ( .C1(n9122), .C2(n9080), .A(n9056), .B(n9055), .ZN(
        P2_U3482) );
  INV_X1 U10460 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n9057) );
  MUX2_X1 U10461 ( .A(n9057), .B(n9123), .S(n10213), .Z(n9059) );
  NAND2_X1 U10462 ( .A1(n9125), .A2(n6647), .ZN(n9058) );
  OAI211_X1 U10463 ( .C1(n9128), .C2(n9080), .A(n9059), .B(n9058), .ZN(
        P2_U3481) );
  INV_X1 U10464 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n9060) );
  MUX2_X1 U10465 ( .A(n9060), .B(n9129), .S(n10213), .Z(n9062) );
  NAND2_X1 U10466 ( .A1(n9131), .A2(n6647), .ZN(n9061) );
  OAI211_X1 U10467 ( .C1(n9080), .C2(n9134), .A(n9062), .B(n9061), .ZN(
        P2_U3480) );
  INV_X1 U10468 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n9063) );
  MUX2_X1 U10469 ( .A(n9063), .B(n9135), .S(n10213), .Z(n9065) );
  NAND2_X1 U10470 ( .A1(n9137), .A2(n6647), .ZN(n9064) );
  OAI211_X1 U10471 ( .C1(n9140), .C2(n9080), .A(n9065), .B(n9064), .ZN(
        P2_U3479) );
  INV_X1 U10472 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n9068) );
  AOI21_X1 U10473 ( .B1(n10198), .B2(n9067), .A(n9066), .ZN(n9141) );
  MUX2_X1 U10474 ( .A(n9068), .B(n9141), .S(n10213), .Z(n9069) );
  OAI21_X1 U10475 ( .B1(n9080), .B2(n9144), .A(n9069), .ZN(P2_U3478) );
  NOR2_X1 U10476 ( .A1(n9070), .A2(n10193), .ZN(n9073) );
  AOI21_X1 U10477 ( .B1(n9073), .B2(n9072), .A(n9071), .ZN(n9145) );
  MUX2_X1 U10478 ( .A(n9074), .B(n9145), .S(n10213), .Z(n9075) );
  OAI21_X1 U10479 ( .B1(n9149), .B2(n9076), .A(n9075), .ZN(P2_U3477) );
  MUX2_X1 U10480 ( .A(n9077), .B(n9150), .S(n10213), .Z(n9079) );
  NAND2_X1 U10481 ( .A1(n9153), .A2(n6647), .ZN(n9078) );
  OAI211_X1 U10482 ( .C1(n9080), .C2(n9157), .A(n9079), .B(n9078), .ZN(
        P2_U3476) );
  NAND2_X1 U10483 ( .A1(n9081), .A2(n9152), .ZN(n9083) );
  NAND2_X1 U10484 ( .A1(n9082), .A2(n10199), .ZN(n9085) );
  OAI211_X1 U10485 ( .C1(n7529), .C2(n10199), .A(n9083), .B(n9085), .ZN(
        P2_U3458) );
  INV_X1 U10486 ( .A(n9084), .ZN(n9087) );
  NAND2_X1 U10487 ( .A1(n10201), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n9086) );
  OAI211_X1 U10488 ( .C1(n9087), .C2(n9148), .A(n9086), .B(n9085), .ZN(
        P2_U3457) );
  OAI22_X1 U10489 ( .A1(n9090), .A2(n9156), .B1(n9089), .B2(n9148), .ZN(n9091)
         );
  OR2_X1 U10490 ( .A1(n9092), .A2(n9091), .ZN(P2_U3455) );
  MUX2_X1 U10491 ( .A(n9093), .B(P2_REG0_REG_27__SCAN_IN), .S(n10201), .Z(
        n9094) );
  INV_X1 U10492 ( .A(n9094), .ZN(n9099) );
  AOI22_X1 U10493 ( .A1(n9097), .A2(n9096), .B1(n9152), .B2(n9095), .ZN(n9098)
         );
  NAND2_X1 U10494 ( .A1(n9099), .A2(n9098), .ZN(P2_U3454) );
  INV_X1 U10495 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n9101) );
  MUX2_X1 U10496 ( .A(n9101), .B(n9100), .S(n10199), .Z(n9104) );
  NAND2_X1 U10497 ( .A1(n9102), .A2(n9152), .ZN(n9103) );
  OAI211_X1 U10498 ( .C1(n9105), .C2(n9156), .A(n9104), .B(n9103), .ZN(
        P2_U3453) );
  MUX2_X1 U10499 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n9106), .S(n10199), .Z(
        n9110) );
  OAI22_X1 U10500 ( .A1(n9108), .A2(n9156), .B1(n9107), .B2(n9148), .ZN(n9109)
         );
  OR2_X1 U10501 ( .A1(n9110), .A2(n9109), .ZN(P2_U3452) );
  INV_X1 U10502 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n9112) );
  MUX2_X1 U10503 ( .A(n9112), .B(n9111), .S(n10199), .Z(n9115) );
  NAND2_X1 U10504 ( .A1(n9113), .A2(n9152), .ZN(n9114) );
  OAI211_X1 U10505 ( .C1(n9116), .C2(n9156), .A(n9115), .B(n9114), .ZN(
        P2_U3451) );
  INV_X1 U10506 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n9118) );
  MUX2_X1 U10507 ( .A(n9118), .B(n9117), .S(n10199), .Z(n9121) );
  NAND2_X1 U10508 ( .A1(n9119), .A2(n9152), .ZN(n9120) );
  OAI211_X1 U10509 ( .C1(n9122), .C2(n9156), .A(n9121), .B(n9120), .ZN(
        P2_U3450) );
  INV_X1 U10510 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n9124) );
  MUX2_X1 U10511 ( .A(n9124), .B(n9123), .S(n10199), .Z(n9127) );
  NAND2_X1 U10512 ( .A1(n9125), .A2(n9152), .ZN(n9126) );
  OAI211_X1 U10513 ( .C1(n9128), .C2(n9156), .A(n9127), .B(n9126), .ZN(
        P2_U3449) );
  INV_X1 U10514 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n9130) );
  MUX2_X1 U10515 ( .A(n9130), .B(n9129), .S(n10199), .Z(n9133) );
  NAND2_X1 U10516 ( .A1(n9131), .A2(n9152), .ZN(n9132) );
  OAI211_X1 U10517 ( .C1(n9134), .C2(n9156), .A(n9133), .B(n9132), .ZN(
        P2_U3448) );
  INV_X1 U10518 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n9136) );
  MUX2_X1 U10519 ( .A(n9136), .B(n9135), .S(n10199), .Z(n9139) );
  NAND2_X1 U10520 ( .A1(n9137), .A2(n9152), .ZN(n9138) );
  OAI211_X1 U10521 ( .C1(n9140), .C2(n9156), .A(n9139), .B(n9138), .ZN(
        P2_U3447) );
  INV_X1 U10522 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n9142) );
  MUX2_X1 U10523 ( .A(n9142), .B(n9141), .S(n10199), .Z(n9143) );
  OAI21_X1 U10524 ( .B1(n9144), .B2(n9156), .A(n9143), .ZN(P2_U3446) );
  INV_X1 U10525 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n9146) );
  MUX2_X1 U10526 ( .A(n9146), .B(n9145), .S(n10199), .Z(n9147) );
  OAI21_X1 U10527 ( .B1(n9149), .B2(n9148), .A(n9147), .ZN(P2_U3444) );
  INV_X1 U10528 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n9151) );
  MUX2_X1 U10529 ( .A(n9151), .B(n9150), .S(n10199), .Z(n9155) );
  NAND2_X1 U10530 ( .A1(n9153), .A2(n9152), .ZN(n9154) );
  OAI211_X1 U10531 ( .C1(n9157), .C2(n9156), .A(n9155), .B(n9154), .ZN(
        P2_U3441) );
  AND2_X1 U10532 ( .A1(n9159), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9162) );
  NAND4_X1 U10533 ( .A1(n9162), .A2(P2_IR_REG_31__SCAN_IN), .A3(n9161), .A4(
        n9160), .ZN(n9164) );
  OAI22_X1 U10534 ( .A1(n9158), .A2(n9164), .B1(n9163), .B2(n8539), .ZN(n9165)
         );
  AOI21_X1 U10535 ( .B1(n9895), .B2(n9166), .A(n9165), .ZN(n9167) );
  INV_X1 U10536 ( .A(n9167), .ZN(P2_U3264) );
  CLKBUF_X1 U10537 ( .A(n9168), .Z(n9169) );
  INV_X1 U10538 ( .A(n9170), .ZN(n9902) );
  OAI222_X1 U10539 ( .A1(n8539), .A2(n9173), .B1(P2_U3151), .B2(n9169), .C1(
        n9902), .C2(n9171), .ZN(P2_U3266) );
  AOI21_X1 U10540 ( .B1(n9176), .B2(n9175), .A(n4583), .ZN(n9184) );
  OR2_X1 U10541 ( .A1(n9177), .A2(n9537), .ZN(n9179) );
  OR2_X1 U10542 ( .A1(n9269), .A2(n9338), .ZN(n9178) );
  NAND2_X1 U10543 ( .A1(n9179), .A2(n9178), .ZN(n9749) );
  NAND2_X1 U10544 ( .A1(n9749), .A2(n4510), .ZN(n9181) );
  OAI211_X1 U10545 ( .C1(n9920), .C2(n9756), .A(n9181), .B(n9180), .ZN(n9182)
         );
  AOI21_X1 U10546 ( .B1(n10073), .B2(n9395), .A(n9182), .ZN(n9183) );
  OAI21_X1 U10547 ( .B1(n9184), .B2(n9916), .A(n9183), .ZN(P1_U3215) );
  AOI21_X1 U10548 ( .B1(n9186), .B2(n9185), .A(n4545), .ZN(n9193) );
  OR2_X1 U10549 ( .A1(n9256), .A2(n9338), .ZN(n9188) );
  NAND2_X1 U10550 ( .A1(n9403), .A2(n9199), .ZN(n9187) );
  NAND2_X1 U10551 ( .A1(n9188), .A2(n9187), .ZN(n9792) );
  INV_X1 U10552 ( .A(n9920), .ZN(n9219) );
  INV_X1 U10553 ( .A(n9219), .ZN(n9951) );
  OAI22_X1 U10554 ( .A1(n9639), .A2(n9951), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9189), .ZN(n9190) );
  AOI21_X1 U10555 ( .B1(n9792), .B2(n4510), .A(n9190), .ZN(n9192) );
  NAND2_X1 U10556 ( .A1(n9791), .A2(n9395), .ZN(n9191) );
  OAI211_X1 U10557 ( .C1(n9193), .C2(n9916), .A(n9192), .B(n9191), .ZN(
        P1_U3216) );
  NAND2_X1 U10558 ( .A1(n9365), .A2(n9194), .ZN(n9360) );
  NAND2_X1 U10559 ( .A1(n4541), .A2(n9195), .ZN(n9362) );
  NAND2_X1 U10560 ( .A1(n9360), .A2(n9362), .ZN(n9359) );
  XOR2_X1 U10561 ( .A(n9197), .B(n9196), .Z(n9198) );
  XNOR2_X1 U10562 ( .A(n9359), .B(n9198), .ZN(n9205) );
  OR2_X1 U10563 ( .A1(n9232), .A2(n9338), .ZN(n9201) );
  NAND2_X1 U10564 ( .A1(n9407), .A2(n9199), .ZN(n9200) );
  NAND2_X1 U10565 ( .A1(n9201), .A2(n9200), .ZN(n9704) );
  AOI22_X1 U10566 ( .A1(n9704), .A2(n4510), .B1(P1_REG3_REG_19__SCAN_IN), .B2(
        P1_U3086), .ZN(n9202) );
  OAI21_X1 U10567 ( .B1(n9698), .B2(n9920), .A(n9202), .ZN(n9203) );
  AOI21_X1 U10568 ( .B1(n9815), .B2(n9395), .A(n9203), .ZN(n9204) );
  OAI21_X1 U10569 ( .B1(n9205), .B2(n9916), .A(n9204), .ZN(P1_U3219) );
  NAND2_X1 U10570 ( .A1(n9556), .A2(n9206), .ZN(n9209) );
  OR2_X1 U10571 ( .A1(n9538), .A2(n9207), .ZN(n9208) );
  NAND2_X1 U10572 ( .A1(n9209), .A2(n9208), .ZN(n9211) );
  XNOR2_X1 U10573 ( .A(n9211), .B(n9210), .ZN(n9216) );
  NAND2_X1 U10574 ( .A1(n9556), .A2(n9212), .ZN(n9213) );
  OAI21_X1 U10575 ( .B1(n9538), .B2(n9214), .A(n9213), .ZN(n9215) );
  XNOR2_X1 U10576 ( .A(n9216), .B(n9215), .ZN(n9225) );
  OR4_X2 U10577 ( .A1(n9218), .A2(n9224), .A3(n9225), .A4(n9916), .ZN(n9229)
         );
  AOI22_X1 U10578 ( .A1(n9555), .A2(n9219), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3086), .ZN(n9220) );
  OAI21_X1 U10579 ( .B1(n9222), .B2(n9221), .A(n9220), .ZN(n9223) );
  AOI21_X1 U10580 ( .B1(n9556), .B2(n9395), .A(n9223), .ZN(n9227) );
  NAND3_X1 U10581 ( .A1(n9225), .A2(n9948), .A3(n9224), .ZN(n9226) );
  NAND4_X1 U10582 ( .A1(n9229), .A2(n9228), .A3(n9227), .A4(n9226), .ZN(
        P1_U3220) );
  XNOR2_X1 U10583 ( .A(n9231), .B(n9230), .ZN(n9237) );
  OAI22_X1 U10584 ( .A1(n9233), .A2(n9338), .B1(n9232), .B2(n9537), .ZN(n9667)
         );
  AOI22_X1 U10585 ( .A1(n9667), .A2(n4510), .B1(P1_REG3_REG_21__SCAN_IN), .B2(
        P1_U3086), .ZN(n9234) );
  OAI21_X1 U10586 ( .B1(n9672), .B2(n9920), .A(n9234), .ZN(n9235) );
  AOI21_X1 U10587 ( .B1(n9671), .B2(n9395), .A(n9235), .ZN(n9236) );
  OAI21_X1 U10588 ( .B1(n9237), .B2(n9916), .A(n9236), .ZN(P1_U3223) );
  INV_X1 U10589 ( .A(n9238), .ZN(n9349) );
  INV_X1 U10590 ( .A(n9239), .ZN(n9241) );
  NOR3_X1 U10591 ( .A1(n9349), .A2(n9241), .A3(n9240), .ZN(n9244) );
  INV_X1 U10592 ( .A(n9242), .ZN(n9243) );
  OAI21_X1 U10593 ( .B1(n9244), .B2(n9243), .A(n9948), .ZN(n9250) );
  NOR2_X1 U10594 ( .A1(n9920), .A2(n9245), .ZN(n9246) );
  AOI211_X1 U10595 ( .C1(n4510), .C2(n9248), .A(n9247), .B(n9246), .ZN(n9249)
         );
  OAI211_X1 U10596 ( .C1(n9251), .C2(n9946), .A(n9250), .B(n9249), .ZN(
        P1_U3224) );
  OAI21_X1 U10597 ( .B1(n9254), .B2(n9252), .A(n9253), .ZN(n9255) );
  NAND2_X1 U10598 ( .A1(n9255), .A2(n9948), .ZN(n9262) );
  OAI22_X1 U10599 ( .A1(n9257), .A2(n9338), .B1(n9256), .B2(n9537), .ZN(n9605)
         );
  INV_X1 U10600 ( .A(n9608), .ZN(n9259) );
  OAI22_X1 U10601 ( .A1(n9259), .A2(n9920), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9258), .ZN(n9260) );
  AOI21_X1 U10602 ( .B1(n9605), .B2(n4510), .A(n9260), .ZN(n9261) );
  OAI211_X1 U10603 ( .C1(n9861), .C2(n9946), .A(n9262), .B(n9261), .ZN(
        P1_U3225) );
  INV_X1 U10604 ( .A(n9263), .ZN(n9268) );
  AOI21_X1 U10605 ( .B1(n9267), .B2(n9265), .A(n9264), .ZN(n9266) );
  AOI21_X1 U10606 ( .B1(n9268), .B2(n9267), .A(n9266), .ZN(n9274) );
  OAI22_X1 U10607 ( .A1(n9269), .A2(n9537), .B1(n9367), .B2(n9338), .ZN(n9836)
         );
  NAND2_X1 U10608 ( .A1(n9836), .A2(n4510), .ZN(n9271) );
  OAI211_X1 U10609 ( .C1(n9920), .C2(n9923), .A(n9271), .B(n9270), .ZN(n9272)
         );
  AOI21_X1 U10610 ( .B1(n9833), .B2(n9395), .A(n9272), .ZN(n9273) );
  OAI21_X1 U10611 ( .B1(n9274), .B2(n9916), .A(n9273), .ZN(P1_U3226) );
  OAI21_X1 U10612 ( .B1(n9277), .B2(n9276), .A(n9275), .ZN(n9278) );
  NAND2_X1 U10613 ( .A1(n9278), .A2(n9948), .ZN(n9284) );
  OR2_X1 U10614 ( .A1(n9279), .A2(n9537), .ZN(n9280) );
  OAI21_X1 U10615 ( .B1(n9281), .B2(n9338), .A(n9280), .ZN(n9731) );
  AND2_X1 U10616 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n9495) );
  NOR2_X1 U10617 ( .A1(n9920), .A2(n9740), .ZN(n9282) );
  AOI211_X1 U10618 ( .C1(n4510), .C2(n9731), .A(n9495), .B(n9282), .ZN(n9283)
         );
  OAI211_X1 U10619 ( .C1(n6494), .C2(n9946), .A(n9284), .B(n9283), .ZN(
        P1_U3228) );
  INV_X1 U10620 ( .A(n9625), .ZN(n9865) );
  INV_X1 U10621 ( .A(n9285), .ZN(n9289) );
  NOR3_X1 U10622 ( .A1(n4545), .A2(n9287), .A3(n9286), .ZN(n9288) );
  OAI21_X1 U10623 ( .B1(n9289), .B2(n9288), .A(n9948), .ZN(n9295) );
  OAI22_X1 U10624 ( .A1(n9290), .A2(n9338), .B1(n9339), .B2(n9537), .ZN(n9620)
         );
  INV_X1 U10625 ( .A(n9626), .ZN(n9292) );
  OAI22_X1 U10626 ( .A1(n9292), .A2(n9951), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9291), .ZN(n9293) );
  AOI21_X1 U10627 ( .B1(n9620), .B2(n4510), .A(n9293), .ZN(n9294) );
  OAI211_X1 U10628 ( .C1(n9865), .C2(n9946), .A(n9295), .B(n9294), .ZN(
        P1_U3229) );
  AND2_X1 U10629 ( .A1(n9297), .A2(n9298), .ZN(n9301) );
  OAI211_X1 U10630 ( .C1(n9301), .C2(n9300), .A(n9948), .B(n9299), .ZN(n9311)
         );
  NAND2_X1 U10631 ( .A1(n9303), .A2(n9302), .ZN(n9305) );
  AOI21_X1 U10632 ( .B1(n9305), .B2(n4510), .A(n9304), .ZN(n9310) );
  NAND2_X1 U10633 ( .A1(n9306), .A2(n9395), .ZN(n9309) );
  OR2_X1 U10634 ( .A1(n9920), .A2(n9307), .ZN(n9308) );
  NAND4_X1 U10635 ( .A1(n9311), .A2(n9310), .A3(n9309), .A4(n9308), .ZN(
        P1_U3231) );
  XNOR2_X1 U10636 ( .A(n9313), .B(n9312), .ZN(n9314) );
  XNOR2_X1 U10637 ( .A(n9315), .B(n9314), .ZN(n9321) );
  INV_X1 U10638 ( .A(n9689), .ZN(n9318) );
  OAI22_X1 U10639 ( .A1(n9337), .A2(n9338), .B1(n9316), .B2(n9537), .ZN(n9683)
         );
  AOI22_X1 U10640 ( .A1(n9683), .A2(n4510), .B1(P1_REG3_REG_20__SCAN_IN), .B2(
        P1_U3086), .ZN(n9317) );
  OAI21_X1 U10641 ( .B1(n9318), .B2(n9920), .A(n9317), .ZN(n9319) );
  AOI21_X1 U10642 ( .B1(n9688), .B2(n9395), .A(n9319), .ZN(n9320) );
  OAI21_X1 U10643 ( .B1(n9321), .B2(n9916), .A(n9320), .ZN(P1_U3233) );
  OAI21_X1 U10644 ( .B1(n9324), .B2(n9322), .A(n9323), .ZN(n9325) );
  NAND2_X1 U10645 ( .A1(n9325), .A2(n9948), .ZN(n9332) );
  INV_X1 U10646 ( .A(n9326), .ZN(n9329) );
  NOR2_X1 U10647 ( .A1(n9951), .A2(n9327), .ZN(n9328) );
  AOI211_X1 U10648 ( .C1(n4510), .C2(n9330), .A(n9329), .B(n9328), .ZN(n9331)
         );
  OAI211_X1 U10649 ( .C1(n4762), .C2(n9946), .A(n9332), .B(n9331), .ZN(
        P1_U3234) );
  XNOR2_X1 U10650 ( .A(n9334), .B(n9333), .ZN(n9335) );
  XNOR2_X1 U10651 ( .A(n9336), .B(n9335), .ZN(n9345) );
  OAI22_X1 U10652 ( .A1(n9339), .A2(n9338), .B1(n9337), .B2(n9537), .ZN(n9657)
         );
  INV_X1 U10653 ( .A(n9652), .ZN(n9341) );
  OAI22_X1 U10654 ( .A1(n9341), .A2(n9951), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9340), .ZN(n9343) );
  NOR2_X1 U10655 ( .A1(n9654), .A2(n9946), .ZN(n9342) );
  AOI211_X1 U10656 ( .C1(n4510), .C2(n9657), .A(n9343), .B(n9342), .ZN(n9344)
         );
  OAI21_X1 U10657 ( .B1(n9345), .B2(n9916), .A(n9344), .ZN(P1_U3235) );
  INV_X1 U10658 ( .A(n9346), .ZN(n9348) );
  NOR3_X1 U10659 ( .A1(n4580), .A2(n9348), .A3(n9347), .ZN(n9350) );
  OAI21_X1 U10660 ( .B1(n9350), .B2(n9349), .A(n9948), .ZN(n9357) );
  INV_X1 U10661 ( .A(n9351), .ZN(n9354) );
  NOR2_X1 U10662 ( .A1(n9951), .A2(n9352), .ZN(n9353) );
  AOI211_X1 U10663 ( .C1(n4510), .C2(n9355), .A(n9354), .B(n9353), .ZN(n9356)
         );
  OAI211_X1 U10664 ( .C1(n9358), .C2(n9946), .A(n9357), .B(n9356), .ZN(
        P1_U3236) );
  INV_X1 U10665 ( .A(n9359), .ZN(n9366) );
  INV_X1 U10666 ( .A(n9360), .ZN(n9363) );
  AOI21_X1 U10667 ( .B1(n9363), .B2(n9362), .A(n9361), .ZN(n9364) );
  AOI21_X1 U10668 ( .B1(n9366), .B2(n9365), .A(n9364), .ZN(n9374) );
  OR2_X1 U10669 ( .A1(n9367), .A2(n9537), .ZN(n9370) );
  NAND2_X1 U10670 ( .A1(n9406), .A2(n9368), .ZN(n9369) );
  NAND2_X1 U10671 ( .A1(n9370), .A2(n9369), .ZN(n9715) );
  AOI22_X1 U10672 ( .A1(n9715), .A2(n4510), .B1(P1_REG3_REG_18__SCAN_IN), .B2(
        P1_U3086), .ZN(n9371) );
  OAI21_X1 U10673 ( .B1(n9720), .B2(n9920), .A(n9371), .ZN(n9372) );
  AOI21_X1 U10674 ( .B1(n9719), .B2(n9395), .A(n9372), .ZN(n9373) );
  OAI21_X1 U10675 ( .B1(n9374), .B2(n9916), .A(n9373), .ZN(P1_U3238) );
  NAND2_X1 U10676 ( .A1(n5148), .A2(n9375), .ZN(n9379) );
  OAI21_X1 U10677 ( .B1(n9377), .B2(n7515), .A(n9376), .ZN(n9378) );
  XOR2_X1 U10678 ( .A(n9379), .B(n9378), .Z(n9380) );
  NAND2_X1 U10679 ( .A1(n9380), .A2(n9948), .ZN(n9386) );
  AOI22_X1 U10680 ( .A1(n9381), .A2(n4510), .B1(P1_REG3_REG_6__SCAN_IN), .B2(
        P1_U3086), .ZN(n9385) );
  OR2_X1 U10681 ( .A1(n9920), .A2(n9382), .ZN(n9384) );
  OR2_X1 U10682 ( .A1(n9946), .A2(n10039), .ZN(n9383) );
  NAND4_X1 U10683 ( .A1(n9386), .A2(n9385), .A3(n9384), .A4(n9383), .ZN(
        P1_U3239) );
  NAND2_X1 U10684 ( .A1(n9388), .A2(n9387), .ZN(n9389) );
  XOR2_X1 U10685 ( .A(n9390), .B(n9389), .Z(n9398) );
  AOI22_X1 U10686 ( .A1(n9391), .A2(n4510), .B1(P1_REG3_REG_15__SCAN_IN), .B2(
        P1_U3086), .ZN(n9392) );
  OAI21_X1 U10687 ( .B1(n9393), .B2(n9920), .A(n9392), .ZN(n9394) );
  AOI21_X1 U10688 ( .B1(n9396), .B2(n9395), .A(n9394), .ZN(n9397) );
  OAI21_X1 U10689 ( .B1(n9398), .B2(n9916), .A(n9397), .ZN(P1_U3241) );
  MUX2_X1 U10690 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n9399), .S(n4511), .Z(
        P1_U3583) );
  INV_X1 U10691 ( .A(n9538), .ZN(n9541) );
  MUX2_X1 U10692 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n9541), .S(n4511), .Z(
        P1_U3582) );
  MUX2_X1 U10693 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n9400), .S(n4511), .Z(
        P1_U3580) );
  MUX2_X1 U10694 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n9401), .S(P1_U3973), .Z(
        P1_U3579) );
  MUX2_X1 U10695 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n4749), .S(P1_U3973), .Z(
        P1_U3578) );
  MUX2_X1 U10696 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n9402), .S(P1_U3973), .Z(
        P1_U3577) );
  MUX2_X1 U10697 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n9403), .S(P1_U3973), .Z(
        P1_U3576) );
  MUX2_X1 U10698 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n9404), .S(P1_U3973), .Z(
        P1_U3575) );
  MUX2_X1 U10699 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n9405), .S(P1_U3973), .Z(
        P1_U3574) );
  MUX2_X1 U10700 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n9406), .S(n4511), .Z(
        P1_U3573) );
  MUX2_X1 U10701 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n9407), .S(n4511), .Z(
        P1_U3572) );
  MUX2_X1 U10702 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n9408), .S(n4511), .Z(
        P1_U3571) );
  MUX2_X1 U10703 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n9409), .S(n4511), .Z(
        P1_U3570) );
  MUX2_X1 U10704 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n9410), .S(n4511), .Z(
        P1_U3569) );
  MUX2_X1 U10705 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n9411), .S(n4511), .Z(
        P1_U3568) );
  MUX2_X1 U10706 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n9412), .S(n4511), .Z(
        P1_U3567) );
  MUX2_X1 U10707 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n9413), .S(n4511), .Z(
        P1_U3566) );
  MUX2_X1 U10708 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n9414), .S(n4511), .Z(
        P1_U3565) );
  MUX2_X1 U10709 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n9415), .S(n4511), .Z(
        P1_U3564) );
  MUX2_X1 U10710 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n9416), .S(n4511), .Z(
        P1_U3563) );
  MUX2_X1 U10711 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n9417), .S(n4511), .Z(
        P1_U3562) );
  MUX2_X1 U10712 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n9418), .S(n4511), .Z(
        P1_U3561) );
  MUX2_X1 U10713 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n9419), .S(n4511), .Z(
        P1_U3560) );
  MUX2_X1 U10714 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n9420), .S(n4511), .Z(
        P1_U3559) );
  MUX2_X1 U10715 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n9421), .S(n4511), .Z(
        P1_U3557) );
  MUX2_X1 U10716 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n5914), .S(n4511), .Z(
        P1_U3555) );
  MUX2_X1 U10717 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(n5927), .S(n4511), .Z(
        P1_U3554) );
  OAI211_X1 U10718 ( .C1(n9424), .C2(n9423), .A(n9499), .B(n9422), .ZN(n9432)
         );
  AOI22_X1 U10719 ( .A1(n9956), .A2(P1_ADDR_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(P1_U3086), .ZN(n9431) );
  NAND2_X1 U10720 ( .A1(n9516), .A2(n9425), .ZN(n9430) );
  OAI211_X1 U10721 ( .C1(n9428), .C2(n9427), .A(n9517), .B(n9426), .ZN(n9429)
         );
  NAND4_X1 U10722 ( .A1(n9432), .A2(n9431), .A3(n9430), .A4(n9429), .ZN(
        P1_U3244) );
  INV_X1 U10723 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n9434) );
  OAI22_X1 U10724 ( .A1(n9507), .A2(n9434), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9433), .ZN(n9435) );
  AOI21_X1 U10725 ( .B1(n9436), .B2(n9516), .A(n9435), .ZN(n9446) );
  OAI21_X1 U10726 ( .B1(n9439), .B2(n9438), .A(n9437), .ZN(n9440) );
  OR2_X1 U10727 ( .A1(n9510), .A2(n9440), .ZN(n9445) );
  OAI211_X1 U10728 ( .C1(n9443), .C2(n9442), .A(n9517), .B(n9441), .ZN(n9444)
         );
  NAND4_X1 U10729 ( .A1(n9447), .A2(n9446), .A3(n9445), .A4(n9444), .ZN(
        P1_U3245) );
  INV_X1 U10730 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n9449) );
  NAND2_X1 U10731 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_U3086), .ZN(n9448) );
  OAI21_X1 U10732 ( .B1(n9507), .B2(n9449), .A(n9448), .ZN(n9450) );
  AOI21_X1 U10733 ( .B1(n9451), .B2(n9516), .A(n9450), .ZN(n9460) );
  OAI211_X1 U10734 ( .C1(n9454), .C2(n9453), .A(n9499), .B(n9452), .ZN(n9459)
         );
  OAI211_X1 U10735 ( .C1(n9457), .C2(n9456), .A(n9517), .B(n9455), .ZN(n9458)
         );
  NAND3_X1 U10736 ( .A1(n9460), .A2(n9459), .A3(n9458), .ZN(P1_U3246) );
  INV_X1 U10737 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n9462) );
  NAND2_X1 U10738 ( .A1(P1_REG3_REG_5__SCAN_IN), .A2(P1_U3086), .ZN(n9461) );
  OAI21_X1 U10739 ( .B1(n9507), .B2(n9462), .A(n9461), .ZN(n9463) );
  AOI21_X1 U10740 ( .B1(n9464), .B2(n9516), .A(n9463), .ZN(n9474) );
  INV_X1 U10741 ( .A(n9465), .ZN(n9466) );
  OAI211_X1 U10742 ( .C1(n9468), .C2(n9467), .A(n9517), .B(n9466), .ZN(n9473)
         );
  OAI211_X1 U10743 ( .C1(n9471), .C2(n9470), .A(n9499), .B(n9469), .ZN(n9472)
         );
  NAND3_X1 U10744 ( .A1(n9474), .A2(n9473), .A3(n9472), .ZN(P1_U3248) );
  INV_X1 U10745 ( .A(n9475), .ZN(n9476) );
  NAND2_X1 U10746 ( .A1(n9517), .A2(n9476), .ZN(n9477) );
  AOI21_X1 U10747 ( .B1(n9478), .B2(n7921), .A(n9477), .ZN(n9479) );
  INV_X1 U10748 ( .A(n9479), .ZN(n9490) );
  INV_X1 U10749 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n9481) );
  NAND2_X1 U10750 ( .A1(P1_REG3_REG_15__SCAN_IN), .A2(P1_U3086), .ZN(n9480) );
  OAI21_X1 U10751 ( .B1(n9507), .B2(n9481), .A(n9480), .ZN(n9482) );
  AOI21_X1 U10752 ( .B1(n9483), .B2(n9516), .A(n9482), .ZN(n9489) );
  NAND2_X1 U10753 ( .A1(n9484), .A2(n6230), .ZN(n9487) );
  INV_X1 U10754 ( .A(n9485), .ZN(n9486) );
  NAND3_X1 U10755 ( .A1(n9499), .A2(n9487), .A3(n9486), .ZN(n9488) );
  NAND3_X1 U10756 ( .A1(n9490), .A2(n9489), .A3(n9488), .ZN(P1_U3258) );
  OAI21_X1 U10757 ( .B1(n9493), .B2(n9492), .A(n9491), .ZN(n9494) );
  NAND2_X1 U10758 ( .A1(n9494), .A2(n9517), .ZN(n9505) );
  AOI21_X1 U10759 ( .B1(n9956), .B2(P1_ADDR_REG_17__SCAN_IN), .A(n9495), .ZN(
        n9504) );
  OAI21_X1 U10760 ( .B1(n9498), .B2(n9497), .A(n9496), .ZN(n9500) );
  NAND2_X1 U10761 ( .A1(n9500), .A2(n9499), .ZN(n9503) );
  NAND2_X1 U10762 ( .A1(n9516), .A2(n9501), .ZN(n9502) );
  NAND4_X1 U10763 ( .A1(n9505), .A2(n9504), .A3(n9503), .A4(n9502), .ZN(
        P1_U3260) );
  INV_X1 U10764 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n10262) );
  NAND2_X1 U10765 ( .A1(P1_REG3_REG_18__SCAN_IN), .A2(P1_U3086), .ZN(n9506) );
  OAI21_X1 U10766 ( .B1(n9507), .B2(n10262), .A(n9506), .ZN(n9514) );
  INV_X1 U10767 ( .A(n9508), .ZN(n9509) );
  AOI211_X1 U10768 ( .C1(n9512), .C2(n9511), .A(n9510), .B(n9509), .ZN(n9513)
         );
  AOI211_X1 U10769 ( .C1(n9516), .C2(n9515), .A(n9514), .B(n9513), .ZN(n9522)
         );
  OAI211_X1 U10770 ( .C1(n9520), .C2(n9519), .A(n9518), .B(n9517), .ZN(n9521)
         );
  NAND2_X1 U10771 ( .A1(n9522), .A2(n9521), .ZN(P1_U3261) );
  NAND2_X1 U10772 ( .A1(n9523), .A2(n9709), .ZN(n9525) );
  AND2_X1 U10773 ( .A1(n9742), .A2(n9935), .ZN(n9528) );
  AOI21_X1 U10774 ( .B1(n9988), .B2(P1_REG2_REG_31__SCAN_IN), .A(n9528), .ZN(
        n9524) );
  OAI211_X1 U10775 ( .C1(n9526), .C2(n9990), .A(n9525), .B(n9524), .ZN(
        P1_U3263) );
  XNOR2_X1 U10776 ( .A(n9933), .B(n9545), .ZN(n9936) );
  NAND2_X1 U10777 ( .A1(n9936), .A2(n9709), .ZN(n9530) );
  AND2_X1 U10778 ( .A1(n10000), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n9527) );
  NOR2_X1 U10779 ( .A1(n9528), .A2(n9527), .ZN(n9529) );
  OAI211_X1 U10780 ( .C1(n9933), .C2(n9990), .A(n9530), .B(n9529), .ZN(
        P1_U3264) );
  XNOR2_X1 U10781 ( .A(n9543), .B(n9534), .ZN(n9540) );
  OAI22_X1 U10782 ( .A1(n9538), .A2(n9537), .B1(n9536), .B2(n9535), .ZN(n9539)
         );
  XNOR2_X1 U10783 ( .A(n9544), .B(n9543), .ZN(n9762) );
  OAI211_X1 U10784 ( .C1(n9852), .C2(n9546), .A(n9993), .B(n9545), .ZN(n9764)
         );
  INV_X1 U10785 ( .A(n9852), .ZN(n9550) );
  INV_X1 U10786 ( .A(P1_REG2_REG_29__SCAN_IN), .ZN(n9547) );
  OAI22_X1 U10787 ( .A1(n9548), .A2(n9970), .B1(n9547), .B2(n9742), .ZN(n9549)
         );
  AOI21_X1 U10788 ( .B1(n9550), .B2(n9633), .A(n9549), .ZN(n9551) );
  OAI21_X1 U10789 ( .B1(n9764), .B2(n9612), .A(n9551), .ZN(n9552) );
  AOI21_X1 U10790 ( .B1(n9762), .B2(n9929), .A(n9552), .ZN(n9553) );
  OAI21_X1 U10791 ( .B1(n9763), .B2(n9988), .A(n9553), .ZN(P1_U3356) );
  INV_X1 U10792 ( .A(n9554), .ZN(n9561) );
  AOI22_X1 U10793 ( .A1(n9555), .A2(n9987), .B1(P1_REG2_REG_28__SCAN_IN), .B2(
        n9988), .ZN(n9558) );
  NAND2_X1 U10794 ( .A1(n9556), .A2(n9633), .ZN(n9557) );
  OAI211_X1 U10795 ( .C1(n9559), .C2(n9612), .A(n9558), .B(n9557), .ZN(n9560)
         );
  AOI21_X1 U10796 ( .B1(n9561), .B2(n9929), .A(n9560), .ZN(n9562) );
  OAI21_X1 U10797 ( .B1(n9988), .B2(n9563), .A(n9562), .ZN(P1_U3265) );
  XNOR2_X1 U10798 ( .A(n9565), .B(n9564), .ZN(n9774) );
  INV_X1 U10799 ( .A(n9566), .ZN(n9567) );
  AOI21_X1 U10800 ( .B1(n9770), .B2(n9590), .A(n9567), .ZN(n9771) );
  AOI22_X1 U10801 ( .A1(n9568), .A2(n9987), .B1(P1_REG2_REG_27__SCAN_IN), .B2(
        n10000), .ZN(n9569) );
  OAI21_X1 U10802 ( .B1(n9570), .B2(n9990), .A(n9569), .ZN(n9580) );
  AOI21_X1 U10803 ( .B1(n9573), .B2(n4625), .A(n9982), .ZN(n9578) );
  INV_X1 U10804 ( .A(n9572), .ZN(n9575) );
  OAI21_X1 U10805 ( .B1(n9575), .B2(n9574), .A(n9573), .ZN(n9577) );
  AOI21_X1 U10806 ( .B1(n9578), .B2(n9577), .A(n9576), .ZN(n9773) );
  NOR2_X1 U10807 ( .A1(n9773), .A2(n10000), .ZN(n9579) );
  AOI211_X1 U10808 ( .C1(n9771), .C2(n9709), .A(n9580), .B(n9579), .ZN(n9581)
         );
  OAI21_X1 U10809 ( .B1(n9726), .B2(n9774), .A(n9581), .ZN(P1_U3266) );
  XNOR2_X1 U10810 ( .A(n9583), .B(n9582), .ZN(n9777) );
  INV_X1 U10811 ( .A(n9777), .ZN(n9598) );
  XNOR2_X1 U10812 ( .A(n9585), .B(n9584), .ZN(n9586) );
  NAND2_X1 U10813 ( .A1(n9586), .A2(n9837), .ZN(n9589) );
  INV_X1 U10814 ( .A(n9587), .ZN(n9588) );
  NAND2_X1 U10815 ( .A1(n9589), .A2(n9588), .ZN(n9775) );
  AOI211_X1 U10816 ( .C1(n9591), .C2(n9607), .A(n9831), .B(n4770), .ZN(n9776)
         );
  NAND2_X1 U10817 ( .A1(n9776), .A2(n9996), .ZN(n9595) );
  INV_X1 U10818 ( .A(n9592), .ZN(n9593) );
  AOI22_X1 U10819 ( .A1(n9593), .A2(n9987), .B1(P1_REG2_REG_26__SCAN_IN), .B2(
        n10000), .ZN(n9594) );
  OAI211_X1 U10820 ( .C1(n9857), .C2(n9990), .A(n9595), .B(n9594), .ZN(n9596)
         );
  AOI21_X1 U10821 ( .B1(n9742), .B2(n9775), .A(n9596), .ZN(n9597) );
  OAI21_X1 U10822 ( .B1(n9598), .B2(n9726), .A(n9597), .ZN(P1_U3267) );
  XNOR2_X1 U10823 ( .A(n9599), .B(n9601), .ZN(n9782) );
  NAND2_X1 U10824 ( .A1(n9619), .A2(n9600), .ZN(n9602) );
  NAND2_X1 U10825 ( .A1(n9602), .A2(n9601), .ZN(n9603) );
  NAND2_X1 U10826 ( .A1(n9604), .A2(n9603), .ZN(n9606) );
  AOI21_X1 U10827 ( .B1(n9606), .B2(n9837), .A(n9605), .ZN(n9781) );
  INV_X1 U10828 ( .A(n9781), .ZN(n9614) );
  OAI211_X1 U10829 ( .C1(n9861), .C2(n9624), .A(n9993), .B(n9607), .ZN(n9780)
         );
  AOI22_X1 U10830 ( .A1(n9608), .A2(n9987), .B1(P1_REG2_REG_25__SCAN_IN), .B2(
        n9988), .ZN(n9611) );
  NAND2_X1 U10831 ( .A1(n9609), .A2(n9633), .ZN(n9610) );
  OAI211_X1 U10832 ( .C1(n9780), .C2(n9612), .A(n9611), .B(n9610), .ZN(n9613)
         );
  AOI21_X1 U10833 ( .B1(n9614), .B2(n9742), .A(n9613), .ZN(n9615) );
  OAI21_X1 U10834 ( .B1(n9782), .B2(n9726), .A(n9615), .ZN(P1_U3268) );
  XOR2_X1 U10835 ( .A(n9617), .B(n9616), .Z(n9788) );
  INV_X1 U10836 ( .A(n9788), .ZN(n9631) );
  AOI21_X1 U10837 ( .B1(n9618), .B2(n9635), .A(n9617), .ZN(n9623) );
  NAND2_X1 U10838 ( .A1(n9619), .A2(n9837), .ZN(n9622) );
  INV_X1 U10839 ( .A(n9620), .ZN(n9621) );
  OAI21_X1 U10840 ( .B1(n9623), .B2(n9622), .A(n9621), .ZN(n9786) );
  AOI211_X1 U10841 ( .C1(n9625), .C2(n4531), .A(n9831), .B(n9624), .ZN(n9787)
         );
  NAND2_X1 U10842 ( .A1(n9787), .A2(n9996), .ZN(n9628) );
  AOI22_X1 U10843 ( .A1(n9626), .A2(n9987), .B1(P1_REG2_REG_24__SCAN_IN), .B2(
        n10000), .ZN(n9627) );
  OAI211_X1 U10844 ( .C1(n9865), .C2(n9990), .A(n9628), .B(n9627), .ZN(n9629)
         );
  AOI21_X1 U10845 ( .B1(n9742), .B2(n9786), .A(n9629), .ZN(n9630) );
  OAI21_X1 U10846 ( .B1(n9631), .B2(n9726), .A(n9630), .ZN(P1_U3269) );
  XNOR2_X1 U10847 ( .A(n9632), .B(n9637), .ZN(n9797) );
  INV_X1 U10848 ( .A(n9797), .ZN(n9646) );
  AOI22_X1 U10849 ( .A1(n9791), .A2(n9633), .B1(P1_REG2_REG_23__SCAN_IN), .B2(
        n9988), .ZN(n9645) );
  AOI21_X1 U10850 ( .B1(n9649), .B2(n9791), .A(n9831), .ZN(n9634) );
  NAND2_X1 U10851 ( .A1(n9634), .A2(n4531), .ZN(n9793) );
  OAI21_X1 U10852 ( .B1(n9637), .B2(n9636), .A(n9635), .ZN(n9638) );
  NAND2_X1 U10853 ( .A1(n9638), .A2(n9837), .ZN(n9795) );
  INV_X1 U10854 ( .A(n9639), .ZN(n9640) );
  AOI21_X1 U10855 ( .B1(n9640), .B2(n9987), .A(n9792), .ZN(n9641) );
  OAI211_X1 U10856 ( .C1(n4509), .C2(n9793), .A(n9795), .B(n9641), .ZN(n9643)
         );
  NAND2_X1 U10857 ( .A1(n9643), .A2(n9742), .ZN(n9644) );
  OAI211_X1 U10858 ( .C1(n9646), .C2(n9726), .A(n9645), .B(n9644), .ZN(
        P1_U3270) );
  XNOR2_X1 U10859 ( .A(n9648), .B(n9647), .ZN(n9804) );
  INV_X1 U10860 ( .A(n9670), .ZN(n9651) );
  INV_X1 U10861 ( .A(n9649), .ZN(n9650) );
  AOI21_X1 U10862 ( .B1(n9800), .B2(n9651), .A(n9650), .ZN(n9801) );
  AOI22_X1 U10863 ( .A1(n9652), .A2(n9987), .B1(P1_REG2_REG_22__SCAN_IN), .B2(
        n9988), .ZN(n9653) );
  OAI21_X1 U10864 ( .B1(n9654), .B2(n9990), .A(n9653), .ZN(n9660) );
  XNOR2_X1 U10865 ( .A(n9656), .B(n9655), .ZN(n9658) );
  AOI21_X1 U10866 ( .B1(n9658), .B2(n9837), .A(n9657), .ZN(n9803) );
  NOR2_X1 U10867 ( .A1(n9803), .A2(n9988), .ZN(n9659) );
  AOI211_X1 U10868 ( .C1(n9801), .C2(n9709), .A(n9660), .B(n9659), .ZN(n9661)
         );
  OAI21_X1 U10869 ( .B1(n9726), .B2(n9804), .A(n9661), .ZN(P1_U3271) );
  XNOR2_X1 U10870 ( .A(n9663), .B(n9662), .ZN(n9807) );
  INV_X1 U10871 ( .A(n9807), .ZN(n9678) );
  XNOR2_X1 U10872 ( .A(n9665), .B(n9664), .ZN(n9666) );
  INV_X1 U10873 ( .A(n9667), .ZN(n9668) );
  NAND2_X1 U10874 ( .A1(n9669), .A2(n9668), .ZN(n9806) );
  INV_X1 U10875 ( .A(n9671), .ZN(n9874) );
  AOI211_X1 U10876 ( .C1(n9671), .C2(n9686), .A(n9831), .B(n9670), .ZN(n9805)
         );
  NAND2_X1 U10877 ( .A1(n9805), .A2(n9996), .ZN(n9675) );
  INV_X1 U10878 ( .A(n9672), .ZN(n9673) );
  AOI22_X1 U10879 ( .A1(n9673), .A2(n9987), .B1(P1_REG2_REG_21__SCAN_IN), .B2(
        n10000), .ZN(n9674) );
  OAI211_X1 U10880 ( .C1(n9874), .C2(n9990), .A(n9675), .B(n9674), .ZN(n9676)
         );
  AOI21_X1 U10881 ( .B1(n9742), .B2(n9806), .A(n9676), .ZN(n9677) );
  OAI21_X1 U10882 ( .B1(n9726), .B2(n9678), .A(n9677), .ZN(P1_U3272) );
  XNOR2_X1 U10883 ( .A(n9679), .B(n9681), .ZN(n9812) );
  INV_X1 U10884 ( .A(n9812), .ZN(n9694) );
  OAI211_X1 U10885 ( .C1(n9682), .C2(n9681), .A(n9680), .B(n9837), .ZN(n9685)
         );
  INV_X1 U10886 ( .A(n9683), .ZN(n9684) );
  NAND2_X1 U10887 ( .A1(n9685), .A2(n9684), .ZN(n9810) );
  INV_X1 U10888 ( .A(n9686), .ZN(n9687) );
  AOI211_X1 U10889 ( .C1(n9688), .C2(n9696), .A(n9831), .B(n9687), .ZN(n9811)
         );
  NAND2_X1 U10890 ( .A1(n9811), .A2(n9996), .ZN(n9691) );
  AOI22_X1 U10891 ( .A1(n9988), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n9689), .B2(
        n9987), .ZN(n9690) );
  OAI211_X1 U10892 ( .C1(n4765), .C2(n9990), .A(n9691), .B(n9690), .ZN(n9692)
         );
  AOI21_X1 U10893 ( .B1(n9742), .B2(n9810), .A(n9692), .ZN(n9693) );
  OAI21_X1 U10894 ( .B1(n9694), .B2(n9726), .A(n9693), .ZN(P1_U3273) );
  XNOR2_X1 U10895 ( .A(n9695), .B(n9702), .ZN(n9819) );
  INV_X1 U10896 ( .A(n9696), .ZN(n9697) );
  AOI21_X1 U10897 ( .B1(n9815), .B2(n4769), .A(n9697), .ZN(n9816) );
  INV_X1 U10898 ( .A(n9698), .ZN(n9699) );
  AOI22_X1 U10899 ( .A1(n9988), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n9699), .B2(
        n9987), .ZN(n9700) );
  OAI21_X1 U10900 ( .B1(n9701), .B2(n9990), .A(n9700), .ZN(n9708) );
  AOI21_X1 U10901 ( .B1(n9703), .B2(n9702), .A(n9982), .ZN(n9706) );
  AOI21_X1 U10902 ( .B1(n9706), .B2(n9705), .A(n9704), .ZN(n9818) );
  NOR2_X1 U10903 ( .A1(n9818), .A2(n10000), .ZN(n9707) );
  AOI211_X1 U10904 ( .C1(n9816), .C2(n9709), .A(n9708), .B(n9707), .ZN(n9710)
         );
  OAI21_X1 U10905 ( .B1(n9726), .B2(n9819), .A(n9710), .ZN(P1_U3274) );
  XNOR2_X1 U10906 ( .A(n9711), .B(n9712), .ZN(n9822) );
  INV_X1 U10907 ( .A(n9822), .ZN(n9727) );
  XNOR2_X1 U10908 ( .A(n9713), .B(n9712), .ZN(n9714) );
  NAND2_X1 U10909 ( .A1(n9714), .A2(n9837), .ZN(n9717) );
  INV_X1 U10910 ( .A(n9715), .ZN(n9716) );
  NAND2_X1 U10911 ( .A1(n9717), .A2(n9716), .ZN(n9820) );
  INV_X1 U10912 ( .A(n9719), .ZN(n9882) );
  AOI211_X1 U10913 ( .C1(n9719), .C2(n9737), .A(n9831), .B(n9718), .ZN(n9821)
         );
  NAND2_X1 U10914 ( .A1(n9821), .A2(n9996), .ZN(n9723) );
  INV_X1 U10915 ( .A(n9720), .ZN(n9721) );
  AOI22_X1 U10916 ( .A1(n9988), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n9721), .B2(
        n9987), .ZN(n9722) );
  OAI211_X1 U10917 ( .C1(n9882), .C2(n9990), .A(n9723), .B(n9722), .ZN(n9724)
         );
  AOI21_X1 U10918 ( .B1(n9742), .B2(n9820), .A(n9724), .ZN(n9725) );
  OAI21_X1 U10919 ( .B1(n9727), .B2(n9726), .A(n9725), .ZN(P1_U3275) );
  NAND3_X1 U10920 ( .A1(n9730), .A2(n9837), .A3(n9729), .ZN(n9733) );
  INV_X1 U10921 ( .A(n9731), .ZN(n9732) );
  NAND2_X1 U10922 ( .A1(n9733), .A2(n9732), .ZN(n9825) );
  INV_X1 U10923 ( .A(n9825), .ZN(n9747) );
  XNOR2_X1 U10924 ( .A(n9735), .B(n9734), .ZN(n9827) );
  NAND2_X1 U10925 ( .A1(n9827), .A2(n9929), .ZN(n9746) );
  INV_X1 U10926 ( .A(n4515), .ZN(n9830) );
  INV_X1 U10927 ( .A(n9737), .ZN(n9738) );
  AOI211_X1 U10928 ( .C1(n9739), .C2(n9830), .A(n9831), .B(n9738), .ZN(n9826)
         );
  NOR2_X1 U10929 ( .A1(n6494), .A2(n9990), .ZN(n9744) );
  OAI22_X1 U10930 ( .A1(n9742), .A2(n9741), .B1(n9740), .B2(n9970), .ZN(n9743)
         );
  AOI211_X1 U10931 ( .C1(n9826), .C2(n9996), .A(n9744), .B(n9743), .ZN(n9745)
         );
  OAI211_X1 U10932 ( .C1(n10000), .C2(n9747), .A(n9746), .B(n9745), .ZN(
        P1_U3276) );
  OAI21_X1 U10933 ( .B1(n4588), .B2(n9752), .A(n9748), .ZN(n9750) );
  AOI21_X1 U10934 ( .B1(n9750), .B2(n9837), .A(n9749), .ZN(n10076) );
  XOR2_X1 U10935 ( .A(n9752), .B(n9751), .Z(n10078) );
  INV_X1 U10936 ( .A(n10078), .ZN(n10080) );
  NAND2_X1 U10937 ( .A1(n10080), .A2(n9929), .ZN(n9761) );
  AOI211_X1 U10938 ( .C1(n10073), .C2(n4764), .A(n9831), .B(n9754), .ZN(n10072) );
  NOR2_X1 U10939 ( .A1(n9755), .A2(n9990), .ZN(n9759) );
  OAI22_X1 U10940 ( .A1(n9742), .A2(n9757), .B1(n9756), .B2(n9970), .ZN(n9758)
         );
  AOI211_X1 U10941 ( .C1(n10072), .C2(n9996), .A(n9759), .B(n9758), .ZN(n9760)
         );
  OAI211_X1 U10942 ( .C1(n9988), .C2(n10076), .A(n9761), .B(n9760), .ZN(
        P1_U3279) );
  NAND2_X1 U10943 ( .A1(n9762), .A2(n10070), .ZN(n9765) );
  NAND2_X1 U10944 ( .A1(n10100), .A2(n9766), .ZN(n9767) );
  NAND2_X1 U10945 ( .A1(n9768), .A2(n9767), .ZN(n9769) );
  OAI21_X1 U10946 ( .B1(n9852), .B2(n9846), .A(n9769), .ZN(P1_U3551) );
  AOI22_X1 U10947 ( .A1(n9771), .A2(n9993), .B1(n10074), .B2(n9770), .ZN(n9772) );
  OAI211_X1 U10948 ( .C1(n9774), .C2(n10034), .A(n9773), .B(n9772), .ZN(n9853)
         );
  MUX2_X1 U10949 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n9853), .S(n10102), .Z(
        P1_U3549) );
  AOI211_X1 U10950 ( .C1(n9777), .C2(n10070), .A(n9776), .B(n9775), .ZN(n9854)
         );
  MUX2_X1 U10951 ( .A(n9778), .B(n9854), .S(n10102), .Z(n9779) );
  OAI21_X1 U10952 ( .B1(n9857), .B2(n9846), .A(n9779), .ZN(P1_U3548) );
  OAI211_X1 U10953 ( .C1(n9782), .C2(n10034), .A(n9781), .B(n9780), .ZN(n9783)
         );
  INV_X1 U10954 ( .A(n9783), .ZN(n9859) );
  MUX2_X1 U10955 ( .A(n9859), .B(n9784), .S(n10100), .Z(n9785) );
  OAI21_X1 U10956 ( .B1(n9861), .B2(n9846), .A(n9785), .ZN(P1_U3547) );
  AOI211_X1 U10957 ( .C1(n9788), .C2(n10070), .A(n9787), .B(n9786), .ZN(n9862)
         );
  MUX2_X1 U10958 ( .A(n9789), .B(n9862), .S(n10102), .Z(n9790) );
  OAI21_X1 U10959 ( .B1(n9865), .B2(n9846), .A(n9790), .ZN(P1_U3546) );
  INV_X1 U10960 ( .A(n9791), .ZN(n9869) );
  INV_X1 U10961 ( .A(n9792), .ZN(n9794) );
  NAND3_X1 U10962 ( .A1(n9795), .A2(n9794), .A3(n9793), .ZN(n9796) );
  AOI21_X1 U10963 ( .B1(n9797), .B2(n10070), .A(n9796), .ZN(n9866) );
  MUX2_X1 U10964 ( .A(n9798), .B(n9866), .S(n10102), .Z(n9799) );
  OAI21_X1 U10965 ( .B1(n9869), .B2(n9846), .A(n9799), .ZN(P1_U3545) );
  AOI22_X1 U10966 ( .A1(n9801), .A2(n9993), .B1(n10074), .B2(n9800), .ZN(n9802) );
  OAI211_X1 U10967 ( .C1(n9804), .C2(n10034), .A(n9803), .B(n9802), .ZN(n9870)
         );
  MUX2_X1 U10968 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n9870), .S(n10102), .Z(
        P1_U3544) );
  INV_X1 U10969 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n9808) );
  AOI211_X1 U10970 ( .C1(n9807), .C2(n10070), .A(n9806), .B(n9805), .ZN(n9871)
         );
  MUX2_X1 U10971 ( .A(n9808), .B(n9871), .S(n10102), .Z(n9809) );
  OAI21_X1 U10972 ( .B1(n9874), .B2(n9846), .A(n9809), .ZN(P1_U3543) );
  INV_X1 U10973 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n9813) );
  AOI211_X1 U10974 ( .C1(n9812), .C2(n10070), .A(n9811), .B(n9810), .ZN(n9875)
         );
  MUX2_X1 U10975 ( .A(n9813), .B(n9875), .S(n10102), .Z(n9814) );
  OAI21_X1 U10976 ( .B1(n4765), .B2(n9846), .A(n9814), .ZN(P1_U3542) );
  AOI22_X1 U10977 ( .A1(n9816), .A2(n9993), .B1(n10074), .B2(n9815), .ZN(n9817) );
  OAI211_X1 U10978 ( .C1(n9819), .C2(n10034), .A(n9818), .B(n9817), .ZN(n9878)
         );
  MUX2_X1 U10979 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n9878), .S(n10102), .Z(
        P1_U3541) );
  AOI211_X1 U10980 ( .C1(n9822), .C2(n10070), .A(n9821), .B(n9820), .ZN(n9879)
         );
  MUX2_X1 U10981 ( .A(n9823), .B(n9879), .S(n10102), .Z(n9824) );
  OAI21_X1 U10982 ( .B1(n9882), .B2(n9846), .A(n9824), .ZN(P1_U3540) );
  AOI211_X1 U10983 ( .C1(n9827), .C2(n10070), .A(n9826), .B(n9825), .ZN(n9883)
         );
  MUX2_X1 U10984 ( .A(n6277), .B(n9883), .S(n10102), .Z(n9828) );
  OAI21_X1 U10985 ( .B1(n6494), .B2(n9846), .A(n9828), .ZN(P1_U3539) );
  XNOR2_X1 U10986 ( .A(n9829), .B(n9834), .ZN(n9930) );
  AOI211_X1 U10987 ( .C1(n9833), .C2(n9832), .A(n9831), .B(n4515), .ZN(n9922)
         );
  XNOR2_X1 U10988 ( .A(n9835), .B(n9834), .ZN(n9838) );
  AOI21_X1 U10989 ( .B1(n9838), .B2(n9837), .A(n9836), .ZN(n9932) );
  INV_X1 U10990 ( .A(n9932), .ZN(n9839) );
  AOI211_X1 U10991 ( .C1(n9930), .C2(n10070), .A(n9922), .B(n9839), .ZN(n9886)
         );
  MUX2_X1 U10992 ( .A(n6254), .B(n9886), .S(n10102), .Z(n9840) );
  OAI21_X1 U10993 ( .B1(n9927), .B2(n9846), .A(n9840), .ZN(P1_U3538) );
  OAI211_X1 U10994 ( .C1(n9843), .C2(n10034), .A(n9842), .B(n9841), .ZN(n9844)
         );
  INV_X1 U10995 ( .A(n9844), .ZN(n9888) );
  MUX2_X1 U10996 ( .A(n6230), .B(n9888), .S(n10102), .Z(n9845) );
  OAI21_X1 U10997 ( .B1(n9892), .B2(n9846), .A(n9845), .ZN(P1_U3537) );
  MUX2_X1 U10998 ( .A(n9847), .B(P1_REG1_REG_0__SCAN_IN), .S(n10100), .Z(
        P1_U3522) );
  OAI21_X1 U10999 ( .B1(n9852), .B2(n9891), .A(n9851), .ZN(P1_U3519) );
  MUX2_X1 U11000 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n9853), .S(n10084), .Z(
        P1_U3517) );
  INV_X1 U11001 ( .A(P1_REG0_REG_26__SCAN_IN), .ZN(n9855) );
  MUX2_X1 U11002 ( .A(n9855), .B(n9854), .S(n10084), .Z(n9856) );
  OAI21_X1 U11003 ( .B1(n9857), .B2(n9891), .A(n9856), .ZN(P1_U3516) );
  INV_X1 U11004 ( .A(P1_REG0_REG_25__SCAN_IN), .ZN(n9858) );
  MUX2_X1 U11005 ( .A(n9859), .B(n9858), .S(n10082), .Z(n9860) );
  OAI21_X1 U11006 ( .B1(n9861), .B2(n9891), .A(n9860), .ZN(P1_U3515) );
  INV_X1 U11007 ( .A(P1_REG0_REG_24__SCAN_IN), .ZN(n9863) );
  MUX2_X1 U11008 ( .A(n9863), .B(n9862), .S(n10084), .Z(n9864) );
  OAI21_X1 U11009 ( .B1(n9865), .B2(n9891), .A(n9864), .ZN(P1_U3514) );
  INV_X1 U11010 ( .A(P1_REG0_REG_23__SCAN_IN), .ZN(n9867) );
  MUX2_X1 U11011 ( .A(n9867), .B(n9866), .S(n10084), .Z(n9868) );
  OAI21_X1 U11012 ( .B1(n9869), .B2(n9891), .A(n9868), .ZN(P1_U3513) );
  MUX2_X1 U11013 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n9870), .S(n10084), .Z(
        P1_U3512) );
  INV_X1 U11014 ( .A(P1_REG0_REG_21__SCAN_IN), .ZN(n9872) );
  MUX2_X1 U11015 ( .A(n9872), .B(n9871), .S(n10084), .Z(n9873) );
  OAI21_X1 U11016 ( .B1(n9874), .B2(n9891), .A(n9873), .ZN(P1_U3511) );
  INV_X1 U11017 ( .A(P1_REG0_REG_20__SCAN_IN), .ZN(n9876) );
  MUX2_X1 U11018 ( .A(n9876), .B(n9875), .S(n10084), .Z(n9877) );
  OAI21_X1 U11019 ( .B1(n4765), .B2(n9891), .A(n9877), .ZN(P1_U3510) );
  MUX2_X1 U11020 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n9878), .S(n10084), .Z(
        P1_U3509) );
  INV_X1 U11021 ( .A(P1_REG0_REG_18__SCAN_IN), .ZN(n9880) );
  MUX2_X1 U11022 ( .A(n9880), .B(n9879), .S(n10084), .Z(n9881) );
  OAI21_X1 U11023 ( .B1(n9882), .B2(n9891), .A(n9881), .ZN(P1_U3507) );
  INV_X1 U11024 ( .A(P1_REG0_REG_17__SCAN_IN), .ZN(n9884) );
  MUX2_X1 U11025 ( .A(n9884), .B(n9883), .S(n10084), .Z(n9885) );
  OAI21_X1 U11026 ( .B1(n6494), .B2(n9891), .A(n9885), .ZN(P1_U3504) );
  MUX2_X1 U11027 ( .A(n6259), .B(n9886), .S(n10084), .Z(n9887) );
  OAI21_X1 U11028 ( .B1(n9927), .B2(n9891), .A(n9887), .ZN(P1_U3501) );
  INV_X1 U11029 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n9889) );
  MUX2_X1 U11030 ( .A(n9889), .B(n9888), .S(n10084), .Z(n9890) );
  OAI21_X1 U11031 ( .B1(n9892), .B2(n9891), .A(n9890), .ZN(P1_U3498) );
  MUX2_X1 U11032 ( .A(n9894), .B(P1_D_REG_0__SCAN_IN), .S(n9893), .Z(P1_U3439)
         );
  INV_X1 U11033 ( .A(n9895), .ZN(n9900) );
  NOR4_X1 U11034 ( .A1(n9896), .A2(P1_IR_REG_30__SCAN_IN), .A3(P1_U3086), .A4(
        n5848), .ZN(n9897) );
  AOI21_X1 U11035 ( .B1(n9898), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n9897), .ZN(
        n9899) );
  OAI21_X1 U11036 ( .B1(n9900), .B2(n9905), .A(n9899), .ZN(P1_U3324) );
  OAI222_X1 U11037 ( .A1(n9905), .A2(n9902), .B1(n9901), .B2(P1_U3086), .C1(
        n10338), .C2(n9903), .ZN(P1_U3326) );
  INV_X1 U11038 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n10571) );
  OAI222_X1 U11039 ( .A1(n9905), .A2(n9904), .B1(n6442), .B2(P1_U3086), .C1(
        n10571), .C2(n9903), .ZN(P1_U3327) );
  INV_X1 U11040 ( .A(n9906), .ZN(n9907) );
  MUX2_X1 U11041 ( .A(n9907), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  AOI21_X1 U11042 ( .B1(n9910), .B2(n9909), .A(n4580), .ZN(n9917) );
  INV_X1 U11043 ( .A(n9911), .ZN(n9913) );
  NOR2_X1 U11044 ( .A1(n10068), .A2(n9946), .ZN(n9912) );
  AOI211_X1 U11045 ( .C1(n4510), .C2(n9914), .A(n9913), .B(n9912), .ZN(n9915)
         );
  OAI21_X1 U11046 ( .B1(n9917), .B2(n9916), .A(n9915), .ZN(n9918) );
  INV_X1 U11047 ( .A(n9918), .ZN(n9919) );
  OAI21_X1 U11048 ( .B1(n9921), .B2(n9920), .A(n9919), .ZN(P1_U3217) );
  NAND2_X1 U11049 ( .A1(n9922), .A2(n9996), .ZN(n9926) );
  INV_X1 U11050 ( .A(n9923), .ZN(n9924) );
  AOI22_X1 U11051 ( .A1(n9988), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n9924), .B2(
        n9987), .ZN(n9925) );
  OAI211_X1 U11052 ( .C1(n9927), .C2(n9990), .A(n9926), .B(n9925), .ZN(n9928)
         );
  AOI21_X1 U11053 ( .B1(n9930), .B2(n9929), .A(n9928), .ZN(n9931) );
  OAI21_X1 U11054 ( .B1(n10000), .B2(n9932), .A(n9931), .ZN(P1_U3277) );
  NOR2_X1 U11055 ( .A1(n9933), .A2(n10067), .ZN(n9934) );
  AOI22_X1 U11056 ( .A1(n10102), .A2(n9938), .B1(n6875), .B2(n10100), .ZN(
        P1_U3552) );
  INV_X1 U11057 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n9937) );
  AOI22_X1 U11058 ( .A1(n10084), .A2(n9938), .B1(n9937), .B2(n10082), .ZN(
        P1_U3520) );
  XNOR2_X1 U11059 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  XNOR2_X1 U11060 ( .A(P1_RD_REG_SCAN_IN), .B(P2_RD_REG_SCAN_IN), .ZN(U126) );
  OAI21_X1 U11061 ( .B1(n9940), .B2(n9939), .A(n9297), .ZN(n9949) );
  INV_X1 U11062 ( .A(n9941), .ZN(n10053) );
  INV_X1 U11063 ( .A(n9942), .ZN(n9943) );
  AOI21_X1 U11064 ( .B1(n9944), .B2(n4510), .A(n9943), .ZN(n9945) );
  OAI21_X1 U11065 ( .B1(n10053), .B2(n9946), .A(n9945), .ZN(n9947) );
  AOI21_X1 U11066 ( .B1(n9949), .B2(n9948), .A(n9947), .ZN(n9950) );
  OAI21_X1 U11067 ( .B1(n9952), .B2(n9951), .A(n9950), .ZN(P1_U3221) );
  AOI21_X1 U11068 ( .B1(n4508), .B2(n9954), .A(n9953), .ZN(n9955) );
  XNOR2_X1 U11069 ( .A(n9955), .B(P1_IR_REG_0__SCAN_IN), .ZN(n9959) );
  AOI22_X1 U11070 ( .A1(n9956), .A2(P1_ADDR_REG_0__SCAN_IN), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(P1_U3086), .ZN(n9957) );
  OAI21_X1 U11071 ( .B1(n9959), .B2(n9958), .A(n9957), .ZN(P1_U3243) );
  INV_X1 U11072 ( .A(n9960), .ZN(n10081) );
  XNOR2_X1 U11073 ( .A(n9961), .B(n9962), .ZN(n10047) );
  NAND3_X1 U11074 ( .A1(n9964), .A2(n9963), .A3(n9962), .ZN(n9965) );
  AOI21_X1 U11075 ( .B1(n9966), .B2(n9965), .A(n9982), .ZN(n9967) );
  AOI211_X1 U11076 ( .C1(n10081), .C2(n10047), .A(n9968), .B(n9967), .ZN(
        n10044) );
  NOR2_X1 U11077 ( .A1(n9970), .A2(n9969), .ZN(n9971) );
  AOI21_X1 U11078 ( .B1(n9988), .B2(P1_REG2_REG_7__SCAN_IN), .A(n9971), .ZN(
        n9972) );
  OAI21_X1 U11079 ( .B1(n9990), .B2(n10043), .A(n9972), .ZN(n9973) );
  INV_X1 U11080 ( .A(n9973), .ZN(n9979) );
  INV_X1 U11081 ( .A(n9974), .ZN(n9997) );
  OAI211_X1 U11082 ( .C1(n9976), .C2(n10043), .A(n9975), .B(n9993), .ZN(n10042) );
  INV_X1 U11083 ( .A(n10042), .ZN(n9977) );
  AOI22_X1 U11084 ( .A1(n10047), .A2(n9997), .B1(n9996), .B2(n9977), .ZN(n9978) );
  OAI211_X1 U11085 ( .C1(n10000), .C2(n10044), .A(n9979), .B(n9978), .ZN(
        P1_U3286) );
  NOR2_X1 U11086 ( .A1(n9983), .A2(n9982), .ZN(n9984) );
  AOI211_X1 U11087 ( .C1(n10081), .C2(n10007), .A(n9985), .B(n9984), .ZN(
        n10004) );
  AOI22_X1 U11088 ( .A1(n9988), .A2(P1_REG2_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(n9987), .ZN(n9989) );
  OAI21_X1 U11089 ( .B1(n9990), .B2(n4998), .A(n9989), .ZN(n9991) );
  INV_X1 U11090 ( .A(n9991), .ZN(n9999) );
  OAI211_X1 U11091 ( .C1(n4998), .C2(n9994), .A(n9993), .B(n9992), .ZN(n10003)
         );
  INV_X1 U11092 ( .A(n10003), .ZN(n9995) );
  AOI22_X1 U11093 ( .A1(n10007), .A2(n9997), .B1(n9996), .B2(n9995), .ZN(n9998) );
  OAI211_X1 U11094 ( .C1(n10000), .C2(n10004), .A(n9999), .B(n9998), .ZN(
        P1_U3292) );
  AND2_X1 U11095 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n10001), .ZN(P1_U3294) );
  AND2_X1 U11096 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n10001), .ZN(P1_U3295) );
  AND2_X1 U11097 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n10001), .ZN(P1_U3296) );
  AND2_X1 U11098 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n10001), .ZN(P1_U3297) );
  AND2_X1 U11099 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n10001), .ZN(P1_U3298) );
  AND2_X1 U11100 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n10001), .ZN(P1_U3299) );
  AND2_X1 U11101 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n10001), .ZN(P1_U3300) );
  AND2_X1 U11102 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n10001), .ZN(P1_U3301) );
  AND2_X1 U11103 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n10001), .ZN(P1_U3302) );
  AND2_X1 U11104 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n10001), .ZN(P1_U3303) );
  AND2_X1 U11105 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n10001), .ZN(P1_U3304) );
  AND2_X1 U11106 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n10001), .ZN(P1_U3305) );
  AND2_X1 U11107 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n10001), .ZN(P1_U3306) );
  AND2_X1 U11108 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n10001), .ZN(P1_U3307) );
  AND2_X1 U11109 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n10001), .ZN(P1_U3308) );
  AND2_X1 U11110 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n10001), .ZN(P1_U3309) );
  AND2_X1 U11111 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n10001), .ZN(P1_U3310) );
  AND2_X1 U11112 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n10001), .ZN(P1_U3311) );
  AND2_X1 U11113 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n10001), .ZN(P1_U3312) );
  AND2_X1 U11114 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n10001), .ZN(P1_U3313) );
  AND2_X1 U11115 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n10001), .ZN(P1_U3314) );
  AND2_X1 U11116 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n10001), .ZN(P1_U3315) );
  AND2_X1 U11117 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n10001), .ZN(P1_U3316) );
  AND2_X1 U11118 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n10001), .ZN(P1_U3317) );
  AND2_X1 U11119 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n10001), .ZN(P1_U3318) );
  AND2_X1 U11120 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n10001), .ZN(P1_U3319) );
  INV_X1 U11121 ( .A(P1_D_REG_5__SCAN_IN), .ZN(n10541) );
  NOR2_X1 U11122 ( .A1(n10002), .A2(n10541), .ZN(P1_U3320) );
  INV_X1 U11123 ( .A(P1_D_REG_4__SCAN_IN), .ZN(n10553) );
  NOR2_X1 U11124 ( .A1(n10002), .A2(n10553), .ZN(P1_U3321) );
  AND2_X1 U11125 ( .A1(n10001), .A2(P1_D_REG_3__SCAN_IN), .ZN(P1_U3322) );
  INV_X1 U11126 ( .A(P1_D_REG_2__SCAN_IN), .ZN(n10597) );
  NOR2_X1 U11127 ( .A1(n10002), .A2(n10597), .ZN(P1_U3323) );
  INV_X1 U11128 ( .A(n10077), .ZN(n10048) );
  OAI21_X1 U11129 ( .B1(n4998), .B2(n10067), .A(n10003), .ZN(n10006) );
  INV_X1 U11130 ( .A(n10004), .ZN(n10005) );
  AOI211_X1 U11131 ( .C1(n10048), .C2(n10007), .A(n10006), .B(n10005), .ZN(
        n10086) );
  INV_X1 U11132 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n10008) );
  AOI22_X1 U11133 ( .A1(n10084), .A2(n10086), .B1(n10008), .B2(n10082), .ZN(
        P1_U3456) );
  INV_X1 U11134 ( .A(n10009), .ZN(n10010) );
  OAI21_X1 U11135 ( .B1(n10011), .B2(n10067), .A(n10010), .ZN(n10014) );
  INV_X1 U11136 ( .A(n10012), .ZN(n10013) );
  AOI211_X1 U11137 ( .C1(n10070), .C2(n10015), .A(n10014), .B(n10013), .ZN(
        n10087) );
  AOI22_X1 U11138 ( .A1(n10084), .A2(n10087), .B1(n5938), .B2(n10082), .ZN(
        P1_U3459) );
  OAI21_X1 U11139 ( .B1(n10017), .B2(n10067), .A(n10016), .ZN(n10020) );
  INV_X1 U11140 ( .A(n10018), .ZN(n10019) );
  AOI211_X1 U11141 ( .C1(n10070), .C2(n10021), .A(n10020), .B(n10019), .ZN(
        n10088) );
  AOI22_X1 U11142 ( .A1(n10084), .A2(n10088), .B1(n5962), .B2(n10082), .ZN(
        P1_U3462) );
  INV_X1 U11143 ( .A(n10022), .ZN(n10028) );
  NOR2_X1 U11144 ( .A1(n10023), .A2(n10034), .ZN(n10027) );
  NOR2_X1 U11145 ( .A1(n10024), .A2(n10067), .ZN(n10025) );
  NOR4_X1 U11146 ( .A1(n10028), .A2(n10027), .A3(n10026), .A4(n10025), .ZN(
        n10089) );
  INV_X1 U11147 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n10029) );
  AOI22_X1 U11148 ( .A1(n10084), .A2(n10089), .B1(n10029), .B2(n10082), .ZN(
        P1_U3465) );
  AOI21_X1 U11149 ( .B1(n10074), .B2(n10031), .A(n10030), .ZN(n10032) );
  OAI21_X1 U11150 ( .B1(n10034), .B2(n10033), .A(n10032), .ZN(n10036) );
  NOR2_X1 U11151 ( .A1(n10036), .A2(n10035), .ZN(n10091) );
  AOI22_X1 U11152 ( .A1(n10084), .A2(n10091), .B1(n5999), .B2(n10082), .ZN(
        P1_U3468) );
  OAI211_X1 U11153 ( .C1(n10039), .C2(n10067), .A(n10038), .B(n10037), .ZN(
        n10040) );
  AOI21_X1 U11154 ( .B1(n10070), .B2(n10041), .A(n10040), .ZN(n10093) );
  AOI22_X1 U11155 ( .A1(n10084), .A2(n10093), .B1(n6022), .B2(n10082), .ZN(
        P1_U3471) );
  OAI21_X1 U11156 ( .B1(n10043), .B2(n10067), .A(n10042), .ZN(n10046) );
  INV_X1 U11157 ( .A(n10044), .ZN(n10045) );
  AOI211_X1 U11158 ( .C1(n10048), .C2(n10047), .A(n10046), .B(n10045), .ZN(
        n10094) );
  INV_X1 U11159 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n10049) );
  AOI22_X1 U11160 ( .A1(n10084), .A2(n10094), .B1(n10049), .B2(n10082), .ZN(
        P1_U3474) );
  INV_X1 U11161 ( .A(n10050), .ZN(n10056) );
  NOR2_X1 U11162 ( .A1(n10050), .A2(n10077), .ZN(n10055) );
  OAI211_X1 U11163 ( .C1(n10053), .C2(n10067), .A(n10052), .B(n10051), .ZN(
        n10054) );
  AOI211_X1 U11164 ( .C1(n10081), .C2(n10056), .A(n10055), .B(n10054), .ZN(
        n10096) );
  AOI22_X1 U11165 ( .A1(n10084), .A2(n10096), .B1(n6082), .B2(n10082), .ZN(
        P1_U3477) );
  AND2_X1 U11166 ( .A1(n10057), .A2(n10070), .ZN(n10062) );
  INV_X1 U11167 ( .A(n10058), .ZN(n10059) );
  OAI21_X1 U11168 ( .B1(n10060), .B2(n10067), .A(n10059), .ZN(n10061) );
  NOR3_X1 U11169 ( .A1(n10063), .A2(n10062), .A3(n10061), .ZN(n10097) );
  INV_X1 U11170 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n10064) );
  AOI22_X1 U11171 ( .A1(n10084), .A2(n10097), .B1(n10064), .B2(n10082), .ZN(
        P1_U3480) );
  OAI211_X1 U11172 ( .C1(n10068), .C2(n10067), .A(n10066), .B(n10065), .ZN(
        n10069) );
  AOI21_X1 U11173 ( .B1(n10071), .B2(n10070), .A(n10069), .ZN(n10099) );
  AOI22_X1 U11174 ( .A1(n10084), .A2(n10099), .B1(n6117), .B2(n10082), .ZN(
        P1_U3483) );
  AOI21_X1 U11175 ( .B1(n10074), .B2(n10073), .A(n10072), .ZN(n10075) );
  OAI211_X1 U11176 ( .C1(n10078), .C2(n10077), .A(n10076), .B(n10075), .ZN(
        n10079) );
  AOI21_X1 U11177 ( .B1(n10081), .B2(n10080), .A(n10079), .ZN(n10101) );
  INV_X1 U11178 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n10083) );
  AOI22_X1 U11179 ( .A1(n10084), .A2(n10101), .B1(n10083), .B2(n10082), .ZN(
        P1_U3495) );
  AOI22_X1 U11180 ( .A1(n10102), .A2(n10086), .B1(n10085), .B2(n10100), .ZN(
        P1_U3523) );
  AOI22_X1 U11181 ( .A1(n10102), .A2(n10087), .B1(n6788), .B2(n10100), .ZN(
        P1_U3524) );
  AOI22_X1 U11182 ( .A1(n10102), .A2(n10088), .B1(n6790), .B2(n10100), .ZN(
        P1_U3525) );
  AOI22_X1 U11183 ( .A1(n10102), .A2(n10089), .B1(n6792), .B2(n10100), .ZN(
        P1_U3526) );
  INV_X1 U11184 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n10090) );
  AOI22_X1 U11185 ( .A1(n10102), .A2(n10091), .B1(n10090), .B2(n10100), .ZN(
        P1_U3527) );
  INV_X1 U11186 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n10092) );
  AOI22_X1 U11187 ( .A1(n10102), .A2(n10093), .B1(n10092), .B2(n10100), .ZN(
        P1_U3528) );
  AOI22_X1 U11188 ( .A1(n10102), .A2(n10094), .B1(n6043), .B2(n10100), .ZN(
        P1_U3529) );
  INV_X1 U11189 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n10095) );
  AOI22_X1 U11190 ( .A1(n10102), .A2(n10096), .B1(n10095), .B2(n10100), .ZN(
        P1_U3530) );
  AOI22_X1 U11191 ( .A1(n10102), .A2(n10097), .B1(n6097), .B2(n10100), .ZN(
        P1_U3531) );
  INV_X1 U11192 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n10098) );
  AOI22_X1 U11193 ( .A1(n10102), .A2(n10099), .B1(n10098), .B2(n10100), .ZN(
        P1_U3532) );
  AOI22_X1 U11194 ( .A1(n10102), .A2(n10101), .B1(n7608), .B2(n10100), .ZN(
        P1_U3536) );
  AOI22_X1 U11195 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(n10118), .B1(
        P2_REG3_REG_13__SCAN_IN), .B2(P2_U3151), .ZN(n10116) );
  AOI21_X1 U11196 ( .B1(n10105), .B2(n10104), .A(n10103), .ZN(n10113) );
  XOR2_X1 U11197 ( .A(n10107), .B(n10106), .Z(n10112) );
  AOI21_X1 U11198 ( .B1(n10110), .B2(n10109), .A(n10108), .ZN(n10111) );
  OAI222_X1 U11199 ( .A1(n10131), .A2(n10113), .B1(n10129), .B2(n10112), .C1(
        n10127), .C2(n10111), .ZN(n10114) );
  INV_X1 U11200 ( .A(n10114), .ZN(n10115) );
  OAI211_X1 U11201 ( .C1(n10136), .C2(n10117), .A(n10116), .B(n10115), .ZN(
        P2_U3195) );
  AOI22_X1 U11202 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(n10118), .B1(
        P2_REG3_REG_14__SCAN_IN), .B2(P2_U3151), .ZN(n10134) );
  AOI21_X1 U11203 ( .B1(n4581), .B2(n10120), .A(n10119), .ZN(n10130) );
  XOR2_X1 U11204 ( .A(n10122), .B(n10121), .Z(n10128) );
  AOI21_X1 U11205 ( .B1(n10125), .B2(n10124), .A(n10123), .ZN(n10126) );
  OAI222_X1 U11206 ( .A1(n10131), .A2(n10130), .B1(n10129), .B2(n10128), .C1(
        n10127), .C2(n10126), .ZN(n10132) );
  INV_X1 U11207 ( .A(n10132), .ZN(n10133) );
  OAI211_X1 U11208 ( .C1(n10136), .C2(n10135), .A(n10134), .B(n10133), .ZN(
        P2_U3196) );
  INV_X1 U11209 ( .A(n10137), .ZN(n10154) );
  OAI21_X1 U11210 ( .B1(n10140), .B2(n10139), .A(n10138), .ZN(n10161) );
  OAI22_X1 U11211 ( .A1(n10143), .A2(n10142), .B1(n10141), .B2(n10583), .ZN(
        n10153) );
  OAI21_X1 U11212 ( .B1(n10146), .B2(n10145), .A(n10144), .ZN(n10150) );
  AOI222_X1 U11213 ( .A1(n10151), .A2(n10150), .B1(n10149), .B2(n10148), .C1(
        n10147), .C2(n9025), .ZN(n10163) );
  INV_X1 U11214 ( .A(n10163), .ZN(n10152) );
  AOI211_X1 U11215 ( .C1(n10154), .C2(n10161), .A(n10153), .B(n10152), .ZN(
        n10158) );
  INV_X1 U11216 ( .A(n10155), .ZN(n10156) );
  AOI22_X1 U11217 ( .A1(n10161), .A2(n10156), .B1(n10159), .B2(
        P2_REG2_REG_2__SCAN_IN), .ZN(n10157) );
  OAI21_X1 U11218 ( .B1(n10159), .B2(n10158), .A(n10157), .ZN(P2_U3231) );
  INV_X1 U11219 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n10164) );
  AOI22_X1 U11220 ( .A1(n10161), .A2(n10192), .B1(n10198), .B2(n10160), .ZN(
        n10162) );
  AND2_X1 U11221 ( .A1(n10163), .A2(n10162), .ZN(n10203) );
  AOI22_X1 U11222 ( .A1(n10201), .A2(n10164), .B1(n10203), .B2(n10199), .ZN(
        P2_U3396) );
  INV_X1 U11223 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n10169) );
  AOI22_X1 U11224 ( .A1(n10166), .A2(n10192), .B1(n10198), .B2(n10165), .ZN(
        n10167) );
  AND2_X1 U11225 ( .A1(n10168), .A2(n10167), .ZN(n10204) );
  AOI22_X1 U11226 ( .A1(n10201), .A2(n10169), .B1(n10204), .B2(n10199), .ZN(
        P2_U3399) );
  INV_X1 U11227 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n10174) );
  NOR2_X1 U11228 ( .A1(n10170), .A2(n10187), .ZN(n10172) );
  AOI211_X1 U11229 ( .C1(n10192), .C2(n10173), .A(n10172), .B(n10171), .ZN(
        n10206) );
  AOI22_X1 U11230 ( .A1(n10201), .A2(n10174), .B1(n10206), .B2(n10199), .ZN(
        P2_U3402) );
  INV_X1 U11231 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n10180) );
  INV_X1 U11232 ( .A(n10175), .ZN(n10179) );
  OAI21_X1 U11233 ( .B1(n10177), .B2(n10187), .A(n10176), .ZN(n10178) );
  AOI21_X1 U11234 ( .B1(n10179), .B2(n10192), .A(n10178), .ZN(n10207) );
  AOI22_X1 U11235 ( .A1(n10201), .A2(n10180), .B1(n10207), .B2(n10199), .ZN(
        P2_U3408) );
  INV_X1 U11236 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n10186) );
  OAI22_X1 U11237 ( .A1(n10183), .A2(n10182), .B1(n10181), .B2(n10187), .ZN(
        n10184) );
  NOR2_X1 U11238 ( .A1(n10185), .A2(n10184), .ZN(n10208) );
  AOI22_X1 U11239 ( .A1(n10201), .A2(n10186), .B1(n10208), .B2(n10199), .ZN(
        P2_U3411) );
  NOR2_X1 U11240 ( .A1(n10188), .A2(n10187), .ZN(n10190) );
  AOI211_X1 U11241 ( .C1(n10192), .C2(n10191), .A(n10190), .B(n10189), .ZN(
        n10210) );
  AOI22_X1 U11242 ( .A1(n10201), .A2(n5444), .B1(n10210), .B2(n10199), .ZN(
        P2_U3414) );
  INV_X1 U11243 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n10200) );
  NOR2_X1 U11244 ( .A1(n10194), .A2(n10193), .ZN(n10196) );
  AOI211_X1 U11245 ( .C1(n10198), .C2(n10197), .A(n10196), .B(n10195), .ZN(
        n10212) );
  AOI22_X1 U11246 ( .A1(n10201), .A2(n10200), .B1(n10212), .B2(n10199), .ZN(
        P2_U3423) );
  AOI22_X1 U11247 ( .A1(n10213), .A2(n10203), .B1(n10202), .B2(n10211), .ZN(
        P2_U3461) );
  AOI22_X1 U11248 ( .A1(n10213), .A2(n10204), .B1(n5347), .B2(n10211), .ZN(
        P2_U3462) );
  AOI22_X1 U11249 ( .A1(n10213), .A2(n10206), .B1(n10205), .B2(n10211), .ZN(
        P2_U3463) );
  AOI22_X1 U11250 ( .A1(n10213), .A2(n10207), .B1(n7146), .B2(n10211), .ZN(
        P2_U3465) );
  AOI22_X1 U11251 ( .A1(n10213), .A2(n10208), .B1(n7136), .B2(n10211), .ZN(
        P2_U3466) );
  AOI22_X1 U11252 ( .A1(n10213), .A2(n10210), .B1(n10209), .B2(n10211), .ZN(
        P2_U3467) );
  AOI22_X1 U11253 ( .A1(n10213), .A2(n10212), .B1(n5497), .B2(n10211), .ZN(
        P2_U3470) );
  NAND3_X1 U11254 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(P1_ADDR_REG_0__SCAN_IN), 
        .A3(P2_ADDR_REG_0__SCAN_IN), .ZN(n10216) );
  AND2_X1 U11255 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .ZN(n10214) );
  NOR2_X1 U11256 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(n10214), .ZN(n10215) );
  INV_X1 U11257 ( .A(n10215), .ZN(n10232) );
  NAND2_X1 U11258 ( .A1(n10217), .A2(n10216), .ZN(n10231) );
  OAI222_X1 U11259 ( .A1(n10217), .A2(n10216), .B1(n10217), .B2(n10232), .C1(
        n10215), .C2(n10231), .ZN(ADD_1068_U5) );
  XOR2_X1 U11260 ( .A(P1_ADDR_REG_0__SCAN_IN), .B(P2_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1068_U46) );
  NOR2_X1 U11261 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n10218) );
  AOI21_X1 U11262 ( .B1(P1_ADDR_REG_17__SCAN_IN), .B2(P2_ADDR_REG_17__SCAN_IN), 
        .A(n10218), .ZN(n10239) );
  NOR2_X1 U11263 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n10219) );
  AOI21_X1 U11264 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(P2_ADDR_REG_16__SCAN_IN), 
        .A(n10219), .ZN(n10242) );
  NOR2_X1 U11265 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n10220) );
  AOI21_X1 U11266 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(P2_ADDR_REG_15__SCAN_IN), 
        .A(n10220), .ZN(n10245) );
  NOR2_X1 U11267 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n10221) );
  AOI21_X1 U11268 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(P2_ADDR_REG_14__SCAN_IN), 
        .A(n10221), .ZN(n10248) );
  NOR2_X1 U11269 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n10222) );
  AOI21_X1 U11270 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(P2_ADDR_REG_13__SCAN_IN), 
        .A(n10222), .ZN(n10251) );
  NOR2_X1 U11271 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n10223) );
  AOI21_X1 U11272 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(P2_ADDR_REG_12__SCAN_IN), 
        .A(n10223), .ZN(n10254) );
  NOR2_X1 U11273 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(P1_ADDR_REG_11__SCAN_IN), 
        .ZN(n10224) );
  AOI21_X1 U11274 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(P2_ADDR_REG_11__SCAN_IN), 
        .A(n10224), .ZN(n10257) );
  NOR2_X1 U11275 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(P1_ADDR_REG_10__SCAN_IN), 
        .ZN(n10225) );
  AOI21_X1 U11276 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(P2_ADDR_REG_10__SCAN_IN), 
        .A(n10225), .ZN(n10260) );
  NOR2_X1 U11277 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(P1_ADDR_REG_9__SCAN_IN), 
        .ZN(n10226) );
  AOI21_X1 U11278 ( .B1(P1_ADDR_REG_9__SCAN_IN), .B2(P2_ADDR_REG_9__SCAN_IN), 
        .A(n10226), .ZN(n10645) );
  NOR2_X1 U11279 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(P1_ADDR_REG_8__SCAN_IN), 
        .ZN(n10227) );
  AOI21_X1 U11280 ( .B1(P1_ADDR_REG_8__SCAN_IN), .B2(P2_ADDR_REG_8__SCAN_IN), 
        .A(n10227), .ZN(n10657) );
  NOR2_X1 U11281 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(P1_ADDR_REG_7__SCAN_IN), 
        .ZN(n10228) );
  AOI21_X1 U11282 ( .B1(P1_ADDR_REG_7__SCAN_IN), .B2(P2_ADDR_REG_7__SCAN_IN), 
        .A(n10228), .ZN(n10654) );
  NOR2_X1 U11283 ( .A1(P1_ADDR_REG_6__SCAN_IN), .A2(P2_ADDR_REG_6__SCAN_IN), 
        .ZN(n10229) );
  AOI21_X1 U11284 ( .B1(P2_ADDR_REG_6__SCAN_IN), .B2(P1_ADDR_REG_6__SCAN_IN), 
        .A(n10229), .ZN(n10660) );
  NOR2_X1 U11285 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(P1_ADDR_REG_5__SCAN_IN), 
        .ZN(n10230) );
  AOI21_X1 U11286 ( .B1(P1_ADDR_REG_5__SCAN_IN), .B2(P2_ADDR_REG_5__SCAN_IN), 
        .A(n10230), .ZN(n10651) );
  NAND2_X1 U11287 ( .A1(n10232), .A2(n10231), .ZN(n10648) );
  NAND2_X1 U11288 ( .A1(P1_ADDR_REG_2__SCAN_IN), .A2(P2_ADDR_REG_2__SCAN_IN), 
        .ZN(n10233) );
  OAI21_X1 U11289 ( .B1(P1_ADDR_REG_2__SCAN_IN), .B2(P2_ADDR_REG_2__SCAN_IN), 
        .A(n10233), .ZN(n10647) );
  NOR2_X1 U11290 ( .A1(n10648), .A2(n10647), .ZN(n10646) );
  AOI21_X1 U11291 ( .B1(P2_ADDR_REG_2__SCAN_IN), .B2(P1_ADDR_REG_2__SCAN_IN), 
        .A(n10646), .ZN(n10663) );
  NAND2_X1 U11292 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n10234) );
  OAI21_X1 U11293 ( .B1(P1_ADDR_REG_3__SCAN_IN), .B2(P2_ADDR_REG_3__SCAN_IN), 
        .A(n10234), .ZN(n10662) );
  NOR2_X1 U11294 ( .A1(n10663), .A2(n10662), .ZN(n10661) );
  AOI21_X1 U11295 ( .B1(P2_ADDR_REG_3__SCAN_IN), .B2(P1_ADDR_REG_3__SCAN_IN), 
        .A(n10661), .ZN(n10666) );
  NOR2_X1 U11296 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n10235) );
  AOI21_X1 U11297 ( .B1(P2_ADDR_REG_4__SCAN_IN), .B2(P1_ADDR_REG_4__SCAN_IN), 
        .A(n10235), .ZN(n10665) );
  NAND2_X1 U11298 ( .A1(n10666), .A2(n10665), .ZN(n10664) );
  OAI21_X1 U11299 ( .B1(P1_ADDR_REG_4__SCAN_IN), .B2(P2_ADDR_REG_4__SCAN_IN), 
        .A(n10664), .ZN(n10650) );
  NAND2_X1 U11300 ( .A1(n10651), .A2(n10650), .ZN(n10649) );
  OAI21_X1 U11301 ( .B1(P2_ADDR_REG_5__SCAN_IN), .B2(P1_ADDR_REG_5__SCAN_IN), 
        .A(n10649), .ZN(n10659) );
  NAND2_X1 U11302 ( .A1(n10660), .A2(n10659), .ZN(n10658) );
  OAI21_X1 U11303 ( .B1(P1_ADDR_REG_6__SCAN_IN), .B2(P2_ADDR_REG_6__SCAN_IN), 
        .A(n10658), .ZN(n10653) );
  NAND2_X1 U11304 ( .A1(n10654), .A2(n10653), .ZN(n10652) );
  OAI21_X1 U11305 ( .B1(P2_ADDR_REG_7__SCAN_IN), .B2(P1_ADDR_REG_7__SCAN_IN), 
        .A(n10652), .ZN(n10656) );
  NAND2_X1 U11306 ( .A1(n10657), .A2(n10656), .ZN(n10655) );
  OAI21_X1 U11307 ( .B1(P2_ADDR_REG_8__SCAN_IN), .B2(P1_ADDR_REG_8__SCAN_IN), 
        .A(n10655), .ZN(n10644) );
  NAND2_X1 U11308 ( .A1(n10645), .A2(n10644), .ZN(n10643) );
  OAI21_X1 U11309 ( .B1(P2_ADDR_REG_9__SCAN_IN), .B2(P1_ADDR_REG_9__SCAN_IN), 
        .A(n10643), .ZN(n10259) );
  NAND2_X1 U11310 ( .A1(n10260), .A2(n10259), .ZN(n10258) );
  OAI21_X1 U11311 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(P1_ADDR_REG_10__SCAN_IN), 
        .A(n10258), .ZN(n10256) );
  NAND2_X1 U11312 ( .A1(n10257), .A2(n10256), .ZN(n10255) );
  OAI21_X1 U11313 ( .B1(P2_ADDR_REG_11__SCAN_IN), .B2(P1_ADDR_REG_11__SCAN_IN), 
        .A(n10255), .ZN(n10253) );
  NAND2_X1 U11314 ( .A1(n10254), .A2(n10253), .ZN(n10252) );
  OAI21_X1 U11315 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(P1_ADDR_REG_12__SCAN_IN), 
        .A(n10252), .ZN(n10250) );
  NAND2_X1 U11316 ( .A1(n10251), .A2(n10250), .ZN(n10249) );
  OAI21_X1 U11317 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(P1_ADDR_REG_13__SCAN_IN), 
        .A(n10249), .ZN(n10247) );
  NAND2_X1 U11318 ( .A1(n10248), .A2(n10247), .ZN(n10246) );
  OAI21_X1 U11319 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(P1_ADDR_REG_14__SCAN_IN), 
        .A(n10246), .ZN(n10244) );
  NAND2_X1 U11320 ( .A1(n10245), .A2(n10244), .ZN(n10243) );
  OAI21_X1 U11321 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(P1_ADDR_REG_15__SCAN_IN), 
        .A(n10243), .ZN(n10241) );
  NAND2_X1 U11322 ( .A1(n10242), .A2(n10241), .ZN(n10240) );
  OAI21_X1 U11323 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(P1_ADDR_REG_16__SCAN_IN), 
        .A(n10240), .ZN(n10238) );
  NAND2_X1 U11324 ( .A1(n10239), .A2(n10238), .ZN(n10237) );
  OAI21_X1 U11325 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(P1_ADDR_REG_17__SCAN_IN), 
        .A(n10237), .ZN(n10261) );
  NAND2_X1 U11326 ( .A1(n10262), .A2(n10261), .ZN(n10263) );
  OAI21_X1 U11327 ( .B1(n10261), .B2(n10262), .A(n10263), .ZN(n10236) );
  XNOR2_X1 U11328 ( .A(n10236), .B(P2_ADDR_REG_18__SCAN_IN), .ZN(ADD_1068_U55)
         );
  OAI21_X1 U11329 ( .B1(n10239), .B2(n10238), .A(n10237), .ZN(ADD_1068_U56) );
  OAI21_X1 U11330 ( .B1(n10242), .B2(n10241), .A(n10240), .ZN(ADD_1068_U57) );
  OAI21_X1 U11331 ( .B1(n10245), .B2(n10244), .A(n10243), .ZN(ADD_1068_U58) );
  OAI21_X1 U11332 ( .B1(n10248), .B2(n10247), .A(n10246), .ZN(ADD_1068_U59) );
  OAI21_X1 U11333 ( .B1(n10251), .B2(n10250), .A(n10249), .ZN(ADD_1068_U60) );
  OAI21_X1 U11334 ( .B1(n10254), .B2(n10253), .A(n10252), .ZN(ADD_1068_U61) );
  OAI21_X1 U11335 ( .B1(n10257), .B2(n10256), .A(n10255), .ZN(ADD_1068_U62) );
  OAI21_X1 U11336 ( .B1(n10260), .B2(n10259), .A(n10258), .ZN(ADD_1068_U63) );
  NOR2_X1 U11337 ( .A1(n10262), .A2(n10261), .ZN(n10264) );
  OAI21_X1 U11338 ( .B1(P2_ADDR_REG_18__SCAN_IN), .B2(n10264), .A(n10263), 
        .ZN(n10642) );
  OAI22_X1 U11339 ( .A1(P1_IR_REG_17__SCAN_IN), .A2(keyinput_g107), .B1(
        P2_REG3_REG_21__SCAN_IN), .B2(keyinput_g45), .ZN(n10265) );
  AOI221_X1 U11340 ( .B1(P1_IR_REG_17__SCAN_IN), .B2(keyinput_g107), .C1(
        keyinput_g45), .C2(P2_REG3_REG_21__SCAN_IN), .A(n10265), .ZN(n10272)
         );
  OAI22_X1 U11341 ( .A1(P1_IR_REG_14__SCAN_IN), .A2(keyinput_g104), .B1(
        keyinput_g6), .B2(SI_26_), .ZN(n10266) );
  AOI221_X1 U11342 ( .B1(P1_IR_REG_14__SCAN_IN), .B2(keyinput_g104), .C1(
        SI_26_), .C2(keyinput_g6), .A(n10266), .ZN(n10271) );
  OAI22_X1 U11343 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(keyinput_g112), .B1(
        P1_IR_REG_3__SCAN_IN), .B2(keyinput_g93), .ZN(n10267) );
  AOI221_X1 U11344 ( .B1(P1_IR_REG_22__SCAN_IN), .B2(keyinput_g112), .C1(
        keyinput_g93), .C2(P1_IR_REG_3__SCAN_IN), .A(n10267), .ZN(n10270) );
  OAI22_X1 U11345 ( .A1(SI_20_), .A2(keyinput_g12), .B1(
        P2_REG3_REG_22__SCAN_IN), .B2(keyinput_g57), .ZN(n10268) );
  AOI221_X1 U11346 ( .B1(SI_20_), .B2(keyinput_g12), .C1(keyinput_g57), .C2(
        P2_REG3_REG_22__SCAN_IN), .A(n10268), .ZN(n10269) );
  NAND4_X1 U11347 ( .A1(n10272), .A2(n10271), .A3(n10270), .A4(n10269), .ZN(
        n10301) );
  OAI22_X1 U11348 ( .A1(P1_IR_REG_18__SCAN_IN), .A2(keyinput_g108), .B1(SI_9_), 
        .B2(keyinput_g23), .ZN(n10273) );
  AOI221_X1 U11349 ( .B1(P1_IR_REG_18__SCAN_IN), .B2(keyinput_g108), .C1(
        keyinput_g23), .C2(SI_9_), .A(n10273), .ZN(n10280) );
  OAI22_X1 U11350 ( .A1(SI_8_), .A2(keyinput_g24), .B1(P2_REG3_REG_20__SCAN_IN), .B2(keyinput_g55), .ZN(n10274) );
  AOI221_X1 U11351 ( .B1(SI_8_), .B2(keyinput_g24), .C1(keyinput_g55), .C2(
        P2_REG3_REG_20__SCAN_IN), .A(n10274), .ZN(n10279) );
  OAI22_X1 U11352 ( .A1(P1_IR_REG_2__SCAN_IN), .A2(keyinput_g92), .B1(
        keyinput_g89), .B2(P2_DATAO_REG_7__SCAN_IN), .ZN(n10275) );
  AOI221_X1 U11353 ( .B1(P1_IR_REG_2__SCAN_IN), .B2(keyinput_g92), .C1(
        P2_DATAO_REG_7__SCAN_IN), .C2(keyinput_g89), .A(n10275), .ZN(n10278)
         );
  OAI22_X1 U11354 ( .A1(SI_19_), .A2(keyinput_g13), .B1(keyinput_g85), .B2(
        P2_DATAO_REG_11__SCAN_IN), .ZN(n10276) );
  AOI221_X1 U11355 ( .B1(SI_19_), .B2(keyinput_g13), .C1(
        P2_DATAO_REG_11__SCAN_IN), .C2(keyinput_g85), .A(n10276), .ZN(n10277)
         );
  NAND4_X1 U11356 ( .A1(n10280), .A2(n10279), .A3(n10278), .A4(n10277), .ZN(
        n10300) );
  OAI22_X1 U11357 ( .A1(P1_IR_REG_12__SCAN_IN), .A2(keyinput_g102), .B1(
        P2_REG3_REG_18__SCAN_IN), .B2(keyinput_g60), .ZN(n10281) );
  AOI221_X1 U11358 ( .B1(P1_IR_REG_12__SCAN_IN), .B2(keyinput_g102), .C1(
        keyinput_g60), .C2(P2_REG3_REG_18__SCAN_IN), .A(n10281), .ZN(n10288)
         );
  OAI22_X1 U11359 ( .A1(SI_25_), .A2(keyinput_g7), .B1(SI_12_), .B2(
        keyinput_g20), .ZN(n10282) );
  AOI221_X1 U11360 ( .B1(SI_25_), .B2(keyinput_g7), .C1(keyinput_g20), .C2(
        SI_12_), .A(n10282), .ZN(n10287) );
  OAI22_X1 U11361 ( .A1(P1_IR_REG_24__SCAN_IN), .A2(keyinput_g114), .B1(SI_13_), .B2(keyinput_g19), .ZN(n10283) );
  AOI221_X1 U11362 ( .B1(P1_IR_REG_24__SCAN_IN), .B2(keyinput_g114), .C1(
        keyinput_g19), .C2(SI_13_), .A(n10283), .ZN(n10286) );
  OAI22_X1 U11363 ( .A1(P2_DATAO_REG_23__SCAN_IN), .A2(keyinput_g73), .B1(
        SI_0_), .B2(keyinput_g32), .ZN(n10284) );
  AOI221_X1 U11364 ( .B1(P2_DATAO_REG_23__SCAN_IN), .B2(keyinput_g73), .C1(
        keyinput_g32), .C2(SI_0_), .A(n10284), .ZN(n10285) );
  NAND4_X1 U11365 ( .A1(n10288), .A2(n10287), .A3(n10286), .A4(n10285), .ZN(
        n10299) );
  OAI22_X1 U11366 ( .A1(SI_16_), .A2(keyinput_g16), .B1(keyinput_g48), .B2(
        P2_REG3_REG_16__SCAN_IN), .ZN(n10289) );
  AOI221_X1 U11367 ( .B1(SI_16_), .B2(keyinput_g16), .C1(
        P2_REG3_REG_16__SCAN_IN), .C2(keyinput_g48), .A(n10289), .ZN(n10297)
         );
  OAI22_X1 U11368 ( .A1(P2_B_REG_SCAN_IN), .A2(keyinput_g64), .B1(keyinput_g42), .B2(P2_REG3_REG_28__SCAN_IN), .ZN(n10290) );
  AOI221_X1 U11369 ( .B1(P2_B_REG_SCAN_IN), .B2(keyinput_g64), .C1(
        P2_REG3_REG_28__SCAN_IN), .C2(keyinput_g42), .A(n10290), .ZN(n10296)
         );
  OAI22_X1 U11370 ( .A1(P1_IR_REG_21__SCAN_IN), .A2(keyinput_g111), .B1(SI_6_), 
        .B2(keyinput_g26), .ZN(n10291) );
  AOI221_X1 U11371 ( .B1(P1_IR_REG_21__SCAN_IN), .B2(keyinput_g111), .C1(
        keyinput_g26), .C2(SI_6_), .A(n10291), .ZN(n10295) );
  OAI22_X1 U11372 ( .A1(n10293), .A2(keyinput_g82), .B1(keyinput_g116), .B2(
        P1_IR_REG_26__SCAN_IN), .ZN(n10292) );
  AOI221_X1 U11373 ( .B1(n10293), .B2(keyinput_g82), .C1(P1_IR_REG_26__SCAN_IN), .C2(keyinput_g116), .A(n10292), .ZN(n10294) );
  NAND4_X1 U11374 ( .A1(n10297), .A2(n10296), .A3(n10295), .A4(n10294), .ZN(
        n10298) );
  NOR4_X1 U11375 ( .A1(n10301), .A2(n10300), .A3(n10299), .A4(n10298), .ZN(
        n10638) );
  OAI22_X1 U11376 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(keyinput_g110), .B1(
        keyinput_g11), .B2(SI_21_), .ZN(n10302) );
  AOI221_X1 U11377 ( .B1(P1_IR_REG_20__SCAN_IN), .B2(keyinput_g110), .C1(
        SI_21_), .C2(keyinput_g11), .A(n10302), .ZN(n10309) );
  OAI22_X1 U11378 ( .A1(P2_DATAO_REG_27__SCAN_IN), .A2(keyinput_g69), .B1(
        P2_DATAO_REG_28__SCAN_IN), .B2(keyinput_g68), .ZN(n10303) );
  AOI221_X1 U11379 ( .B1(P2_DATAO_REG_27__SCAN_IN), .B2(keyinput_g69), .C1(
        keyinput_g68), .C2(P2_DATAO_REG_28__SCAN_IN), .A(n10303), .ZN(n10308)
         );
  OAI22_X1 U11380 ( .A1(P1_IR_REG_23__SCAN_IN), .A2(keyinput_g113), .B1(
        keyinput_g29), .B2(SI_3_), .ZN(n10304) );
  AOI221_X1 U11381 ( .B1(P1_IR_REG_23__SCAN_IN), .B2(keyinput_g113), .C1(SI_3_), .C2(keyinput_g29), .A(n10304), .ZN(n10307) );
  OAI22_X1 U11382 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(keyinput_g61), .B1(
        keyinput_g52), .B2(P2_REG3_REG_4__SCAN_IN), .ZN(n10305) );
  AOI221_X1 U11383 ( .B1(P2_REG3_REG_6__SCAN_IN), .B2(keyinput_g61), .C1(
        P2_REG3_REG_4__SCAN_IN), .C2(keyinput_g52), .A(n10305), .ZN(n10306) );
  NAND4_X1 U11384 ( .A1(n10309), .A2(n10308), .A3(n10307), .A4(n10306), .ZN(
        n10437) );
  OAI22_X1 U11385 ( .A1(SI_23_), .A2(keyinput_g9), .B1(keyinput_g37), .B2(
        P2_REG3_REG_14__SCAN_IN), .ZN(n10310) );
  AOI221_X1 U11386 ( .B1(SI_23_), .B2(keyinput_g9), .C1(
        P2_REG3_REG_14__SCAN_IN), .C2(keyinput_g37), .A(n10310), .ZN(n10335)
         );
  INV_X1 U11387 ( .A(SI_14_), .ZN(n10527) );
  OAI22_X1 U11388 ( .A1(P1_D_REG_5__SCAN_IN), .A2(keyinput_g127), .B1(
        P2_REG3_REG_12__SCAN_IN), .B2(keyinput_g46), .ZN(n10311) );
  AOI221_X1 U11389 ( .B1(P1_D_REG_5__SCAN_IN), .B2(keyinput_g127), .C1(
        keyinput_g46), .C2(P2_REG3_REG_12__SCAN_IN), .A(n10311), .ZN(n10314)
         );
  OAI22_X1 U11390 ( .A1(P2_REG3_REG_26__SCAN_IN), .A2(keyinput_g62), .B1(
        P2_REG3_REG_24__SCAN_IN), .B2(keyinput_g51), .ZN(n10312) );
  AOI221_X1 U11391 ( .B1(P2_REG3_REG_26__SCAN_IN), .B2(keyinput_g62), .C1(
        keyinput_g51), .C2(P2_REG3_REG_24__SCAN_IN), .A(n10312), .ZN(n10313)
         );
  OAI211_X1 U11392 ( .C1(n10527), .C2(keyinput_g18), .A(n10314), .B(n10313), 
        .ZN(n10315) );
  AOI21_X1 U11393 ( .B1(n10527), .B2(keyinput_g18), .A(n10315), .ZN(n10334) );
  AOI22_X1 U11394 ( .A1(SI_30_), .A2(keyinput_g2), .B1(
        P2_DATAO_REG_20__SCAN_IN), .B2(keyinput_g76), .ZN(n10316) );
  OAI221_X1 U11395 ( .B1(SI_30_), .B2(keyinput_g2), .C1(
        P2_DATAO_REG_20__SCAN_IN), .C2(keyinput_g76), .A(n10316), .ZN(n10323)
         );
  AOI22_X1 U11396 ( .A1(P2_REG3_REG_15__SCAN_IN), .A2(keyinput_g63), .B1(
        SI_24_), .B2(keyinput_g8), .ZN(n10317) );
  OAI221_X1 U11397 ( .B1(P2_REG3_REG_15__SCAN_IN), .B2(keyinput_g63), .C1(
        SI_24_), .C2(keyinput_g8), .A(n10317), .ZN(n10322) );
  AOI22_X1 U11398 ( .A1(P2_DATAO_REG_24__SCAN_IN), .A2(keyinput_g72), .B1(
        P1_IR_REG_8__SCAN_IN), .B2(keyinput_g98), .ZN(n10318) );
  OAI221_X1 U11399 ( .B1(P2_DATAO_REG_24__SCAN_IN), .B2(keyinput_g72), .C1(
        P1_IR_REG_8__SCAN_IN), .C2(keyinput_g98), .A(n10318), .ZN(n10321) );
  AOI22_X1 U11400 ( .A1(SI_15_), .A2(keyinput_g17), .B1(P1_IR_REG_11__SCAN_IN), 
        .B2(keyinput_g101), .ZN(n10319) );
  OAI221_X1 U11401 ( .B1(SI_15_), .B2(keyinput_g17), .C1(P1_IR_REG_11__SCAN_IN), .C2(keyinput_g101), .A(n10319), .ZN(n10320) );
  NOR4_X1 U11402 ( .A1(n10323), .A2(n10322), .A3(n10321), .A4(n10320), .ZN(
        n10333) );
  AOI22_X1 U11403 ( .A1(P2_REG3_REG_27__SCAN_IN), .A2(keyinput_g36), .B1(
        P2_STATE_REG_SCAN_IN), .B2(keyinput_g34), .ZN(n10324) );
  OAI221_X1 U11404 ( .B1(P2_REG3_REG_27__SCAN_IN), .B2(keyinput_g36), .C1(
        P2_STATE_REG_SCAN_IN), .C2(keyinput_g34), .A(n10324), .ZN(n10331) );
  AOI22_X1 U11405 ( .A1(P2_REG3_REG_13__SCAN_IN), .A2(keyinput_g56), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(keyinput_g88), .ZN(n10325) );
  OAI221_X1 U11406 ( .B1(P2_REG3_REG_13__SCAN_IN), .B2(keyinput_g56), .C1(
        P2_DATAO_REG_8__SCAN_IN), .C2(keyinput_g88), .A(n10325), .ZN(n10330)
         );
  AOI22_X1 U11407 ( .A1(P2_WR_REG_SCAN_IN), .A2(keyinput_g0), .B1(
        P2_DATAO_REG_31__SCAN_IN), .B2(keyinput_g65), .ZN(n10326) );
  OAI221_X1 U11408 ( .B1(P2_WR_REG_SCAN_IN), .B2(keyinput_g0), .C1(
        P2_DATAO_REG_31__SCAN_IN), .C2(keyinput_g65), .A(n10326), .ZN(n10329)
         );
  AOI22_X1 U11409 ( .A1(P2_DATAO_REG_22__SCAN_IN), .A2(keyinput_g74), .B1(
        P1_IR_REG_15__SCAN_IN), .B2(keyinput_g105), .ZN(n10327) );
  OAI221_X1 U11410 ( .B1(P2_DATAO_REG_22__SCAN_IN), .B2(keyinput_g74), .C1(
        P1_IR_REG_15__SCAN_IN), .C2(keyinput_g105), .A(n10327), .ZN(n10328) );
  NOR4_X1 U11411 ( .A1(n10331), .A2(n10330), .A3(n10329), .A4(n10328), .ZN(
        n10332) );
  NAND4_X1 U11412 ( .A1(n10335), .A2(n10334), .A3(n10333), .A4(n10332), .ZN(
        n10436) );
  AOI22_X1 U11413 ( .A1(n10526), .A2(keyinput_g71), .B1(keyinput_g120), .B2(
        n5869), .ZN(n10336) );
  OAI221_X1 U11414 ( .B1(n10526), .B2(keyinput_g71), .C1(n5869), .C2(
        keyinput_g120), .A(n10336), .ZN(n10345) );
  AOI22_X1 U11415 ( .A1(n10338), .A2(keyinput_g67), .B1(n10511), .B2(
        keyinput_g15), .ZN(n10337) );
  OAI221_X1 U11416 ( .B1(n10338), .B2(keyinput_g67), .C1(n10511), .C2(
        keyinput_g15), .A(n10337), .ZN(n10344) );
  XNOR2_X1 U11417 ( .A(P2_REG3_REG_3__SCAN_IN), .B(keyinput_g40), .ZN(n10342)
         );
  XNOR2_X1 U11418 ( .A(P1_IR_REG_19__SCAN_IN), .B(keyinput_g109), .ZN(n10341)
         );
  XNOR2_X1 U11419 ( .A(P1_IR_REG_9__SCAN_IN), .B(keyinput_g99), .ZN(n10340) );
  XNOR2_X1 U11420 ( .A(P1_IR_REG_4__SCAN_IN), .B(keyinput_g94), .ZN(n10339) );
  NAND4_X1 U11421 ( .A1(n10342), .A2(n10341), .A3(n10340), .A4(n10339), .ZN(
        n10343) );
  NOR3_X1 U11422 ( .A1(n10345), .A2(n10344), .A3(n10343), .ZN(n10382) );
  AOI22_X1 U11423 ( .A1(n10347), .A2(keyinput_g79), .B1(keyinput_g44), .B2(
        n6992), .ZN(n10346) );
  OAI221_X1 U11424 ( .B1(n10347), .B2(keyinput_g79), .C1(n6992), .C2(
        keyinput_g44), .A(n10346), .ZN(n10355) );
  INV_X1 U11425 ( .A(SI_11_), .ZN(n10515) );
  INV_X1 U11426 ( .A(SI_18_), .ZN(n10545) );
  AOI22_X1 U11427 ( .A1(n10515), .A2(keyinput_g21), .B1(n10545), .B2(
        keyinput_g14), .ZN(n10348) );
  OAI221_X1 U11428 ( .B1(n10515), .B2(keyinput_g21), .C1(n10545), .C2(
        keyinput_g14), .A(n10348), .ZN(n10354) );
  INV_X1 U11429 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n10532) );
  AOI22_X1 U11430 ( .A1(n5153), .A2(keyinput_g35), .B1(n10532), .B2(
        keyinput_g122), .ZN(n10349) );
  OAI221_X1 U11431 ( .B1(n5153), .B2(keyinput_g35), .C1(n10532), .C2(
        keyinput_g122), .A(n10349), .ZN(n10353) );
  XNOR2_X1 U11432 ( .A(P2_REG3_REG_25__SCAN_IN), .B(keyinput_g47), .ZN(n10351)
         );
  XNOR2_X1 U11433 ( .A(SI_2_), .B(keyinput_g30), .ZN(n10350) );
  NAND2_X1 U11434 ( .A1(n10351), .A2(n10350), .ZN(n10352) );
  NOR4_X1 U11435 ( .A1(n10355), .A2(n10354), .A3(n10353), .A4(n10352), .ZN(
        n10381) );
  AOI22_X1 U11436 ( .A1(n10553), .A2(keyinput_g126), .B1(keyinput_g49), .B2(
        n5151), .ZN(n10356) );
  OAI221_X1 U11437 ( .B1(n10553), .B2(keyinput_g126), .C1(n5151), .C2(
        keyinput_g49), .A(n10356), .ZN(n10366) );
  AOI22_X1 U11438 ( .A1(n10359), .A2(keyinput_g4), .B1(keyinput_g3), .B2(
        n10358), .ZN(n10357) );
  OAI221_X1 U11439 ( .B1(n10359), .B2(keyinput_g4), .C1(n10358), .C2(
        keyinput_g3), .A(n10357), .ZN(n10365) );
  XOR2_X1 U11440 ( .A(n5155), .B(keyinput_g53), .Z(n10363) );
  XNOR2_X1 U11441 ( .A(SI_4_), .B(keyinput_g28), .ZN(n10362) );
  XNOR2_X1 U11442 ( .A(P2_REG3_REG_8__SCAN_IN), .B(keyinput_g43), .ZN(n10361)
         );
  XNOR2_X1 U11443 ( .A(P1_IR_REG_31__SCAN_IN), .B(keyinput_g121), .ZN(n10360)
         );
  NAND4_X1 U11444 ( .A1(n10363), .A2(n10362), .A3(n10361), .A4(n10360), .ZN(
        n10364) );
  NOR3_X1 U11445 ( .A1(n10366), .A2(n10365), .A3(n10364), .ZN(n10380) );
  AOI22_X1 U11446 ( .A1(n6068), .A2(keyinput_g97), .B1(keyinput_g118), .B2(
        n5033), .ZN(n10367) );
  OAI221_X1 U11447 ( .B1(n6068), .B2(keyinput_g97), .C1(n5033), .C2(
        keyinput_g118), .A(n10367), .ZN(n10378) );
  AOI22_X1 U11448 ( .A1(n10369), .A2(keyinput_g87), .B1(keyinput_g27), .B2(
        n10574), .ZN(n10368) );
  OAI221_X1 U11449 ( .B1(n10369), .B2(keyinput_g87), .C1(n10574), .C2(
        keyinput_g27), .A(n10368), .ZN(n10377) );
  AOI22_X1 U11450 ( .A1(n10372), .A2(keyinput_g66), .B1(n10371), .B2(
        keyinput_g86), .ZN(n10370) );
  OAI221_X1 U11451 ( .B1(n10372), .B2(keyinput_g66), .C1(n10371), .C2(
        keyinput_g86), .A(n10370), .ZN(n10376) );
  XNOR2_X1 U11452 ( .A(P1_IR_REG_5__SCAN_IN), .B(keyinput_g95), .ZN(n10374) );
  XNOR2_X1 U11453 ( .A(SI_22_), .B(keyinput_g10), .ZN(n10373) );
  NAND2_X1 U11454 ( .A1(n10374), .A2(n10373), .ZN(n10375) );
  NOR4_X1 U11455 ( .A1(n10378), .A2(n10377), .A3(n10376), .A4(n10375), .ZN(
        n10379) );
  NAND4_X1 U11456 ( .A1(n10382), .A2(n10381), .A3(n10380), .A4(n10379), .ZN(
        n10435) );
  AOI22_X1 U11457 ( .A1(n5203), .A2(keyinput_g31), .B1(n10586), .B2(
        keyinput_g81), .ZN(n10383) );
  OAI221_X1 U11458 ( .B1(n5203), .B2(keyinput_g31), .C1(n10586), .C2(
        keyinput_g81), .A(n10383), .ZN(n10393) );
  INV_X1 U11459 ( .A(SI_31_), .ZN(n10596) );
  AOI22_X1 U11460 ( .A1(n10596), .A2(keyinput_g1), .B1(n10385), .B2(
        keyinput_g39), .ZN(n10384) );
  OAI221_X1 U11461 ( .B1(n10596), .B2(keyinput_g1), .C1(n10385), .C2(
        keyinput_g39), .A(n10384), .ZN(n10392) );
  INV_X1 U11462 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n10611) );
  AOI22_X1 U11463 ( .A1(n10387), .A2(keyinput_g80), .B1(keyinput_g38), .B2(
        n10611), .ZN(n10386) );
  OAI221_X1 U11464 ( .B1(n10387), .B2(keyinput_g80), .C1(n10611), .C2(
        keyinput_g38), .A(n10386), .ZN(n10391) );
  AOI22_X1 U11465 ( .A1(n6134), .A2(keyinput_g100), .B1(keyinput_g75), .B2(
        n10389), .ZN(n10388) );
  OAI221_X1 U11466 ( .B1(n6134), .B2(keyinput_g100), .C1(n10389), .C2(
        keyinput_g75), .A(n10388), .ZN(n10390) );
  NOR4_X1 U11467 ( .A1(n10393), .A2(n10392), .A3(n10391), .A4(n10390), .ZN(
        n10433) );
  AOI22_X1 U11468 ( .A1(n6067), .A2(keyinput_g96), .B1(keyinput_g78), .B2(
        n10395), .ZN(n10394) );
  OAI221_X1 U11469 ( .B1(n6067), .B2(keyinput_g96), .C1(n10395), .C2(
        keyinput_g78), .A(n10394), .ZN(n10404) );
  AOI22_X1 U11470 ( .A1(n10530), .A2(keyinput_g70), .B1(n10397), .B2(
        keyinput_g90), .ZN(n10396) );
  OAI221_X1 U11471 ( .B1(n10530), .B2(keyinput_g70), .C1(n10397), .C2(
        keyinput_g90), .A(n10396), .ZN(n10403) );
  XOR2_X1 U11472 ( .A(n4731), .B(keyinput_g91), .Z(n10401) );
  XNOR2_X1 U11473 ( .A(P1_IR_REG_13__SCAN_IN), .B(keyinput_g103), .ZN(n10400)
         );
  XNOR2_X1 U11474 ( .A(SI_27_), .B(keyinput_g5), .ZN(n10399) );
  XNOR2_X1 U11475 ( .A(P1_IR_REG_27__SCAN_IN), .B(keyinput_g117), .ZN(n10398)
         );
  NAND4_X1 U11476 ( .A1(n10401), .A2(n10400), .A3(n10399), .A4(n10398), .ZN(
        n10402) );
  NOR3_X1 U11477 ( .A1(n10404), .A2(n10403), .A3(n10402), .ZN(n10432) );
  AOI22_X1 U11478 ( .A1(n10406), .A2(keyinput_g77), .B1(keyinput_g59), .B2(
        n10583), .ZN(n10405) );
  OAI221_X1 U11479 ( .B1(n10406), .B2(keyinput_g77), .C1(n10583), .C2(
        keyinput_g59), .A(n10405), .ZN(n10418) );
  INV_X1 U11480 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n10408) );
  AOI22_X1 U11481 ( .A1(n10408), .A2(keyinput_g106), .B1(keyinput_g124), .B2(
        n10597), .ZN(n10407) );
  OAI221_X1 U11482 ( .B1(n10408), .B2(keyinput_g106), .C1(n10597), .C2(
        keyinput_g124), .A(n10407), .ZN(n10417) );
  AOI22_X1 U11483 ( .A1(n10411), .A2(keyinput_g58), .B1(n10410), .B2(
        keyinput_g84), .ZN(n10409) );
  OAI221_X1 U11484 ( .B1(n10411), .B2(keyinput_g58), .C1(n10410), .C2(
        keyinput_g84), .A(n10409), .ZN(n10416) );
  XOR2_X1 U11485 ( .A(n10412), .B(keyinput_g83), .Z(n10414) );
  XNOR2_X1 U11486 ( .A(P1_IR_REG_25__SCAN_IN), .B(keyinput_g115), .ZN(n10413)
         );
  NAND2_X1 U11487 ( .A1(n10414), .A2(n10413), .ZN(n10415) );
  NOR4_X1 U11488 ( .A1(n10418), .A2(n10417), .A3(n10416), .A4(n10415), .ZN(
        n10431) );
  AOI22_X1 U11489 ( .A1(n5200), .A2(keyinput_g33), .B1(n10420), .B2(
        keyinput_g123), .ZN(n10419) );
  OAI221_X1 U11490 ( .B1(n5200), .B2(keyinput_g33), .C1(n10420), .C2(
        keyinput_g123), .A(n10419), .ZN(n10429) );
  INV_X1 U11491 ( .A(SI_10_), .ZN(n10422) );
  AOI22_X1 U11492 ( .A1(n10422), .A2(keyinput_g22), .B1(keyinput_g50), .B2(
        n10556), .ZN(n10421) );
  OAI221_X1 U11493 ( .B1(n10422), .B2(keyinput_g22), .C1(n10556), .C2(
        keyinput_g50), .A(n10421), .ZN(n10428) );
  INV_X1 U11494 ( .A(SI_7_), .ZN(n10599) );
  AOI22_X1 U11495 ( .A1(n10599), .A2(keyinput_g25), .B1(keyinput_g41), .B2(
        n10602), .ZN(n10423) );
  OAI221_X1 U11496 ( .B1(n10599), .B2(keyinput_g25), .C1(n10602), .C2(
        keyinput_g41), .A(n10423), .ZN(n10427) );
  XNOR2_X1 U11497 ( .A(P1_IR_REG_29__SCAN_IN), .B(keyinput_g119), .ZN(n10425)
         );
  XNOR2_X1 U11498 ( .A(P2_REG3_REG_0__SCAN_IN), .B(keyinput_g54), .ZN(n10424)
         );
  NAND2_X1 U11499 ( .A1(n10425), .A2(n10424), .ZN(n10426) );
  NOR4_X1 U11500 ( .A1(n10429), .A2(n10428), .A3(n10427), .A4(n10426), .ZN(
        n10430) );
  NAND4_X1 U11501 ( .A1(n10433), .A2(n10432), .A3(n10431), .A4(n10430), .ZN(
        n10434) );
  NOR4_X1 U11502 ( .A1(n10437), .A2(n10436), .A3(n10435), .A4(n10434), .ZN(
        n10637) );
  AOI22_X1 U11503 ( .A1(P2_REG3_REG_0__SCAN_IN), .A2(keyinput_f54), .B1(
        P2_REG3_REG_21__SCAN_IN), .B2(keyinput_f45), .ZN(n10438) );
  OAI221_X1 U11504 ( .B1(P2_REG3_REG_0__SCAN_IN), .B2(keyinput_f54), .C1(
        P2_REG3_REG_21__SCAN_IN), .C2(keyinput_f45), .A(n10438), .ZN(n10445)
         );
  AOI22_X1 U11505 ( .A1(SI_19_), .A2(keyinput_f13), .B1(P1_IR_REG_14__SCAN_IN), 
        .B2(keyinput_f104), .ZN(n10439) );
  OAI221_X1 U11506 ( .B1(SI_19_), .B2(keyinput_f13), .C1(P1_IR_REG_14__SCAN_IN), .C2(keyinput_f104), .A(n10439), .ZN(n10444) );
  AOI22_X1 U11507 ( .A1(P2_DATAO_REG_18__SCAN_IN), .A2(keyinput_f78), .B1(
        P2_DATAO_REG_20__SCAN_IN), .B2(keyinput_f76), .ZN(n10440) );
  OAI221_X1 U11508 ( .B1(P2_DATAO_REG_18__SCAN_IN), .B2(keyinput_f78), .C1(
        P2_DATAO_REG_20__SCAN_IN), .C2(keyinput_f76), .A(n10440), .ZN(n10443)
         );
  XNOR2_X1 U11509 ( .A(n10441), .B(keyinput_f114), .ZN(n10442) );
  NOR4_X1 U11510 ( .A1(n10445), .A2(n10444), .A3(n10443), .A4(n10442), .ZN(
        n10473) );
  AOI22_X1 U11511 ( .A1(P2_DATAO_REG_9__SCAN_IN), .A2(keyinput_f87), .B1(
        P1_IR_REG_13__SCAN_IN), .B2(keyinput_f103), .ZN(n10446) );
  OAI221_X1 U11512 ( .B1(P2_DATAO_REG_9__SCAN_IN), .B2(keyinput_f87), .C1(
        P1_IR_REG_13__SCAN_IN), .C2(keyinput_f103), .A(n10446), .ZN(n10453) );
  AOI22_X1 U11513 ( .A1(P2_REG3_REG_24__SCAN_IN), .A2(keyinput_f51), .B1(
        P1_IR_REG_31__SCAN_IN), .B2(keyinput_f121), .ZN(n10447) );
  OAI221_X1 U11514 ( .B1(P2_REG3_REG_24__SCAN_IN), .B2(keyinput_f51), .C1(
        P1_IR_REG_31__SCAN_IN), .C2(keyinput_f121), .A(n10447), .ZN(n10452) );
  AOI22_X1 U11515 ( .A1(P2_DATAO_REG_8__SCAN_IN), .A2(keyinput_f88), .B1(
        SI_26_), .B2(keyinput_f6), .ZN(n10448) );
  OAI221_X1 U11516 ( .B1(P2_DATAO_REG_8__SCAN_IN), .B2(keyinput_f88), .C1(
        SI_26_), .C2(keyinput_f6), .A(n10448), .ZN(n10451) );
  AOI22_X1 U11517 ( .A1(P2_REG3_REG_11__SCAN_IN), .A2(keyinput_f58), .B1(SI_0_), .B2(keyinput_f32), .ZN(n10449) );
  OAI221_X1 U11518 ( .B1(P2_REG3_REG_11__SCAN_IN), .B2(keyinput_f58), .C1(
        SI_0_), .C2(keyinput_f32), .A(n10449), .ZN(n10450) );
  NOR4_X1 U11519 ( .A1(n10453), .A2(n10452), .A3(n10451), .A4(n10450), .ZN(
        n10472) );
  AOI22_X1 U11520 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(keyinput_f98), .B1(
        P1_IR_REG_12__SCAN_IN), .B2(keyinput_f102), .ZN(n10454) );
  OAI221_X1 U11521 ( .B1(P1_IR_REG_8__SCAN_IN), .B2(keyinput_f98), .C1(
        P1_IR_REG_12__SCAN_IN), .C2(keyinput_f102), .A(n10454), .ZN(n10461) );
  AOI22_X1 U11522 ( .A1(SI_10_), .A2(keyinput_f22), .B1(P1_IR_REG_11__SCAN_IN), 
        .B2(keyinput_f101), .ZN(n10455) );
  OAI221_X1 U11523 ( .B1(SI_10_), .B2(keyinput_f22), .C1(P1_IR_REG_11__SCAN_IN), .C2(keyinput_f101), .A(n10455), .ZN(n10460) );
  AOI22_X1 U11524 ( .A1(SI_3_), .A2(keyinput_f29), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(keyinput_f83), .ZN(n10456) );
  OAI221_X1 U11525 ( .B1(SI_3_), .B2(keyinput_f29), .C1(
        P2_DATAO_REG_13__SCAN_IN), .C2(keyinput_f83), .A(n10456), .ZN(n10459)
         );
  AOI22_X1 U11526 ( .A1(SI_28_), .A2(keyinput_f4), .B1(
        P2_DATAO_REG_22__SCAN_IN), .B2(keyinput_f74), .ZN(n10457) );
  OAI221_X1 U11527 ( .B1(SI_28_), .B2(keyinput_f4), .C1(
        P2_DATAO_REG_22__SCAN_IN), .C2(keyinput_f74), .A(n10457), .ZN(n10458)
         );
  NOR4_X1 U11528 ( .A1(n10461), .A2(n10460), .A3(n10459), .A4(n10458), .ZN(
        n10471) );
  AOI22_X1 U11529 ( .A1(P2_REG3_REG_28__SCAN_IN), .A2(keyinput_f42), .B1(
        P1_IR_REG_19__SCAN_IN), .B2(keyinput_f109), .ZN(n10462) );
  OAI221_X1 U11530 ( .B1(P2_REG3_REG_28__SCAN_IN), .B2(keyinput_f42), .C1(
        P1_IR_REG_19__SCAN_IN), .C2(keyinput_f109), .A(n10462), .ZN(n10469) );
  AOI22_X1 U11531 ( .A1(P2_DATAO_REG_17__SCAN_IN), .A2(keyinput_f79), .B1(
        P1_IR_REG_17__SCAN_IN), .B2(keyinput_f107), .ZN(n10463) );
  OAI221_X1 U11532 ( .B1(P2_DATAO_REG_17__SCAN_IN), .B2(keyinput_f79), .C1(
        P1_IR_REG_17__SCAN_IN), .C2(keyinput_f107), .A(n10463), .ZN(n10468) );
  AOI22_X1 U11533 ( .A1(P2_REG3_REG_7__SCAN_IN), .A2(keyinput_f35), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(keyinput_f80), .ZN(n10464) );
  OAI221_X1 U11534 ( .B1(P2_REG3_REG_7__SCAN_IN), .B2(keyinput_f35), .C1(
        P2_DATAO_REG_16__SCAN_IN), .C2(keyinput_f80), .A(n10464), .ZN(n10467)
         );
  AOI22_X1 U11535 ( .A1(SI_13_), .A2(keyinput_f19), .B1(SI_20_), .B2(
        keyinput_f12), .ZN(n10465) );
  OAI221_X1 U11536 ( .B1(SI_13_), .B2(keyinput_f19), .C1(SI_20_), .C2(
        keyinput_f12), .A(n10465), .ZN(n10466) );
  NOR4_X1 U11537 ( .A1(n10469), .A2(n10468), .A3(n10467), .A4(n10466), .ZN(
        n10470) );
  NAND4_X1 U11538 ( .A1(n10473), .A2(n10472), .A3(n10471), .A4(n10470), .ZN(
        n10631) );
  AOI22_X1 U11539 ( .A1(P2_DATAO_REG_31__SCAN_IN), .A2(keyinput_f65), .B1(
        P2_REG3_REG_26__SCAN_IN), .B2(keyinput_f62), .ZN(n10474) );
  OAI221_X1 U11540 ( .B1(P2_DATAO_REG_31__SCAN_IN), .B2(keyinput_f65), .C1(
        P2_REG3_REG_26__SCAN_IN), .C2(keyinput_f62), .A(n10474), .ZN(n10481)
         );
  AOI22_X1 U11541 ( .A1(P2_REG3_REG_25__SCAN_IN), .A2(keyinput_f47), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(keyinput_f86), .ZN(n10475) );
  OAI221_X1 U11542 ( .B1(P2_REG3_REG_25__SCAN_IN), .B2(keyinput_f47), .C1(
        P2_DATAO_REG_10__SCAN_IN), .C2(keyinput_f86), .A(n10475), .ZN(n10480)
         );
  AOI22_X1 U11543 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(keyinput_f53), .B1(
        P1_IR_REG_30__SCAN_IN), .B2(keyinput_f120), .ZN(n10476) );
  OAI221_X1 U11544 ( .B1(P2_REG3_REG_9__SCAN_IN), .B2(keyinput_f53), .C1(
        P1_IR_REG_30__SCAN_IN), .C2(keyinput_f120), .A(n10476), .ZN(n10479) );
  AOI22_X1 U11545 ( .A1(P1_IR_REG_28__SCAN_IN), .A2(keyinput_f118), .B1(
        P1_IR_REG_16__SCAN_IN), .B2(keyinput_f106), .ZN(n10477) );
  OAI221_X1 U11546 ( .B1(P1_IR_REG_28__SCAN_IN), .B2(keyinput_f118), .C1(
        P1_IR_REG_16__SCAN_IN), .C2(keyinput_f106), .A(n10477), .ZN(n10478) );
  NOR4_X1 U11547 ( .A1(n10481), .A2(n10480), .A3(n10479), .A4(n10478), .ZN(
        n10509) );
  AOI22_X1 U11548 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(keyinput_f93), .B1(
        P1_IR_REG_5__SCAN_IN), .B2(keyinput_f95), .ZN(n10482) );
  OAI221_X1 U11549 ( .B1(P1_IR_REG_3__SCAN_IN), .B2(keyinput_f93), .C1(
        P1_IR_REG_5__SCAN_IN), .C2(keyinput_f95), .A(n10482), .ZN(n10489) );
  AOI22_X1 U11550 ( .A1(P1_D_REG_1__SCAN_IN), .A2(keyinput_f123), .B1(
        P1_IR_REG_10__SCAN_IN), .B2(keyinput_f100), .ZN(n10483) );
  OAI221_X1 U11551 ( .B1(P1_D_REG_1__SCAN_IN), .B2(keyinput_f123), .C1(
        P1_IR_REG_10__SCAN_IN), .C2(keyinput_f100), .A(n10483), .ZN(n10488) );
  AOI22_X1 U11552 ( .A1(SI_6_), .A2(keyinput_f26), .B1(
        P2_DATAO_REG_21__SCAN_IN), .B2(keyinput_f75), .ZN(n10484) );
  OAI221_X1 U11553 ( .B1(SI_6_), .B2(keyinput_f26), .C1(
        P2_DATAO_REG_21__SCAN_IN), .C2(keyinput_f75), .A(n10484), .ZN(n10487)
         );
  AOI22_X1 U11554 ( .A1(P2_DATAO_REG_12__SCAN_IN), .A2(keyinput_f84), .B1(
        P1_IR_REG_2__SCAN_IN), .B2(keyinput_f92), .ZN(n10485) );
  OAI221_X1 U11555 ( .B1(P2_DATAO_REG_12__SCAN_IN), .B2(keyinput_f84), .C1(
        P1_IR_REG_2__SCAN_IN), .C2(keyinput_f92), .A(n10485), .ZN(n10486) );
  NOR4_X1 U11556 ( .A1(n10489), .A2(n10488), .A3(n10487), .A4(n10486), .ZN(
        n10508) );
  AOI22_X1 U11557 ( .A1(P2_REG3_REG_15__SCAN_IN), .A2(keyinput_f63), .B1(
        P2_DATAO_REG_19__SCAN_IN), .B2(keyinput_f77), .ZN(n10490) );
  OAI221_X1 U11558 ( .B1(P2_REG3_REG_15__SCAN_IN), .B2(keyinput_f63), .C1(
        P2_DATAO_REG_19__SCAN_IN), .C2(keyinput_f77), .A(n10490), .ZN(n10497)
         );
  AOI22_X1 U11559 ( .A1(P2_RD_REG_SCAN_IN), .A2(keyinput_f33), .B1(
        P1_IR_REG_21__SCAN_IN), .B2(keyinput_f111), .ZN(n10491) );
  OAI221_X1 U11560 ( .B1(P2_RD_REG_SCAN_IN), .B2(keyinput_f33), .C1(
        P1_IR_REG_21__SCAN_IN), .C2(keyinput_f111), .A(n10491), .ZN(n10496) );
  AOI22_X1 U11561 ( .A1(P2_DATAO_REG_29__SCAN_IN), .A2(keyinput_f67), .B1(
        SI_29_), .B2(keyinput_f3), .ZN(n10492) );
  OAI221_X1 U11562 ( .B1(P2_DATAO_REG_29__SCAN_IN), .B2(keyinput_f67), .C1(
        SI_29_), .C2(keyinput_f3), .A(n10492), .ZN(n10495) );
  AOI22_X1 U11563 ( .A1(P2_DATAO_REG_30__SCAN_IN), .A2(keyinput_f66), .B1(
        P2_DATAO_REG_7__SCAN_IN), .B2(keyinput_f89), .ZN(n10493) );
  OAI221_X1 U11564 ( .B1(P2_DATAO_REG_30__SCAN_IN), .B2(keyinput_f66), .C1(
        P2_DATAO_REG_7__SCAN_IN), .C2(keyinput_f89), .A(n10493), .ZN(n10494)
         );
  NOR4_X1 U11565 ( .A1(n10497), .A2(n10496), .A3(n10495), .A4(n10494), .ZN(
        n10507) );
  AOI22_X1 U11566 ( .A1(P2_DATAO_REG_14__SCAN_IN), .A2(keyinput_f82), .B1(
        P1_IR_REG_15__SCAN_IN), .B2(keyinput_f105), .ZN(n10498) );
  OAI221_X1 U11567 ( .B1(P2_DATAO_REG_14__SCAN_IN), .B2(keyinput_f82), .C1(
        P1_IR_REG_15__SCAN_IN), .C2(keyinput_f105), .A(n10498), .ZN(n10505) );
  AOI22_X1 U11568 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(keyinput_f46), .B1(
        P1_IR_REG_23__SCAN_IN), .B2(keyinput_f113), .ZN(n10499) );
  OAI221_X1 U11569 ( .B1(P2_REG3_REG_12__SCAN_IN), .B2(keyinput_f46), .C1(
        P1_IR_REG_23__SCAN_IN), .C2(keyinput_f113), .A(n10499), .ZN(n10504) );
  AOI22_X1 U11570 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(keyinput_f39), .B1(
        P2_DATAO_REG_23__SCAN_IN), .B2(keyinput_f73), .ZN(n10500) );
  OAI221_X1 U11571 ( .B1(P2_REG3_REG_10__SCAN_IN), .B2(keyinput_f39), .C1(
        P2_DATAO_REG_23__SCAN_IN), .C2(keyinput_f73), .A(n10500), .ZN(n10503)
         );
  AOI22_X1 U11572 ( .A1(P2_REG3_REG_27__SCAN_IN), .A2(keyinput_f36), .B1(n5301), .B2(keyinput_f69), .ZN(n10501) );
  OAI221_X1 U11573 ( .B1(P2_REG3_REG_27__SCAN_IN), .B2(keyinput_f36), .C1(
        n5301), .C2(keyinput_f69), .A(n10501), .ZN(n10502) );
  NOR4_X1 U11574 ( .A1(n10505), .A2(n10504), .A3(n10503), .A4(n10502), .ZN(
        n10506) );
  NAND4_X1 U11575 ( .A1(n10509), .A2(n10508), .A3(n10507), .A4(n10506), .ZN(
        n10630) );
  AOI22_X1 U11576 ( .A1(n10511), .A2(keyinput_f15), .B1(keyinput_f64), .B2(
        n5790), .ZN(n10510) );
  OAI221_X1 U11577 ( .B1(n10511), .B2(keyinput_f15), .C1(n5790), .C2(
        keyinput_f64), .A(n10510), .ZN(n10522) );
  INV_X1 U11578 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n10513) );
  AOI22_X1 U11579 ( .A1(n5151), .A2(keyinput_f49), .B1(n10513), .B2(
        keyinput_f56), .ZN(n10512) );
  OAI221_X1 U11580 ( .B1(n5151), .B2(keyinput_f49), .C1(n10513), .C2(
        keyinput_f56), .A(n10512), .ZN(n10521) );
  INV_X1 U11581 ( .A(SI_12_), .ZN(n10516) );
  AOI22_X1 U11582 ( .A1(n10516), .A2(keyinput_f20), .B1(keyinput_f21), .B2(
        n10515), .ZN(n10514) );
  OAI221_X1 U11583 ( .B1(n10516), .B2(keyinput_f20), .C1(n10515), .C2(
        keyinput_f21), .A(n10514), .ZN(n10520) );
  XNOR2_X1 U11584 ( .A(P1_IR_REG_29__SCAN_IN), .B(keyinput_f119), .ZN(n10518)
         );
  XNOR2_X1 U11585 ( .A(SI_30_), .B(keyinput_f2), .ZN(n10517) );
  NAND2_X1 U11586 ( .A1(n10518), .A2(n10517), .ZN(n10519) );
  NOR4_X1 U11587 ( .A1(n10522), .A2(n10521), .A3(n10520), .A4(n10519), .ZN(
        n10569) );
  AOI22_X1 U11588 ( .A1(P2_U3151), .A2(keyinput_f34), .B1(n10524), .B2(
        keyinput_f8), .ZN(n10523) );
  OAI221_X1 U11589 ( .B1(P2_U3151), .B2(keyinput_f34), .C1(n10524), .C2(
        keyinput_f8), .A(n10523), .ZN(n10537) );
  AOI22_X1 U11590 ( .A1(n10527), .A2(keyinput_f18), .B1(n10526), .B2(
        keyinput_f71), .ZN(n10525) );
  OAI221_X1 U11591 ( .B1(n10527), .B2(keyinput_f18), .C1(n10526), .C2(
        keyinput_f71), .A(n10525), .ZN(n10536) );
  AOI22_X1 U11592 ( .A1(n10530), .A2(keyinput_f70), .B1(keyinput_f61), .B2(
        n10529), .ZN(n10528) );
  OAI221_X1 U11593 ( .B1(n10530), .B2(keyinput_f70), .C1(n10529), .C2(
        keyinput_f61), .A(n10528), .ZN(n10535) );
  AOI22_X1 U11594 ( .A1(n10533), .A2(keyinput_f43), .B1(n10532), .B2(
        keyinput_f122), .ZN(n10531) );
  OAI221_X1 U11595 ( .B1(n10533), .B2(keyinput_f43), .C1(n10532), .C2(
        keyinput_f122), .A(n10531), .ZN(n10534) );
  NOR4_X1 U11596 ( .A1(n10537), .A2(n10536), .A3(n10535), .A4(n10534), .ZN(
        n10568) );
  INV_X1 U11597 ( .A(SI_8_), .ZN(n10539) );
  AOI22_X1 U11598 ( .A1(n10539), .A2(keyinput_f24), .B1(n6068), .B2(
        keyinput_f97), .ZN(n10538) );
  OAI221_X1 U11599 ( .B1(n10539), .B2(keyinput_f24), .C1(n6068), .C2(
        keyinput_f97), .A(n10538), .ZN(n10551) );
  AOI22_X1 U11600 ( .A1(n10541), .A2(keyinput_f127), .B1(n6429), .B2(
        keyinput_f112), .ZN(n10540) );
  OAI221_X1 U11601 ( .B1(n10541), .B2(keyinput_f127), .C1(n6429), .C2(
        keyinput_f112), .A(n10540), .ZN(n10550) );
  INV_X1 U11602 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n10544) );
  INV_X1 U11603 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n10543) );
  AOI22_X1 U11604 ( .A1(n10544), .A2(keyinput_f57), .B1(keyinput_f60), .B2(
        n10543), .ZN(n10542) );
  OAI221_X1 U11605 ( .B1(n10544), .B2(keyinput_f57), .C1(n10543), .C2(
        keyinput_f60), .A(n10542), .ZN(n10549) );
  XOR2_X1 U11606 ( .A(n10545), .B(keyinput_f14), .Z(n10547) );
  XNOR2_X1 U11607 ( .A(P1_IR_REG_25__SCAN_IN), .B(keyinput_f115), .ZN(n10546)
         );
  NAND2_X1 U11608 ( .A1(n10547), .A2(n10546), .ZN(n10548) );
  NOR4_X1 U11609 ( .A1(n10551), .A2(n10550), .A3(n10549), .A4(n10548), .ZN(
        n10567) );
  AOI22_X1 U11610 ( .A1(n10554), .A2(keyinput_f16), .B1(n10553), .B2(
        keyinput_f126), .ZN(n10552) );
  OAI221_X1 U11611 ( .B1(n10554), .B2(keyinput_f16), .C1(n10553), .C2(
        keyinput_f126), .A(n10552), .ZN(n10565) );
  AOI22_X1 U11612 ( .A1(n10557), .A2(keyinput_f9), .B1(keyinput_f50), .B2(
        n10556), .ZN(n10555) );
  OAI221_X1 U11613 ( .B1(n10557), .B2(keyinput_f9), .C1(n10556), .C2(
        keyinput_f50), .A(n10555), .ZN(n10564) );
  XNOR2_X1 U11614 ( .A(P1_IR_REG_27__SCAN_IN), .B(keyinput_f117), .ZN(n10560)
         );
  XNOR2_X1 U11615 ( .A(P2_REG3_REG_4__SCAN_IN), .B(keyinput_f52), .ZN(n10559)
         );
  XNOR2_X1 U11616 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(keyinput_f85), .ZN(n10558) );
  NAND3_X1 U11617 ( .A1(n10560), .A2(n10559), .A3(n10558), .ZN(n10563) );
  INV_X1 U11618 ( .A(P2_WR_REG_SCAN_IN), .ZN(n10561) );
  XNOR2_X1 U11619 ( .A(n10561), .B(keyinput_f0), .ZN(n10562) );
  NOR4_X1 U11620 ( .A1(n10565), .A2(n10564), .A3(n10563), .A4(n10562), .ZN(
        n10566) );
  NAND4_X1 U11621 ( .A1(n10569), .A2(n10568), .A3(n10567), .A4(n10566), .ZN(
        n10629) );
  AOI22_X1 U11622 ( .A1(n10572), .A2(keyinput_f5), .B1(keyinput_f68), .B2(
        n10571), .ZN(n10570) );
  OAI221_X1 U11623 ( .B1(n10572), .B2(keyinput_f5), .C1(n10571), .C2(
        keyinput_f68), .A(n10570), .ZN(n10581) );
  AOI22_X1 U11624 ( .A1(n5061), .A2(keyinput_f17), .B1(keyinput_f27), .B2(
        n10574), .ZN(n10573) );
  OAI221_X1 U11625 ( .B1(n5061), .B2(keyinput_f17), .C1(n10574), .C2(
        keyinput_f27), .A(n10573), .ZN(n10580) );
  XOR2_X1 U11626 ( .A(n5849), .B(keyinput_f116), .Z(n10578) );
  XNOR2_X1 U11627 ( .A(SI_2_), .B(keyinput_f30), .ZN(n10577) );
  XNOR2_X1 U11628 ( .A(P1_IR_REG_20__SCAN_IN), .B(keyinput_f110), .ZN(n10576)
         );
  XNOR2_X1 U11629 ( .A(SI_4_), .B(keyinput_f28), .ZN(n10575) );
  NAND4_X1 U11630 ( .A1(n10578), .A2(n10577), .A3(n10576), .A4(n10575), .ZN(
        n10579) );
  NOR3_X1 U11631 ( .A1(n10581), .A2(n10580), .A3(n10579), .ZN(n10627) );
  AOI22_X1 U11632 ( .A1(n10584), .A2(keyinput_f7), .B1(keyinput_f59), .B2(
        n10583), .ZN(n10582) );
  OAI221_X1 U11633 ( .B1(n10584), .B2(keyinput_f7), .C1(n10583), .C2(
        keyinput_f59), .A(n10582), .ZN(n10594) );
  AOI22_X1 U11634 ( .A1(n10586), .A2(keyinput_f81), .B1(n6067), .B2(
        keyinput_f96), .ZN(n10585) );
  OAI221_X1 U11635 ( .B1(n10586), .B2(keyinput_f81), .C1(n6067), .C2(
        keyinput_f96), .A(n10585), .ZN(n10593) );
  AOI22_X1 U11636 ( .A1(n5203), .A2(keyinput_f31), .B1(n10588), .B2(
        keyinput_f72), .ZN(n10587) );
  OAI221_X1 U11637 ( .B1(n5203), .B2(keyinput_f31), .C1(n10588), .C2(
        keyinput_f72), .A(n10587), .ZN(n10592) );
  XNOR2_X1 U11638 ( .A(P1_IR_REG_4__SCAN_IN), .B(keyinput_f94), .ZN(n10590) );
  XNOR2_X1 U11639 ( .A(P1_IR_REG_0__SCAN_IN), .B(keyinput_f90), .ZN(n10589) );
  NAND2_X1 U11640 ( .A1(n10590), .A2(n10589), .ZN(n10591) );
  NOR4_X1 U11641 ( .A1(n10594), .A2(n10593), .A3(n10592), .A4(n10591), .ZN(
        n10626) );
  AOI22_X1 U11642 ( .A1(n10597), .A2(keyinput_f124), .B1(keyinput_f1), .B2(
        n10596), .ZN(n10595) );
  OAI221_X1 U11643 ( .B1(n10597), .B2(keyinput_f124), .C1(n10596), .C2(
        keyinput_f1), .A(n10595), .ZN(n10609) );
  AOI22_X1 U11644 ( .A1(n10600), .A2(keyinput_f10), .B1(keyinput_f25), .B2(
        n10599), .ZN(n10598) );
  OAI221_X1 U11645 ( .B1(n10600), .B2(keyinput_f10), .C1(n10599), .C2(
        keyinput_f25), .A(n10598), .ZN(n10608) );
  INV_X1 U11646 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n10603) );
  AOI22_X1 U11647 ( .A1(n10603), .A2(keyinput_f37), .B1(n10602), .B2(
        keyinput_f41), .ZN(n10601) );
  OAI221_X1 U11648 ( .B1(n10603), .B2(keyinput_f37), .C1(n10602), .C2(
        keyinput_f41), .A(n10601), .ZN(n10607) );
  XNOR2_X1 U11649 ( .A(P1_IR_REG_18__SCAN_IN), .B(keyinput_f108), .ZN(n10605)
         );
  XNOR2_X1 U11650 ( .A(P1_IR_REG_9__SCAN_IN), .B(keyinput_f99), .ZN(n10604) );
  NAND2_X1 U11651 ( .A1(n10605), .A2(n10604), .ZN(n10606) );
  NOR4_X1 U11652 ( .A1(n10609), .A2(n10608), .A3(n10607), .A4(n10606), .ZN(
        n10625) );
  AOI22_X1 U11653 ( .A1(n10611), .A2(keyinput_f38), .B1(n4731), .B2(
        keyinput_f91), .ZN(n10610) );
  OAI221_X1 U11654 ( .B1(n10611), .B2(keyinput_f38), .C1(n4731), .C2(
        keyinput_f91), .A(n10610), .ZN(n10623) );
  AOI22_X1 U11655 ( .A1(n10614), .A2(keyinput_f23), .B1(keyinput_f55), .B2(
        n10613), .ZN(n10612) );
  OAI221_X1 U11656 ( .B1(n10614), .B2(keyinput_f23), .C1(n10613), .C2(
        keyinput_f55), .A(n10612), .ZN(n10622) );
  INV_X1 U11657 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n10617) );
  INV_X1 U11658 ( .A(SI_21_), .ZN(n10616) );
  AOI22_X1 U11659 ( .A1(n10617), .A2(keyinput_f48), .B1(n10616), .B2(
        keyinput_f11), .ZN(n10615) );
  OAI221_X1 U11660 ( .B1(n10617), .B2(keyinput_f48), .C1(n10616), .C2(
        keyinput_f11), .A(n10615), .ZN(n10621) );
  XNOR2_X1 U11661 ( .A(P2_REG3_REG_3__SCAN_IN), .B(keyinput_f40), .ZN(n10619)
         );
  XNOR2_X1 U11662 ( .A(keyinput_f44), .B(P2_REG3_REG_1__SCAN_IN), .ZN(n10618)
         );
  NAND2_X1 U11663 ( .A1(n10619), .A2(n10618), .ZN(n10620) );
  NOR4_X1 U11664 ( .A1(n10623), .A2(n10622), .A3(n10621), .A4(n10620), .ZN(
        n10624) );
  NAND4_X1 U11665 ( .A1(n10627), .A2(n10626), .A3(n10625), .A4(n10624), .ZN(
        n10628) );
  OR4_X1 U11666 ( .A1(n10631), .A2(n10630), .A3(n10629), .A4(n10628), .ZN(
        n10633) );
  AOI21_X1 U11667 ( .B1(keyinput_f125), .B2(n10633), .A(keyinput_g125), .ZN(
        n10635) );
  INV_X1 U11668 ( .A(keyinput_f125), .ZN(n10632) );
  AOI21_X1 U11669 ( .B1(n10633), .B2(n10632), .A(P1_D_REG_3__SCAN_IN), .ZN(
        n10634) );
  AOI22_X1 U11670 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n10635), .B1(keyinput_g125), 
        .B2(n10634), .ZN(n10636) );
  AOI21_X1 U11671 ( .B1(n10638), .B2(n10637), .A(n10636), .ZN(n10640) );
  XNOR2_X1 U11672 ( .A(P1_ADDR_REG_19__SCAN_IN), .B(P2_ADDR_REG_19__SCAN_IN), 
        .ZN(n10639) );
  XNOR2_X1 U11673 ( .A(n10640), .B(n10639), .ZN(n10641) );
  XNOR2_X1 U11674 ( .A(n10642), .B(n10641), .ZN(ADD_1068_U4) );
  OAI21_X1 U11675 ( .B1(n10645), .B2(n10644), .A(n10643), .ZN(ADD_1068_U47) );
  AOI21_X1 U11676 ( .B1(n10648), .B2(n10647), .A(n10646), .ZN(ADD_1068_U54) );
  OAI21_X1 U11677 ( .B1(n10651), .B2(n10650), .A(n10649), .ZN(ADD_1068_U51) );
  OAI21_X1 U11678 ( .B1(n10654), .B2(n10653), .A(n10652), .ZN(ADD_1068_U49) );
  OAI21_X1 U11679 ( .B1(n10657), .B2(n10656), .A(n10655), .ZN(ADD_1068_U48) );
  OAI21_X1 U11680 ( .B1(n10660), .B2(n10659), .A(n10658), .ZN(ADD_1068_U50) );
  AOI21_X1 U11681 ( .B1(n10663), .B2(n10662), .A(n10661), .ZN(ADD_1068_U53) );
  OAI21_X1 U11682 ( .B1(n10666), .B2(n10665), .A(n10664), .ZN(ADD_1068_U52) );
  OR2_X1 U5057 ( .A1(n8899), .A2(n4884), .ZN(n4883) );
  NOR2_X1 U5245 ( .A1(n8899), .A2(n4890), .ZN(n4597) );
  CLKBUF_X1 U5259 ( .A(n5348), .Z(n5775) );
  CLKBUF_X1 U5761 ( .A(n5382), .Z(n5581) );
  CLKBUF_X1 U6335 ( .A(n5341), .Z(n5781) );
  CLKBUF_X2 U6462 ( .A(n5890), .Z(n4513) );
endmodule

