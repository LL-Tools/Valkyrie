

module b17_C_AntiSAT_k_128_1 ( P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, 
        DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, 
        DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, 
        DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, 
        DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, 
        DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, 
        HOLD, NA, BS16, READY1, READY2, P1_READREQUEST_REG_SCAN_IN, 
        P1_ADS_N_REG_SCAN_IN, P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, 
        P1_D_C_N_REG_SCAN_IN, P1_REQUESTPENDING_REG_SCAN_IN, 
        P1_STATEBS16_REG_SCAN_IN, P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, 
        P1_W_R_N_REG_SCAN_IN, P1_BYTEENABLE_REG_0__SCAN_IN, 
        P1_BYTEENABLE_REG_1__SCAN_IN, P1_BYTEENABLE_REG_2__SCAN_IN, 
        P1_BYTEENABLE_REG_3__SCAN_IN, P1_REIP_REG_31__SCAN_IN, 
        P1_REIP_REG_30__SCAN_IN, P1_REIP_REG_29__SCAN_IN, 
        P1_REIP_REG_28__SCAN_IN, P1_REIP_REG_27__SCAN_IN, 
        P1_REIP_REG_26__SCAN_IN, P1_REIP_REG_25__SCAN_IN, 
        P1_REIP_REG_24__SCAN_IN, P1_REIP_REG_23__SCAN_IN, 
        P1_REIP_REG_22__SCAN_IN, P1_REIP_REG_21__SCAN_IN, 
        P1_REIP_REG_20__SCAN_IN, P1_REIP_REG_19__SCAN_IN, 
        P1_REIP_REG_18__SCAN_IN, P1_REIP_REG_17__SCAN_IN, 
        P1_REIP_REG_16__SCAN_IN, P1_REIP_REG_15__SCAN_IN, 
        P1_REIP_REG_14__SCAN_IN, P1_REIP_REG_13__SCAN_IN, 
        P1_REIP_REG_12__SCAN_IN, P1_REIP_REG_11__SCAN_IN, 
        P1_REIP_REG_10__SCAN_IN, P1_REIP_REG_9__SCAN_IN, 
        P1_REIP_REG_8__SCAN_IN, P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN, 
        P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN, P1_REIP_REG_3__SCAN_IN, 
        P1_REIP_REG_2__SCAN_IN, P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN, 
        P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN, P1_EBX_REG_29__SCAN_IN, 
        P1_EBX_REG_28__SCAN_IN, P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN, 
        P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN, P1_EBX_REG_23__SCAN_IN, 
        P1_EBX_REG_22__SCAN_IN, P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN, 
        P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN, P1_EBX_REG_17__SCAN_IN, 
        P1_EBX_REG_16__SCAN_IN, P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN, 
        P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN, P1_EBX_REG_11__SCAN_IN, 
        P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN, P1_EBX_REG_8__SCAN_IN, 
        P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN, P1_EBX_REG_5__SCAN_IN, 
        P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN, P1_EBX_REG_2__SCAN_IN, 
        P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN, P1_EAX_REG_31__SCAN_IN, 
        P1_EAX_REG_30__SCAN_IN, P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN, 
        P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN, P1_EAX_REG_25__SCAN_IN, 
        P1_EAX_REG_24__SCAN_IN, P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN, 
        P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN, P1_EAX_REG_19__SCAN_IN, 
        P1_EAX_REG_18__SCAN_IN, P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN, 
        P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN, P1_EAX_REG_13__SCAN_IN, 
        P1_EAX_REG_12__SCAN_IN, P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, 
        P1_EAX_REG_9__SCAN_IN, P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, 
        P1_EAX_REG_6__SCAN_IN, P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, 
        P1_EAX_REG_3__SCAN_IN, P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, 
        P1_EAX_REG_0__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_UWORD_REG_0__SCAN_IN, 
        P1_UWORD_REG_1__SCAN_IN, P1_UWORD_REG_2__SCAN_IN, 
        P1_UWORD_REG_3__SCAN_IN, P1_UWORD_REG_4__SCAN_IN, 
        P1_UWORD_REG_5__SCAN_IN, P1_UWORD_REG_6__SCAN_IN, 
        P1_UWORD_REG_7__SCAN_IN, P1_UWORD_REG_8__SCAN_IN, 
        P1_UWORD_REG_9__SCAN_IN, P1_UWORD_REG_10__SCAN_IN, 
        P1_UWORD_REG_11__SCAN_IN, P1_UWORD_REG_12__SCAN_IN, 
        P1_UWORD_REG_13__SCAN_IN, P1_UWORD_REG_14__SCAN_IN, 
        P1_LWORD_REG_0__SCAN_IN, P1_LWORD_REG_1__SCAN_IN, 
        P1_LWORD_REG_2__SCAN_IN, P1_LWORD_REG_3__SCAN_IN, 
        P1_LWORD_REG_4__SCAN_IN, P1_LWORD_REG_5__SCAN_IN, 
        P1_LWORD_REG_6__SCAN_IN, P1_LWORD_REG_7__SCAN_IN, 
        P1_LWORD_REG_8__SCAN_IN, P1_LWORD_REG_9__SCAN_IN, 
        P1_LWORD_REG_10__SCAN_IN, P1_LWORD_REG_11__SCAN_IN, 
        P1_LWORD_REG_12__SCAN_IN, P1_LWORD_REG_13__SCAN_IN, 
        P1_LWORD_REG_14__SCAN_IN, P1_LWORD_REG_15__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_31__SCAN_IN, P1_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_29__SCAN_IN, P1_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_27__SCAN_IN, P1_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_25__SCAN_IN, P1_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_23__SCAN_IN, P1_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_21__SCAN_IN, P1_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_19__SCAN_IN, P1_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_17__SCAN_IN, P1_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_13__SCAN_IN, P1_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_11__SCAN_IN, P1_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_9__SCAN_IN, P1_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_7__SCAN_IN, P1_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_5__SCAN_IN, P1_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_3__SCAN_IN, P1_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_1__SCAN_IN, P1_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_31__SCAN_IN, P1_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_29__SCAN_IN, P1_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_27__SCAN_IN, P1_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_25__SCAN_IN, P1_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_23__SCAN_IN, P1_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_21__SCAN_IN, P1_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_19__SCAN_IN, P1_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_17__SCAN_IN, P1_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_15__SCAN_IN, P1_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_13__SCAN_IN, P1_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_11__SCAN_IN, P1_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_9__SCAN_IN, P1_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_7__SCAN_IN, P1_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_5__SCAN_IN, P1_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_3__SCAN_IN, P1_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_1__SCAN_IN, P1_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P1_INSTQUEUE_REG_0__0__SCAN_IN, P1_INSTQUEUE_REG_0__1__SCAN_IN, 
        P1_INSTQUEUE_REG_0__2__SCAN_IN, P1_INSTQUEUE_REG_0__3__SCAN_IN, 
        P1_INSTQUEUE_REG_0__4__SCAN_IN, P1_INSTQUEUE_REG_0__5__SCAN_IN, 
        P1_INSTQUEUE_REG_0__6__SCAN_IN, P1_INSTQUEUE_REG_0__7__SCAN_IN, 
        P1_INSTQUEUE_REG_1__0__SCAN_IN, P1_INSTQUEUE_REG_1__1__SCAN_IN, 
        P1_INSTQUEUE_REG_1__2__SCAN_IN, P1_INSTQUEUE_REG_1__3__SCAN_IN, 
        P1_INSTQUEUE_REG_1__4__SCAN_IN, P1_INSTQUEUE_REG_1__5__SCAN_IN, 
        P1_INSTQUEUE_REG_1__6__SCAN_IN, P1_INSTQUEUE_REG_1__7__SCAN_IN, 
        P1_INSTQUEUE_REG_2__0__SCAN_IN, P1_INSTQUEUE_REG_2__1__SCAN_IN, 
        P1_INSTQUEUE_REG_2__2__SCAN_IN, P1_INSTQUEUE_REG_2__3__SCAN_IN, 
        P1_INSTQUEUE_REG_2__4__SCAN_IN, P1_INSTQUEUE_REG_2__5__SCAN_IN, 
        P1_INSTQUEUE_REG_2__6__SCAN_IN, P1_INSTQUEUE_REG_2__7__SCAN_IN, 
        P1_INSTQUEUE_REG_3__0__SCAN_IN, P1_INSTQUEUE_REG_3__1__SCAN_IN, 
        P1_INSTQUEUE_REG_3__2__SCAN_IN, P1_INSTQUEUE_REG_3__3__SCAN_IN, 
        P1_INSTQUEUE_REG_3__4__SCAN_IN, P1_INSTQUEUE_REG_3__5__SCAN_IN, 
        P1_INSTQUEUE_REG_3__6__SCAN_IN, P1_INSTQUEUE_REG_3__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__0__SCAN_IN, BUF1_REG_0__SCAN_IN, 
        BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN, BUF1_REG_3__SCAN_IN, 
        BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN, BUF1_REG_6__SCAN_IN, 
        BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN, BUF1_REG_9__SCAN_IN, 
        BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN, BUF1_REG_12__SCAN_IN, 
        BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN, BUF1_REG_15__SCAN_IN, 
        BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN, BUF1_REG_18__SCAN_IN, 
        BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN, BUF1_REG_21__SCAN_IN, 
        BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN, BUF1_REG_24__SCAN_IN, 
        BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN, BUF1_REG_27__SCAN_IN, 
        BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN, BUF1_REG_30__SCAN_IN, 
        BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN, BUF2_REG_1__SCAN_IN, 
        BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN, BUF2_REG_4__SCAN_IN, 
        BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN, BUF2_REG_7__SCAN_IN, 
        BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN, BUF2_REG_10__SCAN_IN, 
        BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN, BUF2_REG_13__SCAN_IN, 
        BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN, BUF2_REG_16__SCAN_IN, 
        BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN, BUF2_REG_19__SCAN_IN, 
        BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN, BUF2_REG_22__SCAN_IN, 
        BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN, BUF2_REG_25__SCAN_IN, 
        BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN, BUF2_REG_28__SCAN_IN, 
        BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN, BUF2_REG_31__SCAN_IN, 
        READY12_REG_SCAN_IN, READY21_REG_SCAN_IN, READY22_REG_SCAN_IN, 
        READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN, P3_BE_N_REG_2__SCAN_IN, 
        P3_BE_N_REG_1__SCAN_IN, P3_BE_N_REG_0__SCAN_IN, 
        P3_ADDRESS_REG_29__SCAN_IN, P3_ADDRESS_REG_28__SCAN_IN, 
        P3_ADDRESS_REG_27__SCAN_IN, P3_ADDRESS_REG_26__SCAN_IN, 
        P3_ADDRESS_REG_25__SCAN_IN, P3_ADDRESS_REG_24__SCAN_IN, 
        P3_ADDRESS_REG_23__SCAN_IN, P3_ADDRESS_REG_22__SCAN_IN, 
        P3_ADDRESS_REG_21__SCAN_IN, P3_ADDRESS_REG_20__SCAN_IN, 
        P3_ADDRESS_REG_19__SCAN_IN, P3_ADDRESS_REG_18__SCAN_IN, 
        P3_ADDRESS_REG_17__SCAN_IN, P3_ADDRESS_REG_16__SCAN_IN, 
        P3_ADDRESS_REG_15__SCAN_IN, P3_ADDRESS_REG_14__SCAN_IN, 
        P3_ADDRESS_REG_13__SCAN_IN, P3_ADDRESS_REG_12__SCAN_IN, 
        P3_ADDRESS_REG_11__SCAN_IN, P3_ADDRESS_REG_10__SCAN_IN, 
        P3_ADDRESS_REG_9__SCAN_IN, P3_ADDRESS_REG_8__SCAN_IN, 
        P3_ADDRESS_REG_7__SCAN_IN, P3_ADDRESS_REG_6__SCAN_IN, 
        P3_ADDRESS_REG_5__SCAN_IN, P3_ADDRESS_REG_4__SCAN_IN, 
        P3_ADDRESS_REG_3__SCAN_IN, P3_ADDRESS_REG_2__SCAN_IN, 
        P3_ADDRESS_REG_1__SCAN_IN, P3_ADDRESS_REG_0__SCAN_IN, 
        P3_STATE_REG_2__SCAN_IN, P3_STATE_REG_1__SCAN_IN, 
        P3_STATE_REG_0__SCAN_IN, P3_DATAWIDTH_REG_0__SCAN_IN, 
        P3_DATAWIDTH_REG_1__SCAN_IN, P3_DATAWIDTH_REG_2__SCAN_IN, 
        P3_DATAWIDTH_REG_3__SCAN_IN, P3_DATAWIDTH_REG_4__SCAN_IN, 
        P3_DATAWIDTH_REG_5__SCAN_IN, P3_DATAWIDTH_REG_6__SCAN_IN, 
        P3_DATAWIDTH_REG_7__SCAN_IN, P3_DATAWIDTH_REG_8__SCAN_IN, 
        P3_DATAWIDTH_REG_9__SCAN_IN, P3_DATAWIDTH_REG_10__SCAN_IN, 
        P3_DATAWIDTH_REG_11__SCAN_IN, P3_DATAWIDTH_REG_12__SCAN_IN, 
        P3_DATAWIDTH_REG_13__SCAN_IN, P3_DATAWIDTH_REG_14__SCAN_IN, 
        P3_DATAWIDTH_REG_15__SCAN_IN, P3_DATAWIDTH_REG_16__SCAN_IN, 
        P3_DATAWIDTH_REG_17__SCAN_IN, P3_DATAWIDTH_REG_18__SCAN_IN, 
        P3_DATAWIDTH_REG_19__SCAN_IN, P3_DATAWIDTH_REG_20__SCAN_IN, 
        P3_DATAWIDTH_REG_21__SCAN_IN, P3_DATAWIDTH_REG_22__SCAN_IN, 
        P3_DATAWIDTH_REG_23__SCAN_IN, P3_DATAWIDTH_REG_24__SCAN_IN, 
        P3_DATAWIDTH_REG_25__SCAN_IN, P3_DATAWIDTH_REG_26__SCAN_IN, 
        P3_DATAWIDTH_REG_27__SCAN_IN, P3_DATAWIDTH_REG_28__SCAN_IN, 
        P3_DATAWIDTH_REG_29__SCAN_IN, P3_DATAWIDTH_REG_30__SCAN_IN, 
        P3_DATAWIDTH_REG_31__SCAN_IN, P3_STATE2_REG_3__SCAN_IN, 
        P3_STATE2_REG_2__SCAN_IN, P3_STATE2_REG_1__SCAN_IN, 
        P3_STATE2_REG_0__SCAN_IN, P3_INSTQUEUE_REG_15__7__SCAN_IN, 
        P3_INSTQUEUE_REG_15__6__SCAN_IN, P3_INSTQUEUE_REG_15__5__SCAN_IN, 
        P3_INSTQUEUE_REG_15__4__SCAN_IN, P3_INSTQUEUE_REG_15__3__SCAN_IN, 
        P3_INSTQUEUE_REG_15__2__SCAN_IN, P3_INSTQUEUE_REG_15__1__SCAN_IN, 
        P3_INSTQUEUE_REG_15__0__SCAN_IN, P3_INSTQUEUE_REG_14__7__SCAN_IN, 
        P3_INSTQUEUE_REG_14__6__SCAN_IN, P3_INSTQUEUE_REG_14__5__SCAN_IN, 
        P3_INSTQUEUE_REG_14__4__SCAN_IN, P3_INSTQUEUE_REG_14__3__SCAN_IN, 
        P3_INSTQUEUE_REG_14__2__SCAN_IN, P3_INSTQUEUE_REG_14__1__SCAN_IN, 
        P3_INSTQUEUE_REG_14__0__SCAN_IN, P3_INSTQUEUE_REG_13__7__SCAN_IN, 
        P3_INSTQUEUE_REG_13__6__SCAN_IN, P3_INSTQUEUE_REG_13__5__SCAN_IN, 
        P3_INSTQUEUE_REG_13__4__SCAN_IN, P3_INSTQUEUE_REG_13__3__SCAN_IN, 
        P3_INSTQUEUE_REG_13__2__SCAN_IN, P3_INSTQUEUE_REG_13__1__SCAN_IN, 
        P3_INSTQUEUE_REG_13__0__SCAN_IN, P3_INSTQUEUE_REG_12__7__SCAN_IN, 
        P3_INSTQUEUE_REG_12__6__SCAN_IN, P3_INSTQUEUE_REG_12__5__SCAN_IN, 
        P3_INSTQUEUE_REG_12__4__SCAN_IN, P3_INSTQUEUE_REG_12__3__SCAN_IN, 
        P3_INSTQUEUE_REG_12__2__SCAN_IN, P3_INSTQUEUE_REG_12__1__SCAN_IN, 
        P3_INSTQUEUE_REG_12__0__SCAN_IN, P3_INSTQUEUE_REG_11__7__SCAN_IN, 
        P3_INSTQUEUE_REG_11__6__SCAN_IN, P3_INSTQUEUE_REG_11__5__SCAN_IN, 
        P3_INSTQUEUE_REG_11__4__SCAN_IN, P3_INSTQUEUE_REG_11__3__SCAN_IN, 
        P3_INSTQUEUE_REG_11__2__SCAN_IN, P3_INSTQUEUE_REG_11__1__SCAN_IN, 
        P3_INSTQUEUE_REG_11__0__SCAN_IN, P3_INSTQUEUE_REG_10__7__SCAN_IN, 
        P3_INSTQUEUE_REG_10__6__SCAN_IN, P3_INSTQUEUE_REG_10__5__SCAN_IN, 
        P3_INSTQUEUE_REG_10__4__SCAN_IN, P3_INSTQUEUE_REG_10__3__SCAN_IN, 
        P3_INSTQUEUE_REG_10__2__SCAN_IN, P3_INSTQUEUE_REG_10__1__SCAN_IN, 
        P3_INSTQUEUE_REG_10__0__SCAN_IN, P3_INSTQUEUE_REG_9__7__SCAN_IN, 
        P3_INSTQUEUE_REG_9__6__SCAN_IN, P3_INSTQUEUE_REG_9__5__SCAN_IN, 
        P3_INSTQUEUE_REG_9__4__SCAN_IN, P3_INSTQUEUE_REG_9__3__SCAN_IN, 
        P3_INSTQUEUE_REG_9__2__SCAN_IN, P3_INSTQUEUE_REG_9__1__SCAN_IN, 
        P3_INSTQUEUE_REG_9__0__SCAN_IN, P3_INSTQUEUE_REG_8__7__SCAN_IN, 
        P3_INSTQUEUE_REG_8__6__SCAN_IN, P3_INSTQUEUE_REG_8__5__SCAN_IN, 
        P3_INSTQUEUE_REG_8__4__SCAN_IN, P3_INSTQUEUE_REG_8__3__SCAN_IN, 
        P3_INSTQUEUE_REG_8__2__SCAN_IN, P3_INSTQUEUE_REG_8__1__SCAN_IN, 
        P3_INSTQUEUE_REG_8__0__SCAN_IN, P3_INSTQUEUE_REG_7__7__SCAN_IN, 
        P3_INSTQUEUE_REG_7__6__SCAN_IN, P3_INSTQUEUE_REG_7__5__SCAN_IN, 
        P3_INSTQUEUE_REG_7__4__SCAN_IN, P3_INSTQUEUE_REG_7__3__SCAN_IN, 
        P3_INSTQUEUE_REG_7__2__SCAN_IN, P3_INSTQUEUE_REG_7__1__SCAN_IN, 
        P3_INSTQUEUE_REG_7__0__SCAN_IN, P3_INSTQUEUE_REG_6__7__SCAN_IN, 
        P3_INSTQUEUE_REG_6__6__SCAN_IN, P3_INSTQUEUE_REG_6__5__SCAN_IN, 
        P3_INSTQUEUE_REG_6__4__SCAN_IN, P3_INSTQUEUE_REG_6__3__SCAN_IN, 
        P3_INSTQUEUE_REG_6__2__SCAN_IN, P3_INSTQUEUE_REG_6__1__SCAN_IN, 
        P3_INSTQUEUE_REG_6__0__SCAN_IN, P3_INSTQUEUE_REG_5__7__SCAN_IN, 
        P3_INSTQUEUE_REG_5__6__SCAN_IN, P3_INSTQUEUE_REG_5__5__SCAN_IN, 
        P3_INSTQUEUE_REG_5__4__SCAN_IN, P3_INSTQUEUE_REG_5__3__SCAN_IN, 
        P3_INSTQUEUE_REG_5__2__SCAN_IN, P3_INSTQUEUE_REG_5__1__SCAN_IN, 
        P3_INSTQUEUE_REG_5__0__SCAN_IN, P3_INSTQUEUE_REG_4__7__SCAN_IN, 
        P3_INSTQUEUE_REG_4__6__SCAN_IN, P3_INSTQUEUE_REG_4__5__SCAN_IN, 
        P3_INSTQUEUE_REG_4__4__SCAN_IN, P3_INSTQUEUE_REG_4__3__SCAN_IN, 
        P3_INSTQUEUE_REG_4__2__SCAN_IN, P3_INSTQUEUE_REG_4__1__SCAN_IN, 
        P3_INSTQUEUE_REG_4__0__SCAN_IN, P3_INSTQUEUE_REG_3__7__SCAN_IN, 
        P3_INSTQUEUE_REG_3__6__SCAN_IN, P3_INSTQUEUE_REG_3__5__SCAN_IN, 
        P3_INSTQUEUE_REG_3__4__SCAN_IN, P3_INSTQUEUE_REG_3__3__SCAN_IN, 
        P3_INSTQUEUE_REG_3__2__SCAN_IN, P3_INSTQUEUE_REG_3__1__SCAN_IN, 
        P3_INSTQUEUE_REG_3__0__SCAN_IN, P3_INSTQUEUE_REG_2__7__SCAN_IN, 
        P3_INSTQUEUE_REG_2__6__SCAN_IN, P3_INSTQUEUE_REG_2__5__SCAN_IN, 
        P3_INSTQUEUE_REG_2__4__SCAN_IN, P3_INSTQUEUE_REG_2__3__SCAN_IN, 
        P3_INSTQUEUE_REG_2__2__SCAN_IN, P3_INSTQUEUE_REG_2__1__SCAN_IN, 
        P3_INSTQUEUE_REG_2__0__SCAN_IN, P3_INSTQUEUE_REG_1__7__SCAN_IN, 
        P3_INSTQUEUE_REG_1__6__SCAN_IN, P3_INSTQUEUE_REG_1__5__SCAN_IN, 
        P3_INSTQUEUE_REG_1__4__SCAN_IN, P3_INSTQUEUE_REG_1__3__SCAN_IN, 
        P3_INSTQUEUE_REG_1__2__SCAN_IN, P3_INSTQUEUE_REG_1__1__SCAN_IN, 
        P3_INSTQUEUE_REG_1__0__SCAN_IN, P3_INSTQUEUE_REG_0__7__SCAN_IN, 
        P3_INSTQUEUE_REG_0__6__SCAN_IN, P3_INSTQUEUE_REG_0__5__SCAN_IN, 
        P3_INSTQUEUE_REG_0__4__SCAN_IN, P3_INSTQUEUE_REG_0__3__SCAN_IN, 
        P3_INSTQUEUE_REG_0__2__SCAN_IN, P3_INSTQUEUE_REG_0__1__SCAN_IN, 
        P3_INSTQUEUE_REG_0__0__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_15__SCAN_IN, P3_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_17__SCAN_IN, P3_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_19__SCAN_IN, P3_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_21__SCAN_IN, P3_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_23__SCAN_IN, P3_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_25__SCAN_IN, P3_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_29__SCAN_IN, P3_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN, 
        P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN, 
        P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN, 
        P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN, 
        P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN, 
        P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN, 
        P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN, 
        P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN, 
        P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN, 
        P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN, 
        P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN, 
        P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN, 
        P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN, 
        P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN, 
        P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN, 
        P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN, 
        P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN, 
        P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN, 
        P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN, 
        P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN, P3_EAX_REG_14__SCAN_IN, 
        P3_EAX_REG_15__SCAN_IN, P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN, 
        P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN, P3_EAX_REG_20__SCAN_IN, 
        P3_EAX_REG_21__SCAN_IN, P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN, 
        P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN, P3_EAX_REG_26__SCAN_IN, 
        P3_EAX_REG_27__SCAN_IN, P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN, 
        P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN, 
        P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN, 
        P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN, 
        P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN, 
        P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN, P3_EBX_REG_12__SCAN_IN, 
        P3_EBX_REG_13__SCAN_IN, P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN, 
        P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN, P3_EBX_REG_18__SCAN_IN, 
        P3_EBX_REG_19__SCAN_IN, P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN, 
        P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN, P3_EBX_REG_24__SCAN_IN, 
        P3_EBX_REG_25__SCAN_IN, P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN, 
        P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN, P3_EBX_REG_30__SCAN_IN, 
        P3_EBX_REG_31__SCAN_IN, P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN, 
        P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN, P3_REIP_REG_4__SCAN_IN, 
        P3_REIP_REG_5__SCAN_IN, P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN, 
        P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN, 
        P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN, 
        P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN, 
        P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN, 
        P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN, 
        P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN, 
        P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN, 
        P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN, 
        P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN, 
        P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN, 
        P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN, 
        P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN, 
        P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN, 
        P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN, 
        P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN, 
        P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN, 
        P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN, 
        P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN, 
        P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN, 
        P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN, P2_BE_N_REG_0__SCAN_IN, 
        P2_ADDRESS_REG_29__SCAN_IN, P2_ADDRESS_REG_28__SCAN_IN, 
        P2_ADDRESS_REG_27__SCAN_IN, P2_ADDRESS_REG_26__SCAN_IN, 
        P2_ADDRESS_REG_25__SCAN_IN, P2_ADDRESS_REG_24__SCAN_IN, 
        P2_ADDRESS_REG_23__SCAN_IN, P2_ADDRESS_REG_22__SCAN_IN, 
        P2_ADDRESS_REG_21__SCAN_IN, P2_ADDRESS_REG_20__SCAN_IN, 
        P2_ADDRESS_REG_19__SCAN_IN, P2_ADDRESS_REG_18__SCAN_IN, 
        P2_ADDRESS_REG_17__SCAN_IN, P2_ADDRESS_REG_16__SCAN_IN, 
        P2_ADDRESS_REG_15__SCAN_IN, P2_ADDRESS_REG_14__SCAN_IN, 
        P2_ADDRESS_REG_13__SCAN_IN, P2_ADDRESS_REG_12__SCAN_IN, 
        P2_ADDRESS_REG_11__SCAN_IN, P2_ADDRESS_REG_10__SCAN_IN, 
        P2_ADDRESS_REG_9__SCAN_IN, P2_ADDRESS_REG_8__SCAN_IN, 
        P2_ADDRESS_REG_7__SCAN_IN, P2_ADDRESS_REG_6__SCAN_IN, 
        P2_ADDRESS_REG_5__SCAN_IN, P2_ADDRESS_REG_4__SCAN_IN, 
        P2_ADDRESS_REG_3__SCAN_IN, P2_ADDRESS_REG_2__SCAN_IN, 
        P2_ADDRESS_REG_1__SCAN_IN, P2_ADDRESS_REG_0__SCAN_IN, 
        P2_STATE_REG_2__SCAN_IN, P2_STATE_REG_1__SCAN_IN, 
        P2_STATE_REG_0__SCAN_IN, P2_DATAWIDTH_REG_0__SCAN_IN, 
        P2_DATAWIDTH_REG_1__SCAN_IN, P2_DATAWIDTH_REG_2__SCAN_IN, 
        P2_DATAWIDTH_REG_3__SCAN_IN, P2_DATAWIDTH_REG_4__SCAN_IN, 
        P2_DATAWIDTH_REG_5__SCAN_IN, P2_DATAWIDTH_REG_6__SCAN_IN, 
        P2_DATAWIDTH_REG_7__SCAN_IN, P2_DATAWIDTH_REG_8__SCAN_IN, 
        P2_DATAWIDTH_REG_9__SCAN_IN, P2_DATAWIDTH_REG_10__SCAN_IN, 
        P2_DATAWIDTH_REG_11__SCAN_IN, P2_DATAWIDTH_REG_12__SCAN_IN, 
        P2_DATAWIDTH_REG_13__SCAN_IN, P2_DATAWIDTH_REG_14__SCAN_IN, 
        P2_DATAWIDTH_REG_15__SCAN_IN, P2_DATAWIDTH_REG_16__SCAN_IN, 
        P2_DATAWIDTH_REG_17__SCAN_IN, P2_DATAWIDTH_REG_18__SCAN_IN, 
        P2_DATAWIDTH_REG_19__SCAN_IN, P2_DATAWIDTH_REG_20__SCAN_IN, 
        P2_DATAWIDTH_REG_21__SCAN_IN, P2_DATAWIDTH_REG_22__SCAN_IN, 
        P2_DATAWIDTH_REG_23__SCAN_IN, P2_DATAWIDTH_REG_24__SCAN_IN, 
        P2_DATAWIDTH_REG_25__SCAN_IN, P2_DATAWIDTH_REG_26__SCAN_IN, 
        P2_DATAWIDTH_REG_27__SCAN_IN, P2_DATAWIDTH_REG_28__SCAN_IN, 
        P2_DATAWIDTH_REG_29__SCAN_IN, P2_DATAWIDTH_REG_30__SCAN_IN, 
        P2_DATAWIDTH_REG_31__SCAN_IN, P2_STATE2_REG_3__SCAN_IN, 
        P2_STATE2_REG_2__SCAN_IN, P2_STATE2_REG_1__SCAN_IN, 
        P2_STATE2_REG_0__SCAN_IN, P2_INSTQUEUE_REG_15__7__SCAN_IN, 
        P2_INSTQUEUE_REG_15__6__SCAN_IN, P2_INSTQUEUE_REG_15__5__SCAN_IN, 
        P2_INSTQUEUE_REG_15__4__SCAN_IN, P2_INSTQUEUE_REG_15__3__SCAN_IN, 
        P2_INSTQUEUE_REG_15__2__SCAN_IN, P2_INSTQUEUE_REG_15__1__SCAN_IN, 
        P2_INSTQUEUE_REG_15__0__SCAN_IN, P2_INSTQUEUE_REG_14__7__SCAN_IN, 
        P2_INSTQUEUE_REG_14__6__SCAN_IN, P2_INSTQUEUE_REG_14__5__SCAN_IN, 
        P2_INSTQUEUE_REG_14__4__SCAN_IN, P2_INSTQUEUE_REG_14__3__SCAN_IN, 
        P2_INSTQUEUE_REG_14__2__SCAN_IN, P2_INSTQUEUE_REG_14__1__SCAN_IN, 
        P2_INSTQUEUE_REG_14__0__SCAN_IN, P2_INSTQUEUE_REG_13__7__SCAN_IN, 
        P2_INSTQUEUE_REG_13__6__SCAN_IN, P2_INSTQUEUE_REG_13__5__SCAN_IN, 
        P2_INSTQUEUE_REG_13__4__SCAN_IN, P2_INSTQUEUE_REG_13__3__SCAN_IN, 
        P2_INSTQUEUE_REG_13__2__SCAN_IN, P2_INSTQUEUE_REG_13__1__SCAN_IN, 
        P2_INSTQUEUE_REG_13__0__SCAN_IN, P2_INSTQUEUE_REG_12__7__SCAN_IN, 
        P2_INSTQUEUE_REG_12__6__SCAN_IN, P2_INSTQUEUE_REG_12__5__SCAN_IN, 
        P2_INSTQUEUE_REG_12__4__SCAN_IN, P2_INSTQUEUE_REG_12__3__SCAN_IN, 
        P2_INSTQUEUE_REG_12__2__SCAN_IN, P2_INSTQUEUE_REG_12__1__SCAN_IN, 
        P2_INSTQUEUE_REG_12__0__SCAN_IN, P2_INSTQUEUE_REG_11__7__SCAN_IN, 
        P2_INSTQUEUE_REG_11__6__SCAN_IN, P2_INSTQUEUE_REG_11__5__SCAN_IN, 
        P2_INSTQUEUE_REG_11__4__SCAN_IN, P2_INSTQUEUE_REG_11__3__SCAN_IN, 
        P2_INSTQUEUE_REG_11__2__SCAN_IN, P2_INSTQUEUE_REG_11__1__SCAN_IN, 
        P2_INSTQUEUE_REG_11__0__SCAN_IN, P2_INSTQUEUE_REG_10__7__SCAN_IN, 
        P2_INSTQUEUE_REG_10__6__SCAN_IN, P2_INSTQUEUE_REG_10__5__SCAN_IN, 
        P2_INSTQUEUE_REG_10__4__SCAN_IN, P2_INSTQUEUE_REG_10__3__SCAN_IN, 
        P2_INSTQUEUE_REG_10__2__SCAN_IN, P2_INSTQUEUE_REG_10__1__SCAN_IN, 
        P2_INSTQUEUE_REG_10__0__SCAN_IN, P2_INSTQUEUE_REG_9__7__SCAN_IN, 
        P2_INSTQUEUE_REG_9__6__SCAN_IN, P2_INSTQUEUE_REG_9__5__SCAN_IN, 
        P2_INSTQUEUE_REG_9__4__SCAN_IN, P2_INSTQUEUE_REG_9__3__SCAN_IN, 
        P2_INSTQUEUE_REG_9__2__SCAN_IN, P2_INSTQUEUE_REG_9__1__SCAN_IN, 
        P2_INSTQUEUE_REG_9__0__SCAN_IN, P2_INSTQUEUE_REG_8__7__SCAN_IN, 
        P2_INSTQUEUE_REG_8__6__SCAN_IN, P2_INSTQUEUE_REG_8__5__SCAN_IN, 
        P2_INSTQUEUE_REG_8__4__SCAN_IN, P2_INSTQUEUE_REG_8__3__SCAN_IN, 
        P2_INSTQUEUE_REG_8__2__SCAN_IN, P2_INSTQUEUE_REG_8__1__SCAN_IN, 
        P2_INSTQUEUE_REG_8__0__SCAN_IN, P2_INSTQUEUE_REG_7__7__SCAN_IN, 
        P2_INSTQUEUE_REG_7__6__SCAN_IN, P2_INSTQUEUE_REG_7__5__SCAN_IN, 
        P2_INSTQUEUE_REG_7__4__SCAN_IN, P2_INSTQUEUE_REG_7__3__SCAN_IN, 
        P2_INSTQUEUE_REG_7__2__SCAN_IN, P2_INSTQUEUE_REG_7__1__SCAN_IN, 
        P2_INSTQUEUE_REG_7__0__SCAN_IN, P2_INSTQUEUE_REG_6__7__SCAN_IN, 
        P2_INSTQUEUE_REG_6__6__SCAN_IN, P2_INSTQUEUE_REG_6__5__SCAN_IN, 
        P2_INSTQUEUE_REG_6__4__SCAN_IN, P2_INSTQUEUE_REG_6__3__SCAN_IN, 
        P2_INSTQUEUE_REG_6__2__SCAN_IN, P2_INSTQUEUE_REG_6__1__SCAN_IN, 
        P2_INSTQUEUE_REG_6__0__SCAN_IN, P2_INSTQUEUE_REG_5__7__SCAN_IN, 
        P2_INSTQUEUE_REG_5__6__SCAN_IN, P2_INSTQUEUE_REG_5__5__SCAN_IN, 
        P2_INSTQUEUE_REG_5__4__SCAN_IN, P2_INSTQUEUE_REG_5__3__SCAN_IN, 
        P2_INSTQUEUE_REG_5__2__SCAN_IN, P2_INSTQUEUE_REG_5__1__SCAN_IN, 
        P2_INSTQUEUE_REG_5__0__SCAN_IN, P2_INSTQUEUE_REG_4__7__SCAN_IN, 
        P2_INSTQUEUE_REG_4__6__SCAN_IN, P2_INSTQUEUE_REG_4__5__SCAN_IN, 
        P2_INSTQUEUE_REG_4__4__SCAN_IN, P2_INSTQUEUE_REG_4__3__SCAN_IN, 
        P2_INSTQUEUE_REG_4__2__SCAN_IN, P2_INSTQUEUE_REG_4__1__SCAN_IN, 
        P2_INSTQUEUE_REG_4__0__SCAN_IN, P2_INSTQUEUE_REG_3__7__SCAN_IN, 
        P2_INSTQUEUE_REG_3__6__SCAN_IN, P2_INSTQUEUE_REG_3__5__SCAN_IN, 
        P2_INSTQUEUE_REG_3__4__SCAN_IN, P2_INSTQUEUE_REG_3__3__SCAN_IN, 
        P2_INSTQUEUE_REG_3__2__SCAN_IN, P2_INSTQUEUE_REG_3__1__SCAN_IN, 
        P2_INSTQUEUE_REG_3__0__SCAN_IN, P2_INSTQUEUE_REG_2__7__SCAN_IN, 
        P2_INSTQUEUE_REG_2__6__SCAN_IN, P2_INSTQUEUE_REG_2__5__SCAN_IN, 
        P2_INSTQUEUE_REG_2__4__SCAN_IN, P2_INSTQUEUE_REG_2__3__SCAN_IN, 
        P2_INSTQUEUE_REG_2__2__SCAN_IN, P2_INSTQUEUE_REG_2__1__SCAN_IN, 
        P2_INSTQUEUE_REG_2__0__SCAN_IN, P2_INSTQUEUE_REG_1__7__SCAN_IN, 
        P2_INSTQUEUE_REG_1__6__SCAN_IN, P2_INSTQUEUE_REG_1__5__SCAN_IN, 
        P2_INSTQUEUE_REG_1__4__SCAN_IN, P2_INSTQUEUE_REG_1__3__SCAN_IN, 
        P2_INSTQUEUE_REG_1__2__SCAN_IN, P2_INSTQUEUE_REG_1__1__SCAN_IN, 
        P2_INSTQUEUE_REG_1__0__SCAN_IN, P2_INSTQUEUE_REG_0__7__SCAN_IN, 
        P2_INSTQUEUE_REG_0__6__SCAN_IN, P2_INSTQUEUE_REG_0__5__SCAN_IN, 
        P2_INSTQUEUE_REG_0__4__SCAN_IN, P2_INSTQUEUE_REG_0__3__SCAN_IN, 
        P2_INSTQUEUE_REG_0__2__SCAN_IN, P2_INSTQUEUE_REG_0__1__SCAN_IN, 
        P2_INSTQUEUE_REG_0__0__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_11__SCAN_IN, P2_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_13__SCAN_IN, P2_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_15__SCAN_IN, P2_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_17__SCAN_IN, P2_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_19__SCAN_IN, P2_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_21__SCAN_IN, P2_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_23__SCAN_IN, P2_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_25__SCAN_IN, P2_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_27__SCAN_IN, P2_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_29__SCAN_IN, P2_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN, 
        P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN, 
        P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN, 
        P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN, 
        P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN, 
        P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN, 
        P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN, 
        P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN, 
        P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN, 
        P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN, 
        P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN, 
        P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN, 
        P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN, 
        P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN, 
        P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN, 
        P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN, 
        P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN, 
        P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN, 
        P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN, 
        P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN, 
        P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN, 
        P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN, 
        P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN, P2_EAX_REG_14__SCAN_IN, 
        P2_EAX_REG_15__SCAN_IN, P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN, 
        P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN, P2_EAX_REG_20__SCAN_IN, 
        P2_EAX_REG_21__SCAN_IN, P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN, 
        P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN, P2_EAX_REG_26__SCAN_IN, 
        P2_EAX_REG_27__SCAN_IN, P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN, 
        P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN, 
        P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN, 
        P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN, 
        P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN, 
        P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN, P2_EBX_REG_12__SCAN_IN, 
        P2_EBX_REG_13__SCAN_IN, P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN, 
        P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN, P2_EBX_REG_18__SCAN_IN, 
        P2_EBX_REG_19__SCAN_IN, P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN, 
        P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN, P2_EBX_REG_24__SCAN_IN, 
        P2_EBX_REG_25__SCAN_IN, P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN, 
        P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN, P2_EBX_REG_30__SCAN_IN, 
        P2_EBX_REG_31__SCAN_IN, P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN, 
        P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN, P2_REIP_REG_4__SCAN_IN, 
        P2_REIP_REG_5__SCAN_IN, P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN, 
        P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN, 
        P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN, 
        P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN, 
        P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN, 
        P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN, 
        P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN, 
        P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN, 
        P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN, 
        P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN, 
        P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN, 
        P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN, 
        P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN, 
        P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN, 
        P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN, 
        P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN, 
        P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN, 
        P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN, 
        P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN, 
        P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN, 
        P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN, P1_BE_N_REG_0__SCAN_IN, 
        P1_ADDRESS_REG_29__SCAN_IN, P1_ADDRESS_REG_28__SCAN_IN, 
        P1_ADDRESS_REG_27__SCAN_IN, P1_ADDRESS_REG_26__SCAN_IN, 
        P1_ADDRESS_REG_25__SCAN_IN, P1_ADDRESS_REG_24__SCAN_IN, 
        P1_ADDRESS_REG_23__SCAN_IN, P1_ADDRESS_REG_22__SCAN_IN, 
        P1_ADDRESS_REG_21__SCAN_IN, P1_ADDRESS_REG_20__SCAN_IN, 
        P1_ADDRESS_REG_19__SCAN_IN, P1_ADDRESS_REG_18__SCAN_IN, 
        P1_ADDRESS_REG_17__SCAN_IN, P1_ADDRESS_REG_16__SCAN_IN, 
        P1_ADDRESS_REG_15__SCAN_IN, P1_ADDRESS_REG_14__SCAN_IN, 
        P1_ADDRESS_REG_13__SCAN_IN, P1_ADDRESS_REG_12__SCAN_IN, 
        P1_ADDRESS_REG_11__SCAN_IN, P1_ADDRESS_REG_10__SCAN_IN, 
        P1_ADDRESS_REG_9__SCAN_IN, P1_ADDRESS_REG_8__SCAN_IN, 
        P1_ADDRESS_REG_7__SCAN_IN, P1_ADDRESS_REG_6__SCAN_IN, 
        P1_ADDRESS_REG_5__SCAN_IN, P1_ADDRESS_REG_4__SCAN_IN, 
        P1_ADDRESS_REG_3__SCAN_IN, P1_ADDRESS_REG_2__SCAN_IN, 
        P1_ADDRESS_REG_1__SCAN_IN, P1_ADDRESS_REG_0__SCAN_IN, 
        P1_STATE_REG_2__SCAN_IN, P1_STATE_REG_1__SCAN_IN, 
        P1_STATE_REG_0__SCAN_IN, P1_DATAWIDTH_REG_0__SCAN_IN, 
        P1_DATAWIDTH_REG_1__SCAN_IN, P1_DATAWIDTH_REG_2__SCAN_IN, 
        P1_DATAWIDTH_REG_3__SCAN_IN, P1_DATAWIDTH_REG_4__SCAN_IN, 
        P1_DATAWIDTH_REG_5__SCAN_IN, P1_DATAWIDTH_REG_6__SCAN_IN, 
        P1_DATAWIDTH_REG_7__SCAN_IN, P1_DATAWIDTH_REG_8__SCAN_IN, 
        P1_DATAWIDTH_REG_9__SCAN_IN, P1_DATAWIDTH_REG_10__SCAN_IN, 
        P1_DATAWIDTH_REG_11__SCAN_IN, P1_DATAWIDTH_REG_12__SCAN_IN, 
        P1_DATAWIDTH_REG_13__SCAN_IN, P1_DATAWIDTH_REG_14__SCAN_IN, 
        P1_DATAWIDTH_REG_15__SCAN_IN, P1_DATAWIDTH_REG_16__SCAN_IN, 
        P1_DATAWIDTH_REG_17__SCAN_IN, P1_DATAWIDTH_REG_18__SCAN_IN, 
        P1_DATAWIDTH_REG_19__SCAN_IN, P1_DATAWIDTH_REG_20__SCAN_IN, 
        P1_DATAWIDTH_REG_21__SCAN_IN, P1_DATAWIDTH_REG_22__SCAN_IN, 
        P1_DATAWIDTH_REG_23__SCAN_IN, P1_DATAWIDTH_REG_24__SCAN_IN, 
        P1_DATAWIDTH_REG_25__SCAN_IN, P1_DATAWIDTH_REG_26__SCAN_IN, 
        P1_DATAWIDTH_REG_27__SCAN_IN, P1_DATAWIDTH_REG_28__SCAN_IN, 
        P1_DATAWIDTH_REG_29__SCAN_IN, P1_DATAWIDTH_REG_30__SCAN_IN, 
        P1_DATAWIDTH_REG_31__SCAN_IN, P1_STATE2_REG_3__SCAN_IN, 
        P1_STATE2_REG_2__SCAN_IN, P1_STATE2_REG_1__SCAN_IN, 
        P1_STATE2_REG_0__SCAN_IN, P1_INSTQUEUE_REG_15__7__SCAN_IN, 
        P1_INSTQUEUE_REG_15__6__SCAN_IN, P1_INSTQUEUE_REG_15__5__SCAN_IN, 
        P1_INSTQUEUE_REG_15__4__SCAN_IN, P1_INSTQUEUE_REG_15__3__SCAN_IN, 
        P1_INSTQUEUE_REG_15__2__SCAN_IN, P1_INSTQUEUE_REG_15__1__SCAN_IN, 
        P1_INSTQUEUE_REG_15__0__SCAN_IN, P1_INSTQUEUE_REG_14__7__SCAN_IN, 
        P1_INSTQUEUE_REG_14__6__SCAN_IN, P1_INSTQUEUE_REG_14__5__SCAN_IN, 
        P1_INSTQUEUE_REG_14__4__SCAN_IN, P1_INSTQUEUE_REG_14__3__SCAN_IN, 
        P1_INSTQUEUE_REG_14__2__SCAN_IN, P1_INSTQUEUE_REG_14__1__SCAN_IN, 
        P1_INSTQUEUE_REG_14__0__SCAN_IN, P1_INSTQUEUE_REG_13__7__SCAN_IN, 
        P1_INSTQUEUE_REG_13__6__SCAN_IN, P1_INSTQUEUE_REG_13__5__SCAN_IN, 
        P1_INSTQUEUE_REG_13__4__SCAN_IN, P1_INSTQUEUE_REG_13__3__SCAN_IN, 
        P1_INSTQUEUE_REG_13__2__SCAN_IN, P1_INSTQUEUE_REG_13__1__SCAN_IN, 
        P1_INSTQUEUE_REG_13__0__SCAN_IN, P1_INSTQUEUE_REG_12__7__SCAN_IN, 
        P1_INSTQUEUE_REG_12__6__SCAN_IN, P1_INSTQUEUE_REG_12__5__SCAN_IN, 
        P1_INSTQUEUE_REG_12__4__SCAN_IN, P1_INSTQUEUE_REG_12__3__SCAN_IN, 
        P1_INSTQUEUE_REG_12__2__SCAN_IN, P1_INSTQUEUE_REG_12__1__SCAN_IN, 
        P1_INSTQUEUE_REG_12__0__SCAN_IN, P1_INSTQUEUE_REG_11__7__SCAN_IN, 
        P1_INSTQUEUE_REG_11__6__SCAN_IN, P1_INSTQUEUE_REG_11__5__SCAN_IN, 
        P1_INSTQUEUE_REG_11__4__SCAN_IN, P1_INSTQUEUE_REG_11__3__SCAN_IN, 
        P1_INSTQUEUE_REG_11__2__SCAN_IN, P1_INSTQUEUE_REG_11__1__SCAN_IN, 
        P1_INSTQUEUE_REG_11__0__SCAN_IN, P1_INSTQUEUE_REG_10__7__SCAN_IN, 
        P1_INSTQUEUE_REG_10__6__SCAN_IN, P1_INSTQUEUE_REG_10__5__SCAN_IN, 
        P1_INSTQUEUE_REG_10__4__SCAN_IN, P1_INSTQUEUE_REG_10__3__SCAN_IN, 
        P1_INSTQUEUE_REG_10__2__SCAN_IN, P1_INSTQUEUE_REG_10__1__SCAN_IN, 
        P1_INSTQUEUE_REG_10__0__SCAN_IN, P1_INSTQUEUE_REG_9__7__SCAN_IN, 
        P1_INSTQUEUE_REG_9__6__SCAN_IN, P1_INSTQUEUE_REG_9__5__SCAN_IN, 
        P1_INSTQUEUE_REG_9__4__SCAN_IN, P1_INSTQUEUE_REG_9__3__SCAN_IN, 
        P1_INSTQUEUE_REG_9__2__SCAN_IN, P1_INSTQUEUE_REG_9__1__SCAN_IN, 
        P1_INSTQUEUE_REG_9__0__SCAN_IN, P1_INSTQUEUE_REG_8__7__SCAN_IN, 
        P1_INSTQUEUE_REG_8__6__SCAN_IN, P1_INSTQUEUE_REG_8__5__SCAN_IN, 
        P1_INSTQUEUE_REG_8__4__SCAN_IN, P1_INSTQUEUE_REG_8__3__SCAN_IN, 
        P1_INSTQUEUE_REG_8__2__SCAN_IN, P1_INSTQUEUE_REG_8__1__SCAN_IN, 
        P1_INSTQUEUE_REG_8__0__SCAN_IN, P1_INSTQUEUE_REG_7__7__SCAN_IN, 
        P1_INSTQUEUE_REG_7__6__SCAN_IN, P1_INSTQUEUE_REG_7__5__SCAN_IN, 
        P1_INSTQUEUE_REG_7__4__SCAN_IN, P1_INSTQUEUE_REG_7__3__SCAN_IN, 
        P1_INSTQUEUE_REG_7__2__SCAN_IN, P1_INSTQUEUE_REG_7__1__SCAN_IN, 
        P1_INSTQUEUE_REG_7__0__SCAN_IN, P1_INSTQUEUE_REG_6__7__SCAN_IN, 
        P1_INSTQUEUE_REG_6__6__SCAN_IN, P1_INSTQUEUE_REG_6__5__SCAN_IN, 
        P1_INSTQUEUE_REG_6__4__SCAN_IN, P1_INSTQUEUE_REG_6__3__SCAN_IN, 
        P1_INSTQUEUE_REG_6__2__SCAN_IN, P1_INSTQUEUE_REG_6__1__SCAN_IN, 
        P1_INSTQUEUE_REG_6__0__SCAN_IN, P1_INSTQUEUE_REG_5__7__SCAN_IN, 
        P1_INSTQUEUE_REG_5__6__SCAN_IN, P1_INSTQUEUE_REG_5__5__SCAN_IN, 
        P1_INSTQUEUE_REG_5__4__SCAN_IN, P1_INSTQUEUE_REG_5__3__SCAN_IN, 
        P1_INSTQUEUE_REG_5__2__SCAN_IN, P1_INSTQUEUE_REG_5__1__SCAN_IN, 
        P1_INSTQUEUE_REG_5__0__SCAN_IN, P1_INSTQUEUE_REG_4__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__6__SCAN_IN, P1_INSTQUEUE_REG_4__5__SCAN_IN, 
        P1_INSTQUEUE_REG_4__4__SCAN_IN, P1_INSTQUEUE_REG_4__3__SCAN_IN, 
        P1_INSTQUEUE_REG_4__2__SCAN_IN, P1_INSTQUEUE_REG_4__1__SCAN_IN, 
        keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, 
        keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, 
        keyinput12, keyinput13, keyinput14, keyinput15, keyinput16, keyinput17, 
        keyinput18, keyinput19, keyinput20, keyinput21, keyinput22, keyinput23, 
        keyinput24, keyinput25, keyinput26, keyinput27, keyinput28, keyinput29, 
        keyinput30, keyinput31, keyinput32, keyinput33, keyinput34, keyinput35, 
        keyinput36, keyinput37, keyinput38, keyinput39, keyinput40, keyinput41, 
        keyinput42, keyinput43, keyinput44, keyinput45, keyinput46, keyinput47, 
        keyinput48, keyinput49, keyinput50, keyinput51, keyinput52, keyinput53, 
        keyinput54, keyinput55, keyinput56, keyinput57, keyinput58, keyinput59, 
        keyinput60, keyinput61, keyinput62, keyinput63, keyinput64, keyinput65, 
        keyinput66, keyinput67, keyinput68, keyinput69, keyinput70, keyinput71, 
        keyinput72, keyinput73, keyinput74, keyinput75, keyinput76, keyinput77, 
        keyinput78, keyinput79, keyinput80, keyinput81, keyinput82, keyinput83, 
        keyinput84, keyinput85, keyinput86, keyinput87, keyinput88, keyinput89, 
        keyinput90, keyinput91, keyinput92, keyinput93, keyinput94, keyinput95, 
        keyinput96, keyinput97, keyinput98, keyinput99, keyinput100, 
        keyinput101, keyinput102, keyinput103, keyinput104, keyinput105, 
        keyinput106, keyinput107, keyinput108, keyinput109, keyinput110, 
        keyinput111, keyinput112, keyinput113, keyinput114, keyinput115, 
        keyinput116, keyinput117, keyinput118, keyinput119, keyinput120, 
        keyinput121, keyinput122, keyinput123, keyinput124, keyinput125, 
        keyinput126, keyinput127, U355, U356, U357, U358, U359, U360, U361, 
        U362, U363, U364, U366, U367, U368, U369, U370, U371, U372, U373, U374, 
        U375, U347, U348, U349, U350, U351, U352, U353, U354, U365, U376, U247, 
        U246, U245, U244, U243, U242, U241, U240, U239, U238, U237, U236, U235, 
        U234, U233, U232, U231, U230, U229, U228, U227, U226, U225, U224, U223, 
        U222, U221, U220, U219, U218, U217, U216, U251, U252, U253, U254, U255, 
        U256, U257, U258, U259, U260, U261, U262, U263, U264, U265, U266, U267, 
        U268, U269, U270, U271, U272, U273, U274, U275, U276, U277, U278, U279, 
        U280, U281, U282, U212, U215, U213, U214, P3_U3274, P3_U3275, P3_U3276, 
        P3_U3277, P3_U3061, P3_U3060, P3_U3059, P3_U3058, P3_U3057, P3_U3056, 
        P3_U3055, P3_U3054, P3_U3053, P3_U3052, P3_U3051, P3_U3050, P3_U3049, 
        P3_U3048, P3_U3047, P3_U3046, P3_U3045, P3_U3044, P3_U3043, P3_U3042, 
        P3_U3041, P3_U3040, P3_U3039, P3_U3038, P3_U3037, P3_U3036, P3_U3035, 
        P3_U3034, P3_U3033, P3_U3032, P3_U3031, P3_U3030, P3_U3029, P3_U3280, 
        P3_U3281, P3_U3028, P3_U3027, P3_U3026, P3_U3025, P3_U3024, P3_U3023, 
        P3_U3022, P3_U3021, P3_U3020, P3_U3019, P3_U3018, P3_U3017, P3_U3016, 
        P3_U3015, P3_U3014, P3_U3013, P3_U3012, P3_U3011, P3_U3010, P3_U3009, 
        P3_U3008, P3_U3007, P3_U3006, P3_U3005, P3_U3004, P3_U3003, P3_U3002, 
        P3_U3001, P3_U3000, P3_U2999, P3_U3282, P3_U2998, P3_U2997, P3_U2996, 
        P3_U2995, P3_U2994, P3_U2993, P3_U2992, P3_U2991, P3_U2990, P3_U2989, 
        P3_U2988, P3_U2987, P3_U2986, P3_U2985, P3_U2984, P3_U2983, P3_U2982, 
        P3_U2981, P3_U2980, P3_U2979, P3_U2978, P3_U2977, P3_U2976, P3_U2975, 
        P3_U2974, P3_U2973, P3_U2972, P3_U2971, P3_U2970, P3_U2969, P3_U2968, 
        P3_U2967, P3_U2966, P3_U2965, P3_U2964, P3_U2963, P3_U2962, P3_U2961, 
        P3_U2960, P3_U2959, P3_U2958, P3_U2957, P3_U2956, P3_U2955, P3_U2954, 
        P3_U2953, P3_U2952, P3_U2951, P3_U2950, P3_U2949, P3_U2948, P3_U2947, 
        P3_U2946, P3_U2945, P3_U2944, P3_U2943, P3_U2942, P3_U2941, P3_U2940, 
        P3_U2939, P3_U2938, P3_U2937, P3_U2936, P3_U2935, P3_U2934, P3_U2933, 
        P3_U2932, P3_U2931, P3_U2930, P3_U2929, P3_U2928, P3_U2927, P3_U2926, 
        P3_U2925, P3_U2924, P3_U2923, P3_U2922, P3_U2921, P3_U2920, P3_U2919, 
        P3_U2918, P3_U2917, P3_U2916, P3_U2915, P3_U2914, P3_U2913, P3_U2912, 
        P3_U2911, P3_U2910, P3_U2909, P3_U2908, P3_U2907, P3_U2906, P3_U2905, 
        P3_U2904, P3_U2903, P3_U2902, P3_U2901, P3_U2900, P3_U2899, P3_U2898, 
        P3_U2897, P3_U2896, P3_U2895, P3_U2894, P3_U2893, P3_U2892, P3_U2891, 
        P3_U2890, P3_U2889, P3_U2888, P3_U2887, P3_U2886, P3_U2885, P3_U2884, 
        P3_U2883, P3_U2882, P3_U2881, P3_U2880, P3_U2879, P3_U2878, P3_U2877, 
        P3_U2876, P3_U2875, P3_U2874, P3_U2873, P3_U2872, P3_U2871, P3_U2870, 
        P3_U2869, P3_U2868, P3_U3284, P3_U3285, P3_U3288, P3_U3289, P3_U3290, 
        P3_U2867, P3_U2866, P3_U2865, P3_U2864, P3_U2863, P3_U2862, P3_U2861, 
        P3_U2860, P3_U2859, P3_U2858, P3_U2857, P3_U2856, P3_U2855, P3_U2854, 
        P3_U2853, P3_U2852, P3_U2851, P3_U2850, P3_U2849, P3_U2848, P3_U2847, 
        P3_U2846, P3_U2845, P3_U2844, P3_U2843, P3_U2842, P3_U2841, P3_U2840, 
        P3_U2839, P3_U2838, P3_U2837, P3_U2836, P3_U2835, P3_U2834, P3_U2833, 
        P3_U2832, P3_U2831, P3_U2830, P3_U2829, P3_U2828, P3_U2827, P3_U2826, 
        P3_U2825, P3_U2824, P3_U2823, P3_U2822, P3_U2821, P3_U2820, P3_U2819, 
        P3_U2818, P3_U2817, P3_U2816, P3_U2815, P3_U2814, P3_U2813, P3_U2812, 
        P3_U2811, P3_U2810, P3_U2809, P3_U2808, P3_U2807, P3_U2806, P3_U2805, 
        P3_U2804, P3_U2803, P3_U2802, P3_U2801, P3_U2800, P3_U2799, P3_U2798, 
        P3_U2797, P3_U2796, P3_U2795, P3_U2794, P3_U2793, P3_U2792, P3_U2791, 
        P3_U2790, P3_U2789, P3_U2788, P3_U2787, P3_U2786, P3_U2785, P3_U2784, 
        P3_U2783, P3_U2782, P3_U2781, P3_U2780, P3_U2779, P3_U2778, P3_U2777, 
        P3_U2776, P3_U2775, P3_U2774, P3_U2773, P3_U2772, P3_U2771, P3_U2770, 
        P3_U2769, P3_U2768, P3_U2767, P3_U2766, P3_U2765, P3_U2764, P3_U2763, 
        P3_U2762, P3_U2761, P3_U2760, P3_U2759, P3_U2758, P3_U2757, P3_U2756, 
        P3_U2755, P3_U2754, P3_U2753, P3_U2752, P3_U2751, P3_U2750, P3_U2749, 
        P3_U2748, P3_U2747, P3_U2746, P3_U2745, P3_U2744, P3_U2743, P3_U2742, 
        P3_U2741, P3_U2740, P3_U2739, P3_U2738, P3_U2737, P3_U2736, P3_U2735, 
        P3_U2734, P3_U2733, P3_U2732, P3_U2731, P3_U2730, P3_U2729, P3_U2728, 
        P3_U2727, P3_U2726, P3_U2725, P3_U2724, P3_U2723, P3_U2722, P3_U2721, 
        P3_U2720, P3_U2719, P3_U2718, P3_U2717, P3_U2716, P3_U2715, P3_U2714, 
        P3_U2713, P3_U2712, P3_U2711, P3_U2710, P3_U2709, P3_U2708, P3_U2707, 
        P3_U2706, P3_U2705, P3_U2704, P3_U2703, P3_U2702, P3_U2701, P3_U2700, 
        P3_U2699, P3_U2698, P3_U2697, P3_U2696, P3_U2695, P3_U2694, P3_U2693, 
        P3_U2692, P3_U2691, P3_U2690, P3_U2689, P3_U2688, P3_U2687, P3_U2686, 
        P3_U2685, P3_U2684, P3_U2683, P3_U2682, P3_U2681, P3_U2680, P3_U2679, 
        P3_U2678, P3_U2677, P3_U2676, P3_U2675, P3_U2674, P3_U2673, P3_U2672, 
        P3_U2671, P3_U2670, P3_U2669, P3_U2668, P3_U2667, P3_U2666, P3_U2665, 
        P3_U2664, P3_U2663, P3_U2662, P3_U2661, P3_U2660, P3_U2659, P3_U2658, 
        P3_U2657, P3_U2656, P3_U2655, P3_U2654, P3_U2653, P3_U2652, P3_U2651, 
        P3_U2650, P3_U2649, P3_U2648, P3_U2647, P3_U2646, P3_U2645, P3_U2644, 
        P3_U2643, P3_U2642, P3_U2641, P3_U2640, P3_U2639, P3_U3292, P3_U2638, 
        P3_U3293, P3_U3294, P3_U2637, P3_U3295, P3_U2636, P3_U3296, P3_U2635, 
        P3_U3297, P3_U2634, P3_U2633, P3_U3298, P3_U3299, P2_U3585, P2_U3586, 
        P2_U3587, P2_U3588, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, 
        P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, 
        P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, 
        P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, 
        P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210, P2_U3209, 
        P2_U3591, P2_U3592, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, 
        P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, 
        P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, 
        P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3184, P2_U3183, 
        P2_U3182, P2_U3181, P2_U3180, P2_U3179, P2_U3593, P2_U3178, P2_U3177, 
        P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172, P2_U3171, P2_U3170, 
        P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165, P2_U3164, P2_U3163, 
        P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158, P2_U3157, P2_U3156, 
        P2_U3155, P2_U3154, P2_U3153, P2_U3152, P2_U3151, P2_U3150, P2_U3149, 
        P2_U3148, P2_U3147, P2_U3146, P2_U3145, P2_U3144, P2_U3143, P2_U3142, 
        P2_U3141, P2_U3140, P2_U3139, P2_U3138, P2_U3137, P2_U3136, P2_U3135, 
        P2_U3134, P2_U3133, P2_U3132, P2_U3131, P2_U3130, P2_U3129, P2_U3128, 
        P2_U3127, P2_U3126, P2_U3125, P2_U3124, P2_U3123, P2_U3122, P2_U3121, 
        P2_U3120, P2_U3119, P2_U3118, P2_U3117, P2_U3116, P2_U3115, P2_U3114, 
        P2_U3113, P2_U3112, P2_U3111, P2_U3110, P2_U3109, P2_U3108, P2_U3107, 
        P2_U3106, P2_U3105, P2_U3104, P2_U3103, P2_U3102, P2_U3101, P2_U3100, 
        P2_U3099, P2_U3098, P2_U3097, P2_U3096, P2_U3095, P2_U3094, P2_U3093, 
        P2_U3092, P2_U3091, P2_U3090, P2_U3089, P2_U3088, P2_U3087, P2_U3086, 
        P2_U3085, P2_U3084, P2_U3083, P2_U3082, P2_U3081, P2_U3080, P2_U3079, 
        P2_U3078, P2_U3077, P2_U3076, P2_U3075, P2_U3074, P2_U3073, P2_U3072, 
        P2_U3071, P2_U3070, P2_U3069, P2_U3068, P2_U3067, P2_U3066, P2_U3065, 
        P2_U3064, P2_U3063, P2_U3062, P2_U3061, P2_U3060, P2_U3059, P2_U3058, 
        P2_U3057, P2_U3056, P2_U3055, P2_U3054, P2_U3053, P2_U3052, P2_U3051, 
        P2_U3050, P2_U3049, P2_U3048, P2_U3595, P2_U3596, P2_U3599, P2_U3600, 
        P2_U3601, P2_U3047, P2_U3602, P2_U3603, P2_U3604, P2_U3605, P2_U3046, 
        P2_U3045, P2_U3044, P2_U3043, P2_U3042, P2_U3041, P2_U3040, P2_U3039, 
        P2_U3038, P2_U3037, P2_U3036, P2_U3035, P2_U3034, P2_U3033, P2_U3032, 
        P2_U3031, P2_U3030, P2_U3029, P2_U3028, P2_U3027, P2_U3026, P2_U3025, 
        P2_U3024, P2_U3023, P2_U3022, P2_U3021, P2_U3020, P2_U3019, P2_U3018, 
        P2_U3017, P2_U3016, P2_U3015, P2_U3014, P2_U3013, P2_U3012, P2_U3011, 
        P2_U3010, P2_U3009, P2_U3008, P2_U3007, P2_U3006, P2_U3005, P2_U3004, 
        P2_U3003, P2_U3002, P2_U3001, P2_U3000, P2_U2999, P2_U2998, P2_U2997, 
        P2_U2996, P2_U2995, P2_U2994, P2_U2993, P2_U2992, P2_U2991, P2_U2990, 
        P2_U2989, P2_U2988, P2_U2987, P2_U2986, P2_U2985, P2_U2984, P2_U2983, 
        P2_U2982, P2_U2981, P2_U2980, P2_U2979, P2_U2978, P2_U2977, P2_U2976, 
        P2_U2975, P2_U2974, P2_U2973, P2_U2972, P2_U2971, P2_U2970, P2_U2969, 
        P2_U2968, P2_U2967, P2_U2966, P2_U2965, P2_U2964, P2_U2963, P2_U2962, 
        P2_U2961, P2_U2960, P2_U2959, P2_U2958, P2_U2957, P2_U2956, P2_U2955, 
        P2_U2954, P2_U2953, P2_U2952, P2_U2951, P2_U2950, P2_U2949, P2_U2948, 
        P2_U2947, P2_U2946, P2_U2945, P2_U2944, P2_U2943, P2_U2942, P2_U2941, 
        P2_U2940, P2_U2939, P2_U2938, P2_U2937, P2_U2936, P2_U2935, P2_U2934, 
        P2_U2933, P2_U2932, P2_U2931, P2_U2930, P2_U2929, P2_U2928, P2_U2927, 
        P2_U2926, P2_U2925, P2_U2924, P2_U2923, P2_U2922, P2_U2921, P2_U2920, 
        P2_U2919, P2_U2918, P2_U2917, P2_U2916, P2_U2915, P2_U2914, P2_U2913, 
        P2_U2912, P2_U2911, P2_U2910, P2_U2909, P2_U2908, P2_U2907, P2_U2906, 
        P2_U2905, P2_U2904, P2_U2903, P2_U2902, P2_U2901, P2_U2900, P2_U2899, 
        P2_U2898, P2_U2897, P2_U2896, P2_U2895, P2_U2894, P2_U2893, P2_U2892, 
        P2_U2891, P2_U2890, P2_U2889, P2_U2888, P2_U2887, P2_U2886, P2_U2885, 
        P2_U2884, P2_U2883, P2_U2882, P2_U2881, P2_U2880, P2_U2879, P2_U2878, 
        P2_U2877, P2_U2876, P2_U2875, P2_U2874, P2_U2873, P2_U2872, P2_U2871, 
        P2_U2870, P2_U2869, P2_U2868, P2_U2867, P2_U2866, P2_U2865, P2_U2864, 
        P2_U2863, P2_U2862, P2_U2861, P2_U2860, P2_U2859, P2_U2858, P2_U2857, 
        P2_U2856, P2_U2855, P2_U2854, P2_U2853, P2_U2852, P2_U2851, P2_U2850, 
        P2_U2849, P2_U2848, P2_U2847, P2_U2846, P2_U2845, P2_U2844, P2_U2843, 
        P2_U2842, P2_U2841, P2_U2840, P2_U2839, P2_U2838, P2_U2837, P2_U2836, 
        P2_U2835, P2_U2834, P2_U2833, P2_U2832, P2_U2831, P2_U2830, P2_U2829, 
        P2_U2828, P2_U2827, P2_U2826, P2_U2825, P2_U2824, P2_U2823, P2_U2822, 
        P2_U2821, P2_U2820, P2_U3608, P2_U2819, P2_U3609, P2_U2818, P2_U3610, 
        P2_U2817, P2_U3611, P2_U2816, P2_U2815, P2_U3612, P2_U2814, P1_U3458, 
        P1_U3459, P1_U3460, P1_U3461, P1_U3226, P1_U3225, P1_U3224, P1_U3223, 
        P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, P1_U3216, 
        P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, P1_U3210, P1_U3209, 
        P1_U3208, P1_U3207, P1_U3206, P1_U3205, P1_U3204, P1_U3203, P1_U3202, 
        P1_U3201, P1_U3200, P1_U3199, P1_U3198, P1_U3197, P1_U3196, P1_U3195, 
        P1_U3194, P1_U3464, P1_U3465, P1_U3193, P1_U3192, P1_U3191, P1_U3190, 
        P1_U3189, P1_U3188, P1_U3187, P1_U3186, P1_U3185, P1_U3184, P1_U3183, 
        P1_U3182, P1_U3181, P1_U3180, P1_U3179, P1_U3178, P1_U3177, P1_U3176, 
        P1_U3175, P1_U3174, P1_U3173, P1_U3172, P1_U3171, P1_U3170, P1_U3169, 
        P1_U3168, P1_U3167, P1_U3166, P1_U3165, P1_U3164, P1_U3466, P1_U3163, 
        P1_U3162, P1_U3161, P1_U3160, P1_U3159, P1_U3158, P1_U3157, P1_U3156, 
        P1_U3155, P1_U3154, P1_U3153, P1_U3152, P1_U3151, P1_U3150, P1_U3149, 
        P1_U3148, P1_U3147, P1_U3146, P1_U3145, P1_U3144, P1_U3143, P1_U3142, 
        P1_U3141, P1_U3140, P1_U3139, P1_U3138, P1_U3137, P1_U3136, P1_U3135, 
        P1_U3134, P1_U3133, P1_U3132, P1_U3131, P1_U3130, P1_U3129, P1_U3128, 
        P1_U3127, P1_U3126, P1_U3125, P1_U3124, P1_U3123, P1_U3122, P1_U3121, 
        P1_U3120, P1_U3119, P1_U3118, P1_U3117, P1_U3116, P1_U3115, P1_U3114, 
        P1_U3113, P1_U3112, P1_U3111, P1_U3110, P1_U3109, P1_U3108, P1_U3107, 
        P1_U3106, P1_U3105, P1_U3104, P1_U3103, P1_U3102, P1_U3101, P1_U3100, 
        P1_U3099, P1_U3098, P1_U3097, P1_U3096, P1_U3095, P1_U3094, P1_U3093, 
        P1_U3092, P1_U3091, P1_U3090, P1_U3089, P1_U3088, P1_U3087, P1_U3086, 
        P1_U3085, P1_U3084, P1_U3083, P1_U3082, P1_U3081, P1_U3080, P1_U3079, 
        P1_U3078, P1_U3077, P1_U3076, P1_U3075, P1_U3074, P1_U3073, P1_U3072, 
        P1_U3071, P1_U3070, P1_U3069, P1_U3068, P1_U3067, P1_U3066, P1_U3065, 
        P1_U3064, P1_U3063, P1_U3062, P1_U3061, P1_U3060, P1_U3059, P1_U3058, 
        P1_U3057, P1_U3056, P1_U3055, P1_U3054, P1_U3053, P1_U3052, P1_U3051, 
        P1_U3050, P1_U3049, P1_U3048, P1_U3047, P1_U3046, P1_U3045, P1_U3044, 
        P1_U3043, P1_U3042, P1_U3041, P1_U3040, P1_U3039, P1_U3038, P1_U3037, 
        P1_U3036, P1_U3035, P1_U3034, P1_U3033, P1_U3468, P1_U3469, P1_U3472, 
        P1_U3473, P1_U3474, P1_U3032, P1_U3475, P1_U3476, P1_U3477, P1_U3478, 
        P1_U3031, P1_U3030, P1_U3029, P1_U3028, P1_U3027, P1_U3026, P1_U3025, 
        P1_U3024, P1_U3023, P1_U3022, P1_U3021, P1_U3020, P1_U3019, P1_U3018, 
        P1_U3017, P1_U3016, P1_U3015, P1_U3014, P1_U3013, P1_U3012, P1_U3011, 
        P1_U3010, P1_U3009, P1_U3008, P1_U3007, P1_U3006, P1_U3005, P1_U3004, 
        P1_U3003, P1_U3002, P1_U3001, P1_U3000, P1_U2999, P1_U2998, P1_U2997, 
        P1_U2996, P1_U2995, P1_U2994, P1_U2993, P1_U2992, P1_U2991, P1_U2990, 
        P1_U2989, P1_U2988, P1_U2987, P1_U2986, P1_U2985, P1_U2984, P1_U2983, 
        P1_U2982, P1_U2981, P1_U2980, P1_U2979, P1_U2978, P1_U2977, P1_U2976, 
        P1_U2975, P1_U2974, P1_U2973, P1_U2972, P1_U2971, P1_U2970, P1_U2969, 
        P1_U2968, P1_U2967, P1_U2966, P1_U2965, P1_U2964, P1_U2963, P1_U2962, 
        P1_U2961, P1_U2960, P1_U2959, P1_U2958, P1_U2957, P1_U2956, P1_U2955, 
        P1_U2954, P1_U2953, P1_U2952, P1_U2951, P1_U2950, P1_U2949, P1_U2948, 
        P1_U2947, P1_U2946, P1_U2945, P1_U2944, P1_U2943, P1_U2942, P1_U2941, 
        P1_U2940, P1_U2939, P1_U2938, P1_U2937, P1_U2936, P1_U2935, P1_U2934, 
        P1_U2933, P1_U2932, P1_U2931, P1_U2930, P1_U2929, P1_U2928, P1_U2927, 
        P1_U2926, P1_U2925, P1_U2924, P1_U2923, P1_U2922, P1_U2921, P1_U2920, 
        P1_U2919, P1_U2918, P1_U2917, P1_U2916, P1_U2915, P1_U2914, P1_U2913, 
        P1_U2912, P1_U2911, P1_U2910, P1_U2909, P1_U2908, P1_U2907, P1_U2906, 
        P1_U2905, P1_U2904, P1_U2903, P1_U2902, P1_U2901, P1_U2900, P1_U2899, 
        P1_U2898, P1_U2897, P1_U2896, P1_U2895, P1_U2894, P1_U2893, P1_U2892, 
        P1_U2891, P1_U2890, P1_U2889, P1_U2888, P1_U2887, P1_U2886, P1_U2885, 
        P1_U2884, P1_U2883, P1_U2882, P1_U2881, P1_U2880, P1_U2879, P1_U2878, 
        P1_U2877, P1_U2876, P1_U2875, P1_U2874, P1_U2873, P1_U2872, P1_U2871, 
        P1_U2870, P1_U2869, P1_U2868, P1_U2867, P1_U2866, P1_U2865, P1_U2864, 
        P1_U2863, P1_U2862, P1_U2861, P1_U2860, P1_U2859, P1_U2858, P1_U2857, 
        P1_U2856, P1_U2855, P1_U2854, P1_U2853, P1_U2852, P1_U2851, P1_U2850, 
        P1_U2849, P1_U2848, P1_U2847, P1_U2846, P1_U2845, P1_U2844, P1_U2843, 
        P1_U2842, P1_U2841, P1_U2840, P1_U2839, P1_U2838, P1_U2837, P1_U2836, 
        P1_U2835, P1_U2834, P1_U2833, P1_U2832, P1_U2831, P1_U2830, P1_U2829, 
        P1_U2828, P1_U2827, P1_U2826, P1_U2825, P1_U2824, P1_U2823, P1_U2822, 
        P1_U2821, P1_U2820, P1_U2819, P1_U2818, P1_U2817, P1_U2816, P1_U2815, 
        P1_U2814, P1_U2813, P1_U2812, P1_U2811, P1_U2810, P1_U2809, P1_U2808, 
        P1_U3481, P1_U2807, P1_U3482, P1_U3483, P1_U2806, P1_U3484, P1_U2805, 
        P1_U3485, P1_U2804, P1_U3486, P1_U2803, P1_U2802, P1_U3487, P1_U2801
 );
  input P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_,
         DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_,
         DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_,
         DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_,
         DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_,
         DATAI_2_, DATAI_1_, DATAI_0_, HOLD, NA, BS16, READY1, READY2,
         P1_READREQUEST_REG_SCAN_IN, P1_ADS_N_REG_SCAN_IN,
         P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, P1_D_C_N_REG_SCAN_IN,
         P1_REQUESTPENDING_REG_SCAN_IN, P1_STATEBS16_REG_SCAN_IN,
         P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, P1_W_R_N_REG_SCAN_IN,
         P1_BYTEENABLE_REG_0__SCAN_IN, P1_BYTEENABLE_REG_1__SCAN_IN,
         P1_BYTEENABLE_REG_2__SCAN_IN, P1_BYTEENABLE_REG_3__SCAN_IN,
         P1_REIP_REG_31__SCAN_IN, P1_REIP_REG_30__SCAN_IN,
         P1_REIP_REG_29__SCAN_IN, P1_REIP_REG_28__SCAN_IN,
         P1_REIP_REG_27__SCAN_IN, P1_REIP_REG_26__SCAN_IN,
         P1_REIP_REG_25__SCAN_IN, P1_REIP_REG_24__SCAN_IN,
         P1_REIP_REG_23__SCAN_IN, P1_REIP_REG_22__SCAN_IN,
         P1_REIP_REG_21__SCAN_IN, P1_REIP_REG_20__SCAN_IN,
         P1_REIP_REG_19__SCAN_IN, P1_REIP_REG_18__SCAN_IN,
         P1_REIP_REG_17__SCAN_IN, P1_REIP_REG_16__SCAN_IN,
         P1_REIP_REG_15__SCAN_IN, P1_REIP_REG_14__SCAN_IN,
         P1_REIP_REG_13__SCAN_IN, P1_REIP_REG_12__SCAN_IN,
         P1_REIP_REG_11__SCAN_IN, P1_REIP_REG_10__SCAN_IN,
         P1_REIP_REG_9__SCAN_IN, P1_REIP_REG_8__SCAN_IN,
         P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN,
         P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN,
         P1_REIP_REG_3__SCAN_IN, P1_REIP_REG_2__SCAN_IN,
         P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN,
         P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN,
         P1_EBX_REG_29__SCAN_IN, P1_EBX_REG_28__SCAN_IN,
         P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN,
         P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN,
         P1_EBX_REG_23__SCAN_IN, P1_EBX_REG_22__SCAN_IN,
         P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN,
         P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN,
         P1_EBX_REG_17__SCAN_IN, P1_EBX_REG_16__SCAN_IN,
         P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN,
         P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN,
         P1_EBX_REG_11__SCAN_IN, P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN,
         P1_EBX_REG_8__SCAN_IN, P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN,
         P1_EBX_REG_5__SCAN_IN, P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN,
         P1_EBX_REG_2__SCAN_IN, P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN,
         P1_EAX_REG_31__SCAN_IN, P1_EAX_REG_30__SCAN_IN,
         P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN,
         P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN,
         P1_EAX_REG_25__SCAN_IN, P1_EAX_REG_24__SCAN_IN,
         P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN,
         P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN,
         P1_EAX_REG_19__SCAN_IN, P1_EAX_REG_18__SCAN_IN,
         P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN,
         P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN,
         P1_EAX_REG_13__SCAN_IN, P1_EAX_REG_12__SCAN_IN,
         P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN,
         P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN,
         P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN,
         P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_UWORD_REG_0__SCAN_IN, P1_UWORD_REG_1__SCAN_IN,
         P1_UWORD_REG_2__SCAN_IN, P1_UWORD_REG_3__SCAN_IN,
         P1_UWORD_REG_4__SCAN_IN, P1_UWORD_REG_5__SCAN_IN,
         P1_UWORD_REG_6__SCAN_IN, P1_UWORD_REG_7__SCAN_IN,
         P1_UWORD_REG_8__SCAN_IN, P1_UWORD_REG_9__SCAN_IN,
         P1_UWORD_REG_10__SCAN_IN, P1_UWORD_REG_11__SCAN_IN,
         P1_UWORD_REG_12__SCAN_IN, P1_UWORD_REG_13__SCAN_IN,
         P1_UWORD_REG_14__SCAN_IN, P1_LWORD_REG_0__SCAN_IN,
         P1_LWORD_REG_1__SCAN_IN, P1_LWORD_REG_2__SCAN_IN,
         P1_LWORD_REG_3__SCAN_IN, P1_LWORD_REG_4__SCAN_IN,
         P1_LWORD_REG_5__SCAN_IN, P1_LWORD_REG_6__SCAN_IN,
         P1_LWORD_REG_7__SCAN_IN, P1_LWORD_REG_8__SCAN_IN,
         P1_LWORD_REG_9__SCAN_IN, P1_LWORD_REG_10__SCAN_IN,
         P1_LWORD_REG_11__SCAN_IN, P1_LWORD_REG_12__SCAN_IN,
         P1_LWORD_REG_13__SCAN_IN, P1_LWORD_REG_14__SCAN_IN,
         P1_LWORD_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_31__SCAN_IN,
         P1_PHYADDRPOINTER_REG_30__SCAN_IN, P1_PHYADDRPOINTER_REG_29__SCAN_IN,
         P1_PHYADDRPOINTER_REG_28__SCAN_IN, P1_PHYADDRPOINTER_REG_27__SCAN_IN,
         P1_PHYADDRPOINTER_REG_26__SCAN_IN, P1_PHYADDRPOINTER_REG_25__SCAN_IN,
         P1_PHYADDRPOINTER_REG_24__SCAN_IN, P1_PHYADDRPOINTER_REG_23__SCAN_IN,
         P1_PHYADDRPOINTER_REG_22__SCAN_IN, P1_PHYADDRPOINTER_REG_21__SCAN_IN,
         P1_PHYADDRPOINTER_REG_20__SCAN_IN, P1_PHYADDRPOINTER_REG_19__SCAN_IN,
         P1_PHYADDRPOINTER_REG_18__SCAN_IN, P1_PHYADDRPOINTER_REG_17__SCAN_IN,
         P1_PHYADDRPOINTER_REG_16__SCAN_IN, P1_PHYADDRPOINTER_REG_15__SCAN_IN,
         P1_PHYADDRPOINTER_REG_14__SCAN_IN, P1_PHYADDRPOINTER_REG_13__SCAN_IN,
         P1_PHYADDRPOINTER_REG_12__SCAN_IN, P1_PHYADDRPOINTER_REG_11__SCAN_IN,
         P1_PHYADDRPOINTER_REG_10__SCAN_IN, P1_PHYADDRPOINTER_REG_9__SCAN_IN,
         P1_PHYADDRPOINTER_REG_8__SCAN_IN, P1_PHYADDRPOINTER_REG_7__SCAN_IN,
         P1_PHYADDRPOINTER_REG_6__SCAN_IN, P1_PHYADDRPOINTER_REG_5__SCAN_IN,
         P1_PHYADDRPOINTER_REG_4__SCAN_IN, P1_PHYADDRPOINTER_REG_3__SCAN_IN,
         P1_PHYADDRPOINTER_REG_2__SCAN_IN, P1_PHYADDRPOINTER_REG_1__SCAN_IN,
         P1_PHYADDRPOINTER_REG_0__SCAN_IN, P1_INSTADDRPOINTER_REG_31__SCAN_IN,
         P1_INSTADDRPOINTER_REG_30__SCAN_IN,
         P1_INSTADDRPOINTER_REG_29__SCAN_IN,
         P1_INSTADDRPOINTER_REG_28__SCAN_IN,
         P1_INSTADDRPOINTER_REG_27__SCAN_IN,
         P1_INSTADDRPOINTER_REG_26__SCAN_IN,
         P1_INSTADDRPOINTER_REG_25__SCAN_IN,
         P1_INSTADDRPOINTER_REG_24__SCAN_IN,
         P1_INSTADDRPOINTER_REG_23__SCAN_IN,
         P1_INSTADDRPOINTER_REG_22__SCAN_IN,
         P1_INSTADDRPOINTER_REG_21__SCAN_IN,
         P1_INSTADDRPOINTER_REG_20__SCAN_IN,
         P1_INSTADDRPOINTER_REG_19__SCAN_IN,
         P1_INSTADDRPOINTER_REG_18__SCAN_IN,
         P1_INSTADDRPOINTER_REG_17__SCAN_IN,
         P1_INSTADDRPOINTER_REG_16__SCAN_IN,
         P1_INSTADDRPOINTER_REG_15__SCAN_IN,
         P1_INSTADDRPOINTER_REG_14__SCAN_IN,
         P1_INSTADDRPOINTER_REG_13__SCAN_IN,
         P1_INSTADDRPOINTER_REG_12__SCAN_IN,
         P1_INSTADDRPOINTER_REG_11__SCAN_IN,
         P1_INSTADDRPOINTER_REG_10__SCAN_IN, P1_INSTADDRPOINTER_REG_9__SCAN_IN,
         P1_INSTADDRPOINTER_REG_8__SCAN_IN, P1_INSTADDRPOINTER_REG_7__SCAN_IN,
         P1_INSTADDRPOINTER_REG_6__SCAN_IN, P1_INSTADDRPOINTER_REG_5__SCAN_IN,
         P1_INSTADDRPOINTER_REG_4__SCAN_IN, P1_INSTADDRPOINTER_REG_3__SCAN_IN,
         P1_INSTADDRPOINTER_REG_2__SCAN_IN, P1_INSTADDRPOINTER_REG_1__SCAN_IN,
         P1_INSTADDRPOINTER_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P1_INSTQUEUE_REG_0__0__SCAN_IN,
         P1_INSTQUEUE_REG_0__1__SCAN_IN, P1_INSTQUEUE_REG_0__2__SCAN_IN,
         P1_INSTQUEUE_REG_0__3__SCAN_IN, P1_INSTQUEUE_REG_0__4__SCAN_IN,
         P1_INSTQUEUE_REG_0__5__SCAN_IN, P1_INSTQUEUE_REG_0__6__SCAN_IN,
         P1_INSTQUEUE_REG_0__7__SCAN_IN, P1_INSTQUEUE_REG_1__0__SCAN_IN,
         P1_INSTQUEUE_REG_1__1__SCAN_IN, P1_INSTQUEUE_REG_1__2__SCAN_IN,
         P1_INSTQUEUE_REG_1__3__SCAN_IN, P1_INSTQUEUE_REG_1__4__SCAN_IN,
         P1_INSTQUEUE_REG_1__5__SCAN_IN, P1_INSTQUEUE_REG_1__6__SCAN_IN,
         P1_INSTQUEUE_REG_1__7__SCAN_IN, P1_INSTQUEUE_REG_2__0__SCAN_IN,
         P1_INSTQUEUE_REG_2__1__SCAN_IN, P1_INSTQUEUE_REG_2__2__SCAN_IN,
         P1_INSTQUEUE_REG_2__3__SCAN_IN, P1_INSTQUEUE_REG_2__4__SCAN_IN,
         P1_INSTQUEUE_REG_2__5__SCAN_IN, P1_INSTQUEUE_REG_2__6__SCAN_IN,
         P1_INSTQUEUE_REG_2__7__SCAN_IN, P1_INSTQUEUE_REG_3__0__SCAN_IN,
         P1_INSTQUEUE_REG_3__1__SCAN_IN, P1_INSTQUEUE_REG_3__2__SCAN_IN,
         P1_INSTQUEUE_REG_3__3__SCAN_IN, P1_INSTQUEUE_REG_3__4__SCAN_IN,
         P1_INSTQUEUE_REG_3__5__SCAN_IN, P1_INSTQUEUE_REG_3__6__SCAN_IN,
         P1_INSTQUEUE_REG_3__7__SCAN_IN, P1_INSTQUEUE_REG_4__0__SCAN_IN,
         BUF1_REG_0__SCAN_IN, BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN,
         BUF1_REG_3__SCAN_IN, BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN,
         BUF1_REG_6__SCAN_IN, BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN,
         BUF1_REG_9__SCAN_IN, BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN,
         BUF1_REG_12__SCAN_IN, BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN,
         BUF1_REG_15__SCAN_IN, BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN,
         BUF1_REG_18__SCAN_IN, BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN,
         BUF1_REG_21__SCAN_IN, BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN,
         BUF1_REG_24__SCAN_IN, BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN,
         BUF1_REG_27__SCAN_IN, BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN,
         BUF1_REG_30__SCAN_IN, BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN,
         BUF2_REG_1__SCAN_IN, BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN,
         BUF2_REG_4__SCAN_IN, BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN,
         BUF2_REG_7__SCAN_IN, BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN,
         BUF2_REG_10__SCAN_IN, BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN,
         BUF2_REG_13__SCAN_IN, BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN,
         BUF2_REG_16__SCAN_IN, BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN,
         BUF2_REG_19__SCAN_IN, BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN,
         BUF2_REG_22__SCAN_IN, BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN,
         BUF2_REG_25__SCAN_IN, BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN,
         BUF2_REG_28__SCAN_IN, BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN,
         BUF2_REG_31__SCAN_IN, READY12_REG_SCAN_IN, READY21_REG_SCAN_IN,
         READY22_REG_SCAN_IN, READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN,
         P3_BE_N_REG_2__SCAN_IN, P3_BE_N_REG_1__SCAN_IN,
         P3_BE_N_REG_0__SCAN_IN, P3_ADDRESS_REG_29__SCAN_IN,
         P3_ADDRESS_REG_28__SCAN_IN, P3_ADDRESS_REG_27__SCAN_IN,
         P3_ADDRESS_REG_26__SCAN_IN, P3_ADDRESS_REG_25__SCAN_IN,
         P3_ADDRESS_REG_24__SCAN_IN, P3_ADDRESS_REG_23__SCAN_IN,
         P3_ADDRESS_REG_22__SCAN_IN, P3_ADDRESS_REG_21__SCAN_IN,
         P3_ADDRESS_REG_20__SCAN_IN, P3_ADDRESS_REG_19__SCAN_IN,
         P3_ADDRESS_REG_18__SCAN_IN, P3_ADDRESS_REG_17__SCAN_IN,
         P3_ADDRESS_REG_16__SCAN_IN, P3_ADDRESS_REG_15__SCAN_IN,
         P3_ADDRESS_REG_14__SCAN_IN, P3_ADDRESS_REG_13__SCAN_IN,
         P3_ADDRESS_REG_12__SCAN_IN, P3_ADDRESS_REG_11__SCAN_IN,
         P3_ADDRESS_REG_10__SCAN_IN, P3_ADDRESS_REG_9__SCAN_IN,
         P3_ADDRESS_REG_8__SCAN_IN, P3_ADDRESS_REG_7__SCAN_IN,
         P3_ADDRESS_REG_6__SCAN_IN, P3_ADDRESS_REG_5__SCAN_IN,
         P3_ADDRESS_REG_4__SCAN_IN, P3_ADDRESS_REG_3__SCAN_IN,
         P3_ADDRESS_REG_2__SCAN_IN, P3_ADDRESS_REG_1__SCAN_IN,
         P3_ADDRESS_REG_0__SCAN_IN, P3_STATE_REG_2__SCAN_IN,
         P3_STATE_REG_1__SCAN_IN, P3_STATE_REG_0__SCAN_IN,
         P3_DATAWIDTH_REG_0__SCAN_IN, P3_DATAWIDTH_REG_1__SCAN_IN,
         P3_DATAWIDTH_REG_2__SCAN_IN, P3_DATAWIDTH_REG_3__SCAN_IN,
         P3_DATAWIDTH_REG_4__SCAN_IN, P3_DATAWIDTH_REG_5__SCAN_IN,
         P3_DATAWIDTH_REG_6__SCAN_IN, P3_DATAWIDTH_REG_7__SCAN_IN,
         P3_DATAWIDTH_REG_8__SCAN_IN, P3_DATAWIDTH_REG_9__SCAN_IN,
         P3_DATAWIDTH_REG_10__SCAN_IN, P3_DATAWIDTH_REG_11__SCAN_IN,
         P3_DATAWIDTH_REG_12__SCAN_IN, P3_DATAWIDTH_REG_13__SCAN_IN,
         P3_DATAWIDTH_REG_14__SCAN_IN, P3_DATAWIDTH_REG_15__SCAN_IN,
         P3_DATAWIDTH_REG_16__SCAN_IN, P3_DATAWIDTH_REG_17__SCAN_IN,
         P3_DATAWIDTH_REG_18__SCAN_IN, P3_DATAWIDTH_REG_19__SCAN_IN,
         P3_DATAWIDTH_REG_20__SCAN_IN, P3_DATAWIDTH_REG_21__SCAN_IN,
         P3_DATAWIDTH_REG_22__SCAN_IN, P3_DATAWIDTH_REG_23__SCAN_IN,
         P3_DATAWIDTH_REG_24__SCAN_IN, P3_DATAWIDTH_REG_25__SCAN_IN,
         P3_DATAWIDTH_REG_26__SCAN_IN, P3_DATAWIDTH_REG_27__SCAN_IN,
         P3_DATAWIDTH_REG_28__SCAN_IN, P3_DATAWIDTH_REG_29__SCAN_IN,
         P3_DATAWIDTH_REG_30__SCAN_IN, P3_DATAWIDTH_REG_31__SCAN_IN,
         P3_STATE2_REG_3__SCAN_IN, P3_STATE2_REG_2__SCAN_IN,
         P3_STATE2_REG_1__SCAN_IN, P3_STATE2_REG_0__SCAN_IN,
         P3_INSTQUEUE_REG_15__7__SCAN_IN, P3_INSTQUEUE_REG_15__6__SCAN_IN,
         P3_INSTQUEUE_REG_15__5__SCAN_IN, P3_INSTQUEUE_REG_15__4__SCAN_IN,
         P3_INSTQUEUE_REG_15__3__SCAN_IN, P3_INSTQUEUE_REG_15__2__SCAN_IN,
         P3_INSTQUEUE_REG_15__1__SCAN_IN, P3_INSTQUEUE_REG_15__0__SCAN_IN,
         P3_INSTQUEUE_REG_14__7__SCAN_IN, P3_INSTQUEUE_REG_14__6__SCAN_IN,
         P3_INSTQUEUE_REG_14__5__SCAN_IN, P3_INSTQUEUE_REG_14__4__SCAN_IN,
         P3_INSTQUEUE_REG_14__3__SCAN_IN, P3_INSTQUEUE_REG_14__2__SCAN_IN,
         P3_INSTQUEUE_REG_14__1__SCAN_IN, P3_INSTQUEUE_REG_14__0__SCAN_IN,
         P3_INSTQUEUE_REG_13__7__SCAN_IN, P3_INSTQUEUE_REG_13__6__SCAN_IN,
         P3_INSTQUEUE_REG_13__5__SCAN_IN, P3_INSTQUEUE_REG_13__4__SCAN_IN,
         P3_INSTQUEUE_REG_13__3__SCAN_IN, P3_INSTQUEUE_REG_13__2__SCAN_IN,
         P3_INSTQUEUE_REG_13__1__SCAN_IN, P3_INSTQUEUE_REG_13__0__SCAN_IN,
         P3_INSTQUEUE_REG_12__7__SCAN_IN, P3_INSTQUEUE_REG_12__6__SCAN_IN,
         P3_INSTQUEUE_REG_12__5__SCAN_IN, P3_INSTQUEUE_REG_12__4__SCAN_IN,
         P3_INSTQUEUE_REG_12__3__SCAN_IN, P3_INSTQUEUE_REG_12__2__SCAN_IN,
         P3_INSTQUEUE_REG_12__1__SCAN_IN, P3_INSTQUEUE_REG_12__0__SCAN_IN,
         P3_INSTQUEUE_REG_11__7__SCAN_IN, P3_INSTQUEUE_REG_11__6__SCAN_IN,
         P3_INSTQUEUE_REG_11__5__SCAN_IN, P3_INSTQUEUE_REG_11__4__SCAN_IN,
         P3_INSTQUEUE_REG_11__3__SCAN_IN, P3_INSTQUEUE_REG_11__2__SCAN_IN,
         P3_INSTQUEUE_REG_11__1__SCAN_IN, P3_INSTQUEUE_REG_11__0__SCAN_IN,
         P3_INSTQUEUE_REG_10__7__SCAN_IN, P3_INSTQUEUE_REG_10__6__SCAN_IN,
         P3_INSTQUEUE_REG_10__5__SCAN_IN, P3_INSTQUEUE_REG_10__4__SCAN_IN,
         P3_INSTQUEUE_REG_10__3__SCAN_IN, P3_INSTQUEUE_REG_10__2__SCAN_IN,
         P3_INSTQUEUE_REG_10__1__SCAN_IN, P3_INSTQUEUE_REG_10__0__SCAN_IN,
         P3_INSTQUEUE_REG_9__7__SCAN_IN, P3_INSTQUEUE_REG_9__6__SCAN_IN,
         P3_INSTQUEUE_REG_9__5__SCAN_IN, P3_INSTQUEUE_REG_9__4__SCAN_IN,
         P3_INSTQUEUE_REG_9__3__SCAN_IN, P3_INSTQUEUE_REG_9__2__SCAN_IN,
         P3_INSTQUEUE_REG_9__1__SCAN_IN, P3_INSTQUEUE_REG_9__0__SCAN_IN,
         P3_INSTQUEUE_REG_8__7__SCAN_IN, P3_INSTQUEUE_REG_8__6__SCAN_IN,
         P3_INSTQUEUE_REG_8__5__SCAN_IN, P3_INSTQUEUE_REG_8__4__SCAN_IN,
         P3_INSTQUEUE_REG_8__3__SCAN_IN, P3_INSTQUEUE_REG_8__2__SCAN_IN,
         P3_INSTQUEUE_REG_8__1__SCAN_IN, P3_INSTQUEUE_REG_8__0__SCAN_IN,
         P3_INSTQUEUE_REG_7__7__SCAN_IN, P3_INSTQUEUE_REG_7__6__SCAN_IN,
         P3_INSTQUEUE_REG_7__5__SCAN_IN, P3_INSTQUEUE_REG_7__4__SCAN_IN,
         P3_INSTQUEUE_REG_7__3__SCAN_IN, P3_INSTQUEUE_REG_7__2__SCAN_IN,
         P3_INSTQUEUE_REG_7__1__SCAN_IN, P3_INSTQUEUE_REG_7__0__SCAN_IN,
         P3_INSTQUEUE_REG_6__7__SCAN_IN, P3_INSTQUEUE_REG_6__6__SCAN_IN,
         P3_INSTQUEUE_REG_6__5__SCAN_IN, P3_INSTQUEUE_REG_6__4__SCAN_IN,
         P3_INSTQUEUE_REG_6__3__SCAN_IN, P3_INSTQUEUE_REG_6__2__SCAN_IN,
         P3_INSTQUEUE_REG_6__1__SCAN_IN, P3_INSTQUEUE_REG_6__0__SCAN_IN,
         P3_INSTQUEUE_REG_5__7__SCAN_IN, P3_INSTQUEUE_REG_5__6__SCAN_IN,
         P3_INSTQUEUE_REG_5__5__SCAN_IN, P3_INSTQUEUE_REG_5__4__SCAN_IN,
         P3_INSTQUEUE_REG_5__3__SCAN_IN, P3_INSTQUEUE_REG_5__2__SCAN_IN,
         P3_INSTQUEUE_REG_5__1__SCAN_IN, P3_INSTQUEUE_REG_5__0__SCAN_IN,
         P3_INSTQUEUE_REG_4__7__SCAN_IN, P3_INSTQUEUE_REG_4__6__SCAN_IN,
         P3_INSTQUEUE_REG_4__5__SCAN_IN, P3_INSTQUEUE_REG_4__4__SCAN_IN,
         P3_INSTQUEUE_REG_4__3__SCAN_IN, P3_INSTQUEUE_REG_4__2__SCAN_IN,
         P3_INSTQUEUE_REG_4__1__SCAN_IN, P3_INSTQUEUE_REG_4__0__SCAN_IN,
         P3_INSTQUEUE_REG_3__7__SCAN_IN, P3_INSTQUEUE_REG_3__6__SCAN_IN,
         P3_INSTQUEUE_REG_3__5__SCAN_IN, P3_INSTQUEUE_REG_3__4__SCAN_IN,
         P3_INSTQUEUE_REG_3__3__SCAN_IN, P3_INSTQUEUE_REG_3__2__SCAN_IN,
         P3_INSTQUEUE_REG_3__1__SCAN_IN, P3_INSTQUEUE_REG_3__0__SCAN_IN,
         P3_INSTQUEUE_REG_2__7__SCAN_IN, P3_INSTQUEUE_REG_2__6__SCAN_IN,
         P3_INSTQUEUE_REG_2__5__SCAN_IN, P3_INSTQUEUE_REG_2__4__SCAN_IN,
         P3_INSTQUEUE_REG_2__3__SCAN_IN, P3_INSTQUEUE_REG_2__2__SCAN_IN,
         P3_INSTQUEUE_REG_2__1__SCAN_IN, P3_INSTQUEUE_REG_2__0__SCAN_IN,
         P3_INSTQUEUE_REG_1__7__SCAN_IN, P3_INSTQUEUE_REG_1__6__SCAN_IN,
         P3_INSTQUEUE_REG_1__5__SCAN_IN, P3_INSTQUEUE_REG_1__4__SCAN_IN,
         P3_INSTQUEUE_REG_1__3__SCAN_IN, P3_INSTQUEUE_REG_1__2__SCAN_IN,
         P3_INSTQUEUE_REG_1__1__SCAN_IN, P3_INSTQUEUE_REG_1__0__SCAN_IN,
         P3_INSTQUEUE_REG_0__7__SCAN_IN, P3_INSTQUEUE_REG_0__6__SCAN_IN,
         P3_INSTQUEUE_REG_0__5__SCAN_IN, P3_INSTQUEUE_REG_0__4__SCAN_IN,
         P3_INSTQUEUE_REG_0__3__SCAN_IN, P3_INSTQUEUE_REG_0__2__SCAN_IN,
         P3_INSTQUEUE_REG_0__1__SCAN_IN, P3_INSTQUEUE_REG_0__0__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN,
         P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN,
         P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN,
         P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN,
         P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN,
         P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN,
         P3_INSTADDRPOINTER_REG_11__SCAN_IN,
         P3_INSTADDRPOINTER_REG_12__SCAN_IN,
         P3_INSTADDRPOINTER_REG_13__SCAN_IN,
         P3_INSTADDRPOINTER_REG_14__SCAN_IN,
         P3_INSTADDRPOINTER_REG_15__SCAN_IN,
         P3_INSTADDRPOINTER_REG_16__SCAN_IN,
         P3_INSTADDRPOINTER_REG_17__SCAN_IN,
         P3_INSTADDRPOINTER_REG_18__SCAN_IN,
         P3_INSTADDRPOINTER_REG_19__SCAN_IN,
         P3_INSTADDRPOINTER_REG_20__SCAN_IN,
         P3_INSTADDRPOINTER_REG_21__SCAN_IN,
         P3_INSTADDRPOINTER_REG_22__SCAN_IN,
         P3_INSTADDRPOINTER_REG_23__SCAN_IN,
         P3_INSTADDRPOINTER_REG_24__SCAN_IN,
         P3_INSTADDRPOINTER_REG_25__SCAN_IN,
         P3_INSTADDRPOINTER_REG_26__SCAN_IN,
         P3_INSTADDRPOINTER_REG_27__SCAN_IN,
         P3_INSTADDRPOINTER_REG_28__SCAN_IN,
         P3_INSTADDRPOINTER_REG_29__SCAN_IN,
         P3_INSTADDRPOINTER_REG_30__SCAN_IN,
         P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN,
         P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN,
         P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN,
         P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN,
         P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN,
         P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN,
         P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN,
         P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN,
         P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN,
         P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN,
         P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN,
         P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN,
         P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN,
         P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN,
         P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN,
         P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN,
         P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN,
         P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN,
         P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN,
         P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN,
         P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN,
         P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN,
         P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN,
         P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN,
         P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN,
         P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN,
         P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN,
         P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN,
         P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN,
         P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN,
         P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN,
         P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN,
         P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN,
         P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN,
         P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN,
         P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN,
         P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN,
         P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN,
         P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN,
         P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN,
         P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN,
         P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN,
         P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN,
         P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN,
         P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN,
         P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN,
         P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN,
         P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN,
         P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN,
         P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN,
         P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN,
         P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN,
         P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN,
         P3_EAX_REG_14__SCAN_IN, P3_EAX_REG_15__SCAN_IN,
         P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN,
         P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN,
         P3_EAX_REG_20__SCAN_IN, P3_EAX_REG_21__SCAN_IN,
         P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN,
         P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN,
         P3_EAX_REG_26__SCAN_IN, P3_EAX_REG_27__SCAN_IN,
         P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN,
         P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN,
         P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN,
         P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN,
         P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN,
         P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN,
         P3_EBX_REG_12__SCAN_IN, P3_EBX_REG_13__SCAN_IN,
         P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN,
         P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN,
         P3_EBX_REG_18__SCAN_IN, P3_EBX_REG_19__SCAN_IN,
         P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN,
         P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN,
         P3_EBX_REG_24__SCAN_IN, P3_EBX_REG_25__SCAN_IN,
         P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN,
         P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN,
         P3_EBX_REG_30__SCAN_IN, P3_EBX_REG_31__SCAN_IN,
         P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN,
         P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN,
         P3_REIP_REG_4__SCAN_IN, P3_REIP_REG_5__SCAN_IN,
         P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN,
         P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN,
         P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN,
         P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN,
         P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN,
         P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN,
         P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN,
         P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN,
         P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN,
         P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN,
         P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN,
         P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN,
         P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN,
         P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN,
         P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN,
         P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN,
         P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN,
         P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN,
         P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN,
         P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN,
         P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN,
         P2_BE_N_REG_0__SCAN_IN, P2_ADDRESS_REG_29__SCAN_IN,
         P2_ADDRESS_REG_28__SCAN_IN, P2_ADDRESS_REG_27__SCAN_IN,
         P2_ADDRESS_REG_26__SCAN_IN, P2_ADDRESS_REG_25__SCAN_IN,
         P2_ADDRESS_REG_24__SCAN_IN, P2_ADDRESS_REG_23__SCAN_IN,
         P2_ADDRESS_REG_22__SCAN_IN, P2_ADDRESS_REG_21__SCAN_IN,
         P2_ADDRESS_REG_20__SCAN_IN, P2_ADDRESS_REG_19__SCAN_IN,
         P2_ADDRESS_REG_18__SCAN_IN, P2_ADDRESS_REG_17__SCAN_IN,
         P2_ADDRESS_REG_16__SCAN_IN, P2_ADDRESS_REG_15__SCAN_IN,
         P2_ADDRESS_REG_14__SCAN_IN, P2_ADDRESS_REG_13__SCAN_IN,
         P2_ADDRESS_REG_12__SCAN_IN, P2_ADDRESS_REG_11__SCAN_IN,
         P2_ADDRESS_REG_10__SCAN_IN, P2_ADDRESS_REG_9__SCAN_IN,
         P2_ADDRESS_REG_8__SCAN_IN, P2_ADDRESS_REG_7__SCAN_IN,
         P2_ADDRESS_REG_6__SCAN_IN, P2_ADDRESS_REG_5__SCAN_IN,
         P2_ADDRESS_REG_4__SCAN_IN, P2_ADDRESS_REG_3__SCAN_IN,
         P2_ADDRESS_REG_2__SCAN_IN, P2_ADDRESS_REG_1__SCAN_IN,
         P2_ADDRESS_REG_0__SCAN_IN, P2_STATE_REG_2__SCAN_IN,
         P2_STATE_REG_1__SCAN_IN, P2_STATE_REG_0__SCAN_IN,
         P2_DATAWIDTH_REG_0__SCAN_IN, P2_DATAWIDTH_REG_1__SCAN_IN,
         P2_DATAWIDTH_REG_2__SCAN_IN, P2_DATAWIDTH_REG_3__SCAN_IN,
         P2_DATAWIDTH_REG_4__SCAN_IN, P2_DATAWIDTH_REG_5__SCAN_IN,
         P2_DATAWIDTH_REG_6__SCAN_IN, P2_DATAWIDTH_REG_7__SCAN_IN,
         P2_DATAWIDTH_REG_8__SCAN_IN, P2_DATAWIDTH_REG_9__SCAN_IN,
         P2_DATAWIDTH_REG_10__SCAN_IN, P2_DATAWIDTH_REG_11__SCAN_IN,
         P2_DATAWIDTH_REG_12__SCAN_IN, P2_DATAWIDTH_REG_13__SCAN_IN,
         P2_DATAWIDTH_REG_14__SCAN_IN, P2_DATAWIDTH_REG_15__SCAN_IN,
         P2_DATAWIDTH_REG_16__SCAN_IN, P2_DATAWIDTH_REG_17__SCAN_IN,
         P2_DATAWIDTH_REG_18__SCAN_IN, P2_DATAWIDTH_REG_19__SCAN_IN,
         P2_DATAWIDTH_REG_20__SCAN_IN, P2_DATAWIDTH_REG_21__SCAN_IN,
         P2_DATAWIDTH_REG_22__SCAN_IN, P2_DATAWIDTH_REG_23__SCAN_IN,
         P2_DATAWIDTH_REG_24__SCAN_IN, P2_DATAWIDTH_REG_25__SCAN_IN,
         P2_DATAWIDTH_REG_26__SCAN_IN, P2_DATAWIDTH_REG_27__SCAN_IN,
         P2_DATAWIDTH_REG_28__SCAN_IN, P2_DATAWIDTH_REG_29__SCAN_IN,
         P2_DATAWIDTH_REG_30__SCAN_IN, P2_DATAWIDTH_REG_31__SCAN_IN,
         P2_STATE2_REG_3__SCAN_IN, P2_STATE2_REG_2__SCAN_IN,
         P2_STATE2_REG_1__SCAN_IN, P2_STATE2_REG_0__SCAN_IN,
         P2_INSTQUEUE_REG_15__7__SCAN_IN, P2_INSTQUEUE_REG_15__6__SCAN_IN,
         P2_INSTQUEUE_REG_15__5__SCAN_IN, P2_INSTQUEUE_REG_15__4__SCAN_IN,
         P2_INSTQUEUE_REG_15__3__SCAN_IN, P2_INSTQUEUE_REG_15__2__SCAN_IN,
         P2_INSTQUEUE_REG_15__1__SCAN_IN, P2_INSTQUEUE_REG_15__0__SCAN_IN,
         P2_INSTQUEUE_REG_14__7__SCAN_IN, P2_INSTQUEUE_REG_14__6__SCAN_IN,
         P2_INSTQUEUE_REG_14__5__SCAN_IN, P2_INSTQUEUE_REG_14__4__SCAN_IN,
         P2_INSTQUEUE_REG_14__3__SCAN_IN, P2_INSTQUEUE_REG_14__2__SCAN_IN,
         P2_INSTQUEUE_REG_14__1__SCAN_IN, P2_INSTQUEUE_REG_14__0__SCAN_IN,
         P2_INSTQUEUE_REG_13__7__SCAN_IN, P2_INSTQUEUE_REG_13__6__SCAN_IN,
         P2_INSTQUEUE_REG_13__5__SCAN_IN, P2_INSTQUEUE_REG_13__4__SCAN_IN,
         P2_INSTQUEUE_REG_13__3__SCAN_IN, P2_INSTQUEUE_REG_13__2__SCAN_IN,
         P2_INSTQUEUE_REG_13__1__SCAN_IN, P2_INSTQUEUE_REG_13__0__SCAN_IN,
         P2_INSTQUEUE_REG_12__7__SCAN_IN, P2_INSTQUEUE_REG_12__6__SCAN_IN,
         P2_INSTQUEUE_REG_12__5__SCAN_IN, P2_INSTQUEUE_REG_12__4__SCAN_IN,
         P2_INSTQUEUE_REG_12__3__SCAN_IN, P2_INSTQUEUE_REG_12__2__SCAN_IN,
         P2_INSTQUEUE_REG_12__1__SCAN_IN, P2_INSTQUEUE_REG_12__0__SCAN_IN,
         P2_INSTQUEUE_REG_11__7__SCAN_IN, P2_INSTQUEUE_REG_11__6__SCAN_IN,
         P2_INSTQUEUE_REG_11__5__SCAN_IN, P2_INSTQUEUE_REG_11__4__SCAN_IN,
         P2_INSTQUEUE_REG_11__3__SCAN_IN, P2_INSTQUEUE_REG_11__2__SCAN_IN,
         P2_INSTQUEUE_REG_11__1__SCAN_IN, P2_INSTQUEUE_REG_11__0__SCAN_IN,
         P2_INSTQUEUE_REG_10__7__SCAN_IN, P2_INSTQUEUE_REG_10__6__SCAN_IN,
         P2_INSTQUEUE_REG_10__5__SCAN_IN, P2_INSTQUEUE_REG_10__4__SCAN_IN,
         P2_INSTQUEUE_REG_10__3__SCAN_IN, P2_INSTQUEUE_REG_10__2__SCAN_IN,
         P2_INSTQUEUE_REG_10__1__SCAN_IN, P2_INSTQUEUE_REG_10__0__SCAN_IN,
         P2_INSTQUEUE_REG_9__7__SCAN_IN, P2_INSTQUEUE_REG_9__6__SCAN_IN,
         P2_INSTQUEUE_REG_9__5__SCAN_IN, P2_INSTQUEUE_REG_9__4__SCAN_IN,
         P2_INSTQUEUE_REG_9__3__SCAN_IN, P2_INSTQUEUE_REG_9__2__SCAN_IN,
         P2_INSTQUEUE_REG_9__1__SCAN_IN, P2_INSTQUEUE_REG_9__0__SCAN_IN,
         P2_INSTQUEUE_REG_8__7__SCAN_IN, P2_INSTQUEUE_REG_8__6__SCAN_IN,
         P2_INSTQUEUE_REG_8__5__SCAN_IN, P2_INSTQUEUE_REG_8__4__SCAN_IN,
         P2_INSTQUEUE_REG_8__3__SCAN_IN, P2_INSTQUEUE_REG_8__2__SCAN_IN,
         P2_INSTQUEUE_REG_8__1__SCAN_IN, P2_INSTQUEUE_REG_8__0__SCAN_IN,
         P2_INSTQUEUE_REG_7__7__SCAN_IN, P2_INSTQUEUE_REG_7__6__SCAN_IN,
         P2_INSTQUEUE_REG_7__5__SCAN_IN, P2_INSTQUEUE_REG_7__4__SCAN_IN,
         P2_INSTQUEUE_REG_7__3__SCAN_IN, P2_INSTQUEUE_REG_7__2__SCAN_IN,
         P2_INSTQUEUE_REG_7__1__SCAN_IN, P2_INSTQUEUE_REG_7__0__SCAN_IN,
         P2_INSTQUEUE_REG_6__7__SCAN_IN, P2_INSTQUEUE_REG_6__6__SCAN_IN,
         P2_INSTQUEUE_REG_6__5__SCAN_IN, P2_INSTQUEUE_REG_6__4__SCAN_IN,
         P2_INSTQUEUE_REG_6__3__SCAN_IN, P2_INSTQUEUE_REG_6__2__SCAN_IN,
         P2_INSTQUEUE_REG_6__1__SCAN_IN, P2_INSTQUEUE_REG_6__0__SCAN_IN,
         P2_INSTQUEUE_REG_5__7__SCAN_IN, P2_INSTQUEUE_REG_5__6__SCAN_IN,
         P2_INSTQUEUE_REG_5__5__SCAN_IN, P2_INSTQUEUE_REG_5__4__SCAN_IN,
         P2_INSTQUEUE_REG_5__3__SCAN_IN, P2_INSTQUEUE_REG_5__2__SCAN_IN,
         P2_INSTQUEUE_REG_5__1__SCAN_IN, P2_INSTQUEUE_REG_5__0__SCAN_IN,
         P2_INSTQUEUE_REG_4__7__SCAN_IN, P2_INSTQUEUE_REG_4__6__SCAN_IN,
         P2_INSTQUEUE_REG_4__5__SCAN_IN, P2_INSTQUEUE_REG_4__4__SCAN_IN,
         P2_INSTQUEUE_REG_4__3__SCAN_IN, P2_INSTQUEUE_REG_4__2__SCAN_IN,
         P2_INSTQUEUE_REG_4__1__SCAN_IN, P2_INSTQUEUE_REG_4__0__SCAN_IN,
         P2_INSTQUEUE_REG_3__7__SCAN_IN, P2_INSTQUEUE_REG_3__6__SCAN_IN,
         P2_INSTQUEUE_REG_3__5__SCAN_IN, P2_INSTQUEUE_REG_3__4__SCAN_IN,
         P2_INSTQUEUE_REG_3__3__SCAN_IN, P2_INSTQUEUE_REG_3__2__SCAN_IN,
         P2_INSTQUEUE_REG_3__1__SCAN_IN, P2_INSTQUEUE_REG_3__0__SCAN_IN,
         P2_INSTQUEUE_REG_2__7__SCAN_IN, P2_INSTQUEUE_REG_2__6__SCAN_IN,
         P2_INSTQUEUE_REG_2__5__SCAN_IN, P2_INSTQUEUE_REG_2__4__SCAN_IN,
         P2_INSTQUEUE_REG_2__3__SCAN_IN, P2_INSTQUEUE_REG_2__2__SCAN_IN,
         P2_INSTQUEUE_REG_2__1__SCAN_IN, P2_INSTQUEUE_REG_2__0__SCAN_IN,
         P2_INSTQUEUE_REG_1__7__SCAN_IN, P2_INSTQUEUE_REG_1__6__SCAN_IN,
         P2_INSTQUEUE_REG_1__5__SCAN_IN, P2_INSTQUEUE_REG_1__4__SCAN_IN,
         P2_INSTQUEUE_REG_1__3__SCAN_IN, P2_INSTQUEUE_REG_1__2__SCAN_IN,
         P2_INSTQUEUE_REG_1__1__SCAN_IN, P2_INSTQUEUE_REG_1__0__SCAN_IN,
         P2_INSTQUEUE_REG_0__7__SCAN_IN, P2_INSTQUEUE_REG_0__6__SCAN_IN,
         P2_INSTQUEUE_REG_0__5__SCAN_IN, P2_INSTQUEUE_REG_0__4__SCAN_IN,
         P2_INSTQUEUE_REG_0__3__SCAN_IN, P2_INSTQUEUE_REG_0__2__SCAN_IN,
         P2_INSTQUEUE_REG_0__1__SCAN_IN, P2_INSTQUEUE_REG_0__0__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN,
         P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN,
         P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN,
         P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN,
         P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN,
         P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN,
         P2_INSTADDRPOINTER_REG_11__SCAN_IN,
         P2_INSTADDRPOINTER_REG_12__SCAN_IN,
         P2_INSTADDRPOINTER_REG_13__SCAN_IN,
         P2_INSTADDRPOINTER_REG_14__SCAN_IN,
         P2_INSTADDRPOINTER_REG_15__SCAN_IN,
         P2_INSTADDRPOINTER_REG_16__SCAN_IN,
         P2_INSTADDRPOINTER_REG_17__SCAN_IN,
         P2_INSTADDRPOINTER_REG_18__SCAN_IN,
         P2_INSTADDRPOINTER_REG_19__SCAN_IN,
         P2_INSTADDRPOINTER_REG_20__SCAN_IN,
         P2_INSTADDRPOINTER_REG_21__SCAN_IN,
         P2_INSTADDRPOINTER_REG_22__SCAN_IN,
         P2_INSTADDRPOINTER_REG_23__SCAN_IN,
         P2_INSTADDRPOINTER_REG_24__SCAN_IN,
         P2_INSTADDRPOINTER_REG_25__SCAN_IN,
         P2_INSTADDRPOINTER_REG_26__SCAN_IN,
         P2_INSTADDRPOINTER_REG_27__SCAN_IN,
         P2_INSTADDRPOINTER_REG_28__SCAN_IN,
         P2_INSTADDRPOINTER_REG_29__SCAN_IN,
         P2_INSTADDRPOINTER_REG_30__SCAN_IN,
         P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN,
         P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN,
         P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN,
         P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN,
         P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN,
         P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN,
         P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN,
         P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN,
         P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN,
         P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN,
         P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN,
         P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN,
         P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN,
         P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN,
         P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN,
         P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN,
         P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN,
         P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN,
         P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN,
         P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN,
         P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN,
         P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN,
         P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN,
         P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN,
         P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN,
         P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN,
         P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN,
         P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN,
         P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN,
         P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN,
         P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN,
         P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN,
         P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN,
         P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN,
         P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN,
         P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN,
         P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN,
         P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN,
         P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN,
         P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN,
         P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN,
         P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN,
         P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN,
         P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN,
         P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN,
         P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN,
         P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN,
         P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN,
         P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN,
         P2_EAX_REG_14__SCAN_IN, P2_EAX_REG_15__SCAN_IN,
         P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN,
         P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN,
         P2_EAX_REG_20__SCAN_IN, P2_EAX_REG_21__SCAN_IN,
         P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN,
         P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN,
         P2_EAX_REG_26__SCAN_IN, P2_EAX_REG_27__SCAN_IN,
         P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN,
         P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN,
         P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN,
         P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN,
         P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN,
         P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN,
         P2_EBX_REG_12__SCAN_IN, P2_EBX_REG_13__SCAN_IN,
         P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN,
         P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN,
         P2_EBX_REG_18__SCAN_IN, P2_EBX_REG_19__SCAN_IN,
         P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN,
         P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN,
         P2_EBX_REG_24__SCAN_IN, P2_EBX_REG_25__SCAN_IN,
         P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN,
         P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN,
         P2_EBX_REG_30__SCAN_IN, P2_EBX_REG_31__SCAN_IN,
         P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN,
         P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN,
         P2_REIP_REG_4__SCAN_IN, P2_REIP_REG_5__SCAN_IN,
         P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN,
         P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN,
         P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN,
         P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN,
         P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN,
         P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN,
         P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN,
         P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN,
         P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN,
         P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN,
         P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN,
         P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN,
         P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN,
         P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN,
         P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN,
         P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN,
         P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN,
         P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN,
         P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN,
         P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN,
         P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN,
         P1_BE_N_REG_0__SCAN_IN, P1_ADDRESS_REG_29__SCAN_IN,
         P1_ADDRESS_REG_28__SCAN_IN, P1_ADDRESS_REG_27__SCAN_IN,
         P1_ADDRESS_REG_26__SCAN_IN, P1_ADDRESS_REG_25__SCAN_IN,
         P1_ADDRESS_REG_24__SCAN_IN, P1_ADDRESS_REG_23__SCAN_IN,
         P1_ADDRESS_REG_22__SCAN_IN, P1_ADDRESS_REG_21__SCAN_IN,
         P1_ADDRESS_REG_20__SCAN_IN, P1_ADDRESS_REG_19__SCAN_IN,
         P1_ADDRESS_REG_18__SCAN_IN, P1_ADDRESS_REG_17__SCAN_IN,
         P1_ADDRESS_REG_16__SCAN_IN, P1_ADDRESS_REG_15__SCAN_IN,
         P1_ADDRESS_REG_14__SCAN_IN, P1_ADDRESS_REG_13__SCAN_IN,
         P1_ADDRESS_REG_12__SCAN_IN, P1_ADDRESS_REG_11__SCAN_IN,
         P1_ADDRESS_REG_10__SCAN_IN, P1_ADDRESS_REG_9__SCAN_IN,
         P1_ADDRESS_REG_8__SCAN_IN, P1_ADDRESS_REG_7__SCAN_IN,
         P1_ADDRESS_REG_6__SCAN_IN, P1_ADDRESS_REG_5__SCAN_IN,
         P1_ADDRESS_REG_4__SCAN_IN, P1_ADDRESS_REG_3__SCAN_IN,
         P1_ADDRESS_REG_2__SCAN_IN, P1_ADDRESS_REG_1__SCAN_IN,
         P1_ADDRESS_REG_0__SCAN_IN, P1_STATE_REG_2__SCAN_IN,
         P1_STATE_REG_1__SCAN_IN, P1_STATE_REG_0__SCAN_IN,
         P1_DATAWIDTH_REG_0__SCAN_IN, P1_DATAWIDTH_REG_1__SCAN_IN,
         P1_DATAWIDTH_REG_2__SCAN_IN, P1_DATAWIDTH_REG_3__SCAN_IN,
         P1_DATAWIDTH_REG_4__SCAN_IN, P1_DATAWIDTH_REG_5__SCAN_IN,
         P1_DATAWIDTH_REG_6__SCAN_IN, P1_DATAWIDTH_REG_7__SCAN_IN,
         P1_DATAWIDTH_REG_8__SCAN_IN, P1_DATAWIDTH_REG_9__SCAN_IN,
         P1_DATAWIDTH_REG_10__SCAN_IN, P1_DATAWIDTH_REG_11__SCAN_IN,
         P1_DATAWIDTH_REG_12__SCAN_IN, P1_DATAWIDTH_REG_13__SCAN_IN,
         P1_DATAWIDTH_REG_14__SCAN_IN, P1_DATAWIDTH_REG_15__SCAN_IN,
         P1_DATAWIDTH_REG_16__SCAN_IN, P1_DATAWIDTH_REG_17__SCAN_IN,
         P1_DATAWIDTH_REG_18__SCAN_IN, P1_DATAWIDTH_REG_19__SCAN_IN,
         P1_DATAWIDTH_REG_20__SCAN_IN, P1_DATAWIDTH_REG_21__SCAN_IN,
         P1_DATAWIDTH_REG_22__SCAN_IN, P1_DATAWIDTH_REG_23__SCAN_IN,
         P1_DATAWIDTH_REG_24__SCAN_IN, P1_DATAWIDTH_REG_25__SCAN_IN,
         P1_DATAWIDTH_REG_26__SCAN_IN, P1_DATAWIDTH_REG_27__SCAN_IN,
         P1_DATAWIDTH_REG_28__SCAN_IN, P1_DATAWIDTH_REG_29__SCAN_IN,
         P1_DATAWIDTH_REG_30__SCAN_IN, P1_DATAWIDTH_REG_31__SCAN_IN,
         P1_STATE2_REG_3__SCAN_IN, P1_STATE2_REG_2__SCAN_IN,
         P1_STATE2_REG_1__SCAN_IN, P1_STATE2_REG_0__SCAN_IN,
         P1_INSTQUEUE_REG_15__7__SCAN_IN, P1_INSTQUEUE_REG_15__6__SCAN_IN,
         P1_INSTQUEUE_REG_15__5__SCAN_IN, P1_INSTQUEUE_REG_15__4__SCAN_IN,
         P1_INSTQUEUE_REG_15__3__SCAN_IN, P1_INSTQUEUE_REG_15__2__SCAN_IN,
         P1_INSTQUEUE_REG_15__1__SCAN_IN, P1_INSTQUEUE_REG_15__0__SCAN_IN,
         P1_INSTQUEUE_REG_14__7__SCAN_IN, P1_INSTQUEUE_REG_14__6__SCAN_IN,
         P1_INSTQUEUE_REG_14__5__SCAN_IN, P1_INSTQUEUE_REG_14__4__SCAN_IN,
         P1_INSTQUEUE_REG_14__3__SCAN_IN, P1_INSTQUEUE_REG_14__2__SCAN_IN,
         P1_INSTQUEUE_REG_14__1__SCAN_IN, P1_INSTQUEUE_REG_14__0__SCAN_IN,
         P1_INSTQUEUE_REG_13__7__SCAN_IN, P1_INSTQUEUE_REG_13__6__SCAN_IN,
         P1_INSTQUEUE_REG_13__5__SCAN_IN, P1_INSTQUEUE_REG_13__4__SCAN_IN,
         P1_INSTQUEUE_REG_13__3__SCAN_IN, P1_INSTQUEUE_REG_13__2__SCAN_IN,
         P1_INSTQUEUE_REG_13__1__SCAN_IN, P1_INSTQUEUE_REG_13__0__SCAN_IN,
         P1_INSTQUEUE_REG_12__7__SCAN_IN, P1_INSTQUEUE_REG_12__6__SCAN_IN,
         P1_INSTQUEUE_REG_12__5__SCAN_IN, P1_INSTQUEUE_REG_12__4__SCAN_IN,
         P1_INSTQUEUE_REG_12__3__SCAN_IN, P1_INSTQUEUE_REG_12__2__SCAN_IN,
         P1_INSTQUEUE_REG_12__1__SCAN_IN, P1_INSTQUEUE_REG_12__0__SCAN_IN,
         P1_INSTQUEUE_REG_11__7__SCAN_IN, P1_INSTQUEUE_REG_11__6__SCAN_IN,
         P1_INSTQUEUE_REG_11__5__SCAN_IN, P1_INSTQUEUE_REG_11__4__SCAN_IN,
         P1_INSTQUEUE_REG_11__3__SCAN_IN, P1_INSTQUEUE_REG_11__2__SCAN_IN,
         P1_INSTQUEUE_REG_11__1__SCAN_IN, P1_INSTQUEUE_REG_11__0__SCAN_IN,
         P1_INSTQUEUE_REG_10__7__SCAN_IN, P1_INSTQUEUE_REG_10__6__SCAN_IN,
         P1_INSTQUEUE_REG_10__5__SCAN_IN, P1_INSTQUEUE_REG_10__4__SCAN_IN,
         P1_INSTQUEUE_REG_10__3__SCAN_IN, P1_INSTQUEUE_REG_10__2__SCAN_IN,
         P1_INSTQUEUE_REG_10__1__SCAN_IN, P1_INSTQUEUE_REG_10__0__SCAN_IN,
         P1_INSTQUEUE_REG_9__7__SCAN_IN, P1_INSTQUEUE_REG_9__6__SCAN_IN,
         P1_INSTQUEUE_REG_9__5__SCAN_IN, P1_INSTQUEUE_REG_9__4__SCAN_IN,
         P1_INSTQUEUE_REG_9__3__SCAN_IN, P1_INSTQUEUE_REG_9__2__SCAN_IN,
         P1_INSTQUEUE_REG_9__1__SCAN_IN, P1_INSTQUEUE_REG_9__0__SCAN_IN,
         P1_INSTQUEUE_REG_8__7__SCAN_IN, P1_INSTQUEUE_REG_8__6__SCAN_IN,
         P1_INSTQUEUE_REG_8__5__SCAN_IN, P1_INSTQUEUE_REG_8__4__SCAN_IN,
         P1_INSTQUEUE_REG_8__3__SCAN_IN, P1_INSTQUEUE_REG_8__2__SCAN_IN,
         P1_INSTQUEUE_REG_8__1__SCAN_IN, P1_INSTQUEUE_REG_8__0__SCAN_IN,
         P1_INSTQUEUE_REG_7__7__SCAN_IN, P1_INSTQUEUE_REG_7__6__SCAN_IN,
         P1_INSTQUEUE_REG_7__5__SCAN_IN, P1_INSTQUEUE_REG_7__4__SCAN_IN,
         P1_INSTQUEUE_REG_7__3__SCAN_IN, P1_INSTQUEUE_REG_7__2__SCAN_IN,
         P1_INSTQUEUE_REG_7__1__SCAN_IN, P1_INSTQUEUE_REG_7__0__SCAN_IN,
         P1_INSTQUEUE_REG_6__7__SCAN_IN, P1_INSTQUEUE_REG_6__6__SCAN_IN,
         P1_INSTQUEUE_REG_6__5__SCAN_IN, P1_INSTQUEUE_REG_6__4__SCAN_IN,
         P1_INSTQUEUE_REG_6__3__SCAN_IN, P1_INSTQUEUE_REG_6__2__SCAN_IN,
         P1_INSTQUEUE_REG_6__1__SCAN_IN, P1_INSTQUEUE_REG_6__0__SCAN_IN,
         P1_INSTQUEUE_REG_5__7__SCAN_IN, P1_INSTQUEUE_REG_5__6__SCAN_IN,
         P1_INSTQUEUE_REG_5__5__SCAN_IN, P1_INSTQUEUE_REG_5__4__SCAN_IN,
         P1_INSTQUEUE_REG_5__3__SCAN_IN, P1_INSTQUEUE_REG_5__2__SCAN_IN,
         P1_INSTQUEUE_REG_5__1__SCAN_IN, P1_INSTQUEUE_REG_5__0__SCAN_IN,
         P1_INSTQUEUE_REG_4__7__SCAN_IN, P1_INSTQUEUE_REG_4__6__SCAN_IN,
         P1_INSTQUEUE_REG_4__5__SCAN_IN, P1_INSTQUEUE_REG_4__4__SCAN_IN,
         P1_INSTQUEUE_REG_4__3__SCAN_IN, P1_INSTQUEUE_REG_4__2__SCAN_IN,
         P1_INSTQUEUE_REG_4__1__SCAN_IN, keyinput0, keyinput1, keyinput2,
         keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, keyinput8,
         keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
         keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
         keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
         keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
         keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
         keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
         keyinput90, keyinput91, keyinput92, keyinput93, keyinput94,
         keyinput95, keyinput96, keyinput97, keyinput98, keyinput99,
         keyinput100, keyinput101, keyinput102, keyinput103, keyinput104,
         keyinput105, keyinput106, keyinput107, keyinput108, keyinput109,
         keyinput110, keyinput111, keyinput112, keyinput113, keyinput114,
         keyinput115, keyinput116, keyinput117, keyinput118, keyinput119,
         keyinput120, keyinput121, keyinput122, keyinput123, keyinput124,
         keyinput125, keyinput126, keyinput127;
  output U355, U356, U357, U358, U359, U360, U361, U362, U363, U364, U366,
         U367, U368, U369, U370, U371, U372, U373, U374, U375, U347, U348,
         U349, U350, U351, U352, U353, U354, U365, U376, U247, U246, U245,
         U244, U243, U242, U241, U240, U239, U238, U237, U236, U235, U234,
         U233, U232, U231, U230, U229, U228, U227, U226, U225, U224, U223,
         U222, U221, U220, U219, U218, U217, U216, U251, U252, U253, U254,
         U255, U256, U257, U258, U259, U260, U261, U262, U263, U264, U265,
         U266, U267, U268, U269, U270, U271, U272, U273, U274, U275, U276,
         U277, U278, U279, U280, U281, U282, U212, U215, U213, U214, P3_U3274,
         P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, P3_U3059, P3_U3058,
         P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, P3_U3052, P3_U3051,
         P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, P3_U3045, P3_U3044,
         P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, P3_U3038, P3_U3037,
         P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, P3_U3031, P3_U3030,
         P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, P3_U3026, P3_U3025,
         P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, P3_U3019, P3_U3018,
         P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, P3_U3012, P3_U3011,
         P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, P3_U3005, P3_U3004,
         P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, P3_U3282, P3_U2998,
         P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, P3_U2992, P3_U2991,
         P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, P3_U2985, P3_U2984,
         P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, P3_U2978, P3_U2977,
         P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, P3_U2971, P3_U2970,
         P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, P3_U2964, P3_U2963,
         P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, P3_U2957, P3_U2956,
         P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, P3_U2950, P3_U2949,
         P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, P3_U2943, P3_U2942,
         P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, P3_U2936, P3_U2935,
         P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, P3_U2929, P3_U2928,
         P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, P3_U2922, P3_U2921,
         P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, P3_U2915, P3_U2914,
         P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, P3_U2908, P3_U2907,
         P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, P3_U2901, P3_U2900,
         P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, P3_U2894, P3_U2893,
         P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, P3_U2887, P3_U2886,
         P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, P3_U2880, P3_U2879,
         P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, P3_U2873, P3_U2872,
         P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, P3_U3285, P3_U3288,
         P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, P3_U2864, P3_U2863,
         P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, P3_U2857, P3_U2856,
         P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, P3_U2850, P3_U2849,
         P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, P3_U2843, P3_U2842,
         P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, P3_U2836, P3_U2835,
         P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, P3_U2829, P3_U2828,
         P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, P3_U2822, P3_U2821,
         P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, P3_U2815, P3_U2814,
         P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, P3_U2808, P3_U2807,
         P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, P3_U2801, P3_U2800,
         P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, P3_U2794, P3_U2793,
         P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, P3_U2787, P3_U2786,
         P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, P3_U2780, P3_U2779,
         P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, P3_U2773, P3_U2772,
         P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, P3_U2766, P3_U2765,
         P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, P3_U2759, P3_U2758,
         P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, P3_U2752, P3_U2751,
         P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, P3_U2745, P3_U2744,
         P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, P3_U2738, P3_U2737,
         P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, P3_U2731, P3_U2730,
         P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, P3_U2724, P3_U2723,
         P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, P3_U2717, P3_U2716,
         P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, P3_U2710, P3_U2709,
         P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, P3_U2703, P3_U2702,
         P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, P3_U2696, P3_U2695,
         P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, P3_U2689, P3_U2688,
         P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, P3_U2682, P3_U2681,
         P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, P3_U2675, P3_U2674,
         P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, P3_U2668, P3_U2667,
         P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, P3_U2661, P3_U2660,
         P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, P3_U2654, P3_U2653,
         P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, P3_U2647, P3_U2646,
         P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, P3_U2640, P3_U2639,
         P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, P3_U3295, P3_U2636,
         P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, P3_U3298, P3_U3299,
         P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, P2_U3240, P2_U3239,
         P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232,
         P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225,
         P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218,
         P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, P2_U3207, P2_U3206,
         P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199,
         P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192,
         P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185,
         P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, P2_U3179, P2_U3593,
         P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172,
         P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165,
         P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158,
         P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3152, P2_U3151,
         P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, P2_U3145, P2_U3144,
         P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, P2_U3138, P2_U3137,
         P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, P2_U3131, P2_U3130,
         P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, P2_U3124, P2_U3123,
         P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, P2_U3117, P2_U3116,
         P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, P2_U3110, P2_U3109,
         P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, P2_U3103, P2_U3102,
         P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, P2_U3096, P2_U3095,
         P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, P2_U3089, P2_U3088,
         P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, P2_U3082, P2_U3081,
         P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, P2_U3075, P2_U3074,
         P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, P2_U3068, P2_U3067,
         P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, P2_U3061, P2_U3060,
         P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, P2_U3054, P2_U3053,
         P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, P2_U3595, P2_U3596,
         P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, P2_U3603, P2_U3604,
         P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, P2_U3042, P2_U3041,
         P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, P2_U3035, P2_U3034,
         P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, P2_U3028, P2_U3027,
         P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, P2_U3021, P2_U3020,
         P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, P2_U3014, P2_U3013,
         P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, P2_U3007, P2_U3006,
         P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, P2_U3000, P2_U2999,
         P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, P2_U2993, P2_U2992,
         P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, P2_U2986, P2_U2985,
         P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, P2_U2979, P2_U2978,
         P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, P2_U2972, P2_U2971,
         P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, P2_U2965, P2_U2964,
         P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, P2_U2958, P2_U2957,
         P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, P2_U2951, P2_U2950,
         P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, P2_U2944, P2_U2943,
         P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, P2_U2937, P2_U2936,
         P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, P2_U2930, P2_U2929,
         P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, P2_U2923, P2_U2922,
         P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, P2_U2916, P2_U2915,
         P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, P2_U2909, P2_U2908,
         P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, P2_U2902, P2_U2901,
         P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, P2_U2895, P2_U2894,
         P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, P2_U2888, P2_U2887,
         P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, P2_U2881, P2_U2880,
         P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, P2_U2874, P2_U2873,
         P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, P2_U2867, P2_U2866,
         P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, P2_U2860, P2_U2859,
         P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, P2_U2853, P2_U2852,
         P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, P2_U2846, P2_U2845,
         P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, P2_U2839, P2_U2838,
         P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, P2_U2832, P2_U2831,
         P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, P2_U2825, P2_U2824,
         P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, P2_U2819, P2_U3609,
         P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, P2_U2815, P2_U3612,
         P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211,
         P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, P1_U3205, P1_U3204,
         P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, P1_U3198, P1_U3197,
         P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, P1_U3193, P1_U3192,
         P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, P1_U3186, P1_U3185,
         P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, P1_U3179, P1_U3178,
         P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, P1_U3172, P1_U3171,
         P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, P1_U3165, P1_U3164,
         P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, P1_U3159, P1_U3158,
         P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, P1_U3152, P1_U3151,
         P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, P1_U3145, P1_U3144,
         P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, P1_U3138, P1_U3137,
         P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, P1_U3131, P1_U3130,
         P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, P1_U3124, P1_U3123,
         P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, P1_U3117, P1_U3116,
         P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, P1_U3110, P1_U3109,
         P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, P1_U3103, P1_U3102,
         P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, P1_U3096, P1_U3095,
         P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, P1_U3089, P1_U3088,
         P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, P1_U3082, P1_U3081,
         P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, P1_U3075, P1_U3074,
         P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, P1_U3068, P1_U3067,
         P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, P1_U3061, P1_U3060,
         P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, P1_U3054, P1_U3053,
         P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, P1_U3047, P1_U3046,
         P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, P1_U3040, P1_U3039,
         P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, P1_U3033, P1_U3468,
         P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, P1_U3475, P1_U3476,
         P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, P1_U3028, P1_U3027,
         P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, P1_U3021, P1_U3020,
         P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, P1_U3014, P1_U3013,
         P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, P1_U3007, P1_U3006,
         P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, P1_U3000, P1_U2999,
         P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, P1_U2993, P1_U2992,
         P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, P1_U2986, P1_U2985,
         P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, P1_U2979, P1_U2978,
         P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, P1_U2972, P1_U2971,
         P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, P1_U2965, P1_U2964,
         P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, P1_U2958, P1_U2957,
         P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, P1_U2951, P1_U2950,
         P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, P1_U2944, P1_U2943,
         P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, P1_U2937, P1_U2936,
         P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, P1_U2930, P1_U2929,
         P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, P1_U2923, P1_U2922,
         P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, P1_U2916, P1_U2915,
         P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, P1_U2909, P1_U2908,
         P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, P1_U2902, P1_U2901,
         P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, P1_U2895, P1_U2894,
         P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, P1_U2888, P1_U2887,
         P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, P1_U2881, P1_U2880,
         P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, P1_U2874, P1_U2873,
         P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, P1_U2867, P1_U2866,
         P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, P1_U2860, P1_U2859,
         P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, P1_U2853, P1_U2852,
         P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, P1_U2846, P1_U2845,
         P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, P1_U2839, P1_U2838,
         P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, P1_U2832, P1_U2831,
         P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, P1_U2825, P1_U2824,
         P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, P1_U2818, P1_U2817,
         P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, P1_U2811, P1_U2810,
         P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, P1_U3483, P1_U2806,
         P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, P1_U2803, P1_U2802,
         P1_U3487, P1_U2801;
  wire   n9602, n9603, n9604, n9605, n9606, n9607, n9609, n9610, n9611, n9612,
         n9613, n9614, n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623,
         n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9633, n9634,
         n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644,
         n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654,
         n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664,
         n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674,
         n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684,
         n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694,
         n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704,
         n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714,
         n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724,
         n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734,
         n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744,
         n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754,
         n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764,
         n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774,
         n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784,
         n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794,
         n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804,
         n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814,
         n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824,
         n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834,
         n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844,
         n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854,
         n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864,
         n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874,
         n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884,
         n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894,
         n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904,
         n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914,
         n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924,
         n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934,
         n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944,
         n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954,
         n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964,
         n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974,
         n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984,
         n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994,
         n9995, n9996, n9997, n9998, n9999, n10000, n10001, n10002, n10003,
         n10004, n10005, n10006, n10007, n10008, n10009, n10010, n10011,
         n10012, n10013, n10014, n10015, n10016, n10017, n10018, n10019,
         n10020, n10021, n10022, n10023, n10024, n10025, n10026, n10027,
         n10028, n10029, n10030, n10031, n10032, n10033, n10034, n10035,
         n10036, n10037, n10038, n10039, n10040, n10041, n10042, n10043,
         n10044, n10045, n10046, n10047, n10048, n10049, n10050, n10051,
         n10052, n10053, n10054, n10055, n10056, n10057, n10058, n10059,
         n10060, n10061, n10062, n10063, n10064, n10065, n10066, n10067,
         n10068, n10069, n10070, n10071, n10072, n10073, n10074, n10075,
         n10076, n10077, n10078, n10079, n10080, n10081, n10082, n10083,
         n10084, n10085, n10086, n10087, n10088, n10089, n10090, n10091,
         n10092, n10093, n10094, n10095, n10096, n10097, n10098, n10099,
         n10100, n10101, n10102, n10103, n10104, n10105, n10106, n10107,
         n10108, n10109, n10110, n10111, n10112, n10113, n10114, n10115,
         n10116, n10117, n10118, n10119, n10120, n10121, n10122, n10123,
         n10124, n10125, n10126, n10127, n10128, n10129, n10130, n10131,
         n10132, n10133, n10134, n10135, n10136, n10137, n10138, n10139,
         n10140, n10141, n10142, n10143, n10144, n10145, n10146, n10147,
         n10148, n10149, n10150, n10151, n10152, n10153, n10154, n10155,
         n10156, n10157, n10158, n10159, n10160, n10161, n10162, n10163,
         n10164, n10165, n10166, n10167, n10168, n10169, n10170, n10171,
         n10172, n10173, n10174, n10175, n10176, n10177, n10178, n10179,
         n10180, n10181, n10182, n10183, n10184, n10185, n10186, n10187,
         n10188, n10189, n10190, n10191, n10192, n10193, n10194, n10195,
         n10196, n10197, n10198, n10199, n10200, n10201, n10202, n10203,
         n10204, n10205, n10206, n10207, n10208, n10209, n10210, n10211,
         n10212, n10213, n10214, n10215, n10216, n10217, n10218, n10219,
         n10220, n10221, n10222, n10223, n10224, n10225, n10226, n10227,
         n10228, n10229, n10230, n10231, n10232, n10233, n10234, n10235,
         n10236, n10237, n10238, n10239, n10240, n10241, n10242, n10243,
         n10244, n10245, n10246, n10247, n10248, n10249, n10250, n10251,
         n10252, n10253, n10254, n10255, n10256, n10257, n10258, n10259,
         n10260, n10261, n10262, n10263, n10264, n10265, n10266, n10267,
         n10268, n10269, n10270, n10271, n10272, n10273, n10274, n10275,
         n10276, n10277, n10278, n10279, n10280, n10281, n10282, n10283,
         n10284, n10285, n10286, n10287, n10288, n10289, n10290, n10291,
         n10292, n10293, n10294, n10295, n10296, n10297, n10298, n10299,
         n10300, n10301, n10302, n10303, n10304, n10305, n10306, n10307,
         n10308, n10309, n10310, n10311, n10312, n10313, n10314, n10315,
         n10316, n10317, n10318, n10319, n10320, n10321, n10322, n10323,
         n10324, n10325, n10326, n10327, n10328, n10329, n10330, n10331,
         n10332, n10333, n10334, n10335, n10336, n10337, n10338, n10339,
         n10340, n10341, n10342, n10343, n10344, n10345, n10346, n10347,
         n10348, n10349, n10350, n10351, n10352, n10353, n10354, n10355,
         n10356, n10357, n10358, n10359, n10360, n10361, n10362, n10363,
         n10364, n10365, n10366, n10367, n10368, n10369, n10370, n10371,
         n10372, n10373, n10374, n10375, n10376, n10377, n10378, n10379,
         n10380, n10381, n10382, n10383, n10384, n10385, n10386, n10387,
         n10388, n10389, n10390, n10391, n10392, n10393, n10394, n10395,
         n10396, n10397, n10398, n10399, n10400, n10401, n10402, n10403,
         n10404, n10405, n10406, n10407, n10408, n10409, n10410, n10411,
         n10412, n10413, n10414, n10415, n10416, n10417, n10418, n10419,
         n10420, n10421, n10422, n10423, n10424, n10425, n10426, n10427,
         n10428, n10429, n10430, n10431, n10432, n10433, n10434, n10435,
         n10436, n10437, n10438, n10439, n10440, n10441, n10442, n10443,
         n10444, n10445, n10446, n10447, n10448, n10449, n10450, n10451,
         n10452, n10453, n10454, n10455, n10456, n10457, n10458, n10459,
         n10460, n10461, n10462, n10463, n10464, n10465, n10466, n10467,
         n10468, n10469, n10470, n10471, n10472, n10473, n10474, n10475,
         n10476, n10477, n10478, n10479, n10480, n10481, n10482, n10483,
         n10484, n10485, n10486, n10487, n10488, n10489, n10490, n10491,
         n10492, n10493, n10494, n10495, n10496, n10497, n10498, n10499,
         n10500, n10501, n10502, n10503, n10504, n10505, n10506, n10507,
         n10508, n10509, n10510, n10511, n10512, n10513, n10514, n10515,
         n10516, n10517, n10518, n10519, n10520, n10521, n10522, n10523,
         n10524, n10525, n10526, n10527, n10528, n10529, n10530, n10531,
         n10532, n10533, n10534, n10535, n10536, n10537, n10538, n10539,
         n10540, n10541, n10542, n10543, n10544, n10545, n10546, n10547,
         n10548, n10549, n10550, n10551, n10552, n10553, n10554, n10555,
         n10556, n10557, n10558, n10559, n10560, n10561, n10562, n10563,
         n10564, n10565, n10566, n10567, n10568, n10569, n10570, n10571,
         n10572, n10573, n10574, n10575, n10576, n10577, n10578, n10579,
         n10580, n10581, n10582, n10583, n10584, n10585, n10586, n10587,
         n10588, n10589, n10590, n10591, n10592, n10593, n10594, n10595,
         n10596, n10597, n10598, n10599, n10600, n10601, n10602, n10603,
         n10604, n10605, n10606, n10607, n10608, n10609, n10610, n10611,
         n10612, n10613, n10614, n10615, n10616, n10617, n10618, n10619,
         n10620, n10621, n10622, n10623, n10624, n10625, n10626, n10627,
         n10628, n10629, n10630, n10631, n10632, n10633, n10634, n10635,
         n10636, n10637, n10638, n10639, n10640, n10641, n10642, n10643,
         n10644, n10645, n10646, n10647, n10648, n10649, n10650, n10651,
         n10652, n10653, n10654, n10655, n10656, n10657, n10658, n10659,
         n10660, n10661, n10662, n10663, n10664, n10665, n10666, n10667,
         n10668, n10669, n10670, n10671, n10672, n10673, n10674, n10675,
         n10676, n10677, n10678, n10679, n10680, n10681, n10682, n10683,
         n10684, n10685, n10686, n10687, n10688, n10689, n10690, n10691,
         n10692, n10693, n10694, n10695, n10696, n10697, n10698, n10699,
         n10700, n10701, n10702, n10703, n10704, n10705, n10706, n10707,
         n10708, n10709, n10710, n10711, n10712, n10713, n10714, n10715,
         n10716, n10717, n10718, n10719, n10720, n10721, n10722, n10723,
         n10724, n10725, n10726, n10727, n10728, n10729, n10730, n10731,
         n10732, n10733, n10734, n10735, n10736, n10737, n10738, n10739,
         n10740, n10741, n10742, n10743, n10744, n10745, n10746, n10747,
         n10748, n10749, n10750, n10751, n10752, n10753, n10754, n10755,
         n10756, n10757, n10758, n10759, n10760, n10761, n10762, n10763,
         n10764, n10765, n10766, n10767, n10768, n10769, n10770, n10771,
         n10772, n10773, n10774, n10775, n10776, n10777, n10778, n10779,
         n10780, n10781, n10782, n10783, n10784, n10785, n10786, n10787,
         n10788, n10789, n10790, n10791, n10792, n10793, n10794, n10795,
         n10796, n10797, n10798, n10799, n10800, n10801, n10802, n10803,
         n10804, n10805, n10806, n10807, n10808, n10809, n10810, n10811,
         n10812, n10813, n10814, n10815, n10816, n10817, n10818, n10819,
         n10820, n10821, n10822, n10823, n10824, n10825, n10826, n10827,
         n10828, n10829, n10830, n10831, n10832, n10833, n10834, n10835,
         n10836, n10837, n10838, n10839, n10840, n10841, n10842, n10843,
         n10844, n10845, n10846, n10847, n10848, n10849, n10850, n10851,
         n10852, n10853, n10854, n10855, n10856, n10857, n10858, n10859,
         n10860, n10861, n10862, n10863, n10864, n10865, n10866, n10867,
         n10868, n10869, n10870, n10871, n10872, n10873, n10874, n10875,
         n10876, n10877, n10878, n10879, n10880, n10881, n10882, n10883,
         n10884, n10885, n10886, n10887, n10888, n10889, n10890, n10891,
         n10892, n10893, n10894, n10895, n10896, n10897, n10898, n10899,
         n10900, n10901, n10902, n10903, n10904, n10905, n10906, n10907,
         n10908, n10909, n10910, n10911, n10912, n10913, n10914, n10915,
         n10916, n10917, n10918, n10919, n10920, n10921, n10922, n10923,
         n10924, n10925, n10926, n10927, n10928, n10929, n10930, n10931,
         n10932, n10933, n10934, n10935, n10936, n10937, n10938, n10939,
         n10940, n10941, n10942, n10943, n10944, n10945, n10946, n10947,
         n10948, n10949, n10950, n10951, n10952, n10953, n10954, n10955,
         n10956, n10957, n10958, n10959, n10960, n10961, n10962, n10963,
         n10964, n10965, n10966, n10967, n10968, n10969, n10970, n10971,
         n10972, n10973, n10974, n10975, n10976, n10977, n10978, n10979,
         n10980, n10981, n10982, n10983, n10984, n10985, n10986, n10987,
         n10988, n10989, n10990, n10991, n10992, n10993, n10994, n10995,
         n10996, n10997, n10998, n10999, n11000, n11001, n11002, n11003,
         n11004, n11005, n11006, n11007, n11008, n11009, n11010, n11011,
         n11012, n11013, n11014, n11015, n11016, n11017, n11018, n11019,
         n11020, n11021, n11022, n11023, n11024, n11025, n11026, n11027,
         n11028, n11029, n11030, n11031, n11032, n11033, n11034, n11035,
         n11036, n11037, n11038, n11039, n11040, n11041, n11042, n11044,
         n11045, n11046, n11047, n11048, n11049, n11050, n11051, n11052,
         n11053, n11054, n11055, n11056, n11057, n11058, n11059, n11060,
         n11061, n11062, n11063, n11064, n11065, n11066, n11067, n11068,
         n11069, n11070, n11071, n11072, n11073, n11074, n11075, n11076,
         n11077, n11078, n11079, n11080, n11081, n11082, n11083, n11084,
         n11085, n11086, n11087, n11088, n11089, n11090, n11091, n11092,
         n11093, n11094, n11095, n11096, n11097, n11098, n11099, n11100,
         n11101, n11102, n11103, n11104, n11105, n11106, n11107, n11108,
         n11109, n11110, n11111, n11112, n11113, n11114, n11115, n11116,
         n11117, n11118, n11119, n11120, n11121, n11122, n11123, n11124,
         n11125, n11126, n11127, n11128, n11129, n11130, n11131, n11132,
         n11133, n11134, n11135, n11136, n11137, n11138, n11139, n11140,
         n11141, n11142, n11143, n11144, n11145, n11146, n11147, n11148,
         n11149, n11150, n11151, n11152, n11153, n11154, n11155, n11156,
         n11157, n11158, n11159, n11160, n11161, n11162, n11163, n11164,
         n11165, n11166, n11167, n11168, n11169, n11170, n11171, n11172,
         n11173, n11174, n11175, n11176, n11177, n11178, n11179, n11180,
         n11181, n11182, n11183, n11184, n11185, n11186, n11187, n11188,
         n11189, n11190, n11191, n11192, n11193, n11194, n11195, n11196,
         n11197, n11198, n11199, n11200, n11201, n11202, n11203, n11204,
         n11205, n11206, n11207, n11208, n11209, n11210, n11211, n11212,
         n11213, n11214, n11215, n11216, n11217, n11218, n11219, n11220,
         n11221, n11222, n11223, n11224, n11225, n11226, n11227, n11228,
         n11229, n11230, n11231, n11232, n11233, n11234, n11235, n11236,
         n11237, n11238, n11239, n11240, n11241, n11242, n11243, n11244,
         n11245, n11246, n11247, n11248, n11249, n11250, n11251, n11252,
         n11253, n11254, n11255, n11256, n11257, n11258, n11259, n11260,
         n11261, n11262, n11263, n11264, n11265, n11266, n11267, n11268,
         n11269, n11270, n11271, n11272, n11273, n11274, n11275, n11276,
         n11277, n11278, n11279, n11280, n11281, n11282, n11283, n11284,
         n11285, n11286, n11287, n11288, n11289, n11290, n11291, n11292,
         n11293, n11294, n11295, n11296, n11297, n11298, n11299, n11300,
         n11301, n11302, n11303, n11304, n11305, n11306, n11307, n11308,
         n11309, n11310, n11311, n11312, n11313, n11314, n11315, n11316,
         n11317, n11318, n11319, n11320, n11321, n11322, n11323, n11324,
         n11325, n11326, n11327, n11328, n11329, n11330, n11331, n11332,
         n11333, n11334, n11335, n11336, n11337, n11338, n11339, n11340,
         n11341, n11342, n11343, n11344, n11345, n11346, n11347, n11348,
         n11349, n11350, n11351, n11352, n11353, n11354, n11355, n11356,
         n11357, n11358, n11359, n11360, n11361, n11362, n11363, n11364,
         n11365, n11366, n11367, n11368, n11369, n11370, n11371, n11372,
         n11373, n11374, n11375, n11376, n11377, n11378, n11379, n11380,
         n11381, n11382, n11383, n11384, n11385, n11386, n11387, n11388,
         n11389, n11390, n11391, n11392, n11393, n11394, n11395, n11396,
         n11397, n11398, n11399, n11400, n11401, n11402, n11403, n11404,
         n11405, n11406, n11407, n11408, n11409, n11410, n11411, n11412,
         n11413, n11414, n11415, n11416, n11417, n11418, n11419, n11420,
         n11421, n11422, n11423, n11424, n11425, n11426, n11427, n11428,
         n11429, n11430, n11431, n11432, n11433, n11434, n11435, n11436,
         n11437, n11438, n11439, n11440, n11441, n11442, n11443, n11444,
         n11445, n11446, n11447, n11448, n11449, n11450, n11451, n11452,
         n11453, n11454, n11455, n11456, n11457, n11458, n11459, n11460,
         n11461, n11462, n11463, n11464, n11465, n11466, n11467, n11468,
         n11469, n11470, n11471, n11472, n11473, n11474, n11475, n11476,
         n11477, n11478, n11479, n11480, n11481, n11482, n11483, n11484,
         n11485, n11486, n11487, n11488, n11489, n11490, n11491, n11492,
         n11493, n11494, n11495, n11496, n11497, n11498, n11499, n11500,
         n11501, n11502, n11503, n11504, n11505, n11506, n11507, n11508,
         n11509, n11510, n11511, n11512, n11513, n11514, n11515, n11516,
         n11517, n11518, n11519, n11520, n11521, n11522, n11523, n11524,
         n11525, n11526, n11527, n11528, n11529, n11530, n11531, n11532,
         n11533, n11534, n11535, n11536, n11537, n11538, n11539, n11540,
         n11541, n11542, n11543, n11544, n11545, n11546, n11547, n11548,
         n11549, n11550, n11551, n11552, n11553, n11554, n11555, n11556,
         n11557, n11558, n11559, n11560, n11561, n11562, n11563, n11564,
         n11565, n11566, n11567, n11568, n11569, n11570, n11571, n11572,
         n11573, n11574, n11575, n11576, n11577, n11578, n11579, n11580,
         n11581, n11582, n11583, n11584, n11585, n11586, n11587, n11588,
         n11589, n11590, n11591, n11592, n11593, n11594, n11595, n11596,
         n11597, n11598, n11599, n11600, n11601, n11602, n11603, n11604,
         n11605, n11606, n11607, n11608, n11609, n11610, n11611, n11612,
         n11613, n11614, n11615, n11616, n11617, n11618, n11619, n11620,
         n11621, n11622, n11623, n11624, n11625, n11626, n11627, n11628,
         n11629, n11630, n11631, n11632, n11633, n11634, n11635, n11636,
         n11637, n11638, n11639, n11640, n11641, n11642, n11643, n11644,
         n11645, n11646, n11647, n11648, n11649, n11650, n11651, n11652,
         n11653, n11654, n11656, n11657, n11658, n11659, n11660, n11661,
         n11662, n11663, n11664, n11665, n11666, n11667, n11668, n11669,
         n11670, n11671, n11672, n11673, n11674, n11675, n11676, n11677,
         n11678, n11679, n11680, n11681, n11682, n11683, n11684, n11685,
         n11686, n11687, n11688, n11689, n11690, n11691, n11692, n11693,
         n11694, n11695, n11696, n11697, n11698, n11699, n11700, n11701,
         n11702, n11703, n11704, n11705, n11706, n11707, n11708, n11709,
         n11710, n11711, n11712, n11713, n11714, n11715, n11716, n11717,
         n11718, n11719, n11720, n11721, n11722, n11723, n11724, n11725,
         n11726, n11727, n11728, n11729, n11730, n11731, n11732, n11733,
         n11734, n11735, n11736, n11737, n11738, n11739, n11740, n11741,
         n11742, n11743, n11744, n11745, n11746, n11747, n11748, n11749,
         n11750, n11751, n11752, n11753, n11754, n11755, n11756, n11757,
         n11758, n11759, n11760, n11761, n11762, n11763, n11764, n11765,
         n11766, n11767, n11768, n11769, n11770, n11771, n11772, n11773,
         n11774, n11775, n11776, n11777, n11778, n11779, n11780, n11781,
         n11782, n11783, n11784, n11785, n11786, n11787, n11788, n11789,
         n11790, n11791, n11792, n11793, n11794, n11795, n11796, n11797,
         n11798, n11799, n11800, n11801, n11802, n11803, n11804, n11805,
         n11806, n11807, n11808, n11809, n11810, n11811, n11812, n11813,
         n11814, n11815, n11816, n11817, n11818, n11819, n11820, n11821,
         n11822, n11823, n11824, n11825, n11826, n11827, n11828, n11829,
         n11830, n11831, n11832, n11833, n11834, n11835, n11836, n11837,
         n11838, n11839, n11840, n11841, n11842, n11843, n11844, n11845,
         n11846, n11847, n11848, n11849, n11850, n11851, n11852, n11853,
         n11854, n11855, n11856, n11857, n11858, n11859, n11860, n11861,
         n11862, n11863, n11864, n11865, n11866, n11867, n11868, n11869,
         n11870, n11871, n11872, n11873, n11874, n11875, n11876, n11877,
         n11878, n11879, n11880, n11881, n11882, n11883, n11884, n11885,
         n11886, n11887, n11888, n11889, n11890, n11891, n11892, n11893,
         n11894, n11895, n11896, n11897, n11898, n11899, n11900, n11901,
         n11902, n11903, n11904, n11905, n11906, n11907, n11908, n11909,
         n11910, n11911, n11912, n11913, n11914, n11915, n11916, n11917,
         n11918, n11919, n11920, n11921, n11922, n11923, n11924, n11925,
         n11926, n11927, n11928, n11929, n11930, n11931, n11932, n11933,
         n11934, n11935, n11936, n11937, n11938, n11939, n11940, n11941,
         n11942, n11943, n11944, n11945, n11946, n11947, n11948, n11949,
         n11950, n11951, n11952, n11953, n11954, n11955, n11956, n11957,
         n11958, n11959, n11960, n11961, n11962, n11963, n11964, n11965,
         n11966, n11967, n11968, n11969, n11970, n11971, n11972, n11973,
         n11974, n11975, n11976, n11977, n11978, n11979, n11980, n11981,
         n11982, n11983, n11984, n11985, n11986, n11987, n11988, n11989,
         n11990, n11991, n11992, n11993, n11994, n11995, n11996, n11997,
         n11998, n11999, n12000, n12001, n12002, n12003, n12004, n12005,
         n12006, n12007, n12008, n12009, n12010, n12011, n12012, n12013,
         n12014, n12015, n12016, n12017, n12018, n12019, n12020, n12021,
         n12022, n12023, n12024, n12025, n12026, n12027, n12028, n12029,
         n12030, n12031, n12032, n12033, n12034, n12035, n12036, n12037,
         n12038, n12039, n12040, n12041, n12042, n12043, n12044, n12045,
         n12046, n12047, n12048, n12049, n12050, n12051, n12052, n12053,
         n12054, n12055, n12056, n12057, n12058, n12059, n12060, n12061,
         n12062, n12063, n12064, n12065, n12066, n12067, n12068, n12069,
         n12070, n12071, n12072, n12073, n12074, n12075, n12076, n12077,
         n12078, n12079, n12080, n12081, n12082, n12083, n12084, n12085,
         n12086, n12087, n12088, n12089, n12090, n12091, n12092, n12093,
         n12094, n12095, n12096, n12097, n12098, n12099, n12100, n12101,
         n12102, n12103, n12104, n12105, n12106, n12107, n12108, n12109,
         n12110, n12111, n12112, n12113, n12114, n12115, n12116, n12117,
         n12118, n12119, n12120, n12121, n12122, n12123, n12124, n12125,
         n12126, n12127, n12128, n12129, n12130, n12131, n12132, n12133,
         n12134, n12135, n12136, n12137, n12138, n12139, n12140, n12141,
         n12142, n12143, n12144, n12145, n12146, n12147, n12148, n12149,
         n12150, n12151, n12152, n12153, n12154, n12155, n12156, n12157,
         n12158, n12159, n12160, n12161, n12162, n12163, n12164, n12165,
         n12166, n12167, n12168, n12169, n12170, n12171, n12172, n12173,
         n12174, n12175, n12176, n12177, n12178, n12179, n12180, n12181,
         n12182, n12183, n12184, n12185, n12186, n12187, n12188, n12189,
         n12190, n12191, n12192, n12193, n12194, n12195, n12196, n12197,
         n12198, n12199, n12200, n12201, n12202, n12203, n12204, n12205,
         n12206, n12207, n12208, n12209, n12210, n12211, n12212, n12213,
         n12214, n12215, n12216, n12217, n12218, n12219, n12220, n12221,
         n12222, n12223, n12224, n12225, n12226, n12227, n12228, n12229,
         n12230, n12231, n12232, n12233, n12234, n12235, n12236, n12237,
         n12238, n12239, n12240, n12241, n12242, n12243, n12244, n12245,
         n12246, n12247, n12248, n12249, n12250, n12251, n12252, n12253,
         n12254, n12255, n12256, n12257, n12258, n12259, n12260, n12261,
         n12262, n12263, n12264, n12265, n12266, n12267, n12268, n12269,
         n12270, n12271, n12272, n12273, n12274, n12275, n12276, n12277,
         n12278, n12279, n12280, n12281, n12282, n12283, n12284, n12285,
         n12286, n12287, n12288, n12289, n12290, n12291, n12292, n12293,
         n12294, n12295, n12296, n12297, n12298, n12299, n12300, n12301,
         n12302, n12303, n12304, n12305, n12306, n12307, n12308, n12309,
         n12310, n12311, n12312, n12313, n12314, n12315, n12316, n12317,
         n12318, n12319, n12320, n12321, n12322, n12323, n12324, n12325,
         n12326, n12327, n12328, n12329, n12330, n12331, n12332, n12333,
         n12334, n12335, n12336, n12337, n12338, n12339, n12340, n12341,
         n12342, n12343, n12344, n12345, n12346, n12347, n12348, n12349,
         n12350, n12351, n12352, n12353, n12354, n12355, n12356, n12357,
         n12358, n12359, n12360, n12361, n12362, n12363, n12364, n12365,
         n12366, n12367, n12368, n12369, n12370, n12371, n12372, n12373,
         n12374, n12375, n12376, n12377, n12378, n12379, n12380, n12381,
         n12382, n12383, n12384, n12385, n12386, n12387, n12388, n12389,
         n12390, n12391, n12392, n12393, n12394, n12395, n12396, n12397,
         n12398, n12399, n12400, n12401, n12402, n12403, n12404, n12405,
         n12406, n12407, n12408, n12409, n12410, n12411, n12412, n12413,
         n12414, n12415, n12416, n12417, n12418, n12419, n12420, n12421,
         n12422, n12423, n12424, n12425, n12426, n12427, n12428, n12429,
         n12430, n12431, n12432, n12433, n12434, n12435, n12436, n12437,
         n12438, n12439, n12440, n12441, n12442, n12443, n12444, n12445,
         n12446, n12447, n12448, n12449, n12450, n12451, n12452, n12453,
         n12454, n12455, n12456, n12457, n12458, n12459, n12460, n12461,
         n12462, n12463, n12464, n12465, n12466, n12467, n12468, n12469,
         n12470, n12471, n12472, n12473, n12474, n12475, n12476, n12477,
         n12478, n12479, n12480, n12481, n12482, n12483, n12484, n12485,
         n12486, n12487, n12488, n12489, n12490, n12491, n12492, n12493,
         n12494, n12495, n12496, n12497, n12498, n12499, n12500, n12501,
         n12502, n12503, n12504, n12505, n12506, n12507, n12508, n12509,
         n12510, n12511, n12512, n12513, n12514, n12515, n12516, n12517,
         n12518, n12519, n12520, n12521, n12522, n12523, n12524, n12525,
         n12526, n12527, n12528, n12529, n12530, n12531, n12532, n12533,
         n12534, n12535, n12536, n12537, n12538, n12539, n12540, n12541,
         n12542, n12543, n12544, n12545, n12546, n12547, n12548, n12549,
         n12550, n12551, n12552, n12553, n12554, n12555, n12556, n12557,
         n12558, n12559, n12560, n12561, n12562, n12563, n12564, n12565,
         n12566, n12567, n12568, n12569, n12570, n12571, n12572, n12573,
         n12574, n12575, n12576, n12577, n12578, n12579, n12580, n12581,
         n12582, n12583, n12584, n12585, n12586, n12587, n12588, n12589,
         n12590, n12591, n12592, n12593, n12594, n12595, n12596, n12597,
         n12598, n12599, n12600, n12601, n12602, n12603, n12604, n12605,
         n12606, n12607, n12608, n12609, n12610, n12611, n12612, n12613,
         n12614, n12615, n12616, n12617, n12618, n12619, n12620, n12621,
         n12622, n12623, n12624, n12625, n12626, n12627, n12628, n12629,
         n12630, n12631, n12632, n12633, n12634, n12635, n12636, n12637,
         n12638, n12639, n12640, n12641, n12642, n12643, n12644, n12645,
         n12646, n12647, n12648, n12649, n12650, n12651, n12652, n12653,
         n12654, n12655, n12656, n12657, n12658, n12659, n12660, n12661,
         n12662, n12663, n12664, n12665, n12666, n12667, n12668, n12669,
         n12670, n12671, n12672, n12673, n12674, n12675, n12676, n12677,
         n12678, n12679, n12680, n12681, n12682, n12683, n12684, n12685,
         n12686, n12687, n12688, n12689, n12690, n12691, n12692, n12693,
         n12694, n12695, n12696, n12697, n12698, n12699, n12700, n12701,
         n12702, n12703, n12704, n12705, n12706, n12707, n12708, n12709,
         n12710, n12711, n12712, n12713, n12714, n12715, n12716, n12717,
         n12718, n12719, n12720, n12721, n12722, n12723, n12724, n12725,
         n12726, n12727, n12728, n12729, n12730, n12731, n12732, n12733,
         n12734, n12735, n12736, n12737, n12738, n12739, n12740, n12741,
         n12742, n12743, n12744, n12745, n12746, n12747, n12748, n12749,
         n12750, n12751, n12752, n12753, n12754, n12755, n12756, n12757,
         n12758, n12759, n12760, n12761, n12762, n12763, n12764, n12765,
         n12766, n12767, n12768, n12769, n12770, n12771, n12772, n12773,
         n12774, n12775, n12776, n12777, n12778, n12779, n12780, n12781,
         n12782, n12783, n12784, n12785, n12786, n12787, n12788, n12789,
         n12790, n12791, n12792, n12793, n12794, n12795, n12796, n12797,
         n12798, n12799, n12800, n12801, n12802, n12803, n12804, n12805,
         n12806, n12807, n12808, n12809, n12810, n12811, n12812, n12813,
         n12814, n12815, n12816, n12817, n12818, n12819, n12820, n12821,
         n12822, n12823, n12824, n12825, n12826, n12827, n12828, n12829,
         n12830, n12831, n12832, n12833, n12834, n12835, n12836, n12837,
         n12838, n12839, n12840, n12841, n12842, n12843, n12844, n12845,
         n12846, n12847, n12848, n12849, n12850, n12851, n12852, n12853,
         n12854, n12855, n12856, n12857, n12858, n12859, n12860, n12861,
         n12862, n12863, n12864, n12865, n12866, n12867, n12868, n12869,
         n12870, n12871, n12872, n12873, n12874, n12875, n12876, n12877,
         n12878, n12879, n12880, n12881, n12882, n12883, n12884, n12885,
         n12886, n12887, n12888, n12889, n12890, n12891, n12892, n12893,
         n12894, n12895, n12896, n12897, n12898, n12899, n12900, n12901,
         n12902, n12903, n12904, n12905, n12906, n12907, n12908, n12909,
         n12910, n12911, n12912, n12913, n12914, n12915, n12916, n12917,
         n12918, n12919, n12920, n12921, n12922, n12923, n12924, n12925,
         n12926, n12927, n12928, n12929, n12930, n12931, n12932, n12933,
         n12934, n12935, n12936, n12937, n12938, n12939, n12940, n12941,
         n12942, n12943, n12944, n12945, n12946, n12947, n12948, n12949,
         n12950, n12951, n12952, n12953, n12954, n12955, n12956, n12957,
         n12958, n12959, n12960, n12961, n12962, n12963, n12964, n12965,
         n12966, n12967, n12968, n12969, n12970, n12971, n12972, n12973,
         n12974, n12975, n12976, n12977, n12978, n12979, n12980, n12981,
         n12982, n12983, n12984, n12985, n12986, n12987, n12988, n12989,
         n12990, n12991, n12992, n12993, n12994, n12995, n12996, n12997,
         n12998, n12999, n13000, n13001, n13002, n13003, n13004, n13005,
         n13006, n13007, n13008, n13009, n13010, n13011, n13012, n13013,
         n13014, n13015, n13016, n13017, n13018, n13019, n13020, n13021,
         n13022, n13023, n13024, n13025, n13026, n13027, n13028, n13029,
         n13030, n13031, n13032, n13033, n13034, n13035, n13036, n13037,
         n13038, n13039, n13040, n13041, n13042, n13043, n13044, n13045,
         n13046, n13047, n13048, n13049, n13050, n13051, n13052, n13053,
         n13054, n13055, n13056, n13057, n13058, n13059, n13060, n13061,
         n13062, n13063, n13064, n13065, n13066, n13067, n13068, n13069,
         n13070, n13071, n13072, n13073, n13074, n13075, n13076, n13077,
         n13078, n13079, n13080, n13081, n13082, n13083, n13084, n13085,
         n13086, n13087, n13088, n13089, n13090, n13091, n13092, n13093,
         n13094, n13095, n13096, n13097, n13098, n13099, n13100, n13101,
         n13102, n13103, n13104, n13105, n13106, n13107, n13108, n13109,
         n13110, n13111, n13112, n13113, n13114, n13115, n13116, n13117,
         n13118, n13119, n13120, n13121, n13122, n13123, n13124, n13125,
         n13126, n13127, n13128, n13129, n13130, n13131, n13132, n13133,
         n13134, n13135, n13136, n13137, n13138, n13139, n13140, n13141,
         n13142, n13143, n13144, n13145, n13146, n13147, n13148, n13149,
         n13150, n13151, n13152, n13153, n13154, n13155, n13156, n13157,
         n13158, n13159, n13160, n13161, n13162, n13163, n13164, n13165,
         n13166, n13167, n13168, n13169, n13170, n13171, n13172, n13174,
         n13175, n13176, n13177, n13178, n13179, n13180, n13181, n13182,
         n13183, n13184, n13185, n13186, n13187, n13188, n13189, n13190,
         n13191, n13192, n13193, n13194, n13195, n13196, n13197, n13198,
         n13199, n13200, n13201, n13202, n13203, n13204, n13205, n13206,
         n13207, n13208, n13209, n13210, n13211, n13212, n13213, n13214,
         n13215, n13216, n13217, n13218, n13219, n13220, n13221, n13222,
         n13223, n13224, n13225, n13226, n13227, n13228, n13229, n13230,
         n13231, n13232, n13233, n13234, n13235, n13236, n13237, n13238,
         n13239, n13240, n13241, n13242, n13243, n13244, n13245, n13246,
         n13247, n13248, n13249, n13250, n13251, n13252, n13253, n13254,
         n13255, n13256, n13257, n13258, n13259, n13260, n13261, n13262,
         n13263, n13264, n13265, n13266, n13267, n13268, n13269, n13270,
         n13271, n13272, n13273, n13274, n13275, n13276, n13277, n13278,
         n13279, n13280, n13281, n13282, n13283, n13284, n13285, n13286,
         n13287, n13288, n13289, n13290, n13291, n13292, n13293, n13294,
         n13295, n13296, n13297, n13298, n13299, n13300, n13301, n13302,
         n13303, n13304, n13305, n13306, n13307, n13308, n13309, n13310,
         n13311, n13312, n13313, n13314, n13315, n13316, n13317, n13318,
         n13319, n13320, n13321, n13322, n13323, n13324, n13325, n13326,
         n13327, n13328, n13329, n13330, n13331, n13332, n13333, n13334,
         n13335, n13336, n13337, n13338, n13339, n13340, n13341, n13342,
         n13343, n13344, n13345, n13346, n13347, n13348, n13349, n13350,
         n13351, n13352, n13353, n13354, n13355, n13356, n13357, n13358,
         n13359, n13360, n13361, n13362, n13363, n13364, n13365, n13366,
         n13367, n13368, n13369, n13370, n13371, n13372, n13373, n13374,
         n13375, n13376, n13377, n13378, n13379, n13380, n13381, n13382,
         n13383, n13384, n13385, n13386, n13387, n13388, n13389, n13390,
         n13391, n13392, n13393, n13394, n13395, n13396, n13397, n13398,
         n13399, n13400, n13401, n13402, n13403, n13404, n13405, n13406,
         n13407, n13408, n13409, n13410, n13411, n13412, n13413, n13414,
         n13415, n13416, n13417, n13418, n13419, n13420, n13421, n13422,
         n13423, n13424, n13425, n13426, n13427, n13428, n13429, n13430,
         n13431, n13432, n13433, n13434, n13435, n13436, n13437, n13438,
         n13439, n13440, n13441, n13442, n13443, n13444, n13445, n13446,
         n13447, n13448, n13449, n13450, n13451, n13452, n13453, n13454,
         n13455, n13456, n13457, n13458, n13459, n13460, n13461, n13462,
         n13463, n13464, n13465, n13466, n13467, n13468, n13469, n13470,
         n13471, n13472, n13473, n13474, n13475, n13476, n13477, n13478,
         n13479, n13480, n13481, n13482, n13483, n13484, n13485, n13486,
         n13487, n13488, n13489, n13490, n13491, n13492, n13493, n13494,
         n13495, n13496, n13497, n13498, n13499, n13500, n13501, n13502,
         n13503, n13504, n13505, n13506, n13507, n13508, n13509, n13510,
         n13511, n13512, n13513, n13514, n13515, n13516, n13517, n13518,
         n13519, n13520, n13521, n13522, n13523, n13524, n13525, n13526,
         n13527, n13528, n13529, n13530, n13531, n13532, n13533, n13534,
         n13535, n13536, n13537, n13538, n13539, n13540, n13541, n13542,
         n13543, n13544, n13545, n13546, n13547, n13548, n13549, n13550,
         n13551, n13552, n13553, n13554, n13555, n13556, n13557, n13558,
         n13559, n13560, n13561, n13562, n13563, n13564, n13565, n13566,
         n13567, n13568, n13569, n13570, n13571, n13572, n13573, n13574,
         n13575, n13576, n13577, n13578, n13579, n13580, n13581, n13582,
         n13583, n13584, n13585, n13586, n13587, n13588, n13589, n13590,
         n13591, n13592, n13593, n13594, n13595, n13596, n13597, n13598,
         n13599, n13600, n13601, n13602, n13603, n13604, n13605, n13606,
         n13607, n13608, n13609, n13610, n13611, n13612, n13613, n13614,
         n13615, n13616, n13617, n13618, n13619, n13620, n13621, n13622,
         n13623, n13624, n13625, n13626, n13627, n13628, n13629, n13630,
         n13631, n13632, n13633, n13634, n13635, n13636, n13637, n13638,
         n13639, n13640, n13641, n13642, n13643, n13644, n13645, n13646,
         n13647, n13648, n13649, n13650, n13651, n13652, n13653, n13654,
         n13655, n13656, n13657, n13658, n13659, n13660, n13661, n13662,
         n13663, n13664, n13665, n13666, n13667, n13668, n13669, n13670,
         n13671, n13672, n13673, n13674, n13675, n13676, n13677, n13678,
         n13679, n13680, n13681, n13682, n13683, n13684, n13685, n13686,
         n13687, n13688, n13689, n13690, n13691, n13692, n13693, n13694,
         n13695, n13696, n13697, n13698, n13699, n13700, n13701, n13702,
         n13703, n13704, n13705, n13706, n13707, n13708, n13709, n13710,
         n13711, n13712, n13713, n13714, n13715, n13716, n13717, n13718,
         n13719, n13720, n13721, n13722, n13723, n13724, n13725, n13726,
         n13727, n13728, n13729, n13730, n13731, n13732, n13733, n13734,
         n13735, n13736, n13737, n13738, n13739, n13740, n13741, n13742,
         n13743, n13744, n13745, n13746, n13747, n13748, n13749, n13750,
         n13751, n13752, n13753, n13754, n13755, n13756, n13757, n13758,
         n13759, n13760, n13761, n13762, n13763, n13764, n13765, n13766,
         n13767, n13768, n13769, n13770, n13771, n13772, n13773, n13774,
         n13775, n13776, n13777, n13778, n13779, n13780, n13781, n13783,
         n13784, n13785, n13786, n13787, n13788, n13789, n13790, n13791,
         n13792, n13793, n13794, n13795, n13796, n13797, n13798, n13799,
         n13800, n13801, n13802, n13803, n13804, n13805, n13806, n13807,
         n13808, n13809, n13810, n13811, n13812, n13813, n13814, n13815,
         n13816, n13817, n13818, n13819, n13820, n13821, n13822, n13823,
         n13824, n13825, n13826, n13827, n13828, n13829, n13830, n13831,
         n13832, n13833, n13834, n13835, n13836, n13837, n13838, n13839,
         n13840, n13841, n13842, n13843, n13844, n13845, n13846, n13847,
         n13848, n13849, n13850, n13851, n13852, n13853, n13854, n13855,
         n13856, n13857, n13858, n13859, n13860, n13861, n13862, n13863,
         n13864, n13865, n13866, n13867, n13868, n13869, n13870, n13871,
         n13872, n13873, n13874, n13875, n13876, n13877, n13878, n13879,
         n13880, n13881, n13882, n13883, n13884, n13885, n13886, n13887,
         n13888, n13889, n13890, n13891, n13892, n13893, n13894, n13895,
         n13896, n13897, n13898, n13899, n13900, n13901, n13902, n13903,
         n13904, n13905, n13906, n13907, n13908, n13909, n13910, n13911,
         n13912, n13913, n13914, n13915, n13916, n13917, n13918, n13919,
         n13920, n13921, n13922, n13923, n13924, n13925, n13926, n13927,
         n13928, n13929, n13930, n13931, n13932, n13933, n13934, n13935,
         n13936, n13937, n13938, n13939, n13940, n13941, n13942, n13943,
         n13944, n13945, n13946, n13947, n13948, n13949, n13950, n13951,
         n13952, n13953, n13954, n13955, n13956, n13957, n13958, n13959,
         n13960, n13961, n13962, n13963, n13964, n13965, n13966, n13967,
         n13968, n13969, n13970, n13971, n13972, n13973, n13974, n13975,
         n13976, n13977, n13978, n13979, n13980, n13981, n13982, n13983,
         n13984, n13985, n13986, n13987, n13988, n13989, n13990, n13991,
         n13992, n13993, n13994, n13995, n13996, n13997, n13998, n13999,
         n14000, n14001, n14002, n14003, n14004, n14005, n14006, n14007,
         n14008, n14009, n14010, n14011, n14012, n14013, n14014, n14015,
         n14016, n14017, n14018, n14019, n14020, n14021, n14022, n14023,
         n14024, n14025, n14026, n14027, n14028, n14029, n14030, n14031,
         n14032, n14033, n14034, n14035, n14036, n14037, n14038, n14039,
         n14040, n14041, n14042, n14043, n14044, n14045, n14046, n14047,
         n14048, n14049, n14050, n14051, n14052, n14053, n14054, n14055,
         n14056, n14057, n14058, n14059, n14060, n14061, n14062, n14063,
         n14064, n14065, n14066, n14067, n14068, n14069, n14070, n14071,
         n14072, n14073, n14074, n14075, n14076, n14077, n14078, n14079,
         n14080, n14081, n14082, n14083, n14084, n14085, n14086, n14087,
         n14088, n14089, n14090, n14091, n14092, n14093, n14094, n14095,
         n14096, n14097, n14098, n14099, n14100, n14101, n14102, n14103,
         n14104, n14105, n14106, n14107, n14108, n14109, n14110, n14111,
         n14112, n14113, n14114, n14116, n14117, n14118, n14119, n14120,
         n14121, n14122, n14123, n14124, n14125, n14126, n14127, n14128,
         n14129, n14130, n14131, n14132, n14133, n14134, n14135, n14136,
         n14137, n14138, n14139, n14140, n14141, n14142, n14143, n14144,
         n14145, n14146, n14147, n14148, n14149, n14150, n14151, n14152,
         n14153, n14154, n14155, n14156, n14157, n14158, n14159, n14160,
         n14161, n14162, n14163, n14164, n14165, n14166, n14167, n14168,
         n14169, n14170, n14171, n14172, n14173, n14174, n14175, n14176,
         n14177, n14178, n14179, n14180, n14181, n14182, n14183, n14184,
         n14185, n14186, n14187, n14188, n14189, n14190, n14191, n14192,
         n14193, n14194, n14195, n14196, n14197, n14198, n14199, n14200,
         n14201, n14202, n14203, n14204, n14205, n14206, n14207, n14208,
         n14209, n14210, n14211, n14212, n14213, n14214, n14215, n14216,
         n14217, n14218, n14219, n14220, n14221, n14222, n14223, n14224,
         n14225, n14226, n14227, n14228, n14229, n14230, n14231, n14232,
         n14233, n14234, n14235, n14236, n14237, n14238, n14239, n14240,
         n14241, n14242, n14243, n14244, n14245, n14246, n14247, n14248,
         n14249, n14250, n14251, n14252, n14253, n14254, n14255, n14256,
         n14257, n14258, n14259, n14260, n14261, n14262, n14263, n14264,
         n14265, n14266, n14267, n14268, n14269, n14270, n14271, n14272,
         n14273, n14274, n14275, n14276, n14277, n14278, n14279, n14280,
         n14281, n14282, n14283, n14284, n14285, n14286, n14287, n14288,
         n14289, n14290, n14291, n14292, n14293, n14294, n14295, n14296,
         n14297, n14298, n14299, n14300, n14301, n14302, n14303, n14304,
         n14305, n14306, n14307, n14308, n14309, n14310, n14311, n14312,
         n14313, n14314, n14315, n14316, n14317, n14318, n14319, n14320,
         n14321, n14322, n14323, n14324, n14325, n14326, n14327, n14328,
         n14329, n14330, n14331, n14332, n14333, n14334, n14335, n14336,
         n14337, n14338, n14339, n14340, n14341, n14342, n14343, n14344,
         n14345, n14346, n14347, n14348, n14349, n14350, n14351, n14352,
         n14353, n14354, n14355, n14356, n14357, n14358, n14359, n14360,
         n14361, n14362, n14363, n14364, n14365, n14366, n14367, n14368,
         n14369, n14370, n14371, n14372, n14373, n14374, n14375, n14376,
         n14377, n14378, n14379, n14380, n14381, n14382, n14383, n14384,
         n14385, n14386, n14387, n14388, n14389, n14390, n14391, n14392,
         n14393, n14394, n14395, n14396, n14397, n14398, n14399, n14400,
         n14401, n14402, n14403, n14404, n14405, n14406, n14407, n14408,
         n14409, n14410, n14411, n14412, n14413, n14414, n14415, n14416,
         n14417, n14418, n14419, n14420, n14421, n14422, n14423, n14424,
         n14425, n14426, n14427, n14428, n14429, n14430, n14431, n14432,
         n14433, n14434, n14435, n14436, n14437, n14438, n14439, n14440,
         n14441, n14442, n14443, n14444, n14445, n14446, n14447, n14448,
         n14449, n14450, n14451, n14452, n14453, n14454, n14455, n14456,
         n14457, n14458, n14459, n14460, n14461, n14462, n14463, n14464,
         n14465, n14466, n14467, n14468, n14469, n14470, n14471, n14472,
         n14473, n14474, n14475, n14476, n14477, n14478, n14479, n14480,
         n14481, n14482, n14483, n14484, n14485, n14486, n14487, n14488,
         n14489, n14490, n14491, n14492, n14493, n14494, n14495, n14496,
         n14497, n14498, n14499, n14500, n14501, n14502, n14503, n14504,
         n14505, n14506, n14507, n14508, n14509, n14510, n14511, n14512,
         n14513, n14514, n14515, n14516, n14517, n14518, n14519, n14520,
         n14521, n14522, n14523, n14524, n14525, n14526, n14527, n14528,
         n14529, n14530, n14531, n14532, n14533, n14534, n14535, n14536,
         n14537, n14538, n14539, n14540, n14541, n14542, n14543, n14544,
         n14545, n14546, n14547, n14548, n14549, n14550, n14551, n14552,
         n14553, n14554, n14555, n14556, n14557, n14558, n14559, n14560,
         n14561, n14562, n14563, n14564, n14565, n14566, n14567, n14568,
         n14569, n14570, n14571, n14572, n14573, n14574, n14575, n14576,
         n14577, n14578, n14579, n14580, n14581, n14582, n14583, n14584,
         n14585, n14586, n14587, n14588, n14589, n14590, n14591, n14592,
         n14593, n14594, n14595, n14596, n14597, n14598, n14599, n14600,
         n14601, n14602, n14603, n14604, n14605, n14606, n14607, n14608,
         n14609, n14610, n14611, n14612, n14613, n14614, n14615, n14616,
         n14617, n14618, n14619, n14620, n14621, n14622, n14623, n14624,
         n14625, n14626, n14627, n14628, n14629, n14630, n14631, n14632,
         n14633, n14634, n14635, n14636, n14637, n14638, n14639, n14640,
         n14641, n14642, n14643, n14644, n14645, n14646, n14647, n14648,
         n14649, n14650, n14651, n14652, n14653, n14654, n14655, n14656,
         n14657, n14658, n14659, n14660, n14661, n14662, n14663, n14664,
         n14665, n14666, n14667, n14668, n14669, n14670, n14671, n14672,
         n14673, n14674, n14675, n14676, n14677, n14678, n14679, n14680,
         n14681, n14682, n14683, n14684, n14685, n14686, n14687, n14688,
         n14689, n14690, n14691, n14692, n14693, n14694, n14695, n14696,
         n14697, n14698, n14699, n14700, n14701, n14702, n14703, n14704,
         n14705, n14706, n14707, n14708, n14709, n14710, n14711, n14712,
         n14713, n14714, n14715, n14716, n14717, n14718, n14719, n14720,
         n14721, n14722, n14723, n14724, n14725, n14726, n14727, n14728,
         n14729, n14730, n14731, n14732, n14733, n14734, n14735, n14736,
         n14737, n14738, n14739, n14740, n14741, n14742, n14743, n14744,
         n14745, n14746, n14747, n14748, n14749, n14750, n14751, n14752,
         n14753, n14754, n14755, n14756, n14757, n14758, n14759, n14760,
         n14761, n14762, n14763, n14764, n14765, n14766, n14767, n14768,
         n14769, n14770, n14771, n14772, n14773, n14774, n14775, n14776,
         n14777, n14778, n14779, n14780, n14781, n14782, n14783, n14784,
         n14785, n14786, n14787, n14788, n14789, n14790, n14791, n14792,
         n14793, n14794, n14795, n14796, n14797, n14798, n14799, n14800,
         n14801, n14802, n14803, n14804, n14805, n14806, n14807, n14808,
         n14809, n14810, n14811, n14812, n14813, n14814, n14815, n14816,
         n14817, n14818, n14819, n14820, n14821, n14822, n14823, n14824,
         n14825, n14826, n14827, n14828, n14829, n14830, n14831, n14832,
         n14833, n14834, n14835, n14836, n14837, n14838, n14839, n14840,
         n14841, n14842, n14843, n14844, n14845, n14846, n14847, n14848,
         n14849, n14850, n14851, n14852, n14853, n14854, n14855, n14856,
         n14857, n14858, n14859, n14860, n14861, n14862, n14863, n14864,
         n14865, n14866, n14867, n14868, n14869, n14870, n14871, n14872,
         n14873, n14874, n14875, n14876, n14877, n14878, n14879, n14880,
         n14881, n14882, n14883, n14884, n14885, n14886, n14887, n14888,
         n14889, n14890, n14891, n14892, n14893, n14894, n14895, n14896,
         n14897, n14898, n14899, n14900, n14901, n14902, n14903, n14904,
         n14905, n14906, n14907, n14908, n14909, n14910, n14911, n14912,
         n14913, n14914, n14915, n14916, n14917, n14918, n14919, n14920,
         n14921, n14922, n14923, n14924, n14925, n14926, n14927, n14928,
         n14929, n14930, n14931, n14932, n14933, n14934, n14935, n14936,
         n14937, n14938, n14939, n14940, n14941, n14942, n14943, n14944,
         n14945, n14946, n14947, n14948, n14949, n14950, n14951, n14952,
         n14953, n14954, n14955, n14956, n14957, n14958, n14959, n14960,
         n14961, n14962, n14963, n14964, n14965, n14966, n14967, n14968,
         n14969, n14970, n14971, n14972, n14973, n14974, n14975, n14976,
         n14977, n14978, n14979, n14980, n14981, n14982, n14983, n14984,
         n14985, n14986, n14987, n14988, n14989, n14990, n14991, n14992,
         n14993, n14994, n14995, n14996, n14997, n14998, n14999, n15000,
         n15001, n15002, n15003, n15004, n15005, n15006, n15007, n15008,
         n15009, n15010, n15011, n15012, n15013, n15014, n15015, n15016,
         n15017, n15018, n15019, n15020, n15021, n15022, n15023, n15024,
         n15025, n15026, n15027, n15028, n15029, n15030, n15031, n15032,
         n15033, n15034, n15035, n15036, n15037, n15038, n15039, n15040,
         n15041, n15042, n15043, n15044, n15045, n15046, n15047, n15048,
         n15049, n15050, n15051, n15052, n15053, n15054, n15055, n15056,
         n15057, n15058, n15059, n15060, n15061, n15062, n15063, n15064,
         n15065, n15066, n15067, n15068, n15069, n15070, n15071, n15072,
         n15073, n15074, n15075, n15076, n15077, n15078, n15079, n15080,
         n15081, n15082, n15083, n15084, n15085, n15086, n15087, n15088,
         n15089, n15090, n15091, n15092, n15093, n15094, n15095, n15096,
         n15097, n15098, n15099, n15100, n15101, n15102, n15103, n15104,
         n15105, n15106, n15107, n15108, n15109, n15110, n15111, n15112,
         n15113, n15114, n15115, n15116, n15117, n15118, n15119, n15120,
         n15121, n15122, n15123, n15124, n15125, n15126, n15127, n15128,
         n15129, n15130, n15131, n15132, n15133, n15134, n15135, n15136,
         n15137, n15138, n15139, n15140, n15141, n15142, n15143, n15144,
         n15145, n15146, n15147, n15148, n15149, n15150, n15151, n15152,
         n15153, n15154, n15155, n15156, n15157, n15158, n15159, n15160,
         n15161, n15162, n15163, n15164, n15165, n15166, n15167, n15168,
         n15169, n15170, n15171, n15172, n15173, n15174, n15175, n15176,
         n15177, n15178, n15179, n15180, n15181, n15182, n15183, n15184,
         n15185, n15186, n15187, n15188, n15189, n15190, n15191, n15192,
         n15193, n15194, n15195, n15196, n15197, n15198, n15199, n15200,
         n15201, n15202, n15203, n15204, n15205, n15206, n15207, n15208,
         n15209, n15210, n15211, n15212, n15213, n15214, n15215, n15216,
         n15217, n15218, n15219, n15220, n15221, n15222, n15223, n15224,
         n15225, n15226, n15227, n15228, n15229, n15230, n15231, n15232,
         n15233, n15234, n15235, n15236, n15237, n15238, n15239, n15240,
         n15241, n15242, n15243, n15244, n15245, n15246, n15247, n15248,
         n15249, n15250, n15251, n15252, n15253, n15254, n15255, n15256,
         n15257, n15258, n15259, n15260, n15261, n15262, n15263, n15264,
         n15265, n15266, n15267, n15268, n15269, n15270, n15271, n15272,
         n15273, n15274, n15275, n15276, n15277, n15278, n15279, n15280,
         n15281, n15282, n15283, n15284, n15285, n15286, n15287, n15288,
         n15289, n15290, n15291, n15292, n15293, n15294, n15295, n15296,
         n15297, n15298, n15299, n15300, n15301, n15302, n15303, n15304,
         n15305, n15306, n15307, n15308, n15309, n15310, n15311, n15312,
         n15313, n15314, n15315, n15316, n15317, n15318, n15319, n15320,
         n15321, n15322, n15323, n15324, n15325, n15326, n15327, n15328,
         n15329, n15330, n15331, n15332, n15333, n15334, n15335, n15336,
         n15337, n15338, n15339, n15340, n15341, n15342, n15343, n15344,
         n15345, n15346, n15347, n15348, n15349, n15350, n15351, n15352,
         n15353, n15354, n15355, n15356, n15357, n15358, n15359, n15360,
         n15361, n15362, n15363, n15364, n15365, n15366, n15367, n15368,
         n15369, n15370, n15371, n15372, n15373, n15374, n15375, n15376,
         n15377, n15378, n15379, n15380, n15381, n15382, n15383, n15384,
         n15385, n15386, n15387, n15388, n15389, n15390, n15391, n15392,
         n15393, n15394, n15395, n15396, n15397, n15398, n15399, n15400,
         n15401, n15402, n15403, n15404, n15405, n15406, n15407, n15408,
         n15409, n15410, n15411, n15412, n15413, n15414, n15415, n15416,
         n15417, n15418, n15419, n15420, n15421, n15422, n15423, n15424,
         n15425, n15426, n15427, n15428, n15429, n15430, n15431, n15432,
         n15433, n15434, n15435, n15436, n15437, n15438, n15439, n15440,
         n15441, n15442, n15443, n15444, n15445, n15446, n15447, n15448,
         n15449, n15450, n15451, n15452, n15453, n15454, n15455, n15456,
         n15457, n15458, n15459, n15460, n15461, n15462, n15463, n15464,
         n15465, n15466, n15467, n15468, n15469, n15470, n15471, n15472,
         n15473, n15474, n15475, n15476, n15477, n15478, n15479, n15480,
         n15481, n15482, n15483, n15484, n15485, n15486, n15487, n15488,
         n15489, n15490, n15491, n15492, n15493, n15494, n15495, n15496,
         n15497, n15498, n15499, n15500, n15501, n15502, n15503, n15504,
         n15505, n15506, n15507, n15508, n15509, n15510, n15511, n15512,
         n15513, n15514, n15515, n15516, n15517, n15518, n15519, n15520,
         n15521, n15522, n15523, n15524, n15525, n15526, n15527, n15528,
         n15529, n15530, n15531, n15532, n15533, n15534, n15535, n15536,
         n15537, n15538, n15539, n15540, n15541, n15542, n15543, n15544,
         n15545, n15546, n15547, n15548, n15549, n15550, n15551, n15552,
         n15553, n15554, n15555, n15556, n15557, n15558, n15559, n15560,
         n15561, n15562, n15563, n15564, n15565, n15566, n15567, n15568,
         n15569, n15570, n15571, n15572, n15573, n15574, n15575, n15576,
         n15577, n15578, n15579, n15580, n15581, n15582, n15583, n15584,
         n15585, n15586, n15587, n15588, n15589, n15590, n15591, n15592,
         n15593, n15594, n15595, n15596, n15597, n15598, n15599, n15600,
         n15601, n15602, n15603, n15604, n15605, n15606, n15607, n15608,
         n15609, n15610, n15611, n15612, n15613, n15614, n15615, n15616,
         n15617, n15618, n15619, n15620, n15621, n15622, n15623, n15624,
         n15625, n15626, n15627, n15628, n15629, n15630, n15631, n15632,
         n15633, n15634, n15635, n15636, n15637, n15638, n15639, n15640,
         n15641, n15642, n15643, n15644, n15645, n15646, n15647, n15648,
         n15649, n15650, n15651, n15652, n15653, n15654, n15655, n15656,
         n15657, n15658, n15659, n15660, n15661, n15662, n15663, n15664,
         n15665, n15666, n15667, n15668, n15669, n15670, n15671, n15672,
         n15673, n15674, n15675, n15676, n15677, n15678, n15679, n15680,
         n15681, n15682, n15683, n15684, n15685, n15686, n15687, n15688,
         n15689, n15690, n15691, n15692, n15693, n15694, n15695, n15696,
         n15697, n15698, n15699, n15700, n15701, n15702, n15703, n15704,
         n15705, n15706, n15707, n15708, n15709, n15710, n15711, n15712,
         n15713, n15714, n15715, n15716, n15717, n15718, n15719, n15720,
         n15721, n15722, n15723, n15724, n15725, n15726, n15727, n15728,
         n15729, n15730, n15731, n15732, n15733, n15734, n15735, n15736,
         n15737, n15738, n15739, n15740, n15741, n15742, n15743, n15744,
         n15745, n15746, n15747, n15748, n15749, n15750, n15751, n15752,
         n15753, n15754, n15755, n15756, n15757, n15758, n15759, n15760,
         n15761, n15762, n15763, n15764, n15765, n15766, n15767, n15768,
         n15769, n15770, n15771, n15772, n15773, n15774, n15775, n15776,
         n15777, n15778, n15779, n15780, n15781, n15782, n15783, n15784,
         n15785, n15786, n15787, n15788, n15789, n15790, n15791, n15792,
         n15793, n15794, n15795, n15796, n15797, n15798, n15799, n15800,
         n15801, n15802, n15803, n15804, n15805, n15806, n15807, n15808,
         n15809, n15810, n15811, n15812, n15813, n15814, n15815, n15816,
         n15817, n15818, n15819, n15820, n15821, n15822, n15823, n15824,
         n15825, n15826, n15827, n15828, n15829, n15830, n15831, n15832,
         n15833, n15834, n15835, n15836, n15837, n15838, n15839, n15840,
         n15841, n15842, n15843, n15844, n15845, n15846, n15847, n15848,
         n15849, n15850, n15851, n15852, n15853, n15854, n15855, n15856,
         n15857, n15858, n15859, n15860, n15861, n15862, n15863, n15864,
         n15865, n15866, n15867, n15868, n15869, n15870, n15871, n15872,
         n15873, n15874, n15875, n15876, n15877, n15878, n15879, n15880,
         n15881, n15882, n15883, n15884, n15885, n15886, n15887, n15888,
         n15889, n15890, n15891, n15892, n15893, n15894, n15895, n15896,
         n15897, n15898, n15899, n15900, n15901, n15902, n15903, n15904,
         n15905, n15906, n15907, n15908, n15909, n15910, n15911, n15912,
         n15913, n15914, n15915, n15916, n15917, n15918, n15919, n15920,
         n15921, n15922, n15923, n15924, n15925, n15926, n15927, n15928,
         n15929, n15930, n15931, n15932, n15933, n15934, n15935, n15936,
         n15937, n15938, n15939, n15940, n15941, n15942, n15943, n15944,
         n15945, n15946, n15947, n15948, n15949, n15950, n15951, n15952,
         n15953, n15954, n15955, n15956, n15957, n15958, n15959, n15960,
         n15961, n15962, n15963, n15964, n15965, n15966, n15967, n15968,
         n15969, n15970, n15971, n15972, n15973, n15974, n15975, n15976,
         n15977, n15978, n15979, n15980, n15981, n15982, n15983, n15984,
         n15985, n15986, n15987, n15988, n15989, n15990, n15991, n15992,
         n15993, n15994, n15995, n15996, n15997, n15998, n15999, n16000,
         n16001, n16002, n16003, n16004, n16005, n16006, n16007, n16008,
         n16009, n16010, n16011, n16012, n16013, n16014, n16015, n16016,
         n16017, n16018, n16019, n16020, n16021, n16022, n16023, n16024,
         n16025, n16026, n16027, n16028, n16029, n16030, n16031, n16032,
         n16033, n16034, n16035, n16036, n16037, n16038, n16039, n16040,
         n16041, n16042, n16043, n16044, n16045, n16046, n16047, n16048,
         n16049, n16050, n16051, n16052, n16053, n16054, n16055, n16056,
         n16057, n16058, n16059, n16060, n16061, n16062, n16063, n16064,
         n16065, n16066, n16067, n16068, n16069, n16070, n16071, n16072,
         n16073, n16074, n16075, n16076, n16077, n16078, n16079, n16080,
         n16081, n16082, n16083, n16084, n16085, n16086, n16087, n16088,
         n16089, n16090, n16091, n16092, n16093, n16094, n16095, n16096,
         n16097, n16098, n16099, n16100, n16101, n16102, n16103, n16104,
         n16105, n16106, n16107, n16108, n16109, n16110, n16111, n16112,
         n16113, n16114, n16115, n16116, n16117, n16118, n16119, n16120,
         n16121, n16122, n16123, n16124, n16125, n16126, n16127, n16128,
         n16129, n16130, n16131, n16132, n16133, n16134, n16135, n16136,
         n16137, n16138, n16139, n16140, n16141, n16142, n16143, n16144,
         n16145, n16146, n16147, n16148, n16149, n16150, n16151, n16152,
         n16153, n16154, n16155, n16156, n16157, n16158, n16159, n16160,
         n16161, n16162, n16163, n16164, n16165, n16166, n16167, n16168,
         n16169, n16170, n16171, n16172, n16173, n16174, n16175, n16176,
         n16177, n16178, n16179, n16180, n16181, n16182, n16183, n16184,
         n16185, n16186, n16187, n16188, n16189, n16190, n16191, n16192,
         n16193, n16194, n16195, n16196, n16197, n16198, n16199, n16200,
         n16201, n16202, n16203, n16204, n16205, n16206, n16207, n16208,
         n16209, n16210, n16211, n16212, n16213, n16214, n16215, n16216,
         n16217, n16218, n16219, n16220, n16221, n16222, n16223, n16224,
         n16225, n16226, n16227, n16228, n16229, n16230, n16231, n16232,
         n16233, n16234, n16235, n16236, n16237, n16238, n16239, n16240,
         n16241, n16242, n16243, n16244, n16245, n16246, n16247, n16248,
         n16249, n16250, n16251, n16252, n16253, n16254, n16255, n16256,
         n16257, n16258, n16259, n16260, n16261, n16262, n16263, n16264,
         n16265, n16266, n16267, n16268, n16269, n16270, n16271, n16272,
         n16273, n16274, n16275, n16276, n16277, n16278, n16279, n16280,
         n16281, n16282, n16283, n16284, n16285, n16286, n16287, n16288,
         n16289, n16290, n16291, n16292, n16293, n16294, n16295, n16296,
         n16297, n16298, n16299, n16300, n16301, n16302, n16303, n16304,
         n16305, n16306, n16307, n16308, n16309, n16310, n16311, n16312,
         n16313, n16314, n16315, n16316, n16317, n16318, n16319, n16320,
         n16321, n16322, n16323, n16324, n16325, n16326, n16327, n16328,
         n16329, n16330, n16331, n16332, n16333, n16334, n16335, n16336,
         n16337, n16338, n16339, n16340, n16341, n16342, n16343, n16344,
         n16345, n16346, n16347, n16348, n16349, n16350, n16351, n16352,
         n16353, n16354, n16355, n16356, n16357, n16358, n16359, n16360,
         n16361, n16362, n16363, n16364, n16365, n16366, n16367, n16368,
         n16369, n16370, n16371, n16372, n16373, n16374, n16375, n16376,
         n16377, n16378, n16379, n16380, n16381, n16382, n16383, n16384,
         n16385, n16386, n16387, n16388, n16389, n16390, n16391, n16392,
         n16393, n16394, n16395, n16396, n16397, n16398, n16399, n16400,
         n16401, n16402, n16403, n16404, n16405, n16406, n16407, n16408,
         n16409, n16410, n16411, n16412, n16413, n16414, n16415, n16416,
         n16417, n16418, n16419, n16420, n16421, n16422, n16423, n16424,
         n16425, n16426, n16427, n16428, n16429, n16430, n16431, n16432,
         n16433, n16434, n16435, n16436, n16437, n16438, n16439, n16440,
         n16441, n16442, n16443, n16444, n16445, n16446, n16447, n16448,
         n16449, n16450, n16451, n16452, n16453, n16454, n16455, n16456,
         n16457, n16458, n16459, n16460, n16461, n16462, n16463, n16464,
         n16465, n16466, n16467, n16468, n16469, n16470, n16471, n16472,
         n16473, n16474, n16475, n16476, n16477, n16478, n16479, n16480,
         n16481, n16482, n16483, n16484, n16485, n16486, n16487, n16488,
         n16489, n16490, n16491, n16492, n16493, n16494, n16495, n16496,
         n16497, n16498, n16499, n16500, n16501, n16502, n16503, n16504,
         n16505, n16506, n16507, n16508, n16509, n16510, n16511, n16512,
         n16513, n16514, n16515, n16516, n16517, n16518, n16519, n16520,
         n16521, n16522, n16523, n16524, n16525, n16526, n16527, n16528,
         n16529, n16530, n16531, n16532, n16533, n16534, n16535, n16536,
         n16537, n16538, n16539, n16540, n16541, n16542, n16543, n16544,
         n16545, n16546, n16547, n16548, n16549, n16550, n16551, n16552,
         n16553, n16554, n16555, n16556, n16557, n16558, n16559, n16560,
         n16561, n16562, n16563, n16564, n16565, n16566, n16567, n16568,
         n16569, n16570, n16571, n16572, n16573, n16574, n16575, n16576,
         n16577, n16578, n16579, n16580, n16581, n16582, n16583, n16584,
         n16585, n16586, n16587, n16588, n16589, n16590, n16591, n16592,
         n16593, n16594, n16595, n16596, n16597, n16598, n16599, n16600,
         n16601, n16602, n16603, n16604, n16605, n16606, n16607, n16608,
         n16609, n16610, n16611, n16612, n16613, n16614, n16615, n16616,
         n16617, n16618, n16619, n16620, n16621, n16622, n16623, n16624,
         n16625, n16626, n16627, n16628, n16629, n16630, n16631, n16632,
         n16633, n16634, n16635, n16636, n16637, n16638, n16639, n16640,
         n16641, n16642, n16643, n16644, n16645, n16646, n16647, n16648,
         n16649, n16650, n16651, n16652, n16653, n16654, n16655, n16656,
         n16657, n16658, n16659, n16660, n16661, n16662, n16663, n16664,
         n16665, n16666, n16667, n16668, n16669, n16670, n16671, n16672,
         n16673, n16674, n16675, n16676, n16677, n16678, n16679, n16680,
         n16681, n16682, n16683, n16684, n16685, n16686, n16687, n16688,
         n16689, n16690, n16691, n16692, n16693, n16694, n16695, n16696,
         n16697, n16698, n16699, n16700, n16701, n16702, n16703, n16704,
         n16705, n16706, n16707, n16708, n16709, n16710, n16711, n16712,
         n16713, n16714, n16715, n16716, n16717, n16718, n16719, n16720,
         n16721, n16722, n16723, n16724, n16725, n16726, n16727, n16728,
         n16729, n16730, n16731, n16732, n16733, n16734, n16735, n16736,
         n16737, n16738, n16739, n16740, n16741, n16742, n16743, n16744,
         n16745, n16746, n16747, n16748, n16749, n16750, n16751, n16752,
         n16753, n16754, n16755, n16756, n16757, n16758, n16759, n16760,
         n16761, n16762, n16763, n16764, n16765, n16766, n16767, n16768,
         n16769, n16770, n16771, n16772, n16773, n16774, n16775, n16776,
         n16777, n16778, n16779, n16780, n16781, n16782, n16783, n16784,
         n16785, n16786, n16787, n16788, n16789, n16790, n16791, n16792,
         n16793, n16794, n16795, n16796, n16797, n16798, n16799, n16800,
         n16801, n16802, n16803, n16804, n16805, n16806, n16807, n16808,
         n16809, n16810, n16811, n16812, n16813, n16814, n16815, n16816,
         n16817, n16818, n16819, n16820, n16821, n16822, n16823, n16824,
         n16825, n16826, n16827, n16828, n16829, n16830, n16831, n16832,
         n16833, n16834, n16835, n16836, n16837, n16838, n16839, n16840,
         n16841, n16842, n16843, n16844, n16845, n16846, n16847, n16848,
         n16849, n16850, n16851, n16852, n16853, n16854, n16855, n16856,
         n16857, n16858, n16859, n16860, n16861, n16862, n16863, n16864,
         n16865, n16866, n16867, n16868, n16869, n16870, n16871, n16872,
         n16873, n16874, n16875, n16876, n16877, n16878, n16879, n16880,
         n16881, n16882, n16883, n16884, n16885, n16886, n16887, n16888,
         n16889, n16890, n16891, n16892, n16893, n16894, n16895, n16896,
         n16897, n16898, n16899, n16900, n16901, n16902, n16903, n16904,
         n16905, n16906, n16907, n16908, n16909, n16910, n16911, n16912,
         n16913, n16914, n16915, n16916, n16917, n16918, n16919, n16920,
         n16921, n16922, n16923, n16924, n16925, n16926, n16927, n16928,
         n16929, n16930, n16931, n16932, n16933, n16934, n16935, n16936,
         n16937, n16938, n16939, n16940, n16941, n16942, n16943, n16944,
         n16945, n16946, n16947, n16948, n16949, n16950, n16951, n16952,
         n16953, n16954, n16955, n16956, n16957, n16958, n16959, n16960,
         n16961, n16962, n16963, n16964, n16965, n16966, n16967, n16968,
         n16969, n16970, n16971, n16972, n16973, n16974, n16975, n16976,
         n16977, n16978, n16979, n16980, n16981, n16982, n16983, n16984,
         n16985, n16986, n16987, n16988, n16989, n16990, n16991, n16992,
         n16993, n16994, n16995, n16996, n16997, n16998, n16999, n17000,
         n17001, n17002, n17003, n17004, n17005, n17006, n17007, n17008,
         n17009, n17010, n17011, n17012, n17013, n17014, n17015, n17016,
         n17017, n17018, n17019, n17020, n17021, n17022, n17023, n17024,
         n17025, n17026, n17027, n17028, n17029, n17030, n17031, n17032,
         n17033, n17034, n17035, n17036, n17037, n17038, n17039, n17040,
         n17041, n17042, n17043, n17044, n17045, n17046, n17047, n17048,
         n17049, n17050, n17051, n17052, n17053, n17054, n17055, n17056,
         n17057, n17058, n17059, n17060, n17061, n17062, n17063, n17064,
         n17065, n17066, n17067, n17068, n17069, n17070, n17071, n17072,
         n17073, n17074, n17075, n17076, n17077, n17078, n17079, n17080,
         n17081, n17082, n17083, n17084, n17085, n17086, n17087, n17088,
         n17089, n17090, n17091, n17092, n17093, n17094, n17095, n17096,
         n17097, n17098, n17099, n17100, n17101, n17102, n17103, n17104,
         n17105, n17106, n17107, n17108, n17109, n17110, n17111, n17112,
         n17113, n17114, n17115, n17116, n17117, n17118, n17119, n17120,
         n17121, n17122, n17123, n17124, n17125, n17126, n17127, n17128,
         n17129, n17130, n17131, n17132, n17133, n17134, n17135, n17136,
         n17137, n17138, n17139, n17140, n17141, n17142, n17143, n17144,
         n17145, n17146, n17147, n17148, n17149, n17150, n17151, n17152,
         n17153, n17154, n17155, n17156, n17157, n17158, n17159, n17160,
         n17161, n17162, n17163, n17164, n17165, n17166, n17167, n17168,
         n17169, n17170, n17171, n17172, n17173, n17174, n17175, n17176,
         n17177, n17178, n17179, n17180, n17181, n17182, n17183, n17184,
         n17185, n17186, n17187, n17188, n17189, n17190, n17191, n17192,
         n17193, n17194, n17195, n17196, n17197, n17198, n17199, n17200,
         n17201, n17202, n17203, n17204, n17205, n17206, n17207, n17208,
         n17209, n17210, n17211, n17212, n17213, n17214, n17215, n17216,
         n17217, n17218, n17219, n17220, n17221, n17222, n17223, n17224,
         n17225, n17226, n17227, n17228, n17229, n17230, n17231, n17232,
         n17233, n17234, n17235, n17236, n17237, n17238, n17239, n17240,
         n17241, n17242, n17243, n17244, n17245, n17246, n17247, n17248,
         n17249, n17250, n17251, n17252, n17253, n17254, n17255, n17256,
         n17257, n17258, n17259, n17260, n17261, n17262, n17263, n17264,
         n17265, n17266, n17267, n17268, n17269, n17270, n17271, n17272,
         n17273, n17274, n17275, n17276, n17277, n17278, n17279, n17280,
         n17281, n17282, n17283, n17284, n17285, n17286, n17287, n17288,
         n17289, n17290, n17291, n17292, n17293, n17294, n17295, n17296,
         n17297, n17298, n17299, n17300, n17301, n17302, n17303, n17304,
         n17305, n17306, n17307, n17308, n17309, n17310, n17311, n17312,
         n17313, n17314, n17315, n17316, n17317, n17318, n17319, n17320,
         n17321, n17322, n17323, n17324, n17325, n17326, n17327, n17328,
         n17329, n17330, n17331, n17332, n17333, n17334, n17335, n17336,
         n17337, n17338, n17339, n17340, n17341, n17342, n17343, n17344,
         n17345, n17346, n17347, n17348, n17349, n17350, n17351, n17352,
         n17353, n17354, n17355, n17356, n17357, n17358, n17359, n17360,
         n17361, n17362, n17363, n17364, n17365, n17366, n17367, n17368,
         n17369, n17370, n17371, n17372, n17373, n17374, n17375, n17376,
         n17377, n17378, n17379, n17380, n17381, n17382, n17383, n17384,
         n17385, n17386, n17387, n17388, n17389, n17390, n17391, n17392,
         n17393, n17394, n17395, n17396, n17397, n17398, n17399, n17400,
         n17401, n17402, n17403, n17404, n17405, n17406, n17407, n17408,
         n17409, n17410, n17411, n17412, n17413, n17414, n17415, n17416,
         n17417, n17418, n17419, n17420, n17421, n17422, n17423, n17424,
         n17425, n17426, n17427, n17428, n17429, n17430, n17431, n17432,
         n17433, n17434, n17435, n17436, n17437, n17438, n17439, n17440,
         n17441, n17442, n17443, n17444, n17445, n17446, n17447, n17448,
         n17449, n17450, n17451, n17452, n17453, n17454, n17455, n17456,
         n17457, n17458, n17459, n17460, n17461, n17462, n17463, n17464,
         n17465, n17466, n17467, n17468, n17469, n17470, n17471, n17472,
         n17473, n17474, n17475, n17476, n17477, n17478, n17479, n17480,
         n17481, n17482, n17483, n17484, n17485, n17486, n17487, n17488,
         n17489, n17490, n17491, n17492, n17493, n17494, n17495, n17496,
         n17497, n17498, n17499, n17500, n17501, n17502, n17503, n17504,
         n17505, n17506, n17507, n17508, n17509, n17510, n17511, n17512,
         n17513, n17514, n17515, n17516, n17517, n17518, n17519, n17520,
         n17521, n17522, n17523, n17524, n17525, n17526, n17527, n17528,
         n17529, n17530, n17531, n17532, n17533, n17534, n17535, n17536,
         n17537, n17538, n17539, n17540, n17541, n17542, n17543, n17544,
         n17545, n17546, n17547, n17548, n17549, n17550, n17551, n17552,
         n17553, n17554, n17555, n17556, n17557, n17558, n17559, n17560,
         n17561, n17562, n17563, n17564, n17565, n17566, n17567, n17568,
         n17569, n17570, n17571, n17572, n17573, n17574, n17575, n17576,
         n17577, n17578, n17579, n17580, n17581, n17582, n17583, n17584,
         n17585, n17586, n17587, n17588, n17589, n17590, n17591, n17592,
         n17593, n17594, n17595, n17596, n17597, n17598, n17599, n17600,
         n17601, n17602, n17603, n17604, n17605, n17606, n17607, n17608,
         n17609, n17610, n17611, n17612, n17613, n17614, n17615, n17616,
         n17617, n17618, n17619, n17620, n17621, n17622, n17623, n17624,
         n17625, n17626, n17627, n17628, n17629, n17630, n17631, n17632,
         n17633, n17634, n17635, n17636, n17637, n17638, n17639, n17640,
         n17641, n17642, n17643, n17644, n17645, n17646, n17647, n17648,
         n17649, n17650, n17651, n17652, n17653, n17654, n17655, n17656,
         n17657, n17658, n17659, n17660, n17661, n17662, n17663, n17664,
         n17665, n17666, n17667, n17668, n17669, n17670, n17671, n17672,
         n17673, n17674, n17675, n17676, n17677, n17678, n17679, n17680,
         n17681, n17682, n17683, n17684, n17685, n17686, n17687, n17688,
         n17689, n17690, n17691, n17692, n17693, n17694, n17695, n17696,
         n17697, n17698, n17699, n17700, n17701, n17702, n17703, n17704,
         n17705, n17706, n17707, n17708, n17709, n17710, n17711, n17712,
         n17713, n17714, n17715, n17716, n17717, n17718, n17719, n17720,
         n17721, n17722, n17723, n17724, n17725, n17726, n17727, n17728,
         n17729, n17730, n17731, n17732, n17733, n17734, n17735, n17736,
         n17737, n17738, n17739, n17740, n17741, n17742, n17743, n17744,
         n17745, n17746, n17747, n17748, n17749, n17750, n17751, n17752,
         n17753, n17754, n17755, n17756, n17757, n17758, n17759, n17760,
         n17761, n17762, n17763, n17764, n17765, n17766, n17767, n17768,
         n17769, n17770, n17771, n17772, n17773, n17774, n17775, n17776,
         n17777, n17778, n17779, n17780, n17781, n17782, n17783, n17784,
         n17785, n17786, n17787, n17788, n17789, n17790, n17791, n17792,
         n17793, n17794, n17795, n17796, n17797, n17798, n17799, n17800,
         n17801, n17802, n17803, n17804, n17805, n17806, n17807, n17808,
         n17809, n17810, n17811, n17812, n17813, n17814, n17815, n17816,
         n17817, n17818, n17819, n17820, n17821, n17822, n17823, n17824,
         n17825, n17826, n17827, n17828, n17829, n17830, n17831, n17832,
         n17833, n17834, n17835, n17836, n17837, n17838, n17839, n17840,
         n17841, n17842, n17843, n17844, n17845, n17846, n17847, n17848,
         n17849, n17850, n17851, n17852, n17853, n17854, n17855, n17856,
         n17857, n17858, n17859, n17860, n17861, n17862, n17863, n17864,
         n17865, n17866, n17867, n17868, n17869, n17870, n17871, n17872,
         n17873, n17874, n17875, n17876, n17877, n17878, n17879, n17880,
         n17881, n17882, n17883, n17884, n17885, n17886, n17887, n17888,
         n17889, n17890, n17891, n17892, n17893, n17894, n17895, n17896,
         n17897, n17898, n17899, n17900, n17901, n17902, n17903, n17904,
         n17905, n17906, n17907, n17908, n17909, n17910, n17911, n17912,
         n17913, n17914, n17915, n17916, n17917, n17918, n17919, n17920,
         n17921, n17922, n17923, n17924, n17925, n17926, n17927, n17928,
         n17929, n17930, n17931, n17932, n17933, n17934, n17935, n17936,
         n17937, n17938, n17939, n17940, n17941, n17942, n17943, n17944,
         n17945, n17946, n17947, n17948, n17949, n17950, n17951, n17952,
         n17953, n17954, n17955, n17956, n17957, n17958, n17959, n17960,
         n17961, n17962, n17963, n17964, n17965, n17966, n17967, n17968,
         n17969, n17970, n17971, n17972, n17973, n17974, n17975, n17976,
         n17977, n17978, n17979, n17980, n17981, n17982, n17983, n17984,
         n17985, n17986, n17987, n17988, n17989, n17990, n17991, n17992,
         n17993, n17994, n17995, n17996, n17997, n17998, n17999, n18000,
         n18001, n18002, n18003, n18004, n18005, n18006, n18007, n18008,
         n18009, n18010, n18011, n18012, n18013, n18014, n18015, n18016,
         n18017, n18018, n18019, n18020, n18021, n18022, n18023, n18024,
         n18025, n18026, n18027, n18028, n18029, n18030, n18031, n18032,
         n18033, n18034, n18035, n18036, n18037, n18038, n18039, n18040,
         n18041, n18042, n18043, n18044, n18045, n18046, n18047, n18048,
         n18049, n18050, n18051, n18052, n18053, n18054, n18055, n18056,
         n18057, n18058, n18059, n18060, n18061, n18062, n18063, n18064,
         n18065, n18066, n18067, n18068, n18069, n18070, n18071, n18072,
         n18073, n18074, n18075, n18076, n18077, n18078, n18079, n18080,
         n18081, n18082, n18083, n18084, n18085, n18086, n18087, n18088,
         n18089, n18090, n18091, n18092, n18093, n18094, n18095, n18096,
         n18097, n18098, n18099, n18100, n18101, n18102, n18103, n18104,
         n18105, n18106, n18107, n18108, n18109, n18110, n18111, n18112,
         n18113, n18114, n18115, n18116, n18117, n18118, n18119, n18120,
         n18121, n18122, n18123, n18124, n18125, n18126, n18127, n18128,
         n18129, n18130, n18131, n18132, n18133, n18134, n18135, n18136,
         n18137, n18138, n18139, n18140, n18141, n18142, n18143, n18144,
         n18145, n18146, n18147, n18148, n18149, n18150, n18151, n18152,
         n18153, n18154, n18155, n18156, n18157, n18158, n18159, n18160,
         n18161, n18162, n18163, n18164, n18165, n18166, n18167, n18168,
         n18169, n18170, n18171, n18172, n18173, n18174, n18175, n18176,
         n18177, n18178, n18179, n18180, n18181, n18182, n18183, n18184,
         n18185, n18186, n18187, n18188, n18189, n18190, n18191, n18192,
         n18193, n18194, n18195, n18196, n18197, n18198, n18199, n18200,
         n18201, n18202, n18203, n18204, n18205, n18206, n18207, n18208,
         n18209, n18210, n18211, n18212, n18213, n18214, n18215, n18216,
         n18217, n18218, n18219, n18220, n18221, n18222, n18223, n18224,
         n18225, n18226, n18227, n18228, n18229, n18230, n18231, n18232,
         n18233, n18234, n18235, n18236, n18237, n18238, n18239, n18240,
         n18241, n18242, n18243, n18244, n18245, n18246, n18247, n18248,
         n18249, n18250, n18251, n18252, n18253, n18254, n18255, n18256,
         n18257, n18258, n18259, n18260, n18261, n18262, n18263, n18264,
         n18265, n18266, n18267, n18268, n18269, n18270, n18271, n18272,
         n18273, n18274, n18275, n18276, n18277, n18278, n18279, n18280,
         n18281, n18282, n18283, n18284, n18285, n18286, n18287, n18288,
         n18289, n18290, n18291, n18292, n18293, n18294, n18295, n18296,
         n18297, n18298, n18299, n18300, n18301, n18302, n18303, n18304,
         n18305, n18306, n18307, n18308, n18309, n18310, n18311, n18312,
         n18313, n18314, n18315, n18316, n18317, n18318, n18319, n18320,
         n18321, n18322, n18323, n18324, n18325, n18326, n18327, n18328,
         n18329, n18330, n18331, n18332, n18333, n18334, n18335, n18336,
         n18337, n18338, n18339, n18340, n18341, n18342, n18343, n18344,
         n18345, n18346, n18347, n18348, n18349, n18350, n18351, n18352,
         n18353, n18354, n18355, n18356, n18357, n18358, n18359, n18360,
         n18361, n18362, n18363, n18364, n18365, n18366, n18367, n18368,
         n18369, n18370, n18371, n18372, n18373, n18374, n18375, n18376,
         n18377, n18378, n18379, n18380, n18381, n18382, n18383, n18384,
         n18385, n18386, n18387, n18388, n18389, n18390, n18391, n18392,
         n18393, n18394, n18395, n18396, n18397, n18398, n18399, n18400,
         n18401, n18402, n18403, n18404, n18405, n18406, n18407, n18408,
         n18409, n18410, n18411, n18412, n18413, n18414, n18415, n18416,
         n18417, n18418, n18419, n18420, n18421, n18422, n18423, n18424,
         n18425, n18426, n18427, n18428, n18429, n18430, n18431, n18432,
         n18433, n18434, n18435, n18436, n18437, n18438, n18439, n18440,
         n18441, n18442, n18443, n18444, n18445, n18446, n18447, n18448,
         n18449, n18450, n18451, n18452, n18453, n18454, n18455, n18456,
         n18457, n18458, n18459, n18460, n18461, n18462, n18463, n18464,
         n18465, n18466, n18467, n18468, n18469, n18470, n18471, n18472,
         n18473, n18474, n18475, n18476, n18477, n18478, n18479, n18480,
         n18481, n18482, n18483, n18484, n18485, n18486, n18487, n18488,
         n18489, n18490, n18491, n18492, n18493, n18494, n18495, n18496,
         n18497, n18498, n18499, n18500, n18501, n18502, n18503, n18504,
         n18505, n18506, n18507, n18508, n18509, n18510, n18511, n18512,
         n18513, n18514, n18515, n18516, n18517, n18518, n18519, n18520,
         n18521, n18522, n18523, n18524, n18525, n18526, n18527, n18528,
         n18529, n18530, n18531, n18532, n18533, n18534, n18535, n18536,
         n18537, n18538, n18539, n18540, n18541, n18542, n18543, n18544,
         n18545, n18546, n18547, n18548, n18549, n18550, n18551, n18552,
         n18553, n18554, n18555, n18556, n18557, n18558, n18559, n18560,
         n18561, n18562, n18563, n18564, n18565, n18566, n18567, n18568,
         n18569, n18570, n18571, n18572, n18573, n18574, n18575, n18576,
         n18577, n18578, n18579, n18580, n18581, n18582, n18583, n18584,
         n18585, n18586, n18587, n18588, n18589, n18590, n18591, n18592,
         n18593, n18594, n18595, n18596, n18597, n18598, n18599, n18600,
         n18601, n18602, n18603, n18604, n18605, n18606, n18607, n18608,
         n18609, n18610, n18611, n18612, n18613, n18614, n18615, n18616,
         n18617, n18618, n18619, n18620, n18621, n18622, n18623, n18624,
         n18625, n18626, n18627, n18628, n18629, n18630, n18631, n18632,
         n18633, n18634, n18635, n18636, n18637, n18638, n18639, n18640,
         n18641, n18642, n18643, n18644, n18645, n18646, n18647, n18648,
         n18649, n18650, n18651, n18652, n18653, n18654, n18655, n18656,
         n18657, n18658, n18659, n18660, n18661, n18662, n18663, n18664,
         n18665, n18666, n18667, n18668, n18669, n18670, n18671, n18672,
         n18673, n18674, n18675, n18676, n18677, n18678, n18679, n18680,
         n18681, n18682, n18683, n18684, n18685, n18686, n18687, n18688,
         n18689, n18690, n18691, n18692, n18693, n18694, n18695, n18696,
         n18697, n18698, n18699, n18700, n18701, n18702, n18703, n18704,
         n18705, n18706, n18707, n18708, n18709, n18710, n18711, n18712,
         n18713, n18714, n18715, n18716, n18717, n18718, n18719, n18720,
         n18721, n18722, n18723, n18724, n18725, n18726, n18727, n18728,
         n18729, n18730, n18731, n18732, n18733, n18734, n18735, n18736,
         n18737, n18738, n18739, n18740, n18741, n18742, n18743, n18744,
         n18745, n18746, n18747, n18748, n18749, n18750, n18751, n18752,
         n18753, n18754, n18755, n18756, n18757, n18758, n18759, n18760,
         n18761, n18762, n18763, n18764, n18765, n18766, n18767, n18768,
         n18769, n18770, n18771, n18772, n18773, n18774, n18775, n18776,
         n18777, n18778, n18779, n18780, n18781, n18782, n18783, n18784,
         n18785, n18786, n18787, n18788, n18789, n18790, n18791, n18792,
         n18793, n18794, n18795, n18796, n18797, n18798, n18799, n18800,
         n18801, n18802, n18803, n18804, n18805, n18806, n18807, n18808,
         n18809, n18810, n18811, n18812, n18813, n18814, n18815, n18816,
         n18817, n18818, n18819, n18820, n18821, n18822, n18823, n18824,
         n18825, n18826, n18827, n18828, n18829, n18830, n18831, n18832,
         n18833, n18834, n18835, n18836, n18837, n18838, n18839, n18840,
         n18841, n18842, n18843, n18844, n18845, n18846, n18847, n18848,
         n18849, n18850, n18851, n18852, n18853, n18854, n18855, n18856,
         n18857, n18858, n18859, n18860, n18861, n18862, n18863, n18864,
         n18865, n18866, n18867, n18868, n18869, n18870, n18871, n18872,
         n18873, n18874, n18875, n18876, n18877, n18878, n18879, n18880,
         n18881, n18882, n18883, n18884, n18885, n18886, n18887, n18888,
         n18889, n18890, n18891, n18892, n18893, n18894, n18895, n18896,
         n18897, n18898, n18899, n18900, n18901, n18902, n18903, n18904,
         n18905, n18906, n18907, n18908, n18909, n18910, n18911, n18912,
         n18913, n18914, n18915, n18916, n18917, n18918, n18919, n18920,
         n18921, n18922, n18923, n18924, n18925, n18926, n18927, n18928,
         n18929, n18930, n18931, n18932, n18933, n18934, n18935, n18936,
         n18937, n18938, n18939, n18940, n18941, n18942, n18943, n18944,
         n18945, n18946, n18947, n18948, n18949, n18950, n18951, n18952,
         n18953, n18954, n18955, n18956, n18957, n18958, n18959, n18960,
         n18961, n18962, n18963, n18964, n18965, n18966, n18967, n18968,
         n18969, n18970, n18971, n18972, n18973, n18974, n18975, n18976,
         n18977, n18978, n18979, n18980, n18981, n18982, n18983, n18984,
         n18985, n18986, n18987, n18988, n18989, n18990, n18991, n18992,
         n18993, n18994, n18995, n18996, n18997, n18998, n18999, n19000,
         n19001, n19002, n19003, n19004, n19005, n19006, n19007, n19008,
         n19009, n19010, n19011, n19012, n19013, n19014, n19015, n19016,
         n19017, n19018, n19019, n19020, n19021, n19022, n19023, n19024,
         n19025, n19026, n19027, n19028, n19029, n19030, n19031, n19032,
         n19033, n19034, n19035, n19036, n19037, n19038, n19039, n19040,
         n19041, n19042, n19043, n19044, n19045, n19046, n19047, n19048,
         n19049, n19050, n19051, n19052, n19053, n19054, n19055, n19056,
         n19057, n19058, n19059, n19060, n19061, n19062, n19063, n19064,
         n19065, n19066, n19067, n19068, n19069, n19070, n19071, n19072,
         n19073, n19074, n19075, n19076, n19077, n19078, n19079, n19080,
         n19081, n19082, n19083, n19084, n19085, n19086, n19087, n19088,
         n19089, n19090, n19091, n19092, n19093, n19094, n19095, n19096,
         n19097, n19098, n19099, n19100, n19101, n19102, n19103, n19104,
         n19105, n19106, n19107, n19108, n19109, n19110, n19111, n19112,
         n19113, n19114, n19115, n19116, n19117, n19118, n19119, n19120,
         n19121, n19122, n19123, n19124, n19125, n19126, n19127, n19128,
         n19129, n19130, n19131, n19132, n19133, n19134, n19135, n19136,
         n19137, n19138, n19139, n19140, n19141, n19142, n19143, n19144,
         n19145, n19146, n19147, n19148, n19149, n19150, n19151, n19152,
         n19153, n19154, n19155, n19156, n19157, n19158, n19159, n19160,
         n19161, n19162, n19163, n19164, n19165, n19166, n19167, n19168,
         n19169, n19170, n19171, n19172, n19173, n19174, n19175, n19176,
         n19177, n19178, n19179, n19180, n19181, n19182, n19183, n19184,
         n19185, n19186, n19187, n19188, n19189, n19190, n19191, n19192,
         n19193, n19194, n19195, n19196, n19197, n19198, n19199, n19200,
         n19201, n19202, n19203, n19204, n19205, n19206, n19207, n19208,
         n19209, n19210, n19211, n19212, n19213, n19214, n19215, n19216,
         n19217, n19218, n19219, n19220, n19221, n19222, n19223, n19224,
         n19225, n19226, n19227, n19228, n19229, n19230, n19231, n19232,
         n19233, n19234, n19235, n19236, n19237, n19238, n19239, n19240,
         n19241, n19242, n19243, n19244, n19245, n19246, n19247, n19248,
         n19249, n19250, n19251, n19252, n19253, n19254, n19255, n19256,
         n19257, n19258, n19259, n19260, n19261, n19262, n19263, n19264,
         n19265, n19266, n19267, n19268, n19269, n19270, n19271, n19272,
         n19273, n19274, n19275, n19276, n19277, n19278, n19279, n19280,
         n19281, n19282, n19283, n19284, n19285, n19286, n19287, n19288,
         n19289, n19290, n19291, n19292, n19293, n19294, n19295, n19296,
         n19297, n19298, n19299, n19300, n19301, n19302, n19303, n19304,
         n19305, n19306, n19307, n19308, n19309, n19310, n19311, n19312,
         n19313, n19314, n19315, n19316, n19317, n19318, n19319, n19320,
         n19321, n19322, n19323, n19324, n19325, n19326, n19327, n19328,
         n19329, n19330, n19331, n19332, n19333, n19334, n19335, n19336,
         n19337, n19338, n19339, n19340, n19341, n19342, n19343, n19344,
         n19345, n19346, n19347, n19348, n19349, n19350, n19351, n19352,
         n19353, n19354, n19355, n19356, n19357, n19358, n19359, n19360,
         n19361, n19362, n19363, n19364, n19365, n19366, n19367, n19368,
         n19369, n19370, n19371, n19372, n19373, n19374, n19375, n19376,
         n19377, n19378, n19379, n19380, n19381, n19382, n19383, n19384,
         n19385, n19386, n19387, n19388, n19389, n19390, n19391, n19392,
         n19393, n19394, n19395, n19396, n19397, n19398, n19399, n19400,
         n19401, n19402, n19403, n19404, n19405, n19406, n19407, n19408,
         n19409, n19410, n19411, n19412, n19413, n19414, n19415, n19416,
         n19417, n19418, n19419, n19420, n19421, n19422, n19423, n19424,
         n19425, n19426, n19427, n19428, n19429, n19430, n19431, n19432,
         n19433, n19434, n19435, n19436, n19437, n19438, n19439, n19440,
         n19441, n19442, n19443, n19444, n19445, n19446, n19447, n19448,
         n19449, n19450, n19451, n19452, n19453, n19454, n19455, n19456,
         n19457, n19458, n19459, n19460, n19461, n19462, n19463, n19464,
         n19465, n19466, n19467, n19468, n19469, n19470, n19471, n19472,
         n19473, n19474, n19475, n19476, n19477, n19478, n19479, n19480,
         n19481, n19482, n19483, n19484, n19485, n19486, n19487, n19488,
         n19489, n19490, n19491, n19492, n19493, n19494, n19495, n19496,
         n19497, n19498, n19499, n19500, n19501, n19502, n19503, n19504,
         n19505, n19506, n19507, n19508, n19509, n19510, n19511, n19512,
         n19513, n19514, n19515, n19516, n19517, n19518, n19519, n19520,
         n19521, n19522, n19523, n19524, n19525, n19526, n19527, n19528,
         n19529, n19530, n19531, n19532, n19533, n19534, n19535, n19536,
         n19537, n19538, n19539, n19540, n19541, n19542, n19543, n19544,
         n19545, n19546, n19547, n19548, n19549, n19550, n19551, n19552,
         n19553, n19554, n19555, n19556, n19557, n19558, n19559, n19560,
         n19561, n19562, n19563, n19564, n19565, n19566, n19567, n19568,
         n19569, n19570, n19571, n19572, n19573, n19574, n19575, n19576,
         n19577, n19578, n19579, n19580, n19581, n19582, n19583, n19584,
         n19585, n19586, n19587, n19588, n19589, n19590, n19591, n19592,
         n19593, n19594, n19595, n19596, n19597, n19598, n19599, n19600,
         n19601, n19602, n19603, n19604, n19605, n19606, n19607, n19608,
         n19609, n19610, n19611, n19612, n19613, n19614, n19615, n19616,
         n19617, n19618, n19619, n19620, n19621, n19622, n19623, n19624,
         n19625, n19626, n19627, n19628, n19629, n19630, n19631, n19632,
         n19633, n19634, n19635, n19636, n19637, n19638, n19639, n19640,
         n19641, n19642, n19643, n19644, n19645, n19646, n19647, n19648,
         n19649, n19650, n19651, n19652, n19653, n19654, n19655, n19656,
         n19657, n19658, n19659, n19660, n19661, n19662, n19663, n19664,
         n19665, n19666, n19667, n19668, n19669, n19670, n19671, n19672,
         n19673, n19674, n19675, n19676, n19677, n19678, n19679, n19680,
         n19681, n19682, n19683, n19684, n19685, n19686, n19687, n19688,
         n19689, n19690, n19691, n19692, n19693, n19694, n19695, n19696,
         n19697, n19698, n19699, n19700, n19701, n19702, n19703, n19704,
         n19705, n19706, n19707, n19708, n19709, n19710, n19711, n19712,
         n19713, n19714, n19715, n19716, n19717, n19718, n19719, n19720,
         n19721, n19722, n19723, n19724, n19725, n19726, n19727, n19728,
         n19729, n19730, n19731, n19732, n19733, n19734, n19735, n19736,
         n19737, n19738, n19739, n19740, n19741, n19742, n19743, n19744,
         n19745, n19746, n19747, n19748, n19749, n19750, n19751, n19752,
         n19753, n19754, n19755, n19756, n19757, n19758, n19759, n19760,
         n19761, n19762, n19763, n19764, n19765, n19766, n19767, n19768,
         n19769, n19770, n19771, n19772, n19773, n19774, n19775, n19776,
         n19777, n19778, n19779, n19780, n19781, n19782, n19783, n19784,
         n19785, n19786, n19787, n19788, n19789, n19790, n19791, n19792,
         n19793, n19794, n19795, n19796, n19797, n19798, n19799, n19800,
         n19801, n19802, n19803, n19804, n19805, n19806, n19807, n19808,
         n19809, n19810, n19811, n19812, n19813, n19814, n19815, n19816,
         n19817, n19818, n19819, n19820, n19821, n19822, n19823, n19824,
         n19825, n19826, n19827, n19828, n19829, n19830, n19831, n19832,
         n19833, n19834, n19835, n19836, n19837, n19838, n19839, n19840,
         n19841, n19842, n19843, n19844, n19845, n19846, n19847, n19848,
         n19849, n19850, n19851, n19852, n19853, n19854, n19855, n19856,
         n19857, n19858, n19859, n19860, n19861, n19862, n19863, n19864,
         n19865, n19866, n19867, n19868, n19869, n19870, n19871, n19872,
         n19873, n19874, n19875, n19876, n19877, n19878, n19879, n19880,
         n19881, n19882, n19883, n19884, n19885, n19886, n19887, n19888,
         n19889, n19890, n19891, n19892, n19893, n19894, n19895, n19896,
         n19897, n19898, n19899, n19900, n19901, n19902, n19903, n19904,
         n19905, n19906, n19907, n19908, n19909, n19910, n19911, n19912,
         n19913, n19914, n19915, n19916, n19917, n19918, n19919, n19920,
         n19921, n19922, n19923, n19924, n19925, n19926, n19927, n19928,
         n19929, n19930, n19931, n19932, n19933, n19934, n19935, n19936,
         n19937, n19938, n19939, n19940, n19941, n19942, n19943, n19944,
         n19945, n19946, n19947, n19948, n19949, n19950, n19951, n19952,
         n19953, n19954, n19955, n19956, n19957, n19958, n19959, n19960,
         n19961, n19962, n19963, n19964, n19965, n19966, n19967, n19968,
         n19969, n19970, n19971, n19972, n19973, n19974, n19975, n19976,
         n19977, n19978, n19979, n19980, n19981, n19982, n19983, n19984,
         n19985, n19986, n19987, n19988, n19989, n19990, n19991, n19992,
         n19993, n19994, n19995, n19996, n19997, n19998, n19999, n20000,
         n20001, n20002, n20003, n20004, n20005, n20006, n20007, n20008,
         n20009, n20010, n20011, n20012, n20013, n20014, n20015, n20016,
         n20017, n20018, n20019, n20020, n20021, n20022, n20023, n20024,
         n20025, n20026, n20027, n20028, n20029, n20030, n20031, n20032,
         n20033, n20034, n20035, n20036, n20037, n20038, n20039, n20040,
         n20041, n20042, n20043, n20044, n20045, n20046, n20047, n20048,
         n20049, n20050, n20051, n20052, n20053, n20054, n20055, n20056,
         n20057, n20058, n20059, n20060, n20061, n20062, n20063, n20064,
         n20065, n20066, n20067, n20068, n20069, n20070, n20071, n20072,
         n20073, n20074, n20075, n20076, n20077, n20078, n20079, n20080,
         n20081, n20082, n20083, n20084, n20085, n20086, n20087, n20088,
         n20089, n20090, n20091, n20092, n20093, n20094, n20095, n20096,
         n20097, n20098, n20099, n20100, n20101, n20102, n20103, n20104,
         n20105, n20106, n20107, n20108, n20109, n20110, n20111, n20112,
         n20113, n20114, n20115, n20116, n20117, n20118, n20119, n20120,
         n20121, n20122, n20123, n20124, n20125, n20126, n20127, n20128,
         n20129, n20130, n20131, n20132, n20133, n20134, n20135, n20136,
         n20137, n20138, n20139, n20140, n20141, n20142, n20143, n20144,
         n20145, n20146, n20147, n20148, n20149, n20150, n20151, n20152,
         n20153, n20154, n20155, n20156, n20157, n20158, n20159, n20160,
         n20161, n20162, n20163, n20164, n20165, n20166, n20167, n20168,
         n20169, n20170, n20171, n20172, n20173, n20174, n20175, n20176,
         n20177, n20178, n20179, n20180, n20181, n20182, n20183, n20184,
         n20185, n20186, n20187, n20188, n20189, n20190, n20191, n20192,
         n20193, n20194, n20195, n20196, n20197, n20198, n20199, n20200,
         n20201, n20202, n20203, n20204, n20205, n20206, n20207, n20208,
         n20209, n20210, n20211, n20212, n20213, n20214, n20215, n20216,
         n20217, n20218, n20219, n20220, n20221, n20222, n20223, n20224,
         n20225, n20226, n20227, n20228, n20229, n20230, n20231, n20232,
         n20233, n20234, n20235, n20236, n20237, n20238, n20239, n20240,
         n20241, n20242, n20243, n20244, n20245, n20246, n20247, n20248,
         n20249, n20250, n20251, n20252, n20253, n20254, n20255, n20256,
         n20257, n20258, n20259, n20260, n20261, n20262, n20263, n20264,
         n20265, n20266, n20267, n20268, n20269, n20270, n20271, n20272,
         n20273, n20274, n20275, n20276, n20277, n20278, n20279, n20280,
         n20281, n20282, n20283, n20284, n20285, n20286, n20287, n20288,
         n20289, n20290, n20291, n20292, n20293, n20294, n20295, n20296,
         n20297, n20298, n20299, n20300, n20301, n20302, n20303, n20304,
         n20305, n20306, n20307, n20308, n20309, n20310, n20311, n20312,
         n20313, n20314, n20315, n20316, n20317, n20318, n20319, n20320,
         n20321, n20322, n20323, n20324, n20325, n20326, n20327, n20328,
         n20329, n20330, n20331, n20332, n20333, n20334, n20335, n20336,
         n20337, n20338, n20339, n20340, n20341, n20342, n20343, n20344,
         n20345, n20346, n20347, n20348, n20349, n20350, n20351, n20352,
         n20353, n20354, n20355, n20356, n20357, n20358, n20359, n20360,
         n20361, n20362, n20363, n20364, n20365, n20366, n20367, n20368,
         n20369, n20370, n20371, n20372, n20373, n20374, n20375, n20376,
         n20377, n20378, n20379, n20380, n20381, n20382, n20383, n20384,
         n20385, n20386, n20387, n20388, n20389, n20390, n20391, n20392,
         n20393, n20394, n20395, n20396, n20397, n20398, n20399, n20400,
         n20401, n20402, n20403, n20404, n20405, n20406, n20407, n20408,
         n20409, n20410, n20411, n20412, n20413, n20414, n20415, n20416,
         n20417, n20418, n20419, n20420, n20421, n20422, n20423, n20424,
         n20425, n20426, n20427, n20428, n20429, n20430, n20431, n20432,
         n20433, n20434, n20435, n20436, n20437, n20438, n20439, n20440,
         n20441, n20442, n20443, n20444, n20445, n20446, n20447, n20448,
         n20449, n20450, n20451, n20452, n20453, n20454, n20455, n20456,
         n20457, n20458, n20459, n20460, n20461, n20462, n20463, n20464,
         n20465, n20466, n20467, n20468, n20469, n20470, n20471, n20472,
         n20473, n20474, n20475, n20476, n20477, n20478, n20479, n20480,
         n20481, n20482, n20483, n20484, n20485, n20486, n20487, n20488,
         n20489, n20490, n20491, n20492, n20493, n20494, n20495, n20496,
         n20497, n20498, n20499, n20500, n20501, n20502, n20503, n20504,
         n20505, n20506, n20507, n20508, n20509, n20510, n20511, n20512,
         n20513, n20514, n20515, n20516, n20517, n20518, n20519, n20520,
         n20521, n20522, n20523, n20524, n20525, n20526, n20527, n20528,
         n20529, n20530, n20531, n20532, n20533, n20534, n20535, n20536,
         n20537, n20538, n20539, n20540, n20541, n20542, n20543, n20544,
         n20545, n20546, n20547, n20548, n20549, n20550, n20551, n20552,
         n20553, n20554, n20555, n20556, n20557, n20558, n20559, n20560,
         n20561, n20562, n20563, n20564, n20565, n20566, n20567, n20568,
         n20569, n20570, n20571, n20572, n20573, n20574, n20575, n20576,
         n20577, n20578, n20579, n20580, n20581, n20582, n20583, n20584,
         n20585, n20586, n20587, n20588, n20589, n20590, n20591, n20592,
         n20593, n20594, n20595, n20596, n20597, n20598, n20599, n20600,
         n20601, n20602, n20603, n20604, n20605, n20606, n20607, n20608,
         n20609, n20610, n20611, n20612, n20613, n20614, n20615, n20616,
         n20617, n20618, n20619, n20620, n20621, n20622, n20623, n20624,
         n20625, n20626, n20627, n20628, n20629, n20630, n20631, n20632,
         n20633, n20634, n20635, n20636, n20637, n20638, n20639, n20640,
         n20641, n20642, n20643, n20644, n20645, n20646, n20647, n20648,
         n20649, n20650, n20651, n20652, n20653, n20654, n20655, n20656,
         n20657, n20658, n20659, n20660, n20661, n20662, n20663, n20664,
         n20665, n20666, n20667, n20668, n20669, n20670, n20671, n20672,
         n20673, n20674, n20675, n20676, n20677, n20678, n20679, n20680,
         n20681, n20682, n20683, n20684, n20685, n20686, n20687, n20688,
         n20689, n20690, n20691, n20692, n20693, n20694, n20695, n20696,
         n20697, n20698, n20699, n20700, n20701, n20702, n20703, n20704,
         n20705, n20706, n20707, n20708, n20709, n20710, n20711, n20712,
         n20713, n20714, n20715, n20716, n20717, n20718, n20719, n20720,
         n20721, n20722, n20723, n20724, n20725, n20726, n20727, n20728,
         n20729, n20730, n20731, n20732, n20733, n20734, n20735, n20736,
         n20737, n20738, n20739, n20740, n20741, n20742, n20743, n20744,
         n20745, n20746, n20747, n20748, n20749, n20750, n20751, n20752,
         n20753, n20754, n20755, n20756, n20757, n20758, n20759, n20760,
         n20761, n20762, n20763, n20764, n20765, n20766, n20767, n20768,
         n20769, n20770, n20771, n20772, n20773, n20774, n20775, n20776,
         n20777, n20778, n20779, n20780, n20781, n20782, n20783, n20784,
         n20785, n20786, n20787, n20788, n20789, n20790, n20791, n20792,
         n20793, n20794, n20795, n20796, n20797, n20798, n20799, n20800,
         n20801, n20802, n20803, n20804, n20805, n20806, n20807, n20808,
         n20809, n20810, n20811, n20812, n20813, n20814, n20815, n20816,
         n20817, n20818, n20819, n20820, n20821, n20822, n20823, n20824,
         n20825, n20826, n20827, n20828, n20829, n20830, n20831, n20832,
         n20833, n20834, n20835, n20836, n20837, n20838, n20839, n20840,
         n20841, n20842, n20843, n20844, n20845, n20846, n20847, n20848,
         n20849, n20850, n20851, n20852, n20853, n20854, n20855, n20856,
         n20857, n20858, n20859, n20860, n20861, n20862, n20863, n20864,
         n20865, n20866, n20867, n20868, n20869, n20870, n20871, n20872,
         n20873, n20874, n20875, n20876, n20877, n20878, n20879, n20880,
         n20881, n20882, n20883, n20884, n20885, n20886, n20887, n20888,
         n20889, n20890, n20891, n20892, n20893, n20894, n20895, n20896,
         n20897, n20898, n20899, n20900, n20901, n20902, n20903, n20904,
         n20905, n20906, n20907, n20908, n20909, n20910, n20911, n20912,
         n20913, n20914, n20915, n20916, n20917, n20918, n20919, n20920,
         n20921, n20922, n20923, n20924, n20925, n20926, n20927, n20928,
         n20929, n20930, n20931, n20932, n20933, n20934, n20935, n20936,
         n20937;

  AOI211_X1 U11046 ( .C1(n17884), .C2(n17720), .A(n17734), .B(n17719), .ZN(
        n17728) );
  AND2_X1 U11047 ( .A1(n14326), .A2(n14327), .ZN(n14323) );
  NOR2_X1 U11048 ( .A1(n14220), .A2(n14312), .ZN(n11096) );
  INV_X4 U11049 ( .A(n20042), .ZN(n20031) );
  AND2_X1 U11050 ( .A1(n14252), .A2(n9727), .ZN(n14241) );
  AND2_X1 U11051 ( .A1(n15923), .A2(n9887), .ZN(n14589) );
  NOR2_X1 U11053 ( .A1(n13457), .A2(n10472), .ZN(n13580) );
  INV_X2 U11054 ( .A(n18912), .ZN(n9887) );
  XNOR2_X1 U11055 ( .A(n12205), .B(n14055), .ZN(n13833) );
  OAI211_X1 U11056 ( .C1(n15084), .C2(n15083), .A(n18693), .B(n18482), .ZN(
        n15431) );
  NAND2_X1 U11057 ( .A1(n10353), .A2(n10352), .ZN(n10400) );
  XNOR2_X1 U11058 ( .A(n9812), .B(n10299), .ZN(n10353) );
  NOR2_X1 U11060 ( .A1(n11242), .A2(n11243), .ZN(n11217) );
  OAI21_X2 U11061 ( .B1(n18925), .B2(n12529), .A(n12528), .ZN(n15038) );
  NAND2_X1 U11062 ( .A1(n12060), .A2(n12032), .ZN(n12132) );
  OR2_X2 U11063 ( .A1(n12053), .A2(n12058), .ZN(n19339) );
  AND2_X1 U11064 ( .A1(n13040), .A2(n13039), .ZN(n11683) );
  INV_X1 U11065 ( .A(n15174), .ZN(n16994) );
  NOR2_X1 U11066 ( .A1(n11228), .A2(n18834), .ZN(n11229) );
  CLKBUF_X1 U11067 ( .A(n15173), .Z(n16996) );
  INV_X2 U11068 ( .A(n16777), .ZN(n17023) );
  CLKBUF_X1 U11069 ( .A(n10250), .Z(n13384) );
  INV_X2 U11070 ( .A(n16824), .ZN(n16995) );
  CLKBUF_X2 U11071 ( .A(n10187), .Z(n10484) );
  CLKBUF_X2 U11072 ( .A(n10490), .Z(n10768) );
  CLKBUF_X2 U11073 ( .A(n10291), .Z(n11041) );
  INV_X1 U11074 ( .A(n15343), .ZN(n10249) );
  BUF_X2 U11075 ( .A(n9627), .Z(n16974) );
  INV_X2 U11076 ( .A(n15148), .ZN(n16997) );
  AND2_X1 U11077 ( .A1(n9639), .A2(n9631), .ZN(n12865) );
  NAND2_X1 U11078 ( .A1(n20086), .A2(n20096), .ZN(n15343) );
  BUF_X1 U11079 ( .A(n11742), .Z(n12662) );
  AND2_X1 U11080 ( .A1(n9643), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11694) );
  AND2_X1 U11081 ( .A1(n12690), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11740) );
  INV_X1 U11082 ( .A(n13410), .ZN(n20107) );
  INV_X1 U11083 ( .A(n13389), .ZN(n13172) );
  NAND2_X1 U11084 ( .A1(n12841), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11687) );
  NAND2_X1 U11085 ( .A1(n9642), .A2(n11278), .ZN(n11686) );
  NOR2_X2 U11086 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n15090), .ZN(
        n15174) );
  AND2_X4 U11087 ( .A1(n10142), .A2(n10143), .ZN(n10213) );
  CLKBUF_X2 U11088 ( .A(n17024), .Z(n9627) );
  CLKBUF_X2 U11089 ( .A(n17019), .Z(n9626) );
  CLKBUF_X2 U11090 ( .A(n10207), .Z(n9621) );
  CLKBUF_X2 U11091 ( .A(n10207), .Z(n9620) );
  CLKBUF_X2 U11092 ( .A(n10207), .Z(n9622) );
  INV_X1 U11093 ( .A(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n18647) );
  AND2_X1 U11095 ( .A1(n10038), .A2(n10141), .ZN(n10291) );
  BUF_X1 U11096 ( .A(n10483), .Z(n10458) );
  CLKBUF_X1 U11097 ( .A(n10491), .Z(n10998) );
  AND2_X1 U11098 ( .A1(n11403), .A2(n13152), .ZN(n11459) );
  AND2_X1 U11099 ( .A1(n11454), .A2(n12452), .ZN(n12449) );
  INV_X2 U11100 ( .A(n19796), .ZN(n12068) );
  NAND2_X1 U11101 ( .A1(n11390), .A2(n11389), .ZN(n11458) );
  INV_X1 U11102 ( .A(n12374), .ZN(n11390) );
  INV_X1 U11103 ( .A(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10132) );
  AND3_X1 U11104 ( .A1(n9692), .A2(n11630), .A3(n11450), .ZN(n11454) );
  NAND2_X1 U11105 ( .A1(n11388), .A2(n11387), .ZN(n13728) );
  CLKBUF_X2 U11106 ( .A(n11400), .Z(n11630) );
  AND2_X1 U11107 ( .A1(n11420), .A2(n11640), .ZN(n12375) );
  NAND2_X1 U11108 ( .A1(n11434), .A2(n11640), .ZN(n11470) );
  INV_X1 U11109 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11278) );
  AND2_X4 U11110 ( .A1(n11260), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11281) );
  INV_X1 U11111 ( .A(n11280), .ZN(n9644) );
  INV_X1 U11112 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n11258) );
  AND2_X2 U11113 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n11259) );
  AND2_X1 U11114 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n11650) );
  CLKBUF_X1 U11115 ( .A(n18472), .Z(n9602) );
  NOR2_X1 U11116 ( .A1(n18518), .A2(n18360), .ZN(n18472) );
  OAI21_X2 U11117 ( .B1(n14186), .B2(P2_STATE2_REG_0__SCAN_IN), .A(n12471), 
        .ZN(n18831) );
  AOI21_X4 U11118 ( .B1(n15431), .B2(n15430), .A(n18534), .ZN(n17186) );
  OR2_X2 U11119 ( .A1(n13853), .A2(n13859), .ZN(n15090) );
  NOR2_X1 U11120 ( .A1(n10251), .A2(n13394), .ZN(n10252) );
  NOR2_X2 U11121 ( .A1(n17875), .A2(n17861), .ZN(n17887) );
  NAND2_X2 U11122 ( .A1(n11166), .A2(n15655), .ZN(n15650) );
  NAND2_X2 U11123 ( .A1(n9871), .A2(n12281), .ZN(n14906) );
  OR2_X4 U11124 ( .A1(n12056), .A2(n12058), .ZN(n12122) );
  INV_X1 U11125 ( .A(n9745), .ZN(n9603) );
  AND2_X1 U11126 ( .A1(n9604), .A2(n13781), .ZN(n14271) );
  NOR2_X1 U11127 ( .A1(n10646), .A2(n9603), .ZN(n9604) );
  NOR2_X1 U11128 ( .A1(n13767), .A2(n13783), .ZN(n9605) );
  NOR2_X1 U11129 ( .A1(n11198), .A2(n13410), .ZN(n9606) );
  NOR2_X1 U11130 ( .A1(n13767), .A2(n13783), .ZN(n13781) );
  NAND2_X1 U11131 ( .A1(n10520), .A2(n10519), .ZN(n13767) );
  NOR2_X1 U11132 ( .A1(n11198), .A2(n13410), .ZN(n10253) );
  AND2_X2 U11133 ( .A1(n12441), .A2(n11980), .ZN(n14806) );
  NAND2_X1 U11134 ( .A1(n11465), .A2(n11464), .ZN(n9607) );
  CLKBUF_X1 U11136 ( .A(n14622), .Z(n9609) );
  BUF_X1 U11137 ( .A(n14605), .Z(n9610) );
  CLKBUF_X1 U11138 ( .A(n14624), .Z(n9611) );
  NAND2_X1 U11139 ( .A1(n11465), .A2(n11464), .ZN(n11491) );
  NAND2_X1 U11140 ( .A1(n14622), .A2(n12753), .ZN(n12773) );
  AND2_X1 U11142 ( .A1(n12688), .A2(n11644), .ZN(n9670) );
  OR2_X1 U11143 ( .A1(n11664), .A2(n11663), .ZN(n12399) );
  AND2_X2 U11144 ( .A1(n11259), .A2(n11612), .ZN(n11656) );
  AND2_X1 U11145 ( .A1(n13167), .A2(n10140), .ZN(n10485) );
  AND2_X1 U11146 ( .A1(n12688), .A2(n11645), .ZN(n9652) );
  BUF_X1 U11147 ( .A(n11492), .Z(n11606) );
  INV_X2 U11148 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n13620) );
  NOR2_X1 U11149 ( .A1(n10474), .A2(n10473), .ZN(n11157) );
  AND2_X1 U11150 ( .A1(n14367), .A2(n10256), .ZN(n11154) );
  INV_X1 U11151 ( .A(n11606), .ZN(n12472) );
  INV_X1 U11152 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n11612) );
  NAND2_X1 U11153 ( .A1(n11458), .A2(n11459), .ZN(n13606) );
  AND2_X1 U11154 ( .A1(n12371), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n13591) );
  INV_X1 U11155 ( .A(n16958), .ZN(n14010) );
  NAND2_X2 U11156 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n13859) );
  INV_X2 U11157 ( .A(n20096), .ZN(n10256) );
  AND3_X1 U11158 ( .A1(n9888), .A2(n9887), .A3(n9889), .ZN(n18737) );
  OAI21_X1 U11159 ( .B1(n18912), .B2(n18765), .A(n18764), .ZN(n14072) );
  AND2_X2 U11160 ( .A1(n13711), .A2(n13740), .ZN(n13739) );
  INV_X2 U11161 ( .A(n11558), .ZN(n11592) );
  NAND2_X1 U11162 ( .A1(n12149), .A2(n18907), .ZN(n12167) );
  NAND2_X2 U11163 ( .A1(n11322), .A2(n11321), .ZN(n11450) );
  CLKBUF_X2 U11164 ( .A(n13881), .Z(n16977) );
  INV_X1 U11165 ( .A(n18692), .ZN(n17291) );
  OR2_X1 U11166 ( .A1(n15205), .A2(n17840), .ZN(n9982) );
  INV_X1 U11167 ( .A(n19867), .ZN(n19929) );
  NAND2_X1 U11168 ( .A1(n14363), .A2(n10939), .ZN(n14353) );
  INV_X1 U11169 ( .A(P2_STATE2_REG_3__SCAN_IN), .ZN(n19594) );
  XNOR2_X1 U11170 ( .A(n12167), .B(n12418), .ZN(n13673) );
  INV_X1 U11171 ( .A(n19934), .ZN(n19897) );
  INV_X2 U11172 ( .A(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n9779) );
  AND4_X1 U11173 ( .A1(n10108), .A2(n15133), .A3(n10116), .A4(n15132), .ZN(
        n9612) );
  NOR2_X1 U11174 ( .A1(n13858), .A2(n18504), .ZN(n13926) );
  AND4_X1 U11175 ( .A1(n10155), .A2(n10154), .A3(n10153), .A4(n10152), .ZN(
        n9613) );
  INV_X1 U11176 ( .A(n11021), .ZN(n9614) );
  NAND2_X2 U11177 ( .A1(n11362), .A2(n11361), .ZN(n11434) );
  OR2_X2 U11178 ( .A1(n11801), .A2(n11800), .ZN(n12322) );
  OAI21_X2 U11179 ( .B1(n13024), .B2(n19807), .A(n13347), .ZN(n13250) );
  NOR2_X2 U11180 ( .A1(n14468), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n14476) );
  INV_X2 U11182 ( .A(n9614), .ZN(n9616) );
  INV_X1 U11183 ( .A(n9614), .ZN(n9617) );
  INV_X1 U11184 ( .A(n9614), .ZN(n9618) );
  INV_X1 U11185 ( .A(n9614), .ZN(n9619) );
  AND2_X1 U11186 ( .A1(n10139), .A2(n13167), .ZN(n11021) );
  NOR2_X2 U11187 ( .A1(n17524), .A2(n15204), .ZN(n15205) );
  CLKBUF_X3 U11188 ( .A(n11449), .Z(n9639) );
  NAND2_X2 U11189 ( .A1(n12027), .A2(n12026), .ZN(n18925) );
  NAND2_X2 U11190 ( .A1(n9755), .A2(n9754), .ZN(n12498) );
  BUF_X4 U11191 ( .A(n10491), .Z(n10972) );
  OR2_X2 U11192 ( .A1(n12542), .A2(n12517), .ZN(n12518) );
  NAND2_X2 U11193 ( .A1(n12516), .A2(n12515), .ZN(n12542) );
  NAND2_X2 U11194 ( .A1(n12150), .A2(n12151), .ZN(n12411) );
  AND2_X1 U11195 ( .A1(n12845), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n9623) );
  AND2_X4 U11196 ( .A1(n13593), .A2(n11278), .ZN(n12671) );
  AND2_X4 U11197 ( .A1(n13082), .A2(n12550), .ZN(n13516) );
  OR2_X2 U11199 ( .A1(n12056), .A2(n12055), .ZN(n12128) );
  CLKBUF_X1 U11200 ( .A(n10492), .Z(n9624) );
  CLKBUF_X1 U11201 ( .A(n10492), .Z(n9625) );
  AND2_X1 U11202 ( .A1(n13164), .A2(n10139), .ZN(n10492) );
  AND2_X1 U11203 ( .A1(n13167), .A2(n10142), .ZN(n10207) );
  XNOR2_X2 U11204 ( .A(n15195), .B(n15194), .ZN(n17650) );
  NOR2_X2 U11205 ( .A1(n9985), .A2(n9986), .ZN(n15195) );
  AND2_X1 U11206 ( .A1(n10038), .A2(n13164), .ZN(n10490) );
  NOR2_X2 U11207 ( .A1(n17650), .A2(n17969), .ZN(n17649) );
  NAND2_X2 U11208 ( .A1(n12031), .A2(n12030), .ZN(n12129) );
  NAND2_X2 U11209 ( .A1(n14600), .A2(n12797), .ZN(n14607) );
  NAND2_X2 U11210 ( .A1(n12794), .A2(n12793), .ZN(n14600) );
  NAND2_X2 U11211 ( .A1(n13076), .A2(n13077), .ZN(n13078) );
  NOR2_X4 U11212 ( .A1(n12944), .A2(n14821), .ZN(n14700) );
  NOR2_X1 U11213 ( .A1(n13861), .A2(n18504), .ZN(n17019) );
  NOR2_X2 U11214 ( .A1(n13862), .A2(n16741), .ZN(n15173) );
  NOR2_X4 U11215 ( .A1(n16741), .A2(n13859), .ZN(n16924) );
  NAND2_X2 U11216 ( .A1(n18668), .A2(n13853), .ZN(n16741) );
  OAI21_X2 U11217 ( .B1(n14605), .B2(n12813), .A(n14601), .ZN(n14595) );
  NOR2_X1 U11218 ( .A1(n13862), .A2(n13860), .ZN(n17024) );
  CLKBUF_X1 U11219 ( .A(n14241), .Z(n14242) );
  OR2_X1 U11220 ( .A1(n11196), .A2(n15558), .ZN(n14460) );
  AND2_X1 U11221 ( .A1(n14653), .A2(n12949), .ZN(n14573) );
  NAND2_X1 U11222 ( .A1(n15212), .A2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n16215) );
  NAND3_X1 U11223 ( .A1(n9801), .A2(n9800), .A3(n11175), .ZN(n15639) );
  INV_X1 U11224 ( .A(n15621), .ZN(n15620) );
  INV_X1 U11225 ( .A(n11173), .ZN(n15621) );
  OAI21_X1 U11227 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(n18685), .A(n16349), 
        .ZN(n17707) );
  NOR2_X2 U11228 ( .A1(n17291), .A2(n16349), .ZN(n17697) );
  NAND2_X1 U11229 ( .A1(n18692), .A2(n17947), .ZN(n18486) );
  NOR2_X2 U11230 ( .A1(n17919), .A2(n18510), .ZN(n17947) );
  OAI211_X1 U11231 ( .C1(n10282), .C2(n13329), .A(n10284), .B(n10283), .ZN(
        n10285) );
  NOR2_X2 U11232 ( .A1(n15231), .A2(n15239), .ZN(n18512) );
  NAND2_X1 U11233 ( .A1(n15081), .A2(n18484), .ZN(n15239) );
  OR2_X1 U11234 ( .A1(n17677), .A2(n17678), .ZN(n9987) );
  AND2_X1 U11235 ( .A1(n11067), .A2(n10247), .ZN(n13397) );
  NAND2_X1 U11236 ( .A1(n9696), .A2(n9659), .ZN(n9795) );
  INV_X4 U11237 ( .A(n12475), .ZN(n11558) );
  NAND2_X1 U11238 ( .A1(n12865), .A2(n13044), .ZN(n11974) );
  XOR2_X1 U11239 ( .A(n17205), .B(n15191), .Z(n15192) );
  NAND2_X1 U11240 ( .A1(n10253), .A2(n10246), .ZN(n13185) );
  NAND3_X1 U11241 ( .A1(n13404), .A2(n14298), .A3(n13177), .ZN(n10267) );
  BUF_X1 U11242 ( .A(n10254), .Z(n13490) );
  NOR2_X1 U11243 ( .A1(n17699), .A2(n17705), .ZN(n17698) );
  NAND2_X1 U11244 ( .A1(n11404), .A2(n11991), .ZN(n12861) );
  INV_X2 U11245 ( .A(n12003), .ZN(n12327) );
  BUF_X2 U11246 ( .A(n11640), .Z(n12003) );
  XNOR2_X1 U11247 ( .A(n15248), .B(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n17699) );
  AND2_X1 U11248 ( .A1(n11434), .A2(n11401), .ZN(n12376) );
  INV_X2 U11249 ( .A(n17220), .ZN(n15248) );
  INV_X1 U11250 ( .A(n10832), .ZN(n10248) );
  NAND2_X1 U11251 ( .A1(n9815), .A2(n9680), .ZN(n10869) );
  AND4_X1 U11252 ( .A1(n10159), .A2(n10158), .A3(n10157), .A4(n10156), .ZN(
        n10131) );
  OR2_X1 U11253 ( .A1(n11266), .A2(n11265), .ZN(n11406) );
  CLKBUF_X2 U11254 ( .A(n15173), .Z(n15158) );
  CLKBUF_X2 U11255 ( .A(n10227), .Z(n10682) );
  AND2_X1 U11256 ( .A1(n13164), .A2(n10142), .ZN(n10290) );
  BUF_X4 U11257 ( .A(n10319), .Z(n9628) );
  AND2_X2 U11258 ( .A1(n11650), .A2(n11258), .ZN(n12845) );
  AND2_X2 U11259 ( .A1(n9779), .A2(n9778), .ZN(n10038) );
  NOR2_X2 U11260 ( .A1(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n12688) );
  AND3_X1 U11261 ( .A1(n10102), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A3(
        n12935), .ZN(n14706) );
  AND2_X1 U11262 ( .A1(n12965), .A2(n12964), .ZN(n12966) );
  NAND2_X1 U11263 ( .A1(n16018), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n16017) );
  NOR2_X1 U11264 ( .A1(n16039), .A2(n16084), .ZN(n16018) );
  AOI21_X1 U11265 ( .B1(n14731), .B2(n16009), .A(n14730), .ZN(n15294) );
  OAI21_X1 U11266 ( .B1(n14726), .B2(n9844), .A(n9842), .ZN(n16011) );
  OAI21_X1 U11267 ( .B1(n14467), .B2(n20070), .A(n9817), .ZN(n9816) );
  AOI21_X1 U11268 ( .B1(n14198), .B2(n11098), .A(n14197), .ZN(n14450) );
  XNOR2_X1 U11269 ( .A(n14461), .B(n11193), .ZN(n14467) );
  AND2_X1 U11270 ( .A1(n14222), .A2(n10824), .ZN(n15572) );
  XNOR2_X1 U11271 ( .A(n9929), .B(n9928), .ZN(n12918) );
  NOR2_X1 U11272 ( .A1(n9922), .A2(n9921), .ZN(n9920) );
  AOI21_X1 U11273 ( .B1(n14223), .B2(n14222), .A(n14221), .ZN(n14465) );
  MUX2_X1 U11274 ( .A(n14460), .B(n14459), .S(n15640), .Z(n14461) );
  NOR2_X1 U11275 ( .A1(n14619), .A2(n14618), .ZN(n14617) );
  XNOR2_X1 U11276 ( .A(n12773), .B(n10101), .ZN(n14619) );
  NAND2_X1 U11277 ( .A1(n14323), .A2(n14324), .ZN(n10822) );
  AOI21_X1 U11278 ( .B1(n18959), .B2(n19122), .A(n12468), .ZN(n12495) );
  AND2_X1 U11279 ( .A1(n12921), .A2(n12920), .ZN(n14447) );
  XNOR2_X1 U11280 ( .A(n12441), .B(n12440), .ZN(n18959) );
  INV_X1 U11281 ( .A(n10050), .ZN(n10049) );
  NAND2_X1 U11282 ( .A1(n14571), .A2(n9924), .ZN(n14815) );
  XNOR2_X1 U11283 ( .A(n12505), .B(n12469), .ZN(n14809) );
  NAND2_X1 U11284 ( .A1(n12752), .A2(n12747), .ZN(n12753) );
  NOR2_X1 U11285 ( .A1(n12945), .A2(n12506), .ZN(n12505) );
  NAND2_X1 U11286 ( .A1(n13683), .A2(n13684), .ZN(n13682) );
  NAND2_X1 U11287 ( .A1(n17344), .A2(n16218), .ZN(n17343) );
  AOI21_X1 U11288 ( .B1(n15599), .B2(n15640), .A(n9695), .ZN(n9811) );
  INV_X1 U11289 ( .A(n12420), .ZN(n9629) );
  OR2_X1 U11290 ( .A1(n12977), .A2(n12978), .ZN(n14632) );
  NAND2_X1 U11291 ( .A1(n12419), .A2(n12418), .ZN(n13684) );
  NOR2_X1 U11292 ( .A1(n16215), .A2(n9976), .ZN(n16165) );
  NOR2_X1 U11293 ( .A1(n14059), .A2(n14060), .ZN(n9943) );
  AND2_X2 U11294 ( .A1(n13739), .A2(n10025), .ZN(n9735) );
  AND2_X1 U11295 ( .A1(n12196), .A2(n12195), .ZN(n12199) );
  AND2_X1 U11296 ( .A1(n12144), .A2(n12143), .ZN(n12198) );
  AND2_X2 U11297 ( .A1(n13516), .A2(n10015), .ZN(n13711) );
  NAND2_X1 U11298 ( .A1(n10037), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n10036) );
  NOR2_X1 U11299 ( .A1(n14533), .A2(n14534), .ZN(n9818) );
  NAND2_X1 U11300 ( .A1(n13360), .A2(n14171), .ZN(n14172) );
  NAND2_X1 U11301 ( .A1(n15616), .A2(n9686), .ZN(n14534) );
  NAND2_X1 U11302 ( .A1(n15621), .A2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n15616) );
  NAND2_X1 U11303 ( .A1(n15922), .A2(n15976), .ZN(n15923) );
  NAND2_X1 U11304 ( .A1(n15640), .A2(n10034), .ZN(n10032) );
  OAI22_X1 U11305 ( .A1(n12091), .A2(n12113), .B1(n12114), .B2(n12090), .ZN(
        n12094) );
  AND2_X1 U11306 ( .A1(n11173), .A2(n15803), .ZN(n14533) );
  NAND2_X1 U11307 ( .A1(n10471), .A2(n10470), .ZN(n13749) );
  OAI21_X1 U11308 ( .B1(n11142), .B2(n10580), .A(n10433), .ZN(n13373) );
  NAND2_X1 U11309 ( .A1(n12045), .A2(n12044), .ZN(n12114) );
  OAI21_X1 U11310 ( .B1(n20683), .B2(n10580), .A(n10409), .ZN(n13338) );
  OR2_X2 U11311 ( .A1(n11157), .A2(n11102), .ZN(n11173) );
  OR2_X1 U11312 ( .A1(n12057), .A2(n12043), .ZN(n19425) );
  OR2_X2 U11313 ( .A1(n12047), .A2(n12058), .ZN(n9673) );
  OR2_X1 U11314 ( .A1(n12057), .A2(n12052), .ZN(n12108) );
  NOR2_X1 U11315 ( .A1(n9819), .A2(n10400), .ZN(n10466) );
  NAND2_X1 U11316 ( .A1(n9821), .A2(n9820), .ZN(n10474) );
  NOR2_X1 U11317 ( .A1(n13086), .A2(n13085), .ZN(n13087) );
  AND2_X1 U11318 ( .A1(n15531), .A2(n10930), .ZN(n14363) );
  NOR4_X2 U11319 ( .A1(n20833), .A2(n17154), .A3(n17243), .A4(n17077), .ZN(
        n17118) );
  NOR2_X2 U11320 ( .A1(n14134), .A2(n10923), .ZN(n15531) );
  AND2_X1 U11321 ( .A1(n10401), .A2(n9822), .ZN(n9821) );
  OR2_X1 U11322 ( .A1(n12526), .A2(n12525), .ZN(n12527) );
  NAND2_X1 U11323 ( .A1(n15544), .A2(n9716), .ZN(n14134) );
  OR2_X1 U11324 ( .A1(n19130), .A2(n16141), .ZN(n12055) );
  NAND2_X1 U11325 ( .A1(n12017), .A2(n12021), .ZN(n19130) );
  OR2_X1 U11326 ( .A1(n14072), .A2(n9743), .ZN(n9888) );
  AND2_X1 U11327 ( .A1(n10399), .A2(n10398), .ZN(n20213) );
  INV_X1 U11328 ( .A(n17701), .ZN(n9647) );
  NAND2_X2 U11329 ( .A1(n12016), .A2(n12015), .ZN(n11503) );
  AND2_X1 U11330 ( .A1(n10351), .A2(n10350), .ZN(n10352) );
  NOR2_X2 U11331 ( .A1(n20118), .A2(n20096), .ZN(n9663) );
  NAND2_X1 U11332 ( .A1(n12397), .A2(n12859), .ZN(n12481) );
  NOR2_X2 U11333 ( .A1(n20107), .A2(n20118), .ZN(n20570) );
  INV_X2 U11334 ( .A(n19941), .ZN(n9630) );
  AND2_X1 U11335 ( .A1(n15850), .A2(n10901), .ZN(n13659) );
  NAND2_X1 U11336 ( .A1(n9970), .A2(n9971), .ZN(n9974) );
  NAND2_X1 U11337 ( .A1(n20180), .A2(n10301), .ZN(n20128) );
  NAND2_X1 U11338 ( .A1(n10302), .A2(n10281), .ZN(n9797) );
  NOR2_X2 U11339 ( .A1(n13454), .A2(n10896), .ZN(n15850) );
  NAND2_X1 U11340 ( .A1(n9825), .A2(n9824), .ZN(n13454) );
  AND2_X1 U11341 ( .A1(n10362), .A2(n10361), .ZN(n10364) );
  AND2_X1 U11342 ( .A1(n11509), .A2(n11508), .ZN(n11514) );
  OR2_X1 U11343 ( .A1(n11711), .A2(n11708), .ZN(n13465) );
  NAND2_X1 U11344 ( .A1(n12992), .A2(n12504), .ZN(n19093) );
  AND2_X1 U11345 ( .A1(n11479), .A2(n9684), .ZN(n11489) );
  NAND2_X1 U11346 ( .A1(n13507), .A2(n13506), .ZN(n13508) );
  XNOR2_X1 U11347 ( .A(n11683), .B(n9919), .ZN(n13507) );
  OR2_X1 U11348 ( .A1(n11683), .A2(n11684), .ZN(n11707) );
  NOR2_X1 U11349 ( .A1(n10372), .A2(n9940), .ZN(n9939) );
  AND2_X1 U11350 ( .A1(n10259), .A2(n10261), .ZN(n10029) );
  INV_X1 U11351 ( .A(n11458), .ZN(n11399) );
  NOR2_X1 U11352 ( .A1(n10347), .A2(n11101), .ZN(n10349) );
  AOI211_X1 U11353 ( .C1(n15222), .C2(n15059), .A(n15058), .B(n15057), .ZN(
        n15074) );
  AND2_X1 U11354 ( .A1(n11682), .A2(n11681), .ZN(n13506) );
  XNOR2_X1 U11355 ( .A(n17980), .B(n15192), .ZN(n17666) );
  INV_X2 U11356 ( .A(n11974), .ZN(n11975) );
  OR2_X1 U11357 ( .A1(n13490), .A2(n10255), .ZN(n13165) );
  NAND2_X1 U11358 ( .A1(n11453), .A2(n12383), .ZN(n12457) );
  OR2_X1 U11359 ( .A1(n18068), .A2(n18076), .ZN(n18495) );
  AND3_X1 U11360 ( .A1(n9691), .A2(n11737), .A3(n10068), .ZN(n12412) );
  NAND2_X4 U11361 ( .A1(n19796), .A2(n11389), .ZN(n11991) );
  XNOR2_X1 U11362 ( .A(n9612), .B(n15248), .ZN(n15185) );
  INV_X1 U11363 ( .A(n11639), .ZN(n11969) );
  INV_X1 U11364 ( .A(n10869), .ZN(n10274) );
  AND2_X1 U11365 ( .A1(n19796), .A2(n19594), .ZN(n11639) );
  NOR2_X1 U11366 ( .A1(n13728), .A2(n18715), .ZN(n12355) );
  AND2_X1 U11367 ( .A1(n11635), .A2(n13728), .ZN(n13063) );
  INV_X1 U11368 ( .A(n17078), .ZN(n18076) );
  INV_X1 U11369 ( .A(n12003), .ZN(n9631) );
  INV_X1 U11370 ( .A(n13728), .ZN(n11389) );
  NOR2_X1 U11371 ( .A1(n18087), .A2(n15076), .ZN(n15236) );
  INV_X1 U11372 ( .A(n17208), .ZN(n15244) );
  OR2_X1 U11373 ( .A1(n10325), .A2(n10324), .ZN(n11170) );
  CLKBUF_X1 U11374 ( .A(n11414), .Z(n13574) );
  INV_X1 U11375 ( .A(n20096), .ZN(n9640) );
  NOR2_X2 U11376 ( .A1(n13878), .A2(n13877), .ZN(n18692) );
  CLKBUF_X1 U11377 ( .A(n10832), .Z(n14367) );
  INV_X2 U11378 ( .A(n16296), .ZN(n16300) );
  NAND4_X1 U11379 ( .A1(n15146), .A2(n15145), .A3(n10113), .A4(n15144), .ZN(
        n17220) );
  INV_X2 U11380 ( .A(U212), .ZN(n16293) );
  AND4_X2 U11381 ( .A1(n10243), .A2(n10240), .A3(n10242), .A4(n10241), .ZN(
        n20096) );
  NAND2_X1 U11382 ( .A1(n11409), .A2(n11278), .ZN(n11277) );
  NAND2_X1 U11383 ( .A1(n11374), .A2(n11373), .ZN(n11401) );
  AND4_X1 U11384 ( .A1(n10235), .A2(n10234), .A3(n10233), .A4(n10232), .ZN(
        n10241) );
  AND4_X1 U11385 ( .A1(n10191), .A2(n10190), .A3(n10189), .A4(n10188), .ZN(
        n9657) );
  AND3_X1 U11386 ( .A1(n10138), .A2(n10136), .A3(n10146), .ZN(n9814) );
  AND4_X1 U11387 ( .A1(n10202), .A2(n10201), .A3(n10200), .A4(n10199), .ZN(
        n10221) );
  AND4_X1 U11388 ( .A1(n10212), .A2(n10211), .A3(n10210), .A4(n10209), .ZN(
        n10219) );
  AND4_X1 U11389 ( .A1(n10163), .A2(n10162), .A3(n10161), .A4(n10160), .ZN(
        n10164) );
  AND4_X1 U11390 ( .A1(n10217), .A2(n10216), .A3(n10215), .A4(n10214), .ZN(
        n10218) );
  AND4_X1 U11391 ( .A1(n10225), .A2(n10224), .A3(n10223), .A4(n10222), .ZN(
        n10243) );
  AND4_X1 U11392 ( .A1(n10239), .A2(n10238), .A3(n10237), .A4(n10236), .ZN(
        n10240) );
  AND4_X1 U11393 ( .A1(n10231), .A2(n10230), .A3(n10229), .A4(n10228), .ZN(
        n10242) );
  NOR2_X1 U11394 ( .A1(n11309), .A2(n11308), .ZN(n11405) );
  AND3_X1 U11395 ( .A1(n11398), .A2(n11396), .A3(n11397), .ZN(n9837) );
  BUF_X4 U11396 ( .A(n15127), .Z(n17022) );
  INV_X2 U11397 ( .A(n16331), .ZN(U215) );
  AND2_X1 U11398 ( .A1(n10137), .A2(n10135), .ZN(n9813) );
  NAND2_X2 U11399 ( .A1(n18703), .A2(n18570), .ZN(n18622) );
  NAND2_X2 U11400 ( .A1(n18703), .A2(P3_STATE_REG_2__SCAN_IN), .ZN(n18631) );
  INV_X2 U11401 ( .A(n18687), .ZN(n17285) );
  NAND2_X2 U11402 ( .A1(P2_STATE_REG_2__SCAN_IN), .A2(n19815), .ZN(n19733) );
  INV_X1 U11403 ( .A(n16924), .ZN(n16824) );
  NAND2_X2 U11404 ( .A1(n19815), .A2(n19683), .ZN(n19736) );
  CLKBUF_X2 U11405 ( .A(n13881), .Z(n16990) );
  NAND4_X1 U11406 ( .A1(n11307), .A2(n11306), .A3(n11305), .A4(n11304), .ZN(
        n11308) );
  CLKBUF_X3 U11408 ( .A(n10483), .Z(n10734) );
  BUF_X2 U11409 ( .A(n10485), .Z(n11036) );
  BUF_X2 U11410 ( .A(n9626), .Z(n16923) );
  CLKBUF_X3 U11411 ( .A(n13962), .Z(n17005) );
  AND2_X1 U11412 ( .A1(n11354), .A2(n11347), .ZN(n11360) );
  AND2_X1 U11413 ( .A1(n11349), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11350) );
  OR2_X2 U11415 ( .A1(n13862), .A2(n18504), .ZN(n16777) );
  AND2_X1 U11416 ( .A1(n10140), .A2(n10143), .ZN(n10491) );
  AND2_X1 U11417 ( .A1(n13164), .A2(n10140), .ZN(n10483) );
  NOR2_X1 U11418 ( .A1(n13858), .A2(n9969), .ZN(n13881) );
  INV_X2 U11419 ( .A(n16336), .ZN(n16338) );
  NAND2_X1 U11420 ( .A1(n13943), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13862) );
  AND2_X2 U11421 ( .A1(n10134), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13167) );
  NAND2_X1 U11422 ( .A1(n13853), .A2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n13860) );
  NAND2_X1 U11423 ( .A1(n13943), .A2(n18647), .ZN(n13861) );
  AND2_X1 U11424 ( .A1(n10132), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10140) );
  AND2_X1 U11425 ( .A1(n10134), .A2(n9925), .ZN(n10141) );
  NAND2_X1 U11426 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n18647), .ZN(
        n13858) );
  INV_X2 U11427 ( .A(n19806), .ZN(n9634) );
  AND2_X1 U11428 ( .A1(n10133), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10139) );
  AND3_X2 U11429 ( .A1(n18705), .A2(n18636), .A3(n18704), .ZN(n17971) );
  AND2_X2 U11430 ( .A1(n9925), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13164) );
  INV_X1 U11431 ( .A(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n18668) );
  NAND2_X2 U11432 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n18504) );
  INV_X1 U11433 ( .A(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n13836) );
  AND2_X1 U11434 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10143) );
  AND2_X2 U11435 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10142) );
  NOR2_X1 U11436 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n11260) );
  INV_X1 U11437 ( .A(n17434), .ZN(n9635) );
  NAND2_X1 U11438 ( .A1(n9984), .A2(n17615), .ZN(n17411) );
  INV_X1 U11439 ( .A(n13651), .ZN(n9636) );
  NAND2_X1 U11440 ( .A1(n11399), .A2(n12068), .ZN(n11629) );
  INV_X1 U11441 ( .A(n11280), .ZN(n9637) );
  NAND2_X1 U11442 ( .A1(n13065), .A2(n13728), .ZN(n13152) );
  NOR2_X1 U11443 ( .A1(n11116), .A2(n13389), .ZN(n13174) );
  NOR2_X1 U11444 ( .A1(n12076), .A2(n12075), .ZN(n12083) );
  OR2_X2 U11445 ( .A1(n9650), .A2(n12519), .ZN(n12056) );
  OR2_X4 U11446 ( .A1(n9650), .A2(n13011), .ZN(n12053) );
  NOR2_X1 U11447 ( .A1(n14880), .A2(n14873), .ZN(n14872) );
  AND2_X1 U11448 ( .A1(n10140), .A2(n10141), .ZN(n10227) );
  XNOR2_X1 U11449 ( .A(n12411), .B(n12412), .ZN(n19085) );
  BUF_X1 U11450 ( .A(n13079), .Z(n9649) );
  NAND2_X2 U11451 ( .A1(n13834), .A2(n12425), .ZN(n13818) );
  XNOR2_X2 U11452 ( .A(n12016), .B(n12015), .ZN(n12519) );
  XNOR2_X2 U11453 ( .A(n11499), .B(n11501), .ZN(n12015) );
  OAI21_X2 U11454 ( .B1(n11477), .B2(n12448), .A(n11496), .ZN(n11499) );
  XNOR2_X1 U11455 ( .A(n12431), .B(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n14793) );
  XNOR2_X2 U11456 ( .A(n12429), .B(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n13817) );
  NAND2_X2 U11457 ( .A1(n12431), .A2(n12428), .ZN(n12429) );
  NAND2_X2 U11458 ( .A1(n12207), .A2(n9841), .ZN(n10100) );
  OAI22_X1 U11459 ( .A1(n12085), .A2(n12104), .B1(n19425), .B2(n12084), .ZN(
        n12089) );
  OAI21_X2 U11460 ( .B1(n14486), .B2(n10036), .A(n15569), .ZN(n15568) );
  AND2_X1 U11461 ( .A1(n10141), .A2(n10142), .ZN(n10319) );
  NAND3_X2 U11462 ( .A1(n11490), .A2(n11489), .A3(n11488), .ZN(n12023) );
  NAND2_X2 U11464 ( .A1(n11479), .A2(n11457), .ZN(n11497) );
  NOR2_X2 U11465 ( .A1(n13911), .A2(n13910), .ZN(n17078) );
  AND2_X2 U11466 ( .A1(n14271), .A2(n10665), .ZN(n14252) );
  NOR2_X4 U11467 ( .A1(n14880), .A2(n10053), .ZN(n12943) );
  OR2_X4 U11468 ( .A1(n14901), .A2(n14893), .ZN(n14880) );
  NAND2_X2 U11469 ( .A1(n9867), .A2(n9863), .ZN(n12936) );
  NAND2_X2 U11470 ( .A1(n12294), .A2(n10094), .ZN(n9867) );
  OAI21_X1 U11471 ( .B1(n12398), .B2(n12322), .A(n13555), .ZN(n12161) );
  XNOR2_X2 U11472 ( .A(n10265), .B(n10277), .ZN(n10300) );
  XNOR2_X2 U11473 ( .A(n12169), .B(n12198), .ZN(n12417) );
  NAND2_X2 U11474 ( .A1(n12103), .A2(n12102), .ZN(n12169) );
  NAND2_X2 U11475 ( .A1(n11951), .A2(n15286), .ZN(n13708) );
  OAI21_X2 U11476 ( .B1(n14323), .B2(n14324), .A(n10822), .ZN(n15468) );
  NOR2_X2 U11477 ( .A1(n14595), .A2(n14594), .ZN(n14593) );
  AND2_X2 U11478 ( .A1(n11650), .A2(n11258), .ZN(n9641) );
  INV_X2 U11479 ( .A(n11287), .ZN(n9642) );
  NAND2_X4 U11480 ( .A1(n11657), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11287) );
  OR2_X1 U11481 ( .A1(n11355), .A2(n11278), .ZN(n12675) );
  INV_X2 U11482 ( .A(n11355), .ZN(n12687) );
  OAI21_X2 U11483 ( .B1(n10353), .B2(n10352), .A(n10400), .ZN(n13434) );
  AND2_X4 U11484 ( .A1(n13612), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n9643) );
  NAND2_X4 U11485 ( .A1(n11658), .A2(n13620), .ZN(n11280) );
  AND2_X2 U11486 ( .A1(n11259), .A2(n11612), .ZN(n9645) );
  AND2_X1 U11487 ( .A1(n11259), .A2(n11612), .ZN(n9646) );
  NOR2_X4 U11488 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n11657) );
  NOR2_X1 U11489 ( .A1(n11495), .A2(n11494), .ZN(n11496) );
  NOR2_X2 U11490 ( .A1(n18692), .A2(n16349), .ZN(n17701) );
  BUF_X4 U11491 ( .A(n13079), .Z(n9650) );
  OAI21_X1 U11492 ( .B1(n12934), .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n12940), .ZN(n9754) );
  INV_X1 U11493 ( .A(n12938), .ZN(n9756) );
  AND2_X1 U11494 ( .A1(n9823), .A2(n10465), .ZN(n9822) );
  OR2_X1 U11495 ( .A1(n10849), .A2(n20597), .ZN(n10837) );
  INV_X1 U11496 ( .A(n12169), .ZN(n12201) );
  AND2_X1 U11497 ( .A1(n11621), .A2(n11620), .ZN(n11623) );
  INV_X1 U11498 ( .A(n10823), .ZN(n9938) );
  INV_X1 U11499 ( .A(n14243), .ZN(n9930) );
  INV_X1 U11500 ( .A(n10404), .ZN(n11054) );
  NAND2_X1 U11501 ( .A1(n10274), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n10580) );
  OR2_X1 U11502 ( .A1(n13489), .A2(n20599), .ZN(n11008) );
  NAND2_X1 U11503 ( .A1(n15620), .A2(n11190), .ZN(n10037) );
  NOR2_X1 U11504 ( .A1(n10042), .A2(n9687), .ZN(n10041) );
  INV_X1 U11505 ( .A(n11167), .ZN(n10042) );
  NOR2_X1 U11506 ( .A1(n20107), .A2(n20086), .ZN(n10849) );
  NAND2_X1 U11507 ( .A1(n10067), .A2(n10066), .ZN(n12333) );
  NAND2_X1 U11508 ( .A1(n12352), .A2(n11991), .ZN(n10066) );
  NAND2_X1 U11509 ( .A1(n12412), .A2(n12463), .ZN(n10067) );
  NOR2_X1 U11510 ( .A1(n12001), .A2(n10073), .ZN(n10072) );
  NOR2_X1 U11511 ( .A1(n13574), .A2(n11635), .ZN(n11443) );
  INV_X1 U11512 ( .A(n12412), .ZN(n12102) );
  NAND2_X1 U11513 ( .A1(n12526), .A2(n12525), .ZN(n12539) );
  NAND2_X1 U11514 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(n18668), .ZN(
        n9969) );
  NOR2_X1 U11515 ( .A1(n17201), .A2(n15193), .ZN(n15197) );
  OAI21_X1 U11516 ( .B1(n17666), .B2(n9653), .A(n9689), .ZN(n9986) );
  NOR2_X1 U11517 ( .A1(n9987), .A2(n17666), .ZN(n9985) );
  OAI21_X1 U11518 ( .B1(n15076), .B2(n15075), .A(n15074), .ZN(n15237) );
  NOR2_X1 U11519 ( .A1(n18087), .A2(n17227), .ZN(n15079) );
  OR2_X1 U11520 ( .A1(n20726), .A2(n12885), .ZN(n19922) );
  AND2_X1 U11521 ( .A1(n20599), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n11060) );
  OR3_X2 U11522 ( .A1(n14458), .A2(n11195), .A3(n11194), .ZN(n14446) );
  AOI21_X1 U11523 ( .B1(n13393), .B2(n13392), .A(n19820), .ZN(n13413) );
  NOR2_X1 U11524 ( .A1(n13382), .A2(n13381), .ZN(n13393) );
  NAND2_X1 U11525 ( .A1(n9878), .A2(n9877), .ZN(n9876) );
  NAND2_X1 U11526 ( .A1(n18831), .A2(n9879), .ZN(n9878) );
  OR2_X1 U11527 ( .A1(n9887), .A2(n11252), .ZN(n9877) );
  NAND2_X1 U11528 ( .A1(n15875), .A2(n14565), .ZN(n9879) );
  OR2_X1 U11529 ( .A1(n12209), .A2(n12327), .ZN(n12301) );
  NOR2_X1 U11530 ( .A1(n9688), .A2(n9999), .ZN(n9998) );
  INV_X1 U11531 ( .A(n12541), .ZN(n9999) );
  AND2_X1 U11532 ( .A1(n11250), .A2(n9739), .ZN(n11251) );
  NAND2_X1 U11533 ( .A1(n14580), .A2(n9742), .ZN(n12945) );
  INV_X1 U11534 ( .A(n12947), .ZN(n9965) );
  NOR2_X1 U11535 ( .A1(n9865), .A2(n9763), .ZN(n9863) );
  INV_X1 U11536 ( .A(n14716), .ZN(n9763) );
  INV_X1 U11537 ( .A(n19593), .ZN(n19528) );
  NAND2_X1 U11538 ( .A1(n10854), .A2(n10853), .ZN(n9771) );
  AND2_X1 U11539 ( .A1(n15343), .A2(n10833), .ZN(n10855) );
  OR2_X1 U11540 ( .A1(n10837), .A2(n11069), .ZN(n10856) );
  NAND2_X1 U11541 ( .A1(n11645), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n10077) );
  NAND2_X1 U11542 ( .A1(n11644), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(
        n10076) );
  NOR2_X1 U11543 ( .A1(n11463), .A2(n18715), .ZN(n9840) );
  OAI22_X1 U11544 ( .A1(n11492), .A2(n19685), .B1(n13649), .B2(n13007), .ZN(
        n11462) );
  NAND2_X1 U11545 ( .A1(n10401), .A2(n9823), .ZN(n9819) );
  NAND2_X1 U11546 ( .A1(n10264), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n10277) );
  OAI21_X1 U11547 ( .B1(n11454), .B2(n12451), .A(P2_STATE2_REG_0__SCAN_IN), 
        .ZN(n11481) );
  AND2_X1 U11548 ( .A1(n12199), .A2(n12198), .ZN(n12200) );
  AOI22_X1 U11549 ( .A1(n12841), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n12687), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11398) );
  NAND2_X1 U11550 ( .A1(n11391), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n9869) );
  NAND2_X1 U11551 ( .A1(n9643), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n9868) );
  NAND2_X1 U11552 ( .A1(n11624), .A2(n11617), .ZN(n11621) );
  AND2_X1 U11553 ( .A1(n15244), .A2(n15188), .ZN(n15191) );
  NOR2_X1 U11554 ( .A1(n9612), .A2(n15248), .ZN(n15188) );
  AND2_X1 U11556 ( .A1(n14350), .A2(n14255), .ZN(n9931) );
  INV_X1 U11557 ( .A(n11057), .ZN(n11030) );
  NOR2_X1 U11558 ( .A1(n9934), .A2(n9933), .ZN(n9932) );
  INV_X1 U11559 ( .A(n14101), .ZN(n9933) );
  INV_X1 U11560 ( .A(n9935), .ZN(n9934) );
  INV_X1 U11561 ( .A(n10580), .ZN(n10609) );
  XNOR2_X1 U11562 ( .A(n11157), .B(n10476), .ZN(n11108) );
  NAND2_X1 U11563 ( .A1(n15409), .A2(n13386), .ZN(n13391) );
  NOR2_X1 U11564 ( .A1(n10329), .A2(n10328), .ZN(n10348) );
  INV_X1 U11565 ( .A(n10313), .ZN(n9940) );
  NAND3_X1 U11566 ( .A1(n20128), .A2(n20597), .A3(n10302), .ZN(n9941) );
  XNOR2_X1 U11567 ( .A(n10348), .B(n10349), .ZN(n10372) );
  NAND2_X1 U11568 ( .A1(n9820), .A2(n10401), .ZN(n10424) );
  NAND2_X1 U11569 ( .A1(n9676), .A2(n10302), .ZN(n9798) );
  INV_X1 U11570 ( .A(n10285), .ZN(n10027) );
  AOI221_X1 U11571 ( .B1(n20725), .B2(n14179), .C1(n15412), .C2(n14179), .A(
        P1_STATE2_REG_0__SCAN_IN), .ZN(n20218) );
  AND2_X1 U11572 ( .A1(n10862), .A2(n11154), .ZN(n10867) );
  INV_X1 U11573 ( .A(n10837), .ZN(n10866) );
  NOR2_X1 U11574 ( .A1(n15861), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n9776) );
  OAI22_X1 U11575 ( .A1(n10864), .A2(n10863), .B1(n10862), .B2(n11071), .ZN(
        n10865) );
  AOI21_X1 U11576 ( .B1(n9768), .B2(n9766), .A(n9765), .ZN(n10864) );
  NOR2_X1 U11577 ( .A1(n10862), .A2(n10857), .ZN(n9765) );
  NOR2_X1 U11578 ( .A1(n12289), .A2(n12288), .ZN(n10057) );
  OR2_X1 U11579 ( .A1(n12239), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n12242) );
  OR2_X1 U11580 ( .A1(n14628), .A2(n14688), .ZN(n9995) );
  AND2_X1 U11581 ( .A1(n12567), .A2(n13719), .ZN(n10017) );
  INV_X1 U11582 ( .A(n14612), .ZN(n9966) );
  INV_X1 U11583 ( .A(n9957), .ZN(n9954) );
  NOR2_X1 U11584 ( .A1(n15886), .A2(n12426), .ZN(n12940) );
  AND2_X1 U11585 ( .A1(n12317), .A2(n14715), .ZN(n12938) );
  OR2_X1 U11586 ( .A1(n15901), .A2(n12426), .ZN(n12937) );
  NAND2_X1 U11587 ( .A1(n15909), .A2(n12322), .ZN(n12314) );
  AND3_X1 U11588 ( .A1(n14738), .A2(n10086), .A3(n10085), .ZN(n10084) );
  NOR2_X1 U11589 ( .A1(n14747), .A2(n10087), .ZN(n10086) );
  NAND2_X1 U11590 ( .A1(n10093), .A2(n10089), .ZN(n10087) );
  NAND2_X1 U11591 ( .A1(n15290), .A2(n13720), .ZN(n9957) );
  NOR2_X1 U11592 ( .A1(n9846), .A2(n14729), .ZN(n9845) );
  INV_X1 U11593 ( .A(n9848), .ZN(n9846) );
  NAND2_X1 U11594 ( .A1(n14966), .A2(n9913), .ZN(n9912) );
  INV_X1 U11595 ( .A(n16089), .ZN(n9913) );
  INV_X1 U11596 ( .A(n11609), .ZN(n11608) );
  AND2_X1 U11597 ( .A1(n9963), .A2(n9961), .ZN(n9960) );
  INV_X1 U11598 ( .A(n13233), .ZN(n9961) );
  AND2_X1 U11599 ( .A1(n11739), .A2(n10069), .ZN(n10068) );
  INV_X1 U11600 ( .A(n12398), .ZN(n10046) );
  NAND2_X1 U11601 ( .A1(n9607), .A2(n9783), .ZN(n9782) );
  INV_X1 U11602 ( .A(n11468), .ZN(n9783) );
  NAND3_X1 U11603 ( .A1(n12861), .A2(n11473), .A3(n11472), .ZN(n13600) );
  INV_X1 U11604 ( .A(n12055), .ZN(n12032) );
  NOR2_X1 U11605 ( .A1(n11382), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11386) );
  INV_X1 U11606 ( .A(n11381), .ZN(n11382) );
  NOR2_X1 U11607 ( .A1(n11376), .A2(n11278), .ZN(n11380) );
  INV_X1 U11608 ( .A(n11375), .ZN(n11376) );
  OAI21_X1 U11609 ( .B1(n16348), .B2(n15234), .A(n18481), .ZN(n15080) );
  NOR2_X1 U11610 ( .A1(n16480), .A2(n10009), .ZN(n10007) );
  NAND2_X1 U11611 ( .A1(n17419), .A2(n10010), .ZN(n10009) );
  INV_X1 U11612 ( .A(n15170), .ZN(n15127) );
  INV_X1 U11613 ( .A(n17290), .ZN(n15084) );
  NAND2_X1 U11614 ( .A1(n16217), .A2(n16216), .ZN(n17344) );
  NAND2_X1 U11615 ( .A1(n16215), .A2(n15213), .ZN(n16216) );
  NAND2_X1 U11616 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n15204) );
  NOR2_X1 U11617 ( .A1(n15262), .A2(n17637), .ZN(n15265) );
  OAI21_X1 U11618 ( .B1(n10125), .B2(n17193), .A(n17615), .ZN(n15200) );
  AOI21_X1 U11619 ( .B1(n15196), .B2(n9972), .A(n15199), .ZN(n9971) );
  NOR2_X1 U11620 ( .A1(n15187), .A2(n15186), .ZN(n15190) );
  NOR2_X1 U11621 ( .A1(n17689), .A2(n17690), .ZN(n15187) );
  NOR3_X1 U11622 ( .A1(n18495), .A2(n15067), .A3(n15227), .ZN(n15235) );
  NOR2_X1 U11623 ( .A1(n13932), .A2(n13931), .ZN(n15076) );
  NOR2_X1 U11624 ( .A1(n14228), .A2(n20599), .ZN(n14299) );
  INV_X1 U11625 ( .A(n14299), .ZN(n14296) );
  INV_X1 U11626 ( .A(n13143), .ZN(n9826) );
  INV_X1 U11627 ( .A(n13142), .ZN(n9827) );
  NOR2_X1 U11628 ( .A1(n15409), .A2(n13160), .ZN(n13382) );
  NAND2_X1 U11629 ( .A1(n15409), .A2(n11065), .ZN(n15404) );
  INV_X1 U11630 ( .A(n11008), .ZN(n11061) );
  NOR2_X1 U11631 ( .A1(n14198), .A2(n9927), .ZN(n9926) );
  INV_X1 U11632 ( .A(n11099), .ZN(n9927) );
  NOR2_X1 U11633 ( .A1(n11011), .A2(n14232), .ZN(n11012) );
  AND2_X1 U11634 ( .A1(n9667), .A2(n14327), .ZN(n9937) );
  NOR2_X1 U11635 ( .A1(n10698), .A2(n10697), .ZN(n10699) );
  INV_X1 U11636 ( .A(n10477), .ZN(n10478) );
  NAND2_X1 U11637 ( .A1(n10478), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n10500) );
  OAI21_X1 U11638 ( .B1(n13434), .B2(n10580), .A(n10357), .ZN(n10358) );
  AND2_X1 U11639 ( .A1(n15409), .A2(n13396), .ZN(n15356) );
  NOR2_X1 U11640 ( .A1(n11193), .A2(n9806), .ZN(n9805) );
  INV_X1 U11641 ( .A(n15567), .ZN(n9806) );
  NAND2_X1 U11642 ( .A1(n14468), .A2(n15567), .ZN(n9810) );
  NOR2_X1 U11643 ( .A1(n14225), .A2(n14224), .ZN(n14314) );
  OR2_X1 U11644 ( .A1(n14331), .A2(n14320), .ZN(n14322) );
  NAND2_X1 U11645 ( .A1(n14338), .A2(n14329), .ZN(n14331) );
  AOI21_X1 U11646 ( .B1(n11191), .B2(n10031), .A(n15569), .ZN(n10030) );
  INV_X1 U11647 ( .A(n10034), .ZN(n10031) );
  INV_X1 U11648 ( .A(n15599), .ZN(n11191) );
  XNOR2_X1 U11649 ( .A(n15620), .B(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n15598) );
  INV_X1 U11650 ( .A(n10041), .ZN(n9804) );
  INV_X1 U11651 ( .A(n9674), .ZN(n9803) );
  NAND2_X1 U11652 ( .A1(n9789), .A2(n13494), .ZN(n9788) );
  INV_X1 U11653 ( .A(n11146), .ZN(n9789) );
  AND2_X1 U11654 ( .A1(n15857), .A2(n20597), .ZN(n11205) );
  NAND2_X1 U11655 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n15409), .ZN(n14179) );
  AOI221_X1 U11656 ( .B1(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B2(n11627), 
        .C1(n13643), .C2(n11627), .A(n11618), .ZN(n12365) );
  NAND2_X1 U11657 ( .A1(n12337), .A2(n9759), .ZN(n12360) );
  INV_X1 U11658 ( .A(n9948), .ZN(n9945) );
  NOR2_X1 U11659 ( .A1(n12313), .A2(n12307), .ZN(n12319) );
  NAND2_X1 U11660 ( .A1(n15881), .A2(n12960), .ZN(n15882) );
  NOR2_X1 U11661 ( .A1(n12299), .A2(P2_EBX_REG_25__SCAN_IN), .ZN(n12304) );
  NAND2_X1 U11662 ( .A1(n10057), .A2(n10056), .ZN(n12299) );
  INV_X1 U11663 ( .A(n15977), .ZN(n9886) );
  INV_X1 U11664 ( .A(n10057), .ZN(n12297) );
  NAND2_X1 U11665 ( .A1(n12261), .A2(n9717), .ZN(n12284) );
  OR2_X1 U11666 ( .A1(n9887), .A2(n18754), .ZN(n9889) );
  OR2_X1 U11667 ( .A1(n14072), .A2(n14769), .ZN(n9890) );
  OR2_X1 U11668 ( .A1(n12209), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n11996) );
  NAND2_X1 U11669 ( .A1(n10064), .A2(n10060), .ZN(n12209) );
  NOR2_X1 U11670 ( .A1(n12165), .A2(n10061), .ZN(n10060) );
  INV_X1 U11671 ( .A(n12146), .ZN(n10063) );
  AND2_X1 U11672 ( .A1(n12548), .A2(n13365), .ZN(n13364) );
  NAND2_X1 U11673 ( .A1(n9918), .A2(n9917), .ZN(n14677) );
  INV_X1 U11674 ( .A(n12981), .ZN(n9917) );
  INV_X1 U11675 ( .A(n12980), .ZN(n9918) );
  INV_X1 U11676 ( .A(n13843), .ZN(n9915) );
  AND2_X1 U11677 ( .A1(n12634), .A2(n13845), .ZN(n10025) );
  NOR2_X2 U11678 ( .A1(n19796), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n13044) );
  NAND2_X1 U11679 ( .A1(n12505), .A2(n9950), .ZN(n9946) );
  AND2_X1 U11680 ( .A1(n9951), .A2(n12469), .ZN(n9950) );
  OR2_X1 U11681 ( .A1(n12505), .A2(n9951), .ZN(n9947) );
  NAND2_X1 U11682 ( .A1(n14580), .A2(n9737), .ZN(n14610) );
  AOI21_X1 U11683 ( .B1(n9850), .B2(n10090), .A(n9849), .ZN(n9848) );
  INV_X1 U11684 ( .A(n14959), .ZN(n9849) );
  OR3_X1 U11685 ( .A1(n12272), .A2(n12426), .A3(n12433), .ZN(n16019) );
  INV_X1 U11686 ( .A(n14706), .ZN(n9859) );
  XNOR2_X1 U11687 ( .A(n12314), .B(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n14716) );
  AOI21_X1 U11688 ( .B1(n10097), .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A(
        n10095), .ZN(n10094) );
  INV_X1 U11689 ( .A(n12293), .ZN(n10095) );
  NAND2_X1 U11690 ( .A1(n15019), .A2(n12435), .ZN(n14752) );
  INV_X1 U11691 ( .A(n15285), .ZN(n11951) );
  AND2_X1 U11692 ( .A1(n12206), .A2(n9711), .ZN(n9841) );
  OAI21_X1 U11693 ( .B1(n13817), .B2(n10051), .A(n14793), .ZN(n10050) );
  NAND2_X1 U11694 ( .A1(n13818), .A2(n13817), .ZN(n13816) );
  INV_X1 U11695 ( .A(n13068), .ZN(n12538) );
  OR2_X1 U11696 ( .A1(n19138), .A2(n18999), .ZN(n19459) );
  NAND2_X1 U11697 ( .A1(n19138), .A2(n18999), .ZN(n19533) );
  NAND2_X1 U11698 ( .A1(n19754), .A2(n19779), .ZN(n19555) );
  NAND2_X1 U11699 ( .A1(n19754), .A2(n19137), .ZN(n19534) );
  NAND2_X1 U11700 ( .A1(n13563), .A2(n13562), .ZN(n19593) );
  NAND2_X1 U11701 ( .A1(n19138), .A2(n19767), .ZN(n19587) );
  NOR2_X2 U11702 ( .A1(n15084), .A2(n15080), .ZN(n18484) );
  NAND2_X1 U11703 ( .A1(n10011), .A2(n17419), .ZN(n10008) );
  NOR2_X1 U11704 ( .A1(n16480), .A2(n17431), .ZN(n16479) );
  INV_X2 U11705 ( .A(n14010), .ZN(n17013) );
  INV_X1 U11706 ( .A(n15136), .ZN(n15137) );
  AOI211_X1 U11707 ( .C1(n17005), .C2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .A(
        n13888), .B(n13887), .ZN(n13889) );
  NOR2_X1 U11708 ( .A1(n16693), .A2(n9672), .ZN(n16189) );
  NOR2_X1 U11709 ( .A1(n17489), .A2(n17490), .ZN(n17466) );
  AND2_X1 U11710 ( .A1(n17546), .A2(n10018), .ZN(n17503) );
  INV_X1 U11711 ( .A(n17507), .ZN(n10018) );
  NOR2_X1 U11712 ( .A1(n16606), .A2(n16616), .ZN(n17546) );
  NAND2_X1 U11713 ( .A1(n17363), .A2(n15213), .ZN(n16219) );
  OR2_X1 U11714 ( .A1(n17399), .A2(n15213), .ZN(n17386) );
  AND2_X1 U11715 ( .A1(n17588), .A2(n17948), .ZN(n9991) );
  INV_X1 U11716 ( .A(n17227), .ZN(n18047) );
  AND2_X1 U11717 ( .A1(n19922), .A2(n12889), .ZN(n19872) );
  NAND2_X1 U11718 ( .A1(n20128), .A2(n10302), .ZN(n20438) );
  NAND2_X1 U11719 ( .A1(n9829), .A2(n9828), .ZN(n12899) );
  NAND2_X1 U11720 ( .A1(n14209), .A2(n14201), .ZN(n9828) );
  INV_X1 U11721 ( .A(n19940), .ZN(n14356) );
  INV_X1 U11722 ( .A(n14437), .ZN(n14422) );
  AND2_X1 U11723 ( .A1(n20039), .A2(n11204), .ZN(n15635) );
  INV_X1 U11724 ( .A(n20039), .ZN(n20034) );
  AND2_X1 U11725 ( .A1(n9777), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n15672) );
  OAI21_X1 U11726 ( .B1(n15675), .B2(n15673), .A(n15676), .ZN(n9777) );
  XNOR2_X1 U11727 ( .A(n12923), .B(n11197), .ZN(n15668) );
  NAND2_X1 U11728 ( .A1(n15683), .A2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n9817) );
  NOR2_X1 U11729 ( .A1(n15719), .A2(n9773), .ZN(n15718) );
  AND2_X1 U11730 ( .A1(n15834), .A2(n15722), .ZN(n9773) );
  AND2_X1 U11731 ( .A1(n13413), .A2(n13412), .ZN(n20064) );
  INV_X1 U11732 ( .A(n20064), .ZN(n20081) );
  NOR2_X1 U11733 ( .A1(n9651), .A2(n18890), .ZN(n9873) );
  NAND2_X1 U11734 ( .A1(n9876), .A2(n9880), .ZN(n9875) );
  NAND2_X1 U11735 ( .A1(n9881), .A2(n11252), .ZN(n9880) );
  INV_X1 U11736 ( .A(n14565), .ZN(n9881) );
  AND2_X1 U11737 ( .A1(n15882), .A2(n9887), .ZN(n14566) );
  OR2_X1 U11738 ( .A1(n19804), .A2(n11985), .ZN(n18932) );
  INV_X1 U11739 ( .A(n18924), .ZN(n18916) );
  OR3_X1 U11740 ( .A1(n11987), .A2(n12476), .A3(n11986), .ZN(n18923) );
  NAND2_X1 U11741 ( .A1(n14820), .A2(n9923), .ZN(n9922) );
  AOI21_X1 U11742 ( .B1(n14817), .B2(n19131), .A(n14816), .ZN(n9923) );
  NOR2_X1 U11743 ( .A1(n14822), .A2(n14821), .ZN(n9921) );
  OR2_X1 U11744 ( .A1(n14573), .A2(n14572), .ZN(n9924) );
  XNOR2_X1 U11745 ( .A(n12498), .B(n10103), .ZN(n14826) );
  OR2_X1 U11746 ( .A1(n12481), .A2(n12445), .ZN(n16128) );
  INV_X1 U11747 ( .A(n19125), .ZN(n16122) );
  INV_X1 U11748 ( .A(n16128), .ZN(n19122) );
  INV_X1 U11749 ( .A(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19783) );
  INV_X1 U11750 ( .A(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n19773) );
  NOR2_X1 U11751 ( .A1(n19534), .A2(n19395), .ZN(n19445) );
  XNOR2_X1 U11752 ( .A(n16393), .B(n10024), .ZN(n10023) );
  INV_X1 U11753 ( .A(n16394), .ZN(n10024) );
  NAND2_X1 U11754 ( .A1(P3_STATE2_REG_3__SCAN_IN), .A2(n16752), .ZN(n16739) );
  NAND2_X1 U11755 ( .A1(n18511), .A2(n17186), .ZN(n17214) );
  NOR2_X1 U11756 ( .A1(n18650), .A2(n17700), .ZN(n17565) );
  NAND2_X1 U11757 ( .A1(n9648), .A2(n17193), .ZN(n17617) );
  NAND2_X1 U11758 ( .A1(n17707), .A2(n17668), .ZN(n17700) );
  INV_X1 U11759 ( .A(n17940), .ZN(n17933) );
  INV_X1 U11760 ( .A(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12186) );
  INV_X1 U11761 ( .A(n10423), .ZN(n9823) );
  AND3_X1 U11762 ( .A1(n11364), .A2(n11363), .A3(n11347), .ZN(n11367) );
  OR2_X1 U11763 ( .A1(n11287), .A2(n12074), .ZN(n11274) );
  NAND2_X1 U11764 ( .A1(n9641), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(
        n11255) );
  OR2_X1 U11765 ( .A1(n11280), .A2(n11253), .ZN(n11254) );
  OR2_X1 U11766 ( .A1(n11287), .A2(n11339), .ZN(n11343) );
  AND2_X1 U11767 ( .A1(n10827), .A2(n10826), .ZN(n10835) );
  NAND2_X1 U11768 ( .A1(n9795), .A2(n20086), .ZN(n10259) );
  OR2_X1 U11769 ( .A1(n10312), .A2(n10311), .ZN(n11104) );
  OR2_X1 U11770 ( .A1(n10419), .A2(n10418), .ZN(n11139) );
  NOR2_X1 U11771 ( .A1(n13410), .A2(n20597), .ZN(n10340) );
  AOI22_X1 U11772 ( .A1(n10458), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n10187), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n10151) );
  OR2_X1 U11773 ( .A1(n10854), .A2(n10853), .ZN(n9769) );
  NAND2_X1 U11774 ( .A1(n9771), .A2(n9713), .ZN(n9770) );
  INV_X1 U11775 ( .A(n9767), .ZN(n9766) );
  OAI22_X1 U11776 ( .A1(n10856), .A2(n10855), .B1(n11141), .B2(n10857), .ZN(
        n9767) );
  OAI22_X1 U11777 ( .A1(n11287), .A2(n19175), .B1(n11355), .B2(n12815), .ZN(
        n12816) );
  NAND2_X1 U11778 ( .A1(n11456), .A2(n11455), .ZN(n11480) );
  NAND2_X1 U11779 ( .A1(n19156), .A2(n12453), .ZN(n11455) );
  AND2_X1 U11780 ( .A1(n12266), .A2(n14735), .ZN(n10093) );
  OR2_X1 U11781 ( .A1(n11764), .A2(n11763), .ZN(n12141) );
  NOR2_X1 U11782 ( .A1(n10071), .A2(n10070), .ZN(n10069) );
  INV_X1 U11783 ( .A(n11736), .ZN(n10071) );
  INV_X1 U11784 ( .A(n11738), .ZN(n10070) );
  OAI21_X1 U11785 ( .B1(n12675), .B2(n11734), .A(n10074), .ZN(n11735) );
  NAND2_X1 U11786 ( .A1(n10077), .A2(n10076), .ZN(n10075) );
  AOI22_X1 U11787 ( .A1(n13606), .A2(P2_STATE2_REG_0__SCAN_IN), .B1(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n11510), .ZN(n11460) );
  NAND3_X1 U11788 ( .A1(n9678), .A2(n9839), .A3(n9838), .ZN(n11467) );
  NAND2_X1 U11789 ( .A1(n12470), .A2(n9840), .ZN(n9839) );
  OR2_X1 U11790 ( .A1(n11727), .A2(n11726), .ZN(n12099) );
  INV_X1 U11791 ( .A(n12375), .ZN(n11451) );
  INV_X1 U11792 ( .A(n12052), .ZN(n12030) );
  AOI22_X1 U11793 ( .A1(n11391), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n12846), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n11294) );
  AOI22_X1 U11794 ( .A1(n11391), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n9644), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11283) );
  OR2_X1 U11795 ( .A1(n11287), .A2(n11314), .ZN(n11318) );
  OR2_X1 U11796 ( .A1(n11287), .A2(n11302), .ZN(n11307) );
  NAND2_X2 U11797 ( .A1(n13612), .A2(n11258), .ZN(n11355) );
  NAND2_X1 U11798 ( .A1(n11615), .A2(n11614), .ZN(n11626) );
  OR2_X1 U11799 ( .A1(n12359), .A2(n12154), .ZN(n11615) );
  AND2_X1 U11800 ( .A1(n11617), .A2(n11616), .ZN(n11625) );
  NAND2_X1 U11801 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n19783), .ZN(
        n12154) );
  INV_X1 U11802 ( .A(n17642), .ZN(n9972) );
  OR2_X1 U11803 ( .A1(n15061), .A2(n15060), .ZN(n13944) );
  NOR2_X1 U11804 ( .A1(n10583), .A2(n9936), .ZN(n9935) );
  NOR2_X1 U11805 ( .A1(n14085), .A2(n14089), .ZN(n9936) );
  NAND2_X1 U11806 ( .A1(n9605), .A2(n14085), .ZN(n14090) );
  NAND2_X1 U11807 ( .A1(n15568), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n11196) );
  OR2_X1 U11808 ( .A1(n14224), .A2(n9831), .ZN(n9830) );
  INV_X1 U11809 ( .A(n14313), .ZN(n9831) );
  OR2_X1 U11810 ( .A1(n10036), .A2(n15620), .ZN(n10033) );
  NAND2_X1 U11811 ( .A1(n10107), .A2(n10035), .ZN(n10034) );
  INV_X1 U11812 ( .A(n9671), .ZN(n9793) );
  NAND2_X1 U11813 ( .A1(n9787), .A2(n11129), .ZN(n11135) );
  NAND2_X1 U11814 ( .A1(n13354), .A2(n13355), .ZN(n9787) );
  AOI22_X1 U11815 ( .A1(n9620), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n10208), .B2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n10188) );
  AOI22_X1 U11816 ( .A1(n9616), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n10213), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n10189) );
  AOI22_X1 U11817 ( .A1(n10734), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n10187), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n10191) );
  NAND2_X1 U11818 ( .A1(n9833), .A2(n10873), .ZN(n10877) );
  NOR2_X1 U11819 ( .A1(n13184), .A2(n13384), .ZN(n13394) );
  OR2_X1 U11820 ( .A1(n10339), .A2(n10338), .ZN(n11117) );
  INV_X1 U11821 ( .A(n11117), .ZN(n11109) );
  OR2_X1 U11822 ( .A1(n13423), .A2(n13422), .ZN(n15340) );
  NAND2_X1 U11823 ( .A1(n9795), .A2(n10249), .ZN(n13186) );
  CLKBUF_X1 U11824 ( .A(n12880), .Z(n12881) );
  INV_X1 U11825 ( .A(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20326) );
  NOR2_X1 U11826 ( .A1(n10169), .A2(n10170), .ZN(n9815) );
  NAND2_X1 U11827 ( .A1(n20684), .A2(n20597), .ZN(n10399) );
  NOR2_X1 U11828 ( .A1(n11435), .A2(n11414), .ZN(n11348) );
  NAND2_X1 U11829 ( .A1(n12224), .A2(n9705), .ZN(n12251) );
  NAND2_X1 U11830 ( .A1(n12224), .A2(n12231), .ZN(n12257) );
  AND2_X1 U11831 ( .A1(n11429), .A2(n10059), .ZN(n10058) );
  NOR2_X1 U11832 ( .A1(n12166), .A2(n10065), .ZN(n10064) );
  NAND2_X1 U11833 ( .A1(n12203), .A2(n12146), .ZN(n10065) );
  AND2_X1 U11834 ( .A1(n14581), .A2(n14615), .ZN(n9967) );
  CLKBUF_X1 U11835 ( .A(n12687), .Z(n12842) );
  INV_X1 U11836 ( .A(n12479), .ZN(n9951) );
  AND2_X1 U11837 ( .A1(n9899), .A2(n9726), .ZN(n9898) );
  NAND2_X1 U11838 ( .A1(n9760), .A2(n11698), .ZN(n12404) );
  NOR2_X1 U11839 ( .A1(n11703), .A2(n9761), .ZN(n9760) );
  INV_X1 U11840 ( .A(n12940), .ZN(n9758) );
  INV_X1 U11841 ( .A(n14853), .ZN(n9866) );
  OR2_X1 U11842 ( .A1(n10055), .A2(n11967), .ZN(n10054) );
  NAND2_X1 U11843 ( .A1(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n10055) );
  NAND2_X1 U11844 ( .A1(n9786), .A2(n9785), .ZN(n16039) );
  NOR2_X1 U11845 ( .A1(n15023), .A2(n10099), .ZN(n10098) );
  INV_X1 U11846 ( .A(n12215), .ZN(n10099) );
  NOR2_X1 U11847 ( .A1(n13244), .A2(n9958), .ZN(n13228) );
  NAND2_X1 U11848 ( .A1(n9960), .A2(n9959), .ZN(n9958) );
  INV_X1 U11849 ( .A(n9748), .ZN(n9959) );
  INV_X1 U11850 ( .A(n16113), .ZN(n9914) );
  NOR2_X1 U11851 ( .A1(n9964), .A2(n13245), .ZN(n9963) );
  INV_X1 U11852 ( .A(n13274), .ZN(n9964) );
  INV_X1 U11853 ( .A(n13244), .ZN(n9962) );
  NAND2_X1 U11854 ( .A1(n12205), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n12206) );
  OR2_X1 U11855 ( .A1(n11781), .A2(n11780), .ZN(n12193) );
  INV_X1 U11856 ( .A(n11493), .ZN(n11495) );
  AND2_X1 U11857 ( .A1(n11558), .A2(P2_EBX_REG_2__SCAN_IN), .ZN(n11494) );
  NAND2_X1 U11858 ( .A1(n11512), .A2(n11511), .ZN(n11513) );
  OR2_X1 U11859 ( .A1(n11477), .A2(n12162), .ZN(n11509) );
  NOR2_X1 U11860 ( .A1(n13600), .A2(n11474), .ZN(n13589) );
  NAND2_X2 U11861 ( .A1(n9870), .A2(n9836), .ZN(n11635) );
  NAND2_X1 U11862 ( .A1(n9677), .A2(n9837), .ZN(n9836) );
  OAI21_X2 U11863 ( .B1(n11406), .B2(n11278), .A(n11277), .ZN(n11435) );
  AOI22_X1 U11864 ( .A1(n12841), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n12687), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11353) );
  AND3_X1 U11865 ( .A1(n13643), .A2(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A3(
        n11627), .ZN(n12352) );
  OR2_X1 U11866 ( .A1(n11623), .A2(n11622), .ZN(n12346) );
  INV_X1 U11867 ( .A(n15236), .ZN(n15067) );
  OR2_X1 U11868 ( .A1(n18076), .A2(n15066), .ZN(n15073) );
  OR2_X1 U11869 ( .A1(n16741), .A2(n13858), .ZN(n15170) );
  INV_X1 U11870 ( .A(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n20830) );
  NOR2_X1 U11871 ( .A1(n15257), .A2(n17651), .ZN(n15260) );
  NOR2_X1 U11872 ( .A1(n13942), .A2(n13941), .ZN(n15221) );
  INV_X1 U11873 ( .A(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n18517) );
  INV_X1 U11875 ( .A(n13145), .ZN(n12897) );
  OR2_X1 U11876 ( .A1(n14209), .A2(n10878), .ZN(n9829) );
  INV_X1 U11877 ( .A(n14339), .ZN(n10762) );
  INV_X1 U11878 ( .A(n19996), .ZN(n19947) );
  OR2_X1 U11879 ( .A1(n11014), .A2(n11013), .ZN(n14312) );
  CLKBUF_X1 U11880 ( .A(n11096), .Z(n11097) );
  NOR2_X1 U11881 ( .A1(n10803), .A2(n10802), .ZN(n10804) );
  AOI21_X1 U11882 ( .B1(n10801), .B2(n10800), .A(n10799), .ZN(n14324) );
  AND2_X1 U11883 ( .A1(n11054), .A2(n15470), .ZN(n10799) );
  NOR2_X1 U11884 ( .A1(n10763), .A2(n15496), .ZN(n10764) );
  NAND2_X1 U11885 ( .A1(n10764), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n10803) );
  NOR2_X1 U11886 ( .A1(n10717), .A2(n15506), .ZN(n10718) );
  NAND2_X1 U11887 ( .A1(n10718), .A2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n10763) );
  AND2_X1 U11888 ( .A1(n10716), .A2(n10715), .ZN(n14348) );
  AND2_X1 U11889 ( .A1(n10701), .A2(n10700), .ZN(n14350) );
  AND2_X1 U11890 ( .A1(n10681), .A2(n10680), .ZN(n14255) );
  NOR2_X1 U11891 ( .A1(n10648), .A2(n10647), .ZN(n10649) );
  NAND2_X1 U11892 ( .A1(n10649), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n10698) );
  NOR2_X1 U11893 ( .A1(n10624), .A2(n14290), .ZN(n10643) );
  NAND2_X1 U11894 ( .A1(n10643), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n10648) );
  NAND2_X1 U11896 ( .A1(n10584), .A2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n10600) );
  NOR2_X1 U11897 ( .A1(n10567), .A2(n10551), .ZN(n10584) );
  AND2_X1 U11898 ( .A1(n10537), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n10538) );
  NAND2_X1 U11899 ( .A1(n10538), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n10567) );
  INV_X1 U11901 ( .A(n13769), .ZN(n10519) );
  OAI21_X1 U11902 ( .B1(n11108), .B2(n10580), .A(n10482), .ZN(n13581) );
  NOR2_X1 U11903 ( .A1(n10447), .A2(n15664), .ZN(n10467) );
  NAND2_X1 U11904 ( .A1(n10426), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n10447) );
  NAND2_X1 U11905 ( .A1(n10453), .A2(n10452), .ZN(n13458) );
  NAND2_X1 U11906 ( .A1(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n10403) );
  NOR2_X1 U11907 ( .A1(n10403), .A2(n19908), .ZN(n10426) );
  NAND2_X1 U11908 ( .A1(n15689), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n15675) );
  AND2_X1 U11909 ( .A1(n15718), .A2(n9772), .ZN(n15703) );
  NAND2_X1 U11910 ( .A1(n15798), .A2(n15717), .ZN(n9772) );
  OR2_X1 U11911 ( .A1(n14238), .A2(n9835), .ZN(n9834) );
  INV_X1 U11912 ( .A(n14335), .ZN(n9835) );
  NOR3_X1 U11913 ( .A1(n14353), .A2(n10946), .A3(n14238), .ZN(n14336) );
  AND2_X1 U11914 ( .A1(n9818), .A2(n9714), .ZN(n15618) );
  NAND2_X1 U11915 ( .A1(n15544), .A2(n9703), .ZN(n14132) );
  AND2_X1 U11916 ( .A1(n15544), .A2(n15543), .ZN(n15546) );
  AND2_X1 U11917 ( .A1(n10909), .A2(n10908), .ZN(n13784) );
  NOR2_X1 U11918 ( .A1(n13785), .A2(n13784), .ZN(n15544) );
  INV_X1 U11919 ( .A(n14499), .ZN(n15638) );
  OR2_X1 U11920 ( .A1(n13771), .A2(n13772), .ZN(n13785) );
  NAND2_X1 U11921 ( .A1(n13659), .A2(n13658), .ZN(n13771) );
  AND2_X1 U11922 ( .A1(n10900), .A2(n10899), .ZN(n15849) );
  INV_X1 U11923 ( .A(n13333), .ZN(n9824) );
  XNOR2_X1 U11924 ( .A(n11135), .B(n13409), .ZN(n13350) );
  NOR2_X1 U11925 ( .A1(n15773), .A2(n15376), .ZN(n15819) );
  AND2_X1 U11926 ( .A1(n13413), .A2(n14182), .ZN(n15376) );
  AND2_X1 U11927 ( .A1(n10953), .A2(n14200), .ZN(n13145) );
  AOI21_X1 U11928 ( .B1(n10862), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .A(
        n10298), .ZN(n10299) );
  NAND2_X1 U11929 ( .A1(n9941), .A2(n9939), .ZN(n10351) );
  NAND2_X1 U11930 ( .A1(n10040), .A2(n15358), .ZN(n15366) );
  OR2_X1 U11931 ( .A1(n15340), .A2(n10038), .ZN(n10040) );
  INV_X1 U11932 ( .A(n13165), .ZN(n14177) );
  INV_X1 U11933 ( .A(n10038), .ZN(n13210) );
  INV_X1 U11934 ( .A(n20177), .ZN(n20411) );
  OR2_X1 U11935 ( .A1(n13434), .A2(n20213), .ZN(n20494) );
  AND2_X1 U11936 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20536) );
  AOI21_X1 U11937 ( .B1(P1_STATE2_REG_3__SCAN_IN), .B2(n20703), .A(n20131), 
        .ZN(n20546) );
  INV_X1 U11938 ( .A(n20218), .ZN(n20131) );
  NAND2_X1 U11939 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n20218), .ZN(n20118) );
  NAND2_X1 U11940 ( .A1(n9774), .A2(n9718), .ZN(n15409) );
  NAND2_X1 U11941 ( .A1(n10865), .A2(n9775), .ZN(n9774) );
  AOI21_X1 U11942 ( .B1(n10866), .B2(n11072), .A(n9776), .ZN(n9775) );
  OR2_X1 U11943 ( .A1(n15902), .A2(n18912), .ZN(n15881) );
  INV_X1 U11944 ( .A(n14588), .ZN(n9904) );
  NAND2_X1 U11945 ( .A1(n12304), .A2(n12002), .ZN(n12310) );
  NAND2_X1 U11946 ( .A1(n12305), .A2(n12309), .ZN(n12313) );
  NAND2_X1 U11947 ( .A1(n9904), .A2(n9887), .ZN(n15912) );
  AND2_X1 U11948 ( .A1(n12302), .A2(n12301), .ZN(n14585) );
  NAND2_X1 U11949 ( .A1(n9762), .A2(n12282), .ZN(n12289) );
  AND2_X1 U11950 ( .A1(n12261), .A2(n9709), .ZN(n12264) );
  NAND2_X1 U11951 ( .A1(n12261), .A2(n10072), .ZN(n12245) );
  AND2_X1 U11952 ( .A1(n12240), .A2(n12242), .ZN(n18760) );
  NAND2_X1 U11953 ( .A1(n12247), .A2(n12301), .ZN(n12261) );
  AND2_X1 U11954 ( .A1(n12224), .A2(n9666), .ZN(n12255) );
  NAND2_X1 U11955 ( .A1(n12301), .A2(n12232), .ZN(n12224) );
  AND2_X1 U11956 ( .A1(n12217), .A2(n10058), .ZN(n12223) );
  AND2_X1 U11957 ( .A1(n10064), .A2(n10062), .ZN(n12212) );
  INV_X1 U11958 ( .A(n12165), .ZN(n10062) );
  NOR2_X1 U11959 ( .A1(n12165), .A2(n12166), .ZN(n12147) );
  NOR2_X1 U11960 ( .A1(n12158), .A2(n11993), .ZN(n12153) );
  NAND2_X1 U11961 ( .A1(n12153), .A2(n12152), .ZN(n12165) );
  AND2_X1 U11962 ( .A1(n12547), .A2(n13227), .ZN(n13365) );
  NOR2_X2 U11963 ( .A1(n14663), .A2(n14654), .ZN(n14653) );
  NAND2_X1 U11964 ( .A1(n12710), .A2(n9994), .ZN(n9992) );
  INV_X1 U11965 ( .A(n14628), .ZN(n9994) );
  OR2_X1 U11966 ( .A1(n14689), .A2(n14688), .ZN(n9997) );
  CLKBUF_X1 U11967 ( .A(n14077), .Z(n15936) );
  AND2_X1 U11968 ( .A1(n10017), .A2(n10016), .ZN(n10015) );
  INV_X1 U11969 ( .A(n13710), .ZN(n10016) );
  AND3_X1 U11970 ( .A1(n11930), .A2(n11929), .A3(n11928), .ZN(n16089) );
  NAND2_X1 U11971 ( .A1(n9949), .A2(n12479), .ZN(n9948) );
  INV_X1 U11972 ( .A(n12469), .ZN(n9949) );
  NOR2_X1 U11973 ( .A1(n14759), .A2(n14636), .ZN(n14916) );
  NOR2_X1 U11974 ( .A1(n9907), .A2(n9908), .ZN(n9905) );
  INV_X1 U11975 ( .A(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n9908) );
  NAND2_X1 U11976 ( .A1(n9943), .A2(n9942), .ZN(n14759) );
  INV_X1 U11977 ( .A(n14756), .ZN(n9942) );
  INV_X1 U11978 ( .A(n9943), .ZN(n14757) );
  AND2_X1 U11979 ( .A1(n11223), .A2(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n11224) );
  NAND2_X1 U11980 ( .A1(n11223), .A2(n9665), .ZN(n11222) );
  INV_X1 U11981 ( .A(n14041), .ZN(n9953) );
  INV_X1 U11982 ( .A(n13520), .ZN(n9955) );
  AND2_X1 U11983 ( .A1(n11546), .A2(n11545), .ZN(n13377) );
  NAND2_X1 U11984 ( .A1(n9899), .A2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n9897) );
  NAND2_X1 U11985 ( .A1(n13228), .A2(n15009), .ZN(n15012) );
  INV_X1 U11986 ( .A(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n13017) );
  NAND2_X1 U11987 ( .A1(n11478), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n11490) );
  NAND2_X1 U11988 ( .A1(n12498), .A2(n10081), .ZN(n10080) );
  NOR2_X1 U11989 ( .A1(n14697), .A2(n10082), .ZN(n10081) );
  OR2_X1 U11990 ( .A1(n10054), .A2(n14707), .ZN(n10053) );
  AOI21_X1 U11991 ( .B1(n14585), .B2(n12322), .A(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n14853) );
  NAND2_X1 U11992 ( .A1(n14865), .A2(n14873), .ZN(n10096) );
  OR2_X1 U11993 ( .A1(n12976), .A2(n12292), .ZN(n12293) );
  XNOR2_X1 U11994 ( .A(n12291), .B(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n14879) );
  OR2_X1 U11995 ( .A1(n12976), .A2(n12426), .ZN(n12291) );
  NOR2_X2 U11996 ( .A1(n13708), .A2(n9655), .ZN(n14912) );
  INV_X1 U11997 ( .A(n14078), .ZN(n9916) );
  OR3_X1 U11998 ( .A1(n15306), .A2(n12426), .A3(n14910), .ZN(n14904) );
  NOR2_X1 U11999 ( .A1(n14746), .A2(n14747), .ZN(n14736) );
  NAND2_X1 U12000 ( .A1(n9853), .A2(n9852), .ZN(n9851) );
  INV_X1 U12001 ( .A(n14748), .ZN(n9852) );
  NAND2_X1 U12002 ( .A1(n9855), .A2(n14736), .ZN(n9853) );
  AND2_X1 U12003 ( .A1(n12278), .A2(n15435), .ZN(n14747) );
  NAND2_X1 U12004 ( .A1(n14764), .A2(n14775), .ZN(n14746) );
  NAND2_X1 U12005 ( .A1(n15318), .A2(n14735), .ZN(n14777) );
  NOR2_X1 U12006 ( .A1(n9911), .A2(n9912), .ZN(n9910) );
  INV_X1 U12007 ( .A(n16074), .ZN(n9911) );
  OR3_X1 U12008 ( .A1(n18799), .A2(n12426), .A3(n12269), .ZN(n16009) );
  AOI21_X1 U12009 ( .B1(n9845), .B2(n14728), .A(n9843), .ZN(n9842) );
  INV_X1 U12010 ( .A(n9845), .ZN(n9844) );
  INV_X1 U12011 ( .A(n16019), .ZN(n9843) );
  NOR3_X1 U12012 ( .A1(n14172), .A2(n13520), .A3(n9956), .ZN(n15289) );
  INV_X1 U12013 ( .A(n13720), .ZN(n9956) );
  INV_X1 U12014 ( .A(n16101), .ZN(n9909) );
  NAND2_X1 U12015 ( .A1(n16101), .A2(n14966), .ZN(n16090) );
  AOI21_X1 U12016 ( .B1(n10092), .B2(n10091), .A(n10090), .ZN(n10089) );
  AND3_X1 U12017 ( .A1(n11861), .A2(n11860), .A3(n11859), .ZN(n15003) );
  NAND2_X1 U12018 ( .A1(n16117), .A2(n16115), .ZN(n15028) );
  AOI21_X1 U12019 ( .B1(n10049), .B2(n10051), .A(n9694), .ZN(n10047) );
  AND2_X1 U12020 ( .A1(n12229), .A2(n15029), .ZN(n15023) );
  AND2_X1 U12021 ( .A1(n11538), .A2(n11537), .ZN(n13233) );
  NAND2_X1 U12022 ( .A1(n13825), .A2(n13824), .ZN(n16112) );
  NOR2_X1 U12023 ( .A1(n13244), .A2(n13245), .ZN(n13273) );
  NAND2_X1 U12024 ( .A1(n9962), .A2(n9963), .ZN(n13272) );
  NAND3_X1 U12025 ( .A1(n9781), .A2(n12423), .A3(n9780), .ZN(n13835) );
  NAND2_X1 U12026 ( .A1(n12417), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n13686) );
  AND3_X1 U12027 ( .A1(n11749), .A2(n11748), .A3(n11747), .ZN(n13481) );
  CLKBUF_X1 U12028 ( .A(n13479), .Z(n13549) );
  NAND2_X1 U12029 ( .A1(n10046), .A2(n10045), .ZN(n12410) );
  INV_X1 U12030 ( .A(n13523), .ZN(n10045) );
  AND2_X1 U12031 ( .A1(n11523), .A2(n11522), .ZN(n13085) );
  NAND2_X1 U12032 ( .A1(n12022), .A2(n12023), .ZN(n12027) );
  XNOR2_X1 U12033 ( .A(n15038), .B(n12534), .ZN(n13073) );
  AOI21_X1 U12034 ( .B1(n19130), .B2(n12533), .A(n12532), .ZN(n13072) );
  NAND2_X1 U12035 ( .A1(n12357), .A2(n12356), .ZN(n13635) );
  AND3_X2 U12036 ( .A1(n11402), .A2(n12375), .A3(n11474), .ZN(n13065) );
  AND3_X1 U12037 ( .A1(n9639), .A2(n11450), .A3(n11435), .ZN(n11402) );
  NOR2_X2 U12038 ( .A1(n13571), .A2(n13572), .ZN(n19180) );
  NOR2_X2 U12039 ( .A1(n13118), .A2(n13572), .ZN(n19179) );
  INV_X1 U12040 ( .A(n19180), .ZN(n19163) );
  INV_X1 U12041 ( .A(n19179), .ZN(n19165) );
  NAND2_X1 U12042 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n19593), .ZN(n19176) );
  NOR4_X2 U12043 ( .A1(n15067), .A2(n17082), .A3(n15073), .A4(n18047), .ZN(
        n15069) );
  INV_X1 U12044 ( .A(n18706), .ZN(n18695) );
  NOR2_X1 U12045 ( .A1(n16403), .A2(n16404), .ZN(n16402) );
  NOR2_X1 U12046 ( .A1(n17342), .A2(n16417), .ZN(n16416) );
  NOR2_X1 U12047 ( .A1(n16435), .A2(n10011), .ZN(n16425) );
  NOR2_X1 U12048 ( .A1(n16426), .A2(n16425), .ZN(n16424) );
  NOR2_X1 U12049 ( .A1(n16445), .A2(n16446), .ZN(n16444) );
  NOR2_X1 U12050 ( .A1(n10007), .A2(n10005), .ZN(n16458) );
  NAND2_X1 U12051 ( .A1(n10008), .A2(n10006), .ZN(n10005) );
  OR2_X1 U12052 ( .A1(n16502), .A2(n16679), .ZN(n10003) );
  NOR2_X1 U12053 ( .A1(n16679), .A2(n16381), .ZN(n16503) );
  NOR2_X1 U12054 ( .A1(n16503), .A2(n17458), .ZN(n16502) );
  INV_X1 U12055 ( .A(n17546), .ZN(n17508) );
  OR2_X1 U12056 ( .A1(n17609), .A2(n17532), .ZN(n16606) );
  NOR2_X1 U12057 ( .A1(n17289), .A2(n17226), .ZN(n17255) );
  NAND2_X1 U12058 ( .A1(n10013), .A2(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n10012) );
  INV_X1 U12059 ( .A(n17358), .ZN(n10013) );
  NAND2_X1 U12060 ( .A1(n16369), .A2(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n10014) );
  NOR2_X1 U12061 ( .A1(n17415), .A2(n16471), .ZN(n17389) );
  NAND3_X1 U12062 ( .A1(n17428), .A2(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n17415) );
  NOR2_X1 U12063 ( .A1(n17454), .A2(n17453), .ZN(n17428) );
  NOR2_X1 U12064 ( .A1(n16676), .A2(n16690), .ZN(n17636) );
  NAND2_X1 U12065 ( .A1(n17669), .A2(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n16676) );
  AND2_X1 U12066 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n17669) );
  NAND2_X1 U12067 ( .A1(n17549), .A2(n17707), .ZN(n17427) );
  NOR2_X1 U12068 ( .A1(n15212), .A2(n9975), .ZN(n16163) );
  NAND2_X1 U12069 ( .A1(n9978), .A2(n17711), .ZN(n9975) );
  NOR2_X1 U12070 ( .A1(n9979), .A2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n9978) );
  INV_X1 U12071 ( .A(n15214), .ZN(n9979) );
  NAND2_X1 U12072 ( .A1(n15213), .A2(n9977), .ZN(n9976) );
  INV_X1 U12073 ( .A(n15397), .ZN(n9977) );
  NOR2_X1 U12074 ( .A1(n17347), .A2(n15397), .ZN(n16198) );
  NOR2_X1 U12075 ( .A1(n15397), .A2(n17720), .ZN(n16187) );
  NOR2_X1 U12076 ( .A1(n17751), .A2(n17748), .ZN(n17395) );
  NOR2_X1 U12077 ( .A1(n17748), .A2(n17750), .ZN(n17396) );
  NAND2_X1 U12078 ( .A1(n17411), .A2(n15208), .ZN(n17400) );
  NAND2_X1 U12079 ( .A1(n15207), .A2(n10117), .ZN(n15208) );
  NOR2_X1 U12080 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n15213), .ZN(
        n17482) );
  NAND2_X1 U12081 ( .A1(n15213), .A2(n17840), .ZN(n9981) );
  OR2_X1 U12082 ( .A1(n17501), .A2(n15213), .ZN(n9983) );
  NOR4_X1 U12083 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A4(n17537), .ZN(n17501) );
  NAND2_X1 U12084 ( .A1(n9989), .A2(n9988), .ZN(n17537) );
  NOR2_X1 U12085 ( .A1(n9669), .A2(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n9988) );
  AOI21_X1 U12086 ( .B1(n15238), .B2(n18484), .A(n15237), .ZN(n18493) );
  NOR2_X1 U12087 ( .A1(n15270), .A2(n17612), .ZN(n17875) );
  INV_X1 U12088 ( .A(n16182), .ZN(n17904) );
  NOR2_X1 U12089 ( .A1(n17613), .A2(n17948), .ZN(n17612) );
  INV_X1 U12090 ( .A(n15200), .ZN(n9973) );
  NOR2_X1 U12091 ( .A1(n20912), .A2(n17638), .ZN(n17637) );
  NOR2_X1 U12092 ( .A1(n15253), .A2(n17673), .ZN(n17660) );
  NOR2_X1 U12093 ( .A1(n17675), .A2(n17674), .ZN(n17673) );
  NAND2_X1 U12094 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n17706), .ZN(
        n17705) );
  NAND2_X1 U12095 ( .A1(n15231), .A2(n15082), .ZN(n18483) );
  NOR2_X2 U12096 ( .A1(n13901), .A2(n13900), .ZN(n18068) );
  NOR2_X1 U12097 ( .A1(n13921), .A2(n13920), .ZN(n18071) );
  NOR2_X1 U12098 ( .A1(n15223), .A2(n15087), .ZN(n18520) );
  INV_X1 U12099 ( .A(n19930), .ZN(n15471) );
  NAND2_X1 U12100 ( .A1(n12907), .A2(n12903), .ZN(n19875) );
  INV_X1 U12101 ( .A(n19935), .ZN(n19923) );
  INV_X1 U12102 ( .A(n19875), .ZN(n19920) );
  AND2_X1 U12103 ( .A1(n19922), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n19935) );
  AND2_X1 U12104 ( .A1(n19922), .A2(n13665), .ZN(n19934) );
  AND2_X1 U12105 ( .A1(n19945), .A2(n20117), .ZN(n19940) );
  NAND2_X1 U12106 ( .A1(n14436), .A2(n11090), .ZN(n14437) );
  INV_X1 U12107 ( .A(n15668), .ZN(n15666) );
  OAI21_X1 U12108 ( .B1(n11097), .B2(n11099), .A(n11098), .ZN(n14373) );
  AOI21_X1 U12109 ( .B1(n14312), .B2(n14220), .A(n11097), .ZN(n15563) );
  INV_X1 U12110 ( .A(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n15664) );
  INV_X1 U12111 ( .A(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n19908) );
  NAND2_X1 U12112 ( .A1(n20031), .A2(n11201), .ZN(n20039) );
  AND2_X1 U12113 ( .A1(n15356), .A2(n19826), .ZN(n20042) );
  XNOR2_X1 U12114 ( .A(n12925), .B(n12924), .ZN(n14564) );
  AOI22_X1 U12115 ( .A1(n12923), .A2(n12922), .B1(
        P1_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n14447), .ZN(n12925) );
  OR2_X1 U12116 ( .A1(n14448), .A2(n14447), .ZN(n14449) );
  NAND2_X1 U12117 ( .A1(n9809), .A2(n9807), .ZN(n15561) );
  NOR2_X1 U12118 ( .A1(n15697), .A2(n15559), .ZN(n15689) );
  OAI21_X1 U12119 ( .B1(n14486), .B2(n11190), .A(n15569), .ZN(n15584) );
  INV_X1 U12120 ( .A(n10030), .ZN(n15585) );
  AOI21_X1 U12121 ( .B1(n15418), .B2(n15379), .A(n14559), .ZN(n15719) );
  OR2_X1 U12122 ( .A1(n15650), .A2(n9804), .ZN(n9799) );
  NAND2_X1 U12123 ( .A1(n10043), .A2(n11167), .ZN(n13755) );
  NAND2_X1 U12124 ( .A1(n15650), .A2(n9674), .ZN(n10043) );
  NAND2_X1 U12125 ( .A1(n9790), .A2(n9788), .ZN(n10026) );
  AOI21_X1 U12126 ( .B1(n13494), .B2(n9794), .A(n9671), .ZN(n9790) );
  OAI21_X1 U12127 ( .B1(n20065), .B2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n20073), .ZN(n20046) );
  NAND2_X1 U12128 ( .A1(n15350), .A2(n13413), .ZN(n20066) );
  NOR2_X1 U12129 ( .A1(n15798), .A2(n20047), .ZN(n20060) );
  NAND2_X1 U12130 ( .A1(n9764), .A2(n20050), .ZN(n20073) );
  INV_X1 U12131 ( .A(n13413), .ZN(n9764) );
  INV_X1 U12132 ( .A(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n20703) );
  INV_X1 U12133 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20697) );
  INV_X1 U12134 ( .A(n20702), .ZN(n20706) );
  NOR2_X1 U12135 ( .A1(n14179), .A2(n10039), .ZN(n13215) );
  NAND2_X1 U12136 ( .A1(n13211), .A2(n13210), .ZN(n10039) );
  NOR2_X1 U12137 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n15857) );
  NOR2_X1 U12138 ( .A1(n20494), .A2(n20411), .ZN(n20121) );
  AND2_X1 U12139 ( .A1(n20178), .A2(n20243), .ZN(n20930) );
  INV_X1 U12140 ( .A(n20235), .ZN(n20217) );
  AND2_X1 U12141 ( .A1(n20178), .A2(n20177), .ZN(n20235) );
  OAI211_X1 U12142 ( .C1(n10121), .C2(n20440), .A(n20377), .B(n20331), .ZN(
        n20348) );
  OAI22_X1 U12143 ( .A1(n20382), .A2(n20491), .B1(n20381), .B2(n20380), .ZN(
        n20399) );
  NOR2_X1 U12144 ( .A1(n20681), .A2(n20411), .ZN(n20436) );
  NOR2_X1 U12145 ( .A1(n12988), .A2(n13641), .ZN(n19804) );
  NOR2_X1 U12146 ( .A1(n18924), .A2(n9945), .ZN(n9944) );
  AOI21_X1 U12147 ( .B1(n9904), .B2(n9887), .A(n9900), .ZN(n15902) );
  INV_X1 U12148 ( .A(n9901), .ZN(n9900) );
  AOI21_X1 U12149 ( .B1(n9887), .B2(n9902), .A(n15904), .ZN(n9901) );
  INV_X1 U12150 ( .A(n9903), .ZN(n15903) );
  OAI21_X1 U12151 ( .B1(n9904), .B2(n9902), .A(n9887), .ZN(n9903) );
  AND2_X1 U12152 ( .A1(n12306), .A2(n12329), .ZN(n15909) );
  OR2_X1 U12153 ( .A1(n9887), .A2(n15977), .ZN(n9884) );
  NAND2_X1 U12154 ( .A1(n9886), .A2(n11218), .ZN(n9885) );
  AND2_X1 U12155 ( .A1(n9883), .A2(n9887), .ZN(n12974) );
  OR2_X1 U12156 ( .A1(n18735), .A2(n15985), .ZN(n9883) );
  AND2_X1 U12157 ( .A1(n18735), .A2(n9887), .ZN(n15305) );
  AND2_X1 U12158 ( .A1(n9890), .A2(n18831), .ZN(n18753) );
  NAND2_X1 U12159 ( .A1(n9888), .A2(n9889), .ZN(n18752) );
  NAND2_X1 U12160 ( .A1(n12217), .A2(n11429), .ZN(n12218) );
  NAND2_X1 U12161 ( .A1(n13516), .A2(n13719), .ZN(n18941) );
  INV_X1 U12162 ( .A(n19767), .ZN(n18999) );
  NAND2_X1 U12163 ( .A1(n15948), .A2(n9639), .ZN(n18952) );
  CLKBUF_X1 U12164 ( .A(n15948), .Z(n18958) );
  OR2_X1 U12165 ( .A1(n13708), .A2(n9707), .ZN(n15437) );
  AND2_X1 U12166 ( .A1(n13038), .A2(n13331), .ZN(n18965) );
  AND2_X1 U12167 ( .A1(n13038), .A2(n13571), .ZN(n18964) );
  NOR2_X1 U12168 ( .A1(n19031), .A2(n19027), .ZN(n19006) );
  NOR2_X1 U12169 ( .A1(n10001), .A2(n13234), .ZN(n10000) );
  AND2_X1 U12170 ( .A1(n13078), .A2(n12541), .ZN(n10002) );
  INV_X1 U12171 ( .A(n19002), .ZN(n19031) );
  NAND2_X1 U12172 ( .A1(n9895), .A2(n11220), .ZN(n9891) );
  AOI21_X1 U12173 ( .B1(n12947), .B2(n14610), .A(n12946), .ZN(n15892) );
  OR2_X1 U12174 ( .A1(n12963), .A2(n19087), .ZN(n12964) );
  NAND2_X1 U12175 ( .A1(n9847), .A2(n9848), .ZN(n16022) );
  NAND2_X1 U12176 ( .A1(n14726), .A2(n9850), .ZN(n9847) );
  INV_X1 U12177 ( .A(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n19094) );
  AND2_X1 U12178 ( .A1(n19093), .A2(n14166), .ZN(n19080) );
  INV_X1 U12179 ( .A(n16068), .ZN(n19087) );
  INV_X1 U12180 ( .A(n19088), .ZN(n16066) );
  AND2_X1 U12181 ( .A1(n19093), .A2(n19766), .ZN(n19090) );
  INV_X1 U12182 ( .A(n19090), .ZN(n16072) );
  OAI21_X1 U12183 ( .B1(n12939), .B2(n14706), .A(n9862), .ZN(n9860) );
  OR2_X1 U12184 ( .A1(n14861), .A2(n12489), .ZN(n14836) );
  INV_X1 U12185 ( .A(n12936), .ZN(n14718) );
  INV_X1 U12186 ( .A(n16083), .ZN(n16107) );
  NAND2_X1 U12187 ( .A1(n13816), .A2(n12430), .ZN(n14794) );
  NOR2_X1 U12188 ( .A1(n12481), .A2(n13633), .ZN(n19116) );
  INV_X1 U12189 ( .A(n19112), .ZN(n19131) );
  INV_X1 U12190 ( .A(n19137), .ZN(n19779) );
  INV_X1 U12191 ( .A(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n19764) );
  XNOR2_X1 U12192 ( .A(n13073), .B(n13072), .ZN(n19767) );
  XNOR2_X1 U12193 ( .A(n13068), .B(n10128), .ZN(n19138) );
  INV_X1 U12194 ( .A(n19246), .ZN(n19238) );
  NOR2_X1 U12195 ( .A1(n19342), .A2(n19459), .ZN(n19276) );
  OAI21_X1 U12196 ( .B1(n19327), .B2(n19594), .A(n19311), .ZN(n19329) );
  NOR2_X1 U12197 ( .A1(n19587), .A2(n19307), .ZN(n19360) );
  NOR2_X1 U12198 ( .A1(n19342), .A2(n19587), .ZN(n19386) );
  OAI21_X1 U12199 ( .B1(n19389), .B2(n19368), .A(n19593), .ZN(n19391) );
  NOR2_X1 U12200 ( .A1(n19555), .A2(n19395), .ZN(n19419) );
  OAI21_X1 U12201 ( .B1(n19432), .B2(n19448), .A(n19593), .ZN(n19450) );
  NOR2_X1 U12202 ( .A1(n19534), .A2(n19459), .ZN(n19493) );
  INV_X1 U12203 ( .A(n19515), .ZN(n19634) );
  INV_X1 U12204 ( .A(n19478), .ZN(n19635) );
  INV_X1 U12205 ( .A(n19424), .ZN(n19651) );
  AOI21_X1 U12206 ( .B1(n18484), .B2(n18483), .A(n17289), .ZN(n18707) );
  OR2_X1 U12207 ( .A1(P3_STATE_REG_0__SCAN_IN), .A2(n18559), .ZN(n18701) );
  OAI21_X1 U12208 ( .B1(n16445), .B2(n10020), .A(n10019), .ZN(n16435) );
  NAND2_X1 U12209 ( .A1(n10021), .A2(n17393), .ZN(n10020) );
  NAND2_X1 U12210 ( .A1(n10011), .A2(n10021), .ZN(n10019) );
  INV_X1 U12211 ( .A(n17382), .ZN(n10021) );
  NOR2_X1 U12212 ( .A1(n16444), .A2(n10011), .ZN(n16436) );
  NAND2_X1 U12213 ( .A1(n10004), .A2(n10008), .ZN(n16465) );
  NOR2_X1 U12214 ( .A1(n16479), .A2(n10011), .ZN(n16466) );
  AND2_X1 U12215 ( .A1(n10003), .A2(n17441), .ZN(n16492) );
  INV_X1 U12216 ( .A(n10003), .ZN(n16493) );
  INV_X1 U12217 ( .A(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n16690) );
  INV_X1 U12218 ( .A(n16722), .ZN(n16752) );
  AND2_X1 U12219 ( .A1(P3_EBX_REG_23__SCAN_IN), .A2(n16816), .ZN(n16821) );
  NAND4_X1 U12220 ( .A1(P3_EBX_REG_7__SCAN_IN), .A2(P3_EBX_REG_6__SCAN_IN), 
        .A3(P3_EBX_REG_5__SCAN_IN), .A4(n17044), .ZN(n17032) );
  NOR2_X1 U12221 ( .A1(n17232), .A2(n17097), .ZN(n17092) );
  NAND2_X1 U12222 ( .A1(P3_EAX_REG_27__SCAN_IN), .A2(n17102), .ZN(n17097) );
  NOR2_X1 U12223 ( .A1(n17235), .A2(n17106), .ZN(n17102) );
  NAND2_X1 U12224 ( .A1(P3_EAX_REG_25__SCAN_IN), .A2(n17107), .ZN(n17106) );
  NOR2_X1 U12225 ( .A1(n17123), .A2(n17117), .ZN(n17113) );
  NOR3_X1 U12226 ( .A1(n17123), .A2(n17154), .A3(n17294), .ZN(n17146) );
  NAND2_X1 U12227 ( .A1(P3_EAX_REG_16__SCAN_IN), .A2(n17158), .ZN(n17154) );
  NOR2_X1 U12228 ( .A1(n17339), .A2(n17163), .ZN(n17158) );
  NOR2_X1 U12229 ( .A1(n15112), .A2(n15111), .ZN(n17201) );
  INV_X1 U12230 ( .A(n15254), .ZN(n17205) );
  NOR2_X1 U12231 ( .A1(n15122), .A2(n15121), .ZN(n17208) );
  NAND2_X1 U12232 ( .A1(n13962), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n15144) );
  NOR2_X2 U12233 ( .A1(n13868), .A2(n13867), .ZN(n18087) );
  NOR2_X1 U12234 ( .A1(n17213), .A2(n18511), .ZN(n17222) );
  INV_X1 U12235 ( .A(n17214), .ZN(n17221) );
  NOR2_X1 U12236 ( .A1(n17285), .A2(n17255), .ZN(n17278) );
  CLKBUF_X1 U12237 ( .A(n17278), .Z(n17284) );
  NOR2_X1 U12238 ( .A1(n17291), .A2(n17335), .ZN(n17322) );
  INV_X1 U12239 ( .A(n17322), .ZN(n17338) );
  AOI21_X1 U12240 ( .B1(n17343), .B2(n17356), .A(n17355), .ZN(n17361) );
  INV_X1 U12241 ( .A(n17565), .ZN(n17518) );
  NAND2_X1 U12242 ( .A1(n17503), .A2(n9719), .ZN(n17489) );
  NOR2_X1 U12243 ( .A1(n16182), .A2(n17820), .ZN(n17846) );
  INV_X1 U12244 ( .A(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n17550) );
  INV_X1 U12245 ( .A(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n17568) );
  INV_X1 U12246 ( .A(n17598), .ZN(n17583) );
  INV_X1 U12247 ( .A(n17617), .ZN(n17605) );
  INV_X1 U12248 ( .A(n18078), .ZN(n18426) );
  INV_X1 U12249 ( .A(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n17679) );
  INV_X1 U12250 ( .A(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n17694) );
  INV_X1 U12251 ( .A(n17697), .ZN(n17710) );
  NAND2_X1 U12252 ( .A1(n17364), .A2(n15214), .ZN(n15393) );
  NAND2_X1 U12253 ( .A1(n9989), .A2(n9991), .ZN(n17574) );
  NOR2_X1 U12254 ( .A1(n17649), .A2(n15196), .ZN(n17643) );
  NOR2_X1 U12255 ( .A1(n17667), .A2(n17666), .ZN(n17665) );
  AND2_X1 U12256 ( .A1(n9987), .A2(n9653), .ZN(n17667) );
  NOR2_X1 U12257 ( .A1(n18486), .A2(n18019), .ZN(n17999) );
  INV_X1 U12258 ( .A(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n18522) );
  INV_X1 U12259 ( .A(n20083), .ZN(n20085) );
  NAND2_X1 U12261 ( .A1(n12918), .A2(n19872), .ZN(n12917) );
  NAND2_X1 U12262 ( .A1(n15572), .A2(n19941), .ZN(n10969) );
  AOI22_X1 U12263 ( .A1(n15668), .A2(n20078), .B1(n20064), .B2(n15667), .ZN(
        n15670) );
  INV_X1 U12264 ( .A(n9816), .ZN(n15684) );
  NAND2_X1 U12265 ( .A1(n9875), .A2(n18920), .ZN(n9874) );
  AOI21_X1 U12266 ( .B1(n14566), .B2(n14565), .A(n18890), .ZN(n14567) );
  INV_X1 U12267 ( .A(n12493), .ZN(n12494) );
  OAI21_X1 U12268 ( .B1(n14815), .B2(n16128), .A(n9920), .ZN(n14823) );
  AOI21_X1 U12269 ( .B1(n10023), .B2(n16697), .A(n10022), .ZN(n16400) );
  OR2_X1 U12270 ( .A1(n16397), .A2(n16396), .ZN(n10022) );
  AND2_X1 U12271 ( .A1(n16176), .A2(n16177), .ZN(n9968) );
  NAND2_X1 U12272 ( .A1(n16232), .A2(n18028), .ZN(n16245) );
  INV_X1 U12273 ( .A(n18831), .ZN(n18912) );
  AND2_X1 U12274 ( .A1(n9668), .A2(n9876), .ZN(n9651) );
  CLKBUF_X3 U12275 ( .A(n15106), .Z(n16992) );
  OR2_X1 U12276 ( .A1(n15190), .A2(n15189), .ZN(n9653) );
  AND2_X2 U12277 ( .A1(n12355), .A2(n19796), .ZN(n9654) );
  INV_X1 U12278 ( .A(n11391), .ZN(n11643) );
  INV_X2 U12279 ( .A(n11643), .ZN(n13593) );
  NAND2_X1 U12280 ( .A1(n14252), .A2(n9704), .ZN(n14240) );
  OR2_X1 U12281 ( .A1(n9708), .A2(n9916), .ZN(n9655) );
  NOR2_X1 U12282 ( .A1(n13708), .A2(n9708), .ZN(n9656) );
  AND2_X1 U12283 ( .A1(n9914), .A2(n13824), .ZN(n9658) );
  AOI21_X1 U12284 ( .B1(n10041), .B2(n9803), .A(n9693), .ZN(n9802) );
  NOR2_X1 U12285 ( .A1(n12165), .A2(n9715), .ZN(n12145) );
  AND2_X1 U12286 ( .A1(n10197), .A2(n10196), .ZN(n9659) );
  NAND2_X1 U12287 ( .A1(n15019), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n15021) );
  INV_X1 U12288 ( .A(n15021), .ZN(n9786) );
  AND2_X1 U12289 ( .A1(n15000), .A2(n10098), .ZN(n9660) );
  NAND2_X1 U12290 ( .A1(n15919), .A2(n12322), .ZN(n14865) );
  INV_X1 U12291 ( .A(n14865), .ZN(n10097) );
  NOR3_X1 U12292 ( .A1(n12321), .A2(n12426), .A3(n12490), .ZN(n9661) );
  NAND2_X1 U12293 ( .A1(n9941), .A2(n10313), .ZN(n11115) );
  AND2_X1 U12294 ( .A1(n9658), .A2(n13532), .ZN(n9662) );
  NAND2_X1 U12295 ( .A1(n13424), .A2(n9798), .ZN(n13312) );
  NOR2_X1 U12296 ( .A1(n11214), .A2(n9720), .ZN(n9899) );
  OR2_X1 U12297 ( .A1(n20025), .A2(n20096), .ZN(n9664) );
  NAND2_X1 U12298 ( .A1(n11236), .A2(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n11234) );
  NAND2_X1 U12299 ( .A1(n9896), .A2(n9899), .ZN(n11230) );
  AND2_X1 U12300 ( .A1(n11226), .A2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n11223) );
  AND2_X1 U12301 ( .A1(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n9665) );
  OR2_X1 U12302 ( .A1(n10831), .A2(n10830), .ZN(n11068) );
  AND2_X1 U12303 ( .A1(n12231), .A2(n9738), .ZN(n9666) );
  AND2_X1 U12304 ( .A1(n9938), .A2(n14324), .ZN(n9667) );
  NAND2_X1 U12305 ( .A1(n9887), .A2(n15875), .ZN(n9668) );
  INV_X4 U12306 ( .A(n11635), .ZN(n19796) );
  NOR2_X1 U12307 ( .A1(n11249), .A2(n15895), .ZN(n11250) );
  INV_X1 U12308 ( .A(n14721), .ZN(n9902) );
  NAND2_X1 U12309 ( .A1(n9991), .A2(n9990), .ZN(n9669) );
  NOR2_X2 U12310 ( .A1(n10881), .A2(n10268), .ZN(n9833) );
  AND2_X2 U12311 ( .A1(n12845), .A2(n11278), .ZN(n11788) );
  AND2_X1 U12312 ( .A1(n11153), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n9671) );
  OR3_X1 U12313 ( .A1(n17415), .A2(n10014), .A3(n10012), .ZN(n9672) );
  CLKBUF_X1 U12314 ( .A(n11281), .Z(n12838) );
  AND2_X1 U12315 ( .A1(n9607), .A2(n11468), .ZN(n12018) );
  NAND2_X1 U12316 ( .A1(n12301), .A2(n11996), .ZN(n12217) );
  NAND2_X2 U12317 ( .A1(n12449), .A2(n9654), .ZN(n12475) );
  AND2_X1 U12318 ( .A1(n14252), .A2(n14255), .ZN(n14253) );
  NAND2_X1 U12319 ( .A1(n14678), .A2(n14584), .ZN(n14583) );
  OR2_X1 U12320 ( .A1(n15649), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n9674) );
  NOR2_X1 U12321 ( .A1(n14632), .A2(n14631), .ZN(n14580) );
  INV_X2 U12322 ( .A(n11173), .ZN(n15640) );
  INV_X1 U12323 ( .A(n15621), .ZN(n15569) );
  AND2_X1 U12324 ( .A1(n14241), .A2(n10762), .ZN(n14326) );
  NAND2_X1 U12325 ( .A1(n9856), .A2(n18891), .ZN(n12205) );
  AND2_X1 U12326 ( .A1(n14252), .A2(n9931), .ZN(n14347) );
  NAND2_X1 U12327 ( .A1(n12018), .A2(n12027), .ZN(n12017) );
  AND4_X1 U12328 ( .A1(n10151), .A2(n10150), .A3(n10149), .A4(n10148), .ZN(
        n9675) );
  AND2_X1 U12329 ( .A1(n10027), .A2(n10281), .ZN(n9676) );
  AND2_X1 U12330 ( .A1(n10139), .A2(n10143), .ZN(n10226) );
  AND3_X1 U12331 ( .A1(n9869), .A2(n11347), .A3(n9868), .ZN(n9677) );
  OR2_X1 U12332 ( .A1(n12475), .A2(n11988), .ZN(n9678) );
  OR2_X1 U12333 ( .A1(n14225), .A2(n9830), .ZN(n9679) );
  NAND2_X1 U12334 ( .A1(n10100), .A2(n12215), .ZN(n15022) );
  NAND2_X1 U12335 ( .A1(n12294), .A2(n12293), .ZN(n14864) );
  AND2_X2 U12336 ( .A1(n11658), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11391) );
  AND2_X1 U12337 ( .A1(n14580), .A2(n14581), .ZN(n14579) );
  NAND2_X1 U12338 ( .A1(n11436), .A2(n11435), .ZN(n11474) );
  AND4_X1 U12339 ( .A1(n10175), .A2(n10174), .A3(n10173), .A4(n10172), .ZN(
        n9680) );
  NAND2_X1 U12340 ( .A1(n12045), .A2(n12030), .ZN(n12117) );
  AND4_X1 U12341 ( .A1(n10195), .A2(n10194), .A3(n10193), .A4(n10192), .ZN(
        n9681) );
  AND3_X1 U12342 ( .A1(n10145), .A2(n10147), .A3(n10144), .ZN(n9682) );
  AND2_X1 U12343 ( .A1(n15639), .A2(n11176), .ZN(n14499) );
  OR2_X1 U12344 ( .A1(n18835), .A2(n12235), .ZN(n9683) );
  AND2_X1 U12345 ( .A1(n10100), .A2(n10098), .ZN(n14997) );
  INV_X1 U12346 ( .A(n10400), .ZN(n9820) );
  OR2_X1 U12347 ( .A1(n11482), .A2(n11481), .ZN(n9684) );
  AND2_X1 U12348 ( .A1(n14777), .A2(n9854), .ZN(n9685) );
  INV_X1 U12349 ( .A(n11991), .ZN(n12463) );
  NAND2_X1 U12350 ( .A1(n10100), .A2(n9660), .ZN(n14975) );
  OR2_X1 U12351 ( .A1(n15621), .A2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n9686) );
  AND2_X1 U12352 ( .A1(n13753), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n9687) );
  AND2_X1 U12353 ( .A1(n12542), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n9688) );
  OR2_X1 U12354 ( .A1(n17980), .A2(n15192), .ZN(n9689) );
  NOR2_X1 U12355 ( .A1(n14880), .A2(n10055), .ZN(n14713) );
  OR2_X1 U12356 ( .A1(n15210), .A2(n17615), .ZN(n9690) );
  AND4_X1 U12357 ( .A1(n11746), .A2(n11745), .A3(n11744), .A4(n11743), .ZN(
        n9691) );
  AND2_X1 U12358 ( .A1(n11420), .A2(n11401), .ZN(n9692) );
  INV_X1 U12359 ( .A(n9865), .ZN(n9864) );
  NAND2_X1 U12360 ( .A1(n10096), .A2(n9866), .ZN(n9865) );
  NOR2_X1 U12361 ( .A1(n11320), .A2(n11319), .ZN(n11411) );
  AND2_X1 U12362 ( .A1(n11174), .A2(n15841), .ZN(n9693) );
  INV_X1 U12363 ( .A(n10052), .ZN(n14714) );
  NOR2_X1 U12364 ( .A1(n14880), .A2(n10054), .ZN(n10052) );
  AND2_X1 U12365 ( .A1(n12432), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n9694) );
  NAND2_X1 U12366 ( .A1(n10033), .A2(n10032), .ZN(n9695) );
  NAND2_X1 U12367 ( .A1(n14580), .A2(n9967), .ZN(n14609) );
  NAND2_X1 U12368 ( .A1(n10868), .A2(n13389), .ZN(n9696) );
  NAND2_X1 U12369 ( .A1(n9867), .A2(n10096), .ZN(n14851) );
  NAND2_X1 U12370 ( .A1(n14726), .A2(n14727), .ZN(n16034) );
  AND3_X1 U12371 ( .A1(n11392), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A3(
        n11394), .ZN(n9697) );
  BUF_X1 U12372 ( .A(n11435), .Z(n19156) );
  AND2_X1 U12373 ( .A1(n14777), .A2(n14774), .ZN(n9698) );
  AND2_X1 U12374 ( .A1(n9867), .A2(n9864), .ZN(n9699) );
  INV_X1 U12375 ( .A(n11145), .ZN(n9794) );
  INV_X1 U12376 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10134) );
  AND2_X1 U12377 ( .A1(n14727), .A2(n9683), .ZN(n10092) );
  INV_X1 U12378 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11347) );
  OR2_X2 U12379 ( .A1(n20096), .A2(n20086), .ZN(n10881) );
  NAND2_X1 U12380 ( .A1(n11803), .A2(n11802), .ZN(n13825) );
  NOR2_X1 U12381 ( .A1(n15546), .A2(n15545), .ZN(n9700) );
  NOR2_X1 U12382 ( .A1(n9909), .A2(n9912), .ZN(n16073) );
  AND2_X1 U12383 ( .A1(n13825), .A2(n9658), .ZN(n9701) );
  AND2_X1 U12384 ( .A1(n9605), .A2(n9935), .ZN(n9702) );
  NOR2_X1 U12385 ( .A1(n15230), .A2(n9669), .ZN(n17556) );
  NAND2_X1 U12386 ( .A1(n13739), .A2(n13845), .ZN(n13844) );
  NOR2_X1 U12387 ( .A1(n14172), .A2(n13520), .ZN(n13519) );
  NOR2_X1 U12388 ( .A1(n11234), .A2(n19094), .ZN(n11235) );
  NOR2_X1 U12389 ( .A1(n15230), .A2(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n17585) );
  NOR2_X1 U12390 ( .A1(n9897), .A2(n11233), .ZN(n11231) );
  AND2_X1 U12391 ( .A1(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n11236) );
  NAND2_X1 U12392 ( .A1(n14912), .A2(n14913), .ZN(n12980) );
  INV_X1 U12393 ( .A(n16035), .ZN(n10090) );
  NAND2_X1 U12394 ( .A1(n17193), .A2(n10125), .ZN(n17615) );
  AND2_X1 U12395 ( .A1(n15543), .A2(n14097), .ZN(n9703) );
  AND2_X1 U12396 ( .A1(n9931), .A2(n14348), .ZN(n9704) );
  AND2_X1 U12397 ( .A1(n9666), .A2(n11998), .ZN(n9705) );
  AND2_X1 U12398 ( .A1(n13337), .A2(n13338), .ZN(n13336) );
  AND2_X1 U12399 ( .A1(n13336), .A2(n13373), .ZN(n13372) );
  AND2_X1 U12400 ( .A1(n13580), .A2(n13581), .ZN(n13579) );
  AND2_X1 U12401 ( .A1(n9605), .A2(n9932), .ZN(n9706) );
  NOR2_X1 U12402 ( .A1(n11233), .A2(n11214), .ZN(n11232) );
  OR2_X1 U12403 ( .A1(n11954), .A2(n9915), .ZN(n9707) );
  OR2_X1 U12404 ( .A1(n9707), .A2(n15438), .ZN(n9708) );
  INV_X1 U12405 ( .A(n12211), .ZN(n10061) );
  AND2_X1 U12406 ( .A1(n10072), .A2(n11572), .ZN(n9709) );
  AND2_X1 U12407 ( .A1(n13361), .A2(n13362), .ZN(n13360) );
  NOR2_X1 U12408 ( .A1(n14172), .A2(n9952), .ZN(n14042) );
  OR3_X1 U12409 ( .A1(n14172), .A2(n9957), .A3(n13520), .ZN(n9710) );
  AND2_X1 U12410 ( .A1(n14789), .A2(n14786), .ZN(n9711) );
  AND2_X1 U12411 ( .A1(n15912), .A2(n14721), .ZN(n9712) );
  NOR2_X1 U12412 ( .A1(n13708), .A2(n11954), .ZN(n13734) );
  AND2_X1 U12413 ( .A1(n10861), .A2(n11070), .ZN(n9713) );
  NAND2_X1 U12414 ( .A1(n15620), .A2(n11177), .ZN(n9714) );
  NAND2_X1 U12415 ( .A1(n12527), .A2(n12539), .ZN(n13068) );
  AND2_X1 U12416 ( .A1(n10849), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n10862) );
  INV_X1 U12417 ( .A(n10105), .ZN(n10091) );
  OR2_X1 U12418 ( .A1(n12166), .A2(n10063), .ZN(n9715) );
  NAND2_X1 U12419 ( .A1(n11235), .A2(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n11233) );
  AND2_X1 U12420 ( .A1(n9703), .A2(n9832), .ZN(n9716) );
  AND2_X1 U12421 ( .A1(n9709), .A2(n14637), .ZN(n9717) );
  NAND2_X1 U12422 ( .A1(n11072), .A2(n10867), .ZN(n9718) );
  AND2_X1 U12423 ( .A1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n9719) );
  NAND2_X1 U12424 ( .A1(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n9720) );
  INV_X1 U12425 ( .A(n9907), .ZN(n9906) );
  NAND2_X1 U12426 ( .A1(n9665), .A2(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n9907) );
  NAND2_X1 U12427 ( .A1(n14916), .A2(n14915), .ZN(n12977) );
  AND2_X1 U12428 ( .A1(n10990), .A2(n14327), .ZN(n9721) );
  INV_X1 U12429 ( .A(n9855), .ZN(n9854) );
  NAND2_X1 U12430 ( .A1(n14765), .A2(n14774), .ZN(n9855) );
  OR2_X1 U12431 ( .A1(n11123), .A2(n10839), .ZN(n9722) );
  OR2_X1 U12432 ( .A1(n14353), .A2(n10946), .ZN(n9723) );
  AND2_X1 U12433 ( .A1(n14736), .A2(n14735), .ZN(n9724) );
  NOR2_X1 U12434 ( .A1(n15305), .A2(n15985), .ZN(n9725) );
  AND2_X1 U12435 ( .A1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n9726) );
  AND2_X1 U12436 ( .A1(n9704), .A2(n9930), .ZN(n9727) );
  AND2_X1 U12437 ( .A1(n9997), .A2(n9996), .ZN(n9728) );
  AND2_X1 U12438 ( .A1(n9660), .A2(n10105), .ZN(n9729) );
  AND2_X1 U12439 ( .A1(n9705), .A2(n11557), .ZN(n9730) );
  AND2_X1 U12440 ( .A1(n9981), .A2(n9980), .ZN(n9731) );
  NAND3_X1 U12441 ( .A1(n10855), .A2(n10838), .A3(n10856), .ZN(n9732) );
  AND2_X1 U12442 ( .A1(n9721), .A2(n9667), .ZN(n9733) );
  INV_X1 U12443 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n9778) );
  AND2_X1 U12444 ( .A1(n13413), .A2(n13398), .ZN(n20078) );
  NOR2_X1 U12445 ( .A1(n13479), .A2(n13481), .ZN(n13480) );
  NOR2_X1 U12446 ( .A1(n11227), .A2(n11216), .ZN(n11226) );
  NOR2_X1 U12447 ( .A1(n11219), .A2(n15984), .ZN(n11246) );
  NAND2_X1 U12448 ( .A1(n11250), .A2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n9734) );
  OR3_X1 U12449 ( .A1(n17415), .A2(n10014), .A3(n17358), .ZN(n9736) );
  AND2_X1 U12450 ( .A1(n9967), .A2(n9966), .ZN(n9737) );
  NOR2_X1 U12451 ( .A1(n15012), .A2(n13377), .ZN(n13361) );
  NAND2_X1 U12452 ( .A1(n13516), .A2(n10017), .ZN(n13709) );
  INV_X1 U12453 ( .A(n12260), .ZN(n10073) );
  OR2_X1 U12454 ( .A1(n12003), .A2(n11552), .ZN(n9738) );
  NAND2_X1 U12455 ( .A1(n13675), .A2(n11782), .ZN(n14047) );
  AND2_X1 U12456 ( .A1(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n9739) );
  NOR2_X1 U12457 ( .A1(n12544), .A2(n13241), .ZN(n9740) );
  XNOR2_X1 U12458 ( .A(n9974), .B(n9973), .ZN(n17630) );
  NOR2_X1 U12459 ( .A1(n17643), .A2(n17642), .ZN(n17641) );
  AND2_X1 U12460 ( .A1(n10358), .A2(n10379), .ZN(n9741) );
  AND2_X1 U12461 ( .A1(n9737), .A2(n9965), .ZN(n9742) );
  INV_X1 U12462 ( .A(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n20690) );
  INV_X1 U12463 ( .A(P1_STATE2_REG_0__SCAN_IN), .ZN(n20597) );
  OR2_X1 U12464 ( .A1(n18754), .A2(n14769), .ZN(n9743) );
  INV_X1 U12465 ( .A(n9895), .ZN(n9894) );
  NAND2_X1 U12466 ( .A1(n9739), .A2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n9895) );
  AND2_X1 U12467 ( .A1(n11223), .A2(n9906), .ZN(n9744) );
  AND2_X1 U12468 ( .A1(n9932), .A2(n14116), .ZN(n9745) );
  AND2_X1 U12469 ( .A1(n9962), .A2(n9960), .ZN(n9746) );
  AND2_X1 U12470 ( .A1(n10058), .A2(n11541), .ZN(n9747) );
  INV_X1 U12471 ( .A(P2_EBX_REG_10__SCAN_IN), .ZN(n10059) );
  INV_X1 U12472 ( .A(n17431), .ZN(n10010) );
  NOR2_X1 U12473 ( .A1(n11247), .A2(n15960), .ZN(n11248) );
  INV_X1 U12474 ( .A(n10268), .ZN(n10878) );
  AND2_X1 U12475 ( .A1(n11432), .A2(n11431), .ZN(n9748) );
  NAND2_X1 U12476 ( .A1(n9827), .A2(n9826), .ZN(n13334) );
  INV_X1 U12477 ( .A(n13334), .ZN(n9825) );
  OR2_X1 U12478 ( .A1(n17415), .A2(n10014), .ZN(n9749) );
  INV_X1 U12479 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n9925) );
  NOR2_X1 U12480 ( .A1(n20433), .A2(n20264), .ZN(n9750) );
  NOR2_X1 U12481 ( .A1(n20433), .A2(n20539), .ZN(n9751) );
  INV_X1 U12482 ( .A(n15645), .ZN(n20084) );
  AND2_X1 U12483 ( .A1(n11100), .A2(n20700), .ZN(n15645) );
  INV_X1 U12484 ( .A(n14985), .ZN(n9785) );
  INV_X1 U12485 ( .A(P2_EBX_REG_24__SCAN_IN), .ZN(n10056) );
  INV_X1 U12486 ( .A(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n9990) );
  INV_X1 U12487 ( .A(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n9980) );
  INV_X1 U12488 ( .A(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n10035) );
  NOR3_X2 U12489 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20703), .A3(
        n20539), .ZN(n20486) );
  NOR3_X2 U12490 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20703), .A3(
        n20185), .ZN(n20925) );
  INV_X1 U12491 ( .A(n9664), .ZN(n9752) );
  NOR4_X4 U12492 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(P3_STATE2_REG_0__SCAN_IN), .A3(P3_STATEBS16_REG_SCAN_IN), .A4(n18650), .ZN(n16697) );
  AND2_X1 U12493 ( .A1(n20000), .A2(n20096), .ZN(n9753) );
  NOR2_X2 U12494 ( .A1(n12936), .A2(n12937), .ZN(n12934) );
  AOI21_X1 U12495 ( .B1(n9757), .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n9756), .ZN(n9755) );
  OAI21_X1 U12496 ( .B1(n12936), .B2(n14707), .A(n9758), .ZN(n9757) );
  NAND2_X1 U12497 ( .A1(n12404), .A2(n12463), .ZN(n9759) );
  NAND3_X1 U12498 ( .A1(n11696), .A2(n11697), .A3(n11695), .ZN(n9761) );
  NAND2_X1 U12499 ( .A1(n12284), .A2(n12301), .ZN(n9762) );
  NAND3_X1 U12500 ( .A1(n9770), .A2(n9732), .A3(n9769), .ZN(n9768) );
  NAND2_X2 U12501 ( .A1(n9681), .A2(n9657), .ZN(n13410) );
  NAND2_X1 U12502 ( .A1(n12416), .A2(n12415), .ZN(n13683) );
  NAND3_X1 U12503 ( .A1(n13683), .A2(n13684), .A3(n12420), .ZN(n9780) );
  NAND2_X1 U12504 ( .A1(n10109), .A2(n13682), .ZN(n9781) );
  AND2_X2 U12505 ( .A1(n9784), .A2(n9782), .ZN(n12016) );
  NAND3_X1 U12506 ( .A1(n11491), .A2(n12022), .A3(n12023), .ZN(n9784) );
  AND2_X2 U12507 ( .A1(n12071), .A2(n12070), .ZN(n12151) );
  NAND2_X1 U12508 ( .A1(n12101), .A2(n12100), .ZN(n12150) );
  NOR2_X2 U12509 ( .A1(n16017), .A2(n12269), .ZN(n16013) );
  NAND2_X1 U12510 ( .A1(n13350), .A2(n13349), .ZN(n11137) );
  NAND3_X1 U12511 ( .A1(n9792), .A2(n15656), .A3(n9791), .ZN(n11166) );
  OR2_X1 U12512 ( .A1(n13494), .A2(n9671), .ZN(n9791) );
  NAND3_X1 U12513 ( .A1(n11146), .A2(n11145), .A3(n9793), .ZN(n9792) );
  NAND2_X1 U12514 ( .A1(n11146), .A2(n11145), .ZN(n13495) );
  NAND2_X1 U12515 ( .A1(n9796), .A2(n9722), .ZN(n9812) );
  NAND3_X1 U12516 ( .A1(n13424), .A2(n20597), .A3(n9798), .ZN(n9796) );
  NAND2_X2 U12517 ( .A1(n9797), .A2(n10285), .ZN(n13424) );
  NAND2_X1 U12518 ( .A1(n9799), .A2(n9802), .ZN(n14036) );
  NAND2_X1 U12519 ( .A1(n9802), .A2(n9804), .ZN(n9800) );
  NAND2_X1 U12520 ( .A1(n15650), .A2(n9802), .ZN(n9801) );
  NAND2_X1 U12521 ( .A1(n14468), .A2(n9805), .ZN(n9809) );
  NAND2_X1 U12522 ( .A1(n9810), .A2(n9808), .ZN(n9807) );
  AND2_X1 U12523 ( .A1(n15560), .A2(n15559), .ZN(n9808) );
  OAI21_X2 U12524 ( .B1(n14486), .B2(n10036), .A(n9811), .ZN(n14468) );
  NAND2_X2 U12525 ( .A1(n15599), .A2(n15598), .ZN(n14486) );
  NAND2_X2 U12526 ( .A1(n10044), .A2(n11189), .ZN(n15599) );
  NAND3_X2 U12527 ( .A1(n9814), .A2(n9813), .A3(n9682), .ZN(n10832) );
  NAND2_X1 U12528 ( .A1(n10274), .A2(n10832), .ZN(n10254) );
  NAND3_X1 U12529 ( .A1(n9818), .A2(n9714), .A3(n11178), .ZN(n14515) );
  AND2_X4 U12530 ( .A1(n10038), .A2(n10143), .ZN(n10208) );
  AND2_X2 U12531 ( .A1(n10038), .A2(n13167), .ZN(n10187) );
  NAND2_X1 U12532 ( .A1(n13131), .A2(n10882), .ZN(n13142) );
  NOR3_X4 U12533 ( .A1(n14225), .A2(n14210), .A3(n9830), .ZN(n14209) );
  INV_X1 U12534 ( .A(n14131), .ZN(n9832) );
  NAND2_X1 U12535 ( .A1(n9833), .A2(n10883), .ZN(n10887) );
  NAND2_X1 U12536 ( .A1(n9833), .A2(n15555), .ZN(n10926) );
  NAND2_X1 U12537 ( .A1(n9833), .A2(n10931), .ZN(n10934) );
  NAND2_X1 U12538 ( .A1(n9833), .A2(n14343), .ZN(n10950) );
  NAND2_X1 U12539 ( .A1(n9833), .A2(n10964), .ZN(n10961) );
  NAND2_X1 U12540 ( .A1(n9833), .A2(n13375), .ZN(n10894) );
  NAND2_X1 U12541 ( .A1(n9833), .A2(n19944), .ZN(n10900) );
  NAND2_X1 U12542 ( .A1(n9833), .A2(n10902), .ZN(n10905) );
  NAND2_X1 U12543 ( .A1(n9833), .A2(n13791), .ZN(n10909) );
  NAND2_X1 U12544 ( .A1(n9833), .A2(n15534), .ZN(n10915) );
  NAND2_X1 U12545 ( .A1(n9833), .A2(n14106), .ZN(n10922) );
  NAND2_X1 U12546 ( .A1(n9833), .A2(n10941), .ZN(n10944) );
  NAND2_X1 U12547 ( .A1(n9833), .A2(n14332), .ZN(n10956) );
  NAND2_X1 U12548 ( .A1(n9833), .A2(n14316), .ZN(n12895) );
  NOR3_X2 U12549 ( .A1(n14353), .A2(n10946), .A3(n9834), .ZN(n14338) );
  INV_X1 U12550 ( .A(n11467), .ZN(n11464) );
  INV_X1 U12551 ( .A(n11462), .ZN(n9838) );
  NAND2_X2 U12552 ( .A1(n12470), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n11477) );
  NAND3_X2 U12553 ( .A1(n11459), .A2(n11629), .A3(n11419), .ZN(n12470) );
  NAND2_X1 U12554 ( .A1(n10100), .A2(n9729), .ZN(n14726) );
  INV_X1 U12555 ( .A(n16011), .ZN(n14731) );
  INV_X1 U12556 ( .A(n14728), .ZN(n9850) );
  AOI21_X1 U12557 ( .B1(n15318), .B2(n9724), .A(n9851), .ZN(n14740) );
  NOR2_X4 U12558 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n13612) );
  AND2_X4 U12559 ( .A1(n13612), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11279) );
  NAND2_X1 U12560 ( .A1(n13832), .A2(n13833), .ZN(n12207) );
  NAND2_X1 U12561 ( .A1(n9629), .A2(n12426), .ZN(n9856) );
  NAND2_X1 U12562 ( .A1(n9857), .A2(n12168), .ZN(n13832) );
  NAND2_X1 U12563 ( .A1(n13674), .A2(n13673), .ZN(n9857) );
  INV_X1 U12564 ( .A(n12939), .ZN(n9858) );
  NAND3_X1 U12565 ( .A1(n9859), .A2(n12941), .A3(n9858), .ZN(n9861) );
  NAND2_X1 U12566 ( .A1(n9861), .A2(n9860), .ZN(n12958) );
  NAND2_X1 U12567 ( .A1(n10102), .A2(n12935), .ZN(n14708) );
  INV_X1 U12568 ( .A(n12941), .ZN(n9862) );
  NAND3_X1 U12569 ( .A1(n9697), .A2(n11393), .A3(n11395), .ZN(n9870) );
  NAND2_X1 U12570 ( .A1(n10088), .A2(n10084), .ZN(n9871) );
  NAND2_X1 U12571 ( .A1(n14975), .A2(n10092), .ZN(n10088) );
  NAND2_X1 U12572 ( .A1(n14566), .A2(n9873), .ZN(n9872) );
  OAI211_X1 U12573 ( .C1(n14566), .C2(n9874), .A(n9872), .B(n12012), .ZN(
        P2_U2825) );
  NOR2_X1 U12574 ( .A1(n14566), .A2(n14565), .ZN(n15876) );
  OR2_X1 U12575 ( .A1(n18735), .A2(n9885), .ZN(n9882) );
  NAND2_X1 U12576 ( .A1(n9882), .A2(n9884), .ZN(n12973) );
  INV_X1 U12577 ( .A(n9890), .ZN(n14071) );
  OR2_X1 U12578 ( .A1(n11250), .A2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n9893) );
  NAND3_X1 U12579 ( .A1(n9893), .A2(n9892), .A3(n9891), .ZN(n14186) );
  NAND3_X1 U12580 ( .A1(n11250), .A2(n9894), .A3(
        P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n9892) );
  INV_X1 U12581 ( .A(n11233), .ZN(n9896) );
  NAND2_X1 U12582 ( .A1(n9898), .A2(n9896), .ZN(n11228) );
  NAND2_X1 U12583 ( .A1(n11223), .A2(n9905), .ZN(n11242) );
  NAND2_X1 U12584 ( .A1(n16101), .A2(n9910), .ZN(n15285) );
  NAND2_X1 U12585 ( .A1(n13825), .A2(n9662), .ZN(n15004) );
  OR2_X2 U12586 ( .A1(n14583), .A2(n14661), .ZN(n14663) );
  NOR2_X2 U12587 ( .A1(n14677), .A2(n14676), .ZN(n14678) );
  INV_X1 U12588 ( .A(n11684), .ZN(n9919) );
  NAND2_X1 U12589 ( .A1(n11096), .A2(n9926), .ZN(n9929) );
  INV_X1 U12590 ( .A(n9929), .ZN(n14197) );
  NAND2_X1 U12591 ( .A1(n11096), .A2(n11099), .ZN(n11098) );
  INV_X1 U12592 ( .A(n11062), .ZN(n9928) );
  NAND2_X1 U12593 ( .A1(n9605), .A2(n9745), .ZN(n14114) );
  AND2_X1 U12594 ( .A1(n14326), .A2(n9937), .ZN(n10991) );
  NAND2_X1 U12595 ( .A1(n14326), .A2(n9733), .ZN(n14220) );
  NAND2_X2 U12596 ( .A1(n10300), .A2(n10364), .ZN(n10302) );
  NAND2_X1 U12597 ( .A1(n10252), .A2(n13397), .ZN(n10264) );
  NAND3_X1 U12598 ( .A1(n9947), .A2(n9946), .A3(n9944), .ZN(n15874) );
  NAND3_X1 U12599 ( .A1(n9947), .A2(n9946), .A3(n9948), .ZN(n15932) );
  NAND3_X1 U12600 ( .A1(n9955), .A2(n9954), .A3(n9953), .ZN(n9952) );
  OAI21_X1 U12601 ( .B1(n16214), .B2(n17617), .A(n9968), .ZN(P3_U2799) );
  NOR2_X1 U12602 ( .A1(n9969), .A2(n13862), .ZN(n13962) );
  NOR2_X1 U12603 ( .A1(n13861), .A2(n9969), .ZN(n15172) );
  NAND2_X1 U12604 ( .A1(n17649), .A2(n9972), .ZN(n9970) );
  INV_X1 U12605 ( .A(n9974), .ZN(n15201) );
  NOR2_X1 U12606 ( .A1(n16165), .A2(n16163), .ZN(n15394) );
  INV_X1 U12607 ( .A(n16215), .ZN(n17363) );
  NOR2_X2 U12608 ( .A1(n15212), .A2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n17364) );
  NAND3_X1 U12609 ( .A1(n9983), .A2(n9982), .A3(n9731), .ZN(n9984) );
  NAND3_X1 U12610 ( .A1(n9983), .A2(n9982), .A3(n9981), .ZN(n17491) );
  INV_X1 U12611 ( .A(n9984), .ZN(n17492) );
  INV_X1 U12612 ( .A(n9987), .ZN(n17676) );
  INV_X1 U12613 ( .A(n15230), .ZN(n9989) );
  OR2_X1 U12614 ( .A1(n14689), .A2(n9995), .ZN(n9993) );
  NAND2_X1 U12615 ( .A1(n9993), .A2(n9992), .ZN(n14627) );
  INV_X1 U12616 ( .A(n9997), .ZN(n14687) );
  NOR2_X2 U12617 ( .A1(n14627), .A2(n12730), .ZN(n12750) );
  INV_X1 U12618 ( .A(n12710), .ZN(n9996) );
  NAND2_X1 U12619 ( .A1(n10002), .A2(n10000), .ZN(n13084) );
  INV_X1 U12620 ( .A(n13083), .ZN(n10001) );
  INV_X1 U12621 ( .A(n10007), .ZN(n10004) );
  CLKBUF_X1 U12622 ( .A(n16679), .Z(n10011) );
  NOR2_X1 U12623 ( .A1(n16402), .A2(n16679), .ZN(n16393) );
  XNOR2_X1 U12624 ( .A(n10026), .B(n15657), .ZN(n15852) );
  NAND2_X2 U12625 ( .A1(n10028), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n10282) );
  NAND4_X1 U12626 ( .A1(n10252), .A2(n10029), .A3(n10260), .A4(n13397), .ZN(
        n10028) );
  OAI21_X2 U12627 ( .B1(n10282), .B2(n10133), .A(n10263), .ZN(n10265) );
  NAND2_X1 U12628 ( .A1(n11191), .A2(n10107), .ZN(n14488) );
  NAND3_X1 U12629 ( .A1(n15639), .A2(n11176), .A3(n11183), .ZN(n10044) );
  AOI21_X2 U12630 ( .B1(n14446), .B2(n15640), .A(n12921), .ZN(n12923) );
  NOR2_X2 U12631 ( .A1(n14460), .A2(n15673), .ZN(n12921) );
  XNOR2_X1 U12632 ( .A(n12398), .B(n13523), .ZN(n16131) );
  NAND2_X2 U12633 ( .A1(n10048), .A2(n10047), .ZN(n15019) );
  NAND2_X1 U12634 ( .A1(n13818), .A2(n10049), .ZN(n10048) );
  OAI21_X1 U12635 ( .B1(n13818), .B2(n10051), .A(n10049), .ZN(n14796) );
  INV_X2 U12636 ( .A(n12430), .ZN(n10051) );
  NAND2_X1 U12637 ( .A1(n12217), .A2(n9747), .ZN(n12232) );
  NAND2_X1 U12638 ( .A1(n12261), .A2(n12260), .ZN(n12239) );
  NAND2_X1 U12639 ( .A1(n12224), .A2(n9730), .ZN(n12247) );
  NAND2_X1 U12640 ( .A1(n10075), .A2(n12688), .ZN(n10074) );
  NAND2_X1 U12641 ( .A1(n11334), .A2(n10104), .ZN(n10079) );
  NAND2_X1 U12642 ( .A1(n11346), .A2(n10078), .ZN(n11400) );
  NAND3_X1 U12643 ( .A1(n11334), .A2(n10104), .A3(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10078) );
  NAND4_X1 U12644 ( .A1(n11407), .A2(n11408), .A3(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A4(n10079), .ZN(n11416) );
  NAND2_X1 U12645 ( .A1(n12498), .A2(n12499), .ZN(n10083) );
  NAND2_X1 U12646 ( .A1(n12325), .A2(n10080), .ZN(n12332) );
  INV_X1 U12647 ( .A(n12499), .ZN(n10082) );
  NAND2_X1 U12648 ( .A1(n10083), .A2(n14696), .ZN(n14699) );
  INV_X1 U12649 ( .A(n14746), .ZN(n10085) );
  NAND2_X1 U12650 ( .A1(n10088), .A2(n10089), .ZN(n14960) );
  NAND2_X1 U12651 ( .A1(n12207), .A2(n12206), .ZN(n13819) );
  OAI21_X1 U12652 ( .B1(n14564), .B2(n20031), .A(n12929), .ZN(n12930) );
  INV_X1 U12653 ( .A(n11974), .ZN(n12437) );
  NOR2_X2 U12654 ( .A1(n17375), .A2(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n17374) );
  OAI211_X2 U12655 ( .C1(n15210), .C2(n17738), .A(n17386), .B(n10127), .ZN(
        n17375) );
  NAND2_X1 U12656 ( .A1(n14573), .A2(n14572), .ZN(n14571) );
  NAND2_X1 U12657 ( .A1(n13172), .A2(n11116), .ZN(n11066) );
  NAND2_X1 U12658 ( .A1(n10249), .A2(n10115), .ZN(n13184) );
  AOI22_X1 U12659 ( .A1(n10171), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n10485), .B2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n10190) );
  AOI22_X1 U12660 ( .A1(n10171), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n10208), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n10161) );
  NAND2_X1 U12661 ( .A1(n10869), .A2(n13489), .ZN(n10250) );
  NAND2_X1 U12662 ( .A1(n20107), .A2(n10832), .ZN(n10868) );
  INV_X1 U12663 ( .A(n10300), .ZN(n20180) );
  OAI22_X1 U12664 ( .A1(n12092), .A2(n12117), .B1(n9673), .B2(n19625), .ZN(
        n12093) );
  AND2_X1 U12665 ( .A1(n20000), .A2(n20096), .ZN(n20026) );
  NAND2_X1 U12666 ( .A1(n12201), .A2(n12200), .ZN(n12427) );
  INV_X1 U12667 ( .A(n12519), .ZN(n13011) );
  OAI22_X1 U12668 ( .A1(n11287), .A2(n11289), .B1(n11355), .B2(n11288), .ZN(
        n11290) );
  NAND2_X1 U12669 ( .A1(n12060), .A2(n12059), .ZN(n12125) );
  NOR2_X1 U12670 ( .A1(n12036), .A2(n12035), .ZN(n12067) );
  NAND2_X1 U12671 ( .A1(n10872), .A2(n10871), .ZN(n19945) );
  INV_X1 U12672 ( .A(n19945), .ZN(n10965) );
  AND2_X1 U12673 ( .A1(n19945), .A2(n13489), .ZN(n19941) );
  AND2_X1 U12674 ( .A1(n12770), .A2(n12790), .ZN(n10101) );
  INV_X1 U12675 ( .A(n18958), .ZN(n15938) );
  AOI21_X1 U12676 ( .B1(n13070), .B2(n13069), .A(n16152), .ZN(n15948) );
  NOR2_X1 U12677 ( .A1(n13859), .A2(n18504), .ZN(n15171) );
  INV_X4 U12678 ( .A(n16994), .ZN(n17014) );
  INV_X1 U12679 ( .A(n14436), .ZN(n14421) );
  AND2_X1 U12680 ( .A1(n12933), .A2(n12938), .ZN(n10102) );
  AND2_X1 U12681 ( .A1(n14696), .A2(n12499), .ZN(n10103) );
  AND4_X1 U12682 ( .A1(n11326), .A2(n11325), .A3(n11324), .A4(n11323), .ZN(
        n10104) );
  NAND2_X1 U12683 ( .A1(n12227), .A2(n14988), .ZN(n10105) );
  NAND2_X1 U12684 ( .A1(n15213), .A2(n17715), .ZN(n10106) );
  AND3_X1 U12685 ( .A1(n15413), .A2(n15419), .A3(n15749), .ZN(n10107) );
  AND2_X1 U12686 ( .A1(n15124), .A2(n15123), .ZN(n10108) );
  AND2_X1 U12687 ( .A1(n9629), .A2(n13686), .ZN(n10109) );
  AND2_X1 U12688 ( .A1(n14436), .A2(n20117), .ZN(n10110) );
  OR2_X1 U12689 ( .A1(n12897), .A2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n10111) );
  OR2_X1 U12690 ( .A1(n12897), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n10112) );
  AND4_X1 U12691 ( .A1(n15143), .A2(n15142), .A3(n15141), .A4(n15140), .ZN(
        n10113) );
  OR2_X1 U12692 ( .A1(n12897), .A2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n10114) );
  AND2_X1 U12693 ( .A1(n13174), .A2(n10248), .ZN(n10115) );
  INV_X1 U12694 ( .A(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n11213) );
  INV_X1 U12695 ( .A(n18892), .ZN(n18935) );
  INV_X1 U12696 ( .A(n12729), .ZN(n12708) );
  INV_X1 U12697 ( .A(n13331), .ZN(n13571) );
  AND4_X1 U12698 ( .A1(n15131), .A2(n15130), .A3(n15129), .A4(n15128), .ZN(
        n10116) );
  OR3_X1 U12699 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A3(n17435), .ZN(n10117) );
  OR2_X1 U12700 ( .A1(n12897), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n10118) );
  AND2_X1 U12701 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n10119) );
  OR2_X1 U12702 ( .A1(n12651), .A2(n12650), .ZN(n10120) );
  NAND2_X1 U12703 ( .A1(n9654), .A2(n11390), .ZN(n11492) );
  NOR2_X1 U12704 ( .A1(n20433), .A2(n20404), .ZN(n10121) );
  INV_X1 U12705 ( .A(n12751), .ZN(n12747) );
  OR2_X1 U12706 ( .A1(n12897), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n10122) );
  AND2_X1 U12707 ( .A1(n18995), .A2(n11630), .ZN(n19027) );
  INV_X1 U12708 ( .A(n15139), .ZN(n13880) );
  INV_X1 U12709 ( .A(n15134), .ZN(n13882) );
  OR2_X1 U12710 ( .A1(n12897), .A2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n10123) );
  OR2_X1 U12711 ( .A1(n12897), .A2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n10124) );
  AND2_X1 U12712 ( .A1(n15197), .A2(n15258), .ZN(n10125) );
  INV_X1 U12713 ( .A(n12795), .ZN(n12793) );
  AND2_X2 U12714 ( .A1(n11630), .A2(n19594), .ZN(n11963) );
  XOR2_X1 U12715 ( .A(n15394), .B(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .Z(
        n10126) );
  OR2_X1 U12716 ( .A1(n17615), .A2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n10127) );
  INV_X1 U12717 ( .A(n17615), .ZN(n15213) );
  AND2_X1 U12718 ( .A1(n12537), .A2(n12536), .ZN(n10128) );
  OR3_X1 U12719 ( .A1(n14805), .A2(n14986), .A3(n12492), .ZN(n10129) );
  INV_X1 U12720 ( .A(n19110), .ZN(n12942) );
  NAND2_X1 U12721 ( .A1(n10424), .A2(n10423), .ZN(n10130) );
  INV_X1 U12722 ( .A(n13140), .ZN(n10378) );
  NAND2_X1 U12723 ( .A1(n9650), .A2(n13011), .ZN(n12057) );
  AND2_X1 U12724 ( .A1(n11063), .A2(n12902), .ZN(n10251) );
  OR2_X1 U12725 ( .A1(n11355), .A2(n19161), .ZN(n11273) );
  AND2_X1 U12726 ( .A1(n11471), .A2(n11417), .ZN(n11418) );
  NAND2_X1 U12727 ( .A1(n11420), .A2(n11450), .ZN(n11433) );
  INV_X1 U12728 ( .A(n10862), .ZN(n10858) );
  AND2_X1 U12729 ( .A1(n10422), .A2(n10421), .ZN(n10423) );
  INV_X1 U12730 ( .A(n10868), .ZN(n10198) );
  NOR2_X1 U12731 ( .A1(n10861), .A2(n11071), .ZN(n10863) );
  NAND2_X1 U12732 ( .A1(n12861), .A2(n11418), .ZN(n11419) );
  OAI22_X1 U12733 ( .A1(n12049), .A2(n12122), .B1(n12117), .B2(n12048), .ZN(
        n12050) );
  AND2_X1 U12734 ( .A1(n10829), .A2(n10828), .ZN(n10831) );
  AND2_X1 U12735 ( .A1(n20703), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10848) );
  INV_X1 U12736 ( .A(n13749), .ZN(n10472) );
  INV_X1 U12737 ( .A(n14223), .ZN(n10990) );
  OR2_X1 U12738 ( .A1(n14272), .A2(n14435), .ZN(n10646) );
  AND2_X1 U12739 ( .A1(n14501), .A2(n11182), .ZN(n11183) );
  OR2_X1 U12740 ( .A1(n11213), .A2(n13836), .ZN(n11214) );
  AND2_X1 U12741 ( .A1(n12773), .A2(n10101), .ZN(n12774) );
  INV_X1 U12742 ( .A(n12043), .ZN(n12044) );
  NAND2_X1 U12743 ( .A1(n11626), .A2(n11625), .ZN(n11624) );
  AOI21_X1 U12744 ( .B1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n20690), .A(
        n10831), .ZN(n10859) );
  INV_X1 U12745 ( .A(n10475), .ZN(n10476) );
  NAND2_X1 U12746 ( .A1(n13141), .A2(n10379), .ZN(n13337) );
  INV_X1 U12747 ( .A(n11196), .ZN(n11195) );
  NAND2_X1 U12748 ( .A1(n13128), .A2(n14200), .ZN(n12890) );
  OR2_X1 U12749 ( .A1(n10397), .A2(n10396), .ZN(n11130) );
  OR2_X1 U12750 ( .A1(n10276), .A2(n13401), .ZN(n10361) );
  NAND2_X1 U12751 ( .A1(n10490), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(
        n10211) );
  NOR2_X1 U12752 ( .A1(n11679), .A2(n11678), .ZN(n12400) );
  INV_X1 U12753 ( .A(n11474), .ZN(n12452) );
  INV_X1 U12754 ( .A(n18940), .ZN(n12567) );
  OR2_X1 U12755 ( .A1(n13736), .A2(n13735), .ZN(n11954) );
  AOI21_X1 U12756 ( .B1(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n19757), .A(
        n11623), .ZN(n11627) );
  NOR2_X1 U12757 ( .A1(n13861), .A2(n13860), .ZN(n15134) );
  OAI21_X1 U12758 ( .B1(n16224), .B2(n18486), .A(n16223), .ZN(n16225) );
  INV_X1 U12759 ( .A(n15171), .ZN(n15148) );
  INV_X1 U12760 ( .A(n11064), .ZN(n15346) );
  NAND2_X1 U12761 ( .A1(n10386), .A2(n10385), .ZN(n20214) );
  NAND2_X1 U12762 ( .A1(n14177), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11057) );
  INV_X1 U12763 ( .A(n10500), .ZN(n10503) );
  AND2_X1 U12764 ( .A1(n14529), .A2(n14531), .ZN(n15615) );
  INV_X1 U12765 ( .A(n20066), .ZN(n15798) );
  AND2_X1 U12766 ( .A1(n10340), .A2(n11170), .ZN(n11101) );
  XNOR2_X1 U12767 ( .A(n11115), .B(n10372), .ZN(n13433) );
  AND4_X1 U12768 ( .A1(n10206), .A2(n10205), .A3(n10204), .A4(n10203), .ZN(
        n10220) );
  AND2_X1 U12769 ( .A1(n12549), .A2(n13364), .ZN(n12550) );
  AND2_X1 U12770 ( .A1(n15935), .A2(n12708), .ZN(n12710) );
  INV_X1 U12771 ( .A(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n11220) );
  OR2_X1 U12772 ( .A1(n11609), .A2(n14055), .ZN(n11530) );
  INV_X1 U12773 ( .A(n11487), .ZN(n11488) );
  NOR2_X1 U12774 ( .A1(n14859), .A2(n12488), .ZN(n14829) );
  AND2_X1 U12775 ( .A1(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n14056), .ZN(
        n16115) );
  NAND2_X1 U12776 ( .A1(n12161), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n13524) );
  NAND2_X1 U12777 ( .A1(n12354), .A2(n12353), .ZN(n12357) );
  AND2_X1 U12778 ( .A1(n13560), .A2(n19752), .ZN(n13567) );
  AND2_X1 U12779 ( .A1(n16380), .A2(n16727), .ZN(n16381) );
  NOR2_X1 U12780 ( .A1(n13858), .A2(n13860), .ZN(n15139) );
  OAI21_X1 U12781 ( .B1(n16693), .B2(n17427), .A(n18078), .ZN(n17544) );
  INV_X1 U12782 ( .A(n17411), .ZN(n17434) );
  NAND2_X1 U12783 ( .A1(n18512), .A2(n18509), .ZN(n17919) );
  OAI21_X2 U12784 ( .B1(n18494), .B2(n15239), .A(n18493), .ZN(n18510) );
  NAND2_X1 U12785 ( .A1(n10503), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n10522) );
  INV_X1 U12786 ( .A(n19922), .ZN(n14228) );
  NAND2_X1 U12787 ( .A1(n12910), .A2(n12909), .ZN(n19867) );
  INV_X1 U12788 ( .A(n14271), .ZN(n14360) );
  OR2_X2 U12789 ( .A1(n20086), .A2(n10256), .ZN(n20722) );
  INV_X1 U12790 ( .A(n10991), .ZN(n14222) );
  OR2_X1 U12791 ( .A1(n10600), .A2(n10585), .ZN(n10624) );
  NOR2_X1 U12792 ( .A1(n10522), .A2(n10521), .ZN(n10537) );
  INV_X1 U12793 ( .A(n11154), .ZN(n11141) );
  NOR2_X1 U12794 ( .A1(n20149), .A2(n20693), .ZN(n20177) );
  OR2_X1 U12795 ( .A1(n13434), .A2(n10401), .ZN(n20300) );
  OR2_X1 U12796 ( .A1(n20683), .A2(n20322), .ZN(n20681) );
  INV_X1 U12797 ( .A(n20243), .ZN(n20464) );
  OR2_X1 U12798 ( .A1(n12365), .A2(n11628), .ZN(n13631) );
  AND2_X1 U12799 ( .A1(n12546), .A2(n13234), .ZN(n13227) );
  AND2_X1 U12800 ( .A1(n11530), .A2(n11529), .ZN(n13245) );
  NOR2_X1 U12801 ( .A1(n9661), .A2(n12324), .ZN(n12325) );
  INV_X1 U12802 ( .A(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n14707) );
  AND2_X1 U12803 ( .A1(n12279), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n14748) );
  AND3_X1 U12804 ( .A1(n11824), .A2(n11823), .A3(n11822), .ZN(n16113) );
  NAND2_X1 U12805 ( .A1(n15037), .A2(n18715), .ZN(n13563) );
  AND3_X1 U12806 ( .A1(n13060), .A2(n13070), .A3(n13059), .ZN(n13622) );
  INV_X1 U12807 ( .A(n19185), .ZN(n19342) );
  OR2_X1 U12808 ( .A1(n19138), .A2(n19767), .ZN(n19395) );
  NAND3_X1 U12809 ( .A1(P2_STATEBS16_REG_SCAN_IN), .A2(n19752), .A3(n19593), 
        .ZN(n13572) );
  INV_X1 U12810 ( .A(n16735), .ZN(n16744) );
  NOR3_X1 U12811 ( .A1(n16888), .A2(n16904), .A3(n16892), .ZN(n16874) );
  INV_X1 U12812 ( .A(n18071), .ZN(n17082) );
  INV_X1 U12813 ( .A(n17213), .ZN(n17180) );
  OAI21_X1 U12814 ( .B1(n15065), .B2(n15064), .A(n15063), .ZN(n18482) );
  AND2_X1 U12815 ( .A1(n17352), .A2(n17351), .ZN(n17353) );
  AND2_X1 U12816 ( .A1(n16159), .A2(n16158), .ZN(n16160) );
  AOI21_X1 U12817 ( .B1(n17343), .B2(n16240), .A(n16239), .ZN(n16241) );
  AND2_X1 U12818 ( .A1(n17411), .A2(n17445), .ZN(n17484) );
  NOR2_X1 U12819 ( .A1(n17653), .A2(n17652), .ZN(n17651) );
  OAI21_X1 U12820 ( .B1(n14549), .B2(n19931), .A(n12914), .ZN(n12915) );
  NAND2_X1 U12821 ( .A1(n10699), .A2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n10717) );
  INV_X1 U12822 ( .A(n19879), .ZN(n19891) );
  INV_X1 U12823 ( .A(n19931), .ZN(n19905) );
  INV_X2 U12824 ( .A(n20000), .ZN(n20025) );
  NAND2_X1 U12825 ( .A1(n10804), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n11011) );
  NAND2_X1 U12826 ( .A1(n10467), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n10477) );
  INV_X1 U12827 ( .A(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n12924) );
  AND2_X1 U12828 ( .A1(n13413), .A2(n13405), .ZN(n15773) );
  INV_X1 U12829 ( .A(n20060), .ZN(n15834) );
  INV_X1 U12830 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n13329) );
  AND2_X1 U12831 ( .A1(n20683), .A2(n13434), .ZN(n20178) );
  AND2_X1 U12832 ( .A1(n20178), .A2(n20150), .ZN(n20207) );
  NOR2_X1 U12833 ( .A1(n20300), .A2(n20493), .ZN(n20311) );
  NOR2_X1 U12834 ( .A1(n20701), .A2(n13433), .ZN(n20434) );
  NOR2_X1 U12835 ( .A1(n20681), .A2(n20493), .ZN(n20424) );
  OAI22_X1 U12836 ( .A1(n20492), .A2(n20444), .B1(n20443), .B2(n20442), .ZN(
        n20459) );
  OAI211_X1 U12837 ( .C1(n20528), .C2(n20500), .A(n20499), .B(n20498), .ZN(
        n20530) );
  OR2_X1 U12838 ( .A1(n13631), .A2(n16152), .ZN(n12988) );
  INV_X1 U12839 ( .A(n15875), .ZN(n11252) );
  AND2_X1 U12840 ( .A1(n12226), .A2(n12225), .ZN(n18849) );
  INV_X1 U12841 ( .A(n18932), .ZN(n18910) );
  AOI21_X1 U12842 ( .B1(n14612), .B2(n14609), .A(n14611), .ZN(n15899) );
  INV_X1 U12843 ( .A(n18952), .ZN(n15942) );
  NOR2_X1 U12844 ( .A1(n15038), .A2(n13046), .ZN(n19137) );
  AND2_X1 U12845 ( .A1(n11953), .A2(n11952), .ZN(n13736) );
  OR2_X1 U12846 ( .A1(n18963), .A2(n13038), .ZN(n18997) );
  INV_X1 U12847 ( .A(n13348), .ZN(n13120) );
  AND2_X1 U12848 ( .A1(n12503), .A2(n12068), .ZN(n16068) );
  INV_X1 U12849 ( .A(n15445), .ZN(n18751) );
  INV_X1 U12850 ( .A(n12482), .ZN(n19081) );
  OR2_X1 U12851 ( .A1(n19116), .A2(n14882), .ZN(n19132) );
  INV_X1 U12852 ( .A(n19000), .ZN(n19754) );
  AND2_X1 U12853 ( .A1(n13635), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n15037) );
  OAI21_X1 U12854 ( .B1(n19146), .B2(n19145), .A(n19144), .ZN(n19181) );
  NOR2_X1 U12855 ( .A1(n19395), .A2(n19307), .ZN(n19211) );
  NOR2_X1 U12856 ( .A1(n19754), .A2(n19779), .ZN(n19185) );
  INV_X1 U12857 ( .A(n19261), .ZN(n19263) );
  AND2_X1 U12858 ( .A1(n13808), .A2(n13807), .ZN(n19282) );
  INV_X1 U12859 ( .A(n19293), .ZN(n19299) );
  NOR2_X1 U12860 ( .A1(n19342), .A2(n19533), .ZN(n19324) );
  OAI21_X1 U12861 ( .B1(n19373), .B2(n19372), .A(n19371), .ZN(n19390) );
  NOR2_X1 U12862 ( .A1(n19555), .A2(n19459), .ZN(n19479) );
  OAI21_X1 U12863 ( .B1(n19565), .B2(n19564), .A(n19563), .ZN(n19583) );
  INV_X1 U12864 ( .A(n19518), .ZN(n19641) );
  NAND2_X1 U12865 ( .A1(n18047), .A2(n17291), .ZN(n15234) );
  OAI22_X1 U12866 ( .A1(n16155), .A2(n18486), .B1(n18489), .B2(n16226), .ZN(
        n18491) );
  INV_X1 U12867 ( .A(n16753), .ZN(n16723) );
  INV_X1 U12868 ( .A(n16739), .ZN(n16691) );
  NOR2_X1 U12869 ( .A1(n13956), .A2(n16837), .ZN(n16816) );
  NOR4_X1 U12870 ( .A1(n16593), .A2(n16970), .A3(n17032), .A4(n16946), .ZN(
        n16944) );
  NOR2_X1 U12871 ( .A1(n13955), .A2(n17048), .ZN(n17044) );
  INV_X1 U12872 ( .A(n17112), .ZN(n17107) );
  NOR2_X1 U12873 ( .A1(n20833), .A2(n17142), .ZN(n17137) );
  NAND3_X1 U12874 ( .A1(n13891), .A2(n13890), .A3(n13889), .ZN(n17227) );
  INV_X1 U12875 ( .A(n17338), .ZN(n17329) );
  OR2_X1 U12876 ( .A1(n17354), .A2(n17353), .ZN(n17355) );
  NOR2_X1 U12877 ( .A1(n17608), .A2(n17820), .ZN(n17499) );
  NOR2_X1 U12878 ( .A1(n17193), .A2(n9647), .ZN(n17401) );
  INV_X1 U12879 ( .A(n18083), .ZN(n18388) );
  NAND2_X1 U12880 ( .A1(n16231), .A2(n16230), .ZN(n16232) );
  NAND3_X1 U12881 ( .A1(n15101), .A2(n15100), .A3(n15099), .ZN(n17193) );
  INV_X1 U12882 ( .A(n18012), .ZN(n18021) );
  AOI21_X1 U12883 ( .B1(n15229), .B2(n15228), .A(n18534), .ZN(n18025) );
  INV_X1 U12884 ( .A(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n18515) );
  NAND2_X1 U12885 ( .A1(n15404), .A2(n12996), .ZN(n20726) );
  INV_X1 U12886 ( .A(P1_STATEBS16_REG_SCAN_IN), .ZN(n20891) );
  INV_X1 U12887 ( .A(n12915), .ZN(n12916) );
  NAND2_X1 U12888 ( .A1(n13128), .A2(n12901), .ZN(n19931) );
  INV_X1 U12889 ( .A(n19872), .ZN(n19861) );
  AND2_X1 U12890 ( .A1(n10967), .A2(n10966), .ZN(n10968) );
  INV_X1 U12891 ( .A(n14465), .ZN(n14381) );
  NAND2_X1 U12892 ( .A1(n14436), .A2(n13492), .ZN(n14144) );
  AND2_X1 U12893 ( .A1(n15411), .A2(n15410), .ZN(n19996) );
  NOR2_X1 U12894 ( .A1(n15404), .A2(n13266), .ZN(n20000) );
  NOR2_X1 U12895 ( .A1(n11211), .A2(n11210), .ZN(n11212) );
  INV_X1 U12896 ( .A(n15635), .ZN(n20032) );
  INV_X1 U12897 ( .A(n20078), .ZN(n20070) );
  INV_X1 U12898 ( .A(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n15861) );
  NAND2_X1 U12899 ( .A1(n20178), .A2(n20434), .ZN(n20934) );
  INV_X1 U12900 ( .A(n20930), .ZN(n20176) );
  INV_X1 U12901 ( .A(n20207), .ZN(n20206) );
  NAND2_X1 U12902 ( .A1(n20296), .A2(n20434), .ZN(n20263) );
  INV_X1 U12903 ( .A(n20311), .ZN(n20321) );
  NAND2_X1 U12904 ( .A1(n20323), .A2(n20434), .ZN(n20374) );
  INV_X1 U12905 ( .A(n20424), .ZN(n20432) );
  INV_X1 U12906 ( .A(n20436), .ZN(n20463) );
  INV_X1 U12907 ( .A(n20495), .ZN(n20533) );
  INV_X1 U12908 ( .A(n20121), .ZN(n20595) );
  INV_X1 U12909 ( .A(P2_STATE2_REG_0__SCAN_IN), .ZN(n18715) );
  AND2_X1 U12910 ( .A1(n12011), .A2(n12010), .ZN(n12012) );
  OR3_X1 U12911 ( .A1(n11987), .A2(P2_STATEBS16_REG_SCAN_IN), .A3(n19807), 
        .ZN(n18924) );
  INV_X1 U12912 ( .A(n18958), .ZN(n18945) );
  OAI21_X1 U12913 ( .B1(n13076), .B2(n13077), .A(n13078), .ZN(n19000) );
  AND2_X1 U12914 ( .A1(n12878), .A2(n12877), .ZN(n12879) );
  NAND2_X2 U12915 ( .A1(n12863), .A2(n12862), .ZN(n18995) );
  INV_X1 U12916 ( .A(n18997), .ZN(n19035) );
  OR2_X1 U12917 ( .A1(n19071), .A2(n13156), .ZN(n19037) );
  NAND2_X1 U12918 ( .A1(n13155), .A2(n19795), .ZN(n19071) );
  INV_X1 U12919 ( .A(n19077), .ZN(n13347) );
  INV_X1 U12920 ( .A(n19080), .ZN(n16063) );
  OR2_X1 U12921 ( .A1(n12481), .A2(n19786), .ZN(n19125) );
  OR2_X1 U12922 ( .A1(n12481), .A2(n19791), .ZN(n19110) );
  INV_X1 U12923 ( .A(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19757) );
  AOI211_X2 U12924 ( .C1(n19142), .C2(n19145), .A(n19528), .B(n19141), .ZN(
        n19184) );
  INV_X1 U12925 ( .A(n19211), .ZN(n19208) );
  NAND2_X1 U12926 ( .A1(n19186), .A2(n19185), .ZN(n19246) );
  OR2_X1 U12927 ( .A1(n19307), .A2(n19459), .ZN(n19261) );
  INV_X1 U12928 ( .A(n19276), .ZN(n19286) );
  OR2_X1 U12929 ( .A1(n19307), .A2(n19533), .ZN(n19293) );
  INV_X1 U12930 ( .A(n19324), .ZN(n19332) );
  INV_X1 U12931 ( .A(n19360), .ZN(n19353) );
  INV_X1 U12932 ( .A(n19386), .ZN(n19394) );
  INV_X1 U12933 ( .A(n19419), .ZN(n19418) );
  INV_X1 U12934 ( .A(n19445), .ZN(n19453) );
  INV_X1 U12935 ( .A(n19493), .ZN(n19524) );
  AOI21_X1 U12936 ( .B1(n19561), .B2(n19564), .A(n19560), .ZN(n19586) );
  AOI21_X1 U12937 ( .B1(n19596), .B2(n19597), .A(n19595), .ZN(n19656) );
  NAND2_X1 U12938 ( .A1(n18686), .A2(n18491), .ZN(n16349) );
  INV_X1 U12939 ( .A(n16754), .ZN(n16743) );
  NAND2_X1 U12940 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n16810), .ZN(n16805) );
  INV_X1 U12941 ( .A(n16800), .ZN(n16810) );
  NOR2_X1 U12942 ( .A1(n16563), .A2(n16943), .ZN(n16932) );
  AND2_X1 U12943 ( .A1(n17073), .A2(n17123), .ZN(n17070) );
  OR2_X1 U12944 ( .A1(n17265), .A2(n17182), .ZN(n17176) );
  INV_X1 U12945 ( .A(n15258), .ZN(n17198) );
  INV_X1 U12946 ( .A(n17222), .ZN(n17217) );
  INV_X1 U12947 ( .A(n17255), .ZN(n17287) );
  INV_X1 U12948 ( .A(n17336), .ZN(n17331) );
  INV_X1 U12949 ( .A(n17401), .ZN(n17616) );
  AOI22_X1 U12950 ( .A1(n17697), .A2(n17902), .B1(n17401), .B2(n17904), .ZN(
        n17608) );
  NOR2_X1 U12951 ( .A1(n17376), .A2(n17565), .ZN(n17704) );
  NAND2_X1 U12952 ( .A1(n16242), .A2(n17933), .ZN(n16243) );
  INV_X1 U12953 ( .A(n18025), .ZN(n18019) );
  INV_X1 U12954 ( .A(n17999), .ZN(n18033) );
  INV_X1 U12955 ( .A(P3_STATE2_REG_3__SCAN_IN), .ZN(n18639) );
  NAND2_X1 U12956 ( .A1(n10969), .A2(n10968), .ZN(P1_U2846) );
  OAI21_X1 U12957 ( .B1(n14373), .B2(n20084), .A(n11212), .ZN(P1_U2970) );
  OAI21_X1 U12958 ( .B1(n14826), .B2(n19088), .A(n12511), .ZN(P2_U2985) );
  AOI22_X1 U12959 ( .A1(n10290), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n10291), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n10138) );
  AOI22_X1 U12960 ( .A1(n10490), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n10227), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n10137) );
  INV_X1 U12961 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10133) );
  AOI22_X1 U12962 ( .A1(n10492), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n10226), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n10136) );
  AOI22_X1 U12963 ( .A1(n9616), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n10213), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10135) );
  AOI22_X1 U12964 ( .A1(n10458), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n10187), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n10147) );
  AND2_X2 U12965 ( .A1(n10139), .A2(n10141), .ZN(n10171) );
  AOI22_X1 U12966 ( .A1(n10485), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n10171), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n10146) );
  AOI22_X1 U12967 ( .A1(n10998), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n9638), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10145) );
  AOI22_X1 U12968 ( .A1(n9620), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n10208), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n10144) );
  AOI22_X1 U12969 ( .A1(n10290), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n10291), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n10150) );
  AOI22_X1 U12970 ( .A1(n10972), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n9628), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n10149) );
  AOI22_X1 U12971 ( .A1(n9616), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n10213), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n10148) );
  AOI22_X1 U12972 ( .A1(n10485), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n10227), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n10155) );
  AOI22_X1 U12973 ( .A1(n10492), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n10226), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n10154) );
  AOI22_X1 U12974 ( .A1(n10490), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n9621), .B2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n10153) );
  AOI22_X1 U12975 ( .A1(n10171), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n10208), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n10152) );
  NAND2_X2 U12976 ( .A1(n9675), .A2(n9613), .ZN(n13389) );
  AOI22_X1 U12977 ( .A1(n10290), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n9617), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n10159) );
  AOI22_X1 U12978 ( .A1(n10458), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n10226), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n10158) );
  AOI22_X1 U12979 ( .A1(n10490), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n9622), .B2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n10157) );
  AOI22_X1 U12980 ( .A1(n10972), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n9638), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10156) );
  AOI22_X1 U12981 ( .A1(n10485), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n10227), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n10163) );
  AOI22_X1 U12982 ( .A1(n10492), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n10187), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n10162) );
  AOI22_X1 U12983 ( .A1(n10291), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n10213), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10160) );
  NAND2_X2 U12984 ( .A1(n10131), .A2(n10164), .ZN(n11116) );
  INV_X1 U12985 ( .A(n11116), .ZN(n20103) );
  OAI21_X1 U12986 ( .B1(n10248), .B2(n13389), .A(n20103), .ZN(n10176) );
  AOI22_X1 U12987 ( .A1(n10458), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n10187), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n10166) );
  AOI22_X1 U12988 ( .A1(n9616), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n10213), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10165) );
  NAND2_X1 U12989 ( .A1(n10166), .A2(n10165), .ZN(n10170) );
  AOI22_X1 U12990 ( .A1(n10290), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n10291), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n10168) );
  AOI22_X1 U12991 ( .A1(n10998), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n9628), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n10167) );
  NAND2_X1 U12992 ( .A1(n10168), .A2(n10167), .ZN(n10169) );
  AOI22_X1 U12993 ( .A1(n10490), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n9620), .B2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n10175) );
  AOI22_X1 U12994 ( .A1(n10485), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n10227), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n10174) );
  AOI22_X1 U12995 ( .A1(n10492), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n10226), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n10173) );
  AOI22_X1 U12996 ( .A1(n10171), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n10208), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n10172) );
  NAND2_X1 U12997 ( .A1(n10176), .A2(n10254), .ZN(n10197) );
  AOI22_X1 U12998 ( .A1(n10492), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n10226), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n10180) );
  AOI22_X1 U12999 ( .A1(n10485), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n10227), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n10179) );
  AOI22_X1 U13000 ( .A1(n10490), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n9621), .B2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n10178) );
  AOI22_X1 U13001 ( .A1(n10171), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n10208), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n10177) );
  NAND4_X1 U13002 ( .A1(n10180), .A2(n10179), .A3(n10178), .A4(n10177), .ZN(
        n10186) );
  AOI22_X1 U13003 ( .A1(n10290), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n10291), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n10184) );
  AOI22_X1 U13004 ( .A1(n9618), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n10213), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n10183) );
  AOI22_X1 U13005 ( .A1(n10972), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n9628), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n10182) );
  AOI22_X1 U13006 ( .A1(n10458), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n10187), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n10181) );
  NAND4_X1 U13007 ( .A1(n10184), .A2(n10183), .A3(n10182), .A4(n10181), .ZN(
        n10185) );
  AOI22_X1 U13009 ( .A1(n10492), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n10226), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n10195) );
  AOI22_X1 U13010 ( .A1(n10490), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n10227), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n10194) );
  AOI22_X1 U13011 ( .A1(n10290), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n10291), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n10193) );
  AOI22_X1 U13012 ( .A1(n10998), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n9628), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n10192) );
  NAND2_X1 U13013 ( .A1(n13410), .A2(n13489), .ZN(n10255) );
  NAND2_X1 U13014 ( .A1(n10250), .A2(n10255), .ZN(n10196) );
  NAND2_X1 U13015 ( .A1(n9659), .A2(n10198), .ZN(n12880) );
  INV_X1 U13016 ( .A(n12880), .ZN(n10244) );
  INV_X1 U13017 ( .A(n10290), .ZN(n10318) );
  NAND2_X1 U13018 ( .A1(n10290), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n10202) );
  NAND2_X1 U13019 ( .A1(n10734), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n10201) );
  NAND2_X1 U13020 ( .A1(n10187), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n10200) );
  NAND2_X1 U13021 ( .A1(n10291), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n10199) );
  NAND2_X1 U13022 ( .A1(n10226), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n10206) );
  NAND2_X1 U13023 ( .A1(n10492), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n10205) );
  NAND2_X1 U13024 ( .A1(n10485), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n10204) );
  NAND2_X1 U13025 ( .A1(n10227), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n10203) );
  NAND2_X1 U13026 ( .A1(n10171), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n10212) );
  NAND2_X1 U13027 ( .A1(n9621), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n10210) );
  BUF_X4 U13028 ( .A(n10208), .Z(n11042) );
  NAND2_X1 U13029 ( .A1(n11042), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(
        n10209) );
  NAND2_X1 U13030 ( .A1(n9619), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n10217) );
  NAND2_X1 U13031 ( .A1(n10972), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n10216) );
  NAND2_X1 U13032 ( .A1(n9638), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n10215) );
  NAND2_X1 U13033 ( .A1(n10213), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n10214) );
  AND4_X4 U13034 ( .A1(n10221), .A2(n10220), .A3(n10219), .A4(n10218), .ZN(
        n20086) );
  NAND2_X1 U13035 ( .A1(n10290), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n10225) );
  NAND2_X1 U13036 ( .A1(n10734), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n10224) );
  NAND2_X1 U13037 ( .A1(n10187), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n10223) );
  NAND2_X1 U13038 ( .A1(n10291), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n10222) );
  NAND2_X1 U13039 ( .A1(n10226), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n10231) );
  NAND2_X1 U13040 ( .A1(n10492), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n10230) );
  NAND2_X1 U13041 ( .A1(n10485), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n10229) );
  NAND2_X1 U13042 ( .A1(n10227), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n10228) );
  NAND2_X1 U13043 ( .A1(n9619), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n10235) );
  NAND2_X1 U13044 ( .A1(n10972), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n10234) );
  NAND2_X1 U13045 ( .A1(n9628), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n10233) );
  NAND2_X1 U13046 ( .A1(n10213), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n10232) );
  NAND2_X1 U13047 ( .A1(n10171), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n10239) );
  NAND2_X1 U13048 ( .A1(n10490), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n10238) );
  NAND2_X1 U13049 ( .A1(n9622), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n10237) );
  NAND2_X1 U13050 ( .A1(n11042), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n10236) );
  NAND2_X1 U13051 ( .A1(n10244), .A2(n10249), .ZN(n11067) );
  NAND2_X1 U13052 ( .A1(n10248), .A2(n10869), .ZN(n10245) );
  NAND2_X1 U13053 ( .A1(n10245), .A2(n13489), .ZN(n11198) );
  NOR2_X1 U13054 ( .A1(n11066), .A2(n10832), .ZN(n10246) );
  NOR2_X2 U13055 ( .A1(n13185), .A2(n20086), .ZN(n11063) );
  NAND2_X1 U13056 ( .A1(n11063), .A2(n10256), .ZN(n10247) );
  NOR2_X1 U13057 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(P1_STATE_REG_2__SCAN_IN), 
        .ZN(n20602) );
  AOI21_X1 U13058 ( .B1(P1_STATE_REG_2__SCAN_IN), .B2(P1_STATE_REG_1__SCAN_IN), 
        .A(n20602), .ZN(n12902) );
  NAND2_X1 U13059 ( .A1(n9606), .A2(n13490), .ZN(n13181) );
  NAND2_X1 U13060 ( .A1(n13181), .A2(n13165), .ZN(n10261) );
  NAND2_X1 U13061 ( .A1(n11116), .A2(n9640), .ZN(n10268) );
  OR2_X1 U13062 ( .A1(n10868), .A2(n10268), .ZN(n13404) );
  NAND2_X1 U13063 ( .A1(n20086), .A2(n10256), .ZN(n14298) );
  INV_X1 U13064 ( .A(n20086), .ZN(n19946) );
  NAND2_X1 U13065 ( .A1(n19946), .A2(n13389), .ZN(n13177) );
  INV_X1 U13066 ( .A(n13174), .ZN(n10257) );
  OAI21_X1 U13067 ( .B1(n20722), .B2(n20107), .A(n10257), .ZN(n10258) );
  NOR2_X1 U13068 ( .A1(n10267), .A2(n10258), .ZN(n10260) );
  INV_X1 U13069 ( .A(n20536), .ZN(n10381) );
  NAND2_X1 U13070 ( .A1(n20703), .A2(n20697), .ZN(n20433) );
  NAND2_X1 U13071 ( .A1(n10381), .A2(n20433), .ZN(n20378) );
  INV_X1 U13072 ( .A(n11205), .ZN(n10383) );
  INV_X1 U13073 ( .A(P1_STATE2_REG_1__SCAN_IN), .ZN(n13663) );
  NAND2_X1 U13074 ( .A1(n13663), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n15362) );
  NAND2_X1 U13075 ( .A1(n15362), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n10278) );
  OAI21_X1 U13076 ( .B1(n20378), .B2(n10383), .A(n10278), .ZN(n10262) );
  INV_X1 U13077 ( .A(n10262), .ZN(n10263) );
  MUX2_X1 U13078 ( .A(n15362), .B(n11205), .S(n20703), .Z(n10341) );
  INV_X1 U13079 ( .A(n10341), .ZN(n10266) );
  OAI21_X2 U13080 ( .B1(n10282), .B2(n9779), .A(n10266), .ZN(n10362) );
  NAND3_X1 U13081 ( .A1(n13181), .A2(n13165), .A3(n10256), .ZN(n10273) );
  INV_X1 U13082 ( .A(n10267), .ZN(n10272) );
  AND2_X1 U13083 ( .A1(n15343), .A2(n10268), .ZN(n12998) );
  NAND2_X1 U13084 ( .A1(n13490), .A2(n11116), .ZN(n10269) );
  NAND2_X1 U13085 ( .A1(n15857), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n19822) );
  AOI21_X1 U13086 ( .B1(n12998), .B2(n10269), .A(n19822), .ZN(n10271) );
  OR2_X1 U13087 ( .A1(n9606), .A2(n20722), .ZN(n10270) );
  NAND4_X1 U13088 ( .A1(n10273), .A2(n10272), .A3(n10271), .A4(n10270), .ZN(
        n10276) );
  NAND2_X1 U13089 ( .A1(n13174), .A2(n10274), .ZN(n10275) );
  NAND2_X1 U13090 ( .A1(n13186), .A2(n10275), .ZN(n13401) );
  INV_X1 U13091 ( .A(n10277), .ZN(n10280) );
  NAND2_X1 U13092 ( .A1(n10278), .A2(n9778), .ZN(n10279) );
  NAND2_X1 U13093 ( .A1(n10280), .A2(n10279), .ZN(n10281) );
  NAND2_X1 U13094 ( .A1(n15362), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n10284) );
  XNOR2_X1 U13095 ( .A(n20536), .B(n20326), .ZN(n20091) );
  NAND2_X1 U13096 ( .A1(n20091), .A2(n11205), .ZN(n10283) );
  AOI22_X1 U13097 ( .A1(n9624), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n10504), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n10289) );
  AOI22_X1 U13098 ( .A1(n11036), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n10682), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n10288) );
  AOI22_X1 U13099 ( .A1(n10768), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n9622), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n10287) );
  AOI22_X1 U13100 ( .A1(n11035), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n11042), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n10286) );
  NAND4_X1 U13101 ( .A1(n10289), .A2(n10288), .A3(n10287), .A4(n10286), .ZN(
        n10297) );
  AOI22_X1 U13102 ( .A1(n10458), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n10187), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n10295) );
  INV_X2 U13103 ( .A(n10318), .ZN(n10387) );
  AOI22_X1 U13104 ( .A1(n10387), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n11041), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n10294) );
  AOI22_X1 U13105 ( .A1(n10972), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n9628), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n10293) );
  AOI22_X1 U13106 ( .A1(n9619), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n10213), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n10292) );
  NAND4_X1 U13107 ( .A1(n10295), .A2(n10294), .A3(n10293), .A4(n10292), .ZN(
        n10296) );
  NOR2_X1 U13108 ( .A1(n10297), .A2(n10296), .ZN(n11123) );
  INV_X1 U13109 ( .A(n10340), .ZN(n10839) );
  NAND2_X1 U13110 ( .A1(n20086), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n10327) );
  NOR2_X1 U13111 ( .A1(n10327), .A2(n11123), .ZN(n10298) );
  INV_X1 U13112 ( .A(n10364), .ZN(n10301) );
  AOI22_X1 U13113 ( .A1(n10458), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n9618), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n10306) );
  AOI22_X1 U13114 ( .A1(n9624), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n10504), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n10305) );
  AOI22_X1 U13115 ( .A1(n11036), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n10682), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10304) );
  AOI22_X1 U13116 ( .A1(n9628), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n10213), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n10303) );
  NAND4_X1 U13117 ( .A1(n10306), .A2(n10305), .A3(n10304), .A4(n10303), .ZN(
        n10312) );
  AOI22_X1 U13118 ( .A1(n10387), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n10972), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n10310) );
  AOI22_X1 U13119 ( .A1(n10768), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n9621), .B2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n10309) );
  AOI22_X1 U13120 ( .A1(n10484), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n11041), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n10308) );
  AOI22_X1 U13121 ( .A1(n10171), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n11042), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n10307) );
  NAND4_X1 U13122 ( .A1(n10310), .A2(n10309), .A3(n10308), .A4(n10307), .ZN(
        n10311) );
  NAND2_X1 U13123 ( .A1(n10340), .A2(n11104), .ZN(n10313) );
  INV_X1 U13124 ( .A(n11104), .ZN(n11110) );
  AOI22_X1 U13125 ( .A1(n9625), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n10504), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n10317) );
  AOI22_X1 U13126 ( .A1(n11036), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n10682), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n10316) );
  AOI22_X1 U13127 ( .A1(n10768), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n9620), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n10315) );
  AOI22_X1 U13128 ( .A1(n10171), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n11042), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n10314) );
  NAND4_X1 U13129 ( .A1(n10317), .A2(n10316), .A3(n10315), .A4(n10314), .ZN(
        n10325) );
  AOI22_X1 U13130 ( .A1(n10458), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n10484), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n10323) );
  AOI22_X1 U13131 ( .A1(n10387), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n11041), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n10322) );
  AOI22_X1 U13132 ( .A1(n10998), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n9638), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n10321) );
  AOI22_X1 U13133 ( .A1(n9617), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n10213), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n10320) );
  NAND4_X1 U13134 ( .A1(n10323), .A2(n10322), .A3(n10321), .A4(n10320), .ZN(
        n10324) );
  INV_X1 U13135 ( .A(n11170), .ZN(n10326) );
  NAND2_X1 U13136 ( .A1(n10340), .A2(n10326), .ZN(n10342) );
  OAI21_X1 U13137 ( .B1(n11110), .B2(n10327), .A(n10342), .ZN(n10329) );
  AND2_X1 U13138 ( .A1(n10862), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n10328) );
  AOI22_X1 U13139 ( .A1(n10387), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n10734), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n10333) );
  AOI22_X1 U13140 ( .A1(n9624), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n10504), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n10332) );
  AOI22_X1 U13141 ( .A1(n10682), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n11035), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n10331) );
  AOI22_X1 U13142 ( .A1(n9628), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n10213), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n10330) );
  NAND4_X1 U13143 ( .A1(n10333), .A2(n10332), .A3(n10331), .A4(n10330), .ZN(
        n10339) );
  AOI22_X1 U13144 ( .A1(n9616), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n10972), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n10337) );
  AOI22_X1 U13145 ( .A1(n10768), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n9622), .B2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n10336) );
  AOI22_X1 U13146 ( .A1(n10484), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n11041), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n10335) );
  AOI22_X1 U13147 ( .A1(n11036), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n11042), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n10334) );
  NAND4_X1 U13148 ( .A1(n10337), .A2(n10336), .A3(n10335), .A4(n10334), .ZN(
        n10338) );
  NOR2_X1 U13149 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n10341), .ZN(n10344) );
  NOR2_X1 U13150 ( .A1(n10342), .A2(n11109), .ZN(n10343) );
  AOI211_X1 U13151 ( .C1(n11109), .C2(n11101), .A(n10344), .B(n10343), .ZN(
        n10360) );
  NAND2_X1 U13152 ( .A1(n20107), .A2(n11170), .ZN(n10345) );
  OAI211_X1 U13153 ( .C1(n11109), .C2(n19946), .A(P1_STATE2_REG_0__SCAN_IN), 
        .B(n10345), .ZN(n10346) );
  AOI21_X1 U13154 ( .B1(P1_INSTQUEUE_REG_0__0__SCAN_IN), .B2(n10849), .A(
        n10346), .ZN(n10359) );
  NOR2_X1 U13155 ( .A1(n10360), .A2(n10359), .ZN(n10347) );
  NAND2_X1 U13156 ( .A1(n10349), .A2(n10348), .ZN(n10350) );
  INV_X2 U13157 ( .A(P1_STATE2_REG_2__SCAN_IN), .ZN(n20599) );
  NOR2_X1 U13158 ( .A1(n13384), .A2(n20599), .ZN(n10427) );
  INV_X1 U13159 ( .A(P1_EAX_REG_2__SCAN_IN), .ZN(n10355) );
  NAND2_X1 U13160 ( .A1(n20599), .A2(n20891), .ZN(n10404) );
  XNOR2_X1 U13161 ( .A(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .B(
        P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n14303) );
  AOI21_X1 U13162 ( .B1(n11054), .B2(n14303), .A(n11060), .ZN(n10354) );
  OAI21_X1 U13163 ( .B1(n11008), .B2(n10355), .A(n10354), .ZN(n10356) );
  AOI21_X1 U13164 ( .B1(n10427), .B2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(
        n10356), .ZN(n10357) );
  NAND2_X1 U13165 ( .A1(n11060), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n10379) );
  XOR2_X1 U13166 ( .A(n10360), .B(n10359), .Z(n20701) );
  INV_X1 U13167 ( .A(n20701), .ZN(n20149) );
  AOI21_X1 U13168 ( .B1(n10274), .B2(n20149), .A(n20599), .ZN(n13150) );
  NOR2_X1 U13169 ( .A1(n10362), .A2(n10361), .ZN(n10363) );
  OR2_X1 U13170 ( .A1(n10364), .A2(n10363), .ZN(n20181) );
  OR2_X1 U13171 ( .A1(n20181), .A2(n10580), .ZN(n10369) );
  INV_X1 U13172 ( .A(P1_EAX_REG_0__SCAN_IN), .ZN(n10366) );
  NAND2_X1 U13173 ( .A1(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n20599), .ZN(
        n10365) );
  OAI21_X1 U13174 ( .B1(n11008), .B2(n10366), .A(n10365), .ZN(n10367) );
  AOI21_X1 U13175 ( .B1(n10427), .B2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A(
        n10367), .ZN(n10368) );
  NAND2_X1 U13176 ( .A1(n10369), .A2(n10368), .ZN(n13149) );
  NAND2_X1 U13177 ( .A1(n13150), .A2(n13149), .ZN(n13148) );
  INV_X1 U13178 ( .A(n13149), .ZN(n10370) );
  NAND2_X1 U13179 ( .A1(n10370), .A2(n11054), .ZN(n10371) );
  NAND2_X1 U13180 ( .A1(n13148), .A2(n10371), .ZN(n13127) );
  NAND2_X1 U13181 ( .A1(n13433), .A2(n10609), .ZN(n10377) );
  INV_X1 U13182 ( .A(P1_EAX_REG_1__SCAN_IN), .ZN(n10374) );
  NAND2_X1 U13183 ( .A1(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n20599), .ZN(
        n10373) );
  OAI21_X1 U13184 ( .B1(n11008), .B2(n10374), .A(n10373), .ZN(n10375) );
  AOI21_X1 U13185 ( .B1(n10427), .B2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(
        n10375), .ZN(n10376) );
  NAND2_X1 U13186 ( .A1(n10377), .A2(n10376), .ZN(n13126) );
  NAND2_X1 U13187 ( .A1(n13127), .A2(n13126), .ZN(n13140) );
  NAND2_X1 U13188 ( .A1(n9741), .A2(n10378), .ZN(n13141) );
  INV_X1 U13189 ( .A(n10282), .ZN(n10380) );
  NAND2_X1 U13190 ( .A1(n10380), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10386) );
  NAND2_X1 U13191 ( .A1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n20536), .ZN(
        n10382) );
  NAND2_X1 U13192 ( .A1(n20690), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n20264) );
  NOR2_X1 U13193 ( .A1(n10381), .A2(n20264), .ZN(n20317) );
  AOI21_X1 U13194 ( .B1(n10382), .B2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A(
        n20317), .ZN(n20327) );
  INV_X1 U13195 ( .A(n15362), .ZN(n15371) );
  OAI22_X1 U13196 ( .A1(n20327), .A2(n10383), .B1(n15371), .B2(n20690), .ZN(
        n10384) );
  INV_X1 U13197 ( .A(n10384), .ZN(n10385) );
  XNOR2_X2 U13198 ( .A(n13424), .B(n20214), .ZN(n20684) );
  AOI22_X1 U13199 ( .A1(n9619), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n10972), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10391) );
  AOI22_X1 U13200 ( .A1(n10387), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n10734), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n10390) );
  AOI22_X1 U13201 ( .A1(n11036), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n10682), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10389) );
  AOI22_X1 U13202 ( .A1(n9621), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n10208), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n10388) );
  NAND4_X1 U13203 ( .A1(n10391), .A2(n10390), .A3(n10389), .A4(n10388), .ZN(
        n10397) );
  INV_X1 U13204 ( .A(n10226), .ZN(n10434) );
  AOI22_X1 U13205 ( .A1(n9624), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n10504), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n10395) );
  AOI22_X1 U13206 ( .A1(n10768), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n11035), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n10394) );
  AOI22_X1 U13207 ( .A1(n10484), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n11041), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n10393) );
  AOI22_X1 U13208 ( .A1(n9628), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n10213), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n10392) );
  NAND4_X1 U13209 ( .A1(n10395), .A2(n10394), .A3(n10393), .A4(n10392), .ZN(
        n10396) );
  AOI22_X1 U13210 ( .A1(n10866), .A2(n11130), .B1(n10862), .B2(
        P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n10398) );
  NAND2_X1 U13211 ( .A1(n10400), .A2(n20213), .ZN(n10402) );
  INV_X1 U13212 ( .A(n20213), .ZN(n10401) );
  NAND2_X1 U13213 ( .A1(n10402), .A2(n10424), .ZN(n20683) );
  INV_X1 U13214 ( .A(P1_EAX_REG_3__SCAN_IN), .ZN(n10407) );
  AOI21_X1 U13215 ( .B1(n10403), .B2(n19908), .A(n10426), .ZN(n19911) );
  INV_X1 U13216 ( .A(n11060), .ZN(n10586) );
  OAI22_X1 U13217 ( .A1(n19911), .A2(n10404), .B1(n10586), .B2(n19908), .ZN(
        n10405) );
  INV_X1 U13218 ( .A(n10405), .ZN(n10406) );
  OAI21_X1 U13219 ( .B1(n11008), .B2(n10407), .A(n10406), .ZN(n10408) );
  AOI21_X1 U13220 ( .B1(n10427), .B2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n10408), .ZN(n10409) );
  AOI22_X1 U13221 ( .A1(n9624), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n10504), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n10413) );
  AOI22_X1 U13222 ( .A1(n11036), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n10682), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n10412) );
  AOI22_X1 U13223 ( .A1(n10768), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n9620), .B2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n10411) );
  AOI22_X1 U13224 ( .A1(n11035), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n10208), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n10410) );
  NAND4_X1 U13225 ( .A1(n10413), .A2(n10412), .A3(n10411), .A4(n10410), .ZN(
        n10419) );
  AOI22_X1 U13226 ( .A1(n10458), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n10187), .B2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n10417) );
  AOI22_X1 U13227 ( .A1(n10387), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n11041), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n10416) );
  AOI22_X1 U13228 ( .A1(n10972), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n9638), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n10415) );
  AOI22_X1 U13229 ( .A1(n9619), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n10213), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n10414) );
  NAND4_X1 U13230 ( .A1(n10417), .A2(n10416), .A3(n10415), .A4(n10414), .ZN(
        n10418) );
  INV_X1 U13231 ( .A(n11139), .ZN(n10420) );
  OR2_X1 U13232 ( .A1(n10837), .A2(n10420), .ZN(n10422) );
  NAND2_X1 U13233 ( .A1(n10862), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n10421) );
  INV_X1 U13234 ( .A(n10466), .ZN(n10425) );
  NAND2_X1 U13235 ( .A1(n10425), .A2(n10130), .ZN(n11142) );
  OAI21_X1 U13236 ( .B1(n10426), .B2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n10447), .ZN(n19896) );
  INV_X1 U13237 ( .A(n10427), .ZN(n10431) );
  INV_X1 U13238 ( .A(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n10428) );
  AOI21_X1 U13239 ( .B1(P1_STATEBS16_REG_SCAN_IN), .B2(n10428), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n10429) );
  AOI21_X1 U13240 ( .B1(n11061), .B2(P1_EAX_REG_4__SCAN_IN), .A(n10429), .ZN(
        n10430) );
  OAI21_X1 U13241 ( .B1(n15861), .B2(n10431), .A(n10430), .ZN(n10432) );
  OAI21_X1 U13242 ( .B1(n19896), .B2(n10404), .A(n10432), .ZN(n10433) );
  INV_X2 U13243 ( .A(n10434), .ZN(n10504) );
  AOI22_X1 U13244 ( .A1(n9624), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n10504), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n10438) );
  AOI22_X1 U13245 ( .A1(n11036), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n10682), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10437) );
  AOI22_X1 U13246 ( .A1(P1_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n10171), .B1(
        n9622), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n10436) );
  AOI22_X1 U13247 ( .A1(n10998), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n10213), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n10435) );
  NAND4_X1 U13248 ( .A1(n10438), .A2(n10437), .A3(n10436), .A4(n10435), .ZN(
        n10444) );
  AOI22_X1 U13249 ( .A1(P1_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n10734), .B1(
        n10484), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n10442) );
  AOI22_X1 U13250 ( .A1(n9616), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n9628), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n10441) );
  AOI22_X1 U13251 ( .A1(n10387), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n11041), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n10440) );
  AOI22_X1 U13252 ( .A1(n10768), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n10208), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n10439) );
  NAND4_X1 U13253 ( .A1(n10442), .A2(n10441), .A3(n10440), .A4(n10439), .ZN(
        n10443) );
  NOR2_X1 U13254 ( .A1(n10444), .A2(n10443), .ZN(n11149) );
  INV_X1 U13255 ( .A(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n10445) );
  OAI22_X1 U13256 ( .A1(n11149), .A2(n10837), .B1(n10858), .B2(n10445), .ZN(
        n10465) );
  INV_X1 U13257 ( .A(n10465), .ZN(n10446) );
  XNOR2_X1 U13258 ( .A(n10466), .B(n10446), .ZN(n11147) );
  NAND2_X1 U13259 ( .A1(n11147), .A2(n10609), .ZN(n10453) );
  NAND2_X1 U13260 ( .A1(n10447), .A2(n15664), .ZN(n10449) );
  INV_X1 U13261 ( .A(n10467), .ZN(n10448) );
  NAND2_X1 U13262 ( .A1(n10449), .A2(n10448), .ZN(n19889) );
  NAND2_X1 U13263 ( .A1(n19889), .A2(n11054), .ZN(n10450) );
  OAI21_X1 U13264 ( .B1(n10586), .B2(n15664), .A(n10450), .ZN(n10451) );
  AOI21_X1 U13265 ( .B1(n11061), .B2(P1_EAX_REG_5__SCAN_IN), .A(n10451), .ZN(
        n10452) );
  NAND2_X1 U13266 ( .A1(n13372), .A2(n13458), .ZN(n13457) );
  AOI22_X1 U13267 ( .A1(n9624), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n10504), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n10457) );
  AOI22_X1 U13268 ( .A1(n11036), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n10682), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n10456) );
  AOI22_X1 U13269 ( .A1(n10768), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n9620), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n10455) );
  AOI22_X1 U13270 ( .A1(n10171), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n10208), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n10454) );
  NAND4_X1 U13271 ( .A1(n10457), .A2(n10456), .A3(n10455), .A4(n10454), .ZN(
        n10464) );
  AOI22_X1 U13272 ( .A1(n10458), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n10484), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n10462) );
  AOI22_X1 U13273 ( .A1(n10387), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n11041), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n10461) );
  AOI22_X1 U13274 ( .A1(n10998), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n9638), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n10460) );
  AOI22_X1 U13275 ( .A1(n9617), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n10213), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n10459) );
  NAND4_X1 U13276 ( .A1(n10462), .A2(n10461), .A3(n10460), .A4(n10459), .ZN(
        n10463) );
  OR2_X1 U13277 ( .A1(n10464), .A2(n10463), .ZN(n11158) );
  AOI22_X1 U13278 ( .A1(n10862), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n10866), .B2(n11158), .ZN(n10473) );
  NAND2_X1 U13279 ( .A1(n10473), .A2(n10474), .ZN(n11155) );
  NAND2_X1 U13280 ( .A1(n11155), .A2(n10609), .ZN(n10471) );
  INV_X1 U13281 ( .A(P1_EAX_REG_6__SCAN_IN), .ZN(n13751) );
  OAI21_X1 U13282 ( .B1(n10467), .B2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .A(
        n10477), .ZN(n19874) );
  AOI22_X1 U13283 ( .A1(n11054), .A2(n19874), .B1(n11060), .B2(
        P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n10468) );
  OAI21_X1 U13284 ( .B1(n11008), .B2(n13751), .A(n10468), .ZN(n10469) );
  INV_X1 U13285 ( .A(n10469), .ZN(n10470) );
  AOI22_X1 U13286 ( .A1(n10862), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n10866), .B2(n11170), .ZN(n10475) );
  INV_X1 U13287 ( .A(P1_EAX_REG_7__SCAN_IN), .ZN(n10480) );
  OAI21_X1 U13288 ( .B1(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n10478), .A(
        n10500), .ZN(n19854) );
  AOI22_X1 U13289 ( .A1(n11054), .A2(n19854), .B1(n11060), .B2(
        P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n10479) );
  OAI21_X1 U13290 ( .B1(n11008), .B2(n10480), .A(n10479), .ZN(n10481) );
  INV_X1 U13291 ( .A(n10481), .ZN(n10482) );
  INV_X1 U13292 ( .A(P1_EAX_REG_8__SCAN_IN), .ZN(n13726) );
  AOI22_X1 U13293 ( .A1(n10734), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n10484), .B2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n10489) );
  AOI22_X1 U13294 ( .A1(n11036), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n10504), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n10488) );
  AOI22_X1 U13295 ( .A1(n10682), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n11035), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n10487) );
  AOI22_X1 U13296 ( .A1(n10387), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n11041), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n10486) );
  NAND4_X1 U13297 ( .A1(n10489), .A2(n10488), .A3(n10487), .A4(n10486), .ZN(
        n10498) );
  AOI22_X1 U13298 ( .A1(n10768), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n9622), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n10496) );
  AOI22_X1 U13299 ( .A1(n10972), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n9638), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n10495) );
  AOI22_X1 U13300 ( .A1(n9624), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n11042), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n10494) );
  AOI22_X1 U13301 ( .A1(n9619), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n10213), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n10493) );
  NAND4_X1 U13302 ( .A1(n10496), .A2(n10495), .A3(n10494), .A4(n10493), .ZN(
        n10497) );
  OR2_X1 U13303 ( .A1(n10498), .A2(n10497), .ZN(n10499) );
  NAND2_X1 U13304 ( .A1(n10609), .A2(n10499), .ZN(n10502) );
  XNOR2_X1 U13305 ( .A(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .B(n10503), .ZN(
        n13758) );
  AOI22_X1 U13306 ( .A1(n11054), .A2(n13758), .B1(n11060), .B2(
        P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n10501) );
  OAI211_X1 U13307 ( .C1(n11008), .C2(n13726), .A(n10502), .B(n10501), .ZN(
        n13656) );
  NAND2_X1 U13308 ( .A1(n13579), .A2(n13656), .ZN(n13655) );
  INV_X1 U13309 ( .A(n13655), .ZN(n10520) );
  XNOR2_X1 U13310 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .B(n10522), .ZN(
        n19842) );
  INV_X1 U13311 ( .A(n19842), .ZN(n14038) );
  AOI22_X1 U13312 ( .A1(n9624), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n10734), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n10508) );
  AOI22_X1 U13313 ( .A1(n10504), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n10682), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n10507) );
  AOI22_X1 U13314 ( .A1(n10768), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n11035), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10506) );
  AOI22_X1 U13315 ( .A1(n10484), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n9628), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n10505) );
  NAND4_X1 U13316 ( .A1(n10508), .A2(n10507), .A3(n10506), .A4(n10505), .ZN(
        n10514) );
  AOI22_X1 U13317 ( .A1(n10387), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n9618), .B2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n10512) );
  AOI22_X1 U13318 ( .A1(n11036), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n11041), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n10511) );
  AOI22_X1 U13319 ( .A1(n9621), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n11042), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n10510) );
  AOI22_X1 U13320 ( .A1(n10972), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n10213), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n10509) );
  NAND4_X1 U13321 ( .A1(n10512), .A2(n10511), .A3(n10510), .A4(n10509), .ZN(
        n10513) );
  NOR2_X1 U13322 ( .A1(n10514), .A2(n10513), .ZN(n10517) );
  NAND2_X1 U13323 ( .A1(n11061), .A2(P1_EAX_REG_9__SCAN_IN), .ZN(n10516) );
  NAND2_X1 U13324 ( .A1(n11060), .A2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n10515) );
  OAI211_X1 U13325 ( .C1(n10580), .C2(n10517), .A(n10516), .B(n10515), .ZN(
        n10518) );
  AOI21_X1 U13326 ( .B1(n14038), .B2(n11054), .A(n10518), .ZN(n13769) );
  INV_X1 U13327 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n10521) );
  XNOR2_X1 U13328 ( .A(n10537), .B(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n14544) );
  AOI22_X1 U13329 ( .A1(n10734), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n10484), .B2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n10526) );
  AOI22_X1 U13330 ( .A1(n11036), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n10504), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n10525) );
  AOI22_X1 U13331 ( .A1(n10768), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n11035), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n10524) );
  AOI22_X1 U13332 ( .A1(n10972), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n10213), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n10523) );
  NAND4_X1 U13333 ( .A1(n10526), .A2(n10525), .A3(n10524), .A4(n10523), .ZN(
        n10532) );
  AOI22_X1 U13334 ( .A1(n9624), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n10682), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n10530) );
  AOI22_X1 U13335 ( .A1(n9619), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n9628), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n10529) );
  AOI22_X1 U13336 ( .A1(n10387), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n11041), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n10528) );
  AOI22_X1 U13337 ( .A1(n9622), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n11042), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n10527) );
  NAND4_X1 U13338 ( .A1(n10530), .A2(n10529), .A3(n10528), .A4(n10527), .ZN(
        n10531) );
  NOR2_X1 U13339 ( .A1(n10532), .A2(n10531), .ZN(n10535) );
  NAND2_X1 U13340 ( .A1(n11060), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n10534) );
  NAND2_X1 U13341 ( .A1(n11061), .A2(P1_EAX_REG_10__SCAN_IN), .ZN(n10533) );
  OAI211_X1 U13342 ( .C1(n10580), .C2(n10535), .A(n10534), .B(n10533), .ZN(
        n10536) );
  AOI21_X1 U13343 ( .B1(n14544), .B2(n11054), .A(n10536), .ZN(n13783) );
  INV_X1 U13344 ( .A(P1_EAX_REG_11__SCAN_IN), .ZN(n14087) );
  OAI21_X1 U13345 ( .B1(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n10538), .A(
        n10567), .ZN(n15648) );
  AOI22_X1 U13346 ( .A1(n11054), .A2(n15648), .B1(n11060), .B2(
        P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n10539) );
  OAI21_X1 U13347 ( .B1(n11008), .B2(n14087), .A(n10539), .ZN(n14085) );
  AOI22_X1 U13348 ( .A1(n9619), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n10972), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n10543) );
  AOI22_X1 U13349 ( .A1(n9625), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n10484), .B2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n10542) );
  AOI22_X1 U13350 ( .A1(n11036), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n10682), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n10541) );
  AOI22_X1 U13351 ( .A1(n10768), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n9620), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n10540) );
  NAND4_X1 U13352 ( .A1(n10543), .A2(n10542), .A3(n10541), .A4(n10540), .ZN(
        n10549) );
  AOI22_X1 U13353 ( .A1(n10734), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n10504), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10547) );
  AOI22_X1 U13354 ( .A1(n10387), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n11041), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n10546) );
  AOI22_X1 U13355 ( .A1(n11035), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n11042), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n10545) );
  AOI22_X1 U13356 ( .A1(n9628), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n10213), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n10544) );
  NAND4_X1 U13357 ( .A1(n10547), .A2(n10546), .A3(n10545), .A4(n10544), .ZN(
        n10548) );
  NOR2_X1 U13358 ( .A1(n10549), .A2(n10548), .ZN(n10550) );
  NOR2_X1 U13359 ( .A1(n10580), .A2(n10550), .ZN(n14089) );
  INV_X1 U13360 ( .A(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n10551) );
  XNOR2_X1 U13361 ( .A(n10584), .B(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n14537) );
  NAND2_X1 U13362 ( .A1(n14537), .A2(n11054), .ZN(n10566) );
  AOI22_X1 U13363 ( .A1(n9617), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n10972), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n10555) );
  AOI22_X1 U13364 ( .A1(P1_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n10387), .B1(
        n9624), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n10554) );
  AOI22_X1 U13365 ( .A1(n10768), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n9622), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n10553) );
  AOI22_X1 U13366 ( .A1(P1_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n10682), .B1(
        n11042), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n10552) );
  NAND4_X1 U13367 ( .A1(n10555), .A2(n10554), .A3(n10553), .A4(n10552), .ZN(
        n10561) );
  AOI22_X1 U13368 ( .A1(n10734), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n10504), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10559) );
  AOI22_X1 U13369 ( .A1(n11036), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n11035), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10558) );
  AOI22_X1 U13370 ( .A1(n10484), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n11041), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n10557) );
  AOI22_X1 U13371 ( .A1(n9628), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n10213), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n10556) );
  NAND4_X1 U13372 ( .A1(n10559), .A2(n10558), .A3(n10557), .A4(n10556), .ZN(
        n10560) );
  OR2_X1 U13373 ( .A1(n10561), .A2(n10560), .ZN(n10564) );
  INV_X1 U13374 ( .A(P1_EAX_REG_13__SCAN_IN), .ZN(n14141) );
  INV_X1 U13375 ( .A(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n10562) );
  OAI22_X1 U13376 ( .A1(n11008), .A2(n14141), .B1(n10586), .B2(n10562), .ZN(
        n10563) );
  AOI21_X1 U13377 ( .B1(n10609), .B2(n10564), .A(n10563), .ZN(n10565) );
  NAND2_X1 U13378 ( .A1(n10566), .A2(n10565), .ZN(n14122) );
  XNOR2_X1 U13379 ( .A(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B(n10567), .ZN(
        n15634) );
  OAI22_X1 U13380 ( .A1(n15634), .A2(n10404), .B1(n10586), .B2(n10551), .ZN(
        n10568) );
  AOI21_X1 U13381 ( .B1(n11061), .B2(P1_EAX_REG_12__SCAN_IN), .A(n10568), .ZN(
        n10582) );
  AOI22_X1 U13382 ( .A1(n9624), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n10734), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n10572) );
  AOI22_X1 U13383 ( .A1(n10504), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n10682), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n10571) );
  AOI22_X1 U13384 ( .A1(n10387), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n9628), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n10570) );
  AOI22_X1 U13385 ( .A1(n11035), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n11042), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n10569) );
  NAND4_X1 U13386 ( .A1(n10572), .A2(n10571), .A3(n10570), .A4(n10569), .ZN(
        n10578) );
  AOI22_X1 U13387 ( .A1(n11036), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n10484), .B2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n10576) );
  AOI22_X1 U13388 ( .A1(n10768), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n9621), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n10575) );
  AOI22_X1 U13389 ( .A1(n9618), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n11041), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n10574) );
  AOI22_X1 U13390 ( .A1(n10972), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n10213), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n10573) );
  NAND4_X1 U13391 ( .A1(n10576), .A2(n10575), .A3(n10574), .A4(n10573), .ZN(
        n10577) );
  NOR2_X1 U13392 ( .A1(n10578), .A2(n10577), .ZN(n10579) );
  OR2_X1 U13393 ( .A1(n10580), .A2(n10579), .ZN(n10581) );
  NAND2_X1 U13394 ( .A1(n10582), .A2(n10581), .ZN(n14093) );
  NAND2_X1 U13395 ( .A1(n14122), .A2(n14093), .ZN(n10583) );
  XNOR2_X1 U13396 ( .A(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .B(n10600), .ZN(
        n15625) );
  INV_X1 U13397 ( .A(P1_EAX_REG_14__SCAN_IN), .ZN(n14113) );
  INV_X1 U13398 ( .A(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n10585) );
  OAI22_X1 U13399 ( .A1(n11008), .A2(n14113), .B1(n10586), .B2(n10585), .ZN(
        n10587) );
  INV_X1 U13400 ( .A(n10587), .ZN(n10599) );
  AOI22_X1 U13401 ( .A1(n10768), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n9621), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n10591) );
  AOI22_X1 U13402 ( .A1(n10504), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n11041), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n10590) );
  AOI22_X1 U13403 ( .A1(n11035), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n11042), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n10589) );
  AOI22_X1 U13404 ( .A1(n10387), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n10213), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n10588) );
  NAND4_X1 U13405 ( .A1(n10591), .A2(n10590), .A3(n10589), .A4(n10588), .ZN(
        n10597) );
  AOI22_X1 U13406 ( .A1(n9618), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n10484), .B2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n10595) );
  AOI22_X1 U13407 ( .A1(n9624), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n10734), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n10594) );
  AOI22_X1 U13408 ( .A1(n11036), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n10682), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n10593) );
  AOI22_X1 U13409 ( .A1(n10972), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n9628), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n10592) );
  NAND4_X1 U13410 ( .A1(n10595), .A2(n10594), .A3(n10593), .A4(n10592), .ZN(
        n10596) );
  OAI21_X1 U13411 ( .B1(n10597), .B2(n10596), .A(n10609), .ZN(n10598) );
  OAI211_X1 U13412 ( .C1(n15625), .C2(n10404), .A(n10599), .B(n10598), .ZN(
        n14101) );
  XNOR2_X1 U13413 ( .A(n10624), .B(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n14525) );
  AOI22_X1 U13414 ( .A1(n11061), .A2(P1_EAX_REG_15__SCAN_IN), .B1(n11060), 
        .B2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n10613) );
  AOI22_X1 U13415 ( .A1(n10734), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n10484), .B2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n10604) );
  AOI22_X1 U13416 ( .A1(n9624), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n10682), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n10603) );
  AOI22_X1 U13417 ( .A1(n10171), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n9620), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n10602) );
  AOI22_X1 U13418 ( .A1(n9638), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n10213), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n10601) );
  NAND4_X1 U13419 ( .A1(n10604), .A2(n10603), .A3(n10602), .A4(n10601), .ZN(
        n10611) );
  AOI22_X1 U13420 ( .A1(n9617), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n10972), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n10608) );
  AOI22_X1 U13421 ( .A1(n11036), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n10504), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n10607) );
  AOI22_X1 U13422 ( .A1(n10387), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n11041), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n10606) );
  AOI22_X1 U13423 ( .A1(n10768), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n11042), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n10605) );
  NAND4_X1 U13424 ( .A1(n10608), .A2(n10607), .A3(n10606), .A4(n10605), .ZN(
        n10610) );
  OAI21_X1 U13425 ( .B1(n10611), .B2(n10610), .A(n10609), .ZN(n10612) );
  OAI211_X1 U13426 ( .C1(n14525), .C2(n10404), .A(n10613), .B(n10612), .ZN(
        n14116) );
  AOI22_X1 U13427 ( .A1(n9619), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n10972), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n10617) );
  AOI22_X1 U13428 ( .A1(n10734), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n10682), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n10616) );
  AOI22_X1 U13429 ( .A1(n10768), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n11035), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n10615) );
  AOI22_X1 U13430 ( .A1(n10387), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n11041), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10614) );
  NAND4_X1 U13431 ( .A1(n10617), .A2(n10616), .A3(n10615), .A4(n10614), .ZN(
        n10623) );
  AOI22_X1 U13432 ( .A1(n9624), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n10484), .B2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n10621) );
  AOI22_X1 U13433 ( .A1(n11036), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n10504), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n10620) );
  AOI22_X1 U13434 ( .A1(n9628), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n10213), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n10619) );
  AOI22_X1 U13435 ( .A1(n9622), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n10208), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n10618) );
  NAND4_X1 U13436 ( .A1(n10621), .A2(n10620), .A3(n10619), .A4(n10618), .ZN(
        n10622) );
  OR2_X1 U13437 ( .A1(n10623), .A2(n10622), .ZN(n10628) );
  INV_X1 U13438 ( .A(P1_EAX_REG_17__SCAN_IN), .ZN(n14426) );
  INV_X1 U13439 ( .A(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n14290) );
  INV_X1 U13440 ( .A(n10648), .ZN(n10625) );
  XNOR2_X1 U13441 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .B(n10625), .ZN(
        n14508) );
  AOI22_X1 U13442 ( .A1(n11054), .A2(n14508), .B1(n11060), .B2(
        P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n10626) );
  OAI21_X1 U13443 ( .B1(n11008), .B2(n14426), .A(n10626), .ZN(n10627) );
  AOI21_X1 U13444 ( .B1(n11030), .B2(n10628), .A(n10627), .ZN(n14272) );
  AOI22_X1 U13445 ( .A1(n10387), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n10734), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n10632) );
  AOI22_X1 U13446 ( .A1(n11036), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n10504), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n10631) );
  AOI22_X1 U13447 ( .A1(n10682), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n9622), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n10630) );
  AOI22_X1 U13448 ( .A1(n10972), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n9628), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n10629) );
  NAND4_X1 U13449 ( .A1(n10632), .A2(n10631), .A3(n10630), .A4(n10629), .ZN(
        n10638) );
  AOI22_X1 U13450 ( .A1(n9625), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n10171), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n10636) );
  AOI22_X1 U13451 ( .A1(n10484), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n11041), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n10635) );
  AOI22_X1 U13452 ( .A1(n10768), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n11042), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n10634) );
  AOI22_X1 U13453 ( .A1(n9616), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n10213), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n10633) );
  NAND4_X1 U13454 ( .A1(n10636), .A2(n10635), .A3(n10634), .A4(n10633), .ZN(
        n10637) );
  NOR2_X1 U13455 ( .A1(n10638), .A2(n10637), .ZN(n10642) );
  INV_X1 U13456 ( .A(P1_EAX_REG_16__SCAN_IN), .ZN(n19974) );
  OAI21_X1 U13457 ( .B1(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n20891), .A(
        n20599), .ZN(n10639) );
  OAI21_X1 U13458 ( .B1(n11008), .B2(n19974), .A(n10639), .ZN(n10640) );
  INV_X1 U13459 ( .A(n10640), .ZN(n10641) );
  OAI21_X1 U13460 ( .B1(n11057), .B2(n10642), .A(n10641), .ZN(n10645) );
  OAI21_X1 U13461 ( .B1(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n10643), .A(
        n10648), .ZN(n15610) );
  OR2_X1 U13462 ( .A1(n10404), .A2(n15610), .ZN(n10644) );
  NAND2_X1 U13463 ( .A1(n10645), .A2(n10644), .ZN(n14435) );
  INV_X1 U13464 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n10647) );
  OR2_X1 U13465 ( .A1(n10649), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n10650) );
  NAND2_X1 U13466 ( .A1(n10650), .A2(n10698), .ZN(n15605) );
  AOI22_X1 U13467 ( .A1(n10768), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n9621), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n10654) );
  AOI22_X1 U13468 ( .A1(n10972), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n9638), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n10653) );
  AOI22_X1 U13469 ( .A1(n10171), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n10208), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n10652) );
  AOI22_X1 U13470 ( .A1(n11041), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n10213), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n10651) );
  NAND4_X1 U13471 ( .A1(n10654), .A2(n10653), .A3(n10652), .A4(n10651), .ZN(
        n10660) );
  AOI22_X1 U13472 ( .A1(n10387), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n9617), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n10658) );
  AOI22_X1 U13473 ( .A1(n10734), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n10484), .B2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n10657) );
  AOI22_X1 U13474 ( .A1(n9625), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n10504), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n10656) );
  AOI22_X1 U13475 ( .A1(n11036), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n10682), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n10655) );
  NAND4_X1 U13476 ( .A1(n10658), .A2(n10657), .A3(n10656), .A4(n10655), .ZN(
        n10659) );
  OAI21_X1 U13477 ( .B1(n10660), .B2(n10659), .A(n11030), .ZN(n10663) );
  NAND2_X1 U13478 ( .A1(n11061), .A2(P1_EAX_REG_18__SCAN_IN), .ZN(n10662) );
  NAND2_X1 U13479 ( .A1(n20599), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n10661) );
  NAND4_X1 U13480 ( .A1(n10663), .A2(n10404), .A3(n10662), .A4(n10661), .ZN(
        n10664) );
  OAI21_X1 U13481 ( .B1(n15605), .B2(n10404), .A(n10664), .ZN(n14359) );
  INV_X1 U13482 ( .A(n14359), .ZN(n10665) );
  AOI22_X1 U13483 ( .A1(n9624), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n10768), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n10669) );
  AOI22_X1 U13484 ( .A1(n10734), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n10484), .B2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n10668) );
  AOI22_X1 U13485 ( .A1(n10387), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n11041), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10667) );
  AOI22_X1 U13486 ( .A1(n10972), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n10213), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n10666) );
  NAND4_X1 U13487 ( .A1(n10669), .A2(n10668), .A3(n10667), .A4(n10666), .ZN(
        n10675) );
  AOI22_X1 U13488 ( .A1(n11036), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n10504), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n10673) );
  AOI22_X1 U13489 ( .A1(n10682), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n10171), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n10672) );
  AOI22_X1 U13490 ( .A1(n9619), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n9628), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n10671) );
  AOI22_X1 U13491 ( .A1(n9621), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n11042), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10670) );
  NAND4_X1 U13492 ( .A1(n10673), .A2(n10672), .A3(n10671), .A4(n10670), .ZN(
        n10674) );
  NOR2_X1 U13493 ( .A1(n10675), .A2(n10674), .ZN(n10679) );
  INV_X1 U13494 ( .A(P1_EAX_REG_19__SCAN_IN), .ZN(n14415) );
  NAND2_X1 U13495 ( .A1(n20599), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n10676) );
  OAI211_X1 U13496 ( .C1(n11008), .C2(n14415), .A(n10404), .B(n10676), .ZN(
        n10677) );
  INV_X1 U13497 ( .A(n10677), .ZN(n10678) );
  OAI21_X1 U13498 ( .B1(n11057), .B2(n10679), .A(n10678), .ZN(n10681) );
  XNOR2_X1 U13499 ( .A(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .B(n10698), .ZN(
        n14494) );
  NAND2_X1 U13500 ( .A1(n11054), .A2(n14494), .ZN(n10680) );
  AOI22_X1 U13501 ( .A1(n10504), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n10682), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n10686) );
  AOI22_X1 U13502 ( .A1(n10768), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n9622), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n10685) );
  AOI22_X1 U13503 ( .A1(n9616), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n9628), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n10684) );
  AOI22_X1 U13504 ( .A1(n10171), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n10208), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n10683) );
  NAND4_X1 U13505 ( .A1(n10686), .A2(n10685), .A3(n10684), .A4(n10683), .ZN(
        n10692) );
  AOI22_X1 U13506 ( .A1(n9625), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n10485), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n10690) );
  AOI22_X1 U13507 ( .A1(n10734), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n10484), .B2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n10689) );
  AOI22_X1 U13508 ( .A1(n10387), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n11041), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n10688) );
  AOI22_X1 U13509 ( .A1(n10998), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n10213), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n10687) );
  NAND4_X1 U13510 ( .A1(n10690), .A2(n10689), .A3(n10688), .A4(n10687), .ZN(
        n10691) );
  NOR2_X1 U13511 ( .A1(n10692), .A2(n10691), .ZN(n10696) );
  INV_X1 U13512 ( .A(P1_EAX_REG_20__SCAN_IN), .ZN(n19964) );
  OAI21_X1 U13513 ( .B1(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n20891), .A(
        n20599), .ZN(n10693) );
  OAI21_X1 U13514 ( .B1(n11008), .B2(n19964), .A(n10693), .ZN(n10694) );
  INV_X1 U13515 ( .A(n10694), .ZN(n10695) );
  OAI21_X1 U13516 ( .B1(n11057), .B2(n10696), .A(n10695), .ZN(n10701) );
  INV_X1 U13517 ( .A(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n10697) );
  OAI21_X1 U13518 ( .B1(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n10699), .A(
        n10717), .ZN(n15591) );
  OR2_X1 U13519 ( .A1(n10404), .A2(n15591), .ZN(n10700) );
  AOI22_X1 U13520 ( .A1(P1_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n10734), .B1(
        n9624), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n10705) );
  AOI22_X1 U13521 ( .A1(P1_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n11036), .B1(
        n10504), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n10704) );
  AOI22_X1 U13522 ( .A1(P1_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n10768), .B1(
        n11035), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n10703) );
  AOI22_X1 U13523 ( .A1(n10998), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n11041), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10702) );
  NAND4_X1 U13524 ( .A1(n10705), .A2(n10704), .A3(n10703), .A4(n10702), .ZN(
        n10711) );
  AOI22_X1 U13525 ( .A1(n10387), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n9618), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n10709) );
  AOI22_X1 U13526 ( .A1(P1_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n10682), .B1(
        n10484), .B2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n10708) );
  AOI22_X1 U13527 ( .A1(n9628), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n10213), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n10707) );
  AOI22_X1 U13528 ( .A1(P1_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n9620), .B1(
        n11042), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10706) );
  NAND4_X1 U13529 ( .A1(n10709), .A2(n10708), .A3(n10707), .A4(n10706), .ZN(
        n10710) );
  NOR2_X1 U13530 ( .A1(n10711), .A2(n10710), .ZN(n10714) );
  INV_X1 U13531 ( .A(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n15506) );
  AOI21_X1 U13532 ( .B1(P1_STATEBS16_REG_SCAN_IN), .B2(n15506), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n10712) );
  AOI21_X1 U13533 ( .B1(n11061), .B2(P1_EAX_REG_21__SCAN_IN), .A(n10712), .ZN(
        n10713) );
  OAI21_X1 U13534 ( .B1(n11057), .B2(n10714), .A(n10713), .ZN(n10716) );
  XNOR2_X1 U13535 ( .A(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .B(n10717), .ZN(
        n15497) );
  NAND2_X1 U13536 ( .A1(n11054), .A2(n15497), .ZN(n10715) );
  OR2_X1 U13537 ( .A1(n10718), .A2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n10719) );
  NAND2_X1 U13538 ( .A1(n10719), .A2(n10763), .ZN(n15590) );
  AOI22_X1 U13539 ( .A1(n9624), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n10484), .B2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n10723) );
  AOI22_X1 U13540 ( .A1(n10682), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n10171), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n10722) );
  AOI22_X1 U13541 ( .A1(n10387), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n11041), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n10721) );
  AOI22_X1 U13542 ( .A1(n9620), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n11042), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10720) );
  NAND4_X1 U13543 ( .A1(n10723), .A2(n10722), .A3(n10721), .A4(n10720), .ZN(
        n10729) );
  AOI22_X1 U13544 ( .A1(n10768), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n10485), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n10727) );
  AOI22_X1 U13545 ( .A1(n10734), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n10504), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n10726) );
  AOI22_X1 U13546 ( .A1(n10998), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n9628), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n10725) );
  AOI22_X1 U13547 ( .A1(n9619), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n10213), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n10724) );
  NAND4_X1 U13548 ( .A1(n10727), .A2(n10726), .A3(n10725), .A4(n10724), .ZN(
        n10728) );
  NOR2_X1 U13549 ( .A1(n10729), .A2(n10728), .ZN(n10732) );
  OAI21_X1 U13550 ( .B1(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n20891), .A(
        n20599), .ZN(n10731) );
  NAND2_X1 U13551 ( .A1(n11061), .A2(P1_EAX_REG_22__SCAN_IN), .ZN(n10730) );
  OAI211_X1 U13552 ( .C1(n11057), .C2(n10732), .A(n10731), .B(n10730), .ZN(
        n10733) );
  OAI21_X1 U13553 ( .B1(n15590), .B2(n10404), .A(n10733), .ZN(n14243) );
  AOI22_X1 U13554 ( .A1(n9625), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n10734), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n10738) );
  AOI22_X1 U13555 ( .A1(n10504), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n10682), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n10737) );
  AOI22_X1 U13556 ( .A1(n10768), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n11035), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n10736) );
  AOI22_X1 U13557 ( .A1(n10484), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n10213), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n10735) );
  NAND4_X1 U13558 ( .A1(n10738), .A2(n10737), .A3(n10736), .A4(n10735), .ZN(
        n10744) );
  AOI22_X1 U13559 ( .A1(n10387), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n9616), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n10742) );
  AOI22_X1 U13560 ( .A1(n10972), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n9638), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n10741) );
  AOI22_X1 U13561 ( .A1(n11036), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n11041), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n10740) );
  AOI22_X1 U13562 ( .A1(n9620), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n10208), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n10739) );
  NAND4_X1 U13563 ( .A1(n10742), .A2(n10741), .A3(n10740), .A4(n10739), .ZN(
        n10743) );
  NOR2_X1 U13564 ( .A1(n10744), .A2(n10743), .ZN(n10766) );
  AOI22_X1 U13565 ( .A1(n10387), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n10187), .B2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n10748) );
  AOI22_X1 U13566 ( .A1(n10734), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n10485), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n10747) );
  AOI22_X1 U13567 ( .A1(n10768), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n9621), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n10746) );
  AOI22_X1 U13568 ( .A1(n10972), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n9628), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n10745) );
  NAND4_X1 U13569 ( .A1(n10748), .A2(n10747), .A3(n10746), .A4(n10745), .ZN(
        n10754) );
  AOI22_X1 U13570 ( .A1(n10504), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n10682), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n10752) );
  AOI22_X1 U13571 ( .A1(n9625), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n11041), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n10751) );
  AOI22_X1 U13572 ( .A1(n11035), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n10208), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n10750) );
  AOI22_X1 U13573 ( .A1(n9618), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n10213), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n10749) );
  NAND4_X1 U13574 ( .A1(n10752), .A2(n10751), .A3(n10750), .A4(n10749), .ZN(
        n10753) );
  NOR2_X1 U13575 ( .A1(n10754), .A2(n10753), .ZN(n10767) );
  XOR2_X1 U13576 ( .A(n10766), .B(n10767), .Z(n10755) );
  NAND2_X1 U13577 ( .A1(n10755), .A2(n11030), .ZN(n10759) );
  INV_X1 U13578 ( .A(P1_EAX_REG_23__SCAN_IN), .ZN(n14397) );
  NAND2_X1 U13579 ( .A1(n20599), .A2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n10756) );
  OAI211_X1 U13580 ( .C1(n11008), .C2(n14397), .A(n10404), .B(n10756), .ZN(
        n10757) );
  INV_X1 U13581 ( .A(n10757), .ZN(n10758) );
  NAND2_X1 U13582 ( .A1(n10759), .A2(n10758), .ZN(n10761) );
  XNOR2_X1 U13583 ( .A(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .B(n10763), .ZN(
        n15487) );
  NAND2_X1 U13584 ( .A1(n11054), .A2(n15487), .ZN(n10760) );
  NAND2_X1 U13585 ( .A1(n10761), .A2(n10760), .ZN(n14339) );
  INV_X1 U13586 ( .A(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n15496) );
  OR2_X1 U13587 ( .A1(n10764), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n10765) );
  NAND2_X1 U13588 ( .A1(n10765), .A2(n10803), .ZN(n15583) );
  NOR2_X1 U13589 ( .A1(n10767), .A2(n10766), .ZN(n10785) );
  AOI22_X1 U13590 ( .A1(n9624), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n10504), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n10772) );
  AOI22_X1 U13591 ( .A1(n11036), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n10682), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n10771) );
  AOI22_X1 U13592 ( .A1(n10768), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n9620), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n10770) );
  AOI22_X1 U13593 ( .A1(n11035), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n10208), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n10769) );
  NAND4_X1 U13594 ( .A1(n10772), .A2(n10771), .A3(n10770), .A4(n10769), .ZN(
        n10778) );
  AOI22_X1 U13595 ( .A1(n10734), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n10187), .B2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n10776) );
  AOI22_X1 U13596 ( .A1(n10387), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n11041), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n10775) );
  AOI22_X1 U13597 ( .A1(n10972), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n9638), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n10774) );
  AOI22_X1 U13598 ( .A1(n9618), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n10213), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10773) );
  NAND4_X1 U13599 ( .A1(n10776), .A2(n10775), .A3(n10774), .A4(n10773), .ZN(
        n10777) );
  OR2_X1 U13600 ( .A1(n10778), .A2(n10777), .ZN(n10784) );
  XNOR2_X1 U13601 ( .A(n10785), .B(n10784), .ZN(n10781) );
  OAI21_X1 U13602 ( .B1(n20891), .B2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .A(
        n20599), .ZN(n10780) );
  NAND2_X1 U13603 ( .A1(n11061), .A2(P1_EAX_REG_24__SCAN_IN), .ZN(n10779) );
  OAI211_X1 U13604 ( .C1(n10781), .C2(n11057), .A(n10780), .B(n10779), .ZN(
        n10782) );
  OAI21_X1 U13605 ( .B1(n15583), .B2(n10404), .A(n10782), .ZN(n10783) );
  INV_X1 U13606 ( .A(n10783), .ZN(n14327) );
  NAND2_X1 U13607 ( .A1(n10785), .A2(n10784), .ZN(n10806) );
  AOI22_X1 U13608 ( .A1(n11036), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n10504), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n10789) );
  AOI22_X1 U13609 ( .A1(n10768), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n10682), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n10788) );
  AOI22_X1 U13610 ( .A1(n10972), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n9638), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n10787) );
  AOI22_X1 U13611 ( .A1(n9618), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n10213), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n10786) );
  NAND4_X1 U13612 ( .A1(n10789), .A2(n10788), .A3(n10787), .A4(n10786), .ZN(
        n10795) );
  AOI22_X1 U13613 ( .A1(n10734), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n10187), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n10793) );
  AOI22_X1 U13614 ( .A1(n9625), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n11035), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n10792) );
  AOI22_X1 U13615 ( .A1(n10387), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n11041), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n10791) );
  AOI22_X1 U13616 ( .A1(n9621), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n11042), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n10790) );
  NAND4_X1 U13617 ( .A1(n10793), .A2(n10792), .A3(n10791), .A4(n10790), .ZN(
        n10794) );
  NOR2_X1 U13618 ( .A1(n10795), .A2(n10794), .ZN(n10807) );
  XOR2_X1 U13619 ( .A(n10806), .B(n10807), .Z(n10796) );
  NAND2_X1 U13620 ( .A1(n10796), .A2(n11030), .ZN(n10801) );
  INV_X1 U13621 ( .A(P1_EAX_REG_25__SCAN_IN), .ZN(n14387) );
  NAND2_X1 U13622 ( .A1(n20599), .A2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n10797) );
  OAI211_X1 U13623 ( .C1(n11008), .C2(n14387), .A(n10404), .B(n10797), .ZN(
        n10798) );
  INV_X1 U13624 ( .A(n10798), .ZN(n10800) );
  XNOR2_X1 U13625 ( .A(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .B(n10803), .ZN(
        n15470) );
  INV_X1 U13626 ( .A(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n10802) );
  OR2_X1 U13627 ( .A1(n10804), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n10805) );
  NAND2_X1 U13628 ( .A1(n10805), .A2(n11011), .ZN(n15575) );
  NOR2_X1 U13629 ( .A1(n10807), .A2(n10806), .ZN(n10971) );
  AOI22_X1 U13630 ( .A1(n9624), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n10504), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n10811) );
  AOI22_X1 U13631 ( .A1(n11036), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n10682), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n10810) );
  AOI22_X1 U13632 ( .A1(n10768), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n9620), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10809) );
  AOI22_X1 U13633 ( .A1(n11035), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n11042), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n10808) );
  NAND4_X1 U13634 ( .A1(n10811), .A2(n10810), .A3(n10809), .A4(n10808), .ZN(
        n10817) );
  AOI22_X1 U13635 ( .A1(n10734), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n10187), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n10815) );
  AOI22_X1 U13636 ( .A1(n10387), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n11041), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n10814) );
  AOI22_X1 U13637 ( .A1(n10972), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n9628), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n10813) );
  AOI22_X1 U13638 ( .A1(n9619), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n10213), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10812) );
  NAND4_X1 U13639 ( .A1(n10815), .A2(n10814), .A3(n10813), .A4(n10812), .ZN(
        n10816) );
  OR2_X1 U13640 ( .A1(n10817), .A2(n10816), .ZN(n10970) );
  XNOR2_X1 U13641 ( .A(n10971), .B(n10970), .ZN(n10818) );
  NOR2_X1 U13642 ( .A1(n10818), .A2(n11057), .ZN(n10821) );
  INV_X1 U13643 ( .A(P1_EAX_REG_26__SCAN_IN), .ZN(n14382) );
  NAND2_X1 U13644 ( .A1(n20599), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n10819) );
  OAI211_X1 U13645 ( .C1(n11008), .C2(n14382), .A(n10404), .B(n10819), .ZN(
        n10820) );
  OAI22_X1 U13646 ( .A1(n15575), .A2(n10404), .B1(n10821), .B2(n10820), .ZN(
        n10823) );
  NAND2_X1 U13647 ( .A1(n10822), .A2(n10823), .ZN(n10824) );
  XNOR2_X1 U13648 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n10847) );
  NAND2_X1 U13649 ( .A1(n10848), .A2(n10847), .ZN(n10846) );
  NAND2_X1 U13650 ( .A1(n20697), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10825) );
  NAND2_X1 U13651 ( .A1(n10846), .A2(n10825), .ZN(n10836) );
  NAND2_X1 U13652 ( .A1(n20326), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10827) );
  NAND2_X1 U13653 ( .A1(n13329), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n10826) );
  NAND2_X1 U13654 ( .A1(n10836), .A2(n10835), .ZN(n10834) );
  NAND2_X1 U13655 ( .A1(n10834), .A2(n10827), .ZN(n10829) );
  MUX2_X1 U13656 ( .A(n20690), .B(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .S(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n10828) );
  AOI222_X1 U13657 ( .A1(n10859), .A2(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), 
        .B1(n10859), .B2(n15861), .C1(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), 
        .C2(n15861), .ZN(n11072) );
  NOR2_X1 U13658 ( .A1(n10829), .A2(n10828), .ZN(n10830) );
  INV_X1 U13659 ( .A(n11068), .ZN(n10857) );
  NAND2_X1 U13660 ( .A1(n20096), .A2(n14367), .ZN(n10833) );
  OAI21_X1 U13661 ( .B1(n10836), .B2(n10835), .A(n10834), .ZN(n11069) );
  NAND2_X1 U13662 ( .A1(n10862), .A2(n11069), .ZN(n10838) );
  NOR3_X1 U13663 ( .A1(n10839), .A2(n10248), .A3(n20086), .ZN(n10842) );
  AND2_X1 U13664 ( .A1(n9779), .A2(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n10840) );
  NOR2_X1 U13665 ( .A1(n10848), .A2(n10840), .ZN(n10843) );
  INV_X1 U13666 ( .A(n10843), .ZN(n10841) );
  NOR2_X1 U13667 ( .A1(n10842), .A2(n10841), .ZN(n10845) );
  AOI21_X1 U13668 ( .B1(n10866), .B2(n10843), .A(n10867), .ZN(n10844) );
  AOI21_X1 U13669 ( .B1(n10845), .B2(n10855), .A(n10844), .ZN(n10854) );
  OAI21_X1 U13670 ( .B1(n10848), .B2(n10847), .A(n10846), .ZN(n11070) );
  INV_X1 U13671 ( .A(n11070), .ZN(n10851) );
  OAI21_X1 U13672 ( .B1(n10849), .B2(n20096), .A(n14367), .ZN(n10850) );
  NAND2_X1 U13673 ( .A1(n10850), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n10852) );
  OAI21_X1 U13674 ( .B1(n10851), .B2(n10858), .A(n10852), .ZN(n10853) );
  NAND2_X1 U13675 ( .A1(n10852), .A2(n10256), .ZN(n10861) );
  AND2_X1 U13676 ( .A1(n15861), .A2(n10859), .ZN(n10860) );
  NAND2_X1 U13677 ( .A1(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n10860), .ZN(
        n11071) );
  NAND2_X1 U13678 ( .A1(n14177), .A2(n10256), .ZN(n13160) );
  OR2_X1 U13679 ( .A1(n15362), .A2(n20597), .ZN(n19820) );
  INV_X1 U13680 ( .A(n19820), .ZN(n19826) );
  OR2_X1 U13681 ( .A1(n11116), .A2(n20086), .ZN(n10953) );
  INV_X2 U13682 ( .A(n10878), .ZN(n14200) );
  INV_X1 U13683 ( .A(n11066), .ZN(n11111) );
  OAI22_X1 U13684 ( .A1(n13145), .A2(n11111), .B1(n10198), .B2(n14298), .ZN(
        n13161) );
  INV_X1 U13685 ( .A(n13161), .ZN(n13183) );
  NAND3_X1 U13686 ( .A1(n13382), .A2(n19826), .A3(n13183), .ZN(n10872) );
  INV_X1 U13687 ( .A(n13489), .ZN(n20117) );
  NAND4_X1 U13688 ( .A1(n20107), .A2(n20117), .A3(n19826), .A4(n10869), .ZN(
        n11077) );
  NOR2_X1 U13689 ( .A1(n11077), .A2(n10881), .ZN(n10870) );
  NAND2_X1 U13690 ( .A1(n10115), .A2(n10870), .ZN(n10871) );
  INV_X1 U13691 ( .A(P1_EBX_REG_1__SCAN_IN), .ZN(n10873) );
  INV_X1 U13692 ( .A(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n10874) );
  NAND2_X1 U13693 ( .A1(n10953), .A2(n10874), .ZN(n10875) );
  OAI211_X1 U13694 ( .C1(n10881), .C2(P1_EBX_REG_1__SCAN_IN), .A(n10875), .B(
        n14200), .ZN(n10876) );
  NAND2_X1 U13695 ( .A1(n10877), .A2(n10876), .ZN(n10882) );
  NAND2_X1 U13696 ( .A1(n10953), .A2(P1_EBX_REG_0__SCAN_IN), .ZN(n10880) );
  INV_X1 U13697 ( .A(P1_EBX_REG_0__SCAN_IN), .ZN(n13151) );
  NAND2_X1 U13698 ( .A1(n14200), .A2(n13151), .ZN(n10879) );
  NAND2_X1 U13699 ( .A1(n10880), .A2(n10879), .ZN(n13146) );
  XNOR2_X1 U13700 ( .A(n10882), .B(n13146), .ZN(n13129) );
  INV_X1 U13701 ( .A(n10881), .ZN(n13128) );
  NAND2_X1 U13702 ( .A1(n13129), .A2(n13128), .ZN(n13131) );
  INV_X1 U13703 ( .A(P1_EBX_REG_2__SCAN_IN), .ZN(n10883) );
  NAND2_X1 U13704 ( .A1(n14200), .A2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n10884) );
  NAND2_X1 U13705 ( .A1(n10953), .A2(n10884), .ZN(n10885) );
  OAI21_X1 U13706 ( .B1(n10881), .B2(P1_EBX_REG_2__SCAN_IN), .A(n10885), .ZN(
        n10886) );
  AND2_X1 U13707 ( .A1(n10887), .A2(n10886), .ZN(n13143) );
  MUX2_X1 U13708 ( .A(n12890), .B(n14200), .S(P1_EBX_REG_3__SCAN_IN), .Z(
        n10889) );
  INV_X1 U13709 ( .A(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n13409) );
  NAND2_X1 U13710 ( .A1(n13145), .A2(n13409), .ZN(n10888) );
  NAND2_X1 U13711 ( .A1(n10889), .A2(n10888), .ZN(n13333) );
  MUX2_X1 U13712 ( .A(n12890), .B(n14200), .S(P1_EBX_REG_5__SCAN_IN), .Z(
        n10890) );
  NAND2_X1 U13713 ( .A1(n10890), .A2(n10118), .ZN(n13452) );
  INV_X1 U13714 ( .A(n13452), .ZN(n10895) );
  NAND2_X1 U13715 ( .A1(n14200), .A2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n10891) );
  NAND2_X1 U13716 ( .A1(n10953), .A2(n10891), .ZN(n10892) );
  OAI21_X1 U13717 ( .B1(n10881), .B2(P1_EBX_REG_4__SCAN_IN), .A(n10892), .ZN(
        n10893) );
  NAND2_X1 U13718 ( .A1(n10894), .A2(n10893), .ZN(n13451) );
  NAND2_X1 U13719 ( .A1(n10895), .A2(n13451), .ZN(n10896) );
  MUX2_X1 U13720 ( .A(n12890), .B(n14200), .S(P1_EBX_REG_7__SCAN_IN), .Z(
        n10897) );
  NAND2_X1 U13721 ( .A1(n10897), .A2(n10122), .ZN(n13583) );
  INV_X1 U13722 ( .A(P1_EBX_REG_6__SCAN_IN), .ZN(n19944) );
  INV_X1 U13723 ( .A(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n15835) );
  NAND2_X1 U13724 ( .A1(n10953), .A2(n15835), .ZN(n10898) );
  OAI211_X1 U13725 ( .C1(n10881), .C2(P1_EBX_REG_6__SCAN_IN), .A(n10898), .B(
        n14200), .ZN(n10899) );
  NOR2_X1 U13726 ( .A1(n13583), .A2(n15849), .ZN(n10901) );
  INV_X1 U13727 ( .A(P1_EBX_REG_8__SCAN_IN), .ZN(n10902) );
  INV_X1 U13728 ( .A(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n15841) );
  NAND2_X1 U13729 ( .A1(n10953), .A2(n15841), .ZN(n10903) );
  OAI211_X1 U13730 ( .C1(n10881), .C2(P1_EBX_REG_8__SCAN_IN), .A(n10903), .B(
        n14200), .ZN(n10904) );
  NAND2_X1 U13731 ( .A1(n10905), .A2(n10904), .ZN(n13658) );
  MUX2_X1 U13732 ( .A(n12890), .B(n14200), .S(P1_EBX_REG_9__SCAN_IN), .Z(
        n10906) );
  NAND2_X1 U13733 ( .A1(n10906), .A2(n10123), .ZN(n13772) );
  INV_X1 U13734 ( .A(P1_EBX_REG_10__SCAN_IN), .ZN(n13791) );
  INV_X1 U13735 ( .A(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n11184) );
  NAND2_X1 U13736 ( .A1(n10953), .A2(n11184), .ZN(n10907) );
  OAI211_X1 U13737 ( .C1(n10881), .C2(P1_EBX_REG_10__SCAN_IN), .A(n10907), .B(
        n14200), .ZN(n10908) );
  INV_X1 U13738 ( .A(n12890), .ZN(n10935) );
  INV_X1 U13739 ( .A(P1_EBX_REG_11__SCAN_IN), .ZN(n15557) );
  NAND2_X1 U13740 ( .A1(n10935), .A2(n15557), .ZN(n10912) );
  NAND2_X1 U13741 ( .A1(n14200), .A2(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n10910) );
  OAI211_X1 U13742 ( .C1(n10881), .C2(P1_EBX_REG_11__SCAN_IN), .A(n10953), .B(
        n10910), .ZN(n10911) );
  AND2_X1 U13743 ( .A1(n10912), .A2(n10911), .ZN(n15543) );
  INV_X1 U13744 ( .A(P1_EBX_REG_12__SCAN_IN), .ZN(n15534) );
  INV_X1 U13745 ( .A(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n15803) );
  NAND2_X1 U13746 ( .A1(n10953), .A2(n15803), .ZN(n10913) );
  OAI211_X1 U13747 ( .C1(n10881), .C2(P1_EBX_REG_12__SCAN_IN), .A(n10913), .B(
        n14200), .ZN(n10914) );
  NAND2_X1 U13748 ( .A1(n10915), .A2(n10914), .ZN(n14097) );
  MUX2_X1 U13749 ( .A(n12890), .B(n14200), .S(P1_EBX_REG_13__SCAN_IN), .Z(
        n10916) );
  NAND2_X1 U13750 ( .A1(n10916), .A2(n10124), .ZN(n14131) );
  INV_X1 U13751 ( .A(P1_EBX_REG_15__SCAN_IN), .ZN(n14288) );
  NAND2_X1 U13752 ( .A1(n10935), .A2(n14288), .ZN(n10919) );
  NAND2_X1 U13753 ( .A1(n14200), .A2(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n10917) );
  OAI211_X1 U13754 ( .C1(n10881), .C2(P1_EBX_REG_15__SCAN_IN), .A(n10953), .B(
        n10917), .ZN(n10918) );
  AND2_X1 U13755 ( .A1(n10919), .A2(n10918), .ZN(n14117) );
  INV_X1 U13756 ( .A(P1_EBX_REG_14__SCAN_IN), .ZN(n14106) );
  INV_X1 U13757 ( .A(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n15778) );
  NAND2_X1 U13758 ( .A1(n10953), .A2(n15778), .ZN(n10920) );
  OAI211_X1 U13759 ( .C1(n10881), .C2(P1_EBX_REG_14__SCAN_IN), .A(n10920), .B(
        n14200), .ZN(n10921) );
  NAND2_X1 U13760 ( .A1(n10922), .A2(n10921), .ZN(n14118) );
  NAND2_X1 U13761 ( .A1(n14117), .A2(n14118), .ZN(n10923) );
  INV_X1 U13762 ( .A(P1_EBX_REG_16__SCAN_IN), .ZN(n15555) );
  INV_X1 U13763 ( .A(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n11180) );
  NAND2_X1 U13764 ( .A1(n10953), .A2(n11180), .ZN(n10924) );
  OAI211_X1 U13765 ( .C1(n10881), .C2(P1_EBX_REG_16__SCAN_IN), .A(n10924), .B(
        n14200), .ZN(n10925) );
  AND2_X1 U13766 ( .A1(n10926), .A2(n10925), .ZN(n15530) );
  INV_X1 U13767 ( .A(P1_EBX_REG_17__SCAN_IN), .ZN(n20870) );
  NAND2_X1 U13768 ( .A1(n10935), .A2(n20870), .ZN(n10929) );
  NAND2_X1 U13769 ( .A1(n14200), .A2(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n10927) );
  OAI211_X1 U13770 ( .C1(n10881), .C2(P1_EBX_REG_17__SCAN_IN), .A(n10953), .B(
        n10927), .ZN(n10928) );
  NAND2_X1 U13771 ( .A1(n10929), .A2(n10928), .ZN(n14274) );
  NOR2_X1 U13772 ( .A1(n15530), .A2(n14274), .ZN(n10930) );
  INV_X1 U13773 ( .A(P1_EBX_REG_18__SCAN_IN), .ZN(n10931) );
  INV_X1 U13774 ( .A(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n15749) );
  NAND2_X1 U13775 ( .A1(n10953), .A2(n15749), .ZN(n10932) );
  OAI211_X1 U13776 ( .C1(n10881), .C2(P1_EBX_REG_18__SCAN_IN), .A(n10932), .B(
        n14200), .ZN(n10933) );
  AND2_X1 U13777 ( .A1(n10934), .A2(n10933), .ZN(n14362) );
  INV_X1 U13778 ( .A(P1_EBX_REG_19__SCAN_IN), .ZN(n14355) );
  NAND2_X1 U13779 ( .A1(n10935), .A2(n14355), .ZN(n10938) );
  NAND2_X1 U13780 ( .A1(n14200), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n10936) );
  OAI211_X1 U13781 ( .C1(n10881), .C2(P1_EBX_REG_19__SCAN_IN), .A(n10953), .B(
        n10936), .ZN(n10937) );
  NAND2_X1 U13782 ( .A1(n10938), .A2(n10937), .ZN(n14257) );
  NOR2_X1 U13783 ( .A1(n14362), .A2(n14257), .ZN(n10939) );
  MUX2_X1 U13784 ( .A(n12890), .B(n14200), .S(P1_EBX_REG_21__SCAN_IN), .Z(
        n10940) );
  NAND2_X1 U13785 ( .A1(n10940), .A2(n10111), .ZN(n14344) );
  INV_X1 U13786 ( .A(n14344), .ZN(n10945) );
  INV_X1 U13787 ( .A(P1_EBX_REG_20__SCAN_IN), .ZN(n10941) );
  INV_X1 U13788 ( .A(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n15419) );
  NAND2_X1 U13789 ( .A1(n10953), .A2(n15419), .ZN(n10942) );
  OAI211_X1 U13790 ( .C1(n10881), .C2(P1_EBX_REG_20__SCAN_IN), .A(n10942), .B(
        n14200), .ZN(n10943) );
  NAND2_X1 U13791 ( .A1(n10944), .A2(n10943), .ZN(n14352) );
  NAND2_X1 U13792 ( .A1(n10945), .A2(n14352), .ZN(n10946) );
  INV_X1 U13793 ( .A(P1_EBX_REG_22__SCAN_IN), .ZN(n14343) );
  NAND2_X1 U13794 ( .A1(n14200), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n10947) );
  NAND2_X1 U13795 ( .A1(n10953), .A2(n10947), .ZN(n10948) );
  OAI21_X1 U13796 ( .B1(n10881), .B2(P1_EBX_REG_22__SCAN_IN), .A(n10948), .ZN(
        n10949) );
  AND2_X1 U13797 ( .A1(n10950), .A2(n10949), .ZN(n14238) );
  MUX2_X1 U13798 ( .A(n12890), .B(n14200), .S(P1_EBX_REG_23__SCAN_IN), .Z(
        n10952) );
  INV_X1 U13799 ( .A(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n15717) );
  NAND2_X1 U13800 ( .A1(n13145), .A2(n15717), .ZN(n10951) );
  AND2_X1 U13801 ( .A1(n10952), .A2(n10951), .ZN(n14335) );
  INV_X1 U13802 ( .A(P1_EBX_REG_24__SCAN_IN), .ZN(n14332) );
  INV_X1 U13803 ( .A(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n15577) );
  NAND2_X1 U13804 ( .A1(n10953), .A2(n15577), .ZN(n10954) );
  OAI211_X1 U13805 ( .C1(n10881), .C2(P1_EBX_REG_24__SCAN_IN), .A(n10954), .B(
        n14200), .ZN(n10955) );
  NAND2_X1 U13806 ( .A1(n10956), .A2(n10955), .ZN(n14329) );
  MUX2_X1 U13807 ( .A(n12890), .B(n14200), .S(P1_EBX_REG_25__SCAN_IN), .Z(
        n10957) );
  NAND2_X1 U13808 ( .A1(n10957), .A2(n10112), .ZN(n14320) );
  INV_X1 U13809 ( .A(P1_EBX_REG_26__SCAN_IN), .ZN(n10964) );
  NAND2_X1 U13810 ( .A1(n14200), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n10958) );
  NAND2_X1 U13811 ( .A1(n10953), .A2(n10958), .ZN(n10959) );
  OAI21_X1 U13812 ( .B1(n10881), .B2(P1_EBX_REG_26__SCAN_IN), .A(n10959), .ZN(
        n10960) );
  AND2_X1 U13813 ( .A1(n10961), .A2(n10960), .ZN(n10962) );
  NAND2_X1 U13815 ( .A1(n14322), .A2(n10962), .ZN(n10963) );
  NAND2_X1 U13816 ( .A1(n14225), .A2(n10963), .ZN(n15694) );
  OR2_X1 U13817 ( .A1(n15694), .A2(n14356), .ZN(n10967) );
  NAND2_X1 U13818 ( .A1(n10965), .A2(P1_EBX_REG_26__SCAN_IN), .ZN(n10966) );
  NAND2_X1 U13819 ( .A1(n10971), .A2(n10970), .ZN(n10992) );
  AOI22_X1 U13820 ( .A1(n9618), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n10972), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n10976) );
  AOI22_X1 U13821 ( .A1(n10734), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n10504), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n10975) );
  AOI22_X1 U13822 ( .A1(n11036), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n10682), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n10974) );
  AOI22_X1 U13823 ( .A1(n11035), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n9622), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n10973) );
  NAND4_X1 U13824 ( .A1(n10976), .A2(n10975), .A3(n10974), .A4(n10973), .ZN(
        n10982) );
  AOI22_X1 U13825 ( .A1(n9625), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n10187), .B2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n10980) );
  AOI22_X1 U13826 ( .A1(n10387), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n11041), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n10979) );
  AOI22_X1 U13827 ( .A1(n10768), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n11042), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n10978) );
  AOI22_X1 U13828 ( .A1(n9638), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n10213), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n10977) );
  NAND4_X1 U13829 ( .A1(n10980), .A2(n10979), .A3(n10978), .A4(n10977), .ZN(
        n10981) );
  NOR2_X1 U13830 ( .A1(n10982), .A2(n10981), .ZN(n10993) );
  XOR2_X1 U13831 ( .A(n10992), .B(n10993), .Z(n10983) );
  NAND2_X1 U13832 ( .A1(n10983), .A2(n11030), .ZN(n10987) );
  INV_X1 U13833 ( .A(P1_EAX_REG_27__SCAN_IN), .ZN(n14377) );
  OAI21_X1 U13834 ( .B1(n20891), .B2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .A(
        n20599), .ZN(n10984) );
  OAI21_X1 U13835 ( .B1(n11008), .B2(n14377), .A(n10984), .ZN(n10985) );
  INV_X1 U13836 ( .A(n10985), .ZN(n10986) );
  NAND2_X1 U13837 ( .A1(n10987), .A2(n10986), .ZN(n10989) );
  XNOR2_X1 U13838 ( .A(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .B(n11011), .ZN(
        n14231) );
  NAND2_X1 U13839 ( .A1(n11054), .A2(n14231), .ZN(n10988) );
  NAND2_X1 U13840 ( .A1(n10989), .A2(n10988), .ZN(n14223) );
  NOR2_X1 U13841 ( .A1(n10993), .A2(n10992), .ZN(n11016) );
  AOI22_X1 U13842 ( .A1(P1_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n9625), .B1(
        n10504), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n10997) );
  AOI22_X1 U13843 ( .A1(P1_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n11036), .B1(
        n10682), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n10996) );
  AOI22_X1 U13844 ( .A1(n10768), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n9621), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10995) );
  AOI22_X1 U13845 ( .A1(P1_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n10171), .B1(
        n11042), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n10994) );
  NAND4_X1 U13846 ( .A1(n10997), .A2(n10996), .A3(n10995), .A4(n10994), .ZN(
        n11004) );
  AOI22_X1 U13847 ( .A1(n10734), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n10187), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11002) );
  AOI22_X1 U13848 ( .A1(n10387), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n11041), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11001) );
  AOI22_X1 U13849 ( .A1(P1_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n10998), .B1(
        n9628), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11000) );
  AOI22_X1 U13850 ( .A1(n11021), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n10213), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10999) );
  NAND4_X1 U13851 ( .A1(n11002), .A2(n11001), .A3(n11000), .A4(n10999), .ZN(
        n11003) );
  OR2_X1 U13852 ( .A1(n11004), .A2(n11003), .ZN(n11015) );
  INV_X1 U13853 ( .A(n11015), .ZN(n11005) );
  XNOR2_X1 U13854 ( .A(n11016), .B(n11005), .ZN(n11010) );
  INV_X1 U13855 ( .A(P1_EAX_REG_28__SCAN_IN), .ZN(n11007) );
  NAND2_X1 U13856 ( .A1(n20599), .A2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n11006) );
  OAI211_X1 U13857 ( .C1(n11008), .C2(n11007), .A(n10404), .B(n11006), .ZN(
        n11009) );
  AOI21_X1 U13858 ( .B1(n11010), .B2(n11030), .A(n11009), .ZN(n11014) );
  INV_X1 U13859 ( .A(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n14232) );
  NAND2_X1 U13860 ( .A1(n11012), .A2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n11033) );
  OAI21_X1 U13861 ( .B1(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n11012), .A(
        n11033), .ZN(n15566) );
  NOR2_X1 U13862 ( .A1(n15566), .A2(n10404), .ZN(n11013) );
  XNOR2_X1 U13863 ( .A(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .B(n11033), .ZN(
        n14215) );
  NAND2_X1 U13864 ( .A1(n11016), .A2(n11015), .ZN(n11050) );
  AOI22_X1 U13865 ( .A1(n9624), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n10484), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11020) );
  AOI22_X1 U13866 ( .A1(n11036), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n10504), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11019) );
  AOI22_X1 U13867 ( .A1(n10768), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n9622), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11018) );
  AOI22_X1 U13868 ( .A1(n10972), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n10213), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11017) );
  NAND4_X1 U13869 ( .A1(n11020), .A2(n11019), .A3(n11018), .A4(n11017), .ZN(
        n11027) );
  AOI22_X1 U13870 ( .A1(n10734), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n10682), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11025) );
  AOI22_X1 U13871 ( .A1(n9616), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n9628), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11024) );
  AOI22_X1 U13872 ( .A1(n10387), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n11041), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11023) );
  AOI22_X1 U13873 ( .A1(n11035), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n11042), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11022) );
  NAND4_X1 U13874 ( .A1(n11025), .A2(n11024), .A3(n11023), .A4(n11022), .ZN(
        n11026) );
  NOR2_X1 U13875 ( .A1(n11027), .A2(n11026), .ZN(n11051) );
  XOR2_X1 U13876 ( .A(n11050), .B(n11051), .Z(n11031) );
  INV_X1 U13877 ( .A(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n11206) );
  NAND2_X1 U13878 ( .A1(n11061), .A2(P1_EAX_REG_29__SCAN_IN), .ZN(n11028) );
  OAI211_X1 U13879 ( .C1(P1_STATE2_REG_2__SCAN_IN), .C2(n11206), .A(n11028), 
        .B(n10404), .ZN(n11029) );
  AOI21_X1 U13880 ( .B1(n11031), .B2(n11030), .A(n11029), .ZN(n11032) );
  AOI21_X1 U13881 ( .B1(n11054), .B2(n14215), .A(n11032), .ZN(n11099) );
  INV_X1 U13882 ( .A(n11033), .ZN(n11034) );
  NAND2_X1 U13883 ( .A1(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n11034), .ZN(
        n12886) );
  INV_X1 U13884 ( .A(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n14453) );
  XNOR2_X1 U13885 ( .A(n12886), .B(n14453), .ZN(n14451) );
  AOI22_X1 U13886 ( .A1(n9625), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n10504), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11040) );
  AOI22_X1 U13887 ( .A1(n11036), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n11035), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n11039) );
  AOI22_X1 U13888 ( .A1(n10768), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n9620), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11038) );
  AOI22_X1 U13889 ( .A1(n10972), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n9638), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n11037) );
  NAND4_X1 U13890 ( .A1(n11040), .A2(n11039), .A3(n11038), .A4(n11037), .ZN(
        n11049) );
  AOI22_X1 U13891 ( .A1(n10458), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n10484), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n11047) );
  AOI22_X1 U13892 ( .A1(n10387), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n11041), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11046) );
  AOI22_X1 U13893 ( .A1(n10682), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n11042), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11045) );
  AOI22_X1 U13894 ( .A1(n9617), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n10213), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11044) );
  NAND4_X1 U13895 ( .A1(n11047), .A2(n11046), .A3(n11045), .A4(n11044), .ZN(
        n11048) );
  NOR2_X1 U13896 ( .A1(n11049), .A2(n11048), .ZN(n11053) );
  NOR2_X1 U13897 ( .A1(n11051), .A2(n11050), .ZN(n11052) );
  XOR2_X1 U13898 ( .A(n11053), .B(n11052), .Z(n11058) );
  AOI21_X1 U13899 ( .B1(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n20599), .A(
        n11054), .ZN(n11056) );
  NAND2_X1 U13900 ( .A1(n11061), .A2(P1_EAX_REG_30__SCAN_IN), .ZN(n11055) );
  OAI211_X1 U13901 ( .C1(n11058), .C2(n11057), .A(n11056), .B(n11055), .ZN(
        n11059) );
  OAI21_X1 U13902 ( .B1(n10404), .B2(n14451), .A(n11059), .ZN(n14198) );
  AOI22_X1 U13903 ( .A1(n11061), .A2(P1_EAX_REG_31__SCAN_IN), .B1(n11060), 
        .B2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n11062) );
  AND2_X1 U13904 ( .A1(n11064), .A2(n19826), .ZN(n11065) );
  NAND2_X1 U13905 ( .A1(READY11_REG_SCAN_IN), .A2(READY1), .ZN(n20728) );
  NAND2_X1 U13906 ( .A1(n10256), .A2(n20728), .ZN(n11080) );
  AOI21_X1 U13907 ( .B1(n13165), .B2(n20086), .A(n11066), .ZN(n13198) );
  AND2_X1 U13908 ( .A1(n13198), .A2(n10249), .ZN(n13395) );
  NAND2_X1 U13909 ( .A1(n15409), .A2(n13395), .ZN(n11076) );
  INV_X1 U13910 ( .A(n11067), .ZN(n11074) );
  NOR3_X1 U13911 ( .A1(n11070), .A2(n11069), .A3(n11068), .ZN(n11073) );
  OAI21_X1 U13912 ( .B1(n11073), .B2(n11072), .A(n11071), .ZN(n15349) );
  AND2_X1 U13913 ( .A1(n20728), .A2(n15349), .ZN(n13387) );
  NAND2_X1 U13914 ( .A1(n11074), .A2(n13387), .ZN(n11075) );
  NAND2_X1 U13915 ( .A1(n11076), .A2(n11075), .ZN(n13204) );
  NAND2_X1 U13916 ( .A1(n13204), .A2(n19826), .ZN(n11079) );
  OR2_X1 U13917 ( .A1(n13184), .A2(n11077), .ZN(n11078) );
  OAI211_X4 U13918 ( .C1(n15404), .C2(n11080), .A(n11079), .B(n11078), .ZN(
        n14436) );
  NAND2_X1 U13919 ( .A1(n12918), .A2(n10110), .ZN(n11095) );
  NOR4_X1 U13920 ( .A1(P1_ADDRESS_REG_16__SCAN_IN), .A2(
        P1_ADDRESS_REG_14__SCAN_IN), .A3(P1_ADDRESS_REG_13__SCAN_IN), .A4(
        P1_ADDRESS_REG_12__SCAN_IN), .ZN(n11084) );
  NOR4_X1 U13921 ( .A1(P1_ADDRESS_REG_19__SCAN_IN), .A2(
        P1_ADDRESS_REG_18__SCAN_IN), .A3(P1_ADDRESS_REG_15__SCAN_IN), .A4(
        P1_ADDRESS_REG_17__SCAN_IN), .ZN(n11083) );
  NOR4_X1 U13922 ( .A1(P1_ADDRESS_REG_7__SCAN_IN), .A2(
        P1_ADDRESS_REG_6__SCAN_IN), .A3(P1_ADDRESS_REG_5__SCAN_IN), .A4(
        P1_ADDRESS_REG_4__SCAN_IN), .ZN(n11082) );
  NOR4_X1 U13923 ( .A1(P1_ADDRESS_REG_11__SCAN_IN), .A2(
        P1_ADDRESS_REG_8__SCAN_IN), .A3(P1_ADDRESS_REG_10__SCAN_IN), .A4(
        P1_ADDRESS_REG_9__SCAN_IN), .ZN(n11081) );
  NAND4_X1 U13924 ( .A1(n11084), .A2(n11083), .A3(n11082), .A4(n11081), .ZN(
        n11089) );
  NOR4_X1 U13925 ( .A1(P1_ADDRESS_REG_3__SCAN_IN), .A2(
        P1_ADDRESS_REG_2__SCAN_IN), .A3(P1_ADDRESS_REG_28__SCAN_IN), .A4(
        P1_ADDRESS_REG_1__SCAN_IN), .ZN(n11087) );
  NOR4_X1 U13926 ( .A1(P1_ADDRESS_REG_23__SCAN_IN), .A2(
        P1_ADDRESS_REG_22__SCAN_IN), .A3(P1_ADDRESS_REG_21__SCAN_IN), .A4(
        P1_ADDRESS_REG_20__SCAN_IN), .ZN(n11086) );
  NOR4_X1 U13927 ( .A1(P1_ADDRESS_REG_27__SCAN_IN), .A2(
        P1_ADDRESS_REG_26__SCAN_IN), .A3(P1_ADDRESS_REG_25__SCAN_IN), .A4(
        P1_ADDRESS_REG_24__SCAN_IN), .ZN(n11085) );
  INV_X1 U13928 ( .A(P1_ADDRESS_REG_0__SCAN_IN), .ZN(n20618) );
  NAND4_X1 U13929 ( .A1(n11087), .A2(n11086), .A3(n11085), .A4(n20618), .ZN(
        n11088) );
  OAI21_X1 U13930 ( .B1(n11089), .B2(n11088), .A(P1_ADDRESS_REG_29__SCAN_IN), 
        .ZN(n20083) );
  NOR2_X1 U13931 ( .A1(n13384), .A2(n20083), .ZN(n11090) );
  INV_X1 U13932 ( .A(BUF1_REG_31__SCAN_IN), .ZN(n16249) );
  NOR2_X1 U13933 ( .A1(n14437), .A2(n16249), .ZN(n11093) );
  NOR3_X4 U13934 ( .A1(n14421), .A2(n20085), .A3(n13384), .ZN(n14439) );
  AOI22_X1 U13935 ( .A1(n14439), .A2(DATAI_31_), .B1(P1_EAX_REG_31__SCAN_IN), 
        .B2(n14421), .ZN(n11091) );
  INV_X1 U13936 ( .A(n11091), .ZN(n11092) );
  NOR2_X1 U13937 ( .A1(n11093), .A2(n11092), .ZN(n11094) );
  NAND2_X1 U13938 ( .A1(n11095), .A2(n11094), .ZN(P1_U2873) );
  NAND3_X1 U13939 ( .A1(n20597), .A2(P1_STATE2_REG_1__SCAN_IN), .A3(
        P1_STATEBS16_REG_SCAN_IN), .ZN(n15864) );
  INV_X1 U13940 ( .A(n15864), .ZN(n11100) );
  NOR2_X2 U13941 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20700) );
  NAND2_X1 U13942 ( .A1(n11101), .A2(n11154), .ZN(n11102) );
  INV_X1 U13943 ( .A(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n11103) );
  NAND2_X1 U13944 ( .A1(n15640), .A2(n11103), .ZN(n14445) );
  NAND2_X1 U13945 ( .A1(n15569), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n12919) );
  NAND2_X1 U13946 ( .A1(n14445), .A2(n12919), .ZN(n11197) );
  INV_X1 U13947 ( .A(n20722), .ZN(n11171) );
  INV_X1 U13948 ( .A(n11130), .ZN(n11105) );
  NAND2_X1 U13949 ( .A1(n11104), .A2(n11117), .ZN(n11124) );
  AND2_X1 U13950 ( .A1(n11124), .A2(n11123), .ZN(n11131) );
  NOR2_X1 U13951 ( .A1(n11105), .A2(n11131), .ZN(n11138) );
  NAND2_X1 U13952 ( .A1(n11138), .A2(n11139), .ZN(n11148) );
  NOR2_X1 U13953 ( .A1(n11149), .A2(n11148), .ZN(n11160) );
  NAND2_X1 U13954 ( .A1(n11160), .A2(n11158), .ZN(n11168) );
  XNOR2_X1 U13955 ( .A(n11170), .B(n11168), .ZN(n11106) );
  NAND2_X1 U13956 ( .A1(n11171), .A2(n11106), .ZN(n11107) );
  OAI21_X1 U13957 ( .B1(n11108), .B2(n11141), .A(n11107), .ZN(n15649) );
  XNOR2_X1 U13958 ( .A(n11110), .B(n11109), .ZN(n11112) );
  OAI211_X1 U13959 ( .C1(n20722), .C2(n11112), .A(n11111), .B(n14367), .ZN(
        n11113) );
  INV_X1 U13960 ( .A(n11113), .ZN(n11114) );
  OAI21_X1 U13961 ( .B1(n11115), .B2(n20096), .A(n11114), .ZN(n11120) );
  NAND2_X1 U13962 ( .A1(n20086), .A2(n11116), .ZN(n11127) );
  OAI21_X1 U13963 ( .B1(n20722), .B2(n11117), .A(n11127), .ZN(n11118) );
  AOI21_X1 U13964 ( .B1(n20701), .B2(n11154), .A(n11118), .ZN(n20038) );
  INV_X1 U13965 ( .A(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n20072) );
  OR2_X1 U13966 ( .A1(n20038), .A2(n20072), .ZN(n11119) );
  XNOR2_X1 U13967 ( .A(n11120), .B(n11119), .ZN(n20030) );
  NAND2_X1 U13968 ( .A1(n20030), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n20029) );
  INV_X1 U13969 ( .A(n11119), .ZN(n20037) );
  NAND2_X1 U13970 ( .A1(n11120), .A2(n20037), .ZN(n11121) );
  NAND2_X1 U13971 ( .A1(n20029), .A2(n11121), .ZN(n11128) );
  INV_X1 U13972 ( .A(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n11122) );
  XNOR2_X1 U13973 ( .A(n11128), .B(n11122), .ZN(n13355) );
  NOR2_X1 U13974 ( .A1(n11124), .A2(n11123), .ZN(n11125) );
  OAI21_X1 U13975 ( .B1(n11131), .B2(n11125), .A(n11171), .ZN(n11126) );
  OAI211_X1 U13976 ( .C1(n13434), .C2(n11141), .A(n11127), .B(n11126), .ZN(
        n13354) );
  NAND2_X1 U13977 ( .A1(n11128), .A2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n11129) );
  OR2_X1 U13978 ( .A1(n20683), .A2(n11141), .ZN(n11134) );
  XNOR2_X1 U13979 ( .A(n11131), .B(n11130), .ZN(n11132) );
  NAND2_X1 U13980 ( .A1(n11132), .A2(n11171), .ZN(n11133) );
  NAND2_X1 U13981 ( .A1(n11134), .A2(n11133), .ZN(n13349) );
  NAND2_X1 U13982 ( .A1(n11135), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n11136) );
  NAND2_X1 U13983 ( .A1(n11137), .A2(n11136), .ZN(n13439) );
  XNOR2_X1 U13984 ( .A(n11139), .B(n11138), .ZN(n11140) );
  OAI22_X1 U13985 ( .A1(n11142), .A2(n11141), .B1(n11140), .B2(n20722), .ZN(
        n11144) );
  INV_X1 U13986 ( .A(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n11143) );
  XNOR2_X1 U13987 ( .A(n11144), .B(n11143), .ZN(n13438) );
  NAND2_X1 U13988 ( .A1(n13439), .A2(n13438), .ZN(n11146) );
  NAND2_X1 U13989 ( .A1(n11144), .A2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11145) );
  NAND2_X1 U13990 ( .A1(n11147), .A2(n11154), .ZN(n11152) );
  XOR2_X1 U13991 ( .A(n11149), .B(n11148), .Z(n11150) );
  NAND2_X1 U13992 ( .A1(n11150), .A2(n11171), .ZN(n11151) );
  NAND2_X1 U13993 ( .A1(n11152), .A2(n11151), .ZN(n11153) );
  INV_X1 U13994 ( .A(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n13498) );
  XNOR2_X1 U13995 ( .A(n11153), .B(n13498), .ZN(n13494) );
  NAND2_X1 U13996 ( .A1(n11155), .A2(n11154), .ZN(n11156) );
  OR2_X1 U13997 ( .A1(n11157), .A2(n11156), .ZN(n11163) );
  INV_X1 U13998 ( .A(n11158), .ZN(n11159) );
  XNOR2_X1 U13999 ( .A(n11160), .B(n11159), .ZN(n11161) );
  NAND2_X1 U14000 ( .A1(n11161), .A2(n11171), .ZN(n11162) );
  NAND2_X1 U14001 ( .A1(n11163), .A2(n11162), .ZN(n11165) );
  INV_X1 U14002 ( .A(n11165), .ZN(n11164) );
  NAND2_X1 U14003 ( .A1(n11164), .A2(n15835), .ZN(n15656) );
  NAND2_X1 U14004 ( .A1(n11165), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n15655) );
  NAND2_X1 U14005 ( .A1(n15649), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n11167) );
  INV_X1 U14006 ( .A(n11168), .ZN(n11169) );
  NAND3_X1 U14007 ( .A1(n11171), .A2(n11170), .A3(n11169), .ZN(n11172) );
  NAND2_X1 U14008 ( .A1(n11173), .A2(n11172), .ZN(n13753) );
  INV_X1 U14009 ( .A(n13753), .ZN(n11174) );
  NAND2_X1 U14010 ( .A1(n15640), .A2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n11175) );
  INV_X1 U14011 ( .A(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n15833) );
  NAND2_X1 U14012 ( .A1(n15620), .A2(n15833), .ZN(n11176) );
  NAND2_X1 U14013 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n11177) );
  NAND2_X1 U14014 ( .A1(n15620), .A2(n15778), .ZN(n11178) );
  NAND2_X1 U14015 ( .A1(n15621), .A2(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n14516) );
  INV_X1 U14016 ( .A(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n15793) );
  NAND2_X1 U14017 ( .A1(n15793), .A2(n15778), .ZN(n11179) );
  NAND2_X1 U14018 ( .A1(n15621), .A2(n11179), .ZN(n11186) );
  AND2_X1 U14019 ( .A1(n14516), .A2(n11186), .ZN(n14500) );
  MUX2_X1 U14020 ( .A(n11180), .B(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .S(
        n11173), .Z(n15609) );
  INV_X1 U14021 ( .A(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n11181) );
  NAND2_X1 U14022 ( .A1(n15620), .A2(n11181), .ZN(n14517) );
  NAND2_X1 U14023 ( .A1(n15609), .A2(n14517), .ZN(n15606) );
  AOI21_X1 U14024 ( .B1(n14515), .B2(n14500), .A(n15606), .ZN(n14501) );
  INV_X1 U14025 ( .A(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n14506) );
  NAND2_X1 U14026 ( .A1(n15620), .A2(n14506), .ZN(n11182) );
  NAND2_X1 U14027 ( .A1(n11184), .A2(n15795), .ZN(n11185) );
  NAND2_X1 U14028 ( .A1(n15621), .A2(n11185), .ZN(n14529) );
  NAND2_X1 U14029 ( .A1(n15640), .A2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n14531) );
  NAND2_X1 U14030 ( .A1(n15615), .A2(n11186), .ZN(n14513) );
  NOR2_X1 U14031 ( .A1(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n15757) );
  AND2_X1 U14032 ( .A1(n15757), .A2(n14506), .ZN(n11187) );
  NOR2_X1 U14033 ( .A1(n15620), .A2(n11187), .ZN(n11188) );
  NOR2_X1 U14034 ( .A1(n14513), .A2(n11188), .ZN(n11189) );
  AND2_X1 U14035 ( .A1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n15379) );
  AND2_X1 U14036 ( .A1(n15379), .A2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n14551) );
  INV_X1 U14037 ( .A(n14551), .ZN(n11190) );
  INV_X1 U14038 ( .A(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n15413) );
  NOR2_X1 U14039 ( .A1(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n11192) );
  NAND2_X1 U14040 ( .A1(n14476), .A2(n11192), .ZN(n14458) );
  INV_X1 U14041 ( .A(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n12892) );
  INV_X1 U14042 ( .A(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n11193) );
  NAND2_X1 U14043 ( .A1(n12892), .A2(n11193), .ZN(n11194) );
  INV_X1 U14044 ( .A(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n14471) );
  NAND2_X1 U14045 ( .A1(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n15688) );
  NOR2_X1 U14046 ( .A1(n14471), .A2(n15688), .ZN(n14552) );
  INV_X1 U14047 ( .A(n14552), .ZN(n15558) );
  NAND2_X1 U14048 ( .A1(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n15673) );
  NOR2_X1 U14049 ( .A1(n13490), .A2(n13410), .ZN(n11199) );
  OR2_X1 U14050 ( .A1(n11199), .A2(n11198), .ZN(n13196) );
  NOR2_X1 U14051 ( .A1(n13196), .A2(n10868), .ZN(n11200) );
  AND2_X1 U14052 ( .A1(n11200), .A2(n13198), .ZN(n13396) );
  NOR2_X1 U14053 ( .A1(n15666), .A2(n20031), .ZN(n11211) );
  OR2_X1 U14054 ( .A1(n11205), .A2(n20700), .ZN(n20727) );
  NAND2_X1 U14055 ( .A1(n20727), .A2(n20597), .ZN(n11201) );
  NAND2_X1 U14056 ( .A1(n20597), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n11203) );
  NAND2_X1 U14057 ( .A1(n20891), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n11202) );
  AND2_X1 U14058 ( .A1(n11203), .A2(n11202), .ZN(n20040) );
  INV_X1 U14059 ( .A(n20040), .ZN(n11204) );
  NAND2_X1 U14060 ( .A1(n15635), .A2(n14215), .ZN(n11209) );
  NAND2_X1 U14061 ( .A1(n11205), .A2(n20599), .ZN(n20050) );
  INV_X1 U14062 ( .A(P1_REIP_REG_29__SCAN_IN), .ZN(n14217) );
  OAI22_X1 U14063 ( .A1(n20039), .A2(n11206), .B1(n20050), .B2(n14217), .ZN(
        n11207) );
  INV_X1 U14064 ( .A(n11207), .ZN(n11208) );
  NAND2_X1 U14065 ( .A1(n11209), .A2(n11208), .ZN(n11210) );
  INV_X1 U14066 ( .A(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n16054) );
  INV_X1 U14067 ( .A(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n18834) );
  NAND2_X1 U14068 ( .A1(n11229), .A2(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n11227) );
  INV_X1 U14069 ( .A(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n11215) );
  INV_X1 U14070 ( .A(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n16026) );
  OR2_X1 U14071 ( .A1(n11215), .A2(n16026), .ZN(n11216) );
  INV_X1 U14072 ( .A(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n18789) );
  INV_X1 U14073 ( .A(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n20894) );
  INV_X1 U14074 ( .A(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n11243) );
  NAND2_X1 U14075 ( .A1(n11217), .A2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n11219) );
  OAI21_X1 U14076 ( .B1(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n11217), .A(
        n11219), .ZN(n11218) );
  INV_X1 U14077 ( .A(n11218), .ZN(n15985) );
  INV_X1 U14078 ( .A(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n15984) );
  NAND2_X1 U14079 ( .A1(n11246), .A2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n11247) );
  INV_X1 U14080 ( .A(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n15960) );
  NAND2_X1 U14081 ( .A1(n11248), .A2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n11249) );
  INV_X1 U14082 ( .A(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n15895) );
  INV_X1 U14083 ( .A(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n15888) );
  INV_X1 U14084 ( .A(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n14569) );
  NAND2_X1 U14085 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n12471) );
  AOI21_X1 U14086 ( .B1(n20894), .B2(n11222), .A(n9744), .ZN(n14769) );
  OR2_X1 U14087 ( .A1(n11224), .A2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n11221) );
  NAND2_X1 U14088 ( .A1(n11222), .A2(n11221), .ZN(n18765) );
  INV_X1 U14089 ( .A(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n18771) );
  INV_X1 U14090 ( .A(n11223), .ZN(n11225) );
  AOI21_X1 U14091 ( .B1(n18771), .B2(n11225), .A(n11224), .ZN(n15993) );
  INV_X1 U14092 ( .A(n15993), .ZN(n18781) );
  INV_X1 U14093 ( .A(n11226), .ZN(n11240) );
  AOI21_X1 U14094 ( .B1(n18789), .B2(n11240), .A(n11223), .ZN(n18787) );
  NOR2_X1 U14095 ( .A1(n16026), .A2(n11227), .ZN(n11241) );
  AOI21_X1 U14096 ( .B1(n16026), .B2(n11227), .A(n11241), .ZN(n18807) );
  AOI21_X1 U14097 ( .B1(n18834), .B2(n11228), .A(n11229), .ZN(n18832) );
  AOI21_X1 U14098 ( .B1(n16054), .B2(n11230), .A(n11231), .ZN(n18862) );
  INV_X1 U14099 ( .A(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n14797) );
  INV_X1 U14100 ( .A(n11232), .ZN(n11237) );
  AND2_X1 U14101 ( .A1(n11232), .A2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11239) );
  AOI21_X1 U14102 ( .B1(n14797), .B2(n11237), .A(n11239), .ZN(n18868) );
  NOR2_X1 U14103 ( .A1(n13836), .A2(n11233), .ZN(n11238) );
  AOI21_X1 U14104 ( .B1(n13836), .B2(n11233), .A(n11238), .ZN(n18900) );
  AOI21_X1 U14105 ( .B1(n19094), .B2(n11234), .A(n11235), .ZN(n19079) );
  INV_X1 U14106 ( .A(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n13007) );
  AOI21_X1 U14107 ( .B1(n13017), .B2(n13007), .A(n11236), .ZN(n13462) );
  AOI22_X1 U14108 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n18715), .ZN(n18939) );
  AOI22_X1 U14109 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(n13007), .B2(n18715), .ZN(
        n13504) );
  NAND2_X1 U14110 ( .A1(n18939), .A2(n13504), .ZN(n13503) );
  NOR2_X1 U14111 ( .A1(n13462), .A2(n13503), .ZN(n13543) );
  OAI21_X1 U14112 ( .B1(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n11236), .A(
        n11234), .ZN(n13544) );
  NAND2_X1 U14113 ( .A1(n13543), .A2(n13544), .ZN(n13476) );
  NOR2_X1 U14114 ( .A1(n19079), .A2(n13476), .ZN(n18911) );
  OAI21_X1 U14115 ( .B1(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n11235), .A(
        n11233), .ZN(n18913) );
  NAND2_X1 U14116 ( .A1(n18911), .A2(n18913), .ZN(n18898) );
  NOR2_X1 U14117 ( .A1(n18900), .A2(n18898), .ZN(n18879) );
  OAI21_X1 U14118 ( .B1(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n11238), .A(
        n11237), .ZN(n18881) );
  NAND2_X1 U14119 ( .A1(n18879), .A2(n18881), .ZN(n18866) );
  NOR2_X1 U14120 ( .A1(n18868), .A2(n18866), .ZN(n13533) );
  OAI21_X1 U14121 ( .B1(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n11239), .A(
        n11230), .ZN(n16055) );
  NAND2_X1 U14122 ( .A1(n13533), .A2(n16055), .ZN(n18860) );
  NOR2_X1 U14123 ( .A1(n18862), .A2(n18860), .ZN(n18851) );
  OAI21_X1 U14124 ( .B1(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n11231), .A(
        n11228), .ZN(n18854) );
  NAND2_X1 U14125 ( .A1(n18851), .A2(n18854), .ZN(n18830) );
  NOR2_X1 U14126 ( .A1(n18832), .A2(n18830), .ZN(n18818) );
  OAI21_X1 U14127 ( .B1(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n11229), .A(
        n11227), .ZN(n18823) );
  NAND2_X1 U14128 ( .A1(n18818), .A2(n18823), .ZN(n18806) );
  NOR2_X1 U14129 ( .A1(n18807), .A2(n18806), .ZN(n18796) );
  OAI21_X1 U14130 ( .B1(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n11241), .A(
        n11240), .ZN(n18798) );
  NAND2_X1 U14131 ( .A1(n18796), .A2(n18798), .ZN(n18785) );
  OAI21_X1 U14132 ( .B1(n18787), .B2(n18785), .A(n18831), .ZN(n18780) );
  NAND2_X1 U14133 ( .A1(n18781), .A2(n18780), .ZN(n18779) );
  NAND2_X1 U14134 ( .A1(n18831), .A2(n18779), .ZN(n18764) );
  OAI21_X1 U14135 ( .B1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n9744), .A(
        n11242), .ZN(n14755) );
  INV_X1 U14136 ( .A(n14755), .ZN(n18754) );
  INV_X1 U14137 ( .A(n18737), .ZN(n11245) );
  AOI21_X1 U14138 ( .B1(n11242), .B2(n11243), .A(n11217), .ZN(n18738) );
  INV_X1 U14139 ( .A(n18738), .ZN(n11244) );
  NAND2_X1 U14140 ( .A1(n11245), .A2(n11244), .ZN(n18735) );
  AOI21_X1 U14141 ( .B1(n15984), .B2(n11219), .A(n11246), .ZN(n15977) );
  OR2_X1 U14142 ( .A1(n12973), .A2(n18912), .ZN(n15922) );
  OAI21_X1 U14143 ( .B1(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n11246), .A(
        n11247), .ZN(n15976) );
  INV_X1 U14144 ( .A(n15976), .ZN(n15926) );
  AOI21_X1 U14145 ( .B1(n15960), .B2(n11247), .A(n11248), .ZN(n15962) );
  NOR2_X1 U14146 ( .A1(n14589), .A2(n15962), .ZN(n14588) );
  OAI21_X1 U14147 ( .B1(n11248), .B2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .A(
        n11249), .ZN(n14721) );
  AOI21_X1 U14148 ( .B1(n15895), .B2(n11249), .A(n11250), .ZN(n15904) );
  OAI21_X1 U14149 ( .B1(n11250), .B2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .A(
        n9734), .ZN(n12960) );
  INV_X1 U14150 ( .A(n12960), .ZN(n15885) );
  AOI21_X1 U14151 ( .B1(n9734), .B2(n14569), .A(n11251), .ZN(n14565) );
  XNOR2_X1 U14152 ( .A(n11251), .B(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n15875) );
  NOR3_X1 U14153 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(P2_STATEBS16_REG_SCAN_IN), .ZN(n15425) );
  NAND2_X1 U14154 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(n15425), .ZN(n18890) );
  NAND2_X1 U14155 ( .A1(n9643), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(
        n11257) );
  AND2_X4 U14156 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n11658) );
  NAND2_X1 U14157 ( .A1(n11391), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(
        n11256) );
  INV_X1 U14158 ( .A(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11253) );
  NAND4_X1 U14159 ( .A1(n11257), .A2(n11256), .A3(n11255), .A4(n11254), .ZN(
        n11266) );
  INV_X1 U14160 ( .A(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n12091) );
  OR2_X1 U14161 ( .A1(n11287), .A2(n12091), .ZN(n11264) );
  INV_X1 U14162 ( .A(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12073) );
  OR2_X1 U14163 ( .A1(n11355), .A2(n12073), .ZN(n11263) );
  NAND2_X1 U14164 ( .A1(n9645), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(
        n11262) );
  NAND2_X1 U14165 ( .A1(n11281), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(
        n11261) );
  NAND4_X1 U14166 ( .A1(n11264), .A2(n11263), .A3(n11262), .A4(n11261), .ZN(
        n11265) );
  NAND2_X1 U14167 ( .A1(n9641), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(
        n11270) );
  NAND2_X1 U14168 ( .A1(n11391), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(
        n11269) );
  NAND2_X1 U14169 ( .A1(n11279), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(
        n11268) );
  INV_X2 U14170 ( .A(n11280), .ZN(n12690) );
  NAND2_X1 U14171 ( .A1(n12690), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(
        n11267) );
  NAND4_X1 U14172 ( .A1(n11270), .A2(n11269), .A3(n11268), .A4(n11267), .ZN(
        n11276) );
  INV_X1 U14173 ( .A(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12074) );
  INV_X1 U14174 ( .A(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n19161) );
  NAND2_X1 U14175 ( .A1(n11656), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(
        n11272) );
  NAND2_X1 U14176 ( .A1(n11281), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(
        n11271) );
  NAND4_X1 U14177 ( .A1(n11274), .A2(n11273), .A3(n11272), .A4(n11271), .ZN(
        n11275) );
  NOR2_X1 U14178 ( .A1(n11276), .A2(n11275), .ZN(n11409) );
  AOI22_X1 U14179 ( .A1(n12687), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n9643), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11285) );
  INV_X4 U14180 ( .A(n11287), .ZN(n12841) );
  AOI22_X1 U14181 ( .A1(n9642), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(n9641), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11284) );
  INV_X2 U14182 ( .A(n11280), .ZN(n12846) );
  AOI22_X1 U14183 ( .A1(n11281), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n11656), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11282) );
  NAND4_X1 U14184 ( .A1(n11285), .A2(n11284), .A3(n11283), .A4(n11282), .ZN(
        n11286) );
  NAND2_X1 U14185 ( .A1(n11286), .A2(n11278), .ZN(n11297) );
  AOI22_X1 U14186 ( .A1(n9643), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .B1(n9641), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11293) );
  AOI22_X1 U14187 ( .A1(n11281), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n11656), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11292) );
  INV_X1 U14188 ( .A(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11289) );
  INV_X1 U14189 ( .A(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11288) );
  INV_X1 U14190 ( .A(n11290), .ZN(n11291) );
  NAND4_X1 U14191 ( .A1(n11294), .A2(n11293), .A3(n11292), .A4(n11291), .ZN(
        n11295) );
  NAND2_X1 U14192 ( .A1(n11295), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11296) );
  NAND2_X1 U14193 ( .A1(n11297), .A2(n11296), .ZN(n11414) );
  NAND2_X1 U14194 ( .A1(n11279), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(
        n11301) );
  NAND2_X1 U14195 ( .A1(n11391), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(
        n11300) );
  NAND2_X1 U14196 ( .A1(n9641), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(
        n11299) );
  NAND2_X1 U14197 ( .A1(n12690), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n11298) );
  NAND4_X1 U14198 ( .A1(n11301), .A2(n11300), .A3(n11299), .A4(n11298), .ZN(
        n11309) );
  INV_X1 U14199 ( .A(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n11302) );
  INV_X1 U14200 ( .A(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n11303) );
  OR2_X1 U14201 ( .A1(n11355), .A2(n11303), .ZN(n11306) );
  NAND2_X1 U14202 ( .A1(n9645), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(
        n11305) );
  NAND2_X1 U14203 ( .A1(n11281), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n11304) );
  NAND2_X1 U14204 ( .A1(n11405), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11322) );
  NAND2_X1 U14205 ( .A1(n9643), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n11313) );
  NAND2_X1 U14206 ( .A1(n11391), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(
        n11312) );
  NAND2_X1 U14207 ( .A1(n9641), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(
        n11311) );
  NAND2_X1 U14208 ( .A1(n9644), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(
        n11310) );
  NAND4_X1 U14209 ( .A1(n11313), .A2(n11312), .A3(n11311), .A4(n11310), .ZN(
        n11320) );
  INV_X1 U14210 ( .A(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11314) );
  INV_X1 U14211 ( .A(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12545) );
  OR2_X1 U14212 ( .A1(n11355), .A2(n12545), .ZN(n11317) );
  NAND2_X1 U14213 ( .A1(n11656), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(
        n11316) );
  NAND2_X1 U14214 ( .A1(n11281), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n11315) );
  NAND4_X1 U14215 ( .A1(n11318), .A2(n11317), .A3(n11316), .A4(n11315), .ZN(
        n11319) );
  NAND2_X1 U14216 ( .A1(n11411), .A2(n11347), .ZN(n11321) );
  NAND2_X1 U14217 ( .A1(n11279), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(
        n11326) );
  NAND2_X1 U14218 ( .A1(n11391), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(
        n11325) );
  NAND2_X1 U14219 ( .A1(n9641), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n11324) );
  NAND2_X1 U14220 ( .A1(n12846), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(
        n11323) );
  INV_X1 U14221 ( .A(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n11327) );
  NOR2_X1 U14222 ( .A1(n11287), .A2(n11327), .ZN(n11333) );
  INV_X1 U14223 ( .A(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n11328) );
  OR2_X1 U14224 ( .A1(n11355), .A2(n11328), .ZN(n11331) );
  NAND2_X1 U14225 ( .A1(n11281), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(
        n11330) );
  NAND2_X1 U14226 ( .A1(n9645), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(
        n11329) );
  NAND3_X1 U14227 ( .A1(n11331), .A2(n11330), .A3(n11329), .ZN(n11332) );
  NOR2_X1 U14228 ( .A1(n11333), .A2(n11332), .ZN(n11334) );
  NAND2_X1 U14229 ( .A1(n11279), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(
        n11338) );
  NAND2_X1 U14230 ( .A1(n11391), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(
        n11337) );
  NAND2_X1 U14231 ( .A1(n9641), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(
        n11336) );
  NAND2_X1 U14232 ( .A1(n9637), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(
        n11335) );
  NAND4_X1 U14233 ( .A1(n11338), .A2(n11337), .A3(n11336), .A4(n11335), .ZN(
        n11345) );
  INV_X1 U14234 ( .A(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11339) );
  INV_X1 U14235 ( .A(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12544) );
  OR2_X1 U14236 ( .A1(n11355), .A2(n12544), .ZN(n11342) );
  NAND2_X1 U14237 ( .A1(n9645), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(
        n11341) );
  NAND2_X1 U14238 ( .A1(n11281), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(
        n11340) );
  NAND4_X1 U14239 ( .A1(n11343), .A2(n11342), .A3(n11341), .A4(n11340), .ZN(
        n11344) );
  NOR2_X1 U14240 ( .A1(n11345), .A2(n11344), .ZN(n11410) );
  NAND2_X1 U14241 ( .A1(n11410), .A2(n11347), .ZN(n11346) );
  INV_X1 U14242 ( .A(n11400), .ZN(n11449) );
  AND3_X2 U14243 ( .A1(n11348), .A2(n11450), .A3(n11449), .ZN(n11442) );
  AOI22_X1 U14244 ( .A1(n9643), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n11391), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11352) );
  AOI22_X1 U14245 ( .A1(n12845), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n12846), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n11351) );
  AOI22_X1 U14246 ( .A1(n11281), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n11656), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11349) );
  NAND4_X1 U14247 ( .A1(n11353), .A2(n11352), .A3(n11351), .A4(n11350), .ZN(
        n11362) );
  AOI22_X1 U14248 ( .A1(n11281), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n9645), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11354) );
  AOI22_X1 U14249 ( .A1(n9641), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(n9644), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11359) );
  INV_X1 U14250 ( .A(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12815) );
  INV_X1 U14251 ( .A(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n19175) );
  OAI22_X1 U14252 ( .A1(n11287), .A2(n12815), .B1(n11355), .B2(n19175), .ZN(
        n11356) );
  INV_X1 U14253 ( .A(n11356), .ZN(n11358) );
  AOI22_X1 U14254 ( .A1(n9643), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n11391), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11357) );
  NAND4_X1 U14255 ( .A1(n11360), .A2(n11359), .A3(n11358), .A4(n11357), .ZN(
        n11361) );
  AOI22_X1 U14256 ( .A1(n9641), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n12690), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11364) );
  AOI22_X1 U14257 ( .A1(n11281), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n9645), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11363) );
  AOI22_X1 U14258 ( .A1(n11279), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n11391), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11366) );
  AOI22_X1 U14259 ( .A1(n12841), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n12687), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11365) );
  NAND3_X1 U14260 ( .A1(n11367), .A2(n11366), .A3(n11365), .ZN(n11374) );
  AOI22_X1 U14261 ( .A1(n9641), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n12846), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n11369) );
  AOI22_X1 U14262 ( .A1(n11281), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n11656), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11368) );
  AND3_X1 U14263 ( .A1(n11369), .A2(n11368), .A3(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11372) );
  AOI22_X1 U14264 ( .A1(n9643), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n11391), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11371) );
  AOI22_X1 U14265 ( .A1(n12841), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12687), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11370) );
  NAND3_X1 U14266 ( .A1(n11372), .A2(n11371), .A3(n11370), .ZN(n11373) );
  AOI22_X1 U14267 ( .A1(n11281), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n9645), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n11375) );
  AOI22_X1 U14268 ( .A1(n9643), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n12845), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11379) );
  AOI22_X1 U14269 ( .A1(n11391), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n9644), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n11378) );
  AOI22_X1 U14270 ( .A1(n12841), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12687), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n11377) );
  NAND4_X1 U14271 ( .A1(n11380), .A2(n11379), .A3(n11378), .A4(n11377), .ZN(
        n11388) );
  AOI22_X1 U14272 ( .A1(n11281), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n11656), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11381) );
  AOI22_X1 U14273 ( .A1(n12687), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n11279), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11385) );
  AOI22_X1 U14274 ( .A1(n11391), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n12846), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11384) );
  AOI22_X1 U14275 ( .A1(n12841), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n12845), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n11383) );
  NAND4_X1 U14276 ( .A1(n11386), .A2(n11385), .A3(n11384), .A4(n11383), .ZN(
        n11387) );
  AOI22_X1 U14277 ( .A1(n12841), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n12687), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11395) );
  AOI22_X1 U14278 ( .A1(n11281), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n11656), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11394) );
  AOI22_X1 U14279 ( .A1(n9643), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n11391), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11393) );
  AOI22_X1 U14280 ( .A1(n9641), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n12690), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n11392) );
  AOI22_X1 U14281 ( .A1(n11281), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n9645), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11396) );
  AOI22_X1 U14282 ( .A1(n9641), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n12690), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11397) );
  NOR2_X1 U14283 ( .A1(n11434), .A2(n11630), .ZN(n12876) );
  INV_X1 U14284 ( .A(n11414), .ZN(n11436) );
  INV_X1 U14285 ( .A(n11401), .ZN(n11640) );
  NAND4_X1 U14286 ( .A1(n12876), .A2(n12452), .A3(n9631), .A4(n13063), .ZN(
        n11403) );
  INV_X1 U14287 ( .A(n11434), .ZN(n11420) );
  INV_X1 U14288 ( .A(n13063), .ZN(n11404) );
  AND2_X1 U14289 ( .A1(n12376), .A2(n13728), .ZN(n11471) );
  INV_X1 U14290 ( .A(n11405), .ZN(n11408) );
  INV_X1 U14291 ( .A(n11406), .ZN(n11407) );
  INV_X1 U14292 ( .A(n11410), .ZN(n11413) );
  INV_X1 U14293 ( .A(n11411), .ZN(n11412) );
  NAND4_X1 U14294 ( .A1(n11409), .A2(n11413), .A3(n11412), .A4(n11347), .ZN(
        n11415) );
  AOI21_X1 U14295 ( .B1(n11416), .B2(n11415), .A(n13574), .ZN(n11417) );
  INV_X1 U14296 ( .A(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n12269) );
  OR2_X1 U14297 ( .A1(n11609), .A2(n12269), .ZN(n11426) );
  INV_X1 U14298 ( .A(P2_EBX_REG_15__SCAN_IN), .ZN(n11421) );
  NOR2_X1 U14299 ( .A1(n12475), .A2(n11421), .ZN(n11424) );
  INV_X1 U14300 ( .A(P2_REIP_REG_15__SCAN_IN), .ZN(n11422) );
  INV_X1 U14301 ( .A(P2_STATE2_REG_1__SCAN_IN), .ZN(n13649) );
  OAI22_X1 U14302 ( .A1(n11606), .A2(n11422), .B1(n13649), .B2(n11215), .ZN(
        n11423) );
  NOR2_X1 U14303 ( .A1(n11424), .A2(n11423), .ZN(n11425) );
  NAND2_X1 U14304 ( .A1(n11426), .A2(n11425), .ZN(n13720) );
  INV_X1 U14305 ( .A(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n15029) );
  OR2_X1 U14306 ( .A1(n11609), .A2(n15029), .ZN(n11432) );
  INV_X1 U14307 ( .A(P2_EBX_REG_9__SCAN_IN), .ZN(n11429) );
  NAND2_X1 U14308 ( .A1(n12472), .A2(P2_REIP_REG_9__SCAN_IN), .ZN(n11428) );
  NAND2_X1 U14309 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n11427) );
  OAI211_X1 U14310 ( .C1(n11592), .C2(n11429), .A(n11428), .B(n11427), .ZN(
        n11430) );
  INV_X1 U14311 ( .A(n11430), .ZN(n11431) );
  INV_X1 U14312 ( .A(n13065), .ZN(n11440) );
  OAI21_X1 U14313 ( .B1(n11630), .B2(n11450), .A(n11433), .ZN(n11438) );
  INV_X1 U14314 ( .A(n11435), .ZN(n12459) );
  NAND2_X1 U14315 ( .A1(n11470), .A2(n12459), .ZN(n11437) );
  NAND4_X1 U14316 ( .A1(n11438), .A2(n11437), .A3(n11436), .A4(n11451), .ZN(
        n11439) );
  NAND3_X1 U14317 ( .A1(n11440), .A2(n11439), .A3(n13728), .ZN(n12456) );
  INV_X1 U14318 ( .A(n12456), .ZN(n11441) );
  NAND2_X1 U14319 ( .A1(n11441), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n11448) );
  NAND2_X1 U14320 ( .A1(n11442), .A2(n12375), .ZN(n12367) );
  NAND2_X1 U14321 ( .A1(n12367), .A2(n11443), .ZN(n11444) );
  NAND2_X1 U14322 ( .A1(n11444), .A2(n12374), .ZN(n12442) );
  NAND2_X1 U14323 ( .A1(n12442), .A2(n11389), .ZN(n11446) );
  NAND2_X1 U14324 ( .A1(n11470), .A2(n11635), .ZN(n12451) );
  INV_X1 U14325 ( .A(n12355), .ZN(n13156) );
  NAND2_X1 U14326 ( .A1(n11481), .A2(n13156), .ZN(n11445) );
  NAND2_X1 U14327 ( .A1(n11446), .A2(n11445), .ZN(n11447) );
  AND2_X2 U14328 ( .A1(n11448), .A2(n11447), .ZN(n11479) );
  INV_X1 U14329 ( .A(n11450), .ZN(n12379) );
  NAND2_X1 U14330 ( .A1(n11470), .A2(n12379), .ZN(n12384) );
  AND2_X1 U14331 ( .A1(n12384), .A2(n9639), .ZN(n11453) );
  INV_X1 U14332 ( .A(n12376), .ZN(n11452) );
  NAND3_X1 U14333 ( .A1(n11452), .A2(n11450), .A3(n11451), .ZN(n12383) );
  NAND2_X1 U14334 ( .A1(n12457), .A2(n12459), .ZN(n11456) );
  INV_X1 U14335 ( .A(n11454), .ZN(n12453) );
  NAND2_X1 U14336 ( .A1(n11480), .A2(n9654), .ZN(n11457) );
  NAND2_X1 U14337 ( .A1(n11497), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11461) );
  NOR2_X1 U14338 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n11510) );
  NAND2_X1 U14339 ( .A1(n11461), .A2(n11460), .ZN(n11466) );
  INV_X1 U14340 ( .A(n11466), .ZN(n11465) );
  INV_X1 U14341 ( .A(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n11463) );
  INV_X1 U14342 ( .A(P2_EBX_REG_1__SCAN_IN), .ZN(n11988) );
  NAND2_X1 U14343 ( .A1(n11467), .A2(n11466), .ZN(n11468) );
  AND2_X1 U14344 ( .A1(n9654), .A2(n12452), .ZN(n11469) );
  OAI22_X1 U14345 ( .A1(n11497), .A2(n11469), .B1(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n11558), .ZN(n11476) );
  INV_X1 U14346 ( .A(n11470), .ZN(n12864) );
  MUX2_X1 U14347 ( .A(n12864), .B(n11471), .S(n19156), .Z(n11473) );
  NOR2_X1 U14348 ( .A1(n11450), .A2(n11630), .ZN(n11472) );
  AOI22_X1 U14349 ( .A1(n13589), .A2(P2_STATE2_REG_0__SCAN_IN), .B1(n11510), 
        .B2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n11475) );
  NAND2_X1 U14350 ( .A1(n11476), .A2(n11475), .ZN(n12022) );
  INV_X1 U14351 ( .A(n11477), .ZN(n11478) );
  INV_X1 U14352 ( .A(n11480), .ZN(n11482) );
  INV_X1 U14353 ( .A(P2_EBX_REG_0__SCAN_IN), .ZN(n11989) );
  INV_X1 U14354 ( .A(n11492), .ZN(n11483) );
  NAND2_X1 U14355 ( .A1(n11483), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n11486) );
  INV_X1 U14356 ( .A(n11510), .ZN(n13587) );
  NAND2_X1 U14357 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n11484) );
  AND2_X1 U14358 ( .A1(n13587), .A2(n11484), .ZN(n11485) );
  OAI211_X1 U14359 ( .C1(n11989), .C2(n12475), .A(n11486), .B(n11485), .ZN(
        n11487) );
  INV_X1 U14360 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n12448) );
  AOI22_X1 U14361 ( .A1(n11483), .A2(P2_REIP_REG_2__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n11493) );
  OAI21_X1 U14362 ( .B1(n19764), .B2(P2_STATE2_REG_0__SCAN_IN), .A(n13649), 
        .ZN(n11498) );
  INV_X1 U14364 ( .A(n11499), .ZN(n11500) );
  NAND2_X1 U14365 ( .A1(n11501), .A2(n11500), .ZN(n11502) );
  NAND2_X2 U14366 ( .A1(n11503), .A2(n11502), .ZN(n12014) );
  INV_X1 U14367 ( .A(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n12162) );
  INV_X1 U14368 ( .A(P2_EBX_REG_3__SCAN_IN), .ZN(n13551) );
  NOR2_X1 U14369 ( .A1(n11592), .A2(n13551), .ZN(n11507) );
  INV_X1 U14370 ( .A(P2_REIP_REG_3__SCAN_IN), .ZN(n11505) );
  INV_X1 U14371 ( .A(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n11504) );
  OAI22_X1 U14372 ( .A1(n11606), .A2(n11505), .B1(n13649), .B2(n11504), .ZN(
        n11506) );
  NOR2_X1 U14373 ( .A1(n11507), .A2(n11506), .ZN(n11508) );
  NAND2_X1 U14374 ( .A1(n11497), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11512) );
  NAND2_X1 U14375 ( .A1(n11510), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n11511) );
  XNOR2_X2 U14376 ( .A(n11514), .B(n11513), .ZN(n12013) );
  NAND2_X1 U14377 ( .A1(n12014), .A2(n12013), .ZN(n11517) );
  INV_X1 U14378 ( .A(n11513), .ZN(n11515) );
  NAND2_X1 U14379 ( .A1(n11515), .A2(n11514), .ZN(n11516) );
  NAND2_X1 U14380 ( .A1(n11517), .A2(n11516), .ZN(n13086) );
  INV_X1 U14381 ( .A(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n19101) );
  OR2_X1 U14382 ( .A1(n11609), .A2(n19101), .ZN(n11523) );
  INV_X1 U14383 ( .A(P2_EBX_REG_4__SCAN_IN), .ZN(n11520) );
  NAND2_X1 U14384 ( .A1(n12472), .A2(P2_REIP_REG_4__SCAN_IN), .ZN(n11519) );
  NAND2_X1 U14385 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n11518) );
  OAI211_X1 U14386 ( .C1(n11520), .C2(n12475), .A(n11519), .B(n11518), .ZN(
        n11521) );
  INV_X1 U14387 ( .A(n11521), .ZN(n11522) );
  INV_X1 U14388 ( .A(P2_EBX_REG_5__SCAN_IN), .ZN(n18905) );
  INV_X1 U14389 ( .A(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n12418) );
  OR2_X1 U14390 ( .A1(n11609), .A2(n12418), .ZN(n11525) );
  AOI22_X1 U14391 ( .A1(n12472), .A2(P2_REIP_REG_5__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n11524) );
  OAI211_X1 U14392 ( .C1(n11592), .C2(n18905), .A(n11525), .B(n11524), .ZN(
        n13133) );
  NAND2_X1 U14393 ( .A1(n13087), .A2(n13133), .ZN(n13244) );
  INV_X1 U14394 ( .A(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n14055) );
  INV_X1 U14395 ( .A(P2_EBX_REG_6__SCAN_IN), .ZN(n18894) );
  NOR2_X1 U14396 ( .A1(n11592), .A2(n18894), .ZN(n11528) );
  INV_X1 U14397 ( .A(P2_REIP_REG_6__SCAN_IN), .ZN(n11526) );
  OAI22_X1 U14398 ( .A1(n11606), .A2(n11526), .B1(n13649), .B2(n13836), .ZN(
        n11527) );
  NOR2_X1 U14399 ( .A1(n11528), .A2(n11527), .ZN(n11529) );
  INV_X1 U14400 ( .A(P2_EBX_REG_7__SCAN_IN), .ZN(n11533) );
  INV_X1 U14401 ( .A(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n13822) );
  OR2_X1 U14402 ( .A1(n11609), .A2(n13822), .ZN(n11532) );
  AOI22_X1 U14403 ( .A1(n12472), .A2(P2_REIP_REG_7__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n11531) );
  OAI211_X1 U14404 ( .C1(n11592), .C2(n11533), .A(n11532), .B(n11531), .ZN(
        n13274) );
  INV_X1 U14405 ( .A(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n16118) );
  OR2_X1 U14406 ( .A1(n11609), .A2(n16118), .ZN(n11538) );
  INV_X1 U14407 ( .A(P2_EBX_REG_8__SCAN_IN), .ZN(n18869) );
  NAND2_X1 U14408 ( .A1(n12472), .A2(P2_REIP_REG_8__SCAN_IN), .ZN(n11535) );
  NAND2_X1 U14409 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n11534) );
  OAI211_X1 U14410 ( .C1(n18869), .C2(n12475), .A(n11535), .B(n11534), .ZN(
        n11536) );
  INV_X1 U14411 ( .A(n11536), .ZN(n11537) );
  INV_X1 U14412 ( .A(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n15006) );
  OR2_X1 U14413 ( .A1(n11609), .A2(n15006), .ZN(n11540) );
  AOI22_X1 U14414 ( .A1(n12472), .A2(P2_REIP_REG_10__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), 
        .ZN(n11539) );
  OAI211_X1 U14415 ( .C1(n11592), .C2(n10059), .A(n11540), .B(n11539), .ZN(
        n15009) );
  INV_X1 U14416 ( .A(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n14988) );
  OR2_X1 U14417 ( .A1(n11609), .A2(n14988), .ZN(n11546) );
  INV_X1 U14418 ( .A(P2_EBX_REG_11__SCAN_IN), .ZN(n11541) );
  NOR2_X1 U14419 ( .A1(n11592), .A2(n11541), .ZN(n11544) );
  INV_X1 U14420 ( .A(P2_REIP_REG_11__SCAN_IN), .ZN(n14989) );
  INV_X1 U14421 ( .A(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n11542) );
  OAI22_X1 U14422 ( .A1(n11606), .A2(n14989), .B1(n13649), .B2(n11542), .ZN(
        n11543) );
  NOR2_X1 U14423 ( .A1(n11544), .A2(n11543), .ZN(n11545) );
  INV_X1 U14424 ( .A(P2_EBX_REG_12__SCAN_IN), .ZN(n11549) );
  INV_X1 U14425 ( .A(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n16106) );
  OR2_X1 U14426 ( .A1(n11609), .A2(n16106), .ZN(n11548) );
  AOI22_X1 U14427 ( .A1(n12472), .A2(P2_REIP_REG_12__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), 
        .ZN(n11547) );
  OAI211_X1 U14428 ( .C1(n11592), .C2(n11549), .A(n11548), .B(n11547), .ZN(
        n13362) );
  INV_X1 U14429 ( .A(P2_EBX_REG_13__SCAN_IN), .ZN(n11552) );
  INV_X1 U14430 ( .A(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n16085) );
  OR2_X1 U14431 ( .A1(n11609), .A2(n16085), .ZN(n11551) );
  AOI22_X1 U14432 ( .A1(n12472), .A2(P2_REIP_REG_13__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_13__SCAN_IN), 
        .ZN(n11550) );
  OAI211_X1 U14433 ( .C1(n11552), .C2(n11592), .A(n11551), .B(n11550), .ZN(
        n14171) );
  INV_X1 U14434 ( .A(P2_EBX_REG_14__SCAN_IN), .ZN(n18808) );
  AOI22_X1 U14435 ( .A1(n12472), .A2(P2_REIP_REG_14__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), 
        .ZN(n11553) );
  OAI21_X1 U14436 ( .B1(n11592), .B2(n18808), .A(n11553), .ZN(n11554) );
  AOI21_X1 U14437 ( .B1(n11608), .B2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A(
        n11554), .ZN(n13520) );
  INV_X1 U14438 ( .A(P2_EBX_REG_16__SCAN_IN), .ZN(n11557) );
  INV_X1 U14439 ( .A(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15317) );
  OR2_X1 U14440 ( .A1(n11609), .A2(n15317), .ZN(n11556) );
  AOI22_X1 U14441 ( .A1(n12472), .A2(P2_REIP_REG_16__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), 
        .ZN(n11555) );
  OAI211_X1 U14442 ( .C1(n11592), .C2(n11557), .A(n11556), .B(n11555), .ZN(
        n15290) );
  NAND2_X1 U14443 ( .A1(n11558), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n11560) );
  NAND2_X1 U14444 ( .A1(n12472), .A2(P2_REIP_REG_17__SCAN_IN), .ZN(n11559) );
  OAI211_X1 U14445 ( .C1(n13649), .C2(n18771), .A(n11560), .B(n11559), .ZN(
        n11561) );
  AOI21_X1 U14446 ( .B1(n11608), .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        n11561), .ZN(n14041) );
  INV_X1 U14447 ( .A(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n14952) );
  OR2_X1 U14448 ( .A1(n11609), .A2(n14952), .ZN(n11566) );
  INV_X1 U14449 ( .A(P2_REIP_REG_18__SCAN_IN), .ZN(n19711) );
  NAND2_X1 U14450 ( .A1(n11558), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n11563) );
  NAND2_X1 U14451 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n11562) );
  OAI211_X1 U14452 ( .C1(n11606), .C2(n19711), .A(n11563), .B(n11562), .ZN(
        n11564) );
  INV_X1 U14453 ( .A(n11564), .ZN(n11565) );
  NAND2_X1 U14454 ( .A1(n11566), .A2(n11565), .ZN(n14780) );
  NAND2_X1 U14455 ( .A1(n14042), .A2(n14780), .ZN(n14059) );
  INV_X1 U14456 ( .A(P2_REIP_REG_19__SCAN_IN), .ZN(n19713) );
  NAND2_X1 U14457 ( .A1(n11558), .A2(P2_EBX_REG_19__SCAN_IN), .ZN(n11568) );
  NAND2_X1 U14458 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n11567) );
  OAI211_X1 U14459 ( .C1(n11606), .C2(n19713), .A(n11568), .B(n11567), .ZN(
        n11569) );
  AOI21_X1 U14460 ( .B1(n11608), .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A(
        n11569), .ZN(n14060) );
  INV_X1 U14461 ( .A(P2_EBX_REG_20__SCAN_IN), .ZN(n11572) );
  NAND2_X1 U14462 ( .A1(n12472), .A2(P2_REIP_REG_20__SCAN_IN), .ZN(n11571) );
  NAND2_X1 U14463 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n11570) );
  OAI211_X1 U14464 ( .C1(n11572), .C2(n12475), .A(n11571), .B(n11570), .ZN(
        n11573) );
  AOI21_X1 U14465 ( .B1(n11608), .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A(
        n11573), .ZN(n14756) );
  INV_X1 U14466 ( .A(P2_REIP_REG_21__SCAN_IN), .ZN(n19717) );
  NAND2_X1 U14467 ( .A1(n11558), .A2(P2_EBX_REG_21__SCAN_IN), .ZN(n11575) );
  NAND2_X1 U14468 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n11574) );
  OAI211_X1 U14469 ( .C1(n11606), .C2(n19717), .A(n11575), .B(n11574), .ZN(
        n11576) );
  AOI21_X1 U14470 ( .B1(n11608), .B2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A(
        n11576), .ZN(n14636) );
  INV_X1 U14471 ( .A(P2_EBX_REG_22__SCAN_IN), .ZN(n15307) );
  INV_X1 U14472 ( .A(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n14910) );
  OR2_X1 U14473 ( .A1(n11609), .A2(n14910), .ZN(n11578) );
  AOI22_X1 U14474 ( .A1(n12472), .A2(P2_REIP_REG_22__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), 
        .ZN(n11577) );
  OAI211_X1 U14475 ( .C1(n11592), .C2(n15307), .A(n11578), .B(n11577), .ZN(
        n14915) );
  INV_X1 U14476 ( .A(P2_REIP_REG_23__SCAN_IN), .ZN(n11581) );
  NAND2_X1 U14477 ( .A1(n11558), .A2(P2_EBX_REG_23__SCAN_IN), .ZN(n11580) );
  NAND2_X1 U14478 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n11579) );
  OAI211_X1 U14479 ( .C1(n11606), .C2(n11581), .A(n11580), .B(n11579), .ZN(
        n11582) );
  AOI21_X1 U14480 ( .B1(n11608), .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n11582), .ZN(n12978) );
  NAND2_X1 U14481 ( .A1(n12472), .A2(P2_REIP_REG_24__SCAN_IN), .ZN(n11584) );
  NAND2_X1 U14482 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n11583) );
  OAI211_X1 U14483 ( .C1(n11592), .C2(n10056), .A(n11584), .B(n11583), .ZN(
        n11585) );
  AOI21_X1 U14484 ( .B1(n11608), .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A(
        n11585), .ZN(n14631) );
  INV_X1 U14485 ( .A(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n11586) );
  OR2_X1 U14486 ( .A1(n11609), .A2(n11586), .ZN(n11591) );
  INV_X1 U14487 ( .A(P2_EBX_REG_25__SCAN_IN), .ZN(n11587) );
  NOR2_X1 U14488 ( .A1(n11592), .A2(n11587), .ZN(n11589) );
  INV_X1 U14489 ( .A(P2_REIP_REG_25__SCAN_IN), .ZN(n19724) );
  OAI22_X1 U14490 ( .A1(n11606), .A2(n19724), .B1(n13649), .B2(n15960), .ZN(
        n11588) );
  NOR2_X1 U14491 ( .A1(n11589), .A2(n11588), .ZN(n11590) );
  NAND2_X1 U14492 ( .A1(n11591), .A2(n11590), .ZN(n14581) );
  INV_X1 U14493 ( .A(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n11967) );
  OR2_X1 U14494 ( .A1(n11609), .A2(n11967), .ZN(n11597) );
  INV_X1 U14495 ( .A(P2_EBX_REG_26__SCAN_IN), .ZN(n12002) );
  NOR2_X1 U14496 ( .A1(n11592), .A2(n12002), .ZN(n11595) );
  INV_X1 U14497 ( .A(P2_REIP_REG_26__SCAN_IN), .ZN(n11593) );
  INV_X1 U14498 ( .A(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n14720) );
  OAI22_X1 U14499 ( .A1(n11606), .A2(n11593), .B1(n13649), .B2(n14720), .ZN(
        n11594) );
  NOR2_X1 U14500 ( .A1(n11595), .A2(n11594), .ZN(n11596) );
  NAND2_X1 U14501 ( .A1(n11597), .A2(n11596), .ZN(n14615) );
  INV_X1 U14502 ( .A(P2_REIP_REG_27__SCAN_IN), .ZN(n19728) );
  NAND2_X1 U14503 ( .A1(n11558), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n11599) );
  NAND2_X1 U14504 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n11598) );
  OAI211_X1 U14505 ( .C1(n11606), .C2(n19728), .A(n11599), .B(n11598), .ZN(
        n11600) );
  AOI21_X1 U14506 ( .B1(n11608), .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n11600), .ZN(n14612) );
  INV_X1 U14507 ( .A(P2_REIP_REG_28__SCAN_IN), .ZN(n19729) );
  NAND2_X1 U14508 ( .A1(n11558), .A2(P2_EBX_REG_28__SCAN_IN), .ZN(n11602) );
  NAND2_X1 U14509 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n11601) );
  OAI211_X1 U14510 ( .C1(n11606), .C2(n19729), .A(n11602), .B(n11601), .ZN(
        n11603) );
  AOI21_X1 U14511 ( .B1(n11608), .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n11603), .ZN(n12947) );
  INV_X1 U14512 ( .A(P2_REIP_REG_29__SCAN_IN), .ZN(n19731) );
  NAND2_X1 U14513 ( .A1(n11558), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n11605) );
  NAND2_X1 U14514 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n11604) );
  OAI211_X1 U14515 ( .C1(n11606), .C2(n19731), .A(n11605), .B(n11604), .ZN(
        n11607) );
  AOI21_X1 U14516 ( .B1(n11608), .B2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        n11607), .ZN(n12506) );
  INV_X1 U14517 ( .A(P2_EBX_REG_30__SCAN_IN), .ZN(n12007) );
  INV_X1 U14518 ( .A(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n12490) );
  OR2_X1 U14519 ( .A1(n11609), .A2(n12490), .ZN(n11611) );
  AOI22_X1 U14520 ( .A1(n12472), .A2(P2_REIP_REG_30__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), 
        .ZN(n11610) );
  OAI211_X1 U14521 ( .C1(n12007), .C2(n12475), .A(n11611), .B(n11610), .ZN(
        n12469) );
  NAND2_X1 U14522 ( .A1(n19773), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11614) );
  NAND2_X1 U14523 ( .A1(n11612), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n11613) );
  NAND2_X1 U14524 ( .A1(n11614), .A2(n11613), .ZN(n12359) );
  NAND2_X1 U14525 ( .A1(n19764), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11617) );
  NAND2_X1 U14526 ( .A1(n13620), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n11616) );
  MUX2_X1 U14527 ( .A(n19757), .B(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .S(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n11620) );
  INV_X1 U14528 ( .A(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n13643) );
  INV_X1 U14529 ( .A(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n15428) );
  NOR2_X1 U14530 ( .A1(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n15428), .ZN(
        n11618) );
  INV_X1 U14531 ( .A(n12154), .ZN(n11619) );
  XNOR2_X1 U14532 ( .A(n12359), .B(n11619), .ZN(n12341) );
  NOR2_X1 U14533 ( .A1(n11621), .A2(n11620), .ZN(n11622) );
  OAI21_X1 U14534 ( .B1(n11626), .B2(n11625), .A(n11624), .ZN(n12336) );
  NOR3_X1 U14535 ( .A1(n12346), .A2(n12336), .A3(n12352), .ZN(n12369) );
  AND2_X1 U14536 ( .A1(n12341), .A2(n12369), .ZN(n11628) );
  NAND2_X1 U14537 ( .A1(n13649), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n19658) );
  OR2_X1 U14538 ( .A1(n19658), .A2(n19801), .ZN(n16152) );
  AND2_X1 U14539 ( .A1(n11458), .A2(n13152), .ZN(n13641) );
  NAND2_X1 U14540 ( .A1(n19804), .A2(n12463), .ZN(n11987) );
  NAND2_X1 U14541 ( .A1(READY21_REG_SCAN_IN), .A2(READY12_REG_SCAN_IN), .ZN(
        n15424) );
  INV_X1 U14542 ( .A(n15424), .ZN(n19807) );
  NOR2_X2 U14543 ( .A1(n12988), .A2(n9636), .ZN(n19077) );
  NOR2_X1 U14544 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(P2_STATE_REG_2__SCAN_IN), 
        .ZN(n19667) );
  AOI211_X1 U14545 ( .C1(P2_STATE_REG_1__SCAN_IN), .C2(P2_STATE_REG_2__SCAN_IN), .A(P2_STATE_REG_0__SCAN_IN), .B(n19667), .ZN(n19795) );
  NAND2_X1 U14546 ( .A1(n19795), .A2(n15424), .ZN(n13628) );
  NOR2_X1 U14547 ( .A1(n13628), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n13652) );
  NAND2_X1 U14548 ( .A1(n19077), .A2(n13652), .ZN(n18928) );
  INV_X1 U14549 ( .A(P2_REIP_REG_1__SCAN_IN), .ZN(n19685) );
  NAND2_X1 U14550 ( .A1(n11975), .A2(P2_REIP_REG_1__SCAN_IN), .ZN(n11632) );
  AOI22_X1 U14551 ( .A1(n11963), .A2(P2_EAX_REG_1__SCAN_IN), .B1(n11639), .B2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n11631) );
  NAND2_X1 U14552 ( .A1(n11632), .A2(n11631), .ZN(n11684) );
  INV_X1 U14553 ( .A(P2_REIP_REG_0__SCAN_IN), .ZN(n11633) );
  OR2_X1 U14554 ( .A1(n11974), .A2(n11633), .ZN(n11638) );
  INV_X1 U14555 ( .A(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n13762) );
  NAND2_X1 U14556 ( .A1(n11630), .A2(P2_EAX_REG_0__SCAN_IN), .ZN(n11634) );
  OAI211_X1 U14557 ( .C1(n11635), .C2(n13762), .A(n11634), .B(n19594), .ZN(
        n11636) );
  INV_X1 U14558 ( .A(n11636), .ZN(n11637) );
  NAND2_X1 U14559 ( .A1(n11638), .A2(n11637), .ZN(n13040) );
  OR2_X1 U14560 ( .A1(n11969), .A2(n11470), .ZN(n11704) );
  AND2_X2 U14561 ( .A1(n13044), .A2(n12003), .ZN(n11685) );
  INV_X1 U14562 ( .A(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n13732) );
  INV_X1 U14563 ( .A(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n11641) );
  OAI22_X1 U14564 ( .A1(n13732), .A2(n11686), .B1(n11687), .B2(n11641), .ZN(
        n11642) );
  INV_X1 U14565 ( .A(n11642), .ZN(n11654) );
  AOI22_X1 U14566 ( .A1(P2_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n11788), .B1(
        n12671), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n11653) );
  INV_X1 U14567 ( .A(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n11648) );
  NOR2_X1 U14568 ( .A1(n11612), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11644) );
  NAND2_X1 U14569 ( .A1(n9670), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n11647) );
  AND2_X1 U14570 ( .A1(n11612), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11645) );
  NAND2_X1 U14571 ( .A1(n9652), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n11646) );
  OAI211_X1 U14572 ( .C1(n12675), .C2(n11648), .A(n11647), .B(n11646), .ZN(
        n11649) );
  INV_X1 U14573 ( .A(n11649), .ZN(n11652) );
  INV_X1 U14574 ( .A(n11650), .ZN(n13595) );
  NOR2_X1 U14575 ( .A1(n13595), .A2(n11278), .ZN(n12371) );
  AOI22_X1 U14576 ( .A1(n11694), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n13591), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11651) );
  NAND4_X1 U14577 ( .A1(n11654), .A2(n11653), .A3(n11652), .A4(n11651), .ZN(
        n11664) );
  AND2_X1 U14578 ( .A1(n12845), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11834) );
  AOI22_X1 U14579 ( .A1(P2_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n11740), .B1(
        n9623), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11662) );
  AND2_X2 U14580 ( .A1(n11281), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11741) );
  AND2_X1 U14581 ( .A1(n11656), .A2(n11278), .ZN(n11668) );
  AOI22_X1 U14582 ( .A1(P2_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n11741), .B1(
        n11668), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n11661) );
  AND2_X1 U14583 ( .A1(n11657), .A2(n12688), .ZN(n11720) );
  AND2_X1 U14584 ( .A1(n12688), .A2(n11658), .ZN(n11673) );
  AOI22_X1 U14585 ( .A1(P2_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n11720), .B1(
        n11673), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11660) );
  AND2_X1 U14586 ( .A1(n11656), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11742) );
  NAND2_X1 U14587 ( .A1(n11742), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n11659) );
  NAND4_X1 U14588 ( .A1(n11662), .A2(n11661), .A3(n11660), .A4(n11659), .ZN(
        n11663) );
  NAND2_X1 U14589 ( .A1(n11685), .A2(n12399), .ZN(n11667) );
  AND2_X1 U14590 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n11665) );
  NOR2_X1 U14591 ( .A1(n11963), .A2(n11665), .ZN(n11666) );
  NAND3_X1 U14592 ( .A1(n11704), .A2(n11667), .A3(n11666), .ZN(n13039) );
  INV_X1 U14593 ( .A(n12675), .ZN(n11848) );
  INV_X1 U14594 ( .A(n11694), .ZN(n11829) );
  AOI22_X1 U14595 ( .A1(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n11848), .B1(
        n11694), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n11672) );
  AOI22_X1 U14596 ( .A1(P2_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n11834), .B1(
        n11668), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11671) );
  INV_X1 U14597 ( .A(n11687), .ZN(n11754) );
  AOI22_X1 U14598 ( .A1(n11754), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n13591), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11670) );
  AOI22_X1 U14599 ( .A1(P2_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n11740), .B1(
        n11741), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n11669) );
  NAND4_X1 U14600 ( .A1(n11672), .A2(n11671), .A3(n11670), .A4(n11669), .ZN(
        n11679) );
  AOI22_X1 U14601 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n11720), .B1(
        n9670), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11677) );
  AOI22_X1 U14602 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n9652), .B1(
        n11673), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11676) );
  AOI22_X1 U14603 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n11788), .B1(
        n12671), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11675) );
  INV_X1 U14604 ( .A(n11686), .ZN(n11878) );
  AOI22_X1 U14605 ( .A1(n11878), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_14__1__SCAN_IN), .B2(n12662), .ZN(n11674) );
  NAND4_X1 U14606 ( .A1(n11677), .A2(n11676), .A3(n11675), .A4(n11674), .ZN(
        n11678) );
  INV_X1 U14607 ( .A(n11685), .ZN(n11896) );
  OR2_X1 U14608 ( .A1(n12400), .A2(n11896), .ZN(n11682) );
  NOR2_X1 U14609 ( .A1(n11630), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n11680) );
  AOI22_X1 U14610 ( .A1(n11470), .A2(n11680), .B1(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(P2_STATE2_REG_3__SCAN_IN), 
        .ZN(n11681) );
  INV_X1 U14611 ( .A(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n13707) );
  INV_X1 U14612 ( .A(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11688) );
  OAI22_X1 U14613 ( .A1(n13707), .A2(n11686), .B1(n11687), .B2(n11688), .ZN(
        n11689) );
  INV_X1 U14614 ( .A(n11689), .ZN(n11698) );
  AOI22_X1 U14615 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n11788), .B1(
        n12671), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11697) );
  INV_X1 U14616 ( .A(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11692) );
  NAND2_X1 U14617 ( .A1(n9670), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(
        n11691) );
  NAND2_X1 U14618 ( .A1(n9652), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(
        n11690) );
  OAI211_X1 U14619 ( .C1(n12675), .C2(n11692), .A(n11691), .B(n11690), .ZN(
        n11693) );
  INV_X1 U14620 ( .A(n11693), .ZN(n11696) );
  AOI22_X1 U14621 ( .A1(n11694), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n13591), .B2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11695) );
  AOI22_X1 U14622 ( .A1(P2_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n11740), .B1(
        n11834), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11702) );
  AOI22_X1 U14623 ( .A1(P2_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n11741), .B1(
        n11668), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11701) );
  AOI22_X1 U14624 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n11720), .B1(
        n11673), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11700) );
  NAND2_X1 U14625 ( .A1(n12662), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(
        n11699) );
  NAND4_X1 U14626 ( .A1(n11702), .A2(n11701), .A3(n11700), .A4(n11699), .ZN(
        n11703) );
  NAND2_X1 U14627 ( .A1(n11685), .A2(n12404), .ZN(n11705) );
  OAI211_X1 U14628 ( .C1(n19594), .C2(n19764), .A(n11705), .B(n11704), .ZN(
        n11706) );
  AOI21_X2 U14629 ( .B1(n13508), .B2(n11707), .A(n11706), .ZN(n11711) );
  AND3_X1 U14630 ( .A1(n13508), .A2(n11707), .A3(n11706), .ZN(n11708) );
  NAND2_X1 U14631 ( .A1(n11975), .A2(P2_REIP_REG_2__SCAN_IN), .ZN(n11710) );
  INV_X2 U14632 ( .A(n11969), .ZN(n11976) );
  AOI22_X1 U14633 ( .A1(n11963), .A2(P2_EAX_REG_2__SCAN_IN), .B1(n11976), .B2(
        P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n11709) );
  NAND2_X1 U14634 ( .A1(n11710), .A2(n11709), .ZN(n13464) );
  NOR2_X1 U14635 ( .A1(n13465), .A2(n13464), .ZN(n13466) );
  NOR2_X2 U14636 ( .A1(n13466), .A2(n11711), .ZN(n13547) );
  NAND2_X1 U14637 ( .A1(n11975), .A2(P2_REIP_REG_3__SCAN_IN), .ZN(n11731) );
  AOI22_X1 U14638 ( .A1(n11976), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B1(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(P2_STATE2_REG_3__SCAN_IN), 
        .ZN(n11730) );
  NAND2_X1 U14639 ( .A1(n11963), .A2(P2_EAX_REG_3__SCAN_IN), .ZN(n11729) );
  INV_X1 U14640 ( .A(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n12092) );
  INV_X1 U14641 ( .A(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n12084) );
  OAI22_X1 U14642 ( .A1(n12092), .A2(n11687), .B1(n11829), .B2(n12084), .ZN(
        n11712) );
  INV_X1 U14643 ( .A(n11712), .ZN(n11719) );
  AOI22_X1 U14644 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n11788), .B1(
        n11834), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11718) );
  INV_X1 U14645 ( .A(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12078) );
  NAND2_X1 U14646 ( .A1(n9670), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(
        n11714) );
  NAND2_X1 U14647 ( .A1(n9652), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(
        n11713) );
  OAI211_X1 U14648 ( .C1(n11686), .C2(n12078), .A(n11714), .B(n11713), .ZN(
        n11715) );
  INV_X1 U14649 ( .A(n11715), .ZN(n11717) );
  AOI22_X1 U14650 ( .A1(n11848), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n13591), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11716) );
  NAND4_X1 U14651 ( .A1(n11719), .A2(n11718), .A3(n11717), .A4(n11716), .ZN(
        n11727) );
  AOI22_X1 U14652 ( .A1(P2_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n11740), .B1(
        n12671), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11725) );
  AOI22_X1 U14653 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n11668), .B1(
        n12662), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11724) );
  AOI22_X1 U14654 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n11673), .B1(
        n11720), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11723) );
  INV_X1 U14655 ( .A(n11741), .ZN(n11721) );
  OR2_X1 U14656 ( .A1(n11721), .A2(n11253), .ZN(n11722) );
  NAND4_X1 U14657 ( .A1(n11725), .A2(n11724), .A3(n11723), .A4(n11722), .ZN(
        n11726) );
  NAND2_X1 U14658 ( .A1(n11685), .A2(n12099), .ZN(n11728) );
  NAND4_X1 U14659 ( .A1(n11731), .A2(n11730), .A3(n11729), .A4(n11728), .ZN(
        n13548) );
  NAND2_X1 U14660 ( .A1(n13547), .A2(n13548), .ZN(n13479) );
  NAND2_X1 U14661 ( .A1(n11975), .A2(P2_REIP_REG_4__SCAN_IN), .ZN(n11749) );
  AOI22_X1 U14662 ( .A1(n11963), .A2(P2_EAX_REG_4__SCAN_IN), .B1(n11976), .B2(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n11748) );
  INV_X1 U14663 ( .A(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n11732) );
  INV_X1 U14664 ( .A(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n11880) );
  OAI22_X1 U14665 ( .A1(n11732), .A2(n11687), .B1(n11829), .B2(n11880), .ZN(
        n11733) );
  INV_X1 U14666 ( .A(n11733), .ZN(n11739) );
  AOI22_X1 U14667 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n11788), .B1(
        n11834), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11738) );
  INV_X1 U14668 ( .A(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n11734) );
  INV_X1 U14669 ( .A(n11735), .ZN(n11737) );
  AOI22_X1 U14670 ( .A1(n11878), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n13591), .B2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11736) );
  AOI22_X1 U14671 ( .A1(P2_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n11740), .B1(
        n12671), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n11746) );
  AOI22_X1 U14672 ( .A1(P2_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n11741), .B1(
        n12662), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11745) );
  AOI22_X1 U14673 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n11673), .B1(
        n11720), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11744) );
  NAND2_X1 U14674 ( .A1(n11668), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(
        n11743) );
  NAND2_X1 U14675 ( .A1(n11685), .A2(n12102), .ZN(n11747) );
  INV_X1 U14676 ( .A(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12124) );
  INV_X1 U14677 ( .A(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12105) );
  OAI22_X1 U14678 ( .A1(n12124), .A2(n11686), .B1(n11829), .B2(n12105), .ZN(
        n11750) );
  INV_X1 U14679 ( .A(n11750), .ZN(n11758) );
  AOI22_X1 U14680 ( .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n11788), .B1(
        n11834), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11757) );
  INV_X1 U14681 ( .A(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12109) );
  NAND2_X1 U14682 ( .A1(n11720), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(
        n11752) );
  NAND2_X1 U14683 ( .A1(n9670), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(
        n11751) );
  OAI211_X1 U14684 ( .C1(n12675), .C2(n12109), .A(n11752), .B(n11751), .ZN(
        n11753) );
  INV_X1 U14685 ( .A(n11753), .ZN(n11756) );
  AOI22_X1 U14686 ( .A1(n11754), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n13591), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11755) );
  NAND4_X1 U14687 ( .A1(n11758), .A2(n11757), .A3(n11756), .A4(n11755), .ZN(
        n11764) );
  AOI22_X1 U14688 ( .A1(P2_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n11740), .B1(
        n12671), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11762) );
  AOI22_X1 U14689 ( .A1(P2_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n11741), .B1(
        n12662), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11761) );
  AOI22_X1 U14690 ( .A1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n9652), .B1(
        n11673), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11760) );
  NAND2_X1 U14691 ( .A1(n11668), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(
        n11759) );
  NAND4_X1 U14692 ( .A1(n11762), .A2(n11761), .A3(n11760), .A4(n11759), .ZN(
        n11763) );
  NAND2_X1 U14693 ( .A1(n12141), .A2(n12003), .ZN(n11995) );
  INV_X1 U14694 ( .A(n11995), .ZN(n11765) );
  AOI22_X1 U14695 ( .A1(n12437), .A2(P2_REIP_REG_5__SCAN_IN), .B1(n11765), 
        .B2(n13044), .ZN(n11767) );
  AOI22_X1 U14696 ( .A1(n11963), .A2(P2_EAX_REG_5__SCAN_IN), .B1(n11976), .B2(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n11766) );
  NAND2_X1 U14697 ( .A1(n11767), .A2(n11766), .ZN(n13676) );
  NAND2_X1 U14698 ( .A1(n13480), .A2(n13676), .ZN(n13675) );
  INV_X1 U14699 ( .A(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12182) );
  INV_X1 U14700 ( .A(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12181) );
  OAI22_X1 U14701 ( .A1(n12182), .A2(n11686), .B1(n11687), .B2(n12181), .ZN(
        n11768) );
  INV_X1 U14702 ( .A(n11768), .ZN(n11775) );
  AOI22_X1 U14703 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n11788), .B1(
        n12671), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11774) );
  INV_X1 U14704 ( .A(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12179) );
  NAND2_X1 U14705 ( .A1(n9670), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(
        n11770) );
  NAND2_X1 U14706 ( .A1(n9652), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(
        n11769) );
  OAI211_X1 U14707 ( .C1(n12675), .C2(n12179), .A(n11770), .B(n11769), .ZN(
        n11771) );
  INV_X1 U14708 ( .A(n11771), .ZN(n11773) );
  AOI22_X1 U14709 ( .A1(n11694), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n13591), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11772) );
  NAND4_X1 U14710 ( .A1(n11775), .A2(n11774), .A3(n11773), .A4(n11772), .ZN(
        n11781) );
  AOI22_X1 U14711 ( .A1(P2_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n11740), .B1(
        n11834), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11779) );
  AOI22_X1 U14712 ( .A1(P2_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n11741), .B1(
        n11668), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11778) );
  AOI22_X1 U14713 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n11673), .B1(
        n11720), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11777) );
  NAND2_X1 U14714 ( .A1(n12662), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(
        n11776) );
  NAND4_X1 U14715 ( .A1(n11779), .A2(n11778), .A3(n11777), .A4(n11776), .ZN(
        n11780) );
  NAND2_X1 U14716 ( .A1(n11685), .A2(n12193), .ZN(n11782) );
  NAND2_X1 U14717 ( .A1(n11975), .A2(P2_REIP_REG_6__SCAN_IN), .ZN(n11784) );
  AOI22_X1 U14718 ( .A1(n11963), .A2(P2_EAX_REG_6__SCAN_IN), .B1(n11976), .B2(
        P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n11783) );
  NAND2_X1 U14719 ( .A1(n11784), .A2(n11783), .ZN(n14048) );
  NAND2_X1 U14720 ( .A1(n14047), .A2(n14048), .ZN(n11803) );
  INV_X1 U14721 ( .A(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n11786) );
  INV_X1 U14722 ( .A(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n11785) );
  OAI22_X1 U14723 ( .A1(n11786), .A2(n11686), .B1(n11687), .B2(n11785), .ZN(
        n11787) );
  INV_X1 U14724 ( .A(n11787), .ZN(n11795) );
  AOI22_X1 U14725 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n11788), .B1(
        n12671), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n11794) );
  INV_X1 U14726 ( .A(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n20809) );
  NAND2_X1 U14727 ( .A1(n9670), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(
        n11790) );
  NAND2_X1 U14728 ( .A1(n9652), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(
        n11789) );
  OAI211_X1 U14729 ( .C1(n12675), .C2(n20809), .A(n11790), .B(n11789), .ZN(
        n11791) );
  INV_X1 U14730 ( .A(n11791), .ZN(n11793) );
  AOI22_X1 U14731 ( .A1(n11694), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n13591), .B2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11792) );
  NAND4_X1 U14732 ( .A1(n11795), .A2(n11794), .A3(n11793), .A4(n11792), .ZN(
        n11801) );
  AOI22_X1 U14733 ( .A1(P2_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n11740), .B1(
        n11834), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11799) );
  AOI22_X1 U14734 ( .A1(P2_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n11741), .B1(
        n11668), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n11798) );
  AOI22_X1 U14735 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n11673), .B1(
        n11720), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11797) );
  NAND2_X1 U14736 ( .A1(n12662), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n11796) );
  NAND4_X1 U14737 ( .A1(n11799), .A2(n11798), .A3(n11797), .A4(n11796), .ZN(
        n11800) );
  NAND2_X1 U14738 ( .A1(n11685), .A2(n12322), .ZN(n11802) );
  NAND2_X1 U14739 ( .A1(n11975), .A2(P2_REIP_REG_7__SCAN_IN), .ZN(n11805) );
  AOI22_X1 U14740 ( .A1(n11963), .A2(P2_EAX_REG_7__SCAN_IN), .B1(n11976), .B2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n11804) );
  NAND2_X1 U14741 ( .A1(n11805), .A2(n11804), .ZN(n13824) );
  NAND2_X1 U14742 ( .A1(n11975), .A2(P2_REIP_REG_8__SCAN_IN), .ZN(n11824) );
  AOI22_X1 U14743 ( .A1(n11963), .A2(P2_EAX_REG_8__SCAN_IN), .B1(n11976), .B2(
        P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n11823) );
  INV_X1 U14744 ( .A(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n11806) );
  INV_X1 U14745 ( .A(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n19568) );
  OAI22_X1 U14746 ( .A1(n11806), .A2(n11686), .B1(n11687), .B2(n19568), .ZN(
        n11807) );
  INV_X1 U14747 ( .A(n11807), .ZN(n11815) );
  AOI22_X1 U14748 ( .A1(P2_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n11788), .B1(
        n12671), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n11814) );
  INV_X1 U14749 ( .A(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n11810) );
  NAND2_X1 U14750 ( .A1(n11720), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n11809) );
  NAND2_X1 U14751 ( .A1(n9670), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(
        n11808) );
  OAI211_X1 U14752 ( .C1(n12675), .C2(n11810), .A(n11809), .B(n11808), .ZN(
        n11811) );
  INV_X1 U14753 ( .A(n11811), .ZN(n11813) );
  AOI22_X1 U14754 ( .A1(n11694), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n13591), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11812) );
  NAND4_X1 U14755 ( .A1(n11815), .A2(n11814), .A3(n11813), .A4(n11812), .ZN(
        n11821) );
  AOI22_X1 U14756 ( .A1(P2_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n9623), .B1(
        n11740), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n11819) );
  AOI22_X1 U14757 ( .A1(P2_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n11741), .B1(
        n11668), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n11818) );
  AOI22_X1 U14758 ( .A1(P2_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n11673), .B1(
        n9652), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11817) );
  NAND2_X1 U14759 ( .A1(n12662), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n11816) );
  NAND4_X1 U14760 ( .A1(n11819), .A2(n11818), .A3(n11817), .A4(n11816), .ZN(
        n11820) );
  OR2_X1 U14761 ( .A1(n11821), .A2(n11820), .ZN(n13237) );
  NAND2_X1 U14762 ( .A1(n11685), .A2(n13237), .ZN(n11822) );
  INV_X1 U14763 ( .A(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n12038) );
  INV_X1 U14764 ( .A(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12046) );
  OAI22_X1 U14765 ( .A1(n12038), .A2(n11686), .B1(n11687), .B2(n12046), .ZN(
        n11825) );
  INV_X1 U14766 ( .A(n11825), .ZN(n11833) );
  AOI22_X1 U14767 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n11788), .B1(
        n12671), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n11832) );
  INV_X1 U14768 ( .A(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12037) );
  NAND2_X1 U14769 ( .A1(n9670), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n11827) );
  NAND2_X1 U14770 ( .A1(n9652), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n11826) );
  OAI211_X1 U14771 ( .C1(n12675), .C2(n12037), .A(n11827), .B(n11826), .ZN(
        n11828) );
  INV_X1 U14772 ( .A(n11828), .ZN(n11831) );
  AOI22_X1 U14773 ( .A1(n11694), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n13591), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11830) );
  NAND4_X1 U14774 ( .A1(n11833), .A2(n11832), .A3(n11831), .A4(n11830), .ZN(
        n11840) );
  AOI22_X1 U14775 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n11834), .B1(
        n11740), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11838) );
  AOI22_X1 U14776 ( .A1(P2_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n11741), .B1(
        n11668), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11837) );
  AOI22_X1 U14777 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n11673), .B1(
        n11720), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11836) );
  NAND2_X1 U14778 ( .A1(n12662), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n11835) );
  NAND4_X1 U14779 ( .A1(n11838), .A2(n11837), .A3(n11836), .A4(n11835), .ZN(
        n11839) );
  OR2_X1 U14780 ( .A1(n11840), .A2(n11839), .ZN(n18949) );
  AOI22_X1 U14781 ( .A1(n12437), .A2(P2_REIP_REG_9__SCAN_IN), .B1(n11685), 
        .B2(n18949), .ZN(n11842) );
  AOI22_X1 U14782 ( .A1(n11963), .A2(P2_EAX_REG_9__SCAN_IN), .B1(n11976), .B2(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n11841) );
  NAND2_X1 U14783 ( .A1(n11842), .A2(n11841), .ZN(n13532) );
  NAND2_X1 U14784 ( .A1(n11975), .A2(P2_REIP_REG_10__SCAN_IN), .ZN(n11861) );
  AOI22_X1 U14785 ( .A1(n11963), .A2(P2_EAX_REG_10__SCAN_IN), .B1(n11976), 
        .B2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n11860) );
  INV_X1 U14786 ( .A(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11844) );
  INV_X1 U14787 ( .A(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11843) );
  OAI22_X1 U14788 ( .A1(n11844), .A2(n11686), .B1(n11687), .B2(n11843), .ZN(
        n11845) );
  INV_X1 U14789 ( .A(n11845), .ZN(n11852) );
  AOI22_X1 U14790 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n9670), .B1(n9652), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11847) );
  NAND2_X1 U14791 ( .A1(n11694), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(
        n11846) );
  AND2_X1 U14792 ( .A1(n11847), .A2(n11846), .ZN(n11851) );
  AOI22_X1 U14793 ( .A1(n11848), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n13591), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11850) );
  AOI22_X1 U14794 ( .A1(P2_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n9623), .B1(
        n11788), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11849) );
  NAND4_X1 U14795 ( .A1(n11852), .A2(n11851), .A3(n11850), .A4(n11849), .ZN(
        n11858) );
  AOI22_X1 U14796 ( .A1(P2_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n11740), .B1(
        n12671), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11856) );
  AOI22_X1 U14797 ( .A1(P2_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n11741), .B1(
        n11742), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11855) );
  AOI22_X1 U14798 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n11720), .B1(
        n11673), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11854) );
  NAND2_X1 U14799 ( .A1(n11668), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(
        n11853) );
  NAND4_X1 U14800 ( .A1(n11856), .A2(n11855), .A3(n11854), .A4(n11853), .ZN(
        n11857) );
  OR2_X1 U14801 ( .A1(n11858), .A2(n11857), .ZN(n18948) );
  NAND2_X1 U14802 ( .A1(n11685), .A2(n18948), .ZN(n11859) );
  NOR2_X2 U14803 ( .A1(n15004), .A2(n15003), .ZN(n14984) );
  AOI22_X1 U14804 ( .A1(n12437), .A2(P2_REIP_REG_11__SCAN_IN), .B1(n11963), 
        .B2(P2_EAX_REG_11__SCAN_IN), .ZN(n11877) );
  INV_X1 U14805 ( .A(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12087) );
  INV_X1 U14806 ( .A(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12090) );
  OAI22_X1 U14807 ( .A1(n12087), .A2(n11686), .B1(n11687), .B2(n12090), .ZN(
        n11862) );
  INV_X1 U14808 ( .A(n11862), .ZN(n11869) );
  AOI22_X1 U14809 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n11788), .B1(
        n12671), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n11868) );
  NAND2_X1 U14810 ( .A1(n9670), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(
        n11864) );
  NAND2_X1 U14811 ( .A1(n9652), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(
        n11863) );
  OAI211_X1 U14812 ( .C1(n12675), .C2(n12084), .A(n11864), .B(n11863), .ZN(
        n11865) );
  INV_X1 U14813 ( .A(n11865), .ZN(n11867) );
  AOI22_X1 U14814 ( .A1(n11694), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n13591), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11866) );
  NAND4_X1 U14815 ( .A1(n11869), .A2(n11868), .A3(n11867), .A4(n11866), .ZN(
        n11875) );
  AOI22_X1 U14816 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n11834), .B1(
        n11740), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11873) );
  AOI22_X1 U14817 ( .A1(P2_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n11741), .B1(
        n11668), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11872) );
  AOI22_X1 U14818 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n11673), .B1(
        n11720), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11871) );
  NAND2_X1 U14819 ( .A1(n12662), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(
        n11870) );
  NAND4_X1 U14820 ( .A1(n11873), .A2(n11872), .A3(n11871), .A4(n11870), .ZN(
        n11874) );
  OR2_X1 U14821 ( .A1(n11875), .A2(n11874), .ZN(n13366) );
  AOI22_X1 U14822 ( .A1(n11685), .A2(n13366), .B1(
        P2_INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n11976), .ZN(n11876) );
  NAND2_X1 U14823 ( .A1(n11877), .A2(n11876), .ZN(n14983) );
  NAND2_X1 U14824 ( .A1(n14984), .A2(n14983), .ZN(n14982) );
  AOI22_X1 U14825 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n11878), .B1(
        n11694), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n11888) );
  INV_X1 U14826 ( .A(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11879) );
  OAI22_X1 U14827 ( .A1(n11880), .A2(n12675), .B1(n11687), .B2(n11879), .ZN(
        n11881) );
  INV_X1 U14828 ( .A(n11881), .ZN(n11887) );
  NAND2_X1 U14829 ( .A1(n13591), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n11884) );
  NAND2_X1 U14830 ( .A1(n11720), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n11883) );
  NAND2_X1 U14831 ( .A1(n9670), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(
        n11882) );
  AND3_X1 U14832 ( .A1(n11884), .A2(n11883), .A3(n11882), .ZN(n11886) );
  AOI22_X1 U14833 ( .A1(P2_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n11740), .B1(
        n12671), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n11885) );
  NAND4_X1 U14834 ( .A1(n11888), .A2(n11887), .A3(n11886), .A4(n11885), .ZN(
        n11894) );
  AOI22_X1 U14835 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n9623), .B1(
        n11788), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n11892) );
  AOI22_X1 U14836 ( .A1(P2_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n11741), .B1(
        n12662), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11891) );
  AOI22_X1 U14837 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n11673), .B1(
        n9652), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11890) );
  NAND2_X1 U14838 ( .A1(n11668), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(
        n11889) );
  NAND4_X1 U14839 ( .A1(n11892), .A2(n11891), .A3(n11890), .A4(n11889), .ZN(
        n11893) );
  OR2_X1 U14840 ( .A1(n11894), .A2(n11893), .ZN(n12543) );
  INV_X1 U14841 ( .A(n12543), .ZN(n13367) );
  AOI22_X1 U14842 ( .A1(n11963), .A2(P2_EAX_REG_12__SCAN_IN), .B1(n11976), 
        .B2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n11895) );
  OAI21_X1 U14843 ( .B1(n11896), .B2(n13367), .A(n11895), .ZN(n11897) );
  AOI21_X1 U14844 ( .B1(n11975), .B2(P2_REIP_REG_12__SCAN_IN), .A(n11897), 
        .ZN(n16102) );
  NOR2_X4 U14845 ( .A1(n14982), .A2(n16102), .ZN(n16101) );
  AOI22_X1 U14846 ( .A1(n12437), .A2(P2_REIP_REG_13__SCAN_IN), .B1(n11963), 
        .B2(P2_EAX_REG_13__SCAN_IN), .ZN(n11913) );
  INV_X1 U14847 ( .A(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12110) );
  INV_X1 U14848 ( .A(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12115) );
  OAI22_X1 U14849 ( .A1(n12110), .A2(n11686), .B1(n11687), .B2(n12115), .ZN(
        n11898) );
  INV_X1 U14850 ( .A(n11898), .ZN(n11905) );
  AOI22_X1 U14851 ( .A1(P2_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n11788), .B1(
        n12671), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n11904) );
  NAND2_X1 U14852 ( .A1(n9670), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(
        n11900) );
  NAND2_X1 U14853 ( .A1(n9652), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(
        n11899) );
  OAI211_X1 U14854 ( .C1(n12675), .C2(n12105), .A(n11900), .B(n11899), .ZN(
        n11901) );
  INV_X1 U14855 ( .A(n11901), .ZN(n11903) );
  AOI22_X1 U14856 ( .A1(n11694), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n13591), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11902) );
  NAND4_X1 U14857 ( .A1(n11905), .A2(n11904), .A3(n11903), .A4(n11902), .ZN(
        n11911) );
  INV_X1 U14858 ( .A(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n19171) );
  AOI22_X1 U14859 ( .A1(P2_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n11740), .B1(
        n11834), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11909) );
  AOI22_X1 U14860 ( .A1(P2_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n11741), .B1(
        n11668), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11908) );
  AOI22_X1 U14861 ( .A1(P2_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n11673), .B1(
        n11720), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11907) );
  NAND2_X1 U14862 ( .A1(n11742), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(
        n11906) );
  NAND4_X1 U14863 ( .A1(n11909), .A2(n11908), .A3(n11907), .A4(n11906), .ZN(
        n11910) );
  OR2_X1 U14864 ( .A1(n11911), .A2(n11910), .ZN(n14169) );
  AOI22_X1 U14865 ( .A1(n11685), .A2(n14169), .B1(
        P2_INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n11976), .ZN(n11912) );
  NAND2_X1 U14866 ( .A1(n11913), .A2(n11912), .ZN(n14966) );
  NAND2_X1 U14867 ( .A1(n11975), .A2(P2_REIP_REG_14__SCAN_IN), .ZN(n11930) );
  AOI22_X1 U14868 ( .A1(n11963), .A2(P2_EAX_REG_14__SCAN_IN), .B1(n11976), 
        .B2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n11929) );
  INV_X1 U14869 ( .A(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12170) );
  INV_X1 U14870 ( .A(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12172) );
  OAI22_X1 U14871 ( .A1(n12170), .A2(n11686), .B1(n11687), .B2(n12172), .ZN(
        n11914) );
  INV_X1 U14872 ( .A(n11914), .ZN(n11921) );
  AOI22_X1 U14873 ( .A1(P2_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n11740), .B1(
        n11788), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11920) );
  INV_X1 U14874 ( .A(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12180) );
  NAND2_X1 U14875 ( .A1(n9670), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(
        n11916) );
  NAND2_X1 U14876 ( .A1(n9652), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(
        n11915) );
  OAI211_X1 U14877 ( .C1(n12675), .C2(n12180), .A(n11916), .B(n11915), .ZN(
        n11917) );
  INV_X1 U14878 ( .A(n11917), .ZN(n11919) );
  AOI22_X1 U14879 ( .A1(n11694), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n13591), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11918) );
  NAND4_X1 U14880 ( .A1(n11921), .A2(n11920), .A3(n11919), .A4(n11918), .ZN(
        n11927) );
  AOI22_X1 U14881 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n11834), .B1(
        n12671), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n11925) );
  AOI22_X1 U14882 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n11668), .B1(
        n12662), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11924) );
  AOI22_X1 U14883 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n11673), .B1(
        n11720), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11923) );
  NAND2_X1 U14884 ( .A1(n11741), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(
        n11922) );
  NAND4_X1 U14885 ( .A1(n11925), .A2(n11924), .A3(n11923), .A4(n11922), .ZN(
        n11926) );
  OR2_X1 U14886 ( .A1(n11927), .A2(n11926), .ZN(n13517) );
  NAND2_X1 U14887 ( .A1(n11685), .A2(n13517), .ZN(n11928) );
  INV_X1 U14888 ( .A(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n20836) );
  INV_X1 U14889 ( .A(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11931) );
  OAI22_X1 U14890 ( .A1(n20836), .A2(n11686), .B1(n11687), .B2(n11931), .ZN(
        n11932) );
  INV_X1 U14891 ( .A(n11932), .ZN(n11940) );
  AOI22_X1 U14892 ( .A1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n11788), .B1(
        n12671), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n11939) );
  INV_X1 U14893 ( .A(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n11935) );
  NAND2_X1 U14894 ( .A1(n9670), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(
        n11934) );
  NAND2_X1 U14895 ( .A1(n9652), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(
        n11933) );
  OAI211_X1 U14896 ( .C1(n12675), .C2(n11935), .A(n11934), .B(n11933), .ZN(
        n11936) );
  INV_X1 U14897 ( .A(n11936), .ZN(n11938) );
  AOI22_X1 U14898 ( .A1(n11694), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n13591), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11937) );
  NAND4_X1 U14899 ( .A1(n11940), .A2(n11939), .A3(n11938), .A4(n11937), .ZN(
        n11946) );
  AOI22_X1 U14900 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n9623), .B1(
        n11740), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n11944) );
  AOI22_X1 U14901 ( .A1(P2_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n11741), .B1(
        n11668), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n11943) );
  AOI22_X1 U14902 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n11673), .B1(
        n11720), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11942) );
  NAND2_X1 U14903 ( .A1(n12662), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(
        n11941) );
  NAND4_X1 U14904 ( .A1(n11944), .A2(n11943), .A3(n11942), .A4(n11941), .ZN(
        n11945) );
  OR2_X1 U14905 ( .A1(n11946), .A2(n11945), .ZN(n13719) );
  AOI22_X1 U14906 ( .A1(n12437), .A2(P2_REIP_REG_15__SCAN_IN), .B1(n11685), 
        .B2(n13719), .ZN(n11948) );
  AOI22_X1 U14907 ( .A1(n11963), .A2(P2_EAX_REG_15__SCAN_IN), .B1(n11976), 
        .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n11947) );
  NAND2_X1 U14908 ( .A1(n11948), .A2(n11947), .ZN(n16074) );
  NAND2_X1 U14909 ( .A1(n12437), .A2(P2_REIP_REG_16__SCAN_IN), .ZN(n11950) );
  AOI22_X1 U14910 ( .A1(n11963), .A2(P2_EAX_REG_16__SCAN_IN), .B1(n11976), 
        .B2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n11949) );
  NAND2_X1 U14911 ( .A1(n11950), .A2(n11949), .ZN(n15286) );
  NAND2_X1 U14912 ( .A1(n11975), .A2(P2_REIP_REG_17__SCAN_IN), .ZN(n11953) );
  AOI22_X1 U14913 ( .A1(n11963), .A2(P2_EAX_REG_17__SCAN_IN), .B1(n11976), 
        .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n11952) );
  AOI222_X1 U14914 ( .A1(n12437), .A2(P2_REIP_REG_18__SCAN_IN), .B1(
        P2_INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n11976), .C1(n11963), .C2(
        P2_EAX_REG_18__SCAN_IN), .ZN(n13735) );
  NAND2_X1 U14915 ( .A1(n12437), .A2(P2_REIP_REG_19__SCAN_IN), .ZN(n11956) );
  AOI22_X1 U14916 ( .A1(n11963), .A2(P2_EAX_REG_19__SCAN_IN), .B1(n11976), 
        .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n11955) );
  NAND2_X1 U14917 ( .A1(n11956), .A2(n11955), .ZN(n13843) );
  NAND2_X1 U14918 ( .A1(n12437), .A2(P2_REIP_REG_20__SCAN_IN), .ZN(n11958) );
  AOI22_X1 U14919 ( .A1(n11963), .A2(P2_EAX_REG_20__SCAN_IN), .B1(n11976), 
        .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n11957) );
  AND2_X1 U14920 ( .A1(n11958), .A2(n11957), .ZN(n15438) );
  NAND2_X1 U14921 ( .A1(n12437), .A2(P2_REIP_REG_21__SCAN_IN), .ZN(n11960) );
  AOI22_X1 U14922 ( .A1(n11963), .A2(P2_EAX_REG_21__SCAN_IN), .B1(n11976), 
        .B2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n11959) );
  NAND2_X1 U14923 ( .A1(n11960), .A2(n11959), .ZN(n14078) );
  NAND2_X1 U14924 ( .A1(n12437), .A2(P2_REIP_REG_22__SCAN_IN), .ZN(n11962) );
  AOI22_X1 U14925 ( .A1(n11963), .A2(P2_EAX_REG_22__SCAN_IN), .B1(n11976), 
        .B2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n11961) );
  NAND2_X1 U14926 ( .A1(n11962), .A2(n11961), .ZN(n14913) );
  INV_X1 U14927 ( .A(n11963), .ZN(n11970) );
  INV_X1 U14928 ( .A(P2_EAX_REG_23__SCAN_IN), .ZN(n14690) );
  INV_X1 U14929 ( .A(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n14897) );
  OAI22_X1 U14930 ( .A1(n11970), .A2(n14690), .B1(n11969), .B2(n14897), .ZN(
        n11964) );
  AOI21_X1 U14931 ( .B1(n12437), .B2(P2_REIP_REG_23__SCAN_IN), .A(n11964), 
        .ZN(n12981) );
  INV_X1 U14932 ( .A(P2_EAX_REG_24__SCAN_IN), .ZN(n14680) );
  INV_X1 U14933 ( .A(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n14873) );
  OAI22_X1 U14934 ( .A1(n11970), .A2(n14680), .B1(n11969), .B2(n14873), .ZN(
        n11965) );
  AOI21_X1 U14935 ( .B1(n12437), .B2(P2_REIP_REG_24__SCAN_IN), .A(n11965), 
        .ZN(n14676) );
  AOI22_X1 U14936 ( .A1(n11963), .A2(P2_EAX_REG_25__SCAN_IN), .B1(n11976), 
        .B2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n11966) );
  OAI21_X1 U14937 ( .B1(n11974), .B2(n19724), .A(n11966), .ZN(n14584) );
  INV_X1 U14938 ( .A(P2_EAX_REG_26__SCAN_IN), .ZN(n14664) );
  OAI22_X1 U14939 ( .A1(n11970), .A2(n14664), .B1(n11969), .B2(n11967), .ZN(
        n11968) );
  AOI21_X1 U14940 ( .B1(n11975), .B2(P2_REIP_REG_26__SCAN_IN), .A(n11968), 
        .ZN(n14661) );
  INV_X1 U14941 ( .A(P2_EAX_REG_27__SCAN_IN), .ZN(n14655) );
  OAI22_X1 U14942 ( .A1(n11970), .A2(n14655), .B1(n11969), .B2(n14707), .ZN(
        n11971) );
  AOI21_X1 U14943 ( .B1(n12437), .B2(P2_REIP_REG_27__SCAN_IN), .A(n11971), 
        .ZN(n14654) );
  AOI22_X1 U14944 ( .A1(n11963), .A2(P2_EAX_REG_28__SCAN_IN), .B1(n11976), 
        .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n11972) );
  OAI21_X1 U14945 ( .B1(n11974), .B2(n19729), .A(n11972), .ZN(n12949) );
  AOI22_X1 U14946 ( .A1(n11963), .A2(P2_EAX_REG_29__SCAN_IN), .B1(n11976), 
        .B2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n11973) );
  OAI21_X1 U14947 ( .B1(n11974), .B2(n19731), .A(n11973), .ZN(n14572) );
  NAND2_X1 U14948 ( .A1(n11975), .A2(P2_REIP_REG_30__SCAN_IN), .ZN(n11978) );
  AOI22_X1 U14949 ( .A1(n11963), .A2(P2_EAX_REG_30__SCAN_IN), .B1(n11976), 
        .B2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n11977) );
  AND2_X1 U14950 ( .A1(n11978), .A2(n11977), .ZN(n11979) );
  OR2_X2 U14951 ( .A1(n14571), .A2(n11979), .ZN(n12441) );
  NAND2_X1 U14952 ( .A1(n14571), .A2(n11979), .ZN(n11980) );
  INV_X1 U14953 ( .A(n14806), .ZN(n11981) );
  OAI22_X1 U14954 ( .A1(n14809), .A2(n18924), .B1(n18928), .B2(n11981), .ZN(
        n11982) );
  INV_X1 U14955 ( .A(n11982), .ZN(n12011) );
  NOR2_X1 U14956 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n15042) );
  NOR2_X1 U14957 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n11983) );
  NAND2_X1 U14958 ( .A1(n15042), .A2(n11983), .ZN(n12482) );
  INV_X1 U14959 ( .A(n19081), .ZN(n16114) );
  NOR3_X1 U14960 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n19658), .A3(n19594), 
        .ZN(n16145) );
  INV_X1 U14961 ( .A(n18890), .ZN(n18920) );
  NOR2_X1 U14962 ( .A1(n16145), .A2(n18920), .ZN(n11984) );
  NAND2_X1 U14963 ( .A1(n16114), .A2(n11984), .ZN(n11985) );
  NOR2_X2 U14964 ( .A1(n18910), .A2(n19594), .ZN(n18892) );
  INV_X1 U14965 ( .A(P2_REIP_REG_30__SCAN_IN), .ZN(n12008) );
  INV_X1 U14966 ( .A(P2_EBX_REG_31__SCAN_IN), .ZN(n12476) );
  INV_X1 U14967 ( .A(P2_STATEBS16_REG_SCAN_IN), .ZN(n19221) );
  AND2_X1 U14968 ( .A1(n19221), .A2(n15424), .ZN(n11986) );
  NAND2_X1 U14969 ( .A1(n11989), .A2(n11988), .ZN(n11990) );
  MUX2_X1 U14970 ( .A(n12400), .B(n11990), .S(n12327), .Z(n12158) );
  INV_X1 U14971 ( .A(n12336), .ZN(n12339) );
  NAND2_X1 U14972 ( .A1(n11991), .A2(n12339), .ZN(n12337) );
  INV_X1 U14973 ( .A(P2_EBX_REG_2__SCAN_IN), .ZN(n11992) );
  MUX2_X1 U14974 ( .A(n12360), .B(n11992), .S(n12327), .Z(n12157) );
  INV_X1 U14975 ( .A(n12157), .ZN(n11993) );
  INV_X1 U14976 ( .A(n12346), .ZN(n11994) );
  MUX2_X1 U14977 ( .A(n12099), .B(n11994), .S(n11991), .Z(n12334) );
  MUX2_X1 U14978 ( .A(n13551), .B(n12334), .S(n12003), .Z(n12152) );
  MUX2_X1 U14979 ( .A(P2_EBX_REG_4__SCAN_IN), .B(n12333), .S(n12003), .Z(
        n12166) );
  OAI21_X1 U14980 ( .B1(n12003), .B2(P2_EBX_REG_5__SCAN_IN), .A(n11995), .ZN(
        n12146) );
  MUX2_X1 U14981 ( .A(n18894), .B(n12193), .S(n12003), .Z(n12203) );
  MUX2_X1 U14982 ( .A(n11533), .B(n12322), .S(n12003), .Z(n12211) );
  NAND2_X1 U14983 ( .A1(n12327), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n12231) );
  NAND2_X1 U14984 ( .A1(n18808), .A2(n11421), .ZN(n11997) );
  NAND2_X1 U14985 ( .A1(n12327), .A2(n11997), .ZN(n11998) );
  NAND2_X1 U14986 ( .A1(n12327), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n12260) );
  INV_X1 U14987 ( .A(P2_EBX_REG_18__SCAN_IN), .ZN(n11999) );
  INV_X1 U14988 ( .A(P2_EBX_REG_19__SCAN_IN), .ZN(n14062) );
  NAND2_X1 U14989 ( .A1(n11999), .A2(n14062), .ZN(n12000) );
  AND2_X1 U14990 ( .A1(n12327), .A2(n12000), .ZN(n12001) );
  INV_X1 U14991 ( .A(P2_EBX_REG_21__SCAN_IN), .ZN(n14637) );
  NAND2_X1 U14992 ( .A1(n12327), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n12282) );
  AND2_X1 U14993 ( .A1(n12327), .A2(P2_EBX_REG_23__SCAN_IN), .ZN(n12288) );
  NAND2_X1 U14994 ( .A1(n12301), .A2(n12310), .ZN(n12305) );
  NAND2_X1 U14995 ( .A1(n12327), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n12309) );
  INV_X1 U14996 ( .A(P2_EBX_REG_28__SCAN_IN), .ZN(n15887) );
  NOR2_X1 U14997 ( .A1(n12003), .A2(n15887), .ZN(n12307) );
  NAND2_X1 U14998 ( .A1(n12327), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n12318) );
  NAND2_X1 U14999 ( .A1(n12319), .A2(n12318), .ZN(n12326) );
  NAND2_X1 U15000 ( .A1(n12327), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n12004) );
  XNOR2_X1 U15001 ( .A(n12326), .B(n12004), .ZN(n12320) );
  INV_X1 U15002 ( .A(n12320), .ZN(n12321) );
  NOR2_X1 U15003 ( .A1(n12988), .A2(n11458), .ZN(n13025) );
  OAI21_X1 U15004 ( .B1(P2_STATEBS16_REG_SCAN_IN), .B2(n19807), .A(n12476), 
        .ZN(n12005) );
  AOI21_X1 U15005 ( .B1(n19796), .B2(n12005), .A(n13652), .ZN(n12006) );
  NAND2_X1 U15006 ( .A1(n13025), .A2(n12006), .ZN(n18929) );
  OAI222_X1 U15007 ( .A1(n18932), .A2(n12008), .B1(n18923), .B2(n12321), .C1(
        n12007), .C2(n18929), .ZN(n12009) );
  AOI21_X1 U15008 ( .B1(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n18892), .A(
        n12009), .ZN(n12010) );
  INV_X1 U15009 ( .A(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n20908) );
  XNOR2_X2 U15010 ( .A(n12014), .B(n12013), .ZN(n13079) );
  INV_X1 U15011 ( .A(n12018), .ZN(n12020) );
  INV_X1 U15012 ( .A(n12027), .ZN(n12019) );
  NAND2_X1 U15013 ( .A1(n12020), .A2(n12019), .ZN(n12021) );
  INV_X1 U15014 ( .A(n12022), .ZN(n12025) );
  INV_X1 U15015 ( .A(n12023), .ZN(n12024) );
  NAND2_X1 U15016 ( .A1(n12025), .A2(n12024), .ZN(n12026) );
  NAND2_X1 U15017 ( .A1(n19130), .A2(n18925), .ZN(n12043) );
  OR2_X2 U15018 ( .A1(n12056), .A2(n12043), .ZN(n12104) );
  INV_X1 U15019 ( .A(n18925), .ZN(n16141) );
  OR2_X2 U15020 ( .A1(n12053), .A2(n12055), .ZN(n12131) );
  INV_X1 U15021 ( .A(n12131), .ZN(n12028) );
  NAND2_X1 U15022 ( .A1(n12028), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n12029) );
  OAI211_X1 U15023 ( .C1(n20908), .C2(n12104), .A(n12029), .B(n19796), .ZN(
        n12036) );
  INV_X1 U15024 ( .A(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n12034) );
  INV_X1 U15025 ( .A(n12056), .ZN(n12031) );
  OR2_X1 U15026 ( .A1(n12018), .A2(n18925), .ZN(n12052) );
  INV_X1 U15027 ( .A(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n12033) );
  OAI22_X1 U15028 ( .A1(n12034), .A2(n12129), .B1(n12132), .B2(n12033), .ZN(
        n12035) );
  OR2_X2 U15029 ( .A1(n12053), .A2(n12043), .ZN(n12107) );
  OAI22_X1 U15030 ( .A1(n12038), .A2(n12107), .B1(n19425), .B2(n12037), .ZN(
        n12042) );
  INV_X1 U15031 ( .A(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n12040) );
  NAND2_X1 U15032 ( .A1(n9650), .A2(n12519), .ZN(n12047) );
  OR2_X2 U15033 ( .A1(n12047), .A2(n12055), .ZN(n12113) );
  INV_X1 U15034 ( .A(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n12039) );
  OAI22_X1 U15035 ( .A1(n12040), .A2(n12113), .B1(n12108), .B2(n12039), .ZN(
        n12041) );
  NOR2_X1 U15036 ( .A1(n12042), .A2(n12041), .ZN(n12066) );
  INV_X1 U15037 ( .A(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12568) );
  NAND2_X1 U15038 ( .A1(n16141), .A2(n12018), .ZN(n12058) );
  INV_X1 U15039 ( .A(n12047), .ZN(n12045) );
  OAI22_X1 U15040 ( .A1(n12568), .A2(n9673), .B1(n12114), .B2(n12046), .ZN(
        n12051) );
  INV_X1 U15041 ( .A(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12049) );
  INV_X1 U15042 ( .A(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n12048) );
  NOR2_X1 U15043 ( .A1(n12051), .A2(n12050), .ZN(n12065) );
  INV_X1 U15044 ( .A(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12054) );
  OR2_X2 U15045 ( .A1(n12053), .A2(n12052), .ZN(n12121) );
  INV_X1 U15046 ( .A(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n12569) );
  OAI22_X1 U15047 ( .A1(n12054), .A2(n12121), .B1(n19339), .B2(n12569), .ZN(
        n12063) );
  INV_X1 U15048 ( .A(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n12061) );
  INV_X1 U15049 ( .A(n12057), .ZN(n12060) );
  INV_X1 U15050 ( .A(n12058), .ZN(n12059) );
  INV_X1 U15051 ( .A(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n12573) );
  OAI22_X1 U15052 ( .A1(n12061), .A2(n12128), .B1(n12125), .B2(n12573), .ZN(
        n12062) );
  NOR2_X1 U15053 ( .A1(n12063), .A2(n12062), .ZN(n12064) );
  NAND4_X1 U15054 ( .A1(n12067), .A2(n12066), .A3(n12065), .A4(n12064), .ZN(
        n12071) );
  NAND2_X1 U15055 ( .A1(n12068), .A2(n12399), .ZN(n14160) );
  OR2_X1 U15056 ( .A1(n12400), .A2(n14160), .ZN(n12403) );
  INV_X1 U15057 ( .A(n12404), .ZN(n12069) );
  NAND2_X1 U15058 ( .A1(n12403), .A2(n12069), .ZN(n12070) );
  INV_X1 U15059 ( .A(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12072) );
  OAI22_X1 U15060 ( .A1(n19161), .A2(n12128), .B1(n12129), .B2(n12072), .ZN(
        n12076) );
  OAI22_X1 U15061 ( .A1(n12074), .A2(n12131), .B1(n12132), .B2(n12073), .ZN(
        n12075) );
  INV_X1 U15062 ( .A(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12077) );
  OAI22_X1 U15063 ( .A1(n12078), .A2(n12121), .B1(n12122), .B2(n12077), .ZN(
        n12079) );
  INV_X1 U15064 ( .A(n12079), .ZN(n12082) );
  INV_X1 U15065 ( .A(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12602) );
  OAI22_X1 U15066 ( .A1(n12602), .A2(n19339), .B1(n12125), .B2(n11253), .ZN(
        n12080) );
  INV_X1 U15067 ( .A(n12080), .ZN(n12081) );
  NAND3_X1 U15068 ( .A1(n12083), .A2(n12082), .A3(n12081), .ZN(n12098) );
  INV_X1 U15069 ( .A(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12085) );
  INV_X1 U15070 ( .A(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12086) );
  OAI22_X1 U15071 ( .A1(n12087), .A2(n12107), .B1(n12108), .B2(n12086), .ZN(
        n12088) );
  NOR2_X1 U15072 ( .A1(n12089), .A2(n12088), .ZN(n12096) );
  NOR2_X1 U15073 ( .A1(n12094), .A2(n12093), .ZN(n12095) );
  NAND2_X1 U15074 ( .A1(n12096), .A2(n12095), .ZN(n12097) );
  OAI21_X1 U15075 ( .B1(n12098), .B2(n12097), .A(n19796), .ZN(n12101) );
  NAND2_X1 U15076 ( .A1(n12068), .A2(n12099), .ZN(n12100) );
  INV_X1 U15077 ( .A(n12411), .ZN(n12103) );
  INV_X1 U15078 ( .A(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12106) );
  OAI22_X1 U15079 ( .A1(n12106), .A2(n12104), .B1(n19425), .B2(n12105), .ZN(
        n12112) );
  OAI22_X1 U15080 ( .A1(n12110), .A2(n12107), .B1(n12108), .B2(n12109), .ZN(
        n12111) );
  NOR2_X1 U15081 ( .A1(n12112), .A2(n12111), .ZN(n12140) );
  INV_X1 U15082 ( .A(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n12116) );
  OAI22_X1 U15083 ( .A1(n12116), .A2(n12113), .B1(n12114), .B2(n12115), .ZN(
        n12120) );
  INV_X1 U15084 ( .A(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n12118) );
  INV_X1 U15085 ( .A(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12635) );
  OAI22_X1 U15086 ( .A1(n12118), .A2(n12117), .B1(n9673), .B2(n12635), .ZN(
        n12119) );
  NOR2_X1 U15087 ( .A1(n12120), .A2(n12119), .ZN(n12139) );
  INV_X1 U15088 ( .A(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12123) );
  OAI22_X1 U15089 ( .A1(n12124), .A2(n12121), .B1(n12122), .B2(n12123), .ZN(
        n12127) );
  INV_X1 U15090 ( .A(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12636) );
  INV_X1 U15091 ( .A(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12640) );
  OAI22_X1 U15092 ( .A1(n12636), .A2(n19339), .B1(n12125), .B2(n12640), .ZN(
        n12126) );
  NOR2_X1 U15093 ( .A1(n12127), .A2(n12126), .ZN(n12138) );
  INV_X1 U15094 ( .A(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12130) );
  OAI22_X1 U15095 ( .A1(n19171), .A2(n12128), .B1(n12129), .B2(n12130), .ZN(
        n12136) );
  INV_X1 U15096 ( .A(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12134) );
  INV_X1 U15097 ( .A(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12133) );
  OAI22_X1 U15098 ( .A1(n12134), .A2(n12131), .B1(n12132), .B2(n12133), .ZN(
        n12135) );
  NOR2_X1 U15099 ( .A1(n12136), .A2(n12135), .ZN(n12137) );
  NAND4_X1 U15100 ( .A1(n12140), .A2(n12139), .A3(n12138), .A4(n12137), .ZN(
        n12144) );
  INV_X1 U15101 ( .A(n12141), .ZN(n12142) );
  NAND2_X1 U15102 ( .A1(n12142), .A2(n12068), .ZN(n12143) );
  NAND2_X1 U15103 ( .A1(n12417), .A2(n12426), .ZN(n12149) );
  NOR2_X1 U15104 ( .A1(n12147), .A2(n12146), .ZN(n12148) );
  OR2_X1 U15105 ( .A1(n12145), .A2(n12148), .ZN(n18907) );
  OAI21_X1 U15106 ( .B1(n12151), .B2(n12150), .A(n12411), .ZN(n12398) );
  INV_X1 U15107 ( .A(n12322), .ZN(n12426) );
  OAI21_X1 U15108 ( .B1(n12153), .B2(n12152), .A(n12165), .ZN(n13555) );
  OAI21_X1 U15109 ( .B1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n19783), .A(
        n12154), .ZN(n12340) );
  INV_X1 U15110 ( .A(n12340), .ZN(n12370) );
  MUX2_X1 U15111 ( .A(n12399), .B(n12370), .S(n11991), .Z(n12362) );
  MUX2_X1 U15112 ( .A(n12362), .B(P2_EBX_REG_0__SCAN_IN), .S(n12327), .Z(
        n18921) );
  NAND2_X1 U15113 ( .A1(n18921), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n14163) );
  NAND3_X1 U15114 ( .A1(n12327), .A2(P2_EBX_REG_0__SCAN_IN), .A3(
        P2_EBX_REG_1__SCAN_IN), .ZN(n12155) );
  NAND2_X1 U15115 ( .A1(n12158), .A2(n12155), .ZN(n13512) );
  NOR2_X1 U15116 ( .A1(n14163), .A2(n13512), .ZN(n12156) );
  NAND2_X1 U15117 ( .A1(n14163), .A2(n13512), .ZN(n13000) );
  OAI21_X1 U15118 ( .B1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n12156), .A(
        n13000), .ZN(n13019) );
  XNOR2_X1 U15119 ( .A(n12158), .B(n12157), .ZN(n13469) );
  XNOR2_X1 U15120 ( .A(n13469), .B(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n13018) );
  OR2_X1 U15121 ( .A1(n13019), .A2(n13018), .ZN(n19108) );
  NAND2_X1 U15122 ( .A1(n13469), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n12159) );
  NAND2_X1 U15123 ( .A1(n19108), .A2(n12159), .ZN(n13526) );
  INV_X1 U15124 ( .A(n13526), .ZN(n12160) );
  NAND2_X1 U15125 ( .A1(n13524), .A2(n12160), .ZN(n12164) );
  INV_X1 U15126 ( .A(n12161), .ZN(n12163) );
  NAND2_X1 U15127 ( .A1(n12163), .A2(n12162), .ZN(n13525) );
  NAND2_X1 U15128 ( .A1(n12164), .A2(n13525), .ZN(n19082) );
  XNOR2_X1 U15129 ( .A(n12166), .B(n12165), .ZN(n13485) );
  XNOR2_X1 U15130 ( .A(n13485), .B(n19101), .ZN(n19083) );
  OAI22_X2 U15131 ( .A1(n19082), .A2(n19083), .B1(n13485), .B2(n19101), .ZN(
        n13674) );
  NAND2_X1 U15132 ( .A1(n12167), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n12168) );
  NAND2_X1 U15133 ( .A1(n12201), .A2(n12198), .ZN(n12197) );
  INV_X1 U15134 ( .A(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12171) );
  OAI22_X1 U15135 ( .A1(n12171), .A2(n12104), .B1(n12107), .B2(n12170), .ZN(
        n12175) );
  INV_X1 U15136 ( .A(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12173) );
  OAI22_X1 U15137 ( .A1(n12173), .A2(n12113), .B1(n12114), .B2(n12172), .ZN(
        n12174) );
  NOR2_X1 U15138 ( .A1(n12175), .A2(n12174), .ZN(n12192) );
  OAI22_X1 U15139 ( .A1(n12815), .A2(n12131), .B1(n12128), .B2(n19175), .ZN(
        n12178) );
  INV_X1 U15140 ( .A(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12176) );
  OAI22_X1 U15141 ( .A1(n12176), .A2(n12129), .B1(n9673), .B2(n19644), .ZN(
        n12177) );
  NOR2_X1 U15142 ( .A1(n12178), .A2(n12177), .ZN(n12191) );
  OAI22_X1 U15143 ( .A1(n12180), .A2(n19425), .B1(n12108), .B2(n12179), .ZN(
        n12184) );
  OAI22_X1 U15144 ( .A1(n12182), .A2(n12121), .B1(n12117), .B2(n12181), .ZN(
        n12183) );
  NOR2_X1 U15145 ( .A1(n12184), .A2(n12183), .ZN(n12190) );
  INV_X1 U15146 ( .A(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12185) );
  INV_X1 U15147 ( .A(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12656) );
  OAI22_X1 U15148 ( .A1(n12185), .A2(n12122), .B1(n12125), .B2(n12656), .ZN(
        n12188) );
  INV_X1 U15149 ( .A(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12652) );
  OAI22_X1 U15150 ( .A1(n12652), .A2(n19339), .B1(n12132), .B2(n12186), .ZN(
        n12187) );
  NOR2_X1 U15151 ( .A1(n12188), .A2(n12187), .ZN(n12189) );
  NAND4_X1 U15152 ( .A1(n12192), .A2(n12191), .A3(n12190), .A4(n12189), .ZN(
        n12196) );
  INV_X1 U15153 ( .A(n12193), .ZN(n12194) );
  NAND2_X1 U15154 ( .A1(n12194), .A2(n12068), .ZN(n12195) );
  INV_X1 U15155 ( .A(n12199), .ZN(n12421) );
  NAND2_X1 U15156 ( .A1(n12197), .A2(n12421), .ZN(n12202) );
  NAND2_X1 U15157 ( .A1(n12202), .A2(n12427), .ZN(n12420) );
  NOR2_X1 U15158 ( .A1(n12145), .A2(n12203), .ZN(n12204) );
  OR2_X1 U15159 ( .A1(n12212), .A2(n12204), .ZN(n18891) );
  NAND2_X1 U15160 ( .A1(n12327), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n12208) );
  XNOR2_X1 U15161 ( .A(n12209), .B(n12208), .ZN(n18873) );
  AND2_X1 U15162 ( .A1(n12322), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n12210) );
  NAND2_X1 U15163 ( .A1(n18873), .A2(n12210), .ZN(n14789) );
  XNOR2_X1 U15164 ( .A(n12212), .B(n10061), .ZN(n12214) );
  NAND2_X1 U15165 ( .A1(n12214), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n14786) );
  NAND2_X1 U15166 ( .A1(n18873), .A2(n12322), .ZN(n12213) );
  NAND2_X1 U15167 ( .A1(n12213), .A2(n16118), .ZN(n14790) );
  INV_X1 U15168 ( .A(n12214), .ZN(n18884) );
  NAND2_X1 U15169 ( .A1(n18884), .A2(n13822), .ZN(n14788) );
  AND2_X1 U15170 ( .A1(n14790), .A2(n14788), .ZN(n12215) );
  AND2_X1 U15171 ( .A1(n12327), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n12216) );
  XNOR2_X1 U15172 ( .A(n12217), .B(n12216), .ZN(n13540) );
  NAND2_X1 U15173 ( .A1(n13540), .A2(n12322), .ZN(n12229) );
  NAND2_X1 U15174 ( .A1(n12327), .A2(P2_EBX_REG_10__SCAN_IN), .ZN(n12219) );
  MUX2_X1 U15175 ( .A(P2_EBX_REG_10__SCAN_IN), .B(n12219), .S(n12218), .Z(
        n12220) );
  NAND2_X1 U15176 ( .A1(n12220), .A2(n12301), .ZN(n18858) );
  INV_X1 U15177 ( .A(n18858), .ZN(n12221) );
  NAND2_X1 U15178 ( .A1(n12221), .A2(n12322), .ZN(n12230) );
  NAND2_X1 U15179 ( .A1(n12230), .A2(n15006), .ZN(n15000) );
  NAND2_X1 U15180 ( .A1(n12327), .A2(P2_EBX_REG_11__SCAN_IN), .ZN(n12222) );
  OR2_X1 U15181 ( .A1(n12223), .A2(n12222), .ZN(n12226) );
  INV_X1 U15182 ( .A(n12224), .ZN(n12225) );
  NAND2_X1 U15183 ( .A1(n18849), .A2(n12322), .ZN(n12227) );
  INV_X1 U15184 ( .A(n12227), .ZN(n12228) );
  NAND2_X1 U15185 ( .A1(n12228), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n14977) );
  NOR2_X1 U15186 ( .A1(n12229), .A2(n15029), .ZN(n15024) );
  NOR2_X1 U15187 ( .A1(n15006), .A2(n12230), .ZN(n14998) );
  NOR2_X1 U15188 ( .A1(n15024), .A2(n14998), .ZN(n14976) );
  AND2_X1 U15189 ( .A1(n14977), .A2(n14976), .ZN(n14727) );
  INV_X1 U15190 ( .A(n12231), .ZN(n12233) );
  NAND2_X1 U15191 ( .A1(n12233), .A2(n12232), .ZN(n12234) );
  NAND2_X1 U15192 ( .A1(n12257), .A2(n12234), .ZN(n18835) );
  NAND2_X1 U15193 ( .A1(n12322), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n12235) );
  INV_X1 U15194 ( .A(n18835), .ZN(n12236) );
  NAND2_X1 U15195 ( .A1(n12236), .A2(n12322), .ZN(n12237) );
  NAND2_X1 U15196 ( .A1(n12237), .A2(n16106), .ZN(n16035) );
  NAND2_X1 U15197 ( .A1(n12239), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n12238) );
  MUX2_X1 U15198 ( .A(n12239), .B(n12238), .S(n12327), .Z(n12240) );
  NAND2_X1 U15199 ( .A1(n18760), .A2(n12322), .ZN(n12241) );
  NAND2_X1 U15200 ( .A1(n12241), .A2(n14952), .ZN(n14775) );
  NAND3_X1 U15201 ( .A1(n12242), .A2(n12327), .A3(P2_EBX_REG_19__SCAN_IN), 
        .ZN(n12243) );
  AND2_X1 U15202 ( .A1(n12243), .A2(n12245), .ZN(n14067) );
  NAND2_X1 U15203 ( .A1(n14067), .A2(n12322), .ZN(n12275) );
  INV_X1 U15204 ( .A(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n14943) );
  NAND2_X1 U15205 ( .A1(n12275), .A2(n14943), .ZN(n14764) );
  NAND2_X1 U15206 ( .A1(n12327), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n12244) );
  XNOR2_X1 U15207 ( .A(n12245), .B(n12244), .ZN(n18749) );
  NAND2_X1 U15208 ( .A1(n18749), .A2(n12322), .ZN(n12278) );
  INV_X1 U15209 ( .A(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n15435) );
  AND2_X1 U15210 ( .A1(n12327), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n12246) );
  INV_X1 U15211 ( .A(n12301), .ZN(n12295) );
  AOI21_X1 U15212 ( .B1(n12251), .B2(n12246), .A(n12295), .ZN(n12248) );
  AND2_X1 U15213 ( .A1(n12248), .A2(n12247), .ZN(n18788) );
  NAND2_X1 U15214 ( .A1(n18788), .A2(n12322), .ZN(n12271) );
  XNOR2_X1 U15215 ( .A(n12271), .B(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15295) );
  NAND2_X1 U15216 ( .A1(n12255), .A2(n18808), .ZN(n12250) );
  AND2_X1 U15217 ( .A1(n12327), .A2(P2_EBX_REG_15__SCAN_IN), .ZN(n12249) );
  NAND2_X1 U15218 ( .A1(n12250), .A2(n12249), .ZN(n12252) );
  NAND2_X1 U15219 ( .A1(n12252), .A2(n12251), .ZN(n18799) );
  OR2_X1 U15220 ( .A1(n18799), .A2(n12426), .ZN(n12253) );
  NAND2_X1 U15221 ( .A1(n12253), .A2(n12269), .ZN(n16010) );
  AND2_X1 U15222 ( .A1(n12327), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n12254) );
  XNOR2_X1 U15223 ( .A(n12255), .B(n12254), .ZN(n18813) );
  NAND2_X1 U15224 ( .A1(n18813), .A2(n12322), .ZN(n12256) );
  INV_X1 U15225 ( .A(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n12433) );
  NAND2_X1 U15226 ( .A1(n12256), .A2(n12433), .ZN(n16020) );
  XNOR2_X1 U15227 ( .A(n12257), .B(n9738), .ZN(n18821) );
  NAND2_X1 U15228 ( .A1(n18821), .A2(n12322), .ZN(n12258) );
  NAND2_X1 U15229 ( .A1(n12258), .A2(n16085), .ZN(n14959) );
  AND3_X1 U15230 ( .A1(n16010), .A2(n16020), .A3(n14959), .ZN(n12259) );
  AND2_X1 U15231 ( .A1(n15295), .A2(n12259), .ZN(n12266) );
  XNOR2_X1 U15232 ( .A(n12261), .B(n10073), .ZN(n18775) );
  NAND2_X1 U15233 ( .A1(n18775), .A2(n12322), .ZN(n12262) );
  INV_X1 U15234 ( .A(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n15996) );
  NAND2_X1 U15235 ( .A1(n12262), .A2(n15996), .ZN(n14735) );
  NAND2_X1 U15236 ( .A1(n12327), .A2(P2_EBX_REG_21__SCAN_IN), .ZN(n12263) );
  OAI211_X1 U15237 ( .C1(n12264), .C2(n12263), .A(n12301), .B(n12284), .ZN(
        n18740) );
  OR2_X1 U15238 ( .A1(n18740), .A2(n12426), .ZN(n12265) );
  INV_X1 U15239 ( .A(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n14927) );
  NAND2_X1 U15240 ( .A1(n12265), .A2(n14927), .ZN(n14738) );
  NAND2_X1 U15241 ( .A1(n12322), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n12267) );
  OR2_X1 U15242 ( .A1(n18740), .A2(n12267), .ZN(n14737) );
  AND2_X1 U15243 ( .A1(n12322), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n12268) );
  NAND2_X1 U15244 ( .A1(n18775), .A2(n12268), .ZN(n14734) );
  AND2_X1 U15245 ( .A1(n12322), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n12270) );
  NAND2_X1 U15246 ( .A1(n18821), .A2(n12270), .ZN(n14958) );
  AND2_X1 U15247 ( .A1(n16009), .A2(n14958), .ZN(n12273) );
  OR2_X1 U15248 ( .A1(n12271), .A2(n15317), .ZN(n14732) );
  INV_X1 U15249 ( .A(n18813), .ZN(n12272) );
  AND4_X1 U15250 ( .A1(n14734), .A2(n12273), .A3(n14732), .A4(n16019), .ZN(
        n12277) );
  AND2_X1 U15251 ( .A1(n12322), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n12274) );
  NAND2_X1 U15252 ( .A1(n18760), .A2(n12274), .ZN(n14774) );
  INV_X1 U15253 ( .A(n12275), .ZN(n12276) );
  NAND2_X1 U15254 ( .A1(n12276), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n14765) );
  NAND4_X1 U15255 ( .A1(n14737), .A2(n12277), .A3(n14774), .A4(n14765), .ZN(
        n12280) );
  INV_X1 U15256 ( .A(n12278), .ZN(n12279) );
  NOR2_X1 U15257 ( .A1(n12280), .A2(n14748), .ZN(n12281) );
  INV_X1 U15258 ( .A(n12282), .ZN(n12283) );
  NAND2_X1 U15259 ( .A1(n12284), .A2(n12283), .ZN(n12285) );
  NAND2_X1 U15260 ( .A1(n12289), .A2(n12285), .ZN(n15306) );
  OR2_X1 U15261 ( .A1(n15306), .A2(n12426), .ZN(n12286) );
  NAND2_X1 U15262 ( .A1(n12286), .A2(n14910), .ZN(n14905) );
  NAND2_X1 U15263 ( .A1(n14906), .A2(n14905), .ZN(n12287) );
  NAND2_X1 U15264 ( .A1(n12287), .A2(n14904), .ZN(n14878) );
  NAND2_X1 U15265 ( .A1(n12289), .A2(n12288), .ZN(n12290) );
  NAND2_X1 U15266 ( .A1(n12297), .A2(n12290), .ZN(n12976) );
  NAND2_X1 U15267 ( .A1(n14878), .A2(n14879), .ZN(n12294) );
  NAND2_X1 U15268 ( .A1(n12322), .A2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n12292) );
  AND2_X1 U15269 ( .A1(n12327), .A2(P2_EBX_REG_24__SCAN_IN), .ZN(n12296) );
  AOI21_X1 U15270 ( .B1(n12297), .B2(n12296), .A(n12295), .ZN(n12298) );
  AND2_X1 U15271 ( .A1(n12298), .A2(n12299), .ZN(n15919) );
  NAND2_X1 U15272 ( .A1(n12327), .A2(P2_EBX_REG_25__SCAN_IN), .ZN(n12300) );
  MUX2_X1 U15273 ( .A(P2_EBX_REG_25__SCAN_IN), .B(n12300), .S(n12299), .Z(
        n12302) );
  NAND2_X1 U15274 ( .A1(n12327), .A2(P2_EBX_REG_26__SCAN_IN), .ZN(n12303) );
  OR2_X1 U15275 ( .A1(n12304), .A2(n12303), .ZN(n12306) );
  INV_X1 U15276 ( .A(n12305), .ZN(n12329) );
  AND2_X1 U15277 ( .A1(n12313), .A2(n12307), .ZN(n12308) );
  OR2_X1 U15278 ( .A1(n12319), .A2(n12308), .ZN(n15886) );
  INV_X1 U15279 ( .A(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n12953) );
  INV_X1 U15280 ( .A(n12309), .ZN(n12311) );
  NAND2_X1 U15281 ( .A1(n12311), .A2(n12310), .ZN(n12312) );
  NAND2_X1 U15282 ( .A1(n12313), .A2(n12312), .ZN(n15901) );
  INV_X1 U15283 ( .A(n12314), .ZN(n12315) );
  NAND2_X1 U15284 ( .A1(n12315), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n12317) );
  AND2_X1 U15285 ( .A1(n12322), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n12316) );
  NAND2_X1 U15286 ( .A1(n14585), .A2(n12316), .ZN(n14715) );
  XNOR2_X1 U15287 ( .A(n12319), .B(n12318), .ZN(n14578) );
  INV_X1 U15288 ( .A(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n14821) );
  OAI21_X1 U15289 ( .B1(n14578), .B2(n12426), .A(n14821), .ZN(n12499) );
  AOI21_X1 U15290 ( .B1(n12320), .B2(n12322), .A(
        P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n14697) );
  INV_X1 U15291 ( .A(n14578), .ZN(n12323) );
  NAND3_X1 U15292 ( .A1(n12323), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        n12322), .ZN(n14696) );
  INV_X1 U15293 ( .A(n14696), .ZN(n12324) );
  NOR2_X1 U15294 ( .A1(n12326), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n12328) );
  MUX2_X1 U15295 ( .A(n12329), .B(n12328), .S(n12327), .Z(n15872) );
  NAND2_X1 U15296 ( .A1(n15872), .A2(n12322), .ZN(n12330) );
  XNOR2_X1 U15297 ( .A(n12330), .B(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n12331) );
  XNOR2_X1 U15298 ( .A(n12332), .B(n12331), .ZN(n14193) );
  INV_X1 U15299 ( .A(n12333), .ZN(n12335) );
  NAND2_X1 U15300 ( .A1(n12335), .A2(n12334), .ZN(n12364) );
  OAI21_X1 U15301 ( .B1(n12355), .B2(n12068), .A(n12336), .ZN(n12338) );
  NAND2_X1 U15302 ( .A1(n12338), .A2(n12337), .ZN(n12348) );
  NAND2_X1 U15303 ( .A1(n13063), .A2(n12339), .ZN(n12345) );
  OAI21_X1 U15304 ( .B1(n12340), .B2(n12359), .A(n12463), .ZN(n12344) );
  NAND2_X1 U15305 ( .A1(n12068), .A2(n12340), .ZN(n12342) );
  NAND3_X1 U15306 ( .A1(n12342), .A2(n13728), .A3(n12341), .ZN(n12343) );
  NAND3_X1 U15307 ( .A1(n12345), .A2(n12344), .A3(n12343), .ZN(n12347) );
  AOI21_X1 U15308 ( .B1(n12348), .B2(n12347), .A(n12346), .ZN(n12349) );
  AOI21_X1 U15309 ( .B1(n12364), .B2(n11991), .A(n12349), .ZN(n12350) );
  NOR2_X1 U15310 ( .A1(n12350), .A2(n12365), .ZN(n12351) );
  MUX2_X1 U15311 ( .A(n13643), .B(n12351), .S(P2_STATE2_REG_0__SCAN_IN), .Z(
        n12354) );
  NAND2_X1 U15312 ( .A1(n9654), .A2(n12352), .ZN(n12353) );
  NAND2_X1 U15313 ( .A1(n12365), .A2(n12355), .ZN(n12356) );
  NAND2_X1 U15314 ( .A1(n13635), .A2(n19796), .ZN(n13154) );
  INV_X1 U15315 ( .A(n13628), .ZN(n13056) );
  NAND2_X1 U15316 ( .A1(n13574), .A2(n13056), .ZN(n12396) );
  AOI21_X1 U15317 ( .B1(n12357), .B2(n13728), .A(n11450), .ZN(n12358) );
  NAND2_X1 U15318 ( .A1(n13154), .A2(n12358), .ZN(n12395) );
  INV_X1 U15319 ( .A(n12359), .ZN(n12361) );
  AOI21_X1 U15320 ( .B1(n12362), .B2(n12361), .A(n12360), .ZN(n12363) );
  NOR2_X1 U15321 ( .A1(n12364), .A2(n12363), .ZN(n12366) );
  OR2_X1 U15322 ( .A1(n12366), .A2(n12365), .ZN(n19788) );
  AND2_X1 U15323 ( .A1(n11389), .A2(n12068), .ZN(n12377) );
  INV_X1 U15324 ( .A(n12377), .ZN(n12368) );
  OR2_X1 U15325 ( .A1(n12367), .A2(n12368), .ZN(n19786) );
  AOI21_X1 U15326 ( .B1(n12370), .B2(n12369), .A(n13631), .ZN(n12372) );
  OR2_X1 U15327 ( .A1(n12371), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n13062) );
  INV_X1 U15328 ( .A(P2_FLUSH_REG_SCAN_IN), .ZN(n12993) );
  OAI21_X1 U15329 ( .B1(n12662), .B2(n13062), .A(n12993), .ZN(n19775) );
  MUX2_X1 U15330 ( .A(n12372), .B(n19775), .S(P2_STATE2_REG_1__SCAN_IN), .Z(
        n19792) );
  NAND2_X1 U15331 ( .A1(n19796), .A2(n19792), .ZN(n12373) );
  OAI22_X1 U15332 ( .A1(n19788), .A2(n19786), .B1(n12367), .B2(n12373), .ZN(
        n12502) );
  MUX2_X1 U15333 ( .A(n12374), .B(n11436), .S(n12068), .Z(n12392) );
  NOR2_X1 U15334 ( .A1(n13631), .A2(n19807), .ZN(n12388) );
  INV_X1 U15335 ( .A(n12388), .ZN(n12391) );
  OAI21_X1 U15336 ( .B1(n12376), .B2(n12375), .A(n9639), .ZN(n12378) );
  NAND2_X1 U15337 ( .A1(n12378), .A2(n12377), .ZN(n12458) );
  NAND2_X1 U15338 ( .A1(n12379), .A2(n12068), .ZN(n12446) );
  NAND2_X1 U15339 ( .A1(n12446), .A2(n13728), .ZN(n12380) );
  NAND2_X1 U15340 ( .A1(n12380), .A2(n9639), .ZN(n12381) );
  NAND2_X1 U15341 ( .A1(n12381), .A2(n11436), .ZN(n12382) );
  AND4_X1 U15342 ( .A1(n12458), .A2(n11474), .A3(n12383), .A4(n12382), .ZN(
        n12387) );
  NAND2_X1 U15343 ( .A1(n12384), .A2(n11436), .ZN(n12385) );
  NAND2_X1 U15344 ( .A1(n13152), .A2(n12385), .ZN(n12386) );
  NAND2_X1 U15345 ( .A1(n12387), .A2(n12386), .ZN(n12447) );
  NAND2_X1 U15346 ( .A1(n19795), .A2(n12388), .ZN(n12389) );
  NOR2_X1 U15347 ( .A1(n12374), .A2(n12389), .ZN(n12390) );
  NOR2_X1 U15348 ( .A1(n12447), .A2(n12390), .ZN(n13051) );
  OAI21_X1 U15349 ( .B1(n12392), .B2(n12391), .A(n13051), .ZN(n12393) );
  NOR2_X1 U15350 ( .A1(n12502), .A2(n12393), .ZN(n12394) );
  OAI211_X1 U15351 ( .C1(n13154), .C2(n12396), .A(n12395), .B(n12394), .ZN(
        n12397) );
  INV_X1 U15352 ( .A(n16152), .ZN(n12859) );
  OR2_X1 U15353 ( .A1(n12367), .A2(n11991), .ZN(n19791) );
  AND2_X1 U15354 ( .A1(n14160), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n14162) );
  XNOR2_X1 U15355 ( .A(n12400), .B(n12399), .ZN(n12401) );
  NAND2_X1 U15356 ( .A1(n14162), .A2(n12401), .ZN(n12402) );
  XOR2_X1 U15357 ( .A(n12401), .B(n14162), .Z(n13003) );
  NAND2_X1 U15358 ( .A1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n13003), .ZN(
        n13002) );
  NAND2_X1 U15359 ( .A1(n12402), .A2(n13002), .ZN(n12406) );
  XOR2_X1 U15360 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .B(n12406), .Z(
        n13014) );
  INV_X1 U15361 ( .A(n12403), .ZN(n12405) );
  XNOR2_X1 U15362 ( .A(n12405), .B(n12404), .ZN(n13013) );
  NAND2_X1 U15363 ( .A1(n13014), .A2(n13013), .ZN(n13012) );
  NAND2_X1 U15364 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n12406), .ZN(
        n12407) );
  NAND2_X1 U15365 ( .A1(n13012), .A2(n12407), .ZN(n12408) );
  XNOR2_X1 U15366 ( .A(n12408), .B(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n13523) );
  NAND2_X1 U15367 ( .A1(n12408), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n12409) );
  NAND2_X1 U15368 ( .A1(n12410), .A2(n12409), .ZN(n19084) );
  NAND2_X1 U15369 ( .A1(n19085), .A2(n19101), .ZN(n12413) );
  NAND2_X1 U15370 ( .A1(n19084), .A2(n12413), .ZN(n12416) );
  INV_X1 U15371 ( .A(n19085), .ZN(n12414) );
  NAND2_X1 U15372 ( .A1(n12414), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n12415) );
  INV_X1 U15373 ( .A(n12417), .ZN(n12419) );
  INV_X1 U15374 ( .A(n13686), .ZN(n12422) );
  NAND2_X1 U15375 ( .A1(n12422), .A2(n12421), .ZN(n12423) );
  NAND2_X1 U15376 ( .A1(n13835), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n13834) );
  NAND2_X1 U15377 ( .A1(n13682), .A2(n13686), .ZN(n12424) );
  NAND2_X1 U15378 ( .A1(n12424), .A2(n9629), .ZN(n12425) );
  OR2_X2 U15379 ( .A1(n12427), .A2(n12426), .ZN(n12431) );
  NAND2_X1 U15380 ( .A1(n12427), .A2(n12426), .ZN(n12428) );
  OR2_X2 U15381 ( .A1(n12429), .A2(n13822), .ZN(n12430) );
  INV_X1 U15382 ( .A(n12431), .ZN(n12432) );
  NAND2_X1 U15383 ( .A1(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n14985) );
  NOR2_X1 U15384 ( .A1(n15029), .A2(n14985), .ZN(n14963) );
  NAND2_X1 U15385 ( .A1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n16084) );
  NOR2_X1 U15386 ( .A1(n12433), .A2(n16084), .ZN(n15301) );
  NOR2_X1 U15387 ( .A1(n12269), .A2(n15317), .ZN(n15315) );
  NAND4_X1 U15388 ( .A1(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n14963), .A3(
        n15301), .A4(n15315), .ZN(n14948) );
  INV_X1 U15389 ( .A(n14948), .ZN(n14891) );
  AND3_X1 U15390 ( .A1(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n12434) );
  NAND2_X1 U15391 ( .A1(n14891), .A2(n12434), .ZN(n14883) );
  INV_X1 U15392 ( .A(n14883), .ZN(n12435) );
  OR2_X2 U15393 ( .A1(n14752), .A2(n14927), .ZN(n14901) );
  NAND2_X1 U15394 ( .A1(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n14893) );
  NAND2_X2 U15395 ( .A1(n12943), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n12944) );
  NAND2_X1 U15396 ( .A1(n14700), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n12436) );
  XNOR2_X1 U15397 ( .A(n12436), .B(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n14191) );
  NAND2_X1 U15398 ( .A1(n12437), .A2(P2_REIP_REG_31__SCAN_IN), .ZN(n12439) );
  AOI22_X1 U15399 ( .A1(n11963), .A2(P2_EAX_REG_31__SCAN_IN), .B1(n11976), 
        .B2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n12438) );
  NAND2_X1 U15400 ( .A1(n12439), .A2(n12438), .ZN(n12440) );
  INV_X1 U15401 ( .A(n13600), .ZN(n12443) );
  NAND2_X1 U15402 ( .A1(n12443), .A2(n12442), .ZN(n13630) );
  OAI21_X1 U15403 ( .B1(n12068), .B2(n13641), .A(n13630), .ZN(n12444) );
  INV_X1 U15404 ( .A(n12444), .ZN(n12445) );
  NOR2_X1 U15405 ( .A1(n13822), .A2(n16118), .ZN(n16117) );
  NAND2_X1 U15406 ( .A1(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n13677) );
  NOR2_X1 U15407 ( .A1(n12447), .A2(n12446), .ZN(n12857) );
  INV_X1 U15408 ( .A(n12857), .ZN(n13633) );
  NOR2_X1 U15409 ( .A1(n11463), .A2(n13762), .ZN(n19117) );
  INV_X1 U15410 ( .A(n19117), .ZN(n19133) );
  NOR2_X1 U15411 ( .A1(n12448), .A2(n19133), .ZN(n12465) );
  NAND2_X1 U15412 ( .A1(n12448), .A2(n19133), .ZN(n19105) );
  NAND2_X1 U15413 ( .A1(n12449), .A2(n13063), .ZN(n12858) );
  INV_X1 U15414 ( .A(n12861), .ZN(n19798) );
  NAND2_X1 U15415 ( .A1(n11474), .A2(n11450), .ZN(n12450) );
  AOI22_X1 U15416 ( .A1(n19798), .A2(n12450), .B1(n13574), .B2(n11389), .ZN(
        n12455) );
  NAND3_X1 U15417 ( .A1(n12453), .A2(n12452), .A3(n12451), .ZN(n12454) );
  AND4_X1 U15418 ( .A1(n12456), .A2(n12858), .A3(n12455), .A4(n12454), .ZN(
        n12462) );
  NAND2_X1 U15419 ( .A1(n12457), .A2(n19796), .ZN(n13599) );
  NAND2_X1 U15420 ( .A1(n13599), .A2(n12458), .ZN(n12460) );
  NAND2_X1 U15421 ( .A1(n12460), .A2(n12459), .ZN(n12461) );
  NAND2_X1 U15422 ( .A1(n12462), .A2(n12461), .ZN(n13598) );
  NAND2_X1 U15423 ( .A1(n12449), .A2(n12463), .ZN(n13069) );
  INV_X1 U15424 ( .A(n13069), .ZN(n13588) );
  NOR2_X1 U15425 ( .A1(n13598), .A2(n13588), .ZN(n12464) );
  NOR2_X1 U15426 ( .A1(n12481), .A2(n12464), .ZN(n14882) );
  OAI211_X1 U15427 ( .C1(n19116), .C2(n12465), .A(n19105), .B(n19132), .ZN(
        n16136) );
  NOR2_X1 U15428 ( .A1(n12162), .A2(n16136), .ZN(n19102) );
  INV_X1 U15429 ( .A(n19102), .ZN(n12466) );
  NOR2_X1 U15430 ( .A1(n13677), .A2(n12466), .ZN(n14056) );
  NOR4_X1 U15431 ( .A1(n15028), .A2(n14893), .A3(n14927), .A4(n14883), .ZN(
        n12487) );
  NAND2_X1 U15432 ( .A1(n12487), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n14859) );
  NAND2_X1 U15433 ( .A1(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n12488) );
  NAND2_X1 U15434 ( .A1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n14818) );
  NOR2_X1 U15435 ( .A1(n14821), .A2(n14818), .ZN(n14803) );
  INV_X1 U15436 ( .A(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n12492) );
  NAND4_X1 U15437 ( .A1(n14829), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .A3(
        n14803), .A4(n12492), .ZN(n12467) );
  NAND2_X1 U15438 ( .A1(n19081), .A2(P2_REIP_REG_31__SCAN_IN), .ZN(n14188) );
  NAND2_X1 U15439 ( .A1(n12467), .A2(n14188), .ZN(n12468) );
  INV_X1 U15440 ( .A(n12471), .ZN(n12478) );
  NAND2_X1 U15441 ( .A1(n12472), .A2(P2_REIP_REG_31__SCAN_IN), .ZN(n12474) );
  NAND2_X1 U15442 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n12473) );
  OAI211_X1 U15443 ( .C1(n12476), .C2(n12475), .A(n12474), .B(n12473), .ZN(
        n12477) );
  AOI21_X1 U15444 ( .B1(n12470), .B2(n12478), .A(n12477), .ZN(n12479) );
  NAND2_X1 U15445 ( .A1(n12470), .A2(n12068), .ZN(n12480) );
  OR2_X1 U15446 ( .A1(n12481), .A2(n12480), .ZN(n19112) );
  INV_X1 U15447 ( .A(n14803), .ZN(n12491) );
  INV_X1 U15448 ( .A(n19132), .ZN(n16144) );
  INV_X1 U15449 ( .A(n12481), .ZN(n12483) );
  INV_X1 U15450 ( .A(n12482), .ZN(n18810) );
  NOR2_X1 U15451 ( .A1(n12483), .A2(n18810), .ZN(n19124) );
  INV_X1 U15452 ( .A(n14882), .ZN(n15300) );
  AOI21_X1 U15453 ( .B1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n19117), .A(
        n15300), .ZN(n19106) );
  INV_X1 U15454 ( .A(n19105), .ZN(n12484) );
  AND2_X1 U15455 ( .A1(n19116), .A2(n12484), .ZN(n19113) );
  NOR3_X1 U15456 ( .A1(n19124), .A2(n19106), .A3(n19113), .ZN(n16135) );
  OAI21_X1 U15457 ( .B1(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n16144), .A(
        n16135), .ZN(n19100) );
  AOI21_X1 U15458 ( .B1(n19132), .B2(n13677), .A(n19100), .ZN(n12485) );
  INV_X1 U15459 ( .A(n12485), .ZN(n14049) );
  AOI21_X1 U15460 ( .B1(n14055), .B2(n19132), .A(n14049), .ZN(n16119) );
  OAI21_X1 U15461 ( .B1(n16144), .B2(n16117), .A(n16119), .ZN(n14964) );
  OR3_X1 U15462 ( .A1(n14927), .A2(n14883), .A3(n14893), .ZN(n12486) );
  NAND2_X1 U15463 ( .A1(n12485), .A2(n16144), .ZN(n15296) );
  OAI21_X1 U15464 ( .B1(n14964), .B2(n12486), .A(n15296), .ZN(n14869) );
  NAND2_X1 U15465 ( .A1(n12487), .A2(n14873), .ZN(n14868) );
  NAND2_X1 U15466 ( .A1(n14869), .A2(n14868), .ZN(n14861) );
  AND2_X1 U15467 ( .A1(n19132), .A2(n12488), .ZN(n12489) );
  AOI211_X1 U15468 ( .C1(n19132), .C2(n12491), .A(n12490), .B(n14836), .ZN(
        n14805) );
  INV_X1 U15469 ( .A(n15296), .ZN(n14986) );
  OAI21_X1 U15470 ( .B1(n15932), .B2(n19112), .A(n10129), .ZN(n12493) );
  NAND2_X1 U15471 ( .A1(n12495), .A2(n12494), .ZN(n12496) );
  AOI21_X1 U15472 ( .B1(n14191), .B2(n16122), .A(n12496), .ZN(n12497) );
  OAI21_X1 U15473 ( .B1(n14193), .B2(n19110), .A(n12497), .ZN(P2_U3015) );
  NOR2_X1 U15474 ( .A1(n11991), .A2(n16152), .ZN(n12500) );
  NAND2_X1 U15475 ( .A1(n12502), .A2(n12500), .ZN(n19088) );
  AOI21_X1 U15476 ( .B1(n12944), .B2(n14821), .A(n14700), .ZN(n14824) );
  NOR2_X1 U15477 ( .A1(n13728), .A2(n16152), .ZN(n12501) );
  NAND2_X1 U15478 ( .A1(n12502), .A2(n12501), .ZN(n12992) );
  INV_X1 U15479 ( .A(n12992), .ZN(n12503) );
  NOR2_X2 U15480 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19752) );
  OR2_X1 U15481 ( .A1(n19752), .A2(n15042), .ZN(n19765) );
  NAND2_X1 U15482 ( .A1(n19765), .A2(n18715), .ZN(n12504) );
  AND2_X1 U15483 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19766) );
  AOI21_X1 U15484 ( .B1(n12506), .B2(n12945), .A(n12505), .ZN(n14817) );
  INV_X1 U15485 ( .A(n14817), .ZN(n14598) );
  AND2_X1 U15486 ( .A1(n18715), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n12533) );
  INV_X1 U15487 ( .A(n12533), .ZN(n12529) );
  NAND2_X1 U15488 ( .A1(n19221), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n12507) );
  NAND2_X1 U15489 ( .A1(n12529), .A2(n12507), .ZN(n14166) );
  NAND2_X1 U15490 ( .A1(n14565), .A2(n19080), .ZN(n12509) );
  INV_X1 U15491 ( .A(n19093), .ZN(n16001) );
  NOR2_X1 U15492 ( .A1(n16114), .A2(n19731), .ZN(n14816) );
  AOI21_X1 U15493 ( .B1(n16001), .B2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .A(
        n14816), .ZN(n12508) );
  OAI211_X1 U15494 ( .C1(n16072), .C2(n14598), .A(n12509), .B(n12508), .ZN(
        n12510) );
  AOI21_X1 U15495 ( .B1(n14824), .B2(n16068), .A(n12510), .ZN(n12511) );
  NAND2_X1 U15496 ( .A1(n9649), .A2(n12533), .ZN(n12516) );
  OAI21_X1 U15497 ( .B1(n11434), .B2(n18715), .A(n19594), .ZN(n12530) );
  NAND2_X1 U15498 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n19590) );
  INV_X1 U15499 ( .A(n19590), .ZN(n12512) );
  AND2_X1 U15500 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n12512), .ZN(
        n12513) );
  NAND2_X1 U15501 ( .A1(n12513), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n19591) );
  INV_X1 U15502 ( .A(n12513), .ZN(n12520) );
  NAND2_X1 U15503 ( .A1(n19757), .A2(n12520), .ZN(n12514) );
  AND3_X1 U15504 ( .A1(n19591), .A2(n19752), .A3(n12514), .ZN(n19489) );
  AOI21_X1 U15505 ( .B1(n12530), .B2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n19489), .ZN(n12515) );
  AND2_X1 U15506 ( .A1(n11434), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n13042) );
  NAND2_X1 U15507 ( .A1(n13042), .A2(n19796), .ZN(n12768) );
  NOR2_X1 U15508 ( .A1(n12768), .A2(n19161), .ZN(n12517) );
  NAND2_X1 U15509 ( .A1(n12542), .A2(n12517), .ZN(n13083) );
  AND2_X2 U15510 ( .A1(n12518), .A2(n13083), .ZN(n13076) );
  NAND2_X1 U15511 ( .A1(n12519), .A2(n12533), .ZN(n12523) );
  NAND2_X1 U15512 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19455) );
  NAND2_X1 U15513 ( .A1(n19455), .A2(n19764), .ZN(n12521) );
  AND2_X1 U15514 ( .A1(n12521), .A2(n12520), .ZN(n13801) );
  AOI22_X1 U15515 ( .A1(n12530), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B1(
        n19752), .B2(n13801), .ZN(n12522) );
  NAND2_X1 U15516 ( .A1(n12523), .A2(n12522), .ZN(n12526) );
  INV_X1 U15517 ( .A(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12524) );
  NOR2_X1 U15518 ( .A1(n12768), .A2(n12524), .ZN(n12525) );
  AOI22_X1 U15519 ( .A1(n12530), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B1(
        n19752), .B2(n19783), .ZN(n12528) );
  INV_X1 U15520 ( .A(n12768), .ZN(n12791) );
  NAND2_X1 U15521 ( .A1(n12791), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n12534) );
  NAND2_X1 U15522 ( .A1(n12530), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n12531) );
  NAND2_X1 U15523 ( .A1(n19773), .A2(n19783), .ZN(n19364) );
  AND2_X1 U15524 ( .A1(n19455), .A2(n19364), .ZN(n19304) );
  NAND2_X1 U15525 ( .A1(n19752), .A2(n19304), .ZN(n19427) );
  NAND2_X1 U15526 ( .A1(n12531), .A2(n19427), .ZN(n12532) );
  NAND2_X1 U15527 ( .A1(n13073), .A2(n13072), .ZN(n12537) );
  INV_X1 U15528 ( .A(n15038), .ZN(n12535) );
  NAND2_X1 U15529 ( .A1(n12535), .A2(n12534), .ZN(n12536) );
  NAND2_X1 U15530 ( .A1(n12538), .A2(n10128), .ZN(n12540) );
  NAND2_X1 U15531 ( .A1(n12540), .A2(n12539), .ZN(n13077) );
  NAND2_X1 U15532 ( .A1(n11420), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n12541) );
  AND2_X1 U15533 ( .A1(n14169), .A2(n13517), .ZN(n12549) );
  AND2_X1 U15534 ( .A1(n12543), .A2(n13366), .ZN(n12548) );
  AND2_X1 U15535 ( .A1(n18948), .A2(n18949), .ZN(n12547) );
  NAND2_X1 U15536 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13241) );
  AND2_X1 U15537 ( .A1(n13237), .A2(n9740), .ZN(n12546) );
  NOR2_X1 U15538 ( .A1(n12768), .A2(n12545), .ZN(n13234) );
  INV_X1 U15539 ( .A(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12551) );
  INV_X1 U15540 ( .A(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n19606) );
  OAI22_X1 U15541 ( .A1(n12551), .A2(n11686), .B1(n11687), .B2(n19606), .ZN(
        n12552) );
  INV_X1 U15542 ( .A(n12552), .ZN(n12560) );
  AOI22_X1 U15543 ( .A1(P2_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n12671), .B1(
        n11788), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n12559) );
  INV_X1 U15544 ( .A(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n12555) );
  NAND2_X1 U15545 ( .A1(n9670), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n12554) );
  NAND2_X1 U15546 ( .A1(n9652), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(
        n12553) );
  OAI211_X1 U15547 ( .C1(n12675), .C2(n12555), .A(n12554), .B(n12553), .ZN(
        n12556) );
  INV_X1 U15548 ( .A(n12556), .ZN(n12558) );
  AOI22_X1 U15549 ( .A1(n11694), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n13591), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12557) );
  NAND4_X1 U15550 ( .A1(n12560), .A2(n12559), .A3(n12558), .A4(n12557), .ZN(
        n12566) );
  AOI22_X1 U15551 ( .A1(P2_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n9623), .B1(
        n11740), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n12564) );
  AOI22_X1 U15552 ( .A1(P2_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n11741), .B1(
        n11668), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n12563) );
  AOI22_X1 U15553 ( .A1(P2_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n11673), .B1(
        n11720), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12562) );
  NAND2_X1 U15554 ( .A1(n12662), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n12561) );
  NAND4_X1 U15555 ( .A1(n12564), .A2(n12563), .A3(n12562), .A4(n12561), .ZN(
        n12565) );
  NOR2_X1 U15556 ( .A1(n12566), .A2(n12565), .ZN(n18940) );
  OAI22_X1 U15557 ( .A1(n12569), .A2(n11686), .B1(n11687), .B2(n12568), .ZN(
        n12570) );
  INV_X1 U15558 ( .A(n12570), .ZN(n12578) );
  AOI22_X1 U15559 ( .A1(P2_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n12671), .B1(
        n11788), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n12577) );
  NAND2_X1 U15560 ( .A1(n9670), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n12572) );
  NAND2_X1 U15561 ( .A1(n9652), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n12571) );
  OAI211_X1 U15562 ( .C1(n12675), .C2(n12573), .A(n12572), .B(n12571), .ZN(
        n12574) );
  INV_X1 U15563 ( .A(n12574), .ZN(n12576) );
  AOI22_X1 U15564 ( .A1(n11694), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n13591), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12575) );
  NAND4_X1 U15565 ( .A1(n12578), .A2(n12577), .A3(n12576), .A4(n12575), .ZN(
        n12584) );
  AOI22_X1 U15566 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n11834), .B1(
        n11740), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12582) );
  AOI22_X1 U15567 ( .A1(P2_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n11741), .B1(
        n11668), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n12581) );
  AOI22_X1 U15568 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n11673), .B1(
        n11720), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12580) );
  NAND2_X1 U15569 ( .A1(n12662), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n12579) );
  NAND4_X1 U15570 ( .A1(n12582), .A2(n12581), .A3(n12580), .A4(n12579), .ZN(
        n12583) );
  NOR2_X1 U15571 ( .A1(n12584), .A2(n12583), .ZN(n13710) );
  INV_X1 U15572 ( .A(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n12586) );
  INV_X1 U15573 ( .A(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12585) );
  OAI22_X1 U15574 ( .A1(n12586), .A2(n11686), .B1(n11687), .B2(n12585), .ZN(
        n12587) );
  INV_X1 U15575 ( .A(n12587), .ZN(n12595) );
  AOI22_X1 U15576 ( .A1(P2_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n12671), .B1(
        n11788), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n12594) );
  INV_X1 U15577 ( .A(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n12590) );
  NAND2_X1 U15578 ( .A1(n9670), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(
        n12589) );
  NAND2_X1 U15579 ( .A1(n9652), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(
        n12588) );
  OAI211_X1 U15580 ( .C1(n12675), .C2(n12590), .A(n12589), .B(n12588), .ZN(
        n12591) );
  INV_X1 U15581 ( .A(n12591), .ZN(n12593) );
  AOI22_X1 U15582 ( .A1(n11694), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n13591), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12592) );
  NAND4_X1 U15583 ( .A1(n12595), .A2(n12594), .A3(n12593), .A4(n12592), .ZN(
        n12601) );
  AOI22_X1 U15584 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n9623), .B1(
        n11740), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12599) );
  AOI22_X1 U15585 ( .A1(P2_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n11741), .B1(
        n11668), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n12598) );
  AOI22_X1 U15586 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n11673), .B1(
        n11720), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12597) );
  NAND2_X1 U15587 ( .A1(n11742), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(
        n12596) );
  NAND4_X1 U15588 ( .A1(n12599), .A2(n12598), .A3(n12597), .A4(n12596), .ZN(
        n12600) );
  OR2_X1 U15589 ( .A1(n12601), .A2(n12600), .ZN(n13740) );
  OAI22_X1 U15590 ( .A1(n12602), .A2(n11686), .B1(n11687), .B2(n19625), .ZN(
        n12603) );
  INV_X1 U15591 ( .A(n12603), .ZN(n12610) );
  AOI22_X1 U15592 ( .A1(P2_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n12671), .B1(
        n11788), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12609) );
  NAND2_X1 U15593 ( .A1(n9670), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(
        n12605) );
  NAND2_X1 U15594 ( .A1(n9652), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(
        n12604) );
  OAI211_X1 U15595 ( .C1(n12675), .C2(n11253), .A(n12605), .B(n12604), .ZN(
        n12606) );
  INV_X1 U15596 ( .A(n12606), .ZN(n12608) );
  AOI22_X1 U15597 ( .A1(n11694), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n13591), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12607) );
  NAND4_X1 U15598 ( .A1(n12610), .A2(n12609), .A3(n12608), .A4(n12607), .ZN(
        n12616) );
  AOI22_X1 U15599 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n11834), .B1(
        n11740), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12614) );
  AOI22_X1 U15600 ( .A1(P2_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n11741), .B1(
        n11668), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12613) );
  AOI22_X1 U15601 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n11673), .B1(
        n11720), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12612) );
  NAND2_X1 U15602 ( .A1(n12662), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n12611) );
  NAND4_X1 U15603 ( .A1(n12614), .A2(n12613), .A3(n12612), .A4(n12611), .ZN(
        n12615) );
  OR2_X1 U15604 ( .A1(n12616), .A2(n12615), .ZN(n13845) );
  INV_X1 U15605 ( .A(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12618) );
  INV_X1 U15606 ( .A(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12617) );
  OAI22_X1 U15607 ( .A1(n12618), .A2(n11686), .B1(n11687), .B2(n12617), .ZN(
        n12619) );
  INV_X1 U15608 ( .A(n12619), .ZN(n12627) );
  AOI22_X1 U15609 ( .A1(P2_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n12671), .B1(
        n11788), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n12626) );
  INV_X1 U15610 ( .A(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n12622) );
  NAND2_X1 U15611 ( .A1(n9670), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(
        n12621) );
  NAND2_X1 U15612 ( .A1(n9652), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(
        n12620) );
  OAI211_X1 U15613 ( .C1(n12675), .C2(n12622), .A(n12621), .B(n12620), .ZN(
        n12623) );
  INV_X1 U15614 ( .A(n12623), .ZN(n12625) );
  AOI22_X1 U15615 ( .A1(n11694), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n13591), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12624) );
  NAND4_X1 U15616 ( .A1(n12627), .A2(n12626), .A3(n12625), .A4(n12624), .ZN(
        n12633) );
  AOI22_X1 U15617 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n11834), .B1(
        n11740), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12631) );
  AOI22_X1 U15618 ( .A1(P2_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n11741), .B1(
        n11668), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n12630) );
  AOI22_X1 U15619 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n11673), .B1(
        n11720), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12629) );
  NAND2_X1 U15620 ( .A1(n11742), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n12628) );
  NAND4_X1 U15621 ( .A1(n12631), .A2(n12630), .A3(n12629), .A4(n12628), .ZN(
        n12632) );
  NOR2_X1 U15622 ( .A1(n12633), .A2(n12632), .ZN(n15941) );
  INV_X1 U15623 ( .A(n15941), .ZN(n12634) );
  OAI22_X1 U15624 ( .A1(n12636), .A2(n11686), .B1(n11687), .B2(n12635), .ZN(
        n12637) );
  INV_X1 U15625 ( .A(n12637), .ZN(n12645) );
  AOI22_X1 U15626 ( .A1(P2_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n12671), .B1(
        n11788), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12644) );
  NAND2_X1 U15627 ( .A1(n9670), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(
        n12639) );
  NAND2_X1 U15628 ( .A1(n9652), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(
        n12638) );
  OAI211_X1 U15629 ( .C1(n12675), .C2(n12640), .A(n12639), .B(n12638), .ZN(
        n12641) );
  INV_X1 U15630 ( .A(n12641), .ZN(n12643) );
  AOI22_X1 U15631 ( .A1(n11694), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n13591), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12642) );
  NAND4_X1 U15632 ( .A1(n12645), .A2(n12644), .A3(n12643), .A4(n12642), .ZN(
        n12651) );
  AOI22_X1 U15633 ( .A1(P2_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n9623), .B1(
        n11740), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12649) );
  AOI22_X1 U15634 ( .A1(P2_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n11741), .B1(
        n11668), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12648) );
  AOI22_X1 U15635 ( .A1(P2_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n11673), .B1(
        n11720), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12647) );
  NAND2_X1 U15636 ( .A1(n12662), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n12646) );
  NAND4_X1 U15637 ( .A1(n12649), .A2(n12648), .A3(n12647), .A4(n12646), .ZN(
        n12650) );
  NAND2_X1 U15638 ( .A1(n9735), .A2(n10120), .ZN(n14077) );
  OAI22_X1 U15639 ( .A1(n12652), .A2(n11686), .B1(n11687), .B2(n19644), .ZN(
        n12653) );
  INV_X1 U15640 ( .A(n12653), .ZN(n12661) );
  AOI22_X1 U15641 ( .A1(P2_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n12671), .B1(
        n11788), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12660) );
  NAND2_X1 U15642 ( .A1(n9670), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(
        n12655) );
  NAND2_X1 U15643 ( .A1(n9652), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(
        n12654) );
  OAI211_X1 U15644 ( .C1(n12675), .C2(n12656), .A(n12655), .B(n12654), .ZN(
        n12657) );
  INV_X1 U15645 ( .A(n12657), .ZN(n12659) );
  AOI22_X1 U15646 ( .A1(n11694), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n13591), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12658) );
  NAND4_X1 U15647 ( .A1(n12661), .A2(n12660), .A3(n12659), .A4(n12658), .ZN(
        n12668) );
  AOI22_X1 U15648 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n11834), .B1(
        n11740), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12666) );
  AOI22_X1 U15649 ( .A1(P2_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n11741), .B1(
        n11668), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12665) );
  AOI22_X1 U15650 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n11673), .B1(
        n11720), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12664) );
  NAND2_X1 U15651 ( .A1(n12662), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(
        n12663) );
  NAND4_X1 U15652 ( .A1(n12666), .A2(n12665), .A3(n12664), .A4(n12663), .ZN(
        n12667) );
  NOR2_X1 U15653 ( .A1(n12668), .A2(n12667), .ZN(n15937) );
  NOR2_X2 U15654 ( .A1(n14077), .A2(n15937), .ZN(n15935) );
  INV_X1 U15655 ( .A(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n12669) );
  INV_X1 U15656 ( .A(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n19655) );
  OAI22_X1 U15657 ( .A1(n12669), .A2(n11686), .B1(n11687), .B2(n19655), .ZN(
        n12670) );
  INV_X1 U15658 ( .A(n12670), .ZN(n12680) );
  AOI22_X1 U15659 ( .A1(P2_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n12671), .B1(
        n11740), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n12679) );
  INV_X1 U15660 ( .A(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n12674) );
  NAND2_X1 U15661 ( .A1(n9670), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(
        n12673) );
  NAND2_X1 U15662 ( .A1(n9652), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(
        n12672) );
  OAI211_X1 U15663 ( .C1(n12675), .C2(n12674), .A(n12673), .B(n12672), .ZN(
        n12676) );
  INV_X1 U15664 ( .A(n12676), .ZN(n12678) );
  AOI22_X1 U15665 ( .A1(n11694), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n13591), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12677) );
  NAND4_X1 U15666 ( .A1(n12680), .A2(n12679), .A3(n12678), .A4(n12677), .ZN(
        n12686) );
  AOI22_X1 U15667 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n9623), .B1(
        n11788), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12684) );
  AOI22_X1 U15668 ( .A1(P2_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n11741), .B1(
        n12662), .B2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12683) );
  AOI22_X1 U15669 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n11673), .B1(
        n11720), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12682) );
  NAND2_X1 U15670 ( .A1(n11668), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(
        n12681) );
  NAND4_X1 U15671 ( .A1(n12684), .A2(n12683), .A3(n12682), .A4(n12681), .ZN(
        n12685) );
  NOR2_X1 U15672 ( .A1(n12686), .A2(n12685), .ZN(n12706) );
  INV_X1 U15673 ( .A(n12706), .ZN(n12705) );
  AOI22_X1 U15674 ( .A1(n12841), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n9643), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n12696) );
  AOI22_X1 U15675 ( .A1(n12842), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12838), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n12695) );
  AND2_X1 U15676 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n12689) );
  OR2_X1 U15677 ( .A1(n12689), .A2(n12688), .ZN(n12847) );
  INV_X1 U15678 ( .A(n12847), .ZN(n12825) );
  NAND2_X1 U15679 ( .A1(n9644), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n12692) );
  NAND2_X1 U15680 ( .A1(n9646), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n12691) );
  AND3_X1 U15681 ( .A1(n12825), .A2(n12692), .A3(n12691), .ZN(n12694) );
  AOI22_X1 U15682 ( .A1(n13593), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n12845), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n12693) );
  NAND4_X1 U15683 ( .A1(n12696), .A2(n12695), .A3(n12694), .A4(n12693), .ZN(
        n12704) );
  AOI22_X1 U15684 ( .A1(n12841), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n11279), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12702) );
  AOI22_X1 U15685 ( .A1(n12842), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n12838), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12701) );
  AOI22_X1 U15686 ( .A1(n12845), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n12846), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12700) );
  NAND2_X1 U15687 ( .A1(n13593), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n12698) );
  NAND2_X1 U15688 ( .A1(n11656), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n12697) );
  AND3_X1 U15689 ( .A1(n12698), .A2(n12847), .A3(n12697), .ZN(n12699) );
  NAND4_X1 U15690 ( .A1(n12702), .A2(n12701), .A3(n12700), .A4(n12699), .ZN(
        n12703) );
  NAND2_X1 U15691 ( .A1(n12704), .A2(n12703), .ZN(n12728) );
  INV_X1 U15692 ( .A(n12728), .ZN(n12709) );
  NAND2_X1 U15693 ( .A1(n12705), .A2(n12709), .ZN(n12725) );
  OAI21_X1 U15694 ( .B1(n12068), .B2(n12728), .A(n12706), .ZN(n12707) );
  OAI21_X1 U15695 ( .B1(n12068), .B2(n12725), .A(n12707), .ZN(n12729) );
  XNOR2_X1 U15696 ( .A(n15935), .B(n12708), .ZN(n14689) );
  NAND2_X1 U15697 ( .A1(n12068), .A2(n12709), .ZN(n14688) );
  AOI22_X1 U15698 ( .A1(n12842), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n9643), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n12716) );
  AOI22_X1 U15699 ( .A1(n12841), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n12838), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12715) );
  NAND2_X1 U15700 ( .A1(n9644), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n12712) );
  NAND2_X1 U15701 ( .A1(n9646), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n12711) );
  AND3_X1 U15702 ( .A1(n12825), .A2(n12712), .A3(n12711), .ZN(n12714) );
  AOI22_X1 U15703 ( .A1(n13593), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n12845), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12713) );
  NAND4_X1 U15704 ( .A1(n12716), .A2(n12715), .A3(n12714), .A4(n12713), .ZN(
        n12724) );
  AOI22_X1 U15705 ( .A1(n12842), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n11279), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12722) );
  AOI22_X1 U15706 ( .A1(n12841), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n12838), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n12721) );
  AOI22_X1 U15707 ( .A1(n13593), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n12845), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12720) );
  NAND2_X1 U15708 ( .A1(n12690), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n12718) );
  NAND2_X1 U15709 ( .A1(n9646), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n12717) );
  AND3_X1 U15710 ( .A1(n12718), .A2(n12847), .A3(n12717), .ZN(n12719) );
  NAND4_X1 U15711 ( .A1(n12722), .A2(n12721), .A3(n12720), .A4(n12719), .ZN(
        n12723) );
  AND2_X1 U15712 ( .A1(n12724), .A2(n12723), .ZN(n12727) );
  INV_X1 U15713 ( .A(n12725), .ZN(n12726) );
  NAND2_X1 U15714 ( .A1(n12726), .A2(n12727), .ZN(n12731) );
  OAI211_X1 U15715 ( .C1(n12727), .C2(n12726), .A(n12791), .B(n12731), .ZN(
        n14628) );
  NAND2_X1 U15716 ( .A1(n12068), .A2(n12727), .ZN(n14630) );
  NOR3_X1 U15717 ( .A1(n12729), .A2(n12728), .A3(n14630), .ZN(n12730) );
  INV_X1 U15718 ( .A(n12731), .ZN(n12746) );
  AOI22_X1 U15719 ( .A1(n12842), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n9643), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n12737) );
  AOI22_X1 U15720 ( .A1(n12841), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n12838), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12736) );
  NAND2_X1 U15721 ( .A1(n9637), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(
        n12733) );
  NAND2_X1 U15722 ( .A1(n9646), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(
        n12732) );
  AND3_X1 U15723 ( .A1(n12825), .A2(n12733), .A3(n12732), .ZN(n12735) );
  AOI22_X1 U15724 ( .A1(n13593), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n12845), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n12734) );
  NAND4_X1 U15725 ( .A1(n12737), .A2(n12736), .A3(n12735), .A4(n12734), .ZN(
        n12745) );
  AOI22_X1 U15726 ( .A1(n12842), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n9643), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12743) );
  AOI22_X1 U15727 ( .A1(n9642), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n12838), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12742) );
  AOI22_X1 U15728 ( .A1(n13593), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n12845), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12741) );
  NAND2_X1 U15729 ( .A1(n12846), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(
        n12739) );
  NAND2_X1 U15730 ( .A1(n9646), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(
        n12738) );
  AND3_X1 U15731 ( .A1(n12739), .A2(n12847), .A3(n12738), .ZN(n12740) );
  NAND4_X1 U15732 ( .A1(n12743), .A2(n12742), .A3(n12741), .A4(n12740), .ZN(
        n12744) );
  AND2_X1 U15733 ( .A1(n12745), .A2(n12744), .ZN(n12748) );
  NAND2_X1 U15734 ( .A1(n12746), .A2(n12748), .ZN(n12769) );
  OAI211_X1 U15735 ( .C1(n12746), .C2(n12748), .A(n12791), .B(n12769), .ZN(
        n12751) );
  XNOR2_X1 U15736 ( .A(n12750), .B(n12747), .ZN(n14624) );
  INV_X1 U15737 ( .A(n12748), .ZN(n12749) );
  NOR2_X1 U15738 ( .A1(n19796), .A2(n12749), .ZN(n14623) );
  NAND2_X1 U15739 ( .A1(n14624), .A2(n14623), .ZN(n14622) );
  INV_X1 U15740 ( .A(n12750), .ZN(n12752) );
  AOI22_X1 U15741 ( .A1(n12842), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n9643), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n12759) );
  AOI22_X1 U15742 ( .A1(n12841), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n12838), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12758) );
  NAND2_X1 U15743 ( .A1(n12690), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(
        n12755) );
  NAND2_X1 U15744 ( .A1(n9646), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(
        n12754) );
  AND3_X1 U15745 ( .A1(n12825), .A2(n12755), .A3(n12754), .ZN(n12757) );
  AOI22_X1 U15746 ( .A1(n13593), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n12845), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n12756) );
  NAND4_X1 U15747 ( .A1(n12759), .A2(n12758), .A3(n12757), .A4(n12756), .ZN(
        n12767) );
  AOI22_X1 U15748 ( .A1(n12842), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n11279), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12765) );
  AOI22_X1 U15749 ( .A1(n9642), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n12838), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12764) );
  AOI22_X1 U15750 ( .A1(n13593), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n12845), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12763) );
  NAND2_X1 U15751 ( .A1(n12690), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(
        n12761) );
  NAND2_X1 U15752 ( .A1(n9646), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(
        n12760) );
  AND3_X1 U15753 ( .A1(n12761), .A2(n12847), .A3(n12760), .ZN(n12762) );
  NAND4_X1 U15754 ( .A1(n12765), .A2(n12764), .A3(n12763), .A4(n12762), .ZN(
        n12766) );
  NAND2_X1 U15755 ( .A1(n12767), .A2(n12766), .ZN(n12771) );
  AOI21_X1 U15756 ( .B1(n12769), .B2(n12771), .A(n12768), .ZN(n12770) );
  OR2_X1 U15757 ( .A1(n12769), .A2(n12771), .ZN(n12790) );
  INV_X1 U15758 ( .A(n12771), .ZN(n12772) );
  NAND2_X1 U15759 ( .A1(n12068), .A2(n12772), .ZN(n14618) );
  NOR2_X2 U15760 ( .A1(n14617), .A2(n12774), .ZN(n12796) );
  INV_X1 U15761 ( .A(n12796), .ZN(n12794) );
  AOI22_X1 U15762 ( .A1(n12842), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n11279), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n12780) );
  AOI22_X1 U15763 ( .A1(n9642), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n12838), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12779) );
  NAND2_X1 U15764 ( .A1(n12846), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(
        n12776) );
  NAND2_X1 U15765 ( .A1(n9646), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(
        n12775) );
  AND3_X1 U15766 ( .A1(n12825), .A2(n12776), .A3(n12775), .ZN(n12778) );
  AOI22_X1 U15767 ( .A1(n13593), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n12845), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12777) );
  NAND4_X1 U15768 ( .A1(n12780), .A2(n12779), .A3(n12778), .A4(n12777), .ZN(
        n12788) );
  AOI22_X1 U15769 ( .A1(n12842), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n11279), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12786) );
  AOI22_X1 U15770 ( .A1(n12841), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n12838), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12785) );
  AOI22_X1 U15771 ( .A1(n13593), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n12845), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12784) );
  NAND2_X1 U15772 ( .A1(n9644), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(
        n12782) );
  NAND2_X1 U15773 ( .A1(n9646), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n12781) );
  AND3_X1 U15774 ( .A1(n12782), .A2(n12847), .A3(n12781), .ZN(n12783) );
  NAND4_X1 U15775 ( .A1(n12786), .A2(n12785), .A3(n12784), .A4(n12783), .ZN(
        n12787) );
  NAND2_X1 U15776 ( .A1(n12788), .A2(n12787), .ZN(n12789) );
  INV_X1 U15777 ( .A(n12789), .ZN(n12798) );
  INV_X1 U15778 ( .A(n12790), .ZN(n12792) );
  OR2_X1 U15779 ( .A1(n12790), .A2(n12789), .ZN(n14599) );
  OAI211_X1 U15780 ( .C1(n12798), .C2(n12792), .A(n14599), .B(n12791), .ZN(
        n12795) );
  NAND2_X1 U15781 ( .A1(n12796), .A2(n12795), .ZN(n12797) );
  NAND2_X1 U15782 ( .A1(n12068), .A2(n12798), .ZN(n14606) );
  NOR2_X2 U15783 ( .A1(n14607), .A2(n14606), .ZN(n14605) );
  INV_X1 U15784 ( .A(n14600), .ZN(n12813) );
  AOI22_X1 U15785 ( .A1(n12842), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n11279), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n12804) );
  AOI22_X1 U15786 ( .A1(n9642), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n12838), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12803) );
  NAND2_X1 U15787 ( .A1(n12690), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(
        n12800) );
  NAND2_X1 U15788 ( .A1(n9646), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(
        n12799) );
  AND3_X1 U15789 ( .A1(n12825), .A2(n12800), .A3(n12799), .ZN(n12802) );
  AOI22_X1 U15790 ( .A1(n13593), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n12845), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12801) );
  NAND4_X1 U15791 ( .A1(n12804), .A2(n12803), .A3(n12802), .A4(n12801), .ZN(
        n12812) );
  AOI22_X1 U15792 ( .A1(n12842), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n9643), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12810) );
  AOI22_X1 U15793 ( .A1(n12841), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n12838), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12809) );
  AOI22_X1 U15794 ( .A1(n13593), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n12845), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12808) );
  NAND2_X1 U15795 ( .A1(n12690), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(
        n12806) );
  NAND2_X1 U15796 ( .A1(n9646), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(
        n12805) );
  AND3_X1 U15797 ( .A1(n12806), .A2(n12847), .A3(n12805), .ZN(n12807) );
  NAND4_X1 U15798 ( .A1(n12810), .A2(n12809), .A3(n12808), .A4(n12807), .ZN(
        n12811) );
  AND2_X1 U15799 ( .A1(n12812), .A2(n12811), .ZN(n14601) );
  NAND2_X1 U15800 ( .A1(n19796), .A2(n14601), .ZN(n12814) );
  NOR2_X1 U15801 ( .A1(n14599), .A2(n12814), .ZN(n12833) );
  INV_X1 U15802 ( .A(n12816), .ZN(n12822) );
  AOI22_X1 U15803 ( .A1(n11279), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n12838), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12821) );
  AOI22_X1 U15804 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n12845), .B1(
        n13593), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12820) );
  NAND2_X1 U15805 ( .A1(n12846), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(
        n12818) );
  NAND2_X1 U15806 ( .A1(n9646), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(
        n12817) );
  AND3_X1 U15807 ( .A1(n12818), .A2(n12847), .A3(n12817), .ZN(n12819) );
  NAND4_X1 U15808 ( .A1(n12822), .A2(n12821), .A3(n12820), .A4(n12819), .ZN(
        n12831) );
  AOI22_X1 U15809 ( .A1(n12842), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n9643), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12829) );
  AOI22_X1 U15810 ( .A1(n12841), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n12838), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12828) );
  NAND2_X1 U15811 ( .A1(n9637), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(
        n12824) );
  NAND2_X1 U15812 ( .A1(n9646), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(
        n12823) );
  AND3_X1 U15813 ( .A1(n12825), .A2(n12824), .A3(n12823), .ZN(n12827) );
  AOI22_X1 U15814 ( .A1(n13593), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n12845), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12826) );
  NAND4_X1 U15815 ( .A1(n12829), .A2(n12828), .A3(n12827), .A4(n12826), .ZN(
        n12830) );
  AND2_X1 U15816 ( .A1(n12831), .A2(n12830), .ZN(n12832) );
  NAND2_X1 U15817 ( .A1(n12833), .A2(n12832), .ZN(n12834) );
  OAI21_X1 U15818 ( .B1(n12833), .B2(n12832), .A(n12834), .ZN(n14594) );
  INV_X1 U15819 ( .A(n12834), .ZN(n12835) );
  NOR2_X1 U15820 ( .A1(n14593), .A2(n12835), .ZN(n12856) );
  AOI22_X1 U15821 ( .A1(n9642), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B1(n9643), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n12837) );
  AOI22_X1 U15822 ( .A1(n12842), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n9646), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12836) );
  NAND2_X1 U15823 ( .A1(n12837), .A2(n12836), .ZN(n12854) );
  AOI21_X1 U15824 ( .B1(n12838), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .A(
        n12847), .ZN(n12840) );
  AOI22_X1 U15825 ( .A1(n13593), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n12845), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n12839) );
  OAI211_X1 U15826 ( .C1(n11280), .C2(n19655), .A(n12840), .B(n12839), .ZN(
        n12853) );
  AOI22_X1 U15827 ( .A1(n12841), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n11279), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n12844) );
  AOI22_X1 U15828 ( .A1(n12842), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n12838), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12843) );
  NAND2_X1 U15829 ( .A1(n12844), .A2(n12843), .ZN(n12852) );
  AOI22_X1 U15830 ( .A1(n13593), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n12845), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12850) );
  NAND2_X1 U15831 ( .A1(n9646), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(
        n12849) );
  NAND2_X1 U15832 ( .A1(n12846), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(
        n12848) );
  NAND4_X1 U15833 ( .A1(n12850), .A2(n12849), .A3(n12848), .A4(n12847), .ZN(
        n12851) );
  OAI22_X1 U15834 ( .A1(n12854), .A2(n12853), .B1(n12852), .B2(n12851), .ZN(
        n12855) );
  XNOR2_X1 U15835 ( .A(n12856), .B(n12855), .ZN(n14196) );
  NAND2_X1 U15836 ( .A1(n13635), .A2(n12857), .ZN(n13055) );
  NAND2_X1 U15837 ( .A1(n13055), .A2(n12858), .ZN(n12860) );
  NAND2_X1 U15838 ( .A1(n12860), .A2(n12859), .ZN(n12863) );
  AND2_X1 U15839 ( .A1(n12861), .A2(n15424), .ZN(n13627) );
  NAND2_X1 U15840 ( .A1(n19804), .A2(n13627), .ZN(n12862) );
  NAND2_X1 U15841 ( .A1(n18995), .A2(n12864), .ZN(n19002) );
  NAND2_X1 U15842 ( .A1(n18995), .A2(n12865), .ZN(n14691) );
  NOR4_X1 U15843 ( .A1(P2_ADDRESS_REG_15__SCAN_IN), .A2(
        P2_ADDRESS_REG_14__SCAN_IN), .A3(P2_ADDRESS_REG_12__SCAN_IN), .A4(
        P2_ADDRESS_REG_11__SCAN_IN), .ZN(n12869) );
  NOR4_X1 U15844 ( .A1(P2_ADDRESS_REG_20__SCAN_IN), .A2(
        P2_ADDRESS_REG_18__SCAN_IN), .A3(P2_ADDRESS_REG_17__SCAN_IN), .A4(
        P2_ADDRESS_REG_16__SCAN_IN), .ZN(n12868) );
  NOR4_X1 U15845 ( .A1(P2_ADDRESS_REG_6__SCAN_IN), .A2(
        P2_ADDRESS_REG_5__SCAN_IN), .A3(P2_ADDRESS_REG_4__SCAN_IN), .A4(
        P2_ADDRESS_REG_3__SCAN_IN), .ZN(n12867) );
  NOR4_X1 U15846 ( .A1(P2_ADDRESS_REG_10__SCAN_IN), .A2(
        P2_ADDRESS_REG_9__SCAN_IN), .A3(P2_ADDRESS_REG_8__SCAN_IN), .A4(
        P2_ADDRESS_REG_7__SCAN_IN), .ZN(n12866) );
  NAND4_X1 U15847 ( .A1(n12869), .A2(n12868), .A3(n12867), .A4(n12866), .ZN(
        n12874) );
  NOR4_X1 U15848 ( .A1(P2_ADDRESS_REG_1__SCAN_IN), .A2(
        P2_ADDRESS_REG_0__SCAN_IN), .A3(P2_ADDRESS_REG_19__SCAN_IN), .A4(
        P2_ADDRESS_REG_13__SCAN_IN), .ZN(n12872) );
  NOR4_X1 U15849 ( .A1(P2_ADDRESS_REG_24__SCAN_IN), .A2(
        P2_ADDRESS_REG_23__SCAN_IN), .A3(P2_ADDRESS_REG_22__SCAN_IN), .A4(
        P2_ADDRESS_REG_21__SCAN_IN), .ZN(n12871) );
  NOR4_X1 U15850 ( .A1(P2_ADDRESS_REG_28__SCAN_IN), .A2(
        P2_ADDRESS_REG_27__SCAN_IN), .A3(P2_ADDRESS_REG_26__SCAN_IN), .A4(
        P2_ADDRESS_REG_25__SCAN_IN), .ZN(n12870) );
  INV_X1 U15851 ( .A(P2_ADDRESS_REG_2__SCAN_IN), .ZN(n19687) );
  NAND4_X1 U15852 ( .A1(n12872), .A2(n12871), .A3(n12870), .A4(n19687), .ZN(
        n12873) );
  OAI21_X1 U15853 ( .B1(n12874), .B2(n12873), .A(P2_ADDRESS_REG_29__SCAN_IN), 
        .ZN(n13331) );
  INV_X1 U15854 ( .A(n13571), .ZN(n13118) );
  AOI22_X1 U15855 ( .A1(n13571), .A2(BUF1_REG_14__SCAN_IN), .B1(
        BUF2_REG_14__SCAN_IN), .B2(n13118), .ZN(n18976) );
  INV_X1 U15856 ( .A(P2_EAX_REG_30__SCAN_IN), .ZN(n13158) );
  OAI22_X1 U15857 ( .A1(n14691), .A2(n18976), .B1(n13158), .B2(n18995), .ZN(
        n12875) );
  AOI21_X1 U15858 ( .B1(n14806), .B2(n19027), .A(n12875), .ZN(n12878) );
  AND2_X1 U15859 ( .A1(n18995), .A2(n12876), .ZN(n13038) );
  AOI22_X1 U15860 ( .A1(n18965), .A2(BUF2_REG_30__SCAN_IN), .B1(n18964), .B2(
        BUF1_REG_30__SCAN_IN), .ZN(n12877) );
  OAI21_X1 U15861 ( .B1(n14196), .B2(n19002), .A(n12879), .ZN(P2_U2889) );
  OR2_X1 U15862 ( .A1(n12881), .A2(n19946), .ZN(n15348) );
  NOR2_X1 U15863 ( .A1(n15348), .A2(n19820), .ZN(n12882) );
  NAND2_X1 U15864 ( .A1(n15349), .A2(n12882), .ZN(n12996) );
  NOR2_X1 U15865 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20725) );
  NAND2_X1 U15866 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n20725), .ZN(n15368) );
  NAND2_X1 U15867 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n20597), .ZN(n12883) );
  OAI22_X1 U15868 ( .A1(n20597), .A2(n15368), .B1(n12883), .B2(n10404), .ZN(
        n12884) );
  INV_X2 U15869 ( .A(n20050), .ZN(n20043) );
  OR2_X1 U15870 ( .A1(n12884), .A2(n20043), .ZN(n12885) );
  INV_X1 U15871 ( .A(n12886), .ZN(n12887) );
  NAND2_X1 U15872 ( .A1(n12887), .A2(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n12888) );
  XNOR2_X1 U15873 ( .A(n12888), .B(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n13664) );
  AND2_X1 U15874 ( .A1(n13664), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n12889) );
  AOI22_X1 U15875 ( .A1(n12897), .A2(P1_EBX_REG_30__SCAN_IN), .B1(
        P1_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n10881), .ZN(n14201) );
  MUX2_X1 U15876 ( .A(n12890), .B(n14200), .S(P1_EBX_REG_27__SCAN_IN), .Z(
        n12891) );
  NAND2_X1 U15877 ( .A1(n12891), .A2(n10114), .ZN(n14224) );
  INV_X1 U15878 ( .A(P1_EBX_REG_28__SCAN_IN), .ZN(n14316) );
  NAND2_X1 U15879 ( .A1(n10953), .A2(n12892), .ZN(n12893) );
  OAI211_X1 U15880 ( .C1(n10881), .C2(P1_EBX_REG_28__SCAN_IN), .A(n12893), .B(
        n14200), .ZN(n12894) );
  NAND2_X1 U15881 ( .A1(n12895), .A2(n12894), .ZN(n14313) );
  OR2_X1 U15882 ( .A1(n10881), .A2(P1_EBX_REG_29__SCAN_IN), .ZN(n12896) );
  OAI21_X1 U15883 ( .B1(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n12897), .A(
        n12896), .ZN(n14199) );
  MUX2_X1 U15884 ( .A(n12896), .B(n14199), .S(n14200), .Z(n14210) );
  AOI22_X1 U15885 ( .A1(n12897), .A2(P1_EBX_REG_31__SCAN_IN), .B1(
        P1_INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n10881), .ZN(n12898) );
  XNOR2_X1 U15886 ( .A(n12899), .B(n12898), .ZN(n14549) );
  AND2_X1 U15887 ( .A1(n20728), .A2(n20891), .ZN(n15363) );
  NAND2_X1 U15888 ( .A1(P1_EBX_REG_31__SCAN_IN), .A2(n14299), .ZN(n12900) );
  NOR2_X1 U15889 ( .A1(n15363), .A2(n12900), .ZN(n12901) );
  AND2_X1 U15890 ( .A1(P1_REIP_REG_30__SCAN_IN), .A2(P1_REIP_REG_29__SCAN_IN), 
        .ZN(n12906) );
  INV_X1 U15891 ( .A(P1_STATE_REG_0__SCAN_IN), .ZN(n20604) );
  NAND2_X1 U15892 ( .A1(n20604), .A2(n12902), .ZN(n15405) );
  NAND2_X1 U15893 ( .A1(n20096), .A2(n15405), .ZN(n13383) );
  AND2_X1 U15894 ( .A1(n13383), .A2(n15363), .ZN(n12907) );
  NOR2_X1 U15895 ( .A1(n20086), .A2(n14296), .ZN(n12903) );
  NAND2_X1 U15896 ( .A1(n19922), .A2(n19875), .ZN(n19930) );
  INV_X1 U15897 ( .A(P1_REIP_REG_26__SCAN_IN), .ZN(n20660) );
  INV_X1 U15898 ( .A(P1_REIP_REG_24__SCAN_IN), .ZN(n20656) );
  INV_X1 U15899 ( .A(P1_REIP_REG_14__SCAN_IN), .ZN(n20637) );
  INV_X1 U15900 ( .A(P1_REIP_REG_7__SCAN_IN), .ZN(n20629) );
  INV_X1 U15901 ( .A(P1_REIP_REG_1__SCAN_IN), .ZN(n20707) );
  INV_X1 U15902 ( .A(P1_REIP_REG_4__SCAN_IN), .ZN(n20621) );
  INV_X1 U15903 ( .A(P1_REIP_REG_3__SCAN_IN), .ZN(n20620) );
  INV_X1 U15904 ( .A(P1_REIP_REG_2__SCAN_IN), .ZN(n20824) );
  NOR4_X1 U15905 ( .A1(n20707), .A2(n20621), .A3(n20620), .A4(n20824), .ZN(
        n19876) );
  NAND3_X1 U15906 ( .A1(n19876), .A2(P1_REIP_REG_6__SCAN_IN), .A3(
        P1_REIP_REG_5__SCAN_IN), .ZN(n19852) );
  NOR2_X1 U15907 ( .A1(n20629), .A2(n19852), .ZN(n15537) );
  NAND2_X1 U15908 ( .A1(P1_REIP_REG_8__SCAN_IN), .A2(n15537), .ZN(n13657) );
  NAND4_X1 U15909 ( .A1(P1_REIP_REG_12__SCAN_IN), .A2(P1_REIP_REG_11__SCAN_IN), 
        .A3(P1_REIP_REG_10__SCAN_IN), .A4(P1_REIP_REG_9__SCAN_IN), .ZN(n14125)
         );
  NOR2_X1 U15910 ( .A1(n13657), .A2(n14125), .ZN(n14128) );
  NAND2_X1 U15911 ( .A1(P1_REIP_REG_13__SCAN_IN), .A2(n14128), .ZN(n14104) );
  NOR2_X1 U15912 ( .A1(n20637), .A2(n14104), .ZN(n14285) );
  NAND3_X1 U15913 ( .A1(P1_REIP_REG_17__SCAN_IN), .A2(P1_REIP_REG_16__SCAN_IN), 
        .A3(P1_REIP_REG_15__SCAN_IN), .ZN(n14245) );
  NAND3_X1 U15914 ( .A1(P1_REIP_REG_20__SCAN_IN), .A2(P1_REIP_REG_19__SCAN_IN), 
        .A3(P1_REIP_REG_18__SCAN_IN), .ZN(n14247) );
  NAND3_X1 U15915 ( .A1(P1_REIP_REG_21__SCAN_IN), .A2(P1_REIP_REG_23__SCAN_IN), 
        .A3(P1_REIP_REG_22__SCAN_IN), .ZN(n12904) );
  NOR3_X1 U15916 ( .A1(n14245), .A2(n14247), .A3(n12904), .ZN(n15473) );
  NAND2_X1 U15917 ( .A1(n14285), .A2(n15473), .ZN(n15480) );
  NOR2_X1 U15918 ( .A1(n20656), .A2(n15480), .ZN(n15474) );
  NAND2_X1 U15919 ( .A1(P1_REIP_REG_25__SCAN_IN), .A2(n15474), .ZN(n15461) );
  NOR2_X1 U15920 ( .A1(n20660), .A2(n15461), .ZN(n14227) );
  AND2_X1 U15921 ( .A1(P1_REIP_REG_27__SCAN_IN), .A2(n14227), .ZN(n15450) );
  NAND2_X1 U15922 ( .A1(P1_REIP_REG_28__SCAN_IN), .A2(n15450), .ZN(n15451) );
  INV_X1 U15923 ( .A(n15451), .ZN(n14211) );
  NAND2_X1 U15924 ( .A1(n19922), .A2(n14211), .ZN(n12905) );
  NAND2_X1 U15925 ( .A1(n19930), .A2(n12905), .ZN(n15456) );
  OAI21_X1 U15926 ( .B1(n12906), .B2(n19875), .A(n15456), .ZN(n14203) );
  INV_X1 U15927 ( .A(P1_EBX_REG_31__SCAN_IN), .ZN(n20794) );
  INV_X1 U15928 ( .A(n12907), .ZN(n12910) );
  OR2_X1 U15929 ( .A1(n20086), .A2(P1_EBX_REG_31__SCAN_IN), .ZN(n12908) );
  AOI21_X1 U15930 ( .B1(n20722), .B2(n12908), .A(n14296), .ZN(n12909) );
  NAND2_X1 U15931 ( .A1(n19935), .A2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n12912) );
  NOR3_X1 U15932 ( .A1(n19875), .A2(n15451), .A3(n14217), .ZN(n14204) );
  INV_X1 U15933 ( .A(P1_REIP_REG_31__SCAN_IN), .ZN(n12926) );
  NAND3_X1 U15934 ( .A1(n14204), .A2(P1_REIP_REG_30__SCAN_IN), .A3(n12926), 
        .ZN(n12911) );
  OAI211_X1 U15935 ( .C1(n20794), .C2(n19867), .A(n12912), .B(n12911), .ZN(
        n12913) );
  AOI21_X1 U15936 ( .B1(P1_REIP_REG_31__SCAN_IN), .B2(n14203), .A(n12913), 
        .ZN(n12914) );
  NAND2_X1 U15937 ( .A1(n12917), .A2(n12916), .ZN(P1_U2809) );
  NAND2_X1 U15938 ( .A1(n12918), .A2(n15645), .ZN(n12932) );
  NOR2_X1 U15939 ( .A1(n14445), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n12922) );
  INV_X1 U15940 ( .A(n12919), .ZN(n12920) );
  NOR2_X1 U15941 ( .A1(n20050), .A2(n12926), .ZN(n14554) );
  INV_X1 U15942 ( .A(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n12927) );
  NOR2_X1 U15943 ( .A1(n20039), .A2(n12927), .ZN(n12928) );
  AOI211_X1 U15944 ( .C1(n15635), .C2(n13664), .A(n14554), .B(n12928), .ZN(
        n12929) );
  INV_X1 U15945 ( .A(n12930), .ZN(n12931) );
  NAND2_X1 U15946 ( .A1(n12932), .A2(n12931), .ZN(P1_U2968) );
  NAND2_X1 U15947 ( .A1(n12936), .A2(n12937), .ZN(n12933) );
  INV_X1 U15948 ( .A(n12934), .ZN(n12935) );
  AOI21_X1 U15949 ( .B1(n12936), .B2(n12938), .A(n12937), .ZN(n12939) );
  XOR2_X1 U15950 ( .A(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .B(n12940), .Z(
        n12941) );
  NAND2_X1 U15951 ( .A1(n12958), .A2(n12942), .ZN(n12957) );
  OAI21_X1 U15952 ( .B1(n12943), .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n12944), .ZN(n12963) );
  INV_X1 U15953 ( .A(n12963), .ZN(n12955) );
  AOI21_X1 U15954 ( .B1(n14829), .B2(n14818), .A(n14836), .ZN(n14822) );
  INV_X1 U15955 ( .A(n12945), .ZN(n12946) );
  INV_X1 U15956 ( .A(n14573), .ZN(n12948) );
  OAI21_X1 U15957 ( .B1(n14653), .B2(n12949), .A(n12948), .ZN(n14648) );
  NAND2_X1 U15958 ( .A1(n19081), .A2(P2_REIP_REG_28__SCAN_IN), .ZN(n12959) );
  OAI21_X1 U15959 ( .B1(n16128), .B2(n14648), .A(n12959), .ZN(n12950) );
  AOI21_X1 U15960 ( .B1(n15892), .B2(n19131), .A(n12950), .ZN(n12952) );
  NAND3_X1 U15961 ( .A1(n14818), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A3(
        n14829), .ZN(n12951) );
  OAI211_X1 U15962 ( .C1(n14822), .C2(n12953), .A(n12952), .B(n12951), .ZN(
        n12954) );
  AOI21_X1 U15963 ( .B1(n12955), .B2(n16122), .A(n12954), .ZN(n12956) );
  NAND2_X1 U15964 ( .A1(n12957), .A2(n12956), .ZN(P2_U3018) );
  NAND2_X1 U15965 ( .A1(n12958), .A2(n16066), .ZN(n12967) );
  OAI21_X1 U15966 ( .B1(n19093), .B2(n15888), .A(n12959), .ZN(n12962) );
  NOR2_X1 U15967 ( .A1(n12960), .A2(n16063), .ZN(n12961) );
  AOI211_X1 U15968 ( .C1(n19090), .C2(n15892), .A(n12962), .B(n12961), .ZN(
        n12965) );
  NAND2_X1 U15969 ( .A1(n12967), .A2(n12966), .ZN(P2_U2986) );
  INV_X1 U15970 ( .A(P1_W_R_N_REG_SCAN_IN), .ZN(n20716) );
  NOR3_X1 U15971 ( .A1(P1_BE_N_REG_0__SCAN_IN), .A2(P1_BE_N_REG_1__SCAN_IN), 
        .A3(n20716), .ZN(n12969) );
  NOR4_X1 U15972 ( .A1(P1_BE_N_REG_2__SCAN_IN), .A2(P1_BE_N_REG_3__SCAN_IN), 
        .A3(P1_D_C_N_REG_SCAN_IN), .A4(P1_ADS_N_REG_SCAN_IN), .ZN(n12968) );
  NAND4_X1 U15973 ( .A1(n20085), .A2(P1_M_IO_N_REG_SCAN_IN), .A3(n12969), .A4(
        n12968), .ZN(U214) );
  INV_X1 U15974 ( .A(P2_W_R_N_REG_SCAN_IN), .ZN(n19785) );
  NOR2_X1 U15975 ( .A1(P2_BE_N_REG_1__SCAN_IN), .A2(n19785), .ZN(n12971) );
  NOR4_X1 U15976 ( .A1(P2_BE_N_REG_2__SCAN_IN), .A2(P2_BE_N_REG_3__SCAN_IN), 
        .A3(P2_D_C_N_REG_SCAN_IN), .A4(P2_ADS_N_REG_SCAN_IN), .ZN(n12970) );
  INV_X1 U15977 ( .A(P2_BE_N_REG_0__SCAN_IN), .ZN(n19741) );
  NAND4_X1 U15978 ( .A1(P2_M_IO_N_REG_SCAN_IN), .A2(n12971), .A3(n12970), .A4(
        n19741), .ZN(n12972) );
  NOR2_X1 U15979 ( .A1(n13331), .A2(n12972), .ZN(n16248) );
  NAND2_X1 U15980 ( .A1(n16248), .A2(U214), .ZN(U212) );
  NOR2_X1 U15981 ( .A1(P2_ADDRESS_REG_29__SCAN_IN), .A2(n12972), .ZN(n16332)
         );
  AOI211_X1 U15982 ( .C1(n15977), .C2(n12974), .A(n12973), .B(n18890), .ZN(
        n12987) );
  INV_X1 U15983 ( .A(P2_EBX_REG_23__SCAN_IN), .ZN(n12975) );
  OAI22_X1 U15984 ( .A1(n12976), .A2(n18923), .B1(n12975), .B2(n18929), .ZN(
        n12986) );
  OAI22_X1 U15985 ( .A1(n15984), .A2(n18935), .B1(n11581), .B2(n18932), .ZN(
        n12985) );
  NAND2_X1 U15986 ( .A1(n12977), .A2(n12978), .ZN(n12979) );
  NAND2_X1 U15987 ( .A1(n14632), .A2(n12979), .ZN(n15978) );
  NAND2_X1 U15988 ( .A1(n12980), .A2(n12981), .ZN(n12982) );
  AND2_X1 U15989 ( .A1(n14677), .A2(n12982), .ZN(n14888) );
  INV_X1 U15990 ( .A(n14888), .ZN(n12983) );
  OAI22_X1 U15991 ( .A1(n15978), .A2(n18924), .B1(n18928), .B2(n12983), .ZN(
        n12984) );
  OR4_X1 U15992 ( .A1(n12987), .A2(n12986), .A3(n12985), .A4(n12984), .ZN(
        P2_U2832) );
  INV_X1 U15993 ( .A(n12988), .ZN(n12989) );
  INV_X1 U15994 ( .A(n13152), .ZN(n13057) );
  NAND2_X1 U15995 ( .A1(n12989), .A2(n13057), .ZN(n13559) );
  INV_X1 U15996 ( .A(n13559), .ZN(n18936) );
  INV_X1 U15997 ( .A(P2_MEMORYFETCH_REG_SCAN_IN), .ZN(n19814) );
  INV_X1 U15998 ( .A(n13025), .ZN(n13024) );
  NAND2_X1 U15999 ( .A1(n19752), .A2(n13649), .ZN(n18714) );
  OAI211_X1 U16000 ( .C1(n18936), .C2(n19814), .A(n13024), .B(n18714), .ZN(
        P2_U2814) );
  NOR2_X1 U16001 ( .A1(n19804), .A2(P2_READREQUEST_REG_SCAN_IN), .ZN(n12990)
         );
  AOI22_X1 U16002 ( .A1(n12990), .A2(n18714), .B1(n19798), .B2(n19804), .ZN(
        P2_U3612) );
  NOR4_X1 U16003 ( .A1(n13631), .A2(n13641), .A3(n13627), .A4(n13056), .ZN(
        n12991) );
  NOR2_X1 U16004 ( .A1(n12991), .A2(n16152), .ZN(n19793) );
  OAI21_X1 U16005 ( .B1(n19793), .B2(n12993), .A(n12992), .ZN(P2_U2819) );
  INV_X1 U16006 ( .A(n20700), .ZN(n20541) );
  OAI21_X1 U16007 ( .B1(P1_STATE2_REG_1__SCAN_IN), .B2(n20541), .A(n15404), 
        .ZN(n12995) );
  AOI21_X1 U16008 ( .B1(P1_MEMORYFETCH_REG_SCAN_IN), .B2(n12996), .A(n12995), 
        .ZN(n12994) );
  INV_X1 U16009 ( .A(n12994), .ZN(P1_U2801) );
  NOR2_X1 U16010 ( .A1(P1_READREQUEST_REG_SCAN_IN), .A2(n12995), .ZN(n12997)
         );
  AND2_X1 U16011 ( .A1(n12997), .A2(n12996), .ZN(n12999) );
  OAI22_X1 U16012 ( .A1(n12999), .A2(n12998), .B1(n12997), .B2(n20726), .ZN(
        P1_U3487) );
  OAI21_X1 U16013 ( .B1(n13512), .B2(n14163), .A(n13000), .ZN(n13001) );
  XNOR2_X1 U16014 ( .A(n13001), .B(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n19123) );
  INV_X1 U16015 ( .A(n19123), .ZN(n13010) );
  OAI21_X1 U16016 ( .B1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n13003), .A(
        n13002), .ZN(n19126) );
  INV_X1 U16017 ( .A(n19126), .ZN(n13004) );
  NOR2_X1 U16018 ( .A1(n16114), .A2(n19685), .ZN(n19129) );
  AOI21_X1 U16019 ( .B1(n16068), .B2(n13004), .A(n19129), .ZN(n13006) );
  NAND2_X1 U16020 ( .A1(n19080), .A2(n13007), .ZN(n13005) );
  OAI211_X1 U16021 ( .C1(n13007), .C2(n19093), .A(n13006), .B(n13005), .ZN(
        n13008) );
  AOI21_X1 U16022 ( .B1(n19090), .B2(n19130), .A(n13008), .ZN(n13009) );
  OAI21_X1 U16023 ( .B1(n19088), .B2(n13010), .A(n13009), .ZN(P2_U3013) );
  OAI21_X1 U16024 ( .B1(n13014), .B2(n13013), .A(n13012), .ZN(n19111) );
  INV_X1 U16025 ( .A(n19111), .ZN(n13022) );
  NAND2_X1 U16026 ( .A1(n19080), .A2(n13462), .ZN(n13016) );
  INV_X1 U16027 ( .A(P2_REIP_REG_2__SCAN_IN), .ZN(n13015) );
  OR2_X1 U16028 ( .A1(n16114), .A2(n13015), .ZN(n19118) );
  OAI211_X1 U16029 ( .C1(n13017), .C2(n19093), .A(n13016), .B(n19118), .ZN(
        n13021) );
  NAND2_X1 U16030 ( .A1(n13019), .A2(n13018), .ZN(n19107) );
  AND3_X1 U16031 ( .A1(n19108), .A2(n19107), .A3(n16066), .ZN(n13020) );
  AOI211_X1 U16032 ( .C1(n16068), .C2(n13022), .A(n13021), .B(n13020), .ZN(
        n13023) );
  OAI21_X1 U16033 ( .B1(n13011), .B2(n16072), .A(n13023), .ZN(P2_U3012) );
  INV_X1 U16034 ( .A(P2_LWORD_REG_14__SCAN_IN), .ZN(n13027) );
  NAND3_X1 U16035 ( .A1(n13025), .A2(n19796), .A3(n15424), .ZN(n13348) );
  NOR2_X1 U16036 ( .A1(n13348), .A2(n18976), .ZN(n13030) );
  AOI21_X1 U16037 ( .B1(P2_EAX_REG_14__SCAN_IN), .B2(n19077), .A(n13030), .ZN(
        n13026) );
  OAI21_X1 U16038 ( .B1(n13250), .B2(n13027), .A(n13026), .ZN(P2_U2981) );
  INV_X1 U16039 ( .A(P2_UWORD_REG_1__SCAN_IN), .ZN(n13029) );
  AOI22_X1 U16040 ( .A1(n13571), .A2(BUF1_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n13331), .ZN(n19150) );
  NOR2_X1 U16041 ( .A1(n13348), .A2(n19150), .ZN(n13257) );
  AOI21_X1 U16042 ( .B1(n19077), .B2(P2_EAX_REG_17__SCAN_IN), .A(n13257), .ZN(
        n13028) );
  OAI21_X1 U16043 ( .B1(n13250), .B2(n13029), .A(n13028), .ZN(P2_U2953) );
  INV_X1 U16044 ( .A(P2_UWORD_REG_14__SCAN_IN), .ZN(n13032) );
  AOI21_X1 U16045 ( .B1(n19077), .B2(P2_EAX_REG_30__SCAN_IN), .A(n13030), .ZN(
        n13031) );
  OAI21_X1 U16046 ( .B1(n13250), .B2(n13032), .A(n13031), .ZN(P2_U2966) );
  INV_X1 U16047 ( .A(P2_LWORD_REG_7__SCAN_IN), .ZN(n13034) );
  AOI22_X1 U16048 ( .A1(n13571), .A2(BUF1_REG_7__SCAN_IN), .B1(
        BUF2_REG_7__SCAN_IN), .B2(n13118), .ZN(n19178) );
  NOR2_X1 U16049 ( .A1(n13348), .A2(n19178), .ZN(n13263) );
  AOI21_X1 U16050 ( .B1(n19077), .B2(P2_EAX_REG_7__SCAN_IN), .A(n13263), .ZN(
        n13033) );
  OAI21_X1 U16051 ( .B1(n13250), .B2(n13034), .A(n13033), .ZN(P2_U2974) );
  INV_X1 U16052 ( .A(P2_LWORD_REG_12__SCAN_IN), .ZN(n13037) );
  AOI22_X1 U16053 ( .A1(n13571), .A2(BUF1_REG_12__SCAN_IN), .B1(
        BUF2_REG_12__SCAN_IN), .B2(n13118), .ZN(n18981) );
  INV_X1 U16054 ( .A(n18981), .ZN(n13035) );
  NAND2_X1 U16055 ( .A1(n13120), .A2(n13035), .ZN(n13107) );
  NAND2_X1 U16056 ( .A1(n19077), .A2(P2_EAX_REG_12__SCAN_IN), .ZN(n13036) );
  OAI211_X1 U16057 ( .C1(n13250), .C2(n13037), .A(n13107), .B(n13036), .ZN(
        P2_U2979) );
  INV_X1 U16058 ( .A(n14691), .ZN(n18963) );
  INV_X1 U16059 ( .A(BUF1_REG_0__SCAN_IN), .ZN(n16301) );
  INV_X1 U16060 ( .A(BUF2_REG_0__SCAN_IN), .ZN(n18048) );
  AOI22_X1 U16061 ( .A1(n13571), .A2(n16301), .B1(n18048), .B2(n13331), .ZN(
        n18962) );
  INV_X1 U16062 ( .A(n18962), .ZN(n13727) );
  NOR2_X1 U16063 ( .A1(n13040), .A2(n13039), .ZN(n13041) );
  NOR2_X1 U16064 ( .A1(n11683), .A2(n13041), .ZN(n18926) );
  INV_X1 U16065 ( .A(P2_EAX_REG_0__SCAN_IN), .ZN(n13343) );
  NOR2_X1 U16066 ( .A1(P2_INSTQUEUE_REG_0__0__SCAN_IN), .A2(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n13043) );
  OAI21_X1 U16067 ( .B1(n13044), .B2(n13043), .A(n13042), .ZN(n13045) );
  INV_X1 U16068 ( .A(n13045), .ZN(n13046) );
  NAND2_X1 U16069 ( .A1(n19137), .A2(n18926), .ZN(n19029) );
  OAI211_X1 U16070 ( .C1(n19137), .C2(n18926), .A(n19029), .B(n19031), .ZN(
        n13047) );
  OAI21_X1 U16071 ( .B1(n13343), .B2(n18995), .A(n13047), .ZN(n13048) );
  AOI21_X1 U16072 ( .B1(n19027), .B2(n18926), .A(n13048), .ZN(n13049) );
  OAI21_X1 U16073 ( .B1(n19035), .B2(n13727), .A(n13049), .ZN(P2_U2919) );
  NAND2_X1 U16074 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n19776) );
  NOR2_X1 U16075 ( .A1(n18715), .A2(n19776), .ZN(n16147) );
  INV_X1 U16076 ( .A(n13641), .ZN(n13050) );
  NAND2_X1 U16077 ( .A1(n13050), .A2(n13627), .ZN(n13052) );
  OAI21_X1 U16078 ( .B1(n13631), .B2(n13052), .A(n13051), .ZN(n13053) );
  INV_X1 U16079 ( .A(n13053), .ZN(n13054) );
  AND2_X1 U16080 ( .A1(n13055), .A2(n13054), .ZN(n13060) );
  OR2_X1 U16081 ( .A1(n13635), .A2(n13630), .ZN(n13070) );
  NAND2_X1 U16082 ( .A1(n13057), .A2(n13056), .ZN(n13058) );
  OR2_X1 U16083 ( .A1(n13154), .A2(n13058), .ZN(n13059) );
  OAI22_X1 U16084 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n19594), .B1(n13622), 
        .B2(n16152), .ZN(n13061) );
  AOI21_X1 U16085 ( .B1(P2_FLUSH_REG_SCAN_IN), .B2(n16147), .A(n13061), .ZN(
        n15044) );
  INV_X1 U16086 ( .A(n15044), .ZN(n13067) );
  AND2_X1 U16087 ( .A1(n13063), .A2(n13062), .ZN(n13064) );
  AND2_X1 U16088 ( .A1(n13065), .A2(n13064), .ZN(n13637) );
  NAND3_X1 U16089 ( .A1(n13067), .A2(n15042), .A3(n13637), .ZN(n13066) );
  OAI21_X1 U16090 ( .B1(n13067), .B2(n13643), .A(n13066), .ZN(P2_U3595) );
  INV_X1 U16091 ( .A(n19138), .ZN(n19760) );
  MUX2_X1 U16092 ( .A(n11992), .B(n13011), .S(n18958), .Z(n13071) );
  OAI21_X1 U16093 ( .B1(n19760), .B2(n18952), .A(n13071), .ZN(P2_U2885) );
  INV_X1 U16094 ( .A(n19130), .ZN(n13608) );
  MUX2_X1 U16095 ( .A(n11988), .B(n13608), .S(n18958), .Z(n13074) );
  OAI21_X1 U16096 ( .B1(n18999), .B2(n18952), .A(n13074), .ZN(P2_U2886) );
  MUX2_X1 U16097 ( .A(n11989), .B(n18925), .S(n18958), .Z(n13075) );
  OAI21_X1 U16098 ( .B1(n19779), .B2(n18952), .A(n13075), .ZN(P2_U2887) );
  NAND2_X1 U16099 ( .A1(n15938), .A2(P2_EBX_REG_3__SCAN_IN), .ZN(n13081) );
  NAND2_X1 U16100 ( .A1(n9650), .A2(n18958), .ZN(n13080) );
  OAI211_X1 U16101 ( .C1(n19000), .C2(n18952), .A(n13081), .B(n13080), .ZN(
        P2_U2884) );
  NAND2_X1 U16102 ( .A1(n13082), .A2(n13234), .ZN(n13242) );
  NAND2_X1 U16103 ( .A1(n13242), .A2(n13084), .ZN(n19008) );
  NAND2_X1 U16104 ( .A1(n13086), .A2(n13085), .ZN(n13088) );
  INV_X1 U16105 ( .A(n13087), .ZN(n13134) );
  AND2_X1 U16106 ( .A1(n13088), .A2(n13134), .ZN(n19096) );
  MUX2_X1 U16107 ( .A(P2_EBX_REG_4__SCAN_IN), .B(n19096), .S(n18958), .Z(
        n13089) );
  INV_X1 U16108 ( .A(n13089), .ZN(n13090) );
  OAI21_X1 U16109 ( .B1(n19008), .B2(n18952), .A(n13090), .ZN(P2_U2883) );
  INV_X1 U16110 ( .A(P2_EAX_REG_20__SCAN_IN), .ZN(n13092) );
  INV_X1 U16111 ( .A(n13250), .ZN(n13122) );
  NAND2_X1 U16112 ( .A1(n13122), .A2(P2_UWORD_REG_4__SCAN_IN), .ZN(n13091) );
  OAI22_X1 U16113 ( .A1(n13118), .A2(BUF1_REG_4__SCAN_IN), .B1(
        BUF2_REG_4__SCAN_IN), .B2(n13571), .ZN(n19162) );
  INV_X1 U16114 ( .A(n19162), .ZN(n15955) );
  NAND2_X1 U16115 ( .A1(n13120), .A2(n15955), .ZN(n13123) );
  OAI211_X1 U16116 ( .C1(n13092), .C2(n13347), .A(n13091), .B(n13123), .ZN(
        P2_U2956) );
  INV_X1 U16117 ( .A(P2_EAX_REG_22__SCAN_IN), .ZN(n13094) );
  NAND2_X1 U16118 ( .A1(n13122), .A2(P2_UWORD_REG_6__SCAN_IN), .ZN(n13093) );
  OAI22_X1 U16119 ( .A1(n13331), .A2(BUF1_REG_6__SCAN_IN), .B1(
        BUF2_REG_6__SCAN_IN), .B2(n13571), .ZN(n19172) );
  INV_X1 U16120 ( .A(n19172), .ZN(n15949) );
  NAND2_X1 U16121 ( .A1(n13120), .A2(n15949), .ZN(n13289) );
  OAI211_X1 U16122 ( .C1(n13347), .C2(n13094), .A(n13093), .B(n13289), .ZN(
        P2_U2958) );
  INV_X1 U16123 ( .A(P2_EAX_REG_19__SCAN_IN), .ZN(n13847) );
  NAND2_X1 U16124 ( .A1(n13122), .A2(P2_UWORD_REG_3__SCAN_IN), .ZN(n13096) );
  AOI22_X1 U16125 ( .A1(n13571), .A2(BUF1_REG_3__SCAN_IN), .B1(
        BUF2_REG_3__SCAN_IN), .B2(n13331), .ZN(n19157) );
  INV_X1 U16126 ( .A(n19157), .ZN(n13095) );
  NAND2_X1 U16127 ( .A1(n13120), .A2(n13095), .ZN(n13097) );
  OAI211_X1 U16128 ( .C1(n13847), .C2(n13347), .A(n13096), .B(n13097), .ZN(
        P2_U2955) );
  INV_X1 U16129 ( .A(P2_EAX_REG_3__SCAN_IN), .ZN(n13099) );
  NAND2_X1 U16130 ( .A1(n13122), .A2(P2_LWORD_REG_3__SCAN_IN), .ZN(n13098) );
  OAI211_X1 U16131 ( .C1(n13099), .C2(n13347), .A(n13098), .B(n13097), .ZN(
        P2_U2970) );
  NAND2_X1 U16132 ( .A1(n13122), .A2(P2_UWORD_REG_11__SCAN_IN), .ZN(n13103) );
  INV_X1 U16133 ( .A(BUF2_REG_11__SCAN_IN), .ZN(n13100) );
  NOR2_X1 U16134 ( .A1(n13571), .A2(n13100), .ZN(n13101) );
  AOI21_X1 U16135 ( .B1(BUF1_REG_11__SCAN_IN), .B2(n13571), .A(n13101), .ZN(
        n18983) );
  INV_X1 U16136 ( .A(n18983), .ZN(n13102) );
  NAND2_X1 U16137 ( .A1(n13120), .A2(n13102), .ZN(n13286) );
  OAI211_X1 U16138 ( .C1(n13347), .C2(n14655), .A(n13103), .B(n13286), .ZN(
        P2_U2963) );
  INV_X1 U16139 ( .A(P2_EAX_REG_10__SCAN_IN), .ZN(n19052) );
  NAND2_X1 U16140 ( .A1(n13122), .A2(P2_LWORD_REG_10__SCAN_IN), .ZN(n13106) );
  NAND2_X1 U16141 ( .A1(n13118), .A2(BUF2_REG_10__SCAN_IN), .ZN(n13105) );
  INV_X1 U16142 ( .A(BUF1_REG_10__SCAN_IN), .ZN(n16281) );
  OR2_X1 U16143 ( .A1(n13118), .A2(n16281), .ZN(n13104) );
  NAND2_X1 U16144 ( .A1(n13105), .A2(n13104), .ZN(n18985) );
  NAND2_X1 U16145 ( .A1(n13120), .A2(n18985), .ZN(n19075) );
  OAI211_X1 U16146 ( .C1(n19052), .C2(n13347), .A(n13106), .B(n19075), .ZN(
        P2_U2977) );
  INV_X1 U16147 ( .A(P2_EAX_REG_28__SCAN_IN), .ZN(n20839) );
  NAND2_X1 U16148 ( .A1(n13122), .A2(P2_UWORD_REG_12__SCAN_IN), .ZN(n13108) );
  OAI211_X1 U16149 ( .C1(n13347), .C2(n20839), .A(n13108), .B(n13107), .ZN(
        P2_U2964) );
  INV_X1 U16150 ( .A(P2_EAX_REG_25__SCAN_IN), .ZN(n14670) );
  NAND2_X1 U16151 ( .A1(n13122), .A2(P2_UWORD_REG_9__SCAN_IN), .ZN(n13112) );
  INV_X1 U16152 ( .A(BUF2_REG_9__SCAN_IN), .ZN(n13109) );
  NOR2_X1 U16153 ( .A1(n13571), .A2(n13109), .ZN(n13110) );
  AOI21_X1 U16154 ( .B1(BUF1_REG_9__SCAN_IN), .B2(n13571), .A(n13110), .ZN(
        n18988) );
  INV_X1 U16155 ( .A(n18988), .ZN(n13111) );
  NAND2_X1 U16156 ( .A1(n13120), .A2(n13111), .ZN(n13280) );
  OAI211_X1 U16157 ( .C1(n13347), .C2(n14670), .A(n13112), .B(n13280), .ZN(
        P2_U2961) );
  INV_X1 U16158 ( .A(P2_EAX_REG_8__SCAN_IN), .ZN(n19056) );
  NAND2_X1 U16159 ( .A1(n13122), .A2(P2_LWORD_REG_8__SCAN_IN), .ZN(n13115) );
  NAND2_X1 U16160 ( .A1(n13118), .A2(BUF2_REG_8__SCAN_IN), .ZN(n13114) );
  INV_X1 U16161 ( .A(BUF1_REG_8__SCAN_IN), .ZN(n16285) );
  OR2_X1 U16162 ( .A1(n13331), .A2(n16285), .ZN(n13113) );
  NAND2_X1 U16163 ( .A1(n13114), .A2(n13113), .ZN(n18991) );
  NAND2_X1 U16164 ( .A1(n13120), .A2(n18991), .ZN(n19072) );
  OAI211_X1 U16165 ( .C1(n19056), .C2(n13347), .A(n13115), .B(n19072), .ZN(
        P2_U2975) );
  INV_X1 U16166 ( .A(P2_EAX_REG_29__SCAN_IN), .ZN(n14642) );
  NAND2_X1 U16167 ( .A1(n13122), .A2(P2_UWORD_REG_13__SCAN_IN), .ZN(n13121) );
  INV_X1 U16168 ( .A(BUF1_REG_13__SCAN_IN), .ZN(n13116) );
  NOR2_X1 U16169 ( .A1(n13118), .A2(n13116), .ZN(n13117) );
  AOI21_X1 U16170 ( .B1(n13118), .B2(BUF2_REG_13__SCAN_IN), .A(n13117), .ZN(
        n18978) );
  INV_X1 U16171 ( .A(n18978), .ZN(n13119) );
  NAND2_X1 U16172 ( .A1(n13120), .A2(n13119), .ZN(n13283) );
  OAI211_X1 U16173 ( .C1(n13347), .C2(n14642), .A(n13121), .B(n13283), .ZN(
        P2_U2965) );
  INV_X1 U16174 ( .A(P2_EAX_REG_4__SCAN_IN), .ZN(n13125) );
  NAND2_X1 U16175 ( .A1(n13122), .A2(P2_LWORD_REG_4__SCAN_IN), .ZN(n13124) );
  OAI211_X1 U16176 ( .C1(n13125), .C2(n13347), .A(n13124), .B(n13123), .ZN(
        P2_U2971) );
  OAI21_X1 U16177 ( .B1(n13127), .B2(n13126), .A(n13140), .ZN(n20036) );
  OR2_X1 U16178 ( .A1(n13129), .A2(n13128), .ZN(n13130) );
  NAND2_X1 U16179 ( .A1(n13131), .A2(n13130), .ZN(n20063) );
  AOI22_X1 U16180 ( .A1(n19940), .A2(n20063), .B1(n10965), .B2(
        P1_EBX_REG_1__SCAN_IN), .ZN(n13132) );
  OAI21_X1 U16181 ( .B1(n20036), .B2(n9630), .A(n13132), .ZN(P1_U2871) );
  XOR2_X1 U16182 ( .A(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B(n13242), .Z(n13139)
         );
  NAND2_X1 U16183 ( .A1(n15938), .A2(P2_EBX_REG_5__SCAN_IN), .ZN(n13138) );
  INV_X1 U16184 ( .A(n13133), .ZN(n13135) );
  NAND2_X1 U16185 ( .A1(n13135), .A2(n13134), .ZN(n13136) );
  AND2_X1 U16186 ( .A1(n13136), .A2(n13244), .ZN(n18915) );
  NAND2_X1 U16187 ( .A1(n15948), .A2(n18915), .ZN(n13137) );
  OAI211_X1 U16188 ( .C1(n13139), .C2(n18952), .A(n13138), .B(n13137), .ZN(
        P2_U2882) );
  OAI21_X1 U16189 ( .B1(n9741), .B2(n10378), .A(n13141), .ZN(n14308) );
  AOI21_X1 U16190 ( .B1(n13143), .B2(n13142), .A(n9825), .ZN(n20055) );
  AOI22_X1 U16191 ( .A1(n19940), .A2(n20055), .B1(n10965), .B2(
        P1_EBX_REG_2__SCAN_IN), .ZN(n13144) );
  OAI21_X1 U16192 ( .B1(n14308), .B2(n9630), .A(n13144), .ZN(P1_U2870) );
  NAND2_X1 U16193 ( .A1(n13145), .A2(n20072), .ZN(n13147) );
  NAND2_X1 U16194 ( .A1(n13147), .A2(n13146), .ZN(n20082) );
  OAI21_X1 U16195 ( .B1(n13150), .B2(n13149), .A(n13148), .ZN(n20045) );
  OAI222_X1 U16196 ( .A1(n20082), .A2(n14356), .B1(n19945), .B2(n13151), .C1(
        n9630), .C2(n20045), .ZN(P1_U2872) );
  OR2_X1 U16197 ( .A1(n13152), .A2(n16152), .ZN(n13153) );
  OAI21_X1 U16198 ( .B1(n13154), .B2(n13153), .A(n13347), .ZN(n13155) );
  INV_X1 U16199 ( .A(P2_EAX_REG_21__SCAN_IN), .ZN(n14081) );
  OR2_X1 U16200 ( .A1(n19776), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n19806) );
  AND2_X2 U16201 ( .A1(n19071), .A2(n19806), .ZN(n19067) );
  INV_X1 U16202 ( .A(n19067), .ZN(n19065) );
  INV_X1 U16203 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n20816) );
  INV_X1 U16204 ( .A(P2_UWORD_REG_5__SCAN_IN), .ZN(n13157) );
  OAI222_X1 U16205 ( .A1(n19037), .A2(n14081), .B1(n19065), .B2(n20816), .C1(
        n13157), .C2(n19806), .ZN(P2_U2930) );
  INV_X1 U16206 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n16330) );
  OAI222_X1 U16207 ( .A1(n19037), .A2(n13158), .B1(n19806), .B2(n13032), .C1(
        n19065), .C2(n16330), .ZN(P2_U2921) );
  INV_X1 U16208 ( .A(P2_UWORD_REG_9__SCAN_IN), .ZN(n13159) );
  INV_X1 U16209 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n20802) );
  OAI222_X1 U16210 ( .A1(n19037), .A2(n14670), .B1(n19806), .B2(n13159), .C1(
        n19065), .C2(n20802), .ZN(P2_U2926) );
  OR2_X1 U16211 ( .A1(n12881), .A2(n14298), .ZN(n15328) );
  NOR2_X1 U16212 ( .A1(n15328), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n13314) );
  AOI21_X1 U16213 ( .B1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n13164), .A(
        n13167), .ZN(n13171) );
  MUX2_X1 U16214 ( .A(n13167), .B(n9925), .S(n10142), .Z(n13163) );
  INV_X1 U16215 ( .A(n13395), .ZN(n13162) );
  OR2_X1 U16216 ( .A1(n13161), .A2(n13160), .ZN(n13399) );
  NAND2_X1 U16217 ( .A1(n13162), .A2(n13399), .ZN(n13315) );
  OAI21_X1 U16218 ( .B1(n13164), .B2(n13163), .A(n13315), .ZN(n13170) );
  NAND2_X1 U16219 ( .A1(n10249), .A2(n13174), .ZN(n13166) );
  NOR2_X1 U16220 ( .A1(n13166), .A2(n13165), .ZN(n13317) );
  INV_X1 U16221 ( .A(n10142), .ZN(n13211) );
  AOI21_X1 U16222 ( .B1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n13211), .A(
        n13167), .ZN(n13168) );
  NAND2_X1 U16223 ( .A1(n10318), .A2(n13168), .ZN(n13192) );
  NAND2_X1 U16224 ( .A1(n13317), .A2(n13192), .ZN(n13169) );
  OAI211_X1 U16225 ( .C1(n13171), .C2(n15328), .A(n13170), .B(n13169), .ZN(
        n13190) );
  INV_X1 U16226 ( .A(n20684), .ZN(n20325) );
  NAND2_X1 U16227 ( .A1(n13196), .A2(n10878), .ZN(n13178) );
  OAI21_X1 U16228 ( .B1(n13172), .B2(n10869), .A(n13489), .ZN(n13175) );
  OAI21_X1 U16229 ( .B1(n13175), .B2(n13174), .A(n10256), .ZN(n13176) );
  AND3_X1 U16230 ( .A1(n13178), .A2(n13177), .A3(n13176), .ZN(n13182) );
  INV_X1 U16231 ( .A(n13490), .ZN(n13179) );
  AOI21_X1 U16232 ( .B1(n13179), .B2(n10256), .A(n20086), .ZN(n13180) );
  NAND2_X1 U16233 ( .A1(n13181), .A2(n13180), .ZN(n13199) );
  NAND3_X1 U16234 ( .A1(n13183), .A2(n13182), .A3(n13199), .ZN(n13400) );
  AND2_X1 U16235 ( .A1(n13184), .A2(n13404), .ZN(n13187) );
  NAND4_X1 U16236 ( .A1(n11067), .A2(n13187), .A3(n13185), .A4(n13186), .ZN(
        n13188) );
  NOR2_X1 U16237 ( .A1(n13400), .A2(n13188), .ZN(n14176) );
  NOR2_X1 U16238 ( .A1(n20325), .A2(n14176), .ZN(n13189) );
  AOI211_X1 U16239 ( .C1(n13314), .C2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n13190), .B(n13189), .ZN(n13191) );
  INV_X1 U16240 ( .A(n13191), .ZN(n13419) );
  INV_X1 U16241 ( .A(n14179), .ZN(n13325) );
  AOI22_X1 U16242 ( .A1(n13419), .A2(n15857), .B1(n13192), .B2(n13325), .ZN(
        n13209) );
  INV_X1 U16243 ( .A(n13185), .ZN(n13193) );
  NOR2_X1 U16244 ( .A1(n15328), .A2(n15405), .ZN(n15408) );
  NAND2_X1 U16245 ( .A1(n10881), .A2(n15405), .ZN(n15345) );
  OAI211_X1 U16246 ( .C1(n13193), .C2(n15408), .A(n15345), .B(n20728), .ZN(
        n13194) );
  INV_X1 U16247 ( .A(n13194), .ZN(n13195) );
  NAND2_X1 U16248 ( .A1(n15409), .A2(n13195), .ZN(n13202) );
  INV_X1 U16249 ( .A(n13196), .ZN(n13197) );
  NAND3_X1 U16250 ( .A1(n13199), .A2(n13198), .A3(n13197), .ZN(n13200) );
  AND2_X1 U16251 ( .A1(n13200), .A2(n15348), .ZN(n13381) );
  INV_X1 U16252 ( .A(n13381), .ZN(n13201) );
  OAI211_X1 U16253 ( .C1(n14298), .C2(n13389), .A(n13202), .B(n13201), .ZN(
        n13203) );
  NOR2_X1 U16254 ( .A1(n13382), .A2(n13203), .ZN(n13206) );
  INV_X1 U16255 ( .A(n13204), .ZN(n13205) );
  NAND2_X1 U16256 ( .A1(n13206), .A2(n13205), .ZN(n15331) );
  INV_X1 U16257 ( .A(n15331), .ZN(n13207) );
  NOR2_X1 U16258 ( .A1(n13663), .A2(n20599), .ZN(n15412) );
  NAND2_X1 U16259 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n15412), .ZN(n15870) );
  INV_X1 U16260 ( .A(P1_FLUSH_REG_SCAN_IN), .ZN(n19827) );
  OAI22_X1 U16261 ( .A1(n13207), .A2(n19820), .B1(n15870), .B2(n19827), .ZN(
        n15859) );
  AOI21_X1 U16262 ( .B1(P1_STATE2_REG_3__SCAN_IN), .B2(n20597), .A(n15859), 
        .ZN(n14184) );
  NAND2_X1 U16263 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n14184), .ZN(
        n13208) );
  OAI21_X1 U16264 ( .B1(n13209), .B2(n14184), .A(n13208), .ZN(P1_U3469) );
  INV_X1 U16265 ( .A(n13314), .ZN(n13213) );
  NAND3_X1 U16266 ( .A1(n14177), .A2(n13211), .A3(n13210), .ZN(n13212) );
  OAI211_X1 U16267 ( .C1(n20438), .C2(n14176), .A(n13213), .B(n13212), .ZN(
        n15330) );
  NOR2_X1 U16268 ( .A1(n13663), .A2(n20072), .ZN(n13326) );
  AOI22_X1 U16269 ( .A1(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(n10874), .B2(n12924), .ZN(
        n13327) );
  INV_X1 U16270 ( .A(n13327), .ZN(n13214) );
  AND2_X1 U16271 ( .A1(n13326), .A2(n13214), .ZN(n13216) );
  AOI211_X1 U16272 ( .C1(n15330), .C2(n15857), .A(n13216), .B(n13215), .ZN(
        n13218) );
  NAND2_X1 U16273 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(n14184), .ZN(
        n13217) );
  OAI21_X1 U16274 ( .B1(n13218), .B2(n14184), .A(n13217), .ZN(P1_U3473) );
  INV_X1 U16275 ( .A(P2_EAX_REG_16__SCAN_IN), .ZN(n13346) );
  AOI22_X1 U16276 ( .A1(n9634), .A2(P2_UWORD_REG_0__SCAN_IN), .B1(n19067), 
        .B2(P2_DATAO_REG_16__SCAN_IN), .ZN(n13219) );
  OAI21_X1 U16277 ( .B1(n13346), .B2(n19037), .A(n13219), .ZN(P2_U2935) );
  INV_X1 U16278 ( .A(P2_EAX_REG_18__SCAN_IN), .ZN(n13742) );
  AOI22_X1 U16279 ( .A1(n9634), .A2(P2_UWORD_REG_2__SCAN_IN), .B1(n19067), 
        .B2(P2_DATAO_REG_18__SCAN_IN), .ZN(n13220) );
  OAI21_X1 U16280 ( .B1(n13742), .B2(n19037), .A(n13220), .ZN(P2_U2933) );
  AOI22_X1 U16281 ( .A1(n9634), .A2(P2_UWORD_REG_11__SCAN_IN), .B1(n19067), 
        .B2(P2_DATAO_REG_27__SCAN_IN), .ZN(n13221) );
  OAI21_X1 U16282 ( .B1(n14655), .B2(n19037), .A(n13221), .ZN(P2_U2924) );
  AOI22_X1 U16283 ( .A1(n9634), .A2(P2_UWORD_REG_6__SCAN_IN), .B1(n19067), 
        .B2(P2_DATAO_REG_22__SCAN_IN), .ZN(n13222) );
  OAI21_X1 U16284 ( .B1(n13094), .B2(n19037), .A(n13222), .ZN(P2_U2929) );
  AOI22_X1 U16285 ( .A1(n9634), .A2(P2_UWORD_REG_7__SCAN_IN), .B1(n19067), 
        .B2(P2_DATAO_REG_23__SCAN_IN), .ZN(n13223) );
  OAI21_X1 U16286 ( .B1(n14690), .B2(n19037), .A(n13223), .ZN(P2_U2928) );
  AOI22_X1 U16287 ( .A1(n9634), .A2(P2_UWORD_REG_4__SCAN_IN), .B1(n19067), 
        .B2(P2_DATAO_REG_20__SCAN_IN), .ZN(n13224) );
  OAI21_X1 U16288 ( .B1(n13092), .B2(n19037), .A(n13224), .ZN(P2_U2931) );
  INV_X1 U16289 ( .A(P2_EAX_REG_17__SCAN_IN), .ZN(n13713) );
  AOI22_X1 U16290 ( .A1(n9634), .A2(P2_UWORD_REG_1__SCAN_IN), .B1(n19067), 
        .B2(P2_DATAO_REG_17__SCAN_IN), .ZN(n13225) );
  OAI21_X1 U16291 ( .B1(n13713), .B2(n19037), .A(n13225), .ZN(P2_U2934) );
  AOI22_X1 U16292 ( .A1(n9634), .A2(P2_UWORD_REG_3__SCAN_IN), .B1(n19067), 
        .B2(P2_DATAO_REG_19__SCAN_IN), .ZN(n13226) );
  OAI21_X1 U16293 ( .B1(n13847), .B2(n19037), .A(n13226), .ZN(P2_U2932) );
  NAND2_X1 U16294 ( .A1(n13082), .A2(n13227), .ZN(n13236) );
  INV_X1 U16295 ( .A(n13236), .ZN(n18950) );
  XNOR2_X1 U16296 ( .A(n18950), .B(n18949), .ZN(n13232) );
  INV_X1 U16297 ( .A(n13228), .ZN(n15011) );
  INV_X1 U16298 ( .A(n9746), .ZN(n13229) );
  NAND2_X1 U16299 ( .A1(n9748), .A2(n13229), .ZN(n13230) );
  NAND2_X1 U16300 ( .A1(n15011), .A2(n13230), .ZN(n16062) );
  MUX2_X1 U16301 ( .A(n11429), .B(n16062), .S(n18958), .Z(n13231) );
  OAI21_X1 U16302 ( .B1(n13232), .B2(n18952), .A(n13231), .ZN(P2_U2878) );
  AOI21_X1 U16303 ( .B1(n13233), .B2(n13272), .A(n9746), .ZN(n18875) );
  INV_X1 U16304 ( .A(n18875), .ZN(n14798) );
  AND2_X1 U16305 ( .A1(n13082), .A2(n13234), .ZN(n13235) );
  AND2_X1 U16306 ( .A1(n13235), .A2(n9740), .ZN(n13238) );
  OAI211_X1 U16307 ( .C1(n13238), .C2(n13237), .A(n13236), .B(n15942), .ZN(
        n13240) );
  NAND2_X1 U16308 ( .A1(n15938), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n13239) );
  OAI211_X1 U16309 ( .C1(n14798), .C2(n15938), .A(n13240), .B(n13239), .ZN(
        P2_U2879) );
  NOR2_X1 U16310 ( .A1(n13242), .A2(n19171), .ZN(n13243) );
  OR2_X1 U16311 ( .A1(n13242), .A2(n13241), .ZN(n13271) );
  OAI211_X1 U16312 ( .C1(n13243), .C2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A(
        n15942), .B(n13271), .ZN(n13249) );
  NAND2_X1 U16313 ( .A1(n13245), .A2(n13244), .ZN(n13247) );
  INV_X1 U16314 ( .A(n13273), .ZN(n13246) );
  NAND2_X1 U16315 ( .A1(n13247), .A2(n13246), .ZN(n13837) );
  INV_X1 U16316 ( .A(n13837), .ZN(n18901) );
  NAND2_X1 U16317 ( .A1(n15948), .A2(n18901), .ZN(n13248) );
  OAI211_X1 U16318 ( .C1(n18958), .C2(n18894), .A(n13249), .B(n13248), .ZN(
        P2_U2881) );
  INV_X1 U16319 ( .A(P2_LWORD_REG_5__SCAN_IN), .ZN(n13252) );
  AOI22_X1 U16320 ( .A1(n13571), .A2(BUF1_REG_5__SCAN_IN), .B1(
        BUF2_REG_5__SCAN_IN), .B2(n13331), .ZN(n19168) );
  NOR2_X1 U16321 ( .A1(n13348), .A2(n19168), .ZN(n13255) );
  AOI21_X1 U16322 ( .B1(n19077), .B2(P2_EAX_REG_5__SCAN_IN), .A(n13255), .ZN(
        n13251) );
  OAI21_X1 U16323 ( .B1(n13250), .B2(n13252), .A(n13251), .ZN(P2_U2972) );
  INV_X1 U16324 ( .A(P2_LWORD_REG_2__SCAN_IN), .ZN(n13254) );
  AOI22_X1 U16325 ( .A1(n13571), .A2(BUF1_REG_2__SCAN_IN), .B1(
        BUF2_REG_2__SCAN_IN), .B2(n13331), .ZN(n19025) );
  NOR2_X1 U16326 ( .A1(n13348), .A2(n19025), .ZN(n13260) );
  AOI21_X1 U16327 ( .B1(P2_EAX_REG_2__SCAN_IN), .B2(n19077), .A(n13260), .ZN(
        n13253) );
  OAI21_X1 U16328 ( .B1(n13250), .B2(n13254), .A(n13253), .ZN(P2_U2969) );
  AOI21_X1 U16329 ( .B1(n19077), .B2(P2_EAX_REG_21__SCAN_IN), .A(n13255), .ZN(
        n13256) );
  OAI21_X1 U16330 ( .B1(n13250), .B2(n13157), .A(n13256), .ZN(P2_U2957) );
  INV_X1 U16331 ( .A(P2_LWORD_REG_1__SCAN_IN), .ZN(n13259) );
  AOI21_X1 U16332 ( .B1(P2_EAX_REG_1__SCAN_IN), .B2(n19077), .A(n13257), .ZN(
        n13258) );
  OAI21_X1 U16333 ( .B1(n13250), .B2(n13259), .A(n13258), .ZN(P2_U2968) );
  INV_X1 U16334 ( .A(P2_UWORD_REG_2__SCAN_IN), .ZN(n13262) );
  AOI21_X1 U16335 ( .B1(P2_EAX_REG_18__SCAN_IN), .B2(n19077), .A(n13260), .ZN(
        n13261) );
  OAI21_X1 U16336 ( .B1(n13250), .B2(n13262), .A(n13261), .ZN(P2_U2954) );
  INV_X1 U16337 ( .A(P2_UWORD_REG_7__SCAN_IN), .ZN(n13265) );
  AOI21_X1 U16338 ( .B1(n19077), .B2(P2_EAX_REG_23__SCAN_IN), .A(n13263), .ZN(
        n13264) );
  OAI21_X1 U16339 ( .B1(n13250), .B2(n13265), .A(n13264), .ZN(P2_U2959) );
  INV_X1 U16340 ( .A(n20728), .ZN(n20607) );
  AND2_X1 U16341 ( .A1(n20722), .A2(n20607), .ZN(n13266) );
  MUX2_X1 U16342 ( .A(DATAI_2_), .B(BUF1_REG_2__SCAN_IN), .S(n20085), .Z(
        n14423) );
  NAND2_X1 U16343 ( .A1(n9752), .A2(n14423), .ZN(n13300) );
  AOI22_X1 U16344 ( .A1(n20026), .A2(P1_EAX_REG_18__SCAN_IN), .B1(n20025), 
        .B2(P1_UWORD_REG_2__SCAN_IN), .ZN(n13267) );
  NAND2_X1 U16345 ( .A1(n13300), .A2(n13267), .ZN(P1_U2939) );
  MUX2_X1 U16346 ( .A(DATAI_0_), .B(BUF1_REG_0__SCAN_IN), .S(n20085), .Z(
        n14440) );
  NAND2_X1 U16347 ( .A1(n9752), .A2(n14440), .ZN(n13293) );
  AOI22_X1 U16348 ( .A1(n20026), .A2(P1_EAX_REG_16__SCAN_IN), .B1(n20025), 
        .B2(P1_UWORD_REG_0__SCAN_IN), .ZN(n13268) );
  NAND2_X1 U16349 ( .A1(n13293), .A2(n13268), .ZN(P1_U2937) );
  MUX2_X1 U16350 ( .A(DATAI_3_), .B(BUF1_REG_3__SCAN_IN), .S(n20085), .Z(
        n14418) );
  NAND2_X1 U16351 ( .A1(n9752), .A2(n14418), .ZN(n13302) );
  AOI22_X1 U16352 ( .A1(n20026), .A2(P1_EAX_REG_19__SCAN_IN), .B1(n20025), 
        .B2(P1_UWORD_REG_3__SCAN_IN), .ZN(n13269) );
  NAND2_X1 U16353 ( .A1(n13302), .A2(n13269), .ZN(P1_U2940) );
  MUX2_X1 U16354 ( .A(DATAI_1_), .B(BUF1_REG_1__SCAN_IN), .S(n20085), .Z(
        n14429) );
  NAND2_X1 U16355 ( .A1(n9752), .A2(n14429), .ZN(n13295) );
  AOI22_X1 U16356 ( .A1(n20026), .A2(P1_EAX_REG_17__SCAN_IN), .B1(n20025), 
        .B2(P1_UWORD_REG_1__SCAN_IN), .ZN(n13270) );
  NAND2_X1 U16357 ( .A1(n13295), .A2(n13270), .ZN(P1_U2938) );
  XOR2_X1 U16358 ( .A(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B(n13271), .Z(n13276)
         );
  OAI21_X1 U16359 ( .B1(n13274), .B2(n13273), .A(n13272), .ZN(n18885) );
  MUX2_X1 U16360 ( .A(n11533), .B(n18885), .S(n18958), .Z(n13275) );
  OAI21_X1 U16361 ( .B1(n13276), .B2(n18952), .A(n13275), .ZN(P2_U2880) );
  INV_X1 U16362 ( .A(n9753), .ZN(n13291) );
  INV_X1 U16363 ( .A(P1_EAX_REG_15__SCAN_IN), .ZN(n13278) );
  AOI22_X1 U16364 ( .A1(n20085), .A2(BUF1_REG_15__SCAN_IN), .B1(DATAI_15_), 
        .B2(n20083), .ZN(n14143) );
  INV_X1 U16365 ( .A(P1_LWORD_REG_15__SCAN_IN), .ZN(n13277) );
  OAI222_X1 U16366 ( .A1(n13291), .A2(n13278), .B1(n9664), .B2(n14143), .C1(
        n13277), .C2(n20000), .ZN(P1_U2967) );
  INV_X1 U16367 ( .A(P2_LWORD_REG_9__SCAN_IN), .ZN(n13281) );
  NAND2_X1 U16368 ( .A1(n19077), .A2(P2_EAX_REG_9__SCAN_IN), .ZN(n13279) );
  OAI211_X1 U16369 ( .C1(n13250), .C2(n13281), .A(n13280), .B(n13279), .ZN(
        P2_U2976) );
  INV_X1 U16370 ( .A(P2_LWORD_REG_13__SCAN_IN), .ZN(n13284) );
  NAND2_X1 U16371 ( .A1(n19077), .A2(P2_EAX_REG_13__SCAN_IN), .ZN(n13282) );
  OAI211_X1 U16372 ( .C1(n13250), .C2(n13284), .A(n13283), .B(n13282), .ZN(
        P2_U2980) );
  INV_X1 U16373 ( .A(P2_LWORD_REG_11__SCAN_IN), .ZN(n13287) );
  NAND2_X1 U16374 ( .A1(n19077), .A2(P2_EAX_REG_11__SCAN_IN), .ZN(n13285) );
  OAI211_X1 U16375 ( .C1(n13250), .C2(n13287), .A(n13286), .B(n13285), .ZN(
        P2_U2978) );
  INV_X1 U16376 ( .A(P2_LWORD_REG_6__SCAN_IN), .ZN(n13290) );
  NAND2_X1 U16377 ( .A1(n19077), .A2(P2_EAX_REG_6__SCAN_IN), .ZN(n13288) );
  OAI211_X1 U16378 ( .C1(n13250), .C2(n13290), .A(n13289), .B(n13288), .ZN(
        P2_U2973) );
  AOI22_X1 U16379 ( .A1(n20026), .A2(P1_EAX_REG_0__SCAN_IN), .B1(n20025), .B2(
        P1_LWORD_REG_0__SCAN_IN), .ZN(n13292) );
  NAND2_X1 U16380 ( .A1(n13293), .A2(n13292), .ZN(P1_U2952) );
  AOI22_X1 U16381 ( .A1(n20026), .A2(P1_EAX_REG_1__SCAN_IN), .B1(n20025), .B2(
        P1_LWORD_REG_1__SCAN_IN), .ZN(n13294) );
  NAND2_X1 U16382 ( .A1(n13295), .A2(n13294), .ZN(P1_U2953) );
  MUX2_X1 U16383 ( .A(DATAI_4_), .B(BUF1_REG_4__SCAN_IN), .S(n20085), .Z(
        n14412) );
  NAND2_X1 U16384 ( .A1(n9752), .A2(n14412), .ZN(n13304) );
  AOI22_X1 U16385 ( .A1(n20026), .A2(P1_EAX_REG_20__SCAN_IN), .B1(n20025), 
        .B2(P1_UWORD_REG_4__SCAN_IN), .ZN(n13296) );
  NAND2_X1 U16386 ( .A1(n13304), .A2(n13296), .ZN(P1_U2941) );
  MUX2_X1 U16387 ( .A(DATAI_6_), .B(BUF1_REG_6__SCAN_IN), .S(n20085), .Z(
        n14403) );
  NAND2_X1 U16388 ( .A1(n9752), .A2(n14403), .ZN(n13307) );
  AOI22_X1 U16389 ( .A1(n20026), .A2(P1_EAX_REG_6__SCAN_IN), .B1(n20025), .B2(
        P1_LWORD_REG_6__SCAN_IN), .ZN(n13297) );
  NAND2_X1 U16390 ( .A1(n13307), .A2(n13297), .ZN(P1_U2958) );
  MUX2_X1 U16391 ( .A(DATAI_5_), .B(BUF1_REG_5__SCAN_IN), .S(n20085), .Z(
        n14407) );
  NAND2_X1 U16392 ( .A1(n9752), .A2(n14407), .ZN(n13309) );
  AOI22_X1 U16393 ( .A1(n20026), .A2(P1_EAX_REG_21__SCAN_IN), .B1(n20025), 
        .B2(P1_UWORD_REG_5__SCAN_IN), .ZN(n13298) );
  NAND2_X1 U16394 ( .A1(n13309), .A2(n13298), .ZN(P1_U2942) );
  AOI22_X1 U16395 ( .A1(n20026), .A2(P1_EAX_REG_2__SCAN_IN), .B1(n20025), .B2(
        P1_LWORD_REG_2__SCAN_IN), .ZN(n13299) );
  NAND2_X1 U16396 ( .A1(n13300), .A2(n13299), .ZN(P1_U2954) );
  AOI22_X1 U16397 ( .A1(n20026), .A2(P1_EAX_REG_3__SCAN_IN), .B1(n20025), .B2(
        P1_LWORD_REG_3__SCAN_IN), .ZN(n13301) );
  NAND2_X1 U16398 ( .A1(n13302), .A2(n13301), .ZN(P1_U2955) );
  AOI22_X1 U16399 ( .A1(n20026), .A2(P1_EAX_REG_4__SCAN_IN), .B1(n20025), .B2(
        P1_LWORD_REG_4__SCAN_IN), .ZN(n13303) );
  NAND2_X1 U16400 ( .A1(n13304), .A2(n13303), .ZN(P1_U2956) );
  MUX2_X1 U16401 ( .A(DATAI_7_), .B(BUF1_REG_7__SCAN_IN), .S(n20085), .Z(
        n14399) );
  NAND2_X1 U16402 ( .A1(n9752), .A2(n14399), .ZN(n13311) );
  AOI22_X1 U16403 ( .A1(n20026), .A2(P1_EAX_REG_23__SCAN_IN), .B1(n20025), 
        .B2(P1_UWORD_REG_7__SCAN_IN), .ZN(n13305) );
  NAND2_X1 U16404 ( .A1(n13311), .A2(n13305), .ZN(P1_U2944) );
  AOI22_X1 U16405 ( .A1(n20026), .A2(P1_EAX_REG_22__SCAN_IN), .B1(n20025), 
        .B2(P1_UWORD_REG_6__SCAN_IN), .ZN(n13306) );
  NAND2_X1 U16406 ( .A1(n13307), .A2(n13306), .ZN(P1_U2943) );
  AOI22_X1 U16407 ( .A1(n20026), .A2(P1_EAX_REG_5__SCAN_IN), .B1(n20025), .B2(
        P1_LWORD_REG_5__SCAN_IN), .ZN(n13308) );
  NAND2_X1 U16408 ( .A1(n13309), .A2(n13308), .ZN(P1_U2957) );
  AOI22_X1 U16409 ( .A1(n20026), .A2(P1_EAX_REG_7__SCAN_IN), .B1(n20025), .B2(
        P1_LWORD_REG_7__SCAN_IN), .ZN(n13310) );
  NAND2_X1 U16410 ( .A1(n13311), .A2(n13310), .ZN(P1_U2959) );
  OR2_X1 U16411 ( .A1(n13312), .A2(n14176), .ZN(n13323) );
  NOR2_X1 U16412 ( .A1(n15328), .A2(n9778), .ZN(n13313) );
  MUX2_X1 U16413 ( .A(n13314), .B(n13313), .S(n13329), .Z(n13321) );
  XNOR2_X1 U16414 ( .A(n10142), .B(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13316) );
  NAND2_X1 U16415 ( .A1(n13315), .A2(n13316), .ZN(n13319) );
  INV_X1 U16416 ( .A(n13316), .ZN(n13324) );
  NAND2_X1 U16417 ( .A1(n13317), .A2(n13324), .ZN(n13318) );
  NAND2_X1 U16418 ( .A1(n13319), .A2(n13318), .ZN(n13320) );
  NOR2_X1 U16419 ( .A1(n13321), .A2(n13320), .ZN(n13322) );
  NAND2_X1 U16420 ( .A1(n13323), .A2(n13322), .ZN(n13420) );
  AOI222_X1 U16421 ( .A1(n13420), .A2(n15857), .B1(n13327), .B2(n13326), .C1(
        n13325), .C2(n13324), .ZN(n13328) );
  INV_X1 U16422 ( .A(n14184), .ZN(n15862) );
  MUX2_X1 U16423 ( .A(n13329), .B(n13328), .S(n15862), .Z(n13330) );
  INV_X1 U16424 ( .A(n13330), .ZN(P1_U3472) );
  INV_X1 U16425 ( .A(P2_LWORD_REG_15__SCAN_IN), .ZN(n13332) );
  AOI22_X1 U16426 ( .A1(n13571), .A2(BUF1_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n13331), .ZN(n18973) );
  INV_X1 U16427 ( .A(P2_EAX_REG_15__SCAN_IN), .ZN(n19042) );
  OAI222_X1 U16428 ( .A1(n13250), .A2(n13332), .B1(n13348), .B2(n18973), .C1(
        n13347), .C2(n19042), .ZN(P2_U2982) );
  NAND2_X1 U16429 ( .A1(n13334), .A2(n13333), .ZN(n13335) );
  NAND2_X1 U16430 ( .A1(n13454), .A2(n13335), .ZN(n13414) );
  INV_X1 U16431 ( .A(P1_EBX_REG_3__SCAN_IN), .ZN(n13340) );
  NOR2_X1 U16432 ( .A1(n13337), .A2(n13338), .ZN(n13339) );
  OR2_X1 U16433 ( .A1(n13336), .A2(n13339), .ZN(n13493) );
  OAI222_X1 U16434 ( .A1(n13414), .A2(n14356), .B1(n13340), .B2(n19945), .C1(
        n13493), .C2(n9630), .ZN(P1_U2869) );
  AOI22_X1 U16435 ( .A1(n9634), .A2(P2_UWORD_REG_12__SCAN_IN), .B1(n19067), 
        .B2(P2_DATAO_REG_28__SCAN_IN), .ZN(n13341) );
  OAI21_X1 U16436 ( .B1(n20839), .B2(n19037), .A(n13341), .ZN(P2_U2923) );
  AOI22_X1 U16437 ( .A1(n9634), .A2(P2_UWORD_REG_13__SCAN_IN), .B1(n19067), 
        .B2(P2_DATAO_REG_29__SCAN_IN), .ZN(n13342) );
  OAI21_X1 U16438 ( .B1(n14642), .B2(n19037), .A(n13342), .ZN(P2_U2922) );
  INV_X1 U16439 ( .A(P2_LWORD_REG_0__SCAN_IN), .ZN(n13344) );
  OAI222_X1 U16440 ( .A1(n13344), .A2(n13250), .B1(n13348), .B2(n13727), .C1(
        n13347), .C2(n13343), .ZN(P2_U2967) );
  INV_X1 U16441 ( .A(P2_UWORD_REG_0__SCAN_IN), .ZN(n13345) );
  OAI222_X1 U16442 ( .A1(n13348), .A2(n13727), .B1(n13347), .B2(n13346), .C1(
        n13250), .C2(n13345), .ZN(P2_U2952) );
  XNOR2_X1 U16443 ( .A(n13350), .B(n13349), .ZN(n13418) );
  NOR2_X1 U16444 ( .A1(n20050), .A2(n20620), .ZN(n13415) );
  NOR2_X1 U16445 ( .A1(n20039), .A2(n19908), .ZN(n13351) );
  AOI211_X1 U16446 ( .C1(n15635), .C2(n19911), .A(n13415), .B(n13351), .ZN(
        n13353) );
  INV_X1 U16447 ( .A(n13493), .ZN(n19913) );
  NAND2_X1 U16448 ( .A1(n19913), .A2(n15645), .ZN(n13352) );
  OAI211_X1 U16449 ( .C1(n13418), .C2(n20031), .A(n13353), .B(n13352), .ZN(
        P1_U2996) );
  XNOR2_X1 U16450 ( .A(n13355), .B(n13354), .ZN(n20052) );
  INV_X1 U16451 ( .A(n14308), .ZN(n13358) );
  AOI22_X1 U16452 ( .A1(n20034), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B1(
        n20043), .B2(P1_REIP_REG_2__SCAN_IN), .ZN(n13356) );
  OAI21_X1 U16453 ( .B1(n20032), .B2(n14303), .A(n13356), .ZN(n13357) );
  AOI21_X1 U16454 ( .B1(n13358), .B2(n15645), .A(n13357), .ZN(n13359) );
  OAI21_X1 U16455 ( .B1(n20031), .B2(n20052), .A(n13359), .ZN(P1_U2997) );
  NOR2_X1 U16456 ( .A1(n13361), .A2(n13362), .ZN(n13363) );
  OR2_X1 U16457 ( .A1(n13360), .A2(n13363), .ZN(n16033) );
  AND2_X1 U16458 ( .A1(n13082), .A2(n13364), .ZN(n14170) );
  INV_X1 U16459 ( .A(n14170), .ZN(n13369) );
  NAND2_X1 U16460 ( .A1(n13082), .A2(n13365), .ZN(n18951) );
  INV_X1 U16461 ( .A(n13366), .ZN(n13376) );
  OAI21_X1 U16462 ( .B1(n18951), .B2(n13376), .A(n13367), .ZN(n13368) );
  NAND3_X1 U16463 ( .A1(n13369), .A2(n15942), .A3(n13368), .ZN(n13371) );
  NAND2_X1 U16464 ( .A1(n15938), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n13370) );
  OAI211_X1 U16465 ( .C1(n16033), .C2(n15938), .A(n13371), .B(n13370), .ZN(
        P2_U2875) );
  NOR2_X1 U16466 ( .A1(n13336), .A2(n13373), .ZN(n13374) );
  OR2_X1 U16467 ( .A1(n13372), .A2(n13374), .ZN(n19892) );
  XOR2_X1 U16468 ( .A(n13451), .B(n13454), .Z(n19893) );
  INV_X1 U16469 ( .A(P1_EBX_REG_4__SCAN_IN), .ZN(n13375) );
  OAI222_X1 U16470 ( .A1(n19892), .A2(n9630), .B1(n14356), .B2(n19893), .C1(
        n19945), .C2(n13375), .ZN(P1_U2868) );
  XNOR2_X1 U16471 ( .A(n18951), .B(n13376), .ZN(n13380) );
  AND2_X1 U16472 ( .A1(n15012), .A2(n13377), .ZN(n13378) );
  OR2_X1 U16473 ( .A1(n13378), .A2(n13361), .ZN(n18846) );
  MUX2_X1 U16474 ( .A(n11541), .B(n18846), .S(n18958), .Z(n13379) );
  OAI21_X1 U16475 ( .B1(n13380), .B2(n18952), .A(n13379), .ZN(P2_U2876) );
  NAND2_X1 U16476 ( .A1(n13383), .A2(n20728), .ZN(n13385) );
  OAI211_X1 U16477 ( .C1(n13185), .C2(n13385), .A(n19946), .B(n13384), .ZN(
        n13386) );
  NAND2_X1 U16478 ( .A1(n10256), .A2(n15405), .ZN(n13388) );
  NAND2_X1 U16479 ( .A1(n13388), .A2(n13387), .ZN(n13390) );
  MUX2_X1 U16480 ( .A(n13391), .B(n13390), .S(n13389), .Z(n13392) );
  INV_X1 U16481 ( .A(n13394), .ZN(n13411) );
  NOR2_X1 U16482 ( .A1(n13396), .A2(n13395), .ZN(n15347) );
  OAI211_X1 U16483 ( .C1(n20107), .C2(n13411), .A(n13397), .B(n15347), .ZN(
        n13398) );
  INV_X1 U16484 ( .A(n13399), .ZN(n15350) );
  AOI21_X1 U16485 ( .B1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n20048) );
  INV_X1 U16486 ( .A(n13400), .ZN(n13403) );
  INV_X1 U16487 ( .A(n13401), .ZN(n13402) );
  OAI211_X1 U16488 ( .C1(n13404), .C2(n14298), .A(n13403), .B(n13402), .ZN(
        n13405) );
  INV_X1 U16489 ( .A(n15328), .ZN(n14182) );
  INV_X1 U16490 ( .A(n15773), .ZN(n20065) );
  INV_X1 U16491 ( .A(n20046), .ZN(n15739) );
  OAI221_X1 U16492 ( .B1(n15819), .B2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .C1(
        n15819), .C2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A(n15739), .ZN(
        n13406) );
  AOI21_X1 U16493 ( .B1(n15798), .B2(n20048), .A(n13406), .ZN(n13407) );
  INV_X1 U16494 ( .A(n13407), .ZN(n13496) );
  NOR2_X1 U16495 ( .A1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n15376), .ZN(
        n20059) );
  NOR2_X1 U16496 ( .A1(n15819), .A2(n20059), .ZN(n15802) );
  NAND2_X1 U16497 ( .A1(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n15802), .ZN(
        n20058) );
  OAI21_X1 U16498 ( .B1(n11122), .B2(n20058), .A(n20066), .ZN(n15811) );
  INV_X1 U16499 ( .A(n15811), .ZN(n13408) );
  NOR2_X1 U16500 ( .A1(n20048), .A2(n13408), .ZN(n13499) );
  AOI22_X1 U16501 ( .A1(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n13496), .B1(
        n13499), .B2(n13409), .ZN(n13417) );
  NAND2_X1 U16502 ( .A1(n11064), .A2(n20096), .ZN(n15360) );
  OAI21_X1 U16503 ( .B1(n13411), .B2(n13410), .A(n15360), .ZN(n13412) );
  INV_X1 U16504 ( .A(n13414), .ZN(n19906) );
  AOI21_X1 U16505 ( .B1(n20064), .B2(n19906), .A(n13415), .ZN(n13416) );
  OAI211_X1 U16506 ( .C1(n20070), .C2(n13418), .A(n13417), .B(n13416), .ZN(
        P1_U3028) );
  NOR2_X1 U16507 ( .A1(P1_FLUSH_REG_SCAN_IN), .A2(n13663), .ZN(n13421) );
  MUX2_X1 U16508 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n13419), .S(
        n15331), .Z(n15339) );
  AOI22_X1 U16509 ( .A1(n13421), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B1(
        n15339), .B2(n13663), .ZN(n13423) );
  MUX2_X1 U16510 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n13420), .S(
        n15331), .Z(n15335) );
  AOI22_X1 U16511 ( .A1(n15335), .A2(n13663), .B1(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B2(n13421), .ZN(n13422) );
  NAND2_X1 U16512 ( .A1(n13663), .A2(n15331), .ZN(n13426) );
  OAI21_X1 U16513 ( .B1(n15861), .B2(P1_FLUSH_REG_SCAN_IN), .A(n13426), .ZN(
        n13429) );
  INV_X1 U16514 ( .A(n20214), .ZN(n20437) );
  OR2_X1 U16515 ( .A1(n13424), .A2(n20437), .ZN(n13425) );
  XNOR2_X1 U16516 ( .A(n13425), .B(n15861), .ZN(n19904) );
  OR2_X1 U16517 ( .A1(n19904), .A2(n11067), .ZN(n15856) );
  INV_X1 U16518 ( .A(n13426), .ZN(n13427) );
  NAND2_X1 U16519 ( .A1(n15856), .A2(n13427), .ZN(n13428) );
  NAND2_X1 U16520 ( .A1(n13429), .A2(n13428), .ZN(n15358) );
  OR2_X1 U16521 ( .A1(n15366), .A2(P1_FLUSH_REG_SCAN_IN), .ZN(n13431) );
  INV_X1 U16522 ( .A(n15870), .ZN(n13430) );
  NAND2_X1 U16523 ( .A1(n13431), .A2(n13430), .ZN(n13432) );
  NAND2_X1 U16524 ( .A1(n13432), .A2(n20131), .ZN(n20702) );
  NAND2_X1 U16525 ( .A1(P1_STATEBS16_REG_SCAN_IN), .A2(n13433), .ZN(n20691) );
  XOR2_X1 U16526 ( .A(n20691), .B(n13434), .Z(n13435) );
  INV_X1 U16527 ( .A(n13312), .ZN(n20324) );
  INV_X1 U16528 ( .A(P1_STATE2_REG_3__SCAN_IN), .ZN(n20440) );
  NAND2_X1 U16529 ( .A1(n20440), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n20698) );
  AOI22_X1 U16530 ( .A1(n13435), .A2(n20700), .B1(n20324), .B2(n20698), .ZN(
        n13437) );
  NAND2_X1 U16531 ( .A1(n20706), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n13436) );
  OAI21_X1 U16532 ( .B1(n20706), .B2(n13437), .A(n13436), .ZN(P1_U3476) );
  XNOR2_X1 U16533 ( .A(n13439), .B(n13438), .ZN(n13450) );
  NAND2_X1 U16534 ( .A1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n13440) );
  OAI211_X1 U16535 ( .C1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .C2(
        P1_INSTADDRPOINTER_REG_3__SCAN_IN), .A(n13499), .B(n13440), .ZN(n13443) );
  NOR2_X1 U16536 ( .A1(n20050), .A2(n20621), .ZN(n13444) );
  NOR2_X1 U16537 ( .A1(n20081), .A2(n19893), .ZN(n13441) );
  AOI211_X1 U16538 ( .C1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .C2(n13496), .A(
        n13444), .B(n13441), .ZN(n13442) );
  OAI211_X1 U16539 ( .C1(n20070), .C2(n13450), .A(n13443), .B(n13442), .ZN(
        P1_U3027) );
  AOI21_X1 U16540 ( .B1(n20034), .B2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n13444), .ZN(n13447) );
  INV_X1 U16541 ( .A(n19896), .ZN(n13445) );
  NAND2_X1 U16542 ( .A1(n15635), .A2(n13445), .ZN(n13446) );
  OAI211_X1 U16543 ( .C1(n19892), .C2(n20084), .A(n13447), .B(n13446), .ZN(
        n13448) );
  INV_X1 U16544 ( .A(n13448), .ZN(n13449) );
  OAI21_X1 U16545 ( .B1(n13450), .B2(n20031), .A(n13449), .ZN(P1_U2995) );
  INV_X1 U16546 ( .A(n15850), .ZN(n13456) );
  INV_X1 U16547 ( .A(n13451), .ZN(n13453) );
  OAI21_X1 U16548 ( .B1(n13454), .B2(n13453), .A(n13452), .ZN(n13455) );
  NAND2_X1 U16549 ( .A1(n13456), .A2(n13455), .ZN(n19882) );
  INV_X1 U16550 ( .A(P1_EBX_REG_5__SCAN_IN), .ZN(n13460) );
  INV_X1 U16551 ( .A(n13457), .ZN(n13750) );
  NOR2_X1 U16552 ( .A1(n13372), .A2(n13458), .ZN(n13459) );
  OR2_X1 U16553 ( .A1(n13750), .A2(n13459), .ZN(n19885) );
  OAI222_X1 U16554 ( .A1(n19882), .A2(n14356), .B1(n13460), .B2(n19945), .C1(
        n19885), .C2(n9630), .ZN(P1_U2867) );
  NAND2_X1 U16555 ( .A1(n9887), .A2(n13503), .ZN(n13461) );
  XNOR2_X1 U16556 ( .A(n13462), .B(n13461), .ZN(n13463) );
  NAND2_X1 U16557 ( .A1(n13463), .A2(n18920), .ZN(n13475) );
  INV_X1 U16558 ( .A(n18928), .ZN(n18874) );
  NAND2_X1 U16559 ( .A1(n13465), .A2(n13464), .ZN(n13468) );
  INV_X1 U16560 ( .A(n13466), .ZN(n13467) );
  NAND2_X1 U16561 ( .A1(n13468), .A2(n13467), .ZN(n19762) );
  INV_X1 U16562 ( .A(n18923), .ZN(n18896) );
  NAND2_X1 U16563 ( .A1(n18896), .A2(n13469), .ZN(n13471) );
  INV_X1 U16564 ( .A(n18929), .ZN(n18842) );
  AOI22_X1 U16565 ( .A1(n18842), .A2(P2_EBX_REG_2__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n18892), .ZN(n13470) );
  OAI211_X1 U16566 ( .C1(n13015), .C2(n18932), .A(n13471), .B(n13470), .ZN(
        n13473) );
  NOR2_X1 U16567 ( .A1(n13011), .A2(n18924), .ZN(n13472) );
  AOI211_X1 U16568 ( .C1(n18874), .C2(n19762), .A(n13473), .B(n13472), .ZN(
        n13474) );
  OAI211_X1 U16569 ( .C1(n13559), .C2(n19760), .A(n13475), .B(n13474), .ZN(
        P2_U2853) );
  AND2_X1 U16570 ( .A1(n18831), .A2(n13476), .ZN(n13478) );
  AOI21_X1 U16571 ( .B1(n19079), .B2(n13478), .A(n18890), .ZN(n13477) );
  OAI21_X1 U16572 ( .B1(n19079), .B2(n13478), .A(n13477), .ZN(n13488) );
  AOI21_X1 U16573 ( .B1(n13481), .B2(n13549), .A(n13480), .ZN(n19095) );
  AOI22_X1 U16574 ( .A1(n18910), .A2(P2_REIP_REG_4__SCAN_IN), .B1(n18874), 
        .B2(n19095), .ZN(n13484) );
  OAI21_X1 U16575 ( .B1(n19094), .B2(n18935), .A(n12482), .ZN(n13482) );
  AOI21_X1 U16576 ( .B1(n18842), .B2(P2_EBX_REG_4__SCAN_IN), .A(n13482), .ZN(
        n13483) );
  OAI211_X1 U16577 ( .C1(n13485), .C2(n18923), .A(n13484), .B(n13483), .ZN(
        n13486) );
  AOI21_X1 U16578 ( .B1(n19096), .B2(n18916), .A(n13486), .ZN(n13487) );
  OAI211_X1 U16579 ( .C1(n13559), .C2(n19008), .A(n13488), .B(n13487), .ZN(
        P2_U2851) );
  NAND2_X1 U16580 ( .A1(n13490), .A2(n13489), .ZN(n13491) );
  NAND2_X2 U16581 ( .A1(n14436), .A2(n13491), .ZN(n14396) );
  INV_X1 U16582 ( .A(n13491), .ZN(n13492) );
  INV_X1 U16583 ( .A(n14429), .ZN(n20097) );
  OAI222_X1 U16584 ( .A1(n20036), .A2(n14396), .B1(n14144), .B2(n20097), .C1(
        n14436), .C2(n10374), .ZN(P1_U2903) );
  INV_X1 U16585 ( .A(n14418), .ZN(n20104) );
  OAI222_X1 U16586 ( .A1(n13493), .A2(n14396), .B1(n14144), .B2(n20104), .C1(
        n14436), .C2(n10407), .ZN(P1_U2901) );
  INV_X1 U16587 ( .A(n14407), .ZN(n20111) );
  INV_X1 U16588 ( .A(P1_EAX_REG_5__SCAN_IN), .ZN(n19989) );
  OAI222_X1 U16589 ( .A1(n19885), .A2(n14396), .B1(n14144), .B2(n20111), .C1(
        n14436), .C2(n19989), .ZN(P1_U2899) );
  INV_X1 U16590 ( .A(n14423), .ZN(n20100) );
  OAI222_X1 U16591 ( .A1(n14308), .A2(n14396), .B1(n14144), .B2(n20100), .C1(
        n14436), .C2(n10355), .ZN(P1_U2902) );
  XNOR2_X1 U16592 ( .A(n13495), .B(n13494), .ZN(n15660) );
  INV_X1 U16593 ( .A(n15819), .ZN(n20047) );
  NAND3_X1 U16594 ( .A1(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_4__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n14550) );
  AOI21_X1 U16595 ( .B1(n15834), .B2(n14550), .A(n13496), .ZN(n13497) );
  INV_X1 U16596 ( .A(n13497), .ZN(n15851) );
  NAND4_X1 U16597 ( .A1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_3__SCAN_IN), .A3(n13499), .A4(n13498), .ZN(
        n13500) );
  NAND2_X1 U16598 ( .A1(n20043), .A2(P1_REIP_REG_5__SCAN_IN), .ZN(n15662) );
  OAI211_X1 U16599 ( .C1(n20081), .C2(n19882), .A(n13500), .B(n15662), .ZN(
        n13501) );
  AOI21_X1 U16600 ( .B1(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n15851), .A(
        n13501), .ZN(n13502) );
  OAI21_X1 U16601 ( .B1(n20070), .B2(n15660), .A(n13502), .ZN(P1_U3026) );
  NAND2_X1 U16602 ( .A1(n18920), .A2(n18912), .ZN(n18855) );
  OAI211_X1 U16603 ( .C1(n18939), .C2(n13504), .A(n9887), .B(n13503), .ZN(
        n13763) );
  OAI22_X1 U16604 ( .A1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n18855), .B1(
        n13763), .B2(n18890), .ZN(n13505) );
  INV_X1 U16605 ( .A(n13505), .ZN(n13515) );
  OR2_X1 U16606 ( .A1(n13507), .A2(n13506), .ZN(n13509) );
  NAND2_X1 U16607 ( .A1(n13509), .A2(n13508), .ZN(n19771) );
  AOI22_X1 U16608 ( .A1(n18910), .A2(P2_REIP_REG_1__SCAN_IN), .B1(n18874), 
        .B2(n19771), .ZN(n13511) );
  AOI22_X1 U16609 ( .A1(n18842), .A2(P2_EBX_REG_1__SCAN_IN), .B1(n18892), .B2(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n13510) );
  OAI211_X1 U16610 ( .C1(n18923), .C2(n13512), .A(n13511), .B(n13510), .ZN(
        n13513) );
  AOI21_X1 U16611 ( .B1(n18916), .B2(n19130), .A(n13513), .ZN(n13514) );
  OAI211_X1 U16612 ( .C1(n13559), .C2(n18999), .A(n13515), .B(n13514), .ZN(
        P2_U2854) );
  AOI21_X1 U16613 ( .B1(n14170), .B2(n14169), .A(n13517), .ZN(n13518) );
  OR3_X1 U16614 ( .A1(n13516), .A2(n13518), .A3(n18952), .ZN(n13522) );
  AOI21_X1 U16615 ( .B1(n13520), .B2(n14172), .A(n13519), .ZN(n18814) );
  NAND2_X1 U16616 ( .A1(n15948), .A2(n18814), .ZN(n13521) );
  OAI211_X1 U16617 ( .C1(n15948), .C2(n18808), .A(n13522), .B(n13521), .ZN(
        P2_U2873) );
  NAND2_X1 U16618 ( .A1(n13525), .A2(n13524), .ZN(n13527) );
  XNOR2_X1 U16619 ( .A(n13527), .B(n13526), .ZN(n16133) );
  NAND2_X1 U16620 ( .A1(n16133), .A2(n16066), .ZN(n13531) );
  NAND2_X1 U16621 ( .A1(n19081), .A2(P2_REIP_REG_3__SCAN_IN), .ZN(n16127) );
  OAI21_X1 U16622 ( .B1(n19093), .B2(n11504), .A(n16127), .ZN(n13529) );
  NOR2_X1 U16623 ( .A1(n16063), .A2(n13544), .ZN(n13528) );
  AOI211_X1 U16624 ( .C1(n9650), .C2(n19090), .A(n13529), .B(n13528), .ZN(
        n13530) );
  OAI211_X1 U16625 ( .C1(n16131), .C2(n19087), .A(n13531), .B(n13530), .ZN(
        P2_U3011) );
  XOR2_X1 U16626 ( .A(n9701), .B(n13532), .Z(n15026) );
  INV_X1 U16627 ( .A(n15026), .ZN(n18989) );
  NOR2_X1 U16628 ( .A1(n18912), .A2(n13533), .ZN(n13534) );
  XNOR2_X1 U16629 ( .A(n13534), .B(n16055), .ZN(n13535) );
  NAND2_X1 U16630 ( .A1(n13535), .A2(n18920), .ZN(n13542) );
  AOI21_X1 U16631 ( .B1(n18892), .B2(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .A(
        n19081), .ZN(n13536) );
  OAI21_X1 U16632 ( .B1(n18929), .B2(n11429), .A(n13536), .ZN(n13537) );
  AOI21_X1 U16633 ( .B1(n18910), .B2(P2_REIP_REG_9__SCAN_IN), .A(n13537), .ZN(
        n13538) );
  OAI21_X1 U16634 ( .B1(n18924), .B2(n16062), .A(n13538), .ZN(n13539) );
  AOI21_X1 U16635 ( .B1(n13540), .B2(n18896), .A(n13539), .ZN(n13541) );
  OAI211_X1 U16636 ( .C1(n18989), .C2(n18928), .A(n13542), .B(n13541), .ZN(
        P2_U2846) );
  NOR2_X1 U16637 ( .A1(n18912), .A2(n13543), .ZN(n13545) );
  XNOR2_X1 U16638 ( .A(n13545), .B(n13544), .ZN(n13546) );
  NAND2_X1 U16639 ( .A1(n13546), .A2(n18920), .ZN(n13558) );
  OR2_X1 U16640 ( .A1(n13548), .A2(n13547), .ZN(n13550) );
  NAND2_X1 U16641 ( .A1(n13550), .A2(n13549), .ZN(n19012) );
  OAI22_X1 U16642 ( .A1(n11505), .A2(n18932), .B1(n18928), .B2(n19012), .ZN(
        n13553) );
  OAI22_X1 U16643 ( .A1(n18929), .A2(n13551), .B1(n11504), .B2(n18935), .ZN(
        n13552) );
  NOR2_X1 U16644 ( .A1(n13553), .A2(n13552), .ZN(n13554) );
  OAI21_X1 U16645 ( .B1(n13555), .B2(n18923), .A(n13554), .ZN(n13556) );
  AOI21_X1 U16646 ( .B1(n9650), .B2(n18916), .A(n13556), .ZN(n13557) );
  OAI211_X1 U16647 ( .C1(n13559), .C2(n19000), .A(n13558), .B(n13557), .ZN(
        P2_U2852) );
  NAND2_X1 U16648 ( .A1(n19000), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19338) );
  OR2_X1 U16649 ( .A1(n19338), .A2(n19459), .ZN(n13560) );
  NAND2_X1 U16650 ( .A1(n19757), .A2(n19764), .ZN(n19217) );
  OR2_X1 U16651 ( .A1(n19773), .A2(n19217), .ZN(n19215) );
  NAND2_X1 U16652 ( .A1(n13567), .A2(n19215), .ZN(n13566) );
  INV_X1 U16653 ( .A(n19752), .ZN(n19747) );
  NOR2_X1 U16654 ( .A1(n19455), .A2(n19217), .ZN(n19262) );
  INV_X1 U16655 ( .A(n19262), .ZN(n13561) );
  OAI211_X1 U16656 ( .C1(n12122), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19747), 
        .B(n13561), .ZN(n13564) );
  INV_X1 U16657 ( .A(P2_STATE2_REG_2__SCAN_IN), .ZN(n19801) );
  AOI21_X1 U16658 ( .B1(n19801), .B2(n13649), .A(P2_STATE2_REG_0__SCAN_IN), 
        .ZN(n19799) );
  NAND2_X1 U16659 ( .A1(n19799), .A2(n19776), .ZN(n13562) );
  AND2_X1 U16660 ( .A1(n13564), .A2(n19593), .ZN(n13565) );
  NAND2_X1 U16661 ( .A1(n13566), .A2(n13565), .ZN(n19265) );
  INV_X1 U16662 ( .A(n19265), .ZN(n19250) );
  INV_X1 U16663 ( .A(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n13578) );
  NOR2_X2 U16664 ( .A1(n19025), .A2(n19528), .ZN(n19614) );
  INV_X1 U16665 ( .A(n13567), .ZN(n13570) );
  INV_X1 U16666 ( .A(n12122), .ZN(n13568) );
  OAI21_X1 U16667 ( .B1(n13568), .B2(n19262), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n13569) );
  OAI21_X1 U16668 ( .B1(n13570), .B2(n19215), .A(n13569), .ZN(n19264) );
  NAND2_X1 U16669 ( .A1(n19000), .A2(n19779), .ZN(n19307) );
  INV_X1 U16670 ( .A(BUF2_REG_26__SCAN_IN), .ZN(n18060) );
  INV_X1 U16671 ( .A(BUF1_REG_26__SCAN_IN), .ZN(n16257) );
  OAI22_X2 U16672 ( .A1(n18060), .A2(n19163), .B1(n16257), .B2(n19165), .ZN(
        n19616) );
  INV_X1 U16673 ( .A(n19616), .ZN(n19506) );
  AOI22_X1 U16674 ( .A1(BUF1_REG_18__SCAN_IN), .A2(n19179), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n19180), .ZN(n19471) );
  INV_X1 U16675 ( .A(n19471), .ZN(n19615) );
  INV_X1 U16676 ( .A(n19176), .ZN(n13573) );
  AND2_X1 U16677 ( .A1(n13574), .A2(n13573), .ZN(n19613) );
  AOI22_X1 U16678 ( .A1(n19276), .A2(n19615), .B1(n19613), .B2(n19262), .ZN(
        n13575) );
  OAI21_X1 U16679 ( .B1(n19261), .B2(n19506), .A(n13575), .ZN(n13576) );
  AOI21_X1 U16680 ( .B1(n19614), .B2(n19264), .A(n13576), .ZN(n13577) );
  OAI21_X1 U16681 ( .B1(n19250), .B2(n13578), .A(n13577), .ZN(P2_U3074) );
  NOR2_X1 U16682 ( .A1(n13581), .A2(n13580), .ZN(n13582) );
  OR2_X1 U16683 ( .A1(n13579), .A2(n13582), .ZN(n19862) );
  INV_X1 U16684 ( .A(n14399), .ZN(n20123) );
  OAI222_X1 U16685 ( .A1(n19862), .A2(n14396), .B1(n14144), .B2(n20123), .C1(
        n14436), .C2(n10480), .ZN(P1_U2897) );
  INV_X1 U16686 ( .A(n15849), .ZN(n13585) );
  INV_X1 U16687 ( .A(n13583), .ZN(n13584) );
  AOI21_X1 U16688 ( .B1(n15850), .B2(n13585), .A(n13584), .ZN(n13586) );
  OR2_X1 U16689 ( .A1(n13659), .A2(n13586), .ZN(n19856) );
  INV_X1 U16690 ( .A(P1_EBX_REG_7__SCAN_IN), .ZN(n19855) );
  OAI222_X1 U16691 ( .A1(n19856), .A2(n14356), .B1(n19855), .B2(n19945), .C1(
        n19862), .C2(n9630), .ZN(P1_U2865) );
  INV_X1 U16692 ( .A(n11629), .ZN(n13651) );
  NAND2_X1 U16693 ( .A1(n13587), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n19809) );
  NOR2_X1 U16694 ( .A1(n13589), .A2(n13588), .ZN(n13614) );
  AND2_X1 U16695 ( .A1(n13614), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13592) );
  NAND2_X1 U16696 ( .A1(n13606), .A2(n13595), .ZN(n13613) );
  INV_X1 U16697 ( .A(n11658), .ZN(n13590) );
  NAND2_X1 U16698 ( .A1(n13590), .A2(n13620), .ZN(n13611) );
  OAI211_X1 U16699 ( .C1(n13592), .C2(n13591), .A(n13613), .B(n13611), .ZN(
        n13597) );
  INV_X1 U16700 ( .A(n13606), .ZN(n13601) );
  NAND2_X1 U16701 ( .A1(n13633), .A2(n13630), .ZN(n13617) );
  OAI21_X1 U16702 ( .B1(n13617), .B2(n13593), .A(n13611), .ZN(n13594) );
  OAI211_X1 U16703 ( .C1(n13601), .C2(n13595), .A(n13594), .B(n11278), .ZN(
        n13596) );
  AOI22_X1 U16704 ( .A1(n9650), .A2(n13598), .B1(n13597), .B2(n13596), .ZN(
        n15043) );
  INV_X1 U16705 ( .A(n13622), .ZN(n13642) );
  MUX2_X1 U16706 ( .A(n11347), .B(n15043), .S(n13642), .Z(n13645) );
  INV_X1 U16707 ( .A(n13598), .ZN(n13619) );
  NAND2_X1 U16708 ( .A1(n13600), .A2(n13599), .ZN(n13605) );
  INV_X1 U16709 ( .A(n13605), .ZN(n13602) );
  MUX2_X1 U16710 ( .A(n13602), .B(n13601), .S(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .Z(n13603) );
  OAI21_X1 U16711 ( .B1(n18925), .B2(n13619), .A(n13603), .ZN(n15036) );
  NOR2_X1 U16712 ( .A1(n11657), .A2(n11658), .ZN(n13604) );
  AOI22_X1 U16713 ( .A1(n13606), .A2(n11612), .B1(n13605), .B2(n13604), .ZN(
        n13607) );
  OAI21_X1 U16714 ( .B1(n13608), .B2(n13619), .A(n13607), .ZN(n13778) );
  OAI21_X1 U16715 ( .B1(n15036), .B2(n19455), .A(n13778), .ZN(n13610) );
  OAI21_X1 U16716 ( .B1(n15036), .B2(n19783), .A(n19773), .ZN(n13609) );
  AOI21_X1 U16717 ( .B1(n13610), .B2(n13609), .A(n13622), .ZN(n13625) );
  NAND2_X1 U16718 ( .A1(n11643), .A2(n13611), .ZN(n13616) );
  OAI22_X1 U16719 ( .A1(n13614), .A2(n13616), .B1(n13612), .B2(n13613), .ZN(
        n13615) );
  AOI21_X1 U16720 ( .B1(n13617), .B2(n13616), .A(n13615), .ZN(n13618) );
  OAI21_X1 U16721 ( .B1(n13011), .B2(n13619), .A(n13618), .ZN(n13764) );
  NAND2_X1 U16722 ( .A1(n13622), .A2(n13620), .ZN(n13621) );
  OAI21_X1 U16723 ( .B1(n13764), .B2(n13622), .A(n13621), .ZN(n13644) );
  NOR2_X1 U16724 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n13644), .ZN(
        n13624) );
  AOI21_X1 U16725 ( .B1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n13645), .A(
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n13623) );
  AOI222_X1 U16726 ( .A1(n13625), .A2(n13624), .B1(n13625), .B2(n13623), .C1(
        n13624), .C2(n19764), .ZN(n13626) );
  OAI21_X1 U16727 ( .B1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n13645), .A(
        n13626), .ZN(n13648) );
  INV_X1 U16728 ( .A(n13627), .ZN(n13629) );
  OAI211_X1 U16729 ( .C1(P2_MORE_REG_SCAN_IN), .C2(P2_FLUSH_REG_SCAN_IN), .A(
        n13629), .B(n13628), .ZN(n13640) );
  INV_X1 U16730 ( .A(n13630), .ZN(n13636) );
  INV_X1 U16731 ( .A(n13631), .ZN(n13632) );
  OAI22_X1 U16732 ( .A1(n13635), .A2(n13633), .B1(n13641), .B2(n13632), .ZN(
        n13634) );
  AOI21_X1 U16733 ( .B1(n13636), .B2(n13635), .A(n13634), .ZN(n19790) );
  INV_X1 U16734 ( .A(n12367), .ZN(n13638) );
  AOI21_X1 U16735 ( .B1(n13638), .B2(n11389), .A(n13637), .ZN(n13639) );
  OAI211_X1 U16736 ( .C1(n13641), .C2(n13640), .A(n19790), .B(n13639), .ZN(
        n13647) );
  OAI22_X1 U16737 ( .A1(n13645), .A2(n13644), .B1(n13643), .B2(n13642), .ZN(
        n13646) );
  AOI211_X1 U16738 ( .C1(n15428), .C2(n13648), .A(n13647), .B(n13646), .ZN(
        n16153) );
  AOI21_X1 U16739 ( .B1(n16153), .B2(n13649), .A(n18715), .ZN(n13650) );
  AOI211_X1 U16740 ( .C1(n13652), .C2(n13651), .A(n19809), .B(n13650), .ZN(
        n19657) );
  OAI21_X1 U16741 ( .B1(n19657), .B2(n18715), .A(P2_STATE2_REG_3__SCAN_IN), 
        .ZN(n13654) );
  INV_X1 U16742 ( .A(n16147), .ZN(n13653) );
  NAND2_X1 U16743 ( .A1(n13654), .A2(n13653), .ZN(P2_U3593) );
  OAI21_X1 U16744 ( .B1(n13579), .B2(n13656), .A(n13655), .ZN(n13756) );
  NOR2_X1 U16745 ( .A1(n14228), .A2(n13657), .ZN(n14126) );
  NOR2_X1 U16746 ( .A1(n15471), .A2(n14126), .ZN(n13669) );
  OAI21_X1 U16747 ( .B1(n13659), .B2(n13658), .A(n13771), .ZN(n15837) );
  AND2_X1 U16748 ( .A1(n20700), .A2(n13663), .ZN(n13660) );
  NAND2_X1 U16749 ( .A1(n19922), .A2(n13660), .ZN(n19879) );
  NOR2_X1 U16750 ( .A1(n19875), .A2(P1_REIP_REG_8__SCAN_IN), .ZN(n13661) );
  AOI22_X1 U16751 ( .A1(n19929), .A2(P1_EBX_REG_8__SCAN_IN), .B1(n13661), .B2(
        n15537), .ZN(n13662) );
  OAI211_X1 U16752 ( .C1(n19931), .C2(n15837), .A(n19879), .B(n13662), .ZN(
        n13668) );
  NOR2_X1 U16753 ( .A1(n13664), .A2(n13663), .ZN(n13665) );
  INV_X1 U16754 ( .A(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n13666) );
  OAI22_X1 U16755 ( .A1(n13758), .A2(n19897), .B1(n19923), .B2(n13666), .ZN(
        n13667) );
  AOI211_X1 U16756 ( .C1(n13669), .C2(P1_REIP_REG_8__SCAN_IN), .A(n13668), .B(
        n13667), .ZN(n13670) );
  OAI21_X1 U16757 ( .B1(n13756), .B2(n19861), .A(n13670), .ZN(P1_U2832) );
  INV_X1 U16758 ( .A(n15837), .ZN(n13671) );
  AOI22_X1 U16759 ( .A1(n19940), .A2(n13671), .B1(n10965), .B2(
        P1_EBX_REG_8__SCAN_IN), .ZN(n13672) );
  OAI21_X1 U16760 ( .B1(n13756), .B2(n9630), .A(n13672), .ZN(P1_U2864) );
  XNOR2_X1 U16761 ( .A(n13674), .B(n13673), .ZN(n13695) );
  OAI21_X1 U16762 ( .B1(n13480), .B2(n13676), .A(n13675), .ZN(n19005) );
  OAI211_X1 U16763 ( .C1(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .A(n19102), .B(n13677), .ZN(n13680) );
  INV_X1 U16764 ( .A(P2_REIP_REG_5__SCAN_IN), .ZN(n13678) );
  NOR2_X1 U16765 ( .A1(n12482), .A2(n13678), .ZN(n13691) );
  AOI21_X1 U16766 ( .B1(n19131), .B2(n18915), .A(n13691), .ZN(n13679) );
  OAI211_X1 U16767 ( .C1(n19005), .C2(n16128), .A(n13680), .B(n13679), .ZN(
        n13681) );
  AOI21_X1 U16768 ( .B1(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n19100), .A(
        n13681), .ZN(n13689) );
  INV_X1 U16769 ( .A(n13682), .ZN(n13687) );
  AOI21_X1 U16770 ( .B1(n13686), .B2(n13684), .A(n13683), .ZN(n13685) );
  AOI21_X1 U16771 ( .B1(n13687), .B2(n13686), .A(n13685), .ZN(n13692) );
  NAND2_X1 U16772 ( .A1(n13692), .A2(n16122), .ZN(n13688) );
  OAI211_X1 U16773 ( .C1(n13695), .C2(n19110), .A(n13689), .B(n13688), .ZN(
        P2_U3041) );
  INV_X1 U16774 ( .A(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n18906) );
  OAI22_X1 U16775 ( .A1(n18906), .A2(n19093), .B1(n16063), .B2(n18913), .ZN(
        n13690) );
  AOI211_X1 U16776 ( .C1(n19090), .C2(n18915), .A(n13691), .B(n13690), .ZN(
        n13694) );
  NAND2_X1 U16777 ( .A1(n13692), .A2(n16068), .ZN(n13693) );
  OAI211_X1 U16778 ( .C1(n13695), .C2(n19088), .A(n13694), .B(n13693), .ZN(
        P2_U3009) );
  NOR2_X1 U16779 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n19764), .ZN(
        n19333) );
  NAND2_X1 U16780 ( .A1(n19333), .A2(n19773), .ZN(n13702) );
  NOR2_X1 U16781 ( .A1(n19783), .A2(n13702), .ZN(n19298) );
  AOI21_X1 U16782 ( .B1(n12121), .B2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n13698) );
  INV_X1 U16783 ( .A(n19338), .ZN(n13696) );
  INV_X1 U16784 ( .A(n19533), .ZN(n19526) );
  AOI21_X1 U16785 ( .B1(n13696), .B2(n19526), .A(n19747), .ZN(n13699) );
  NAND2_X1 U16786 ( .A1(n13699), .A2(n13702), .ZN(n13697) );
  OAI211_X1 U16787 ( .C1(n19298), .C2(n13698), .A(n13697), .B(n19593), .ZN(
        n19301) );
  INV_X1 U16788 ( .A(n19301), .ZN(n13733) );
  INV_X1 U16789 ( .A(n13699), .ZN(n13703) );
  INV_X1 U16790 ( .A(n12121), .ZN(n13700) );
  OAI21_X1 U16791 ( .B1(n13700), .B2(n19298), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n13701) );
  OAI21_X1 U16792 ( .B1(n13703), .B2(n13702), .A(n13701), .ZN(n19300) );
  AOI22_X1 U16793 ( .A1(n19324), .A2(n19615), .B1(n19298), .B2(n19613), .ZN(
        n13704) );
  OAI21_X1 U16794 ( .B1(n19293), .B2(n19506), .A(n13704), .ZN(n13705) );
  AOI21_X1 U16795 ( .B1(n19614), .B2(n19300), .A(n13705), .ZN(n13706) );
  OAI21_X1 U16796 ( .B1(n13733), .B2(n13707), .A(n13706), .ZN(P2_U3090) );
  XNOR2_X1 U16797 ( .A(n13708), .B(n13736), .ZN(n18777) );
  INV_X1 U16798 ( .A(n19027), .ZN(n13748) );
  AND2_X1 U16799 ( .A1(n13709), .A2(n13710), .ZN(n13712) );
  OR2_X1 U16800 ( .A1(n13712), .A2(n13711), .ZN(n14046) );
  OAI22_X1 U16801 ( .A1(n14691), .A2(n19150), .B1(n13713), .B2(n18995), .ZN(
        n13714) );
  AOI21_X1 U16802 ( .B1(n18965), .B2(BUF2_REG_17__SCAN_IN), .A(n13714), .ZN(
        n13716) );
  NAND2_X1 U16803 ( .A1(n18964), .A2(BUF1_REG_17__SCAN_IN), .ZN(n13715) );
  OAI211_X1 U16804 ( .C1(n14046), .C2(n19002), .A(n13716), .B(n13715), .ZN(
        n13717) );
  INV_X1 U16805 ( .A(n13717), .ZN(n13718) );
  OAI21_X1 U16806 ( .B1(n18777), .B2(n13748), .A(n13718), .ZN(P2_U2902) );
  XNOR2_X1 U16807 ( .A(n13516), .B(n13719), .ZN(n13724) );
  NOR2_X1 U16808 ( .A1(n13720), .A2(n13519), .ZN(n13721) );
  NOR2_X1 U16809 ( .A1(n15289), .A2(n13721), .ZN(n18802) );
  NOR2_X1 U16810 ( .A1(n18958), .A2(n11421), .ZN(n13722) );
  AOI21_X1 U16811 ( .B1(n18802), .B2(n18958), .A(n13722), .ZN(n13723) );
  OAI21_X1 U16812 ( .B1(n13724), .B2(n18952), .A(n13723), .ZN(P2_U2872) );
  MUX2_X1 U16813 ( .A(DATAI_8_), .B(BUF1_REG_8__SCAN_IN), .S(n20085), .Z(
        n19997) );
  INV_X1 U16814 ( .A(n19997), .ZN(n13725) );
  OAI222_X1 U16815 ( .A1(n13756), .A2(n14396), .B1(n14436), .B2(n13726), .C1(
        n14144), .C2(n13725), .ZN(P1_U2896) );
  NOR2_X2 U16816 ( .A1(n13727), .A2(n19528), .ZN(n19601) );
  INV_X1 U16817 ( .A(BUF1_REG_16__SCAN_IN), .ZN(n20909) );
  INV_X1 U16818 ( .A(BUF2_REG_16__SCAN_IN), .ZN(n18052) );
  OAI22_X2 U16819 ( .A1(n20909), .A2(n19165), .B1(n18052), .B2(n19163), .ZN(
        n19603) );
  INV_X1 U16820 ( .A(n19603), .ZN(n19466) );
  AOI22_X1 U16821 ( .A1(BUF1_REG_24__SCAN_IN), .A2(n19179), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n19180), .ZN(n19500) );
  INV_X1 U16822 ( .A(n19500), .ZN(n19602) );
  NOR2_X2 U16823 ( .A1(n13728), .A2(n19176), .ZN(n19600) );
  AOI22_X1 U16824 ( .A1(n19602), .A2(n19299), .B1(n19600), .B2(n19298), .ZN(
        n13729) );
  OAI21_X1 U16825 ( .B1(n19332), .B2(n19466), .A(n13729), .ZN(n13730) );
  AOI21_X1 U16826 ( .B1(n19601), .B2(n19300), .A(n13730), .ZN(n13731) );
  OAI21_X1 U16827 ( .B1(n13733), .B2(n13732), .A(n13731), .ZN(P2_U3088) );
  INV_X1 U16828 ( .A(n13734), .ZN(n13738) );
  OAI21_X1 U16829 ( .B1(n13708), .B2(n13736), .A(n13735), .ZN(n13737) );
  NAND2_X1 U16830 ( .A1(n13738), .A2(n13737), .ZN(n18770) );
  NOR2_X1 U16831 ( .A1(n13711), .A2(n13740), .ZN(n13741) );
  OR2_X1 U16832 ( .A1(n13739), .A2(n13741), .ZN(n15945) );
  OAI22_X1 U16833 ( .A1(n14691), .A2(n19025), .B1(n13742), .B2(n18995), .ZN(
        n13743) );
  AOI21_X1 U16834 ( .B1(n18965), .B2(BUF2_REG_18__SCAN_IN), .A(n13743), .ZN(
        n13745) );
  NAND2_X1 U16835 ( .A1(n18964), .A2(BUF1_REG_18__SCAN_IN), .ZN(n13744) );
  OAI211_X1 U16836 ( .C1(n15945), .C2(n19002), .A(n13745), .B(n13744), .ZN(
        n13746) );
  INV_X1 U16837 ( .A(n13746), .ZN(n13747) );
  OAI21_X1 U16838 ( .B1(n18770), .B2(n13748), .A(n13747), .ZN(P2_U2901) );
  INV_X1 U16839 ( .A(P1_EAX_REG_4__SCAN_IN), .ZN(n19991) );
  INV_X1 U16840 ( .A(n14412), .ZN(n20108) );
  OAI222_X1 U16841 ( .A1(n14396), .A2(n19892), .B1(n14436), .B2(n19991), .C1(
        n14144), .C2(n20108), .ZN(P1_U2900) );
  INV_X1 U16842 ( .A(n14440), .ZN(n20089) );
  OAI222_X1 U16843 ( .A1(n14396), .A2(n20045), .B1(n14144), .B2(n20089), .C1(
        n14436), .C2(n10366), .ZN(P1_U2904) );
  INV_X1 U16844 ( .A(n14403), .ZN(n20114) );
  XOR2_X1 U16845 ( .A(n13750), .B(n13749), .Z(n19942) );
  INV_X1 U16846 ( .A(n19942), .ZN(n13752) );
  OAI222_X1 U16847 ( .A1(n14144), .A2(n20114), .B1(n14396), .B2(n13752), .C1(
        n13751), .C2(n14436), .ZN(P1_U2898) );
  XNOR2_X1 U16848 ( .A(n13753), .B(n15841), .ZN(n13754) );
  XNOR2_X1 U16849 ( .A(n13755), .B(n13754), .ZN(n15836) );
  INV_X1 U16850 ( .A(n13756), .ZN(n13760) );
  AOI22_X1 U16851 ( .A1(n20034), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .B1(
        n20043), .B2(P1_REIP_REG_8__SCAN_IN), .ZN(n13757) );
  OAI21_X1 U16852 ( .B1(n20032), .B2(n13758), .A(n13757), .ZN(n13759) );
  AOI21_X1 U16853 ( .B1(n13760), .B2(n15645), .A(n13759), .ZN(n13761) );
  OAI21_X1 U16854 ( .B1(n20031), .B2(n15836), .A(n13761), .ZN(P1_U2991) );
  AOI221_X1 U16855 ( .B1(n18939), .B2(n9887), .C1(n13762), .C2(n18912), .A(
        n13649), .ZN(n15040) );
  OAI21_X1 U16856 ( .B1(n9887), .B2(n11463), .A(n13763), .ZN(n13776) );
  AOI222_X1 U16857 ( .A1(n13764), .A2(n15042), .B1(n15040), .B2(n13776), .C1(
        n15037), .C2(n19138), .ZN(n13766) );
  NAND2_X1 U16858 ( .A1(n15044), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13765) );
  OAI21_X1 U16859 ( .B1(n13766), .B2(n15044), .A(n13765), .ZN(P2_U3599) );
  INV_X1 U16860 ( .A(n13767), .ZN(n13768) );
  AOI21_X1 U16861 ( .B1(n13769), .B2(n13655), .A(n13768), .ZN(n19843) );
  INV_X1 U16862 ( .A(n19843), .ZN(n13775) );
  INV_X1 U16863 ( .A(n13785), .ZN(n13770) );
  AOI21_X1 U16864 ( .B1(n13772), .B2(n13771), .A(n13770), .ZN(n19841) );
  AOI22_X1 U16865 ( .A1(n19940), .A2(n19841), .B1(n10965), .B2(
        P1_EBX_REG_9__SCAN_IN), .ZN(n13773) );
  OAI21_X1 U16866 ( .B1(n13775), .B2(n9630), .A(n13773), .ZN(P1_U2863) );
  INV_X1 U16867 ( .A(n14144), .ZN(n14095) );
  MUX2_X1 U16868 ( .A(DATAI_9_), .B(BUF1_REG_9__SCAN_IN), .S(n20085), .Z(
        n20001) );
  AOI22_X1 U16869 ( .A1(n14095), .A2(n20001), .B1(P1_EAX_REG_9__SCAN_IN), .B2(
        n14421), .ZN(n13774) );
  OAI21_X1 U16870 ( .B1(n13775), .B2(n14396), .A(n13774), .ZN(P1_U2895) );
  INV_X1 U16871 ( .A(n13776), .ZN(n13777) );
  AOI222_X1 U16872 ( .A1(n13778), .A2(n15042), .B1(n15037), .B2(n19767), .C1(
        n13777), .C2(n15040), .ZN(n13780) );
  NAND2_X1 U16873 ( .A1(n15044), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n13779) );
  OAI21_X1 U16874 ( .B1(n13780), .B2(n15044), .A(n13779), .ZN(P2_U3600) );
  AOI21_X1 U16875 ( .B1(n13783), .B2(n13767), .A(n9605), .ZN(n14546) );
  INV_X1 U16876 ( .A(n14546), .ZN(n13798) );
  AND2_X1 U16877 ( .A1(n13785), .A2(n13784), .ZN(n13786) );
  OR2_X1 U16878 ( .A1(n13786), .A2(n15544), .ZN(n15822) );
  INV_X1 U16879 ( .A(n15822), .ZN(n13789) );
  AOI22_X1 U16880 ( .A1(n19940), .A2(n13789), .B1(n10965), .B2(
        P1_EBX_REG_10__SCAN_IN), .ZN(n13787) );
  OAI21_X1 U16881 ( .B1(n13798), .B2(n9630), .A(n13787), .ZN(P1_U2862) );
  NAND2_X1 U16882 ( .A1(P1_REIP_REG_10__SCAN_IN), .A2(P1_REIP_REG_9__SCAN_IN), 
        .ZN(n15538) );
  INV_X1 U16883 ( .A(n15538), .ZN(n13788) );
  AOI21_X1 U16884 ( .B1(n13788), .B2(n14126), .A(n15471), .ZN(n15551) );
  INV_X1 U16885 ( .A(P1_REIP_REG_10__SCAN_IN), .ZN(n20633) );
  OAI21_X1 U16886 ( .B1(n15471), .B2(n14126), .A(P1_REIP_REG_9__SCAN_IN), .ZN(
        n19845) );
  NAND2_X1 U16887 ( .A1(n20633), .A2(n19845), .ZN(n13795) );
  NAND2_X1 U16888 ( .A1(n13789), .A2(n19905), .ZN(n13790) );
  OAI211_X1 U16889 ( .C1(n13791), .C2(n19867), .A(n19879), .B(n13790), .ZN(
        n13794) );
  INV_X1 U16890 ( .A(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n13792) );
  OAI22_X1 U16891 ( .A1(n14544), .A2(n19897), .B1(n19923), .B2(n13792), .ZN(
        n13793) );
  AOI211_X1 U16892 ( .C1(n15551), .C2(n13795), .A(n13794), .B(n13793), .ZN(
        n13796) );
  OAI21_X1 U16893 ( .B1(n13798), .B2(n19861), .A(n13796), .ZN(P1_U2830) );
  MUX2_X1 U16894 ( .A(DATAI_10_), .B(BUF1_REG_10__SCAN_IN), .S(n20085), .Z(
        n20003) );
  AOI22_X1 U16895 ( .A1(n14095), .A2(n20003), .B1(P1_EAX_REG_10__SCAN_IN), 
        .B2(n14421), .ZN(n13797) );
  OAI21_X1 U16896 ( .B1(n13798), .B2(n14396), .A(n13797), .ZN(P1_U2894) );
  INV_X1 U16897 ( .A(n19333), .ZN(n13799) );
  NOR2_X1 U16898 ( .A1(n19364), .A2(n13799), .ZN(n19281) );
  NOR2_X1 U16899 ( .A1(n19801), .A2(n19281), .ZN(n13800) );
  NAND2_X1 U16900 ( .A1(n12131), .A2(n13800), .ZN(n13808) );
  INV_X1 U16901 ( .A(n19281), .ZN(n13810) );
  NAND2_X1 U16902 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n13810), .ZN(n13805) );
  OAI21_X1 U16903 ( .B1(n19276), .B2(n19299), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n13803) );
  INV_X1 U16904 ( .A(n19304), .ZN(n13802) );
  NAND2_X1 U16905 ( .A1(n13802), .A2(n13801), .ZN(n19495) );
  OR2_X1 U16906 ( .A1(n19495), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n13806) );
  NAND2_X1 U16907 ( .A1(n13803), .A2(n13806), .ZN(n13804) );
  NAND4_X1 U16908 ( .A1(n13808), .A2(n19593), .A3(n13805), .A4(n13804), .ZN(
        n19283) );
  INV_X1 U16909 ( .A(n19283), .ZN(n13815) );
  INV_X1 U16910 ( .A(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n13814) );
  OAI21_X1 U16911 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n13806), .A(n19801), 
        .ZN(n13807) );
  INV_X1 U16912 ( .A(n19600), .ZN(n13811) );
  AOI22_X1 U16913 ( .A1(n19299), .A2(n19603), .B1(n19276), .B2(n19602), .ZN(
        n13809) );
  OAI21_X1 U16914 ( .B1(n13811), .B2(n13810), .A(n13809), .ZN(n13812) );
  AOI21_X1 U16915 ( .B1(n19282), .B2(n19601), .A(n13812), .ZN(n13813) );
  OAI21_X1 U16916 ( .B1(n13815), .B2(n13814), .A(n13813), .ZN(P2_U3080) );
  OAI21_X1 U16917 ( .B1(n13818), .B2(n13817), .A(n13816), .ZN(n16065) );
  NAND2_X1 U16918 ( .A1(n14786), .A2(n14788), .ZN(n13820) );
  XNOR2_X1 U16919 ( .A(n13819), .B(n13820), .ZN(n16067) );
  NAND2_X1 U16920 ( .A1(n16067), .A2(n12942), .ZN(n13831) );
  INV_X1 U16921 ( .A(n18885), .ZN(n13829) );
  INV_X1 U16922 ( .A(P2_REIP_REG_7__SCAN_IN), .ZN(n19692) );
  NOR2_X1 U16923 ( .A1(n13822), .A2(n16119), .ZN(n13821) );
  AOI21_X1 U16924 ( .B1(n16115), .B2(n13822), .A(n13821), .ZN(n13823) );
  OAI21_X1 U16925 ( .B1(n19692), .B2(n12482), .A(n13823), .ZN(n13828) );
  OR2_X1 U16926 ( .A1(n13825), .A2(n13824), .ZN(n13826) );
  NAND2_X1 U16927 ( .A1(n13826), .A2(n16112), .ZN(n18994) );
  NOR2_X1 U16928 ( .A1(n18994), .A2(n16128), .ZN(n13827) );
  AOI211_X1 U16929 ( .C1(n19131), .C2(n13829), .A(n13828), .B(n13827), .ZN(
        n13830) );
  OAI211_X1 U16930 ( .C1(n16065), .C2(n19125), .A(n13831), .B(n13830), .ZN(
        P2_U3039) );
  XNOR2_X1 U16931 ( .A(n13833), .B(n13832), .ZN(n14058) );
  OAI21_X1 U16932 ( .B1(n13835), .B2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A(
        n13834), .ZN(n14052) );
  INV_X1 U16933 ( .A(n14052), .ZN(n13841) );
  OAI22_X1 U16934 ( .A1(n13836), .A2(n19093), .B1(n11526), .B2(n12482), .ZN(
        n13840) );
  INV_X1 U16935 ( .A(n18900), .ZN(n13838) );
  OAI22_X1 U16936 ( .A1(n16063), .A2(n13838), .B1(n16072), .B2(n13837), .ZN(
        n13839) );
  AOI211_X1 U16937 ( .C1(n13841), .C2(n16068), .A(n13840), .B(n13839), .ZN(
        n13842) );
  OAI21_X1 U16938 ( .B1(n19088), .B2(n14058), .A(n13842), .ZN(P2_U3008) );
  XOR2_X1 U16939 ( .A(n13843), .B(n13734), .Z(n14937) );
  OR2_X1 U16940 ( .A1(n13739), .A2(n13845), .ZN(n13846) );
  NAND2_X1 U16941 ( .A1(n13844), .A2(n13846), .ZN(n14064) );
  OAI22_X1 U16942 ( .A1(n14691), .A2(n19157), .B1(n18995), .B2(n13847), .ZN(
        n13848) );
  AOI21_X1 U16943 ( .B1(n18965), .B2(BUF2_REG_19__SCAN_IN), .A(n13848), .ZN(
        n13850) );
  NAND2_X1 U16944 ( .A1(n18964), .A2(BUF1_REG_19__SCAN_IN), .ZN(n13849) );
  OAI211_X1 U16945 ( .C1(n14064), .C2(n19002), .A(n13850), .B(n13849), .ZN(
        n13851) );
  AOI21_X1 U16946 ( .B1(n14937), .B2(n19027), .A(n13851), .ZN(n13852) );
  INV_X1 U16947 ( .A(n13852), .ZN(P2_U2900) );
  AND2_X1 U16948 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(P3_EBX_REG_27__SCAN_IN), 
        .ZN(n16794) );
  INV_X2 U16949 ( .A(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n13943) );
  INV_X2 U16950 ( .A(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13853) );
  AOI22_X1 U16951 ( .A1(n17005), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n16974), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n13857) );
  NOR2_X2 U16952 ( .A1(n13861), .A2(n16741), .ZN(n15106) );
  AOI22_X1 U16953 ( .A1(n16992), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n17020), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n13856) );
  AOI22_X1 U16954 ( .A1(n16990), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n16923), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n13855) );
  NOR2_X2 U16955 ( .A1(n13859), .A2(n13860), .ZN(n16958) );
  INV_X2 U16956 ( .A(n14010), .ZN(n16998) );
  AOI22_X1 U16957 ( .A1(n16998), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n17014), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n13854) );
  NAND4_X1 U16958 ( .A1(n13857), .A2(n13856), .A3(n13855), .A4(n13854), .ZN(
        n13868) );
  INV_X4 U16959 ( .A(n13880), .ZN(n16989) );
  AOI22_X1 U16960 ( .A1(n16989), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n16975), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n13866) );
  AOI22_X1 U16961 ( .A1(n9633), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n17022), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n13865) );
  AOI22_X1 U16962 ( .A1(n16997), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n16995), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n13864) );
  INV_X2 U16963 ( .A(n13882), .ZN(n16991) );
  INV_X2 U16964 ( .A(n13882), .ZN(n17021) );
  AOI22_X1 U16965 ( .A1(n17021), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n16996), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n13863) );
  NAND4_X1 U16966 ( .A1(n13866), .A2(n13865), .A3(n13864), .A4(n13863), .ZN(
        n13867) );
  INV_X1 U16967 ( .A(P3_STATE2_REG_1__SCAN_IN), .ZN(n18650) );
  NAND2_X1 U16968 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n18650), .ZN(n18543) );
  INV_X1 U16969 ( .A(P3_STATE2_REG_2__SCAN_IN), .ZN(n18704) );
  NOR2_X1 U16970 ( .A1(n18543), .A2(n18704), .ZN(n18686) );
  BUF_X4 U16971 ( .A(n16825), .Z(n17020) );
  AOI22_X1 U16972 ( .A1(n17021), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n17020), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n13872) );
  AOI22_X1 U16973 ( .A1(n9633), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(n9626), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n13871) );
  AOI22_X1 U16975 ( .A1(n17023), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n17022), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n13870) );
  AOI22_X1 U16976 ( .A1(n17014), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n15158), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n13869) );
  NAND4_X1 U16977 ( .A1(n13872), .A2(n13871), .A3(n13870), .A4(n13869), .ZN(
        n13878) );
  AOI22_X1 U16978 ( .A1(n16977), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n16997), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n13876) );
  AOI22_X1 U16979 ( .A1(n17005), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n16992), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n13875) );
  AOI22_X1 U16980 ( .A1(n16974), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n16958), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n13874) );
  AOI22_X1 U16981 ( .A1(n16989), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n16995), .B2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n13873) );
  NAND4_X1 U16982 ( .A1(n13876), .A2(n13875), .A3(n13874), .A4(n13873), .ZN(
        n13877) );
  AOI22_X1 U16983 ( .A1(n16995), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n15158), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n13891) );
  AOI22_X1 U16984 ( .A1(n16997), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n17023), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n13890) );
  AOI22_X1 U16985 ( .A1(n16992), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n17020), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n13879) );
  OAI21_X1 U16986 ( .B1(n13880), .B2(n20830), .A(n13879), .ZN(n13888) );
  AOI22_X1 U16987 ( .A1(n9633), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n16923), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n13886) );
  AOI22_X1 U16988 ( .A1(n16977), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n16974), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n13885) );
  AOI22_X1 U16989 ( .A1(n16998), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n17022), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n13884) );
  AOI22_X1 U16990 ( .A1(n17021), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n17014), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n13883) );
  NAND4_X1 U16991 ( .A1(n13886), .A2(n13885), .A3(n13884), .A4(n13883), .ZN(
        n13887) );
  AOI22_X1 U16992 ( .A1(n16992), .A2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n16923), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n13895) );
  AOI22_X1 U16993 ( .A1(n16977), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n16989), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n13894) );
  AOI22_X1 U16994 ( .A1(n17005), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n15158), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n13893) );
  AOI22_X1 U16995 ( .A1(n16995), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n17014), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n13892) );
  NAND4_X1 U16996 ( .A1(n13895), .A2(n13894), .A3(n13893), .A4(n13892), .ZN(
        n13901) );
  AOI22_X1 U16997 ( .A1(n16998), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n17022), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n13899) );
  AOI22_X1 U16998 ( .A1(n9633), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n16975), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n13898) );
  AOI22_X1 U16999 ( .A1(n17021), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n17020), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n13897) );
  AOI22_X1 U17000 ( .A1(n16997), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n16974), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n13896) );
  NAND4_X1 U17001 ( .A1(n13899), .A2(n13898), .A3(n13897), .A4(n13896), .ZN(
        n13900) );
  AOI22_X1 U17002 ( .A1(n16989), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n17020), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n13905) );
  AOI22_X1 U17003 ( .A1(n17021), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n16975), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n13904) );
  AOI22_X1 U17004 ( .A1(n16995), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n17022), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n13903) );
  AOI22_X1 U17005 ( .A1(n16998), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n15174), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n13902) );
  NAND4_X1 U17006 ( .A1(n13905), .A2(n13904), .A3(n13903), .A4(n13902), .ZN(
        n13911) );
  AOI22_X1 U17007 ( .A1(n9633), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n16923), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n13909) );
  AOI22_X1 U17008 ( .A1(n16992), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n16974), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n13908) );
  AOI22_X1 U17009 ( .A1(n16977), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n16997), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n13907) );
  AOI22_X1 U17010 ( .A1(n17005), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n15158), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n13906) );
  NAND4_X1 U17011 ( .A1(n13909), .A2(n13908), .A3(n13907), .A4(n13906), .ZN(
        n13910) );
  AOI22_X1 U17012 ( .A1(n16997), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n16825), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n13915) );
  AOI22_X1 U17013 ( .A1(n17005), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n16992), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13914) );
  AOI22_X1 U17014 ( .A1(n16995), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n17022), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n13913) );
  AOI22_X1 U17015 ( .A1(n16974), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n17014), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n13912) );
  NAND4_X1 U17016 ( .A1(n13915), .A2(n13914), .A3(n13913), .A4(n13912), .ZN(
        n13921) );
  AOI22_X1 U17017 ( .A1(n16989), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n16991), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n13919) );
  AOI22_X1 U17018 ( .A1(n9633), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(n9626), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n13918) );
  AOI22_X1 U17019 ( .A1(n16977), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n15158), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n13917) );
  AOI22_X1 U17020 ( .A1(n16998), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n17023), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n13916) );
  NAND4_X1 U17021 ( .A1(n13919), .A2(n13918), .A3(n13917), .A4(n13916), .ZN(
        n13920) );
  NOR2_X1 U17022 ( .A1(n17078), .A2(n17082), .ZN(n15052) );
  INV_X1 U17023 ( .A(n15052), .ZN(n15050) );
  AOI22_X1 U17024 ( .A1(n16996), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n17023), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n13925) );
  AOI22_X1 U17025 ( .A1(n16974), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n17022), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n13924) );
  AOI22_X1 U17026 ( .A1(n16977), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n16825), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n13923) );
  AOI22_X1 U17027 ( .A1(n16923), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n17014), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n13922) );
  NAND4_X1 U17028 ( .A1(n13925), .A2(n13924), .A3(n13923), .A4(n13922), .ZN(
        n13932) );
  AOI22_X1 U17029 ( .A1(n16992), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n17021), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n13930) );
  AOI22_X1 U17030 ( .A1(n16989), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n16995), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n13929) );
  AOI22_X1 U17031 ( .A1(n16998), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n9633), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n13928) );
  AOI22_X1 U17032 ( .A1(n17005), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n16997), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n13927) );
  NAND4_X1 U17033 ( .A1(n13930), .A2(n13929), .A3(n13928), .A4(n13927), .ZN(
        n13931) );
  AOI22_X1 U17034 ( .A1(n16974), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n17021), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n13936) );
  AOI22_X1 U17035 ( .A1(n16977), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n9626), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n13935) );
  AOI22_X1 U17036 ( .A1(n16992), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n16989), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n13934) );
  AOI22_X1 U17037 ( .A1(n17020), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n17014), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n13933) );
  NAND4_X1 U17038 ( .A1(n13936), .A2(n13935), .A3(n13934), .A4(n13933), .ZN(
        n13942) );
  AOI22_X1 U17039 ( .A1(n16995), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n17022), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n13940) );
  AOI22_X1 U17040 ( .A1(n9633), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n15158), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n13939) );
  AOI22_X1 U17041 ( .A1(n17005), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n16997), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n13938) );
  AOI22_X1 U17042 ( .A1(n16998), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n17023), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n13937) );
  NAND4_X1 U17043 ( .A1(n13940), .A2(n13939), .A3(n13938), .A4(n13937), .ZN(
        n13941) );
  NAND2_X1 U17044 ( .A1(n15076), .A2(n15221), .ZN(n18494) );
  NOR2_X1 U17045 ( .A1(n15050), .A2(n18494), .ZN(n15078) );
  NAND3_X1 U17046 ( .A1(n18068), .A2(n15078), .A3(n18087), .ZN(n13954) );
  AOI22_X1 U17047 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B1(n18517), .B2(n13853), .ZN(
        n15061) );
  INV_X1 U17048 ( .A(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n18044) );
  AOI22_X1 U17049 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n18522), .B1(
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n13943), .ZN(n13948) );
  NAND2_X1 U17050 ( .A1(n18515), .A2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n15060) );
  OAI21_X1 U17051 ( .B1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n13853), .A(
        n13944), .ZN(n13949) );
  NAND2_X1 U17052 ( .A1(n13948), .A2(n13949), .ZN(n13945) );
  OAI21_X1 U17053 ( .B1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n13943), .A(
        n13945), .ZN(n13946) );
  OAI22_X1 U17054 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n18044), .B1(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n13946), .ZN(n13951) );
  NOR2_X1 U17055 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n18044), .ZN(
        n13947) );
  NAND2_X1 U17056 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n13946), .ZN(
        n13950) );
  AOI22_X1 U17057 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n13951), .B1(
        n13947), .B2(n13950), .ZN(n13953) );
  OAI211_X1 U17058 ( .C1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .C2(n18515), .A(
        n13953), .B(n15060), .ZN(n15218) );
  XOR2_X1 U17059 ( .A(n13949), .B(n13948), .Z(n15219) );
  INV_X1 U17060 ( .A(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n16701) );
  AND2_X1 U17061 ( .A1(n13950), .A2(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n13952) );
  OAI22_X1 U17062 ( .A1(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n16701), .B1(
        n13952), .B2(n13951), .ZN(n15064) );
  AOI21_X1 U17063 ( .B1(n13953), .B2(n15219), .A(n15064), .ZN(n15062) );
  OAI21_X1 U17064 ( .B1(n15061), .B2(n15218), .A(n15062), .ZN(n16155) );
  INV_X1 U17065 ( .A(n16155), .ZN(n18485) );
  NAND2_X1 U17066 ( .A1(n15221), .A2(n17082), .ZN(n15227) );
  NAND2_X1 U17067 ( .A1(n18485), .A2(n15235), .ZN(n15085) );
  NAND2_X1 U17068 ( .A1(n13954), .A2(n15085), .ZN(n15429) );
  NAND4_X1 U17069 ( .A1(n18686), .A2(n17291), .A3(n17227), .A4(n15429), .ZN(
        n13955) );
  INV_X1 U17070 ( .A(n13955), .ZN(n17073) );
  NAND2_X1 U17071 ( .A1(n18087), .A2(n17073), .ZN(n17067) );
  INV_X1 U17072 ( .A(n18087), .ZN(n17123) );
  INV_X2 U17073 ( .A(n17070), .ZN(n17064) );
  INV_X1 U17074 ( .A(P3_EBX_REG_22__SCAN_IN), .ZN(n13956) );
  INV_X1 U17075 ( .A(P3_EBX_REG_18__SCAN_IN), .ZN(n16888) );
  INV_X1 U17076 ( .A(P3_EBX_REG_17__SCAN_IN), .ZN(n16904) );
  INV_X1 U17077 ( .A(P3_EBX_REG_15__SCAN_IN), .ZN(n16563) );
  INV_X1 U17078 ( .A(P3_EBX_REG_13__SCAN_IN), .ZN(n16593) );
  INV_X1 U17079 ( .A(P3_EBX_REG_12__SCAN_IN), .ZN(n16970) );
  INV_X1 U17080 ( .A(P3_EBX_REG_2__SCAN_IN), .ZN(n16725) );
  NAND2_X1 U17081 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .ZN(n17062) );
  NOR2_X1 U17082 ( .A1(n16725), .A2(n17062), .ZN(n17049) );
  NAND3_X1 U17083 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(P3_EBX_REG_3__SCAN_IN), 
        .A3(n17049), .ZN(n17048) );
  NAND4_X1 U17084 ( .A1(P3_EBX_REG_11__SCAN_IN), .A2(P3_EBX_REG_10__SCAN_IN), 
        .A3(P3_EBX_REG_9__SCAN_IN), .A4(P3_EBX_REG_8__SCAN_IN), .ZN(n16946) );
  NAND2_X1 U17085 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n16944), .ZN(n16943) );
  NAND2_X1 U17086 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n16932), .ZN(n16892) );
  NAND3_X1 U17087 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(P3_EBX_REG_19__SCAN_IN), 
        .A3(n16874), .ZN(n16848) );
  NOR2_X1 U17088 ( .A1(n17123), .A2(n16848), .ZN(n16850) );
  NAND2_X1 U17089 ( .A1(P3_EBX_REG_21__SCAN_IN), .A2(n16850), .ZN(n16837) );
  NAND3_X1 U17090 ( .A1(P3_EBX_REG_25__SCAN_IN), .A2(P3_EBX_REG_24__SCAN_IN), 
        .A3(n16821), .ZN(n16800) );
  NAND2_X1 U17091 ( .A1(n17064), .A2(n16805), .ZN(n13957) );
  OAI21_X1 U17092 ( .B1(n16794), .B2(n17067), .A(n13957), .ZN(n16795) );
  AOI22_X1 U17093 ( .A1(n16992), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n16974), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n13961) );
  AOI22_X1 U17094 ( .A1(n16995), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n9633), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n13960) );
  AOI22_X1 U17095 ( .A1(n16997), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n16998), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n13959) );
  AOI22_X1 U17096 ( .A1(n17021), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n17014), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n13958) );
  NAND4_X1 U17097 ( .A1(n13961), .A2(n13960), .A3(n13959), .A4(n13958), .ZN(
        n13968) );
  AOI22_X1 U17098 ( .A1(n17020), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n15158), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n13966) );
  AOI22_X1 U17099 ( .A1(n16923), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n17022), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n13965) );
  AOI22_X1 U17100 ( .A1(n17005), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n17023), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n13964) );
  AOI22_X1 U17101 ( .A1(n16977), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n16989), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n13963) );
  NAND4_X1 U17102 ( .A1(n13966), .A2(n13965), .A3(n13964), .A4(n13963), .ZN(
        n13967) );
  NOR2_X1 U17103 ( .A1(n13968), .A2(n13967), .ZN(n14030) );
  AOI22_X1 U17104 ( .A1(n16974), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n17022), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n13972) );
  AOI22_X1 U17105 ( .A1(n16995), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n17021), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n13971) );
  AOI22_X1 U17106 ( .A1(n16992), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n16998), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n13970) );
  AOI22_X1 U17107 ( .A1(n17014), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n17023), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n13969) );
  NAND4_X1 U17108 ( .A1(n13972), .A2(n13971), .A3(n13970), .A4(n13969), .ZN(
        n13978) );
  AOI22_X1 U17109 ( .A1(n16977), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n9633), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n13976) );
  AOI22_X1 U17110 ( .A1(n16997), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n9626), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n13975) );
  AOI22_X1 U17111 ( .A1(n17005), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n15158), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n13974) );
  AOI22_X1 U17112 ( .A1(n16989), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n16825), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n13973) );
  NAND4_X1 U17113 ( .A1(n13976), .A2(n13975), .A3(n13974), .A4(n13973), .ZN(
        n13977) );
  NOR2_X1 U17114 ( .A1(n13978), .A2(n13977), .ZN(n16803) );
  AOI22_X1 U17115 ( .A1(n16992), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_12__1__SCAN_IN), .B2(n16996), .ZN(n13982) );
  AOI22_X1 U17116 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n17020), .B1(
        P3_INSTQUEUE_REG_5__1__SCAN_IN), .B2(n17021), .ZN(n13981) );
  AOI22_X1 U17117 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n16923), .B1(
        P3_INSTQUEUE_REG_8__1__SCAN_IN), .B2(n17022), .ZN(n13980) );
  AOI22_X1 U17118 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n16977), .B1(
        P3_INSTQUEUE_REG_2__1__SCAN_IN), .B2(n17014), .ZN(n13979) );
  NAND4_X1 U17119 ( .A1(n13982), .A2(n13981), .A3(n13980), .A4(n13979), .ZN(
        n13988) );
  AOI22_X1 U17120 ( .A1(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n17023), .B1(
        n9633), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n13986) );
  AOI22_X1 U17121 ( .A1(P3_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n16924), .B1(
        n16997), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n13985) );
  AOI22_X1 U17122 ( .A1(n17005), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n16998), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n13984) );
  AOI22_X1 U17123 ( .A1(n16989), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n16974), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n13983) );
  NAND4_X1 U17124 ( .A1(n13986), .A2(n13985), .A3(n13984), .A4(n13983), .ZN(
        n13987) );
  NOR2_X1 U17125 ( .A1(n13988), .A2(n13987), .ZN(n16812) );
  AOI22_X1 U17126 ( .A1(n16977), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n16998), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n13998) );
  AOI22_X1 U17127 ( .A1(n17005), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n16825), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n13997) );
  AOI22_X1 U17128 ( .A1(n16923), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n17023), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n13989) );
  OAI21_X1 U17129 ( .B1(n13882), .B2(n20830), .A(n13989), .ZN(n13995) );
  AOI22_X1 U17130 ( .A1(n16989), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n15158), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n13993) );
  AOI22_X1 U17131 ( .A1(n16997), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n16974), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n13992) );
  AOI22_X1 U17132 ( .A1(n16995), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n17022), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n13991) );
  AOI22_X1 U17133 ( .A1(n16992), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n17014), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n13990) );
  NAND4_X1 U17134 ( .A1(n13993), .A2(n13992), .A3(n13991), .A4(n13990), .ZN(
        n13994) );
  AOI211_X1 U17135 ( .C1(n9633), .C2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .A(
        n13995), .B(n13994), .ZN(n13996) );
  NAND3_X1 U17136 ( .A1(n13998), .A2(n13997), .A3(n13996), .ZN(n16818) );
  AOI22_X1 U17137 ( .A1(n16997), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n16825), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n14008) );
  AOI22_X1 U17138 ( .A1(n16996), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n17023), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n14007) );
  INV_X1 U17139 ( .A(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n17039) );
  AOI22_X1 U17140 ( .A1(n17021), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n17022), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n13999) );
  OAI21_X1 U17141 ( .B1(n14010), .B2(n17039), .A(n13999), .ZN(n14005) );
  AOI22_X1 U17142 ( .A1(n17005), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n16977), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n14003) );
  AOI22_X1 U17143 ( .A1(n16989), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n9626), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n14002) );
  AOI22_X1 U17144 ( .A1(n16995), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n9633), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n14001) );
  AOI22_X1 U17145 ( .A1(n9627), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n17014), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n14000) );
  NAND4_X1 U17146 ( .A1(n14003), .A2(n14002), .A3(n14001), .A4(n14000), .ZN(
        n14004) );
  AOI211_X1 U17147 ( .C1(n16992), .C2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A(
        n14005), .B(n14004), .ZN(n14006) );
  NAND3_X1 U17148 ( .A1(n14008), .A2(n14007), .A3(n14006), .ZN(n16819) );
  NAND2_X1 U17149 ( .A1(n16818), .A2(n16819), .ZN(n16817) );
  NOR2_X1 U17150 ( .A1(n16812), .A2(n16817), .ZN(n16811) );
  AOI22_X1 U17151 ( .A1(n16992), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n16974), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n14019) );
  AOI22_X1 U17152 ( .A1(n16997), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n17021), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n14018) );
  INV_X1 U17153 ( .A(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n17061) );
  AOI22_X1 U17154 ( .A1(n16923), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n17022), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n14009) );
  OAI21_X1 U17155 ( .B1(n16824), .B2(n17061), .A(n14009), .ZN(n14016) );
  AOI22_X1 U17156 ( .A1(n16977), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n16989), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n14014) );
  AOI22_X1 U17157 ( .A1(n17020), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n17023), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n14013) );
  AOI22_X1 U17158 ( .A1(n17005), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n17013), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n14012) );
  AOI22_X1 U17159 ( .A1(n17014), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n15158), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n14011) );
  NAND4_X1 U17160 ( .A1(n14014), .A2(n14013), .A3(n14012), .A4(n14011), .ZN(
        n14015) );
  AOI211_X1 U17161 ( .C1(n9633), .C2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .A(
        n14016), .B(n14015), .ZN(n14017) );
  NAND3_X1 U17162 ( .A1(n14019), .A2(n14018), .A3(n14017), .ZN(n16808) );
  NAND2_X1 U17163 ( .A1(n16811), .A2(n16808), .ZN(n16807) );
  NOR2_X1 U17164 ( .A1(n16803), .A2(n16807), .ZN(n16802) );
  AOI22_X1 U17165 ( .A1(n16923), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n15158), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n14029) );
  AOI22_X1 U17166 ( .A1(n16997), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n16974), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n14028) );
  INV_X1 U17167 ( .A(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n17051) );
  AOI22_X1 U17168 ( .A1(n17014), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n17022), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n14020) );
  OAI21_X1 U17169 ( .B1(n16824), .B2(n17051), .A(n14020), .ZN(n14026) );
  AOI22_X1 U17170 ( .A1(n16977), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n9633), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n14024) );
  AOI22_X1 U17171 ( .A1(n17021), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n16825), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n14023) );
  AOI22_X1 U17172 ( .A1(n17005), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n17013), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n14022) );
  AOI22_X1 U17173 ( .A1(n16989), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n17023), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n14021) );
  NAND4_X1 U17174 ( .A1(n14024), .A2(n14023), .A3(n14022), .A4(n14021), .ZN(
        n14025) );
  AOI211_X1 U17175 ( .C1(n16992), .C2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .A(
        n14026), .B(n14025), .ZN(n14027) );
  NAND3_X1 U17176 ( .A1(n14029), .A2(n14028), .A3(n14027), .ZN(n16798) );
  NAND2_X1 U17177 ( .A1(n16802), .A2(n16798), .ZN(n16797) );
  NOR2_X1 U17178 ( .A1(n14030), .A2(n16797), .ZN(n16792) );
  AOI21_X1 U17179 ( .B1(n14030), .B2(n16797), .A(n16792), .ZN(n17091) );
  AOI22_X1 U17180 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n16795), .B1(n17091), 
        .B2(n17070), .ZN(n14034) );
  INV_X1 U17181 ( .A(P3_EBX_REG_28__SCAN_IN), .ZN(n14032) );
  INV_X1 U17182 ( .A(n16805), .ZN(n14031) );
  NAND3_X1 U17183 ( .A1(P3_EBX_REG_27__SCAN_IN), .A2(n14032), .A3(n14031), 
        .ZN(n14033) );
  NAND2_X1 U17184 ( .A1(n14034), .A2(n14033), .ZN(P3_U2675) );
  XNOR2_X1 U17185 ( .A(n15569), .B(n15833), .ZN(n14035) );
  XNOR2_X1 U17186 ( .A(n14036), .B(n14035), .ZN(n15828) );
  AOI22_X1 U17187 ( .A1(n20034), .A2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .B1(
        n20043), .B2(P1_REIP_REG_9__SCAN_IN), .ZN(n14037) );
  OAI21_X1 U17188 ( .B1(n20032), .B2(n14038), .A(n14037), .ZN(n14039) );
  AOI21_X1 U17189 ( .B1(n19843), .B2(n15645), .A(n14039), .ZN(n14040) );
  OAI21_X1 U17190 ( .B1(n20031), .B2(n15828), .A(n14040), .ZN(P1_U2990) );
  AND2_X1 U17191 ( .A1(n9710), .A2(n14041), .ZN(n14043) );
  OR2_X1 U17192 ( .A1(n14043), .A2(n14042), .ZN(n18776) );
  NOR2_X1 U17193 ( .A1(n15938), .A2(n18776), .ZN(n14044) );
  AOI21_X1 U17194 ( .B1(P2_EBX_REG_17__SCAN_IN), .B2(n15938), .A(n14044), .ZN(
        n14045) );
  OAI21_X1 U17195 ( .B1(n14046), .B2(n18952), .A(n14045), .ZN(P2_U2870) );
  XNOR2_X1 U17196 ( .A(n14047), .B(n14048), .ZN(n18996) );
  NAND2_X1 U17197 ( .A1(n14049), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n14051) );
  AOI22_X1 U17198 ( .A1(n19131), .A2(n18901), .B1(n19081), .B2(
        P2_REIP_REG_6__SCAN_IN), .ZN(n14050) );
  OAI211_X1 U17199 ( .C1(n16128), .C2(n18996), .A(n14051), .B(n14050), .ZN(
        n14054) );
  NOR2_X1 U17200 ( .A1(n14052), .A2(n19125), .ZN(n14053) );
  AOI211_X1 U17201 ( .C1(n14056), .C2(n14055), .A(n14054), .B(n14053), .ZN(
        n14057) );
  OAI21_X1 U17202 ( .B1(n19110), .B2(n14058), .A(n14057), .ZN(P2_U3040) );
  NAND2_X1 U17203 ( .A1(n14059), .A2(n14060), .ZN(n14061) );
  NAND2_X1 U17204 ( .A1(n14757), .A2(n14061), .ZN(n14938) );
  MUX2_X1 U17205 ( .A(n14062), .B(n14938), .S(n18958), .Z(n14063) );
  OAI21_X1 U17206 ( .B1(n14064), .B2(n18952), .A(n14063), .ZN(P2_U2868) );
  INV_X1 U17207 ( .A(n14937), .ZN(n14076) );
  INV_X1 U17208 ( .A(n14938), .ZN(n14070) );
  NAND2_X1 U17209 ( .A1(P2_EBX_REG_19__SCAN_IN), .A2(n18842), .ZN(n14065) );
  OAI211_X1 U17210 ( .C1(n20894), .C2(n18935), .A(n16114), .B(n14065), .ZN(
        n14066) );
  AOI21_X1 U17211 ( .B1(n14067), .B2(n18896), .A(n14066), .ZN(n14068) );
  OAI21_X1 U17212 ( .B1(n19713), .B2(n18932), .A(n14068), .ZN(n14069) );
  AOI21_X1 U17213 ( .B1(n14070), .B2(n18916), .A(n14069), .ZN(n14075) );
  AOI211_X1 U17214 ( .C1(n14769), .C2(n14072), .A(n14071), .B(n18890), .ZN(
        n14073) );
  INV_X1 U17215 ( .A(n14073), .ZN(n14074) );
  OAI211_X1 U17216 ( .C1(n14076), .C2(n18928), .A(n14075), .B(n14074), .ZN(
        P2_U2836) );
  OAI21_X1 U17217 ( .B1(n9735), .B2(n10120), .A(n15936), .ZN(n14639) );
  OR2_X1 U17218 ( .A1(n14078), .A2(n9656), .ZN(n14080) );
  INV_X1 U17219 ( .A(n14912), .ZN(n14079) );
  AND2_X1 U17220 ( .A1(n14080), .A2(n14079), .ZN(n18743) );
  OAI22_X1 U17221 ( .A1(n14691), .A2(n19168), .B1(n14081), .B2(n18995), .ZN(
        n14082) );
  AOI21_X1 U17222 ( .B1(n19027), .B2(n18743), .A(n14082), .ZN(n14084) );
  AOI22_X1 U17223 ( .A1(n18965), .A2(BUF2_REG_21__SCAN_IN), .B1(n18964), .B2(
        BUF1_REG_21__SCAN_IN), .ZN(n14083) );
  OAI211_X1 U17224 ( .C1(n14639), .C2(n19002), .A(n14084), .B(n14083), .ZN(
        P2_U2898) );
  OAI21_X1 U17225 ( .B1(n9605), .B2(n14085), .A(n14090), .ZN(n14092) );
  XNOR2_X1 U17226 ( .A(n14092), .B(n14089), .ZN(n15644) );
  INV_X1 U17227 ( .A(n15644), .ZN(n14088) );
  MUX2_X1 U17228 ( .A(DATAI_11_), .B(BUF1_REG_11__SCAN_IN), .S(n20085), .Z(
        n20005) );
  INV_X1 U17229 ( .A(n20005), .ZN(n14086) );
  OAI222_X1 U17230 ( .A1(n14088), .A2(n14396), .B1(n14436), .B2(n14087), .C1(
        n14086), .C2(n14144), .ZN(P1_U2893) );
  INV_X1 U17231 ( .A(n14089), .ZN(n14091) );
  OAI21_X1 U17232 ( .B1(n14092), .B2(n14091), .A(n14090), .ZN(n14094) );
  NAND2_X1 U17233 ( .A1(n14094), .A2(n14093), .ZN(n14124) );
  OAI21_X1 U17234 ( .B1(n14094), .B2(n14093), .A(n14124), .ZN(n15536) );
  MUX2_X1 U17235 ( .A(DATAI_12_), .B(BUF1_REG_12__SCAN_IN), .S(n20085), .Z(
        n20007) );
  AOI22_X1 U17236 ( .A1(n14095), .A2(n20007), .B1(P1_EAX_REG_12__SCAN_IN), 
        .B2(n14421), .ZN(n14096) );
  OAI21_X1 U17237 ( .B1(n15536), .B2(n14396), .A(n14096), .ZN(P1_U2892) );
  OR2_X1 U17238 ( .A1(n15546), .A2(n14097), .ZN(n14098) );
  NAND2_X1 U17239 ( .A1(n14132), .A2(n14098), .ZN(n15810) );
  INV_X1 U17240 ( .A(n15810), .ZN(n14099) );
  AOI22_X1 U17241 ( .A1(n19940), .A2(n14099), .B1(n10965), .B2(
        P1_EBX_REG_12__SCAN_IN), .ZN(n14100) );
  OAI21_X1 U17242 ( .B1(n15536), .B2(n9630), .A(n14100), .ZN(P1_U2860) );
  NOR2_X1 U17243 ( .A1(n9702), .A2(n14101), .ZN(n14102) );
  OR2_X1 U17244 ( .A1(n9706), .A2(n14102), .ZN(n15624) );
  XNOR2_X1 U17245 ( .A(n14134), .B(n14118), .ZN(n15777) );
  AOI22_X1 U17246 ( .A1(n19940), .A2(n15777), .B1(n10965), .B2(
        P1_EBX_REG_14__SCAN_IN), .ZN(n14103) );
  OAI21_X1 U17247 ( .B1(n15624), .B2(n9630), .A(n14103), .ZN(P1_U2858) );
  AND2_X1 U17248 ( .A1(n19922), .A2(n14285), .ZN(n15472) );
  AOI221_X1 U17249 ( .B1(n19875), .B2(n20637), .C1(n14104), .C2(n20637), .A(
        n15472), .ZN(n14110) );
  NAND2_X1 U17250 ( .A1(n15777), .A2(n19905), .ZN(n14105) );
  OAI211_X1 U17251 ( .C1(n14106), .C2(n19867), .A(n14105), .B(n19879), .ZN(
        n14109) );
  INV_X1 U17252 ( .A(n15625), .ZN(n14107) );
  OAI22_X1 U17253 ( .A1(n10585), .A2(n19923), .B1(n19897), .B2(n14107), .ZN(
        n14108) );
  AOI211_X1 U17254 ( .C1(n14110), .C2(n19930), .A(n14109), .B(n14108), .ZN(
        n14111) );
  OAI21_X1 U17255 ( .B1(n15624), .B2(n19861), .A(n14111), .ZN(P1_U2826) );
  MUX2_X1 U17256 ( .A(DATAI_14_), .B(BUF1_REG_14__SCAN_IN), .S(n20085), .Z(
        n20011) );
  INV_X1 U17257 ( .A(n20011), .ZN(n14112) );
  OAI222_X1 U17258 ( .A1(n15624), .A2(n14396), .B1(n14436), .B2(n14113), .C1(
        n14144), .C2(n14112), .ZN(P1_U2890) );
  OAI21_X1 U17259 ( .B1(n9706), .B2(n14116), .A(n14114), .ZN(n14528) );
  INV_X1 U17260 ( .A(n14134), .ZN(n14119) );
  AOI21_X1 U17261 ( .B1(n14119), .B2(n14118), .A(n14117), .ZN(n14120) );
  OR2_X1 U17262 ( .A1(n14120), .A2(n15531), .ZN(n14289) );
  INV_X1 U17263 ( .A(n14289), .ZN(n15766) );
  AOI22_X1 U17264 ( .A1(n15766), .A2(n19940), .B1(n10965), .B2(
        P1_EBX_REG_15__SCAN_IN), .ZN(n14121) );
  OAI21_X1 U17265 ( .B1(n14528), .B2(n9630), .A(n14121), .ZN(P1_U2857) );
  INV_X1 U17266 ( .A(n14122), .ZN(n14123) );
  AOI21_X1 U17267 ( .B1(n14124), .B2(n14123), .A(n9702), .ZN(n14539) );
  INV_X1 U17268 ( .A(n14539), .ZN(n14142) );
  INV_X1 U17269 ( .A(n14125), .ZN(n14127) );
  AOI21_X1 U17270 ( .B1(n14127), .B2(n14126), .A(n15471), .ZN(n15539) );
  NAND2_X1 U17271 ( .A1(n19920), .A2(n14128), .ZN(n14130) );
  AOI22_X1 U17272 ( .A1(n19935), .A2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .B1(
        n19929), .B2(P1_EBX_REG_13__SCAN_IN), .ZN(n14129) );
  OAI21_X1 U17273 ( .B1(P1_REIP_REG_13__SCAN_IN), .B2(n14130), .A(n14129), 
        .ZN(n14137) );
  NAND2_X1 U17274 ( .A1(n14132), .A2(n14131), .ZN(n14133) );
  AND2_X1 U17275 ( .A1(n14134), .A2(n14133), .ZN(n15790) );
  AOI21_X1 U17276 ( .B1(n19905), .B2(n15790), .A(n19891), .ZN(n14135) );
  OAI21_X1 U17277 ( .B1(n14537), .B2(n19897), .A(n14135), .ZN(n14136) );
  AOI211_X1 U17278 ( .C1(n15539), .C2(P1_REIP_REG_13__SCAN_IN), .A(n14137), 
        .B(n14136), .ZN(n14138) );
  OAI21_X1 U17279 ( .B1(n14142), .B2(n19861), .A(n14138), .ZN(P1_U2827) );
  AOI22_X1 U17280 ( .A1(n19940), .A2(n15790), .B1(n10965), .B2(
        P1_EBX_REG_13__SCAN_IN), .ZN(n14139) );
  OAI21_X1 U17281 ( .B1(n14142), .B2(n9630), .A(n14139), .ZN(P1_U2859) );
  MUX2_X1 U17282 ( .A(DATAI_13_), .B(BUF1_REG_13__SCAN_IN), .S(n20085), .Z(
        n20009) );
  INV_X1 U17283 ( .A(n20009), .ZN(n14140) );
  OAI222_X1 U17284 ( .A1(n14142), .A2(n14396), .B1(n14436), .B2(n14141), .C1(
        n14140), .C2(n14144), .ZN(P1_U2891) );
  OAI222_X1 U17285 ( .A1(n14528), .A2(n14396), .B1(n14144), .B2(n14143), .C1(
        n14436), .C2(n13278), .ZN(P1_U2889) );
  AOI22_X1 U17286 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n17022), .B1(
        P3_INSTQUEUE_REG_3__1__SCAN_IN), .B2(n17021), .ZN(n14154) );
  AOI22_X1 U17287 ( .A1(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n17013), .B1(
        P3_INSTQUEUE_REG_5__1__SCAN_IN), .B2(n16923), .ZN(n14153) );
  INV_X1 U17288 ( .A(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n17065) );
  AOI22_X1 U17289 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n16996), .B1(
        n16995), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n14145) );
  OAI21_X1 U17290 ( .B1(n17065), .B2(n16994), .A(n14145), .ZN(n14151) );
  AOI22_X1 U17291 ( .A1(n16997), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_13__1__SCAN_IN), .B2(n17023), .ZN(n14149) );
  AOI22_X1 U17292 ( .A1(n16992), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n16974), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n14148) );
  AOI22_X1 U17293 ( .A1(n16990), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n16989), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n14147) );
  AOI22_X1 U17294 ( .A1(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n9633), .B1(
        n17020), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n14146) );
  NAND4_X1 U17295 ( .A1(n14149), .A2(n14148), .A3(n14147), .A4(n14146), .ZN(
        n14150) );
  AOI211_X1 U17296 ( .C1(n17005), .C2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A(
        n14151), .B(n14150), .ZN(n14152) );
  NAND3_X1 U17297 ( .A1(n14154), .A2(n14153), .A3(n14152), .ZN(n17184) );
  INV_X1 U17298 ( .A(P3_EBX_REG_9__SCAN_IN), .ZN(n16640) );
  INV_X1 U17299 ( .A(P3_EBX_REG_8__SCAN_IN), .ZN(n17033) );
  NOR3_X1 U17300 ( .A1(n17032), .A2(n16640), .A3(n17033), .ZN(n17009) );
  INV_X1 U17301 ( .A(n17032), .ZN(n17031) );
  AOI21_X1 U17302 ( .B1(P3_EBX_REG_8__SCAN_IN), .B2(n17031), .A(
        P3_EBX_REG_9__SCAN_IN), .ZN(n14155) );
  NOR2_X1 U17303 ( .A1(n17009), .A2(n14155), .ZN(n14156) );
  MUX2_X1 U17304 ( .A(n17184), .B(n14156), .S(n17064), .Z(P3_U2694) );
  NAND3_X1 U17305 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_STATE2_REG_0__SCAN_IN), .A3(P3_STATE2_REG_2__SCAN_IN), .ZN(n18638)
         );
  NAND2_X1 U17306 ( .A1(n15090), .A2(n16701), .ZN(n14157) );
  NOR2_X1 U17307 ( .A1(n16958), .A2(n14157), .ZN(n18036) );
  INV_X1 U17308 ( .A(P3_FLUSH_REG_SCAN_IN), .ZN(n16350) );
  INV_X1 U17309 ( .A(P3_STATE2_REG_0__SCAN_IN), .ZN(n18636) );
  NOR2_X1 U17310 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n18639), .ZN(
        n18663) );
  NOR2_X1 U17311 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n18696) );
  AOI21_X1 U17312 ( .B1(P3_STATE2_REG_2__SCAN_IN), .B2(
        P3_STATE2_REG_1__SCAN_IN), .A(n18696), .ZN(n18550) );
  OR2_X1 U17313 ( .A1(n18663), .A2(n18550), .ZN(n18045) );
  NAND2_X1 U17314 ( .A1(n18636), .A2(n18045), .ZN(n18083) );
  OAI221_X1 U17315 ( .B1(n18638), .B2(n18036), .C1(n18638), .C2(n16350), .A(
        n18083), .ZN(n18043) );
  INV_X1 U17316 ( .A(n18043), .ZN(n18039) );
  NAND2_X1 U17317 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_STATEBS16_REG_SCAN_IN), .ZN(n17668) );
  INV_X1 U17318 ( .A(n17668), .ZN(n17464) );
  NOR2_X1 U17319 ( .A1(n18650), .A2(n18704), .ZN(n18035) );
  NOR2_X1 U17320 ( .A1(P3_STATE2_REG_3__SCAN_IN), .A2(n18035), .ZN(n18037) );
  INV_X1 U17321 ( .A(n18037), .ZN(n18685) );
  NOR2_X1 U17322 ( .A1(n17464), .A2(n18685), .ZN(n15047) );
  AOI21_X1 U17323 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(n15047), .ZN(n15048) );
  NOR2_X1 U17324 ( .A1(n18039), .A2(n15048), .ZN(n14159) );
  INV_X1 U17325 ( .A(P3_STATEBS16_REG_SCAN_IN), .ZN(n18691) );
  NOR3_X1 U17326 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(P3_STATE2_REG_3__SCAN_IN), .A3(n18691), .ZN(n16171) );
  NAND2_X1 U17327 ( .A1(P3_STATE2_REG_3__SCAN_IN), .A2(n18515), .ZN(n18091) );
  NAND2_X1 U17328 ( .A1(n18091), .A2(n18043), .ZN(n15046) );
  OR2_X1 U17329 ( .A1(n16171), .A2(n15046), .ZN(n14158) );
  MUX2_X1 U17330 ( .A(n14159), .B(n14158), .S(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .Z(P3_U2864) );
  NOR2_X1 U17331 ( .A1(n14160), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n14161) );
  OR2_X1 U17332 ( .A1(n14162), .A2(n14161), .ZN(n16137) );
  INV_X1 U17333 ( .A(n16137), .ZN(n14165) );
  NOR2_X1 U17334 ( .A1(n16114), .A2(n11633), .ZN(n16140) );
  OAI21_X1 U17335 ( .B1(n18921), .B2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n14163), .ZN(n16138) );
  NOR2_X1 U17336 ( .A1(n19088), .A2(n16138), .ZN(n14164) );
  AOI211_X1 U17337 ( .C1(n16068), .C2(n14165), .A(n16140), .B(n14164), .ZN(
        n14168) );
  OAI21_X1 U17338 ( .B1(n16001), .B2(n14166), .A(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n14167) );
  OAI211_X1 U17339 ( .C1(n16072), .C2(n18925), .A(n14168), .B(n14167), .ZN(
        P2_U3014) );
  XNOR2_X1 U17340 ( .A(n14170), .B(n14169), .ZN(n14175) );
  OR2_X1 U17341 ( .A1(n13360), .A2(n14171), .ZN(n14173) );
  NAND2_X1 U17342 ( .A1(n14173), .A2(n14172), .ZN(n18824) );
  MUX2_X1 U17343 ( .A(n11552), .B(n18824), .S(n18958), .Z(n14174) );
  OAI21_X1 U17344 ( .B1(n14175), .B2(n18952), .A(n14174), .ZN(P2_U2874) );
  INV_X1 U17345 ( .A(n20181), .ZN(n20699) );
  INV_X1 U17346 ( .A(n14176), .ZN(n14178) );
  AOI22_X1 U17347 ( .A1(n20699), .A2(n14178), .B1(n14177), .B2(n10132), .ZN(
        n15327) );
  INV_X1 U17348 ( .A(n15327), .ZN(n14181) );
  OAI22_X1 U17349 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n14179), .B1(
        P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n13663), .ZN(n14180) );
  AOI21_X1 U17350 ( .B1(n14181), .B2(n15857), .A(n14180), .ZN(n14185) );
  AOI21_X1 U17351 ( .B1(n14182), .B2(n15857), .A(n14184), .ZN(n14183) );
  OAI22_X1 U17352 ( .A1(n14185), .A2(n14184), .B1(n14183), .B2(n9779), .ZN(
        P1_U3474) );
  NOR2_X1 U17353 ( .A1(n14186), .A2(n16063), .ZN(n14190) );
  NAND2_X1 U17354 ( .A1(n16001), .A2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n14187) );
  OAI211_X1 U17355 ( .C1(n15932), .C2(n16072), .A(n14188), .B(n14187), .ZN(
        n14189) );
  AOI211_X2 U17356 ( .C1(n14191), .C2(n16068), .A(n14190), .B(n14189), .ZN(
        n14192) );
  OAI21_X1 U17357 ( .B1(n14193), .B2(n19088), .A(n14192), .ZN(P2_U2983) );
  NOR2_X1 U17358 ( .A1(n14809), .A2(n15938), .ZN(n14194) );
  AOI21_X1 U17359 ( .B1(P2_EBX_REG_30__SCAN_IN), .B2(n15938), .A(n14194), .ZN(
        n14195) );
  OAI21_X1 U17360 ( .B1(n14196), .B2(n18952), .A(n14195), .ZN(P2_U2857) );
  INV_X1 U17361 ( .A(n14450), .ZN(n14370) );
  OAI22_X1 U17362 ( .A1(n14209), .A2(n14200), .B1(n9679), .B2(n14199), .ZN(
        n14202) );
  XNOR2_X1 U17363 ( .A(n14202), .B(n14201), .ZN(n15389) );
  OAI21_X1 U17364 ( .B1(P1_REIP_REG_30__SCAN_IN), .B2(n14204), .A(n14203), 
        .ZN(n14206) );
  AOI22_X1 U17365 ( .A1(n19935), .A2(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .B1(
        P1_EBX_REG_30__SCAN_IN), .B2(n19929), .ZN(n14205) );
  OAI211_X1 U17366 ( .C1(n14451), .C2(n19897), .A(n14206), .B(n14205), .ZN(
        n14207) );
  AOI21_X1 U17367 ( .B1(n15389), .B2(n19905), .A(n14207), .ZN(n14208) );
  OAI21_X1 U17368 ( .B1(n14370), .B2(n19861), .A(n14208), .ZN(P1_U2810) );
  AOI21_X1 U17369 ( .B1(n9679), .B2(n14210), .A(n14209), .ZN(n15667) );
  INV_X1 U17370 ( .A(P1_EBX_REG_29__SCAN_IN), .ZN(n14310) );
  NAND2_X1 U17371 ( .A1(n19935), .A2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n14213) );
  NAND3_X1 U17372 ( .A1(n19920), .A2(n14217), .A3(n14211), .ZN(n14212) );
  OAI211_X1 U17373 ( .C1(n14310), .C2(n19867), .A(n14213), .B(n14212), .ZN(
        n14214) );
  AOI21_X1 U17374 ( .B1(n19934), .B2(n14215), .A(n14214), .ZN(n14216) );
  OAI21_X1 U17375 ( .B1(n15456), .B2(n14217), .A(n14216), .ZN(n14218) );
  AOI21_X1 U17376 ( .B1(n15667), .B2(n19905), .A(n14218), .ZN(n14219) );
  OAI21_X1 U17377 ( .B1(n14373), .B2(n19861), .A(n14219), .ZN(P1_U2811) );
  INV_X1 U17378 ( .A(n14220), .ZN(n14221) );
  AND2_X1 U17379 ( .A1(n14225), .A2(n14224), .ZN(n14226) );
  OR2_X1 U17380 ( .A1(n14226), .A2(n14314), .ZN(n15686) );
  NOR2_X1 U17381 ( .A1(n15686), .A2(n19931), .ZN(n14236) );
  INV_X1 U17382 ( .A(n14227), .ZN(n14229) );
  NOR3_X1 U17383 ( .A1(P1_REIP_REG_27__SCAN_IN), .A2(n19875), .A3(n14229), 
        .ZN(n14235) );
  AOI21_X1 U17384 ( .B1(n19920), .B2(n14229), .A(n14228), .ZN(n15460) );
  INV_X1 U17385 ( .A(P1_REIP_REG_27__SCAN_IN), .ZN(n14230) );
  INV_X1 U17386 ( .A(P1_EBX_REG_27__SCAN_IN), .ZN(n14319) );
  OAI22_X1 U17387 ( .A1(n15460), .A2(n14230), .B1(n14319), .B2(n19867), .ZN(
        n14234) );
  INV_X1 U17388 ( .A(n14231), .ZN(n14463) );
  OAI22_X1 U17389 ( .A1(n14463), .A2(n19897), .B1(n19923), .B2(n14232), .ZN(
        n14233) );
  NOR4_X1 U17390 ( .A1(n14236), .A2(n14235), .A3(n14234), .A4(n14233), .ZN(
        n14237) );
  OAI21_X1 U17391 ( .B1(n14381), .B2(n19861), .A(n14237), .ZN(P1_U2813) );
  AND2_X1 U17392 ( .A1(n9723), .A2(n14238), .ZN(n14239) );
  OR2_X1 U17393 ( .A1(n14239), .A2(n14336), .ZN(n15727) );
  INV_X1 U17394 ( .A(n14242), .ZN(n14340) );
  AOI21_X1 U17395 ( .B1(n14243), .B2(n14240), .A(n14242), .ZN(n15587) );
  NAND2_X1 U17396 ( .A1(n15587), .A2(n19872), .ZN(n14251) );
  INV_X1 U17397 ( .A(P1_REIP_REG_21__SCAN_IN), .ZN(n20650) );
  NAND2_X1 U17398 ( .A1(P1_REIP_REG_19__SCAN_IN), .A2(P1_REIP_REG_18__SCAN_IN), 
        .ZN(n14244) );
  INV_X1 U17399 ( .A(P1_REIP_REG_16__SCAN_IN), .ZN(n20643) );
  NAND3_X1 U17400 ( .A1(n19920), .A2(n14285), .A3(P1_REIP_REG_15__SCAN_IN), 
        .ZN(n15528) );
  NOR2_X1 U17401 ( .A1(n20643), .A2(n15528), .ZN(n14273) );
  NAND2_X1 U17402 ( .A1(P1_REIP_REG_17__SCAN_IN), .A2(n14273), .ZN(n14261) );
  NOR2_X1 U17403 ( .A1(n14244), .A2(n14261), .ZN(n15507) );
  NAND2_X1 U17404 ( .A1(P1_REIP_REG_20__SCAN_IN), .A2(n15507), .ZN(n15498) );
  NOR2_X1 U17405 ( .A1(n20650), .A2(n15498), .ZN(n15488) );
  INV_X1 U17406 ( .A(P1_REIP_REG_22__SCAN_IN), .ZN(n20653) );
  INV_X1 U17407 ( .A(n14245), .ZN(n14246) );
  NAND2_X1 U17408 ( .A1(n14246), .A2(n15472), .ZN(n14260) );
  OAI21_X1 U17409 ( .B1(n14247), .B2(n14260), .A(n19930), .ZN(n15510) );
  OAI21_X1 U17410 ( .B1(P1_REIP_REG_21__SCAN_IN), .B2(n15471), .A(n15510), 
        .ZN(n15503) );
  AOI22_X1 U17411 ( .A1(n19935), .A2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .B1(
        n19929), .B2(P1_EBX_REG_22__SCAN_IN), .ZN(n14248) );
  OAI21_X1 U17412 ( .B1(n15590), .B2(n19897), .A(n14248), .ZN(n14249) );
  AOI221_X1 U17413 ( .B1(n15488), .B2(n20653), .C1(n15503), .C2(
        P1_REIP_REG_22__SCAN_IN), .A(n14249), .ZN(n14250) );
  OAI211_X1 U17414 ( .C1(n19931), .C2(n15727), .A(n14251), .B(n14250), .ZN(
        P1_U2818) );
  INV_X1 U17415 ( .A(n14253), .ZN(n14254) );
  OAI21_X1 U17416 ( .B1(n14255), .B2(n14252), .A(n14254), .ZN(n14498) );
  INV_X1 U17417 ( .A(n14498), .ZN(n14269) );
  INV_X1 U17418 ( .A(P1_REIP_REG_18__SCAN_IN), .ZN(n20646) );
  NOR3_X1 U17419 ( .A1(P1_REIP_REG_19__SCAN_IN), .A2(n20646), .A3(n14261), 
        .ZN(n14268) );
  INV_X1 U17420 ( .A(n14362), .ZN(n14256) );
  NAND2_X1 U17421 ( .A1(n14363), .A2(n14256), .ZN(n14258) );
  NAND2_X1 U17422 ( .A1(n14258), .A2(n14257), .ZN(n14259) );
  NAND2_X1 U17423 ( .A1(n14259), .A2(n14353), .ZN(n15736) );
  OR2_X1 U17424 ( .A1(n15736), .A2(n19931), .ZN(n14266) );
  AND2_X1 U17425 ( .A1(n19930), .A2(n14260), .ZN(n15516) );
  NOR2_X1 U17426 ( .A1(P1_REIP_REG_18__SCAN_IN), .A2(n14261), .ZN(n15522) );
  OAI21_X1 U17427 ( .B1(n15516), .B2(n15522), .A(P1_REIP_REG_19__SCAN_IN), 
        .ZN(n14262) );
  OAI21_X1 U17428 ( .B1(n19867), .B2(n14355), .A(n14262), .ZN(n14263) );
  INV_X1 U17429 ( .A(n14263), .ZN(n14265) );
  AOI22_X1 U17430 ( .A1(n19935), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .B1(
        n19934), .B2(n14494), .ZN(n14264) );
  NAND4_X1 U17431 ( .A1(n14266), .A2(n14265), .A3(n14264), .A4(n19879), .ZN(
        n14267) );
  AOI211_X1 U17432 ( .C1(n14269), .C2(n19872), .A(n14268), .B(n14267), .ZN(
        n14270) );
  INV_X1 U17433 ( .A(n14270), .ZN(P1_U2821) );
  OR2_X1 U17434 ( .A1(n14114), .A2(n14435), .ZN(n14433) );
  AOI21_X1 U17435 ( .B1(n14272), .B2(n14433), .A(n14271), .ZN(n14510) );
  OAI21_X1 U17436 ( .B1(P1_REIP_REG_17__SCAN_IN), .B2(n14273), .A(n15516), 
        .ZN(n14282) );
  INV_X1 U17437 ( .A(n15530), .ZN(n14276) );
  INV_X1 U17438 ( .A(n14274), .ZN(n14275) );
  AOI21_X1 U17439 ( .B1(n15531), .B2(n14276), .A(n14275), .ZN(n14277) );
  OR2_X1 U17440 ( .A1(n14363), .A2(n14277), .ZN(n14365) );
  OAI22_X1 U17441 ( .A1(n14365), .A2(n19931), .B1(n20870), .B2(n19867), .ZN(
        n14278) );
  INV_X1 U17442 ( .A(n14278), .ZN(n14281) );
  INV_X1 U17443 ( .A(n14508), .ZN(n14279) );
  AOI22_X1 U17444 ( .A1(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .A2(n19935), .B1(
        n19934), .B2(n14279), .ZN(n14280) );
  NAND4_X1 U17445 ( .A1(n14282), .A2(n14281), .A3(n14280), .A4(n19879), .ZN(
        n14283) );
  AOI21_X1 U17446 ( .B1(n14510), .B2(n19872), .A(n14283), .ZN(n14284) );
  INV_X1 U17447 ( .A(n14284), .ZN(P1_U2823) );
  AOI21_X1 U17448 ( .B1(P1_REIP_REG_15__SCAN_IN), .B2(n15472), .A(n15471), 
        .ZN(n15526) );
  INV_X1 U17449 ( .A(n15526), .ZN(n14287) );
  AOI21_X1 U17450 ( .B1(n14285), .B2(n19920), .A(P1_REIP_REG_15__SCAN_IN), 
        .ZN(n14286) );
  NOR2_X1 U17451 ( .A1(n14287), .A2(n14286), .ZN(n14294) );
  OAI22_X1 U17452 ( .A1(n14289), .A2(n19931), .B1(n14288), .B2(n19867), .ZN(
        n14293) );
  INV_X1 U17453 ( .A(n14525), .ZN(n14291) );
  OAI22_X1 U17454 ( .A1(n14291), .A2(n19897), .B1(n19923), .B2(n14290), .ZN(
        n14292) );
  NOR4_X1 U17455 ( .A1(n14294), .A2(n19891), .A3(n14293), .A4(n14292), .ZN(
        n14295) );
  OAI21_X1 U17456 ( .B1(n14528), .B2(n19861), .A(n14295), .ZN(P1_U2825) );
  NOR2_X1 U17457 ( .A1(n15343), .A2(n14296), .ZN(n14297) );
  NOR2_X1 U17458 ( .A1(n19872), .A2(n14297), .ZN(n19938) );
  NAND2_X1 U17459 ( .A1(n19920), .A2(P1_REIP_REG_1__SCAN_IN), .ZN(n19907) );
  NOR2_X1 U17460 ( .A1(P1_REIP_REG_2__SCAN_IN), .A2(n19907), .ZN(n19915) );
  INV_X1 U17461 ( .A(n19915), .ZN(n14307) );
  OAI21_X1 U17462 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(n19875), .A(n19922), .ZN(
        n19914) );
  INV_X1 U17463 ( .A(n14298), .ZN(n14300) );
  NAND2_X1 U17464 ( .A1(n14300), .A2(n14299), .ZN(n19932) );
  AOI22_X1 U17465 ( .A1(n20055), .A2(n19905), .B1(n19929), .B2(
        P1_EBX_REG_2__SCAN_IN), .ZN(n14301) );
  OAI21_X1 U17466 ( .B1(n13312), .B2(n19932), .A(n14301), .ZN(n14305) );
  INV_X1 U17467 ( .A(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n14302) );
  OAI22_X1 U17468 ( .A1(n14303), .A2(n19897), .B1(n19923), .B2(n14302), .ZN(
        n14304) );
  AOI211_X1 U17469 ( .C1(P1_REIP_REG_2__SCAN_IN), .C2(n19914), .A(n14305), .B(
        n14304), .ZN(n14306) );
  OAI211_X1 U17470 ( .C1(n19938), .C2(n14308), .A(n14307), .B(n14306), .ZN(
        P1_U2838) );
  OAI22_X1 U17471 ( .A1(n14549), .A2(n14356), .B1(n20794), .B2(n19945), .ZN(
        P1_U2841) );
  AOI22_X1 U17472 ( .A1(n15389), .A2(n19940), .B1(P1_EBX_REG_30__SCAN_IN), 
        .B2(n10965), .ZN(n14309) );
  OAI21_X1 U17473 ( .B1(n14370), .B2(n9630), .A(n14309), .ZN(P1_U2842) );
  INV_X1 U17474 ( .A(n15667), .ZN(n14311) );
  OAI222_X1 U17475 ( .A1(n14311), .A2(n14356), .B1(n19945), .B2(n14310), .C1(
        n9630), .C2(n14373), .ZN(P1_U2843) );
  INV_X1 U17476 ( .A(n15563), .ZN(n14376) );
  OR2_X1 U17477 ( .A1(n14314), .A2(n14313), .ZN(n14315) );
  NAND2_X1 U17478 ( .A1(n9679), .A2(n14315), .ZN(n15680) );
  OAI22_X1 U17479 ( .A1(n15680), .A2(n14356), .B1(n14316), .B2(n19945), .ZN(
        n14317) );
  INV_X1 U17480 ( .A(n14317), .ZN(n14318) );
  OAI21_X1 U17481 ( .B1(n14376), .B2(n9630), .A(n14318), .ZN(P1_U2844) );
  OAI222_X1 U17482 ( .A1(n15686), .A2(n14356), .B1(n19945), .B2(n14319), .C1(
        n9630), .C2(n14381), .ZN(P1_U2845) );
  NAND2_X1 U17483 ( .A1(n14331), .A2(n14320), .ZN(n14321) );
  NAND2_X1 U17484 ( .A1(n14322), .A2(n14321), .ZN(n15700) );
  INV_X1 U17485 ( .A(P1_EBX_REG_25__SCAN_IN), .ZN(n14325) );
  OAI222_X1 U17486 ( .A1(n15700), .A2(n14356), .B1(n19945), .B2(n14325), .C1(
        n9630), .C2(n15468), .ZN(P1_U2847) );
  NOR2_X1 U17487 ( .A1(n14326), .A2(n14327), .ZN(n14328) );
  OR2_X1 U17488 ( .A1(n14323), .A2(n14328), .ZN(n15479) );
  OR2_X1 U17489 ( .A1(n14338), .A2(n14329), .ZN(n14330) );
  NAND2_X1 U17490 ( .A1(n14331), .A2(n14330), .ZN(n15709) );
  OAI22_X1 U17491 ( .A1(n15709), .A2(n14356), .B1(n14332), .B2(n19945), .ZN(
        n14333) );
  INV_X1 U17492 ( .A(n14333), .ZN(n14334) );
  OAI21_X1 U17493 ( .B1(n15479), .B2(n9630), .A(n14334), .ZN(P1_U2848) );
  NOR2_X1 U17494 ( .A1(n14336), .A2(n14335), .ZN(n14337) );
  OR2_X1 U17495 ( .A1(n14338), .A2(n14337), .ZN(n15712) );
  INV_X1 U17496 ( .A(P1_EBX_REG_23__SCAN_IN), .ZN(n14342) );
  AND2_X1 U17497 ( .A1(n14340), .A2(n14339), .ZN(n14341) );
  OR2_X1 U17498 ( .A1(n14341), .A2(n14326), .ZN(n14480) );
  OAI222_X1 U17499 ( .A1(n15712), .A2(n14356), .B1(n14342), .B2(n19945), .C1(
        n14480), .C2(n9630), .ZN(P1_U2849) );
  INV_X1 U17500 ( .A(n15587), .ZN(n14406) );
  OAI222_X1 U17501 ( .A1(n15727), .A2(n14356), .B1(n14343), .B2(n19945), .C1(
        n14406), .C2(n9630), .ZN(P1_U2850) );
  INV_X1 U17502 ( .A(n14352), .ZN(n14345) );
  OAI21_X1 U17503 ( .B1(n14353), .B2(n14345), .A(n14344), .ZN(n14346) );
  AND2_X1 U17504 ( .A1(n14346), .A2(n9723), .ZN(n15381) );
  INV_X1 U17505 ( .A(n15381), .ZN(n15499) );
  INV_X1 U17506 ( .A(P1_EBX_REG_21__SCAN_IN), .ZN(n14349) );
  OAI21_X1 U17507 ( .B1(n14347), .B2(n14348), .A(n14240), .ZN(n15500) );
  OAI222_X1 U17508 ( .A1(n15499), .A2(n14356), .B1(n19945), .B2(n14349), .C1(
        n9630), .C2(n15500), .ZN(P1_U2851) );
  NOR2_X1 U17509 ( .A1(n14253), .A2(n14350), .ZN(n14351) );
  OR2_X1 U17510 ( .A1(n14347), .A2(n14351), .ZN(n15592) );
  XNOR2_X1 U17511 ( .A(n14353), .B(n14352), .ZN(n15508) );
  AOI22_X1 U17512 ( .A1(n15508), .A2(n19940), .B1(n10965), .B2(
        P1_EBX_REG_20__SCAN_IN), .ZN(n14354) );
  OAI21_X1 U17513 ( .B1(n15592), .B2(n9630), .A(n14354), .ZN(P1_U2852) );
  OAI22_X1 U17514 ( .A1(n15736), .A2(n14356), .B1(n14355), .B2(n19945), .ZN(
        n14357) );
  INV_X1 U17515 ( .A(n14357), .ZN(n14358) );
  OAI21_X1 U17516 ( .B1(n14498), .B2(n9630), .A(n14358), .ZN(P1_U2853) );
  AND2_X1 U17517 ( .A1(n14360), .A2(n14359), .ZN(n14361) );
  OR2_X1 U17518 ( .A1(n14361), .A2(n14252), .ZN(n15601) );
  XNOR2_X1 U17519 ( .A(n14363), .B(n14362), .ZN(n15741) );
  AOI22_X1 U17520 ( .A1(n15741), .A2(n19940), .B1(n10965), .B2(
        P1_EBX_REG_18__SCAN_IN), .ZN(n14364) );
  OAI21_X1 U17521 ( .B1(n15601), .B2(n9630), .A(n14364), .ZN(P1_U2854) );
  INV_X1 U17522 ( .A(n14510), .ZN(n14432) );
  INV_X1 U17523 ( .A(n14365), .ZN(n15751) );
  AOI22_X1 U17524 ( .A1(n15751), .A2(n19940), .B1(n10965), .B2(
        P1_EBX_REG_17__SCAN_IN), .ZN(n14366) );
  OAI21_X1 U17525 ( .B1(n14432), .B2(n9630), .A(n14366), .ZN(P1_U2855) );
  AOI22_X1 U17526 ( .A1(n14422), .A2(BUF1_REG_30__SCAN_IN), .B1(
        P1_EAX_REG_30__SCAN_IN), .B2(n14421), .ZN(n14369) );
  NOR3_X4 U17527 ( .A1(n14421), .A2(n20117), .A3(n14367), .ZN(n14441) );
  AOI22_X1 U17528 ( .A1(n20011), .A2(n14441), .B1(n14439), .B2(DATAI_30_), 
        .ZN(n14368) );
  OAI211_X1 U17529 ( .C1(n14370), .C2(n14396), .A(n14369), .B(n14368), .ZN(
        P1_U2874) );
  AOI22_X1 U17530 ( .A1(n14422), .A2(BUF1_REG_29__SCAN_IN), .B1(
        P1_EAX_REG_29__SCAN_IN), .B2(n14421), .ZN(n14372) );
  AOI22_X1 U17531 ( .A1(n14441), .A2(n20009), .B1(n14439), .B2(DATAI_29_), 
        .ZN(n14371) );
  OAI211_X1 U17532 ( .C1(n14373), .C2(n14396), .A(n14372), .B(n14371), .ZN(
        P1_U2875) );
  AOI22_X1 U17533 ( .A1(n14422), .A2(BUF1_REG_28__SCAN_IN), .B1(
        P1_EAX_REG_28__SCAN_IN), .B2(n14421), .ZN(n14375) );
  AOI22_X1 U17534 ( .A1(n14441), .A2(n20007), .B1(n14439), .B2(DATAI_28_), 
        .ZN(n14374) );
  OAI211_X1 U17535 ( .C1(n14376), .C2(n14396), .A(n14375), .B(n14374), .ZN(
        P1_U2876) );
  OAI22_X1 U17536 ( .A1(n14437), .A2(n16255), .B1(n14377), .B2(n14436), .ZN(
        n14378) );
  INV_X1 U17537 ( .A(n14378), .ZN(n14380) );
  AOI22_X1 U17538 ( .A1(n14441), .A2(n20005), .B1(n14439), .B2(DATAI_27_), 
        .ZN(n14379) );
  OAI211_X1 U17539 ( .C1(n14381), .C2(n14396), .A(n14380), .B(n14379), .ZN(
        P1_U2877) );
  INV_X1 U17540 ( .A(n15572), .ZN(n14386) );
  OAI22_X1 U17541 ( .A1(n14437), .A2(n16257), .B1(n14382), .B2(n14436), .ZN(
        n14383) );
  INV_X1 U17542 ( .A(n14383), .ZN(n14385) );
  AOI22_X1 U17543 ( .A1(n14441), .A2(n20003), .B1(n14439), .B2(DATAI_26_), 
        .ZN(n14384) );
  OAI211_X1 U17544 ( .C1(n14386), .C2(n14396), .A(n14385), .B(n14384), .ZN(
        P1_U2878) );
  INV_X1 U17545 ( .A(BUF1_REG_25__SCAN_IN), .ZN(n14388) );
  OAI22_X1 U17546 ( .A1(n14437), .A2(n14388), .B1(n14387), .B2(n14436), .ZN(
        n14389) );
  INV_X1 U17547 ( .A(n14389), .ZN(n14391) );
  AOI22_X1 U17548 ( .A1(n14441), .A2(n20001), .B1(n14439), .B2(DATAI_25_), 
        .ZN(n14390) );
  OAI211_X1 U17549 ( .C1(n15468), .C2(n14396), .A(n14391), .B(n14390), .ZN(
        P1_U2879) );
  INV_X1 U17550 ( .A(BUF1_REG_24__SCAN_IN), .ZN(n14392) );
  INV_X1 U17551 ( .A(P1_EAX_REG_24__SCAN_IN), .ZN(n19957) );
  OAI22_X1 U17552 ( .A1(n14437), .A2(n14392), .B1(n19957), .B2(n14436), .ZN(
        n14393) );
  INV_X1 U17553 ( .A(n14393), .ZN(n14395) );
  AOI22_X1 U17554 ( .A1(n14441), .A2(n19997), .B1(n14439), .B2(DATAI_24_), 
        .ZN(n14394) );
  OAI211_X1 U17555 ( .C1(n15479), .C2(n14396), .A(n14395), .B(n14394), .ZN(
        P1_U2880) );
  OAI22_X1 U17556 ( .A1(n14437), .A2(n16261), .B1(n14397), .B2(n14436), .ZN(
        n14398) );
  INV_X1 U17557 ( .A(n14398), .ZN(n14401) );
  AOI22_X1 U17558 ( .A1(n14441), .A2(n14399), .B1(n14439), .B2(DATAI_23_), 
        .ZN(n14400) );
  OAI211_X1 U17559 ( .C1(n14480), .C2(n14396), .A(n14401), .B(n14400), .ZN(
        P1_U2881) );
  INV_X1 U17560 ( .A(BUF1_REG_22__SCAN_IN), .ZN(n16263) );
  INV_X1 U17561 ( .A(P1_EAX_REG_22__SCAN_IN), .ZN(n19960) );
  OAI22_X1 U17562 ( .A1(n14437), .A2(n16263), .B1(n19960), .B2(n14436), .ZN(
        n14402) );
  INV_X1 U17563 ( .A(n14402), .ZN(n14405) );
  AOI22_X1 U17564 ( .A1(n14441), .A2(n14403), .B1(n14439), .B2(DATAI_22_), 
        .ZN(n14404) );
  OAI211_X1 U17565 ( .C1(n14406), .C2(n14396), .A(n14405), .B(n14404), .ZN(
        P1_U2882) );
  AOI22_X1 U17566 ( .A1(n14422), .A2(BUF1_REG_21__SCAN_IN), .B1(
        P1_EAX_REG_21__SCAN_IN), .B2(n14421), .ZN(n14409) );
  AOI22_X1 U17567 ( .A1(n14441), .A2(n14407), .B1(n14439), .B2(DATAI_21_), 
        .ZN(n14408) );
  OAI211_X1 U17568 ( .C1(n15500), .C2(n14396), .A(n14409), .B(n14408), .ZN(
        P1_U2883) );
  INV_X1 U17569 ( .A(BUF1_REG_20__SCAN_IN), .ZN(n14410) );
  OAI22_X1 U17570 ( .A1(n14437), .A2(n14410), .B1(n19964), .B2(n14436), .ZN(
        n14411) );
  INV_X1 U17571 ( .A(n14411), .ZN(n14414) );
  AOI22_X1 U17572 ( .A1(n14441), .A2(n14412), .B1(n14439), .B2(DATAI_20_), 
        .ZN(n14413) );
  OAI211_X1 U17573 ( .C1(n15592), .C2(n14396), .A(n14414), .B(n14413), .ZN(
        P1_U2884) );
  INV_X1 U17574 ( .A(BUF1_REG_19__SCAN_IN), .ZN(n14416) );
  OAI22_X1 U17575 ( .A1(n14437), .A2(n14416), .B1(n14415), .B2(n14436), .ZN(
        n14417) );
  INV_X1 U17576 ( .A(n14417), .ZN(n14420) );
  AOI22_X1 U17577 ( .A1(n14441), .A2(n14418), .B1(n14439), .B2(DATAI_19_), 
        .ZN(n14419) );
  OAI211_X1 U17578 ( .C1(n14498), .C2(n14396), .A(n14420), .B(n14419), .ZN(
        P1_U2885) );
  AOI22_X1 U17579 ( .A1(n14422), .A2(BUF1_REG_18__SCAN_IN), .B1(
        P1_EAX_REG_18__SCAN_IN), .B2(n14421), .ZN(n14425) );
  AOI22_X1 U17580 ( .A1(n14441), .A2(n14423), .B1(n14439), .B2(DATAI_18_), 
        .ZN(n14424) );
  OAI211_X1 U17581 ( .C1(n15601), .C2(n14396), .A(n14425), .B(n14424), .ZN(
        P1_U2886) );
  INV_X1 U17582 ( .A(BUF1_REG_17__SCAN_IN), .ZN(n14427) );
  OAI22_X1 U17583 ( .A1(n14437), .A2(n14427), .B1(n14426), .B2(n14436), .ZN(
        n14428) );
  INV_X1 U17584 ( .A(n14428), .ZN(n14431) );
  AOI22_X1 U17585 ( .A1(n14441), .A2(n14429), .B1(n14439), .B2(DATAI_17_), 
        .ZN(n14430) );
  OAI211_X1 U17586 ( .C1(n14432), .C2(n14396), .A(n14431), .B(n14430), .ZN(
        P1_U2887) );
  INV_X1 U17587 ( .A(n14433), .ZN(n14434) );
  AOI21_X1 U17588 ( .B1(n14435), .B2(n14114), .A(n14434), .ZN(n15612) );
  INV_X1 U17589 ( .A(n15612), .ZN(n14444) );
  OAI22_X1 U17590 ( .A1(n14437), .A2(n20909), .B1(n19974), .B2(n14436), .ZN(
        n14438) );
  INV_X1 U17591 ( .A(n14438), .ZN(n14443) );
  AOI22_X1 U17592 ( .A1(n14441), .A2(n14440), .B1(n14439), .B2(DATAI_16_), 
        .ZN(n14442) );
  OAI211_X1 U17593 ( .C1(n14444), .C2(n14396), .A(n14443), .B(n14442), .ZN(
        P1_U2888) );
  NOR2_X1 U17594 ( .A1(n14446), .A2(n14445), .ZN(n14448) );
  XNOR2_X1 U17595 ( .A(n14449), .B(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n15392) );
  NAND2_X1 U17596 ( .A1(n14450), .A2(n15645), .ZN(n14457) );
  INV_X1 U17597 ( .A(n14451), .ZN(n14455) );
  INV_X1 U17598 ( .A(P1_REIP_REG_30__SCAN_IN), .ZN(n14452) );
  OR2_X1 U17599 ( .A1(n20050), .A2(n14452), .ZN(n15390) );
  OAI21_X1 U17600 ( .B1(n20039), .B2(n14453), .A(n15390), .ZN(n14454) );
  AOI21_X1 U17601 ( .B1(n14455), .B2(n15635), .A(n14454), .ZN(n14456) );
  OAI211_X1 U17602 ( .C1(n15392), .C2(n20031), .A(n14457), .B(n14456), .ZN(
        P1_U2969) );
  INV_X1 U17603 ( .A(n14458), .ZN(n15570) );
  NAND2_X1 U17604 ( .A1(n15570), .A2(n15559), .ZN(n14459) );
  AOI22_X1 U17605 ( .A1(n20034), .A2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .B1(
        n20043), .B2(P1_REIP_REG_27__SCAN_IN), .ZN(n14462) );
  OAI21_X1 U17606 ( .B1(n20032), .B2(n14463), .A(n14462), .ZN(n14464) );
  AOI21_X1 U17607 ( .B1(n14465), .B2(n15645), .A(n14464), .ZN(n14466) );
  OAI21_X1 U17608 ( .B1(n14467), .B2(n20031), .A(n14466), .ZN(P1_U2972) );
  MUX2_X1 U17609 ( .A(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .B(n15640), .S(
        P1_INSTADDRPOINTER_REG_23__SCAN_IN), .Z(n14470) );
  INV_X1 U17610 ( .A(n15568), .ZN(n14469) );
  AOI211_X1 U17611 ( .C1(n15577), .C2(n14468), .A(n14470), .B(n14469), .ZN(
        n14472) );
  XNOR2_X1 U17612 ( .A(n14472), .B(n14471), .ZN(n15696) );
  AOI22_X1 U17613 ( .A1(n20042), .A2(n15696), .B1(n20043), .B2(
        P1_REIP_REG_25__SCAN_IN), .ZN(n14473) );
  OAI21_X1 U17614 ( .B1(n20039), .B2(n10802), .A(n14473), .ZN(n14474) );
  AOI21_X1 U17615 ( .B1(n15635), .B2(n15470), .A(n14474), .ZN(n14475) );
  OAI21_X1 U17616 ( .B1(n15468), .B2(n20084), .A(n14475), .ZN(P1_U2974) );
  NOR2_X1 U17617 ( .A1(n15640), .A2(n15717), .ZN(n14478) );
  MUX2_X1 U17618 ( .A(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .B(n15717), .S(
        n15569), .Z(n14477) );
  MUX2_X1 U17619 ( .A(n14478), .B(n14477), .S(n14468), .Z(n14479) );
  AOI21_X1 U17620 ( .B1(n14476), .B2(n15640), .A(n14479), .ZN(n15711) );
  INV_X1 U17621 ( .A(n14480), .ZN(n15493) );
  INV_X1 U17622 ( .A(n15487), .ZN(n14482) );
  AOI22_X1 U17623 ( .A1(n20034), .A2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .B1(
        n20043), .B2(P1_REIP_REG_23__SCAN_IN), .ZN(n14481) );
  OAI21_X1 U17624 ( .B1(n20032), .B2(n14482), .A(n14481), .ZN(n14483) );
  AOI21_X1 U17625 ( .B1(n15493), .B2(n15645), .A(n14483), .ZN(n14484) );
  OAI21_X1 U17626 ( .B1(n15711), .B2(n20031), .A(n14484), .ZN(P1_U2976) );
  OAI22_X1 U17627 ( .A1(n20039), .A2(n15506), .B1(n20050), .B2(n20650), .ZN(
        n14485) );
  AOI21_X1 U17628 ( .B1(n15635), .B2(n15497), .A(n14485), .ZN(n14491) );
  INV_X1 U17629 ( .A(n14486), .ZN(n14487) );
  NAND3_X1 U17630 ( .A1(n14487), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A3(
        n15569), .ZN(n15415) );
  OAI22_X1 U17631 ( .A1(n15415), .A2(n15419), .B1(n15569), .B2(n14488), .ZN(
        n14489) );
  XOR2_X1 U17632 ( .A(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .B(n14489), .Z(
        n15380) );
  NAND2_X1 U17633 ( .A1(n15380), .A2(n20042), .ZN(n14490) );
  OAI211_X1 U17634 ( .C1(n15500), .C2(n20084), .A(n14491), .B(n14490), .ZN(
        P1_U2978) );
  INV_X1 U17635 ( .A(P1_REIP_REG_19__SCAN_IN), .ZN(n14492) );
  OAI22_X1 U17636 ( .A1(n20039), .A2(n10697), .B1(n20050), .B2(n14492), .ZN(
        n14493) );
  AOI21_X1 U17637 ( .B1(n15635), .B2(n14494), .A(n14493), .ZN(n14497) );
  NOR2_X1 U17638 ( .A1(n15569), .A2(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n15414) );
  MUX2_X1 U17639 ( .A(n15569), .B(n15414), .S(n14486), .Z(n14495) );
  XNOR2_X1 U17640 ( .A(n14495), .B(n15413), .ZN(n15733) );
  NAND2_X1 U17641 ( .A1(n15733), .A2(n20042), .ZN(n14496) );
  OAI211_X1 U17642 ( .C1(n14498), .C2(n20084), .A(n14497), .B(n14496), .ZN(
        P1_U2980) );
  NAND3_X1 U17643 ( .A1(n15638), .A2(n14500), .A3(n15615), .ZN(n14502) );
  NAND2_X1 U17644 ( .A1(n14502), .A2(n14501), .ZN(n14503) );
  NAND2_X1 U17645 ( .A1(n15640), .A2(n14503), .ZN(n14504) );
  OAI22_X1 U17646 ( .A1(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n14504), .B1(
        n15640), .B2(n14503), .ZN(n14505) );
  XNOR2_X1 U17647 ( .A(n14506), .B(n14505), .ZN(n15750) );
  INV_X1 U17648 ( .A(n15750), .ZN(n14512) );
  AOI22_X1 U17649 ( .A1(n20034), .A2(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .B1(
        n20043), .B2(P1_REIP_REG_17__SCAN_IN), .ZN(n14507) );
  OAI21_X1 U17650 ( .B1(n20032), .B2(n14508), .A(n14507), .ZN(n14509) );
  AOI21_X1 U17651 ( .B1(n14510), .B2(n15645), .A(n14509), .ZN(n14511) );
  OAI21_X1 U17652 ( .B1(n14512), .B2(n20031), .A(n14511), .ZN(P1_U2982) );
  INV_X1 U17653 ( .A(n14513), .ZN(n14514) );
  OAI21_X1 U17654 ( .B1(n15638), .B2(n14515), .A(n14514), .ZN(n14518) );
  INV_X1 U17655 ( .A(n14516), .ZN(n14519) );
  NOR2_X1 U17656 ( .A1(n14518), .A2(n14519), .ZN(n15607) );
  INV_X1 U17657 ( .A(n15607), .ZN(n14522) );
  INV_X1 U17658 ( .A(n14517), .ZN(n14521) );
  OAI21_X1 U17659 ( .B1(n14519), .B2(n14521), .A(n14518), .ZN(n14520) );
  OAI21_X1 U17660 ( .B1(n14522), .B2(n14521), .A(n14520), .ZN(n15765) );
  NAND2_X1 U17661 ( .A1(n15765), .A2(n20042), .ZN(n14527) );
  INV_X1 U17662 ( .A(P1_REIP_REG_15__SCAN_IN), .ZN(n14523) );
  OAI22_X1 U17663 ( .A1(n20039), .A2(n14290), .B1(n20050), .B2(n14523), .ZN(
        n14524) );
  AOI21_X1 U17664 ( .B1(n15635), .B2(n14525), .A(n14524), .ZN(n14526) );
  OAI211_X1 U17665 ( .C1(n20084), .C2(n14528), .A(n14527), .B(n14526), .ZN(
        P1_U2984) );
  INV_X1 U17666 ( .A(n14529), .ZN(n14530) );
  AOI21_X1 U17667 ( .B1(n14499), .B2(n9714), .A(n14530), .ZN(n15630) );
  INV_X1 U17668 ( .A(n14533), .ZN(n14532) );
  AND2_X1 U17669 ( .A1(n14532), .A2(n14531), .ZN(n15629) );
  AND2_X1 U17670 ( .A1(n15630), .A2(n15629), .ZN(n15632) );
  NOR2_X1 U17671 ( .A1(n15632), .A2(n14533), .ZN(n14535) );
  XNOR2_X1 U17672 ( .A(n14535), .B(n14534), .ZN(n15789) );
  INV_X1 U17673 ( .A(n15789), .ZN(n14541) );
  AOI22_X1 U17674 ( .A1(n20034), .A2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .B1(
        n20043), .B2(P1_REIP_REG_13__SCAN_IN), .ZN(n14536) );
  OAI21_X1 U17675 ( .B1(n20032), .B2(n14537), .A(n14536), .ZN(n14538) );
  AOI21_X1 U17676 ( .B1(n14539), .B2(n15645), .A(n14538), .ZN(n14540) );
  OAI21_X1 U17677 ( .B1(n14541), .B2(n20031), .A(n14540), .ZN(P1_U2986) );
  MUX2_X1 U17678 ( .A(n15638), .B(n15639), .S(n15640), .Z(n14542) );
  XOR2_X1 U17679 ( .A(n11184), .B(n14542), .Z(n15825) );
  INV_X1 U17680 ( .A(n15825), .ZN(n14548) );
  AOI22_X1 U17681 ( .A1(n20034), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .B1(
        n20043), .B2(P1_REIP_REG_10__SCAN_IN), .ZN(n14543) );
  OAI21_X1 U17682 ( .B1(n20032), .B2(n14544), .A(n14543), .ZN(n14545) );
  AOI21_X1 U17683 ( .B1(n14546), .B2(n15645), .A(n14545), .ZN(n14547) );
  OAI21_X1 U17684 ( .B1(n14548), .B2(n20031), .A(n14547), .ZN(P1_U2989) );
  INV_X1 U17685 ( .A(n14549), .ZN(n14555) );
  NOR2_X1 U17686 ( .A1(n11181), .A2(n11180), .ZN(n15756) );
  NAND2_X1 U17687 ( .A1(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n15756), .ZN(
        n15743) );
  NOR3_X1 U17688 ( .A1(n15749), .A2(n15778), .A3(n15743), .ZN(n14557) );
  NAND3_X1 U17689 ( .A1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n15820) );
  NOR3_X1 U17690 ( .A1(n11184), .A2(n15833), .A3(n15820), .ZN(n15796) );
  NOR2_X1 U17691 ( .A1(n20048), .A2(n14550), .ZN(n15818) );
  NAND3_X1 U17692 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n15796), .A3(
        n15818), .ZN(n15797) );
  NOR2_X1 U17693 ( .A1(n15803), .A2(n15797), .ZN(n15770) );
  NAND2_X1 U17694 ( .A1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n15770), .ZN(
        n15737) );
  NOR3_X1 U17695 ( .A1(n11122), .A2(n10874), .A3(n14550), .ZN(n15817) );
  AND2_X1 U17696 ( .A1(n15817), .A2(n15796), .ZN(n15800) );
  NAND3_X1 U17697 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A3(n15800), .ZN(n14556) );
  NOR2_X1 U17698 ( .A1(n15793), .A2(n14556), .ZN(n15783) );
  NAND2_X1 U17699 ( .A1(n15802), .A2(n15783), .ZN(n15704) );
  OAI21_X1 U17700 ( .B1(n15737), .B2(n20066), .A(n15704), .ZN(n15740) );
  NAND4_X1 U17701 ( .A1(n14551), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .A3(
        n14557), .A4(n15740), .ZN(n15701) );
  INV_X1 U17702 ( .A(n15701), .ZN(n15710) );
  AND2_X1 U17703 ( .A1(n14552), .A2(n15710), .ZN(n15691) );
  NAND2_X1 U17704 ( .A1(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n15691), .ZN(
        n15681) );
  NOR2_X1 U17705 ( .A1(n15673), .A2(n15681), .ZN(n15665) );
  NAND2_X1 U17706 ( .A1(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(n15665), .ZN(
        n15385) );
  INV_X1 U17707 ( .A(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n15386) );
  NOR3_X1 U17708 ( .A1(n15385), .A2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n15386), .ZN(n14553) );
  AOI211_X1 U17709 ( .C1(n20064), .C2(n14555), .A(n14554), .B(n14553), .ZN(
        n14563) );
  INV_X1 U17710 ( .A(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n15559) );
  INV_X1 U17711 ( .A(n15688), .ZN(n14560) );
  NAND2_X1 U17712 ( .A1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n15722) );
  INV_X1 U17713 ( .A(n14556), .ZN(n15788) );
  AND2_X1 U17714 ( .A1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n14557), .ZN(
        n15378) );
  NAND2_X1 U17715 ( .A1(n15788), .A2(n15378), .ZN(n15730) );
  INV_X1 U17716 ( .A(n15737), .ZN(n15779) );
  AOI21_X1 U17717 ( .B1(n14557), .B2(n15779), .A(n20066), .ZN(n14558) );
  AOI211_X1 U17718 ( .C1(n20047), .C2(n15730), .A(n14558), .B(n20046), .ZN(
        n15418) );
  NOR2_X1 U17719 ( .A1(n15834), .A2(n20046), .ZN(n14559) );
  OAI21_X1 U17720 ( .B1(n14560), .B2(n20060), .A(n15703), .ZN(n15697) );
  NAND2_X1 U17721 ( .A1(n15718), .A2(n20060), .ZN(n15676) );
  INV_X1 U17722 ( .A(n15672), .ZN(n14561) );
  OAI211_X1 U17723 ( .C1(n14561), .C2(n15386), .A(
        P1_INSTADDRPOINTER_REG_31__SCAN_IN), .B(n15676), .ZN(n14562) );
  OAI211_X1 U17724 ( .C1(n14564), .C2(n20070), .A(n14563), .B(n14562), .ZN(
        P1_U3000) );
  INV_X1 U17725 ( .A(n15876), .ZN(n14568) );
  NAND2_X1 U17726 ( .A1(n14568), .A2(n14567), .ZN(n14577) );
  INV_X1 U17727 ( .A(P2_EBX_REG_29__SCAN_IN), .ZN(n14570) );
  OAI22_X1 U17728 ( .A1(n18929), .A2(n14570), .B1(n14569), .B2(n18935), .ZN(
        n14575) );
  OAI22_X1 U17729 ( .A1(n14815), .A2(n18928), .B1(n19731), .B2(n18932), .ZN(
        n14574) );
  AOI211_X1 U17730 ( .C1(n14817), .C2(n18916), .A(n14575), .B(n14574), .ZN(
        n14576) );
  OAI211_X1 U17731 ( .C1(n14578), .C2(n18923), .A(n14577), .B(n14576), .ZN(
        P2_U2826) );
  NOR2_X1 U17732 ( .A1(n14580), .A2(n14581), .ZN(n14582) );
  OR2_X1 U17733 ( .A1(n14579), .A2(n14582), .ZN(n15968) );
  OAI21_X1 U17734 ( .B1(n14678), .B2(n14584), .A(n14583), .ZN(n14855) );
  AOI22_X1 U17735 ( .A1(n14585), .A2(n18896), .B1(P2_EBX_REG_25__SCAN_IN), 
        .B2(n18842), .ZN(n14587) );
  AOI22_X1 U17736 ( .A1(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n18892), .B1(
        P2_REIP_REG_25__SCAN_IN), .B2(n18910), .ZN(n14586) );
  OAI211_X1 U17737 ( .C1(n14855), .C2(n18928), .A(n14587), .B(n14586), .ZN(
        n14591) );
  AOI211_X1 U17738 ( .C1(n15962), .C2(n14589), .A(n14588), .B(n18890), .ZN(
        n14590) );
  NOR2_X1 U17739 ( .A1(n14591), .A2(n14590), .ZN(n14592) );
  OAI21_X1 U17740 ( .B1(n18924), .B2(n15968), .A(n14592), .ZN(P2_U2830) );
  INV_X1 U17741 ( .A(n14593), .ZN(n14641) );
  NAND2_X1 U17742 ( .A1(n14595), .A2(n14594), .ZN(n14640) );
  NAND3_X1 U17743 ( .A1(n14641), .A2(n15942), .A3(n14640), .ZN(n14597) );
  NAND2_X1 U17744 ( .A1(n18945), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n14596) );
  OAI211_X1 U17745 ( .C1(n14598), .C2(n18945), .A(n14597), .B(n14596), .ZN(
        P2_U2858) );
  NAND2_X1 U17746 ( .A1(n14600), .A2(n14599), .ZN(n14602) );
  XNOR2_X1 U17747 ( .A(n14602), .B(n14601), .ZN(n14652) );
  NAND2_X1 U17748 ( .A1(n18945), .A2(P2_EBX_REG_28__SCAN_IN), .ZN(n14604) );
  NAND2_X1 U17749 ( .A1(n15892), .A2(n15948), .ZN(n14603) );
  OAI211_X1 U17750 ( .C1(n14652), .C2(n18952), .A(n14604), .B(n14603), .ZN(
        P2_U2859) );
  AOI21_X1 U17751 ( .B1(n14607), .B2(n14606), .A(n9610), .ZN(n14608) );
  INV_X1 U17752 ( .A(n14608), .ZN(n14659) );
  NAND2_X1 U17753 ( .A1(n18945), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n14614) );
  INV_X1 U17754 ( .A(n14610), .ZN(n14611) );
  NAND2_X1 U17755 ( .A1(n15899), .A2(n15948), .ZN(n14613) );
  OAI211_X1 U17756 ( .C1(n14659), .C2(n18952), .A(n14614), .B(n14613), .ZN(
        P2_U2860) );
  OR2_X1 U17757 ( .A1(n14579), .A2(n14615), .ZN(n14616) );
  NAND2_X1 U17758 ( .A1(n14609), .A2(n14616), .ZN(n14843) );
  AOI21_X1 U17759 ( .B1(n14619), .B2(n14618), .A(n14617), .ZN(n14660) );
  NAND2_X1 U17760 ( .A1(n14660), .A2(n15942), .ZN(n14621) );
  NAND2_X1 U17761 ( .A1(n15938), .A2(P2_EBX_REG_26__SCAN_IN), .ZN(n14620) );
  OAI211_X1 U17762 ( .C1(n14843), .C2(n15938), .A(n14621), .B(n14620), .ZN(
        P2_U2861) );
  OAI21_X1 U17763 ( .B1(n9611), .B2(n14623), .A(n9609), .ZN(n14675) );
  NOR2_X1 U17764 ( .A1(n15968), .A2(n15938), .ZN(n14625) );
  AOI21_X1 U17765 ( .B1(P2_EBX_REG_25__SCAN_IN), .B2(n15938), .A(n14625), .ZN(
        n14626) );
  OAI21_X1 U17766 ( .B1(n14675), .B2(n18952), .A(n14626), .ZN(P2_U2862) );
  AOI21_X1 U17767 ( .B1(n9728), .B2(n14628), .A(n14627), .ZN(n14629) );
  XOR2_X1 U17768 ( .A(n14630), .B(n14629), .Z(n14686) );
  AND2_X1 U17769 ( .A1(n14632), .A2(n14631), .ZN(n14633) );
  OR2_X1 U17770 ( .A1(n14633), .A2(n14580), .ZN(n15969) );
  NOR2_X1 U17771 ( .A1(n15969), .A2(n15938), .ZN(n14634) );
  AOI21_X1 U17772 ( .B1(P2_EBX_REG_24__SCAN_IN), .B2(n15938), .A(n14634), .ZN(
        n14635) );
  OAI21_X1 U17773 ( .B1(n14686), .B2(n18952), .A(n14635), .ZN(P2_U2863) );
  XNOR2_X1 U17774 ( .A(n14759), .B(n14636), .ZN(n18742) );
  MUX2_X1 U17775 ( .A(n18742), .B(n14637), .S(n18945), .Z(n14638) );
  OAI21_X1 U17776 ( .B1(n14639), .B2(n18952), .A(n14638), .ZN(P2_U2866) );
  NAND3_X1 U17777 ( .A1(n14641), .A2(n19031), .A3(n14640), .ZN(n14647) );
  INV_X1 U17778 ( .A(n14815), .ZN(n14644) );
  OAI22_X1 U17779 ( .A1(n14691), .A2(n18978), .B1(n14642), .B2(n18995), .ZN(
        n14643) );
  AOI21_X1 U17780 ( .B1(n19027), .B2(n14644), .A(n14643), .ZN(n14646) );
  AOI22_X1 U17781 ( .A1(n18965), .A2(BUF2_REG_29__SCAN_IN), .B1(n18964), .B2(
        BUF1_REG_29__SCAN_IN), .ZN(n14645) );
  NAND3_X1 U17782 ( .A1(n14647), .A2(n14646), .A3(n14645), .ZN(P2_U2890) );
  INV_X1 U17783 ( .A(n14648), .ZN(n15891) );
  OAI22_X1 U17784 ( .A1(n14691), .A2(n18981), .B1(n20839), .B2(n18995), .ZN(
        n14649) );
  AOI21_X1 U17785 ( .B1(n15891), .B2(n19027), .A(n14649), .ZN(n14651) );
  AOI22_X1 U17786 ( .A1(n18965), .A2(BUF2_REG_28__SCAN_IN), .B1(n18964), .B2(
        BUF1_REG_28__SCAN_IN), .ZN(n14650) );
  OAI211_X1 U17787 ( .C1(n14652), .C2(n19002), .A(n14651), .B(n14650), .ZN(
        P2_U2891) );
  AOI21_X1 U17788 ( .B1(n14654), .B2(n14663), .A(n14653), .ZN(n14830) );
  OAI22_X1 U17789 ( .A1(n14691), .A2(n18983), .B1(n14655), .B2(n18995), .ZN(
        n14656) );
  AOI21_X1 U17790 ( .B1(n19027), .B2(n14830), .A(n14656), .ZN(n14658) );
  AOI22_X1 U17791 ( .A1(n18965), .A2(BUF2_REG_27__SCAN_IN), .B1(n18964), .B2(
        BUF1_REG_27__SCAN_IN), .ZN(n14657) );
  OAI211_X1 U17792 ( .C1(n14659), .C2(n19002), .A(n14658), .B(n14657), .ZN(
        P2_U2892) );
  INV_X1 U17793 ( .A(n14660), .ZN(n14669) );
  NAND2_X1 U17794 ( .A1(n14583), .A2(n14661), .ZN(n14662) );
  AND2_X1 U17795 ( .A1(n14663), .A2(n14662), .ZN(n15910) );
  INV_X1 U17796 ( .A(n18985), .ZN(n14665) );
  OAI22_X1 U17797 ( .A1(n14691), .A2(n14665), .B1(n14664), .B2(n18995), .ZN(
        n14666) );
  AOI21_X1 U17798 ( .B1(n19027), .B2(n15910), .A(n14666), .ZN(n14668) );
  AOI22_X1 U17799 ( .A1(n18965), .A2(BUF2_REG_26__SCAN_IN), .B1(n18964), .B2(
        BUF1_REG_26__SCAN_IN), .ZN(n14667) );
  OAI211_X1 U17800 ( .C1(n14669), .C2(n19002), .A(n14668), .B(n14667), .ZN(
        P2_U2893) );
  INV_X1 U17801 ( .A(n14855), .ZN(n14672) );
  OAI22_X1 U17802 ( .A1(n14691), .A2(n18988), .B1(n14670), .B2(n18995), .ZN(
        n14671) );
  AOI21_X1 U17803 ( .B1(n19027), .B2(n14672), .A(n14671), .ZN(n14674) );
  AOI22_X1 U17804 ( .A1(n18965), .A2(BUF2_REG_25__SCAN_IN), .B1(n18964), .B2(
        BUF1_REG_25__SCAN_IN), .ZN(n14673) );
  OAI211_X1 U17805 ( .C1(n14675), .C2(n19002), .A(n14674), .B(n14673), .ZN(
        P2_U2894) );
  AND2_X1 U17806 ( .A1(n14677), .A2(n14676), .ZN(n14679) );
  OR2_X1 U17807 ( .A1(n14679), .A2(n14678), .ZN(n15920) );
  INV_X1 U17808 ( .A(n15920), .ZN(n14683) );
  INV_X1 U17809 ( .A(n18991), .ZN(n14681) );
  OAI22_X1 U17810 ( .A1(n14691), .A2(n14681), .B1(n14680), .B2(n18995), .ZN(
        n14682) );
  AOI21_X1 U17811 ( .B1(n19027), .B2(n14683), .A(n14682), .ZN(n14685) );
  AOI22_X1 U17812 ( .A1(n18965), .A2(BUF2_REG_24__SCAN_IN), .B1(n18964), .B2(
        BUF1_REG_24__SCAN_IN), .ZN(n14684) );
  OAI211_X1 U17813 ( .C1(n14686), .C2(n19002), .A(n14685), .B(n14684), .ZN(
        P2_U2895) );
  AOI21_X1 U17814 ( .B1(n14689), .B2(n14688), .A(n14687), .ZN(n15933) );
  INV_X1 U17815 ( .A(n15933), .ZN(n14695) );
  OAI22_X1 U17816 ( .A1(n14691), .A2(n19178), .B1(n14690), .B2(n18995), .ZN(
        n14692) );
  AOI21_X1 U17817 ( .B1(n19027), .B2(n14888), .A(n14692), .ZN(n14694) );
  AOI22_X1 U17818 ( .A1(n18965), .A2(BUF2_REG_23__SCAN_IN), .B1(n18964), .B2(
        BUF1_REG_23__SCAN_IN), .ZN(n14693) );
  OAI211_X1 U17819 ( .C1(n14695), .C2(n19002), .A(n14694), .B(n14693), .ZN(
        P2_U2896) );
  NOR2_X1 U17820 ( .A1(n14697), .A2(n9661), .ZN(n14698) );
  XNOR2_X1 U17821 ( .A(n14699), .B(n14698), .ZN(n14814) );
  XOR2_X1 U17822 ( .A(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .B(n14700), .Z(
        n14812) );
  NOR2_X1 U17823 ( .A1(n15875), .A2(n16063), .ZN(n14703) );
  NAND2_X1 U17824 ( .A1(n19081), .A2(P2_REIP_REG_30__SCAN_IN), .ZN(n14808) );
  NAND2_X1 U17825 ( .A1(n16001), .A2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14701) );
  OAI211_X1 U17826 ( .C1(n14809), .C2(n16072), .A(n14808), .B(n14701), .ZN(
        n14702) );
  AOI211_X1 U17827 ( .C1(n14812), .C2(n16068), .A(n14703), .B(n14702), .ZN(
        n14704) );
  OAI21_X1 U17828 ( .B1(n14814), .B2(n19088), .A(n14704), .ZN(P2_U2984) );
  INV_X1 U17829 ( .A(n12943), .ZN(n14705) );
  OAI21_X1 U17830 ( .B1(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n10052), .A(
        n14705), .ZN(n14839) );
  INV_X1 U17831 ( .A(n14706), .ZN(n14828) );
  NAND2_X1 U17832 ( .A1(n14708), .A2(n14707), .ZN(n14827) );
  NAND3_X1 U17833 ( .A1(n14828), .A2(n16066), .A3(n14827), .ZN(n14712) );
  NAND2_X1 U17834 ( .A1(n15899), .A2(n19090), .ZN(n14709) );
  NAND2_X1 U17835 ( .A1(n19081), .A2(P2_REIP_REG_27__SCAN_IN), .ZN(n14831) );
  OAI211_X1 U17836 ( .C1(n15895), .C2(n19093), .A(n14709), .B(n14831), .ZN(
        n14710) );
  AOI21_X1 U17837 ( .B1(n19080), .B2(n15904), .A(n14710), .ZN(n14711) );
  OAI211_X1 U17838 ( .C1(n19087), .C2(n14839), .A(n14712), .B(n14711), .ZN(
        P2_U2987) );
  OAI21_X1 U17839 ( .B1(n14713), .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n14714), .ZN(n14849) );
  INV_X1 U17840 ( .A(n14715), .ZN(n14852) );
  NOR2_X1 U17841 ( .A1(n9699), .A2(n14852), .ZN(n14717) );
  MUX2_X1 U17842 ( .A(n14717), .B(n14852), .S(n14716), .Z(n14719) );
  NOR2_X1 U17843 ( .A1(n14719), .A2(n14718), .ZN(n14840) );
  NAND2_X1 U17844 ( .A1(n14840), .A2(n16066), .ZN(n14725) );
  INV_X1 U17845 ( .A(n14843), .ZN(n15911) );
  NAND2_X1 U17846 ( .A1(n19081), .A2(P2_REIP_REG_26__SCAN_IN), .ZN(n14842) );
  OAI21_X1 U17847 ( .B1(n19093), .B2(n14720), .A(n14842), .ZN(n14723) );
  NOR2_X1 U17848 ( .A1(n14721), .A2(n16063), .ZN(n14722) );
  AOI211_X1 U17849 ( .C1(n19090), .C2(n15911), .A(n14723), .B(n14722), .ZN(
        n14724) );
  OAI211_X1 U17850 ( .C1(n19087), .C2(n14849), .A(n14725), .B(n14724), .ZN(
        P2_U2988) );
  NAND3_X1 U17851 ( .A1(n14727), .A2(n9683), .A3(n14958), .ZN(n14728) );
  INV_X1 U17852 ( .A(n16020), .ZN(n14729) );
  INV_X1 U17853 ( .A(n16010), .ZN(n14730) );
  INV_X1 U17854 ( .A(n14732), .ZN(n14733) );
  AOI21_X1 U17855 ( .B1(n15294), .B2(n15295), .A(n14733), .ZN(n15320) );
  AND2_X1 U17856 ( .A1(n14735), .A2(n14734), .ZN(n15319) );
  NAND2_X1 U17857 ( .A1(n15320), .A2(n15319), .ZN(n15318) );
  NAND2_X1 U17858 ( .A1(n14738), .A2(n14737), .ZN(n14739) );
  XNOR2_X1 U17859 ( .A(n14740), .B(n14739), .ZN(n14935) );
  NOR2_X1 U17860 ( .A1(n16114), .A2(n19717), .ZN(n14923) );
  AOI21_X1 U17861 ( .B1(n16001), .B2(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .A(
        n14923), .ZN(n14741) );
  OAI21_X1 U17862 ( .B1(n18742), .B2(n16072), .A(n14741), .ZN(n14744) );
  NAND2_X1 U17863 ( .A1(n14752), .A2(n14927), .ZN(n14742) );
  NAND2_X1 U17864 ( .A1(n14901), .A2(n14742), .ZN(n14932) );
  NOR2_X1 U17865 ( .A1(n14932), .A2(n19087), .ZN(n14743) );
  AOI211_X1 U17866 ( .C1(n19080), .C2(n18738), .A(n14744), .B(n14743), .ZN(
        n14745) );
  OAI21_X1 U17867 ( .B1(n14935), .B2(n19088), .A(n14745), .ZN(P2_U2993) );
  NOR2_X1 U17868 ( .A1(n9685), .A2(n14746), .ZN(n14750) );
  NOR2_X1 U17869 ( .A1(n14748), .A2(n14747), .ZN(n14749) );
  XNOR2_X1 U17870 ( .A(n14750), .B(n14749), .ZN(n15449) );
  INV_X1 U17871 ( .A(n15019), .ZN(n14751) );
  NOR2_X1 U17872 ( .A1(n14751), .A2(n14948), .ZN(n15995) );
  INV_X1 U17873 ( .A(n15995), .ZN(n14779) );
  NOR2_X1 U17874 ( .A1(n14779), .A2(n14952), .ZN(n14778) );
  AOI21_X1 U17875 ( .B1(n14778), .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A(
        P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n14754) );
  INV_X1 U17876 ( .A(n14752), .ZN(n14753) );
  NOR2_X1 U17877 ( .A1(n14754), .A2(n14753), .ZN(n15446) );
  NOR2_X1 U17878 ( .A1(n16063), .A2(n14755), .ZN(n14762) );
  NAND2_X1 U17879 ( .A1(n14757), .A2(n14756), .ZN(n14758) );
  NAND2_X1 U17880 ( .A1(n14759), .A2(n14758), .ZN(n15445) );
  INV_X1 U17881 ( .A(P2_REIP_REG_20__SCAN_IN), .ZN(n19715) );
  NOR2_X1 U17882 ( .A1(n16114), .A2(n19715), .ZN(n15439) );
  AOI21_X1 U17883 ( .B1(n16001), .B2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .A(
        n15439), .ZN(n14760) );
  OAI21_X1 U17884 ( .B1(n15445), .B2(n16072), .A(n14760), .ZN(n14761) );
  AOI211_X1 U17885 ( .C1(n15446), .C2(n16068), .A(n14762), .B(n14761), .ZN(
        n14763) );
  OAI21_X1 U17886 ( .B1(n15449), .B2(n19088), .A(n14763), .ZN(P2_U2994) );
  NAND2_X1 U17887 ( .A1(n14765), .A2(n14764), .ZN(n14768) );
  INV_X1 U17888 ( .A(n14775), .ZN(n14766) );
  NOR2_X1 U17889 ( .A1(n9698), .A2(n14766), .ZN(n14767) );
  XOR2_X1 U17890 ( .A(n14768), .B(n14767), .Z(n14947) );
  XNOR2_X1 U17891 ( .A(n14778), .B(n14943), .ZN(n14945) );
  NAND2_X1 U17892 ( .A1(n14769), .A2(n19080), .ZN(n14771) );
  NOR2_X1 U17893 ( .A1(n16114), .A2(n19713), .ZN(n14939) );
  AOI21_X1 U17894 ( .B1(n16001), .B2(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .A(
        n14939), .ZN(n14770) );
  OAI211_X1 U17895 ( .C1(n16072), .C2(n14938), .A(n14771), .B(n14770), .ZN(
        n14772) );
  AOI21_X1 U17896 ( .B1(n14945), .B2(n16068), .A(n14772), .ZN(n14773) );
  OAI21_X1 U17897 ( .B1(n14947), .B2(n19088), .A(n14773), .ZN(P2_U2995) );
  NAND2_X1 U17898 ( .A1(n14775), .A2(n14774), .ZN(n14776) );
  XNOR2_X1 U17899 ( .A(n14777), .B(n14776), .ZN(n14957) );
  AOI21_X1 U17900 ( .B1(n14952), .B2(n14779), .A(n14778), .ZN(n14955) );
  NOR2_X1 U17901 ( .A1(n16114), .A2(n19711), .ZN(n14950) );
  OR2_X1 U17902 ( .A1(n14042), .A2(n14780), .ZN(n14781) );
  NAND2_X1 U17903 ( .A1(n14059), .A2(n14781), .ZN(n15944) );
  NOR2_X1 U17904 ( .A1(n15944), .A2(n16072), .ZN(n14782) );
  AOI211_X1 U17905 ( .C1(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .C2(n16001), .A(
        n14950), .B(n14782), .ZN(n14783) );
  OAI21_X1 U17906 ( .B1(n16063), .B2(n18765), .A(n14783), .ZN(n14784) );
  AOI21_X1 U17907 ( .B1(n14955), .B2(n16068), .A(n14784), .ZN(n14785) );
  OAI21_X1 U17908 ( .B1(n14957), .B2(n19088), .A(n14785), .ZN(P2_U2996) );
  INV_X1 U17909 ( .A(n14786), .ZN(n14787) );
  AOI21_X1 U17910 ( .B1(n13819), .B2(n14788), .A(n14787), .ZN(n14792) );
  NAND2_X1 U17911 ( .A1(n14790), .A2(n14789), .ZN(n14791) );
  XNOR2_X1 U17912 ( .A(n14792), .B(n14791), .ZN(n16126) );
  OR2_X1 U17913 ( .A1(n14794), .A2(n14793), .ZN(n14795) );
  AND2_X1 U17914 ( .A1(n14796), .A2(n14795), .ZN(n16123) );
  INV_X1 U17915 ( .A(P2_REIP_REG_8__SCAN_IN), .ZN(n19694) );
  OAI22_X1 U17916 ( .A1(n14797), .A2(n19093), .B1(n19694), .B2(n16114), .ZN(
        n14801) );
  INV_X1 U17917 ( .A(n18868), .ZN(n14799) );
  OAI22_X1 U17918 ( .A1(n16063), .A2(n14799), .B1(n16072), .B2(n14798), .ZN(
        n14800) );
  AOI211_X1 U17919 ( .C1(n16123), .C2(n16068), .A(n14801), .B(n14800), .ZN(
        n14802) );
  OAI21_X1 U17920 ( .B1(n16126), .B2(n19088), .A(n14802), .ZN(P2_U3006) );
  AOI21_X1 U17921 ( .B1(n14829), .B2(n14803), .A(
        P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n14804) );
  NOR2_X1 U17922 ( .A1(n14805), .A2(n14804), .ZN(n14811) );
  NAND2_X1 U17923 ( .A1(n19122), .A2(n14806), .ZN(n14807) );
  OAI211_X1 U17924 ( .C1(n14809), .C2(n19112), .A(n14808), .B(n14807), .ZN(
        n14810) );
  AOI211_X1 U17925 ( .C1(n14812), .C2(n16122), .A(n14811), .B(n14810), .ZN(
        n14813) );
  OAI21_X1 U17926 ( .B1(n14814), .B2(n19110), .A(n14813), .ZN(P2_U3016) );
  INV_X1 U17927 ( .A(n14818), .ZN(n14819) );
  NAND3_X1 U17928 ( .A1(n14829), .A2(n14819), .A3(n14821), .ZN(n14820) );
  AOI21_X1 U17929 ( .B1(n14824), .B2(n16122), .A(n14823), .ZN(n14825) );
  OAI21_X1 U17930 ( .B1(n14826), .B2(n19110), .A(n14825), .ZN(P2_U3017) );
  NAND3_X1 U17931 ( .A1(n14828), .A2(n12942), .A3(n14827), .ZN(n14838) );
  INV_X1 U17932 ( .A(n14829), .ZN(n14834) );
  INV_X1 U17933 ( .A(n14830), .ZN(n15908) );
  OAI21_X1 U17934 ( .B1(n16128), .B2(n15908), .A(n14831), .ZN(n14832) );
  AOI21_X1 U17935 ( .B1(n15899), .B2(n19131), .A(n14832), .ZN(n14833) );
  OAI21_X1 U17936 ( .B1(n14834), .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n14833), .ZN(n14835) );
  AOI21_X1 U17937 ( .B1(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n14836), .A(
        n14835), .ZN(n14837) );
  OAI211_X1 U17938 ( .C1(n14839), .C2(n19125), .A(n14838), .B(n14837), .ZN(
        P2_U3019) );
  NAND2_X1 U17939 ( .A1(n14840), .A2(n12942), .ZN(n14848) );
  NAND2_X1 U17940 ( .A1(n19122), .A2(n15910), .ZN(n14841) );
  OAI211_X1 U17941 ( .C1(n14843), .C2(n19112), .A(n14842), .B(n14841), .ZN(
        n14846) );
  XNOR2_X1 U17942 ( .A(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .B(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n14844) );
  NOR2_X1 U17943 ( .A1(n14859), .A2(n14844), .ZN(n14845) );
  AOI211_X1 U17944 ( .C1(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .C2(n14861), .A(
        n14846), .B(n14845), .ZN(n14847) );
  OAI211_X1 U17945 ( .C1(n14849), .C2(n19125), .A(n14848), .B(n14847), .ZN(
        P2_U3020) );
  NOR2_X1 U17946 ( .A1(n14872), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n14850) );
  OR2_X1 U17947 ( .A1(n14713), .A2(n14850), .ZN(n15963) );
  NOR2_X1 U17948 ( .A1(n14853), .A2(n14852), .ZN(n14854) );
  XNOR2_X1 U17949 ( .A(n14851), .B(n14854), .ZN(n15965) );
  NAND2_X1 U17950 ( .A1(n15965), .A2(n12942), .ZN(n14863) );
  INV_X1 U17951 ( .A(n15968), .ZN(n14857) );
  OAI22_X1 U17952 ( .A1(n16128), .A2(n14855), .B1(n19724), .B2(n12482), .ZN(
        n14856) );
  AOI21_X1 U17953 ( .B1(n14857), .B2(n19131), .A(n14856), .ZN(n14858) );
  OAI21_X1 U17954 ( .B1(n14859), .B2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n14858), .ZN(n14860) );
  AOI21_X1 U17955 ( .B1(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n14861), .A(
        n14860), .ZN(n14862) );
  OAI211_X1 U17956 ( .C1(n15963), .C2(n19125), .A(n14863), .B(n14862), .ZN(
        P2_U3021) );
  XNOR2_X1 U17957 ( .A(n14865), .B(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n14866) );
  XNOR2_X1 U17958 ( .A(n14864), .B(n14866), .ZN(n15971) );
  NAND2_X1 U17959 ( .A1(P2_REIP_REG_24__SCAN_IN), .A2(n18810), .ZN(n14867) );
  OAI211_X1 U17960 ( .C1(n14869), .C2(n14873), .A(n14868), .B(n14867), .ZN(
        n14871) );
  OAI22_X1 U17961 ( .A1(n15969), .A2(n19112), .B1(n16128), .B2(n15920), .ZN(
        n14870) );
  NOR2_X1 U17962 ( .A1(n14871), .A2(n14870), .ZN(n14877) );
  INV_X1 U17963 ( .A(n14872), .ZN(n14875) );
  NAND2_X1 U17964 ( .A1(n14880), .A2(n14873), .ZN(n14874) );
  NAND2_X1 U17965 ( .A1(n14875), .A2(n14874), .ZN(n15970) );
  OR2_X1 U17966 ( .A1(n15970), .A2(n19125), .ZN(n14876) );
  OAI211_X1 U17967 ( .C1(n15971), .C2(n19110), .A(n14877), .B(n14876), .ZN(
        P2_U3022) );
  XOR2_X1 U17968 ( .A(n14878), .B(n14879), .Z(n15981) );
  INV_X1 U17969 ( .A(n15981), .ZN(n14900) );
  OR2_X1 U17970 ( .A1(n14901), .A2(n14910), .ZN(n14903) );
  NAND2_X1 U17971 ( .A1(n14903), .A2(n14897), .ZN(n14881) );
  AND2_X1 U17972 ( .A1(n14881), .A2(n14880), .ZN(n15979) );
  INV_X1 U17973 ( .A(n14964), .ZN(n14885) );
  AOI22_X1 U17974 ( .A1(n19132), .A2(n14883), .B1(n14882), .B2(n14927), .ZN(
        n14884) );
  NAND2_X1 U17975 ( .A1(n14885), .A2(n14884), .ZN(n14929) );
  AND2_X1 U17976 ( .A1(n19116), .A2(n14927), .ZN(n14886) );
  NOR2_X1 U17977 ( .A1(n14929), .A2(n14886), .ZN(n14909) );
  NOR2_X1 U17978 ( .A1(n11581), .A2(n16114), .ZN(n14887) );
  AOI21_X1 U17979 ( .B1(n19122), .B2(n14888), .A(n14887), .ZN(n14889) );
  OAI21_X1 U17980 ( .B1(n15978), .B2(n19112), .A(n14889), .ZN(n14890) );
  INV_X1 U17981 ( .A(n14890), .ZN(n14896) );
  NAND2_X1 U17982 ( .A1(n14891), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n14936) );
  NOR2_X1 U17983 ( .A1(n15028), .A2(n14936), .ZN(n15434) );
  NAND2_X1 U17984 ( .A1(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n15433) );
  INV_X1 U17985 ( .A(n15433), .ZN(n14892) );
  AND2_X1 U17986 ( .A1(n15434), .A2(n14892), .ZN(n14928) );
  NAND2_X1 U17987 ( .A1(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n14928), .ZN(
        n14911) );
  AOI21_X1 U17988 ( .B1(n14910), .B2(n14897), .A(n14911), .ZN(n14894) );
  NAND2_X1 U17989 ( .A1(n14894), .A2(n14893), .ZN(n14895) );
  OAI211_X1 U17990 ( .C1(n14909), .C2(n14897), .A(n14896), .B(n14895), .ZN(
        n14898) );
  AOI21_X1 U17991 ( .B1(n15979), .B2(n16122), .A(n14898), .ZN(n14899) );
  OAI21_X1 U17992 ( .B1(n14900), .B2(n19110), .A(n14899), .ZN(P2_U3023) );
  NAND2_X1 U17993 ( .A1(n14901), .A2(n14910), .ZN(n14902) );
  NAND2_X1 U17994 ( .A1(n14903), .A2(n14902), .ZN(n15986) );
  NAND2_X1 U17995 ( .A1(n14905), .A2(n14904), .ZN(n14907) );
  XOR2_X1 U17996 ( .A(n14907), .B(n14906), .Z(n15987) );
  OR2_X1 U17997 ( .A1(n15987), .A2(n19110), .ZN(n14922) );
  NAND2_X1 U17998 ( .A1(P2_REIP_REG_22__SCAN_IN), .A2(n19081), .ZN(n14908) );
  OAI221_X1 U17999 ( .B1(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n14911), 
        .C1(n14910), .C2(n14909), .A(n14908), .ZN(n14920) );
  OR2_X1 U18000 ( .A1(n14913), .A2(n14912), .ZN(n14914) );
  NAND2_X1 U18001 ( .A1(n12980), .A2(n14914), .ZN(n15311) );
  OR2_X1 U18002 ( .A1(n14916), .A2(n14915), .ZN(n14917) );
  AND2_X1 U18003 ( .A1(n12977), .A2(n14917), .ZN(n15989) );
  NAND2_X1 U18004 ( .A1(n15989), .A2(n19131), .ZN(n14918) );
  OAI21_X1 U18005 ( .B1(n16128), .B2(n15311), .A(n14918), .ZN(n14919) );
  NOR2_X1 U18006 ( .A1(n14920), .A2(n14919), .ZN(n14921) );
  OAI211_X1 U18007 ( .C1(n15986), .C2(n19125), .A(n14922), .B(n14921), .ZN(
        P2_U3024) );
  INV_X1 U18008 ( .A(n14923), .ZN(n14925) );
  NAND2_X1 U18009 ( .A1(n19122), .A2(n18743), .ZN(n14924) );
  OAI211_X1 U18010 ( .C1(n18742), .C2(n19112), .A(n14925), .B(n14924), .ZN(
        n14926) );
  AOI21_X1 U18011 ( .B1(n14928), .B2(n14927), .A(n14926), .ZN(n14931) );
  NAND2_X1 U18012 ( .A1(n14929), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n14930) );
  OAI211_X1 U18013 ( .C1(n14932), .C2(n19125), .A(n14931), .B(n14930), .ZN(
        n14933) );
  INV_X1 U18014 ( .A(n14933), .ZN(n14934) );
  OAI21_X1 U18015 ( .B1(n14935), .B2(n19110), .A(n14934), .ZN(P2_U3025) );
  OAI21_X1 U18016 ( .B1(n14964), .B2(n14936), .A(n15296), .ZN(n15436) );
  NAND2_X1 U18017 ( .A1(n14937), .A2(n19122), .ZN(n14942) );
  NOR2_X1 U18018 ( .A1(n19112), .A2(n14938), .ZN(n14940) );
  AOI211_X1 U18019 ( .C1(n15434), .C2(n14943), .A(n14940), .B(n14939), .ZN(
        n14941) );
  OAI211_X1 U18020 ( .C1(n14943), .C2(n15436), .A(n14942), .B(n14941), .ZN(
        n14944) );
  AOI21_X1 U18021 ( .B1(n14945), .B2(n16122), .A(n14944), .ZN(n14946) );
  OAI21_X1 U18022 ( .B1(n14947), .B2(n19110), .A(n14946), .ZN(P2_U3027) );
  NOR2_X1 U18023 ( .A1(n18770), .A2(n16128), .ZN(n14954) );
  INV_X1 U18024 ( .A(n15944), .ZN(n18766) );
  NOR3_X1 U18025 ( .A1(n15028), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A3(
        n14948), .ZN(n14949) );
  AOI211_X1 U18026 ( .C1(n18766), .C2(n19131), .A(n14950), .B(n14949), .ZN(
        n14951) );
  OAI21_X1 U18027 ( .B1(n14952), .B2(n15436), .A(n14951), .ZN(n14953) );
  AOI211_X1 U18028 ( .C1(n14955), .C2(n16122), .A(n14954), .B(n14953), .ZN(
        n14956) );
  OAI21_X1 U18029 ( .B1(n14957), .B2(n19110), .A(n14956), .ZN(P2_U3028) );
  INV_X1 U18030 ( .A(n16039), .ZN(n14980) );
  NAND2_X1 U18031 ( .A1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n14980), .ZN(
        n16037) );
  AOI21_X1 U18032 ( .B1(n16085), .B2(n16037), .A(n16018), .ZN(n16030) );
  INV_X1 U18033 ( .A(n16030), .ZN(n14974) );
  NAND2_X1 U18034 ( .A1(n14959), .A2(n14958), .ZN(n14961) );
  XOR2_X1 U18035 ( .A(n14961), .B(n14960), .Z(n16029) );
  INV_X1 U18036 ( .A(n15028), .ZN(n14962) );
  NAND2_X1 U18037 ( .A1(n14963), .A2(n14962), .ZN(n16083) );
  NOR2_X1 U18038 ( .A1(n15029), .A2(n14964), .ZN(n15027) );
  AOI21_X1 U18039 ( .B1(n9785), .B2(n15027), .A(n14986), .ZN(n16103) );
  AOI21_X1 U18040 ( .B1(n16107), .B2(n16106), .A(n16103), .ZN(n14965) );
  NOR2_X1 U18041 ( .A1(n14965), .A2(n16085), .ZN(n14972) );
  OAI21_X1 U18042 ( .B1(n16101), .B2(n14966), .A(n16090), .ZN(n18979) );
  NOR2_X1 U18043 ( .A1(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n16083), .ZN(
        n14969) );
  INV_X1 U18044 ( .A(P2_REIP_REG_13__SCAN_IN), .ZN(n19703) );
  NOR2_X1 U18045 ( .A1(n19703), .A2(n16114), .ZN(n14968) );
  NOR2_X1 U18046 ( .A1(n18824), .A2(n19112), .ZN(n14967) );
  AOI211_X1 U18047 ( .C1(n14969), .C2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n14968), .B(n14967), .ZN(n14970) );
  OAI21_X1 U18048 ( .B1(n18979), .B2(n16128), .A(n14970), .ZN(n14971) );
  AOI211_X1 U18049 ( .C1(n16029), .C2(n12942), .A(n14972), .B(n14971), .ZN(
        n14973) );
  OAI21_X1 U18050 ( .B1(n14974), .B2(n19125), .A(n14973), .ZN(P2_U3033) );
  NAND2_X1 U18051 ( .A1(n14975), .A2(n14976), .ZN(n14979) );
  NAND2_X1 U18052 ( .A1(n10105), .A2(n14977), .ZN(n14978) );
  XNOR2_X1 U18053 ( .A(n14979), .B(n14978), .ZN(n16045) );
  INV_X1 U18054 ( .A(n16045), .ZN(n14996) );
  NAND2_X1 U18055 ( .A1(n9786), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n14981) );
  AOI21_X1 U18056 ( .B1(n14988), .B2(n14981), .A(n14980), .ZN(n16046) );
  OAI21_X1 U18057 ( .B1(n14984), .B2(n14983), .A(n14982), .ZN(n18984) );
  NOR2_X1 U18058 ( .A1(n15029), .A2(n15028), .ZN(n15007) );
  OAI211_X1 U18059 ( .C1(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A(n15007), .B(n14985), .ZN(
        n14993) );
  INV_X1 U18060 ( .A(n18846), .ZN(n14991) );
  NOR2_X1 U18061 ( .A1(n14986), .A2(n15027), .ZN(n15008) );
  INV_X1 U18062 ( .A(n15008), .ZN(n14987) );
  OAI22_X1 U18063 ( .A1(n16114), .A2(n14989), .B1(n14988), .B2(n14987), .ZN(
        n14990) );
  AOI21_X1 U18064 ( .B1(n19131), .B2(n14991), .A(n14990), .ZN(n14992) );
  OAI211_X1 U18065 ( .C1(n18984), .C2(n16128), .A(n14993), .B(n14992), .ZN(
        n14994) );
  AOI21_X1 U18066 ( .B1(n16046), .B2(n16122), .A(n14994), .ZN(n14995) );
  OAI21_X1 U18067 ( .B1(n14996), .B2(n19110), .A(n14995), .ZN(P2_U3035) );
  XNOR2_X1 U18068 ( .A(n15021), .B(n15006), .ZN(n16049) );
  NOR2_X1 U18069 ( .A1(n14997), .A2(n15024), .ZN(n15002) );
  INV_X1 U18070 ( .A(n14998), .ZN(n14999) );
  NAND2_X1 U18071 ( .A1(n15000), .A2(n14999), .ZN(n15001) );
  XNOR2_X1 U18072 ( .A(n15002), .B(n15001), .ZN(n16050) );
  INV_X1 U18073 ( .A(n16050), .ZN(n15017) );
  XNOR2_X1 U18074 ( .A(n15004), .B(n15003), .ZN(n18987) );
  INV_X1 U18075 ( .A(P2_REIP_REG_10__SCAN_IN), .ZN(n19698) );
  NOR2_X1 U18076 ( .A1(n19698), .A2(n16114), .ZN(n15005) );
  AOI221_X1 U18077 ( .B1(n15008), .B2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), 
        .C1(n15007), .C2(n15006), .A(n15005), .ZN(n15015) );
  INV_X1 U18078 ( .A(n15009), .ZN(n15010) );
  NAND2_X1 U18079 ( .A1(n15011), .A2(n15010), .ZN(n15013) );
  AND2_X1 U18080 ( .A1(n15013), .A2(n15012), .ZN(n18956) );
  NAND2_X1 U18081 ( .A1(n19131), .A2(n18956), .ZN(n15014) );
  OAI211_X1 U18082 ( .C1(n16128), .C2(n18987), .A(n15015), .B(n15014), .ZN(
        n15016) );
  AOI21_X1 U18083 ( .B1(n15017), .B2(n12942), .A(n15016), .ZN(n15018) );
  OAI21_X1 U18084 ( .B1(n19125), .B2(n16049), .A(n15018), .ZN(P2_U3036) );
  OR2_X1 U18085 ( .A1(n15019), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n15020) );
  AND2_X1 U18086 ( .A1(n15021), .A2(n15020), .ZN(n16059) );
  INV_X1 U18087 ( .A(n16059), .ZN(n15035) );
  NOR2_X1 U18088 ( .A1(n15024), .A2(n15023), .ZN(n15025) );
  XNOR2_X1 U18089 ( .A(n15022), .B(n15025), .ZN(n16058) );
  NAND2_X1 U18090 ( .A1(n15026), .A2(n19122), .ZN(n15032) );
  AOI21_X1 U18091 ( .B1(n15029), .B2(n15028), .A(n15027), .ZN(n15030) );
  AOI21_X1 U18092 ( .B1(n19081), .B2(P2_REIP_REG_9__SCAN_IN), .A(n15030), .ZN(
        n15031) );
  OAI211_X1 U18093 ( .C1(n19112), .C2(n16062), .A(n15032), .B(n15031), .ZN(
        n15033) );
  AOI21_X1 U18094 ( .B1(n16058), .B2(n12942), .A(n15033), .ZN(n15034) );
  OAI21_X1 U18095 ( .B1(n15035), .B2(n19125), .A(n15034), .ZN(P2_U3037) );
  AOI21_X1 U18096 ( .B1(n15036), .B2(n19594), .A(P2_STATE2_REG_1__SCAN_IN), 
        .ZN(n15039) );
  INV_X1 U18097 ( .A(n15037), .ZN(n16148) );
  OAI22_X1 U18098 ( .A1(n15040), .A2(n15039), .B1(n15038), .B2(n16148), .ZN(
        n15041) );
  MUX2_X1 U18099 ( .A(n15041), .B(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .S(
        n15044), .Z(P2_U3601) );
  INV_X1 U18100 ( .A(n15042), .ZN(n19749) );
  OAI22_X1 U18101 ( .A1(n19000), .A2(n16148), .B1(n15043), .B2(n19749), .ZN(
        n15045) );
  MUX2_X1 U18102 ( .A(n15045), .B(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(
        n15044), .Z(P2_U3596) );
  NAND2_X1 U18103 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n18198) );
  AOI221_X1 U18104 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(n18198), .C1(n15047), 
        .C2(n18198), .A(n15046), .ZN(n18042) );
  INV_X1 U18105 ( .A(n15048), .ZN(n15049) );
  INV_X1 U18106 ( .A(n16171), .ZN(n18385) );
  NAND2_X1 U18107 ( .A1(n18517), .A2(n18385), .ZN(n18223) );
  OAI211_X1 U18108 ( .C1(n16171), .C2(n15049), .A(n18043), .B(n18223), .ZN(
        n18040) );
  AOI22_X1 U18109 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n18042), .B1(
        n18040), .B2(n18522), .ZN(P3_U2865) );
  NOR2_X1 U18110 ( .A1(n17078), .A2(n18071), .ZN(n15053) );
  NAND4_X1 U18111 ( .A1(n18068), .A2(n15076), .A3(n15079), .A4(n15053), .ZN(
        n15077) );
  NOR2_X1 U18112 ( .A1(n15221), .A2(n15077), .ZN(n15068) );
  NAND2_X1 U18113 ( .A1(n15221), .A2(n15234), .ZN(n15059) );
  NOR2_X1 U18114 ( .A1(n18076), .A2(n18071), .ZN(n18511) );
  OAI211_X1 U18115 ( .C1(n18068), .C2(n18511), .A(n15236), .B(n15050), .ZN(
        n15051) );
  NOR2_X1 U18116 ( .A1(n15059), .A2(n15051), .ZN(n15217) );
  INV_X1 U18117 ( .A(n15053), .ZN(n15222) );
  NAND2_X1 U18118 ( .A1(n18495), .A2(n15221), .ZN(n15066) );
  NOR3_X1 U18119 ( .A1(n15052), .A2(n15066), .A3(n17227), .ZN(n15058) );
  NOR2_X1 U18120 ( .A1(n18087), .A2(n15053), .ZN(n15056) );
  INV_X1 U18121 ( .A(n15076), .ZN(n18063) );
  OR2_X1 U18122 ( .A1(n18063), .A2(n15079), .ZN(n15055) );
  NAND2_X1 U18123 ( .A1(n18068), .A2(n18511), .ZN(n15054) );
  OAI211_X1 U18124 ( .C1(n18068), .C2(n15056), .A(n15055), .B(n15054), .ZN(
        n15057) );
  NOR2_X1 U18125 ( .A1(n17291), .A2(n18047), .ZN(n15232) );
  OAI21_X1 U18126 ( .B1(n18087), .B2(n18511), .A(n15232), .ZN(n15071) );
  OAI211_X1 U18127 ( .C1(n15068), .C2(n15217), .A(n15074), .B(n15071), .ZN(
        n15223) );
  XOR2_X1 U18128 ( .A(n15061), .B(n15060), .Z(n15065) );
  INV_X1 U18129 ( .A(n15062), .ZN(n15063) );
  NAND2_X1 U18130 ( .A1(READY22_REG_SCAN_IN), .A2(READY2), .ZN(n18693) );
  NAND2_X1 U18131 ( .A1(n18482), .A2(n18693), .ZN(n15086) );
  INV_X1 U18132 ( .A(P3_STATE_REG_0__SCAN_IN), .ZN(n18567) );
  INV_X1 U18133 ( .A(P3_STATE_REG_1__SCAN_IN), .ZN(n18559) );
  INV_X2 U18134 ( .A(n18701), .ZN(n18703) );
  OAI211_X1 U18135 ( .C1(P3_STATE_REG_1__SCAN_IN), .C2(P3_STATE_REG_2__SCAN_IN), .A(n18567), .B(n18631), .ZN(n18690) );
  INV_X1 U18136 ( .A(n18690), .ZN(n16364) );
  NOR2_X1 U18137 ( .A1(n15069), .A2(n15068), .ZN(n16348) );
  NAND2_X1 U18138 ( .A1(n18692), .A2(n15069), .ZN(n18481) );
  NAND2_X1 U18139 ( .A1(n16364), .A2(n15080), .ZN(n17226) );
  XNOR2_X1 U18140 ( .A(n18692), .B(n15221), .ZN(n15226) );
  INV_X1 U18141 ( .A(n15226), .ZN(n15070) );
  NAND2_X1 U18142 ( .A1(n15070), .A2(n15069), .ZN(n17290) );
  INV_X1 U18143 ( .A(n15071), .ZN(n15072) );
  AOI21_X1 U18144 ( .B1(n15227), .B2(n15073), .A(n15072), .ZN(n15075) );
  NOR2_X2 U18145 ( .A1(n15077), .A2(n15237), .ZN(n15231) );
  NAND3_X1 U18146 ( .A1(n15079), .A2(n15078), .A3(n18692), .ZN(n15081) );
  INV_X1 U18147 ( .A(n15239), .ZN(n15082) );
  INV_X1 U18148 ( .A(n18483), .ZN(n15083) );
  OAI211_X1 U18149 ( .C1(n15086), .C2(n17226), .A(n15085), .B(n15431), .ZN(
        n15087) );
  INV_X1 U18150 ( .A(n18520), .ZN(n15089) );
  NOR2_X1 U18151 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n18639), .ZN(n18046) );
  NOR2_X1 U18152 ( .A1(n16350), .A2(n18638), .ZN(n15088) );
  AOI211_X1 U18153 ( .C1(n18686), .C2(n15089), .A(n18046), .B(n15088), .ZN(
        n18669) );
  INV_X1 U18154 ( .A(n18669), .ZN(n18666) );
  NOR2_X1 U18155 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n18705) );
  AOI21_X1 U18156 ( .B1(n15090), .B2(n16701), .A(n18483), .ZN(n18492) );
  NAND3_X1 U18157 ( .A1(n18666), .A2(n18705), .A3(n18492), .ZN(n15091) );
  OAI21_X1 U18158 ( .B1(n18666), .B2(n16701), .A(n15091), .ZN(P3_U3284) );
  INV_X1 U18159 ( .A(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n17349) );
  AOI22_X1 U18160 ( .A1(n16977), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n17023), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n15101) );
  AOI22_X1 U18161 ( .A1(n9633), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n17022), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n15100) );
  AOI22_X1 U18162 ( .A1(n9627), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n17021), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n15092) );
  OAI21_X1 U18163 ( .B1(n15148), .B2(n17039), .A(n15092), .ZN(n15098) );
  AOI22_X1 U18164 ( .A1(n17005), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n16995), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n15096) );
  AOI22_X1 U18165 ( .A1(n17020), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n15158), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n15095) );
  AOI22_X1 U18166 ( .A1(n16998), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n9626), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n15094) );
  AOI22_X1 U18167 ( .A1(n16992), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n17014), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n15093) );
  NAND4_X1 U18168 ( .A1(n15096), .A2(n15095), .A3(n15094), .A4(n15093), .ZN(
        n15097) );
  AOI211_X1 U18169 ( .C1(n16989), .C2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A(
        n15098), .B(n15097), .ZN(n15099) );
  AOI22_X1 U18170 ( .A1(n16958), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n17023), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n15105) );
  AOI22_X1 U18171 ( .A1(n17020), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n15158), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n15104) );
  AOI22_X1 U18172 ( .A1(n16989), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n17021), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n15103) );
  AOI22_X1 U18173 ( .A1(n9627), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n15174), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n15102) );
  NAND4_X1 U18174 ( .A1(n15105), .A2(n15104), .A3(n15103), .A4(n15102), .ZN(
        n15112) );
  AOI22_X1 U18175 ( .A1(n16992), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n17022), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n15110) );
  AOI22_X1 U18176 ( .A1(n16997), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n9633), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n15109) );
  AOI22_X1 U18177 ( .A1(n16924), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n9626), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n15108) );
  AOI22_X1 U18178 ( .A1(n17005), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n16977), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n15107) );
  NAND4_X1 U18179 ( .A1(n15110), .A2(n15109), .A3(n15108), .A4(n15107), .ZN(
        n15111) );
  AOI22_X1 U18180 ( .A1(n16977), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n17022), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n15116) );
  AOI22_X1 U18181 ( .A1(n17020), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n15158), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n15115) );
  AOI22_X1 U18182 ( .A1(n16997), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n17013), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n15114) );
  AOI22_X1 U18183 ( .A1(n17021), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n15174), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n15113) );
  NAND4_X1 U18184 ( .A1(n15116), .A2(n15115), .A3(n15114), .A4(n15113), .ZN(
        n15122) );
  AOI22_X1 U18185 ( .A1(n17005), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n9633), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n15120) );
  AOI22_X1 U18186 ( .A1(n16989), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n16995), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n15119) );
  AOI22_X1 U18187 ( .A1(n15106), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n16974), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n15118) );
  AOI22_X1 U18188 ( .A1(n16923), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n16975), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n15117) );
  NAND4_X1 U18189 ( .A1(n15120), .A2(n15119), .A3(n15118), .A4(n15117), .ZN(
        n15121) );
  AOI22_X1 U18190 ( .A1(n16825), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n15158), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n15124) );
  AOI22_X1 U18191 ( .A1(n9627), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n9626), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n15123) );
  AOI22_X1 U18192 ( .A1(n16924), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n16975), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n15125) );
  OAI21_X1 U18193 ( .B1(n15148), .B2(n17061), .A(n15125), .ZN(n15126) );
  INV_X1 U18194 ( .A(n15126), .ZN(n15133) );
  AOI22_X1 U18195 ( .A1(n13962), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n15127), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n15131) );
  AOI22_X1 U18196 ( .A1(n16958), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n13926), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n15130) );
  AOI22_X1 U18197 ( .A1(n15106), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n15139), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n15129) );
  AOI22_X1 U18198 ( .A1(n15134), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n15174), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n15128) );
  NAND2_X1 U18199 ( .A1(n16977), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(
        n15132) );
  AOI22_X1 U18200 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n9627), .B1(
        n15134), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n15135) );
  OAI21_X1 U18201 ( .B1(n17065), .B2(n15148), .A(n15135), .ZN(n15138) );
  AOI22_X1 U18202 ( .A1(n13881), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n9626), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n15136) );
  NOR2_X1 U18203 ( .A1(n15138), .A2(n15137), .ZN(n15146) );
  AOI22_X1 U18204 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n15139), .B1(
        n16958), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n15145) );
  AOI22_X1 U18205 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n15127), .B1(
        P3_INSTQUEUE_REG_3__1__SCAN_IN), .B2(n15172), .ZN(n15143) );
  AOI22_X1 U18206 ( .A1(n15106), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n13926), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n15142) );
  AOI22_X1 U18207 ( .A1(n16924), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_12__1__SCAN_IN), .B2(n16975), .ZN(n15141) );
  AOI22_X1 U18208 ( .A1(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n15174), .B1(
        P3_INSTQUEUE_REG_9__1__SCAN_IN), .B2(n15173), .ZN(n15140) );
  AOI22_X1 U18209 ( .A1(n16923), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n17023), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n15157) );
  AOI22_X1 U18210 ( .A1(n16996), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n17022), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n15156) );
  AOI22_X1 U18211 ( .A1(n15106), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n17013), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n15147) );
  OAI21_X1 U18212 ( .B1(n15148), .B2(n17051), .A(n15147), .ZN(n15154) );
  AOI22_X1 U18213 ( .A1(n16977), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n16995), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n15152) );
  AOI22_X1 U18214 ( .A1(n9633), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n16991), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n15151) );
  AOI22_X1 U18215 ( .A1(n9627), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n16825), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n15150) );
  AOI22_X1 U18216 ( .A1(n16989), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n15174), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n15149) );
  NAND4_X1 U18217 ( .A1(n15152), .A2(n15151), .A3(n15150), .A4(n15149), .ZN(
        n15153) );
  AOI211_X1 U18218 ( .C1(n17005), .C2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .A(
        n15154), .B(n15153), .ZN(n15155) );
  NAND3_X1 U18219 ( .A1(n15157), .A2(n15156), .A3(n15155), .ZN(n15254) );
  NAND2_X1 U18220 ( .A1(n15191), .A2(n15254), .ZN(n15193) );
  AOI22_X1 U18221 ( .A1(n16997), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n16974), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n15168) );
  AOI22_X1 U18222 ( .A1(n16992), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n17023), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n15167) );
  INV_X1 U18223 ( .A(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n16823) );
  AOI22_X1 U18224 ( .A1(n17020), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n15158), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n15159) );
  OAI21_X1 U18225 ( .B1(n16994), .B2(n16823), .A(n15159), .ZN(n15165) );
  AOI22_X1 U18226 ( .A1(n16989), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n17022), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n15163) );
  AOI22_X1 U18227 ( .A1(n17005), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n17013), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n15162) );
  AOI22_X1 U18228 ( .A1(n16977), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n17021), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n15161) );
  AOI22_X1 U18229 ( .A1(n16924), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n9633), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n15160) );
  NAND4_X1 U18230 ( .A1(n15163), .A2(n15162), .A3(n15161), .A4(n15160), .ZN(
        n15164) );
  AOI211_X1 U18231 ( .C1(n16923), .C2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .A(
        n15165), .B(n15164), .ZN(n15166) );
  NAND3_X1 U18232 ( .A1(n15168), .A2(n15167), .A3(n15166), .ZN(n15258) );
  INV_X1 U18233 ( .A(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n17632) );
  INV_X1 U18234 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n17678) );
  AOI22_X1 U18235 ( .A1(n15139), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n16958), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n15183) );
  AOI22_X1 U18236 ( .A1(n15106), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n16991), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n15182) );
  AOI22_X1 U18237 ( .A1(n9627), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n16975), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n15169) );
  OAI21_X1 U18238 ( .B1(n15170), .B2(n20830), .A(n15169), .ZN(n15180) );
  AOI22_X1 U18239 ( .A1(n13926), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n9626), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n15178) );
  AOI22_X1 U18240 ( .A1(n13962), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n15171), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n15177) );
  AOI22_X1 U18241 ( .A1(n16990), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n15172), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n15176) );
  AOI22_X1 U18242 ( .A1(n15174), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n15173), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n15175) );
  NAND4_X1 U18243 ( .A1(n15178), .A2(n15177), .A3(n15176), .A4(n15175), .ZN(
        n15179) );
  AOI211_X1 U18244 ( .C1(n16924), .C2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .A(
        n15180), .B(n15179), .ZN(n15181) );
  NAND3_X1 U18245 ( .A1(n15183), .A2(n15182), .A3(n15181), .ZN(n17706) );
  INV_X1 U18246 ( .A(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n18652) );
  NOR2_X1 U18247 ( .A1(n17220), .A2(n18652), .ZN(n15184) );
  NOR2_X2 U18248 ( .A1(n17698), .A2(n15184), .ZN(n17689) );
  INV_X1 U18249 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n18011) );
  XNOR2_X1 U18250 ( .A(n15185), .B(n18011), .ZN(n17690) );
  NOR2_X1 U18251 ( .A1(n18011), .A2(n15185), .ZN(n15186) );
  XNOR2_X1 U18252 ( .A(n15244), .B(n15188), .ZN(n15189) );
  XNOR2_X1 U18253 ( .A(n15190), .B(n15189), .ZN(n17677) );
  INV_X1 U18254 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n17980) );
  INV_X1 U18255 ( .A(n17201), .ZN(n15240) );
  XOR2_X1 U18256 ( .A(n15240), .B(n15193), .Z(n15194) );
  INV_X1 U18257 ( .A(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n17969) );
  NOR2_X1 U18258 ( .A1(n15195), .A2(n15194), .ZN(n15196) );
  XNOR2_X1 U18259 ( .A(n17198), .B(n15197), .ZN(n15198) );
  XNOR2_X1 U18260 ( .A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .B(n15198), .ZN(
        n17642) );
  AND2_X1 U18261 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n15198), .ZN(
        n15199) );
  NOR2_X1 U18262 ( .A1(n17632), .A2(n17630), .ZN(n17631) );
  NOR2_X1 U18263 ( .A1(n15201), .A2(n15200), .ZN(n15202) );
  NOR2_X2 U18264 ( .A1(n17631), .A2(n15202), .ZN(n17500) );
  NAND2_X1 U18265 ( .A1(n17500), .A2(n17615), .ZN(n15230) );
  NOR2_X1 U18266 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n17588) );
  INV_X1 U18267 ( .A(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n17543) );
  INV_X1 U18268 ( .A(n17500), .ZN(n15203) );
  XNOR2_X2 U18269 ( .A(n15203), .B(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n17939) );
  NOR2_X1 U18270 ( .A1(n17615), .A2(n17939), .ZN(n17614) );
  INV_X1 U18271 ( .A(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n17936) );
  INV_X1 U18272 ( .A(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n17922) );
  NOR2_X1 U18273 ( .A1(n17936), .A2(n17922), .ZN(n17910) );
  NAND2_X1 U18274 ( .A1(n17910), .A2(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n17895) );
  NOR3_X1 U18275 ( .A1(n17500), .A2(n17614), .A3(n17895), .ZN(n17559) );
  NAND2_X1 U18276 ( .A1(n17559), .A2(n10119), .ZN(n17524) );
  INV_X1 U18277 ( .A(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n17894) );
  INV_X1 U18278 ( .A(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n17845) );
  INV_X1 U18279 ( .A(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n17840) );
  NAND2_X1 U18280 ( .A1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n17485) );
  INV_X1 U18281 ( .A(n17485), .ZN(n17818) );
  NAND2_X1 U18282 ( .A1(n17818), .A2(n15205), .ZN(n17445) );
  INV_X1 U18283 ( .A(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n17810) );
  INV_X1 U18284 ( .A(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n17451) );
  NOR2_X1 U18285 ( .A1(n17810), .A2(n17451), .ZN(n17791) );
  NAND3_X1 U18286 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A3(n17791), .ZN(n17766) );
  INV_X1 U18287 ( .A(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n17436) );
  NOR2_X1 U18288 ( .A1(n17766), .A2(n17436), .ZN(n16237) );
  NAND2_X1 U18289 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(n16237), .ZN(
        n15209) );
  NOR2_X1 U18290 ( .A1(n17485), .A2(n15209), .ZN(n15271) );
  NAND2_X1 U18291 ( .A1(n15205), .A2(n15271), .ZN(n15207) );
  NAND2_X1 U18292 ( .A1(n17482), .A2(n17810), .ZN(n15206) );
  NOR2_X1 U18293 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n15206), .ZN(
        n17446) );
  INV_X1 U18294 ( .A(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n17774) );
  NAND2_X1 U18295 ( .A1(n17446), .A2(n17774), .ZN(n17435) );
  NOR2_X2 U18296 ( .A1(n17400), .A2(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n17399) );
  NOR3_X1 U18297 ( .A1(n17484), .A2(n17399), .A3(n15209), .ZN(n15210) );
  NAND2_X1 U18298 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n17715) );
  NAND2_X1 U18299 ( .A1(n9690), .A2(n10106), .ZN(n15211) );
  INV_X1 U18300 ( .A(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n17738) );
  NOR2_X2 U18301 ( .A1(n15211), .A2(n17374), .ZN(n15212) );
  NOR2_X1 U18302 ( .A1(n15213), .A2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n15214) );
  OAI21_X1 U18303 ( .B1(n17349), .B2(n16219), .A(n15393), .ZN(n15215) );
  XNOR2_X1 U18304 ( .A(n15215), .B(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n16202) );
  NAND2_X1 U18305 ( .A1(n15221), .A2(n17291), .ZN(n15216) );
  NOR2_X1 U18306 ( .A1(n17078), .A2(n15216), .ZN(n15225) );
  NAND2_X1 U18307 ( .A1(n15225), .A2(n15217), .ZN(n16226) );
  INV_X1 U18308 ( .A(n16226), .ZN(n18490) );
  INV_X1 U18309 ( .A(n15218), .ZN(n15220) );
  INV_X1 U18310 ( .A(n18482), .ZN(n16347) );
  AOI21_X1 U18311 ( .B1(n15220), .B2(n15219), .A(n16347), .ZN(n16154) );
  INV_X1 U18312 ( .A(n15221), .ZN(n18058) );
  AOI211_X1 U18313 ( .C1(n18068), .C2(n15222), .A(n18058), .B(n16155), .ZN(
        n15224) );
  AOI211_X1 U18314 ( .C1(n15225), .C2(n16154), .A(n15224), .B(n15223), .ZN(
        n15229) );
  INV_X1 U18315 ( .A(n18693), .ZN(n18688) );
  AOI21_X1 U18316 ( .B1(n15226), .B2(n18690), .A(n18688), .ZN(n16346) );
  NAND3_X1 U18317 ( .A1(n16346), .A2(n15227), .A3(n18482), .ZN(n15228) );
  INV_X1 U18318 ( .A(n18686), .ZN(n18534) );
  NAND3_X1 U18319 ( .A1(n18490), .A2(n18025), .A3(n17193), .ZN(n17940) );
  NAND2_X1 U18320 ( .A1(n18490), .A2(n18025), .ZN(n18031) );
  NOR2_X1 U18321 ( .A1(n17193), .A2(n18031), .ZN(n17877) );
  INV_X1 U18322 ( .A(n17877), .ZN(n17938) );
  INV_X1 U18323 ( .A(n17715), .ZN(n15274) );
  INV_X1 U18324 ( .A(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n17748) );
  NAND2_X1 U18325 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n15230), .ZN(
        n16182) );
  INV_X1 U18326 ( .A(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n17867) );
  INV_X1 U18327 ( .A(n17895), .ZN(n17882) );
  NAND2_X1 U18328 ( .A1(n17882), .A2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n17861) );
  INV_X1 U18329 ( .A(n17861), .ZN(n17554) );
  NAND2_X1 U18330 ( .A1(n17554), .A2(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n17536) );
  NOR2_X1 U18331 ( .A1(n17867), .A2(n17536), .ZN(n17836) );
  NAND2_X1 U18332 ( .A1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n17836), .ZN(
        n17820) );
  NAND2_X1 U18333 ( .A1(n15271), .A2(n17846), .ZN(n17750) );
  NAND2_X1 U18334 ( .A1(n15274), .A2(n17396), .ZN(n17720) );
  INV_X1 U18335 ( .A(n17720), .ZN(n17348) );
  NAND3_X1 U18336 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A3(n17348), .ZN(n16227) );
  INV_X1 U18337 ( .A(n15232), .ZN(n15233) );
  NAND2_X1 U18338 ( .A1(n15234), .A2(n15233), .ZN(n18706) );
  NAND2_X1 U18339 ( .A1(n18695), .A2(n15235), .ZN(n18509) );
  NOR2_X1 U18340 ( .A1(n18692), .A2(n15236), .ZN(n15238) );
  NAND2_X1 U18341 ( .A1(n17706), .A2(n17220), .ZN(n15245) );
  NAND2_X1 U18342 ( .A1(n9612), .A2(n15245), .ZN(n15243) );
  NAND2_X1 U18343 ( .A1(n15243), .A2(n15244), .ZN(n15255) );
  NOR2_X1 U18344 ( .A1(n17205), .A2(n15255), .ZN(n15241) );
  NAND2_X1 U18345 ( .A1(n15241), .A2(n15240), .ZN(n15259) );
  NOR2_X1 U18346 ( .A1(n17198), .A2(n15259), .ZN(n15263) );
  NAND2_X1 U18347 ( .A1(n15263), .A2(n17193), .ZN(n15264) );
  XNOR2_X1 U18348 ( .A(n15241), .B(n17201), .ZN(n15242) );
  AND2_X1 U18349 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n15242), .ZN(
        n15257) );
  XNOR2_X1 U18350 ( .A(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .B(n15242), .ZN(
        n17653) );
  XNOR2_X1 U18351 ( .A(n15244), .B(n15243), .ZN(n15252) );
  NOR2_X1 U18352 ( .A1(n15252), .A2(n17678), .ZN(n15253) );
  XOR2_X1 U18353 ( .A(n9612), .B(n15245), .Z(n15246) );
  NOR2_X1 U18354 ( .A1(n15246), .A2(n18011), .ZN(n15251) );
  XNOR2_X1 U18355 ( .A(n18011), .B(n15246), .ZN(n17688) );
  INV_X1 U18356 ( .A(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n18665) );
  NOR2_X1 U18357 ( .A1(n15248), .A2(n18665), .ZN(n15250) );
  INV_X1 U18358 ( .A(n17706), .ZN(n15249) );
  NAND3_X1 U18359 ( .A1(n15249), .A2(n15248), .A3(n18665), .ZN(n15247) );
  OAI221_X1 U18360 ( .B1(n15250), .B2(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .C1(
        n15249), .C2(n15248), .A(n15247), .ZN(n17687) );
  NOR2_X1 U18361 ( .A1(n17688), .A2(n17687), .ZN(n17686) );
  NOR2_X1 U18362 ( .A1(n15251), .A2(n17686), .ZN(n17675) );
  XNOR2_X1 U18363 ( .A(n15252), .B(n17678), .ZN(n17674) );
  XOR2_X1 U18364 ( .A(n15255), .B(n15254), .Z(n17661) );
  NOR2_X1 U18365 ( .A1(n17660), .A2(n17661), .ZN(n15256) );
  NAND2_X1 U18366 ( .A1(n17660), .A2(n17661), .ZN(n17659) );
  OAI21_X1 U18367 ( .B1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n15256), .A(
        n17659), .ZN(n17652) );
  XOR2_X1 U18368 ( .A(n15259), .B(n15258), .Z(n15261) );
  NOR2_X1 U18369 ( .A1(n15260), .A2(n15261), .ZN(n15262) );
  INV_X1 U18370 ( .A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n20912) );
  XNOR2_X1 U18371 ( .A(n15261), .B(n15260), .ZN(n17638) );
  XNOR2_X1 U18372 ( .A(n15263), .B(n17193), .ZN(n15266) );
  NAND2_X1 U18373 ( .A1(n15265), .A2(n15266), .ZN(n17627) );
  NAND2_X1 U18374 ( .A1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(n17627), .ZN(
        n15268) );
  NOR2_X1 U18375 ( .A1(n15264), .A2(n15268), .ZN(n15270) );
  INV_X1 U18376 ( .A(n15264), .ZN(n15269) );
  OR2_X1 U18377 ( .A1(n15266), .A2(n15265), .ZN(n17628) );
  OAI21_X1 U18378 ( .B1(n15269), .B2(n15268), .A(n17628), .ZN(n15267) );
  AOI21_X1 U18379 ( .B1(n15269), .B2(n15268), .A(n15267), .ZN(n17613) );
  INV_X1 U18380 ( .A(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n17948) );
  NAND3_X1 U18381 ( .A1(n17887), .A2(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n17539) );
  NOR2_X2 U18382 ( .A1(n17539), .A2(n17845), .ZN(n17847) );
  NAND2_X1 U18383 ( .A1(n17847), .A2(n15271), .ZN(n17751) );
  NAND2_X1 U18384 ( .A1(n17395), .A2(n15274), .ZN(n17347) );
  NAND2_X1 U18385 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n15272) );
  NOR2_X1 U18386 ( .A1(n17347), .A2(n15272), .ZN(n16224) );
  NAND3_X1 U18387 ( .A1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n15273) );
  INV_X1 U18388 ( .A(n15273), .ZN(n17844) );
  NAND3_X1 U18389 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n17946) );
  NAND2_X1 U18390 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n17977) );
  NOR2_X1 U18391 ( .A1(n17946), .A2(n17977), .ZN(n17944) );
  NAND2_X1 U18392 ( .A1(n17844), .A2(n17944), .ZN(n17879) );
  NOR2_X1 U18393 ( .A1(n17820), .A2(n17879), .ZN(n17813) );
  NOR2_X1 U18394 ( .A1(n17485), .A2(n17766), .ZN(n17772) );
  NAND2_X1 U18395 ( .A1(n17813), .A2(n17772), .ZN(n17714) );
  OR2_X1 U18396 ( .A1(n17436), .A2(n17714), .ZN(n15278) );
  INV_X1 U18397 ( .A(n18509), .ZN(n18003) );
  INV_X1 U18398 ( .A(n17820), .ZN(n17833) );
  AOI21_X1 U18399 ( .B1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n18000) );
  NOR3_X1 U18400 ( .A1(n18000), .A2(n17946), .A3(n15273), .ZN(n17859) );
  NAND2_X1 U18401 ( .A1(n17833), .A2(n17859), .ZN(n17768) );
  NOR2_X1 U18402 ( .A1(n17485), .A2(n17768), .ZN(n17812) );
  NAND2_X1 U18403 ( .A1(n18003), .A2(n17812), .ZN(n16235) );
  INV_X1 U18404 ( .A(n16237), .ZN(n17412) );
  INV_X1 U18405 ( .A(n18510), .ZN(n17929) );
  NOR2_X1 U18406 ( .A1(n18665), .A2(n15278), .ZN(n17713) );
  INV_X1 U18407 ( .A(n17713), .ZN(n15277) );
  OAI222_X1 U18408 ( .A1(n18512), .A2(n15278), .B1(n16235), .B2(n17412), .C1(
        n17929), .C2(n15277), .ZN(n17736) );
  INV_X1 U18409 ( .A(n17736), .ZN(n15275) );
  INV_X1 U18410 ( .A(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n17711) );
  INV_X1 U18411 ( .A(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n17760) );
  NOR2_X1 U18412 ( .A1(n17760), .A2(n17748), .ZN(n17737) );
  NAND2_X1 U18413 ( .A1(n15274), .A2(n17737), .ZN(n17712) );
  OR2_X1 U18414 ( .A1(n17711), .A2(n17712), .ZN(n16238) );
  NOR4_X1 U18415 ( .A1(n15275), .A2(n18019), .A3(n17349), .A4(n16238), .ZN(
        n16203) );
  AOI21_X1 U18416 ( .B1(n17999), .B2(n16224), .A(n16203), .ZN(n15276) );
  OAI21_X1 U18417 ( .B1(n17938), .B2(n16227), .A(n15276), .ZN(n15395) );
  INV_X1 U18418 ( .A(n15395), .ZN(n15283) );
  NAND3_X1 U18419 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n15397) );
  OAI22_X1 U18420 ( .A1(n16187), .A2(n17938), .B1(n16198), .B2(n18033), .ZN(
        n15398) );
  NAND2_X1 U18421 ( .A1(n18013), .A2(n18019), .ZN(n18012) );
  NAND2_X1 U18422 ( .A1(n16237), .A2(n17812), .ZN(n17754) );
  OAI21_X1 U18423 ( .B1(n17754), .B2(n17712), .A(n18003), .ZN(n17716) );
  OAI21_X1 U18424 ( .B1(n15277), .B2(n16238), .A(n18510), .ZN(n15280) );
  INV_X1 U18425 ( .A(n18512), .ZN(n18499) );
  OAI21_X1 U18426 ( .B1(n17712), .B2(n15278), .A(n18499), .ZN(n15279) );
  NAND4_X1 U18427 ( .A1(n18012), .A2(n17716), .A3(n15280), .A4(n15279), .ZN(
        n15396) );
  AOI21_X1 U18428 ( .B1(n17919), .B2(n17711), .A(n15396), .ZN(n16223) );
  NOR2_X1 U18429 ( .A1(n17947), .A2(n18019), .ZN(n17979) );
  INV_X1 U18430 ( .A(n17979), .ZN(n18014) );
  OAI22_X1 U18431 ( .A1(n17971), .A2(n16223), .B1(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .B2(n18014), .ZN(n15281) );
  NOR2_X1 U18432 ( .A1(n15398), .A2(n15281), .ZN(n15282) );
  MUX2_X1 U18433 ( .A(n15283), .B(n15282), .S(
        P3_INSTADDRPOINTER_REG_29__SCAN_IN), .Z(n15284) );
  NAND2_X1 U18434 ( .A1(n17971), .A2(P3_REIP_REG_29__SCAN_IN), .ZN(n16193) );
  OAI211_X1 U18435 ( .C1(n16202), .C2(n17940), .A(n15284), .B(n16193), .ZN(
        P3_U2833) );
  INV_X1 U18436 ( .A(n15286), .ZN(n15287) );
  NAND2_X1 U18437 ( .A1(n15285), .A2(n15287), .ZN(n15288) );
  AND2_X1 U18438 ( .A1(n13708), .A2(n15288), .ZN(n18968) );
  INV_X1 U18439 ( .A(n15289), .ZN(n15292) );
  INV_X1 U18440 ( .A(n15290), .ZN(n15291) );
  NAND2_X1 U18441 ( .A1(n15292), .A2(n15291), .ZN(n15293) );
  AND2_X1 U18442 ( .A1(n15293), .A2(n9710), .ZN(n18943) );
  AOI22_X1 U18443 ( .A1(n18968), .A2(n19122), .B1(n19131), .B2(n18943), .ZN(
        n15304) );
  XOR2_X1 U18444 ( .A(n15295), .B(n15294), .Z(n16002) );
  INV_X1 U18445 ( .A(n15301), .ZN(n15297) );
  AOI21_X1 U18446 ( .B1(n15297), .B2(n15296), .A(n16103), .ZN(n16076) );
  INV_X1 U18447 ( .A(n16017), .ZN(n15298) );
  NAND2_X1 U18448 ( .A1(n15315), .A2(n15298), .ZN(n16003) );
  OAI21_X1 U18449 ( .B1(n16122), .B2(n19116), .A(n16003), .ZN(n15299) );
  OAI211_X1 U18450 ( .C1(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .C2(n15300), .A(
        n16076), .B(n15299), .ZN(n15316) );
  AOI22_X1 U18451 ( .A1(n16002), .A2(n12942), .B1(
        P2_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n15316), .ZN(n15303) );
  NAND2_X1 U18452 ( .A1(n15301), .A2(n16107), .ZN(n16077) );
  OAI21_X1 U18453 ( .B1(n16017), .B2(n19125), .A(n16077), .ZN(n15314) );
  NAND3_X1 U18454 ( .A1(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n15317), .A3(
        n15314), .ZN(n15302) );
  NAND2_X1 U18455 ( .A1(P2_REIP_REG_16__SCAN_IN), .A2(n18810), .ZN(n16005) );
  NAND4_X1 U18456 ( .A1(n15304), .A2(n15303), .A3(n15302), .A4(n16005), .ZN(
        P2_U3030) );
  AOI211_X1 U18457 ( .C1(n15985), .C2(n15305), .A(n9725), .B(n18890), .ZN(
        n15310) );
  INV_X1 U18458 ( .A(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n15308) );
  OAI222_X1 U18459 ( .A1(n18935), .A2(n15308), .B1(n18929), .B2(n15307), .C1(
        n18923), .C2(n15306), .ZN(n15309) );
  AOI211_X1 U18460 ( .C1(n18910), .C2(P2_REIP_REG_22__SCAN_IN), .A(n15310), 
        .B(n15309), .ZN(n15313) );
  INV_X1 U18461 ( .A(n15311), .ZN(n15950) );
  AOI22_X1 U18462 ( .A1(n15989), .A2(n18916), .B1(n18874), .B2(n15950), .ZN(
        n15312) );
  NAND2_X1 U18463 ( .A1(n15313), .A2(n15312), .ZN(P2_U2833) );
  NAND2_X1 U18464 ( .A1(n15315), .A2(n15314), .ZN(n15326) );
  AOI21_X1 U18465 ( .B1(n15317), .B2(n19132), .A(n15316), .ZN(n15325) );
  OAI21_X1 U18466 ( .B1(n15320), .B2(n15319), .A(n15318), .ZN(n15999) );
  INV_X1 U18467 ( .A(n18776), .ZN(n15321) );
  INV_X1 U18468 ( .A(P2_REIP_REG_17__SCAN_IN), .ZN(n19709) );
  NOR2_X1 U18469 ( .A1(n16114), .A2(n19709), .ZN(n15992) );
  AOI21_X1 U18470 ( .B1(n19131), .B2(n15321), .A(n15992), .ZN(n15322) );
  OAI21_X1 U18471 ( .B1(n18777), .B2(n16128), .A(n15322), .ZN(n15323) );
  AOI21_X1 U18472 ( .B1(n15999), .B2(n12942), .A(n15323), .ZN(n15324) );
  OAI221_X1 U18473 ( .B1(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n15326), 
        .C1(n15996), .C2(n15325), .A(n15324), .ZN(P2_U3029) );
  INV_X1 U18474 ( .A(n15409), .ZN(n15344) );
  NOR2_X1 U18475 ( .A1(n15344), .A2(n15368), .ZN(n15375) );
  INV_X1 U18476 ( .A(n15335), .ZN(n15337) );
  OAI211_X1 U18477 ( .C1(n9779), .C2(n15328), .A(n15327), .B(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n15329) );
  INV_X1 U18478 ( .A(n15329), .ZN(n15333) );
  AOI22_X1 U18479 ( .A1(n15331), .A2(n15330), .B1(n20697), .B2(n15329), .ZN(
        n15332) );
  AOI21_X1 U18480 ( .B1(n15333), .B2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A(
        n15332), .ZN(n15334) );
  OAI21_X1 U18481 ( .B1(n15335), .B2(n20326), .A(n15334), .ZN(n15336) );
  OAI21_X1 U18482 ( .B1(n15337), .B2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A(
        n15336), .ZN(n15338) );
  AOI222_X1 U18483 ( .A1(n15339), .A2(n15338), .B1(n15339), .B2(n20690), .C1(
        n15338), .C2(n20690), .ZN(n15359) );
  INV_X1 U18484 ( .A(n15340), .ZN(n15355) );
  INV_X1 U18485 ( .A(P1_MORE_REG_SCAN_IN), .ZN(n20719) );
  INV_X1 U18486 ( .A(n15348), .ZN(n15341) );
  AOI21_X1 U18487 ( .B1(n15349), .B2(n15341), .A(n11064), .ZN(n15342) );
  AOI21_X1 U18488 ( .B1(n15344), .B2(n15343), .A(n15342), .ZN(n19818) );
  OAI21_X1 U18489 ( .B1(n15345), .B2(n10249), .A(n20728), .ZN(n20723) );
  NAND2_X1 U18490 ( .A1(n19818), .A2(n20723), .ZN(n19825) );
  AOI21_X1 U18491 ( .B1(n19827), .B2(n20719), .A(n19825), .ZN(n15354) );
  AND2_X1 U18492 ( .A1(n15347), .A2(n15346), .ZN(n15353) );
  OR2_X1 U18493 ( .A1(n15349), .A2(n15348), .ZN(n15352) );
  NAND2_X1 U18494 ( .A1(n15409), .A2(n15350), .ZN(n15351) );
  OAI211_X1 U18495 ( .C1(n15409), .C2(n15353), .A(n15352), .B(n15351), .ZN(
        n20717) );
  NOR4_X1 U18496 ( .A1(n15356), .A2(n15355), .A3(n15354), .A4(n20717), .ZN(
        n15357) );
  OAI211_X1 U18497 ( .C1(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .C2(n15359), .A(
        n15358), .B(n15357), .ZN(n15370) );
  INV_X1 U18498 ( .A(n15370), .ZN(n15365) );
  NOR2_X1 U18499 ( .A1(n15360), .A2(n15405), .ZN(n15364) );
  NAND3_X1 U18500 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n20607), .A3(n20597), 
        .ZN(n15361) );
  AOI22_X1 U18501 ( .A1(n15364), .A2(n15363), .B1(n15362), .B2(n15361), .ZN(
        n15865) );
  OAI221_X1 U18502 ( .B1(P1_STATE2_REG_1__SCAN_IN), .B2(
        P1_STATE2_REG_0__SCAN_IN), .C1(P1_STATE2_REG_1__SCAN_IN), .C2(n15365), 
        .A(n15865), .ZN(n15871) );
  NAND2_X1 U18503 ( .A1(n15871), .A2(n20597), .ZN(n15374) );
  INV_X1 U18504 ( .A(n15366), .ZN(n15367) );
  NAND2_X1 U18505 ( .A1(n15367), .A2(n15412), .ZN(n20704) );
  OAI211_X1 U18506 ( .C1(P1_STATE2_REG_2__SCAN_IN), .C2(n20728), .A(n20704), 
        .B(n15368), .ZN(n15369) );
  AOI21_X1 U18507 ( .B1(n15371), .B2(n15370), .A(n15369), .ZN(n15372) );
  AND2_X1 U18508 ( .A1(n15871), .A2(n15372), .ZN(n15373) );
  OAI22_X1 U18509 ( .A1(n15375), .A2(n15374), .B1(n15373), .B2(n20597), .ZN(
        P1_U3161) );
  INV_X1 U18510 ( .A(n15376), .ZN(n20074) );
  INV_X1 U18511 ( .A(n15770), .ZN(n15377) );
  NAND2_X1 U18512 ( .A1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n15788), .ZN(
        n15772) );
  OAI22_X1 U18513 ( .A1(n20066), .A2(n15377), .B1(n20065), .B2(n15772), .ZN(
        n15774) );
  NAND2_X1 U18514 ( .A1(n15378), .A2(n15774), .ZN(n15729) );
  OAI21_X1 U18515 ( .B1(n20074), .B2(n15730), .A(n15729), .ZN(n15420) );
  NAND2_X1 U18516 ( .A1(n15379), .A2(n15420), .ZN(n15720) );
  AOI22_X1 U18517 ( .A1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n15719), .B1(
        n20043), .B2(P1_REIP_REG_21__SCAN_IN), .ZN(n15383) );
  AOI22_X1 U18518 ( .A1(n20064), .A2(n15381), .B1(n20078), .B2(n15380), .ZN(
        n15382) );
  OAI211_X1 U18519 ( .C1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .C2(n15720), .A(
        n15383), .B(n15382), .ZN(P1_U3010) );
  INV_X1 U18520 ( .A(n15676), .ZN(n15384) );
  OAI21_X1 U18521 ( .B1(n15672), .B2(n15384), .A(
        P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n15388) );
  NAND2_X1 U18522 ( .A1(n15386), .A2(n15385), .ZN(n15387) );
  AOI22_X1 U18523 ( .A1(n15389), .A2(n20064), .B1(n15388), .B2(n15387), .ZN(
        n15391) );
  OAI211_X1 U18524 ( .C1(n15392), .C2(n20070), .A(n15391), .B(n15390), .ZN(
        P1_U3001) );
  NOR2_X1 U18525 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n15397), .ZN(
        n16183) );
  AOI22_X1 U18526 ( .A1(n17971), .A2(P3_REIP_REG_30__SCAN_IN), .B1(n16183), 
        .B2(n15395), .ZN(n15401) );
  AOI22_X1 U18527 ( .A1(n17979), .A2(n15397), .B1(n18013), .B2(n15396), .ZN(
        n16206) );
  INV_X1 U18528 ( .A(n16206), .ZN(n15399) );
  OAI21_X1 U18529 ( .B1(n15399), .B2(n15398), .A(
        P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n15400) );
  OAI211_X1 U18530 ( .C1(n10126), .C2(n17940), .A(n15401), .B(n15400), .ZN(
        P3_U2832) );
  INV_X1 U18531 ( .A(HOLD), .ZN(n20601) );
  INV_X1 U18532 ( .A(P1_STATE_REG_2__SCAN_IN), .ZN(n20617) );
  NAND2_X1 U18533 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(n20617), .ZN(n20606) );
  INV_X1 U18534 ( .A(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n20608) );
  NOR2_X1 U18535 ( .A1(n20604), .A2(n20608), .ZN(n20611) );
  INV_X1 U18536 ( .A(P1_STATE_REG_1__SCAN_IN), .ZN(n20609) );
  NOR2_X1 U18537 ( .A1(n20609), .A2(n20728), .ZN(n15402) );
  AOI221_X1 U18538 ( .B1(n20601), .B2(n20611), .C1(n20617), .C2(n20611), .A(
        n15402), .ZN(n15403) );
  OAI211_X1 U18539 ( .C1(n20601), .C2(n20606), .A(n15403), .B(n15405), .ZN(
        P1_U3195) );
  INV_X1 U18540 ( .A(n15404), .ZN(n15407) );
  NOR2_X1 U18541 ( .A1(n10256), .A2(n15405), .ZN(n15406) );
  NAND2_X1 U18542 ( .A1(n15407), .A2(n15406), .ZN(n15411) );
  NAND3_X1 U18543 ( .A1(n15409), .A2(n19826), .A3(n15408), .ZN(n15410) );
  INV_X1 U18544 ( .A(n15412), .ZN(n15866) );
  OR2_X1 U18545 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n15866), .ZN(n19967) );
  INV_X2 U18546 ( .A(n19967), .ZN(n20729) );
  NOR2_X4 U18547 ( .A1(n19947), .A2(n20729), .ZN(n19970) );
  AND2_X1 U18548 ( .A1(n19970), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(P1_U2905)
         );
  NAND2_X1 U18549 ( .A1(n15414), .A2(n15413), .ZN(n15416) );
  OAI21_X1 U18550 ( .B1(n15599), .B2(n15416), .A(n15415), .ZN(n15417) );
  XNOR2_X1 U18551 ( .A(n15417), .B(n15419), .ZN(n15594) );
  AOI22_X1 U18552 ( .A1(n20064), .A2(n15508), .B1(n20078), .B2(n15594), .ZN(
        n15423) );
  AOI21_X1 U18553 ( .B1(n20074), .B2(n15729), .A(
        P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n15732) );
  INV_X1 U18554 ( .A(n15418), .ZN(n15728) );
  OAI21_X1 U18555 ( .B1(n15732), .B2(n15728), .A(
        P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n15422) );
  NAND2_X1 U18556 ( .A1(n20043), .A2(P1_REIP_REG_20__SCAN_IN), .ZN(n15595) );
  NAND3_X1 U18557 ( .A1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n15420), .A3(
        n15419), .ZN(n15421) );
  NAND4_X1 U18558 ( .A1(n15423), .A2(n15422), .A3(n15595), .A4(n15421), .ZN(
        P1_U3011) );
  NOR3_X1 U18559 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n18715), .A3(n15424), 
        .ZN(n16146) );
  NOR2_X1 U18560 ( .A1(n15425), .A2(n16146), .ZN(n19665) );
  INV_X1 U18561 ( .A(n19665), .ZN(n15426) );
  AOI211_X1 U18562 ( .C1(n19801), .C2(n13649), .A(n16147), .B(n15426), .ZN(
        P2_U3178) );
  INV_X1 U18563 ( .A(n19792), .ZN(n15427) );
  AOI221_X1 U18564 ( .B1(P2_FLUSH_REG_SCAN_IN), .B2(n16147), .C1(n15427), .C2(
        n16147), .A(n19593), .ZN(n19774) );
  INV_X1 U18565 ( .A(n19774), .ZN(n19784) );
  NOR2_X1 U18566 ( .A1(n15428), .A2(n19784), .ZN(P2_U3047) );
  NAND3_X1 U18567 ( .A1(n18047), .A2(n18692), .A3(n15429), .ZN(n15430) );
  NAND2_X1 U18568 ( .A1(n18087), .A2(n17186), .ZN(n17211) );
  INV_X1 U18569 ( .A(P3_EAX_REG_0__SCAN_IN), .ZN(n17288) );
  NAND2_X2 U18570 ( .A1(n17186), .A2(n17123), .ZN(n17213) );
  AOI22_X1 U18571 ( .A1(n17222), .A2(BUF2_REG_0__SCAN_IN), .B1(n17221), .B2(
        n17706), .ZN(n15432) );
  OAI221_X1 U18572 ( .B1(P3_EAX_REG_0__SCAN_IN), .B2(n17211), .C1(n17288), 
        .C2(n17186), .A(n15432), .ZN(P3_U2735) );
  OAI21_X1 U18573 ( .B1(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A(n15433), .ZN(n15443) );
  INV_X1 U18574 ( .A(n15434), .ZN(n15442) );
  OR2_X1 U18575 ( .A1(n15436), .A2(n15435), .ZN(n15441) );
  AOI21_X1 U18576 ( .B1(n15438), .B2(n15437), .A(n9656), .ZN(n18750) );
  AOI21_X1 U18577 ( .B1(n19122), .B2(n18750), .A(n15439), .ZN(n15440) );
  OAI211_X1 U18578 ( .C1(n15443), .C2(n15442), .A(n15441), .B(n15440), .ZN(
        n15444) );
  INV_X1 U18579 ( .A(n15444), .ZN(n15448) );
  AOI22_X1 U18580 ( .A1(n15446), .A2(n16122), .B1(n19131), .B2(n18751), .ZN(
        n15447) );
  OAI211_X1 U18581 ( .C1(n19110), .C2(n15449), .A(n15448), .B(n15447), .ZN(
        P2_U3026) );
  NOR2_X1 U18582 ( .A1(n15680), .A2(n19931), .ZN(n15458) );
  INV_X1 U18583 ( .A(P1_REIP_REG_28__SCAN_IN), .ZN(n15455) );
  AND3_X1 U18584 ( .A1(n19920), .A2(n15451), .A3(n15450), .ZN(n15452) );
  AOI21_X1 U18585 ( .B1(P1_EBX_REG_28__SCAN_IN), .B2(n19929), .A(n15452), .ZN(
        n15454) );
  NAND2_X1 U18586 ( .A1(n19935), .A2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n15453) );
  OAI211_X1 U18587 ( .C1(n15456), .C2(n15455), .A(n15454), .B(n15453), .ZN(
        n15457) );
  AOI211_X1 U18588 ( .C1(n15563), .C2(n19872), .A(n15458), .B(n15457), .ZN(
        n15459) );
  OAI21_X1 U18589 ( .B1(n15566), .B2(n19897), .A(n15459), .ZN(P1_U2812) );
  INV_X1 U18590 ( .A(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n15467) );
  INV_X1 U18591 ( .A(n15460), .ZN(n15463) );
  OAI21_X1 U18592 ( .B1(n15461), .B2(n19875), .A(n20660), .ZN(n15462) );
  AOI22_X1 U18593 ( .A1(n15463), .A2(n15462), .B1(n19929), .B2(
        P1_EBX_REG_26__SCAN_IN), .ZN(n15466) );
  OAI22_X1 U18594 ( .A1(n15694), .A2(n19931), .B1(n15575), .B2(n19897), .ZN(
        n15464) );
  AOI21_X1 U18595 ( .B1(n15572), .B2(n19872), .A(n15464), .ZN(n15465) );
  OAI211_X1 U18596 ( .C1(n15467), .C2(n19923), .A(n15466), .B(n15465), .ZN(
        P1_U2814) );
  AOI22_X1 U18597 ( .A1(n19935), .A2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .B1(
        P1_EBX_REG_25__SCAN_IN), .B2(n19929), .ZN(n15478) );
  OAI22_X1 U18598 ( .A1(n15468), .A2(n19861), .B1(n19931), .B2(n15700), .ZN(
        n15469) );
  AOI21_X1 U18599 ( .B1(n15470), .B2(n19934), .A(n15469), .ZN(n15477) );
  AOI21_X1 U18600 ( .B1(n15473), .B2(n15472), .A(n15471), .ZN(n15489) );
  NOR2_X1 U18601 ( .A1(P1_REIP_REG_24__SCAN_IN), .A2(n19875), .ZN(n15481) );
  OAI21_X1 U18602 ( .B1(n15489), .B2(n15481), .A(P1_REIP_REG_25__SCAN_IN), 
        .ZN(n15476) );
  INV_X1 U18603 ( .A(P1_REIP_REG_25__SCAN_IN), .ZN(n20657) );
  NAND3_X1 U18604 ( .A1(n19920), .A2(n15474), .A3(n20657), .ZN(n15475) );
  NAND4_X1 U18605 ( .A1(n15478), .A2(n15477), .A3(n15476), .A4(n15475), .ZN(
        P1_U2815) );
  INV_X1 U18606 ( .A(n15479), .ZN(n15580) );
  INV_X1 U18607 ( .A(n15480), .ZN(n15482) );
  AOI22_X1 U18608 ( .A1(P1_REIP_REG_24__SCAN_IN), .A2(n15489), .B1(n15482), 
        .B2(n15481), .ZN(n15484) );
  AOI22_X1 U18609 ( .A1(n19935), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .B1(
        n19929), .B2(P1_EBX_REG_24__SCAN_IN), .ZN(n15483) );
  OAI211_X1 U18610 ( .C1(n19931), .C2(n15709), .A(n15484), .B(n15483), .ZN(
        n15485) );
  AOI21_X1 U18611 ( .B1(n15580), .B2(n19872), .A(n15485), .ZN(n15486) );
  OAI21_X1 U18612 ( .B1(n15583), .B2(n19897), .A(n15486), .ZN(P1_U2816) );
  AOI22_X1 U18613 ( .A1(n19934), .A2(n15487), .B1(P1_EBX_REG_23__SCAN_IN), 
        .B2(n19929), .ZN(n15495) );
  AOI21_X1 U18614 ( .B1(P1_REIP_REG_22__SCAN_IN), .B2(n15488), .A(
        P1_REIP_REG_23__SCAN_IN), .ZN(n15491) );
  INV_X1 U18615 ( .A(n15489), .ZN(n15490) );
  OAI22_X1 U18616 ( .A1(n15491), .A2(n15490), .B1(n19931), .B2(n15712), .ZN(
        n15492) );
  AOI21_X1 U18617 ( .B1(n15493), .B2(n19872), .A(n15492), .ZN(n15494) );
  OAI211_X1 U18618 ( .C1(n15496), .C2(n19923), .A(n15495), .B(n15494), .ZN(
        P1_U2817) );
  AOI22_X1 U18619 ( .A1(n19934), .A2(n15497), .B1(n19929), .B2(
        P1_EBX_REG_21__SCAN_IN), .ZN(n15505) );
  NAND2_X1 U18620 ( .A1(n15498), .A2(n20650), .ZN(n15502) );
  OAI22_X1 U18621 ( .A1(n15500), .A2(n19861), .B1(n19931), .B2(n15499), .ZN(
        n15501) );
  AOI21_X1 U18622 ( .B1(n15503), .B2(n15502), .A(n15501), .ZN(n15504) );
  OAI211_X1 U18623 ( .C1(n15506), .C2(n19923), .A(n15505), .B(n15504), .ZN(
        P1_U2819) );
  AOI22_X1 U18624 ( .A1(n19935), .A2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .B1(
        n19929), .B2(P1_EBX_REG_20__SCAN_IN), .ZN(n15515) );
  INV_X1 U18625 ( .A(n15592), .ZN(n15513) );
  NOR2_X1 U18626 ( .A1(P1_REIP_REG_20__SCAN_IN), .A2(n15507), .ZN(n15511) );
  INV_X1 U18627 ( .A(n15508), .ZN(n15509) );
  OAI22_X1 U18628 ( .A1(n15511), .A2(n15510), .B1(n15509), .B2(n19931), .ZN(
        n15512) );
  AOI21_X1 U18629 ( .B1(n15513), .B2(n19872), .A(n15512), .ZN(n15514) );
  OAI211_X1 U18630 ( .C1(n15591), .C2(n19897), .A(n15515), .B(n15514), .ZN(
        P1_U2820) );
  NAND2_X1 U18631 ( .A1(n15516), .A2(P1_REIP_REG_18__SCAN_IN), .ZN(n15520) );
  OAI21_X1 U18632 ( .B1(n19867), .B2(n10931), .A(n19879), .ZN(n15517) );
  INV_X1 U18633 ( .A(n15517), .ZN(n15519) );
  AOI22_X1 U18634 ( .A1(n15741), .A2(n19905), .B1(
        P1_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n19935), .ZN(n15518) );
  NAND3_X1 U18635 ( .A1(n15520), .A2(n15519), .A3(n15518), .ZN(n15521) );
  NOR2_X1 U18636 ( .A1(n15522), .A2(n15521), .ZN(n15523) );
  OAI21_X1 U18637 ( .B1(n15601), .B2(n19861), .A(n15523), .ZN(n15524) );
  INV_X1 U18638 ( .A(n15524), .ZN(n15525) );
  OAI21_X1 U18639 ( .B1(n15605), .B2(n19897), .A(n15525), .ZN(P1_U2822) );
  AOI22_X1 U18640 ( .A1(n15526), .A2(P1_REIP_REG_16__SCAN_IN), .B1(n19929), 
        .B2(P1_EBX_REG_16__SCAN_IN), .ZN(n15527) );
  OAI21_X1 U18641 ( .B1(P1_REIP_REG_16__SCAN_IN), .B2(n15528), .A(n15527), 
        .ZN(n15529) );
  AOI211_X1 U18642 ( .C1(n19935), .C2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .A(
        n19891), .B(n15529), .ZN(n15533) );
  XNOR2_X1 U18643 ( .A(n15531), .B(n15530), .ZN(n15760) );
  AOI22_X1 U18644 ( .A1(n15612), .A2(n19872), .B1(n19905), .B2(n15760), .ZN(
        n15532) );
  OAI211_X1 U18645 ( .C1(n15610), .C2(n19897), .A(n15533), .B(n15532), .ZN(
        P1_U2824) );
  OAI22_X1 U18646 ( .A1(n15810), .A2(n19931), .B1(n15534), .B2(n19867), .ZN(
        n15535) );
  AOI211_X1 U18647 ( .C1(n19935), .C2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .A(
        n19891), .B(n15535), .ZN(n15542) );
  INV_X1 U18648 ( .A(n15536), .ZN(n15633) );
  AOI22_X1 U18649 ( .A1(n15634), .A2(n19934), .B1(n19872), .B2(n15633), .ZN(
        n15541) );
  NAND3_X1 U18650 ( .A1(n19920), .A2(P1_REIP_REG_8__SCAN_IN), .A3(n15537), 
        .ZN(n19844) );
  NOR2_X1 U18651 ( .A1(n15538), .A2(n19844), .ZN(n15550) );
  OAI221_X1 U18652 ( .B1(P1_REIP_REG_12__SCAN_IN), .B2(P1_REIP_REG_11__SCAN_IN), .C1(P1_REIP_REG_12__SCAN_IN), .C2(n15550), .A(n15539), .ZN(n15540) );
  NAND3_X1 U18653 ( .A1(n15542), .A2(n15541), .A3(n15540), .ZN(P1_U2828) );
  INV_X1 U18654 ( .A(P1_REIP_REG_11__SCAN_IN), .ZN(n20635) );
  INV_X1 U18655 ( .A(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n15548) );
  NOR2_X1 U18656 ( .A1(n15544), .A2(n15543), .ZN(n15545) );
  AOI22_X1 U18657 ( .A1(n9700), .A2(n19905), .B1(n19929), .B2(
        P1_EBX_REG_11__SCAN_IN), .ZN(n15547) );
  OAI211_X1 U18658 ( .C1(n19923), .C2(n15548), .A(n15547), .B(n19879), .ZN(
        n15549) );
  AOI221_X1 U18659 ( .B1(n15551), .B2(P1_REIP_REG_11__SCAN_IN), .C1(n15550), 
        .C2(n20635), .A(n15549), .ZN(n15553) );
  NAND2_X1 U18660 ( .A1(n19872), .A2(n15644), .ZN(n15552) );
  OAI211_X1 U18661 ( .C1(n19897), .C2(n15648), .A(n15553), .B(n15552), .ZN(
        P1_U2829) );
  AOI22_X1 U18662 ( .A1(n15612), .A2(n19941), .B1(n19940), .B2(n15760), .ZN(
        n15554) );
  OAI21_X1 U18663 ( .B1(n19945), .B2(n15555), .A(n15554), .ZN(P1_U2856) );
  AOI22_X1 U18664 ( .A1(n15644), .A2(n19941), .B1(n19940), .B2(n9700), .ZN(
        n15556) );
  OAI21_X1 U18665 ( .B1(n19945), .B2(n15557), .A(n15556), .ZN(P1_U2861) );
  AOI22_X1 U18666 ( .A1(n20034), .A2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .B1(
        n20043), .B2(P1_REIP_REG_28__SCAN_IN), .ZN(n15565) );
  NAND2_X1 U18667 ( .A1(n15569), .A2(n15558), .ZN(n15567) );
  NOR3_X1 U18668 ( .A1(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n15560) );
  OAI221_X1 U18669 ( .B1(n15640), .B2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), 
        .C1(n15569), .C2(n11193), .A(n15561), .ZN(n15562) );
  XOR2_X1 U18670 ( .A(n12892), .B(n15562), .Z(n15677) );
  AOI22_X1 U18671 ( .A1(n15563), .A2(n15645), .B1(n20042), .B2(n15677), .ZN(
        n15564) );
  OAI211_X1 U18672 ( .C1(n20032), .C2(n15566), .A(n15565), .B(n15564), .ZN(
        P1_U2971) );
  AOI22_X1 U18673 ( .A1(n20034), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .B1(
        n20043), .B2(P1_REIP_REG_26__SCAN_IN), .ZN(n15574) );
  OAI211_X1 U18674 ( .C1(n15570), .C2(n15569), .A(n15568), .B(n15567), .ZN(
        n15571) );
  XNOR2_X1 U18675 ( .A(n15571), .B(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n15687) );
  AOI22_X1 U18676 ( .A1(n15572), .A2(n15645), .B1(n20042), .B2(n15687), .ZN(
        n15573) );
  OAI211_X1 U18677 ( .C1(n20032), .C2(n15575), .A(n15574), .B(n15573), .ZN(
        P1_U2973) );
  AOI22_X1 U18678 ( .A1(n20034), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .B1(
        n20043), .B2(P1_REIP_REG_24__SCAN_IN), .ZN(n15582) );
  AOI21_X1 U18679 ( .B1(n14468), .B2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n15640), .ZN(n15576) );
  OR2_X1 U18680 ( .A1(n14476), .A2(n15576), .ZN(n15579) );
  MUX2_X1 U18681 ( .A(n15577), .B(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .S(
        n15569), .Z(n15578) );
  XNOR2_X1 U18682 ( .A(n15579), .B(n15578), .ZN(n15705) );
  AOI22_X1 U18683 ( .A1(n15580), .A2(n15645), .B1(n20042), .B2(n15705), .ZN(
        n15581) );
  OAI211_X1 U18684 ( .C1(n20032), .C2(n15583), .A(n15582), .B(n15581), .ZN(
        P1_U2975) );
  AOI22_X1 U18685 ( .A1(n20034), .A2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .B1(
        n20043), .B2(P1_REIP_REG_22__SCAN_IN), .ZN(n15589) );
  NAND2_X1 U18686 ( .A1(n15585), .A2(n15584), .ZN(n15586) );
  XNOR2_X1 U18687 ( .A(n15586), .B(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n15724) );
  AOI22_X1 U18688 ( .A1(n15587), .A2(n15645), .B1(n20042), .B2(n15724), .ZN(
        n15588) );
  OAI211_X1 U18689 ( .C1(n20032), .C2(n15590), .A(n15589), .B(n15588), .ZN(
        P1_U2977) );
  INV_X1 U18690 ( .A(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n15597) );
  OAI22_X1 U18691 ( .A1(n15592), .A2(n20084), .B1(n15591), .B2(n20032), .ZN(
        n15593) );
  AOI21_X1 U18692 ( .B1(n20042), .B2(n15594), .A(n15593), .ZN(n15596) );
  OAI211_X1 U18693 ( .C1(n15597), .C2(n20039), .A(n15596), .B(n15595), .ZN(
        P1_U2979) );
  AOI22_X1 U18694 ( .A1(n20034), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .B1(
        n20043), .B2(P1_REIP_REG_18__SCAN_IN), .ZN(n15604) );
  OR2_X1 U18695 ( .A1(n15599), .A2(n15598), .ZN(n15600) );
  NAND2_X1 U18696 ( .A1(n14486), .A2(n15600), .ZN(n15745) );
  OAI22_X1 U18697 ( .A1(n15601), .A2(n20084), .B1(n20031), .B2(n15745), .ZN(
        n15602) );
  INV_X1 U18698 ( .A(n15602), .ZN(n15603) );
  OAI211_X1 U18699 ( .C1(n20032), .C2(n15605), .A(n15604), .B(n15603), .ZN(
        P1_U2981) );
  NOR2_X1 U18700 ( .A1(n15757), .A2(n15607), .ZN(n15608) );
  OAI22_X1 U18701 ( .A1(n15609), .A2(n15608), .B1(n15607), .B2(n15606), .ZN(
        n15763) );
  AOI22_X1 U18702 ( .A1(n20034), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .B1(
        n20043), .B2(P1_REIP_REG_16__SCAN_IN), .ZN(n15614) );
  INV_X1 U18703 ( .A(n15610), .ZN(n15611) );
  AOI22_X1 U18704 ( .A1(n15612), .A2(n15645), .B1(n15611), .B2(n15635), .ZN(
        n15613) );
  OAI211_X1 U18705 ( .C1(n20031), .C2(n15763), .A(n15614), .B(n15613), .ZN(
        P1_U2983) );
  NAND2_X1 U18706 ( .A1(n15638), .A2(n15615), .ZN(n15619) );
  INV_X1 U18707 ( .A(n15616), .ZN(n15617) );
  AOI21_X1 U18708 ( .B1(n15619), .B2(n15618), .A(n15617), .ZN(n15623) );
  AOI22_X1 U18709 ( .A1(n15640), .A2(n15778), .B1(
        P1_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n15569), .ZN(n15622) );
  XNOR2_X1 U18710 ( .A(n15623), .B(n15622), .ZN(n15782) );
  AOI22_X1 U18711 ( .A1(n20034), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .B1(
        n20043), .B2(P1_REIP_REG_14__SCAN_IN), .ZN(n15628) );
  INV_X1 U18712 ( .A(n15624), .ZN(n15626) );
  AOI22_X1 U18713 ( .A1(n15626), .A2(n15645), .B1(n15635), .B2(n15625), .ZN(
        n15627) );
  OAI211_X1 U18714 ( .C1(n15782), .C2(n20031), .A(n15628), .B(n15627), .ZN(
        P1_U2985) );
  NOR2_X1 U18715 ( .A1(n15630), .A2(n15629), .ZN(n15631) );
  NOR2_X1 U18716 ( .A1(n15632), .A2(n15631), .ZN(n15805) );
  AOI22_X1 U18717 ( .A1(n20034), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B1(
        n20043), .B2(P1_REIP_REG_12__SCAN_IN), .ZN(n15637) );
  AOI22_X1 U18718 ( .A1(n15635), .A2(n15634), .B1(n15645), .B2(n15633), .ZN(
        n15636) );
  OAI211_X1 U18719 ( .C1(n15805), .C2(n20031), .A(n15637), .B(n15636), .ZN(
        P1_U2987) );
  AOI22_X1 U18720 ( .A1(n20034), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .B1(
        n20043), .B2(P1_REIP_REG_11__SCAN_IN), .ZN(n15647) );
  NOR2_X1 U18721 ( .A1(n15638), .A2(n11184), .ZN(n15642) );
  NOR2_X1 U18722 ( .A1(n15639), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n15641) );
  MUX2_X1 U18723 ( .A(n15642), .B(n15641), .S(n15640), .Z(n15643) );
  INV_X1 U18724 ( .A(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n15795) );
  XNOR2_X1 U18725 ( .A(n15643), .B(n15795), .ZN(n15812) );
  AOI22_X1 U18726 ( .A1(n20042), .A2(n15812), .B1(n15645), .B2(n15644), .ZN(
        n15646) );
  OAI211_X1 U18727 ( .C1(n20032), .C2(n15648), .A(n15647), .B(n15646), .ZN(
        P1_U2988) );
  AOI22_X1 U18728 ( .A1(n20034), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .B1(
        n20043), .B2(P1_REIP_REG_7__SCAN_IN), .ZN(n15654) );
  XNOR2_X1 U18729 ( .A(n15649), .B(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n15651) );
  XNOR2_X1 U18730 ( .A(n15651), .B(n15650), .ZN(n15844) );
  INV_X1 U18731 ( .A(n19862), .ZN(n15652) );
  AOI22_X1 U18732 ( .A1(n15844), .A2(n20042), .B1(n15652), .B2(n15645), .ZN(
        n15653) );
  OAI211_X1 U18733 ( .C1(n20032), .C2(n19854), .A(n15654), .B(n15653), .ZN(
        P1_U2992) );
  AOI22_X1 U18734 ( .A1(n20034), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .B1(
        n20043), .B2(P1_REIP_REG_6__SCAN_IN), .ZN(n15659) );
  NAND2_X1 U18735 ( .A1(n15656), .A2(n15655), .ZN(n15657) );
  AOI22_X1 U18736 ( .A1(n15852), .A2(n20042), .B1(n15645), .B2(n19942), .ZN(
        n15658) );
  OAI211_X1 U18737 ( .C1(n20032), .C2(n19874), .A(n15659), .B(n15658), .ZN(
        P1_U2993) );
  OAI222_X1 U18738 ( .A1(n15660), .A2(n20031), .B1(n19885), .B2(n20084), .C1(
        n20032), .C2(n19889), .ZN(n15661) );
  INV_X1 U18739 ( .A(n15661), .ZN(n15663) );
  OAI211_X1 U18740 ( .C1(n15664), .C2(n20039), .A(n15663), .B(n15662), .ZN(
        P1_U2994) );
  NOR2_X1 U18741 ( .A1(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(n15665), .ZN(
        n15671) );
  NAND2_X1 U18742 ( .A1(n20043), .A2(P1_REIP_REG_29__SCAN_IN), .ZN(n15669) );
  OAI211_X1 U18743 ( .C1(n15672), .C2(n15671), .A(n15670), .B(n15669), .ZN(
        P1_U3002) );
  AOI21_X1 U18744 ( .B1(n12892), .B2(n11193), .A(n15681), .ZN(n15674) );
  AOI22_X1 U18745 ( .A1(P1_REIP_REG_28__SCAN_IN), .A2(n20043), .B1(n15674), 
        .B2(n15673), .ZN(n15679) );
  AND2_X1 U18746 ( .A1(n15676), .A2(n15675), .ZN(n15683) );
  AOI22_X1 U18747 ( .A1(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n15683), .B1(
        n20078), .B2(n15677), .ZN(n15678) );
  OAI211_X1 U18748 ( .C1(n20081), .C2(n15680), .A(n15679), .B(n15678), .ZN(
        P1_U3003) );
  INV_X1 U18749 ( .A(n15681), .ZN(n15682) );
  AOI22_X1 U18750 ( .A1(P1_REIP_REG_27__SCAN_IN), .A2(n20043), .B1(n15682), 
        .B2(n11193), .ZN(n15685) );
  OAI211_X1 U18751 ( .C1(n20081), .C2(n15686), .A(n15685), .B(n15684), .ZN(
        P1_U3004) );
  AOI22_X1 U18752 ( .A1(n20043), .A2(P1_REIP_REG_26__SCAN_IN), .B1(n20078), 
        .B2(n15687), .ZN(n15693) );
  NOR3_X1 U18753 ( .A1(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(n15688), .A3(
        n15701), .ZN(n15695) );
  INV_X1 U18754 ( .A(n15689), .ZN(n15690) );
  OAI22_X1 U18755 ( .A1(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n15691), .B1(
        n15695), .B2(n15690), .ZN(n15692) );
  OAI211_X1 U18756 ( .C1(n20081), .C2(n15694), .A(n15693), .B(n15692), .ZN(
        P1_U3005) );
  AOI21_X1 U18757 ( .B1(P1_REIP_REG_25__SCAN_IN), .B2(n20043), .A(n15695), 
        .ZN(n15699) );
  AOI22_X1 U18758 ( .A1(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(n15697), .B1(
        n20078), .B2(n15696), .ZN(n15698) );
  OAI211_X1 U18759 ( .C1(n20081), .C2(n15700), .A(n15699), .B(n15698), .ZN(
        P1_U3006) );
  NOR3_X1 U18760 ( .A1(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n15717), .A3(
        n15701), .ZN(n15702) );
  AOI21_X1 U18761 ( .B1(P1_REIP_REG_24__SCAN_IN), .B2(n20043), .A(n15702), 
        .ZN(n15708) );
  OAI21_X1 U18762 ( .B1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n15704), .A(
        n15703), .ZN(n15706) );
  AOI22_X1 U18763 ( .A1(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n15706), .B1(
        n20078), .B2(n15705), .ZN(n15707) );
  OAI211_X1 U18764 ( .C1(n20081), .C2(n15709), .A(n15708), .B(n15707), .ZN(
        P1_U3007) );
  AOI22_X1 U18765 ( .A1(P1_REIP_REG_23__SCAN_IN), .A2(n20043), .B1(n15710), 
        .B2(n15717), .ZN(n15716) );
  INV_X1 U18766 ( .A(n15711), .ZN(n15714) );
  INV_X1 U18767 ( .A(n15712), .ZN(n15713) );
  AOI22_X1 U18768 ( .A1(n15714), .A2(n20078), .B1(n20064), .B2(n15713), .ZN(
        n15715) );
  OAI211_X1 U18769 ( .C1(n15718), .C2(n15717), .A(n15716), .B(n15715), .ZN(
        P1_U3008) );
  AOI22_X1 U18770 ( .A1(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n15719), .B1(
        n20043), .B2(P1_REIP_REG_22__SCAN_IN), .ZN(n15726) );
  INV_X1 U18771 ( .A(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n15721) );
  AOI21_X1 U18772 ( .B1(n10035), .B2(n15721), .A(n15720), .ZN(n15723) );
  AOI22_X1 U18773 ( .A1(n15724), .A2(n20078), .B1(n15723), .B2(n15722), .ZN(
        n15725) );
  OAI211_X1 U18774 ( .C1(n20081), .C2(n15727), .A(n15726), .B(n15725), .ZN(
        P1_U3009) );
  AOI22_X1 U18775 ( .A1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n15728), .B1(
        n20043), .B2(P1_REIP_REG_19__SCAN_IN), .ZN(n15735) );
  NAND2_X1 U18776 ( .A1(n15730), .A2(n15729), .ZN(n15731) );
  AOI22_X1 U18777 ( .A1(n20078), .A2(n15733), .B1(n15732), .B2(n15731), .ZN(
        n15734) );
  OAI211_X1 U18778 ( .C1(n20081), .C2(n15736), .A(n15735), .B(n15734), .ZN(
        P1_U3012) );
  OAI21_X1 U18779 ( .B1(n15778), .B2(n15737), .A(n15834), .ZN(n15738) );
  OAI211_X1 U18780 ( .C1(n15819), .C2(n15783), .A(n15739), .B(n15738), .ZN(
        n15764) );
  AOI21_X1 U18781 ( .B1(n15834), .B2(n15743), .A(n15764), .ZN(n15755) );
  NAND2_X1 U18782 ( .A1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n15740), .ZN(
        n15769) );
  INV_X1 U18783 ( .A(n15769), .ZN(n15759) );
  NAND2_X1 U18784 ( .A1(n15759), .A2(n15749), .ZN(n15744) );
  INV_X1 U18785 ( .A(n15741), .ZN(n15742) );
  OAI222_X1 U18786 ( .A1(n15745), .A2(n20070), .B1(n15744), .B2(n15743), .C1(
        n20081), .C2(n15742), .ZN(n15746) );
  INV_X1 U18787 ( .A(n15746), .ZN(n15748) );
  NAND2_X1 U18788 ( .A1(n20043), .A2(P1_REIP_REG_18__SCAN_IN), .ZN(n15747) );
  OAI211_X1 U18789 ( .C1(n15755), .C2(n15749), .A(n15748), .B(n15747), .ZN(
        P1_U3013) );
  AOI21_X1 U18790 ( .B1(n15756), .B2(n15759), .A(
        P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n15754) );
  AOI22_X1 U18791 ( .A1(n20064), .A2(n15751), .B1(n20078), .B2(n15750), .ZN(
        n15753) );
  NAND2_X1 U18792 ( .A1(n20043), .A2(P1_REIP_REG_17__SCAN_IN), .ZN(n15752) );
  OAI211_X1 U18793 ( .C1(n15755), .C2(n15754), .A(n15753), .B(n15752), .ZN(
        P1_U3014) );
  AOI22_X1 U18794 ( .A1(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n15764), .B1(
        n20043), .B2(P1_REIP_REG_16__SCAN_IN), .ZN(n15762) );
  NOR2_X1 U18795 ( .A1(n15757), .A2(n15756), .ZN(n15758) );
  AOI22_X1 U18796 ( .A1(n20064), .A2(n15760), .B1(n15759), .B2(n15758), .ZN(
        n15761) );
  OAI211_X1 U18797 ( .C1(n20070), .C2(n15763), .A(n15762), .B(n15761), .ZN(
        P1_U3015) );
  AOI22_X1 U18798 ( .A1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n15764), .B1(
        n20043), .B2(P1_REIP_REG_15__SCAN_IN), .ZN(n15768) );
  AOI22_X1 U18799 ( .A1(n20064), .A2(n15766), .B1(n20078), .B2(n15765), .ZN(
        n15767) );
  OAI211_X1 U18800 ( .C1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .C2(n15769), .A(
        n15768), .B(n15767), .ZN(P1_U3016) );
  NOR2_X1 U18801 ( .A1(n20050), .A2(n20637), .ZN(n15776) );
  INV_X1 U18802 ( .A(n20073), .ZN(n20067) );
  OAI22_X1 U18803 ( .A1(n15770), .A2(n20066), .B1(n15783), .B2(n20074), .ZN(
        n15771) );
  AOI211_X1 U18804 ( .C1(n15773), .C2(n15772), .A(n20067), .B(n15771), .ZN(
        n15794) );
  NAND2_X1 U18805 ( .A1(n15793), .A2(n15774), .ZN(n15784) );
  AOI21_X1 U18806 ( .B1(n15794), .B2(n15784), .A(n15778), .ZN(n15775) );
  AOI211_X1 U18807 ( .C1(n20064), .C2(n15777), .A(n15776), .B(n15775), .ZN(
        n15781) );
  NAND3_X1 U18808 ( .A1(n15779), .A2(n15778), .A3(n15811), .ZN(n15780) );
  OAI211_X1 U18809 ( .C1(n15782), .C2(n20070), .A(n15781), .B(n15780), .ZN(
        P1_U3017) );
  NOR2_X1 U18810 ( .A1(n15783), .A2(n20074), .ZN(n15787) );
  INV_X1 U18811 ( .A(P1_REIP_REG_13__SCAN_IN), .ZN(n20639) );
  NOR2_X1 U18812 ( .A1(n20050), .A2(n20639), .ZN(n15786) );
  INV_X1 U18813 ( .A(n15784), .ZN(n15785) );
  AOI211_X1 U18814 ( .C1(n15788), .C2(n15787), .A(n15786), .B(n15785), .ZN(
        n15792) );
  AOI22_X1 U18815 ( .A1(n20064), .A2(n15790), .B1(n20078), .B2(n15789), .ZN(
        n15791) );
  OAI211_X1 U18816 ( .C1(n15794), .C2(n15793), .A(n15792), .B(n15791), .ZN(
        P1_U3018) );
  NOR2_X1 U18817 ( .A1(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n15797), .ZN(
        n15807) );
  NAND2_X1 U18818 ( .A1(n15796), .A2(n15795), .ZN(n15816) );
  INV_X1 U18819 ( .A(n15816), .ZN(n15801) );
  AOI21_X1 U18820 ( .B1(n15798), .B2(n15797), .A(n20046), .ZN(n15799) );
  OAI21_X1 U18821 ( .B1(n15819), .B2(n15800), .A(n15799), .ZN(n15813) );
  AOI21_X1 U18822 ( .B1(n15802), .B2(n15801), .A(n15813), .ZN(n15804) );
  OAI22_X1 U18823 ( .A1(n15805), .A2(n20070), .B1(n15804), .B2(n15803), .ZN(
        n15806) );
  AOI21_X1 U18824 ( .B1(n15807), .B2(n15811), .A(n15806), .ZN(n15809) );
  NAND2_X1 U18825 ( .A1(n20043), .A2(P1_REIP_REG_12__SCAN_IN), .ZN(n15808) );
  OAI211_X1 U18826 ( .C1(n20081), .C2(n15810), .A(n15809), .B(n15808), .ZN(
        P1_U3019) );
  NAND2_X1 U18827 ( .A1(n15818), .A2(n15811), .ZN(n15855) );
  AOI22_X1 U18828 ( .A1(n20043), .A2(P1_REIP_REG_11__SCAN_IN), .B1(n20064), 
        .B2(n9700), .ZN(n15815) );
  AOI22_X1 U18829 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n15813), .B1(
        n20078), .B2(n15812), .ZN(n15814) );
  OAI211_X1 U18830 ( .C1(n15855), .C2(n15816), .A(n15815), .B(n15814), .ZN(
        P1_U3020) );
  AOI21_X1 U18831 ( .B1(n15819), .B2(n15818), .A(n15817), .ZN(n15821) );
  AOI221_X1 U18832 ( .B1(n15821), .B2(n15834), .C1(n15820), .C2(n15834), .A(
        n20046), .ZN(n15832) );
  NOR2_X1 U18833 ( .A1(n15835), .A2(n15855), .ZN(n15843) );
  NAND3_X1 U18834 ( .A1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .A3(n15843), .ZN(n15827) );
  AOI221_X1 U18835 ( .B1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_9__SCAN_IN), .C1(n11184), .C2(n15833), .A(
        n15827), .ZN(n15824) );
  OAI22_X1 U18836 ( .A1(n20050), .A2(n20633), .B1(n20081), .B2(n15822), .ZN(
        n15823) );
  AOI211_X1 U18837 ( .C1(n15825), .C2(n20078), .A(n15824), .B(n15823), .ZN(
        n15826) );
  OAI21_X1 U18838 ( .B1(n11184), .B2(n15832), .A(n15826), .ZN(P1_U3021) );
  AND2_X1 U18839 ( .A1(n20043), .A2(P1_REIP_REG_9__SCAN_IN), .ZN(n15830) );
  OAI22_X1 U18840 ( .A1(n15828), .A2(n20070), .B1(
        P1_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n15827), .ZN(n15829) );
  AOI211_X1 U18841 ( .C1(n20064), .C2(n19841), .A(n15830), .B(n15829), .ZN(
        n15831) );
  OAI21_X1 U18842 ( .B1(n15833), .B2(n15832), .A(n15831), .ZN(P1_U3022) );
  AOI21_X1 U18843 ( .B1(n15835), .B2(n15834), .A(n15851), .ZN(n15848) );
  INV_X1 U18844 ( .A(P1_REIP_REG_8__SCAN_IN), .ZN(n20627) );
  OAI222_X1 U18845 ( .A1(n15837), .A2(n20081), .B1(n20050), .B2(n20627), .C1(
        n20070), .C2(n15836), .ZN(n15838) );
  INV_X1 U18846 ( .A(n15838), .ZN(n15840) );
  INV_X1 U18847 ( .A(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n15847) );
  OAI221_X1 U18848 ( .B1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .C1(n15841), .C2(n15847), .A(
        n15843), .ZN(n15839) );
  OAI211_X1 U18849 ( .C1(n15848), .C2(n15841), .A(n15840), .B(n15839), .ZN(
        P1_U3023) );
  INV_X1 U18850 ( .A(n19856), .ZN(n15842) );
  AOI22_X1 U18851 ( .A1(n20043), .A2(P1_REIP_REG_7__SCAN_IN), .B1(n20064), 
        .B2(n15842), .ZN(n15846) );
  AOI22_X1 U18852 ( .A1(n15844), .A2(n20078), .B1(n15847), .B2(n15843), .ZN(
        n15845) );
  OAI211_X1 U18853 ( .C1(n15848), .C2(n15847), .A(n15846), .B(n15845), .ZN(
        P1_U3024) );
  XNOR2_X1 U18854 ( .A(n15850), .B(n15849), .ZN(n19939) );
  AOI22_X1 U18855 ( .A1(n20043), .A2(P1_REIP_REG_6__SCAN_IN), .B1(n20064), 
        .B2(n19939), .ZN(n15854) );
  AOI22_X1 U18856 ( .A1(n15852), .A2(n20078), .B1(
        P1_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n15851), .ZN(n15853) );
  OAI211_X1 U18857 ( .C1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .C2(n15855), .A(
        n15854), .B(n15853), .ZN(P1_U3025) );
  INV_X1 U18858 ( .A(n15856), .ZN(n15858) );
  NAND3_X1 U18859 ( .A1(n15859), .A2(n15858), .A3(n15857), .ZN(n15860) );
  OAI21_X1 U18860 ( .B1(n15862), .B2(n15861), .A(n15860), .ZN(P1_U3468) );
  NAND2_X1 U18861 ( .A1(n20440), .A2(n20728), .ZN(n15869) );
  AOI21_X1 U18862 ( .B1(P1_STATE2_REG_0__SCAN_IN), .B2(n15871), .A(
        P1_STATE2_REG_1__SCAN_IN), .ZN(n15868) );
  NAND4_X1 U18863 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(
        P1_STATE2_REG_0__SCAN_IN), .A3(n20599), .A4(n20728), .ZN(n15863) );
  AND2_X1 U18864 ( .A1(n15864), .A2(n15863), .ZN(n20598) );
  AOI21_X1 U18865 ( .B1(n20598), .B2(n15866), .A(n15865), .ZN(n15867) );
  AOI211_X1 U18866 ( .C1(n20725), .C2(n15869), .A(n15868), .B(n15867), .ZN(
        P1_U3162) );
  OAI221_X1 U18867 ( .B1(n20440), .B2(P1_STATE2_REG_0__SCAN_IN), .C1(n20440), 
        .C2(n15871), .A(n15870), .ZN(P1_U3466) );
  AOI22_X1 U18868 ( .A1(n15872), .A2(n18896), .B1(P2_REIP_REG_31__SCAN_IN), 
        .B2(n18910), .ZN(n15880) );
  AOI22_X1 U18869 ( .A1(n18842), .A2(P2_EBX_REG_31__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_31__SCAN_IN), .B2(n18892), .ZN(n15879) );
  NAND2_X1 U18870 ( .A1(n18959), .A2(n18874), .ZN(n15873) );
  AND2_X1 U18871 ( .A1(n15874), .A2(n15873), .ZN(n15878) );
  NAND4_X1 U18872 ( .A1(n18920), .A2(n15876), .A3(n15875), .A4(n18831), .ZN(
        n15877) );
  NAND4_X1 U18873 ( .A1(n15880), .A2(n15879), .A3(n15878), .A4(n15877), .ZN(
        P2_U2824) );
  INV_X1 U18874 ( .A(n15881), .ZN(n15884) );
  INV_X1 U18875 ( .A(n15882), .ZN(n15883) );
  AOI211_X1 U18876 ( .C1(n15885), .C2(n15884), .A(n15883), .B(n18890), .ZN(
        n15890) );
  OAI222_X1 U18877 ( .A1(n18935), .A2(n15888), .B1(n18929), .B2(n15887), .C1(
        n18923), .C2(n15886), .ZN(n15889) );
  AOI211_X1 U18878 ( .C1(n18910), .C2(P2_REIP_REG_28__SCAN_IN), .A(n15890), 
        .B(n15889), .ZN(n15894) );
  AOI22_X1 U18879 ( .A1(n15892), .A2(n18916), .B1(n15891), .B2(n18874), .ZN(
        n15893) );
  NAND2_X1 U18880 ( .A1(n15894), .A2(n15893), .ZN(P2_U2827) );
  NOR2_X1 U18881 ( .A1(n18932), .A2(n19728), .ZN(n15898) );
  INV_X1 U18882 ( .A(P2_EBX_REG_27__SCAN_IN), .ZN(n15896) );
  OAI22_X1 U18883 ( .A1(n18929), .A2(n15896), .B1(n15895), .B2(n18935), .ZN(
        n15897) );
  AOI211_X1 U18884 ( .C1(n15899), .C2(n18916), .A(n15898), .B(n15897), .ZN(
        n15900) );
  OAI21_X1 U18885 ( .B1(n15901), .B2(n18923), .A(n15900), .ZN(n15906) );
  AOI211_X1 U18886 ( .C1(n15904), .C2(n15903), .A(n15902), .B(n18890), .ZN(
        n15905) );
  NOR2_X1 U18887 ( .A1(n15906), .A2(n15905), .ZN(n15907) );
  OAI21_X1 U18888 ( .B1(n15908), .B2(n18928), .A(n15907), .ZN(P2_U2828) );
  AOI22_X1 U18889 ( .A1(n15909), .A2(n18896), .B1(P2_REIP_REG_26__SCAN_IN), 
        .B2(n18910), .ZN(n15918) );
  AOI22_X1 U18890 ( .A1(n18842), .A2(P2_EBX_REG_26__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n18892), .ZN(n15917) );
  AOI22_X1 U18891 ( .A1(n15911), .A2(n18916), .B1(n18874), .B2(n15910), .ZN(
        n15916) );
  INV_X1 U18892 ( .A(n15912), .ZN(n15913) );
  AOI21_X1 U18893 ( .B1(n9902), .B2(n15913), .A(n9712), .ZN(n15914) );
  NAND2_X1 U18894 ( .A1(n18920), .A2(n15914), .ZN(n15915) );
  NAND4_X1 U18895 ( .A1(n15918), .A2(n15917), .A3(n15916), .A4(n15915), .ZN(
        P2_U2829) );
  AOI22_X1 U18896 ( .A1(n15919), .A2(n18896), .B1(P2_EBX_REG_24__SCAN_IN), 
        .B2(n18842), .ZN(n15931) );
  AOI22_X1 U18897 ( .A1(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n18892), .B1(
        P2_REIP_REG_24__SCAN_IN), .B2(n18910), .ZN(n15930) );
  OAI22_X1 U18898 ( .A1(n15969), .A2(n18924), .B1(n18928), .B2(n15920), .ZN(
        n15921) );
  INV_X1 U18899 ( .A(n15921), .ZN(n15929) );
  INV_X1 U18900 ( .A(n15922), .ZN(n15925) );
  INV_X1 U18901 ( .A(n15923), .ZN(n15924) );
  AOI21_X1 U18902 ( .B1(n15926), .B2(n15925), .A(n15924), .ZN(n15927) );
  NAND2_X1 U18903 ( .A1(n18920), .A2(n15927), .ZN(n15928) );
  NAND4_X1 U18904 ( .A1(n15931), .A2(n15930), .A3(n15929), .A4(n15928), .ZN(
        P2_U2831) );
  AOI22_X1 U18905 ( .A1(n18958), .A2(n15932), .B1(n12476), .B2(n18945), .ZN(
        P2_U2856) );
  AOI22_X1 U18906 ( .A1(n15933), .A2(n15942), .B1(P2_EBX_REG_23__SCAN_IN), 
        .B2(n15938), .ZN(n15934) );
  OAI21_X1 U18907 ( .B1(n18945), .B2(n15978), .A(n15934), .ZN(P2_U2864) );
  INV_X1 U18908 ( .A(n15989), .ZN(n15940) );
  AOI21_X1 U18909 ( .B1(n15937), .B2(n15936), .A(n15935), .ZN(n15951) );
  AOI22_X1 U18910 ( .A1(n15951), .A2(n15942), .B1(P2_EBX_REG_22__SCAN_IN), 
        .B2(n15938), .ZN(n15939) );
  OAI21_X1 U18911 ( .B1(n18945), .B2(n15940), .A(n15939), .ZN(P2_U2865) );
  AOI21_X1 U18912 ( .B1(n15941), .B2(n13844), .A(n9735), .ZN(n15956) );
  AOI22_X1 U18913 ( .A1(n15956), .A2(n15942), .B1(n18958), .B2(n18751), .ZN(
        n15943) );
  OAI21_X1 U18914 ( .B1(n15948), .B2(n11572), .A(n15943), .ZN(P2_U2867) );
  OAI22_X1 U18915 ( .A1(n15945), .A2(n18952), .B1(n18945), .B2(n15944), .ZN(
        n15946) );
  INV_X1 U18916 ( .A(n15946), .ZN(n15947) );
  OAI21_X1 U18917 ( .B1(n15948), .B2(n11999), .A(n15947), .ZN(P2_U2869) );
  INV_X1 U18918 ( .A(n18995), .ZN(n19026) );
  AOI22_X1 U18919 ( .A1(n18963), .A2(n15949), .B1(P2_EAX_REG_22__SCAN_IN), 
        .B2(n19026), .ZN(n15954) );
  AOI22_X1 U18920 ( .A1(n18965), .A2(BUF2_REG_22__SCAN_IN), .B1(n18964), .B2(
        BUF1_REG_22__SCAN_IN), .ZN(n15953) );
  AOI22_X1 U18921 ( .A1(n15951), .A2(n19031), .B1(n19027), .B2(n15950), .ZN(
        n15952) );
  NAND3_X1 U18922 ( .A1(n15954), .A2(n15953), .A3(n15952), .ZN(P2_U2897) );
  AOI22_X1 U18923 ( .A1(n18963), .A2(n15955), .B1(n19026), .B2(
        P2_EAX_REG_20__SCAN_IN), .ZN(n15959) );
  AOI22_X1 U18924 ( .A1(n18965), .A2(BUF2_REG_20__SCAN_IN), .B1(n18964), .B2(
        BUF1_REG_20__SCAN_IN), .ZN(n15958) );
  AOI22_X1 U18925 ( .A1(n15956), .A2(n19031), .B1(n19027), .B2(n18750), .ZN(
        n15957) );
  NAND3_X1 U18926 ( .A1(n15959), .A2(n15958), .A3(n15957), .ZN(P2_U2899) );
  OAI22_X1 U18927 ( .A1(n15960), .A2(n19093), .B1(n19724), .B2(n12482), .ZN(
        n15961) );
  AOI21_X1 U18928 ( .B1(n19080), .B2(n15962), .A(n15961), .ZN(n15967) );
  INV_X1 U18929 ( .A(n15963), .ZN(n15964) );
  AOI22_X1 U18930 ( .A1(n15965), .A2(n16066), .B1(n16068), .B2(n15964), .ZN(
        n15966) );
  OAI211_X1 U18931 ( .C1(n16072), .C2(n15968), .A(n15967), .B(n15966), .ZN(
        P2_U2989) );
  AOI22_X1 U18932 ( .A1(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n16001), .B1(
        P2_REIP_REG_24__SCAN_IN), .B2(n18810), .ZN(n15975) );
  INV_X1 U18933 ( .A(n15969), .ZN(n15973) );
  OAI22_X1 U18934 ( .A1(n15971), .A2(n19088), .B1(n19087), .B2(n15970), .ZN(
        n15972) );
  AOI21_X1 U18935 ( .B1(n19090), .B2(n15973), .A(n15972), .ZN(n15974) );
  OAI211_X1 U18936 ( .C1(n16063), .C2(n15976), .A(n15975), .B(n15974), .ZN(
        P2_U2990) );
  AOI22_X1 U18937 ( .A1(P2_REIP_REG_23__SCAN_IN), .A2(n19081), .B1(n19080), 
        .B2(n15977), .ZN(n15983) );
  INV_X1 U18938 ( .A(n15978), .ZN(n15980) );
  AOI222_X1 U18939 ( .A1(n15981), .A2(n16066), .B1(n19090), .B2(n15980), .C1(
        n16068), .C2(n15979), .ZN(n15982) );
  OAI211_X1 U18940 ( .C1(n15984), .C2(n19093), .A(n15983), .B(n15982), .ZN(
        P2_U2991) );
  AOI22_X1 U18941 ( .A1(P2_REIP_REG_22__SCAN_IN), .A2(n19081), .B1(n19080), 
        .B2(n15985), .ZN(n15991) );
  OAI22_X1 U18942 ( .A1(n15987), .A2(n19088), .B1(n19087), .B2(n15986), .ZN(
        n15988) );
  AOI21_X1 U18943 ( .B1(n19090), .B2(n15989), .A(n15988), .ZN(n15990) );
  OAI211_X1 U18944 ( .C1(n15308), .C2(n19093), .A(n15991), .B(n15990), .ZN(
        P2_U2992) );
  AOI21_X1 U18945 ( .B1(n19080), .B2(n15993), .A(n15992), .ZN(n15994) );
  OAI21_X1 U18946 ( .B1(n19093), .B2(n18771), .A(n15994), .ZN(n15998) );
  AOI211_X1 U18947 ( .C1(n16003), .C2(n15996), .A(n15995), .B(n19087), .ZN(
        n15997) );
  AOI211_X1 U18948 ( .C1(n16066), .C2(n15999), .A(n15998), .B(n15997), .ZN(
        n16000) );
  OAI21_X1 U18949 ( .B1(n16072), .B2(n18776), .A(n16000), .ZN(P2_U2997) );
  AOI22_X1 U18950 ( .A1(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(n16001), .B1(
        n19080), .B2(n18787), .ZN(n16007) );
  AOI22_X1 U18951 ( .A1(n16002), .A2(n16066), .B1(n19090), .B2(n18943), .ZN(
        n16006) );
  OAI211_X1 U18952 ( .C1(n16013), .C2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A(
        n16068), .B(n16003), .ZN(n16004) );
  NAND4_X1 U18953 ( .A1(n16007), .A2(n16006), .A3(n16005), .A4(n16004), .ZN(
        P2_U2998) );
  INV_X1 U18954 ( .A(n18798), .ZN(n16008) );
  AOI22_X1 U18955 ( .A1(P2_REIP_REG_15__SCAN_IN), .A2(n18810), .B1(n19080), 
        .B2(n16008), .ZN(n16016) );
  NAND2_X1 U18956 ( .A1(n16010), .A2(n16009), .ZN(n16012) );
  XOR2_X1 U18957 ( .A(n16012), .B(n16011), .Z(n16082) );
  INV_X1 U18958 ( .A(n16082), .ZN(n16014) );
  AOI21_X1 U18959 ( .B1(n12269), .B2(n16017), .A(n16013), .ZN(n16079) );
  AOI222_X1 U18960 ( .A1(n16014), .A2(n16066), .B1(n19090), .B2(n18802), .C1(
        n16068), .C2(n16079), .ZN(n16015) );
  OAI211_X1 U18961 ( .C1(n11215), .C2(n19093), .A(n16016), .B(n16015), .ZN(
        P2_U2999) );
  AOI22_X1 U18962 ( .A1(P2_REIP_REG_14__SCAN_IN), .A2(n18810), .B1(n19080), 
        .B2(n18807), .ZN(n16025) );
  OAI21_X1 U18963 ( .B1(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n16018), .A(
        n16017), .ZN(n16100) );
  NAND2_X1 U18964 ( .A1(n16020), .A2(n16019), .ZN(n16021) );
  XNOR2_X1 U18965 ( .A(n16022), .B(n16021), .ZN(n16096) );
  OAI22_X1 U18966 ( .A1(n16100), .A2(n19087), .B1(n19088), .B2(n16096), .ZN(
        n16023) );
  AOI21_X1 U18967 ( .B1(n19090), .B2(n18814), .A(n16023), .ZN(n16024) );
  OAI211_X1 U18968 ( .C1(n16026), .C2(n19093), .A(n16025), .B(n16024), .ZN(
        P2_U3000) );
  INV_X1 U18969 ( .A(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n16027) );
  OAI22_X1 U18970 ( .A1(n16027), .A2(n19093), .B1(n16063), .B2(n18823), .ZN(
        n16028) );
  AOI21_X1 U18971 ( .B1(P2_REIP_REG_13__SCAN_IN), .B2(n18810), .A(n16028), 
        .ZN(n16032) );
  AOI22_X1 U18972 ( .A1(n16030), .A2(n16068), .B1(n16066), .B2(n16029), .ZN(
        n16031) );
  OAI211_X1 U18973 ( .C1(n16072), .C2(n18824), .A(n16032), .B(n16031), .ZN(
        P2_U3001) );
  AOI22_X1 U18974 ( .A1(P2_REIP_REG_12__SCAN_IN), .A2(n19081), .B1(n19080), 
        .B2(n18832), .ZN(n16043) );
  INV_X1 U18975 ( .A(n16033), .ZN(n18838) );
  NAND2_X1 U18976 ( .A1(n9683), .A2(n16035), .ZN(n16036) );
  XNOR2_X1 U18977 ( .A(n16034), .B(n16036), .ZN(n16105) );
  INV_X1 U18978 ( .A(n16037), .ZN(n16038) );
  AOI21_X1 U18979 ( .B1(n16039), .B2(n16106), .A(n16038), .ZN(n16104) );
  AOI22_X1 U18980 ( .A1(n16105), .A2(n16066), .B1(n16104), .B2(n16068), .ZN(
        n16040) );
  INV_X1 U18981 ( .A(n16040), .ZN(n16041) );
  AOI21_X1 U18982 ( .B1(n19090), .B2(n18838), .A(n16041), .ZN(n16042) );
  OAI211_X1 U18983 ( .C1(n18834), .C2(n19093), .A(n16043), .B(n16042), .ZN(
        P2_U3002) );
  OAI22_X1 U18984 ( .A1(n11542), .A2(n19093), .B1(n16063), .B2(n18854), .ZN(
        n16044) );
  AOI21_X1 U18985 ( .B1(P2_REIP_REG_11__SCAN_IN), .B2(n18810), .A(n16044), 
        .ZN(n16048) );
  AOI22_X1 U18986 ( .A1(n16046), .A2(n16068), .B1(n16066), .B2(n16045), .ZN(
        n16047) );
  OAI211_X1 U18987 ( .C1(n16072), .C2(n18846), .A(n16048), .B(n16047), .ZN(
        P2_U3003) );
  AOI22_X1 U18988 ( .A1(P2_REIP_REG_10__SCAN_IN), .A2(n19081), .B1(n19080), 
        .B2(n18862), .ZN(n16053) );
  OAI22_X1 U18989 ( .A1(n16050), .A2(n19088), .B1(n16049), .B2(n19087), .ZN(
        n16051) );
  AOI21_X1 U18990 ( .B1(n19090), .B2(n18956), .A(n16051), .ZN(n16052) );
  OAI211_X1 U18991 ( .C1(n16054), .C2(n19093), .A(n16053), .B(n16052), .ZN(
        P2_U3004) );
  INV_X1 U18992 ( .A(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n16056) );
  OAI22_X1 U18993 ( .A1(n16056), .A2(n19093), .B1(n16063), .B2(n16055), .ZN(
        n16057) );
  AOI21_X1 U18994 ( .B1(P2_REIP_REG_9__SCAN_IN), .B2(n18810), .A(n16057), .ZN(
        n16061) );
  AOI22_X1 U18995 ( .A1(n16059), .A2(n16068), .B1(n16066), .B2(n16058), .ZN(
        n16060) );
  OAI211_X1 U18996 ( .C1(n16072), .C2(n16062), .A(n16061), .B(n16060), .ZN(
        P2_U3005) );
  OAI22_X1 U18997 ( .A1(n11213), .A2(n19093), .B1(n16063), .B2(n18881), .ZN(
        n16064) );
  AOI21_X1 U18998 ( .B1(P2_REIP_REG_7__SCAN_IN), .B2(n18810), .A(n16064), .ZN(
        n16071) );
  INV_X1 U18999 ( .A(n16065), .ZN(n16069) );
  AOI22_X1 U19000 ( .A1(n16069), .A2(n16068), .B1(n16067), .B2(n16066), .ZN(
        n16070) );
  OAI211_X1 U19001 ( .C1(n16072), .C2(n18885), .A(n16071), .B(n16070), .ZN(
        P2_U3007) );
  XOR2_X1 U19002 ( .A(n16073), .B(n16074), .Z(n18972) );
  NAND2_X1 U19003 ( .A1(P2_REIP_REG_15__SCAN_IN), .A2(n19081), .ZN(n16075) );
  OAI221_X1 U19004 ( .B1(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n16077), 
        .C1(n12269), .C2(n16076), .A(n16075), .ZN(n16078) );
  AOI21_X1 U19005 ( .B1(n19122), .B2(n18972), .A(n16078), .ZN(n16081) );
  AOI22_X1 U19006 ( .A1(n16079), .A2(n16122), .B1(n19131), .B2(n18802), .ZN(
        n16080) );
  OAI211_X1 U19007 ( .C1(n16082), .C2(n19110), .A(n16081), .B(n16080), .ZN(
        P2_U3031) );
  NOR2_X1 U19008 ( .A1(n16084), .A2(n16083), .ZN(n16088) );
  AOI221_X1 U19009 ( .B1(n16085), .B2(n16107), .C1(n16106), .C2(n16107), .A(
        n16103), .ZN(n16086) );
  INV_X1 U19010 ( .A(n16086), .ZN(n16087) );
  MUX2_X1 U19011 ( .A(n16088), .B(n16087), .S(
        P2_INSTADDRPOINTER_REG_14__SCAN_IN), .Z(n16095) );
  INV_X1 U19012 ( .A(P2_REIP_REG_14__SCAN_IN), .ZN(n19705) );
  NAND2_X1 U19013 ( .A1(n16090), .A2(n16089), .ZN(n16092) );
  INV_X1 U19014 ( .A(n16073), .ZN(n16091) );
  AND2_X1 U19015 ( .A1(n16092), .A2(n16091), .ZN(n18975) );
  NAND2_X1 U19016 ( .A1(n18975), .A2(n19122), .ZN(n16093) );
  OAI21_X1 U19017 ( .B1(n19705), .B2(n12482), .A(n16093), .ZN(n16094) );
  NOR2_X1 U19018 ( .A1(n16095), .A2(n16094), .ZN(n16099) );
  INV_X1 U19019 ( .A(n16096), .ZN(n16097) );
  AOI22_X1 U19020 ( .A1(n16097), .A2(n12942), .B1(n19131), .B2(n18814), .ZN(
        n16098) );
  OAI211_X1 U19021 ( .C1(n19125), .C2(n16100), .A(n16099), .B(n16098), .ZN(
        P2_U3032) );
  AOI21_X1 U19022 ( .B1(n14982), .B2(n16102), .A(n16101), .ZN(n18980) );
  AOI22_X1 U19023 ( .A1(n16103), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .B1(
        n18980), .B2(n19122), .ZN(n16111) );
  AOI222_X1 U19024 ( .A1(n16105), .A2(n12942), .B1(n19131), .B2(n18838), .C1(
        n16122), .C2(n16104), .ZN(n16110) );
  NAND2_X1 U19025 ( .A1(n16107), .A2(n16106), .ZN(n16109) );
  NAND2_X1 U19026 ( .A1(P2_REIP_REG_12__SCAN_IN), .A2(n19081), .ZN(n16108) );
  NAND4_X1 U19027 ( .A1(n16111), .A2(n16110), .A3(n16109), .A4(n16108), .ZN(
        P2_U3034) );
  AOI21_X1 U19028 ( .B1(n16113), .B2(n16112), .A(n9701), .ZN(n18990) );
  NOR2_X1 U19029 ( .A1(n16114), .A2(n19694), .ZN(n16121) );
  OAI21_X1 U19030 ( .B1(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A(n16115), .ZN(n16116) );
  OAI22_X1 U19031 ( .A1(n16119), .A2(n16118), .B1(n16117), .B2(n16116), .ZN(
        n16120) );
  AOI211_X1 U19032 ( .C1(n19122), .C2(n18990), .A(n16121), .B(n16120), .ZN(
        n16125) );
  AOI22_X1 U19033 ( .A1(n16123), .A2(n16122), .B1(n19131), .B2(n18875), .ZN(
        n16124) );
  OAI211_X1 U19034 ( .C1(n16126), .C2(n19110), .A(n16125), .B(n16124), .ZN(
        P2_U3038) );
  OAI21_X1 U19035 ( .B1(n16128), .B2(n19012), .A(n16127), .ZN(n16129) );
  AOI21_X1 U19036 ( .B1(n9650), .B2(n19131), .A(n16129), .ZN(n16130) );
  OAI21_X1 U19037 ( .B1(n16131), .B2(n19125), .A(n16130), .ZN(n16132) );
  AOI21_X1 U19038 ( .B1(n16133), .B2(n12942), .A(n16132), .ZN(n16134) );
  OAI221_X1 U19039 ( .B1(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n16136), .C1(
        n12162), .C2(n16135), .A(n16134), .ZN(P2_U3043) );
  AOI22_X1 U19040 ( .A1(n19124), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        n19122), .B2(n18926), .ZN(n16143) );
  OAI22_X1 U19041 ( .A1(n19110), .A2(n16138), .B1(n19125), .B2(n16137), .ZN(
        n16139) );
  AOI211_X1 U19042 ( .C1(n19131), .C2(n16141), .A(n16140), .B(n16139), .ZN(
        n16142) );
  OAI211_X1 U19043 ( .C1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .C2(n16144), .A(
        n16143), .B(n16142), .ZN(P2_U3046) );
  AOI211_X1 U19044 ( .C1(n19792), .C2(n16147), .A(n16146), .B(n16145), .ZN(
        n16151) );
  MUX2_X1 U19045 ( .A(n16148), .B(n19657), .S(P2_STATE2_REG_0__SCAN_IN), .Z(
        n16149) );
  NAND2_X1 U19046 ( .A1(n19657), .A2(n19807), .ZN(n19664) );
  OAI22_X1 U19047 ( .A1(n16149), .A2(n19799), .B1(n19664), .B2(
        P2_STATE2_REG_0__SCAN_IN), .ZN(n16150) );
  OAI211_X1 U19048 ( .C1(n16153), .C2(n16152), .A(n16151), .B(n16150), .ZN(
        P2_U3176) );
  INV_X1 U19049 ( .A(n16154), .ZN(n18489) );
  INV_X1 U19050 ( .A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n18651) );
  NAND2_X1 U19051 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n18651), .ZN(
        n16205) );
  INV_X1 U19052 ( .A(n16165), .ZN(n16156) );
  OAI211_X1 U19053 ( .C1(n15213), .C2(n16163), .A(n16205), .B(n16156), .ZN(
        n16161) );
  AOI21_X1 U19054 ( .B1(n15213), .B2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A(
        n18651), .ZN(n16157) );
  INV_X1 U19055 ( .A(n16157), .ZN(n16159) );
  NOR2_X1 U19056 ( .A1(n17615), .A2(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n16162) );
  INV_X1 U19057 ( .A(n16162), .ZN(n16158) );
  NAND2_X1 U19058 ( .A1(n16161), .A2(n16160), .ZN(n16169) );
  NOR2_X1 U19059 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n18651), .ZN(
        n16209) );
  AOI21_X1 U19060 ( .B1(n16209), .B2(n16163), .A(n16162), .ZN(n16164) );
  INV_X1 U19061 ( .A(n16164), .ZN(n16167) );
  NAND2_X1 U19062 ( .A1(n16165), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n16166) );
  NAND2_X1 U19063 ( .A1(n16167), .A2(n16166), .ZN(n16168) );
  NAND2_X1 U19064 ( .A1(n16169), .A2(n16168), .ZN(n16214) );
  INV_X1 U19065 ( .A(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n16693) );
  NAND2_X1 U19066 ( .A1(n17636), .A2(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n17609) );
  NAND2_X1 U19067 ( .A1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n17619) );
  INV_X1 U19068 ( .A(n17619), .ZN(n17599) );
  NAND2_X1 U19069 ( .A1(n17599), .A2(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n17598) );
  NAND2_X1 U19070 ( .A1(n17583), .A2(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n17532) );
  INV_X1 U19071 ( .A(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n16616) );
  NOR2_X1 U19072 ( .A1(n17568), .A2(n17550), .ZN(n17545) );
  NAND2_X1 U19073 ( .A1(n17545), .A2(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n17507) );
  INV_X1 U19074 ( .A(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n17490) );
  NAND3_X1 U19075 ( .A1(n17466), .A2(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n17454) );
  INV_X1 U19076 ( .A(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n17453) );
  INV_X1 U19077 ( .A(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n16471) );
  NAND2_X1 U19078 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n17391) );
  INV_X1 U19079 ( .A(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n17380) );
  NOR2_X1 U19080 ( .A1(n17391), .A2(n17380), .ZN(n16369) );
  NAND2_X1 U19081 ( .A1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n17358) );
  NAND2_X1 U19082 ( .A1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n16189), .ZN(
        n16170) );
  XOR2_X2 U19083 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .B(n16170), .Z(
        n16679) );
  INV_X1 U19084 ( .A(P3_REIP_REG_31__SCAN_IN), .ZN(n18628) );
  INV_X1 U19085 ( .A(n17971), .ZN(n18028) );
  NOR2_X1 U19086 ( .A1(n18628), .A2(n18028), .ZN(n16208) );
  NOR2_X1 U19087 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n18704), .ZN(n17549) );
  NAND2_X1 U19088 ( .A1(n18388), .A2(n16171), .ZN(n18078) );
  INV_X1 U19089 ( .A(n17544), .ZN(n17509) );
  OR2_X1 U19090 ( .A1(n9672), .A2(n17509), .ZN(n16180) );
  INV_X1 U19091 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n16391) );
  XOR2_X1 U19092 ( .A(n16391), .B(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .Z(
        n16172) );
  NOR2_X1 U19093 ( .A1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n17427), .ZN(
        n16191) );
  NOR2_X1 U19094 ( .A1(n16693), .A2(n9736), .ZN(n16370) );
  INV_X1 U19095 ( .A(n17549), .ZN(n18554) );
  NAND2_X1 U19096 ( .A1(n18426), .A2(n9672), .ZN(n16194) );
  OAI211_X1 U19097 ( .C1(n16370), .C2(n18554), .A(n16194), .B(n17707), .ZN(
        n16197) );
  NOR2_X1 U19098 ( .A1(n16191), .A2(n16197), .ZN(n16179) );
  OAI22_X1 U19099 ( .A1(n16180), .A2(n16172), .B1(n16179), .B2(n16391), .ZN(
        n16173) );
  AOI211_X1 U19100 ( .C1(n17565), .C2(n10006), .A(n16208), .B(n16173), .ZN(
        n16177) );
  NAND2_X1 U19101 ( .A1(n16198), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n16174) );
  XNOR2_X1 U19102 ( .A(n16174), .B(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n16211) );
  NAND2_X1 U19103 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n16187), .ZN(
        n16175) );
  XNOR2_X1 U19104 ( .A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B(n16175), .ZN(
        n16210) );
  AOI22_X1 U19105 ( .A1(n17697), .A2(n16211), .B1(n17401), .B2(n16210), .ZN(
        n16176) );
  XOR2_X1 U19106 ( .A(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .B(n16189), .Z(
        n16394) );
  INV_X1 U19107 ( .A(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n16395) );
  NAND2_X1 U19108 ( .A1(n17971), .A2(P3_REIP_REG_30__SCAN_IN), .ZN(n16178) );
  OAI221_X1 U19109 ( .B1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n16180), .C1(
        n16395), .C2(n16179), .A(n16178), .ZN(n16181) );
  AOI21_X1 U19110 ( .B1(n17565), .B2(n16394), .A(n16181), .ZN(n16186) );
  OAI22_X1 U19111 ( .A1(n16198), .A2(n17710), .B1(n16187), .B2(n17616), .ZN(
        n16184) );
  INV_X1 U19112 ( .A(n17875), .ZN(n17902) );
  NAND2_X1 U19113 ( .A1(n17772), .A2(n17499), .ZN(n17440) );
  NOR2_X1 U19114 ( .A1(n17436), .A2(n17440), .ZN(n17352) );
  INV_X1 U19115 ( .A(n17352), .ZN(n17424) );
  NOR2_X1 U19116 ( .A1(n17712), .A2(n17424), .ZN(n17371) );
  AOI22_X1 U19117 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n16184), .B1(
        n16183), .B2(n17371), .ZN(n16185) );
  OAI211_X1 U19118 ( .C1(n10126), .C2(n17617), .A(n16186), .B(n16185), .ZN(
        P3_U2800) );
  INV_X1 U19119 ( .A(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n16188) );
  AOI211_X1 U19120 ( .C1(n16188), .C2(n16227), .A(n16187), .B(n17616), .ZN(
        n16196) );
  INV_X1 U19121 ( .A(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n16405) );
  INV_X1 U19122 ( .A(n16370), .ZN(n16190) );
  AOI21_X1 U19123 ( .B1(n16405), .B2(n16190), .A(n16189), .ZN(n16404) );
  OAI21_X1 U19124 ( .B1(n16191), .B2(n17565), .A(n16404), .ZN(n16192) );
  OAI211_X1 U19125 ( .C1(n16194), .C2(n9736), .A(n16193), .B(n16192), .ZN(
        n16195) );
  AOI211_X1 U19126 ( .C1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .C2(n16197), .A(
        n16196), .B(n16195), .ZN(n16201) );
  NOR2_X1 U19127 ( .A1(n16198), .A2(n17710), .ZN(n16199) );
  OAI21_X1 U19128 ( .B1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n16224), .A(
        n16199), .ZN(n16200) );
  OAI211_X1 U19129 ( .C1(n16202), .C2(n17617), .A(n16201), .B(n16200), .ZN(
        P3_U2801) );
  NAND2_X1 U19130 ( .A1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(n16203), .ZN(
        n16204) );
  OAI22_X1 U19131 ( .A1(n16206), .A2(n18651), .B1(n16205), .B2(n16204), .ZN(
        n16207) );
  AOI211_X1 U19132 ( .C1(n16209), .C2(n17979), .A(n16208), .B(n16207), .ZN(
        n16213) );
  AOI22_X1 U19133 ( .A1(n16211), .A2(n17999), .B1(n16210), .B2(n17877), .ZN(
        n16212) );
  OAI211_X1 U19134 ( .C1(n16214), .C2(n17940), .A(n16213), .B(n16212), .ZN(
        P3_U2831) );
  INV_X1 U19135 ( .A(n17364), .ZN(n16217) );
  OAI22_X1 U19136 ( .A1(n17349), .A2(n17615), .B1(n15213), .B2(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n17345) );
  INV_X1 U19137 ( .A(n17345), .ZN(n16218) );
  INV_X1 U19138 ( .A(n16219), .ZN(n16221) );
  NAND2_X1 U19139 ( .A1(n18490), .A2(n17193), .ZN(n16220) );
  NOR2_X1 U19140 ( .A1(n16221), .A2(n16220), .ZN(n16222) );
  NAND2_X1 U19141 ( .A1(n17343), .A2(n16222), .ZN(n16231) );
  INV_X1 U19142 ( .A(n16225), .ZN(n16229) );
  NOR2_X1 U19143 ( .A1(n16226), .A2(n17193), .ZN(n17884) );
  NAND2_X1 U19144 ( .A1(n16227), .A2(n17884), .ZN(n16228) );
  AND2_X1 U19145 ( .A1(n16229), .A2(n16228), .ZN(n16230) );
  INV_X1 U19146 ( .A(n17813), .ZN(n16233) );
  AOI21_X1 U19147 ( .B1(n18510), .B2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n18499), .ZN(n18002) );
  INV_X1 U19148 ( .A(n18486), .ZN(n17771) );
  AOI22_X1 U19149 ( .A1(n17771), .A2(n17847), .B1(n17846), .B2(n17884), .ZN(
        n17821) );
  OAI21_X1 U19150 ( .B1(n16233), .B2(n18002), .A(n17821), .ZN(n16234) );
  INV_X1 U19151 ( .A(n16234), .ZN(n16236) );
  OAI21_X1 U19152 ( .B1(n16236), .B2(n17485), .A(n16235), .ZN(n17784) );
  NAND2_X1 U19153 ( .A1(n16237), .A2(n17784), .ZN(n17761) );
  NOR2_X1 U19154 ( .A1(n18019), .A2(n17761), .ZN(n17726) );
  NOR2_X1 U19155 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n16238), .ZN(
        n17351) );
  AOI22_X1 U19156 ( .A1(n17971), .A2(P3_REIP_REG_28__SCAN_IN), .B1(n17726), 
        .B2(n17351), .ZN(n16244) );
  AND2_X1 U19157 ( .A1(n10125), .A2(n17349), .ZN(n16240) );
  AND2_X1 U19158 ( .A1(n17364), .A2(n17345), .ZN(n16239) );
  INV_X1 U19159 ( .A(n16241), .ZN(n16242) );
  OAI211_X1 U19160 ( .C1(n17349), .C2(n16245), .A(n16244), .B(n16243), .ZN(
        P3_U2834) );
  NOR3_X1 U19161 ( .A1(P3_W_R_N_REG_SCAN_IN), .A2(P3_BE_N_REG_0__SCAN_IN), 
        .A3(P3_BE_N_REG_1__SCAN_IN), .ZN(n16247) );
  NOR4_X1 U19162 ( .A1(P3_BE_N_REG_2__SCAN_IN), .A2(P3_BE_N_REG_3__SCAN_IN), 
        .A3(P3_D_C_N_REG_SCAN_IN), .A4(P3_ADS_N_REG_SCAN_IN), .ZN(n16246) );
  NAND4_X1 U19163 ( .A1(P3_M_IO_N_REG_SCAN_IN), .A2(n16247), .A3(n16246), .A4(
        U215), .ZN(U213) );
  INV_X1 U19164 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n16335) );
  INV_X2 U19165 ( .A(U214), .ZN(n16298) );
  NOR2_X1 U19166 ( .A1(n16298), .A2(n16248), .ZN(n16296) );
  INV_X1 U19167 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n19036) );
  OAI222_X1 U19168 ( .A1(U214), .A2(n16335), .B1(n16300), .B2(n16249), .C1(
        U212), .C2(n19036), .ZN(U216) );
  AOI222_X1 U19169 ( .A1(n16298), .A2(P1_DATAO_REG_30__SCAN_IN), .B1(n16296), 
        .B2(BUF1_REG_30__SCAN_IN), .C1(n16293), .C2(P2_DATAO_REG_30__SCAN_IN), 
        .ZN(n16250) );
  INV_X1 U19170 ( .A(n16250), .ZN(U217) );
  INV_X1 U19171 ( .A(BUF1_REG_29__SCAN_IN), .ZN(n16252) );
  AOI22_X1 U19172 ( .A1(P2_DATAO_REG_29__SCAN_IN), .A2(n16293), .B1(
        P1_DATAO_REG_29__SCAN_IN), .B2(n16298), .ZN(n16251) );
  OAI21_X1 U19173 ( .B1(n16252), .B2(n16300), .A(n16251), .ZN(U218) );
  INV_X1 U19174 ( .A(BUF1_REG_28__SCAN_IN), .ZN(n20837) );
  AOI22_X1 U19175 ( .A1(P2_DATAO_REG_28__SCAN_IN), .A2(n16293), .B1(
        P1_DATAO_REG_28__SCAN_IN), .B2(n16298), .ZN(n16253) );
  OAI21_X1 U19176 ( .B1(n20837), .B2(n16300), .A(n16253), .ZN(U219) );
  INV_X1 U19177 ( .A(BUF1_REG_27__SCAN_IN), .ZN(n16255) );
  AOI22_X1 U19178 ( .A1(P2_DATAO_REG_27__SCAN_IN), .A2(n16293), .B1(
        P1_DATAO_REG_27__SCAN_IN), .B2(n16298), .ZN(n16254) );
  OAI21_X1 U19179 ( .B1(n16255), .B2(n16300), .A(n16254), .ZN(U220) );
  AOI22_X1 U19180 ( .A1(P2_DATAO_REG_26__SCAN_IN), .A2(n16293), .B1(
        P1_DATAO_REG_26__SCAN_IN), .B2(n16298), .ZN(n16256) );
  OAI21_X1 U19181 ( .B1(n16257), .B2(n16300), .A(n16256), .ZN(U221) );
  INV_X1 U19182 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n16258) );
  OAI222_X1 U19183 ( .A1(U214), .A2(n16258), .B1(n16300), .B2(n14388), .C1(
        U212), .C2(n20802), .ZN(U222) );
  AOI22_X1 U19184 ( .A1(P2_DATAO_REG_24__SCAN_IN), .A2(n16293), .B1(
        P1_DATAO_REG_24__SCAN_IN), .B2(n16298), .ZN(n16259) );
  OAI21_X1 U19185 ( .B1(n14392), .B2(n16300), .A(n16259), .ZN(U223) );
  INV_X1 U19186 ( .A(BUF1_REG_23__SCAN_IN), .ZN(n16261) );
  AOI22_X1 U19187 ( .A1(P2_DATAO_REG_23__SCAN_IN), .A2(n16293), .B1(
        P1_DATAO_REG_23__SCAN_IN), .B2(n16298), .ZN(n16260) );
  OAI21_X1 U19188 ( .B1(n16261), .B2(n16300), .A(n16260), .ZN(U224) );
  AOI22_X1 U19189 ( .A1(P2_DATAO_REG_22__SCAN_IN), .A2(n16293), .B1(
        P1_DATAO_REG_22__SCAN_IN), .B2(n16298), .ZN(n16262) );
  OAI21_X1 U19190 ( .B1(n16263), .B2(n16300), .A(n16262), .ZN(U225) );
  AOI222_X1 U19191 ( .A1(n16298), .A2(P1_DATAO_REG_21__SCAN_IN), .B1(n16296), 
        .B2(BUF1_REG_21__SCAN_IN), .C1(n16293), .C2(P2_DATAO_REG_21__SCAN_IN), 
        .ZN(n16264) );
  INV_X1 U19192 ( .A(n16264), .ZN(U226) );
  AOI22_X1 U19193 ( .A1(P2_DATAO_REG_20__SCAN_IN), .A2(n16293), .B1(
        P1_DATAO_REG_20__SCAN_IN), .B2(n16298), .ZN(n16265) );
  OAI21_X1 U19194 ( .B1(n14410), .B2(n16300), .A(n16265), .ZN(U227) );
  AOI22_X1 U19195 ( .A1(P2_DATAO_REG_19__SCAN_IN), .A2(n16293), .B1(
        P1_DATAO_REG_19__SCAN_IN), .B2(n16298), .ZN(n16266) );
  OAI21_X1 U19196 ( .B1(n14416), .B2(n16300), .A(n16266), .ZN(U228) );
  INV_X1 U19197 ( .A(BUF1_REG_18__SCAN_IN), .ZN(n16268) );
  AOI22_X1 U19198 ( .A1(P2_DATAO_REG_18__SCAN_IN), .A2(n16293), .B1(
        P1_DATAO_REG_18__SCAN_IN), .B2(n16298), .ZN(n16267) );
  OAI21_X1 U19199 ( .B1(n16268), .B2(n16300), .A(n16267), .ZN(U229) );
  AOI22_X1 U19200 ( .A1(P2_DATAO_REG_17__SCAN_IN), .A2(n16293), .B1(
        P1_DATAO_REG_17__SCAN_IN), .B2(n16298), .ZN(n16269) );
  OAI21_X1 U19201 ( .B1(n14427), .B2(n16300), .A(n16269), .ZN(U230) );
  AOI22_X1 U19202 ( .A1(P2_DATAO_REG_16__SCAN_IN), .A2(n16293), .B1(
        P1_DATAO_REG_16__SCAN_IN), .B2(n16298), .ZN(n16270) );
  OAI21_X1 U19203 ( .B1(n20909), .B2(n16300), .A(n16270), .ZN(U231) );
  INV_X1 U19204 ( .A(BUF1_REG_15__SCAN_IN), .ZN(n16272) );
  AOI22_X1 U19205 ( .A1(P2_DATAO_REG_15__SCAN_IN), .A2(n16293), .B1(
        P1_DATAO_REG_15__SCAN_IN), .B2(n16298), .ZN(n16271) );
  OAI21_X1 U19206 ( .B1(n16272), .B2(n16300), .A(n16271), .ZN(U232) );
  INV_X1 U19207 ( .A(BUF1_REG_14__SCAN_IN), .ZN(n16274) );
  AOI22_X1 U19208 ( .A1(P2_DATAO_REG_14__SCAN_IN), .A2(n16293), .B1(
        P1_DATAO_REG_14__SCAN_IN), .B2(n16298), .ZN(n16273) );
  OAI21_X1 U19209 ( .B1(n16274), .B2(n16300), .A(n16273), .ZN(U233) );
  AOI22_X1 U19210 ( .A1(P2_DATAO_REG_13__SCAN_IN), .A2(n16293), .B1(
        P1_DATAO_REG_13__SCAN_IN), .B2(n16298), .ZN(n16275) );
  OAI21_X1 U19211 ( .B1(n13116), .B2(n16300), .A(n16275), .ZN(U234) );
  INV_X1 U19212 ( .A(BUF1_REG_12__SCAN_IN), .ZN(n16277) );
  AOI22_X1 U19213 ( .A1(P2_DATAO_REG_12__SCAN_IN), .A2(n16293), .B1(
        P1_DATAO_REG_12__SCAN_IN), .B2(n16298), .ZN(n16276) );
  OAI21_X1 U19214 ( .B1(n16277), .B2(n16300), .A(n16276), .ZN(U235) );
  INV_X1 U19215 ( .A(BUF1_REG_11__SCAN_IN), .ZN(n16279) );
  AOI22_X1 U19216 ( .A1(P2_DATAO_REG_11__SCAN_IN), .A2(n16293), .B1(
        P1_DATAO_REG_11__SCAN_IN), .B2(n16298), .ZN(n16278) );
  OAI21_X1 U19217 ( .B1(n16279), .B2(n16300), .A(n16278), .ZN(U236) );
  AOI22_X1 U19218 ( .A1(P2_DATAO_REG_10__SCAN_IN), .A2(n16293), .B1(
        P1_DATAO_REG_10__SCAN_IN), .B2(n16298), .ZN(n16280) );
  OAI21_X1 U19219 ( .B1(n16281), .B2(n16300), .A(n16280), .ZN(U237) );
  INV_X1 U19220 ( .A(BUF1_REG_9__SCAN_IN), .ZN(n16283) );
  AOI22_X1 U19221 ( .A1(P2_DATAO_REG_9__SCAN_IN), .A2(n16293), .B1(
        P1_DATAO_REG_9__SCAN_IN), .B2(n16298), .ZN(n16282) );
  OAI21_X1 U19222 ( .B1(n16283), .B2(n16300), .A(n16282), .ZN(U238) );
  AOI22_X1 U19223 ( .A1(P2_DATAO_REG_8__SCAN_IN), .A2(n16293), .B1(
        P1_DATAO_REG_8__SCAN_IN), .B2(n16298), .ZN(n16284) );
  OAI21_X1 U19224 ( .B1(n16285), .B2(n16300), .A(n16284), .ZN(U239) );
  INV_X1 U19225 ( .A(BUF1_REG_7__SCAN_IN), .ZN(n16287) );
  AOI22_X1 U19226 ( .A1(P2_DATAO_REG_7__SCAN_IN), .A2(n16293), .B1(
        P1_DATAO_REG_7__SCAN_IN), .B2(n16298), .ZN(n16286) );
  OAI21_X1 U19227 ( .B1(n16287), .B2(n16300), .A(n16286), .ZN(U240) );
  INV_X1 U19228 ( .A(BUF1_REG_6__SCAN_IN), .ZN(n16289) );
  AOI22_X1 U19229 ( .A1(P2_DATAO_REG_6__SCAN_IN), .A2(n16293), .B1(
        P1_DATAO_REG_6__SCAN_IN), .B2(n16298), .ZN(n16288) );
  OAI21_X1 U19230 ( .B1(n16289), .B2(n16300), .A(n16288), .ZN(U241) );
  INV_X1 U19231 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n20905) );
  AOI22_X1 U19232 ( .A1(BUF1_REG_5__SCAN_IN), .A2(n16296), .B1(
        P2_DATAO_REG_5__SCAN_IN), .B2(n16293), .ZN(n16290) );
  OAI21_X1 U19233 ( .B1(n20905), .B2(U214), .A(n16290), .ZN(U242) );
  INV_X1 U19234 ( .A(BUF1_REG_4__SCAN_IN), .ZN(n16292) );
  AOI22_X1 U19235 ( .A1(P2_DATAO_REG_4__SCAN_IN), .A2(n16293), .B1(
        P1_DATAO_REG_4__SCAN_IN), .B2(n16298), .ZN(n16291) );
  OAI21_X1 U19236 ( .B1(n16292), .B2(n16300), .A(n16291), .ZN(U243) );
  INV_X1 U19237 ( .A(BUF1_REG_3__SCAN_IN), .ZN(n20911) );
  AOI22_X1 U19238 ( .A1(P2_DATAO_REG_3__SCAN_IN), .A2(n16293), .B1(
        P1_DATAO_REG_3__SCAN_IN), .B2(n16298), .ZN(n16294) );
  OAI21_X1 U19239 ( .B1(n20911), .B2(n16300), .A(n16294), .ZN(U244) );
  INV_X1 U19240 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n19064) );
  AOI22_X1 U19241 ( .A1(BUF1_REG_2__SCAN_IN), .A2(n16296), .B1(
        P1_DATAO_REG_2__SCAN_IN), .B2(n16298), .ZN(n16295) );
  OAI21_X1 U19242 ( .B1(n19064), .B2(U212), .A(n16295), .ZN(U245) );
  INV_X1 U19243 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n16303) );
  AOI22_X1 U19244 ( .A1(BUF1_REG_1__SCAN_IN), .A2(n16296), .B1(
        P1_DATAO_REG_1__SCAN_IN), .B2(n16298), .ZN(n16297) );
  OAI21_X1 U19245 ( .B1(n16303), .B2(U212), .A(n16297), .ZN(U246) );
  AOI22_X1 U19246 ( .A1(P2_DATAO_REG_0__SCAN_IN), .A2(n16293), .B1(
        P1_DATAO_REG_0__SCAN_IN), .B2(n16298), .ZN(n16299) );
  OAI21_X1 U19247 ( .B1(n16301), .B2(n16300), .A(n16299), .ZN(U247) );
  INV_X1 U19248 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n16302) );
  AOI22_X1 U19249 ( .A1(n16331), .A2(n16302), .B1(n18048), .B2(U215), .ZN(U251) );
  INV_X1 U19250 ( .A(BUF2_REG_1__SCAN_IN), .ZN(n18055) );
  AOI22_X1 U19251 ( .A1(n16331), .A2(n16303), .B1(n18055), .B2(U215), .ZN(U252) );
  INV_X1 U19252 ( .A(BUF2_REG_2__SCAN_IN), .ZN(n18059) );
  AOI22_X1 U19253 ( .A1(n16331), .A2(n19064), .B1(n18059), .B2(U215), .ZN(U253) );
  INV_X1 U19254 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n16304) );
  INV_X1 U19255 ( .A(BUF2_REG_3__SCAN_IN), .ZN(n18064) );
  AOI22_X1 U19256 ( .A1(n16331), .A2(n16304), .B1(n18064), .B2(U215), .ZN(U254) );
  INV_X1 U19257 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n16305) );
  INV_X1 U19258 ( .A(BUF2_REG_4__SCAN_IN), .ZN(n18067) );
  AOI22_X1 U19259 ( .A1(n16331), .A2(n16305), .B1(n18067), .B2(U215), .ZN(U255) );
  INV_X1 U19260 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n16306) );
  INV_X1 U19261 ( .A(BUF2_REG_5__SCAN_IN), .ZN(n18072) );
  AOI22_X1 U19262 ( .A1(n16332), .A2(n16306), .B1(n18072), .B2(U215), .ZN(U256) );
  INV_X1 U19263 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n16307) );
  INV_X1 U19264 ( .A(BUF2_REG_6__SCAN_IN), .ZN(n18080) );
  AOI22_X1 U19265 ( .A1(n16332), .A2(n16307), .B1(n18080), .B2(U215), .ZN(U257) );
  INV_X1 U19266 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n16308) );
  INV_X1 U19267 ( .A(BUF2_REG_7__SCAN_IN), .ZN(n18084) );
  AOI22_X1 U19268 ( .A1(n16331), .A2(n16308), .B1(n18084), .B2(U215), .ZN(U258) );
  INV_X1 U19269 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n16309) );
  INV_X1 U19270 ( .A(BUF2_REG_8__SCAN_IN), .ZN(n17320) );
  AOI22_X1 U19271 ( .A1(n16332), .A2(n16309), .B1(n17320), .B2(U215), .ZN(U259) );
  INV_X1 U19272 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n16310) );
  AOI22_X1 U19273 ( .A1(n16331), .A2(n16310), .B1(n13109), .B2(U215), .ZN(U260) );
  INV_X1 U19274 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n16311) );
  INV_X1 U19275 ( .A(BUF2_REG_10__SCAN_IN), .ZN(n17324) );
  AOI22_X1 U19276 ( .A1(n16332), .A2(n16311), .B1(n17324), .B2(U215), .ZN(U261) );
  OAI22_X1 U19277 ( .A1(U215), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(
        BUF2_REG_11__SCAN_IN), .B2(n16331), .ZN(n16312) );
  INV_X1 U19278 ( .A(n16312), .ZN(U262) );
  INV_X1 U19279 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n16313) );
  INV_X1 U19280 ( .A(BUF2_REG_12__SCAN_IN), .ZN(n17328) );
  AOI22_X1 U19281 ( .A1(n16331), .A2(n16313), .B1(n17328), .B2(U215), .ZN(U263) );
  INV_X1 U19282 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n16314) );
  INV_X1 U19283 ( .A(BUF2_REG_13__SCAN_IN), .ZN(n17332) );
  AOI22_X1 U19284 ( .A1(n16332), .A2(n16314), .B1(n17332), .B2(U215), .ZN(U264) );
  OAI22_X1 U19285 ( .A1(U215), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(
        BUF2_REG_14__SCAN_IN), .B2(n16331), .ZN(n16315) );
  INV_X1 U19286 ( .A(n16315), .ZN(U265) );
  OAI22_X1 U19287 ( .A1(U215), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n16331), .ZN(n16316) );
  INV_X1 U19288 ( .A(n16316), .ZN(U266) );
  INV_X1 U19289 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n16317) );
  AOI22_X1 U19290 ( .A1(n16332), .A2(n16317), .B1(n18052), .B2(U215), .ZN(U267) );
  INV_X1 U19291 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n16318) );
  INV_X1 U19292 ( .A(BUF2_REG_17__SCAN_IN), .ZN(n19151) );
  AOI22_X1 U19293 ( .A1(n16331), .A2(n16318), .B1(n19151), .B2(U215), .ZN(U268) );
  OAI22_X1 U19294 ( .A1(U215), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n16331), .ZN(n16319) );
  INV_X1 U19295 ( .A(n16319), .ZN(U269) );
  INV_X1 U19296 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n16320) );
  INV_X1 U19297 ( .A(BUF2_REG_19__SCAN_IN), .ZN(n19158) );
  AOI22_X1 U19298 ( .A1(n16331), .A2(n16320), .B1(n19158), .B2(U215), .ZN(U270) );
  INV_X1 U19299 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n16321) );
  INV_X1 U19300 ( .A(BUF2_REG_20__SCAN_IN), .ZN(n19164) );
  AOI22_X1 U19301 ( .A1(n16331), .A2(n16321), .B1(n19164), .B2(U215), .ZN(U271) );
  INV_X1 U19302 ( .A(BUF2_REG_21__SCAN_IN), .ZN(n18073) );
  AOI22_X1 U19303 ( .A1(n16331), .A2(n20816), .B1(n18073), .B2(U215), .ZN(U272) );
  OAI22_X1 U19304 ( .A1(U215), .A2(P2_DATAO_REG_22__SCAN_IN), .B1(
        BUF2_REG_22__SCAN_IN), .B2(n16331), .ZN(n16322) );
  INV_X1 U19305 ( .A(n16322), .ZN(U273) );
  OAI22_X1 U19306 ( .A1(U215), .A2(P2_DATAO_REG_23__SCAN_IN), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n16332), .ZN(n16323) );
  INV_X1 U19307 ( .A(n16323), .ZN(U274) );
  OAI22_X1 U19308 ( .A1(U215), .A2(P2_DATAO_REG_24__SCAN_IN), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n16332), .ZN(n16324) );
  INV_X1 U19309 ( .A(n16324), .ZN(U275) );
  OAI22_X1 U19310 ( .A1(U215), .A2(P2_DATAO_REG_25__SCAN_IN), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n16331), .ZN(n16325) );
  INV_X1 U19311 ( .A(n16325), .ZN(U276) );
  INV_X1 U19312 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n16326) );
  AOI22_X1 U19313 ( .A1(n16331), .A2(n16326), .B1(n18060), .B2(U215), .ZN(U277) );
  OAI22_X1 U19314 ( .A1(U215), .A2(P2_DATAO_REG_27__SCAN_IN), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n16331), .ZN(n16327) );
  INV_X1 U19315 ( .A(n16327), .ZN(U278) );
  INV_X1 U19316 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n16328) );
  INV_X1 U19317 ( .A(BUF2_REG_28__SCAN_IN), .ZN(n17096) );
  AOI22_X1 U19318 ( .A1(n16332), .A2(n16328), .B1(n17096), .B2(U215), .ZN(U279) );
  OAI22_X1 U19319 ( .A1(U215), .A2(P2_DATAO_REG_29__SCAN_IN), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n16331), .ZN(n16329) );
  INV_X1 U19320 ( .A(n16329), .ZN(U280) );
  INV_X1 U19321 ( .A(BUF2_REG_30__SCAN_IN), .ZN(n18079) );
  AOI22_X1 U19322 ( .A1(n16331), .A2(n16330), .B1(n18079), .B2(U215), .ZN(U281) );
  OAI22_X1 U19323 ( .A1(U215), .A2(P2_DATAO_REG_31__SCAN_IN), .B1(
        BUF2_REG_31__SCAN_IN), .B2(n16332), .ZN(n16333) );
  INV_X1 U19324 ( .A(n16333), .ZN(U282) );
  INV_X1 U19325 ( .A(P3_DATAO_REG_31__SCAN_IN), .ZN(n16334) );
  AOI222_X1 U19326 ( .A1(n19036), .A2(P2_DATAO_REG_30__SCAN_IN), .B1(n16335), 
        .B2(P1_DATAO_REG_30__SCAN_IN), .C1(n16334), .C2(
        P3_DATAO_REG_30__SCAN_IN), .ZN(n16336) );
  INV_X1 U19327 ( .A(n16338), .ZN(n16337) );
  INV_X1 U19328 ( .A(P3_ADDRESS_REG_9__SCAN_IN), .ZN(n18589) );
  INV_X1 U19329 ( .A(P2_ADDRESS_REG_9__SCAN_IN), .ZN(n19699) );
  AOI22_X1 U19330 ( .A1(n16337), .A2(n18589), .B1(n19699), .B2(n16338), .ZN(
        U347) );
  INV_X1 U19331 ( .A(n16338), .ZN(n16339) );
  INV_X1 U19332 ( .A(P3_ADDRESS_REG_8__SCAN_IN), .ZN(n18587) );
  INV_X1 U19333 ( .A(P2_ADDRESS_REG_8__SCAN_IN), .ZN(n19697) );
  AOI22_X1 U19334 ( .A1(n16339), .A2(n18587), .B1(n19697), .B2(n16338), .ZN(
        U348) );
  INV_X1 U19335 ( .A(P3_ADDRESS_REG_7__SCAN_IN), .ZN(n18584) );
  INV_X1 U19336 ( .A(P2_ADDRESS_REG_7__SCAN_IN), .ZN(n19695) );
  AOI22_X1 U19337 ( .A1(n16337), .A2(n18584), .B1(n19695), .B2(n16338), .ZN(
        U349) );
  INV_X1 U19338 ( .A(P3_ADDRESS_REG_6__SCAN_IN), .ZN(n18583) );
  INV_X1 U19339 ( .A(P2_ADDRESS_REG_6__SCAN_IN), .ZN(n19693) );
  AOI22_X1 U19340 ( .A1(n16337), .A2(n18583), .B1(n19693), .B2(n16338), .ZN(
        U350) );
  INV_X1 U19341 ( .A(P3_ADDRESS_REG_5__SCAN_IN), .ZN(n18581) );
  INV_X1 U19342 ( .A(P2_ADDRESS_REG_5__SCAN_IN), .ZN(n19691) );
  AOI22_X1 U19343 ( .A1(n16337), .A2(n18581), .B1(n19691), .B2(n16338), .ZN(
        U351) );
  INV_X1 U19344 ( .A(P3_ADDRESS_REG_4__SCAN_IN), .ZN(n18579) );
  INV_X1 U19345 ( .A(P2_ADDRESS_REG_4__SCAN_IN), .ZN(n19690) );
  AOI22_X1 U19346 ( .A1(n16337), .A2(n18579), .B1(n19690), .B2(n16338), .ZN(
        U352) );
  INV_X1 U19347 ( .A(P3_ADDRESS_REG_3__SCAN_IN), .ZN(n18577) );
  INV_X1 U19348 ( .A(P2_ADDRESS_REG_3__SCAN_IN), .ZN(n19689) );
  AOI22_X1 U19349 ( .A1(n16339), .A2(n18577), .B1(n19689), .B2(n16338), .ZN(
        U353) );
  INV_X1 U19350 ( .A(P3_ADDRESS_REG_2__SCAN_IN), .ZN(n18575) );
  AOI22_X1 U19351 ( .A1(n16337), .A2(n18575), .B1(n19687), .B2(n16338), .ZN(
        U354) );
  INV_X1 U19352 ( .A(P3_ADDRESS_REG_29__SCAN_IN), .ZN(n18629) );
  INV_X1 U19353 ( .A(P2_ADDRESS_REG_29__SCAN_IN), .ZN(n19734) );
  AOI22_X1 U19354 ( .A1(n16337), .A2(n18629), .B1(n19734), .B2(n16338), .ZN(
        U355) );
  INV_X1 U19355 ( .A(P3_ADDRESS_REG_28__SCAN_IN), .ZN(n18627) );
  INV_X1 U19356 ( .A(P2_ADDRESS_REG_28__SCAN_IN), .ZN(n19732) );
  AOI22_X1 U19357 ( .A1(n16337), .A2(n18627), .B1(n19732), .B2(n16338), .ZN(
        U356) );
  INV_X1 U19358 ( .A(P3_ADDRESS_REG_27__SCAN_IN), .ZN(n18625) );
  INV_X1 U19359 ( .A(P2_ADDRESS_REG_27__SCAN_IN), .ZN(n19730) );
  AOI22_X1 U19360 ( .A1(n16337), .A2(n18625), .B1(n19730), .B2(n16338), .ZN(
        U357) );
  INV_X1 U19361 ( .A(P3_ADDRESS_REG_26__SCAN_IN), .ZN(n18624) );
  INV_X1 U19362 ( .A(P2_ADDRESS_REG_26__SCAN_IN), .ZN(n19727) );
  AOI22_X1 U19363 ( .A1(n16337), .A2(n18624), .B1(n19727), .B2(n16338), .ZN(
        U358) );
  INV_X1 U19364 ( .A(P3_ADDRESS_REG_25__SCAN_IN), .ZN(n18621) );
  INV_X1 U19365 ( .A(P2_ADDRESS_REG_25__SCAN_IN), .ZN(n19726) );
  AOI22_X1 U19366 ( .A1(n16337), .A2(n18621), .B1(n19726), .B2(n16338), .ZN(
        U359) );
  INV_X1 U19367 ( .A(P3_ADDRESS_REG_24__SCAN_IN), .ZN(n18619) );
  INV_X1 U19368 ( .A(P2_ADDRESS_REG_24__SCAN_IN), .ZN(n19725) );
  AOI22_X1 U19369 ( .A1(n16337), .A2(n18619), .B1(n19725), .B2(n16338), .ZN(
        U360) );
  INV_X1 U19370 ( .A(P3_ADDRESS_REG_23__SCAN_IN), .ZN(n18617) );
  INV_X1 U19371 ( .A(P2_ADDRESS_REG_23__SCAN_IN), .ZN(n19723) );
  AOI22_X1 U19372 ( .A1(n16337), .A2(n18617), .B1(n19723), .B2(n16338), .ZN(
        U361) );
  INV_X1 U19373 ( .A(P3_ADDRESS_REG_22__SCAN_IN), .ZN(n18614) );
  INV_X1 U19374 ( .A(P2_ADDRESS_REG_22__SCAN_IN), .ZN(n19721) );
  AOI22_X1 U19375 ( .A1(n16337), .A2(n18614), .B1(n19721), .B2(n16338), .ZN(
        U362) );
  INV_X1 U19376 ( .A(P3_ADDRESS_REG_21__SCAN_IN), .ZN(n18613) );
  INV_X1 U19377 ( .A(P2_ADDRESS_REG_21__SCAN_IN), .ZN(n19720) );
  AOI22_X1 U19378 ( .A1(n16337), .A2(n18613), .B1(n19720), .B2(n16338), .ZN(
        U363) );
  INV_X1 U19379 ( .A(P3_ADDRESS_REG_20__SCAN_IN), .ZN(n18610) );
  INV_X1 U19380 ( .A(P2_ADDRESS_REG_20__SCAN_IN), .ZN(n19718) );
  AOI22_X1 U19381 ( .A1(n16337), .A2(n18610), .B1(n19718), .B2(n16338), .ZN(
        U364) );
  INV_X1 U19382 ( .A(P3_ADDRESS_REG_1__SCAN_IN), .ZN(n18573) );
  INV_X1 U19383 ( .A(P2_ADDRESS_REG_1__SCAN_IN), .ZN(n19686) );
  AOI22_X1 U19384 ( .A1(n16337), .A2(n18573), .B1(n19686), .B2(n16338), .ZN(
        U365) );
  INV_X1 U19385 ( .A(P3_ADDRESS_REG_19__SCAN_IN), .ZN(n18609) );
  INV_X1 U19386 ( .A(P2_ADDRESS_REG_19__SCAN_IN), .ZN(n19716) );
  AOI22_X1 U19387 ( .A1(n16337), .A2(n18609), .B1(n19716), .B2(n16338), .ZN(
        U366) );
  INV_X1 U19388 ( .A(P3_ADDRESS_REG_18__SCAN_IN), .ZN(n18606) );
  INV_X1 U19389 ( .A(P2_ADDRESS_REG_18__SCAN_IN), .ZN(n19714) );
  AOI22_X1 U19390 ( .A1(n16337), .A2(n18606), .B1(n19714), .B2(n16338), .ZN(
        U367) );
  INV_X1 U19391 ( .A(P3_ADDRESS_REG_17__SCAN_IN), .ZN(n18605) );
  INV_X1 U19392 ( .A(P2_ADDRESS_REG_17__SCAN_IN), .ZN(n19712) );
  AOI22_X1 U19393 ( .A1(n16337), .A2(n18605), .B1(n19712), .B2(n16338), .ZN(
        U368) );
  INV_X1 U19394 ( .A(P3_ADDRESS_REG_16__SCAN_IN), .ZN(n18603) );
  INV_X1 U19395 ( .A(P2_ADDRESS_REG_16__SCAN_IN), .ZN(n19710) );
  AOI22_X1 U19396 ( .A1(n16337), .A2(n18603), .B1(n19710), .B2(n16338), .ZN(
        U369) );
  INV_X1 U19397 ( .A(P3_ADDRESS_REG_15__SCAN_IN), .ZN(n18601) );
  INV_X1 U19398 ( .A(P2_ADDRESS_REG_15__SCAN_IN), .ZN(n19708) );
  AOI22_X1 U19399 ( .A1(n16337), .A2(n18601), .B1(n19708), .B2(n16338), .ZN(
        U370) );
  INV_X1 U19400 ( .A(P3_ADDRESS_REG_14__SCAN_IN), .ZN(n18599) );
  INV_X1 U19401 ( .A(P2_ADDRESS_REG_14__SCAN_IN), .ZN(n19706) );
  AOI22_X1 U19402 ( .A1(n16339), .A2(n18599), .B1(n19706), .B2(n16338), .ZN(
        U371) );
  INV_X1 U19403 ( .A(P3_ADDRESS_REG_13__SCAN_IN), .ZN(n18596) );
  INV_X1 U19404 ( .A(P2_ADDRESS_REG_13__SCAN_IN), .ZN(n20739) );
  AOI22_X1 U19405 ( .A1(n16339), .A2(n18596), .B1(n20739), .B2(n16338), .ZN(
        U372) );
  INV_X1 U19406 ( .A(P3_ADDRESS_REG_12__SCAN_IN), .ZN(n18595) );
  INV_X1 U19407 ( .A(P2_ADDRESS_REG_12__SCAN_IN), .ZN(n19704) );
  AOI22_X1 U19408 ( .A1(n16339), .A2(n18595), .B1(n19704), .B2(n16338), .ZN(
        U373) );
  INV_X1 U19409 ( .A(P3_ADDRESS_REG_11__SCAN_IN), .ZN(n18593) );
  INV_X1 U19410 ( .A(P2_ADDRESS_REG_11__SCAN_IN), .ZN(n19702) );
  AOI22_X1 U19411 ( .A1(n16339), .A2(n18593), .B1(n19702), .B2(n16338), .ZN(
        U374) );
  INV_X1 U19412 ( .A(P3_ADDRESS_REG_10__SCAN_IN), .ZN(n18591) );
  INV_X1 U19413 ( .A(P2_ADDRESS_REG_10__SCAN_IN), .ZN(n19700) );
  AOI22_X1 U19414 ( .A1(n16339), .A2(n18591), .B1(n19700), .B2(n16338), .ZN(
        U375) );
  INV_X1 U19415 ( .A(P3_ADDRESS_REG_0__SCAN_IN), .ZN(n18571) );
  INV_X1 U19416 ( .A(P2_ADDRESS_REG_0__SCAN_IN), .ZN(n19684) );
  AOI22_X1 U19417 ( .A1(n16339), .A2(n18571), .B1(n19684), .B2(n16338), .ZN(
        U376) );
  INV_X1 U19418 ( .A(P3_ADS_N_REG_SCAN_IN), .ZN(n16341) );
  INV_X1 U19419 ( .A(P3_STATE_REG_2__SCAN_IN), .ZN(n18570) );
  NAND3_X1 U19420 ( .A1(n18570), .A2(P3_STATE_REG_0__SCAN_IN), .A3(
        P3_STATE_REG_1__SCAN_IN), .ZN(n16340) );
  NAND2_X1 U19421 ( .A1(n18567), .A2(n18559), .ZN(n18555) );
  NAND2_X1 U19422 ( .A1(n16340), .A2(n18555), .ZN(n18635) );
  INV_X1 U19423 ( .A(n18635), .ZN(n18633) );
  OAI21_X1 U19424 ( .B1(n18567), .B2(n16341), .A(n18633), .ZN(P3_U2633) );
  NAND2_X1 U19425 ( .A1(n18704), .A2(n18639), .ZN(n16343) );
  NAND2_X1 U19426 ( .A1(n18686), .A2(n18482), .ZN(n17289) );
  OAI21_X1 U19427 ( .B1(n16348), .B2(n17289), .A(P3_CODEFETCH_REG_SCAN_IN), 
        .ZN(n16342) );
  OAI21_X1 U19428 ( .B1(n16343), .B2(n18543), .A(n16342), .ZN(P3_U2634) );
  AOI221_X1 U19429 ( .B1(P3_STATE_REG_1__SCAN_IN), .B2(n18567), .C1(n18570), 
        .C2(n18567), .A(P3_D_C_N_REG_SCAN_IN), .ZN(n16344) );
  AOI21_X1 U19430 ( .B1(P3_CODEFETCH_REG_SCAN_IN), .B2(n18703), .A(n16344), 
        .ZN(P3_U2635) );
  NOR2_X1 U19431 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(P3_STATE_REG_2__SCAN_IN), 
        .ZN(n16345) );
  OAI21_X1 U19432 ( .B1(n16345), .B2(BS16), .A(n18635), .ZN(n18634) );
  OAI21_X1 U19433 ( .B1(n18635), .B2(n18691), .A(n18634), .ZN(P3_U2636) );
  NOR3_X1 U19434 ( .A1(n16348), .A2(n16347), .A3(n16346), .ZN(n18530) );
  NOR2_X1 U19435 ( .A1(n18530), .A2(n18534), .ZN(n18681) );
  OAI21_X1 U19436 ( .B1(n18681), .B2(n16350), .A(n16349), .ZN(P3_U2637) );
  INV_X1 U19437 ( .A(P3_REIP_REG_1__SCAN_IN), .ZN(n18679) );
  NOR4_X1 U19438 ( .A1(P3_DATAWIDTH_REG_12__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_13__SCAN_IN), .A3(P3_DATAWIDTH_REG_14__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_15__SCAN_IN), .ZN(n16360) );
  NOR4_X1 U19439 ( .A1(P3_DATAWIDTH_REG_8__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_9__SCAN_IN), .A3(P3_DATAWIDTH_REG_10__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_11__SCAN_IN), .ZN(n16359) );
  INV_X1 U19440 ( .A(P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(n20823) );
  INV_X1 U19441 ( .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(n18671) );
  NOR4_X1 U19442 ( .A1(P3_DATAWIDTH_REG_3__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_4__SCAN_IN), .A3(P3_DATAWIDTH_REG_5__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_7__SCAN_IN), .ZN(n16351) );
  OAI21_X1 U19443 ( .B1(n20823), .B2(n18671), .A(n16351), .ZN(n16357) );
  NOR4_X1 U19444 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_21__SCAN_IN), .A3(P3_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_23__SCAN_IN), .ZN(n16355) );
  NOR4_X1 U19445 ( .A1(P3_DATAWIDTH_REG_16__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_17__SCAN_IN), .A3(P3_DATAWIDTH_REG_18__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_19__SCAN_IN), .ZN(n16354) );
  NOR4_X1 U19446 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_29__SCAN_IN), .A3(P3_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_31__SCAN_IN), .ZN(n16353) );
  NOR4_X1 U19447 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_25__SCAN_IN), .A3(P3_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_27__SCAN_IN), .ZN(n16352) );
  NAND4_X1 U19448 ( .A1(n16355), .A2(n16354), .A3(n16353), .A4(n16352), .ZN(
        n16356) );
  NOR4_X1 U19449 ( .A1(P3_DATAWIDTH_REG_6__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_2__SCAN_IN), .A3(n16357), .A4(n16356), .ZN(n16358) );
  NAND3_X1 U19450 ( .A1(n16360), .A2(n16359), .A3(n16358), .ZN(n18678) );
  INV_X1 U19451 ( .A(n18678), .ZN(n18676) );
  INV_X1 U19452 ( .A(P3_REIP_REG_0__SCAN_IN), .ZN(n18672) );
  NAND2_X1 U19453 ( .A1(n18676), .A2(n18672), .ZN(n18675) );
  NOR3_X1 U19454 ( .A1(P3_DATAWIDTH_REG_0__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_1__SCAN_IN), .A3(n18675), .ZN(n16362) );
  AOI21_X1 U19455 ( .B1(P3_BYTEENABLE_REG_1__SCAN_IN), .B2(n18678), .A(n16362), 
        .ZN(n16361) );
  OAI21_X1 U19456 ( .B1(n18679), .B2(n18678), .A(n16361), .ZN(P3_U2638) );
  NAND2_X1 U19457 ( .A1(n18676), .A2(n18679), .ZN(n18670) );
  AOI21_X1 U19458 ( .B1(P3_BYTEENABLE_REG_3__SCAN_IN), .B2(n18678), .A(n16362), 
        .ZN(n16363) );
  OAI21_X1 U19459 ( .B1(P3_DATAWIDTH_REG_1__SCAN_IN), .B2(n18670), .A(n16363), 
        .ZN(P3_U2639) );
  NAND2_X1 U19460 ( .A1(P3_STATE2_REG_3__SCAN_IN), .A2(n18704), .ZN(n18544) );
  NOR2_X1 U19461 ( .A1(n18543), .A2(n18544), .ZN(n18538) );
  NOR4_X4 U19462 ( .A1(n17971), .A2(n18707), .A3(n16697), .A4(n18538), .ZN(
        n16722) );
  OAI211_X1 U19463 ( .C1(n17291), .C2(n16364), .A(n18693), .B(n18691), .ZN(
        n16365) );
  INV_X1 U19464 ( .A(n16365), .ZN(n18536) );
  NAND2_X1 U19465 ( .A1(n18707), .A2(n17227), .ZN(n16368) );
  AOI211_X4 U19466 ( .C1(P3_EBX_REG_31__SCAN_IN), .C2(n17291), .A(n18536), .B(
        n16368), .ZN(n16754) );
  INV_X1 U19467 ( .A(P3_REIP_REG_30__SCAN_IN), .ZN(n18630) );
  INV_X1 U19468 ( .A(P3_REIP_REG_26__SCAN_IN), .ZN(n18620) );
  NOR2_X2 U19469 ( .A1(n16365), .A2(n16368), .ZN(n16735) );
  INV_X1 U19470 ( .A(P3_REIP_REG_23__SCAN_IN), .ZN(n18615) );
  INV_X1 U19471 ( .A(P3_REIP_REG_21__SCAN_IN), .ZN(n18611) );
  INV_X1 U19472 ( .A(P3_REIP_REG_14__SCAN_IN), .ZN(n18597) );
  INV_X1 U19473 ( .A(P3_REIP_REG_13__SCAN_IN), .ZN(n18594) );
  INV_X1 U19474 ( .A(P3_REIP_REG_11__SCAN_IN), .ZN(n18590) );
  INV_X1 U19475 ( .A(P3_REIP_REG_7__SCAN_IN), .ZN(n18582) );
  INV_X1 U19476 ( .A(P3_REIP_REG_6__SCAN_IN), .ZN(n18580) );
  INV_X1 U19477 ( .A(P3_REIP_REG_4__SCAN_IN), .ZN(n18576) );
  NAND3_X1 U19478 ( .A1(P3_REIP_REG_3__SCAN_IN), .A2(P3_REIP_REG_1__SCAN_IN), 
        .A3(P3_REIP_REG_2__SCAN_IN), .ZN(n16712) );
  NOR2_X1 U19479 ( .A1(n18576), .A2(n16712), .ZN(n16680) );
  NAND2_X1 U19480 ( .A1(P3_REIP_REG_5__SCAN_IN), .A2(n16680), .ZN(n16653) );
  NOR3_X1 U19481 ( .A1(n18582), .A2(n18580), .A3(n16653), .ZN(n16642) );
  NAND2_X1 U19482 ( .A1(P3_REIP_REG_8__SCAN_IN), .A2(n16642), .ZN(n16618) );
  NAND2_X1 U19483 ( .A1(P3_REIP_REG_10__SCAN_IN), .A2(P3_REIP_REG_9__SCAN_IN), 
        .ZN(n16619) );
  NOR3_X1 U19484 ( .A1(n18590), .A2(n16618), .A3(n16619), .ZN(n16579) );
  NAND2_X1 U19485 ( .A1(P3_REIP_REG_12__SCAN_IN), .A2(n16579), .ZN(n16567) );
  NOR3_X1 U19486 ( .A1(n18597), .A2(n18594), .A3(n16567), .ZN(n16510) );
  INV_X1 U19487 ( .A(P3_REIP_REG_17__SCAN_IN), .ZN(n18602) );
  INV_X1 U19488 ( .A(P3_REIP_REG_16__SCAN_IN), .ZN(n18600) );
  INV_X1 U19489 ( .A(P3_REIP_REG_15__SCAN_IN), .ZN(n18598) );
  NOR3_X1 U19490 ( .A1(n18602), .A2(n18600), .A3(n18598), .ZN(n16511) );
  INV_X1 U19491 ( .A(P3_REIP_REG_19__SCAN_IN), .ZN(n18607) );
  INV_X1 U19492 ( .A(P3_REIP_REG_18__SCAN_IN), .ZN(n18604) );
  NOR2_X1 U19493 ( .A1(n18607), .A2(n18604), .ZN(n16512) );
  NAND4_X1 U19494 ( .A1(P3_REIP_REG_20__SCAN_IN), .A2(n16510), .A3(n16511), 
        .A4(n16512), .ZN(n16491) );
  NOR2_X1 U19495 ( .A1(n18611), .A2(n16491), .ZN(n16484) );
  NAND2_X1 U19496 ( .A1(P3_REIP_REG_22__SCAN_IN), .A2(n16484), .ZN(n16470) );
  NOR2_X1 U19497 ( .A1(n18615), .A2(n16470), .ZN(n16468) );
  NAND2_X1 U19498 ( .A1(P3_REIP_REG_24__SCAN_IN), .A2(n16468), .ZN(n16382) );
  NOR2_X1 U19499 ( .A1(n16744), .A2(n16382), .ZN(n16448) );
  NAND2_X1 U19500 ( .A1(P3_REIP_REG_25__SCAN_IN), .A2(n16448), .ZN(n16439) );
  NOR2_X1 U19501 ( .A1(n18620), .A2(n16439), .ZN(n16414) );
  NAND4_X1 U19502 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_29__SCAN_IN), 
        .A3(P3_REIP_REG_27__SCAN_IN), .A4(n16414), .ZN(n16385) );
  NOR3_X1 U19503 ( .A1(P3_REIP_REG_31__SCAN_IN), .A2(n18630), .A3(n16385), 
        .ZN(n16366) );
  AOI21_X1 U19504 ( .B1(n16754), .B2(P3_EBX_REG_31__SCAN_IN), .A(n16366), .ZN(
        n16390) );
  NAND2_X1 U19505 ( .A1(P3_EBX_REG_31__SCAN_IN), .A2(n17291), .ZN(n16367) );
  AOI211_X4 U19506 ( .C1(n18691), .C2(n18693), .A(n16368), .B(n16367), .ZN(
        n16753) );
  NOR3_X1 U19507 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .A3(P3_EBX_REG_2__SCAN_IN), .ZN(n16724) );
  INV_X1 U19508 ( .A(P3_EBX_REG_3__SCAN_IN), .ZN(n17050) );
  NAND2_X1 U19509 ( .A1(n16724), .A2(n17050), .ZN(n16718) );
  NOR2_X1 U19510 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(n16718), .ZN(n16692) );
  INV_X1 U19511 ( .A(P3_EBX_REG_5__SCAN_IN), .ZN(n17040) );
  NAND2_X1 U19512 ( .A1(n16692), .A2(n17040), .ZN(n16684) );
  NOR2_X1 U19513 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(n16684), .ZN(n16669) );
  INV_X1 U19514 ( .A(P3_EBX_REG_7__SCAN_IN), .ZN(n16660) );
  NAND2_X1 U19515 ( .A1(n16669), .A2(n16660), .ZN(n16659) );
  NOR2_X1 U19516 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n16659), .ZN(n16641) );
  NAND2_X1 U19517 ( .A1(n16641), .A2(n16640), .ZN(n16637) );
  NOR2_X1 U19518 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n16637), .ZN(n16617) );
  INV_X1 U19519 ( .A(P3_EBX_REG_11__SCAN_IN), .ZN(n16613) );
  NAND2_X1 U19520 ( .A1(n16617), .A2(n16613), .ZN(n16612) );
  NOR2_X1 U19521 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n16612), .ZN(n16594) );
  NAND2_X1 U19522 ( .A1(n16594), .A2(n16593), .ZN(n16590) );
  NOR2_X1 U19523 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n16590), .ZN(n16566) );
  NAND2_X1 U19524 ( .A1(n16566), .A2(n16563), .ZN(n16562) );
  NOR2_X1 U19525 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n16562), .ZN(n16543) );
  NAND2_X1 U19526 ( .A1(n16543), .A2(n16904), .ZN(n16540) );
  NOR2_X1 U19527 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n16540), .ZN(n16523) );
  INV_X1 U19528 ( .A(P3_EBX_REG_19__SCAN_IN), .ZN(n16875) );
  NAND2_X1 U19529 ( .A1(n16523), .A2(n16875), .ZN(n16519) );
  NOR2_X1 U19530 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n16519), .ZN(n16501) );
  INV_X1 U19531 ( .A(P3_EBX_REG_21__SCAN_IN), .ZN(n16849) );
  NAND2_X1 U19532 ( .A1(n16501), .A2(n16849), .ZN(n16489) );
  NOR2_X1 U19533 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(n16489), .ZN(n16478) );
  INV_X1 U19534 ( .A(P3_EBX_REG_23__SCAN_IN), .ZN(n16759) );
  NAND2_X1 U19535 ( .A1(n16478), .A2(n16759), .ZN(n16474) );
  NOR2_X1 U19536 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(n16474), .ZN(n16456) );
  INV_X1 U19537 ( .A(P3_EBX_REG_25__SCAN_IN), .ZN(n16451) );
  NAND2_X1 U19538 ( .A1(n16456), .A2(n16451), .ZN(n16450) );
  NOR2_X1 U19539 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n16450), .ZN(n16434) );
  INV_X1 U19540 ( .A(P3_EBX_REG_27__SCAN_IN), .ZN(n16430) );
  NAND2_X1 U19541 ( .A1(n16434), .A2(n16430), .ZN(n16429) );
  NOR2_X1 U19542 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n16429), .ZN(n16415) );
  INV_X1 U19543 ( .A(P3_EBX_REG_29__SCAN_IN), .ZN(n16401) );
  NAND2_X1 U19544 ( .A1(n16415), .A2(n16401), .ZN(n16392) );
  NOR2_X1 U19545 ( .A1(n16723), .A2(n16392), .ZN(n16398) );
  INV_X1 U19546 ( .A(P3_EBX_REG_30__SCAN_IN), .ZN(n16764) );
  INV_X1 U19547 ( .A(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n16371) );
  INV_X1 U19548 ( .A(n16369), .ZN(n17357) );
  NAND2_X1 U19549 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17389), .ZN(
        n16376) );
  NOR2_X1 U19550 ( .A1(n17357), .A2(n16376), .ZN(n16373) );
  NAND2_X1 U19551 ( .A1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n16373), .ZN(
        n16372) );
  AOI21_X1 U19552 ( .B1(n16371), .B2(n16372), .A(n16370), .ZN(n17342) );
  OAI21_X1 U19553 ( .B1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n16373), .A(
        n16372), .ZN(n17366) );
  INV_X1 U19554 ( .A(n17366), .ZN(n16426) );
  NOR2_X1 U19555 ( .A1(n17391), .A2(n16376), .ZN(n17340) );
  INV_X1 U19556 ( .A(n17340), .ZN(n16374) );
  AOI21_X1 U19557 ( .B1(n17380), .B2(n16374), .A(n16373), .ZN(n17382) );
  INV_X1 U19558 ( .A(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n16463) );
  NOR2_X1 U19559 ( .A1(n16463), .A2(n16376), .ZN(n16375) );
  OAI21_X1 U19560 ( .B1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n16375), .A(
        n16374), .ZN(n17393) );
  INV_X1 U19561 ( .A(n17393), .ZN(n16446) );
  AOI21_X1 U19562 ( .B1(n16463), .B2(n16376), .A(n16375), .ZN(n17402) );
  NOR2_X1 U19563 ( .A1(n16693), .A2(n17415), .ZN(n17388) );
  OAI21_X1 U19564 ( .B1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n17388), .A(
        n16376), .ZN(n17419) );
  INV_X1 U19565 ( .A(n17419), .ZN(n16467) );
  INV_X1 U19566 ( .A(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n17429) );
  INV_X1 U19567 ( .A(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n17430) );
  NAND2_X1 U19568 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17428), .ZN(
        n16378) );
  OR2_X1 U19569 ( .A1(n17430), .A2(n16378), .ZN(n16377) );
  AOI21_X1 U19570 ( .B1(n17429), .B2(n16377), .A(n17388), .ZN(n17431) );
  XOR2_X1 U19571 ( .A(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .B(n16378), .Z(
        n17441) );
  INV_X1 U19572 ( .A(n17441), .ZN(n16494) );
  NAND2_X1 U19573 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n17467) );
  NOR2_X1 U19574 ( .A1(n16693), .A2(n17489), .ZN(n16545) );
  NAND2_X1 U19575 ( .A1(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .A2(n16545), .ZN(
        n16533) );
  NOR2_X1 U19576 ( .A1(n17467), .A2(n16533), .ZN(n17425) );
  OAI21_X1 U19577 ( .B1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n17425), .A(
        n16378), .ZN(n16379) );
  INV_X1 U19578 ( .A(n16379), .ZN(n17458) );
  INV_X1 U19579 ( .A(n17454), .ZN(n16380) );
  NOR2_X1 U19580 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n16693), .ZN(
        n16727) );
  NOR2_X1 U19581 ( .A1(n16492), .A2(n16679), .ZN(n16480) );
  NOR2_X1 U19582 ( .A1(n17402), .A2(n16458), .ZN(n16457) );
  NOR2_X1 U19583 ( .A1(n16457), .A2(n16679), .ZN(n16445) );
  NOR2_X1 U19584 ( .A1(n16424), .A2(n16679), .ZN(n16417) );
  NOR2_X1 U19585 ( .A1(n16416), .A2(n16679), .ZN(n16403) );
  NAND2_X1 U19586 ( .A1(n10006), .A2(n16697), .ZN(n16730) );
  NOR3_X1 U19587 ( .A1(n16394), .A2(n16393), .A3(n16730), .ZN(n16388) );
  NAND3_X1 U19588 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_29__SCAN_IN), 
        .A3(P3_REIP_REG_27__SCAN_IN), .ZN(n16384) );
  NOR2_X1 U19589 ( .A1(n16722), .A2(n16382), .ZN(n16443) );
  INV_X1 U19590 ( .A(P3_REIP_REG_25__SCAN_IN), .ZN(n18618) );
  NOR2_X1 U19591 ( .A1(n18620), .A2(n18618), .ZN(n16383) );
  NOR2_X1 U19592 ( .A1(n16735), .A2(n16722), .ZN(n16681) );
  AOI21_X1 U19593 ( .B1(n16443), .B2(n16383), .A(n16681), .ZN(n16413) );
  AOI21_X1 U19594 ( .B1(n16735), .B2(n16384), .A(n16413), .ZN(n16406) );
  NOR2_X1 U19595 ( .A1(P3_REIP_REG_30__SCAN_IN), .A2(n16385), .ZN(n16397) );
  INV_X1 U19596 ( .A(n16397), .ZN(n16386) );
  AOI21_X1 U19597 ( .B1(n16406), .B2(n16386), .A(n18628), .ZN(n16387) );
  AOI211_X1 U19598 ( .C1(n16398), .C2(n16764), .A(n16388), .B(n16387), .ZN(
        n16389) );
  OAI211_X1 U19599 ( .C1(n16391), .C2(n16739), .A(n16390), .B(n16389), .ZN(
        P3_U2640) );
  NAND2_X1 U19600 ( .A1(n16753), .A2(n16392), .ZN(n16411) );
  OAI22_X1 U19601 ( .A1(n16406), .A2(n18630), .B1(n16395), .B2(n16739), .ZN(
        n16396) );
  OAI21_X1 U19602 ( .B1(n16754), .B2(n16398), .A(P3_EBX_REG_30__SCAN_IN), .ZN(
        n16399) );
  OAI211_X1 U19603 ( .C1(P3_EBX_REG_30__SCAN_IN), .C2(n16411), .A(n16400), .B(
        n16399), .ZN(P3_U2641) );
  NOR2_X1 U19604 ( .A1(n16415), .A2(n16401), .ZN(n16412) );
  INV_X1 U19605 ( .A(n16697), .ZN(n18549) );
  AOI211_X1 U19606 ( .C1(n16404), .C2(n16403), .A(n16402), .B(n18549), .ZN(
        n16408) );
  INV_X1 U19607 ( .A(P3_REIP_REG_29__SCAN_IN), .ZN(n20840) );
  OAI22_X1 U19608 ( .A1(n16406), .A2(n20840), .B1(n16405), .B2(n16739), .ZN(
        n16407) );
  AOI211_X1 U19609 ( .C1(P3_EBX_REG_29__SCAN_IN), .C2(n16754), .A(n16408), .B(
        n16407), .ZN(n16410) );
  NAND4_X1 U19610 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_27__SCAN_IN), 
        .A3(n16414), .A4(n20840), .ZN(n16409) );
  OAI211_X1 U19611 ( .C1(n16412), .C2(n16411), .A(n16410), .B(n16409), .ZN(
        P3_U2642) );
  NAND2_X1 U19612 ( .A1(P3_REIP_REG_27__SCAN_IN), .A2(n16414), .ZN(n16423) );
  AOI22_X1 U19613 ( .A1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n16691), .B1(
        n16754), .B2(P3_EBX_REG_28__SCAN_IN), .ZN(n16422) );
  INV_X1 U19614 ( .A(n16413), .ZN(n16438) );
  INV_X1 U19615 ( .A(P3_REIP_REG_27__SCAN_IN), .ZN(n18623) );
  NAND2_X1 U19616 ( .A1(n16414), .A2(n18623), .ZN(n16432) );
  NAND2_X1 U19617 ( .A1(n16438), .A2(n16432), .ZN(n16420) );
  AOI211_X1 U19618 ( .C1(P3_EBX_REG_28__SCAN_IN), .C2(n16429), .A(n16415), .B(
        n16723), .ZN(n16419) );
  AOI211_X1 U19619 ( .C1(n17342), .C2(n16417), .A(n16416), .B(n18549), .ZN(
        n16418) );
  AOI211_X1 U19620 ( .C1(P3_REIP_REG_28__SCAN_IN), .C2(n16420), .A(n16419), 
        .B(n16418), .ZN(n16421) );
  OAI211_X1 U19621 ( .C1(P3_REIP_REG_28__SCAN_IN), .C2(n16423), .A(n16422), 
        .B(n16421), .ZN(P3_U2643) );
  AOI211_X1 U19622 ( .C1(n16426), .C2(n16425), .A(n16424), .B(n18549), .ZN(
        n16428) );
  INV_X1 U19623 ( .A(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n17369) );
  OAI22_X1 U19624 ( .A1(n17369), .A2(n16739), .B1(n18623), .B2(n16438), .ZN(
        n16427) );
  AOI211_X1 U19625 ( .C1(P3_EBX_REG_27__SCAN_IN), .C2(n16754), .A(n16428), .B(
        n16427), .ZN(n16433) );
  OAI211_X1 U19626 ( .C1(n16434), .C2(n16430), .A(n16753), .B(n16429), .ZN(
        n16431) );
  NAND3_X1 U19627 ( .A1(n16433), .A2(n16432), .A3(n16431), .ZN(P3_U2644) );
  AOI211_X1 U19628 ( .C1(P3_EBX_REG_26__SCAN_IN), .C2(n16450), .A(n16434), .B(
        n16723), .ZN(n16442) );
  AOI211_X1 U19629 ( .C1(n17382), .C2(n16436), .A(n16435), .B(n18549), .ZN(
        n16441) );
  AOI22_X1 U19630 ( .A1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n16691), .B1(
        n16754), .B2(P3_EBX_REG_26__SCAN_IN), .ZN(n16437) );
  OAI221_X1 U19631 ( .B1(P3_REIP_REG_26__SCAN_IN), .B2(n16439), .C1(n18620), 
        .C2(n16438), .A(n16437), .ZN(n16440) );
  OR3_X1 U19632 ( .A1(n16442), .A2(n16441), .A3(n16440), .ZN(P3_U2645) );
  AOI22_X1 U19633 ( .A1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n16691), .B1(
        n16754), .B2(P3_EBX_REG_25__SCAN_IN), .ZN(n16454) );
  NOR2_X1 U19634 ( .A1(n16681), .A2(n16443), .ZN(n16449) );
  AOI211_X1 U19635 ( .C1(n16446), .C2(n16445), .A(n16444), .B(n18549), .ZN(
        n16447) );
  AOI221_X1 U19636 ( .B1(n16449), .B2(P3_REIP_REG_25__SCAN_IN), .C1(n16448), 
        .C2(n18618), .A(n16447), .ZN(n16453) );
  OAI211_X1 U19637 ( .C1(n16456), .C2(n16451), .A(n16753), .B(n16450), .ZN(
        n16452) );
  NAND3_X1 U19638 ( .A1(n16454), .A2(n16453), .A3(n16452), .ZN(P3_U2646) );
  NOR2_X1 U19639 ( .A1(P3_REIP_REG_24__SCAN_IN), .A2(n16744), .ZN(n16455) );
  AOI22_X1 U19640 ( .A1(n16754), .A2(P3_EBX_REG_24__SCAN_IN), .B1(n16468), 
        .B2(n16455), .ZN(n16462) );
  OAI21_X1 U19641 ( .B1(n16468), .B2(n16744), .A(n16752), .ZN(n16464) );
  AOI211_X1 U19642 ( .C1(P3_EBX_REG_24__SCAN_IN), .C2(n16474), .A(n16456), .B(
        n16723), .ZN(n16460) );
  AOI211_X1 U19643 ( .C1(n17402), .C2(n16458), .A(n16457), .B(n18549), .ZN(
        n16459) );
  AOI211_X1 U19644 ( .C1(P3_REIP_REG_24__SCAN_IN), .C2(n16464), .A(n16460), 
        .B(n16459), .ZN(n16461) );
  OAI211_X1 U19645 ( .C1(n16463), .C2(n16739), .A(n16462), .B(n16461), .ZN(
        P3_U2647) );
  INV_X1 U19646 ( .A(n16464), .ZN(n16477) );
  AOI211_X1 U19647 ( .C1(n16467), .C2(n16466), .A(n16465), .B(n18549), .ZN(
        n16473) );
  OR2_X1 U19648 ( .A1(n16744), .A2(n16468), .ZN(n16469) );
  OAI22_X1 U19649 ( .A1(n16471), .A2(n16739), .B1(n16470), .B2(n16469), .ZN(
        n16472) );
  AOI211_X1 U19650 ( .C1(P3_EBX_REG_23__SCAN_IN), .C2(n16754), .A(n16473), .B(
        n16472), .ZN(n16476) );
  OAI211_X1 U19651 ( .C1(n16478), .C2(n16759), .A(n16753), .B(n16474), .ZN(
        n16475) );
  OAI211_X1 U19652 ( .C1(n16477), .C2(n18615), .A(n16476), .B(n16475), .ZN(
        P3_U2648) );
  AOI221_X1 U19653 ( .B1(n18611), .B2(n16735), .C1(n16491), .C2(n16735), .A(
        n16722), .ZN(n16487) );
  INV_X1 U19654 ( .A(P3_REIP_REG_22__SCAN_IN), .ZN(n18612) );
  AOI22_X1 U19655 ( .A1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n16691), .B1(
        n16754), .B2(P3_EBX_REG_22__SCAN_IN), .ZN(n16486) );
  NOR2_X1 U19656 ( .A1(P3_REIP_REG_22__SCAN_IN), .A2(n16744), .ZN(n16483) );
  AOI211_X1 U19657 ( .C1(P3_EBX_REG_22__SCAN_IN), .C2(n16489), .A(n16478), .B(
        n16723), .ZN(n16482) );
  AOI211_X1 U19658 ( .C1(n17431), .C2(n16480), .A(n16479), .B(n18549), .ZN(
        n16481) );
  AOI211_X1 U19659 ( .C1(n16484), .C2(n16483), .A(n16482), .B(n16481), .ZN(
        n16485) );
  OAI211_X1 U19660 ( .C1(n16487), .C2(n18612), .A(n16486), .B(n16485), .ZN(
        P3_U2649) );
  AOI21_X1 U19661 ( .B1(n16735), .B2(n16491), .A(n16722), .ZN(n16508) );
  INV_X1 U19662 ( .A(n16501), .ZN(n16488) );
  AOI21_X1 U19663 ( .B1(P3_EBX_REG_21__SCAN_IN), .B2(n16488), .A(n16723), .ZN(
        n16490) );
  AOI22_X1 U19664 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n16691), .B1(
        n16490), .B2(n16489), .ZN(n16498) );
  NOR3_X1 U19665 ( .A1(P3_REIP_REG_21__SCAN_IN), .A2(n16744), .A3(n16491), 
        .ZN(n16496) );
  AOI211_X1 U19666 ( .C1(n16494), .C2(n16493), .A(n16492), .B(n18549), .ZN(
        n16495) );
  AOI211_X1 U19667 ( .C1(P3_EBX_REG_21__SCAN_IN), .C2(n16754), .A(n16496), .B(
        n16495), .ZN(n16497) );
  OAI211_X1 U19668 ( .C1(n18611), .C2(n16508), .A(n16498), .B(n16497), .ZN(
        P3_U2650) );
  NAND2_X1 U19669 ( .A1(n16735), .A2(n16510), .ZN(n16553) );
  INV_X1 U19670 ( .A(n16553), .ZN(n16499) );
  NAND2_X1 U19671 ( .A1(n16511), .A2(n16499), .ZN(n16532) );
  INV_X1 U19672 ( .A(n16532), .ZN(n16500) );
  AOI21_X1 U19673 ( .B1(n16512), .B2(n16500), .A(P3_REIP_REG_20__SCAN_IN), 
        .ZN(n16509) );
  AOI22_X1 U19674 ( .A1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n16691), .B1(
        n16754), .B2(P3_EBX_REG_20__SCAN_IN), .ZN(n16507) );
  AOI211_X1 U19675 ( .C1(P3_EBX_REG_20__SCAN_IN), .C2(n16519), .A(n16501), .B(
        n16723), .ZN(n16505) );
  AOI211_X1 U19676 ( .C1(n17458), .C2(n16503), .A(n16502), .B(n18549), .ZN(
        n16504) );
  NOR2_X1 U19677 ( .A1(n16505), .A2(n16504), .ZN(n16506) );
  OAI211_X1 U19678 ( .C1(n16509), .C2(n16508), .A(n16507), .B(n16506), .ZN(
        P3_U2651) );
  INV_X1 U19679 ( .A(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n16522) );
  AND2_X1 U19680 ( .A1(n16752), .A2(n16510), .ZN(n16568) );
  AOI21_X1 U19681 ( .B1(n16511), .B2(n16568), .A(n16681), .ZN(n16539) );
  AOI211_X1 U19682 ( .C1(n18607), .C2(n18604), .A(n16512), .B(n16532), .ZN(
        n16518) );
  INV_X1 U19683 ( .A(n16533), .ZN(n17465) );
  NAND2_X1 U19684 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n17465), .ZN(
        n16524) );
  AOI21_X1 U19685 ( .B1(n16522), .B2(n16524), .A(n17425), .ZN(n16513) );
  INV_X1 U19686 ( .A(n16513), .ZN(n17469) );
  NAND2_X1 U19687 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17503), .ZN(
        n16573) );
  INV_X1 U19688 ( .A(n16573), .ZN(n17505) );
  NAND2_X1 U19689 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n17505), .ZN(
        n16554) );
  OR2_X1 U19690 ( .A1(n16554), .A2(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n16555) );
  OAI21_X1 U19691 ( .B1(n16524), .B2(n16555), .A(n10006), .ZN(n16515) );
  AOI21_X1 U19692 ( .B1(n17469), .B2(n16515), .A(n18549), .ZN(n16514) );
  OAI21_X1 U19693 ( .B1(n17469), .B2(n16515), .A(n16514), .ZN(n16516) );
  OAI211_X1 U19694 ( .C1(n16743), .C2(n16875), .A(n18028), .B(n16516), .ZN(
        n16517) );
  AOI211_X1 U19695 ( .C1(P3_REIP_REG_19__SCAN_IN), .C2(n16539), .A(n16518), 
        .B(n16517), .ZN(n16521) );
  OAI211_X1 U19696 ( .C1(n16523), .C2(n16875), .A(n16753), .B(n16519), .ZN(
        n16520) );
  OAI211_X1 U19697 ( .C1(n16739), .C2(n16522), .A(n16521), .B(n16520), .ZN(
        P3_U2652) );
  INV_X1 U19698 ( .A(n16539), .ZN(n16531) );
  AOI211_X1 U19699 ( .C1(P3_EBX_REG_18__SCAN_IN), .C2(n16540), .A(n16523), .B(
        n16723), .ZN(n16529) );
  OAI21_X1 U19700 ( .B1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n17465), .A(
        n16524), .ZN(n17478) );
  INV_X1 U19701 ( .A(n17466), .ZN(n17463) );
  INV_X1 U19702 ( .A(n16727), .ZN(n16696) );
  OAI21_X1 U19703 ( .B1(n17463), .B2(n16696), .A(n10006), .ZN(n16526) );
  AOI21_X1 U19704 ( .B1(n17478), .B2(n16526), .A(n18549), .ZN(n16525) );
  OAI21_X1 U19705 ( .B1(n17478), .B2(n16526), .A(n16525), .ZN(n16527) );
  OAI211_X1 U19706 ( .C1(n16743), .C2(n16888), .A(n18028), .B(n16527), .ZN(
        n16528) );
  AOI211_X1 U19707 ( .C1(n16691), .C2(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n16529), .B(n16528), .ZN(n16530) );
  OAI221_X1 U19708 ( .B1(P3_REIP_REG_18__SCAN_IN), .B2(n16532), .C1(n18604), 
        .C2(n16531), .A(n16530), .ZN(P3_U2653) );
  NOR3_X1 U19709 ( .A1(n18600), .A2(n18598), .A3(n16553), .ZN(n16538) );
  OAI21_X1 U19710 ( .B1(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n16545), .A(
        n16533), .ZN(n17493) );
  OAI21_X1 U19711 ( .B1(n17489), .B2(n16696), .A(n10006), .ZN(n16535) );
  AOI21_X1 U19712 ( .B1(n17493), .B2(n16535), .A(n18549), .ZN(n16534) );
  OAI21_X1 U19713 ( .B1(n17493), .B2(n16535), .A(n16534), .ZN(n16536) );
  OAI211_X1 U19714 ( .C1(n16743), .C2(n16904), .A(n18028), .B(n16536), .ZN(
        n16537) );
  AOI221_X1 U19715 ( .B1(n16539), .B2(P3_REIP_REG_17__SCAN_IN), .C1(n16538), 
        .C2(n18602), .A(n16537), .ZN(n16542) );
  OAI211_X1 U19716 ( .C1(n16543), .C2(n16904), .A(n16753), .B(n16540), .ZN(
        n16541) );
  OAI211_X1 U19717 ( .C1(n16739), .C2(n17490), .A(n16542), .B(n16541), .ZN(
        P3_U2654) );
  AOI211_X1 U19718 ( .C1(P3_EBX_REG_16__SCAN_IN), .C2(n16562), .A(n16543), .B(
        n16723), .ZN(n16544) );
  AOI21_X1 U19719 ( .B1(n16691), .B2(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A(
        n16544), .ZN(n16552) );
  INV_X1 U19720 ( .A(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n16546) );
  AOI21_X1 U19721 ( .B1(n16546), .B2(n16554), .A(n16545), .ZN(n17506) );
  NAND2_X1 U19722 ( .A1(n10006), .A2(n16555), .ZN(n16547) );
  XNOR2_X1 U19723 ( .A(n17506), .B(n16547), .ZN(n16548) );
  AOI22_X1 U19724 ( .A1(n16754), .A2(P3_EBX_REG_16__SCAN_IN), .B1(n16697), 
        .B2(n16548), .ZN(n16551) );
  AOI21_X1 U19725 ( .B1(P3_REIP_REG_15__SCAN_IN), .B2(n16568), .A(n16681), 
        .ZN(n16561) );
  NOR2_X1 U19726 ( .A1(n18598), .A2(n16553), .ZN(n16549) );
  AOI22_X1 U19727 ( .A1(P3_REIP_REG_16__SCAN_IN), .A2(n16561), .B1(n16549), 
        .B2(n18600), .ZN(n16550) );
  NAND4_X1 U19728 ( .A1(n16552), .A2(n16551), .A3(n16550), .A4(n18028), .ZN(
        P3_U2655) );
  INV_X1 U19729 ( .A(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n17521) );
  NAND2_X1 U19730 ( .A1(n18598), .A2(n16553), .ZN(n16560) );
  NAND2_X1 U19731 ( .A1(n16697), .A2(n16679), .ZN(n16728) );
  OAI21_X1 U19732 ( .B1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n17505), .A(
        n16554), .ZN(n17517) );
  AOI21_X1 U19733 ( .B1(n10006), .B2(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A(
        n18549), .ZN(n16584) );
  INV_X1 U19734 ( .A(n16584), .ZN(n16750) );
  AOI211_X1 U19735 ( .C1(n16573), .C2(n16728), .A(n17517), .B(n16750), .ZN(
        n16559) );
  INV_X1 U19736 ( .A(n16730), .ZN(n16556) );
  NAND3_X1 U19737 ( .A1(n16556), .A2(n17517), .A3(n16555), .ZN(n16557) );
  OAI211_X1 U19738 ( .C1(n16743), .C2(n16563), .A(n18028), .B(n16557), .ZN(
        n16558) );
  AOI211_X1 U19739 ( .C1(n16561), .C2(n16560), .A(n16559), .B(n16558), .ZN(
        n16565) );
  OAI211_X1 U19740 ( .C1(n16566), .C2(n16563), .A(n16753), .B(n16562), .ZN(
        n16564) );
  OAI211_X1 U19741 ( .C1(n16739), .C2(n17521), .A(n16565), .B(n16564), .ZN(
        P3_U2656) );
  AOI211_X1 U19742 ( .C1(P3_EBX_REG_14__SCAN_IN), .C2(n16590), .A(n16566), .B(
        n16723), .ZN(n16571) );
  OR2_X1 U19743 ( .A1(n16744), .A2(n16567), .ZN(n16586) );
  INV_X1 U19744 ( .A(n16681), .ZN(n16751) );
  NAND2_X1 U19745 ( .A1(P3_REIP_REG_14__SCAN_IN), .A2(n16751), .ZN(n16569) );
  AOI221_X1 U19746 ( .B1(n16586), .B2(n16569), .C1(n18594), .C2(n16569), .A(
        n16568), .ZN(n16570) );
  AOI211_X1 U19747 ( .C1(n16691), .C2(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .A(
        n16571), .B(n16570), .ZN(n16578) );
  INV_X1 U19748 ( .A(n17545), .ZN(n16572) );
  NAND2_X1 U19749 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17546), .ZN(
        n17548) );
  NOR2_X1 U19750 ( .A1(n16572), .A2(n17548), .ZN(n16580) );
  OAI21_X1 U19751 ( .B1(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n16580), .A(
        n16573), .ZN(n17533) );
  INV_X1 U19752 ( .A(n17533), .ZN(n16575) );
  OAI21_X1 U19753 ( .B1(n17508), .B2(n16696), .A(n10006), .ZN(n16597) );
  OAI21_X1 U19754 ( .B1(n17545), .B2(n16679), .A(n16597), .ZN(n16582) );
  INV_X1 U19755 ( .A(n16582), .ZN(n16574) );
  AOI221_X1 U19756 ( .B1(n16575), .B2(n16582), .C1(n17533), .C2(n16574), .A(
        n18549), .ZN(n16576) );
  AOI211_X1 U19757 ( .C1(n16754), .C2(P3_EBX_REG_14__SCAN_IN), .A(n17971), .B(
        n16576), .ZN(n16577) );
  NAND2_X1 U19758 ( .A1(n16578), .A2(n16577), .ZN(P3_U2657) );
  INV_X1 U19759 ( .A(n16579), .ZN(n16595) );
  AOI21_X1 U19760 ( .B1(n16735), .B2(n16595), .A(n16722), .ZN(n16609) );
  OAI21_X1 U19761 ( .B1(P3_REIP_REG_12__SCAN_IN), .B2(n16744), .A(n16609), 
        .ZN(n16589) );
  INV_X1 U19762 ( .A(n17548), .ZN(n16596) );
  NAND2_X1 U19763 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n16596), .ZN(
        n16581) );
  AOI21_X1 U19764 ( .B1(n17550), .B2(n16581), .A(n16580), .ZN(n17553) );
  NAND2_X1 U19765 ( .A1(n16697), .A2(n16582), .ZN(n16583) );
  OAI22_X1 U19766 ( .A1(n17553), .A2(n16583), .B1(n17550), .B2(n16739), .ZN(
        n16588) );
  OAI211_X1 U19767 ( .C1(n17550), .C2(n16679), .A(n17553), .B(n16584), .ZN(
        n16585) );
  OAI211_X1 U19768 ( .C1(P3_REIP_REG_13__SCAN_IN), .C2(n16586), .A(n18028), 
        .B(n16585), .ZN(n16587) );
  AOI211_X1 U19769 ( .C1(P3_REIP_REG_13__SCAN_IN), .C2(n16589), .A(n16588), 
        .B(n16587), .ZN(n16592) );
  OAI211_X1 U19770 ( .C1(n16594), .C2(n16593), .A(n16753), .B(n16590), .ZN(
        n16591) );
  OAI211_X1 U19771 ( .C1(n16593), .C2(n16743), .A(n16592), .B(n16591), .ZN(
        P3_U2658) );
  INV_X1 U19772 ( .A(P3_REIP_REG_12__SCAN_IN), .ZN(n18592) );
  AOI22_X1 U19773 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n16691), .B1(
        n16754), .B2(P3_EBX_REG_12__SCAN_IN), .ZN(n16604) );
  AOI211_X1 U19774 ( .C1(P3_EBX_REG_12__SCAN_IN), .C2(n16612), .A(n16594), .B(
        n16723), .ZN(n16602) );
  NOR3_X1 U19775 ( .A1(P3_REIP_REG_12__SCAN_IN), .A2(n16744), .A3(n16595), 
        .ZN(n16601) );
  AOI22_X1 U19776 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n16596), .B1(
        n17548), .B2(n17568), .ZN(n17564) );
  INV_X1 U19777 ( .A(n16597), .ZN(n16599) );
  INV_X1 U19778 ( .A(n17564), .ZN(n16598) );
  AOI221_X1 U19779 ( .B1(n17564), .B2(n16599), .C1(n16598), .C2(n16597), .A(
        n18549), .ZN(n16600) );
  NOR4_X1 U19780 ( .A1(n17971), .A2(n16602), .A3(n16601), .A4(n16600), .ZN(
        n16603) );
  OAI211_X1 U19781 ( .C1(n18592), .C2(n16609), .A(n16604), .B(n16603), .ZN(
        P3_U2659) );
  INV_X1 U19782 ( .A(n16619), .ZN(n16605) );
  NOR2_X1 U19783 ( .A1(n16744), .A2(n16618), .ZN(n16635) );
  AOI21_X1 U19784 ( .B1(n16605), .B2(n16635), .A(P3_REIP_REG_11__SCAN_IN), 
        .ZN(n16610) );
  NOR2_X1 U19785 ( .A1(n16693), .A2(n16606), .ZN(n16620) );
  OAI21_X1 U19786 ( .B1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n16620), .A(
        n17548), .ZN(n17577) );
  OAI21_X1 U19787 ( .B1(n16606), .B2(n16696), .A(n10006), .ZN(n16607) );
  XNOR2_X1 U19788 ( .A(n17577), .B(n16607), .ZN(n16608) );
  OAI22_X1 U19789 ( .A1(n16610), .A2(n16609), .B1(n18549), .B2(n16608), .ZN(
        n16611) );
  AOI211_X1 U19790 ( .C1(n16754), .C2(P3_EBX_REG_11__SCAN_IN), .A(n17971), .B(
        n16611), .ZN(n16615) );
  OAI211_X1 U19791 ( .C1(n16617), .C2(n16613), .A(n16753), .B(n16612), .ZN(
        n16614) );
  OAI211_X1 U19792 ( .C1(n16739), .C2(n16616), .A(n16615), .B(n16614), .ZN(
        P3_U2660) );
  INV_X1 U19793 ( .A(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n16628) );
  AOI211_X1 U19794 ( .C1(P3_EBX_REG_10__SCAN_IN), .C2(n16637), .A(n16617), .B(
        n16723), .ZN(n16626) );
  AOI21_X1 U19795 ( .B1(n16735), .B2(n16618), .A(n16722), .ZN(n16648) );
  INV_X1 U19796 ( .A(P3_REIP_REG_10__SCAN_IN), .ZN(n18588) );
  OAI211_X1 U19797 ( .C1(P3_REIP_REG_10__SCAN_IN), .C2(P3_REIP_REG_9__SCAN_IN), 
        .A(n16635), .B(n16619), .ZN(n16624) );
  INV_X1 U19798 ( .A(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n17647) );
  NAND2_X1 U19799 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17636), .ZN(
        n16677) );
  NOR2_X1 U19800 ( .A1(n17647), .A2(n16677), .ZN(n16664) );
  NAND2_X1 U19801 ( .A1(n17583), .A2(n16664), .ZN(n16629) );
  AOI21_X1 U19802 ( .B1(n16628), .B2(n16629), .A(n16620), .ZN(n17590) );
  OAI21_X1 U19803 ( .B1(n16629), .B2(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A(
        n10006), .ZN(n16621) );
  INV_X1 U19804 ( .A(n16621), .ZN(n16632) );
  AOI21_X1 U19805 ( .B1(n17590), .B2(n16632), .A(n18549), .ZN(n16622) );
  OAI21_X1 U19806 ( .B1(n17590), .B2(n16632), .A(n16622), .ZN(n16623) );
  OAI211_X1 U19807 ( .C1(n16648), .C2(n18588), .A(n16624), .B(n16623), .ZN(
        n16625) );
  AOI211_X1 U19808 ( .C1(P3_EBX_REG_10__SCAN_IN), .C2(n16754), .A(n16626), .B(
        n16625), .ZN(n16627) );
  OAI211_X1 U19809 ( .C1(n16628), .C2(n16739), .A(n16627), .B(n18028), .ZN(
        P3_U2661) );
  INV_X1 U19810 ( .A(n16648), .ZN(n16636) );
  INV_X1 U19811 ( .A(P3_REIP_REG_9__SCAN_IN), .ZN(n18586) );
  INV_X1 U19812 ( .A(n16664), .ZN(n16654) );
  NOR2_X1 U19813 ( .A1(n17619), .A2(n16654), .ZN(n16643) );
  OAI21_X1 U19814 ( .B1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n16643), .A(
        n16629), .ZN(n17600) );
  INV_X1 U19815 ( .A(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n16644) );
  INV_X1 U19816 ( .A(n17600), .ZN(n16630) );
  INV_X1 U19817 ( .A(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n17624) );
  NOR2_X1 U19818 ( .A1(n17609), .A2(n17624), .ZN(n17620) );
  NAND2_X1 U19819 ( .A1(n16727), .A2(n17620), .ZN(n16645) );
  AOI221_X1 U19820 ( .B1(n16644), .B2(n16630), .C1(n16645), .C2(n16630), .A(
        n18549), .ZN(n16631) );
  AOI22_X1 U19821 ( .A1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n16691), .B1(
        n16632), .B2(n16631), .ZN(n16633) );
  OAI211_X1 U19822 ( .C1(n17600), .C2(n16728), .A(n16633), .B(n18028), .ZN(
        n16634) );
  AOI221_X1 U19823 ( .B1(n16636), .B2(P3_REIP_REG_9__SCAN_IN), .C1(n16635), 
        .C2(n18586), .A(n16634), .ZN(n16639) );
  OAI211_X1 U19824 ( .C1(n16641), .C2(n16640), .A(n16753), .B(n16637), .ZN(
        n16638) );
  OAI211_X1 U19825 ( .C1(n16640), .C2(n16743), .A(n16639), .B(n16638), .ZN(
        P3_U2662) );
  AOI211_X1 U19826 ( .C1(P3_EBX_REG_8__SCAN_IN), .C2(n16659), .A(n16641), .B(
        n16723), .ZN(n16651) );
  AOI21_X1 U19827 ( .B1(n16735), .B2(n16642), .A(P3_REIP_REG_8__SCAN_IN), .ZN(
        n16649) );
  NAND2_X1 U19828 ( .A1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(n16664), .ZN(
        n16655) );
  AOI21_X1 U19829 ( .B1(n16644), .B2(n16655), .A(n16643), .ZN(n17611) );
  NAND2_X1 U19830 ( .A1(n10006), .A2(n16645), .ZN(n16646) );
  XOR2_X1 U19831 ( .A(n17611), .B(n16646), .Z(n16647) );
  OAI22_X1 U19832 ( .A1(n16649), .A2(n16648), .B1(n18549), .B2(n16647), .ZN(
        n16650) );
  AOI211_X1 U19833 ( .C1(n16691), .C2(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A(
        n16651), .B(n16650), .ZN(n16652) );
  OAI211_X1 U19834 ( .C1(n16743), .C2(n17033), .A(n16652), .B(n18028), .ZN(
        P3_U2663) );
  AOI22_X1 U19835 ( .A1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(n16691), .B1(
        n16754), .B2(P3_EBX_REG_7__SCAN_IN), .ZN(n16663) );
  NOR2_X1 U19836 ( .A1(n16722), .A2(n16653), .ZN(n16682) );
  AOI21_X1 U19837 ( .B1(P3_REIP_REG_6__SCAN_IN), .B2(n16682), .A(n16681), .ZN(
        n16666) );
  NAND3_X1 U19838 ( .A1(n16735), .A2(P3_REIP_REG_5__SCAN_IN), .A3(n16680), 
        .ZN(n16668) );
  NOR2_X1 U19839 ( .A1(n18580), .A2(n16668), .ZN(n16658) );
  OAI21_X1 U19840 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n16654), .A(
        n10006), .ZN(n16672) );
  OAI21_X1 U19841 ( .B1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n16664), .A(
        n16655), .ZN(n17635) );
  OAI21_X1 U19842 ( .B1(n16672), .B2(n17635), .A(n16697), .ZN(n16656) );
  AOI21_X1 U19843 ( .B1(n16672), .B2(n17635), .A(n16656), .ZN(n16657) );
  AOI221_X1 U19844 ( .B1(n16666), .B2(P3_REIP_REG_7__SCAN_IN), .C1(n16658), 
        .C2(n18582), .A(n16657), .ZN(n16662) );
  OAI211_X1 U19845 ( .C1(n16669), .C2(n16660), .A(n16753), .B(n16659), .ZN(
        n16661) );
  NAND4_X1 U19846 ( .A1(n16663), .A2(n16662), .A3(n18028), .A4(n16661), .ZN(
        P3_U2664) );
  AOI21_X1 U19847 ( .B1(n17647), .B2(n16677), .A(n16664), .ZN(n17644) );
  AOI21_X1 U19848 ( .B1(n10006), .B2(n16677), .A(n16750), .ZN(n16665) );
  AOI22_X1 U19849 ( .A1(n16754), .A2(P3_EBX_REG_6__SCAN_IN), .B1(n17644), .B2(
        n16665), .ZN(n16675) );
  INV_X1 U19850 ( .A(n16666), .ZN(n16667) );
  AOI21_X1 U19851 ( .B1(n18580), .B2(n16668), .A(n16667), .ZN(n16671) );
  AOI211_X1 U19852 ( .C1(P3_EBX_REG_6__SCAN_IN), .C2(n16684), .A(n16669), .B(
        n16723), .ZN(n16670) );
  AOI211_X1 U19853 ( .C1(n16691), .C2(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A(
        n16671), .B(n16670), .ZN(n16674) );
  OR3_X1 U19854 ( .A1(n17644), .A2(n16672), .A3(n18549), .ZN(n16673) );
  NAND4_X1 U19855 ( .A1(n16675), .A2(n16674), .A3(n18028), .A4(n16673), .ZN(
        P3_U2665) );
  INV_X1 U19856 ( .A(n16676), .ZN(n17648) );
  NAND2_X1 U19857 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17648), .ZN(
        n16694) );
  INV_X1 U19858 ( .A(n16677), .ZN(n16678) );
  AOI21_X1 U19859 ( .B1(n16690), .B2(n16694), .A(n16678), .ZN(n17654) );
  AOI21_X1 U19860 ( .B1(n17648), .B2(n16727), .A(n16679), .ZN(n16698) );
  XOR2_X1 U19861 ( .A(n17654), .B(n16698), .Z(n16688) );
  INV_X1 U19862 ( .A(P3_REIP_REG_5__SCAN_IN), .ZN(n18578) );
  NAND2_X1 U19863 ( .A1(n16735), .A2(n16680), .ZN(n16683) );
  AOI211_X1 U19864 ( .C1(n18578), .C2(n16683), .A(n16682), .B(n16681), .ZN(
        n16687) );
  OAI211_X1 U19865 ( .C1(n16692), .C2(n17040), .A(n16753), .B(n16684), .ZN(
        n16685) );
  OAI21_X1 U19866 ( .B1(n17040), .B2(n16743), .A(n16685), .ZN(n16686) );
  AOI211_X1 U19867 ( .C1(n16697), .C2(n16688), .A(n16687), .B(n16686), .ZN(
        n16689) );
  INV_X1 U19868 ( .A(n17971), .ZN(n18013) );
  OAI211_X1 U19869 ( .C1(n16690), .C2(n16739), .A(n16689), .B(n18013), .ZN(
        P3_U2666) );
  AOI21_X1 U19870 ( .B1(n16735), .B2(n16712), .A(n16722), .ZN(n16707) );
  AOI22_X1 U19871 ( .A1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n16691), .B1(
        n16754), .B2(P3_EBX_REG_4__SCAN_IN), .ZN(n16706) );
  AOI211_X1 U19872 ( .C1(P3_EBX_REG_4__SCAN_IN), .C2(n16718), .A(n16692), .B(
        n16723), .ZN(n16704) );
  NOR3_X1 U19873 ( .A1(P3_REIP_REG_4__SCAN_IN), .A2(n16744), .A3(n16712), .ZN(
        n16703) );
  NAND2_X1 U19874 ( .A1(n18047), .A2(n18707), .ZN(n16742) );
  INV_X1 U19875 ( .A(n17669), .ZN(n16695) );
  NOR2_X1 U19876 ( .A1(n16693), .A2(n16695), .ZN(n16709) );
  OAI21_X1 U19877 ( .B1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n16709), .A(
        n16694), .ZN(n17672) );
  OR2_X1 U19878 ( .A1(n16695), .A2(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n17663) );
  OAI22_X1 U19879 ( .A1(n10006), .A2(n17672), .B1(n17663), .B2(n16696), .ZN(
        n16699) );
  OAI221_X1 U19880 ( .B1(n16699), .B2(n16698), .C1(n16699), .C2(n17672), .A(
        n16697), .ZN(n16700) );
  OAI221_X1 U19881 ( .B1(n16742), .B2(n15148), .C1(n16742), .C2(n16701), .A(
        n16700), .ZN(n16702) );
  NOR4_X1 U19882 ( .A1(n17971), .A2(n16704), .A3(n16703), .A4(n16702), .ZN(
        n16705) );
  OAI211_X1 U19883 ( .C1(n16707), .C2(n18576), .A(n16706), .B(n16705), .ZN(
        P3_U2667) );
  INV_X1 U19884 ( .A(n16707), .ZN(n16717) );
  NAND2_X1 U19885 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n18505) );
  INV_X1 U19886 ( .A(n18505), .ZN(n16708) );
  NAND2_X1 U19887 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n16708), .ZN(
        n18496) );
  INV_X1 U19888 ( .A(n18496), .ZN(n16721) );
  OAI21_X1 U19889 ( .B1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n16721), .A(
        n15148), .ZN(n18641) );
  OAI22_X1 U19890 ( .A1(n16743), .A2(n17050), .B1(n16742), .B2(n18641), .ZN(
        n16716) );
  NAND2_X1 U19891 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n16726) );
  AOI21_X1 U19892 ( .B1(n17679), .B2(n16726), .A(n16709), .ZN(n16710) );
  INV_X1 U19893 ( .A(n16710), .ZN(n17685) );
  OAI21_X1 U19894 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n16726), .A(
        n10006), .ZN(n16711) );
  XNOR2_X1 U19895 ( .A(n17685), .B(n16711), .ZN(n16714) );
  NAND2_X1 U19896 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(P3_REIP_REG_2__SCAN_IN), 
        .ZN(n16734) );
  NAND2_X1 U19897 ( .A1(n16735), .A2(n16712), .ZN(n16713) );
  OAI22_X1 U19898 ( .A1(n18549), .A2(n16714), .B1(n16734), .B2(n16713), .ZN(
        n16715) );
  AOI211_X1 U19899 ( .C1(P3_REIP_REG_3__SCAN_IN), .C2(n16717), .A(n16716), .B(
        n16715), .ZN(n16720) );
  OAI211_X1 U19900 ( .C1(n16724), .C2(n17050), .A(n16753), .B(n16718), .ZN(
        n16719) );
  OAI211_X1 U19901 ( .C1(n16739), .C2(n17679), .A(n16720), .B(n16719), .ZN(
        P3_U2668) );
  AOI21_X1 U19902 ( .B1(n13943), .B2(n18504), .A(n16721), .ZN(n18653) );
  INV_X1 U19903 ( .A(n16742), .ZN(n18709) );
  AOI22_X1 U19904 ( .A1(P3_REIP_REG_2__SCAN_IN), .A2(n16722), .B1(n18653), 
        .B2(n18709), .ZN(n16738) );
  INV_X1 U19905 ( .A(P3_EBX_REG_0__SCAN_IN), .ZN(n17072) );
  INV_X1 U19906 ( .A(P3_EBX_REG_1__SCAN_IN), .ZN(n17066) );
  NAND2_X1 U19907 ( .A1(n17072), .A2(n17066), .ZN(n17063) );
  AOI211_X1 U19908 ( .C1(P3_EBX_REG_2__SCAN_IN), .C2(n17063), .A(n16724), .B(
        n16723), .ZN(n16733) );
  OAI22_X1 U19909 ( .A1(n17694), .A2(n16739), .B1(n16743), .B2(n16725), .ZN(
        n16732) );
  OAI21_X1 U19910 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A(n16726), .ZN(n17691) );
  OAI22_X1 U19911 ( .A1(n16727), .A2(n17691), .B1(
        P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n16726), .ZN(n16729) );
  OAI22_X1 U19912 ( .A1(n16730), .A2(n16729), .B1(n17691), .B2(n16728), .ZN(
        n16731) );
  NOR3_X1 U19913 ( .A1(n16733), .A2(n16732), .A3(n16731), .ZN(n16737) );
  OAI211_X1 U19914 ( .C1(P3_REIP_REG_1__SCAN_IN), .C2(P3_REIP_REG_2__SCAN_IN), 
        .A(n16735), .B(n16734), .ZN(n16736) );
  NAND3_X1 U19915 ( .A1(n16738), .A2(n16737), .A3(n16736), .ZN(P3_U2669) );
  NAND2_X1 U19916 ( .A1(n10006), .A2(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n16740) );
  OAI21_X1 U19917 ( .B1(n18549), .B2(n16740), .A(n16739), .ZN(n16747) );
  NAND2_X1 U19918 ( .A1(n16741), .A2(n18504), .ZN(n18656) );
  OAI22_X1 U19919 ( .A1(n18679), .A2(n16752), .B1(n18656), .B2(n16742), .ZN(
        n16746) );
  OAI22_X1 U19920 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(n16744), .B1(n16743), 
        .B2(n17066), .ZN(n16745) );
  AOI211_X1 U19921 ( .C1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .C2(n16747), .A(
        n16746), .B(n16745), .ZN(n16749) );
  NAND3_X1 U19922 ( .A1(n16753), .A2(n17063), .A3(n17062), .ZN(n16748) );
  OAI211_X1 U19923 ( .C1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .C2(n16750), .A(
        n16749), .B(n16748), .ZN(P3_U2670) );
  AOI22_X1 U19924 ( .A1(P3_REIP_REG_0__SCAN_IN), .A2(n16751), .B1(n18709), 
        .B2(n18668), .ZN(n16757) );
  INV_X1 U19925 ( .A(n18705), .ZN(n18642) );
  NAND3_X1 U19926 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n18642), .A3(
        n16752), .ZN(n16756) );
  OAI21_X1 U19927 ( .B1(n16754), .B2(n16753), .A(P3_EBX_REG_0__SCAN_IN), .ZN(
        n16755) );
  NAND3_X1 U19928 ( .A1(n16757), .A2(n16756), .A3(n16755), .ZN(P3_U2671) );
  INV_X1 U19929 ( .A(P3_EBX_REG_26__SCAN_IN), .ZN(n16801) );
  NAND3_X1 U19930 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(P3_EBX_REG_21__SCAN_IN), 
        .A3(n16794), .ZN(n16758) );
  NOR4_X1 U19931 ( .A1(n16801), .A2(n16759), .A3(n16848), .A4(n16758), .ZN(
        n16760) );
  NAND4_X1 U19932 ( .A1(P3_EBX_REG_29__SCAN_IN), .A2(P3_EBX_REG_25__SCAN_IN), 
        .A3(P3_EBX_REG_24__SCAN_IN), .A4(n16760), .ZN(n16763) );
  NOR2_X1 U19933 ( .A1(n16764), .A2(n16763), .ZN(n16789) );
  NAND2_X1 U19934 ( .A1(n17064), .A2(P3_EBX_REG_31__SCAN_IN), .ZN(n16762) );
  NAND2_X1 U19935 ( .A1(n16789), .A2(n18087), .ZN(n16761) );
  OAI22_X1 U19936 ( .A1(n16789), .A2(n16762), .B1(P3_EBX_REG_31__SCAN_IN), 
        .B2(n16761), .ZN(P3_U2672) );
  NAND2_X1 U19937 ( .A1(n16764), .A2(n16763), .ZN(n16765) );
  NAND2_X1 U19938 ( .A1(n16765), .A2(n17064), .ZN(n16788) );
  AOI22_X1 U19939 ( .A1(n16992), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n16995), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n16769) );
  AOI22_X1 U19940 ( .A1(n17005), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n16977), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n16768) );
  AOI22_X1 U19941 ( .A1(n9633), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n17022), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n16767) );
  AOI22_X1 U19942 ( .A1(n16997), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n17014), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n16766) );
  NAND4_X1 U19943 ( .A1(n16769), .A2(n16768), .A3(n16767), .A4(n16766), .ZN(
        n16775) );
  AOI22_X1 U19944 ( .A1(n16989), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n16825), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n16773) );
  AOI22_X1 U19945 ( .A1(n9627), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n16991), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n16772) );
  AOI22_X1 U19946 ( .A1(n16923), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n17023), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n16771) );
  AOI22_X1 U19947 ( .A1(n16958), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n16996), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n16770) );
  NAND4_X1 U19948 ( .A1(n16773), .A2(n16772), .A3(n16771), .A4(n16770), .ZN(
        n16774) );
  NOR2_X1 U19949 ( .A1(n16775), .A2(n16774), .ZN(n16787) );
  AOI22_X1 U19950 ( .A1(n16989), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n9633), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n16786) );
  AOI22_X1 U19951 ( .A1(n16992), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n16991), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n16785) );
  AOI22_X1 U19952 ( .A1(n9627), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n17013), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n16776) );
  OAI21_X1 U19953 ( .B1(n16777), .B2(n16823), .A(n16776), .ZN(n16783) );
  AOI22_X1 U19954 ( .A1(n16923), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n17022), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n16781) );
  AOI22_X1 U19955 ( .A1(n17005), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n16995), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n16780) );
  AOI22_X1 U19956 ( .A1(n16997), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n16825), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n16779) );
  AOI22_X1 U19957 ( .A1(n17014), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n16996), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n16778) );
  NAND4_X1 U19958 ( .A1(n16781), .A2(n16780), .A3(n16779), .A4(n16778), .ZN(
        n16782) );
  AOI211_X1 U19959 ( .C1(n16977), .C2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .A(
        n16783), .B(n16782), .ZN(n16784) );
  NAND3_X1 U19960 ( .A1(n16786), .A2(n16785), .A3(n16784), .ZN(n16791) );
  NAND2_X1 U19961 ( .A1(n16792), .A2(n16791), .ZN(n16790) );
  XNOR2_X1 U19962 ( .A(n16787), .B(n16790), .ZN(n17083) );
  OAI22_X1 U19963 ( .A1(n16789), .A2(n16788), .B1(n17083), .B2(n17064), .ZN(
        P3_U2673) );
  OAI21_X1 U19964 ( .B1(n16792), .B2(n16791), .A(n16790), .ZN(n17090) );
  NOR2_X1 U19965 ( .A1(P3_EBX_REG_29__SCAN_IN), .A2(n16805), .ZN(n16793) );
  AOI22_X1 U19966 ( .A1(P3_EBX_REG_29__SCAN_IN), .A2(n16795), .B1(n16794), 
        .B2(n16793), .ZN(n16796) );
  OAI21_X1 U19967 ( .B1(n17090), .B2(n17064), .A(n16796), .ZN(P3_U2674) );
  OAI21_X1 U19968 ( .B1(n16802), .B2(n16798), .A(n16797), .ZN(n17100) );
  NAND3_X1 U19969 ( .A1(n16805), .A2(P3_EBX_REG_27__SCAN_IN), .A3(n17064), 
        .ZN(n16799) );
  OAI221_X1 U19970 ( .B1(n16805), .B2(P3_EBX_REG_27__SCAN_IN), .C1(n17064), 
        .C2(n17100), .A(n16799), .ZN(P3_U2676) );
  OAI21_X1 U19971 ( .B1(n16801), .B2(n17070), .A(n16800), .ZN(n16804) );
  AOI21_X1 U19972 ( .B1(n16803), .B2(n16807), .A(n16802), .ZN(n17101) );
  AOI22_X1 U19973 ( .A1(n16805), .A2(n16804), .B1(n17070), .B2(n17101), .ZN(
        n16806) );
  INV_X1 U19974 ( .A(n16806), .ZN(P3_U2677) );
  AND2_X1 U19975 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(n16821), .ZN(n16815) );
  AOI21_X1 U19976 ( .B1(P3_EBX_REG_25__SCAN_IN), .B2(n17064), .A(n16815), .ZN(
        n16809) );
  OAI21_X1 U19977 ( .B1(n16811), .B2(n16808), .A(n16807), .ZN(n17110) );
  OAI22_X1 U19978 ( .A1(n16810), .A2(n16809), .B1(n17064), .B2(n17110), .ZN(
        P3_U2678) );
  AOI21_X1 U19979 ( .B1(P3_EBX_REG_24__SCAN_IN), .B2(n17064), .A(n16821), .ZN(
        n16814) );
  AOI21_X1 U19980 ( .B1(n16812), .B2(n16817), .A(n16811), .ZN(n17111) );
  INV_X1 U19981 ( .A(n17111), .ZN(n16813) );
  OAI22_X1 U19982 ( .A1(n16815), .A2(n16814), .B1(n17064), .B2(n16813), .ZN(
        P3_U2679) );
  AOI21_X1 U19983 ( .B1(P3_EBX_REG_23__SCAN_IN), .B2(n17064), .A(n16816), .ZN(
        n16820) );
  OAI21_X1 U19984 ( .B1(n16819), .B2(n16818), .A(n16817), .ZN(n17121) );
  OAI22_X1 U19985 ( .A1(n16821), .A2(n16820), .B1(n17064), .B2(n17121), .ZN(
        P3_U2680) );
  AOI22_X1 U19986 ( .A1(n16958), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n17022), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n16834) );
  AOI22_X1 U19987 ( .A1(n17005), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n17023), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n16833) );
  AOI22_X1 U19988 ( .A1(n17021), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n16996), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n16822) );
  OAI21_X1 U19989 ( .B1(n16824), .B2(n16823), .A(n16822), .ZN(n16831) );
  AOI22_X1 U19990 ( .A1(n16997), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n16974), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n16829) );
  AOI22_X1 U19991 ( .A1(n16992), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n16989), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n16828) );
  AOI22_X1 U19992 ( .A1(n16923), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n16825), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n16827) );
  AOI22_X1 U19993 ( .A1(n16990), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n17014), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n16826) );
  NAND4_X1 U19994 ( .A1(n16829), .A2(n16828), .A3(n16827), .A4(n16826), .ZN(
        n16830) );
  AOI211_X1 U19995 ( .C1(n9633), .C2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .A(
        n16831), .B(n16830), .ZN(n16832) );
  NAND3_X1 U19996 ( .A1(n16834), .A2(n16833), .A3(n16832), .ZN(n17122) );
  INV_X1 U19997 ( .A(n17122), .ZN(n16836) );
  NAND3_X1 U19998 ( .A1(n16837), .A2(P3_EBX_REG_22__SCAN_IN), .A3(n17064), 
        .ZN(n16835) );
  OAI221_X1 U19999 ( .B1(n16837), .B2(P3_EBX_REG_22__SCAN_IN), .C1(n17064), 
        .C2(n16836), .A(n16835), .ZN(P3_U2681) );
  AOI22_X1 U20000 ( .A1(n16992), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n16991), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n16841) );
  AOI22_X1 U20001 ( .A1(n9627), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n16923), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n16840) );
  AOI22_X1 U20002 ( .A1(n16990), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n17014), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n16839) );
  AOI22_X1 U20003 ( .A1(n17005), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n16996), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n16838) );
  NAND4_X1 U20004 ( .A1(n16841), .A2(n16840), .A3(n16839), .A4(n16838), .ZN(
        n16847) );
  AOI22_X1 U20005 ( .A1(n16924), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n17022), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n16845) );
  AOI22_X1 U20006 ( .A1(n17020), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n17023), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n16844) );
  AOI22_X1 U20007 ( .A1(n16989), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n17013), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n16843) );
  AOI22_X1 U20008 ( .A1(n16997), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n9633), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n16842) );
  NAND4_X1 U20009 ( .A1(n16845), .A2(n16844), .A3(n16843), .A4(n16842), .ZN(
        n16846) );
  NOR2_X1 U20010 ( .A1(n16847), .A2(n16846), .ZN(n17129) );
  AND2_X1 U20011 ( .A1(n17064), .A2(n16848), .ZN(n16862) );
  AOI22_X1 U20012 ( .A1(P3_EBX_REG_21__SCAN_IN), .A2(n16862), .B1(n16850), 
        .B2(n16849), .ZN(n16851) );
  OAI21_X1 U20013 ( .B1(n17129), .B2(n17064), .A(n16851), .ZN(P3_U2682) );
  AOI22_X1 U20014 ( .A1(n17005), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n17022), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n16855) );
  AOI22_X1 U20015 ( .A1(n16997), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n17023), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n16854) );
  AOI22_X1 U20016 ( .A1(n17013), .A2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n16996), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n16853) );
  AOI22_X1 U20017 ( .A1(n9633), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n17014), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n16852) );
  NAND4_X1 U20018 ( .A1(n16855), .A2(n16854), .A3(n16853), .A4(n16852), .ZN(
        n16861) );
  AOI22_X1 U20019 ( .A1(n16995), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n16923), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n16859) );
  AOI22_X1 U20020 ( .A1(n16989), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n17020), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n16858) );
  AOI22_X1 U20021 ( .A1(n16992), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n16977), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n16857) );
  AOI22_X1 U20022 ( .A1(n16974), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n16991), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n16856) );
  NAND4_X1 U20023 ( .A1(n16859), .A2(n16858), .A3(n16857), .A4(n16856), .ZN(
        n16860) );
  NOR2_X1 U20024 ( .A1(n16861), .A2(n16860), .ZN(n17136) );
  AND2_X1 U20025 ( .A1(n18087), .A2(n16874), .ZN(n16876) );
  OAI221_X1 U20026 ( .B1(P3_EBX_REG_20__SCAN_IN), .B2(P3_EBX_REG_19__SCAN_IN), 
        .C1(P3_EBX_REG_20__SCAN_IN), .C2(n16876), .A(n16862), .ZN(n16863) );
  OAI21_X1 U20027 ( .B1(n17136), .B2(n17064), .A(n16863), .ZN(P3_U2683) );
  AOI22_X1 U20028 ( .A1(n17005), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n16974), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n16867) );
  AOI22_X1 U20029 ( .A1(n16924), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n9633), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n16866) );
  AOI22_X1 U20030 ( .A1(n16989), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n17022), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n16865) );
  AOI22_X1 U20031 ( .A1(n16923), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n17014), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n16864) );
  NAND4_X1 U20032 ( .A1(n16867), .A2(n16866), .A3(n16865), .A4(n16864), .ZN(
        n16873) );
  AOI22_X1 U20033 ( .A1(n16996), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n17023), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n16871) );
  AOI22_X1 U20034 ( .A1(n16992), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n16977), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n16870) );
  AOI22_X1 U20035 ( .A1(n16997), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n17020), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n16869) );
  AOI22_X1 U20036 ( .A1(n16958), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n16991), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n16868) );
  NAND4_X1 U20037 ( .A1(n16871), .A2(n16870), .A3(n16869), .A4(n16868), .ZN(
        n16872) );
  NOR2_X1 U20038 ( .A1(n16873), .A2(n16872), .ZN(n17141) );
  NOR2_X1 U20039 ( .A1(n17070), .A2(n16874), .ZN(n16890) );
  AOI22_X1 U20040 ( .A1(P3_EBX_REG_19__SCAN_IN), .A2(n16890), .B1(n16876), 
        .B2(n16875), .ZN(n16877) );
  OAI21_X1 U20041 ( .B1(n17141), .B2(n17064), .A(n16877), .ZN(P3_U2684) );
  AOI22_X1 U20042 ( .A1(n9633), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n17023), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n16881) );
  AOI22_X1 U20043 ( .A1(n17020), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n17022), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n16880) );
  AOI22_X1 U20044 ( .A1(n16990), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n16923), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n16879) );
  AOI22_X1 U20045 ( .A1(n17005), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n17014), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n16878) );
  NAND4_X1 U20046 ( .A1(n16881), .A2(n16880), .A3(n16879), .A4(n16878), .ZN(
        n16887) );
  AOI22_X1 U20047 ( .A1(n16924), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n16996), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n16885) );
  AOI22_X1 U20048 ( .A1(n16974), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n17013), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n16884) );
  AOI22_X1 U20049 ( .A1(n16997), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n16991), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n16883) );
  AOI22_X1 U20050 ( .A1(n16992), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n16989), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n16882) );
  NAND4_X1 U20051 ( .A1(n16885), .A2(n16884), .A3(n16883), .A4(n16882), .ZN(
        n16886) );
  NOR2_X1 U20052 ( .A1(n16887), .A2(n16886), .ZN(n17145) );
  NAND3_X1 U20053 ( .A1(n18087), .A2(P3_EBX_REG_16__SCAN_IN), .A3(n16932), 
        .ZN(n16905) );
  NOR2_X1 U20054 ( .A1(n16904), .A2(n16905), .ZN(n16889) );
  AOI22_X1 U20055 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n16890), .B1(n16889), 
        .B2(n16888), .ZN(n16891) );
  OAI21_X1 U20056 ( .B1(n17145), .B2(n17064), .A(n16891), .ZN(P3_U2685) );
  NAND2_X1 U20057 ( .A1(n17064), .A2(n16892), .ZN(n16916) );
  AOI22_X1 U20058 ( .A1(n16997), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n16989), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n16896) );
  AOI22_X1 U20059 ( .A1(n16992), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_15__1__SCAN_IN), .B2(n16924), .ZN(n16895) );
  AOI22_X1 U20060 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n9633), .B1(
        P3_INSTQUEUE_REG_7__1__SCAN_IN), .B2(n17022), .ZN(n16894) );
  AOI22_X1 U20061 ( .A1(n17005), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_1__1__SCAN_IN), .B2(n17014), .ZN(n16893) );
  NAND4_X1 U20062 ( .A1(n16896), .A2(n16895), .A3(n16894), .A4(n16893), .ZN(
        n16902) );
  AOI22_X1 U20063 ( .A1(P3_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n16958), .B1(
        n16996), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n16900) );
  AOI22_X1 U20064 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n17020), .B1(
        P3_INSTQUEUE_REG_12__1__SCAN_IN), .B2(n9627), .ZN(n16899) );
  AOI22_X1 U20065 ( .A1(n16990), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_6__1__SCAN_IN), .B2(n16923), .ZN(n16898) );
  AOI22_X1 U20066 ( .A1(n17021), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_14__1__SCAN_IN), .B2(n17023), .ZN(n16897) );
  NAND4_X1 U20067 ( .A1(n16900), .A2(n16899), .A3(n16898), .A4(n16897), .ZN(
        n16901) );
  NOR2_X1 U20068 ( .A1(n16902), .A2(n16901), .ZN(n17151) );
  OR2_X1 U20069 ( .A1(n17151), .A2(n17064), .ZN(n16903) );
  OAI221_X1 U20070 ( .B1(P3_EBX_REG_17__SCAN_IN), .B2(n16905), .C1(n16904), 
        .C2(n16916), .A(n16903), .ZN(P3_U2686) );
  AOI22_X1 U20071 ( .A1(n16974), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n17020), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n16909) );
  AOI22_X1 U20072 ( .A1(n9633), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n16991), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n16908) );
  AOI22_X1 U20073 ( .A1(n16958), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n17022), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n16907) );
  AOI22_X1 U20074 ( .A1(n17014), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n17023), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n16906) );
  NAND4_X1 U20075 ( .A1(n16909), .A2(n16908), .A3(n16907), .A4(n16906), .ZN(
        n16915) );
  AOI22_X1 U20076 ( .A1(n16989), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n16995), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n16913) );
  AOI22_X1 U20077 ( .A1(n16992), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n16977), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n16912) );
  AOI22_X1 U20078 ( .A1(n16997), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n16923), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n16911) );
  AOI22_X1 U20079 ( .A1(n17005), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n16996), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n16910) );
  NAND4_X1 U20080 ( .A1(n16913), .A2(n16912), .A3(n16911), .A4(n16910), .ZN(
        n16914) );
  NOR2_X1 U20081 ( .A1(n16915), .A2(n16914), .ZN(n17157) );
  NOR2_X1 U20082 ( .A1(n16932), .A2(P3_EBX_REG_16__SCAN_IN), .ZN(n16917) );
  OAI22_X1 U20083 ( .A1(n17157), .A2(n17064), .B1(n16917), .B2(n16916), .ZN(
        P3_U2687) );
  INV_X1 U20084 ( .A(n16943), .ZN(n16918) );
  OAI21_X1 U20085 ( .B1(P3_EBX_REG_15__SCAN_IN), .B2(n16918), .A(n17064), .ZN(
        n16931) );
  AOI22_X1 U20086 ( .A1(n17020), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n17023), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n16922) );
  AOI22_X1 U20087 ( .A1(n17005), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n17013), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n16921) );
  AOI22_X1 U20088 ( .A1(n16990), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n9633), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n16920) );
  AOI22_X1 U20089 ( .A1(n16974), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n17014), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n16919) );
  NAND4_X1 U20090 ( .A1(n16922), .A2(n16921), .A3(n16920), .A4(n16919), .ZN(
        n16930) );
  AOI22_X1 U20091 ( .A1(n16992), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n16991), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n16928) );
  AOI22_X1 U20092 ( .A1(n16997), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n16989), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n16927) );
  AOI22_X1 U20093 ( .A1(n16923), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n17022), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n16926) );
  AOI22_X1 U20094 ( .A1(n16924), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n16996), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n16925) );
  NAND4_X1 U20095 ( .A1(n16928), .A2(n16927), .A3(n16926), .A4(n16925), .ZN(
        n16929) );
  NOR2_X1 U20096 ( .A1(n16930), .A2(n16929), .ZN(n17161) );
  OAI22_X1 U20097 ( .A1(n16932), .A2(n16931), .B1(n17161), .B2(n17064), .ZN(
        P3_U2688) );
  AOI22_X1 U20098 ( .A1(n16992), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n16995), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n16936) );
  AOI22_X1 U20099 ( .A1(n16989), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n17021), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n16935) );
  AOI22_X1 U20100 ( .A1(n16998), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n17014), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n16934) );
  AOI22_X1 U20101 ( .A1(n17023), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n17022), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n16933) );
  NAND4_X1 U20102 ( .A1(n16936), .A2(n16935), .A3(n16934), .A4(n16933), .ZN(
        n16942) );
  AOI22_X1 U20103 ( .A1(n17005), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n9633), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n16940) );
  AOI22_X1 U20104 ( .A1(n16974), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n17020), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n16939) );
  AOI22_X1 U20105 ( .A1(n16990), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n16997), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n16938) );
  AOI22_X1 U20106 ( .A1(n9626), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n16996), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n16937) );
  NAND4_X1 U20107 ( .A1(n16940), .A2(n16939), .A3(n16938), .A4(n16937), .ZN(
        n16941) );
  NOR2_X1 U20108 ( .A1(n16942), .A2(n16941), .ZN(n17166) );
  OAI21_X1 U20109 ( .B1(P3_EBX_REG_14__SCAN_IN), .B2(n16944), .A(n16943), .ZN(
        n16945) );
  AOI22_X1 U20110 ( .A1(n17070), .A2(n17166), .B1(n16945), .B2(n17064), .ZN(
        P3_U2689) );
  NOR3_X1 U20111 ( .A1(n17123), .A2(n17032), .A3(n16946), .ZN(n16988) );
  NAND2_X1 U20112 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n16988), .ZN(n16972) );
  AOI22_X1 U20113 ( .A1(n17005), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n16992), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n16950) );
  AOI22_X1 U20114 ( .A1(n16995), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n16991), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n16949) );
  AOI22_X1 U20115 ( .A1(n16998), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n16923), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n16948) );
  AOI22_X1 U20116 ( .A1(n17014), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n17022), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n16947) );
  NAND4_X1 U20117 ( .A1(n16950), .A2(n16949), .A3(n16948), .A4(n16947), .ZN(
        n16956) );
  AOI22_X1 U20118 ( .A1(n16989), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n16974), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n16954) );
  AOI22_X1 U20119 ( .A1(n16990), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n16996), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n16953) );
  AOI22_X1 U20120 ( .A1(n16997), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n17023), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n16952) );
  AOI22_X1 U20121 ( .A1(n9633), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n17020), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n16951) );
  NAND4_X1 U20122 ( .A1(n16954), .A2(n16953), .A3(n16952), .A4(n16951), .ZN(
        n16955) );
  NOR2_X1 U20123 ( .A1(n16956), .A2(n16955), .ZN(n17167) );
  NAND3_X1 U20124 ( .A1(n16972), .A2(P3_EBX_REG_13__SCAN_IN), .A3(n17064), 
        .ZN(n16957) );
  OAI221_X1 U20125 ( .B1(n16972), .B2(P3_EBX_REG_13__SCAN_IN), .C1(n17064), 
        .C2(n17167), .A(n16957), .ZN(P3_U2690) );
  AOI22_X1 U20126 ( .A1(n16974), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n9626), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n16962) );
  AOI22_X1 U20127 ( .A1(n16995), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n17020), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n16961) );
  AOI22_X1 U20128 ( .A1(n16989), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n16958), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n16960) );
  AOI22_X1 U20129 ( .A1(n17021), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n17014), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n16959) );
  NAND4_X1 U20130 ( .A1(n16962), .A2(n16961), .A3(n16960), .A4(n16959), .ZN(
        n16968) );
  AOI22_X1 U20131 ( .A1(n17023), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n17022), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n16966) );
  AOI22_X1 U20132 ( .A1(n16992), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n16997), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n16965) );
  AOI22_X1 U20133 ( .A1(n17005), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n16996), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n16964) );
  AOI22_X1 U20134 ( .A1(n16990), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n9633), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n16963) );
  NAND4_X1 U20135 ( .A1(n16966), .A2(n16965), .A3(n16964), .A4(n16963), .ZN(
        n16967) );
  NOR2_X1 U20136 ( .A1(n16968), .A2(n16967), .ZN(n17171) );
  INV_X1 U20137 ( .A(n16988), .ZN(n16969) );
  OAI221_X1 U20138 ( .B1(n17070), .B2(n16970), .C1(n17064), .C2(n17171), .A(
        n16969), .ZN(n16971) );
  AND2_X1 U20139 ( .A1(n16972), .A2(n16971), .ZN(P3_U2691) );
  NAND3_X1 U20140 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(P3_EBX_REG_9__SCAN_IN), 
        .A3(P3_EBX_REG_8__SCAN_IN), .ZN(n16973) );
  OAI21_X1 U20141 ( .B1(n17032), .B2(n16973), .A(n17064), .ZN(n17010) );
  AOI22_X1 U20142 ( .A1(n16995), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n9633), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n16986) );
  AOI22_X1 U20143 ( .A1(n16974), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n17020), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n16985) );
  INV_X1 U20144 ( .A(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n20815) );
  AOI22_X1 U20145 ( .A1(n17014), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n17023), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n16976) );
  OAI21_X1 U20146 ( .B1(n13882), .B2(n20815), .A(n16976), .ZN(n16983) );
  AOI22_X1 U20147 ( .A1(n16989), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n17022), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n16981) );
  AOI22_X1 U20148 ( .A1(n16992), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n16977), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n16980) );
  AOI22_X1 U20149 ( .A1(n16998), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n16996), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n16979) );
  AOI22_X1 U20150 ( .A1(n16997), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n16923), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n16978) );
  NAND4_X1 U20151 ( .A1(n16981), .A2(n16980), .A3(n16979), .A4(n16978), .ZN(
        n16982) );
  AOI211_X1 U20152 ( .C1(n17005), .C2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .A(
        n16983), .B(n16982), .ZN(n16984) );
  NAND3_X1 U20153 ( .A1(n16986), .A2(n16985), .A3(n16984), .ZN(n17174) );
  OAI22_X1 U20154 ( .A1(P3_EBX_REG_11__SCAN_IN), .A2(n17010), .B1(n17174), 
        .B2(n17064), .ZN(n16987) );
  NOR2_X1 U20155 ( .A1(n16988), .A2(n16987), .ZN(P3_U2692) );
  AOI22_X1 U20156 ( .A1(n16989), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n17023), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n17008) );
  AOI22_X1 U20157 ( .A1(n16990), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n17022), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n17007) );
  AOI22_X1 U20158 ( .A1(n16992), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n16991), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n16993) );
  OAI21_X1 U20159 ( .B1(n16994), .B2(n17061), .A(n16993), .ZN(n17004) );
  AOI22_X1 U20160 ( .A1(n16995), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n16974), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n17002) );
  AOI22_X1 U20161 ( .A1(n16997), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n16996), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n17001) );
  AOI22_X1 U20162 ( .A1(n9633), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n17020), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n17000) );
  AOI22_X1 U20163 ( .A1(n16998), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n16923), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n16999) );
  NAND4_X1 U20164 ( .A1(n17002), .A2(n17001), .A3(n17000), .A4(n16999), .ZN(
        n17003) );
  AOI211_X1 U20165 ( .C1(n17005), .C2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .A(
        n17004), .B(n17003), .ZN(n17006) );
  NAND3_X1 U20166 ( .A1(n17008), .A2(n17007), .A3(n17006), .ZN(n17177) );
  INV_X1 U20167 ( .A(n17177), .ZN(n17012) );
  NOR2_X1 U20168 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n17009), .ZN(n17011) );
  OAI22_X1 U20169 ( .A1(n17012), .A2(n17064), .B1(n17011), .B2(n17010), .ZN(
        P3_U2693) );
  AOI22_X1 U20170 ( .A1(n16997), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n16996), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n17018) );
  AOI22_X1 U20171 ( .A1(n17005), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n17013), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n17017) );
  AOI22_X1 U20172 ( .A1(n16977), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n16995), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n17016) );
  AOI22_X1 U20173 ( .A1(n16992), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n17014), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n17015) );
  NAND4_X1 U20174 ( .A1(n17018), .A2(n17017), .A3(n17016), .A4(n17015), .ZN(
        n17030) );
  AOI22_X1 U20175 ( .A1(n16989), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n9626), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n17028) );
  AOI22_X1 U20176 ( .A1(n17021), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n17020), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n17027) );
  AOI22_X1 U20177 ( .A1(n17023), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n17022), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n17026) );
  AOI22_X1 U20178 ( .A1(n9627), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n9633), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n17025) );
  NAND4_X1 U20179 ( .A1(n17028), .A2(n17027), .A3(n17026), .A4(n17025), .ZN(
        n17029) );
  NOR2_X1 U20180 ( .A1(n17030), .A2(n17029), .ZN(n17191) );
  NOR2_X1 U20181 ( .A1(n17070), .A2(n17031), .ZN(n17037) );
  NOR2_X1 U20182 ( .A1(n17123), .A2(n17032), .ZN(n17034) );
  AOI22_X1 U20183 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n17037), .B1(n17034), .B2(
        n17033), .ZN(n17035) );
  OAI21_X1 U20184 ( .B1(n17191), .B2(n17064), .A(n17035), .ZN(P3_U2695) );
  INV_X1 U20185 ( .A(P3_EBX_REG_6__SCAN_IN), .ZN(n17036) );
  NOR4_X1 U20186 ( .A1(n17036), .A2(n17040), .A3(n17048), .A4(n17067), .ZN(
        n17043) );
  OAI21_X1 U20187 ( .B1(P3_EBX_REG_7__SCAN_IN), .B2(n17043), .A(n17037), .ZN(
        n17038) );
  OAI21_X1 U20188 ( .B1(n17064), .B2(n17039), .A(n17038), .ZN(P3_U2696) );
  NOR3_X1 U20189 ( .A1(n17040), .A2(n17048), .A3(n17067), .ZN(n17047) );
  AOI21_X1 U20190 ( .B1(P3_EBX_REG_6__SCAN_IN), .B2(n17064), .A(n17047), .ZN(
        n17042) );
  INV_X1 U20191 ( .A(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n17041) );
  OAI22_X1 U20192 ( .A1(n17043), .A2(n17042), .B1(n17041), .B2(n17064), .ZN(
        P3_U2697) );
  OAI21_X1 U20193 ( .B1(P3_EBX_REG_5__SCAN_IN), .B2(n17044), .A(n17064), .ZN(
        n17046) );
  INV_X1 U20194 ( .A(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n17045) );
  OAI22_X1 U20195 ( .A1(n17047), .A2(n17046), .B1(n17045), .B2(n17064), .ZN(
        P3_U2698) );
  NOR2_X1 U20196 ( .A1(n17048), .A2(n17067), .ZN(n17053) );
  INV_X1 U20197 ( .A(n17067), .ZN(n17069) );
  NAND2_X1 U20198 ( .A1(n17049), .A2(n17069), .ZN(n17058) );
  NOR2_X1 U20199 ( .A1(n17050), .A2(n17058), .ZN(n17057) );
  AOI21_X1 U20200 ( .B1(P3_EBX_REG_4__SCAN_IN), .B2(n17064), .A(n17057), .ZN(
        n17052) );
  OAI22_X1 U20201 ( .A1(n17053), .A2(n17052), .B1(n17051), .B2(n17064), .ZN(
        P3_U2699) );
  INV_X1 U20202 ( .A(n17058), .ZN(n17054) );
  AOI21_X1 U20203 ( .B1(P3_EBX_REG_3__SCAN_IN), .B2(n17064), .A(n17054), .ZN(
        n17056) );
  INV_X1 U20204 ( .A(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n17055) );
  OAI22_X1 U20205 ( .A1(n17057), .A2(n17056), .B1(n17055), .B2(n17064), .ZN(
        P3_U2700) );
  INV_X1 U20206 ( .A(n17062), .ZN(n17059) );
  OAI221_X1 U20207 ( .B1(P3_EBX_REG_2__SCAN_IN), .B2(n17073), .C1(
        P3_EBX_REG_2__SCAN_IN), .C2(n17059), .A(n17058), .ZN(n17060) );
  AOI22_X1 U20208 ( .A1(n17070), .A2(n17061), .B1(n17060), .B2(n17064), .ZN(
        P3_U2701) );
  NAND2_X1 U20209 ( .A1(n17063), .A2(n17062), .ZN(n17068) );
  OAI222_X1 U20210 ( .A1(n17068), .A2(n17067), .B1(n17066), .B2(n17073), .C1(
        n17065), .C2(n17064), .ZN(P3_U2702) );
  AOI22_X1 U20211 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n17070), .B1(
        n17069), .B2(n17072), .ZN(n17071) );
  OAI21_X1 U20212 ( .B1(n17073), .B2(n17072), .A(n17071), .ZN(P3_U2703) );
  INV_X1 U20213 ( .A(P3_EAX_REG_28__SCAN_IN), .ZN(n17232) );
  INV_X1 U20214 ( .A(P3_EAX_REG_26__SCAN_IN), .ZN(n17235) );
  INV_X1 U20215 ( .A(P3_EAX_REG_19__SCAN_IN), .ZN(n20833) );
  INV_X1 U20216 ( .A(P3_EAX_REG_15__SCAN_IN), .ZN(n17339) );
  INV_X1 U20217 ( .A(P3_EAX_REG_8__SCAN_IN), .ZN(n17269) );
  INV_X1 U20218 ( .A(P3_EAX_REG_1__SCAN_IN), .ZN(n17312) );
  NAND4_X1 U20219 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(P3_EAX_REG_4__SCAN_IN), 
        .A3(P3_EAX_REG_3__SCAN_IN), .A4(P3_EAX_REG_2__SCAN_IN), .ZN(n17074) );
  NOR3_X1 U20220 ( .A1(n17312), .A2(n17288), .A3(n17074), .ZN(n17075) );
  NAND3_X1 U20221 ( .A1(P3_EAX_REG_7__SCAN_IN), .A2(P3_EAX_REG_6__SCAN_IN), 
        .A3(n17075), .ZN(n17192) );
  NOR2_X1 U20222 ( .A1(n17269), .A2(n17192), .ZN(n17187) );
  NAND2_X1 U20223 ( .A1(n17186), .A2(n17187), .ZN(n17181) );
  NAND3_X1 U20224 ( .A1(P3_EAX_REG_13__SCAN_IN), .A2(P3_EAX_REG_12__SCAN_IN), 
        .A3(P3_EAX_REG_11__SCAN_IN), .ZN(n17162) );
  NOR2_X1 U20225 ( .A1(n17181), .A2(n17162), .ZN(n17076) );
  NAND4_X1 U20226 ( .A1(P3_EAX_REG_9__SCAN_IN), .A2(P3_EAX_REG_14__SCAN_IN), 
        .A3(P3_EAX_REG_10__SCAN_IN), .A4(n17076), .ZN(n17163) );
  INV_X1 U20227 ( .A(P3_EAX_REG_22__SCAN_IN), .ZN(n17243) );
  NAND4_X1 U20228 ( .A1(P3_EAX_REG_21__SCAN_IN), .A2(P3_EAX_REG_20__SCAN_IN), 
        .A3(P3_EAX_REG_18__SCAN_IN), .A4(P3_EAX_REG_17__SCAN_IN), .ZN(n17077)
         );
  NAND2_X1 U20229 ( .A1(P3_EAX_REG_23__SCAN_IN), .A2(n17118), .ZN(n17117) );
  NAND2_X1 U20230 ( .A1(P3_EAX_REG_24__SCAN_IN), .A2(n17113), .ZN(n17112) );
  NAND2_X1 U20231 ( .A1(P3_EAX_REG_29__SCAN_IN), .A2(n17092), .ZN(n17087) );
  INV_X1 U20232 ( .A(P3_EAX_REG_30__SCAN_IN), .ZN(n17309) );
  OR2_X1 U20233 ( .A1(n17087), .A2(n17309), .ZN(n17081) );
  NOR2_X2 U20234 ( .A1(n17078), .A2(n17213), .ZN(n17152) );
  NAND2_X1 U20235 ( .A1(n17213), .A2(n17087), .ZN(n17086) );
  OAI21_X1 U20236 ( .B1(P3_EAX_REG_30__SCAN_IN), .B2(n17211), .A(n17086), .ZN(
        n17079) );
  AOI22_X1 U20237 ( .A1(BUF2_REG_31__SCAN_IN), .A2(n17152), .B1(
        P3_EAX_REG_31__SCAN_IN), .B2(n17079), .ZN(n17080) );
  OAI21_X1 U20238 ( .B1(P3_EAX_REG_31__SCAN_IN), .B2(n17081), .A(n17080), .ZN(
        P3_U2704) );
  NOR2_X2 U20239 ( .A1(n17082), .A2(n17213), .ZN(n17153) );
  INV_X1 U20240 ( .A(n17152), .ZN(n17128) );
  OAI22_X1 U20241 ( .A1(n17083), .A2(n17214), .B1(n18079), .B2(n17128), .ZN(
        n17084) );
  AOI21_X1 U20242 ( .B1(BUF2_REG_14__SCAN_IN), .B2(n17153), .A(n17084), .ZN(
        n17085) );
  OAI221_X1 U20243 ( .B1(P3_EAX_REG_30__SCAN_IN), .B2(n17087), .C1(n17309), 
        .C2(n17086), .A(n17085), .ZN(P3_U2705) );
  AOI22_X1 U20244 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17153), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n17152), .ZN(n17089) );
  OAI211_X1 U20245 ( .C1(n17092), .C2(P3_EAX_REG_29__SCAN_IN), .A(n17213), .B(
        n17087), .ZN(n17088) );
  OAI211_X1 U20246 ( .C1(n17090), .C2(n17214), .A(n17089), .B(n17088), .ZN(
        P3_U2706) );
  AOI22_X1 U20247 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n17153), .B1(n17221), .B2(
        n17091), .ZN(n17095) );
  AOI211_X1 U20248 ( .C1(n17232), .C2(n17097), .A(n17092), .B(n17180), .ZN(
        n17093) );
  INV_X1 U20249 ( .A(n17093), .ZN(n17094) );
  OAI211_X1 U20250 ( .C1(n17128), .C2(n17096), .A(n17095), .B(n17094), .ZN(
        P3_U2707) );
  AOI22_X1 U20251 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17153), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n17152), .ZN(n17099) );
  OAI211_X1 U20252 ( .C1(n17102), .C2(P3_EAX_REG_27__SCAN_IN), .A(n17213), .B(
        n17097), .ZN(n17098) );
  OAI211_X1 U20253 ( .C1(n17100), .C2(n17214), .A(n17099), .B(n17098), .ZN(
        P3_U2708) );
  AOI22_X1 U20254 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17153), .B1(n17221), .B2(
        n17101), .ZN(n17105) );
  AOI211_X1 U20255 ( .C1(n17235), .C2(n17106), .A(n17102), .B(n17180), .ZN(
        n17103) );
  INV_X1 U20256 ( .A(n17103), .ZN(n17104) );
  OAI211_X1 U20257 ( .C1(n17128), .C2(n18060), .A(n17105), .B(n17104), .ZN(
        P3_U2709) );
  AOI22_X1 U20258 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n17153), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n17152), .ZN(n17109) );
  OAI211_X1 U20259 ( .C1(n17107), .C2(P3_EAX_REG_25__SCAN_IN), .A(n17213), .B(
        n17106), .ZN(n17108) );
  OAI211_X1 U20260 ( .C1(n17110), .C2(n17214), .A(n17109), .B(n17108), .ZN(
        P3_U2710) );
  INV_X1 U20261 ( .A(n17153), .ZN(n17116) );
  AOI22_X1 U20262 ( .A1(BUF2_REG_24__SCAN_IN), .A2(n17152), .B1(n17221), .B2(
        n17111), .ZN(n17115) );
  OAI211_X1 U20263 ( .C1(n17113), .C2(P3_EAX_REG_24__SCAN_IN), .A(n17213), .B(
        n17112), .ZN(n17114) );
  OAI211_X1 U20264 ( .C1(n17116), .C2(n17320), .A(n17115), .B(n17114), .ZN(
        P3_U2711) );
  AOI22_X1 U20265 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n17153), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n17152), .ZN(n17120) );
  OAI211_X1 U20266 ( .C1(P3_EAX_REG_23__SCAN_IN), .C2(n17118), .A(n17213), .B(
        n17117), .ZN(n17119) );
  OAI211_X1 U20267 ( .C1(n17121), .C2(n17214), .A(n17120), .B(n17119), .ZN(
        P3_U2712) );
  AOI22_X1 U20268 ( .A1(BUF2_REG_22__SCAN_IN), .A2(n17152), .B1(n17221), .B2(
        n17122), .ZN(n17127) );
  INV_X1 U20269 ( .A(P3_EAX_REG_17__SCAN_IN), .ZN(n17294) );
  NAND2_X1 U20270 ( .A1(P3_EAX_REG_18__SCAN_IN), .A2(n17146), .ZN(n17142) );
  NAND2_X1 U20271 ( .A1(P3_EAX_REG_20__SCAN_IN), .A2(n17137), .ZN(n17133) );
  NAND2_X1 U20272 ( .A1(n17213), .A2(n17133), .ZN(n17132) );
  OAI21_X1 U20273 ( .B1(P3_EAX_REG_21__SCAN_IN), .B2(n17211), .A(n17132), .ZN(
        n17124) );
  AOI22_X1 U20274 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n17153), .B1(
        P3_EAX_REG_22__SCAN_IN), .B2(n17124), .ZN(n17126) );
  NAND4_X1 U20275 ( .A1(P3_EAX_REG_20__SCAN_IN), .A2(P3_EAX_REG_21__SCAN_IN), 
        .A3(n17137), .A4(n17243), .ZN(n17125) );
  NAND3_X1 U20276 ( .A1(n17127), .A2(n17126), .A3(n17125), .ZN(P3_U2713) );
  INV_X1 U20277 ( .A(P3_EAX_REG_21__SCAN_IN), .ZN(n17245) );
  OAI22_X1 U20278 ( .A1(n17129), .A2(n17214), .B1(n18073), .B2(n17128), .ZN(
        n17130) );
  AOI21_X1 U20279 ( .B1(BUF2_REG_5__SCAN_IN), .B2(n17153), .A(n17130), .ZN(
        n17131) );
  OAI221_X1 U20280 ( .B1(P3_EAX_REG_21__SCAN_IN), .B2(n17133), .C1(n17245), 
        .C2(n17132), .A(n17131), .ZN(P3_U2714) );
  AOI22_X1 U20281 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n17153), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n17152), .ZN(n17135) );
  OAI211_X1 U20282 ( .C1(n17137), .C2(P3_EAX_REG_20__SCAN_IN), .A(n17213), .B(
        n17133), .ZN(n17134) );
  OAI211_X1 U20283 ( .C1(n17136), .C2(n17214), .A(n17135), .B(n17134), .ZN(
        P3_U2715) );
  AOI22_X1 U20284 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n17153), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n17152), .ZN(n17140) );
  AOI211_X1 U20285 ( .C1(n20833), .C2(n17142), .A(n17137), .B(n17180), .ZN(
        n17138) );
  INV_X1 U20286 ( .A(n17138), .ZN(n17139) );
  OAI211_X1 U20287 ( .C1(n17141), .C2(n17214), .A(n17140), .B(n17139), .ZN(
        P3_U2716) );
  AOI22_X1 U20288 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n17153), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n17152), .ZN(n17144) );
  OAI211_X1 U20289 ( .C1(n17146), .C2(P3_EAX_REG_18__SCAN_IN), .A(n17213), .B(
        n17142), .ZN(n17143) );
  OAI211_X1 U20290 ( .C1(n17145), .C2(n17214), .A(n17144), .B(n17143), .ZN(
        P3_U2717) );
  AOI22_X1 U20291 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17153), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n17152), .ZN(n17150) );
  INV_X1 U20292 ( .A(n17154), .ZN(n17148) );
  INV_X1 U20293 ( .A(n17146), .ZN(n17147) );
  OAI211_X1 U20294 ( .C1(n17148), .C2(P3_EAX_REG_17__SCAN_IN), .A(n17213), .B(
        n17147), .ZN(n17149) );
  OAI211_X1 U20295 ( .C1(n17151), .C2(n17214), .A(n17150), .B(n17149), .ZN(
        P3_U2718) );
  AOI22_X1 U20296 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n17153), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n17152), .ZN(n17156) );
  OAI211_X1 U20297 ( .C1(P3_EAX_REG_16__SCAN_IN), .C2(n17158), .A(n17213), .B(
        n17154), .ZN(n17155) );
  OAI211_X1 U20298 ( .C1(n17157), .C2(n17214), .A(n17156), .B(n17155), .ZN(
        P3_U2719) );
  AOI211_X1 U20299 ( .C1(n17339), .C2(n17163), .A(n17180), .B(n17158), .ZN(
        n17159) );
  AOI21_X1 U20300 ( .B1(n17222), .B2(BUF2_REG_15__SCAN_IN), .A(n17159), .ZN(
        n17160) );
  OAI21_X1 U20301 ( .B1(n17161), .B2(n17214), .A(n17160), .ZN(P3_U2720) );
  INV_X1 U20302 ( .A(P3_EAX_REG_10__SCAN_IN), .ZN(n17265) );
  INV_X1 U20303 ( .A(n17211), .ZN(n17218) );
  NAND3_X1 U20304 ( .A1(P3_EAX_REG_9__SCAN_IN), .A2(n17187), .A3(n17218), .ZN(
        n17182) );
  NOR2_X1 U20305 ( .A1(n17162), .A2(n17176), .ZN(n17168) );
  INV_X1 U20306 ( .A(P3_EAX_REG_14__SCAN_IN), .ZN(n17334) );
  AOI22_X1 U20307 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17222), .B1(n17168), .B2(
        n17334), .ZN(n17165) );
  NAND3_X1 U20308 ( .A1(P3_EAX_REG_14__SCAN_IN), .A2(n17213), .A3(n17163), 
        .ZN(n17164) );
  OAI211_X1 U20309 ( .C1(n17166), .C2(n17214), .A(n17165), .B(n17164), .ZN(
        P3_U2721) );
  INV_X1 U20310 ( .A(P3_EAX_REG_11__SCAN_IN), .ZN(n17263) );
  NOR2_X1 U20311 ( .A1(n17263), .A2(n17176), .ZN(n17170) );
  AND2_X1 U20312 ( .A1(P3_EAX_REG_12__SCAN_IN), .A2(n17170), .ZN(n17173) );
  AOI21_X1 U20313 ( .B1(P3_EAX_REG_13__SCAN_IN), .B2(n17213), .A(n17173), .ZN(
        n17169) );
  OAI222_X1 U20314 ( .A1(n17217), .A2(n17332), .B1(n17169), .B2(n17168), .C1(
        n17214), .C2(n17167), .ZN(P3_U2722) );
  AOI21_X1 U20315 ( .B1(P3_EAX_REG_12__SCAN_IN), .B2(n17213), .A(n17170), .ZN(
        n17172) );
  OAI222_X1 U20316 ( .A1(n17217), .A2(n17328), .B1(n17173), .B2(n17172), .C1(
        n17214), .C2(n17171), .ZN(P3_U2723) );
  NAND2_X1 U20317 ( .A1(n17213), .A2(n17176), .ZN(n17179) );
  AOI22_X1 U20318 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17222), .B1(n17221), .B2(
        n17174), .ZN(n17175) );
  OAI221_X1 U20319 ( .B1(P3_EAX_REG_11__SCAN_IN), .B2(n17176), .C1(n17263), 
        .C2(n17179), .A(n17175), .ZN(P3_U2724) );
  AOI22_X1 U20320 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17222), .B1(n17221), .B2(
        n17177), .ZN(n17178) );
  OAI221_X1 U20321 ( .B1(n17179), .B2(n17265), .C1(n17179), .C2(n17182), .A(
        n17178), .ZN(P3_U2725) );
  INV_X1 U20322 ( .A(P3_EAX_REG_9__SCAN_IN), .ZN(n17267) );
  AOI21_X1 U20323 ( .B1(n17267), .B2(n17181), .A(n17180), .ZN(n17183) );
  AOI22_X1 U20324 ( .A1(n17221), .A2(n17184), .B1(n17183), .B2(n17182), .ZN(
        n17185) );
  OAI21_X1 U20325 ( .B1(n13109), .B2(n17217), .A(n17185), .ZN(P3_U2726) );
  INV_X1 U20326 ( .A(n17186), .ZN(n17219) );
  AOI22_X1 U20327 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17222), .B1(
        P3_EAX_REG_8__SCAN_IN), .B2(n17219), .ZN(n17190) );
  AOI211_X1 U20328 ( .C1(n17269), .C2(n17192), .A(n17211), .B(n17187), .ZN(
        n17188) );
  INV_X1 U20329 ( .A(n17188), .ZN(n17189) );
  OAI211_X1 U20330 ( .C1(n17191), .C2(n17214), .A(n17190), .B(n17189), .ZN(
        P3_U2727) );
  NOR2_X1 U20331 ( .A1(n17192), .A2(n17211), .ZN(n17196) );
  INV_X1 U20332 ( .A(P3_EAX_REG_6__SCAN_IN), .ZN(n17273) );
  INV_X1 U20333 ( .A(P3_EAX_REG_4__SCAN_IN), .ZN(n17277) );
  INV_X1 U20334 ( .A(P3_EAX_REG_2__SCAN_IN), .ZN(n17282) );
  NOR4_X1 U20335 ( .A1(n17282), .A2(n17312), .A3(n17288), .A4(n17211), .ZN(
        n17216) );
  NAND2_X1 U20336 ( .A1(P3_EAX_REG_3__SCAN_IN), .A2(n17216), .ZN(n17204) );
  NOR2_X1 U20337 ( .A1(n17277), .A2(n17204), .ZN(n17207) );
  NAND2_X1 U20338 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(n17207), .ZN(n17197) );
  NOR2_X1 U20339 ( .A1(n17273), .A2(n17197), .ZN(n17200) );
  AOI21_X1 U20340 ( .B1(P3_EAX_REG_7__SCAN_IN), .B2(n17213), .A(n17200), .ZN(
        n17195) );
  INV_X1 U20341 ( .A(n17193), .ZN(n17194) );
  OAI222_X1 U20342 ( .A1(n17217), .A2(n18084), .B1(n17196), .B2(n17195), .C1(
        n17214), .C2(n17194), .ZN(P3_U2728) );
  INV_X1 U20343 ( .A(n17197), .ZN(n17203) );
  AOI21_X1 U20344 ( .B1(P3_EAX_REG_6__SCAN_IN), .B2(n17213), .A(n17203), .ZN(
        n17199) );
  OAI222_X1 U20345 ( .A1(n18080), .A2(n17217), .B1(n17200), .B2(n17199), .C1(
        n17214), .C2(n17198), .ZN(P3_U2729) );
  AOI21_X1 U20346 ( .B1(P3_EAX_REG_5__SCAN_IN), .B2(n17213), .A(n17207), .ZN(
        n17202) );
  OAI222_X1 U20347 ( .A1(n18072), .A2(n17217), .B1(n17203), .B2(n17202), .C1(
        n17214), .C2(n17201), .ZN(P3_U2730) );
  INV_X1 U20348 ( .A(n17204), .ZN(n17210) );
  AOI21_X1 U20349 ( .B1(P3_EAX_REG_4__SCAN_IN), .B2(n17213), .A(n17210), .ZN(
        n17206) );
  OAI222_X1 U20350 ( .A1(n18067), .A2(n17217), .B1(n17207), .B2(n17206), .C1(
        n17214), .C2(n17205), .ZN(P3_U2731) );
  AOI21_X1 U20351 ( .B1(P3_EAX_REG_3__SCAN_IN), .B2(n17213), .A(n17216), .ZN(
        n17209) );
  OAI222_X1 U20352 ( .A1(n18064), .A2(n17217), .B1(n17210), .B2(n17209), .C1(
        n17214), .C2(n17208), .ZN(P3_U2732) );
  NOR3_X1 U20353 ( .A1(n17312), .A2(n17288), .A3(n17211), .ZN(n17212) );
  AOI21_X1 U20354 ( .B1(P3_EAX_REG_2__SCAN_IN), .B2(n17213), .A(n17212), .ZN(
        n17215) );
  OAI222_X1 U20355 ( .A1(n18059), .A2(n17217), .B1(n17216), .B2(n17215), .C1(
        n17214), .C2(n9612), .ZN(P3_U2733) );
  NAND2_X1 U20356 ( .A1(P3_EAX_REG_0__SCAN_IN), .A2(n17218), .ZN(n17225) );
  AOI21_X1 U20357 ( .B1(n18087), .B2(n17288), .A(n17219), .ZN(n17224) );
  AOI22_X1 U20358 ( .A1(n17222), .A2(BUF2_REG_1__SCAN_IN), .B1(n17221), .B2(
        n17220), .ZN(n17223) );
  OAI221_X1 U20359 ( .B1(P3_EAX_REG_1__SCAN_IN), .B2(n17225), .C1(n17312), 
        .C2(n17224), .A(n17223), .ZN(P3_U2734) );
  NAND2_X1 U20360 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(n17549), .ZN(n18687) );
  AND2_X1 U20361 ( .A1(n17278), .A2(P3_DATAO_REG_31__SCAN_IN), .ZN(P3_U2736)
         );
  NAND2_X1 U20362 ( .A1(n17255), .A2(n17227), .ZN(n17253) );
  AOI22_X1 U20363 ( .A1(n17285), .A2(P3_UWORD_REG_14__SCAN_IN), .B1(n17284), 
        .B2(P3_DATAO_REG_30__SCAN_IN), .ZN(n17228) );
  OAI21_X1 U20364 ( .B1(n17309), .B2(n17253), .A(n17228), .ZN(P3_U2737) );
  INV_X1 U20365 ( .A(P3_EAX_REG_29__SCAN_IN), .ZN(n17230) );
  AOI22_X1 U20366 ( .A1(n17285), .A2(P3_UWORD_REG_13__SCAN_IN), .B1(n17284), 
        .B2(P3_DATAO_REG_29__SCAN_IN), .ZN(n17229) );
  OAI21_X1 U20367 ( .B1(n17230), .B2(n17253), .A(n17229), .ZN(P3_U2738) );
  AOI22_X1 U20368 ( .A1(n17285), .A2(P3_UWORD_REG_12__SCAN_IN), .B1(n17278), 
        .B2(P3_DATAO_REG_28__SCAN_IN), .ZN(n17231) );
  OAI21_X1 U20369 ( .B1(n17232), .B2(n17253), .A(n17231), .ZN(P3_U2739) );
  INV_X1 U20370 ( .A(P3_EAX_REG_27__SCAN_IN), .ZN(n17305) );
  AOI22_X1 U20371 ( .A1(P3_UWORD_REG_11__SCAN_IN), .A2(n17285), .B1(n17278), 
        .B2(P3_DATAO_REG_27__SCAN_IN), .ZN(n17233) );
  OAI21_X1 U20372 ( .B1(n17305), .B2(n17253), .A(n17233), .ZN(P3_U2740) );
  AOI22_X1 U20373 ( .A1(P3_UWORD_REG_10__SCAN_IN), .A2(n17285), .B1(n17278), 
        .B2(P3_DATAO_REG_26__SCAN_IN), .ZN(n17234) );
  OAI21_X1 U20374 ( .B1(n17235), .B2(n17253), .A(n17234), .ZN(P3_U2741) );
  INV_X1 U20375 ( .A(P3_EAX_REG_25__SCAN_IN), .ZN(n17237) );
  AOI22_X1 U20376 ( .A1(n17285), .A2(P3_UWORD_REG_9__SCAN_IN), .B1(n17284), 
        .B2(P3_DATAO_REG_25__SCAN_IN), .ZN(n17236) );
  OAI21_X1 U20377 ( .B1(n17237), .B2(n17253), .A(n17236), .ZN(P3_U2742) );
  INV_X1 U20378 ( .A(P3_EAX_REG_24__SCAN_IN), .ZN(n17239) );
  AOI22_X1 U20379 ( .A1(n17285), .A2(P3_UWORD_REG_8__SCAN_IN), .B1(n17278), 
        .B2(P3_DATAO_REG_24__SCAN_IN), .ZN(n17238) );
  OAI21_X1 U20380 ( .B1(n17239), .B2(n17253), .A(n17238), .ZN(P3_U2743) );
  INV_X1 U20381 ( .A(P3_EAX_REG_23__SCAN_IN), .ZN(n17241) );
  AOI22_X1 U20382 ( .A1(n17285), .A2(P3_UWORD_REG_7__SCAN_IN), .B1(n17284), 
        .B2(P3_DATAO_REG_23__SCAN_IN), .ZN(n17240) );
  OAI21_X1 U20383 ( .B1(n17241), .B2(n17253), .A(n17240), .ZN(P3_U2744) );
  AOI22_X1 U20384 ( .A1(n17285), .A2(P3_UWORD_REG_6__SCAN_IN), .B1(n17284), 
        .B2(P3_DATAO_REG_22__SCAN_IN), .ZN(n17242) );
  OAI21_X1 U20385 ( .B1(n17243), .B2(n17253), .A(n17242), .ZN(P3_U2745) );
  AOI22_X1 U20386 ( .A1(n17285), .A2(P3_UWORD_REG_5__SCAN_IN), .B1(n17284), 
        .B2(P3_DATAO_REG_21__SCAN_IN), .ZN(n17244) );
  OAI21_X1 U20387 ( .B1(n17245), .B2(n17253), .A(n17244), .ZN(P3_U2746) );
  INV_X1 U20388 ( .A(P3_EAX_REG_20__SCAN_IN), .ZN(n17247) );
  AOI22_X1 U20389 ( .A1(n17285), .A2(P3_UWORD_REG_4__SCAN_IN), .B1(n17284), 
        .B2(P3_DATAO_REG_20__SCAN_IN), .ZN(n17246) );
  OAI21_X1 U20390 ( .B1(n17247), .B2(n17253), .A(n17246), .ZN(P3_U2747) );
  AOI22_X1 U20391 ( .A1(n17285), .A2(P3_UWORD_REG_3__SCAN_IN), .B1(n17284), 
        .B2(P3_DATAO_REG_19__SCAN_IN), .ZN(n17248) );
  OAI21_X1 U20392 ( .B1(n20833), .B2(n17253), .A(n17248), .ZN(P3_U2748) );
  INV_X1 U20393 ( .A(P3_EAX_REG_18__SCAN_IN), .ZN(n17250) );
  AOI22_X1 U20394 ( .A1(n17285), .A2(P3_UWORD_REG_2__SCAN_IN), .B1(n17284), 
        .B2(P3_DATAO_REG_18__SCAN_IN), .ZN(n17249) );
  OAI21_X1 U20395 ( .B1(n17250), .B2(n17253), .A(n17249), .ZN(P3_U2749) );
  AOI22_X1 U20396 ( .A1(P3_UWORD_REG_1__SCAN_IN), .A2(n17285), .B1(n17284), 
        .B2(P3_DATAO_REG_17__SCAN_IN), .ZN(n17251) );
  OAI21_X1 U20397 ( .B1(n17294), .B2(n17253), .A(n17251), .ZN(P3_U2750) );
  INV_X1 U20398 ( .A(P3_EAX_REG_16__SCAN_IN), .ZN(n17254) );
  AOI22_X1 U20399 ( .A1(n17285), .A2(P3_UWORD_REG_0__SCAN_IN), .B1(n17284), 
        .B2(P3_DATAO_REG_16__SCAN_IN), .ZN(n17252) );
  OAI21_X1 U20400 ( .B1(n17254), .B2(n17253), .A(n17252), .ZN(P3_U2751) );
  AOI22_X1 U20401 ( .A1(n17285), .A2(P3_LWORD_REG_15__SCAN_IN), .B1(n17284), 
        .B2(P3_DATAO_REG_15__SCAN_IN), .ZN(n17256) );
  OAI21_X1 U20402 ( .B1(n17339), .B2(n17287), .A(n17256), .ZN(P3_U2752) );
  AOI22_X1 U20403 ( .A1(n17285), .A2(P3_LWORD_REG_14__SCAN_IN), .B1(n17284), 
        .B2(P3_DATAO_REG_14__SCAN_IN), .ZN(n17257) );
  OAI21_X1 U20404 ( .B1(n17334), .B2(n17287), .A(n17257), .ZN(P3_U2753) );
  INV_X1 U20405 ( .A(P3_EAX_REG_13__SCAN_IN), .ZN(n17259) );
  AOI22_X1 U20406 ( .A1(n17285), .A2(P3_LWORD_REG_13__SCAN_IN), .B1(n17284), 
        .B2(P3_DATAO_REG_13__SCAN_IN), .ZN(n17258) );
  OAI21_X1 U20407 ( .B1(n17259), .B2(n17287), .A(n17258), .ZN(P3_U2754) );
  INV_X1 U20408 ( .A(P3_EAX_REG_12__SCAN_IN), .ZN(n17261) );
  AOI22_X1 U20409 ( .A1(n17285), .A2(P3_LWORD_REG_12__SCAN_IN), .B1(n17278), 
        .B2(P3_DATAO_REG_12__SCAN_IN), .ZN(n17260) );
  OAI21_X1 U20410 ( .B1(n17261), .B2(n17287), .A(n17260), .ZN(P3_U2755) );
  AOI22_X1 U20411 ( .A1(P3_LWORD_REG_11__SCAN_IN), .A2(n17285), .B1(n17284), 
        .B2(P3_DATAO_REG_11__SCAN_IN), .ZN(n17262) );
  OAI21_X1 U20412 ( .B1(n17263), .B2(n17287), .A(n17262), .ZN(P3_U2756) );
  AOI22_X1 U20413 ( .A1(n17285), .A2(P3_LWORD_REG_10__SCAN_IN), .B1(n17278), 
        .B2(P3_DATAO_REG_10__SCAN_IN), .ZN(n17264) );
  OAI21_X1 U20414 ( .B1(n17265), .B2(n17287), .A(n17264), .ZN(P3_U2757) );
  AOI22_X1 U20415 ( .A1(P3_LWORD_REG_9__SCAN_IN), .A2(n17285), .B1(n17284), 
        .B2(P3_DATAO_REG_9__SCAN_IN), .ZN(n17266) );
  OAI21_X1 U20416 ( .B1(n17267), .B2(n17287), .A(n17266), .ZN(P3_U2758) );
  AOI22_X1 U20417 ( .A1(P3_DATAO_REG_8__SCAN_IN), .A2(n17284), .B1(n17285), 
        .B2(P3_LWORD_REG_8__SCAN_IN), .ZN(n17268) );
  OAI21_X1 U20418 ( .B1(n17269), .B2(n17287), .A(n17268), .ZN(P3_U2759) );
  INV_X1 U20419 ( .A(P3_EAX_REG_7__SCAN_IN), .ZN(n17271) );
  AOI22_X1 U20420 ( .A1(n17285), .A2(P3_LWORD_REG_7__SCAN_IN), .B1(n17278), 
        .B2(P3_DATAO_REG_7__SCAN_IN), .ZN(n17270) );
  OAI21_X1 U20421 ( .B1(n17271), .B2(n17287), .A(n17270), .ZN(P3_U2760) );
  AOI22_X1 U20422 ( .A1(n17285), .A2(P3_LWORD_REG_6__SCAN_IN), .B1(n17278), 
        .B2(P3_DATAO_REG_6__SCAN_IN), .ZN(n17272) );
  OAI21_X1 U20423 ( .B1(n17273), .B2(n17287), .A(n17272), .ZN(P3_U2761) );
  INV_X1 U20424 ( .A(P3_EAX_REG_5__SCAN_IN), .ZN(n17275) );
  AOI22_X1 U20425 ( .A1(n17285), .A2(P3_LWORD_REG_5__SCAN_IN), .B1(n17278), 
        .B2(P3_DATAO_REG_5__SCAN_IN), .ZN(n17274) );
  OAI21_X1 U20426 ( .B1(n17275), .B2(n17287), .A(n17274), .ZN(P3_U2762) );
  AOI22_X1 U20427 ( .A1(P3_DATAO_REG_4__SCAN_IN), .A2(n17284), .B1(n17285), 
        .B2(P3_LWORD_REG_4__SCAN_IN), .ZN(n17276) );
  OAI21_X1 U20428 ( .B1(n17277), .B2(n17287), .A(n17276), .ZN(P3_U2763) );
  INV_X1 U20429 ( .A(P3_EAX_REG_3__SCAN_IN), .ZN(n17280) );
  AOI22_X1 U20430 ( .A1(n17285), .A2(P3_LWORD_REG_3__SCAN_IN), .B1(n17278), 
        .B2(P3_DATAO_REG_3__SCAN_IN), .ZN(n17279) );
  OAI21_X1 U20431 ( .B1(n17280), .B2(n17287), .A(n17279), .ZN(P3_U2764) );
  AOI22_X1 U20432 ( .A1(n17285), .A2(P3_LWORD_REG_2__SCAN_IN), .B1(n17284), 
        .B2(P3_DATAO_REG_2__SCAN_IN), .ZN(n17281) );
  OAI21_X1 U20433 ( .B1(n17282), .B2(n17287), .A(n17281), .ZN(P3_U2765) );
  AOI22_X1 U20434 ( .A1(n17285), .A2(P3_LWORD_REG_1__SCAN_IN), .B1(n17284), 
        .B2(P3_DATAO_REG_1__SCAN_IN), .ZN(n17283) );
  OAI21_X1 U20435 ( .B1(n17312), .B2(n17287), .A(n17283), .ZN(P3_U2766) );
  AOI22_X1 U20436 ( .A1(n17285), .A2(P3_LWORD_REG_0__SCAN_IN), .B1(n17284), 
        .B2(P3_DATAO_REG_0__SCAN_IN), .ZN(n17286) );
  OAI21_X1 U20437 ( .B1(n17288), .B2(n17287), .A(n17286), .ZN(P3_U2767) );
  AOI221_X1 U20438 ( .B1(n18688), .B2(n18481), .C1(n17290), .C2(n18481), .A(
        n17289), .ZN(n17326) );
  AND2_X1 U20439 ( .A1(n17326), .A2(n17291), .ZN(n17336) );
  INV_X2 U20440 ( .A(n17326), .ZN(n17335) );
  AOI22_X1 U20441 ( .A1(P3_EAX_REG_16__SCAN_IN), .A2(n17329), .B1(
        P3_UWORD_REG_0__SCAN_IN), .B2(n17335), .ZN(n17292) );
  OAI21_X1 U20442 ( .B1(n18048), .B2(n17331), .A(n17292), .ZN(P3_U2768) );
  AOI22_X1 U20443 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17336), .B1(
        P3_UWORD_REG_1__SCAN_IN), .B2(n17335), .ZN(n17293) );
  OAI21_X1 U20444 ( .B1(n17294), .B2(n17338), .A(n17293), .ZN(P3_U2769) );
  AOI22_X1 U20445 ( .A1(P3_EAX_REG_18__SCAN_IN), .A2(n17329), .B1(
        P3_UWORD_REG_2__SCAN_IN), .B2(n17335), .ZN(n17295) );
  OAI21_X1 U20446 ( .B1(n18059), .B2(n17331), .A(n17295), .ZN(P3_U2770) );
  AOI22_X1 U20447 ( .A1(P3_EAX_REG_19__SCAN_IN), .A2(n17329), .B1(
        P3_UWORD_REG_3__SCAN_IN), .B2(n17335), .ZN(n17296) );
  OAI21_X1 U20448 ( .B1(n18064), .B2(n17331), .A(n17296), .ZN(P3_U2771) );
  AOI22_X1 U20449 ( .A1(P3_EAX_REG_20__SCAN_IN), .A2(n17329), .B1(
        P3_UWORD_REG_4__SCAN_IN), .B2(n17335), .ZN(n17297) );
  OAI21_X1 U20450 ( .B1(n18067), .B2(n17331), .A(n17297), .ZN(P3_U2772) );
  AOI22_X1 U20451 ( .A1(P3_EAX_REG_21__SCAN_IN), .A2(n17329), .B1(
        P3_UWORD_REG_5__SCAN_IN), .B2(n17335), .ZN(n17298) );
  OAI21_X1 U20452 ( .B1(n18072), .B2(n17331), .A(n17298), .ZN(P3_U2773) );
  AOI22_X1 U20453 ( .A1(P3_EAX_REG_22__SCAN_IN), .A2(n17329), .B1(
        P3_UWORD_REG_6__SCAN_IN), .B2(n17335), .ZN(n17299) );
  OAI21_X1 U20454 ( .B1(n18080), .B2(n17331), .A(n17299), .ZN(P3_U2774) );
  AOI22_X1 U20455 ( .A1(P3_EAX_REG_23__SCAN_IN), .A2(n17329), .B1(
        P3_UWORD_REG_7__SCAN_IN), .B2(n17335), .ZN(n17300) );
  OAI21_X1 U20456 ( .B1(n18084), .B2(n17331), .A(n17300), .ZN(P3_U2775) );
  AOI22_X1 U20457 ( .A1(P3_EAX_REG_24__SCAN_IN), .A2(n17329), .B1(
        P3_UWORD_REG_8__SCAN_IN), .B2(n17335), .ZN(n17301) );
  OAI21_X1 U20458 ( .B1(n17320), .B2(n17331), .A(n17301), .ZN(P3_U2776) );
  AOI22_X1 U20459 ( .A1(P3_EAX_REG_25__SCAN_IN), .A2(n17329), .B1(
        P3_UWORD_REG_9__SCAN_IN), .B2(n17335), .ZN(n17302) );
  OAI21_X1 U20460 ( .B1(n13109), .B2(n17331), .A(n17302), .ZN(P3_U2777) );
  AOI22_X1 U20461 ( .A1(P3_UWORD_REG_10__SCAN_IN), .A2(n17335), .B1(
        P3_EAX_REG_26__SCAN_IN), .B2(n17329), .ZN(n17303) );
  OAI21_X1 U20462 ( .B1(n17324), .B2(n17331), .A(n17303), .ZN(P3_U2778) );
  AOI22_X1 U20463 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17336), .B1(
        P3_UWORD_REG_11__SCAN_IN), .B2(n17335), .ZN(n17304) );
  OAI21_X1 U20464 ( .B1(n17305), .B2(n17338), .A(n17304), .ZN(P3_U2779) );
  AOI22_X1 U20465 ( .A1(P3_EAX_REG_28__SCAN_IN), .A2(n17329), .B1(
        P3_UWORD_REG_12__SCAN_IN), .B2(n17335), .ZN(n17306) );
  OAI21_X1 U20466 ( .B1(n17328), .B2(n17331), .A(n17306), .ZN(P3_U2780) );
  AOI22_X1 U20467 ( .A1(P3_EAX_REG_29__SCAN_IN), .A2(n17329), .B1(
        P3_UWORD_REG_13__SCAN_IN), .B2(n17335), .ZN(n17307) );
  OAI21_X1 U20468 ( .B1(n17332), .B2(n17331), .A(n17307), .ZN(P3_U2781) );
  AOI22_X1 U20469 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17336), .B1(
        P3_UWORD_REG_14__SCAN_IN), .B2(n17335), .ZN(n17308) );
  OAI21_X1 U20470 ( .B1(n17309), .B2(n17338), .A(n17308), .ZN(P3_U2782) );
  AOI22_X1 U20471 ( .A1(P3_EAX_REG_0__SCAN_IN), .A2(n17329), .B1(
        P3_LWORD_REG_0__SCAN_IN), .B2(n17335), .ZN(n17310) );
  OAI21_X1 U20472 ( .B1(n18048), .B2(n17331), .A(n17310), .ZN(P3_U2783) );
  AOI22_X1 U20473 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17336), .B1(
        P3_LWORD_REG_1__SCAN_IN), .B2(n17335), .ZN(n17311) );
  OAI21_X1 U20474 ( .B1(n17312), .B2(n17338), .A(n17311), .ZN(P3_U2784) );
  AOI22_X1 U20475 ( .A1(P3_EAX_REG_2__SCAN_IN), .A2(n17322), .B1(
        P3_LWORD_REG_2__SCAN_IN), .B2(n17335), .ZN(n17313) );
  OAI21_X1 U20476 ( .B1(n18059), .B2(n17331), .A(n17313), .ZN(P3_U2785) );
  AOI22_X1 U20477 ( .A1(P3_EAX_REG_3__SCAN_IN), .A2(n17322), .B1(
        P3_LWORD_REG_3__SCAN_IN), .B2(n17335), .ZN(n17314) );
  OAI21_X1 U20478 ( .B1(n18064), .B2(n17331), .A(n17314), .ZN(P3_U2786) );
  AOI22_X1 U20479 ( .A1(P3_EAX_REG_4__SCAN_IN), .A2(n17322), .B1(
        P3_LWORD_REG_4__SCAN_IN), .B2(n17335), .ZN(n17315) );
  OAI21_X1 U20480 ( .B1(n18067), .B2(n17331), .A(n17315), .ZN(P3_U2787) );
  AOI22_X1 U20481 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(n17322), .B1(
        P3_LWORD_REG_5__SCAN_IN), .B2(n17335), .ZN(n17316) );
  OAI21_X1 U20482 ( .B1(n18072), .B2(n17331), .A(n17316), .ZN(P3_U2788) );
  AOI22_X1 U20483 ( .A1(P3_EAX_REG_6__SCAN_IN), .A2(n17322), .B1(
        P3_LWORD_REG_6__SCAN_IN), .B2(n17335), .ZN(n17317) );
  OAI21_X1 U20484 ( .B1(n18080), .B2(n17331), .A(n17317), .ZN(P3_U2789) );
  AOI22_X1 U20485 ( .A1(P3_EAX_REG_7__SCAN_IN), .A2(n17322), .B1(
        P3_LWORD_REG_7__SCAN_IN), .B2(n17335), .ZN(n17318) );
  OAI21_X1 U20486 ( .B1(n18084), .B2(n17331), .A(n17318), .ZN(P3_U2790) );
  AOI22_X1 U20487 ( .A1(P3_EAX_REG_8__SCAN_IN), .A2(n17322), .B1(
        P3_LWORD_REG_8__SCAN_IN), .B2(n17335), .ZN(n17319) );
  OAI21_X1 U20488 ( .B1(n17320), .B2(n17331), .A(n17319), .ZN(P3_U2791) );
  AOI22_X1 U20489 ( .A1(P3_LWORD_REG_9__SCAN_IN), .A2(n17335), .B1(
        P3_EAX_REG_9__SCAN_IN), .B2(n17329), .ZN(n17321) );
  OAI21_X1 U20490 ( .B1(n13109), .B2(n17331), .A(n17321), .ZN(P3_U2792) );
  AOI22_X1 U20491 ( .A1(P3_EAX_REG_10__SCAN_IN), .A2(n17322), .B1(
        P3_LWORD_REG_10__SCAN_IN), .B2(n17335), .ZN(n17323) );
  OAI21_X1 U20492 ( .B1(n17324), .B2(n17331), .A(n17323), .ZN(P3_U2793) );
  INV_X1 U20493 ( .A(P3_LWORD_REG_11__SCAN_IN), .ZN(n20889) );
  AOI22_X1 U20494 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17336), .B1(
        P3_EAX_REG_11__SCAN_IN), .B2(n17329), .ZN(n17325) );
  OAI21_X1 U20495 ( .B1(n17326), .B2(n20889), .A(n17325), .ZN(P3_U2794) );
  AOI22_X1 U20496 ( .A1(P3_EAX_REG_12__SCAN_IN), .A2(n17329), .B1(
        P3_LWORD_REG_12__SCAN_IN), .B2(n17335), .ZN(n17327) );
  OAI21_X1 U20497 ( .B1(n17328), .B2(n17331), .A(n17327), .ZN(P3_U2795) );
  AOI22_X1 U20498 ( .A1(P3_EAX_REG_13__SCAN_IN), .A2(n17329), .B1(
        P3_LWORD_REG_13__SCAN_IN), .B2(n17335), .ZN(n17330) );
  OAI21_X1 U20499 ( .B1(n17332), .B2(n17331), .A(n17330), .ZN(P3_U2796) );
  AOI22_X1 U20500 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17336), .B1(
        P3_LWORD_REG_14__SCAN_IN), .B2(n17335), .ZN(n17333) );
  OAI21_X1 U20501 ( .B1(n17334), .B2(n17338), .A(n17333), .ZN(P3_U2797) );
  AOI22_X1 U20502 ( .A1(BUF2_REG_15__SCAN_IN), .A2(n17336), .B1(
        P3_LWORD_REG_15__SCAN_IN), .B2(n17335), .ZN(n17337) );
  OAI21_X1 U20503 ( .B1(n17339), .B2(n17338), .A(n17337), .ZN(P3_U2798) );
  INV_X1 U20504 ( .A(n17707), .ZN(n17680) );
  NOR2_X1 U20505 ( .A1(n17340), .A2(n18554), .ZN(n17341) );
  AOI211_X1 U20506 ( .C1(n17464), .C2(n9749), .A(n17680), .B(n17341), .ZN(
        n17378) );
  OAI21_X1 U20507 ( .B1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n17427), .A(
        n17378), .ZN(n17368) );
  AOI22_X1 U20508 ( .A1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n17368), .B1(
        n17565), .B2(n17342), .ZN(n17362) );
  INV_X1 U20509 ( .A(n17344), .ZN(n17346) );
  AOI21_X1 U20510 ( .B1(n17346), .B2(n17345), .A(n17617), .ZN(n17356) );
  NOR2_X1 U20511 ( .A1(n17697), .A2(n17401), .ZN(n17459) );
  INV_X1 U20512 ( .A(n17347), .ZN(n17718) );
  OAI22_X1 U20513 ( .A1(n17718), .A2(n17710), .B1(n17348), .B2(n17616), .ZN(
        n17383) );
  NOR2_X1 U20514 ( .A1(n17711), .A2(n17383), .ZN(n17350) );
  NOR3_X1 U20515 ( .A1(n17459), .A2(n17350), .A3(n17349), .ZN(n17354) );
  NAND2_X1 U20516 ( .A1(n17971), .A2(P3_REIP_REG_28__SCAN_IN), .ZN(n17360) );
  NAND2_X1 U20517 ( .A1(n17389), .A2(n17544), .ZN(n17406) );
  NOR2_X1 U20518 ( .A1(n17357), .A2(n17406), .ZN(n17370) );
  OAI211_X1 U20519 ( .C1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A(n17370), .B(n17358), .ZN(n17359) );
  NAND4_X1 U20520 ( .A1(n17362), .A2(n17361), .A3(n17360), .A4(n17359), .ZN(
        P3_U2802) );
  NOR2_X1 U20521 ( .A1(n17363), .A2(n17364), .ZN(n17365) );
  XNOR2_X1 U20522 ( .A(n17365), .B(n17615), .ZN(n17725) );
  OAI22_X1 U20523 ( .A1(n18028), .A2(n18623), .B1(n17518), .B2(n17366), .ZN(
        n17367) );
  AOI221_X1 U20524 ( .B1(n17370), .B2(n17369), .C1(n17368), .C2(
        P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A(n17367), .ZN(n17373) );
  AOI22_X1 U20525 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n17383), .B1(
        n17371), .B2(n17711), .ZN(n17372) );
  OAI211_X1 U20526 ( .C1(n17725), .C2(n17617), .A(n17373), .B(n17372), .ZN(
        P3_U2803) );
  AOI21_X1 U20527 ( .B1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n17375), .A(
        n17374), .ZN(n17733) );
  INV_X1 U20528 ( .A(n17427), .ZN(n17376) );
  INV_X1 U20529 ( .A(n17704), .ZN(n17457) );
  NOR2_X1 U20530 ( .A1(n18028), .A2(n18620), .ZN(n17729) );
  INV_X1 U20531 ( .A(n17391), .ZN(n17377) );
  NAND3_X1 U20532 ( .A1(n18426), .A2(n17389), .A3(n17377), .ZN(n17379) );
  AOI21_X1 U20533 ( .B1(n17380), .B2(n17379), .A(n17378), .ZN(n17381) );
  AOI211_X1 U20534 ( .C1(n17382), .C2(n17457), .A(n17729), .B(n17381), .ZN(
        n17385) );
  NOR3_X1 U20535 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n17738), .A3(
        n17748), .ZN(n17731) );
  NOR2_X1 U20536 ( .A1(n17760), .A2(n17424), .ZN(n17409) );
  AOI22_X1 U20537 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n17383), .B1(
        n17731), .B2(n17409), .ZN(n17384) );
  OAI211_X1 U20538 ( .C1(n17733), .C2(n17617), .A(n17385), .B(n17384), .ZN(
        P3_U2804) );
  OAI21_X1 U20539 ( .B1(n17615), .B2(n15210), .A(n17386), .ZN(n17387) );
  XNOR2_X1 U20540 ( .A(n17387), .B(n17738), .ZN(n17747) );
  OAI22_X1 U20541 ( .A1(n17389), .A2(n18078), .B1(n17388), .B2(n18554), .ZN(
        n17390) );
  NOR2_X1 U20542 ( .A1(n17680), .A2(n17390), .ZN(n17416) );
  OAI21_X1 U20543 ( .B1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n18554), .A(
        n17416), .ZN(n17403) );
  NOR2_X1 U20544 ( .A1(n18013), .A2(n18618), .ZN(n17742) );
  OAI21_X1 U20545 ( .B1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A(n17391), .ZN(n17392) );
  OAI22_X1 U20546 ( .A1(n17518), .A2(n17393), .B1(n17406), .B2(n17392), .ZN(
        n17394) );
  AOI211_X1 U20547 ( .C1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .C2(n17403), .A(
        n17742), .B(n17394), .ZN(n17398) );
  XNOR2_X1 U20548 ( .A(n17395), .B(n17738), .ZN(n17743) );
  XNOR2_X1 U20549 ( .A(n17396), .B(n17738), .ZN(n17744) );
  AOI22_X1 U20550 ( .A1(n17697), .A2(n17743), .B1(n17401), .B2(n17744), .ZN(
        n17397) );
  OAI211_X1 U20551 ( .C1(n17617), .C2(n17747), .A(n17398), .B(n17397), .ZN(
        P3_U2805) );
  AOI21_X1 U20552 ( .B1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n17400), .A(
        n17399), .ZN(n17759) );
  AOI22_X1 U20553 ( .A1(n17697), .A2(n17751), .B1(n17401), .B2(n17750), .ZN(
        n17423) );
  INV_X1 U20554 ( .A(n17423), .ZN(n17408) );
  AOI22_X1 U20555 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n17403), .B1(
        n17565), .B2(n17402), .ZN(n17405) );
  NAND2_X1 U20556 ( .A1(n17971), .A2(P3_REIP_REG_24__SCAN_IN), .ZN(n17404) );
  OAI211_X1 U20557 ( .C1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .C2(n17406), .A(
        n17405), .B(n17404), .ZN(n17407) );
  AOI221_X1 U20558 ( .B1(n17409), .B2(n17748), .C1(n17408), .C2(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A(n17407), .ZN(n17410) );
  OAI21_X1 U20559 ( .B1(n17759), .B2(n17617), .A(n17410), .ZN(P3_U2806) );
  OAI21_X1 U20560 ( .B1(n17484), .B2(n17412), .A(n17435), .ZN(n17413) );
  OAI211_X1 U20561 ( .C1(n15213), .C2(n17436), .A(n9635), .B(n17413), .ZN(
        n17414) );
  XNOR2_X1 U20562 ( .A(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .B(n17414), .ZN(
        n17764) );
  NOR2_X1 U20563 ( .A1(n17509), .A2(n17415), .ZN(n17418) );
  INV_X1 U20564 ( .A(n17416), .ZN(n17417) );
  MUX2_X1 U20565 ( .A(n17418), .B(n17417), .S(
        P3_PHYADDRPOINTER_REG_23__SCAN_IN), .Z(n17421) );
  OAI22_X1 U20566 ( .A1(n18028), .A2(n18615), .B1(n17518), .B2(n17419), .ZN(
        n17420) );
  AOI211_X1 U20567 ( .C1(n17605), .C2(n17764), .A(n17421), .B(n17420), .ZN(
        n17422) );
  OAI221_X1 U20568 ( .B1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n17424), 
        .C1(n17760), .C2(n17423), .A(n17422), .ZN(P3_U2807) );
  OAI22_X1 U20569 ( .A1(n17428), .A2(n17668), .B1(n17425), .B2(n18554), .ZN(
        n17426) );
  NOR2_X1 U20570 ( .A1(n17680), .A2(n17426), .ZN(n17452) );
  OAI21_X1 U20571 ( .B1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n17427), .A(
        n17452), .ZN(n17444) );
  NAND2_X1 U20572 ( .A1(n17428), .A2(n17544), .ZN(n17442) );
  AOI221_X1 U20573 ( .B1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .C1(n17430), .C2(n17429), .A(
        n17442), .ZN(n17433) );
  NAND2_X1 U20574 ( .A1(n17971), .A2(P3_REIP_REG_22__SCAN_IN), .ZN(n17781) );
  OAI21_X1 U20575 ( .B1(n17518), .B2(n10010), .A(n17781), .ZN(n17432) );
  AOI211_X1 U20576 ( .C1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .C2(n17444), .A(
        n17433), .B(n17432), .ZN(n17439) );
  OAI22_X1 U20577 ( .A1(n17710), .A2(n17847), .B1(n17616), .B2(n17846), .ZN(
        n17477) );
  INV_X1 U20578 ( .A(n17477), .ZN(n17515) );
  OAI21_X1 U20579 ( .B1(n17772), .B2(n17459), .A(n17515), .ZN(n17448) );
  AOI221_X1 U20580 ( .B1(n17766), .B2(n17435), .C1(n17445), .C2(n17435), .A(
        n17434), .ZN(n17437) );
  XNOR2_X1 U20581 ( .A(n17437), .B(n17436), .ZN(n17780) );
  AOI22_X1 U20582 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n17448), .B1(
        n17605), .B2(n17780), .ZN(n17438) );
  OAI211_X1 U20583 ( .C1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .C2(n17440), .A(
        n17439), .B(n17438), .ZN(P3_U2808) );
  NAND2_X1 U20584 ( .A1(n17791), .A2(n17774), .ZN(n17796) );
  INV_X1 U20585 ( .A(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n17828) );
  NOR2_X1 U20586 ( .A1(n17485), .A2(n17828), .ZN(n17787) );
  NAND2_X1 U20587 ( .A1(n17499), .A2(n17787), .ZN(n17476) );
  NOR2_X1 U20588 ( .A1(n18013), .A2(n18611), .ZN(n17785) );
  OAI22_X1 U20589 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n17442), .B1(
        n17441), .B2(n17518), .ZN(n17443) );
  AOI211_X1 U20590 ( .C1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .C2(n17444), .A(
        n17785), .B(n17443), .ZN(n17450) );
  NOR3_X1 U20591 ( .A1(n17828), .A2(n17615), .A3(n17445), .ZN(n17471) );
  AOI22_X1 U20592 ( .A1(n17791), .A2(n17471), .B1(n17484), .B2(n17446), .ZN(
        n17447) );
  XNOR2_X1 U20593 ( .A(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .B(n17447), .ZN(
        n17786) );
  AOI22_X1 U20594 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n17448), .B1(
        n17605), .B2(n17786), .ZN(n17449) );
  OAI211_X1 U20595 ( .C1(n17796), .C2(n17476), .A(n17450), .B(n17449), .ZN(
        P3_U2809) );
  NAND2_X1 U20596 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n17451), .ZN(
        n17805) );
  NAND2_X1 U20597 ( .A1(n17971), .A2(P3_REIP_REG_20__SCAN_IN), .ZN(n17803) );
  INV_X1 U20598 ( .A(n17803), .ZN(n17456) );
  AOI221_X1 U20599 ( .B1(n17454), .B2(n17453), .C1(n18078), .C2(n17453), .A(
        n17452), .ZN(n17455) );
  AOI211_X1 U20600 ( .C1(n17458), .C2(n17457), .A(n17456), .B(n17455), .ZN(
        n17462) );
  INV_X1 U20601 ( .A(n17787), .ZN(n17767) );
  NOR2_X1 U20602 ( .A1(n17810), .A2(n17767), .ZN(n17798) );
  OAI21_X1 U20603 ( .B1(n17459), .B2(n17798), .A(n17515), .ZN(n17473) );
  OAI221_X1 U20604 ( .B1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n17482), 
        .C1(n17810), .C2(n17471), .A(n9635), .ZN(n17460) );
  XNOR2_X1 U20605 ( .A(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .B(n17460), .ZN(
        n17801) );
  AOI22_X1 U20606 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n17473), .B1(
        n17605), .B2(n17801), .ZN(n17461) );
  OAI211_X1 U20607 ( .C1(n17476), .C2(n17805), .A(n17462), .B(n17461), .ZN(
        P3_U2810) );
  AOI21_X1 U20608 ( .B1(n17464), .B2(n17463), .A(n17680), .ZN(n17488) );
  OAI21_X1 U20609 ( .B1(n17465), .B2(n18554), .A(n17488), .ZN(n17481) );
  NOR2_X1 U20610 ( .A1(n18013), .A2(n18607), .ZN(n17806) );
  NAND2_X1 U20611 ( .A1(n17466), .A2(n17544), .ZN(n17479) );
  OAI21_X1 U20612 ( .B1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A(n17467), .ZN(n17468) );
  OAI22_X1 U20613 ( .A1(n17518), .A2(n17469), .B1(n17479), .B2(n17468), .ZN(
        n17470) );
  AOI211_X1 U20614 ( .C1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .C2(n17481), .A(
        n17806), .B(n17470), .ZN(n17475) );
  AOI21_X1 U20615 ( .B1(n17482), .B2(n17484), .A(n17471), .ZN(n17472) );
  XNOR2_X1 U20616 ( .A(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B(n17472), .ZN(
        n17807) );
  AOI22_X1 U20617 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n17473), .B1(
        n17605), .B2(n17807), .ZN(n17474) );
  OAI211_X1 U20618 ( .C1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n17476), .A(
        n17475), .B(n17474), .ZN(P3_U2811) );
  AOI21_X1 U20619 ( .B1(n17499), .B2(n17485), .A(n17477), .ZN(n17498) );
  NOR2_X1 U20620 ( .A1(n18013), .A2(n18604), .ZN(n17824) );
  OAI22_X1 U20621 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n17479), .B1(
        n17478), .B2(n17518), .ZN(n17480) );
  AOI211_X1 U20622 ( .C1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .C2(n17481), .A(
        n17824), .B(n17480), .ZN(n17487) );
  AOI21_X1 U20623 ( .B1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n15213), .A(
        n17482), .ZN(n17483) );
  XOR2_X1 U20624 ( .A(n17484), .B(n17483), .Z(n17823) );
  NOR2_X1 U20625 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n17485), .ZN(
        n17822) );
  AOI22_X1 U20626 ( .A1(n17605), .A2(n17823), .B1(n17499), .B2(n17822), .ZN(
        n17486) );
  OAI211_X1 U20627 ( .C1(n17498), .C2(n17828), .A(n17487), .B(n17486), .ZN(
        P3_U2812) );
  AOI21_X1 U20628 ( .B1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n17499), .A(
        P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n17497) );
  AOI221_X1 U20629 ( .B1(n18078), .B2(n17490), .C1(n17489), .C2(n17490), .A(
        n17488), .ZN(n17495) );
  AOI21_X1 U20630 ( .B1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n17491), .A(
        n17492), .ZN(n17832) );
  OAI22_X1 U20631 ( .A1(n17832), .A2(n17617), .B1(n17704), .B2(n17493), .ZN(
        n17494) );
  AOI211_X1 U20632 ( .C1(P3_REIP_REG_17__SCAN_IN), .C2(n17971), .A(n17495), 
        .B(n17494), .ZN(n17496) );
  OAI21_X1 U20633 ( .B1(n17498), .B2(n17497), .A(n17496), .ZN(P3_U2813) );
  INV_X1 U20634 ( .A(n17499), .ZN(n17516) );
  NOR3_X1 U20635 ( .A1(n17500), .A2(n17615), .A3(n17948), .ZN(n17595) );
  AOI21_X1 U20636 ( .B1(n17833), .B2(n17595), .A(n17501), .ZN(n17502) );
  XNOR2_X1 U20637 ( .A(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B(n17502), .ZN(
        n17841) );
  OAI21_X1 U20638 ( .B1(n17668), .B2(n17503), .A(n17707), .ZN(n17504) );
  INV_X1 U20639 ( .A(n17504), .ZN(n17535) );
  OAI21_X1 U20640 ( .B1(n17505), .B2(n18554), .A(n17535), .ZN(n17520) );
  AOI22_X1 U20641 ( .A1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(n17520), .B1(
        n17565), .B2(n17506), .ZN(n17512) );
  NOR3_X1 U20642 ( .A1(n17509), .A2(n17508), .A3(n17507), .ZN(n17522) );
  NAND2_X1 U20643 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n17510) );
  OAI211_X1 U20644 ( .C1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A(n17522), .B(n17510), .ZN(n17511) );
  OAI211_X1 U20645 ( .C1(n18600), .C2(n18013), .A(n17512), .B(n17511), .ZN(
        n17513) );
  AOI21_X1 U20646 ( .B1(n17605), .B2(n17841), .A(n17513), .ZN(n17514) );
  OAI221_X1 U20647 ( .B1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n17516), 
        .C1(n17840), .C2(n17515), .A(n17514), .ZN(P3_U2814) );
  NAND2_X1 U20648 ( .A1(n17904), .A2(n17836), .ZN(n17531) );
  NAND2_X1 U20649 ( .A1(n17845), .A2(n17531), .ZN(n17851) );
  INV_X1 U20650 ( .A(n17851), .ZN(n17530) );
  OR2_X1 U20651 ( .A1(n17616), .A2(n17846), .ZN(n17529) );
  NAND2_X1 U20652 ( .A1(n17971), .A2(P3_REIP_REG_15__SCAN_IN), .ZN(n17855) );
  OAI21_X1 U20653 ( .B1(n17518), .B2(n17517), .A(n17855), .ZN(n17519) );
  AOI221_X1 U20654 ( .B1(n17522), .B2(n17521), .C1(n17520), .C2(
        P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A(n17519), .ZN(n17528) );
  NAND2_X1 U20655 ( .A1(n17894), .A2(n17867), .ZN(n17523) );
  NAND2_X1 U20656 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n15213), .ZN(
        n17557) );
  AOI22_X1 U20657 ( .A1(n17524), .A2(n17537), .B1(n17523), .B2(n17557), .ZN(
        n17525) );
  XNOR2_X1 U20658 ( .A(n17525), .B(n17845), .ZN(n17854) );
  NOR2_X1 U20659 ( .A1(n17847), .A2(n17710), .ZN(n17526) );
  NAND2_X1 U20660 ( .A1(n17539), .A2(n17845), .ZN(n17849) );
  AOI22_X1 U20661 ( .A1(n17605), .A2(n17854), .B1(n17526), .B2(n17849), .ZN(
        n17527) );
  OAI211_X1 U20662 ( .C1(n17530), .C2(n17529), .A(n17528), .B(n17527), .ZN(
        P3_U2815) );
  INV_X1 U20663 ( .A(n17536), .ZN(n17858) );
  OAI221_X1 U20664 ( .B1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n17904), 
        .C1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .C2(n17858), .A(n17531), .ZN(
        n17868) );
  NAND3_X1 U20665 ( .A1(n18426), .A2(n17636), .A3(
        P3_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n17597) );
  NOR2_X1 U20666 ( .A1(n17532), .A2(n17597), .ZN(n17593) );
  AND2_X1 U20667 ( .A1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .A2(n17593), .ZN(
        n17579) );
  AOI21_X1 U20668 ( .B1(n17545), .B2(n17579), .A(
        P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n17534) );
  OAI22_X1 U20669 ( .A1(n17535), .A2(n17534), .B1(n17704), .B2(n17533), .ZN(
        n17541) );
  INV_X1 U20670 ( .A(n17595), .ZN(n17575) );
  OAI22_X1 U20671 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n17537), .B1(
        n17575), .B2(n17536), .ZN(n17538) );
  XNOR2_X1 U20672 ( .A(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B(n17538), .ZN(
        n17869) );
  OAI221_X1 U20673 ( .B1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .C1(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .C2(n17887), .A(n17539), .ZN(
        n17873) );
  OAI22_X1 U20674 ( .A1(n17869), .A2(n17617), .B1(n17710), .B2(n17873), .ZN(
        n17540) );
  AOI211_X1 U20675 ( .C1(n17971), .C2(P3_REIP_REG_14__SCAN_IN), .A(n17541), 
        .B(n17540), .ZN(n17542) );
  OAI21_X1 U20676 ( .B1(n17616), .B2(n17868), .A(n17542), .ZN(P3_U2816) );
  NAND2_X1 U20677 ( .A1(n17554), .A2(n17543), .ZN(n17893) );
  NAND2_X1 U20678 ( .A1(n17546), .A2(n17544), .ZN(n17569) );
  AOI211_X1 U20679 ( .C1(n17568), .C2(n17550), .A(n17545), .B(n17569), .ZN(
        n17552) );
  OAI21_X1 U20680 ( .B1(n17546), .B2(n17668), .A(n17707), .ZN(n17547) );
  AOI21_X1 U20681 ( .B1(n17549), .B2(n17548), .A(n17547), .ZN(n17567) );
  OAI22_X1 U20682 ( .A1(n17567), .A2(n17550), .B1(n18028), .B2(n18594), .ZN(
        n17551) );
  AOI211_X1 U20683 ( .C1(n17565), .C2(n17553), .A(n17552), .B(n17551), .ZN(
        n17562) );
  NAND2_X1 U20684 ( .A1(n17554), .A2(n17904), .ZN(n17883) );
  INV_X1 U20685 ( .A(n17883), .ZN(n17555) );
  OAI22_X1 U20686 ( .A1(n17887), .A2(n17710), .B1(n17555), .B2(n17616), .ZN(
        n17571) );
  INV_X1 U20687 ( .A(n17557), .ZN(n17558) );
  OAI22_X1 U20688 ( .A1(n17559), .A2(n17894), .B1(n17556), .B2(n17558), .ZN(
        n17560) );
  XNOR2_X1 U20689 ( .A(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .B(n17560), .ZN(
        n17878) );
  AOI22_X1 U20690 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n17571), .B1(
        n17605), .B2(n17878), .ZN(n17561) );
  OAI211_X1 U20691 ( .C1(n17608), .C2(n17893), .A(n17562), .B(n17561), .ZN(
        P3_U2817) );
  AOI21_X1 U20692 ( .B1(n17595), .B2(n17882), .A(n17556), .ZN(n17563) );
  XNOR2_X1 U20693 ( .A(n17563), .B(n17894), .ZN(n17901) );
  NOR2_X1 U20694 ( .A1(n17608), .A2(n17895), .ZN(n17572) );
  AOI22_X1 U20695 ( .A1(n17971), .A2(P3_REIP_REG_12__SCAN_IN), .B1(n17565), 
        .B2(n17564), .ZN(n17566) );
  OAI221_X1 U20696 ( .B1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n17569), .C1(
        n17568), .C2(n17567), .A(n17566), .ZN(n17570) );
  AOI221_X1 U20697 ( .B1(n17572), .B2(n17894), .C1(n17571), .C2(
        P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A(n17570), .ZN(n17573) );
  OAI21_X1 U20698 ( .B1(n17901), .B2(n17617), .A(n17573), .ZN(P3_U2818) );
  NAND2_X1 U20699 ( .A1(n17910), .A2(n9990), .ZN(n17917) );
  INV_X1 U20700 ( .A(n17910), .ZN(n17880) );
  OAI21_X1 U20701 ( .B1(n17880), .B2(n17575), .A(n17574), .ZN(n17576) );
  XNOR2_X1 U20702 ( .A(n17576), .B(n9990), .ZN(n17915) );
  NOR2_X1 U20703 ( .A1(n18013), .A2(n18590), .ZN(n17914) );
  AOI21_X1 U20704 ( .B1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n17700), .A(
        n17593), .ZN(n17578) );
  OAI22_X1 U20705 ( .A1(n17579), .A2(n17578), .B1(n17704), .B2(n17577), .ZN(
        n17580) );
  AOI211_X1 U20706 ( .C1(n17605), .C2(n17915), .A(n17914), .B(n17580), .ZN(
        n17582) );
  NOR2_X1 U20707 ( .A1(n17910), .A2(n17608), .ZN(n17584) );
  OAI22_X1 U20708 ( .A1(n17904), .A2(n17616), .B1(n17710), .B2(n17902), .ZN(
        n17594) );
  OAI21_X1 U20709 ( .B1(n17584), .B2(n17594), .A(
        P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n17581) );
  OAI211_X1 U20710 ( .C1(n17608), .C2(n17917), .A(n17582), .B(n17581), .ZN(
        P3_U2819) );
  INV_X1 U20711 ( .A(n17597), .ZN(n17625) );
  AOI22_X1 U20712 ( .A1(n17583), .A2(n17625), .B1(
        P3_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n17700), .ZN(n17592) );
  AOI21_X1 U20713 ( .B1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n17594), .A(
        n17584), .ZN(n17587) );
  AOI22_X1 U20714 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n17595), .B1(
        n17585), .B2(n17936), .ZN(n17586) );
  XNOR2_X1 U20715 ( .A(n17586), .B(n17922), .ZN(n17926) );
  OAI22_X1 U20716 ( .A1(n17588), .A2(n17587), .B1(n17926), .B2(n17617), .ZN(
        n17589) );
  AOI21_X1 U20717 ( .B1(n17590), .B2(n17457), .A(n17589), .ZN(n17591) );
  NAND2_X1 U20718 ( .A1(n17971), .A2(P3_REIP_REG_10__SCAN_IN), .ZN(n17924) );
  OAI211_X1 U20719 ( .C1(n17593), .C2(n17592), .A(n17591), .B(n17924), .ZN(
        P3_U2820) );
  INV_X1 U20720 ( .A(n17594), .ZN(n17607) );
  NOR2_X1 U20721 ( .A1(n17595), .A2(n17585), .ZN(n17596) );
  XNOR2_X1 U20722 ( .A(n17596), .B(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n17932) );
  NOR2_X1 U20723 ( .A1(n18013), .A2(n18586), .ZN(n17604) );
  NOR2_X1 U20724 ( .A1(n17598), .A2(n17597), .ZN(n17602) );
  AOI22_X1 U20725 ( .A1(n17599), .A2(n17625), .B1(
        P3_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n17700), .ZN(n17601) );
  OAI22_X1 U20726 ( .A1(n17602), .A2(n17601), .B1(n17704), .B2(n17600), .ZN(
        n17603) );
  AOI211_X1 U20727 ( .C1(n17605), .C2(n17932), .A(n17604), .B(n17603), .ZN(
        n17606) );
  OAI221_X1 U20728 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n17608), .C1(
        n17936), .C2(n17607), .A(n17606), .ZN(P3_U2821) );
  INV_X1 U20729 ( .A(n17609), .ZN(n17610) );
  OAI21_X1 U20730 ( .B1(n17610), .B2(n17668), .A(n17707), .ZN(n17626) );
  AOI22_X1 U20731 ( .A1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n17626), .B1(
        n17611), .B2(n17457), .ZN(n17623) );
  AOI21_X1 U20732 ( .B1(n17613), .B2(n17948), .A(n17612), .ZN(n17943) );
  AOI21_X1 U20733 ( .B1(n17615), .B2(n17939), .A(n17614), .ZN(n17941) );
  OAI22_X1 U20734 ( .A1(n17941), .A2(n17617), .B1(n17616), .B2(n17939), .ZN(
        n17618) );
  AOI21_X1 U20735 ( .B1(n17697), .B2(n17943), .A(n17618), .ZN(n17622) );
  NAND2_X1 U20736 ( .A1(n17971), .A2(P3_REIP_REG_8__SCAN_IN), .ZN(n17951) );
  OAI211_X1 U20737 ( .C1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .C2(n17620), .A(
        n18426), .B(n17619), .ZN(n17621) );
  NAND4_X1 U20738 ( .A1(n17623), .A2(n17622), .A3(n17951), .A4(n17621), .ZN(
        P3_U2822) );
  NOR2_X1 U20739 ( .A1(n18013), .A2(n18582), .ZN(n17956) );
  AOI221_X1 U20740 ( .B1(n17626), .B2(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .C1(
        n17625), .C2(n17624), .A(n17956), .ZN(n17634) );
  NAND2_X1 U20741 ( .A1(n17628), .A2(n17627), .ZN(n17629) );
  XNOR2_X1 U20742 ( .A(n17629), .B(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n17957) );
  AOI21_X1 U20743 ( .B1(n17632), .B2(n17630), .A(n17631), .ZN(n17958) );
  AOI22_X1 U20744 ( .A1(n17697), .A2(n17957), .B1(n9648), .B2(n17958), .ZN(
        n17633) );
  OAI211_X1 U20745 ( .C1(n17704), .C2(n17635), .A(n17634), .B(n17633), .ZN(
        P3_U2823) );
  NAND2_X1 U20746 ( .A1(n18426), .A2(n17636), .ZN(n17639) );
  NAND2_X1 U20747 ( .A1(n17700), .A2(n17639), .ZN(n17657) );
  AOI21_X1 U20748 ( .B1(n20912), .B2(n17638), .A(n17637), .ZN(n17965) );
  OAI22_X1 U20749 ( .A1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n17639), .B1(
        n18013), .B2(n18580), .ZN(n17640) );
  AOI21_X1 U20750 ( .B1(n17697), .B2(n17965), .A(n17640), .ZN(n17646) );
  AOI21_X1 U20751 ( .B1(n17643), .B2(n17642), .A(n17641), .ZN(n17966) );
  AOI22_X1 U20752 ( .A1(n9648), .A2(n17966), .B1(n17644), .B2(n17457), .ZN(
        n17645) );
  OAI211_X1 U20753 ( .C1(n17647), .C2(n17657), .A(n17646), .B(n17645), .ZN(
        P3_U2824) );
  AOI21_X1 U20754 ( .B1(n17648), .B2(n17707), .A(
        P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n17658) );
  AOI21_X1 U20755 ( .B1(n17969), .B2(n17650), .A(n17649), .ZN(n17972) );
  AOI22_X1 U20756 ( .A1(n9648), .A2(n17972), .B1(n17971), .B2(
        P3_REIP_REG_5__SCAN_IN), .ZN(n17656) );
  AOI21_X1 U20757 ( .B1(n17653), .B2(n17652), .A(n17651), .ZN(n17970) );
  AOI22_X1 U20758 ( .A1(n17697), .A2(n17970), .B1(n17654), .B2(n17457), .ZN(
        n17655) );
  OAI211_X1 U20759 ( .C1(n17658), .C2(n17657), .A(n17656), .B(n17655), .ZN(
        P3_U2825) );
  OAI21_X1 U20760 ( .B1(n17661), .B2(n17660), .A(n17659), .ZN(n17662) );
  XNOR2_X1 U20761 ( .A(n17662), .B(n17980), .ZN(n17987) );
  OAI22_X1 U20762 ( .A1(n17710), .A2(n17987), .B1(n18078), .B2(n17663), .ZN(
        n17664) );
  AOI21_X1 U20763 ( .B1(n17971), .B2(P3_REIP_REG_4__SCAN_IN), .A(n17664), .ZN(
        n17671) );
  AOI21_X1 U20764 ( .B1(n17667), .B2(n17666), .A(n17665), .ZN(n17985) );
  OAI21_X1 U20765 ( .B1(n17669), .B2(n17668), .A(n17707), .ZN(n17682) );
  AOI22_X1 U20766 ( .A1(n9648), .A2(n17985), .B1(
        P3_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n17682), .ZN(n17670) );
  OAI211_X1 U20767 ( .C1(n17704), .C2(n17672), .A(n17671), .B(n17670), .ZN(
        P3_U2826) );
  AOI21_X1 U20768 ( .B1(n17675), .B2(n17674), .A(n17673), .ZN(n17989) );
  AOI22_X1 U20769 ( .A1(n17697), .A2(n17989), .B1(n17971), .B2(
        P3_REIP_REG_3__SCAN_IN), .ZN(n17684) );
  AOI21_X1 U20770 ( .B1(n17678), .B2(n17677), .A(n17676), .ZN(n17988) );
  OAI21_X1 U20771 ( .B1(n17680), .B2(n17694), .A(n17679), .ZN(n17681) );
  AOI22_X1 U20772 ( .A1(n9648), .A2(n17988), .B1(n17682), .B2(n17681), .ZN(
        n17683) );
  OAI211_X1 U20773 ( .C1(n17704), .C2(n17685), .A(n17684), .B(n17683), .ZN(
        P3_U2827) );
  AOI21_X1 U20774 ( .B1(n17688), .B2(n17687), .A(n17686), .ZN(n17998) );
  INV_X1 U20775 ( .A(P3_REIP_REG_2__SCAN_IN), .ZN(n18572) );
  NOR2_X1 U20776 ( .A1(n18013), .A2(n18572), .ZN(n17997) );
  XNOR2_X1 U20777 ( .A(n17690), .B(n17689), .ZN(n17995) );
  OAI22_X1 U20778 ( .A1(n17704), .A2(n17691), .B1(n9647), .B2(n17995), .ZN(
        n17692) );
  AOI211_X1 U20779 ( .C1(n17697), .C2(n17998), .A(n17997), .B(n17692), .ZN(
        n17693) );
  OAI221_X1 U20780 ( .B1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n18078), .C1(
        n17694), .C2(n17707), .A(n17693), .ZN(P3_U2828) );
  NOR2_X1 U20781 ( .A1(n17706), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n17695) );
  XOR2_X1 U20782 ( .A(n17699), .B(n17695), .Z(n18024) );
  INV_X1 U20783 ( .A(n18024), .ZN(n17696) );
  AOI22_X1 U20784 ( .A1(n17697), .A2(n17696), .B1(n17971), .B2(
        P3_REIP_REG_1__SCAN_IN), .ZN(n17703) );
  AOI21_X1 U20785 ( .B1(n17699), .B2(n17705), .A(n17698), .ZN(n18018) );
  AOI22_X1 U20786 ( .A1(n9648), .A2(n18018), .B1(
        P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n17700), .ZN(n17702) );
  OAI211_X1 U20787 ( .C1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .C2(n17704), .A(
        n17703), .B(n17702), .ZN(P3_U2829) );
  OAI21_X1 U20788 ( .B1(n17706), .B2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n17705), .ZN(n18032) );
  INV_X1 U20789 ( .A(n18032), .ZN(n18034) );
  NAND3_X1 U20790 ( .A1(n18650), .A2(n18554), .A3(n17707), .ZN(n17708) );
  AOI22_X1 U20791 ( .A1(n17971), .A2(P3_REIP_REG_0__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n17708), .ZN(n17709) );
  OAI221_X1 U20792 ( .B1(n18034), .B2(n17710), .C1(n18032), .C2(n9647), .A(
        n17709), .ZN(P3_U2830) );
  AOI221_X1 U20793 ( .B1(n17712), .B2(n17711), .C1(n17761), .C2(n17711), .A(
        n18019), .ZN(n17722) );
  NOR2_X1 U20794 ( .A1(n18499), .A2(n18510), .ZN(n18006) );
  AOI21_X1 U20795 ( .B1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n17929), .A(
        n17713), .ZN(n17773) );
  INV_X1 U20796 ( .A(n18006), .ZN(n17819) );
  OAI21_X1 U20797 ( .B1(n17773), .B2(n17714), .A(n17819), .ZN(n17752) );
  OAI21_X1 U20798 ( .B1(n17737), .B2(n18006), .A(n17752), .ZN(n17734) );
  AOI22_X1 U20799 ( .A1(n18499), .A2(n17738), .B1(n18510), .B2(n17715), .ZN(
        n17717) );
  OAI211_X1 U20800 ( .C1(n17718), .C2(n18486), .A(n17717), .B(n17716), .ZN(
        n17719) );
  OAI211_X1 U20801 ( .C1(n18512), .C2(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        P3_INSTADDRPOINTER_REG_27__SCAN_IN), .B(n17728), .ZN(n17721) );
  AOI22_X1 U20802 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n18021), .B1(
        n17722), .B2(n17721), .ZN(n17724) );
  NAND2_X1 U20803 ( .A1(n17971), .A2(P3_REIP_REG_27__SCAN_IN), .ZN(n17723) );
  OAI211_X1 U20804 ( .C1(n17725), .C2(n17940), .A(n17724), .B(n17723), .ZN(
        P3_U2835) );
  AND2_X1 U20805 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(n17726), .ZN(
        n17749) );
  INV_X1 U20806 ( .A(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n17727) );
  AOI211_X1 U20807 ( .C1(n18025), .C2(n17728), .A(n17971), .B(n17727), .ZN(
        n17730) );
  AOI211_X1 U20808 ( .C1(n17731), .C2(n17749), .A(n17730), .B(n17729), .ZN(
        n17732) );
  OAI21_X1 U20809 ( .B1(n17733), .B2(n17940), .A(n17732), .ZN(P3_U2836) );
  INV_X1 U20810 ( .A(n17737), .ZN(n17735) );
  AOI221_X1 U20811 ( .B1(n17754), .B2(n18003), .C1(n17735), .C2(n18003), .A(
        n17734), .ZN(n17740) );
  NAND2_X1 U20812 ( .A1(n17737), .A2(n17736), .ZN(n17739) );
  AOI221_X1 U20813 ( .B1(n17740), .B2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), 
        .C1(n17739), .C2(n17738), .A(n18019), .ZN(n17741) );
  AOI211_X1 U20814 ( .C1(n18021), .C2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n17742), .B(n17741), .ZN(n17746) );
  AOI22_X1 U20815 ( .A1(n17877), .A2(n17744), .B1(n17999), .B2(n17743), .ZN(
        n17745) );
  OAI211_X1 U20816 ( .C1(n17940), .C2(n17747), .A(n17746), .B(n17745), .ZN(
        P3_U2837) );
  AOI22_X1 U20817 ( .A1(P3_REIP_REG_24__SCAN_IN), .A2(n17971), .B1(n17749), 
        .B2(n17748), .ZN(n17758) );
  INV_X1 U20818 ( .A(n17947), .ZN(n17837) );
  AOI22_X1 U20819 ( .A1(n17771), .A2(n17751), .B1(n17884), .B2(n17750), .ZN(
        n17753) );
  NAND3_X1 U20820 ( .A1(n17753), .A2(n18012), .A3(n17752), .ZN(n17756) );
  AOI211_X1 U20821 ( .C1(n18003), .C2(n17754), .A(n17760), .B(n17756), .ZN(
        n17755) );
  NOR2_X1 U20822 ( .A1(n17971), .A2(n17755), .ZN(n17763) );
  OAI211_X1 U20823 ( .C1(n17837), .C2(n17756), .A(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .B(n17763), .ZN(n17757) );
  OAI211_X1 U20824 ( .C1(n17759), .C2(n17940), .A(n17758), .B(n17757), .ZN(
        P3_U2838) );
  OAI21_X1 U20825 ( .B1(n18021), .B2(n17761), .A(n17760), .ZN(n17762) );
  AOI22_X1 U20826 ( .A1(n17933), .A2(n17764), .B1(n17763), .B2(n17762), .ZN(
        n17765) );
  OAI21_X1 U20827 ( .B1(n18028), .B2(n18615), .A(n17765), .ZN(P3_U2839) );
  INV_X1 U20828 ( .A(n17766), .ZN(n17779) );
  INV_X1 U20829 ( .A(n17884), .ZN(n17903) );
  OAI22_X1 U20830 ( .A1(n18486), .A2(n17847), .B1(n17903), .B2(n17846), .ZN(
        n17788) );
  INV_X1 U20831 ( .A(n17788), .ZN(n17777) );
  INV_X1 U20832 ( .A(n17791), .ZN(n17770) );
  OAI21_X1 U20833 ( .B1(n17768), .B2(n17767), .A(n18003), .ZN(n17769) );
  OAI221_X1 U20834 ( .B1(n18512), .B2(n17813), .C1(n18512), .C2(n17798), .A(
        n17769), .ZN(n17789) );
  AOI21_X1 U20835 ( .B1(n18003), .B2(n17770), .A(n17789), .ZN(n17776) );
  NOR2_X1 U20836 ( .A1(n17771), .A2(n17884), .ZN(n17909) );
  OAI22_X1 U20837 ( .A1(n18512), .A2(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .B1(
        n17772), .B2(n17909), .ZN(n17793) );
  AOI211_X1 U20838 ( .C1(n17919), .C2(n17774), .A(n17773), .B(n17793), .ZN(
        n17775) );
  NAND3_X1 U20839 ( .A1(n17777), .A2(n17776), .A3(n17775), .ZN(n17778) );
  OAI221_X1 U20840 ( .B1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n17779), 
        .C1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .C2(n17784), .A(n17778), .ZN(
        n17783) );
  AOI22_X1 U20841 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n18021), .B1(
        n17933), .B2(n17780), .ZN(n17782) );
  OAI211_X1 U20842 ( .C1(n18019), .C2(n17783), .A(n17782), .B(n17781), .ZN(
        P3_U2840) );
  NAND3_X1 U20843 ( .A1(n18025), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A3(
        n17784), .ZN(n17811) );
  AOI21_X1 U20844 ( .B1(n17933), .B2(n17786), .A(n17785), .ZN(n17795) );
  NOR2_X1 U20845 ( .A1(n18003), .A2(n18510), .ZN(n18020) );
  NOR2_X1 U20846 ( .A1(n18665), .A2(n17879), .ZN(n17930) );
  NAND3_X1 U20847 ( .A1(n17833), .A2(n17787), .A3(n17930), .ZN(n17790) );
  NOR2_X1 U20848 ( .A1(n18019), .A2(n17788), .ZN(n17817) );
  INV_X1 U20849 ( .A(n17817), .ZN(n17838) );
  AOI211_X1 U20850 ( .C1(n18510), .C2(n17790), .A(n17838), .B(n17789), .ZN(
        n17797) );
  OAI21_X1 U20851 ( .B1(n17791), .B2(n18020), .A(n17797), .ZN(n17792) );
  OAI211_X1 U20852 ( .C1(n17793), .C2(n17792), .A(
        P3_INSTADDRPOINTER_REG_21__SCAN_IN), .B(n18028), .ZN(n17794) );
  OAI211_X1 U20853 ( .C1(n17796), .C2(n17811), .A(n17795), .B(n17794), .ZN(
        P3_U2841) );
  NAND2_X1 U20854 ( .A1(n17810), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n17800) );
  OAI21_X1 U20855 ( .B1(n17798), .B2(n17909), .A(n17797), .ZN(n17799) );
  NAND2_X1 U20856 ( .A1(n17799), .A2(n18028), .ZN(n17809) );
  OAI21_X1 U20857 ( .B1(n18020), .B2(n17800), .A(n17809), .ZN(n17802) );
  AOI22_X1 U20858 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n17802), .B1(
        n17933), .B2(n17801), .ZN(n17804) );
  OAI211_X1 U20859 ( .C1(n17811), .C2(n17805), .A(n17804), .B(n17803), .ZN(
        P3_U2842) );
  AOI21_X1 U20860 ( .B1(n17933), .B2(n17807), .A(n17806), .ZN(n17808) );
  OAI221_X1 U20861 ( .B1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n17811), 
        .C1(n17810), .C2(n17809), .A(n17808), .ZN(P3_U2843) );
  INV_X1 U20862 ( .A(n17812), .ZN(n17815) );
  OAI211_X1 U20863 ( .C1(n17929), .C2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B(n17813), .ZN(n17814) );
  AOI22_X1 U20864 ( .A1(n18003), .A2(n17815), .B1(n17819), .B2(n17814), .ZN(
        n17816) );
  OAI211_X1 U20865 ( .C1(n17818), .C2(n17909), .A(n17817), .B(n17816), .ZN(
        n17829) );
  OAI221_X1 U20866 ( .B1(n17829), .B2(n9980), .C1(n17829), .C2(n17819), .A(
        n18028), .ZN(n17827) );
  OAI22_X1 U20867 ( .A1(n18000), .A2(n18509), .B1(n17977), .B2(n18002), .ZN(
        n17991) );
  NAND3_X1 U20868 ( .A1(n18025), .A2(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A3(
        n17991), .ZN(n17981) );
  NOR3_X1 U20869 ( .A1(n17969), .A2(n17980), .A3(n17981), .ZN(n17964) );
  NAND2_X1 U20870 ( .A1(n17844), .A2(n17964), .ZN(n17874) );
  OAI22_X1 U20871 ( .A1(n17821), .A2(n18019), .B1(n17820), .B2(n17874), .ZN(
        n17839) );
  AOI22_X1 U20872 ( .A1(n17933), .A2(n17823), .B1(n17822), .B2(n17839), .ZN(
        n17826) );
  INV_X1 U20873 ( .A(n17824), .ZN(n17825) );
  OAI211_X1 U20874 ( .C1(n17828), .C2(n17827), .A(n17826), .B(n17825), .ZN(
        P3_U2844) );
  OAI221_X1 U20875 ( .B1(P3_REIP_REG_17__SCAN_IN), .B2(n18013), .C1(
        P3_INSTADDRPOINTER_REG_17__SCAN_IN), .C2(n17971), .A(n17829), .ZN(
        n17831) );
  NAND3_X1 U20876 ( .A1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n9980), .A3(
        n17839), .ZN(n17830) );
  OAI211_X1 U20877 ( .C1(n17832), .C2(n17940), .A(n17831), .B(n17830), .ZN(
        P3_U2845) );
  INV_X1 U20878 ( .A(n17919), .ZN(n17889) );
  NAND2_X1 U20879 ( .A1(n17833), .A2(n17930), .ZN(n17834) );
  NOR2_X1 U20880 ( .A1(n17859), .A2(n18509), .ZN(n17906) );
  AOI211_X1 U20881 ( .C1(n17834), .C2(n18510), .A(n17845), .B(n17906), .ZN(
        n17835) );
  NAND2_X1 U20882 ( .A1(n18499), .A2(n17879), .ZN(n17928) );
  OAI211_X1 U20883 ( .C1(n17889), .C2(n17836), .A(n17835), .B(n17928), .ZN(
        n17852) );
  OAI221_X1 U20884 ( .B1(n17838), .B2(n17837), .C1(n17838), .C2(n17852), .A(
        P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n17843) );
  AOI22_X1 U20885 ( .A1(n17933), .A2(n17841), .B1(n17840), .B2(n17839), .ZN(
        n17842) );
  OAI221_X1 U20886 ( .B1(n17971), .B2(n17843), .C1(n18013), .C2(n18600), .A(
        n17842), .ZN(P3_U2846) );
  INV_X1 U20887 ( .A(n17946), .ZN(n17953) );
  NAND4_X1 U20888 ( .A1(n17953), .A2(n17858), .A3(n17844), .A4(n17991), .ZN(
        n17865) );
  OAI21_X1 U20889 ( .B1(n17867), .B2(n17865), .A(n17845), .ZN(n17853) );
  NOR2_X1 U20890 ( .A1(n17846), .A2(n17903), .ZN(n17850) );
  NOR2_X1 U20891 ( .A1(n17847), .A2(n18486), .ZN(n17848) );
  AOI222_X1 U20892 ( .A1(n17853), .A2(n17852), .B1(n17851), .B2(n17850), .C1(
        n17849), .C2(n17848), .ZN(n17857) );
  AOI22_X1 U20893 ( .A1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n18021), .B1(
        n17933), .B2(n17854), .ZN(n17856) );
  OAI211_X1 U20894 ( .C1(n17857), .C2(n18019), .A(n17856), .B(n17855), .ZN(
        P3_U2847) );
  OAI22_X1 U20895 ( .A1(n18512), .A2(n17858), .B1(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n18020), .ZN(n17864) );
  INV_X1 U20896 ( .A(n17930), .ZN(n17907) );
  OAI21_X1 U20897 ( .B1(n17861), .B2(n17907), .A(n18510), .ZN(n17885) );
  INV_X1 U20898 ( .A(n17859), .ZN(n17860) );
  OAI21_X1 U20899 ( .B1(n17861), .B2(n17860), .A(n18003), .ZN(n17862) );
  NAND4_X1 U20900 ( .A1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n17885), .A3(
        n17928), .A4(n17862), .ZN(n17863) );
  OAI21_X1 U20901 ( .B1(n17864), .B2(n17863), .A(n18025), .ZN(n17866) );
  AOI222_X1 U20902 ( .A1(n17867), .A2(n17866), .B1(n17867), .B2(n17865), .C1(
        n17866), .C2(n18012), .ZN(n17871) );
  OAI22_X1 U20903 ( .A1(n17869), .A2(n17940), .B1(n17938), .B2(n17868), .ZN(
        n17870) );
  AOI211_X1 U20904 ( .C1(n17971), .C2(P3_REIP_REG_14__SCAN_IN), .A(n17871), 
        .B(n17870), .ZN(n17872) );
  OAI21_X1 U20905 ( .B1(n18033), .B2(n17873), .A(n17872), .ZN(P3_U2848) );
  OAI21_X1 U20906 ( .B1(n17875), .B2(n18033), .A(n17874), .ZN(n17876) );
  AOI21_X1 U20907 ( .B1(n17904), .B2(n17877), .A(n17876), .ZN(n17937) );
  AOI22_X1 U20908 ( .A1(n17971), .A2(P3_REIP_REG_13__SCAN_IN), .B1(n17933), 
        .B2(n17878), .ZN(n17892) );
  OAI21_X1 U20909 ( .B1(n17880), .B2(n17879), .A(n18499), .ZN(n17881) );
  OAI21_X1 U20910 ( .B1(n17882), .B2(n18509), .A(n17881), .ZN(n17911) );
  AOI211_X1 U20911 ( .C1(n17884), .C2(n17883), .A(n17906), .B(n17911), .ZN(
        n17886) );
  OAI211_X1 U20912 ( .C1(n17887), .C2(n18486), .A(n17886), .B(n17885), .ZN(
        n17897) );
  OAI21_X1 U20913 ( .B1(n18512), .B2(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A(
        P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n17898) );
  INV_X1 U20914 ( .A(n17898), .ZN(n17888) );
  OAI21_X1 U20915 ( .B1(n17889), .B2(n17888), .A(n18025), .ZN(n17890) );
  OAI211_X1 U20916 ( .C1(n17897), .C2(n17890), .A(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .B(n18028), .ZN(n17891) );
  OAI211_X1 U20917 ( .C1(n17937), .C2(n17893), .A(n17892), .B(n17891), .ZN(
        P3_U2849) );
  AOI22_X1 U20918 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n18021), .B1(
        n17971), .B2(P3_REIP_REG_12__SCAN_IN), .ZN(n17900) );
  OAI22_X1 U20919 ( .A1(n17937), .A2(n17895), .B1(n17894), .B2(n18019), .ZN(
        n17896) );
  OAI21_X1 U20920 ( .B1(n17898), .B2(n17897), .A(n17896), .ZN(n17899) );
  OAI211_X1 U20921 ( .C1(n17901), .C2(n17940), .A(n17900), .B(n17899), .ZN(
        P3_U2850) );
  OAI22_X1 U20922 ( .A1(n17904), .A2(n17903), .B1(n18486), .B2(n17902), .ZN(
        n17905) );
  NOR3_X1 U20923 ( .A1(n17906), .A2(n18019), .A3(n17905), .ZN(n17927) );
  OAI21_X1 U20924 ( .B1(n17936), .B2(n17907), .A(n18510), .ZN(n17908) );
  OAI211_X1 U20925 ( .C1(n17910), .C2(n17909), .A(n17927), .B(n17908), .ZN(
        n17918) );
  AOI211_X1 U20926 ( .C1(n18510), .C2(n17922), .A(n17911), .B(n17918), .ZN(
        n17912) );
  NOR3_X1 U20927 ( .A1(n17971), .A2(n17912), .A3(n9990), .ZN(n17913) );
  AOI211_X1 U20928 ( .C1(n17933), .C2(n17915), .A(n17914), .B(n17913), .ZN(
        n17916) );
  OAI21_X1 U20929 ( .B1(n17937), .B2(n17917), .A(n17916), .ZN(P3_U2851) );
  AOI21_X1 U20930 ( .B1(n17919), .B2(n17936), .A(n17918), .ZN(n17920) );
  AOI21_X1 U20931 ( .B1(n17920), .B2(n17928), .A(n17971), .ZN(n17923) );
  OAI21_X1 U20932 ( .B1(n17936), .B2(n17937), .A(n17922), .ZN(n17921) );
  OAI21_X1 U20933 ( .B1(n17923), .B2(n17922), .A(n17921), .ZN(n17925) );
  OAI211_X1 U20934 ( .C1(n17926), .C2(n17940), .A(n17925), .B(n17924), .ZN(
        P3_U2852) );
  OAI211_X1 U20935 ( .C1(n17930), .C2(n17929), .A(n17928), .B(n17927), .ZN(
        n17931) );
  NAND2_X1 U20936 ( .A1(n18013), .A2(n17931), .ZN(n17935) );
  AOI22_X1 U20937 ( .A1(n17971), .A2(P3_REIP_REG_9__SCAN_IN), .B1(n17933), 
        .B2(n17932), .ZN(n17934) );
  OAI221_X1 U20938 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n17937), .C1(
        n17936), .C2(n17935), .A(n17934), .ZN(P3_U2853) );
  OAI22_X1 U20939 ( .A1(n17941), .A2(n17940), .B1(n17939), .B2(n17938), .ZN(
        n17942) );
  AOI21_X1 U20940 ( .B1(n17999), .B2(n17943), .A(n17942), .ZN(n17952) );
  AOI22_X1 U20941 ( .A1(n18003), .A2(n18000), .B1(n18510), .B2(n18665), .ZN(
        n18005) );
  OAI21_X1 U20942 ( .B1(n17944), .B2(n18006), .A(n18005), .ZN(n17945) );
  AOI21_X1 U20943 ( .B1(n18003), .B2(n17946), .A(n17945), .ZN(n17962) );
  OAI211_X1 U20944 ( .C1(n17947), .C2(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A(
        P3_INSTADDRPOINTER_REG_7__SCAN_IN), .B(n17962), .ZN(n17954) );
  OAI221_X1 U20945 ( .B1(n18021), .B2(n17979), .C1(n18021), .C2(n17954), .A(
        P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n17950) );
  NAND4_X1 U20946 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A3(n17964), .A4(n17948), .ZN(
        n17949) );
  NAND4_X1 U20947 ( .A1(n17952), .A2(n17951), .A3(n17950), .A4(n17949), .ZN(
        P3_U2854) );
  AND2_X1 U20948 ( .A1(n17991), .A2(n17953), .ZN(n17955) );
  OAI221_X1 U20949 ( .B1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_6__SCAN_IN), .C1(
        P3_INSTADDRPOINTER_REG_7__SCAN_IN), .C2(n17955), .A(n17954), .ZN(
        n17961) );
  AOI21_X1 U20950 ( .B1(n18021), .B2(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A(
        n17956), .ZN(n17960) );
  INV_X1 U20951 ( .A(n18031), .ZN(n18017) );
  AOI22_X1 U20952 ( .A1(n18017), .A2(n17958), .B1(n17999), .B2(n17957), .ZN(
        n17959) );
  OAI211_X1 U20953 ( .C1(n18019), .C2(n17961), .A(n17960), .B(n17959), .ZN(
        P3_U2855) );
  OAI21_X1 U20954 ( .B1(n17962), .B2(n18019), .A(n18012), .ZN(n17973) );
  NOR2_X1 U20955 ( .A1(n18013), .A2(n18580), .ZN(n17963) );
  AOI221_X1 U20956 ( .B1(n17964), .B2(n20912), .C1(n17973), .C2(
        P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A(n17963), .ZN(n17968) );
  AOI22_X1 U20957 ( .A1(n18017), .A2(n17966), .B1(n17999), .B2(n17965), .ZN(
        n17967) );
  NAND2_X1 U20958 ( .A1(n17968), .A2(n17967), .ZN(P3_U2856) );
  NAND2_X1 U20959 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n17969), .ZN(
        n17976) );
  AOI22_X1 U20960 ( .A1(n17971), .A2(P3_REIP_REG_5__SCAN_IN), .B1(n17999), 
        .B2(n17970), .ZN(n17975) );
  AOI22_X1 U20961 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n17973), .B1(
        n18017), .B2(n17972), .ZN(n17974) );
  OAI211_X1 U20962 ( .C1(n17981), .C2(n17976), .A(n17975), .B(n17974), .ZN(
        P3_U2857) );
  NOR2_X1 U20963 ( .A1(n18013), .A2(n18576), .ZN(n17984) );
  INV_X1 U20964 ( .A(n17977), .ZN(n17978) );
  OAI211_X1 U20965 ( .C1(n17978), .C2(n18006), .A(
        P3_INSTADDRPOINTER_REG_3__SCAN_IN), .B(n18005), .ZN(n17990) );
  AOI21_X1 U20966 ( .B1(n17979), .B2(n17990), .A(n18021), .ZN(n17982) );
  AOI22_X1 U20967 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n17982), .B1(
        n17981), .B2(n17980), .ZN(n17983) );
  AOI211_X1 U20968 ( .C1(n17985), .C2(n18017), .A(n17984), .B(n17983), .ZN(
        n17986) );
  OAI21_X1 U20969 ( .B1(n18033), .B2(n17987), .A(n17986), .ZN(P3_U2858) );
  AOI22_X1 U20970 ( .A1(n17971), .A2(P3_REIP_REG_3__SCAN_IN), .B1(n18017), 
        .B2(n17988), .ZN(n17994) );
  AOI22_X1 U20971 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n18021), .B1(
        n17999), .B2(n17989), .ZN(n17993) );
  OAI211_X1 U20972 ( .C1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .C2(n17991), .A(
        n18025), .B(n17990), .ZN(n17992) );
  NAND3_X1 U20973 ( .A1(n17994), .A2(n17993), .A3(n17992), .ZN(P3_U2859) );
  NOR2_X1 U20974 ( .A1(n18031), .A2(n17995), .ZN(n17996) );
  AOI211_X1 U20975 ( .C1(n17999), .C2(n17998), .A(n17997), .B(n17996), .ZN(
        n18010) );
  NAND2_X1 U20976 ( .A1(n18003), .A2(n18000), .ZN(n18001) );
  OAI21_X1 U20977 ( .B1(n18002), .B2(n18652), .A(n18001), .ZN(n18008) );
  NAND3_X1 U20978 ( .A1(n18003), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n18004) );
  OAI211_X1 U20979 ( .C1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .C2(n18006), .A(
        n18005), .B(n18004), .ZN(n18007) );
  OAI221_X1 U20980 ( .B1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n18008), .C1(
        n18011), .C2(n18007), .A(n18025), .ZN(n18009) );
  OAI211_X1 U20981 ( .C1(n18012), .C2(n18011), .A(n18010), .B(n18009), .ZN(
        P3_U2860) );
  NOR2_X1 U20982 ( .A1(n18013), .A2(n18679), .ZN(n18016) );
  AOI211_X1 U20983 ( .C1(n18512), .C2(n18665), .A(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B(n18014), .ZN(n18015) );
  AOI211_X1 U20984 ( .C1(n18018), .C2(n18017), .A(n18016), .B(n18015), .ZN(
        n18023) );
  NOR3_X1 U20985 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n18020), .A3(
        n18019), .ZN(n18027) );
  OAI21_X1 U20986 ( .B1(n18021), .B2(n18027), .A(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n18022) );
  OAI211_X1 U20987 ( .C1(n18024), .C2(n18033), .A(n18023), .B(n18022), .ZN(
        P3_U2861) );
  AOI21_X1 U20988 ( .B1(n18512), .B2(n18025), .A(n18665), .ZN(n18026) );
  NOR2_X1 U20989 ( .A1(n18027), .A2(n18026), .ZN(n18029) );
  MUX2_X1 U20990 ( .A(n18672), .B(n18029), .S(n18028), .Z(n18030) );
  OAI221_X1 U20991 ( .B1(n18034), .B2(n18033), .C1(n18032), .C2(n18031), .A(
        n18030), .ZN(P3_U2862) );
  OAI21_X1 U20992 ( .B1(P3_FLUSH_REG_SCAN_IN), .B2(n18036), .A(n18035), .ZN(
        n18541) );
  OAI21_X1 U20993 ( .B1(n18037), .B2(n18039), .A(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n18038) );
  OAI221_X1 U20994 ( .B1(n18039), .B2(n18541), .C1(n18039), .C2(n18091), .A(
        n18038), .ZN(P3_U2863) );
  INV_X1 U20995 ( .A(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n18049) );
  NOR2_X1 U20996 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n18522), .ZN(
        n18224) );
  NOR2_X1 U20997 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n18049), .ZN(
        n18290) );
  NOR2_X1 U20998 ( .A1(n18224), .A2(n18290), .ZN(n18041) );
  OAI22_X1 U20999 ( .A1(n18042), .A2(n18049), .B1(n18041), .B2(n18040), .ZN(
        P3_U2866) );
  NOR2_X1 U21000 ( .A1(n18044), .A2(n18043), .ZN(P3_U2867) );
  NAND2_X1 U21001 ( .A1(n18046), .A2(n18045), .ZN(n18086) );
  NOR2_X1 U21002 ( .A1(n18047), .A2(n18086), .ZN(n18337) );
  INV_X1 U21003 ( .A(n18337), .ZN(n18430) );
  NAND2_X1 U21004 ( .A1(n18517), .A2(n18515), .ZN(n18518) );
  NOR2_X1 U21005 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n18110) );
  INV_X1 U21006 ( .A(n18110), .ZN(n18133) );
  NOR2_X2 U21007 ( .A1(n18518), .A2(n18133), .ZN(n18151) );
  INV_X1 U21008 ( .A(n18151), .ZN(n18131) );
  NAND2_X1 U21009 ( .A1(BUF2_REG_24__SCAN_IN), .A2(n18426), .ZN(n18340) );
  INV_X1 U21010 ( .A(n18340), .ZN(n18422) );
  NOR2_X1 U21011 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18515), .ZN(
        n18269) );
  NOR2_X1 U21012 ( .A1(n18522), .A2(n18049), .ZN(n18362) );
  NAND2_X1 U21013 ( .A1(n18269), .A2(n18362), .ZN(n18479) );
  INV_X1 U21014 ( .A(n18479), .ZN(n18464) );
  NOR2_X2 U21015 ( .A1(n18083), .A2(n18048), .ZN(n18421) );
  INV_X1 U21016 ( .A(n18544), .ZN(n18420) );
  NOR2_X1 U21017 ( .A1(n18049), .A2(n18198), .ZN(n18424) );
  INV_X1 U21018 ( .A(n18424), .ZN(n18419) );
  NOR2_X2 U21019 ( .A1(n18515), .A2(n18419), .ZN(n18474) );
  NOR2_X1 U21020 ( .A1(n18474), .A2(n18151), .ZN(n18111) );
  NOR2_X1 U21021 ( .A1(n18420), .A2(n18111), .ZN(n18085) );
  AOI22_X1 U21022 ( .A1(n18422), .A2(n18464), .B1(n18421), .B2(n18085), .ZN(
        n18054) );
  NAND2_X1 U21023 ( .A1(n18424), .A2(n18515), .ZN(n18410) );
  NAND2_X1 U21024 ( .A1(n18410), .A2(n18479), .ZN(n18383) );
  AOI21_X1 U21025 ( .B1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(
        P3_STATE2_REG_3__SCAN_IN), .A(n18083), .ZN(n18051) );
  INV_X1 U21026 ( .A(n18111), .ZN(n18050) );
  AOI22_X1 U21027 ( .A1(n18426), .A2(n18383), .B1(n18051), .B2(n18050), .ZN(
        n18088) );
  NOR2_X2 U21028 ( .A1(n18078), .A2(n18052), .ZN(n18427) );
  INV_X1 U21029 ( .A(n18410), .ZN(n18413) );
  AOI22_X1 U21030 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n18088), .B1(
        n18427), .B2(n18413), .ZN(n18053) );
  OAI211_X1 U21031 ( .C1(n18430), .C2(n18131), .A(n18054), .B(n18053), .ZN(
        P3_U2868) );
  NOR2_X1 U21032 ( .A1(n18692), .A2(n18086), .ZN(n18433) );
  INV_X1 U21033 ( .A(n18433), .ZN(n18394) );
  NAND2_X1 U21034 ( .A1(BUF2_REG_25__SCAN_IN), .A2(n18426), .ZN(n18437) );
  INV_X1 U21035 ( .A(n18437), .ZN(n18391) );
  NOR2_X2 U21036 ( .A1(n18083), .A2(n18055), .ZN(n18432) );
  AOI22_X1 U21037 ( .A1(n18391), .A2(n18464), .B1(n18432), .B2(n18085), .ZN(
        n18057) );
  NOR2_X2 U21038 ( .A1(n18078), .A2(n19151), .ZN(n18431) );
  AOI22_X1 U21039 ( .A1(P3_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n18088), .B1(
        n18431), .B2(n18413), .ZN(n18056) );
  OAI211_X1 U21040 ( .C1(n18394), .C2(n18131), .A(n18057), .B(n18056), .ZN(
        P3_U2869) );
  INV_X1 U21041 ( .A(n18086), .ZN(n18077) );
  NAND2_X1 U21042 ( .A1(n18077), .A2(n18058), .ZN(n18443) );
  AND2_X1 U21043 ( .A1(n18426), .A2(BUF2_REG_18__SCAN_IN), .ZN(n18440) );
  NOR2_X2 U21044 ( .A1(n18083), .A2(n18059), .ZN(n18438) );
  AOI22_X1 U21045 ( .A1(n18440), .A2(n18413), .B1(n18438), .B2(n18085), .ZN(
        n18062) );
  NOR2_X2 U21046 ( .A1(n18060), .A2(n18078), .ZN(n18439) );
  AOI22_X1 U21047 ( .A1(P3_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n18088), .B1(
        n18439), .B2(n18464), .ZN(n18061) );
  OAI211_X1 U21048 ( .C1(n18443), .C2(n18131), .A(n18062), .B(n18061), .ZN(
        P3_U2870) );
  NAND2_X1 U21049 ( .A1(n18077), .A2(n18063), .ZN(n18449) );
  NOR2_X2 U21050 ( .A1(n18078), .A2(n19158), .ZN(n18446) );
  NOR2_X2 U21051 ( .A1(n18083), .A2(n18064), .ZN(n18444) );
  AOI22_X1 U21052 ( .A1(n18446), .A2(n18413), .B1(n18444), .B2(n18085), .ZN(
        n18066) );
  AND2_X1 U21053 ( .A1(BUF2_REG_27__SCAN_IN), .A2(n18426), .ZN(n18445) );
  AOI22_X1 U21054 ( .A1(P3_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n18088), .B1(
        n18445), .B2(n18464), .ZN(n18065) );
  OAI211_X1 U21055 ( .C1(n18449), .C2(n18131), .A(n18066), .B(n18065), .ZN(
        P3_U2871) );
  NAND2_X1 U21056 ( .A1(BUF2_REG_28__SCAN_IN), .A2(n18426), .ZN(n18402) );
  NOR2_X2 U21057 ( .A1(n18078), .A2(n19164), .ZN(n18452) );
  NOR2_X2 U21058 ( .A1(n18083), .A2(n18067), .ZN(n18450) );
  AOI22_X1 U21059 ( .A1(n18452), .A2(n18413), .B1(n18450), .B2(n18085), .ZN(
        n18070) );
  NOR2_X1 U21060 ( .A1(n18068), .A2(n18086), .ZN(n18399) );
  AOI22_X1 U21061 ( .A1(P3_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n18088), .B1(
        n18399), .B2(n18151), .ZN(n18069) );
  OAI211_X1 U21062 ( .C1(n18402), .C2(n18479), .A(n18070), .B(n18069), .ZN(
        P3_U2872) );
  NOR2_X1 U21063 ( .A1(n18071), .A2(n18086), .ZN(n18403) );
  INV_X1 U21064 ( .A(n18403), .ZN(n18461) );
  NAND2_X1 U21065 ( .A1(BUF2_REG_29__SCAN_IN), .A2(n18426), .ZN(n18406) );
  INV_X1 U21066 ( .A(n18406), .ZN(n18457) );
  NOR2_X2 U21067 ( .A1(n18083), .A2(n18072), .ZN(n18456) );
  AOI22_X1 U21068 ( .A1(n18457), .A2(n18464), .B1(n18456), .B2(n18085), .ZN(
        n18075) );
  NOR2_X2 U21069 ( .A1(n18078), .A2(n18073), .ZN(n18458) );
  AOI22_X1 U21070 ( .A1(P3_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n18088), .B1(
        n18458), .B2(n18413), .ZN(n18074) );
  OAI211_X1 U21071 ( .C1(n18461), .C2(n18131), .A(n18075), .B(n18074), .ZN(
        P3_U2873) );
  NAND2_X1 U21072 ( .A1(n18077), .A2(n18076), .ZN(n18469) );
  NOR2_X2 U21073 ( .A1(n18079), .A2(n18078), .ZN(n18463) );
  NOR2_X2 U21074 ( .A1(n18083), .A2(n18080), .ZN(n18462) );
  AOI22_X1 U21075 ( .A1(n18463), .A2(n18464), .B1(n18462), .B2(n18085), .ZN(
        n18082) );
  AND2_X1 U21076 ( .A1(n18426), .A2(BUF2_REG_22__SCAN_IN), .ZN(n18465) );
  AOI22_X1 U21077 ( .A1(P3_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n18088), .B1(
        n18465), .B2(n18413), .ZN(n18081) );
  OAI211_X1 U21078 ( .C1(n18469), .C2(n18131), .A(n18082), .B(n18081), .ZN(
        P3_U2874) );
  NAND2_X1 U21079 ( .A1(BUF2_REG_23__SCAN_IN), .A2(n18426), .ZN(n18480) );
  NAND2_X1 U21080 ( .A1(n18426), .A2(BUF2_REG_31__SCAN_IN), .ZN(n18418) );
  INV_X1 U21081 ( .A(n18418), .ZN(n18473) );
  NOR2_X2 U21082 ( .A1(n18084), .A2(n18083), .ZN(n18471) );
  AOI22_X1 U21083 ( .A1(n18473), .A2(n18464), .B1(n18471), .B2(n18085), .ZN(
        n18090) );
  NOR2_X2 U21084 ( .A1(n18087), .A2(n18086), .ZN(n18475) );
  AOI22_X1 U21085 ( .A1(P3_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n18088), .B1(
        n18475), .B2(n18151), .ZN(n18089) );
  OAI211_X1 U21086 ( .C1(n18480), .C2(n18410), .A(n18090), .B(n18089), .ZN(
        P3_U2875) );
  NAND2_X1 U21087 ( .A1(n18269), .A2(n18110), .ZN(n18175) );
  NAND2_X1 U21088 ( .A1(n18517), .A2(n18544), .ZN(n18359) );
  NOR2_X1 U21089 ( .A1(n18133), .A2(n18359), .ZN(n18106) );
  AOI22_X1 U21090 ( .A1(n18422), .A2(n18413), .B1(n18421), .B2(n18106), .ZN(
        n18093) );
  NAND2_X1 U21091 ( .A1(n18388), .A2(n18091), .ZN(n18222) );
  NOR2_X1 U21092 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18222), .ZN(
        n18361) );
  AOI22_X1 U21093 ( .A1(n18426), .A2(n18424), .B1(n18110), .B2(n18361), .ZN(
        n18107) );
  AOI22_X1 U21094 ( .A1(P3_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n18107), .B1(
        n18427), .B2(n18474), .ZN(n18092) );
  OAI211_X1 U21095 ( .C1(n18175), .C2(n18430), .A(n18093), .B(n18092), .ZN(
        P3_U2876) );
  AOI22_X1 U21096 ( .A1(n18391), .A2(n18413), .B1(n18432), .B2(n18106), .ZN(
        n18095) );
  AOI22_X1 U21097 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n18107), .B1(
        n18431), .B2(n18474), .ZN(n18094) );
  OAI211_X1 U21098 ( .C1(n18175), .C2(n18394), .A(n18095), .B(n18094), .ZN(
        P3_U2877) );
  AOI22_X1 U21099 ( .A1(n18440), .A2(n18474), .B1(n18438), .B2(n18106), .ZN(
        n18097) );
  AOI22_X1 U21100 ( .A1(P3_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n18107), .B1(
        n18439), .B2(n18413), .ZN(n18096) );
  OAI211_X1 U21101 ( .C1(n18175), .C2(n18443), .A(n18097), .B(n18096), .ZN(
        P3_U2878) );
  AOI22_X1 U21102 ( .A1(n18445), .A2(n18413), .B1(n18444), .B2(n18106), .ZN(
        n18099) );
  AOI22_X1 U21103 ( .A1(P3_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n18107), .B1(
        n18446), .B2(n18474), .ZN(n18098) );
  OAI211_X1 U21104 ( .C1(n18175), .C2(n18449), .A(n18099), .B(n18098), .ZN(
        P3_U2879) );
  AOI22_X1 U21105 ( .A1(n18452), .A2(n18474), .B1(n18450), .B2(n18106), .ZN(
        n18101) );
  INV_X1 U21106 ( .A(n18175), .ZN(n18168) );
  AOI22_X1 U21107 ( .A1(P3_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n18107), .B1(
        n18168), .B2(n18399), .ZN(n18100) );
  OAI211_X1 U21108 ( .C1(n18402), .C2(n18410), .A(n18101), .B(n18100), .ZN(
        P3_U2880) );
  AOI22_X1 U21109 ( .A1(n18457), .A2(n18413), .B1(n18456), .B2(n18106), .ZN(
        n18103) );
  AOI22_X1 U21110 ( .A1(P3_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n18107), .B1(
        n18458), .B2(n18474), .ZN(n18102) );
  OAI211_X1 U21111 ( .C1(n18175), .C2(n18461), .A(n18103), .B(n18102), .ZN(
        P3_U2881) );
  AOI22_X1 U21112 ( .A1(n18463), .A2(n18413), .B1(n18462), .B2(n18106), .ZN(
        n18105) );
  AOI22_X1 U21113 ( .A1(P3_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n18107), .B1(
        n18465), .B2(n18474), .ZN(n18104) );
  OAI211_X1 U21114 ( .C1(n18175), .C2(n18469), .A(n18105), .B(n18104), .ZN(
        P3_U2882) );
  INV_X1 U21115 ( .A(n18474), .ZN(n18468) );
  AOI22_X1 U21116 ( .A1(n18473), .A2(n18413), .B1(n18471), .B2(n18106), .ZN(
        n18109) );
  AOI22_X1 U21117 ( .A1(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n18107), .B1(
        n18168), .B2(n18475), .ZN(n18108) );
  OAI211_X1 U21118 ( .C1(n18480), .C2(n18468), .A(n18109), .B(n18108), .ZN(
        P3_U2883) );
  NAND2_X1 U21119 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18110), .ZN(
        n18132) );
  NOR2_X2 U21120 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18132), .ZN(
        n18190) );
  NOR2_X1 U21121 ( .A1(n18168), .A2(n18190), .ZN(n18154) );
  NOR2_X1 U21122 ( .A1(n18420), .A2(n18154), .ZN(n18127) );
  AOI22_X1 U21123 ( .A1(n18427), .A2(n18151), .B1(n18421), .B2(n18127), .ZN(
        n18114) );
  OAI21_X1 U21124 ( .B1(n18111), .B2(n18385), .A(n18154), .ZN(n18112) );
  OAI211_X1 U21125 ( .C1(n18190), .C2(n18639), .A(n18388), .B(n18112), .ZN(
        n18128) );
  AOI22_X1 U21126 ( .A1(P3_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n18128), .B1(
        n18190), .B2(n18337), .ZN(n18113) );
  OAI211_X1 U21127 ( .C1(n18340), .C2(n18468), .A(n18114), .B(n18113), .ZN(
        P3_U2884) );
  AOI22_X1 U21128 ( .A1(n18432), .A2(n18127), .B1(n18431), .B2(n18151), .ZN(
        n18116) );
  AOI22_X1 U21129 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n18128), .B1(
        n18190), .B2(n18433), .ZN(n18115) );
  OAI211_X1 U21130 ( .C1(n18437), .C2(n18468), .A(n18116), .B(n18115), .ZN(
        P3_U2885) );
  INV_X1 U21131 ( .A(n18190), .ZN(n18197) );
  AOI22_X1 U21132 ( .A1(n18440), .A2(n18151), .B1(n18438), .B2(n18127), .ZN(
        n18118) );
  AOI22_X1 U21133 ( .A1(P3_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n18128), .B1(
        n18439), .B2(n18474), .ZN(n18117) );
  OAI211_X1 U21134 ( .C1(n18197), .C2(n18443), .A(n18118), .B(n18117), .ZN(
        P3_U2886) );
  AOI22_X1 U21135 ( .A1(n18446), .A2(n18151), .B1(n18444), .B2(n18127), .ZN(
        n18120) );
  AOI22_X1 U21136 ( .A1(P3_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n18128), .B1(
        n18445), .B2(n18474), .ZN(n18119) );
  OAI211_X1 U21137 ( .C1(n18197), .C2(n18449), .A(n18120), .B(n18119), .ZN(
        P3_U2887) );
  AOI22_X1 U21138 ( .A1(n18452), .A2(n18151), .B1(n18450), .B2(n18127), .ZN(
        n18122) );
  AOI22_X1 U21139 ( .A1(P3_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n18128), .B1(
        n18190), .B2(n18399), .ZN(n18121) );
  OAI211_X1 U21140 ( .C1(n18402), .C2(n18468), .A(n18122), .B(n18121), .ZN(
        P3_U2888) );
  AOI22_X1 U21141 ( .A1(n18456), .A2(n18127), .B1(n18458), .B2(n18151), .ZN(
        n18124) );
  AOI22_X1 U21142 ( .A1(P3_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n18128), .B1(
        n18190), .B2(n18403), .ZN(n18123) );
  OAI211_X1 U21143 ( .C1(n18406), .C2(n18468), .A(n18124), .B(n18123), .ZN(
        P3_U2889) );
  AOI22_X1 U21144 ( .A1(n18465), .A2(n18151), .B1(n18462), .B2(n18127), .ZN(
        n18126) );
  AOI22_X1 U21145 ( .A1(P3_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n18128), .B1(
        n18463), .B2(n18474), .ZN(n18125) );
  OAI211_X1 U21146 ( .C1(n18197), .C2(n18469), .A(n18126), .B(n18125), .ZN(
        P3_U2890) );
  AOI22_X1 U21147 ( .A1(n18473), .A2(n18474), .B1(n18471), .B2(n18127), .ZN(
        n18130) );
  AOI22_X1 U21148 ( .A1(P3_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n18128), .B1(
        n18190), .B2(n18475), .ZN(n18129) );
  OAI211_X1 U21149 ( .C1(n18480), .C2(n18131), .A(n18130), .B(n18129), .ZN(
        P3_U2891) );
  INV_X1 U21150 ( .A(n18132), .ZN(n18177) );
  NAND2_X1 U21151 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18177), .ZN(
        n18221) );
  NOR2_X1 U21152 ( .A1(n18420), .A2(n18132), .ZN(n18149) );
  AOI22_X1 U21153 ( .A1(n18422), .A2(n18151), .B1(n18421), .B2(n18149), .ZN(
        n18136) );
  OAI21_X1 U21154 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(n18133), .A(n18221), 
        .ZN(n18134) );
  NAND3_X1 U21155 ( .A1(n18388), .A2(n18223), .A3(n18134), .ZN(n18150) );
  AOI22_X1 U21156 ( .A1(P3_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n18150), .B1(
        n18168), .B2(n18427), .ZN(n18135) );
  OAI211_X1 U21157 ( .C1(n18221), .C2(n18430), .A(n18136), .B(n18135), .ZN(
        P3_U2892) );
  AOI22_X1 U21158 ( .A1(n18168), .A2(n18431), .B1(n18432), .B2(n18149), .ZN(
        n18138) );
  AOI22_X1 U21159 ( .A1(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n18150), .B1(
        n18391), .B2(n18151), .ZN(n18137) );
  OAI211_X1 U21160 ( .C1(n18221), .C2(n18394), .A(n18138), .B(n18137), .ZN(
        P3_U2893) );
  AOI22_X1 U21161 ( .A1(P3_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n18150), .B1(
        n18438), .B2(n18149), .ZN(n18140) );
  AOI22_X1 U21162 ( .A1(n18168), .A2(n18440), .B1(n18439), .B2(n18151), .ZN(
        n18139) );
  OAI211_X1 U21163 ( .C1(n18221), .C2(n18443), .A(n18140), .B(n18139), .ZN(
        P3_U2894) );
  AOI22_X1 U21164 ( .A1(n18445), .A2(n18151), .B1(n18444), .B2(n18149), .ZN(
        n18142) );
  AOI22_X1 U21165 ( .A1(P3_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n18150), .B1(
        n18168), .B2(n18446), .ZN(n18141) );
  OAI211_X1 U21166 ( .C1(n18221), .C2(n18449), .A(n18142), .B(n18141), .ZN(
        P3_U2895) );
  INV_X1 U21167 ( .A(n18399), .ZN(n18455) );
  INV_X1 U21168 ( .A(n18402), .ZN(n18451) );
  AOI22_X1 U21169 ( .A1(n18451), .A2(n18151), .B1(n18450), .B2(n18149), .ZN(
        n18144) );
  AOI22_X1 U21170 ( .A1(P3_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n18150), .B1(
        n18168), .B2(n18452), .ZN(n18143) );
  OAI211_X1 U21171 ( .C1(n18221), .C2(n18455), .A(n18144), .B(n18143), .ZN(
        P3_U2896) );
  AOI22_X1 U21172 ( .A1(n18168), .A2(n18458), .B1(n18456), .B2(n18149), .ZN(
        n18146) );
  AOI22_X1 U21173 ( .A1(P3_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n18150), .B1(
        n18457), .B2(n18151), .ZN(n18145) );
  OAI211_X1 U21174 ( .C1(n18221), .C2(n18461), .A(n18146), .B(n18145), .ZN(
        P3_U2897) );
  AOI22_X1 U21175 ( .A1(n18463), .A2(n18151), .B1(n18462), .B2(n18149), .ZN(
        n18148) );
  AOI22_X1 U21176 ( .A1(P3_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n18150), .B1(
        n18168), .B2(n18465), .ZN(n18147) );
  OAI211_X1 U21177 ( .C1(n18221), .C2(n18469), .A(n18148), .B(n18147), .ZN(
        P3_U2898) );
  AOI22_X1 U21178 ( .A1(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n18150), .B1(
        n18471), .B2(n18149), .ZN(n18153) );
  INV_X1 U21179 ( .A(n18221), .ZN(n18213) );
  AOI22_X1 U21180 ( .A1(n18213), .A2(n18475), .B1(n18473), .B2(n18151), .ZN(
        n18152) );
  OAI211_X1 U21181 ( .C1(n18175), .C2(n18480), .A(n18153), .B(n18152), .ZN(
        P3_U2899) );
  INV_X1 U21182 ( .A(n18224), .ZN(n18176) );
  NOR2_X1 U21183 ( .A1(n18518), .A2(n18176), .ZN(n18239) );
  INV_X1 U21184 ( .A(n18239), .ZN(n18246) );
  AOI21_X1 U21185 ( .B1(n18246), .B2(n18221), .A(n18420), .ZN(n18171) );
  AOI22_X1 U21186 ( .A1(n18190), .A2(n18427), .B1(n18421), .B2(n18171), .ZN(
        n18157) );
  CLKBUF_X1 U21187 ( .A(n18239), .Z(n18236) );
  AOI221_X1 U21188 ( .B1(n18154), .B2(n18221), .C1(n18385), .C2(n18221), .A(
        P3_STATE2_REG_3__SCAN_IN), .ZN(n18155) );
  OAI21_X1 U21189 ( .B1(n18236), .B2(n18155), .A(n18388), .ZN(n18172) );
  AOI22_X1 U21190 ( .A1(P3_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n18172), .B1(
        n18239), .B2(n18337), .ZN(n18156) );
  OAI211_X1 U21191 ( .C1(n18340), .C2(n18175), .A(n18157), .B(n18156), .ZN(
        P3_U2900) );
  AOI22_X1 U21192 ( .A1(n18190), .A2(n18431), .B1(n18171), .B2(n18432), .ZN(
        n18159) );
  AOI22_X1 U21193 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n18172), .B1(
        n18236), .B2(n18433), .ZN(n18158) );
  OAI211_X1 U21194 ( .C1(n18175), .C2(n18437), .A(n18159), .B(n18158), .ZN(
        P3_U2901) );
  AOI22_X1 U21195 ( .A1(n18168), .A2(n18439), .B1(n18171), .B2(n18438), .ZN(
        n18161) );
  AOI22_X1 U21196 ( .A1(P3_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n18172), .B1(
        n18190), .B2(n18440), .ZN(n18160) );
  OAI211_X1 U21197 ( .C1(n18246), .C2(n18443), .A(n18161), .B(n18160), .ZN(
        P3_U2902) );
  AOI22_X1 U21198 ( .A1(n18168), .A2(n18445), .B1(n18171), .B2(n18444), .ZN(
        n18163) );
  AOI22_X1 U21199 ( .A1(P3_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n18172), .B1(
        n18190), .B2(n18446), .ZN(n18162) );
  OAI211_X1 U21200 ( .C1(n18246), .C2(n18449), .A(n18163), .B(n18162), .ZN(
        P3_U2903) );
  AOI22_X1 U21201 ( .A1(n18190), .A2(n18452), .B1(n18171), .B2(n18450), .ZN(
        n18165) );
  AOI22_X1 U21202 ( .A1(P3_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n18172), .B1(
        n18239), .B2(n18399), .ZN(n18164) );
  OAI211_X1 U21203 ( .C1(n18175), .C2(n18402), .A(n18165), .B(n18164), .ZN(
        P3_U2904) );
  AOI22_X1 U21204 ( .A1(n18190), .A2(n18458), .B1(n18171), .B2(n18456), .ZN(
        n18167) );
  AOI22_X1 U21205 ( .A1(P3_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n18172), .B1(
        n18239), .B2(n18403), .ZN(n18166) );
  OAI211_X1 U21206 ( .C1(n18175), .C2(n18406), .A(n18167), .B(n18166), .ZN(
        P3_U2905) );
  AOI22_X1 U21207 ( .A1(n18168), .A2(n18463), .B1(n18171), .B2(n18462), .ZN(
        n18170) );
  AOI22_X1 U21208 ( .A1(P3_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n18172), .B1(
        n18190), .B2(n18465), .ZN(n18169) );
  OAI211_X1 U21209 ( .C1(n18246), .C2(n18469), .A(n18170), .B(n18169), .ZN(
        P3_U2906) );
  INV_X1 U21210 ( .A(n18480), .ZN(n18412) );
  AOI22_X1 U21211 ( .A1(n18190), .A2(n18412), .B1(n18171), .B2(n18471), .ZN(
        n18174) );
  AOI22_X1 U21212 ( .A1(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n18172), .B1(
        n18239), .B2(n18475), .ZN(n18173) );
  OAI211_X1 U21213 ( .C1(n18175), .C2(n18418), .A(n18174), .B(n18173), .ZN(
        P3_U2907) );
  NOR2_X1 U21214 ( .A1(n18176), .A2(n18359), .ZN(n18193) );
  AOI22_X1 U21215 ( .A1(n18213), .A2(n18427), .B1(n18421), .B2(n18193), .ZN(
        n18179) );
  AOI22_X1 U21216 ( .A1(n18426), .A2(n18177), .B1(n18224), .B2(n18361), .ZN(
        n18194) );
  NAND2_X1 U21217 ( .A1(n18269), .A2(n18224), .ZN(n18268) );
  INV_X1 U21218 ( .A(n18268), .ZN(n18261) );
  AOI22_X1 U21219 ( .A1(P3_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n18194), .B1(
        n18337), .B2(n18261), .ZN(n18178) );
  OAI211_X1 U21220 ( .C1(n18340), .C2(n18197), .A(n18179), .B(n18178), .ZN(
        P3_U2908) );
  AOI22_X1 U21221 ( .A1(n18213), .A2(n18431), .B1(n18432), .B2(n18193), .ZN(
        n18181) );
  AOI22_X1 U21222 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n18194), .B1(
        n18433), .B2(n18261), .ZN(n18180) );
  OAI211_X1 U21223 ( .C1(n18197), .C2(n18437), .A(n18181), .B(n18180), .ZN(
        P3_U2909) );
  AOI22_X1 U21224 ( .A1(n18213), .A2(n18440), .B1(n18438), .B2(n18193), .ZN(
        n18183) );
  AOI22_X1 U21225 ( .A1(P3_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n18194), .B1(
        n18190), .B2(n18439), .ZN(n18182) );
  OAI211_X1 U21226 ( .C1(n18443), .C2(n18268), .A(n18183), .B(n18182), .ZN(
        P3_U2910) );
  AOI22_X1 U21227 ( .A1(n18190), .A2(n18445), .B1(n18444), .B2(n18193), .ZN(
        n18185) );
  AOI22_X1 U21228 ( .A1(P3_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n18194), .B1(
        n18213), .B2(n18446), .ZN(n18184) );
  OAI211_X1 U21229 ( .C1(n18449), .C2(n18268), .A(n18185), .B(n18184), .ZN(
        P3_U2911) );
  AOI22_X1 U21230 ( .A1(n18190), .A2(n18451), .B1(n18450), .B2(n18193), .ZN(
        n18187) );
  AOI22_X1 U21231 ( .A1(P3_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n18194), .B1(
        n18213), .B2(n18452), .ZN(n18186) );
  OAI211_X1 U21232 ( .C1(n18455), .C2(n18268), .A(n18187), .B(n18186), .ZN(
        P3_U2912) );
  AOI22_X1 U21233 ( .A1(n18213), .A2(n18458), .B1(n18456), .B2(n18193), .ZN(
        n18189) );
  AOI22_X1 U21234 ( .A1(P3_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n18194), .B1(
        n18403), .B2(n18261), .ZN(n18188) );
  OAI211_X1 U21235 ( .C1(n18197), .C2(n18406), .A(n18189), .B(n18188), .ZN(
        P3_U2913) );
  AOI22_X1 U21236 ( .A1(n18213), .A2(n18465), .B1(n18462), .B2(n18193), .ZN(
        n18192) );
  AOI22_X1 U21237 ( .A1(P3_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n18194), .B1(
        n18190), .B2(n18463), .ZN(n18191) );
  OAI211_X1 U21238 ( .C1(n18469), .C2(n18268), .A(n18192), .B(n18191), .ZN(
        P3_U2914) );
  AOI22_X1 U21239 ( .A1(n18213), .A2(n18412), .B1(n18471), .B2(n18193), .ZN(
        n18196) );
  AOI22_X1 U21240 ( .A1(P3_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n18194), .B1(
        n18475), .B2(n18261), .ZN(n18195) );
  OAI211_X1 U21241 ( .C1(n18197), .C2(n18418), .A(n18196), .B(n18195), .ZN(
        P3_U2915) );
  NOR2_X1 U21242 ( .A1(n18198), .A2(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n18271) );
  INV_X1 U21243 ( .A(n18271), .ZN(n18225) );
  OR2_X1 U21244 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18225), .ZN(
        n18216) );
  INV_X1 U21245 ( .A(n18216), .ZN(n18286) );
  NOR2_X1 U21246 ( .A1(n18261), .A2(n18286), .ZN(n18247) );
  NOR2_X1 U21247 ( .A1(n18420), .A2(n18247), .ZN(n18217) );
  AOI22_X1 U21248 ( .A1(n18236), .A2(n18427), .B1(n18421), .B2(n18217), .ZN(
        n18202) );
  NOR2_X1 U21249 ( .A1(n18236), .A2(n18213), .ZN(n18199) );
  OAI21_X1 U21250 ( .B1(n18199), .B2(n18385), .A(n18247), .ZN(n18200) );
  OAI211_X1 U21251 ( .C1(n18286), .C2(n18639), .A(n18388), .B(n18200), .ZN(
        n18218) );
  AOI22_X1 U21252 ( .A1(P3_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n18218), .B1(
        n18337), .B2(n18286), .ZN(n18201) );
  OAI211_X1 U21253 ( .C1(n18340), .C2(n18221), .A(n18202), .B(n18201), .ZN(
        P3_U2916) );
  AOI22_X1 U21254 ( .A1(n18236), .A2(n18431), .B1(n18432), .B2(n18217), .ZN(
        n18204) );
  AOI22_X1 U21255 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n18218), .B1(
        n18433), .B2(n18286), .ZN(n18203) );
  OAI211_X1 U21256 ( .C1(n18221), .C2(n18437), .A(n18204), .B(n18203), .ZN(
        P3_U2917) );
  AOI22_X1 U21257 ( .A1(n18213), .A2(n18439), .B1(n18438), .B2(n18217), .ZN(
        n18206) );
  AOI22_X1 U21258 ( .A1(P3_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n18218), .B1(
        n18239), .B2(n18440), .ZN(n18205) );
  OAI211_X1 U21259 ( .C1(n18443), .C2(n18216), .A(n18206), .B(n18205), .ZN(
        P3_U2918) );
  AOI22_X1 U21260 ( .A1(n18213), .A2(n18445), .B1(n18444), .B2(n18217), .ZN(
        n18208) );
  AOI22_X1 U21261 ( .A1(P3_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n18218), .B1(
        n18236), .B2(n18446), .ZN(n18207) );
  OAI211_X1 U21262 ( .C1(n18449), .C2(n18216), .A(n18208), .B(n18207), .ZN(
        P3_U2919) );
  AOI22_X1 U21263 ( .A1(n18236), .A2(n18452), .B1(n18450), .B2(n18217), .ZN(
        n18210) );
  AOI22_X1 U21264 ( .A1(P3_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n18218), .B1(
        n18399), .B2(n18286), .ZN(n18209) );
  OAI211_X1 U21265 ( .C1(n18221), .C2(n18402), .A(n18210), .B(n18209), .ZN(
        P3_U2920) );
  AOI22_X1 U21266 ( .A1(n18239), .A2(n18458), .B1(n18456), .B2(n18217), .ZN(
        n18212) );
  AOI22_X1 U21267 ( .A1(P3_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n18218), .B1(
        n18403), .B2(n18286), .ZN(n18211) );
  OAI211_X1 U21268 ( .C1(n18221), .C2(n18406), .A(n18212), .B(n18211), .ZN(
        P3_U2921) );
  AOI22_X1 U21269 ( .A1(n18213), .A2(n18463), .B1(n18462), .B2(n18217), .ZN(
        n18215) );
  AOI22_X1 U21270 ( .A1(P3_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n18218), .B1(
        n18239), .B2(n18465), .ZN(n18214) );
  OAI211_X1 U21271 ( .C1(n18469), .C2(n18216), .A(n18215), .B(n18214), .ZN(
        P3_U2922) );
  AOI22_X1 U21272 ( .A1(n18239), .A2(n18412), .B1(n18471), .B2(n18217), .ZN(
        n18220) );
  AOI22_X1 U21273 ( .A1(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n18218), .B1(
        n18475), .B2(n18286), .ZN(n18219) );
  OAI211_X1 U21274 ( .C1(n18221), .C2(n18418), .A(n18220), .B(n18219), .ZN(
        P3_U2923) );
  NAND2_X1 U21275 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18271), .ZN(
        n18305) );
  INV_X1 U21276 ( .A(n18222), .ZN(n18423) );
  NAND3_X1 U21277 ( .A1(n18423), .A2(n18224), .A3(n18223), .ZN(n18243) );
  NOR2_X1 U21278 ( .A1(n18420), .A2(n18225), .ZN(n18242) );
  AOI22_X1 U21279 ( .A1(P3_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n18243), .B1(
        n18421), .B2(n18242), .ZN(n18227) );
  AOI22_X1 U21280 ( .A1(n18422), .A2(n18239), .B1(n18427), .B2(n18261), .ZN(
        n18226) );
  OAI211_X1 U21281 ( .C1(n18430), .C2(n18305), .A(n18227), .B(n18226), .ZN(
        P3_U2924) );
  AOI22_X1 U21282 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n18243), .B1(
        n18432), .B2(n18242), .ZN(n18229) );
  AOI22_X1 U21283 ( .A1(n18236), .A2(n18391), .B1(n18431), .B2(n18261), .ZN(
        n18228) );
  OAI211_X1 U21284 ( .C1(n18394), .C2(n18305), .A(n18229), .B(n18228), .ZN(
        P3_U2925) );
  AOI22_X1 U21285 ( .A1(P3_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n18243), .B1(
        n18438), .B2(n18242), .ZN(n18231) );
  AOI22_X1 U21286 ( .A1(n18236), .A2(n18439), .B1(n18440), .B2(n18261), .ZN(
        n18230) );
  OAI211_X1 U21287 ( .C1(n18443), .C2(n18305), .A(n18231), .B(n18230), .ZN(
        P3_U2926) );
  AOI22_X1 U21288 ( .A1(P3_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n18243), .B1(
        n18444), .B2(n18242), .ZN(n18233) );
  AOI22_X1 U21289 ( .A1(n18236), .A2(n18445), .B1(n18446), .B2(n18261), .ZN(
        n18232) );
  OAI211_X1 U21290 ( .C1(n18449), .C2(n18305), .A(n18233), .B(n18232), .ZN(
        P3_U2927) );
  AOI22_X1 U21291 ( .A1(n18236), .A2(n18451), .B1(n18450), .B2(n18242), .ZN(
        n18235) );
  AOI22_X1 U21292 ( .A1(P3_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n18243), .B1(
        n18452), .B2(n18261), .ZN(n18234) );
  OAI211_X1 U21293 ( .C1(n18455), .C2(n18305), .A(n18235), .B(n18234), .ZN(
        P3_U2928) );
  AOI22_X1 U21294 ( .A1(n18456), .A2(n18242), .B1(n18458), .B2(n18261), .ZN(
        n18238) );
  AOI22_X1 U21295 ( .A1(P3_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n18243), .B1(
        n18236), .B2(n18457), .ZN(n18237) );
  OAI211_X1 U21296 ( .C1(n18461), .C2(n18305), .A(n18238), .B(n18237), .ZN(
        P3_U2929) );
  AOI22_X1 U21297 ( .A1(P3_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n18243), .B1(
        n18462), .B2(n18242), .ZN(n18241) );
  AOI22_X1 U21298 ( .A1(n18239), .A2(n18463), .B1(n18465), .B2(n18261), .ZN(
        n18240) );
  OAI211_X1 U21299 ( .C1(n18469), .C2(n18305), .A(n18241), .B(n18240), .ZN(
        P3_U2930) );
  AOI22_X1 U21300 ( .A1(n18412), .A2(n18261), .B1(n18471), .B2(n18242), .ZN(
        n18245) );
  INV_X1 U21301 ( .A(n18305), .ZN(n18309) );
  AOI22_X1 U21302 ( .A1(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n18243), .B1(
        n18475), .B2(n18309), .ZN(n18244) );
  OAI211_X1 U21303 ( .C1(n18246), .C2(n18418), .A(n18245), .B(n18244), .ZN(
        P3_U2931) );
  INV_X1 U21304 ( .A(n18290), .ZN(n18270) );
  NOR2_X2 U21305 ( .A1(n18518), .A2(n18270), .ZN(n18327) );
  INV_X1 U21306 ( .A(n18327), .ZN(n18334) );
  AOI21_X1 U21307 ( .B1(n18334), .B2(n18305), .A(n18420), .ZN(n18264) );
  AOI22_X1 U21308 ( .A1(n18427), .A2(n18286), .B1(n18421), .B2(n18264), .ZN(
        n18250) );
  AOI221_X1 U21309 ( .B1(n18247), .B2(n18305), .C1(n18385), .C2(n18305), .A(
        P3_STATE2_REG_3__SCAN_IN), .ZN(n18248) );
  OAI21_X1 U21310 ( .B1(n18327), .B2(n18248), .A(n18388), .ZN(n18265) );
  AOI22_X1 U21311 ( .A1(P3_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n18265), .B1(
        n18337), .B2(n18327), .ZN(n18249) );
  OAI211_X1 U21312 ( .C1(n18340), .C2(n18268), .A(n18250), .B(n18249), .ZN(
        P3_U2932) );
  AOI22_X1 U21313 ( .A1(n18391), .A2(n18261), .B1(n18432), .B2(n18264), .ZN(
        n18252) );
  AOI22_X1 U21314 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n18265), .B1(
        n18431), .B2(n18286), .ZN(n18251) );
  OAI211_X1 U21315 ( .C1(n18394), .C2(n18334), .A(n18252), .B(n18251), .ZN(
        P3_U2933) );
  AOI22_X1 U21316 ( .A1(n18440), .A2(n18286), .B1(n18438), .B2(n18264), .ZN(
        n18254) );
  AOI22_X1 U21317 ( .A1(P3_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n18265), .B1(
        n18439), .B2(n18261), .ZN(n18253) );
  OAI211_X1 U21318 ( .C1(n18443), .C2(n18334), .A(n18254), .B(n18253), .ZN(
        P3_U2934) );
  AOI22_X1 U21319 ( .A1(n18445), .A2(n18261), .B1(n18444), .B2(n18264), .ZN(
        n18256) );
  AOI22_X1 U21320 ( .A1(P3_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n18265), .B1(
        n18446), .B2(n18286), .ZN(n18255) );
  OAI211_X1 U21321 ( .C1(n18449), .C2(n18334), .A(n18256), .B(n18255), .ZN(
        P3_U2935) );
  AOI22_X1 U21322 ( .A1(n18451), .A2(n18261), .B1(n18450), .B2(n18264), .ZN(
        n18258) );
  AOI22_X1 U21323 ( .A1(P3_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n18265), .B1(
        n18452), .B2(n18286), .ZN(n18257) );
  OAI211_X1 U21324 ( .C1(n18455), .C2(n18334), .A(n18258), .B(n18257), .ZN(
        P3_U2936) );
  AOI22_X1 U21325 ( .A1(n18457), .A2(n18261), .B1(n18456), .B2(n18264), .ZN(
        n18260) );
  AOI22_X1 U21326 ( .A1(P3_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n18265), .B1(
        n18458), .B2(n18286), .ZN(n18259) );
  OAI211_X1 U21327 ( .C1(n18461), .C2(n18334), .A(n18260), .B(n18259), .ZN(
        P3_U2937) );
  AOI22_X1 U21328 ( .A1(n18465), .A2(n18286), .B1(n18462), .B2(n18264), .ZN(
        n18263) );
  AOI22_X1 U21329 ( .A1(P3_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n18265), .B1(
        n18463), .B2(n18261), .ZN(n18262) );
  OAI211_X1 U21330 ( .C1(n18469), .C2(n18334), .A(n18263), .B(n18262), .ZN(
        P3_U2938) );
  AOI22_X1 U21331 ( .A1(n18412), .A2(n18286), .B1(n18471), .B2(n18264), .ZN(
        n18267) );
  AOI22_X1 U21332 ( .A1(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n18265), .B1(
        n18475), .B2(n18327), .ZN(n18266) );
  OAI211_X1 U21333 ( .C1(n18418), .C2(n18268), .A(n18267), .B(n18266), .ZN(
        P3_U2939) );
  NAND2_X1 U21334 ( .A1(n18269), .A2(n18290), .ZN(n18358) );
  NOR2_X1 U21335 ( .A1(n18270), .A2(n18359), .ZN(n18314) );
  AOI22_X1 U21336 ( .A1(n18422), .A2(n18286), .B1(n18421), .B2(n18314), .ZN(
        n18273) );
  AOI22_X1 U21337 ( .A1(n18426), .A2(n18271), .B1(n18290), .B2(n18361), .ZN(
        n18287) );
  AOI22_X1 U21338 ( .A1(P3_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n18287), .B1(
        n18427), .B2(n18309), .ZN(n18272) );
  OAI211_X1 U21339 ( .C1(n18430), .C2(n18358), .A(n18273), .B(n18272), .ZN(
        P3_U2940) );
  AOI22_X1 U21340 ( .A1(n18391), .A2(n18286), .B1(n18432), .B2(n18314), .ZN(
        n18275) );
  AOI22_X1 U21341 ( .A1(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n18287), .B1(
        n18431), .B2(n18309), .ZN(n18274) );
  OAI211_X1 U21342 ( .C1(n18394), .C2(n18358), .A(n18275), .B(n18274), .ZN(
        P3_U2941) );
  AOI22_X1 U21343 ( .A1(n18439), .A2(n18286), .B1(n18438), .B2(n18314), .ZN(
        n18277) );
  AOI22_X1 U21344 ( .A1(P3_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n18287), .B1(
        n18440), .B2(n18309), .ZN(n18276) );
  OAI211_X1 U21345 ( .C1(n18443), .C2(n18358), .A(n18277), .B(n18276), .ZN(
        P3_U2942) );
  AOI22_X1 U21346 ( .A1(n18445), .A2(n18286), .B1(n18444), .B2(n18314), .ZN(
        n18279) );
  AOI22_X1 U21347 ( .A1(P3_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n18287), .B1(
        n18446), .B2(n18309), .ZN(n18278) );
  OAI211_X1 U21348 ( .C1(n18449), .C2(n18358), .A(n18279), .B(n18278), .ZN(
        P3_U2943) );
  AOI22_X1 U21349 ( .A1(n18451), .A2(n18286), .B1(n18450), .B2(n18314), .ZN(
        n18281) );
  AOI22_X1 U21350 ( .A1(P3_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n18287), .B1(
        n18452), .B2(n18309), .ZN(n18280) );
  OAI211_X1 U21351 ( .C1(n18455), .C2(n18358), .A(n18281), .B(n18280), .ZN(
        P3_U2944) );
  AOI22_X1 U21352 ( .A1(n18457), .A2(n18286), .B1(n18456), .B2(n18314), .ZN(
        n18283) );
  AOI22_X1 U21353 ( .A1(P3_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n18287), .B1(
        n18458), .B2(n18309), .ZN(n18282) );
  OAI211_X1 U21354 ( .C1(n18461), .C2(n18358), .A(n18283), .B(n18282), .ZN(
        P3_U2945) );
  AOI22_X1 U21355 ( .A1(n18463), .A2(n18286), .B1(n18462), .B2(n18314), .ZN(
        n18285) );
  AOI22_X1 U21356 ( .A1(P3_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n18287), .B1(
        n18465), .B2(n18309), .ZN(n18284) );
  OAI211_X1 U21357 ( .C1(n18469), .C2(n18358), .A(n18285), .B(n18284), .ZN(
        P3_U2946) );
  AOI22_X1 U21358 ( .A1(n18473), .A2(n18286), .B1(n18471), .B2(n18314), .ZN(
        n18289) );
  INV_X1 U21359 ( .A(n18358), .ZN(n18351) );
  AOI22_X1 U21360 ( .A1(P3_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n18287), .B1(
        n18475), .B2(n18351), .ZN(n18288) );
  OAI211_X1 U21361 ( .C1(n18480), .C2(n18305), .A(n18289), .B(n18288), .ZN(
        P3_U2947) );
  NAND2_X1 U21362 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18290), .ZN(
        n18313) );
  NOR2_X2 U21363 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18313), .ZN(
        n18376) );
  INV_X1 U21364 ( .A(n18376), .ZN(n18382) );
  NOR2_X1 U21365 ( .A1(n18351), .A2(n18376), .ZN(n18335) );
  NOR2_X1 U21366 ( .A1(n18420), .A2(n18335), .ZN(n18308) );
  AOI22_X1 U21367 ( .A1(n18422), .A2(n18309), .B1(n18421), .B2(n18308), .ZN(
        n18294) );
  NOR2_X1 U21368 ( .A1(n18327), .A2(n18309), .ZN(n18291) );
  OAI21_X1 U21369 ( .B1(n18291), .B2(n18385), .A(n18335), .ZN(n18292) );
  OAI211_X1 U21370 ( .C1(n18376), .C2(n18639), .A(n18388), .B(n18292), .ZN(
        n18310) );
  AOI22_X1 U21371 ( .A1(P3_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n18310), .B1(
        n18427), .B2(n18327), .ZN(n18293) );
  OAI211_X1 U21372 ( .C1(n18430), .C2(n18382), .A(n18294), .B(n18293), .ZN(
        P3_U2948) );
  AOI22_X1 U21373 ( .A1(n18432), .A2(n18308), .B1(n18431), .B2(n18327), .ZN(
        n18296) );
  AOI22_X1 U21374 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n18310), .B1(
        n18433), .B2(n18376), .ZN(n18295) );
  OAI211_X1 U21375 ( .C1(n18437), .C2(n18305), .A(n18296), .B(n18295), .ZN(
        P3_U2949) );
  AOI22_X1 U21376 ( .A1(n18440), .A2(n18327), .B1(n18438), .B2(n18308), .ZN(
        n18298) );
  AOI22_X1 U21377 ( .A1(P3_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n18310), .B1(
        n18439), .B2(n18309), .ZN(n18297) );
  OAI211_X1 U21378 ( .C1(n18443), .C2(n18382), .A(n18298), .B(n18297), .ZN(
        P3_U2950) );
  AOI22_X1 U21379 ( .A1(n18445), .A2(n18309), .B1(n18444), .B2(n18308), .ZN(
        n18300) );
  AOI22_X1 U21380 ( .A1(P3_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n18310), .B1(
        n18446), .B2(n18327), .ZN(n18299) );
  OAI211_X1 U21381 ( .C1(n18449), .C2(n18382), .A(n18300), .B(n18299), .ZN(
        P3_U2951) );
  AOI22_X1 U21382 ( .A1(n18451), .A2(n18309), .B1(n18450), .B2(n18308), .ZN(
        n18302) );
  AOI22_X1 U21383 ( .A1(P3_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n18310), .B1(
        n18452), .B2(n18327), .ZN(n18301) );
  OAI211_X1 U21384 ( .C1(n18455), .C2(n18382), .A(n18302), .B(n18301), .ZN(
        P3_U2952) );
  AOI22_X1 U21385 ( .A1(n18456), .A2(n18308), .B1(n18458), .B2(n18327), .ZN(
        n18304) );
  AOI22_X1 U21386 ( .A1(P3_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n18310), .B1(
        n18403), .B2(n18376), .ZN(n18303) );
  OAI211_X1 U21387 ( .C1(n18406), .C2(n18305), .A(n18304), .B(n18303), .ZN(
        P3_U2953) );
  AOI22_X1 U21388 ( .A1(n18463), .A2(n18309), .B1(n18462), .B2(n18308), .ZN(
        n18307) );
  AOI22_X1 U21389 ( .A1(P3_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n18310), .B1(
        n18465), .B2(n18327), .ZN(n18306) );
  OAI211_X1 U21390 ( .C1(n18469), .C2(n18382), .A(n18307), .B(n18306), .ZN(
        P3_U2954) );
  AOI22_X1 U21391 ( .A1(n18473), .A2(n18309), .B1(n18471), .B2(n18308), .ZN(
        n18312) );
  AOI22_X1 U21392 ( .A1(P3_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n18310), .B1(
        n18475), .B2(n18376), .ZN(n18311) );
  OAI211_X1 U21393 ( .C1(n18480), .C2(n18334), .A(n18312), .B(n18311), .ZN(
        P3_U2955) );
  INV_X1 U21394 ( .A(n18313), .ZN(n18363) );
  NAND2_X1 U21395 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18363), .ZN(
        n18417) );
  NOR2_X1 U21396 ( .A1(n18420), .A2(n18313), .ZN(n18330) );
  AOI22_X1 U21397 ( .A1(n18422), .A2(n18327), .B1(n18421), .B2(n18330), .ZN(
        n18316) );
  AOI22_X1 U21398 ( .A1(n18426), .A2(n18314), .B1(n18363), .B2(n18423), .ZN(
        n18331) );
  AOI22_X1 U21399 ( .A1(P3_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n18331), .B1(
        n18427), .B2(n18351), .ZN(n18315) );
  OAI211_X1 U21400 ( .C1(n18430), .C2(n18417), .A(n18316), .B(n18315), .ZN(
        P3_U2956) );
  AOI22_X1 U21401 ( .A1(n18391), .A2(n18327), .B1(n18432), .B2(n18330), .ZN(
        n18318) );
  AOI22_X1 U21402 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n18331), .B1(
        n18431), .B2(n18351), .ZN(n18317) );
  OAI211_X1 U21403 ( .C1(n18394), .C2(n18417), .A(n18318), .B(n18317), .ZN(
        P3_U2957) );
  AOI22_X1 U21404 ( .A1(n18440), .A2(n18351), .B1(n18438), .B2(n18330), .ZN(
        n18320) );
  AOI22_X1 U21405 ( .A1(P3_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n18331), .B1(
        n18439), .B2(n18327), .ZN(n18319) );
  OAI211_X1 U21406 ( .C1(n18443), .C2(n18417), .A(n18320), .B(n18319), .ZN(
        P3_U2958) );
  AOI22_X1 U21407 ( .A1(n18445), .A2(n18327), .B1(n18444), .B2(n18330), .ZN(
        n18322) );
  AOI22_X1 U21408 ( .A1(P3_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n18331), .B1(
        n18446), .B2(n18351), .ZN(n18321) );
  OAI211_X1 U21409 ( .C1(n18449), .C2(n18417), .A(n18322), .B(n18321), .ZN(
        P3_U2959) );
  AOI22_X1 U21410 ( .A1(n18452), .A2(n18351), .B1(n18450), .B2(n18330), .ZN(
        n18324) );
  AOI22_X1 U21411 ( .A1(P3_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n18331), .B1(
        n18451), .B2(n18327), .ZN(n18323) );
  OAI211_X1 U21412 ( .C1(n18455), .C2(n18417), .A(n18324), .B(n18323), .ZN(
        P3_U2960) );
  AOI22_X1 U21413 ( .A1(n18457), .A2(n18327), .B1(n18456), .B2(n18330), .ZN(
        n18326) );
  AOI22_X1 U21414 ( .A1(P3_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n18331), .B1(
        n18458), .B2(n18351), .ZN(n18325) );
  OAI211_X1 U21415 ( .C1(n18461), .C2(n18417), .A(n18326), .B(n18325), .ZN(
        P3_U2961) );
  AOI22_X1 U21416 ( .A1(n18463), .A2(n18327), .B1(n18462), .B2(n18330), .ZN(
        n18329) );
  AOI22_X1 U21417 ( .A1(P3_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n18331), .B1(
        n18465), .B2(n18351), .ZN(n18328) );
  OAI211_X1 U21418 ( .C1(n18469), .C2(n18417), .A(n18329), .B(n18328), .ZN(
        P3_U2962) );
  AOI22_X1 U21419 ( .A1(n18412), .A2(n18351), .B1(n18471), .B2(n18330), .ZN(
        n18333) );
  INV_X1 U21420 ( .A(n18417), .ZN(n18407) );
  AOI22_X1 U21421 ( .A1(P3_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n18331), .B1(
        n18475), .B2(n18407), .ZN(n18332) );
  OAI211_X1 U21422 ( .C1(n18418), .C2(n18334), .A(n18333), .B(n18332), .ZN(
        P3_U2963) );
  INV_X1 U21423 ( .A(n18362), .ZN(n18360) );
  INV_X1 U21424 ( .A(n9602), .ZN(n18436) );
  AOI21_X1 U21425 ( .B1(n18436), .B2(n18417), .A(n18420), .ZN(n18354) );
  AOI22_X1 U21426 ( .A1(n18427), .A2(n18376), .B1(n18421), .B2(n18354), .ZN(
        n18339) );
  AOI221_X1 U21427 ( .B1(n18335), .B2(n18417), .C1(n18385), .C2(n18417), .A(
        P3_STATE2_REG_3__SCAN_IN), .ZN(n18336) );
  OAI21_X1 U21428 ( .B1(n9602), .B2(n18336), .A(n18388), .ZN(n18355) );
  AOI22_X1 U21429 ( .A1(P3_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n18355), .B1(
        n18337), .B2(n9602), .ZN(n18338) );
  OAI211_X1 U21430 ( .C1(n18340), .C2(n18358), .A(n18339), .B(n18338), .ZN(
        P3_U2964) );
  AOI22_X1 U21431 ( .A1(n18432), .A2(n18354), .B1(n18431), .B2(n18376), .ZN(
        n18342) );
  AOI22_X1 U21432 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n18355), .B1(
        n18433), .B2(n9602), .ZN(n18341) );
  OAI211_X1 U21433 ( .C1(n18437), .C2(n18358), .A(n18342), .B(n18341), .ZN(
        P3_U2965) );
  AOI22_X1 U21434 ( .A1(n18439), .A2(n18351), .B1(n18438), .B2(n18354), .ZN(
        n18344) );
  AOI22_X1 U21435 ( .A1(P3_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n18355), .B1(
        n18440), .B2(n18376), .ZN(n18343) );
  OAI211_X1 U21436 ( .C1(n18443), .C2(n18436), .A(n18344), .B(n18343), .ZN(
        P3_U2966) );
  AOI22_X1 U21437 ( .A1(n18445), .A2(n18351), .B1(n18444), .B2(n18354), .ZN(
        n18346) );
  AOI22_X1 U21438 ( .A1(P3_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n18355), .B1(
        n18446), .B2(n18376), .ZN(n18345) );
  OAI211_X1 U21439 ( .C1(n18449), .C2(n18436), .A(n18346), .B(n18345), .ZN(
        P3_U2967) );
  AOI22_X1 U21440 ( .A1(n18452), .A2(n18376), .B1(n18450), .B2(n18354), .ZN(
        n18348) );
  AOI22_X1 U21441 ( .A1(P3_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n18355), .B1(
        n18399), .B2(n9602), .ZN(n18347) );
  OAI211_X1 U21442 ( .C1(n18402), .C2(n18358), .A(n18348), .B(n18347), .ZN(
        P3_U2968) );
  AOI22_X1 U21443 ( .A1(n18457), .A2(n18351), .B1(n18456), .B2(n18354), .ZN(
        n18350) );
  AOI22_X1 U21444 ( .A1(P3_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n18355), .B1(
        n18458), .B2(n18376), .ZN(n18349) );
  OAI211_X1 U21445 ( .C1(n18461), .C2(n18436), .A(n18350), .B(n18349), .ZN(
        P3_U2969) );
  AOI22_X1 U21446 ( .A1(n18465), .A2(n18376), .B1(n18462), .B2(n18354), .ZN(
        n18353) );
  AOI22_X1 U21447 ( .A1(P3_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n18355), .B1(
        n18463), .B2(n18351), .ZN(n18352) );
  OAI211_X1 U21448 ( .C1(n18469), .C2(n18436), .A(n18353), .B(n18352), .ZN(
        P3_U2970) );
  AOI22_X1 U21449 ( .A1(n18412), .A2(n18376), .B1(n18471), .B2(n18354), .ZN(
        n18357) );
  AOI22_X1 U21450 ( .A1(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n18355), .B1(
        n18475), .B2(n9602), .ZN(n18356) );
  OAI211_X1 U21451 ( .C1(n18418), .C2(n18358), .A(n18357), .B(n18356), .ZN(
        P3_U2971) );
  NOR2_X1 U21452 ( .A1(n18360), .A2(n18359), .ZN(n18425) );
  AOI22_X1 U21453 ( .A1(n18422), .A2(n18376), .B1(n18421), .B2(n18425), .ZN(
        n18365) );
  AOI22_X1 U21454 ( .A1(n18426), .A2(n18363), .B1(n18362), .B2(n18361), .ZN(
        n18379) );
  AOI22_X1 U21455 ( .A1(P3_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n18379), .B1(
        n18427), .B2(n18407), .ZN(n18364) );
  OAI211_X1 U21456 ( .C1(n18430), .C2(n18479), .A(n18365), .B(n18364), .ZN(
        P3_U2972) );
  AOI22_X1 U21457 ( .A1(n18391), .A2(n18376), .B1(n18432), .B2(n18425), .ZN(
        n18367) );
  AOI22_X1 U21458 ( .A1(P3_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n18379), .B1(
        n18431), .B2(n18407), .ZN(n18366) );
  OAI211_X1 U21459 ( .C1(n18394), .C2(n18479), .A(n18367), .B(n18366), .ZN(
        P3_U2973) );
  AOI22_X1 U21460 ( .A1(n18440), .A2(n18407), .B1(n18438), .B2(n18425), .ZN(
        n18369) );
  AOI22_X1 U21461 ( .A1(P3_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n18379), .B1(
        n18439), .B2(n18376), .ZN(n18368) );
  OAI211_X1 U21462 ( .C1(n18443), .C2(n18479), .A(n18369), .B(n18368), .ZN(
        P3_U2974) );
  AOI22_X1 U21463 ( .A1(n18445), .A2(n18376), .B1(n18444), .B2(n18425), .ZN(
        n18371) );
  AOI22_X1 U21464 ( .A1(P3_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n18379), .B1(
        n18446), .B2(n18407), .ZN(n18370) );
  OAI211_X1 U21465 ( .C1(n18449), .C2(n18479), .A(n18371), .B(n18370), .ZN(
        P3_U2975) );
  AOI22_X1 U21466 ( .A1(n18452), .A2(n18407), .B1(n18450), .B2(n18425), .ZN(
        n18373) );
  AOI22_X1 U21467 ( .A1(P3_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n18379), .B1(
        n18399), .B2(n18464), .ZN(n18372) );
  OAI211_X1 U21468 ( .C1(n18402), .C2(n18382), .A(n18373), .B(n18372), .ZN(
        P3_U2976) );
  AOI22_X1 U21469 ( .A1(n18457), .A2(n18376), .B1(n18456), .B2(n18425), .ZN(
        n18375) );
  AOI22_X1 U21470 ( .A1(P3_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n18379), .B1(
        n18458), .B2(n18407), .ZN(n18374) );
  OAI211_X1 U21471 ( .C1(n18461), .C2(n18479), .A(n18375), .B(n18374), .ZN(
        P3_U2977) );
  AOI22_X1 U21472 ( .A1(n18463), .A2(n18376), .B1(n18462), .B2(n18425), .ZN(
        n18378) );
  AOI22_X1 U21473 ( .A1(P3_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n18379), .B1(
        n18465), .B2(n18407), .ZN(n18377) );
  OAI211_X1 U21474 ( .C1(n18469), .C2(n18479), .A(n18378), .B(n18377), .ZN(
        P3_U2978) );
  AOI22_X1 U21475 ( .A1(n18412), .A2(n18407), .B1(n18471), .B2(n18425), .ZN(
        n18381) );
  AOI22_X1 U21476 ( .A1(P3_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n18379), .B1(
        n18475), .B2(n18464), .ZN(n18380) );
  OAI211_X1 U21477 ( .C1(n18418), .C2(n18382), .A(n18381), .B(n18380), .ZN(
        P3_U2979) );
  INV_X1 U21478 ( .A(n18383), .ZN(n18384) );
  NOR2_X1 U21479 ( .A1(n18420), .A2(n18384), .ZN(n18411) );
  AOI22_X1 U21480 ( .A1(n18422), .A2(n18407), .B1(n18421), .B2(n18411), .ZN(
        n18390) );
  NOR2_X1 U21481 ( .A1(n9602), .A2(n18407), .ZN(n18386) );
  OAI21_X1 U21482 ( .B1(n18386), .B2(n18385), .A(n18384), .ZN(n18387) );
  OAI211_X1 U21483 ( .C1(n18413), .C2(n18639), .A(n18388), .B(n18387), .ZN(
        n18414) );
  AOI22_X1 U21484 ( .A1(P3_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n18414), .B1(
        n18427), .B2(n9602), .ZN(n18389) );
  OAI211_X1 U21485 ( .C1(n18430), .C2(n18410), .A(n18390), .B(n18389), .ZN(
        P3_U2980) );
  AOI22_X1 U21486 ( .A1(n18391), .A2(n18407), .B1(n18432), .B2(n18411), .ZN(
        n18393) );
  AOI22_X1 U21487 ( .A1(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n18414), .B1(
        n18431), .B2(n9602), .ZN(n18392) );
  OAI211_X1 U21488 ( .C1(n18394), .C2(n18410), .A(n18393), .B(n18392), .ZN(
        P3_U2981) );
  AOI22_X1 U21489 ( .A1(n18440), .A2(n9602), .B1(n18438), .B2(n18411), .ZN(
        n18396) );
  AOI22_X1 U21490 ( .A1(P3_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n18414), .B1(
        n18439), .B2(n18407), .ZN(n18395) );
  OAI211_X1 U21491 ( .C1(n18443), .C2(n18410), .A(n18396), .B(n18395), .ZN(
        P3_U2982) );
  AOI22_X1 U21492 ( .A1(n18445), .A2(n18407), .B1(n18444), .B2(n18411), .ZN(
        n18398) );
  AOI22_X1 U21493 ( .A1(P3_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n18414), .B1(
        n18446), .B2(n9602), .ZN(n18397) );
  OAI211_X1 U21494 ( .C1(n18449), .C2(n18410), .A(n18398), .B(n18397), .ZN(
        P3_U2983) );
  AOI22_X1 U21495 ( .A1(n18452), .A2(n9602), .B1(n18450), .B2(n18411), .ZN(
        n18401) );
  AOI22_X1 U21496 ( .A1(P3_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n18414), .B1(
        n18399), .B2(n18413), .ZN(n18400) );
  OAI211_X1 U21497 ( .C1(n18402), .C2(n18417), .A(n18401), .B(n18400), .ZN(
        P3_U2984) );
  AOI22_X1 U21498 ( .A1(n18456), .A2(n18411), .B1(n18458), .B2(n9602), .ZN(
        n18405) );
  AOI22_X1 U21499 ( .A1(P3_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n18414), .B1(
        n18403), .B2(n18413), .ZN(n18404) );
  OAI211_X1 U21500 ( .C1(n18406), .C2(n18417), .A(n18405), .B(n18404), .ZN(
        P3_U2985) );
  AOI22_X1 U21501 ( .A1(n18463), .A2(n18407), .B1(n18462), .B2(n18411), .ZN(
        n18409) );
  AOI22_X1 U21502 ( .A1(P3_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n18414), .B1(
        n18465), .B2(n9602), .ZN(n18408) );
  OAI211_X1 U21503 ( .C1(n18469), .C2(n18410), .A(n18409), .B(n18408), .ZN(
        P3_U2986) );
  AOI22_X1 U21504 ( .A1(n18412), .A2(n9602), .B1(n18471), .B2(n18411), .ZN(
        n18416) );
  AOI22_X1 U21505 ( .A1(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n18414), .B1(
        n18475), .B2(n18413), .ZN(n18415) );
  OAI211_X1 U21506 ( .C1(n18418), .C2(n18417), .A(n18416), .B(n18415), .ZN(
        P3_U2987) );
  NOR2_X1 U21507 ( .A1(n18420), .A2(n18419), .ZN(n18470) );
  AOI22_X1 U21508 ( .A1(n18422), .A2(n9602), .B1(n18421), .B2(n18470), .ZN(
        n18429) );
  AOI22_X1 U21509 ( .A1(n18426), .A2(n18425), .B1(n18424), .B2(n18423), .ZN(
        n18476) );
  AOI22_X1 U21510 ( .A1(P3_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n18476), .B1(
        n18427), .B2(n18464), .ZN(n18428) );
  OAI211_X1 U21511 ( .C1(n18430), .C2(n18468), .A(n18429), .B(n18428), .ZN(
        P3_U2988) );
  AOI22_X1 U21512 ( .A1(n18432), .A2(n18470), .B1(n18431), .B2(n18464), .ZN(
        n18435) );
  AOI22_X1 U21513 ( .A1(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n18476), .B1(
        n18433), .B2(n18474), .ZN(n18434) );
  OAI211_X1 U21514 ( .C1(n18437), .C2(n18436), .A(n18435), .B(n18434), .ZN(
        P3_U2989) );
  AOI22_X1 U21515 ( .A1(n18439), .A2(n9602), .B1(n18438), .B2(n18470), .ZN(
        n18442) );
  AOI22_X1 U21516 ( .A1(P3_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n18476), .B1(
        n18440), .B2(n18464), .ZN(n18441) );
  OAI211_X1 U21517 ( .C1(n18443), .C2(n18468), .A(n18442), .B(n18441), .ZN(
        P3_U2990) );
  AOI22_X1 U21518 ( .A1(n18445), .A2(n9602), .B1(n18444), .B2(n18470), .ZN(
        n18448) );
  AOI22_X1 U21519 ( .A1(P3_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n18476), .B1(
        n18446), .B2(n18464), .ZN(n18447) );
  OAI211_X1 U21520 ( .C1(n18449), .C2(n18468), .A(n18448), .B(n18447), .ZN(
        P3_U2991) );
  AOI22_X1 U21521 ( .A1(n18451), .A2(n9602), .B1(n18450), .B2(n18470), .ZN(
        n18454) );
  AOI22_X1 U21522 ( .A1(P3_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n18476), .B1(
        n18452), .B2(n18464), .ZN(n18453) );
  OAI211_X1 U21523 ( .C1(n18455), .C2(n18468), .A(n18454), .B(n18453), .ZN(
        P3_U2992) );
  AOI22_X1 U21524 ( .A1(n18457), .A2(n9602), .B1(n18456), .B2(n18470), .ZN(
        n18460) );
  AOI22_X1 U21525 ( .A1(P3_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n18476), .B1(
        n18458), .B2(n18464), .ZN(n18459) );
  OAI211_X1 U21526 ( .C1(n18461), .C2(n18468), .A(n18460), .B(n18459), .ZN(
        P3_U2993) );
  AOI22_X1 U21527 ( .A1(n18463), .A2(n9602), .B1(n18462), .B2(n18470), .ZN(
        n18467) );
  AOI22_X1 U21528 ( .A1(P3_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n18476), .B1(
        n18465), .B2(n18464), .ZN(n18466) );
  OAI211_X1 U21529 ( .C1(n18469), .C2(n18468), .A(n18467), .B(n18466), .ZN(
        P3_U2994) );
  AOI22_X1 U21530 ( .A1(n18473), .A2(n9602), .B1(n18471), .B2(n18470), .ZN(
        n18478) );
  AOI22_X1 U21531 ( .A1(P3_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n18476), .B1(
        n18475), .B2(n18474), .ZN(n18477) );
  OAI211_X1 U21532 ( .C1(n18480), .C2(n18479), .A(n18478), .B(n18477), .ZN(
        P3_U2995) );
  INV_X1 U21533 ( .A(n18481), .ZN(n18535) );
  AOI21_X1 U21534 ( .B1(n18484), .B2(n18483), .A(n18482), .ZN(n18488) );
  AOI21_X1 U21535 ( .B1(n18509), .B2(n18486), .A(n18485), .ZN(n18487) );
  AOI211_X1 U21536 ( .C1(n18490), .C2(n18489), .A(n18488), .B(n18487), .ZN(
        n18683) );
  AOI211_X1 U21537 ( .C1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .C2(n18520), .A(
        n18492), .B(n18491), .ZN(n18533) );
  OAI21_X1 U21538 ( .B1(n18495), .B2(n18494), .A(n18493), .ZN(n18503) );
  AOI22_X1 U21539 ( .A1(n18499), .A2(n18505), .B1(n18503), .B2(n18496), .ZN(
        n18497) );
  NAND2_X1 U21540 ( .A1(n13943), .A2(n18504), .ZN(n18498) );
  NAND2_X1 U21541 ( .A1(n18497), .A2(n18498), .ZN(n18646) );
  NOR2_X1 U21542 ( .A1(n18520), .A2(n18646), .ZN(n18502) );
  INV_X1 U21543 ( .A(n18498), .ZN(n18500) );
  AOI21_X1 U21544 ( .B1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n18510), .A(
        n18499), .ZN(n18513) );
  OAI22_X1 U21545 ( .A1(n18500), .A2(n18509), .B1(n18513), .B2(n18505), .ZN(
        n18643) );
  NAND2_X1 U21546 ( .A1(n18647), .A2(n18643), .ZN(n18501) );
  OAI22_X1 U21547 ( .A1(n18502), .A2(n18647), .B1(n18520), .B2(n18501), .ZN(
        n18529) );
  NAND3_X1 U21548 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n18504), .A3(
        n18503), .ZN(n18508) );
  INV_X1 U21549 ( .A(n18513), .ZN(n18506) );
  OAI211_X1 U21550 ( .C1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .C2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(n18506), .B(n18505), .ZN(
        n18507) );
  OAI211_X1 U21551 ( .C1(n18653), .C2(n18509), .A(n18508), .B(n18507), .ZN(
        n18654) );
  MUX2_X1 U21552 ( .A(n18654), .B(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .S(
        n18520), .Z(n18523) );
  NOR2_X1 U21553 ( .A1(n18511), .A2(n18510), .ZN(n18514) );
  AOI22_X1 U21554 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18512), .B1(
        n18514), .B2(n18668), .ZN(n18664) );
  OAI22_X1 U21555 ( .A1(n18514), .A2(n18656), .B1(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n18513), .ZN(n18661) );
  OR3_X1 U21556 ( .A1(n18664), .A2(n18517), .A3(n18515), .ZN(n18516) );
  AOI22_X1 U21557 ( .A1(n18664), .A2(n18517), .B1(n18661), .B2(n18516), .ZN(
        n18519) );
  OAI21_X1 U21558 ( .B1(n18520), .B2(n18519), .A(n18518), .ZN(n18521) );
  OAI21_X1 U21559 ( .B1(n18523), .B2(n18522), .A(n18521), .ZN(n18524) );
  INV_X1 U21560 ( .A(n18523), .ZN(n18525) );
  OAI221_X1 U21561 ( .B1(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .C1(
        P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .C2(n18524), .A(n18525), .ZN(
        n18528) );
  NOR2_X1 U21562 ( .A1(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n18527) );
  OAI21_X1 U21563 ( .B1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n18525), .A(
        n18524), .ZN(n18526) );
  AOI22_X1 U21564 ( .A1(n18529), .A2(n18528), .B1(n18527), .B2(n18526), .ZN(
        n18532) );
  OAI21_X1 U21565 ( .B1(P3_MORE_REG_SCAN_IN), .B2(P3_FLUSH_REG_SCAN_IN), .A(
        n18530), .ZN(n18531) );
  NAND4_X1 U21566 ( .A1(n18683), .A2(n18533), .A3(n18532), .A4(n18531), .ZN(
        n18539) );
  AOI211_X1 U21567 ( .C1(n18536), .C2(n18535), .A(n18534), .B(n18539), .ZN(
        n18637) );
  AOI21_X1 U21568 ( .B1(n18688), .B2(n18704), .A(n18637), .ZN(n18545) );
  NOR2_X1 U21569 ( .A1(n18693), .A2(n18687), .ZN(n18542) );
  AOI211_X1 U21570 ( .C1(n18663), .C2(n18696), .A(P3_STATE2_REG_0__SCAN_IN), 
        .B(n18542), .ZN(n18537) );
  AOI211_X1 U21571 ( .C1(n18686), .C2(n18539), .A(n18538), .B(n18537), .ZN(
        n18540) );
  OAI221_X1 U21572 ( .B1(n18636), .B2(n18545), .C1(n18636), .C2(n18541), .A(
        n18540), .ZN(P3_U2996) );
  INV_X1 U21573 ( .A(n18542), .ZN(n18548) );
  NAND4_X1 U21574 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(
        P3_STATE2_REG_1__SCAN_IN), .A3(n18688), .A4(n18704), .ZN(n18551) );
  INV_X1 U21575 ( .A(n18543), .ZN(n18546) );
  NAND3_X1 U21576 ( .A1(n18546), .A2(n18545), .A3(n18544), .ZN(n18547) );
  NAND4_X1 U21577 ( .A1(n18549), .A2(n18548), .A3(n18551), .A4(n18547), .ZN(
        P3_U2997) );
  OAI21_X1 U21578 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(
        P3_STATEBS16_REG_SCAN_IN), .A(n18550), .ZN(n18553) );
  INV_X1 U21579 ( .A(n18551), .ZN(n18552) );
  AOI21_X1 U21580 ( .B1(n18554), .B2(n18553), .A(n18552), .ZN(P3_U2998) );
  AND2_X1 U21581 ( .A1(P3_DATAWIDTH_REG_31__SCAN_IN), .A2(n18633), .ZN(
        P3_U2999) );
  AND2_X1 U21582 ( .A1(P3_DATAWIDTH_REG_30__SCAN_IN), .A2(n18633), .ZN(
        P3_U3000) );
  AND2_X1 U21583 ( .A1(P3_DATAWIDTH_REG_29__SCAN_IN), .A2(n18633), .ZN(
        P3_U3001) );
  AND2_X1 U21584 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(n18633), .ZN(
        P3_U3002) );
  AND2_X1 U21585 ( .A1(P3_DATAWIDTH_REG_27__SCAN_IN), .A2(n18633), .ZN(
        P3_U3003) );
  AND2_X1 U21586 ( .A1(P3_DATAWIDTH_REG_26__SCAN_IN), .A2(n18633), .ZN(
        P3_U3004) );
  AND2_X1 U21587 ( .A1(P3_DATAWIDTH_REG_25__SCAN_IN), .A2(n18633), .ZN(
        P3_U3005) );
  AND2_X1 U21588 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(n18633), .ZN(
        P3_U3006) );
  AND2_X1 U21589 ( .A1(P3_DATAWIDTH_REG_23__SCAN_IN), .A2(n18633), .ZN(
        P3_U3007) );
  AND2_X1 U21590 ( .A1(P3_DATAWIDTH_REG_22__SCAN_IN), .A2(n18633), .ZN(
        P3_U3008) );
  AND2_X1 U21591 ( .A1(P3_DATAWIDTH_REG_21__SCAN_IN), .A2(n18633), .ZN(
        P3_U3009) );
  AND2_X1 U21592 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(n18633), .ZN(
        P3_U3010) );
  AND2_X1 U21593 ( .A1(P3_DATAWIDTH_REG_19__SCAN_IN), .A2(n18633), .ZN(
        P3_U3011) );
  AND2_X1 U21594 ( .A1(P3_DATAWIDTH_REG_18__SCAN_IN), .A2(n18633), .ZN(
        P3_U3012) );
  AND2_X1 U21595 ( .A1(P3_DATAWIDTH_REG_17__SCAN_IN), .A2(n18633), .ZN(
        P3_U3013) );
  AND2_X1 U21596 ( .A1(P3_DATAWIDTH_REG_16__SCAN_IN), .A2(n18633), .ZN(
        P3_U3014) );
  AND2_X1 U21597 ( .A1(P3_DATAWIDTH_REG_15__SCAN_IN), .A2(n18633), .ZN(
        P3_U3015) );
  AND2_X1 U21598 ( .A1(P3_DATAWIDTH_REG_14__SCAN_IN), .A2(n18633), .ZN(
        P3_U3016) );
  AND2_X1 U21599 ( .A1(P3_DATAWIDTH_REG_13__SCAN_IN), .A2(n18633), .ZN(
        P3_U3017) );
  AND2_X1 U21600 ( .A1(P3_DATAWIDTH_REG_12__SCAN_IN), .A2(n18633), .ZN(
        P3_U3018) );
  AND2_X1 U21601 ( .A1(P3_DATAWIDTH_REG_11__SCAN_IN), .A2(n18633), .ZN(
        P3_U3019) );
  AND2_X1 U21602 ( .A1(P3_DATAWIDTH_REG_10__SCAN_IN), .A2(n18633), .ZN(
        P3_U3020) );
  AND2_X1 U21603 ( .A1(P3_DATAWIDTH_REG_9__SCAN_IN), .A2(n18633), .ZN(P3_U3021) );
  AND2_X1 U21604 ( .A1(P3_DATAWIDTH_REG_8__SCAN_IN), .A2(n18633), .ZN(P3_U3022) );
  AND2_X1 U21605 ( .A1(P3_DATAWIDTH_REG_7__SCAN_IN), .A2(n18633), .ZN(P3_U3023) );
  INV_X1 U21606 ( .A(P3_DATAWIDTH_REG_6__SCAN_IN), .ZN(n20895) );
  NOR2_X1 U21607 ( .A1(n20895), .A2(n18635), .ZN(P3_U3024) );
  AND2_X1 U21608 ( .A1(P3_DATAWIDTH_REG_5__SCAN_IN), .A2(n18633), .ZN(P3_U3025) );
  AND2_X1 U21609 ( .A1(P3_DATAWIDTH_REG_4__SCAN_IN), .A2(n18633), .ZN(P3_U3026) );
  AND2_X1 U21610 ( .A1(P3_DATAWIDTH_REG_3__SCAN_IN), .A2(n18633), .ZN(P3_U3027) );
  AND2_X1 U21611 ( .A1(P3_DATAWIDTH_REG_2__SCAN_IN), .A2(n18633), .ZN(P3_U3028) );
  NOR2_X1 U21612 ( .A1(n18570), .A2(n20601), .ZN(n18565) );
  INV_X1 U21613 ( .A(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n18558) );
  AOI211_X1 U21614 ( .C1(P3_STATE_REG_1__SCAN_IN), .C2(HOLD), .A(n18565), .B(
        n18558), .ZN(n18557) );
  NAND2_X1 U21615 ( .A1(n18688), .A2(P3_STATE_REG_1__SCAN_IN), .ZN(n18563) );
  AND2_X1 U21616 ( .A1(n18563), .A2(P3_STATE_REG_0__SCAN_IN), .ZN(n18569) );
  INV_X1 U21617 ( .A(NA), .ZN(n20612) );
  OAI21_X1 U21618 ( .B1(n20612), .B2(n18555), .A(P3_STATE_REG_2__SCAN_IN), 
        .ZN(n18568) );
  INV_X1 U21619 ( .A(n18568), .ZN(n18556) );
  OAI22_X1 U21620 ( .A1(n18703), .A2(n18557), .B1(n18569), .B2(n18556), .ZN(
        P3_U3029) );
  NOR2_X1 U21621 ( .A1(n18565), .A2(n18558), .ZN(n18561) );
  NOR2_X1 U21622 ( .A1(n18559), .A2(n20601), .ZN(n18560) );
  AOI22_X1 U21623 ( .A1(P3_STATE_REG_0__SCAN_IN), .A2(n18561), .B1(n18560), 
        .B2(n18570), .ZN(n18562) );
  NAND3_X1 U21624 ( .A1(n18562), .A2(n18690), .A3(n18563), .ZN(P3_U3030) );
  OAI22_X1 U21625 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(
        P3_REQUESTPENDING_REG_SCAN_IN), .B1(NA), .B2(n18563), .ZN(n18564) );
  OAI22_X1 U21626 ( .A1(n18565), .A2(n18564), .B1(
        P3_REQUESTPENDING_REG_SCAN_IN), .B2(HOLD), .ZN(n18566) );
  OAI22_X1 U21627 ( .A1(n18569), .A2(n18568), .B1(n18567), .B2(n18566), .ZN(
        P3_U3031) );
  OAI222_X1 U21628 ( .A1(n18679), .A2(n18631), .B1(n18571), .B2(n18703), .C1(
        n18572), .C2(n18622), .ZN(P3_U3032) );
  INV_X1 U21629 ( .A(P3_REIP_REG_3__SCAN_IN), .ZN(n18574) );
  OAI222_X1 U21630 ( .A1(n18622), .A2(n18574), .B1(n18573), .B2(n18703), .C1(
        n18572), .C2(n18631), .ZN(P3_U3033) );
  OAI222_X1 U21631 ( .A1(n18622), .A2(n18576), .B1(n18575), .B2(n18703), .C1(
        n18574), .C2(n18631), .ZN(P3_U3034) );
  OAI222_X1 U21632 ( .A1(n18622), .A2(n18578), .B1(n18577), .B2(n18703), .C1(
        n18576), .C2(n18631), .ZN(P3_U3035) );
  OAI222_X1 U21633 ( .A1(n18622), .A2(n18580), .B1(n18579), .B2(n18703), .C1(
        n18578), .C2(n18631), .ZN(P3_U3036) );
  OAI222_X1 U21634 ( .A1(n18622), .A2(n18582), .B1(n18581), .B2(n18703), .C1(
        n18580), .C2(n18631), .ZN(P3_U3037) );
  INV_X1 U21635 ( .A(P3_REIP_REG_8__SCAN_IN), .ZN(n18585) );
  OAI222_X1 U21636 ( .A1(n18622), .A2(n18585), .B1(n18583), .B2(n18703), .C1(
        n18582), .C2(n18631), .ZN(P3_U3038) );
  OAI222_X1 U21637 ( .A1(n18585), .A2(n18631), .B1(n18584), .B2(n18703), .C1(
        n18586), .C2(n18622), .ZN(P3_U3039) );
  OAI222_X1 U21638 ( .A1(n18622), .A2(n18588), .B1(n18587), .B2(n18703), .C1(
        n18586), .C2(n18631), .ZN(P3_U3040) );
  OAI222_X1 U21639 ( .A1(n18622), .A2(n18590), .B1(n18589), .B2(n18703), .C1(
        n18588), .C2(n18631), .ZN(P3_U3041) );
  OAI222_X1 U21640 ( .A1(n18622), .A2(n18592), .B1(n18591), .B2(n18703), .C1(
        n18590), .C2(n18631), .ZN(P3_U3042) );
  OAI222_X1 U21641 ( .A1(n18622), .A2(n18594), .B1(n18593), .B2(n18703), .C1(
        n18592), .C2(n18631), .ZN(P3_U3043) );
  OAI222_X1 U21642 ( .A1(n18622), .A2(n18597), .B1(n18595), .B2(n18703), .C1(
        n18594), .C2(n18631), .ZN(P3_U3044) );
  OAI222_X1 U21643 ( .A1(n18597), .A2(n18631), .B1(n18596), .B2(n18703), .C1(
        n18598), .C2(n18622), .ZN(P3_U3045) );
  OAI222_X1 U21644 ( .A1(n18622), .A2(n18600), .B1(n18599), .B2(n18703), .C1(
        n18598), .C2(n18631), .ZN(P3_U3046) );
  OAI222_X1 U21645 ( .A1(n18622), .A2(n18602), .B1(n18601), .B2(n18703), .C1(
        n18600), .C2(n18631), .ZN(P3_U3047) );
  OAI222_X1 U21646 ( .A1(n18622), .A2(n18604), .B1(n18603), .B2(n18703), .C1(
        n18602), .C2(n18631), .ZN(P3_U3048) );
  OAI222_X1 U21647 ( .A1(n18622), .A2(n18607), .B1(n18605), .B2(n18703), .C1(
        n18604), .C2(n18631), .ZN(P3_U3049) );
  INV_X1 U21648 ( .A(P3_REIP_REG_20__SCAN_IN), .ZN(n18608) );
  OAI222_X1 U21649 ( .A1(n18607), .A2(n18631), .B1(n18606), .B2(n18703), .C1(
        n18608), .C2(n18622), .ZN(P3_U3050) );
  OAI222_X1 U21650 ( .A1(n18622), .A2(n18611), .B1(n18609), .B2(n18703), .C1(
        n18608), .C2(n18631), .ZN(P3_U3051) );
  OAI222_X1 U21651 ( .A1(n18611), .A2(n18631), .B1(n18610), .B2(n18703), .C1(
        n18612), .C2(n18622), .ZN(P3_U3052) );
  OAI222_X1 U21652 ( .A1(n18622), .A2(n18615), .B1(n18613), .B2(n18703), .C1(
        n18612), .C2(n18631), .ZN(P3_U3053) );
  INV_X1 U21653 ( .A(P3_REIP_REG_24__SCAN_IN), .ZN(n18616) );
  OAI222_X1 U21654 ( .A1(n18615), .A2(n18631), .B1(n18614), .B2(n18703), .C1(
        n18616), .C2(n18622), .ZN(P3_U3054) );
  OAI222_X1 U21655 ( .A1(n18622), .A2(n18618), .B1(n18617), .B2(n18703), .C1(
        n18616), .C2(n18631), .ZN(P3_U3055) );
  OAI222_X1 U21656 ( .A1(n18622), .A2(n18620), .B1(n18619), .B2(n18703), .C1(
        n18618), .C2(n18631), .ZN(P3_U3056) );
  OAI222_X1 U21657 ( .A1(n18622), .A2(n18623), .B1(n18621), .B2(n18703), .C1(
        n18620), .C2(n18631), .ZN(P3_U3057) );
  INV_X1 U21658 ( .A(P3_REIP_REG_28__SCAN_IN), .ZN(n18626) );
  OAI222_X1 U21659 ( .A1(n18622), .A2(n18626), .B1(n18624), .B2(n18703), .C1(
        n18623), .C2(n18631), .ZN(P3_U3058) );
  OAI222_X1 U21660 ( .A1(n18626), .A2(n18631), .B1(n18625), .B2(n18703), .C1(
        n20840), .C2(n18622), .ZN(P3_U3059) );
  OAI222_X1 U21661 ( .A1(n20840), .A2(n18631), .B1(n18627), .B2(n18703), .C1(
        n18630), .C2(n18622), .ZN(P3_U3060) );
  OAI222_X1 U21662 ( .A1(n18631), .A2(n18630), .B1(n18629), .B2(n18703), .C1(
        n18628), .C2(n18622), .ZN(P3_U3061) );
  MUX2_X1 U21663 ( .A(P3_BE_N_REG_3__SCAN_IN), .B(P3_BYTEENABLE_REG_3__SCAN_IN), .S(n18703), .Z(P3_U3274) );
  MUX2_X1 U21664 ( .A(P3_BE_N_REG_2__SCAN_IN), .B(P3_BYTEENABLE_REG_2__SCAN_IN), .S(n18703), .Z(P3_U3275) );
  MUX2_X1 U21665 ( .A(P3_BE_N_REG_1__SCAN_IN), .B(P3_BYTEENABLE_REG_1__SCAN_IN), .S(n18703), .Z(P3_U3276) );
  MUX2_X1 U21666 ( .A(P3_BE_N_REG_0__SCAN_IN), .B(P3_BYTEENABLE_REG_0__SCAN_IN), .S(n18703), .Z(P3_U3277) );
  INV_X1 U21667 ( .A(n18634), .ZN(n18632) );
  AOI21_X1 U21668 ( .B1(n18633), .B2(n20823), .A(n18632), .ZN(P3_U3280) );
  OAI21_X1 U21669 ( .B1(n18635), .B2(n18671), .A(n18634), .ZN(P3_U3281) );
  NOR2_X1 U21670 ( .A1(n18637), .A2(n18636), .ZN(n18640) );
  OAI21_X1 U21671 ( .B1(n18640), .B2(n18639), .A(n18638), .ZN(P3_U3282) );
  INV_X1 U21672 ( .A(n18641), .ZN(n18645) );
  NOR2_X1 U21673 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n18642), .ZN(
        n18644) );
  AOI22_X1 U21674 ( .A1(n18663), .A2(n18645), .B1(n18644), .B2(n18643), .ZN(
        n18649) );
  AOI21_X1 U21675 ( .B1(n18705), .B2(n18646), .A(n18669), .ZN(n18648) );
  OAI22_X1 U21676 ( .A1(n18669), .A2(n18649), .B1(n18648), .B2(n18647), .ZN(
        P3_U3285) );
  NOR2_X1 U21677 ( .A1(n18650), .A2(n18665), .ZN(n18658) );
  AOI22_X1 U21678 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(n18652), .B2(n18651), .ZN(
        n18657) );
  AOI222_X1 U21679 ( .A1(n18654), .A2(n18705), .B1(n18658), .B2(n18657), .C1(
        n18663), .C2(n18653), .ZN(n18655) );
  AOI22_X1 U21680 ( .A1(n18669), .A2(n13943), .B1(n18655), .B2(n18666), .ZN(
        P3_U3288) );
  INV_X1 U21681 ( .A(n18656), .ZN(n18660) );
  INV_X1 U21682 ( .A(n18657), .ZN(n18659) );
  AOI222_X1 U21683 ( .A1(n18661), .A2(n18705), .B1(n18663), .B2(n18660), .C1(
        n18659), .C2(n18658), .ZN(n18662) );
  AOI22_X1 U21684 ( .A1(n18669), .A2(n13853), .B1(n18662), .B2(n18666), .ZN(
        P3_U3289) );
  AOI222_X1 U21685 ( .A1(n18665), .A2(P3_STATE2_REG_1__SCAN_IN), .B1(n18705), 
        .B2(n18664), .C1(n18668), .C2(n18663), .ZN(n18667) );
  AOI22_X1 U21686 ( .A1(n18669), .A2(n18668), .B1(n18667), .B2(n18666), .ZN(
        P3_U3290) );
  AOI221_X1 U21687 ( .B1(P3_DATAWIDTH_REG_0__SCAN_IN), .B2(n18672), .C1(n20823), .C2(n18671), .A(n18670), .ZN(n18674) );
  OAI22_X1 U21688 ( .A1(n18676), .A2(P3_BYTEENABLE_REG_2__SCAN_IN), .B1(n18679), .B2(n18675), .ZN(n18673) );
  NOR2_X1 U21689 ( .A1(n18674), .A2(n18673), .ZN(P3_U3292) );
  OAI21_X1 U21690 ( .B1(n18676), .B2(P3_BYTEENABLE_REG_0__SCAN_IN), .A(n18675), 
        .ZN(n18677) );
  OAI21_X1 U21691 ( .B1(n18679), .B2(n18678), .A(n18677), .ZN(P3_U3293) );
  INV_X1 U21692 ( .A(P3_W_R_N_REG_SCAN_IN), .ZN(n18680) );
  AOI22_X1 U21693 ( .A1(n18703), .A2(P3_READREQUEST_REG_SCAN_IN), .B1(n18680), 
        .B2(n18701), .ZN(P3_U3294) );
  INV_X1 U21694 ( .A(n18681), .ZN(n18684) );
  NAND2_X1 U21695 ( .A1(n18684), .A2(P3_MORE_REG_SCAN_IN), .ZN(n18682) );
  OAI21_X1 U21696 ( .B1(n18684), .B2(n18683), .A(n18682), .ZN(P3_U3295) );
  OAI22_X1 U21697 ( .A1(n18688), .A2(n18687), .B1(n18686), .B2(n18685), .ZN(
        n18689) );
  NOR2_X1 U21698 ( .A1(n18707), .A2(n18689), .ZN(n18700) );
  AOI21_X1 U21699 ( .B1(n18692), .B2(n18691), .A(n18690), .ZN(n18694) );
  OAI211_X1 U21700 ( .C1(n18695), .C2(n18694), .A(P3_STATE2_REG_2__SCAN_IN), 
        .B(n18693), .ZN(n18697) );
  AOI21_X1 U21701 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(n18697), .A(n18696), 
        .ZN(n18699) );
  NAND2_X1 U21702 ( .A1(n18700), .A2(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(
        n18698) );
  OAI21_X1 U21703 ( .B1(n18700), .B2(n18699), .A(n18698), .ZN(P3_U3296) );
  INV_X1 U21704 ( .A(P3_MEMORYFETCH_REG_SCAN_IN), .ZN(n18710) );
  INV_X1 U21705 ( .A(P3_M_IO_N_REG_SCAN_IN), .ZN(n18702) );
  AOI22_X1 U21706 ( .A1(n18703), .A2(n18710), .B1(n18702), .B2(n18701), .ZN(
        P3_U3297) );
  AOI21_X1 U21707 ( .B1(n18705), .B2(n18704), .A(n18707), .ZN(n18711) );
  INV_X1 U21708 ( .A(P3_READREQUEST_REG_SCAN_IN), .ZN(n18708) );
  AOI22_X1 U21709 ( .A1(n18711), .A2(n18708), .B1(n18707), .B2(n18706), .ZN(
        P3_U3298) );
  AOI21_X1 U21710 ( .B1(n18711), .B2(n18710), .A(n18709), .ZN(P3_U3299) );
  INV_X1 U21711 ( .A(P2_STATE_REG_0__SCAN_IN), .ZN(n18713) );
  INV_X1 U21712 ( .A(P2_ADS_N_REG_SCAN_IN), .ZN(n18712) );
  INV_X1 U21713 ( .A(P2_STATE_REG_2__SCAN_IN), .ZN(n19683) );
  NAND2_X1 U21714 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(n19683), .ZN(n19673) );
  AOI22_X1 U21715 ( .A1(P2_STATE_REG_0__SCAN_IN), .A2(n19673), .B1(
        P2_STATE_REG_1__SCAN_IN), .B2(n18713), .ZN(n19746) );
  INV_X1 U21716 ( .A(n19746), .ZN(n19666) );
  OAI21_X1 U21717 ( .B1(n18713), .B2(n18712), .A(n19666), .ZN(P2_U2815) );
  INV_X1 U21718 ( .A(P2_CODEFETCH_REG_SCAN_IN), .ZN(n18716) );
  OAI22_X1 U21719 ( .A1(n19804), .A2(n18716), .B1(n18715), .B2(n18714), .ZN(
        P2_U2816) );
  INV_X1 U21720 ( .A(n19667), .ZN(n19678) );
  INV_X1 U21721 ( .A(P2_STATE_REG_1__SCAN_IN), .ZN(n19674) );
  OR2_X1 U21722 ( .A1(P2_STATE_REG_0__SCAN_IN), .A2(n19674), .ZN(n19812) );
  INV_X2 U21723 ( .A(n19812), .ZN(n19815) );
  AOI22_X1 U21724 ( .A1(n19815), .A2(n18716), .B1(P2_D_C_N_REG_SCAN_IN), .B2(
        n19812), .ZN(n18717) );
  OAI21_X1 U21725 ( .B1(P2_STATE_REG_0__SCAN_IN), .B2(n19678), .A(n18717), 
        .ZN(P2_U2817) );
  OAI21_X1 U21726 ( .B1(n19667), .B2(BS16), .A(n19746), .ZN(n19744) );
  OAI21_X1 U21727 ( .B1(n19746), .B2(n19221), .A(n19744), .ZN(P2_U2818) );
  NOR4_X1 U21728 ( .A1(P2_DATAWIDTH_REG_10__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_11__SCAN_IN), .A3(P2_DATAWIDTH_REG_12__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_13__SCAN_IN), .ZN(n18727) );
  NOR4_X1 U21729 ( .A1(P2_DATAWIDTH_REG_6__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_7__SCAN_IN), .A3(P2_DATAWIDTH_REG_8__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_9__SCAN_IN), .ZN(n18726) );
  AOI211_X1 U21730 ( .C1(P2_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P2_DATAWIDTH_REG_1__SCAN_IN), .A(P2_DATAWIDTH_REG_2__SCAN_IN), .B(
        P2_DATAWIDTH_REG_4__SCAN_IN), .ZN(n18718) );
  INV_X1 U21731 ( .A(P2_DATAWIDTH_REG_20__SCAN_IN), .ZN(n20737) );
  INV_X1 U21732 ( .A(P2_DATAWIDTH_REG_3__SCAN_IN), .ZN(n20807) );
  NAND3_X1 U21733 ( .A1(n18718), .A2(n20737), .A3(n20807), .ZN(n18724) );
  NOR4_X1 U21734 ( .A1(P2_DATAWIDTH_REG_19__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_21__SCAN_IN), .A3(P2_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_23__SCAN_IN), .ZN(n18722) );
  NOR4_X1 U21735 ( .A1(P2_DATAWIDTH_REG_14__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_16__SCAN_IN), .A3(P2_DATAWIDTH_REG_17__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_18__SCAN_IN), .ZN(n18721) );
  NOR4_X1 U21736 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_29__SCAN_IN), .A3(P2_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_31__SCAN_IN), .ZN(n18720) );
  NOR4_X1 U21737 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_25__SCAN_IN), .A3(P2_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_27__SCAN_IN), .ZN(n18719) );
  NAND4_X1 U21738 ( .A1(n18722), .A2(n18721), .A3(n18720), .A4(n18719), .ZN(
        n18723) );
  NOR4_X1 U21739 ( .A1(P2_DATAWIDTH_REG_5__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_15__SCAN_IN), .A3(n18724), .A4(n18723), .ZN(n18725)
         );
  NAND3_X1 U21740 ( .A1(n18727), .A2(n18726), .A3(n18725), .ZN(n18733) );
  NOR2_X1 U21741 ( .A1(P2_REIP_REG_1__SCAN_IN), .A2(n18733), .ZN(n18728) );
  INV_X1 U21742 ( .A(P2_BYTEENABLE_REG_0__SCAN_IN), .ZN(n19742) );
  AOI22_X1 U21743 ( .A1(n18728), .A2(n11633), .B1(n18733), .B2(n19742), .ZN(
        P2_U2820) );
  OR3_X1 U21744 ( .A1(P2_REIP_REG_0__SCAN_IN), .A2(P2_DATAWIDTH_REG_1__SCAN_IN), .A3(P2_DATAWIDTH_REG_0__SCAN_IN), .ZN(n18732) );
  INV_X1 U21745 ( .A(P2_BYTEENABLE_REG_1__SCAN_IN), .ZN(n19740) );
  AOI22_X1 U21746 ( .A1(n18728), .A2(n18732), .B1(n18733), .B2(n19740), .ZN(
        P2_U2821) );
  INV_X1 U21747 ( .A(P2_DATAWIDTH_REG_1__SCAN_IN), .ZN(n19745) );
  NAND2_X1 U21748 ( .A1(n18728), .A2(n19745), .ZN(n18731) );
  INV_X1 U21749 ( .A(n18733), .ZN(n18734) );
  OAI21_X1 U21750 ( .B1(n11633), .B2(n19685), .A(n18734), .ZN(n18729) );
  OAI21_X1 U21751 ( .B1(P2_BYTEENABLE_REG_2__SCAN_IN), .B2(n18734), .A(n18729), 
        .ZN(n18730) );
  OAI221_X1 U21752 ( .B1(n18731), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .C1(n18731), .C2(P2_REIP_REG_0__SCAN_IN), .A(n18730), .ZN(P2_U2822) );
  INV_X1 U21753 ( .A(P2_BYTEENABLE_REG_3__SCAN_IN), .ZN(n19738) );
  OAI221_X1 U21754 ( .B1(n18734), .B2(n19738), .C1(n18733), .C2(n18732), .A(
        n18731), .ZN(P2_U2823) );
  INV_X1 U21755 ( .A(n18735), .ZN(n18736) );
  AOI211_X1 U21756 ( .C1(n18738), .C2(n18737), .A(n18736), .B(n18890), .ZN(
        n18739) );
  INV_X1 U21757 ( .A(n18739), .ZN(n18748) );
  OAI22_X1 U21758 ( .A1(n18740), .A2(n18923), .B1(n19717), .B2(n18932), .ZN(
        n18741) );
  INV_X1 U21759 ( .A(n18741), .ZN(n18747) );
  AOI22_X1 U21760 ( .A1(n18842), .A2(P2_EBX_REG_21__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n18892), .ZN(n18746) );
  INV_X1 U21761 ( .A(n18742), .ZN(n18744) );
  AOI22_X1 U21762 ( .A1(n18744), .A2(n18916), .B1(n18874), .B2(n18743), .ZN(
        n18745) );
  NAND4_X1 U21763 ( .A1(n18748), .A2(n18747), .A3(n18746), .A4(n18745), .ZN(
        P2_U2834) );
  AOI22_X1 U21764 ( .A1(n18749), .A2(n18896), .B1(P2_EBX_REG_20__SCAN_IN), 
        .B2(n18842), .ZN(n18759) );
  AOI22_X1 U21765 ( .A1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n18892), .B1(
        P2_REIP_REG_20__SCAN_IN), .B2(n18910), .ZN(n18758) );
  AOI22_X1 U21766 ( .A1(n18751), .A2(n18916), .B1(n18874), .B2(n18750), .ZN(
        n18757) );
  AOI21_X1 U21767 ( .B1(n18754), .B2(n18753), .A(n18752), .ZN(n18755) );
  NAND2_X1 U21768 ( .A1(n18920), .A2(n18755), .ZN(n18756) );
  NAND4_X1 U21769 ( .A1(n18759), .A2(n18758), .A3(n18757), .A4(n18756), .ZN(
        P2_U2835) );
  OAI21_X1 U21770 ( .B1(n18929), .B2(n11999), .A(n12482), .ZN(n18763) );
  INV_X1 U21771 ( .A(n18760), .ZN(n18761) );
  OAI22_X1 U21772 ( .A1(n18761), .A2(n18923), .B1(n19711), .B2(n18932), .ZN(
        n18762) );
  AOI211_X1 U21773 ( .C1(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .C2(n18892), .A(
        n18763), .B(n18762), .ZN(n18769) );
  XOR2_X1 U21774 ( .A(n18765), .B(n18764), .Z(n18767) );
  AOI22_X1 U21775 ( .A1(n18767), .A2(n18920), .B1(n18916), .B2(n18766), .ZN(
        n18768) );
  OAI211_X1 U21776 ( .C1(n18770), .C2(n18928), .A(n18769), .B(n18768), .ZN(
        P2_U2837) );
  OAI21_X1 U21777 ( .B1(n18771), .B2(n18935), .A(n12482), .ZN(n18772) );
  AOI21_X1 U21778 ( .B1(n18842), .B2(P2_EBX_REG_17__SCAN_IN), .A(n18772), .ZN(
        n18773) );
  OAI21_X1 U21779 ( .B1(n19709), .B2(n18932), .A(n18773), .ZN(n18774) );
  AOI21_X1 U21780 ( .B1(n18775), .B2(n18896), .A(n18774), .ZN(n18784) );
  OAI22_X1 U21781 ( .A1(n18777), .A2(n18928), .B1(n18924), .B2(n18776), .ZN(
        n18778) );
  INV_X1 U21782 ( .A(n18778), .ZN(n18783) );
  OAI211_X1 U21783 ( .C1(n18781), .C2(n18780), .A(n18920), .B(n18779), .ZN(
        n18782) );
  NAND3_X1 U21784 ( .A1(n18784), .A2(n18783), .A3(n18782), .ZN(P2_U2838) );
  NAND2_X1 U21785 ( .A1(n9887), .A2(n18785), .ZN(n18786) );
  XOR2_X1 U21786 ( .A(n18787), .B(n18786), .Z(n18795) );
  OAI21_X1 U21787 ( .B1(n18929), .B2(n11557), .A(n12482), .ZN(n18792) );
  INV_X1 U21788 ( .A(n18788), .ZN(n18790) );
  OAI22_X1 U21789 ( .A1(n18790), .A2(n18923), .B1(n18789), .B2(n18935), .ZN(
        n18791) );
  AOI211_X1 U21790 ( .C1(P2_REIP_REG_16__SCAN_IN), .C2(n18910), .A(n18792), 
        .B(n18791), .ZN(n18794) );
  AOI22_X1 U21791 ( .A1(n18968), .A2(n18874), .B1(n18916), .B2(n18943), .ZN(
        n18793) );
  OAI211_X1 U21792 ( .C1(n18890), .C2(n18795), .A(n18794), .B(n18793), .ZN(
        P2_U2839) );
  NOR2_X1 U21793 ( .A1(n18912), .A2(n18796), .ZN(n18797) );
  XOR2_X1 U21794 ( .A(n18798), .B(n18797), .Z(n18805) );
  OAI21_X1 U21795 ( .B1(n18929), .B2(n11421), .A(n12482), .ZN(n18801) );
  OAI22_X1 U21796 ( .A1(n18799), .A2(n18923), .B1(n11215), .B2(n18935), .ZN(
        n18800) );
  AOI211_X1 U21797 ( .C1(P2_REIP_REG_15__SCAN_IN), .C2(n18910), .A(n18801), 
        .B(n18800), .ZN(n18804) );
  AOI22_X1 U21798 ( .A1(n18972), .A2(n18874), .B1(n18916), .B2(n18802), .ZN(
        n18803) );
  OAI211_X1 U21799 ( .C1(n18890), .C2(n18805), .A(n18804), .B(n18803), .ZN(
        P2_U2840) );
  NAND2_X1 U21800 ( .A1(n9887), .A2(n18806), .ZN(n18829) );
  XOR2_X1 U21801 ( .A(n18807), .B(n18829), .Z(n18817) );
  NOR2_X1 U21802 ( .A1(n18929), .A2(n18808), .ZN(n18809) );
  AOI211_X1 U21803 ( .C1(n18892), .C2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .A(
        n18810), .B(n18809), .ZN(n18811) );
  OAI21_X1 U21804 ( .B1(n19705), .B2(n18932), .A(n18811), .ZN(n18812) );
  AOI21_X1 U21805 ( .B1(n18813), .B2(n18896), .A(n18812), .ZN(n18816) );
  AOI22_X1 U21806 ( .A1(n18975), .A2(n18874), .B1(n18916), .B2(n18814), .ZN(
        n18815) );
  OAI211_X1 U21807 ( .C1(n18890), .C2(n18817), .A(n18816), .B(n18815), .ZN(
        P2_U2841) );
  OAI21_X1 U21808 ( .B1(n18818), .B2(n18823), .A(n18920), .ZN(n18828) );
  NOR2_X1 U21809 ( .A1(n18932), .A2(n19703), .ZN(n18820) );
  OAI21_X1 U21810 ( .B1(n18929), .B2(n11552), .A(n16114), .ZN(n18819) );
  AOI211_X1 U21811 ( .C1(n18821), .C2(n18896), .A(n18820), .B(n18819), .ZN(
        n18822) );
  OAI21_X1 U21812 ( .B1(n18823), .B2(n18855), .A(n18822), .ZN(n18826) );
  OAI22_X1 U21813 ( .A1(n18979), .A2(n18928), .B1(n18924), .B2(n18824), .ZN(
        n18825) );
  AOI211_X1 U21814 ( .C1(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .C2(n18892), .A(
        n18826), .B(n18825), .ZN(n18827) );
  OAI21_X1 U21815 ( .B1(n18829), .B2(n18828), .A(n18827), .ZN(P2_U2842) );
  AND2_X1 U21816 ( .A1(n9887), .A2(n18830), .ZN(n18850) );
  XNOR2_X1 U21817 ( .A(n18832), .B(n18850), .ZN(n18841) );
  NAND2_X1 U21818 ( .A1(n18842), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n18833) );
  OAI211_X1 U21819 ( .C1(n18834), .C2(n18935), .A(n18833), .B(n12482), .ZN(
        n18837) );
  NOR2_X1 U21820 ( .A1(n18835), .A2(n18923), .ZN(n18836) );
  AOI211_X1 U21821 ( .C1(P2_REIP_REG_12__SCAN_IN), .C2(n18910), .A(n18837), 
        .B(n18836), .ZN(n18840) );
  AOI22_X1 U21822 ( .A1(n18980), .A2(n18874), .B1(n18916), .B2(n18838), .ZN(
        n18839) );
  OAI211_X1 U21823 ( .C1(n18890), .C2(n18841), .A(n18840), .B(n18839), .ZN(
        P2_U2843) );
  NAND2_X1 U21824 ( .A1(n18842), .A2(P2_EBX_REG_11__SCAN_IN), .ZN(n18843) );
  OAI211_X1 U21825 ( .C1(n11542), .C2(n18935), .A(n18843), .B(n16114), .ZN(
        n18844) );
  AOI21_X1 U21826 ( .B1(n18910), .B2(P2_REIP_REG_11__SCAN_IN), .A(n18844), 
        .ZN(n18845) );
  OAI21_X1 U21827 ( .B1(n18924), .B2(n18846), .A(n18845), .ZN(n18848) );
  NOR2_X1 U21828 ( .A1(n18984), .A2(n18928), .ZN(n18847) );
  AOI211_X1 U21829 ( .C1(n18896), .C2(n18849), .A(n18848), .B(n18847), .ZN(
        n18853) );
  OAI211_X1 U21830 ( .C1(n18851), .C2(n18854), .A(n18920), .B(n18850), .ZN(
        n18852) );
  OAI211_X1 U21831 ( .C1(n18855), .C2(n18854), .A(n18853), .B(n18852), .ZN(
        P2_U2844) );
  NOR2_X1 U21832 ( .A1(n18929), .A2(n10059), .ZN(n18856) );
  AOI211_X1 U21833 ( .C1(n18892), .C2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .A(
        n19081), .B(n18856), .ZN(n18857) );
  OAI21_X1 U21834 ( .B1(n18858), .B2(n18923), .A(n18857), .ZN(n18859) );
  AOI21_X1 U21835 ( .B1(P2_REIP_REG_10__SCAN_IN), .B2(n18910), .A(n18859), 
        .ZN(n18865) );
  NAND2_X1 U21836 ( .A1(n9887), .A2(n18860), .ZN(n18861) );
  XNOR2_X1 U21837 ( .A(n18862), .B(n18861), .ZN(n18863) );
  AOI22_X1 U21838 ( .A1(n18863), .A2(n18920), .B1(n18916), .B2(n18956), .ZN(
        n18864) );
  OAI211_X1 U21839 ( .C1(n18928), .C2(n18987), .A(n18865), .B(n18864), .ZN(
        P2_U2845) );
  NAND2_X1 U21840 ( .A1(n9887), .A2(n18866), .ZN(n18867) );
  XOR2_X1 U21841 ( .A(n18868), .B(n18867), .Z(n18878) );
  NOR2_X1 U21842 ( .A1(n18929), .A2(n18869), .ZN(n18870) );
  AOI211_X1 U21843 ( .C1(n18892), .C2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .A(
        n19081), .B(n18870), .ZN(n18871) );
  OAI21_X1 U21844 ( .B1(n19694), .B2(n18932), .A(n18871), .ZN(n18872) );
  AOI21_X1 U21845 ( .B1(n18896), .B2(n18873), .A(n18872), .ZN(n18877) );
  AOI22_X1 U21846 ( .A1(n18916), .A2(n18875), .B1(n18874), .B2(n18990), .ZN(
        n18876) );
  OAI211_X1 U21847 ( .C1(n18890), .C2(n18878), .A(n18877), .B(n18876), .ZN(
        P2_U2847) );
  NOR2_X1 U21848 ( .A1(n18912), .A2(n18879), .ZN(n18880) );
  XOR2_X1 U21849 ( .A(n18881), .B(n18880), .Z(n18889) );
  NOR2_X1 U21850 ( .A1(n18929), .A2(n11533), .ZN(n18882) );
  AOI211_X1 U21851 ( .C1(n18892), .C2(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .A(
        n19081), .B(n18882), .ZN(n18883) );
  OAI21_X1 U21852 ( .B1(n18884), .B2(n18923), .A(n18883), .ZN(n18887) );
  OAI22_X1 U21853 ( .A1(n18994), .A2(n18928), .B1(n18924), .B2(n18885), .ZN(
        n18886) );
  AOI211_X1 U21854 ( .C1(P2_REIP_REG_7__SCAN_IN), .C2(n18910), .A(n18887), .B(
        n18886), .ZN(n18888) );
  OAI21_X1 U21855 ( .B1(n18890), .B2(n18889), .A(n18888), .ZN(P2_U2848) );
  INV_X1 U21856 ( .A(n18891), .ZN(n18897) );
  AOI22_X1 U21857 ( .A1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n18892), .B1(
        P2_REIP_REG_6__SCAN_IN), .B2(n18910), .ZN(n18893) );
  OAI211_X1 U21858 ( .C1(n18929), .C2(n18894), .A(n18893), .B(n12482), .ZN(
        n18895) );
  AOI21_X1 U21859 ( .B1(n18897), .B2(n18896), .A(n18895), .ZN(n18904) );
  NAND2_X1 U21860 ( .A1(n18831), .A2(n18898), .ZN(n18899) );
  XNOR2_X1 U21861 ( .A(n18900), .B(n18899), .ZN(n18902) );
  AOI22_X1 U21862 ( .A1(n18902), .A2(n18920), .B1(n18916), .B2(n18901), .ZN(
        n18903) );
  OAI211_X1 U21863 ( .C1(n18928), .C2(n18996), .A(n18904), .B(n18903), .ZN(
        P2_U2849) );
  OAI21_X1 U21864 ( .B1(n18929), .B2(n18905), .A(n12482), .ZN(n18909) );
  OAI22_X1 U21865 ( .A1(n18923), .A2(n18907), .B1(n18906), .B2(n18935), .ZN(
        n18908) );
  AOI211_X1 U21866 ( .C1(P2_REIP_REG_5__SCAN_IN), .C2(n18910), .A(n18909), .B(
        n18908), .ZN(n18919) );
  NOR2_X1 U21867 ( .A1(n18912), .A2(n18911), .ZN(n18914) );
  XNOR2_X1 U21868 ( .A(n18914), .B(n18913), .ZN(n18917) );
  AOI22_X1 U21869 ( .A1(n18917), .A2(n18920), .B1(n18916), .B2(n18915), .ZN(
        n18918) );
  OAI211_X1 U21870 ( .C1(n18928), .C2(n19005), .A(n18919), .B(n18918), .ZN(
        P2_U2850) );
  INV_X1 U21871 ( .A(n18921), .ZN(n18922) );
  OAI22_X1 U21872 ( .A1(n18925), .A2(n18924), .B1(n18923), .B2(n18922), .ZN(
        n18934) );
  INV_X1 U21873 ( .A(n18926), .ZN(n18927) );
  OR2_X1 U21874 ( .A1(n18928), .A2(n18927), .ZN(n18931) );
  OR2_X1 U21875 ( .A1(n18929), .A2(n11989), .ZN(n18930) );
  OAI211_X1 U21876 ( .C1(n18932), .C2(n11633), .A(n18931), .B(n18930), .ZN(
        n18933) );
  NOR2_X1 U21877 ( .A1(n18934), .A2(n18933), .ZN(n18938) );
  AOI22_X1 U21878 ( .A1(n18892), .A2(P2_PHYADDRPOINTER_REG_0__SCAN_IN), .B1(
        n18936), .B2(n19137), .ZN(n18937) );
  OAI211_X1 U21879 ( .C1(n18939), .C2(n18890), .A(n18938), .B(n18937), .ZN(
        P2_U2855) );
  NAND2_X1 U21880 ( .A1(n18941), .A2(n18940), .ZN(n18942) );
  NAND2_X1 U21881 ( .A1(n13709), .A2(n18942), .ZN(n18966) );
  INV_X1 U21882 ( .A(n18943), .ZN(n18944) );
  OAI22_X1 U21883 ( .A1(n18966), .A2(n18952), .B1(n18945), .B2(n18944), .ZN(
        n18946) );
  INV_X1 U21884 ( .A(n18946), .ZN(n18947) );
  OAI21_X1 U21885 ( .B1(n18958), .B2(n11557), .A(n18947), .ZN(P2_U2871) );
  AOI21_X1 U21886 ( .B1(n18950), .B2(n18949), .A(n18948), .ZN(n18954) );
  INV_X1 U21887 ( .A(n18951), .ZN(n18953) );
  NOR3_X1 U21888 ( .A1(n18954), .A2(n18953), .A3(n18952), .ZN(n18955) );
  AOI21_X1 U21889 ( .B1(n18956), .B2(n18958), .A(n18955), .ZN(n18957) );
  OAI21_X1 U21890 ( .B1(n18958), .B2(n10059), .A(n18957), .ZN(P2_U2877) );
  AOI22_X1 U21891 ( .A1(n18965), .A2(BUF2_REG_31__SCAN_IN), .B1(n18959), .B2(
        n19027), .ZN(n18961) );
  AOI22_X1 U21892 ( .A1(P2_EAX_REG_31__SCAN_IN), .A2(n19026), .B1(n18964), 
        .B2(BUF1_REG_31__SCAN_IN), .ZN(n18960) );
  NAND2_X1 U21893 ( .A1(n18961), .A2(n18960), .ZN(P2_U2888) );
  AOI22_X1 U21894 ( .A1(n18963), .A2(n18962), .B1(n19026), .B2(
        P2_EAX_REG_16__SCAN_IN), .ZN(n18971) );
  AOI22_X1 U21895 ( .A1(n18965), .A2(BUF2_REG_16__SCAN_IN), .B1(n18964), .B2(
        BUF1_REG_16__SCAN_IN), .ZN(n18970) );
  NOR2_X1 U21896 ( .A1(n18966), .A2(n19002), .ZN(n18967) );
  AOI21_X1 U21897 ( .B1(n18968), .B2(n19027), .A(n18967), .ZN(n18969) );
  NAND3_X1 U21898 ( .A1(n18971), .A2(n18970), .A3(n18969), .ZN(P2_U2903) );
  INV_X1 U21899 ( .A(n18972), .ZN(n18974) );
  OAI222_X1 U21900 ( .A1(n18974), .A2(n19006), .B1(n19042), .B2(n18995), .C1(
        n18973), .C2(n19035), .ZN(P2_U2904) );
  INV_X1 U21901 ( .A(n18975), .ZN(n18977) );
  INV_X1 U21902 ( .A(P2_EAX_REG_14__SCAN_IN), .ZN(n19044) );
  OAI222_X1 U21903 ( .A1(n18977), .A2(n19006), .B1(n19044), .B2(n18995), .C1(
        n19035), .C2(n18976), .ZN(P2_U2905) );
  INV_X1 U21904 ( .A(P2_EAX_REG_13__SCAN_IN), .ZN(n19046) );
  OAI222_X1 U21905 ( .A1(n18979), .A2(n19006), .B1(n19046), .B2(n18995), .C1(
        n19035), .C2(n18978), .ZN(P2_U2906) );
  INV_X1 U21906 ( .A(n18980), .ZN(n18982) );
  INV_X1 U21907 ( .A(P2_EAX_REG_12__SCAN_IN), .ZN(n19048) );
  OAI222_X1 U21908 ( .A1(n18982), .A2(n19006), .B1(n19048), .B2(n18995), .C1(
        n19035), .C2(n18981), .ZN(P2_U2907) );
  INV_X1 U21909 ( .A(P2_EAX_REG_11__SCAN_IN), .ZN(n19050) );
  OAI222_X1 U21910 ( .A1(n18984), .A2(n19006), .B1(n19050), .B2(n18995), .C1(
        n19035), .C2(n18983), .ZN(P2_U2908) );
  AOI22_X1 U21911 ( .A1(P2_EAX_REG_10__SCAN_IN), .A2(n19026), .B1(n18985), 
        .B2(n18997), .ZN(n18986) );
  OAI21_X1 U21912 ( .B1(n19006), .B2(n18987), .A(n18986), .ZN(P2_U2909) );
  INV_X1 U21913 ( .A(P2_EAX_REG_9__SCAN_IN), .ZN(n19054) );
  OAI222_X1 U21914 ( .A1(n18989), .A2(n19006), .B1(n19054), .B2(n18995), .C1(
        n19035), .C2(n18988), .ZN(P2_U2910) );
  INV_X1 U21915 ( .A(n18990), .ZN(n18993) );
  AOI22_X1 U21916 ( .A1(P2_EAX_REG_8__SCAN_IN), .A2(n19026), .B1(n18991), .B2(
        n18997), .ZN(n18992) );
  OAI21_X1 U21917 ( .B1(n19006), .B2(n18993), .A(n18992), .ZN(P2_U2911) );
  INV_X1 U21918 ( .A(P2_EAX_REG_7__SCAN_IN), .ZN(n20789) );
  OAI222_X1 U21919 ( .A1(n18994), .A2(n19006), .B1(n20789), .B2(n18995), .C1(
        n19035), .C2(n19178), .ZN(P2_U2912) );
  INV_X1 U21920 ( .A(P2_EAX_REG_6__SCAN_IN), .ZN(n19059) );
  OAI222_X1 U21921 ( .A1(n18996), .A2(n19006), .B1(n19059), .B2(n18995), .C1(
        n19035), .C2(n19172), .ZN(P2_U2913) );
  INV_X1 U21922 ( .A(n19168), .ZN(n18998) );
  AOI22_X1 U21923 ( .A1(P2_EAX_REG_5__SCAN_IN), .A2(n19026), .B1(n18998), .B2(
        n18997), .ZN(n19004) );
  XNOR2_X1 U21924 ( .A(n19760), .B(n19762), .ZN(n19021) );
  XNOR2_X1 U21925 ( .A(n18999), .B(n19771), .ZN(n19030) );
  NAND2_X1 U21926 ( .A1(n19030), .A2(n19029), .ZN(n19028) );
  OAI21_X1 U21927 ( .B1(n19767), .B2(n19771), .A(n19028), .ZN(n19020) );
  NAND2_X1 U21928 ( .A1(n19021), .A2(n19020), .ZN(n19019) );
  OAI21_X1 U21929 ( .B1(n19138), .B2(n19762), .A(n19019), .ZN(n19014) );
  XNOR2_X1 U21930 ( .A(n19754), .B(n19012), .ZN(n19015) );
  NAND2_X1 U21931 ( .A1(n19014), .A2(n19015), .ZN(n19013) );
  NAND2_X1 U21932 ( .A1(n19000), .A2(n19012), .ZN(n19001) );
  AOI21_X1 U21933 ( .B1(n19013), .B2(n19001), .A(n19095), .ZN(n19007) );
  OR3_X1 U21934 ( .A1(n19007), .A2(n19008), .A3(n19002), .ZN(n19003) );
  OAI211_X1 U21935 ( .C1(n19006), .C2(n19005), .A(n19004), .B(n19003), .ZN(
        P2_U2914) );
  AOI22_X1 U21936 ( .A1(n19027), .A2(n19095), .B1(n19026), .B2(
        P2_EAX_REG_4__SCAN_IN), .ZN(n19011) );
  XOR2_X1 U21937 ( .A(n19008), .B(n19007), .Z(n19009) );
  NAND2_X1 U21938 ( .A1(n19009), .A2(n19031), .ZN(n19010) );
  OAI211_X1 U21939 ( .C1(n19162), .C2(n19035), .A(n19011), .B(n19010), .ZN(
        P2_U2915) );
  INV_X1 U21940 ( .A(n19012), .ZN(n19753) );
  AOI22_X1 U21941 ( .A1(n19027), .A2(n19753), .B1(n19026), .B2(
        P2_EAX_REG_3__SCAN_IN), .ZN(n19018) );
  OAI21_X1 U21942 ( .B1(n19015), .B2(n19014), .A(n19013), .ZN(n19016) );
  NAND2_X1 U21943 ( .A1(n19016), .A2(n19031), .ZN(n19017) );
  OAI211_X1 U21944 ( .C1(n19157), .C2(n19035), .A(n19018), .B(n19017), .ZN(
        P2_U2916) );
  AOI22_X1 U21945 ( .A1(n19027), .A2(n19762), .B1(n19026), .B2(
        P2_EAX_REG_2__SCAN_IN), .ZN(n19024) );
  OAI21_X1 U21946 ( .B1(n19021), .B2(n19020), .A(n19019), .ZN(n19022) );
  NAND2_X1 U21947 ( .A1(n19022), .A2(n19031), .ZN(n19023) );
  OAI211_X1 U21948 ( .C1(n19025), .C2(n19035), .A(n19024), .B(n19023), .ZN(
        P2_U2917) );
  AOI22_X1 U21949 ( .A1(n19027), .A2(n19771), .B1(n19026), .B2(
        P2_EAX_REG_1__SCAN_IN), .ZN(n19034) );
  OAI21_X1 U21950 ( .B1(n19030), .B2(n19029), .A(n19028), .ZN(n19032) );
  NAND2_X1 U21951 ( .A1(n19032), .A2(n19031), .ZN(n19033) );
  OAI211_X1 U21952 ( .C1(n19150), .C2(n19035), .A(n19034), .B(n19033), .ZN(
        P2_U2918) );
  NOR2_X1 U21953 ( .A1(n19065), .A2(n19036), .ZN(P2_U2920) );
  INV_X1 U21954 ( .A(P2_UWORD_REG_10__SCAN_IN), .ZN(n20806) );
  INV_X1 U21955 ( .A(n19037), .ZN(n19039) );
  AOI22_X1 U21956 ( .A1(n19039), .A2(P2_EAX_REG_26__SCAN_IN), .B1(n19067), 
        .B2(P2_DATAO_REG_26__SCAN_IN), .ZN(n19038) );
  OAI21_X1 U21957 ( .B1(n20806), .B2(n19806), .A(n19038), .ZN(P2_U2925) );
  INV_X1 U21958 ( .A(P2_UWORD_REG_8__SCAN_IN), .ZN(n20892) );
  AOI22_X1 U21959 ( .A1(n19039), .A2(P2_EAX_REG_24__SCAN_IN), .B1(n19067), 
        .B2(P2_DATAO_REG_24__SCAN_IN), .ZN(n19040) );
  OAI21_X1 U21960 ( .B1(n20892), .B2(n19806), .A(n19040), .ZN(P2_U2927) );
  AOI22_X1 U21961 ( .A1(n9634), .A2(P2_LWORD_REG_15__SCAN_IN), .B1(n19067), 
        .B2(P2_DATAO_REG_15__SCAN_IN), .ZN(n19041) );
  OAI21_X1 U21962 ( .B1(n19042), .B2(n19071), .A(n19041), .ZN(P2_U2936) );
  AOI22_X1 U21963 ( .A1(n9634), .A2(P2_LWORD_REG_14__SCAN_IN), .B1(n19067), 
        .B2(P2_DATAO_REG_14__SCAN_IN), .ZN(n19043) );
  OAI21_X1 U21964 ( .B1(n19044), .B2(n19071), .A(n19043), .ZN(P2_U2937) );
  AOI22_X1 U21965 ( .A1(n9634), .A2(P2_LWORD_REG_13__SCAN_IN), .B1(n19067), 
        .B2(P2_DATAO_REG_13__SCAN_IN), .ZN(n19045) );
  OAI21_X1 U21966 ( .B1(n19046), .B2(n19071), .A(n19045), .ZN(P2_U2938) );
  AOI22_X1 U21967 ( .A1(n9634), .A2(P2_LWORD_REG_12__SCAN_IN), .B1(n19067), 
        .B2(P2_DATAO_REG_12__SCAN_IN), .ZN(n19047) );
  OAI21_X1 U21968 ( .B1(n19048), .B2(n19071), .A(n19047), .ZN(P2_U2939) );
  AOI22_X1 U21969 ( .A1(n9634), .A2(P2_LWORD_REG_11__SCAN_IN), .B1(n19067), 
        .B2(P2_DATAO_REG_11__SCAN_IN), .ZN(n19049) );
  OAI21_X1 U21970 ( .B1(n19050), .B2(n19071), .A(n19049), .ZN(P2_U2940) );
  AOI22_X1 U21971 ( .A1(n9634), .A2(P2_LWORD_REG_10__SCAN_IN), .B1(n19067), 
        .B2(P2_DATAO_REG_10__SCAN_IN), .ZN(n19051) );
  OAI21_X1 U21972 ( .B1(n19052), .B2(n19071), .A(n19051), .ZN(P2_U2941) );
  AOI22_X1 U21973 ( .A1(n9634), .A2(P2_LWORD_REG_9__SCAN_IN), .B1(n19067), 
        .B2(P2_DATAO_REG_9__SCAN_IN), .ZN(n19053) );
  OAI21_X1 U21974 ( .B1(n19054), .B2(n19071), .A(n19053), .ZN(P2_U2942) );
  AOI22_X1 U21975 ( .A1(n9634), .A2(P2_LWORD_REG_8__SCAN_IN), .B1(n19067), 
        .B2(P2_DATAO_REG_8__SCAN_IN), .ZN(n19055) );
  OAI21_X1 U21976 ( .B1(n19056), .B2(n19071), .A(n19055), .ZN(P2_U2943) );
  AOI22_X1 U21977 ( .A1(n9634), .A2(P2_LWORD_REG_7__SCAN_IN), .B1(n19067), 
        .B2(P2_DATAO_REG_7__SCAN_IN), .ZN(n19057) );
  OAI21_X1 U21978 ( .B1(n20789), .B2(n19071), .A(n19057), .ZN(P2_U2944) );
  AOI22_X1 U21979 ( .A1(n9634), .A2(P2_LWORD_REG_6__SCAN_IN), .B1(n19067), 
        .B2(P2_DATAO_REG_6__SCAN_IN), .ZN(n19058) );
  OAI21_X1 U21980 ( .B1(n19059), .B2(n19071), .A(n19058), .ZN(P2_U2945) );
  INV_X1 U21981 ( .A(P2_EAX_REG_5__SCAN_IN), .ZN(n19061) );
  AOI22_X1 U21982 ( .A1(n9634), .A2(P2_LWORD_REG_5__SCAN_IN), .B1(n19067), 
        .B2(P2_DATAO_REG_5__SCAN_IN), .ZN(n19060) );
  OAI21_X1 U21983 ( .B1(n19061), .B2(n19071), .A(n19060), .ZN(P2_U2946) );
  AOI22_X1 U21984 ( .A1(n9634), .A2(P2_LWORD_REG_4__SCAN_IN), .B1(n19067), 
        .B2(P2_DATAO_REG_4__SCAN_IN), .ZN(n19062) );
  OAI21_X1 U21985 ( .B1(n13125), .B2(n19071), .A(n19062), .ZN(P2_U2947) );
  AOI22_X1 U21986 ( .A1(n9634), .A2(P2_LWORD_REG_3__SCAN_IN), .B1(n19067), 
        .B2(P2_DATAO_REG_3__SCAN_IN), .ZN(n19063) );
  OAI21_X1 U21987 ( .B1(n13099), .B2(n19071), .A(n19063), .ZN(P2_U2948) );
  INV_X1 U21988 ( .A(P2_EAX_REG_2__SCAN_IN), .ZN(n19066) );
  OAI222_X1 U21989 ( .A1(n19806), .A2(n13254), .B1(n19071), .B2(n19066), .C1(
        n19065), .C2(n19064), .ZN(P2_U2949) );
  INV_X1 U21990 ( .A(P2_EAX_REG_1__SCAN_IN), .ZN(n19069) );
  AOI22_X1 U21991 ( .A1(n9634), .A2(P2_LWORD_REG_1__SCAN_IN), .B1(n19067), 
        .B2(P2_DATAO_REG_1__SCAN_IN), .ZN(n19068) );
  OAI21_X1 U21992 ( .B1(n19069), .B2(n19071), .A(n19068), .ZN(P2_U2950) );
  AOI22_X1 U21993 ( .A1(n9634), .A2(P2_LWORD_REG_0__SCAN_IN), .B1(n19067), 
        .B2(P2_DATAO_REG_0__SCAN_IN), .ZN(n19070) );
  OAI21_X1 U21994 ( .B1(n13343), .B2(n19071), .A(n19070), .ZN(P2_U2951) );
  INV_X1 U21995 ( .A(n19072), .ZN(n19073) );
  AOI21_X1 U21996 ( .B1(n19077), .B2(P2_EAX_REG_24__SCAN_IN), .A(n19073), .ZN(
        n19074) );
  OAI21_X1 U21997 ( .B1(n20892), .B2(n13250), .A(n19074), .ZN(P2_U2960) );
  INV_X1 U21998 ( .A(n19075), .ZN(n19076) );
  AOI21_X1 U21999 ( .B1(n19077), .B2(P2_EAX_REG_26__SCAN_IN), .A(n19076), .ZN(
        n19078) );
  OAI21_X1 U22000 ( .B1(n20806), .B2(n13250), .A(n19078), .ZN(P2_U2962) );
  AOI22_X1 U22001 ( .A1(P2_REIP_REG_4__SCAN_IN), .A2(n19081), .B1(n19080), 
        .B2(n19079), .ZN(n19092) );
  XNOR2_X1 U22002 ( .A(n19082), .B(n19083), .ZN(n19098) );
  XNOR2_X1 U22003 ( .A(n19084), .B(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n19086) );
  XNOR2_X1 U22004 ( .A(n19086), .B(n19085), .ZN(n19097) );
  OAI22_X1 U22005 ( .A1(n19098), .A2(n19088), .B1(n19097), .B2(n19087), .ZN(
        n19089) );
  AOI21_X1 U22006 ( .B1(n19090), .B2(n19096), .A(n19089), .ZN(n19091) );
  OAI211_X1 U22007 ( .C1(n19094), .C2(n19093), .A(n19092), .B(n19091), .ZN(
        P2_U3010) );
  INV_X1 U22008 ( .A(P2_REIP_REG_4__SCAN_IN), .ZN(n19688) );
  AOI22_X1 U22009 ( .A1(n19096), .A2(n19131), .B1(n19122), .B2(n19095), .ZN(
        n19104) );
  OAI22_X1 U22010 ( .A1(n19098), .A2(n19110), .B1(n19097), .B2(n19125), .ZN(
        n19099) );
  AOI221_X1 U22011 ( .B1(n19102), .B2(n19101), .C1(n19100), .C2(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .A(n19099), .ZN(n19103) );
  OAI211_X1 U22012 ( .C1(n19688), .C2(n12482), .A(n19104), .B(n19103), .ZN(
        P2_U3042) );
  AOI22_X1 U22013 ( .A1(n19106), .A2(n19105), .B1(n19122), .B2(n19762), .ZN(
        n19121) );
  NAND2_X1 U22014 ( .A1(n19108), .A2(n19107), .ZN(n19109) );
  NOR2_X1 U22015 ( .A1(n19110), .A2(n19109), .ZN(n19115) );
  OAI22_X1 U22016 ( .A1(n13011), .A2(n19112), .B1(n19125), .B2(n19111), .ZN(
        n19114) );
  NOR3_X1 U22017 ( .A1(n19115), .A2(n19114), .A3(n19113), .ZN(n19120) );
  OAI221_X1 U22018 ( .B1(n19124), .B2(n19117), .C1(n19124), .C2(n19116), .A(
        P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n19119) );
  NAND4_X1 U22019 ( .A1(n19121), .A2(n19120), .A3(n19119), .A4(n19118), .ZN(
        P2_U3044) );
  AOI22_X1 U22020 ( .A1(n12942), .A2(n19123), .B1(n19122), .B2(n19771), .ZN(
        n19136) );
  INV_X1 U22021 ( .A(n19124), .ZN(n19127) );
  OAI22_X1 U22022 ( .A1(n19127), .A2(n11463), .B1(n19126), .B2(n19125), .ZN(
        n19128) );
  AOI211_X1 U22023 ( .C1(n19131), .C2(n19130), .A(n19129), .B(n19128), .ZN(
        n19135) );
  OAI211_X1 U22024 ( .C1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(n19133), .B(n19132), .ZN(n19134) );
  NAND3_X1 U22025 ( .A1(n19136), .A2(n19135), .A3(n19134), .ZN(P2_U3045) );
  NOR2_X2 U22026 ( .A1(n19534), .A2(n19587), .ZN(n19652) );
  NAND2_X1 U22027 ( .A1(n19752), .A2(n19208), .ZN(n19139) );
  NAND2_X1 U22028 ( .A1(n19752), .A2(n19221), .ZN(n19556) );
  OAI21_X1 U22029 ( .B1(n19652), .B2(n19139), .A(n19556), .ZN(n19142) );
  NOR2_X1 U22030 ( .A1(n19364), .A2(n19217), .ZN(n19177) );
  INV_X1 U22031 ( .A(n19177), .ZN(n19140) );
  AND2_X1 U22032 ( .A1(n19591), .A2(n19140), .ZN(n19145) );
  INV_X1 U22033 ( .A(n12128), .ZN(n19143) );
  AOI211_X1 U22034 ( .C1(n19143), .C2(n19594), .A(n19752), .B(n19177), .ZN(
        n19141) );
  INV_X1 U22035 ( .A(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n19149) );
  AOI22_X1 U22036 ( .A1(n19602), .A2(n19652), .B1(n19600), .B2(n19177), .ZN(
        n19148) );
  INV_X1 U22037 ( .A(n19142), .ZN(n19146) );
  OAI21_X1 U22038 ( .B1(n19143), .B2(n19177), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19144) );
  AOI22_X1 U22039 ( .A1(n19601), .A2(n19181), .B1(n19211), .B2(n19603), .ZN(
        n19147) );
  OAI211_X1 U22040 ( .C1(n19184), .C2(n19149), .A(n19148), .B(n19147), .ZN(
        P2_U3048) );
  AOI22_X2 U22041 ( .A1(BUF2_REG_25__SCAN_IN), .A2(n19180), .B1(
        BUF1_REG_25__SCAN_IN), .B2(n19179), .ZN(n19503) );
  INV_X1 U22042 ( .A(n19503), .ZN(n19609) );
  NOR2_X2 U22043 ( .A1(n12068), .A2(n19176), .ZN(n19607) );
  AOI22_X1 U22044 ( .A1(n19609), .A2(n19652), .B1(n19177), .B2(n19607), .ZN(
        n19153) );
  NOR2_X2 U22045 ( .A1(n19150), .A2(n19528), .ZN(n19608) );
  OAI22_X2 U22046 ( .A1(n14427), .A2(n19165), .B1(n19151), .B2(n19163), .ZN(
        n19610) );
  AOI22_X1 U22047 ( .A1(n19608), .A2(n19181), .B1(n19211), .B2(n19610), .ZN(
        n19152) );
  OAI211_X1 U22048 ( .C1(n19184), .C2(n12061), .A(n19153), .B(n19152), .ZN(
        P2_U3049) );
  AOI22_X1 U22049 ( .A1(n19616), .A2(n19652), .B1(n19613), .B2(n19177), .ZN(
        n19155) );
  AOI22_X1 U22050 ( .A1(n19614), .A2(n19181), .B1(n19211), .B2(n19615), .ZN(
        n19154) );
  OAI211_X1 U22051 ( .C1(n19184), .C2(n12524), .A(n19155), .B(n19154), .ZN(
        P2_U3050) );
  AOI22_X2 U22052 ( .A1(BUF2_REG_27__SCAN_IN), .A2(n19180), .B1(
        BUF1_REG_27__SCAN_IN), .B2(n19179), .ZN(n19509) );
  INV_X1 U22053 ( .A(n19509), .ZN(n19621) );
  NOR2_X2 U22054 ( .A1(n19156), .A2(n19176), .ZN(n19619) );
  AOI22_X1 U22055 ( .A1(n19621), .A2(n19652), .B1(n19177), .B2(n19619), .ZN(
        n19160) );
  NOR2_X2 U22056 ( .A1(n19157), .A2(n19528), .ZN(n19620) );
  OAI22_X2 U22057 ( .A1(n14416), .A2(n19165), .B1(n19158), .B2(n19163), .ZN(
        n19622) );
  AOI22_X1 U22058 ( .A1(n19620), .A2(n19181), .B1(n19211), .B2(n19622), .ZN(
        n19159) );
  OAI211_X1 U22059 ( .C1(n19184), .C2(n19161), .A(n19160), .B(n19159), .ZN(
        P2_U3051) );
  AOI22_X2 U22060 ( .A1(BUF1_REG_28__SCAN_IN), .A2(n19179), .B1(
        BUF2_REG_28__SCAN_IN), .B2(n19180), .ZN(n19512) );
  INV_X1 U22061 ( .A(n19512), .ZN(n19628) );
  NOR2_X2 U22062 ( .A1(n11450), .A2(n19176), .ZN(n19626) );
  AOI22_X1 U22063 ( .A1(n19628), .A2(n19652), .B1(n19177), .B2(n19626), .ZN(
        n19167) );
  NOR2_X2 U22064 ( .A1(n19162), .A2(n19528), .ZN(n19627) );
  OAI22_X2 U22065 ( .A1(n14410), .A2(n19165), .B1(n19164), .B2(n19163), .ZN(
        n19629) );
  AOI22_X1 U22066 ( .A1(n19627), .A2(n19181), .B1(n19211), .B2(n19629), .ZN(
        n19166) );
  OAI211_X1 U22067 ( .C1(n19184), .C2(n12545), .A(n19167), .B(n19166), .ZN(
        P2_U3052) );
  AOI22_X1 U22068 ( .A1(BUF1_REG_29__SCAN_IN), .A2(n19179), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n19180), .ZN(n19515) );
  NOR2_X2 U22069 ( .A1(n12327), .A2(n19176), .ZN(n19632) );
  AOI22_X1 U22070 ( .A1(n19634), .A2(n19652), .B1(n19177), .B2(n19632), .ZN(
        n19170) );
  NOR2_X2 U22071 ( .A1(n19168), .A2(n19528), .ZN(n19633) );
  AOI22_X1 U22072 ( .A1(BUF1_REG_21__SCAN_IN), .A2(n19179), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n19180), .ZN(n19478) );
  AOI22_X1 U22073 ( .A1(n19633), .A2(n19181), .B1(n19211), .B2(n19635), .ZN(
        n19169) );
  OAI211_X1 U22074 ( .C1(n19184), .C2(n19171), .A(n19170), .B(n19169), .ZN(
        P2_U3053) );
  AOI22_X1 U22075 ( .A1(BUF2_REG_30__SCAN_IN), .A2(n19180), .B1(
        BUF1_REG_30__SCAN_IN), .B2(n19179), .ZN(n19518) );
  NOR2_X2 U22076 ( .A1(n11434), .A2(n19176), .ZN(n19638) );
  AOI22_X1 U22077 ( .A1(n19652), .A2(n19641), .B1(n19177), .B2(n19638), .ZN(
        n19174) );
  NOR2_X2 U22078 ( .A1(n19172), .A2(n19528), .ZN(n19639) );
  AOI22_X1 U22079 ( .A1(BUF1_REG_22__SCAN_IN), .A2(n19179), .B1(
        BUF2_REG_22__SCAN_IN), .B2(n19180), .ZN(n19482) );
  INV_X1 U22080 ( .A(n19482), .ZN(n19640) );
  AOI22_X1 U22081 ( .A1(n19639), .A2(n19181), .B1(n19211), .B2(n19640), .ZN(
        n19173) );
  OAI211_X1 U22082 ( .C1(n19184), .C2(n19175), .A(n19174), .B(n19173), .ZN(
        P2_U3054) );
  AOI22_X1 U22083 ( .A1(BUF1_REG_31__SCAN_IN), .A2(n19179), .B1(
        BUF2_REG_31__SCAN_IN), .B2(n19180), .ZN(n19525) );
  INV_X1 U22084 ( .A(n19525), .ZN(n19649) );
  NOR2_X2 U22085 ( .A1(n11630), .A2(n19176), .ZN(n19645) );
  AOI22_X1 U22086 ( .A1(n19649), .A2(n19652), .B1(n19177), .B2(n19645), .ZN(
        n19183) );
  NOR2_X2 U22087 ( .A1(n19178), .A2(n19528), .ZN(n19647) );
  AOI22_X1 U22088 ( .A1(BUF2_REG_23__SCAN_IN), .A2(n19180), .B1(
        BUF1_REG_23__SCAN_IN), .B2(n19179), .ZN(n19424) );
  AOI22_X1 U22089 ( .A1(n19647), .A2(n19181), .B1(n19211), .B2(n19651), .ZN(
        n19182) );
  OAI211_X1 U22090 ( .C1(n19184), .C2(n12544), .A(n19183), .B(n19182), .ZN(
        P2_U3055) );
  INV_X1 U22091 ( .A(n19395), .ZN(n19186) );
  OR2_X1 U22092 ( .A1(n19217), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n19191) );
  NAND2_X1 U22093 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n19801), .ZN(n19659) );
  INV_X1 U22094 ( .A(n19659), .ZN(n19189) );
  NOR3_X2 U22095 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19783), .A3(
        n19217), .ZN(n19209) );
  INV_X1 U22096 ( .A(n19209), .ZN(n19187) );
  NAND3_X1 U22097 ( .A1(n12129), .A2(P2_STATE2_REG_2__SCAN_IN), .A3(n19187), 
        .ZN(n19192) );
  INV_X1 U22098 ( .A(n19192), .ZN(n19188) );
  AOI211_X2 U22099 ( .C1(n19801), .C2(n19191), .A(n19189), .B(n19188), .ZN(
        n19210) );
  AOI22_X1 U22100 ( .A1(n19210), .A2(n19601), .B1(n19600), .B2(n19209), .ZN(
        n19195) );
  NOR2_X1 U22101 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19594), .ZN(
        n19780) );
  OR3_X1 U22102 ( .A1(n19395), .A2(n19338), .A3(P2_STATE2_REG_3__SCAN_IN), 
        .ZN(n19190) );
  OAI21_X1 U22103 ( .B1(n19780), .B2(n19191), .A(n19190), .ZN(n19193) );
  NAND3_X1 U22104 ( .A1(n19193), .A2(n19593), .A3(n19192), .ZN(n19212) );
  AOI22_X1 U22105 ( .A1(P2_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n19212), .B1(
        n19211), .B2(n19602), .ZN(n19194) );
  OAI211_X1 U22106 ( .C1(n19466), .C2(n19246), .A(n19195), .B(n19194), .ZN(
        P2_U3056) );
  AOI22_X1 U22107 ( .A1(n19210), .A2(n19608), .B1(n19607), .B2(n19209), .ZN(
        n19197) );
  AOI22_X1 U22108 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n19212), .B1(
        n19238), .B2(n19610), .ZN(n19196) );
  OAI211_X1 U22109 ( .C1(n19503), .C2(n19208), .A(n19197), .B(n19196), .ZN(
        P2_U3057) );
  AOI22_X1 U22110 ( .A1(n19210), .A2(n19614), .B1(n19613), .B2(n19209), .ZN(
        n19199) );
  AOI22_X1 U22111 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n19212), .B1(
        n19211), .B2(n19616), .ZN(n19198) );
  OAI211_X1 U22112 ( .C1(n19471), .C2(n19246), .A(n19199), .B(n19198), .ZN(
        P2_U3058) );
  AOI22_X1 U22113 ( .A1(n19210), .A2(n19620), .B1(n19619), .B2(n19209), .ZN(
        n19201) );
  AOI22_X1 U22114 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n19212), .B1(
        n19238), .B2(n19622), .ZN(n19200) );
  OAI211_X1 U22115 ( .C1(n19509), .C2(n19208), .A(n19201), .B(n19200), .ZN(
        P2_U3059) );
  AOI22_X1 U22116 ( .A1(n19210), .A2(n19627), .B1(n19626), .B2(n19209), .ZN(
        n19203) );
  AOI22_X1 U22117 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n19212), .B1(
        n19238), .B2(n19629), .ZN(n19202) );
  OAI211_X1 U22118 ( .C1(n19512), .C2(n19208), .A(n19203), .B(n19202), .ZN(
        P2_U3060) );
  AOI22_X1 U22119 ( .A1(n19210), .A2(n19633), .B1(n19632), .B2(n19209), .ZN(
        n19205) );
  AOI22_X1 U22120 ( .A1(P2_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n19212), .B1(
        n19238), .B2(n19635), .ZN(n19204) );
  OAI211_X1 U22121 ( .C1(n19515), .C2(n19208), .A(n19205), .B(n19204), .ZN(
        P2_U3061) );
  AOI22_X1 U22122 ( .A1(n19210), .A2(n19639), .B1(n19638), .B2(n19209), .ZN(
        n19207) );
  AOI22_X1 U22123 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n19212), .B1(
        n19238), .B2(n19640), .ZN(n19206) );
  OAI211_X1 U22124 ( .C1(n19518), .C2(n19208), .A(n19207), .B(n19206), .ZN(
        P2_U3062) );
  AOI22_X1 U22125 ( .A1(n19210), .A2(n19647), .B1(n19645), .B2(n19209), .ZN(
        n19214) );
  AOI22_X1 U22126 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n19212), .B1(
        n19211), .B2(n19649), .ZN(n19213) );
  OAI211_X1 U22127 ( .C1(n19424), .C2(n19246), .A(n19214), .B(n19213), .ZN(
        P2_U3063) );
  INV_X1 U22128 ( .A(n12104), .ZN(n19216) );
  NOR2_X1 U22129 ( .A1(n19215), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n19241) );
  OAI21_X1 U22130 ( .B1(n19216), .B2(n19241), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19218) );
  OR2_X1 U22131 ( .A1(n19427), .A2(n19217), .ZN(n19220) );
  NAND2_X1 U22132 ( .A1(n19218), .A2(n19220), .ZN(n19242) );
  AOI22_X1 U22133 ( .A1(n19242), .A2(n19601), .B1(n19600), .B2(n19241), .ZN(
        n19227) );
  INV_X1 U22134 ( .A(n19241), .ZN(n19219) );
  OAI21_X1 U22135 ( .B1(n12104), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n19219), 
        .ZN(n19224) );
  NOR2_X1 U22136 ( .A1(n19263), .A2(n19238), .ZN(n19222) );
  OAI21_X1 U22137 ( .B1(n19222), .B2(n19221), .A(n19220), .ZN(n19223) );
  MUX2_X1 U22138 ( .A(n19224), .B(n19223), .S(n19752), .Z(n19225) );
  NAND2_X1 U22139 ( .A1(n19225), .A2(n19593), .ZN(n19243) );
  AOI22_X1 U22140 ( .A1(P2_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n19243), .B1(
        n19263), .B2(n19603), .ZN(n19226) );
  OAI211_X1 U22141 ( .C1(n19500), .C2(n19246), .A(n19227), .B(n19226), .ZN(
        P2_U3064) );
  AOI22_X1 U22142 ( .A1(n19242), .A2(n19608), .B1(n19607), .B2(n19241), .ZN(
        n19229) );
  AOI22_X1 U22143 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n19243), .B1(
        n19263), .B2(n19610), .ZN(n19228) );
  OAI211_X1 U22144 ( .C1(n19503), .C2(n19246), .A(n19229), .B(n19228), .ZN(
        P2_U3065) );
  AOI22_X1 U22145 ( .A1(n19242), .A2(n19614), .B1(n19613), .B2(n19241), .ZN(
        n19231) );
  AOI22_X1 U22146 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n19243), .B1(
        n19238), .B2(n19616), .ZN(n19230) );
  OAI211_X1 U22147 ( .C1(n19471), .C2(n19261), .A(n19231), .B(n19230), .ZN(
        P2_U3066) );
  AOI22_X1 U22148 ( .A1(n19242), .A2(n19620), .B1(n19619), .B2(n19241), .ZN(
        n19233) );
  AOI22_X1 U22149 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n19243), .B1(
        n19263), .B2(n19622), .ZN(n19232) );
  OAI211_X1 U22150 ( .C1(n19509), .C2(n19246), .A(n19233), .B(n19232), .ZN(
        P2_U3067) );
  AOI22_X1 U22151 ( .A1(n19242), .A2(n19627), .B1(n19626), .B2(n19241), .ZN(
        n19235) );
  AOI22_X1 U22152 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n19243), .B1(
        n19263), .B2(n19629), .ZN(n19234) );
  OAI211_X1 U22153 ( .C1(n19512), .C2(n19246), .A(n19235), .B(n19234), .ZN(
        P2_U3068) );
  AOI22_X1 U22154 ( .A1(n19242), .A2(n19633), .B1(n19632), .B2(n19241), .ZN(
        n19237) );
  AOI22_X1 U22155 ( .A1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n19243), .B1(
        n19263), .B2(n19635), .ZN(n19236) );
  OAI211_X1 U22156 ( .C1(n19515), .C2(n19246), .A(n19237), .B(n19236), .ZN(
        P2_U3069) );
  AOI22_X1 U22157 ( .A1(n19242), .A2(n19639), .B1(n19638), .B2(n19241), .ZN(
        n19240) );
  AOI22_X1 U22158 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n19243), .B1(
        n19238), .B2(n19641), .ZN(n19239) );
  OAI211_X1 U22159 ( .C1(n19482), .C2(n19261), .A(n19240), .B(n19239), .ZN(
        P2_U3070) );
  AOI22_X1 U22160 ( .A1(n19242), .A2(n19647), .B1(n19645), .B2(n19241), .ZN(
        n19245) );
  AOI22_X1 U22161 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n19243), .B1(
        n19263), .B2(n19651), .ZN(n19244) );
  OAI211_X1 U22162 ( .C1(n19525), .C2(n19246), .A(n19245), .B(n19244), .ZN(
        P2_U3071) );
  INV_X1 U22163 ( .A(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n19249) );
  AOI22_X1 U22164 ( .A1(n19602), .A2(n19263), .B1(n19600), .B2(n19262), .ZN(
        n19248) );
  AOI22_X1 U22165 ( .A1(n19601), .A2(n19264), .B1(n19276), .B2(n19603), .ZN(
        n19247) );
  OAI211_X1 U22166 ( .C1(n19250), .C2(n19249), .A(n19248), .B(n19247), .ZN(
        P2_U3072) );
  AOI22_X1 U22167 ( .A1(n19276), .A2(n19610), .B1(n19262), .B2(n19607), .ZN(
        n19252) );
  AOI22_X1 U22168 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n19265), .B1(
        n19608), .B2(n19264), .ZN(n19251) );
  OAI211_X1 U22169 ( .C1(n19503), .C2(n19261), .A(n19252), .B(n19251), .ZN(
        P2_U3073) );
  AOI22_X1 U22170 ( .A1(n19276), .A2(n19622), .B1(n19262), .B2(n19619), .ZN(
        n19254) );
  AOI22_X1 U22171 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n19265), .B1(
        n19620), .B2(n19264), .ZN(n19253) );
  OAI211_X1 U22172 ( .C1(n19509), .C2(n19261), .A(n19254), .B(n19253), .ZN(
        P2_U3075) );
  AOI22_X1 U22173 ( .A1(n19276), .A2(n19629), .B1(n19262), .B2(n19626), .ZN(
        n19256) );
  AOI22_X1 U22174 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n19265), .B1(
        n19627), .B2(n19264), .ZN(n19255) );
  OAI211_X1 U22175 ( .C1(n19512), .C2(n19261), .A(n19256), .B(n19255), .ZN(
        P2_U3076) );
  AOI22_X1 U22176 ( .A1(n19634), .A2(n19263), .B1(n19262), .B2(n19632), .ZN(
        n19258) );
  AOI22_X1 U22177 ( .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n19265), .B1(
        n19633), .B2(n19264), .ZN(n19257) );
  OAI211_X1 U22178 ( .C1(n19478), .C2(n19286), .A(n19258), .B(n19257), .ZN(
        P2_U3077) );
  AOI22_X1 U22179 ( .A1(n19276), .A2(n19640), .B1(n19262), .B2(n19638), .ZN(
        n19260) );
  AOI22_X1 U22180 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n19265), .B1(
        n19639), .B2(n19264), .ZN(n19259) );
  OAI211_X1 U22181 ( .C1(n19518), .C2(n19261), .A(n19260), .B(n19259), .ZN(
        P2_U3078) );
  AOI22_X1 U22182 ( .A1(n19649), .A2(n19263), .B1(n19262), .B2(n19645), .ZN(
        n19267) );
  AOI22_X1 U22183 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n19265), .B1(
        n19647), .B2(n19264), .ZN(n19266) );
  OAI211_X1 U22184 ( .C1(n19424), .C2(n19286), .A(n19267), .B(n19266), .ZN(
        P2_U3079) );
  AOI22_X1 U22185 ( .A1(n19282), .A2(n19608), .B1(n19607), .B2(n19281), .ZN(
        n19269) );
  AOI22_X1 U22186 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n19283), .B1(
        n19299), .B2(n19610), .ZN(n19268) );
  OAI211_X1 U22187 ( .C1(n19503), .C2(n19286), .A(n19269), .B(n19268), .ZN(
        P2_U3081) );
  AOI22_X1 U22188 ( .A1(n19282), .A2(n19614), .B1(n19613), .B2(n19281), .ZN(
        n19271) );
  AOI22_X1 U22189 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n19283), .B1(
        n19276), .B2(n19616), .ZN(n19270) );
  OAI211_X1 U22190 ( .C1(n19471), .C2(n19293), .A(n19271), .B(n19270), .ZN(
        P2_U3082) );
  AOI22_X1 U22191 ( .A1(n19282), .A2(n19620), .B1(n19619), .B2(n19281), .ZN(
        n19273) );
  AOI22_X1 U22192 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n19283), .B1(
        n19299), .B2(n19622), .ZN(n19272) );
  OAI211_X1 U22193 ( .C1(n19509), .C2(n19286), .A(n19273), .B(n19272), .ZN(
        P2_U3083) );
  AOI22_X1 U22194 ( .A1(n19282), .A2(n19627), .B1(n19626), .B2(n19281), .ZN(
        n19275) );
  AOI22_X1 U22195 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n19283), .B1(
        n19299), .B2(n19629), .ZN(n19274) );
  OAI211_X1 U22196 ( .C1(n19512), .C2(n19286), .A(n19275), .B(n19274), .ZN(
        P2_U3084) );
  AOI22_X1 U22197 ( .A1(n19282), .A2(n19633), .B1(n19632), .B2(n19281), .ZN(
        n19278) );
  AOI22_X1 U22198 ( .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n19283), .B1(
        n19276), .B2(n19634), .ZN(n19277) );
  OAI211_X1 U22199 ( .C1(n19478), .C2(n19293), .A(n19278), .B(n19277), .ZN(
        P2_U3085) );
  AOI22_X1 U22200 ( .A1(n19282), .A2(n19639), .B1(n19638), .B2(n19281), .ZN(
        n19280) );
  AOI22_X1 U22201 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n19283), .B1(
        n19299), .B2(n19640), .ZN(n19279) );
  OAI211_X1 U22202 ( .C1(n19518), .C2(n19286), .A(n19280), .B(n19279), .ZN(
        P2_U3086) );
  AOI22_X1 U22203 ( .A1(n19282), .A2(n19647), .B1(n19645), .B2(n19281), .ZN(
        n19285) );
  AOI22_X1 U22204 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n19283), .B1(
        n19299), .B2(n19651), .ZN(n19284) );
  OAI211_X1 U22205 ( .C1(n19525), .C2(n19286), .A(n19285), .B(n19284), .ZN(
        P2_U3087) );
  AOI22_X1 U22206 ( .A1(n19324), .A2(n19610), .B1(n19298), .B2(n19607), .ZN(
        n19288) );
  AOI22_X1 U22207 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n19301), .B1(
        n19608), .B2(n19300), .ZN(n19287) );
  OAI211_X1 U22208 ( .C1(n19503), .C2(n19293), .A(n19288), .B(n19287), .ZN(
        P2_U3089) );
  AOI22_X1 U22209 ( .A1(n19324), .A2(n19622), .B1(n19298), .B2(n19619), .ZN(
        n19290) );
  AOI22_X1 U22210 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n19301), .B1(
        n19620), .B2(n19300), .ZN(n19289) );
  OAI211_X1 U22211 ( .C1(n19509), .C2(n19293), .A(n19290), .B(n19289), .ZN(
        P2_U3091) );
  AOI22_X1 U22212 ( .A1(n19324), .A2(n19629), .B1(n19298), .B2(n19626), .ZN(
        n19292) );
  AOI22_X1 U22213 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n19301), .B1(
        n19627), .B2(n19300), .ZN(n19291) );
  OAI211_X1 U22214 ( .C1(n19512), .C2(n19293), .A(n19292), .B(n19291), .ZN(
        P2_U3092) );
  AOI22_X1 U22215 ( .A1(n19634), .A2(n19299), .B1(n19298), .B2(n19632), .ZN(
        n19295) );
  AOI22_X1 U22216 ( .A1(P2_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n19301), .B1(
        n19633), .B2(n19300), .ZN(n19294) );
  OAI211_X1 U22217 ( .C1(n19478), .C2(n19332), .A(n19295), .B(n19294), .ZN(
        P2_U3093) );
  AOI22_X1 U22218 ( .A1(n19641), .A2(n19299), .B1(n19298), .B2(n19638), .ZN(
        n19297) );
  AOI22_X1 U22219 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n19301), .B1(
        n19639), .B2(n19300), .ZN(n19296) );
  OAI211_X1 U22220 ( .C1(n19482), .C2(n19332), .A(n19297), .B(n19296), .ZN(
        P2_U3094) );
  AOI22_X1 U22221 ( .A1(n19649), .A2(n19299), .B1(n19298), .B2(n19645), .ZN(
        n19303) );
  AOI22_X1 U22222 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n19301), .B1(
        n19647), .B2(n19300), .ZN(n19302) );
  OAI211_X1 U22223 ( .C1(n19424), .C2(n19332), .A(n19303), .B(n19302), .ZN(
        P2_U3095) );
  NAND2_X1 U22224 ( .A1(n19304), .A2(n19333), .ZN(n19309) );
  OR2_X1 U22225 ( .A1(n19309), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19306) );
  INV_X1 U22226 ( .A(n12107), .ZN(n19305) );
  NOR3_X2 U22227 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A3(n19590), .ZN(n19327) );
  NOR3_X1 U22228 ( .A1(n19305), .A2(n19801), .A3(n19327), .ZN(n19308) );
  AOI21_X1 U22229 ( .B1(n19801), .B2(n19306), .A(n19308), .ZN(n19328) );
  AOI22_X1 U22230 ( .A1(n19328), .A2(n19601), .B1(n19600), .B2(n19327), .ZN(
        n19313) );
  OAI21_X1 U22231 ( .B1(n19324), .B2(n19360), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19310) );
  AOI211_X1 U22232 ( .C1(n19310), .C2(n19309), .A(n19528), .B(n19308), .ZN(
        n19311) );
  AOI22_X1 U22233 ( .A1(P2_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n19329), .B1(
        n19360), .B2(n19603), .ZN(n19312) );
  OAI211_X1 U22234 ( .C1(n19500), .C2(n19332), .A(n19313), .B(n19312), .ZN(
        P2_U3096) );
  AOI22_X1 U22235 ( .A1(n19328), .A2(n19608), .B1(n19607), .B2(n19327), .ZN(
        n19315) );
  AOI22_X1 U22236 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n19329), .B1(
        n19360), .B2(n19610), .ZN(n19314) );
  OAI211_X1 U22237 ( .C1(n19503), .C2(n19332), .A(n19315), .B(n19314), .ZN(
        P2_U3097) );
  AOI22_X1 U22238 ( .A1(n19328), .A2(n19614), .B1(n19613), .B2(n19327), .ZN(
        n19317) );
  AOI22_X1 U22239 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n19329), .B1(
        n19324), .B2(n19616), .ZN(n19316) );
  OAI211_X1 U22240 ( .C1(n19471), .C2(n19353), .A(n19317), .B(n19316), .ZN(
        P2_U3098) );
  AOI22_X1 U22241 ( .A1(n19328), .A2(n19620), .B1(n19619), .B2(n19327), .ZN(
        n19319) );
  AOI22_X1 U22242 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n19329), .B1(
        n19360), .B2(n19622), .ZN(n19318) );
  OAI211_X1 U22243 ( .C1(n19509), .C2(n19332), .A(n19319), .B(n19318), .ZN(
        P2_U3099) );
  AOI22_X1 U22244 ( .A1(n19328), .A2(n19627), .B1(n19626), .B2(n19327), .ZN(
        n19321) );
  AOI22_X1 U22245 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n19329), .B1(
        n19360), .B2(n19629), .ZN(n19320) );
  OAI211_X1 U22246 ( .C1(n19512), .C2(n19332), .A(n19321), .B(n19320), .ZN(
        P2_U3100) );
  AOI22_X1 U22247 ( .A1(n19328), .A2(n19633), .B1(n19632), .B2(n19327), .ZN(
        n19323) );
  AOI22_X1 U22248 ( .A1(P2_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n19329), .B1(
        n19324), .B2(n19634), .ZN(n19322) );
  OAI211_X1 U22249 ( .C1(n19478), .C2(n19353), .A(n19323), .B(n19322), .ZN(
        P2_U3101) );
  AOI22_X1 U22250 ( .A1(n19328), .A2(n19639), .B1(n19638), .B2(n19327), .ZN(
        n19326) );
  AOI22_X1 U22251 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n19329), .B1(
        n19324), .B2(n19641), .ZN(n19325) );
  OAI211_X1 U22252 ( .C1(n19482), .C2(n19353), .A(n19326), .B(n19325), .ZN(
        P2_U3102) );
  AOI22_X1 U22253 ( .A1(n19328), .A2(n19647), .B1(n19645), .B2(n19327), .ZN(
        n19331) );
  AOI22_X1 U22254 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n19329), .B1(
        n19360), .B2(n19651), .ZN(n19330) );
  OAI211_X1 U22255 ( .C1(n19525), .C2(n19332), .A(n19331), .B(n19330), .ZN(
        P2_U3103) );
  NOR2_X1 U22256 ( .A1(n19590), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n19341) );
  INV_X1 U22257 ( .A(n19341), .ZN(n19337) );
  INV_X1 U22258 ( .A(n19339), .ZN(n19335) );
  INV_X1 U22259 ( .A(n19455), .ZN(n19334) );
  NAND2_X1 U22260 ( .A1(n19334), .A2(n19333), .ZN(n19372) );
  INV_X1 U22261 ( .A(n19372), .ZN(n19358) );
  OAI21_X1 U22262 ( .B1(n19335), .B2(n19358), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19336) );
  OAI21_X1 U22263 ( .B1(n19337), .B2(n19747), .A(n19336), .ZN(n19359) );
  AOI22_X1 U22264 ( .A1(n19359), .A2(n19601), .B1(n19358), .B2(n19600), .ZN(
        n19344) );
  NOR2_X1 U22265 ( .A1(n19338), .A2(n19587), .ZN(n19751) );
  OAI211_X1 U22266 ( .C1(n19339), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19747), 
        .B(n19372), .ZN(n19340) );
  OAI211_X1 U22267 ( .C1(n19751), .C2(n19341), .A(n19593), .B(n19340), .ZN(
        n19361) );
  AOI22_X1 U22268 ( .A1(P2_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n19361), .B1(
        n19386), .B2(n19603), .ZN(n19343) );
  OAI211_X1 U22269 ( .C1(n19500), .C2(n19353), .A(n19344), .B(n19343), .ZN(
        P2_U3104) );
  AOI22_X1 U22270 ( .A1(n19359), .A2(n19608), .B1(n19358), .B2(n19607), .ZN(
        n19346) );
  AOI22_X1 U22271 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n19361), .B1(
        n19386), .B2(n19610), .ZN(n19345) );
  OAI211_X1 U22272 ( .C1(n19503), .C2(n19353), .A(n19346), .B(n19345), .ZN(
        P2_U3105) );
  AOI22_X1 U22273 ( .A1(n19359), .A2(n19614), .B1(n19358), .B2(n19613), .ZN(
        n19348) );
  AOI22_X1 U22274 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n19361), .B1(
        n19386), .B2(n19615), .ZN(n19347) );
  OAI211_X1 U22275 ( .C1(n19506), .C2(n19353), .A(n19348), .B(n19347), .ZN(
        P2_U3106) );
  AOI22_X1 U22276 ( .A1(n19359), .A2(n19620), .B1(n19358), .B2(n19619), .ZN(
        n19350) );
  AOI22_X1 U22277 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n19361), .B1(
        n19386), .B2(n19622), .ZN(n19349) );
  OAI211_X1 U22278 ( .C1(n19509), .C2(n19353), .A(n19350), .B(n19349), .ZN(
        P2_U3107) );
  AOI22_X1 U22279 ( .A1(n19359), .A2(n19627), .B1(n19358), .B2(n19626), .ZN(
        n19352) );
  AOI22_X1 U22280 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n19361), .B1(
        n19386), .B2(n19629), .ZN(n19351) );
  OAI211_X1 U22281 ( .C1(n19512), .C2(n19353), .A(n19352), .B(n19351), .ZN(
        P2_U3108) );
  AOI22_X1 U22282 ( .A1(n19359), .A2(n19633), .B1(n19358), .B2(n19632), .ZN(
        n19355) );
  AOI22_X1 U22283 ( .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n19361), .B1(
        n19360), .B2(n19634), .ZN(n19354) );
  OAI211_X1 U22284 ( .C1(n19478), .C2(n19394), .A(n19355), .B(n19354), .ZN(
        P2_U3109) );
  AOI22_X1 U22285 ( .A1(n19359), .A2(n19639), .B1(n19358), .B2(n19638), .ZN(
        n19357) );
  AOI22_X1 U22286 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n19361), .B1(
        n19360), .B2(n19641), .ZN(n19356) );
  OAI211_X1 U22287 ( .C1(n19482), .C2(n19394), .A(n19357), .B(n19356), .ZN(
        P2_U3110) );
  AOI22_X1 U22288 ( .A1(n19359), .A2(n19647), .B1(n19358), .B2(n19645), .ZN(
        n19363) );
  AOI22_X1 U22289 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n19361), .B1(
        n19360), .B2(n19649), .ZN(n19362) );
  OAI211_X1 U22290 ( .C1(n19424), .C2(n19394), .A(n19363), .B(n19362), .ZN(
        P2_U3111) );
  NAND2_X1 U22291 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n19764), .ZN(
        n19454) );
  NOR2_X1 U22292 ( .A1(n19364), .A2(n19454), .ZN(n19389) );
  AOI22_X1 U22293 ( .A1(n19603), .A2(n19419), .B1(n19600), .B2(n19389), .ZN(
        n19375) );
  NAND2_X1 U22294 ( .A1(n19394), .A2(n19752), .ZN(n19365) );
  OAI21_X1 U22295 ( .B1(n19365), .B2(n19419), .A(n19556), .ZN(n19370) );
  INV_X1 U22296 ( .A(n12132), .ZN(n19366) );
  AOI21_X1 U22297 ( .B1(n19366), .B2(n19594), .A(n19752), .ZN(n19367) );
  AOI21_X1 U22298 ( .B1(n19370), .B2(n19372), .A(n19367), .ZN(n19368) );
  INV_X1 U22299 ( .A(n19370), .ZN(n19373) );
  NOR2_X1 U22300 ( .A1(n12132), .A2(n19801), .ZN(n19369) );
  OAI22_X1 U22301 ( .A1(n19370), .A2(P2_STATE2_REG_2__SCAN_IN), .B1(n19389), 
        .B2(n19369), .ZN(n19371) );
  AOI22_X1 U22302 ( .A1(P2_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n19391), .B1(
        n19601), .B2(n19390), .ZN(n19374) );
  OAI211_X1 U22303 ( .C1(n19500), .C2(n19394), .A(n19375), .B(n19374), .ZN(
        P2_U3112) );
  AOI22_X1 U22304 ( .A1(n19610), .A2(n19419), .B1(n19389), .B2(n19607), .ZN(
        n19377) );
  AOI22_X1 U22305 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n19391), .B1(
        n19390), .B2(n19608), .ZN(n19376) );
  OAI211_X1 U22306 ( .C1(n19503), .C2(n19394), .A(n19377), .B(n19376), .ZN(
        P2_U3113) );
  AOI22_X1 U22307 ( .A1(n19386), .A2(n19616), .B1(n19613), .B2(n19389), .ZN(
        n19379) );
  AOI22_X1 U22308 ( .A1(P2_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n19391), .B1(
        n19390), .B2(n19614), .ZN(n19378) );
  OAI211_X1 U22309 ( .C1(n19471), .C2(n19418), .A(n19379), .B(n19378), .ZN(
        P2_U3114) );
  AOI22_X1 U22310 ( .A1(n19622), .A2(n19419), .B1(n19389), .B2(n19619), .ZN(
        n19381) );
  AOI22_X1 U22311 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n19391), .B1(
        n19390), .B2(n19620), .ZN(n19380) );
  OAI211_X1 U22312 ( .C1(n19509), .C2(n19394), .A(n19381), .B(n19380), .ZN(
        P2_U3115) );
  AOI22_X1 U22313 ( .A1(n19629), .A2(n19419), .B1(n19389), .B2(n19626), .ZN(
        n19383) );
  AOI22_X1 U22314 ( .A1(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n19391), .B1(
        n19390), .B2(n19627), .ZN(n19382) );
  OAI211_X1 U22315 ( .C1(n19512), .C2(n19394), .A(n19383), .B(n19382), .ZN(
        P2_U3116) );
  AOI22_X1 U22316 ( .A1(n19635), .A2(n19419), .B1(n19389), .B2(n19632), .ZN(
        n19385) );
  AOI22_X1 U22317 ( .A1(P2_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n19391), .B1(
        n19390), .B2(n19633), .ZN(n19384) );
  OAI211_X1 U22318 ( .C1(n19515), .C2(n19394), .A(n19385), .B(n19384), .ZN(
        P2_U3117) );
  AOI22_X1 U22319 ( .A1(n19386), .A2(n19641), .B1(n19389), .B2(n19638), .ZN(
        n19388) );
  AOI22_X1 U22320 ( .A1(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n19391), .B1(
        n19390), .B2(n19639), .ZN(n19387) );
  OAI211_X1 U22321 ( .C1(n19482), .C2(n19418), .A(n19388), .B(n19387), .ZN(
        P2_U3118) );
  AOI22_X1 U22322 ( .A1(n19419), .A2(n19651), .B1(n19389), .B2(n19645), .ZN(
        n19393) );
  AOI22_X1 U22323 ( .A1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n19391), .B1(
        n19390), .B2(n19647), .ZN(n19392) );
  OAI211_X1 U22324 ( .C1(n19525), .C2(n19394), .A(n19393), .B(n19392), .ZN(
        P2_U3119) );
  NOR3_X2 U22325 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19783), .A3(
        n19454), .ZN(n19428) );
  AOI22_X1 U22326 ( .A1(n19603), .A2(n19445), .B1(n19600), .B2(n19428), .ZN(
        n19405) );
  NAND2_X1 U22327 ( .A1(n19754), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19458) );
  OAI21_X1 U22328 ( .B1(n19458), .B2(n19395), .A(n19752), .ZN(n19403) );
  NOR2_X1 U22329 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19454), .ZN(
        n19399) );
  INV_X1 U22330 ( .A(n12108), .ZN(n19400) );
  OAI21_X1 U22331 ( .B1(n19400), .B2(n19801), .A(n19594), .ZN(n19397) );
  INV_X1 U22332 ( .A(n19428), .ZN(n19396) );
  AOI21_X1 U22333 ( .B1(n19397), .B2(n19396), .A(n19528), .ZN(n19398) );
  OAI21_X1 U22334 ( .B1(n19403), .B2(n19399), .A(n19398), .ZN(n19421) );
  INV_X1 U22335 ( .A(n19399), .ZN(n19402) );
  OAI21_X1 U22336 ( .B1(n19400), .B2(n19428), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19401) );
  OAI21_X1 U22337 ( .B1(n19403), .B2(n19402), .A(n19401), .ZN(n19420) );
  AOI22_X1 U22338 ( .A1(P2_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n19421), .B1(
        n19601), .B2(n19420), .ZN(n19404) );
  OAI211_X1 U22339 ( .C1(n19500), .C2(n19418), .A(n19405), .B(n19404), .ZN(
        P2_U3120) );
  AOI22_X1 U22340 ( .A1(n19610), .A2(n19445), .B1(n19428), .B2(n19607), .ZN(
        n19407) );
  AOI22_X1 U22341 ( .A1(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n19421), .B1(
        n19608), .B2(n19420), .ZN(n19406) );
  OAI211_X1 U22342 ( .C1(n19503), .C2(n19418), .A(n19407), .B(n19406), .ZN(
        P2_U3121) );
  AOI22_X1 U22343 ( .A1(n19615), .A2(n19445), .B1(n19613), .B2(n19428), .ZN(
        n19409) );
  AOI22_X1 U22344 ( .A1(P2_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n19421), .B1(
        n19614), .B2(n19420), .ZN(n19408) );
  OAI211_X1 U22345 ( .C1(n19506), .C2(n19418), .A(n19409), .B(n19408), .ZN(
        P2_U3122) );
  AOI22_X1 U22346 ( .A1(n19622), .A2(n19445), .B1(n19428), .B2(n19619), .ZN(
        n19411) );
  AOI22_X1 U22347 ( .A1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n19421), .B1(
        n19620), .B2(n19420), .ZN(n19410) );
  OAI211_X1 U22348 ( .C1(n19509), .C2(n19418), .A(n19411), .B(n19410), .ZN(
        P2_U3123) );
  AOI22_X1 U22349 ( .A1(n19629), .A2(n19445), .B1(n19428), .B2(n19626), .ZN(
        n19413) );
  AOI22_X1 U22350 ( .A1(P2_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n19421), .B1(
        n19627), .B2(n19420), .ZN(n19412) );
  OAI211_X1 U22351 ( .C1(n19512), .C2(n19418), .A(n19413), .B(n19412), .ZN(
        P2_U3124) );
  AOI22_X1 U22352 ( .A1(n19635), .A2(n19445), .B1(n19428), .B2(n19632), .ZN(
        n19415) );
  AOI22_X1 U22353 ( .A1(P2_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n19421), .B1(
        n19633), .B2(n19420), .ZN(n19414) );
  OAI211_X1 U22354 ( .C1(n19515), .C2(n19418), .A(n19415), .B(n19414), .ZN(
        P2_U3125) );
  AOI22_X1 U22355 ( .A1(n19640), .A2(n19445), .B1(n19428), .B2(n19638), .ZN(
        n19417) );
  AOI22_X1 U22356 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n19421), .B1(
        n19639), .B2(n19420), .ZN(n19416) );
  OAI211_X1 U22357 ( .C1(n19518), .C2(n19418), .A(n19417), .B(n19416), .ZN(
        P2_U3126) );
  AOI22_X1 U22358 ( .A1(n19649), .A2(n19419), .B1(n19428), .B2(n19645), .ZN(
        n19423) );
  AOI22_X1 U22359 ( .A1(P2_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n19421), .B1(
        n19647), .B2(n19420), .ZN(n19422) );
  OAI211_X1 U22360 ( .C1(n19424), .C2(n19453), .A(n19423), .B(n19422), .ZN(
        P2_U3127) );
  INV_X1 U22361 ( .A(n19425), .ZN(n19429) );
  NOR3_X2 U22362 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19773), .A3(
        n19454), .ZN(n19448) );
  OAI21_X1 U22363 ( .B1(n19429), .B2(n19448), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19426) );
  OAI21_X1 U22364 ( .B1(n19454), .B2(n19427), .A(n19426), .ZN(n19449) );
  AOI22_X1 U22365 ( .A1(n19449), .A2(n19601), .B1(n19600), .B2(n19448), .ZN(
        n19434) );
  AOI221_X1 U22366 ( .B1(n19479), .B2(P2_STATEBS16_REG_SCAN_IN), .C1(n19445), 
        .C2(P2_STATEBS16_REG_SCAN_IN), .A(n19428), .ZN(n19431) );
  OAI21_X1 U22367 ( .B1(n19429), .B2(n19801), .A(n19594), .ZN(n19430) );
  NOR2_X1 U22368 ( .A1(n19431), .A2(n19430), .ZN(n19432) );
  AOI22_X1 U22369 ( .A1(P2_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n19450), .B1(
        n19479), .B2(n19603), .ZN(n19433) );
  OAI211_X1 U22370 ( .C1(n19500), .C2(n19453), .A(n19434), .B(n19433), .ZN(
        P2_U3128) );
  AOI22_X1 U22371 ( .A1(n19449), .A2(n19608), .B1(n19607), .B2(n19448), .ZN(
        n19436) );
  AOI22_X1 U22372 ( .A1(P2_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n19450), .B1(
        n19479), .B2(n19610), .ZN(n19435) );
  OAI211_X1 U22373 ( .C1(n19503), .C2(n19453), .A(n19436), .B(n19435), .ZN(
        P2_U3129) );
  INV_X1 U22374 ( .A(n19479), .ZN(n19488) );
  AOI22_X1 U22375 ( .A1(n19449), .A2(n19614), .B1(n19613), .B2(n19448), .ZN(
        n19438) );
  AOI22_X1 U22376 ( .A1(P2_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n19450), .B1(
        n19445), .B2(n19616), .ZN(n19437) );
  OAI211_X1 U22377 ( .C1(n19471), .C2(n19488), .A(n19438), .B(n19437), .ZN(
        P2_U3130) );
  AOI22_X1 U22378 ( .A1(n19449), .A2(n19620), .B1(n19619), .B2(n19448), .ZN(
        n19440) );
  AOI22_X1 U22379 ( .A1(P2_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n19450), .B1(
        n19479), .B2(n19622), .ZN(n19439) );
  OAI211_X1 U22380 ( .C1(n19509), .C2(n19453), .A(n19440), .B(n19439), .ZN(
        P2_U3131) );
  AOI22_X1 U22381 ( .A1(n19449), .A2(n19627), .B1(n19626), .B2(n19448), .ZN(
        n19442) );
  AOI22_X1 U22382 ( .A1(P2_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n19450), .B1(
        n19479), .B2(n19629), .ZN(n19441) );
  OAI211_X1 U22383 ( .C1(n19512), .C2(n19453), .A(n19442), .B(n19441), .ZN(
        P2_U3132) );
  AOI22_X1 U22384 ( .A1(n19449), .A2(n19633), .B1(n19632), .B2(n19448), .ZN(
        n19444) );
  AOI22_X1 U22385 ( .A1(P2_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n19450), .B1(
        n19479), .B2(n19635), .ZN(n19443) );
  OAI211_X1 U22386 ( .C1(n19515), .C2(n19453), .A(n19444), .B(n19443), .ZN(
        P2_U3133) );
  AOI22_X1 U22387 ( .A1(n19449), .A2(n19639), .B1(n19638), .B2(n19448), .ZN(
        n19447) );
  AOI22_X1 U22388 ( .A1(P2_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n19450), .B1(
        n19445), .B2(n19641), .ZN(n19446) );
  OAI211_X1 U22389 ( .C1(n19482), .C2(n19488), .A(n19447), .B(n19446), .ZN(
        P2_U3134) );
  AOI22_X1 U22390 ( .A1(n19449), .A2(n19647), .B1(n19645), .B2(n19448), .ZN(
        n19452) );
  AOI22_X1 U22391 ( .A1(P2_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n19450), .B1(
        n19479), .B2(n19651), .ZN(n19451) );
  OAI211_X1 U22392 ( .C1(n19525), .C2(n19453), .A(n19452), .B(n19451), .ZN(
        P2_U3135) );
  OR2_X1 U22393 ( .A1(n19773), .A2(n19454), .ZN(n19461) );
  OR2_X1 U22394 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n19461), .ZN(n19457) );
  INV_X1 U22395 ( .A(n12125), .ZN(n19456) );
  NOR2_X1 U22396 ( .A1(n19455), .A2(n19454), .ZN(n19483) );
  NOR3_X1 U22397 ( .A1(n19456), .A2(n19801), .A3(n19483), .ZN(n19460) );
  AOI21_X1 U22398 ( .B1(n19801), .B2(n19457), .A(n19460), .ZN(n19484) );
  AOI22_X1 U22399 ( .A1(n19484), .A2(n19601), .B1(n19600), .B2(n19483), .ZN(
        n19465) );
  INV_X1 U22400 ( .A(n19458), .ZN(n19589) );
  INV_X1 U22401 ( .A(n19459), .ZN(n19748) );
  NAND2_X1 U22402 ( .A1(n19589), .A2(n19748), .ZN(n19462) );
  AOI21_X1 U22403 ( .B1(n19462), .B2(n19461), .A(n19460), .ZN(n19463) );
  OAI211_X1 U22404 ( .C1(n19483), .C2(n19594), .A(n19463), .B(n19593), .ZN(
        n19485) );
  AOI22_X1 U22405 ( .A1(P2_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n19485), .B1(
        n19479), .B2(n19602), .ZN(n19464) );
  OAI211_X1 U22406 ( .C1(n19466), .C2(n19524), .A(n19465), .B(n19464), .ZN(
        P2_U3136) );
  AOI22_X1 U22407 ( .A1(n19484), .A2(n19608), .B1(n19607), .B2(n19483), .ZN(
        n19468) );
  AOI22_X1 U22408 ( .A1(P2_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n19485), .B1(
        n19493), .B2(n19610), .ZN(n19467) );
  OAI211_X1 U22409 ( .C1(n19503), .C2(n19488), .A(n19468), .B(n19467), .ZN(
        P2_U3137) );
  AOI22_X1 U22410 ( .A1(n19484), .A2(n19614), .B1(n19613), .B2(n19483), .ZN(
        n19470) );
  AOI22_X1 U22411 ( .A1(P2_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n19485), .B1(
        n19479), .B2(n19616), .ZN(n19469) );
  OAI211_X1 U22412 ( .C1(n19471), .C2(n19524), .A(n19470), .B(n19469), .ZN(
        P2_U3138) );
  AOI22_X1 U22413 ( .A1(n19484), .A2(n19620), .B1(n19619), .B2(n19483), .ZN(
        n19473) );
  AOI22_X1 U22414 ( .A1(P2_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n19485), .B1(
        n19493), .B2(n19622), .ZN(n19472) );
  OAI211_X1 U22415 ( .C1(n19509), .C2(n19488), .A(n19473), .B(n19472), .ZN(
        P2_U3139) );
  AOI22_X1 U22416 ( .A1(n19484), .A2(n19627), .B1(n19626), .B2(n19483), .ZN(
        n19475) );
  AOI22_X1 U22417 ( .A1(P2_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n19485), .B1(
        n19493), .B2(n19629), .ZN(n19474) );
  OAI211_X1 U22418 ( .C1(n19512), .C2(n19488), .A(n19475), .B(n19474), .ZN(
        P2_U3140) );
  AOI22_X1 U22419 ( .A1(n19484), .A2(n19633), .B1(n19632), .B2(n19483), .ZN(
        n19477) );
  AOI22_X1 U22420 ( .A1(P2_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n19485), .B1(
        n19479), .B2(n19634), .ZN(n19476) );
  OAI211_X1 U22421 ( .C1(n19478), .C2(n19524), .A(n19477), .B(n19476), .ZN(
        P2_U3141) );
  AOI22_X1 U22422 ( .A1(n19484), .A2(n19639), .B1(n19638), .B2(n19483), .ZN(
        n19481) );
  AOI22_X1 U22423 ( .A1(P2_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n19485), .B1(
        n19479), .B2(n19641), .ZN(n19480) );
  OAI211_X1 U22424 ( .C1(n19482), .C2(n19524), .A(n19481), .B(n19480), .ZN(
        P2_U3142) );
  AOI22_X1 U22425 ( .A1(n19484), .A2(n19647), .B1(n19645), .B2(n19483), .ZN(
        n19487) );
  AOI22_X1 U22426 ( .A1(P2_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n19485), .B1(
        n19493), .B2(n19651), .ZN(n19486) );
  OAI211_X1 U22427 ( .C1(n19525), .C2(n19488), .A(n19487), .B(n19486), .ZN(
        P2_U3143) );
  INV_X1 U22428 ( .A(n19489), .ZN(n19492) );
  INV_X1 U22429 ( .A(n12113), .ZN(n19490) );
  NAND3_X1 U22430 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(n19773), .ZN(n19532) );
  NOR2_X1 U22431 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19532), .ZN(
        n19519) );
  OAI21_X1 U22432 ( .B1(n19490), .B2(n19519), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19491) );
  OAI21_X1 U22433 ( .B1(n19492), .B2(n19495), .A(n19491), .ZN(n19520) );
  AOI22_X1 U22434 ( .A1(n19520), .A2(n19601), .B1(n19600), .B2(n19519), .ZN(
        n19499) );
  AOI21_X1 U22435 ( .B1(n12113), .B2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n19497) );
  NOR2_X2 U22436 ( .A1(n19555), .A2(n19533), .ZN(n19550) );
  OAI21_X1 U22437 ( .B1(n19493), .B2(n19550), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19494) );
  OAI21_X1 U22438 ( .B1(n19495), .B2(n19757), .A(n19494), .ZN(n19496) );
  OAI211_X1 U22439 ( .C1(n19519), .C2(n19497), .A(n19496), .B(n19593), .ZN(
        n19521) );
  AOI22_X1 U22440 ( .A1(P2_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n19521), .B1(
        n19550), .B2(n19603), .ZN(n19498) );
  OAI211_X1 U22441 ( .C1(n19500), .C2(n19524), .A(n19499), .B(n19498), .ZN(
        P2_U3144) );
  AOI22_X1 U22442 ( .A1(n19520), .A2(n19608), .B1(n19607), .B2(n19519), .ZN(
        n19502) );
  AOI22_X1 U22443 ( .A1(P2_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n19521), .B1(
        n19550), .B2(n19610), .ZN(n19501) );
  OAI211_X1 U22444 ( .C1(n19503), .C2(n19524), .A(n19502), .B(n19501), .ZN(
        P2_U3145) );
  AOI22_X1 U22445 ( .A1(n19520), .A2(n19614), .B1(n19613), .B2(n19519), .ZN(
        n19505) );
  AOI22_X1 U22446 ( .A1(P2_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n19521), .B1(
        n19550), .B2(n19615), .ZN(n19504) );
  OAI211_X1 U22447 ( .C1(n19506), .C2(n19524), .A(n19505), .B(n19504), .ZN(
        P2_U3146) );
  AOI22_X1 U22448 ( .A1(n19520), .A2(n19620), .B1(n19619), .B2(n19519), .ZN(
        n19508) );
  AOI22_X1 U22449 ( .A1(P2_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n19521), .B1(
        n19550), .B2(n19622), .ZN(n19507) );
  OAI211_X1 U22450 ( .C1(n19509), .C2(n19524), .A(n19508), .B(n19507), .ZN(
        P2_U3147) );
  AOI22_X1 U22451 ( .A1(n19520), .A2(n19627), .B1(n19626), .B2(n19519), .ZN(
        n19511) );
  AOI22_X1 U22452 ( .A1(P2_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n19521), .B1(
        n19550), .B2(n19629), .ZN(n19510) );
  OAI211_X1 U22453 ( .C1(n19512), .C2(n19524), .A(n19511), .B(n19510), .ZN(
        P2_U3148) );
  AOI22_X1 U22454 ( .A1(n19520), .A2(n19633), .B1(n19632), .B2(n19519), .ZN(
        n19514) );
  AOI22_X1 U22455 ( .A1(P2_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n19521), .B1(
        n19550), .B2(n19635), .ZN(n19513) );
  OAI211_X1 U22456 ( .C1(n19515), .C2(n19524), .A(n19514), .B(n19513), .ZN(
        P2_U3149) );
  AOI22_X1 U22457 ( .A1(n19520), .A2(n19639), .B1(n19638), .B2(n19519), .ZN(
        n19517) );
  AOI22_X1 U22458 ( .A1(P2_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n19521), .B1(
        n19550), .B2(n19640), .ZN(n19516) );
  OAI211_X1 U22459 ( .C1(n19518), .C2(n19524), .A(n19517), .B(n19516), .ZN(
        P2_U3150) );
  AOI22_X1 U22460 ( .A1(n19520), .A2(n19647), .B1(n19645), .B2(n19519), .ZN(
        n19523) );
  AOI22_X1 U22461 ( .A1(P2_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n19521), .B1(
        n19550), .B2(n19651), .ZN(n19522) );
  OAI211_X1 U22462 ( .C1(n19525), .C2(n19524), .A(n19523), .B(n19522), .ZN(
        P2_U3151) );
  NAND2_X1 U22463 ( .A1(n19589), .A2(n19526), .ZN(n19529) );
  INV_X1 U22464 ( .A(n12117), .ZN(n19530) );
  NOR2_X1 U22465 ( .A1(n19783), .A2(n19532), .ZN(n19558) );
  AOI211_X1 U22466 ( .C1(n19530), .C2(n19594), .A(n19752), .B(n19558), .ZN(
        n19527) );
  AOI211_X2 U22467 ( .C1(n19529), .C2(n19532), .A(n19528), .B(n19527), .ZN(
        n19553) );
  OAI21_X1 U22468 ( .B1(n19530), .B2(n19558), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19531) );
  OAI21_X1 U22469 ( .B1(n19532), .B2(n19747), .A(n19531), .ZN(n19549) );
  AOI22_X1 U22470 ( .A1(n19549), .A2(n19601), .B1(n19600), .B2(n19558), .ZN(
        n19536) );
  NOR2_X2 U22471 ( .A1(n19534), .A2(n19533), .ZN(n19582) );
  AOI22_X1 U22472 ( .A1(n19582), .A2(n19603), .B1(n19550), .B2(n19602), .ZN(
        n19535) );
  OAI211_X1 U22473 ( .C1(n19553), .C2(n11641), .A(n19536), .B(n19535), .ZN(
        P2_U3152) );
  AOI22_X1 U22474 ( .A1(n19549), .A2(n19608), .B1(n19607), .B2(n19558), .ZN(
        n19538) );
  AOI22_X1 U22475 ( .A1(n19582), .A2(n19610), .B1(n19550), .B2(n19609), .ZN(
        n19537) );
  OAI211_X1 U22476 ( .C1(n19553), .C2(n12048), .A(n19538), .B(n19537), .ZN(
        P2_U3153) );
  AOI22_X1 U22477 ( .A1(n19549), .A2(n19614), .B1(n19613), .B2(n19558), .ZN(
        n19540) );
  AOI22_X1 U22478 ( .A1(n19550), .A2(n19616), .B1(n19582), .B2(n19615), .ZN(
        n19539) );
  OAI211_X1 U22479 ( .C1(n19553), .C2(n11688), .A(n19540), .B(n19539), .ZN(
        P2_U3154) );
  AOI22_X1 U22480 ( .A1(n19549), .A2(n19620), .B1(n19619), .B2(n19558), .ZN(
        n19542) );
  AOI22_X1 U22481 ( .A1(n19582), .A2(n19622), .B1(n19550), .B2(n19621), .ZN(
        n19541) );
  OAI211_X1 U22482 ( .C1(n19553), .C2(n12092), .A(n19542), .B(n19541), .ZN(
        P2_U3155) );
  AOI22_X1 U22483 ( .A1(n19549), .A2(n19627), .B1(n19626), .B2(n19558), .ZN(
        n19544) );
  AOI22_X1 U22484 ( .A1(n19582), .A2(n19629), .B1(n19550), .B2(n19628), .ZN(
        n19543) );
  OAI211_X1 U22485 ( .C1(n19553), .C2(n11732), .A(n19544), .B(n19543), .ZN(
        P2_U3156) );
  AOI22_X1 U22486 ( .A1(n19549), .A2(n19633), .B1(n19632), .B2(n19558), .ZN(
        n19546) );
  AOI22_X1 U22487 ( .A1(n19582), .A2(n19635), .B1(n19550), .B2(n19634), .ZN(
        n19545) );
  OAI211_X1 U22488 ( .C1(n19553), .C2(n12118), .A(n19546), .B(n19545), .ZN(
        P2_U3157) );
  AOI22_X1 U22489 ( .A1(n19549), .A2(n19639), .B1(n19638), .B2(n19558), .ZN(
        n19548) );
  AOI22_X1 U22490 ( .A1(n19550), .A2(n19641), .B1(n19582), .B2(n19640), .ZN(
        n19547) );
  OAI211_X1 U22491 ( .C1(n19553), .C2(n12181), .A(n19548), .B(n19547), .ZN(
        P2_U3158) );
  AOI22_X1 U22492 ( .A1(n19549), .A2(n19647), .B1(n19645), .B2(n19558), .ZN(
        n19552) );
  AOI22_X1 U22493 ( .A1(n19582), .A2(n19651), .B1(n19550), .B2(n19649), .ZN(
        n19551) );
  OAI211_X1 U22494 ( .C1(n19553), .C2(n11785), .A(n19552), .B(n19551), .ZN(
        P2_U3159) );
  INV_X1 U22495 ( .A(n19582), .ZN(n19554) );
  NAND2_X1 U22496 ( .A1(n19554), .A2(n19752), .ZN(n19557) );
  NOR2_X2 U22497 ( .A1(n19555), .A2(n19587), .ZN(n19650) );
  OAI21_X1 U22498 ( .B1(n19557), .B2(n19650), .A(n19556), .ZN(n19561) );
  NOR3_X2 U22499 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19757), .A3(
        n19590), .ZN(n19581) );
  NOR2_X1 U22500 ( .A1(n19581), .A2(n19558), .ZN(n19564) );
  AOI21_X1 U22501 ( .B1(n12114), .B2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n19559) );
  OAI21_X1 U22502 ( .B1(n19559), .B2(n19581), .A(n19593), .ZN(n19560) );
  AOI22_X1 U22503 ( .A1(n19603), .A2(n19650), .B1(n19600), .B2(n19581), .ZN(
        n19567) );
  INV_X1 U22504 ( .A(n19561), .ZN(n19565) );
  INV_X1 U22505 ( .A(n12114), .ZN(n19562) );
  OAI21_X1 U22506 ( .B1(n19562), .B2(n19581), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19563) );
  AOI22_X1 U22507 ( .A1(n19601), .A2(n19583), .B1(n19582), .B2(n19602), .ZN(
        n19566) );
  OAI211_X1 U22508 ( .C1(n19586), .C2(n19568), .A(n19567), .B(n19566), .ZN(
        P2_U3160) );
  AOI22_X1 U22509 ( .A1(n19610), .A2(n19650), .B1(n19581), .B2(n19607), .ZN(
        n19570) );
  AOI22_X1 U22510 ( .A1(n19608), .A2(n19583), .B1(n19582), .B2(n19609), .ZN(
        n19569) );
  OAI211_X1 U22511 ( .C1(n19586), .C2(n12046), .A(n19570), .B(n19569), .ZN(
        P2_U3161) );
  AOI22_X1 U22512 ( .A1(n19615), .A2(n19650), .B1(n19613), .B2(n19581), .ZN(
        n19572) );
  AOI22_X1 U22513 ( .A1(n19614), .A2(n19583), .B1(n19582), .B2(n19616), .ZN(
        n19571) );
  OAI211_X1 U22514 ( .C1(n19586), .C2(n11843), .A(n19572), .B(n19571), .ZN(
        P2_U3162) );
  AOI22_X1 U22515 ( .A1(n19621), .A2(n19582), .B1(n19581), .B2(n19619), .ZN(
        n19574) );
  AOI22_X1 U22516 ( .A1(n19620), .A2(n19583), .B1(n19650), .B2(n19622), .ZN(
        n19573) );
  OAI211_X1 U22517 ( .C1(n19586), .C2(n12090), .A(n19574), .B(n19573), .ZN(
        P2_U3163) );
  AOI22_X1 U22518 ( .A1(n19628), .A2(n19582), .B1(n19581), .B2(n19626), .ZN(
        n19576) );
  AOI22_X1 U22519 ( .A1(n19627), .A2(n19583), .B1(n19650), .B2(n19629), .ZN(
        n19575) );
  OAI211_X1 U22520 ( .C1(n19586), .C2(n11879), .A(n19576), .B(n19575), .ZN(
        P2_U3164) );
  AOI22_X1 U22521 ( .A1(n19634), .A2(n19582), .B1(n19581), .B2(n19632), .ZN(
        n19578) );
  AOI22_X1 U22522 ( .A1(n19633), .A2(n19583), .B1(n19650), .B2(n19635), .ZN(
        n19577) );
  OAI211_X1 U22523 ( .C1(n19586), .C2(n12115), .A(n19578), .B(n19577), .ZN(
        P2_U3165) );
  AOI22_X1 U22524 ( .A1(n19582), .A2(n19641), .B1(n19581), .B2(n19638), .ZN(
        n19580) );
  AOI22_X1 U22525 ( .A1(n19639), .A2(n19583), .B1(n19650), .B2(n19640), .ZN(
        n19579) );
  OAI211_X1 U22526 ( .C1(n19586), .C2(n12172), .A(n19580), .B(n19579), .ZN(
        P2_U3166) );
  AOI22_X1 U22527 ( .A1(n19649), .A2(n19582), .B1(n19581), .B2(n19645), .ZN(
        n19585) );
  AOI22_X1 U22528 ( .A1(n19647), .A2(n19583), .B1(n19650), .B2(n19651), .ZN(
        n19584) );
  OAI211_X1 U22529 ( .C1(n19586), .C2(n11931), .A(n19585), .B(n19584), .ZN(
        P2_U3167) );
  INV_X1 U22530 ( .A(n19587), .ZN(n19588) );
  NAND2_X1 U22531 ( .A1(n19589), .A2(n19588), .ZN(n19596) );
  OR2_X1 U22532 ( .A1(n19757), .A2(n19590), .ZN(n19597) );
  INV_X1 U22533 ( .A(n19591), .ZN(n19646) );
  AND2_X1 U22534 ( .A1(n19591), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n19592) );
  NAND2_X1 U22535 ( .A1(n9673), .A2(n19592), .ZN(n19599) );
  OAI211_X1 U22536 ( .C1(n19646), .C2(n19594), .A(n19599), .B(n19593), .ZN(
        n19595) );
  OAI21_X1 U22537 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n19597), .A(n19801), 
        .ZN(n19598) );
  AND2_X1 U22538 ( .A1(n19599), .A2(n19598), .ZN(n19648) );
  AOI22_X1 U22539 ( .A1(n19648), .A2(n19601), .B1(n19646), .B2(n19600), .ZN(
        n19605) );
  AOI22_X1 U22540 ( .A1(n19652), .A2(n19603), .B1(n19650), .B2(n19602), .ZN(
        n19604) );
  OAI211_X1 U22541 ( .C1(n19656), .C2(n19606), .A(n19605), .B(n19604), .ZN(
        P2_U3168) );
  AOI22_X1 U22542 ( .A1(n19648), .A2(n19608), .B1(n19646), .B2(n19607), .ZN(
        n19612) );
  AOI22_X1 U22543 ( .A1(n19652), .A2(n19610), .B1(n19650), .B2(n19609), .ZN(
        n19611) );
  OAI211_X1 U22544 ( .C1(n19656), .C2(n12568), .A(n19612), .B(n19611), .ZN(
        P2_U3169) );
  AOI22_X1 U22545 ( .A1(n19648), .A2(n19614), .B1(n19646), .B2(n19613), .ZN(
        n19618) );
  AOI22_X1 U22546 ( .A1(n19650), .A2(n19616), .B1(n19652), .B2(n19615), .ZN(
        n19617) );
  OAI211_X1 U22547 ( .C1(n19656), .C2(n12585), .A(n19618), .B(n19617), .ZN(
        P2_U3170) );
  INV_X1 U22548 ( .A(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n19625) );
  AOI22_X1 U22549 ( .A1(n19648), .A2(n19620), .B1(n19646), .B2(n19619), .ZN(
        n19624) );
  AOI22_X1 U22550 ( .A1(n19652), .A2(n19622), .B1(n19650), .B2(n19621), .ZN(
        n19623) );
  OAI211_X1 U22551 ( .C1(n19656), .C2(n19625), .A(n19624), .B(n19623), .ZN(
        P2_U3171) );
  AOI22_X1 U22552 ( .A1(n19648), .A2(n19627), .B1(n19646), .B2(n19626), .ZN(
        n19631) );
  AOI22_X1 U22553 ( .A1(n19652), .A2(n19629), .B1(n19650), .B2(n19628), .ZN(
        n19630) );
  OAI211_X1 U22554 ( .C1(n19656), .C2(n12617), .A(n19631), .B(n19630), .ZN(
        P2_U3172) );
  AOI22_X1 U22555 ( .A1(n19648), .A2(n19633), .B1(n19646), .B2(n19632), .ZN(
        n19637) );
  AOI22_X1 U22556 ( .A1(n19652), .A2(n19635), .B1(n19650), .B2(n19634), .ZN(
        n19636) );
  OAI211_X1 U22557 ( .C1(n19656), .C2(n12635), .A(n19637), .B(n19636), .ZN(
        P2_U3173) );
  INV_X1 U22558 ( .A(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n19644) );
  AOI22_X1 U22559 ( .A1(n19648), .A2(n19639), .B1(n19646), .B2(n19638), .ZN(
        n19643) );
  AOI22_X1 U22560 ( .A1(n19650), .A2(n19641), .B1(n19652), .B2(n19640), .ZN(
        n19642) );
  OAI211_X1 U22561 ( .C1(n19656), .C2(n19644), .A(n19643), .B(n19642), .ZN(
        P2_U3174) );
  AOI22_X1 U22562 ( .A1(n19648), .A2(n19647), .B1(n19646), .B2(n19645), .ZN(
        n19654) );
  AOI22_X1 U22563 ( .A1(n19652), .A2(n19651), .B1(n19650), .B2(n19649), .ZN(
        n19653) );
  OAI211_X1 U22564 ( .C1(n19656), .C2(n19655), .A(n19654), .B(n19653), .ZN(
        P2_U3175) );
  INV_X1 U22565 ( .A(n19657), .ZN(n19662) );
  INV_X1 U22566 ( .A(n19658), .ZN(n19661) );
  NAND2_X1 U22567 ( .A1(n19807), .A2(n19801), .ZN(n19660) );
  NAND4_X1 U22568 ( .A1(n19662), .A2(n19661), .A3(n19660), .A4(n19659), .ZN(
        n19663) );
  OAI221_X1 U22569 ( .B1(n13649), .B2(n19665), .C1(n13649), .C2(n19664), .A(
        n19663), .ZN(P2_U3177) );
  AND2_X1 U22570 ( .A1(P2_DATAWIDTH_REG_31__SCAN_IN), .A2(n19666), .ZN(
        P2_U3179) );
  AND2_X1 U22571 ( .A1(P2_DATAWIDTH_REG_30__SCAN_IN), .A2(n19666), .ZN(
        P2_U3180) );
  AND2_X1 U22572 ( .A1(P2_DATAWIDTH_REG_29__SCAN_IN), .A2(n19666), .ZN(
        P2_U3181) );
  AND2_X1 U22573 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(n19666), .ZN(
        P2_U3182) );
  AND2_X1 U22574 ( .A1(P2_DATAWIDTH_REG_27__SCAN_IN), .A2(n19666), .ZN(
        P2_U3183) );
  AND2_X1 U22575 ( .A1(P2_DATAWIDTH_REG_26__SCAN_IN), .A2(n19666), .ZN(
        P2_U3184) );
  AND2_X1 U22576 ( .A1(P2_DATAWIDTH_REG_25__SCAN_IN), .A2(n19666), .ZN(
        P2_U3185) );
  AND2_X1 U22577 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(n19666), .ZN(
        P2_U3186) );
  AND2_X1 U22578 ( .A1(P2_DATAWIDTH_REG_23__SCAN_IN), .A2(n19666), .ZN(
        P2_U3187) );
  AND2_X1 U22579 ( .A1(P2_DATAWIDTH_REG_22__SCAN_IN), .A2(n19666), .ZN(
        P2_U3188) );
  AND2_X1 U22580 ( .A1(P2_DATAWIDTH_REG_21__SCAN_IN), .A2(n19666), .ZN(
        P2_U3189) );
  NOR2_X1 U22581 ( .A1(n20737), .A2(n19746), .ZN(P2_U3190) );
  AND2_X1 U22582 ( .A1(P2_DATAWIDTH_REG_19__SCAN_IN), .A2(n19666), .ZN(
        P2_U3191) );
  AND2_X1 U22583 ( .A1(P2_DATAWIDTH_REG_18__SCAN_IN), .A2(n19666), .ZN(
        P2_U3192) );
  AND2_X1 U22584 ( .A1(P2_DATAWIDTH_REG_17__SCAN_IN), .A2(n19666), .ZN(
        P2_U3193) );
  AND2_X1 U22585 ( .A1(P2_DATAWIDTH_REG_16__SCAN_IN), .A2(n19666), .ZN(
        P2_U3194) );
  INV_X1 U22586 ( .A(P2_DATAWIDTH_REG_15__SCAN_IN), .ZN(n20868) );
  NOR2_X1 U22587 ( .A1(n20868), .A2(n19746), .ZN(P2_U3195) );
  AND2_X1 U22588 ( .A1(P2_DATAWIDTH_REG_14__SCAN_IN), .A2(n19666), .ZN(
        P2_U3196) );
  AND2_X1 U22589 ( .A1(P2_DATAWIDTH_REG_13__SCAN_IN), .A2(n19666), .ZN(
        P2_U3197) );
  AND2_X1 U22590 ( .A1(P2_DATAWIDTH_REG_12__SCAN_IN), .A2(n19666), .ZN(
        P2_U3198) );
  AND2_X1 U22591 ( .A1(P2_DATAWIDTH_REG_11__SCAN_IN), .A2(n19666), .ZN(
        P2_U3199) );
  AND2_X1 U22592 ( .A1(P2_DATAWIDTH_REG_10__SCAN_IN), .A2(n19666), .ZN(
        P2_U3200) );
  AND2_X1 U22593 ( .A1(P2_DATAWIDTH_REG_9__SCAN_IN), .A2(n19666), .ZN(P2_U3201) );
  AND2_X1 U22594 ( .A1(P2_DATAWIDTH_REG_8__SCAN_IN), .A2(n19666), .ZN(P2_U3202) );
  AND2_X1 U22595 ( .A1(P2_DATAWIDTH_REG_7__SCAN_IN), .A2(n19666), .ZN(P2_U3203) );
  AND2_X1 U22596 ( .A1(P2_DATAWIDTH_REG_6__SCAN_IN), .A2(n19666), .ZN(P2_U3204) );
  AND2_X1 U22597 ( .A1(P2_DATAWIDTH_REG_5__SCAN_IN), .A2(n19666), .ZN(P2_U3205) );
  AND2_X1 U22598 ( .A1(P2_DATAWIDTH_REG_4__SCAN_IN), .A2(n19666), .ZN(P2_U3206) );
  NOR2_X1 U22599 ( .A1(n20807), .A2(n19746), .ZN(P2_U3207) );
  AND2_X1 U22600 ( .A1(P2_DATAWIDTH_REG_2__SCAN_IN), .A2(n19666), .ZN(P2_U3208) );
  NAND2_X1 U22601 ( .A1(n19807), .A2(P2_STATE_REG_1__SCAN_IN), .ZN(n19677) );
  NAND3_X1 U22602 ( .A1(P2_REQUESTPENDING_REG_SCAN_IN), .A2(
        P2_STATE_REG_0__SCAN_IN), .A3(n19677), .ZN(n19669) );
  AOI211_X1 U22603 ( .C1(P2_REQUESTPENDING_REG_SCAN_IN), .C2(n20601), .A(
        n19667), .B(n19815), .ZN(n19668) );
  NOR3_X1 U22604 ( .A1(P2_STATE_REG_0__SCAN_IN), .A2(P2_STATE_REG_1__SCAN_IN), 
        .A3(n20612), .ZN(n19682) );
  AOI211_X1 U22605 ( .C1(n19683), .C2(n19669), .A(n19668), .B(n19682), .ZN(
        n19670) );
  INV_X1 U22606 ( .A(n19670), .ZN(P2_U3209) );
  AOI21_X1 U22607 ( .B1(P2_STATE_REG_0__SCAN_IN), .B2(n20601), .A(n19683), 
        .ZN(n19675) );
  NOR2_X1 U22608 ( .A1(n18713), .A2(n19675), .ZN(n19671) );
  AOI21_X1 U22609 ( .B1(n19671), .B2(P2_REQUESTPENDING_REG_SCAN_IN), .A(n19795), .ZN(n19672) );
  OAI211_X1 U22610 ( .C1(n20601), .C2(n19673), .A(n19672), .B(n19677), .ZN(
        P2_U3210) );
  NOR2_X1 U22611 ( .A1(n19674), .A2(n19683), .ZN(n19676) );
  AOI21_X1 U22612 ( .B1(n19676), .B2(n19807), .A(n19675), .ZN(n19681) );
  OAI22_X1 U22613 ( .A1(P2_REQUESTPENDING_REG_SCAN_IN), .A2(n19678), .B1(NA), 
        .B2(n19677), .ZN(n19679) );
  OAI211_X1 U22614 ( .C1(P2_REQUESTPENDING_REG_SCAN_IN), .C2(HOLD), .A(
        P2_STATE_REG_0__SCAN_IN), .B(n19679), .ZN(n19680) );
  OAI21_X1 U22615 ( .B1(n19682), .B2(n19681), .A(n19680), .ZN(P2_U3211) );
  OAI222_X1 U22616 ( .A1(n19733), .A2(n19685), .B1(n19684), .B2(n19815), .C1(
        n13015), .C2(n19736), .ZN(P2_U3212) );
  OAI222_X1 U22617 ( .A1(n19733), .A2(n13015), .B1(n19686), .B2(n19815), .C1(
        n11505), .C2(n19736), .ZN(P2_U3213) );
  OAI222_X1 U22618 ( .A1(n19733), .A2(n11505), .B1(n19687), .B2(n19815), .C1(
        n19688), .C2(n19736), .ZN(P2_U3214) );
  OAI222_X1 U22619 ( .A1(n19736), .A2(n13678), .B1(n19689), .B2(n19815), .C1(
        n19688), .C2(n19733), .ZN(P2_U3215) );
  OAI222_X1 U22620 ( .A1(n19736), .A2(n11526), .B1(n19690), .B2(n19815), .C1(
        n13678), .C2(n19733), .ZN(P2_U3216) );
  OAI222_X1 U22621 ( .A1(n19736), .A2(n19692), .B1(n19691), .B2(n19815), .C1(
        n11526), .C2(n19733), .ZN(P2_U3217) );
  OAI222_X1 U22622 ( .A1(n19736), .A2(n19694), .B1(n19693), .B2(n19815), .C1(
        n19692), .C2(n19733), .ZN(P2_U3218) );
  INV_X1 U22623 ( .A(P2_REIP_REG_9__SCAN_IN), .ZN(n19696) );
  OAI222_X1 U22624 ( .A1(n19736), .A2(n19696), .B1(n19695), .B2(n19815), .C1(
        n19694), .C2(n19733), .ZN(P2_U3219) );
  OAI222_X1 U22625 ( .A1(n19736), .A2(n19698), .B1(n19697), .B2(n19815), .C1(
        n19696), .C2(n19733), .ZN(P2_U3220) );
  OAI222_X1 U22626 ( .A1(n19736), .A2(n14989), .B1(n19699), .B2(n19815), .C1(
        n19698), .C2(n19733), .ZN(P2_U3221) );
  INV_X1 U22627 ( .A(P2_REIP_REG_12__SCAN_IN), .ZN(n19701) );
  OAI222_X1 U22628 ( .A1(n19736), .A2(n19701), .B1(n19700), .B2(n19815), .C1(
        n14989), .C2(n19733), .ZN(P2_U3222) );
  OAI222_X1 U22629 ( .A1(n19736), .A2(n19703), .B1(n19702), .B2(n19815), .C1(
        n19701), .C2(n19733), .ZN(P2_U3223) );
  OAI222_X1 U22630 ( .A1(n19736), .A2(n19705), .B1(n19704), .B2(n19815), .C1(
        n19703), .C2(n19733), .ZN(P2_U3224) );
  OAI222_X1 U22631 ( .A1(n19736), .A2(n11422), .B1(n20739), .B2(n19815), .C1(
        n19705), .C2(n19733), .ZN(P2_U3225) );
  INV_X1 U22632 ( .A(P2_REIP_REG_16__SCAN_IN), .ZN(n19707) );
  OAI222_X1 U22633 ( .A1(n19736), .A2(n19707), .B1(n19706), .B2(n19815), .C1(
        n11422), .C2(n19733), .ZN(P2_U3226) );
  OAI222_X1 U22634 ( .A1(n19736), .A2(n19709), .B1(n19708), .B2(n19815), .C1(
        n19707), .C2(n19733), .ZN(P2_U3227) );
  OAI222_X1 U22635 ( .A1(n19736), .A2(n19711), .B1(n19710), .B2(n19815), .C1(
        n19709), .C2(n19733), .ZN(P2_U3228) );
  OAI222_X1 U22636 ( .A1(n19736), .A2(n19713), .B1(n19712), .B2(n19815), .C1(
        n19711), .C2(n19733), .ZN(P2_U3229) );
  OAI222_X1 U22637 ( .A1(n19736), .A2(n19715), .B1(n19714), .B2(n19815), .C1(
        n19713), .C2(n19733), .ZN(P2_U3230) );
  OAI222_X1 U22638 ( .A1(n19736), .A2(n19717), .B1(n19716), .B2(n19815), .C1(
        n19715), .C2(n19733), .ZN(P2_U3231) );
  INV_X1 U22639 ( .A(P2_REIP_REG_22__SCAN_IN), .ZN(n19719) );
  OAI222_X1 U22640 ( .A1(n19736), .A2(n19719), .B1(n19718), .B2(n19815), .C1(
        n19717), .C2(n19733), .ZN(P2_U3232) );
  OAI222_X1 U22641 ( .A1(n19736), .A2(n11581), .B1(n19720), .B2(n19815), .C1(
        n19719), .C2(n19733), .ZN(P2_U3233) );
  INV_X1 U22642 ( .A(P2_REIP_REG_24__SCAN_IN), .ZN(n19722) );
  OAI222_X1 U22643 ( .A1(n19736), .A2(n19722), .B1(n19721), .B2(n19815), .C1(
        n11581), .C2(n19733), .ZN(P2_U3234) );
  OAI222_X1 U22644 ( .A1(n19736), .A2(n19724), .B1(n19723), .B2(n19815), .C1(
        n19722), .C2(n19733), .ZN(P2_U3235) );
  OAI222_X1 U22645 ( .A1(n19736), .A2(n11593), .B1(n19725), .B2(n19815), .C1(
        n19724), .C2(n19733), .ZN(P2_U3236) );
  OAI222_X1 U22646 ( .A1(n19736), .A2(n19728), .B1(n19726), .B2(n19815), .C1(
        n11593), .C2(n19733), .ZN(P2_U3237) );
  OAI222_X1 U22647 ( .A1(n19733), .A2(n19728), .B1(n19727), .B2(n19815), .C1(
        n19729), .C2(n19736), .ZN(P2_U3238) );
  OAI222_X1 U22648 ( .A1(n19736), .A2(n19731), .B1(n19730), .B2(n19815), .C1(
        n19729), .C2(n19733), .ZN(P2_U3239) );
  OAI222_X1 U22649 ( .A1(n19736), .A2(n12008), .B1(n19732), .B2(n19815), .C1(
        n19731), .C2(n19733), .ZN(P2_U3240) );
  INV_X1 U22650 ( .A(P2_REIP_REG_31__SCAN_IN), .ZN(n19735) );
  OAI222_X1 U22651 ( .A1(n19736), .A2(n19735), .B1(n19734), .B2(n19815), .C1(
        n12008), .C2(n19733), .ZN(P2_U3241) );
  INV_X1 U22652 ( .A(P2_BE_N_REG_3__SCAN_IN), .ZN(n19737) );
  AOI22_X1 U22653 ( .A1(n19815), .A2(n19738), .B1(n19737), .B2(n19812), .ZN(
        P2_U3585) );
  MUX2_X1 U22654 ( .A(P2_BE_N_REG_2__SCAN_IN), .B(P2_BYTEENABLE_REG_2__SCAN_IN), .S(n19815), .Z(P2_U3586) );
  INV_X1 U22655 ( .A(P2_BE_N_REG_1__SCAN_IN), .ZN(n19739) );
  AOI22_X1 U22656 ( .A1(n19815), .A2(n19740), .B1(n19739), .B2(n19812), .ZN(
        P2_U3587) );
  AOI22_X1 U22657 ( .A1(n19815), .A2(n19742), .B1(n19741), .B2(n19812), .ZN(
        P2_U3588) );
  OAI21_X1 U22658 ( .B1(n19746), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .A(n19744), 
        .ZN(n19743) );
  INV_X1 U22659 ( .A(n19743), .ZN(P2_U3591) );
  OAI21_X1 U22660 ( .B1(n19746), .B2(n19745), .A(n19744), .ZN(P2_U3592) );
  NOR2_X1 U22661 ( .A1(n19747), .A2(n19221), .ZN(n19769) );
  NAND2_X1 U22662 ( .A1(n19748), .A2(n19769), .ZN(n19758) );
  NAND3_X1 U22663 ( .A1(n19767), .A2(n19749), .A3(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19750) );
  NAND2_X1 U22664 ( .A1(n19750), .A2(n19765), .ZN(n19759) );
  NAND2_X1 U22665 ( .A1(n19758), .A2(n19759), .ZN(n19755) );
  AOI222_X1 U22666 ( .A1(n19755), .A2(n19754), .B1(P2_STATE2_REG_3__SCAN_IN), 
        .B2(n19753), .C1(n19752), .C2(n19751), .ZN(n19756) );
  AOI22_X1 U22667 ( .A1(n19774), .A2(n19757), .B1(n19756), .B2(n19784), .ZN(
        P2_U3602) );
  OAI21_X1 U22668 ( .B1(n19760), .B2(n19759), .A(n19758), .ZN(n19761) );
  AOI21_X1 U22669 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n19762), .A(n19761), 
        .ZN(n19763) );
  AOI22_X1 U22670 ( .A1(n19774), .A2(n19764), .B1(n19763), .B2(n19784), .ZN(
        P2_U3603) );
  INV_X1 U22671 ( .A(n19765), .ZN(n19778) );
  NOR2_X1 U22672 ( .A1(n19778), .A2(n19766), .ZN(n19768) );
  MUX2_X1 U22673 ( .A(n19769), .B(n19768), .S(n19767), .Z(n19770) );
  AOI21_X1 U22674 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n19771), .A(n19770), 
        .ZN(n19772) );
  AOI22_X1 U22675 ( .A1(n19774), .A2(n19773), .B1(n19772), .B2(n19784), .ZN(
        P2_U3604) );
  INV_X1 U22676 ( .A(n19775), .ZN(n19777) );
  OAI22_X1 U22677 ( .A1(n19779), .A2(n19778), .B1(n19777), .B2(n19776), .ZN(
        n19781) );
  OAI21_X1 U22678 ( .B1(n19781), .B2(n19780), .A(n19784), .ZN(n19782) );
  OAI21_X1 U22679 ( .B1(n19784), .B2(n19783), .A(n19782), .ZN(P2_U3605) );
  AOI22_X1 U22680 ( .A1(n19815), .A2(P2_READREQUEST_REG_SCAN_IN), .B1(n19785), 
        .B2(n19812), .ZN(P2_U3608) );
  INV_X1 U22681 ( .A(n19786), .ZN(n19787) );
  NAND2_X1 U22682 ( .A1(n19788), .A2(n19787), .ZN(n19789) );
  OAI211_X1 U22683 ( .C1(n19792), .C2(n19791), .A(n19790), .B(n19789), .ZN(
        n19794) );
  MUX2_X1 U22684 ( .A(P2_MORE_REG_SCAN_IN), .B(n19794), .S(n19793), .Z(
        P2_U3609) );
  OAI21_X1 U22685 ( .B1(n19796), .B2(P2_STATEBS16_REG_SCAN_IN), .A(n19795), 
        .ZN(n19797) );
  NAND3_X1 U22686 ( .A1(n19798), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(n19797), 
        .ZN(n19803) );
  INV_X1 U22687 ( .A(n19799), .ZN(n19800) );
  OAI21_X1 U22688 ( .B1(n19807), .B2(n19801), .A(n19800), .ZN(n19802) );
  NAND2_X1 U22689 ( .A1(n19803), .A2(n19802), .ZN(n19811) );
  INV_X1 U22690 ( .A(n19804), .ZN(n19805) );
  OAI21_X1 U22691 ( .B1(n19807), .B2(n19806), .A(n19805), .ZN(n19808) );
  AOI21_X1 U22692 ( .B1(n19594), .B2(n19809), .A(n19808), .ZN(n19810) );
  MUX2_X1 U22693 ( .A(n19811), .B(P2_REQUESTPENDING_REG_SCAN_IN), .S(n19810), 
        .Z(P2_U3610) );
  INV_X1 U22694 ( .A(P2_M_IO_N_REG_SCAN_IN), .ZN(n19813) );
  AOI22_X1 U22695 ( .A1(n19815), .A2(n19814), .B1(n19813), .B2(n19812), .ZN(
        P2_U3611) );
  AND2_X1 U22696 ( .A1(n20606), .A2(P1_STATE_REG_0__SCAN_IN), .ZN(n19817) );
  INV_X1 U22697 ( .A(P1_ADS_N_REG_SCAN_IN), .ZN(n19816) );
  OR2_X1 U22698 ( .A1(P1_STATE_REG_0__SCAN_IN), .A2(n20609), .ZN(n20715) );
  INV_X2 U22699 ( .A(n20715), .ZN(n20733) );
  AOI21_X1 U22700 ( .B1(n19817), .B2(n19816), .A(n20733), .ZN(P1_U2802) );
  INV_X1 U22701 ( .A(n19818), .ZN(n19819) );
  OAI21_X1 U22702 ( .B1(n19820), .B2(n19819), .A(P1_CODEFETCH_REG_SCAN_IN), 
        .ZN(n19821) );
  OAI21_X1 U22703 ( .B1(P1_STATE2_REG_2__SCAN_IN), .B2(n19822), .A(n19821), 
        .ZN(P1_U2803) );
  NOR2_X1 U22704 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(P1_STATE_REG_0__SCAN_IN), 
        .ZN(n19824) );
  OAI21_X1 U22705 ( .B1(n19824), .B2(P1_D_C_N_REG_SCAN_IN), .A(n20715), .ZN(
        n19823) );
  OAI21_X1 U22706 ( .B1(P1_CODEFETCH_REG_SCAN_IN), .B2(n20715), .A(n19823), 
        .ZN(P1_U2804) );
  AOI21_X1 U22707 ( .B1(P1_STATE_REG_0__SCAN_IN), .B2(n20606), .A(n20733), 
        .ZN(n20680) );
  OAI21_X1 U22708 ( .B1(BS16), .B2(n19824), .A(n20680), .ZN(n20678) );
  OAI21_X1 U22709 ( .B1(n20680), .B2(n20891), .A(n20678), .ZN(P1_U2805) );
  NAND2_X1 U22710 ( .A1(n19826), .A2(n19825), .ZN(n20718) );
  INV_X1 U22711 ( .A(n20718), .ZN(n20721) );
  OAI21_X1 U22712 ( .B1(n20721), .B2(n19827), .A(n20031), .ZN(P1_U2806) );
  NOR4_X1 U22713 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_21__SCAN_IN), .A3(P1_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_23__SCAN_IN), .ZN(n19831) );
  NOR4_X1 U22714 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_17__SCAN_IN), .A3(P1_DATAWIDTH_REG_18__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_19__SCAN_IN), .ZN(n19830) );
  NOR4_X1 U22715 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_29__SCAN_IN), .A3(P1_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_31__SCAN_IN), .ZN(n19829) );
  NOR4_X1 U22716 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_25__SCAN_IN), .A3(P1_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_27__SCAN_IN), .ZN(n19828) );
  NAND4_X1 U22717 ( .A1(n19831), .A2(n19830), .A3(n19829), .A4(n19828), .ZN(
        n19837) );
  NOR4_X1 U22718 ( .A1(P1_DATAWIDTH_REG_3__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_4__SCAN_IN), .A3(P1_DATAWIDTH_REG_5__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_6__SCAN_IN), .ZN(n19835) );
  AOI211_X1 U22719 ( .C1(P1_DATAWIDTH_REG_1__SCAN_IN), .C2(
        P1_DATAWIDTH_REG_0__SCAN_IN), .A(P1_DATAWIDTH_REG_8__SCAN_IN), .B(
        P1_DATAWIDTH_REG_2__SCAN_IN), .ZN(n19834) );
  NOR4_X1 U22720 ( .A1(P1_DATAWIDTH_REG_12__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_13__SCAN_IN), .A3(P1_DATAWIDTH_REG_14__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_15__SCAN_IN), .ZN(n19833) );
  NOR4_X1 U22721 ( .A1(P1_DATAWIDTH_REG_7__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_9__SCAN_IN), .A3(P1_DATAWIDTH_REG_10__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_11__SCAN_IN), .ZN(n19832) );
  NAND4_X1 U22722 ( .A1(n19835), .A2(n19834), .A3(n19833), .A4(n19832), .ZN(
        n19836) );
  NOR2_X1 U22723 ( .A1(n19837), .A2(n19836), .ZN(n20714) );
  INV_X1 U22724 ( .A(P1_BYTEENABLE_REG_1__SCAN_IN), .ZN(n20673) );
  NOR3_X1 U22725 ( .A1(P1_REIP_REG_0__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .A3(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n19839) );
  OAI21_X1 U22726 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(n19839), .A(n20714), .ZN(
        n19838) );
  OAI21_X1 U22727 ( .B1(n20714), .B2(n20673), .A(n19838), .ZN(P1_U2807) );
  INV_X1 U22728 ( .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(n20679) );
  AOI21_X1 U22729 ( .B1(n20707), .B2(n20679), .A(n19839), .ZN(n19840) );
  INV_X1 U22730 ( .A(P1_BYTEENABLE_REG_3__SCAN_IN), .ZN(n20670) );
  INV_X1 U22731 ( .A(n20714), .ZN(n20709) );
  AOI22_X1 U22732 ( .A1(n20714), .A2(n19840), .B1(n20670), .B2(n20709), .ZN(
        P1_U2808) );
  AOI22_X1 U22733 ( .A1(n19841), .A2(n19905), .B1(n19929), .B2(
        P1_EBX_REG_9__SCAN_IN), .ZN(n19850) );
  AOI21_X1 U22734 ( .B1(n19935), .B2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .A(
        n19891), .ZN(n19849) );
  AOI22_X1 U22735 ( .A1(n19843), .A2(n19872), .B1(n19934), .B2(n19842), .ZN(
        n19848) );
  INV_X1 U22736 ( .A(n19844), .ZN(n19846) );
  OAI21_X1 U22737 ( .B1(P1_REIP_REG_9__SCAN_IN), .B2(n19846), .A(n19845), .ZN(
        n19847) );
  NAND4_X1 U22738 ( .A1(n19850), .A2(n19849), .A3(n19848), .A4(n19847), .ZN(
        P1_U2831) );
  NAND2_X1 U22739 ( .A1(P1_REIP_REG_6__SCAN_IN), .A2(P1_REIP_REG_5__SCAN_IN), 
        .ZN(n19851) );
  NAND2_X1 U22740 ( .A1(n19876), .A2(n19922), .ZN(n19878) );
  OAI21_X1 U22741 ( .B1(n19851), .B2(n19878), .A(n19930), .ZN(n19870) );
  NOR3_X1 U22742 ( .A1(P1_REIP_REG_7__SCAN_IN), .A2(n19875), .A3(n19852), .ZN(
        n19853) );
  AOI211_X1 U22743 ( .C1(n19935), .C2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .A(
        n19891), .B(n19853), .ZN(n19860) );
  INV_X1 U22744 ( .A(n19854), .ZN(n19858) );
  OAI22_X1 U22745 ( .A1(n19856), .A2(n19931), .B1(n19867), .B2(n19855), .ZN(
        n19857) );
  AOI21_X1 U22746 ( .B1(n19934), .B2(n19858), .A(n19857), .ZN(n19859) );
  OAI211_X1 U22747 ( .C1(n19862), .C2(n19861), .A(n19860), .B(n19859), .ZN(
        n19863) );
  INV_X1 U22748 ( .A(n19863), .ZN(n19864) );
  OAI21_X1 U22749 ( .B1(n20629), .B2(n19870), .A(n19864), .ZN(P1_U2833) );
  INV_X1 U22750 ( .A(P1_REIP_REG_6__SCAN_IN), .ZN(n20626) );
  NAND2_X1 U22751 ( .A1(n19939), .A2(n19905), .ZN(n19866) );
  NAND4_X1 U22752 ( .A1(n19920), .A2(n19876), .A3(P1_REIP_REG_5__SCAN_IN), 
        .A4(n20626), .ZN(n19865) );
  OAI211_X1 U22753 ( .C1(n19944), .C2(n19867), .A(n19866), .B(n19865), .ZN(
        n19868) );
  AOI211_X1 U22754 ( .C1(n19935), .C2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .A(
        n19868), .B(n19891), .ZN(n19869) );
  OAI21_X1 U22755 ( .B1(n19870), .B2(n20626), .A(n19869), .ZN(n19871) );
  AOI21_X1 U22756 ( .B1(n19942), .B2(n19872), .A(n19871), .ZN(n19873) );
  OAI21_X1 U22757 ( .B1(n19874), .B2(n19897), .A(n19873), .ZN(P1_U2834) );
  NOR2_X1 U22758 ( .A1(n19875), .A2(P1_REIP_REG_5__SCAN_IN), .ZN(n19877) );
  AOI22_X1 U22759 ( .A1(n19929), .A2(P1_EBX_REG_5__SCAN_IN), .B1(n19877), .B2(
        n19876), .ZN(n19888) );
  INV_X1 U22760 ( .A(P1_REIP_REG_5__SCAN_IN), .ZN(n20624) );
  NAND2_X1 U22761 ( .A1(n19930), .A2(n19878), .ZN(n19898) );
  OAI21_X1 U22762 ( .B1(n20624), .B2(n19898), .A(n19879), .ZN(n19880) );
  INV_X1 U22763 ( .A(n19880), .ZN(n19881) );
  OAI21_X1 U22764 ( .B1(n19882), .B2(n19931), .A(n19881), .ZN(n19883) );
  AOI21_X1 U22765 ( .B1(n19935), .B2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .A(
        n19883), .ZN(n19884) );
  OAI21_X1 U22766 ( .B1(n19885), .B2(n19938), .A(n19884), .ZN(n19886) );
  INV_X1 U22767 ( .A(n19886), .ZN(n19887) );
  OAI211_X1 U22768 ( .C1(n19889), .C2(n19897), .A(n19888), .B(n19887), .ZN(
        P1_U2835) );
  NOR4_X1 U22769 ( .A1(P1_REIP_REG_4__SCAN_IN), .A2(n20620), .A3(n20824), .A4(
        n19907), .ZN(n19890) );
  AOI211_X1 U22770 ( .C1(n19935), .C2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n19891), .B(n19890), .ZN(n19903) );
  INV_X1 U22771 ( .A(n19892), .ZN(n19901) );
  INV_X1 U22772 ( .A(n19938), .ZN(n19912) );
  INV_X1 U22773 ( .A(n19893), .ZN(n19894) );
  AOI22_X1 U22774 ( .A1(n19894), .A2(n19905), .B1(P1_EBX_REG_4__SCAN_IN), .B2(
        n19929), .ZN(n19895) );
  OAI21_X1 U22775 ( .B1(n19897), .B2(n19896), .A(n19895), .ZN(n19900) );
  NOR2_X1 U22776 ( .A1(n19898), .A2(n20621), .ZN(n19899) );
  AOI211_X1 U22777 ( .C1(n19901), .C2(n19912), .A(n19900), .B(n19899), .ZN(
        n19902) );
  OAI211_X1 U22778 ( .C1(n19904), .C2(n19932), .A(n19903), .B(n19902), .ZN(
        P1_U2836) );
  AOI22_X1 U22779 ( .A1(n19906), .A2(n19905), .B1(n19929), .B2(
        P1_EBX_REG_3__SCAN_IN), .ZN(n19919) );
  NOR2_X1 U22780 ( .A1(n19907), .A2(P1_REIP_REG_3__SCAN_IN), .ZN(n19910) );
  OAI22_X1 U22781 ( .A1(n19923), .A2(n19908), .B1(n20325), .B2(n19932), .ZN(
        n19909) );
  AOI21_X1 U22782 ( .B1(n19910), .B2(P1_REIP_REG_2__SCAN_IN), .A(n19909), .ZN(
        n19918) );
  AOI22_X1 U22783 ( .A1(n19913), .A2(n19912), .B1(n19934), .B2(n19911), .ZN(
        n19917) );
  OAI21_X1 U22784 ( .B1(n19915), .B2(n19914), .A(P1_REIP_REG_3__SCAN_IN), .ZN(
        n19916) );
  NAND4_X1 U22785 ( .A1(n19919), .A2(n19918), .A3(n19917), .A4(n19916), .ZN(
        P1_U2837) );
  AOI22_X1 U22786 ( .A1(n19929), .A2(P1_EBX_REG_1__SCAN_IN), .B1(n19920), .B2(
        n20707), .ZN(n19928) );
  INV_X1 U22787 ( .A(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n19926) );
  INV_X1 U22788 ( .A(n20063), .ZN(n19921) );
  OAI22_X1 U22789 ( .A1(n19922), .A2(n20707), .B1(n19921), .B2(n19931), .ZN(
        n19925) );
  OAI22_X1 U22790 ( .A1(n19923), .A2(n19926), .B1(n20438), .B2(n19932), .ZN(
        n19924) );
  AOI211_X1 U22791 ( .C1(n19934), .C2(n19926), .A(n19925), .B(n19924), .ZN(
        n19927) );
  OAI211_X1 U22792 ( .C1(n19938), .C2(n20036), .A(n19928), .B(n19927), .ZN(
        P1_U2839) );
  AOI22_X1 U22793 ( .A1(n19930), .A2(P1_REIP_REG_0__SCAN_IN), .B1(
        P1_EBX_REG_0__SCAN_IN), .B2(n19929), .ZN(n19937) );
  OAI22_X1 U22794 ( .A1(n20181), .A2(n19932), .B1(n19931), .B2(n20082), .ZN(
        n19933) );
  AOI221_X1 U22795 ( .B1(n19935), .B2(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .C1(
        n19934), .C2(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .A(n19933), .ZN(n19936) );
  OAI211_X1 U22796 ( .C1(n19938), .C2(n20045), .A(n19937), .B(n19936), .ZN(
        P1_U2840) );
  AOI22_X1 U22797 ( .A1(n19942), .A2(n19941), .B1(n19940), .B2(n19939), .ZN(
        n19943) );
  OAI21_X1 U22798 ( .B1(n19945), .B2(n19944), .A(n19943), .ZN(P1_U2866) );
  INV_X1 U22799 ( .A(P1_EAX_REG_30__SCAN_IN), .ZN(n19949) );
  NAND2_X1 U22800 ( .A1(n19947), .A2(n19946), .ZN(n19973) );
  AOI22_X1 U22801 ( .A1(P1_UWORD_REG_14__SCAN_IN), .A2(n20729), .B1(n19970), 
        .B2(P1_DATAO_REG_30__SCAN_IN), .ZN(n19948) );
  OAI21_X1 U22802 ( .B1(n19949), .B2(n19973), .A(n19948), .ZN(P1_U2906) );
  INV_X1 U22803 ( .A(P1_EAX_REG_29__SCAN_IN), .ZN(n19951) );
  AOI22_X1 U22804 ( .A1(P1_UWORD_REG_13__SCAN_IN), .A2(n20729), .B1(n19970), 
        .B2(P1_DATAO_REG_29__SCAN_IN), .ZN(n19950) );
  OAI21_X1 U22805 ( .B1(n19951), .B2(n19973), .A(n19950), .ZN(P1_U2907) );
  AOI22_X1 U22806 ( .A1(P1_UWORD_REG_12__SCAN_IN), .A2(n20729), .B1(n19970), 
        .B2(P1_DATAO_REG_28__SCAN_IN), .ZN(n19952) );
  OAI21_X1 U22807 ( .B1(n11007), .B2(n19973), .A(n19952), .ZN(P1_U2908) );
  AOI22_X1 U22808 ( .A1(P1_UWORD_REG_11__SCAN_IN), .A2(n20729), .B1(n19970), 
        .B2(P1_DATAO_REG_27__SCAN_IN), .ZN(n19953) );
  OAI21_X1 U22809 ( .B1(n14377), .B2(n19973), .A(n19953), .ZN(P1_U2909) );
  AOI22_X1 U22810 ( .A1(P1_UWORD_REG_10__SCAN_IN), .A2(n20729), .B1(n19970), 
        .B2(P1_DATAO_REG_26__SCAN_IN), .ZN(n19954) );
  OAI21_X1 U22811 ( .B1(n14382), .B2(n19973), .A(n19954), .ZN(P1_U2910) );
  AOI22_X1 U22812 ( .A1(P1_UWORD_REG_9__SCAN_IN), .A2(n20729), .B1(n19970), 
        .B2(P1_DATAO_REG_25__SCAN_IN), .ZN(n19955) );
  OAI21_X1 U22813 ( .B1(n14387), .B2(n19973), .A(n19955), .ZN(P1_U2911) );
  AOI22_X1 U22814 ( .A1(P1_UWORD_REG_8__SCAN_IN), .A2(n20729), .B1(n19970), 
        .B2(P1_DATAO_REG_24__SCAN_IN), .ZN(n19956) );
  OAI21_X1 U22815 ( .B1(n19957), .B2(n19973), .A(n19956), .ZN(P1_U2912) );
  AOI22_X1 U22816 ( .A1(P1_UWORD_REG_7__SCAN_IN), .A2(n20729), .B1(n19970), 
        .B2(P1_DATAO_REG_23__SCAN_IN), .ZN(n19958) );
  OAI21_X1 U22817 ( .B1(n14397), .B2(n19973), .A(n19958), .ZN(P1_U2913) );
  AOI22_X1 U22818 ( .A1(P1_UWORD_REG_6__SCAN_IN), .A2(n20729), .B1(n19970), 
        .B2(P1_DATAO_REG_22__SCAN_IN), .ZN(n19959) );
  OAI21_X1 U22819 ( .B1(n19960), .B2(n19973), .A(n19959), .ZN(P1_U2914) );
  INV_X1 U22820 ( .A(P1_EAX_REG_21__SCAN_IN), .ZN(n19962) );
  AOI22_X1 U22821 ( .A1(P1_UWORD_REG_5__SCAN_IN), .A2(n20729), .B1(n19970), 
        .B2(P1_DATAO_REG_21__SCAN_IN), .ZN(n19961) );
  OAI21_X1 U22822 ( .B1(n19962), .B2(n19973), .A(n19961), .ZN(P1_U2915) );
  AOI22_X1 U22823 ( .A1(P1_UWORD_REG_4__SCAN_IN), .A2(n20729), .B1(n19970), 
        .B2(P1_DATAO_REG_20__SCAN_IN), .ZN(n19963) );
  OAI21_X1 U22824 ( .B1(n19964), .B2(n19973), .A(n19963), .ZN(P1_U2916) );
  INV_X1 U22825 ( .A(P1_UWORD_REG_3__SCAN_IN), .ZN(n20903) );
  INV_X1 U22826 ( .A(n19973), .ZN(n19965) );
  AOI22_X1 U22827 ( .A1(P1_EAX_REG_19__SCAN_IN), .A2(n19965), .B1(n19970), 
        .B2(P1_DATAO_REG_19__SCAN_IN), .ZN(n19966) );
  OAI21_X1 U22828 ( .B1(n20903), .B2(n19967), .A(n19966), .ZN(P1_U2917) );
  INV_X1 U22829 ( .A(P1_EAX_REG_18__SCAN_IN), .ZN(n19969) );
  AOI22_X1 U22830 ( .A1(P1_UWORD_REG_2__SCAN_IN), .A2(n20729), .B1(n19970), 
        .B2(P1_DATAO_REG_18__SCAN_IN), .ZN(n19968) );
  OAI21_X1 U22831 ( .B1(n19969), .B2(n19973), .A(n19968), .ZN(P1_U2918) );
  AOI22_X1 U22832 ( .A1(P1_UWORD_REG_1__SCAN_IN), .A2(n20729), .B1(n19970), 
        .B2(P1_DATAO_REG_17__SCAN_IN), .ZN(n19971) );
  OAI21_X1 U22833 ( .B1(n14426), .B2(n19973), .A(n19971), .ZN(P1_U2919) );
  AOI22_X1 U22834 ( .A1(P1_UWORD_REG_0__SCAN_IN), .A2(n20729), .B1(n19970), 
        .B2(P1_DATAO_REG_16__SCAN_IN), .ZN(n19972) );
  OAI21_X1 U22835 ( .B1(n19974), .B2(n19973), .A(n19972), .ZN(P1_U2920) );
  AOI22_X1 U22836 ( .A1(P1_LWORD_REG_15__SCAN_IN), .A2(n20729), .B1(n19970), 
        .B2(P1_DATAO_REG_15__SCAN_IN), .ZN(n19975) );
  OAI21_X1 U22837 ( .B1(n13278), .B2(n19996), .A(n19975), .ZN(P1_U2921) );
  AOI22_X1 U22838 ( .A1(P1_LWORD_REG_14__SCAN_IN), .A2(n20729), .B1(n19970), 
        .B2(P1_DATAO_REG_14__SCAN_IN), .ZN(n19976) );
  OAI21_X1 U22839 ( .B1(n14113), .B2(n19996), .A(n19976), .ZN(P1_U2922) );
  AOI22_X1 U22840 ( .A1(P1_LWORD_REG_13__SCAN_IN), .A2(n20729), .B1(n19970), 
        .B2(P1_DATAO_REG_13__SCAN_IN), .ZN(n19977) );
  OAI21_X1 U22841 ( .B1(n14141), .B2(n19996), .A(n19977), .ZN(P1_U2923) );
  INV_X1 U22842 ( .A(P1_EAX_REG_12__SCAN_IN), .ZN(n19979) );
  AOI22_X1 U22843 ( .A1(P1_LWORD_REG_12__SCAN_IN), .A2(n20729), .B1(n19970), 
        .B2(P1_DATAO_REG_12__SCAN_IN), .ZN(n19978) );
  OAI21_X1 U22844 ( .B1(n19979), .B2(n19996), .A(n19978), .ZN(P1_U2924) );
  AOI22_X1 U22845 ( .A1(P1_LWORD_REG_11__SCAN_IN), .A2(n20729), .B1(n19970), 
        .B2(P1_DATAO_REG_11__SCAN_IN), .ZN(n19980) );
  OAI21_X1 U22846 ( .B1(n14087), .B2(n19996), .A(n19980), .ZN(P1_U2925) );
  INV_X1 U22847 ( .A(P1_EAX_REG_10__SCAN_IN), .ZN(n19982) );
  AOI22_X1 U22848 ( .A1(P1_LWORD_REG_10__SCAN_IN), .A2(n20729), .B1(n19970), 
        .B2(P1_DATAO_REG_10__SCAN_IN), .ZN(n19981) );
  OAI21_X1 U22849 ( .B1(n19982), .B2(n19996), .A(n19981), .ZN(P1_U2926) );
  INV_X1 U22850 ( .A(P1_EAX_REG_9__SCAN_IN), .ZN(n19984) );
  AOI22_X1 U22851 ( .A1(P1_LWORD_REG_9__SCAN_IN), .A2(n20729), .B1(n19970), 
        .B2(P1_DATAO_REG_9__SCAN_IN), .ZN(n19983) );
  OAI21_X1 U22852 ( .B1(n19984), .B2(n19996), .A(n19983), .ZN(P1_U2927) );
  AOI22_X1 U22853 ( .A1(P1_LWORD_REG_8__SCAN_IN), .A2(n20729), .B1(n19970), 
        .B2(P1_DATAO_REG_8__SCAN_IN), .ZN(n19985) );
  OAI21_X1 U22854 ( .B1(n13726), .B2(n19996), .A(n19985), .ZN(P1_U2928) );
  AOI22_X1 U22855 ( .A1(P1_LWORD_REG_7__SCAN_IN), .A2(n20729), .B1(n19970), 
        .B2(P1_DATAO_REG_7__SCAN_IN), .ZN(n19986) );
  OAI21_X1 U22856 ( .B1(n10480), .B2(n19996), .A(n19986), .ZN(P1_U2929) );
  AOI22_X1 U22857 ( .A1(P1_LWORD_REG_6__SCAN_IN), .A2(n20729), .B1(n19970), 
        .B2(P1_DATAO_REG_6__SCAN_IN), .ZN(n19987) );
  OAI21_X1 U22858 ( .B1(n13751), .B2(n19996), .A(n19987), .ZN(P1_U2930) );
  AOI22_X1 U22859 ( .A1(P1_DATAO_REG_5__SCAN_IN), .A2(n19970), .B1(
        P1_LWORD_REG_5__SCAN_IN), .B2(n20729), .ZN(n19988) );
  OAI21_X1 U22860 ( .B1(n19989), .B2(n19996), .A(n19988), .ZN(P1_U2931) );
  AOI22_X1 U22861 ( .A1(P1_LWORD_REG_4__SCAN_IN), .A2(n20729), .B1(n19970), 
        .B2(P1_DATAO_REG_4__SCAN_IN), .ZN(n19990) );
  OAI21_X1 U22862 ( .B1(n19991), .B2(n19996), .A(n19990), .ZN(P1_U2932) );
  AOI22_X1 U22863 ( .A1(P1_LWORD_REG_3__SCAN_IN), .A2(n20729), .B1(n19970), 
        .B2(P1_DATAO_REG_3__SCAN_IN), .ZN(n19992) );
  OAI21_X1 U22864 ( .B1(n10407), .B2(n19996), .A(n19992), .ZN(P1_U2933) );
  AOI22_X1 U22865 ( .A1(P1_LWORD_REG_2__SCAN_IN), .A2(n20729), .B1(n19970), 
        .B2(P1_DATAO_REG_2__SCAN_IN), .ZN(n19993) );
  OAI21_X1 U22866 ( .B1(n10355), .B2(n19996), .A(n19993), .ZN(P1_U2934) );
  AOI22_X1 U22867 ( .A1(P1_LWORD_REG_1__SCAN_IN), .A2(n20729), .B1(n19970), 
        .B2(P1_DATAO_REG_1__SCAN_IN), .ZN(n19994) );
  OAI21_X1 U22868 ( .B1(n10374), .B2(n19996), .A(n19994), .ZN(P1_U2935) );
  AOI22_X1 U22869 ( .A1(P1_LWORD_REG_0__SCAN_IN), .A2(n20729), .B1(n19970), 
        .B2(P1_DATAO_REG_0__SCAN_IN), .ZN(n19995) );
  OAI21_X1 U22870 ( .B1(n10366), .B2(n19996), .A(n19995), .ZN(P1_U2936) );
  INV_X1 U22871 ( .A(P1_UWORD_REG_8__SCAN_IN), .ZN(n20871) );
  NAND2_X1 U22872 ( .A1(n9752), .A2(n19997), .ZN(n20013) );
  INV_X1 U22873 ( .A(n20013), .ZN(n19998) );
  AOI21_X1 U22874 ( .B1(n9753), .B2(P1_EAX_REG_24__SCAN_IN), .A(n19998), .ZN(
        n19999) );
  OAI21_X1 U22875 ( .B1(n20000), .B2(n20871), .A(n19999), .ZN(P1_U2945) );
  AOI22_X1 U22876 ( .A1(n9753), .A2(P1_EAX_REG_25__SCAN_IN), .B1(n20025), .B2(
        P1_UWORD_REG_9__SCAN_IN), .ZN(n20002) );
  NAND2_X1 U22877 ( .A1(n9752), .A2(n20001), .ZN(n20015) );
  NAND2_X1 U22878 ( .A1(n20002), .A2(n20015), .ZN(P1_U2946) );
  AOI22_X1 U22879 ( .A1(n9753), .A2(P1_EAX_REG_26__SCAN_IN), .B1(n20025), .B2(
        P1_UWORD_REG_10__SCAN_IN), .ZN(n20004) );
  NAND2_X1 U22880 ( .A1(n9752), .A2(n20003), .ZN(n20017) );
  NAND2_X1 U22881 ( .A1(n20004), .A2(n20017), .ZN(P1_U2947) );
  AOI22_X1 U22882 ( .A1(n9753), .A2(P1_EAX_REG_27__SCAN_IN), .B1(n20025), .B2(
        P1_UWORD_REG_11__SCAN_IN), .ZN(n20006) );
  NAND2_X1 U22883 ( .A1(n9752), .A2(n20005), .ZN(n20019) );
  NAND2_X1 U22884 ( .A1(n20006), .A2(n20019), .ZN(P1_U2948) );
  AOI22_X1 U22885 ( .A1(n9753), .A2(P1_EAX_REG_28__SCAN_IN), .B1(n20025), .B2(
        P1_UWORD_REG_12__SCAN_IN), .ZN(n20008) );
  NAND2_X1 U22886 ( .A1(n9752), .A2(n20007), .ZN(n20021) );
  NAND2_X1 U22887 ( .A1(n20008), .A2(n20021), .ZN(P1_U2949) );
  AOI22_X1 U22888 ( .A1(n9753), .A2(P1_EAX_REG_29__SCAN_IN), .B1(n20025), .B2(
        P1_UWORD_REG_13__SCAN_IN), .ZN(n20010) );
  NAND2_X1 U22889 ( .A1(n9752), .A2(n20009), .ZN(n20023) );
  NAND2_X1 U22890 ( .A1(n20010), .A2(n20023), .ZN(P1_U2950) );
  AOI22_X1 U22891 ( .A1(n9753), .A2(P1_EAX_REG_30__SCAN_IN), .B1(n20025), .B2(
        P1_UWORD_REG_14__SCAN_IN), .ZN(n20012) );
  NAND2_X1 U22892 ( .A1(n9752), .A2(n20011), .ZN(n20027) );
  NAND2_X1 U22893 ( .A1(n20012), .A2(n20027), .ZN(P1_U2951) );
  AOI22_X1 U22894 ( .A1(n9753), .A2(P1_EAX_REG_8__SCAN_IN), .B1(n20025), .B2(
        P1_LWORD_REG_8__SCAN_IN), .ZN(n20014) );
  NAND2_X1 U22895 ( .A1(n20014), .A2(n20013), .ZN(P1_U2960) );
  AOI22_X1 U22896 ( .A1(n9753), .A2(P1_EAX_REG_9__SCAN_IN), .B1(n20025), .B2(
        P1_LWORD_REG_9__SCAN_IN), .ZN(n20016) );
  NAND2_X1 U22897 ( .A1(n20016), .A2(n20015), .ZN(P1_U2961) );
  AOI22_X1 U22898 ( .A1(n9753), .A2(P1_EAX_REG_10__SCAN_IN), .B1(n20025), .B2(
        P1_LWORD_REG_10__SCAN_IN), .ZN(n20018) );
  NAND2_X1 U22899 ( .A1(n20018), .A2(n20017), .ZN(P1_U2962) );
  AOI22_X1 U22900 ( .A1(n9753), .A2(P1_EAX_REG_11__SCAN_IN), .B1(n20025), .B2(
        P1_LWORD_REG_11__SCAN_IN), .ZN(n20020) );
  NAND2_X1 U22901 ( .A1(n20020), .A2(n20019), .ZN(P1_U2963) );
  AOI22_X1 U22902 ( .A1(n9753), .A2(P1_EAX_REG_12__SCAN_IN), .B1(n20025), .B2(
        P1_LWORD_REG_12__SCAN_IN), .ZN(n20022) );
  NAND2_X1 U22903 ( .A1(n20022), .A2(n20021), .ZN(P1_U2964) );
  AOI22_X1 U22904 ( .A1(n9753), .A2(P1_EAX_REG_13__SCAN_IN), .B1(n20025), .B2(
        P1_LWORD_REG_13__SCAN_IN), .ZN(n20024) );
  NAND2_X1 U22905 ( .A1(n20024), .A2(n20023), .ZN(P1_U2965) );
  AOI22_X1 U22906 ( .A1(n9753), .A2(P1_EAX_REG_14__SCAN_IN), .B1(n20025), .B2(
        P1_LWORD_REG_14__SCAN_IN), .ZN(n20028) );
  NAND2_X1 U22907 ( .A1(n20028), .A2(n20027), .ZN(P1_U2966) );
  NOR2_X1 U22908 ( .A1(n20050), .A2(n20707), .ZN(n20062) );
  OAI21_X1 U22909 ( .B1(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n20030), .A(
        n20029), .ZN(n20071) );
  OAI22_X1 U22910 ( .A1(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n20032), .B1(
        n20031), .B2(n20071), .ZN(n20033) );
  AOI211_X1 U22911 ( .C1(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .C2(n20034), .A(
        n20062), .B(n20033), .ZN(n20035) );
  OAI21_X1 U22912 ( .B1(n20084), .B2(n20036), .A(n20035), .ZN(P1_U2998) );
  AOI21_X1 U22913 ( .B1(n20038), .B2(n20072), .A(n20037), .ZN(n20077) );
  NAND2_X1 U22914 ( .A1(n20040), .A2(n20039), .ZN(n20041) );
  AOI22_X1 U22915 ( .A1(n20042), .A2(n20077), .B1(
        P1_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n20041), .ZN(n20044) );
  NAND2_X1 U22916 ( .A1(n20043), .A2(P1_REIP_REG_0__SCAN_IN), .ZN(n20079) );
  OAI211_X1 U22917 ( .C1(n20045), .C2(n20084), .A(n20044), .B(n20079), .ZN(
        P1_U2999) );
  AOI21_X1 U22918 ( .B1(n10874), .B2(n20047), .A(n20046), .ZN(n20057) );
  NOR2_X1 U22919 ( .A1(n20072), .A2(n10874), .ZN(n20049) );
  AOI21_X1 U22920 ( .B1(n20049), .B2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A(
        n20048), .ZN(n20051) );
  OAI22_X1 U22921 ( .A1(n20051), .A2(n20066), .B1(n20824), .B2(n20050), .ZN(
        n20054) );
  NOR2_X1 U22922 ( .A1(n20052), .A2(n20070), .ZN(n20053) );
  AOI211_X1 U22923 ( .C1(n20055), .C2(n20064), .A(n20054), .B(n20053), .ZN(
        n20056) );
  OAI221_X1 U22924 ( .B1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n20058), .C1(
        n11122), .C2(n20057), .A(n20056), .ZN(P1_U3029) );
  NOR3_X1 U22925 ( .A1(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n20060), .A3(
        n20059), .ZN(n20061) );
  AOI211_X1 U22926 ( .C1(n20064), .C2(n20063), .A(n20062), .B(n20061), .ZN(
        n20069) );
  AOI21_X1 U22927 ( .B1(n20066), .B2(n20065), .A(
        P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n20075) );
  OAI21_X1 U22928 ( .B1(n20067), .B2(n20075), .A(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n20068) );
  OAI211_X1 U22929 ( .C1(n20071), .C2(n20070), .A(n20069), .B(n20068), .ZN(
        P1_U3030) );
  AOI21_X1 U22930 ( .B1(n20074), .B2(n20073), .A(n20072), .ZN(n20076) );
  AOI211_X1 U22931 ( .C1(n20078), .C2(n20077), .A(n20076), .B(n20075), .ZN(
        n20080) );
  OAI211_X1 U22932 ( .C1(n20082), .C2(n20081), .A(n20080), .B(n20079), .ZN(
        P1_U3031) );
  AND2_X1 U22933 ( .A1(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n20706), .ZN(
        P1_U3032) );
  NOR2_X2 U22934 ( .A1(n20084), .A2(n20083), .ZN(n20120) );
  NOR2_X2 U22935 ( .A1(n20085), .A2(n20084), .ZN(n20119) );
  AOI22_X1 U22936 ( .A1(BUF1_REG_16__SCAN_IN), .A2(n20120), .B1(DATAI_16_), 
        .B2(n20119), .ZN(n20552) );
  INV_X1 U22937 ( .A(n13433), .ZN(n20693) );
  AOI22_X1 U22938 ( .A1(BUF1_REG_24__SCAN_IN), .A2(n20120), .B1(DATAI_24_), 
        .B2(n20119), .ZN(n20504) );
  INV_X1 U22939 ( .A(n20504), .ZN(n20549) );
  NAND2_X1 U22940 ( .A1(n20690), .A2(n20326), .ZN(n20185) );
  OR2_X1 U22941 ( .A1(n20433), .A2(n20185), .ZN(n20087) );
  INV_X1 U22942 ( .A(n20087), .ZN(n20122) );
  NOR2_X2 U22943 ( .A1(n20086), .A2(n20118), .ZN(n20543) );
  AOI22_X1 U22944 ( .A1(n20121), .A2(n20549), .B1(n20122), .B2(n20543), .ZN(
        n20095) );
  OR2_X1 U22945 ( .A1(n20684), .A2(n20324), .ZN(n20182) );
  INV_X1 U22946 ( .A(n20438), .ZN(n20695) );
  NOR2_X1 U22947 ( .A1(n20182), .A2(n20695), .ZN(n20090) );
  OAI221_X1 U22948 ( .B1(n20891), .B2(n20934), .C1(n20891), .C2(n20595), .A(
        n20700), .ZN(n20093) );
  NAND2_X1 U22949 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n20091), .ZN(n20492) );
  AND2_X1 U22950 ( .A1(n20218), .A2(n20492), .ZN(n20377) );
  NAND2_X1 U22951 ( .A1(n20327), .A2(n20378), .ZN(n20215) );
  AOI22_X1 U22952 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n20215), .B1(
        P1_STATE2_REG_3__SCAN_IN), .B2(n20087), .ZN(n20088) );
  OAI211_X1 U22953 ( .C1(n20090), .C2(n20093), .A(n20377), .B(n20088), .ZN(
        n20125) );
  NOR2_X2 U22954 ( .A1(n20089), .A2(n20131), .ZN(n20544) );
  INV_X1 U22955 ( .A(n20090), .ZN(n20092) );
  OR2_X1 U22956 ( .A1(n20599), .A2(n20091), .ZN(n20382) );
  OAI22_X1 U22957 ( .A1(n20093), .A2(n20092), .B1(n20382), .B2(n20215), .ZN(
        n20124) );
  AOI22_X1 U22958 ( .A1(P1_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n20125), .B1(
        n20544), .B2(n20124), .ZN(n20094) );
  OAI211_X1 U22959 ( .C1(n20552), .C2(n20934), .A(n20095), .B(n20094), .ZN(
        P1_U3033) );
  AOI22_X1 U22960 ( .A1(DATAI_17_), .A2(n20119), .B1(BUF1_REG_17__SCAN_IN), 
        .B2(n20120), .ZN(n20557) );
  AOI22_X1 U22961 ( .A1(BUF1_REG_25__SCAN_IN), .A2(n20120), .B1(DATAI_25_), 
        .B2(n20119), .ZN(n20508) );
  INV_X1 U22962 ( .A(n20508), .ZN(n20554) );
  AOI22_X1 U22963 ( .A1(n9663), .A2(n20122), .B1(n20121), .B2(n20554), .ZN(
        n20099) );
  NOR2_X2 U22964 ( .A1(n20097), .A2(n20131), .ZN(n20553) );
  AOI22_X1 U22965 ( .A1(P1_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n20125), .B1(
        n20553), .B2(n20124), .ZN(n20098) );
  OAI211_X1 U22966 ( .C1(n20557), .C2(n20934), .A(n20099), .B(n20098), .ZN(
        P1_U3034) );
  AOI22_X1 U22967 ( .A1(DATAI_18_), .A2(n20119), .B1(BUF1_REG_18__SCAN_IN), 
        .B2(n20120), .ZN(n20563) );
  AOI22_X1 U22968 ( .A1(BUF1_REG_26__SCAN_IN), .A2(n20120), .B1(DATAI_26_), 
        .B2(n20119), .ZN(n20512) );
  INV_X1 U22969 ( .A(n20512), .ZN(n20560) );
  NOR2_X2 U22970 ( .A1(n13172), .A2(n20118), .ZN(n20558) );
  AOI22_X1 U22971 ( .A1(n20121), .A2(n20560), .B1(n20122), .B2(n20558), .ZN(
        n20102) );
  NOR2_X2 U22972 ( .A1(n20100), .A2(n20131), .ZN(n20559) );
  AOI22_X1 U22973 ( .A1(P1_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n20125), .B1(
        n20559), .B2(n20124), .ZN(n20101) );
  OAI211_X1 U22974 ( .C1(n20563), .C2(n20934), .A(n20102), .B(n20101), .ZN(
        P1_U3035) );
  AOI22_X1 U22975 ( .A1(BUF1_REG_19__SCAN_IN), .A2(n20120), .B1(DATAI_19_), 
        .B2(n20119), .ZN(n20569) );
  AOI22_X1 U22976 ( .A1(BUF1_REG_27__SCAN_IN), .A2(n20120), .B1(DATAI_27_), 
        .B2(n20119), .ZN(n20516) );
  INV_X1 U22977 ( .A(n20516), .ZN(n20566) );
  NOR2_X2 U22978 ( .A1(n20103), .A2(n20118), .ZN(n20564) );
  AOI22_X1 U22979 ( .A1(n20121), .A2(n20566), .B1(n20122), .B2(n20564), .ZN(
        n20106) );
  NOR2_X2 U22980 ( .A1(n20104), .A2(n20131), .ZN(n20565) );
  AOI22_X1 U22981 ( .A1(P1_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n20125), .B1(
        n20565), .B2(n20124), .ZN(n20105) );
  OAI211_X1 U22982 ( .C1(n20569), .C2(n20934), .A(n20106), .B(n20105), .ZN(
        P1_U3036) );
  AOI22_X1 U22983 ( .A1(BUF1_REG_20__SCAN_IN), .A2(n20120), .B1(DATAI_20_), 
        .B2(n20119), .ZN(n20575) );
  AOI22_X1 U22984 ( .A1(BUF1_REG_28__SCAN_IN), .A2(n20120), .B1(DATAI_28_), 
        .B2(n20119), .ZN(n20520) );
  INV_X1 U22985 ( .A(n20520), .ZN(n20572) );
  AOI22_X1 U22986 ( .A1(n20121), .A2(n20572), .B1(n20122), .B2(n20570), .ZN(
        n20110) );
  NOR2_X2 U22987 ( .A1(n20108), .A2(n20131), .ZN(n20571) );
  AOI22_X1 U22988 ( .A1(P1_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n20125), .B1(
        n20571), .B2(n20124), .ZN(n20109) );
  OAI211_X1 U22989 ( .C1(n20575), .C2(n20934), .A(n20110), .B(n20109), .ZN(
        P1_U3037) );
  AOI22_X1 U22990 ( .A1(BUF1_REG_21__SCAN_IN), .A2(n20120), .B1(DATAI_21_), 
        .B2(n20119), .ZN(n20581) );
  AOI22_X1 U22991 ( .A1(BUF1_REG_29__SCAN_IN), .A2(n20120), .B1(DATAI_29_), 
        .B2(n20119), .ZN(n20524) );
  INV_X1 U22992 ( .A(n20524), .ZN(n20578) );
  NOR2_X2 U22993 ( .A1(n10248), .A2(n20118), .ZN(n20576) );
  AOI22_X1 U22994 ( .A1(n20121), .A2(n20578), .B1(n20122), .B2(n20576), .ZN(
        n20113) );
  NOR2_X2 U22995 ( .A1(n20111), .A2(n20131), .ZN(n20577) );
  AOI22_X1 U22996 ( .A1(P1_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n20125), .B1(
        n20577), .B2(n20124), .ZN(n20112) );
  OAI211_X1 U22997 ( .C1(n20581), .C2(n20934), .A(n20113), .B(n20112), .ZN(
        P1_U3038) );
  AOI22_X1 U22998 ( .A1(BUF1_REG_22__SCAN_IN), .A2(n20120), .B1(DATAI_22_), 
        .B2(n20119), .ZN(n20585) );
  AOI22_X1 U22999 ( .A1(BUF1_REG_30__SCAN_IN), .A2(n20120), .B1(DATAI_30_), 
        .B2(n20119), .ZN(n20935) );
  INV_X1 U23000 ( .A(n20935), .ZN(n20582) );
  NOR2_X2 U23001 ( .A1(n10274), .A2(n20118), .ZN(n20926) );
  AOI22_X1 U23002 ( .A1(n20121), .A2(n20582), .B1(n20122), .B2(n20926), .ZN(
        n20116) );
  NOR2_X2 U23003 ( .A1(n20114), .A2(n20131), .ZN(n20928) );
  AOI22_X1 U23004 ( .A1(P1_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n20125), .B1(
        n20928), .B2(n20124), .ZN(n20115) );
  OAI211_X1 U23005 ( .C1(n20585), .C2(n20934), .A(n20116), .B(n20115), .ZN(
        P1_U3039) );
  AOI22_X1 U23006 ( .A1(BUF1_REG_23__SCAN_IN), .A2(n20120), .B1(DATAI_23_), 
        .B2(n20119), .ZN(n20596) );
  NOR2_X2 U23007 ( .A1(n20118), .A2(n20117), .ZN(n20589) );
  AOI22_X1 U23008 ( .A1(BUF1_REG_31__SCAN_IN), .A2(n20120), .B1(DATAI_31_), 
        .B2(n20119), .ZN(n20534) );
  INV_X1 U23009 ( .A(n20534), .ZN(n20590) );
  AOI22_X1 U23010 ( .A1(n20589), .A2(n20122), .B1(n20121), .B2(n20590), .ZN(
        n20127) );
  NOR2_X2 U23011 ( .A1(n20123), .A2(n20131), .ZN(n20587) );
  AOI22_X1 U23012 ( .A1(P1_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n20125), .B1(
        n20587), .B2(n20124), .ZN(n20126) );
  OAI211_X1 U23013 ( .C1(n20596), .C2(n20934), .A(n20127), .B(n20126), .ZN(
        P1_U3040) );
  INV_X1 U23014 ( .A(n20182), .ZN(n20129) );
  INV_X1 U23015 ( .A(n20128), .ZN(n20465) );
  AOI21_X1 U23016 ( .B1(n20129), .B2(n20465), .A(n20925), .ZN(n20132) );
  INV_X1 U23017 ( .A(n20185), .ZN(n20188) );
  NAND2_X1 U23018 ( .A1(n20188), .A2(n20697), .ZN(n20130) );
  OAI22_X1 U23019 ( .A1(n20132), .A2(n20541), .B1(n20130), .B2(n20599), .ZN(
        n20927) );
  AOI22_X1 U23020 ( .A1(n20544), .A2(n20927), .B1(n20543), .B2(n20925), .ZN(
        n20136) );
  INV_X1 U23021 ( .A(n20130), .ZN(n20134) );
  INV_X1 U23022 ( .A(n20178), .ZN(n20179) );
  NAND2_X1 U23023 ( .A1(P1_STATEBS16_REG_SCAN_IN), .A2(n20693), .ZN(n20469) );
  OAI211_X1 U23024 ( .C1(n20179), .C2(n20469), .A(n20700), .B(n20132), .ZN(
        n20133) );
  OAI211_X1 U23025 ( .C1(n20700), .C2(n20134), .A(n20546), .B(n20133), .ZN(
        n20931) );
  NOR2_X1 U23026 ( .A1(n20149), .A2(n13433), .ZN(n20243) );
  INV_X1 U23027 ( .A(n20552), .ZN(n20501) );
  AOI22_X1 U23028 ( .A1(P1_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n20931), .B1(
        n20930), .B2(n20501), .ZN(n20135) );
  OAI211_X1 U23029 ( .C1(n20504), .C2(n20934), .A(n20136), .B(n20135), .ZN(
        P1_U3041) );
  AOI22_X1 U23030 ( .A1(n9663), .A2(n20925), .B1(n20553), .B2(n20927), .ZN(
        n20138) );
  INV_X1 U23031 ( .A(n20557), .ZN(n20505) );
  AOI22_X1 U23032 ( .A1(P1_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n20931), .B1(
        n20930), .B2(n20505), .ZN(n20137) );
  OAI211_X1 U23033 ( .C1(n20508), .C2(n20934), .A(n20138), .B(n20137), .ZN(
        P1_U3042) );
  AOI22_X1 U23034 ( .A1(n20559), .A2(n20927), .B1(n20558), .B2(n20925), .ZN(
        n20140) );
  INV_X1 U23035 ( .A(n20563), .ZN(n20509) );
  AOI22_X1 U23036 ( .A1(P1_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n20931), .B1(
        n20930), .B2(n20509), .ZN(n20139) );
  OAI211_X1 U23037 ( .C1(n20512), .C2(n20934), .A(n20140), .B(n20139), .ZN(
        P1_U3043) );
  AOI22_X1 U23038 ( .A1(n20565), .A2(n20927), .B1(n20564), .B2(n20925), .ZN(
        n20142) );
  INV_X1 U23039 ( .A(n20569), .ZN(n20513) );
  AOI22_X1 U23040 ( .A1(P1_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n20931), .B1(
        n20930), .B2(n20513), .ZN(n20141) );
  OAI211_X1 U23041 ( .C1(n20516), .C2(n20934), .A(n20142), .B(n20141), .ZN(
        P1_U3044) );
  AOI22_X1 U23042 ( .A1(n20571), .A2(n20927), .B1(n20570), .B2(n20925), .ZN(
        n20144) );
  INV_X1 U23043 ( .A(n20575), .ZN(n20517) );
  AOI22_X1 U23044 ( .A1(P1_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n20931), .B1(
        n20930), .B2(n20517), .ZN(n20143) );
  OAI211_X1 U23045 ( .C1(n20520), .C2(n20934), .A(n20144), .B(n20143), .ZN(
        P1_U3045) );
  AOI22_X1 U23046 ( .A1(n20577), .A2(n20927), .B1(n20576), .B2(n20925), .ZN(
        n20146) );
  INV_X1 U23047 ( .A(n20581), .ZN(n20521) );
  AOI22_X1 U23048 ( .A1(P1_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n20931), .B1(
        n20930), .B2(n20521), .ZN(n20145) );
  OAI211_X1 U23049 ( .C1(n20524), .C2(n20934), .A(n20146), .B(n20145), .ZN(
        P1_U3046) );
  AOI22_X1 U23050 ( .A1(n20589), .A2(n20925), .B1(n20587), .B2(n20927), .ZN(
        n20148) );
  INV_X1 U23051 ( .A(n20596), .ZN(n20529) );
  AOI22_X1 U23052 ( .A1(P1_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n20931), .B1(
        n20930), .B2(n20529), .ZN(n20147) );
  OAI211_X1 U23053 ( .C1(n20534), .C2(n20934), .A(n20148), .B(n20147), .ZN(
        P1_U3048) );
  NOR3_X2 U23054 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20697), .A3(
        n20185), .ZN(n20171) );
  NAND2_X1 U23055 ( .A1(n20149), .A2(n13433), .ZN(n20493) );
  INV_X1 U23056 ( .A(n20493), .ZN(n20150) );
  AOI22_X1 U23057 ( .A1(n20171), .A2(n20543), .B1(n20207), .B2(n20501), .ZN(
        n20158) );
  NOR2_X1 U23058 ( .A1(n20182), .A2(n20438), .ZN(n20154) );
  OAI221_X1 U23059 ( .B1(n20891), .B2(n20176), .C1(n20891), .C2(n20206), .A(
        n20700), .ZN(n20155) );
  INV_X1 U23060 ( .A(n20171), .ZN(n20151) );
  NOR2_X1 U23061 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n20378), .ZN(
        n20153) );
  NOR2_X1 U23062 ( .A1(n20153), .A2(n20599), .ZN(n20265) );
  AOI21_X1 U23063 ( .B1(P1_STATE2_REG_3__SCAN_IN), .B2(n20151), .A(n20265), 
        .ZN(n20152) );
  OAI211_X1 U23064 ( .C1(n20154), .C2(n20155), .A(n20377), .B(n20152), .ZN(
        n20173) );
  INV_X1 U23065 ( .A(n20153), .ZN(n20270) );
  INV_X1 U23066 ( .A(n20154), .ZN(n20156) );
  OAI22_X1 U23067 ( .A1(n20382), .A2(n20270), .B1(n20156), .B2(n20155), .ZN(
        n20172) );
  AOI22_X1 U23068 ( .A1(P1_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n20173), .B1(
        n20544), .B2(n20172), .ZN(n20157) );
  OAI211_X1 U23069 ( .C1(n20504), .C2(n20176), .A(n20158), .B(n20157), .ZN(
        P1_U3049) );
  AOI22_X1 U23070 ( .A1(n9663), .A2(n20171), .B1(n20930), .B2(n20554), .ZN(
        n20160) );
  AOI22_X1 U23071 ( .A1(P1_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n20173), .B1(
        n20553), .B2(n20172), .ZN(n20159) );
  OAI211_X1 U23072 ( .C1(n20557), .C2(n20206), .A(n20160), .B(n20159), .ZN(
        P1_U3050) );
  AOI22_X1 U23073 ( .A1(n20171), .A2(n20558), .B1(n20207), .B2(n20509), .ZN(
        n20162) );
  AOI22_X1 U23074 ( .A1(P1_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n20173), .B1(
        n20559), .B2(n20172), .ZN(n20161) );
  OAI211_X1 U23075 ( .C1(n20512), .C2(n20176), .A(n20162), .B(n20161), .ZN(
        P1_U3051) );
  AOI22_X1 U23076 ( .A1(n20171), .A2(n20564), .B1(n20930), .B2(n20566), .ZN(
        n20164) );
  AOI22_X1 U23077 ( .A1(P1_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n20173), .B1(
        n20565), .B2(n20172), .ZN(n20163) );
  OAI211_X1 U23078 ( .C1(n20569), .C2(n20206), .A(n20164), .B(n20163), .ZN(
        P1_U3052) );
  AOI22_X1 U23079 ( .A1(n20171), .A2(n20570), .B1(n20207), .B2(n20517), .ZN(
        n20166) );
  AOI22_X1 U23080 ( .A1(P1_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n20173), .B1(
        n20571), .B2(n20172), .ZN(n20165) );
  OAI211_X1 U23081 ( .C1(n20520), .C2(n20176), .A(n20166), .B(n20165), .ZN(
        P1_U3053) );
  AOI22_X1 U23082 ( .A1(n20171), .A2(n20576), .B1(n20207), .B2(n20521), .ZN(
        n20168) );
  AOI22_X1 U23083 ( .A1(P1_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n20173), .B1(
        n20577), .B2(n20172), .ZN(n20167) );
  OAI211_X1 U23084 ( .C1(n20524), .C2(n20176), .A(n20168), .B(n20167), .ZN(
        P1_U3054) );
  AOI22_X1 U23085 ( .A1(n20926), .A2(n20171), .B1(n20930), .B2(n20582), .ZN(
        n20170) );
  AOI22_X1 U23086 ( .A1(P1_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n20173), .B1(
        n20928), .B2(n20172), .ZN(n20169) );
  OAI211_X1 U23087 ( .C1(n20585), .C2(n20206), .A(n20170), .B(n20169), .ZN(
        P1_U3055) );
  AOI22_X1 U23088 ( .A1(n20589), .A2(n20171), .B1(n20207), .B2(n20529), .ZN(
        n20175) );
  AOI22_X1 U23089 ( .A1(P1_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n20173), .B1(
        n20587), .B2(n20172), .ZN(n20174) );
  OAI211_X1 U23090 ( .C1(n20534), .C2(n20176), .A(n20175), .B(n20174), .ZN(
        P1_U3056) );
  AND2_X1 U23091 ( .A1(n20536), .A2(n20188), .ZN(n20208) );
  AOI22_X1 U23092 ( .A1(n20543), .A2(n20208), .B1(n20207), .B2(n20549), .ZN(
        n20193) );
  OAI21_X1 U23093 ( .B1(n20179), .B2(n20691), .A(n20700), .ZN(n20191) );
  OR2_X1 U23094 ( .A1(n20181), .A2(n20180), .ZN(n20292) );
  OR2_X1 U23095 ( .A1(n20182), .A2(n20292), .ZN(n20184) );
  INV_X1 U23096 ( .A(n20208), .ZN(n20183) );
  AND2_X1 U23097 ( .A1(n20184), .A2(n20183), .ZN(n20190) );
  INV_X1 U23098 ( .A(n20190), .ZN(n20187) );
  OAI21_X1 U23099 ( .B1(n20697), .B2(n20185), .A(n20541), .ZN(n20186) );
  OAI211_X1 U23100 ( .C1(n20191), .C2(n20187), .A(n20546), .B(n20186), .ZN(
        n20210) );
  NAND2_X1 U23101 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20188), .ZN(
        n20189) );
  OAI22_X1 U23102 ( .A1(n20191), .A2(n20190), .B1(n20599), .B2(n20189), .ZN(
        n20209) );
  AOI22_X1 U23103 ( .A1(P1_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n20210), .B1(
        n20544), .B2(n20209), .ZN(n20192) );
  OAI211_X1 U23104 ( .C1(n20552), .C2(n20217), .A(n20193), .B(n20192), .ZN(
        P1_U3057) );
  AOI22_X1 U23105 ( .A1(n9663), .A2(n20208), .B1(n20235), .B2(n20505), .ZN(
        n20195) );
  AOI22_X1 U23106 ( .A1(P1_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n20210), .B1(
        n20553), .B2(n20209), .ZN(n20194) );
  OAI211_X1 U23107 ( .C1(n20508), .C2(n20206), .A(n20195), .B(n20194), .ZN(
        P1_U3058) );
  AOI22_X1 U23108 ( .A1(n20208), .A2(n20558), .B1(n20235), .B2(n20509), .ZN(
        n20197) );
  AOI22_X1 U23109 ( .A1(P1_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n20210), .B1(
        n20559), .B2(n20209), .ZN(n20196) );
  OAI211_X1 U23110 ( .C1(n20512), .C2(n20206), .A(n20197), .B(n20196), .ZN(
        P1_U3059) );
  AOI22_X1 U23111 ( .A1(n20208), .A2(n20564), .B1(n20207), .B2(n20566), .ZN(
        n20199) );
  AOI22_X1 U23112 ( .A1(P1_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n20210), .B1(
        n20565), .B2(n20209), .ZN(n20198) );
  OAI211_X1 U23113 ( .C1(n20569), .C2(n20217), .A(n20199), .B(n20198), .ZN(
        P1_U3060) );
  AOI22_X1 U23114 ( .A1(n20208), .A2(n20570), .B1(n20207), .B2(n20572), .ZN(
        n20201) );
  AOI22_X1 U23115 ( .A1(P1_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n20210), .B1(
        n20571), .B2(n20209), .ZN(n20200) );
  OAI211_X1 U23116 ( .C1(n20575), .C2(n20217), .A(n20201), .B(n20200), .ZN(
        P1_U3061) );
  AOI22_X1 U23117 ( .A1(n20208), .A2(n20576), .B1(n20235), .B2(n20521), .ZN(
        n20203) );
  AOI22_X1 U23118 ( .A1(P1_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n20210), .B1(
        n20577), .B2(n20209), .ZN(n20202) );
  OAI211_X1 U23119 ( .C1(n20524), .C2(n20206), .A(n20203), .B(n20202), .ZN(
        P1_U3062) );
  INV_X1 U23120 ( .A(n20585), .ZN(n20929) );
  AOI22_X1 U23121 ( .A1(n20208), .A2(n20926), .B1(n20235), .B2(n20929), .ZN(
        n20205) );
  AOI22_X1 U23122 ( .A1(P1_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n20210), .B1(
        n20928), .B2(n20209), .ZN(n20204) );
  OAI211_X1 U23123 ( .C1(n20935), .C2(n20206), .A(n20205), .B(n20204), .ZN(
        P1_U3063) );
  AOI22_X1 U23124 ( .A1(n20589), .A2(n20208), .B1(n20207), .B2(n20590), .ZN(
        n20212) );
  AOI22_X1 U23125 ( .A1(P1_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n20210), .B1(
        n20587), .B2(n20209), .ZN(n20211) );
  OAI211_X1 U23126 ( .C1(n20596), .C2(n20217), .A(n20212), .B(n20211), .ZN(
        P1_U3064) );
  INV_X1 U23127 ( .A(n20300), .ZN(n20296) );
  NOR2_X1 U23128 ( .A1(n13312), .A2(n20214), .ZN(n20293) );
  NAND2_X1 U23129 ( .A1(n20293), .A2(n20438), .ZN(n20216) );
  OAI22_X1 U23130 ( .A1(n20216), .A2(n20541), .B1(n20492), .B2(n20215), .ZN(
        n20234) );
  AOI22_X1 U23131 ( .A1(n20544), .A2(n20234), .B1(n20543), .B2(n9750), .ZN(
        n20221) );
  OAI221_X1 U23132 ( .B1(n20891), .B2(n20217), .C1(n20891), .C2(n20263), .A(
        n20216), .ZN(n20219) );
  AND2_X1 U23133 ( .A1(n20218), .A2(n20382), .ZN(n20499) );
  OAI221_X1 U23134 ( .B1(n9750), .B2(n20440), .C1(n9750), .C2(n20219), .A(
        n20499), .ZN(n20236) );
  AOI22_X1 U23135 ( .A1(P1_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n20236), .B1(
        n20235), .B2(n20549), .ZN(n20220) );
  OAI211_X1 U23136 ( .C1(n20552), .C2(n20263), .A(n20221), .B(n20220), .ZN(
        P1_U3065) );
  AOI22_X1 U23137 ( .A1(n9663), .A2(n9750), .B1(n20553), .B2(n20234), .ZN(
        n20223) );
  AOI22_X1 U23138 ( .A1(P1_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n20236), .B1(
        n20235), .B2(n20554), .ZN(n20222) );
  OAI211_X1 U23139 ( .C1(n20557), .C2(n20263), .A(n20223), .B(n20222), .ZN(
        P1_U3066) );
  AOI22_X1 U23140 ( .A1(n20559), .A2(n20234), .B1(n20558), .B2(n9750), .ZN(
        n20225) );
  AOI22_X1 U23141 ( .A1(P1_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n20236), .B1(
        n20235), .B2(n20560), .ZN(n20224) );
  OAI211_X1 U23142 ( .C1(n20563), .C2(n20263), .A(n20225), .B(n20224), .ZN(
        P1_U3067) );
  AOI22_X1 U23143 ( .A1(n20565), .A2(n20234), .B1(n20564), .B2(n9750), .ZN(
        n20227) );
  AOI22_X1 U23144 ( .A1(P1_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n20236), .B1(
        n20235), .B2(n20566), .ZN(n20226) );
  OAI211_X1 U23145 ( .C1(n20569), .C2(n20263), .A(n20227), .B(n20226), .ZN(
        P1_U3068) );
  AOI22_X1 U23146 ( .A1(n20571), .A2(n20234), .B1(n20570), .B2(n9750), .ZN(
        n20229) );
  AOI22_X1 U23147 ( .A1(P1_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n20236), .B1(
        n20235), .B2(n20572), .ZN(n20228) );
  OAI211_X1 U23148 ( .C1(n20575), .C2(n20263), .A(n20229), .B(n20228), .ZN(
        P1_U3069) );
  AOI22_X1 U23149 ( .A1(n20577), .A2(n20234), .B1(n20576), .B2(n9750), .ZN(
        n20231) );
  AOI22_X1 U23150 ( .A1(P1_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n20236), .B1(
        n20235), .B2(n20578), .ZN(n20230) );
  OAI211_X1 U23151 ( .C1(n20581), .C2(n20263), .A(n20231), .B(n20230), .ZN(
        P1_U3070) );
  AOI22_X1 U23152 ( .A1(n20928), .A2(n20234), .B1(n20926), .B2(n9750), .ZN(
        n20233) );
  AOI22_X1 U23153 ( .A1(P1_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n20236), .B1(
        n20235), .B2(n20582), .ZN(n20232) );
  OAI211_X1 U23154 ( .C1(n20585), .C2(n20263), .A(n20233), .B(n20232), .ZN(
        P1_U3071) );
  AOI22_X1 U23155 ( .A1(n20589), .A2(n9750), .B1(n20587), .B2(n20234), .ZN(
        n20238) );
  AOI22_X1 U23156 ( .A1(P1_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n20236), .B1(
        n20235), .B2(n20590), .ZN(n20237) );
  OAI211_X1 U23157 ( .C1(n20596), .C2(n20263), .A(n20238), .B(n20237), .ZN(
        P1_U3072) );
  NOR2_X1 U23158 ( .A1(n20264), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n20242) );
  INV_X1 U23159 ( .A(n20242), .ZN(n20239) );
  NOR2_X1 U23160 ( .A1(n20703), .A2(n20239), .ZN(n20259) );
  AOI21_X1 U23161 ( .B1(n20293), .B2(n20465), .A(n20259), .ZN(n20240) );
  OAI22_X1 U23162 ( .A1(n20240), .A2(n20541), .B1(n20239), .B2(n20599), .ZN(
        n20258) );
  AOI22_X1 U23163 ( .A1(n20544), .A2(n20258), .B1(n20543), .B2(n20259), .ZN(
        n20245) );
  OAI21_X1 U23164 ( .B1(n20300), .B2(n20469), .A(n20240), .ZN(n20241) );
  OAI221_X1 U23165 ( .B1(n20700), .B2(n20242), .C1(n20541), .C2(n20241), .A(
        n20546), .ZN(n20260) );
  NOR2_X2 U23166 ( .A1(n20300), .A2(n20464), .ZN(n20286) );
  AOI22_X1 U23167 ( .A1(P1_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n20260), .B1(
        n20286), .B2(n20501), .ZN(n20244) );
  OAI211_X1 U23168 ( .C1(n20504), .C2(n20263), .A(n20245), .B(n20244), .ZN(
        P1_U3073) );
  AOI22_X1 U23169 ( .A1(n9663), .A2(n20259), .B1(n20553), .B2(n20258), .ZN(
        n20247) );
  AOI22_X1 U23170 ( .A1(P1_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n20260), .B1(
        n20286), .B2(n20505), .ZN(n20246) );
  OAI211_X1 U23171 ( .C1(n20508), .C2(n20263), .A(n20247), .B(n20246), .ZN(
        P1_U3074) );
  AOI22_X1 U23172 ( .A1(n20559), .A2(n20258), .B1(n20558), .B2(n20259), .ZN(
        n20249) );
  AOI22_X1 U23173 ( .A1(P1_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n20260), .B1(
        n20286), .B2(n20509), .ZN(n20248) );
  OAI211_X1 U23174 ( .C1(n20512), .C2(n20263), .A(n20249), .B(n20248), .ZN(
        P1_U3075) );
  AOI22_X1 U23175 ( .A1(n20565), .A2(n20258), .B1(n20564), .B2(n20259), .ZN(
        n20251) );
  AOI22_X1 U23176 ( .A1(P1_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n20260), .B1(
        n20286), .B2(n20513), .ZN(n20250) );
  OAI211_X1 U23177 ( .C1(n20516), .C2(n20263), .A(n20251), .B(n20250), .ZN(
        P1_U3076) );
  AOI22_X1 U23178 ( .A1(n20571), .A2(n20258), .B1(n20570), .B2(n20259), .ZN(
        n20253) );
  AOI22_X1 U23179 ( .A1(P1_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n20260), .B1(
        n20286), .B2(n20517), .ZN(n20252) );
  OAI211_X1 U23180 ( .C1(n20520), .C2(n20263), .A(n20253), .B(n20252), .ZN(
        P1_U3077) );
  AOI22_X1 U23181 ( .A1(n20577), .A2(n20258), .B1(n20576), .B2(n20259), .ZN(
        n20255) );
  AOI22_X1 U23182 ( .A1(P1_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n20260), .B1(
        n20286), .B2(n20521), .ZN(n20254) );
  OAI211_X1 U23183 ( .C1(n20524), .C2(n20263), .A(n20255), .B(n20254), .ZN(
        P1_U3078) );
  AOI22_X1 U23184 ( .A1(n20928), .A2(n20258), .B1(n20926), .B2(n20259), .ZN(
        n20257) );
  AOI22_X1 U23185 ( .A1(P1_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n20260), .B1(
        n20286), .B2(n20929), .ZN(n20256) );
  OAI211_X1 U23186 ( .C1(n20935), .C2(n20263), .A(n20257), .B(n20256), .ZN(
        P1_U3079) );
  AOI22_X1 U23187 ( .A1(n20589), .A2(n20259), .B1(n20587), .B2(n20258), .ZN(
        n20262) );
  AOI22_X1 U23188 ( .A1(P1_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n20260), .B1(
        n20286), .B2(n20529), .ZN(n20261) );
  OAI211_X1 U23189 ( .C1(n20534), .C2(n20263), .A(n20262), .B(n20261), .ZN(
        P1_U3080) );
  INV_X1 U23190 ( .A(n20286), .ZN(n20279) );
  NOR2_X1 U23191 ( .A1(n20697), .A2(n20264), .ZN(n20299) );
  INV_X1 U23192 ( .A(n20299), .ZN(n20294) );
  NOR2_X1 U23193 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20294), .ZN(
        n20287) );
  AOI22_X1 U23194 ( .A1(n20287), .A2(n20543), .B1(n20311), .B2(n20501), .ZN(
        n20272) );
  AOI221_X1 U23195 ( .B1(n20286), .B2(P1_STATEBS16_REG_SCAN_IN), .C1(n20311), 
        .C2(P1_STATEBS16_REG_SCAN_IN), .A(n20541), .ZN(n20267) );
  NAND2_X1 U23196 ( .A1(n20293), .A2(n20695), .ZN(n20268) );
  AOI21_X1 U23197 ( .B1(n20267), .B2(n20268), .A(n20265), .ZN(n20266) );
  OAI211_X1 U23198 ( .C1(n20287), .C2(n20440), .A(n20499), .B(n20266), .ZN(
        n20289) );
  INV_X1 U23199 ( .A(n20267), .ZN(n20269) );
  OAI22_X1 U23200 ( .A1(n20492), .A2(n20270), .B1(n20269), .B2(n20268), .ZN(
        n20288) );
  AOI22_X1 U23201 ( .A1(P1_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n20289), .B1(
        n20544), .B2(n20288), .ZN(n20271) );
  OAI211_X1 U23202 ( .C1(n20504), .C2(n20279), .A(n20272), .B(n20271), .ZN(
        P1_U3081) );
  AOI22_X1 U23203 ( .A1(n9663), .A2(n20287), .B1(n20311), .B2(n20505), .ZN(
        n20274) );
  AOI22_X1 U23204 ( .A1(P1_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n20289), .B1(
        n20553), .B2(n20288), .ZN(n20273) );
  OAI211_X1 U23205 ( .C1(n20508), .C2(n20279), .A(n20274), .B(n20273), .ZN(
        P1_U3082) );
  AOI22_X1 U23206 ( .A1(n20287), .A2(n20558), .B1(n20311), .B2(n20509), .ZN(
        n20276) );
  AOI22_X1 U23207 ( .A1(P1_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n20289), .B1(
        n20559), .B2(n20288), .ZN(n20275) );
  OAI211_X1 U23208 ( .C1(n20512), .C2(n20279), .A(n20276), .B(n20275), .ZN(
        P1_U3083) );
  AOI22_X1 U23209 ( .A1(n20287), .A2(n20564), .B1(n20311), .B2(n20513), .ZN(
        n20278) );
  AOI22_X1 U23210 ( .A1(P1_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n20289), .B1(
        n20565), .B2(n20288), .ZN(n20277) );
  OAI211_X1 U23211 ( .C1(n20516), .C2(n20279), .A(n20278), .B(n20277), .ZN(
        P1_U3084) );
  AOI22_X1 U23212 ( .A1(n20287), .A2(n20570), .B1(n20286), .B2(n20572), .ZN(
        n20281) );
  AOI22_X1 U23213 ( .A1(P1_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n20289), .B1(
        n20571), .B2(n20288), .ZN(n20280) );
  OAI211_X1 U23214 ( .C1(n20575), .C2(n20321), .A(n20281), .B(n20280), .ZN(
        P1_U3085) );
  AOI22_X1 U23215 ( .A1(n20287), .A2(n20576), .B1(n20286), .B2(n20578), .ZN(
        n20283) );
  AOI22_X1 U23216 ( .A1(P1_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n20289), .B1(
        n20577), .B2(n20288), .ZN(n20282) );
  OAI211_X1 U23217 ( .C1(n20581), .C2(n20321), .A(n20283), .B(n20282), .ZN(
        P1_U3086) );
  AOI22_X1 U23218 ( .A1(n20926), .A2(n20287), .B1(n20286), .B2(n20582), .ZN(
        n20285) );
  AOI22_X1 U23219 ( .A1(P1_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n20289), .B1(
        n20928), .B2(n20288), .ZN(n20284) );
  OAI211_X1 U23220 ( .C1(n20585), .C2(n20321), .A(n20285), .B(n20284), .ZN(
        P1_U3087) );
  AOI22_X1 U23221 ( .A1(n20589), .A2(n20287), .B1(n20286), .B2(n20590), .ZN(
        n20291) );
  AOI22_X1 U23222 ( .A1(P1_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n20289), .B1(
        n20587), .B2(n20288), .ZN(n20290) );
  OAI211_X1 U23223 ( .C1(n20596), .C2(n20321), .A(n20291), .B(n20290), .ZN(
        P1_U3088) );
  INV_X1 U23224 ( .A(n20292), .ZN(n20537) );
  AOI21_X1 U23225 ( .B1(n20293), .B2(n20537), .A(n20317), .ZN(n20297) );
  OAI22_X1 U23226 ( .A1(n20297), .A2(n20541), .B1(n20294), .B2(n20599), .ZN(
        n20316) );
  AOI22_X1 U23227 ( .A1(n20317), .A2(n20543), .B1(n20544), .B2(n20316), .ZN(
        n20302) );
  INV_X1 U23228 ( .A(n20691), .ZN(n20295) );
  NAND2_X1 U23229 ( .A1(n20296), .A2(n20295), .ZN(n20682) );
  NAND2_X1 U23230 ( .A1(n20297), .A2(n20682), .ZN(n20298) );
  OAI221_X1 U23231 ( .B1(n20700), .B2(n20299), .C1(n20541), .C2(n20298), .A(
        n20546), .ZN(n20318) );
  NOR2_X2 U23232 ( .A1(n20300), .A2(n20411), .ZN(n20347) );
  AOI22_X1 U23233 ( .A1(P1_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n20318), .B1(
        n20347), .B2(n20501), .ZN(n20301) );
  OAI211_X1 U23234 ( .C1(n20504), .C2(n20321), .A(n20302), .B(n20301), .ZN(
        P1_U3089) );
  AOI22_X1 U23235 ( .A1(n9663), .A2(n20317), .B1(n20553), .B2(n20316), .ZN(
        n20304) );
  AOI22_X1 U23236 ( .A1(P1_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n20318), .B1(
        n20347), .B2(n20505), .ZN(n20303) );
  OAI211_X1 U23237 ( .C1(n20508), .C2(n20321), .A(n20304), .B(n20303), .ZN(
        P1_U3090) );
  INV_X1 U23238 ( .A(n20347), .ZN(n20330) );
  AOI22_X1 U23239 ( .A1(n20317), .A2(n20558), .B1(n20559), .B2(n20316), .ZN(
        n20306) );
  AOI22_X1 U23240 ( .A1(P1_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n20318), .B1(
        n20311), .B2(n20560), .ZN(n20305) );
  OAI211_X1 U23241 ( .C1(n20563), .C2(n20330), .A(n20306), .B(n20305), .ZN(
        P1_U3091) );
  AOI22_X1 U23242 ( .A1(n20317), .A2(n20564), .B1(n20565), .B2(n20316), .ZN(
        n20308) );
  AOI22_X1 U23243 ( .A1(P1_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n20318), .B1(
        n20311), .B2(n20566), .ZN(n20307) );
  OAI211_X1 U23244 ( .C1(n20569), .C2(n20330), .A(n20308), .B(n20307), .ZN(
        P1_U3092) );
  AOI22_X1 U23245 ( .A1(n20317), .A2(n20570), .B1(n20571), .B2(n20316), .ZN(
        n20310) );
  AOI22_X1 U23246 ( .A1(P1_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n20318), .B1(
        n20311), .B2(n20572), .ZN(n20309) );
  OAI211_X1 U23247 ( .C1(n20575), .C2(n20330), .A(n20310), .B(n20309), .ZN(
        P1_U3093) );
  AOI22_X1 U23248 ( .A1(n20317), .A2(n20576), .B1(n20577), .B2(n20316), .ZN(
        n20313) );
  AOI22_X1 U23249 ( .A1(P1_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n20318), .B1(
        n20311), .B2(n20578), .ZN(n20312) );
  OAI211_X1 U23250 ( .C1(n20581), .C2(n20330), .A(n20313), .B(n20312), .ZN(
        P1_U3094) );
  AOI22_X1 U23251 ( .A1(n20317), .A2(n20926), .B1(n20928), .B2(n20316), .ZN(
        n20315) );
  AOI22_X1 U23252 ( .A1(P1_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n20318), .B1(
        n20347), .B2(n20929), .ZN(n20314) );
  OAI211_X1 U23253 ( .C1(n20935), .C2(n20321), .A(n20315), .B(n20314), .ZN(
        P1_U3095) );
  AOI22_X1 U23254 ( .A1(n20589), .A2(n20317), .B1(n20587), .B2(n20316), .ZN(
        n20320) );
  AOI22_X1 U23255 ( .A1(P1_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n20318), .B1(
        n20347), .B2(n20529), .ZN(n20319) );
  OAI211_X1 U23256 ( .C1(n20534), .C2(n20321), .A(n20320), .B(n20319), .ZN(
        P1_U3096) );
  INV_X1 U23257 ( .A(n13434), .ZN(n20322) );
  INV_X1 U23258 ( .A(n20681), .ZN(n20323) );
  NOR2_X1 U23259 ( .A1(n20325), .A2(n20324), .ZN(n20406) );
  NAND2_X1 U23260 ( .A1(n20326), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n20404) );
  AOI21_X1 U23261 ( .B1(n20406), .B2(n20438), .A(n10121), .ZN(n20329) );
  INV_X1 U23262 ( .A(n20327), .ZN(n20328) );
  NAND2_X1 U23263 ( .A1(n20378), .A2(n20328), .ZN(n20444) );
  OAI22_X1 U23264 ( .A1(n20329), .A2(n20541), .B1(n20444), .B2(n20382), .ZN(
        n20346) );
  AOI22_X1 U23265 ( .A1(n20544), .A2(n20346), .B1(n20543), .B2(n10121), .ZN(
        n20333) );
  OAI221_X1 U23266 ( .B1(n20891), .B2(n20374), .C1(n20891), .C2(n20330), .A(
        n20329), .ZN(n20331) );
  AOI22_X1 U23267 ( .A1(P1_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n20348), .B1(
        n20347), .B2(n20549), .ZN(n20332) );
  OAI211_X1 U23268 ( .C1(n20552), .C2(n20374), .A(n20333), .B(n20332), .ZN(
        P1_U3097) );
  AOI22_X1 U23269 ( .A1(n9663), .A2(n10121), .B1(n20553), .B2(n20346), .ZN(
        n20335) );
  AOI22_X1 U23270 ( .A1(P1_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n20348), .B1(
        n20347), .B2(n20554), .ZN(n20334) );
  OAI211_X1 U23271 ( .C1(n20557), .C2(n20374), .A(n20335), .B(n20334), .ZN(
        P1_U3098) );
  AOI22_X1 U23272 ( .A1(n20559), .A2(n20346), .B1(n20558), .B2(n10121), .ZN(
        n20337) );
  AOI22_X1 U23273 ( .A1(P1_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n20348), .B1(
        n20347), .B2(n20560), .ZN(n20336) );
  OAI211_X1 U23274 ( .C1(n20563), .C2(n20374), .A(n20337), .B(n20336), .ZN(
        P1_U3099) );
  AOI22_X1 U23275 ( .A1(n20565), .A2(n20346), .B1(n20564), .B2(n10121), .ZN(
        n20339) );
  AOI22_X1 U23276 ( .A1(P1_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n20348), .B1(
        n20347), .B2(n20566), .ZN(n20338) );
  OAI211_X1 U23277 ( .C1(n20569), .C2(n20374), .A(n20339), .B(n20338), .ZN(
        P1_U3100) );
  AOI22_X1 U23278 ( .A1(n20571), .A2(n20346), .B1(n20570), .B2(n10121), .ZN(
        n20341) );
  AOI22_X1 U23279 ( .A1(P1_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n20348), .B1(
        n20347), .B2(n20572), .ZN(n20340) );
  OAI211_X1 U23280 ( .C1(n20575), .C2(n20374), .A(n20341), .B(n20340), .ZN(
        P1_U3101) );
  AOI22_X1 U23281 ( .A1(n20577), .A2(n20346), .B1(n20576), .B2(n10121), .ZN(
        n20343) );
  AOI22_X1 U23282 ( .A1(P1_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n20348), .B1(
        n20347), .B2(n20578), .ZN(n20342) );
  OAI211_X1 U23283 ( .C1(n20581), .C2(n20374), .A(n20343), .B(n20342), .ZN(
        P1_U3102) );
  AOI22_X1 U23284 ( .A1(n20928), .A2(n20346), .B1(n20926), .B2(n10121), .ZN(
        n20345) );
  AOI22_X1 U23285 ( .A1(P1_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n20348), .B1(
        n20347), .B2(n20582), .ZN(n20344) );
  OAI211_X1 U23286 ( .C1(n20585), .C2(n20374), .A(n20345), .B(n20344), .ZN(
        P1_U3103) );
  AOI22_X1 U23287 ( .A1(n20589), .A2(n10121), .B1(n20587), .B2(n20346), .ZN(
        n20350) );
  AOI22_X1 U23288 ( .A1(P1_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n20348), .B1(
        n20347), .B2(n20590), .ZN(n20349) );
  OAI211_X1 U23289 ( .C1(n20596), .C2(n20374), .A(n20350), .B(n20349), .ZN(
        P1_U3104) );
  NOR2_X1 U23290 ( .A1(n20404), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n20354) );
  INV_X1 U23291 ( .A(n20354), .ZN(n20351) );
  NOR2_X1 U23292 ( .A1(n20703), .A2(n20351), .ZN(n20370) );
  AOI21_X1 U23293 ( .B1(n20406), .B2(n20465), .A(n20370), .ZN(n20352) );
  OAI22_X1 U23294 ( .A1(n20352), .A2(n20541), .B1(n20351), .B2(n20599), .ZN(
        n20369) );
  AOI22_X1 U23295 ( .A1(n20544), .A2(n20369), .B1(n20543), .B2(n20370), .ZN(
        n20356) );
  OAI211_X1 U23296 ( .C1(n20681), .C2(n20469), .A(n20700), .B(n20352), .ZN(
        n20353) );
  OAI211_X1 U23297 ( .C1(n20700), .C2(n20354), .A(n20546), .B(n20353), .ZN(
        n20371) );
  NOR2_X2 U23298 ( .A1(n20681), .A2(n20464), .ZN(n20389) );
  AOI22_X1 U23299 ( .A1(P1_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n20371), .B1(
        n20389), .B2(n20501), .ZN(n20355) );
  OAI211_X1 U23300 ( .C1(n20504), .C2(n20374), .A(n20356), .B(n20355), .ZN(
        P1_U3105) );
  AOI22_X1 U23301 ( .A1(n9663), .A2(n20370), .B1(n20553), .B2(n20369), .ZN(
        n20358) );
  AOI22_X1 U23302 ( .A1(P1_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n20371), .B1(
        n20389), .B2(n20505), .ZN(n20357) );
  OAI211_X1 U23303 ( .C1(n20508), .C2(n20374), .A(n20358), .B(n20357), .ZN(
        P1_U3106) );
  AOI22_X1 U23304 ( .A1(n20559), .A2(n20369), .B1(n20558), .B2(n20370), .ZN(
        n20360) );
  AOI22_X1 U23305 ( .A1(P1_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n20371), .B1(
        n20389), .B2(n20509), .ZN(n20359) );
  OAI211_X1 U23306 ( .C1(n20512), .C2(n20374), .A(n20360), .B(n20359), .ZN(
        P1_U3107) );
  AOI22_X1 U23307 ( .A1(n20565), .A2(n20369), .B1(n20564), .B2(n20370), .ZN(
        n20362) );
  AOI22_X1 U23308 ( .A1(P1_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n20371), .B1(
        n20389), .B2(n20513), .ZN(n20361) );
  OAI211_X1 U23309 ( .C1(n20516), .C2(n20374), .A(n20362), .B(n20361), .ZN(
        P1_U3108) );
  AOI22_X1 U23310 ( .A1(n20571), .A2(n20369), .B1(n20570), .B2(n20370), .ZN(
        n20364) );
  AOI22_X1 U23311 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n20371), .B1(
        n20389), .B2(n20517), .ZN(n20363) );
  OAI211_X1 U23312 ( .C1(n20520), .C2(n20374), .A(n20364), .B(n20363), .ZN(
        P1_U3109) );
  AOI22_X1 U23313 ( .A1(n20577), .A2(n20369), .B1(n20576), .B2(n20370), .ZN(
        n20366) );
  AOI22_X1 U23314 ( .A1(P1_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n20371), .B1(
        n20389), .B2(n20521), .ZN(n20365) );
  OAI211_X1 U23315 ( .C1(n20524), .C2(n20374), .A(n20366), .B(n20365), .ZN(
        P1_U3110) );
  AOI22_X1 U23316 ( .A1(n20928), .A2(n20369), .B1(n20926), .B2(n20370), .ZN(
        n20368) );
  AOI22_X1 U23317 ( .A1(P1_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n20371), .B1(
        n20389), .B2(n20929), .ZN(n20367) );
  OAI211_X1 U23318 ( .C1(n20935), .C2(n20374), .A(n20368), .B(n20367), .ZN(
        P1_U3111) );
  AOI22_X1 U23319 ( .A1(n20589), .A2(n20370), .B1(n20587), .B2(n20369), .ZN(
        n20373) );
  AOI22_X1 U23320 ( .A1(P1_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n20371), .B1(
        n20389), .B2(n20529), .ZN(n20372) );
  OAI211_X1 U23321 ( .C1(n20534), .C2(n20374), .A(n20373), .B(n20372), .ZN(
        P1_U3112) );
  INV_X1 U23322 ( .A(n20389), .ZN(n20403) );
  NOR2_X1 U23323 ( .A1(n20697), .A2(n20404), .ZN(n20410) );
  INV_X1 U23324 ( .A(n20410), .ZN(n20407) );
  NOR2_X1 U23325 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20407), .ZN(
        n20398) );
  AOI22_X1 U23326 ( .A1(n20398), .A2(n20543), .B1(n20424), .B2(n20501), .ZN(
        n20384) );
  INV_X1 U23327 ( .A(n20398), .ZN(n20375) );
  AOI221_X1 U23328 ( .B1(n20389), .B2(P1_STATEBS16_REG_SCAN_IN), .C1(n20424), 
        .C2(P1_STATEBS16_REG_SCAN_IN), .A(n20541), .ZN(n20379) );
  NAND2_X1 U23329 ( .A1(n20406), .A2(n20695), .ZN(n20381) );
  AOI22_X1 U23330 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n20375), .B1(n20379), 
        .B2(n20381), .ZN(n20376) );
  OAI21_X1 U23331 ( .B1(n20690), .B2(n20378), .A(P1_STATE2_REG_2__SCAN_IN), 
        .ZN(n20498) );
  NAND3_X1 U23332 ( .A1(n20377), .A2(n20376), .A3(n20498), .ZN(n20400) );
  OR2_X1 U23333 ( .A1(n20690), .A2(n20378), .ZN(n20491) );
  INV_X1 U23334 ( .A(n20379), .ZN(n20380) );
  AOI22_X1 U23335 ( .A1(P1_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n20400), .B1(
        n20544), .B2(n20399), .ZN(n20383) );
  OAI211_X1 U23336 ( .C1(n20504), .C2(n20403), .A(n20384), .B(n20383), .ZN(
        P1_U3113) );
  AOI22_X1 U23337 ( .A1(n9663), .A2(n20398), .B1(n20389), .B2(n20554), .ZN(
        n20386) );
  AOI22_X1 U23338 ( .A1(P1_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n20400), .B1(
        n20553), .B2(n20399), .ZN(n20385) );
  OAI211_X1 U23339 ( .C1(n20557), .C2(n20432), .A(n20386), .B(n20385), .ZN(
        P1_U3114) );
  AOI22_X1 U23340 ( .A1(n20398), .A2(n20558), .B1(n20389), .B2(n20560), .ZN(
        n20388) );
  AOI22_X1 U23341 ( .A1(P1_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n20400), .B1(
        n20559), .B2(n20399), .ZN(n20387) );
  OAI211_X1 U23342 ( .C1(n20563), .C2(n20432), .A(n20388), .B(n20387), .ZN(
        P1_U3115) );
  AOI22_X1 U23343 ( .A1(n20398), .A2(n20564), .B1(n20389), .B2(n20566), .ZN(
        n20391) );
  AOI22_X1 U23344 ( .A1(P1_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n20400), .B1(
        n20565), .B2(n20399), .ZN(n20390) );
  OAI211_X1 U23345 ( .C1(n20569), .C2(n20432), .A(n20391), .B(n20390), .ZN(
        P1_U3116) );
  AOI22_X1 U23346 ( .A1(n20398), .A2(n20570), .B1(n20424), .B2(n20517), .ZN(
        n20393) );
  AOI22_X1 U23347 ( .A1(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n20400), .B1(
        n20571), .B2(n20399), .ZN(n20392) );
  OAI211_X1 U23348 ( .C1(n20520), .C2(n20403), .A(n20393), .B(n20392), .ZN(
        P1_U3117) );
  AOI22_X1 U23349 ( .A1(n20398), .A2(n20576), .B1(n20424), .B2(n20521), .ZN(
        n20395) );
  AOI22_X1 U23350 ( .A1(P1_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n20400), .B1(
        n20577), .B2(n20399), .ZN(n20394) );
  OAI211_X1 U23351 ( .C1(n20524), .C2(n20403), .A(n20395), .B(n20394), .ZN(
        P1_U3118) );
  AOI22_X1 U23352 ( .A1(n20398), .A2(n20926), .B1(n20424), .B2(n20929), .ZN(
        n20397) );
  AOI22_X1 U23353 ( .A1(P1_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n20400), .B1(
        n20928), .B2(n20399), .ZN(n20396) );
  OAI211_X1 U23354 ( .C1(n20935), .C2(n20403), .A(n20397), .B(n20396), .ZN(
        P1_U3119) );
  AOI22_X1 U23355 ( .A1(n20589), .A2(n20398), .B1(n20424), .B2(n20529), .ZN(
        n20402) );
  AOI22_X1 U23356 ( .A1(P1_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n20400), .B1(
        n20587), .B2(n20399), .ZN(n20401) );
  OAI211_X1 U23357 ( .C1(n20534), .C2(n20403), .A(n20402), .B(n20401), .ZN(
        P1_U3120) );
  INV_X1 U23358 ( .A(n20404), .ZN(n20405) );
  AND2_X1 U23359 ( .A1(n20536), .A2(n20405), .ZN(n20428) );
  AOI21_X1 U23360 ( .B1(n20406), .B2(n20537), .A(n20428), .ZN(n20408) );
  OAI22_X1 U23361 ( .A1(n20408), .A2(n20541), .B1(n20407), .B2(n20599), .ZN(
        n20427) );
  AOI22_X1 U23362 ( .A1(n20544), .A2(n20427), .B1(n20543), .B2(n20428), .ZN(
        n20413) );
  OAI211_X1 U23363 ( .C1(n20681), .C2(n20691), .A(n20700), .B(n20408), .ZN(
        n20409) );
  OAI211_X1 U23364 ( .C1(n20700), .C2(n20410), .A(n20546), .B(n20409), .ZN(
        n20429) );
  AOI22_X1 U23365 ( .A1(P1_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n20429), .B1(
        n20436), .B2(n20501), .ZN(n20412) );
  OAI211_X1 U23366 ( .C1(n20504), .C2(n20432), .A(n20413), .B(n20412), .ZN(
        P1_U3121) );
  AOI22_X1 U23367 ( .A1(n9663), .A2(n20428), .B1(n20553), .B2(n20427), .ZN(
        n20415) );
  AOI22_X1 U23368 ( .A1(P1_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n20429), .B1(
        n20424), .B2(n20554), .ZN(n20414) );
  OAI211_X1 U23369 ( .C1(n20557), .C2(n20463), .A(n20415), .B(n20414), .ZN(
        P1_U3122) );
  AOI22_X1 U23370 ( .A1(n20559), .A2(n20427), .B1(n20558), .B2(n20428), .ZN(
        n20417) );
  AOI22_X1 U23371 ( .A1(P1_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n20429), .B1(
        n20424), .B2(n20560), .ZN(n20416) );
  OAI211_X1 U23372 ( .C1(n20563), .C2(n20463), .A(n20417), .B(n20416), .ZN(
        P1_U3123) );
  AOI22_X1 U23373 ( .A1(n20565), .A2(n20427), .B1(n20564), .B2(n20428), .ZN(
        n20419) );
  AOI22_X1 U23374 ( .A1(P1_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n20429), .B1(
        n20424), .B2(n20566), .ZN(n20418) );
  OAI211_X1 U23375 ( .C1(n20569), .C2(n20463), .A(n20419), .B(n20418), .ZN(
        P1_U3124) );
  AOI22_X1 U23376 ( .A1(n20571), .A2(n20427), .B1(n20570), .B2(n20428), .ZN(
        n20421) );
  AOI22_X1 U23377 ( .A1(P1_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n20429), .B1(
        n20436), .B2(n20517), .ZN(n20420) );
  OAI211_X1 U23378 ( .C1(n20520), .C2(n20432), .A(n20421), .B(n20420), .ZN(
        P1_U3125) );
  AOI22_X1 U23379 ( .A1(n20577), .A2(n20427), .B1(n20576), .B2(n20428), .ZN(
        n20423) );
  AOI22_X1 U23380 ( .A1(P1_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n20429), .B1(
        n20436), .B2(n20521), .ZN(n20422) );
  OAI211_X1 U23381 ( .C1(n20524), .C2(n20432), .A(n20423), .B(n20422), .ZN(
        P1_U3126) );
  AOI22_X1 U23382 ( .A1(n20928), .A2(n20427), .B1(n20926), .B2(n20428), .ZN(
        n20426) );
  AOI22_X1 U23383 ( .A1(P1_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n20429), .B1(
        n20424), .B2(n20582), .ZN(n20425) );
  OAI211_X1 U23384 ( .C1(n20585), .C2(n20463), .A(n20426), .B(n20425), .ZN(
        P1_U3127) );
  AOI22_X1 U23385 ( .A1(n20589), .A2(n20428), .B1(n20587), .B2(n20427), .ZN(
        n20431) );
  AOI22_X1 U23386 ( .A1(P1_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n20429), .B1(
        n20436), .B2(n20529), .ZN(n20430) );
  OAI211_X1 U23387 ( .C1(n20534), .C2(n20432), .A(n20431), .B(n20430), .ZN(
        P1_U3128) );
  NAND2_X1 U23388 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20539) );
  INV_X1 U23389 ( .A(n20434), .ZN(n20435) );
  NOR2_X2 U23390 ( .A1(n20494), .A2(n20435), .ZN(n20487) );
  AOI22_X1 U23391 ( .A1(n9751), .A2(n20543), .B1(n20487), .B2(n20501), .ZN(
        n20446) );
  AOI221_X1 U23392 ( .B1(n20436), .B2(P1_STATEBS16_REG_SCAN_IN), .C1(n20487), 
        .C2(P1_STATEBS16_REG_SCAN_IN), .A(n20541), .ZN(n20441) );
  NOR2_X1 U23393 ( .A1(n13312), .A2(n20437), .ZN(n20538) );
  NAND2_X1 U23394 ( .A1(n20538), .A2(n20438), .ZN(n20443) );
  AOI22_X1 U23395 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n20444), .B1(n20441), 
        .B2(n20443), .ZN(n20439) );
  OAI211_X1 U23396 ( .C1(n9751), .C2(n20440), .A(n20499), .B(n20439), .ZN(
        n20460) );
  INV_X1 U23397 ( .A(n20441), .ZN(n20442) );
  AOI22_X1 U23398 ( .A1(P1_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n20460), .B1(
        n20544), .B2(n20459), .ZN(n20445) );
  OAI211_X1 U23399 ( .C1(n20504), .C2(n20463), .A(n20446), .B(n20445), .ZN(
        P1_U3129) );
  AOI22_X1 U23400 ( .A1(n9663), .A2(n9751), .B1(n20487), .B2(n20505), .ZN(
        n20448) );
  AOI22_X1 U23401 ( .A1(P1_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n20460), .B1(
        n20553), .B2(n20459), .ZN(n20447) );
  OAI211_X1 U23402 ( .C1(n20508), .C2(n20463), .A(n20448), .B(n20447), .ZN(
        P1_U3130) );
  AOI22_X1 U23403 ( .A1(n9751), .A2(n20558), .B1(n20487), .B2(n20509), .ZN(
        n20450) );
  AOI22_X1 U23404 ( .A1(P1_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n20460), .B1(
        n20559), .B2(n20459), .ZN(n20449) );
  OAI211_X1 U23405 ( .C1(n20512), .C2(n20463), .A(n20450), .B(n20449), .ZN(
        P1_U3131) );
  AOI22_X1 U23406 ( .A1(n9751), .A2(n20564), .B1(n20487), .B2(n20513), .ZN(
        n20452) );
  AOI22_X1 U23407 ( .A1(P1_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n20460), .B1(
        n20565), .B2(n20459), .ZN(n20451) );
  OAI211_X1 U23408 ( .C1(n20516), .C2(n20463), .A(n20452), .B(n20451), .ZN(
        P1_U3132) );
  AOI22_X1 U23409 ( .A1(n9751), .A2(n20570), .B1(n20487), .B2(n20517), .ZN(
        n20454) );
  AOI22_X1 U23410 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n20460), .B1(
        n20571), .B2(n20459), .ZN(n20453) );
  OAI211_X1 U23411 ( .C1(n20520), .C2(n20463), .A(n20454), .B(n20453), .ZN(
        P1_U3133) );
  AOI22_X1 U23412 ( .A1(n9751), .A2(n20576), .B1(n20487), .B2(n20521), .ZN(
        n20456) );
  AOI22_X1 U23413 ( .A1(P1_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n20460), .B1(
        n20577), .B2(n20459), .ZN(n20455) );
  OAI211_X1 U23414 ( .C1(n20524), .C2(n20463), .A(n20456), .B(n20455), .ZN(
        P1_U3134) );
  AOI22_X1 U23415 ( .A1(n9751), .A2(n20926), .B1(n20487), .B2(n20929), .ZN(
        n20458) );
  AOI22_X1 U23416 ( .A1(P1_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n20460), .B1(
        n20928), .B2(n20459), .ZN(n20457) );
  OAI211_X1 U23417 ( .C1(n20935), .C2(n20463), .A(n20458), .B(n20457), .ZN(
        P1_U3135) );
  AOI22_X1 U23418 ( .A1(n20589), .A2(n9751), .B1(n20487), .B2(n20529), .ZN(
        n20462) );
  AOI22_X1 U23419 ( .A1(P1_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n20460), .B1(
        n20587), .B2(n20459), .ZN(n20461) );
  OAI211_X1 U23420 ( .C1(n20534), .C2(n20463), .A(n20462), .B(n20461), .ZN(
        P1_U3136) );
  NOR2_X1 U23421 ( .A1(n20494), .A2(n20464), .ZN(n20495) );
  AOI21_X1 U23422 ( .B1(n20538), .B2(n20465), .A(n20486), .ZN(n20467) );
  NOR2_X1 U23423 ( .A1(n20539), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n20470) );
  INV_X1 U23424 ( .A(n20470), .ZN(n20466) );
  OAI22_X1 U23425 ( .A1(n20467), .A2(n20541), .B1(n20466), .B2(n20599), .ZN(
        n20485) );
  AOI22_X1 U23426 ( .A1(n20544), .A2(n20485), .B1(n20543), .B2(n20486), .ZN(
        n20472) );
  INV_X1 U23427 ( .A(n20494), .ZN(n20468) );
  NAND2_X1 U23428 ( .A1(n20468), .A2(n20700), .ZN(n20545) );
  NOR2_X1 U23429 ( .A1(n20545), .A2(n20469), .ZN(n20687) );
  OAI21_X1 U23430 ( .B1(n20687), .B2(n20470), .A(n20546), .ZN(n20488) );
  AOI22_X1 U23431 ( .A1(P1_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n20488), .B1(
        n20487), .B2(n20549), .ZN(n20471) );
  OAI211_X1 U23432 ( .C1(n20552), .C2(n20533), .A(n20472), .B(n20471), .ZN(
        P1_U3137) );
  AOI22_X1 U23433 ( .A1(n9663), .A2(n20486), .B1(n20553), .B2(n20485), .ZN(
        n20474) );
  AOI22_X1 U23434 ( .A1(P1_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n20488), .B1(
        n20487), .B2(n20554), .ZN(n20473) );
  OAI211_X1 U23435 ( .C1(n20557), .C2(n20533), .A(n20474), .B(n20473), .ZN(
        P1_U3138) );
  AOI22_X1 U23436 ( .A1(n20559), .A2(n20485), .B1(n20558), .B2(n20486), .ZN(
        n20476) );
  AOI22_X1 U23437 ( .A1(P1_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n20488), .B1(
        n20487), .B2(n20560), .ZN(n20475) );
  OAI211_X1 U23438 ( .C1(n20563), .C2(n20533), .A(n20476), .B(n20475), .ZN(
        P1_U3139) );
  AOI22_X1 U23439 ( .A1(n20565), .A2(n20485), .B1(n20564), .B2(n20486), .ZN(
        n20478) );
  AOI22_X1 U23440 ( .A1(P1_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n20488), .B1(
        n20487), .B2(n20566), .ZN(n20477) );
  OAI211_X1 U23441 ( .C1(n20569), .C2(n20533), .A(n20478), .B(n20477), .ZN(
        P1_U3140) );
  AOI22_X1 U23442 ( .A1(n20571), .A2(n20485), .B1(n20570), .B2(n20486), .ZN(
        n20480) );
  AOI22_X1 U23443 ( .A1(P1_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n20488), .B1(
        n20487), .B2(n20572), .ZN(n20479) );
  OAI211_X1 U23444 ( .C1(n20575), .C2(n20533), .A(n20480), .B(n20479), .ZN(
        P1_U3141) );
  AOI22_X1 U23445 ( .A1(n20577), .A2(n20485), .B1(n20576), .B2(n20486), .ZN(
        n20482) );
  AOI22_X1 U23446 ( .A1(P1_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n20488), .B1(
        n20487), .B2(n20578), .ZN(n20481) );
  OAI211_X1 U23447 ( .C1(n20581), .C2(n20533), .A(n20482), .B(n20481), .ZN(
        P1_U3142) );
  AOI22_X1 U23448 ( .A1(n20928), .A2(n20485), .B1(n20926), .B2(n20486), .ZN(
        n20484) );
  AOI22_X1 U23449 ( .A1(P1_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n20488), .B1(
        n20487), .B2(n20582), .ZN(n20483) );
  OAI211_X1 U23450 ( .C1(n20585), .C2(n20533), .A(n20484), .B(n20483), .ZN(
        P1_U3143) );
  AOI22_X1 U23451 ( .A1(n20589), .A2(n20486), .B1(n20587), .B2(n20485), .ZN(
        n20490) );
  AOI22_X1 U23452 ( .A1(P1_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n20488), .B1(
        n20487), .B2(n20590), .ZN(n20489) );
  OAI211_X1 U23453 ( .C1(n20596), .C2(n20533), .A(n20490), .B(n20489), .ZN(
        P1_U3144) );
  NAND2_X1 U23454 ( .A1(n20538), .A2(n20695), .ZN(n20497) );
  OAI22_X1 U23455 ( .A1(n20497), .A2(n20541), .B1(n20492), .B2(n20491), .ZN(
        n20527) );
  NOR3_X2 U23456 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20697), .A3(
        n20539), .ZN(n20528) );
  AOI22_X1 U23457 ( .A1(n20544), .A2(n20527), .B1(n20543), .B2(n20528), .ZN(
        n20503) );
  NOR2_X2 U23458 ( .A1(n20494), .A2(n20493), .ZN(n20591) );
  OAI21_X1 U23459 ( .B1(n20495), .B2(n20591), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20496) );
  AOI21_X1 U23460 ( .B1(n20497), .B2(n20496), .A(P1_STATE2_REG_3__SCAN_IN), 
        .ZN(n20500) );
  AOI22_X1 U23461 ( .A1(P1_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n20530), .B1(
        n20591), .B2(n20501), .ZN(n20502) );
  OAI211_X1 U23462 ( .C1(n20504), .C2(n20533), .A(n20503), .B(n20502), .ZN(
        P1_U3145) );
  AOI22_X1 U23463 ( .A1(n9663), .A2(n20528), .B1(n20553), .B2(n20527), .ZN(
        n20507) );
  AOI22_X1 U23464 ( .A1(P1_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n20530), .B1(
        n20591), .B2(n20505), .ZN(n20506) );
  OAI211_X1 U23465 ( .C1(n20508), .C2(n20533), .A(n20507), .B(n20506), .ZN(
        P1_U3146) );
  AOI22_X1 U23466 ( .A1(n20559), .A2(n20527), .B1(n20558), .B2(n20528), .ZN(
        n20511) );
  AOI22_X1 U23467 ( .A1(P1_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n20530), .B1(
        n20591), .B2(n20509), .ZN(n20510) );
  OAI211_X1 U23468 ( .C1(n20512), .C2(n20533), .A(n20511), .B(n20510), .ZN(
        P1_U3147) );
  AOI22_X1 U23469 ( .A1(n20565), .A2(n20527), .B1(n20564), .B2(n20528), .ZN(
        n20515) );
  AOI22_X1 U23470 ( .A1(P1_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n20530), .B1(
        n20591), .B2(n20513), .ZN(n20514) );
  OAI211_X1 U23471 ( .C1(n20516), .C2(n20533), .A(n20515), .B(n20514), .ZN(
        P1_U3148) );
  AOI22_X1 U23472 ( .A1(n20571), .A2(n20527), .B1(n20570), .B2(n20528), .ZN(
        n20519) );
  AOI22_X1 U23473 ( .A1(P1_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n20530), .B1(
        n20591), .B2(n20517), .ZN(n20518) );
  OAI211_X1 U23474 ( .C1(n20520), .C2(n20533), .A(n20519), .B(n20518), .ZN(
        P1_U3149) );
  AOI22_X1 U23475 ( .A1(n20577), .A2(n20527), .B1(n20576), .B2(n20528), .ZN(
        n20523) );
  AOI22_X1 U23476 ( .A1(P1_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n20530), .B1(
        n20591), .B2(n20521), .ZN(n20522) );
  OAI211_X1 U23477 ( .C1(n20524), .C2(n20533), .A(n20523), .B(n20522), .ZN(
        P1_U3150) );
  AOI22_X1 U23478 ( .A1(n20928), .A2(n20527), .B1(n20926), .B2(n20528), .ZN(
        n20526) );
  AOI22_X1 U23479 ( .A1(P1_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n20530), .B1(
        n20591), .B2(n20929), .ZN(n20525) );
  OAI211_X1 U23480 ( .C1(n20935), .C2(n20533), .A(n20526), .B(n20525), .ZN(
        P1_U3151) );
  AOI22_X1 U23481 ( .A1(n20589), .A2(n20528), .B1(n20587), .B2(n20527), .ZN(
        n20532) );
  AOI22_X1 U23482 ( .A1(P1_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n20530), .B1(
        n20591), .B2(n20529), .ZN(n20531) );
  OAI211_X1 U23483 ( .C1(n20534), .C2(n20533), .A(n20532), .B(n20531), .ZN(
        P1_U3152) );
  INV_X1 U23484 ( .A(n20539), .ZN(n20535) );
  AND2_X1 U23485 ( .A1(n20536), .A2(n20535), .ZN(n20588) );
  AOI21_X1 U23486 ( .B1(n20538), .B2(n20537), .A(n20588), .ZN(n20542) );
  NOR2_X1 U23487 ( .A1(n20697), .A2(n20539), .ZN(n20547) );
  INV_X1 U23488 ( .A(n20547), .ZN(n20540) );
  OAI22_X1 U23489 ( .A1(n20542), .A2(n20541), .B1(n20540), .B2(n20599), .ZN(
        n20586) );
  AOI22_X1 U23490 ( .A1(n20544), .A2(n20586), .B1(n20543), .B2(n20588), .ZN(
        n20551) );
  NOR2_X1 U23491 ( .A1(n20545), .A2(n20691), .ZN(n20548) );
  OAI21_X1 U23492 ( .B1(n20548), .B2(n20547), .A(n20546), .ZN(n20592) );
  AOI22_X1 U23493 ( .A1(P1_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n20592), .B1(
        n20591), .B2(n20549), .ZN(n20550) );
  OAI211_X1 U23494 ( .C1(n20552), .C2(n20595), .A(n20551), .B(n20550), .ZN(
        P1_U3153) );
  AOI22_X1 U23495 ( .A1(n9663), .A2(n20588), .B1(n20553), .B2(n20586), .ZN(
        n20556) );
  AOI22_X1 U23496 ( .A1(P1_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n20592), .B1(
        n20591), .B2(n20554), .ZN(n20555) );
  OAI211_X1 U23497 ( .C1(n20557), .C2(n20595), .A(n20556), .B(n20555), .ZN(
        P1_U3154) );
  AOI22_X1 U23498 ( .A1(n20559), .A2(n20586), .B1(n20558), .B2(n20588), .ZN(
        n20562) );
  AOI22_X1 U23499 ( .A1(P1_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n20592), .B1(
        n20591), .B2(n20560), .ZN(n20561) );
  OAI211_X1 U23500 ( .C1(n20563), .C2(n20595), .A(n20562), .B(n20561), .ZN(
        P1_U3155) );
  AOI22_X1 U23501 ( .A1(n20565), .A2(n20586), .B1(n20564), .B2(n20588), .ZN(
        n20568) );
  AOI22_X1 U23502 ( .A1(P1_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n20592), .B1(
        n20591), .B2(n20566), .ZN(n20567) );
  OAI211_X1 U23503 ( .C1(n20569), .C2(n20595), .A(n20568), .B(n20567), .ZN(
        P1_U3156) );
  AOI22_X1 U23504 ( .A1(n20571), .A2(n20586), .B1(n20570), .B2(n20588), .ZN(
        n20574) );
  AOI22_X1 U23505 ( .A1(P1_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n20592), .B1(
        n20591), .B2(n20572), .ZN(n20573) );
  OAI211_X1 U23506 ( .C1(n20575), .C2(n20595), .A(n20574), .B(n20573), .ZN(
        P1_U3157) );
  AOI22_X1 U23507 ( .A1(n20577), .A2(n20586), .B1(n20576), .B2(n20588), .ZN(
        n20580) );
  AOI22_X1 U23508 ( .A1(P1_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n20592), .B1(
        n20591), .B2(n20578), .ZN(n20579) );
  OAI211_X1 U23509 ( .C1(n20581), .C2(n20595), .A(n20580), .B(n20579), .ZN(
        P1_U3158) );
  AOI22_X1 U23510 ( .A1(n20928), .A2(n20586), .B1(n20926), .B2(n20588), .ZN(
        n20584) );
  AOI22_X1 U23511 ( .A1(P1_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n20592), .B1(
        n20591), .B2(n20582), .ZN(n20583) );
  OAI211_X1 U23512 ( .C1(n20585), .C2(n20595), .A(n20584), .B(n20583), .ZN(
        P1_U3159) );
  AOI22_X1 U23513 ( .A1(n20589), .A2(n20588), .B1(n20587), .B2(n20586), .ZN(
        n20594) );
  AOI22_X1 U23514 ( .A1(P1_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n20592), .B1(
        n20591), .B2(n20590), .ZN(n20593) );
  OAI211_X1 U23515 ( .C1(n20596), .C2(n20595), .A(n20594), .B(n20593), .ZN(
        P1_U3160) );
  NOR2_X1 U23516 ( .A1(n20597), .A2(n13663), .ZN(n20600) );
  OAI21_X1 U23517 ( .B1(n20600), .B2(n20599), .A(n20598), .ZN(P1_U3163) );
  INV_X1 U23518 ( .A(n20680), .ZN(n20676) );
  AND2_X1 U23519 ( .A1(P1_DATAWIDTH_REG_31__SCAN_IN), .A2(n20676), .ZN(
        P1_U3164) );
  AND2_X1 U23520 ( .A1(P1_DATAWIDTH_REG_30__SCAN_IN), .A2(n20676), .ZN(
        P1_U3165) );
  AND2_X1 U23521 ( .A1(P1_DATAWIDTH_REG_29__SCAN_IN), .A2(n20676), .ZN(
        P1_U3166) );
  AND2_X1 U23522 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(n20676), .ZN(
        P1_U3167) );
  AND2_X1 U23523 ( .A1(P1_DATAWIDTH_REG_27__SCAN_IN), .A2(n20676), .ZN(
        P1_U3168) );
  AND2_X1 U23524 ( .A1(P1_DATAWIDTH_REG_26__SCAN_IN), .A2(n20676), .ZN(
        P1_U3169) );
  AND2_X1 U23525 ( .A1(P1_DATAWIDTH_REG_25__SCAN_IN), .A2(n20676), .ZN(
        P1_U3170) );
  AND2_X1 U23526 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(n20676), .ZN(
        P1_U3171) );
  AND2_X1 U23527 ( .A1(P1_DATAWIDTH_REG_23__SCAN_IN), .A2(n20676), .ZN(
        P1_U3172) );
  AND2_X1 U23528 ( .A1(P1_DATAWIDTH_REG_22__SCAN_IN), .A2(n20676), .ZN(
        P1_U3173) );
  AND2_X1 U23529 ( .A1(P1_DATAWIDTH_REG_21__SCAN_IN), .A2(n20676), .ZN(
        P1_U3174) );
  AND2_X1 U23530 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(n20676), .ZN(
        P1_U3175) );
  AND2_X1 U23531 ( .A1(P1_DATAWIDTH_REG_19__SCAN_IN), .A2(n20676), .ZN(
        P1_U3176) );
  AND2_X1 U23532 ( .A1(P1_DATAWIDTH_REG_18__SCAN_IN), .A2(n20676), .ZN(
        P1_U3177) );
  AND2_X1 U23533 ( .A1(P1_DATAWIDTH_REG_17__SCAN_IN), .A2(n20676), .ZN(
        P1_U3178) );
  AND2_X1 U23534 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(n20676), .ZN(
        P1_U3179) );
  AND2_X1 U23535 ( .A1(P1_DATAWIDTH_REG_15__SCAN_IN), .A2(n20676), .ZN(
        P1_U3180) );
  AND2_X1 U23536 ( .A1(P1_DATAWIDTH_REG_14__SCAN_IN), .A2(n20676), .ZN(
        P1_U3181) );
  AND2_X1 U23537 ( .A1(P1_DATAWIDTH_REG_13__SCAN_IN), .A2(n20676), .ZN(
        P1_U3182) );
  AND2_X1 U23538 ( .A1(P1_DATAWIDTH_REG_12__SCAN_IN), .A2(n20676), .ZN(
        P1_U3183) );
  AND2_X1 U23539 ( .A1(P1_DATAWIDTH_REG_11__SCAN_IN), .A2(n20676), .ZN(
        P1_U3184) );
  AND2_X1 U23540 ( .A1(P1_DATAWIDTH_REG_10__SCAN_IN), .A2(n20676), .ZN(
        P1_U3185) );
  AND2_X1 U23541 ( .A1(P1_DATAWIDTH_REG_9__SCAN_IN), .A2(n20676), .ZN(P1_U3186) );
  INV_X1 U23542 ( .A(P1_DATAWIDTH_REG_8__SCAN_IN), .ZN(n20793) );
  NOR2_X1 U23543 ( .A1(n20680), .A2(n20793), .ZN(P1_U3187) );
  AND2_X1 U23544 ( .A1(P1_DATAWIDTH_REG_7__SCAN_IN), .A2(n20676), .ZN(P1_U3188) );
  AND2_X1 U23545 ( .A1(P1_DATAWIDTH_REG_6__SCAN_IN), .A2(n20676), .ZN(P1_U3189) );
  AND2_X1 U23546 ( .A1(P1_DATAWIDTH_REG_5__SCAN_IN), .A2(n20676), .ZN(P1_U3190) );
  AND2_X1 U23547 ( .A1(P1_DATAWIDTH_REG_4__SCAN_IN), .A2(n20676), .ZN(P1_U3191) );
  AND2_X1 U23548 ( .A1(P1_DATAWIDTH_REG_3__SCAN_IN), .A2(n20676), .ZN(P1_U3192) );
  AND2_X1 U23549 ( .A1(P1_DATAWIDTH_REG_2__SCAN_IN), .A2(n20676), .ZN(P1_U3193) );
  AOI21_X1 U23550 ( .B1(P1_STATE_REG_1__SCAN_IN), .B2(n20607), .A(n20604), 
        .ZN(n20614) );
  NOR2_X1 U23551 ( .A1(n20602), .A2(n20601), .ZN(n20603) );
  AOI211_X1 U23552 ( .C1(NA), .C2(n20604), .A(n20603), .B(n20608), .ZN(n20605)
         );
  OAI22_X1 U23553 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n20614), .B1(n20733), 
        .B2(n20605), .ZN(P1_U3194) );
  AOI21_X1 U23554 ( .B1(n20607), .B2(n20612), .A(n20606), .ZN(n20616) );
  OAI211_X1 U23555 ( .C1(P1_STATE_REG_2__SCAN_IN), .C2(n20608), .A(
        P1_STATE_REG_0__SCAN_IN), .B(HOLD), .ZN(n20615) );
  NOR2_X1 U23556 ( .A1(n20609), .A2(n20617), .ZN(n20610) );
  AOI221_X1 U23557 ( .B1(P1_STATE_REG_2__SCAN_IN), .B2(n20612), .C1(n20611), 
        .C2(n20612), .A(n20610), .ZN(n20613) );
  OAI22_X1 U23558 ( .A1(n20616), .A2(n20615), .B1(n20614), .B2(n20613), .ZN(
        P1_U3196) );
  NAND2_X1 U23559 ( .A1(n20733), .A2(n20617), .ZN(n20662) );
  NAND2_X1 U23560 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n20733), .ZN(n20664) );
  OAI222_X1 U23561 ( .A1(n20662), .A2(n20824), .B1(n20618), .B2(n20733), .C1(
        n20707), .C2(n20664), .ZN(P1_U3197) );
  INV_X1 U23562 ( .A(P1_ADDRESS_REG_1__SCAN_IN), .ZN(n20803) );
  OAI222_X1 U23563 ( .A1(n20664), .A2(n20824), .B1(n20803), .B2(n20733), .C1(
        n20620), .C2(n20662), .ZN(P1_U3198) );
  INV_X1 U23564 ( .A(P1_ADDRESS_REG_2__SCAN_IN), .ZN(n20619) );
  OAI222_X1 U23565 ( .A1(n20664), .A2(n20620), .B1(n20619), .B2(n20733), .C1(
        n20621), .C2(n20662), .ZN(P1_U3199) );
  INV_X1 U23566 ( .A(P1_ADDRESS_REG_3__SCAN_IN), .ZN(n20622) );
  OAI222_X1 U23567 ( .A1(n20662), .A2(n20624), .B1(n20622), .B2(n20733), .C1(
        n20621), .C2(n20664), .ZN(P1_U3200) );
  INV_X1 U23568 ( .A(P1_ADDRESS_REG_4__SCAN_IN), .ZN(n20623) );
  OAI222_X1 U23569 ( .A1(n20664), .A2(n20624), .B1(n20623), .B2(n20733), .C1(
        n20626), .C2(n20662), .ZN(P1_U3201) );
  INV_X1 U23570 ( .A(P1_ADDRESS_REG_5__SCAN_IN), .ZN(n20625) );
  OAI222_X1 U23571 ( .A1(n20664), .A2(n20626), .B1(n20625), .B2(n20733), .C1(
        n20629), .C2(n20662), .ZN(P1_U3202) );
  INV_X1 U23572 ( .A(P1_ADDRESS_REG_6__SCAN_IN), .ZN(n20628) );
  OAI222_X1 U23573 ( .A1(n20664), .A2(n20629), .B1(n20628), .B2(n20733), .C1(
        n20627), .C2(n20662), .ZN(P1_U3203) );
  INV_X1 U23574 ( .A(n20662), .ZN(n20666) );
  INV_X1 U23575 ( .A(n20664), .ZN(n20667) );
  AOI222_X1 U23576 ( .A1(n20666), .A2(P1_REIP_REG_9__SCAN_IN), .B1(
        P1_ADDRESS_REG_7__SCAN_IN), .B2(n20715), .C1(P1_REIP_REG_8__SCAN_IN), 
        .C2(n20667), .ZN(n20630) );
  INV_X1 U23577 ( .A(n20630), .ZN(P1_U3204) );
  AOI222_X1 U23578 ( .A1(n20667), .A2(P1_REIP_REG_9__SCAN_IN), .B1(
        P1_ADDRESS_REG_8__SCAN_IN), .B2(n20715), .C1(P1_REIP_REG_10__SCAN_IN), 
        .C2(n20666), .ZN(n20631) );
  INV_X1 U23579 ( .A(n20631), .ZN(P1_U3205) );
  INV_X1 U23580 ( .A(P1_ADDRESS_REG_9__SCAN_IN), .ZN(n20632) );
  OAI222_X1 U23581 ( .A1(n20664), .A2(n20633), .B1(n20632), .B2(n20733), .C1(
        n20635), .C2(n20662), .ZN(P1_U3206) );
  AOI22_X1 U23582 ( .A1(P1_ADDRESS_REG_10__SCAN_IN), .A2(n20715), .B1(
        P1_REIP_REG_12__SCAN_IN), .B2(n20666), .ZN(n20634) );
  OAI21_X1 U23583 ( .B1(n20635), .B2(n20664), .A(n20634), .ZN(P1_U3207) );
  AOI22_X1 U23584 ( .A1(P1_ADDRESS_REG_11__SCAN_IN), .A2(n20715), .B1(
        P1_REIP_REG_12__SCAN_IN), .B2(n20667), .ZN(n20636) );
  OAI21_X1 U23585 ( .B1(n20639), .B2(n20662), .A(n20636), .ZN(P1_U3208) );
  INV_X1 U23586 ( .A(P1_ADDRESS_REG_12__SCAN_IN), .ZN(n20638) );
  OAI222_X1 U23587 ( .A1(n20664), .A2(n20639), .B1(n20638), .B2(n20733), .C1(
        n20637), .C2(n20662), .ZN(P1_U3209) );
  AOI222_X1 U23588 ( .A1(n20666), .A2(P1_REIP_REG_15__SCAN_IN), .B1(
        P1_ADDRESS_REG_13__SCAN_IN), .B2(n20715), .C1(P1_REIP_REG_14__SCAN_IN), 
        .C2(n20667), .ZN(n20640) );
  INV_X1 U23589 ( .A(n20640), .ZN(P1_U3210) );
  AOI222_X1 U23590 ( .A1(n20667), .A2(P1_REIP_REG_15__SCAN_IN), .B1(
        P1_ADDRESS_REG_14__SCAN_IN), .B2(n20715), .C1(P1_REIP_REG_16__SCAN_IN), 
        .C2(n20666), .ZN(n20641) );
  INV_X1 U23591 ( .A(n20641), .ZN(P1_U3211) );
  INV_X1 U23592 ( .A(P1_ADDRESS_REG_15__SCAN_IN), .ZN(n20642) );
  INV_X1 U23593 ( .A(P1_REIP_REG_17__SCAN_IN), .ZN(n20821) );
  OAI222_X1 U23594 ( .A1(n20664), .A2(n20643), .B1(n20642), .B2(n20733), .C1(
        n20821), .C2(n20662), .ZN(P1_U3212) );
  INV_X1 U23595 ( .A(P1_ADDRESS_REG_16__SCAN_IN), .ZN(n20644) );
  OAI222_X1 U23596 ( .A1(n20662), .A2(n20646), .B1(n20644), .B2(n20733), .C1(
        n20821), .C2(n20664), .ZN(P1_U3213) );
  AOI22_X1 U23597 ( .A1(P1_ADDRESS_REG_17__SCAN_IN), .A2(n20715), .B1(
        P1_REIP_REG_19__SCAN_IN), .B2(n20666), .ZN(n20645) );
  OAI21_X1 U23598 ( .B1(n20646), .B2(n20664), .A(n20645), .ZN(P1_U3214) );
  INV_X1 U23599 ( .A(P1_REIP_REG_20__SCAN_IN), .ZN(n20649) );
  AOI22_X1 U23600 ( .A1(P1_ADDRESS_REG_18__SCAN_IN), .A2(n20715), .B1(
        P1_REIP_REG_19__SCAN_IN), .B2(n20667), .ZN(n20647) );
  OAI21_X1 U23601 ( .B1(n20649), .B2(n20662), .A(n20647), .ZN(P1_U3215) );
  INV_X1 U23602 ( .A(P1_ADDRESS_REG_19__SCAN_IN), .ZN(n20648) );
  OAI222_X1 U23603 ( .A1(n20664), .A2(n20649), .B1(n20648), .B2(n20733), .C1(
        n20650), .C2(n20662), .ZN(P1_U3216) );
  INV_X1 U23604 ( .A(P1_ADDRESS_REG_20__SCAN_IN), .ZN(n20651) );
  OAI222_X1 U23605 ( .A1(n20662), .A2(n20653), .B1(n20651), .B2(n20733), .C1(
        n20650), .C2(n20664), .ZN(P1_U3217) );
  AOI22_X1 U23606 ( .A1(P1_ADDRESS_REG_21__SCAN_IN), .A2(n20715), .B1(
        P1_REIP_REG_23__SCAN_IN), .B2(n20666), .ZN(n20652) );
  OAI21_X1 U23607 ( .B1(n20653), .B2(n20664), .A(n20652), .ZN(P1_U3218) );
  AOI22_X1 U23608 ( .A1(P1_ADDRESS_REG_22__SCAN_IN), .A2(n20715), .B1(
        P1_REIP_REG_23__SCAN_IN), .B2(n20667), .ZN(n20654) );
  OAI21_X1 U23609 ( .B1(n20656), .B2(n20662), .A(n20654), .ZN(P1_U3219) );
  INV_X1 U23610 ( .A(P1_ADDRESS_REG_23__SCAN_IN), .ZN(n20655) );
  OAI222_X1 U23611 ( .A1(n20664), .A2(n20656), .B1(n20655), .B2(n20733), .C1(
        n20657), .C2(n20662), .ZN(P1_U3220) );
  INV_X1 U23612 ( .A(P1_ADDRESS_REG_24__SCAN_IN), .ZN(n20658) );
  OAI222_X1 U23613 ( .A1(n20662), .A2(n20660), .B1(n20658), .B2(n20733), .C1(
        n20657), .C2(n20664), .ZN(P1_U3221) );
  AOI22_X1 U23614 ( .A1(P1_REIP_REG_27__SCAN_IN), .A2(n20666), .B1(
        P1_ADDRESS_REG_25__SCAN_IN), .B2(n20715), .ZN(n20659) );
  OAI21_X1 U23615 ( .B1(n20660), .B2(n20664), .A(n20659), .ZN(P1_U3222) );
  AOI22_X1 U23616 ( .A1(P1_REIP_REG_27__SCAN_IN), .A2(n20667), .B1(
        P1_ADDRESS_REG_26__SCAN_IN), .B2(n20715), .ZN(n20661) );
  OAI21_X1 U23617 ( .B1(n15455), .B2(n20662), .A(n20661), .ZN(P1_U3223) );
  INV_X1 U23618 ( .A(P1_ADDRESS_REG_27__SCAN_IN), .ZN(n20663) );
  OAI222_X1 U23619 ( .A1(n20664), .A2(n15455), .B1(n20663), .B2(n20733), .C1(
        n14217), .C2(n20662), .ZN(P1_U3224) );
  AOI222_X1 U23620 ( .A1(n20666), .A2(P1_REIP_REG_30__SCAN_IN), .B1(
        P1_ADDRESS_REG_28__SCAN_IN), .B2(n20715), .C1(P1_REIP_REG_29__SCAN_IN), 
        .C2(n20667), .ZN(n20665) );
  INV_X1 U23621 ( .A(n20665), .ZN(P1_U3225) );
  AOI222_X1 U23622 ( .A1(n20667), .A2(P1_REIP_REG_30__SCAN_IN), .B1(
        P1_ADDRESS_REG_29__SCAN_IN), .B2(n20715), .C1(P1_REIP_REG_31__SCAN_IN), 
        .C2(n20666), .ZN(n20668) );
  INV_X1 U23623 ( .A(n20668), .ZN(P1_U3226) );
  INV_X1 U23624 ( .A(P1_BE_N_REG_3__SCAN_IN), .ZN(n20669) );
  AOI22_X1 U23625 ( .A1(n20733), .A2(n20670), .B1(n20669), .B2(n20715), .ZN(
        P1_U3458) );
  INV_X1 U23626 ( .A(P1_BYTEENABLE_REG_2__SCAN_IN), .ZN(n20710) );
  INV_X1 U23627 ( .A(P1_BE_N_REG_2__SCAN_IN), .ZN(n20671) );
  AOI22_X1 U23628 ( .A1(n20733), .A2(n20710), .B1(n20671), .B2(n20715), .ZN(
        P1_U3459) );
  INV_X1 U23629 ( .A(P1_BE_N_REG_1__SCAN_IN), .ZN(n20672) );
  AOI22_X1 U23630 ( .A1(n20733), .A2(n20673), .B1(n20672), .B2(n20715), .ZN(
        P1_U3460) );
  INV_X1 U23631 ( .A(P1_BYTEENABLE_REG_0__SCAN_IN), .ZN(n20713) );
  INV_X1 U23632 ( .A(P1_BE_N_REG_0__SCAN_IN), .ZN(n20674) );
  AOI22_X1 U23633 ( .A1(n20733), .A2(n20713), .B1(n20674), .B2(n20715), .ZN(
        P1_U3461) );
  INV_X1 U23634 ( .A(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(n20677) );
  INV_X1 U23635 ( .A(n20678), .ZN(n20675) );
  AOI21_X1 U23636 ( .B1(n20677), .B2(n20676), .A(n20675), .ZN(P1_U3464) );
  OAI21_X1 U23637 ( .B1(n20680), .B2(n20679), .A(n20678), .ZN(P1_U3465) );
  OAI211_X1 U23638 ( .C1(P1_STATEBS16_REG_SCAN_IN), .C2(n20683), .A(n20682), 
        .B(n20681), .ZN(n20685) );
  AOI22_X1 U23639 ( .A1(n20685), .A2(n20700), .B1(n20698), .B2(n20684), .ZN(
        n20686) );
  INV_X1 U23640 ( .A(n20686), .ZN(n20688) );
  OAI21_X1 U23641 ( .B1(n20688), .B2(n20687), .A(n20702), .ZN(n20689) );
  OAI21_X1 U23642 ( .B1(n20702), .B2(n20690), .A(n20689), .ZN(P1_U3475) );
  NAND2_X1 U23643 ( .A1(n20700), .A2(n20691), .ZN(n20692) );
  AOI21_X1 U23644 ( .B1(n20693), .B2(n20891), .A(n20692), .ZN(n20694) );
  AOI21_X1 U23645 ( .B1(n20698), .B2(n20695), .A(n20694), .ZN(n20696) );
  AOI22_X1 U23646 ( .A1(n20706), .A2(n20697), .B1(n20696), .B2(n20702), .ZN(
        P1_U3477) );
  AOI22_X1 U23647 ( .A1(n20701), .A2(n20700), .B1(n20699), .B2(n20698), .ZN(
        n20705) );
  OAI222_X1 U23648 ( .A1(n20706), .A2(n20705), .B1(n20706), .B2(n20704), .C1(
        n20703), .C2(n20702), .ZN(P1_U3478) );
  AOI21_X1 U23649 ( .B1(P1_REIP_REG_0__SCAN_IN), .B2(
        P1_DATAWIDTH_REG_0__SCAN_IN), .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(
        n20708) );
  AOI22_X1 U23650 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_REIP_REG_0__SCAN_IN), 
        .B1(n20708), .B2(n20707), .ZN(n20711) );
  AOI22_X1 U23651 ( .A1(n20714), .A2(n20711), .B1(n20710), .B2(n20709), .ZN(
        P1_U3481) );
  OAI21_X1 U23652 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(P1_REIP_REG_0__SCAN_IN), 
        .A(n20714), .ZN(n20712) );
  OAI21_X1 U23653 ( .B1(n20714), .B2(n20713), .A(n20712), .ZN(P1_U3482) );
  AOI22_X1 U23654 ( .A1(n20733), .A2(P1_READREQUEST_REG_SCAN_IN), .B1(n20716), 
        .B2(n20715), .ZN(P1_U3483) );
  INV_X1 U23655 ( .A(n20717), .ZN(n20720) );
  AOI22_X1 U23656 ( .A1(n20721), .A2(n20720), .B1(n20719), .B2(n20718), .ZN(
        P1_U3484) );
  OAI21_X1 U23657 ( .B1(n20722), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n20724) );
  OAI22_X1 U23658 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n20725), .B1(n20724), 
        .B2(n20723), .ZN(n20732) );
  AOI211_X1 U23659 ( .C1(n20729), .C2(n20728), .A(n20727), .B(n20726), .ZN(
        n20731) );
  NAND2_X1 U23660 ( .A1(n20731), .A2(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(
        n20730) );
  OAI21_X1 U23661 ( .B1(n20732), .B2(n20731), .A(n20730), .ZN(P1_U3485) );
  MUX2_X1 U23662 ( .A(P1_M_IO_N_REG_SCAN_IN), .B(P1_MEMORYFETCH_REG_SCAN_IN), 
        .S(n20733), .Z(P1_U3486) );
  INV_X1 U23663 ( .A(P3_DATAO_REG_4__SCAN_IN), .ZN(n20818) );
  OAI22_X1 U23664 ( .A1(n14388), .A2(keyinput24), .B1(n20818), .B2(keyinput51), 
        .ZN(n20734) );
  AOI221_X1 U23665 ( .B1(n14388), .B2(keyinput24), .C1(keyinput51), .C2(n20818), .A(n20734), .ZN(n20743) );
  OAI22_X1 U23666 ( .A1(n20837), .A2(keyinput45), .B1(n20823), .B2(keyinput22), 
        .ZN(n20735) );
  AOI221_X1 U23667 ( .B1(n20837), .B2(keyinput45), .C1(keyinput22), .C2(n20823), .A(n20735), .ZN(n20742) );
  OAI22_X1 U23668 ( .A1(n20870), .A2(keyinput41), .B1(n20737), .B2(keyinput18), 
        .ZN(n20736) );
  AOI221_X1 U23669 ( .B1(n20870), .B2(keyinput41), .C1(keyinput18), .C2(n20737), .A(n20736), .ZN(n20741) );
  OAI22_X1 U23670 ( .A1(n20739), .A2(keyinput37), .B1(n20807), .B2(keyinput54), 
        .ZN(n20738) );
  AOI221_X1 U23671 ( .B1(n20739), .B2(keyinput37), .C1(keyinput54), .C2(n20807), .A(n20738), .ZN(n20740) );
  NAND4_X1 U23672 ( .A1(n20743), .A2(n20742), .A3(n20741), .A4(n20740), .ZN(
        n20924) );
  OAI22_X1 U23673 ( .A1(P2_INSTQUEUE_REG_15__7__SCAN_IN), .A2(keyinput31), 
        .B1(keyinput29), .B2(P1_ADDRESS_REG_1__SCAN_IN), .ZN(n20744) );
  AOI221_X1 U23674 ( .B1(P2_INSTQUEUE_REG_15__7__SCAN_IN), .B2(keyinput31), 
        .C1(P1_ADDRESS_REG_1__SCAN_IN), .C2(keyinput29), .A(n20744), .ZN(
        n20751) );
  OAI22_X1 U23675 ( .A1(P3_ADDRESS_REG_28__SCAN_IN), .A2(keyinput32), .B1(
        keyinput16), .B2(P2_DATAWIDTH_REG_15__SCAN_IN), .ZN(n20745) );
  AOI221_X1 U23676 ( .B1(P3_ADDRESS_REG_28__SCAN_IN), .B2(keyinput32), .C1(
        P2_DATAWIDTH_REG_15__SCAN_IN), .C2(keyinput16), .A(n20745), .ZN(n20750) );
  OAI22_X1 U23677 ( .A1(n20809), .A2(keyinput53), .B1(keyinput55), .B2(
        P3_REIP_REG_29__SCAN_IN), .ZN(n20746) );
  AOI221_X1 U23678 ( .B1(n20809), .B2(keyinput53), .C1(P3_REIP_REG_29__SCAN_IN), .C2(keyinput55), .A(n20746), .ZN(n20749) );
  OAI22_X1 U23679 ( .A1(P2_DATAWIDTH_REG_5__SCAN_IN), .A2(keyinput13), .B1(
        P2_BE_N_REG_0__SCAN_IN), .B2(keyinput9), .ZN(n20747) );
  AOI221_X1 U23680 ( .B1(P2_DATAWIDTH_REG_5__SCAN_IN), .B2(keyinput13), .C1(
        keyinput9), .C2(P2_BE_N_REG_0__SCAN_IN), .A(n20747), .ZN(n20748) );
  NAND4_X1 U23681 ( .A1(n20751), .A2(n20750), .A3(n20749), .A4(n20748), .ZN(
        n20923) );
  AOI22_X1 U23682 ( .A1(P2_LWORD_REG_2__SCAN_IN), .A2(keyinput3), .B1(
        P3_UWORD_REG_10__SCAN_IN), .B2(keyinput6), .ZN(n20752) );
  OAI221_X1 U23683 ( .B1(P2_LWORD_REG_2__SCAN_IN), .B2(keyinput3), .C1(
        P3_UWORD_REG_10__SCAN_IN), .C2(keyinput6), .A(n20752), .ZN(n20759) );
  AOI22_X1 U23684 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(keyinput1), .B1(
        P1_EBX_REG_31__SCAN_IN), .B2(keyinput40), .ZN(n20753) );
  OAI221_X1 U23685 ( .B1(P3_EBX_REG_14__SCAN_IN), .B2(keyinput1), .C1(
        P1_EBX_REG_31__SCAN_IN), .C2(keyinput40), .A(n20753), .ZN(n20758) );
  AOI22_X1 U23686 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(keyinput2), .B1(
        P2_INSTQUEUE_REG_8__7__SCAN_IN), .B2(keyinput7), .ZN(n20754) );
  OAI221_X1 U23687 ( .B1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .B2(keyinput2), .C1(
        P2_INSTQUEUE_REG_8__7__SCAN_IN), .C2(keyinput7), .A(n20754), .ZN(
        n20757) );
  AOI22_X1 U23688 ( .A1(P1_DATAWIDTH_REG_8__SCAN_IN), .A2(keyinput12), .B1(
        P3_INSTQUEUE_REG_15__6__SCAN_IN), .B2(keyinput39), .ZN(n20755) );
  OAI221_X1 U23689 ( .B1(P1_DATAWIDTH_REG_8__SCAN_IN), .B2(keyinput12), .C1(
        P3_INSTQUEUE_REG_15__6__SCAN_IN), .C2(keyinput39), .A(n20755), .ZN(
        n20756) );
  NOR4_X1 U23690 ( .A1(n20759), .A2(n20758), .A3(n20757), .A4(n20756), .ZN(
        n20787) );
  AOI22_X1 U23691 ( .A1(P3_INSTQUEUE_REG_3__3__SCAN_IN), .A2(keyinput21), .B1(
        P2_INSTQUEUE_REG_3__4__SCAN_IN), .B2(keyinput17), .ZN(n20760) );
  OAI221_X1 U23692 ( .B1(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B2(keyinput21), 
        .C1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .C2(keyinput17), .A(n20760), .ZN(
        n20767) );
  AOI22_X1 U23693 ( .A1(P1_REIP_REG_17__SCAN_IN), .A2(keyinput5), .B1(
        P2_EAX_REG_7__SCAN_IN), .B2(keyinput10), .ZN(n20761) );
  OAI221_X1 U23694 ( .B1(P1_REIP_REG_17__SCAN_IN), .B2(keyinput5), .C1(
        P2_EAX_REG_7__SCAN_IN), .C2(keyinput10), .A(n20761), .ZN(n20766) );
  AOI22_X1 U23695 ( .A1(P3_EAX_REG_19__SCAN_IN), .A2(keyinput48), .B1(
        P3_REIP_REG_17__SCAN_IN), .B2(keyinput25), .ZN(n20762) );
  OAI221_X1 U23696 ( .B1(P3_EAX_REG_19__SCAN_IN), .B2(keyinput48), .C1(
        P3_REIP_REG_17__SCAN_IN), .C2(keyinput25), .A(n20762), .ZN(n20765) );
  AOI22_X1 U23697 ( .A1(P2_DATAO_REG_25__SCAN_IN), .A2(keyinput44), .B1(
        P3_INSTQUEUE_REG_5__0__SCAN_IN), .B2(keyinput49), .ZN(n20763) );
  OAI221_X1 U23698 ( .B1(P2_DATAO_REG_25__SCAN_IN), .B2(keyinput44), .C1(
        P3_INSTQUEUE_REG_5__0__SCAN_IN), .C2(keyinput49), .A(n20763), .ZN(
        n20764) );
  NOR4_X1 U23699 ( .A1(n20767), .A2(n20766), .A3(n20765), .A4(n20764), .ZN(
        n20786) );
  AOI22_X1 U23700 ( .A1(BUF2_REG_9__SCAN_IN), .A2(keyinput28), .B1(
        P1_INSTQUEUE_REG_10__5__SCAN_IN), .B2(keyinput57), .ZN(n20768) );
  OAI221_X1 U23701 ( .B1(BUF2_REG_9__SCAN_IN), .B2(keyinput28), .C1(
        P1_INSTQUEUE_REG_10__5__SCAN_IN), .C2(keyinput57), .A(n20768), .ZN(
        n20775) );
  AOI22_X1 U23702 ( .A1(P2_UWORD_REG_10__SCAN_IN), .A2(keyinput33), .B1(
        P1_UWORD_REG_8__SCAN_IN), .B2(keyinput43), .ZN(n20769) );
  OAI221_X1 U23703 ( .B1(P2_UWORD_REG_10__SCAN_IN), .B2(keyinput33), .C1(
        P1_UWORD_REG_8__SCAN_IN), .C2(keyinput43), .A(n20769), .ZN(n20774) );
  AOI22_X1 U23704 ( .A1(P2_DATAO_REG_21__SCAN_IN), .A2(keyinput4), .B1(
        P1_ADDRESS_REG_12__SCAN_IN), .B2(keyinput61), .ZN(n20770) );
  OAI221_X1 U23705 ( .B1(P2_DATAO_REG_21__SCAN_IN), .B2(keyinput4), .C1(
        P1_ADDRESS_REG_12__SCAN_IN), .C2(keyinput61), .A(n20770), .ZN(n20773)
         );
  AOI22_X1 U23706 ( .A1(P2_UWORD_REG_14__SCAN_IN), .A2(keyinput20), .B1(
        P2_EAX_REG_28__SCAN_IN), .B2(keyinput23), .ZN(n20771) );
  OAI221_X1 U23707 ( .B1(P2_UWORD_REG_14__SCAN_IN), .B2(keyinput20), .C1(
        P2_EAX_REG_28__SCAN_IN), .C2(keyinput23), .A(n20771), .ZN(n20772) );
  NOR4_X1 U23708 ( .A1(n20775), .A2(n20774), .A3(n20773), .A4(n20772), .ZN(
        n20785) );
  AOI22_X1 U23709 ( .A1(BUF2_REG_3__SCAN_IN), .A2(keyinput42), .B1(
        P1_REIP_REG_3__SCAN_IN), .B2(keyinput38), .ZN(n20776) );
  OAI221_X1 U23710 ( .B1(BUF2_REG_3__SCAN_IN), .B2(keyinput42), .C1(
        P1_REIP_REG_3__SCAN_IN), .C2(keyinput38), .A(n20776), .ZN(n20783) );
  AOI22_X1 U23711 ( .A1(P3_DATAO_REG_8__SCAN_IN), .A2(keyinput14), .B1(
        P3_LWORD_REG_9__SCAN_IN), .B2(keyinput35), .ZN(n20777) );
  OAI221_X1 U23712 ( .B1(P3_DATAO_REG_8__SCAN_IN), .B2(keyinput14), .C1(
        P3_LWORD_REG_9__SCAN_IN), .C2(keyinput35), .A(n20777), .ZN(n20782) );
  AOI22_X1 U23713 ( .A1(P1_REIP_REG_2__SCAN_IN), .A2(keyinput36), .B1(
        P2_ADDRESS_REG_19__SCAN_IN), .B2(keyinput52), .ZN(n20778) );
  OAI221_X1 U23714 ( .B1(P1_REIP_REG_2__SCAN_IN), .B2(keyinput36), .C1(
        P2_ADDRESS_REG_19__SCAN_IN), .C2(keyinput52), .A(n20778), .ZN(n20781)
         );
  AOI22_X1 U23715 ( .A1(P3_UWORD_REG_1__SCAN_IN), .A2(keyinput59), .B1(
        P1_EAX_REG_0__SCAN_IN), .B2(keyinput62), .ZN(n20779) );
  OAI221_X1 U23716 ( .B1(P3_UWORD_REG_1__SCAN_IN), .B2(keyinput59), .C1(
        P1_EAX_REG_0__SCAN_IN), .C2(keyinput62), .A(n20779), .ZN(n20780) );
  NOR4_X1 U23717 ( .A1(n20783), .A2(n20782), .A3(n20781), .A4(n20780), .ZN(
        n20784) );
  NAND4_X1 U23718 ( .A1(n20787), .A2(n20786), .A3(n20785), .A4(n20784), .ZN(
        n20922) );
  AOI22_X1 U23719 ( .A1(n20892), .A2(keyinput94), .B1(n20789), .B2(keyinput74), 
        .ZN(n20788) );
  OAI221_X1 U23720 ( .B1(n20892), .B2(keyinput94), .C1(n20789), .C2(keyinput74), .A(n20788), .ZN(n20800) );
  INV_X1 U23721 ( .A(P3_DATAO_REG_8__SCAN_IN), .ZN(n20791) );
  AOI22_X1 U23722 ( .A1(n20791), .A2(keyinput78), .B1(n13109), .B2(keyinput92), 
        .ZN(n20790) );
  OAI221_X1 U23723 ( .B1(n20791), .B2(keyinput78), .C1(n13109), .C2(keyinput92), .A(n20790), .ZN(n20799) );
  AOI22_X1 U23724 ( .A1(n20794), .A2(keyinput104), .B1(keyinput76), .B2(n20793), .ZN(n20792) );
  OAI221_X1 U23725 ( .B1(n20794), .B2(keyinput104), .C1(n20793), .C2(
        keyinput76), .A(n20792), .ZN(n20798) );
  XOR2_X1 U23726 ( .A(n13254), .B(keyinput67), .Z(n20796) );
  XNOR2_X1 U23727 ( .A(P2_INSTQUEUE_REG_3__2__SCAN_IN), .B(keyinput90), .ZN(
        n20795) );
  NAND2_X1 U23728 ( .A1(n20796), .A2(n20795), .ZN(n20797) );
  NOR4_X1 U23729 ( .A1(n20800), .A2(n20799), .A3(n20798), .A4(n20797), .ZN(
        n20848) );
  AOI22_X1 U23730 ( .A1(n20803), .A2(keyinput93), .B1(keyinput108), .B2(n20802), .ZN(n20801) );
  OAI221_X1 U23731 ( .B1(n20803), .B2(keyinput93), .C1(n20802), .C2(
        keyinput108), .A(n20801), .ZN(n20813) );
  AOI22_X1 U23732 ( .A1(n20889), .A2(keyinput110), .B1(n14388), .B2(keyinput88), .ZN(n20804) );
  OAI221_X1 U23733 ( .B1(n20889), .B2(keyinput110), .C1(n14388), .C2(
        keyinput88), .A(n20804), .ZN(n20812) );
  AOI22_X1 U23734 ( .A1(n20807), .A2(keyinput118), .B1(keyinput97), .B2(n20806), .ZN(n20805) );
  OAI221_X1 U23735 ( .B1(n20807), .B2(keyinput118), .C1(n20806), .C2(
        keyinput97), .A(n20805), .ZN(n20811) );
  AOI22_X1 U23736 ( .A1(n20909), .A2(keyinput120), .B1(n20809), .B2(
        keyinput117), .ZN(n20808) );
  OAI221_X1 U23737 ( .B1(n20909), .B2(keyinput120), .C1(n20809), .C2(
        keyinput117), .A(n20808), .ZN(n20810) );
  NOR4_X1 U23738 ( .A1(n20813), .A2(n20812), .A3(n20811), .A4(n20810), .ZN(
        n20847) );
  AOI22_X1 U23739 ( .A1(n20816), .A2(keyinput68), .B1(n20815), .B2(keyinput85), 
        .ZN(n20814) );
  OAI221_X1 U23740 ( .B1(n20816), .B2(keyinput68), .C1(n20815), .C2(keyinput85), .A(n20814), .ZN(n20828) );
  INV_X1 U23741 ( .A(P3_EBX_REG_14__SCAN_IN), .ZN(n20819) );
  AOI22_X1 U23742 ( .A1(n20819), .A2(keyinput65), .B1(keyinput115), .B2(n20818), .ZN(n20817) );
  OAI221_X1 U23743 ( .B1(n20819), .B2(keyinput65), .C1(n20818), .C2(
        keyinput115), .A(n20817), .ZN(n20827) );
  AOI22_X1 U23744 ( .A1(n20894), .A2(keyinput79), .B1(keyinput69), .B2(n20821), 
        .ZN(n20820) );
  OAI221_X1 U23745 ( .B1(n20894), .B2(keyinput79), .C1(n20821), .C2(keyinput69), .A(n20820), .ZN(n20826) );
  AOI22_X1 U23746 ( .A1(n20824), .A2(keyinput100), .B1(keyinput86), .B2(n20823), .ZN(n20822) );
  OAI221_X1 U23747 ( .B1(n20824), .B2(keyinput100), .C1(n20823), .C2(
        keyinput86), .A(n20822), .ZN(n20825) );
  NOR4_X1 U23748 ( .A1(n20828), .A2(n20827), .A3(n20826), .A4(n20825), .ZN(
        n20846) );
  INV_X1 U23749 ( .A(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n20831) );
  AOI22_X1 U23750 ( .A1(n20831), .A2(keyinput121), .B1(keyinput113), .B2(
        n20830), .ZN(n20829) );
  OAI221_X1 U23751 ( .B1(n20831), .B2(keyinput121), .C1(n20830), .C2(
        keyinput113), .A(n20829), .ZN(n20844) );
  INV_X1 U23752 ( .A(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n20834) );
  AOI22_X1 U23753 ( .A1(n20834), .A2(keyinput81), .B1(keyinput112), .B2(n20833), .ZN(n20832) );
  OAI221_X1 U23754 ( .B1(n20834), .B2(keyinput81), .C1(n20833), .C2(
        keyinput112), .A(n20832), .ZN(n20843) );
  AOI22_X1 U23755 ( .A1(n20837), .A2(keyinput109), .B1(n20836), .B2(keyinput66), .ZN(n20835) );
  OAI221_X1 U23756 ( .B1(n20837), .B2(keyinput109), .C1(n20836), .C2(
        keyinput66), .A(n20835), .ZN(n20842) );
  AOI22_X1 U23757 ( .A1(n20840), .A2(keyinput119), .B1(n20839), .B2(keyinput87), .ZN(n20838) );
  OAI221_X1 U23758 ( .B1(n20840), .B2(keyinput119), .C1(n20839), .C2(
        keyinput87), .A(n20838), .ZN(n20841) );
  NOR4_X1 U23759 ( .A1(n20844), .A2(n20843), .A3(n20842), .A4(n20841), .ZN(
        n20845) );
  NAND4_X1 U23760 ( .A1(n20848), .A2(n20847), .A3(n20846), .A4(n20845), .ZN(
        n20920) );
  AOI22_X1 U23761 ( .A1(P3_UWORD_REG_11__SCAN_IN), .A2(keyinput127), .B1(
        BUF1_REG_3__SCAN_IN), .B2(keyinput122), .ZN(n20849) );
  OAI221_X1 U23762 ( .B1(P3_UWORD_REG_11__SCAN_IN), .B2(keyinput127), .C1(
        BUF1_REG_3__SCAN_IN), .C2(keyinput122), .A(n20849), .ZN(n20856) );
  AOI22_X1 U23763 ( .A1(P2_UWORD_REG_14__SCAN_IN), .A2(keyinput84), .B1(
        P2_INSTQUEUE_REG_15__7__SCAN_IN), .B2(keyinput95), .ZN(n20850) );
  OAI221_X1 U23764 ( .B1(P2_UWORD_REG_14__SCAN_IN), .B2(keyinput84), .C1(
        P2_INSTQUEUE_REG_15__7__SCAN_IN), .C2(keyinput95), .A(n20850), .ZN(
        n20855) );
  AOI22_X1 U23765 ( .A1(P3_UWORD_REG_1__SCAN_IN), .A2(keyinput123), .B1(
        P3_INSTQUEUE_REG_15__6__SCAN_IN), .B2(keyinput103), .ZN(n20851) );
  OAI221_X1 U23766 ( .B1(P3_UWORD_REG_1__SCAN_IN), .B2(keyinput123), .C1(
        P3_INSTQUEUE_REG_15__6__SCAN_IN), .C2(keyinput103), .A(n20851), .ZN(
        n20854) );
  AOI22_X1 U23767 ( .A1(P3_DATAWIDTH_REG_6__SCAN_IN), .A2(keyinput114), .B1(
        P2_PHYADDRPOINTER_REG_31__SCAN_IN), .B2(keyinput124), .ZN(n20852) );
  OAI221_X1 U23768 ( .B1(P3_DATAWIDTH_REG_6__SCAN_IN), .B2(keyinput114), .C1(
        P2_PHYADDRPOINTER_REG_31__SCAN_IN), .C2(keyinput124), .A(n20852), .ZN(
        n20853) );
  NOR4_X1 U23769 ( .A1(n20856), .A2(n20855), .A3(n20854), .A4(n20853), .ZN(
        n20887) );
  AOI22_X1 U23770 ( .A1(P1_UWORD_REG_3__SCAN_IN), .A2(keyinput91), .B1(
        P2_DATAWIDTH_REG_5__SCAN_IN), .B2(keyinput77), .ZN(n20857) );
  OAI221_X1 U23771 ( .B1(P1_UWORD_REG_3__SCAN_IN), .B2(keyinput91), .C1(
        P2_DATAWIDTH_REG_5__SCAN_IN), .C2(keyinput77), .A(n20857), .ZN(n20864)
         );
  AOI22_X1 U23772 ( .A1(P3_UWORD_REG_10__SCAN_IN), .A2(keyinput70), .B1(
        BUF2_REG_3__SCAN_IN), .B2(keyinput106), .ZN(n20858) );
  OAI221_X1 U23773 ( .B1(P3_UWORD_REG_10__SCAN_IN), .B2(keyinput70), .C1(
        BUF2_REG_3__SCAN_IN), .C2(keyinput106), .A(n20858), .ZN(n20863) );
  AOI22_X1 U23774 ( .A1(P1_REIP_REG_3__SCAN_IN), .A2(keyinput102), .B1(
        P2_ADDRESS_REG_19__SCAN_IN), .B2(keyinput116), .ZN(n20859) );
  OAI221_X1 U23775 ( .B1(P1_REIP_REG_3__SCAN_IN), .B2(keyinput102), .C1(
        P2_ADDRESS_REG_19__SCAN_IN), .C2(keyinput116), .A(n20859), .ZN(n20862)
         );
  AOI22_X1 U23776 ( .A1(P2_ADDRESS_REG_13__SCAN_IN), .A2(keyinput101), .B1(
        P2_INSTQUEUE_REG_8__7__SCAN_IN), .B2(keyinput71), .ZN(n20860) );
  OAI221_X1 U23777 ( .B1(P2_ADDRESS_REG_13__SCAN_IN), .B2(keyinput101), .C1(
        P2_INSTQUEUE_REG_8__7__SCAN_IN), .C2(keyinput71), .A(n20860), .ZN(
        n20861) );
  NOR4_X1 U23778 ( .A1(n20864), .A2(n20863), .A3(n20862), .A4(n20861), .ZN(
        n20886) );
  AOI22_X1 U23779 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(keyinput82), .B1(
        P3_ADDRESS_REG_28__SCAN_IN), .B2(keyinput96), .ZN(n20865) );
  OAI221_X1 U23780 ( .B1(P2_DATAWIDTH_REG_20__SCAN_IN), .B2(keyinput82), .C1(
        P3_ADDRESS_REG_28__SCAN_IN), .C2(keyinput96), .A(n20865), .ZN(n20875)
         );
  AOI22_X1 U23781 ( .A1(P3_LWORD_REG_9__SCAN_IN), .A2(keyinput99), .B1(
        P3_REIP_REG_17__SCAN_IN), .B2(keyinput89), .ZN(n20866) );
  OAI221_X1 U23782 ( .B1(P3_LWORD_REG_9__SCAN_IN), .B2(keyinput99), .C1(
        P3_REIP_REG_17__SCAN_IN), .C2(keyinput89), .A(n20866), .ZN(n20874) );
  AOI22_X1 U23783 ( .A1(n20868), .A2(keyinput80), .B1(n13751), .B2(keyinput72), 
        .ZN(n20867) );
  OAI221_X1 U23784 ( .B1(n20868), .B2(keyinput80), .C1(n13751), .C2(keyinput72), .A(n20867), .ZN(n20873) );
  AOI22_X1 U23785 ( .A1(n20871), .A2(keyinput107), .B1(n20870), .B2(
        keyinput105), .ZN(n20869) );
  OAI221_X1 U23786 ( .B1(n20871), .B2(keyinput107), .C1(n20870), .C2(
        keyinput105), .A(n20869), .ZN(n20872) );
  NOR4_X1 U23787 ( .A1(n20875), .A2(n20874), .A3(n20873), .A4(n20872), .ZN(
        n20885) );
  AOI22_X1 U23788 ( .A1(P1_DATAO_REG_5__SCAN_IN), .A2(keyinput98), .B1(
        P3_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(keyinput83), .ZN(n20876) );
  OAI221_X1 U23789 ( .B1(P1_DATAO_REG_5__SCAN_IN), .B2(keyinput98), .C1(
        P3_INSTADDRPOINTER_REG_6__SCAN_IN), .C2(keyinput83), .A(n20876), .ZN(
        n20883) );
  AOI22_X1 U23790 ( .A1(P2_BE_N_REG_0__SCAN_IN), .A2(keyinput73), .B1(
        P1_ADDRESS_REG_12__SCAN_IN), .B2(keyinput125), .ZN(n20877) );
  OAI221_X1 U23791 ( .B1(P2_BE_N_REG_0__SCAN_IN), .B2(keyinput73), .C1(
        P1_ADDRESS_REG_12__SCAN_IN), .C2(keyinput125), .A(n20877), .ZN(n20882)
         );
  AOI22_X1 U23792 ( .A1(P1_EAX_REG_0__SCAN_IN), .A2(keyinput126), .B1(
        P1_STATEBS16_REG_SCAN_IN), .B2(keyinput75), .ZN(n20878) );
  OAI221_X1 U23793 ( .B1(P1_EAX_REG_0__SCAN_IN), .B2(keyinput126), .C1(
        P1_STATEBS16_REG_SCAN_IN), .C2(keyinput75), .A(n20878), .ZN(n20881) );
  AOI22_X1 U23794 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(keyinput64), .B1(
        P2_INSTQUEUE_REG_10__6__SCAN_IN), .B2(keyinput111), .ZN(n20879) );
  OAI221_X1 U23795 ( .B1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B2(keyinput64), 
        .C1(P2_INSTQUEUE_REG_10__6__SCAN_IN), .C2(keyinput111), .A(n20879), 
        .ZN(n20880) );
  NOR4_X1 U23796 ( .A1(n20883), .A2(n20882), .A3(n20881), .A4(n20880), .ZN(
        n20884) );
  NAND4_X1 U23797 ( .A1(n20887), .A2(n20886), .A3(n20885), .A4(n20884), .ZN(
        n20919) );
  AOI22_X1 U23798 ( .A1(n20889), .A2(keyinput46), .B1(n11220), .B2(keyinput60), 
        .ZN(n20888) );
  OAI221_X1 U23799 ( .B1(n20889), .B2(keyinput46), .C1(n11220), .C2(keyinput60), .A(n20888), .ZN(n20901) );
  AOI22_X1 U23800 ( .A1(n20892), .A2(keyinput30), .B1(n20891), .B2(keyinput11), 
        .ZN(n20890) );
  OAI221_X1 U23801 ( .B1(n20892), .B2(keyinput30), .C1(n20891), .C2(keyinput11), .A(n20890), .ZN(n20900) );
  AOI22_X1 U23802 ( .A1(n20895), .A2(keyinput50), .B1(n20894), .B2(keyinput15), 
        .ZN(n20893) );
  OAI221_X1 U23803 ( .B1(n20895), .B2(keyinput50), .C1(n20894), .C2(keyinput15), .A(n20893), .ZN(n20899) );
  XOR2_X1 U23804 ( .A(n13751), .B(keyinput8), .Z(n20897) );
  XNOR2_X1 U23805 ( .A(P2_INSTQUEUE_REG_3__2__SCAN_IN), .B(keyinput26), .ZN(
        n20896) );
  NAND2_X1 U23806 ( .A1(n20897), .A2(n20896), .ZN(n20898) );
  NOR4_X1 U23807 ( .A1(n20901), .A2(n20900), .A3(n20899), .A4(n20898), .ZN(
        n20918) );
  AOI22_X1 U23808 ( .A1(n20903), .A2(keyinput27), .B1(n12180), .B2(keyinput47), 
        .ZN(n20902) );
  OAI221_X1 U23809 ( .B1(n20903), .B2(keyinput27), .C1(n12180), .C2(keyinput47), .A(n20902), .ZN(n20916) );
  INV_X1 U23810 ( .A(P3_UWORD_REG_11__SCAN_IN), .ZN(n20906) );
  AOI22_X1 U23811 ( .A1(n20906), .A2(keyinput63), .B1(keyinput34), .B2(n20905), 
        .ZN(n20904) );
  OAI221_X1 U23812 ( .B1(n20906), .B2(keyinput63), .C1(n20905), .C2(keyinput34), .A(n20904), .ZN(n20915) );
  AOI22_X1 U23813 ( .A1(n20909), .A2(keyinput56), .B1(n20908), .B2(keyinput0), 
        .ZN(n20907) );
  OAI221_X1 U23814 ( .B1(n20909), .B2(keyinput56), .C1(n20908), .C2(keyinput0), 
        .A(n20907), .ZN(n20914) );
  AOI22_X1 U23815 ( .A1(n20912), .A2(keyinput19), .B1(keyinput58), .B2(n20911), 
        .ZN(n20910) );
  OAI221_X1 U23816 ( .B1(n20912), .B2(keyinput19), .C1(n20911), .C2(keyinput58), .A(n20910), .ZN(n20913) );
  NOR4_X1 U23817 ( .A1(n20916), .A2(n20915), .A3(n20914), .A4(n20913), .ZN(
        n20917) );
  OAI211_X1 U23818 ( .C1(n20920), .C2(n20919), .A(n20918), .B(n20917), .ZN(
        n20921) );
  NOR4_X1 U23819 ( .A1(n20924), .A2(n20923), .A3(n20922), .A4(n20921), .ZN(
        n20937) );
  AOI22_X1 U23820 ( .A1(n20928), .A2(n20927), .B1(n20926), .B2(n20925), .ZN(
        n20933) );
  AOI22_X1 U23821 ( .A1(P1_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n20931), .B1(
        n20930), .B2(n20929), .ZN(n20932) );
  OAI211_X1 U23822 ( .C1(n20935), .C2(n20934), .A(n20933), .B(n20932), .ZN(
        n20936) );
  XOR2_X1 U23823 ( .A(n20937), .B(n20936), .Z(P1_U3047) );
  INV_X1 U16974 ( .A(n16777), .ZN(n16975) );
  OR2_X1 U13008 ( .A1(n10186), .A2(n10185), .ZN(n13489) );
  BUF_X2 U11414 ( .A(n13926), .Z(n9633) );
  INV_X1 U11052 ( .A(n10011), .ZN(n10006) );
  OR2_X1 U13814 ( .A1(n14322), .A2(n10962), .ZN(n14225) );
  CLKBUF_X1 U11059 ( .A(n10171), .Z(n11035) );
  CLKBUF_X3 U11094 ( .A(n10319), .Z(n9638) );
  NAND2_X1 U11135 ( .A1(n11442), .A2(n12376), .ZN(n12374) );
  CLKBUF_X1 U11141 ( .A(n11063), .Z(n11064) );
  CLKBUF_X1 U11181 ( .A(n11477), .Z(n11609) );
  AOI21_X1 U11198 ( .B1(n11497), .B2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(
        n11498), .ZN(n11501) );
  CLKBUF_X2 U11226 ( .A(n15172), .Z(n16825) );
  NAND2_X2 U11407 ( .A1(n13078), .A2(n9998), .ZN(n13082) );
  CLKBUF_X1 U11463 ( .A(n17701), .Z(n9648) );
  CLKBUF_X1 U11555 ( .A(n16332), .Z(n16331) );
endmodule

