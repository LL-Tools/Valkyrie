

module b15_C_gen_AntiSAT_k_128_8 ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, 
        READY_N, HOLD, READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, 
        CODEFETCH_REG_SCAN_IN, M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, 
        REQUESTPENDING_REG_SCAN_IN, STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, 
        FLUSH_REG_SCAN_IN, W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN, 
        BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN, 
        BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN, 
        REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN, 
        REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN, 
        REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN, 
        REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN, 
        REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN, 
        BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN, 
        ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN, 
        ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN, 
        ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN, 
        ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN, 
        ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN, 
        ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN, 
        ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN, 
        ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN, 
        ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN, 
        ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN, 
        ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN, ADDRESS_REG_7__SCAN_IN, 
        ADDRESS_REG_6__SCAN_IN, ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN, 
        ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN, ADDRESS_REG_1__SCAN_IN, 
        ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN, STATE_REG_1__SCAN_IN, 
        STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN, 
        DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN, 
        DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN, 
        DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN, 
        DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN, 
        DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN, 
        DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN, 
        DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN, 
        DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN, 
        DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN, 
        DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN, 
        DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN, 
        DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN, 
        DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN, 
        DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN, 
        DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN, 
        DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN, 
        STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN, 
        INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN, 
        INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN, 
        INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN, 
        INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN, 
        INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN, 
        INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN, 
        INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN, 
        INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN, 
        INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN, 
        INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN, 
        INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN, 
        INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN, 
        INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN, 
        INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN, 
        INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN, 
        INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN, 
        INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN, 
        INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN, 
        INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN, 
        INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN, 
        INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN, 
        INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN, 
        INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN, 
        INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN, 
        INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN, 
        INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN, 
        INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN, 
        INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN, 
        INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN, 
        INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN, 
        INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN, 
        INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN, 
        INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN, 
        INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN, 
        INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN, 
        INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN, 
        INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN, 
        INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN, 
        INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN, 
        INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN, 
        INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN, 
        INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN, 
        INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN, 
        INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN, 
        INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN, 
        INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN, 
        INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN, 
        INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN, 
        INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN, 
        INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN, 
        INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN, 
        INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN, 
        INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN, 
        INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN, 
        INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN, 
        INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN, 
        INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN, 
        INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN, 
        INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN, 
        INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN, 
        INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN, 
        INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN, 
        INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN, 
        INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN, 
        INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN, 
        INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN, 
        INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN, 
        INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN, 
        INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN, 
        INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN, 
        INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN, 
        INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN, 
        INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN, 
        INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN, 
        INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN, 
        INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN, 
        INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN, 
        INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN, 
        INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN, 
        INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN, 
        PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN, 
        PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN, 
        PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN, 
        PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN, 
        PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN, 
        PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN, 
        PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN, 
        PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN, 
        PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN, 
        PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN, 
        PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN, 
        PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN, 
        PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN, 
        PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN, 
        PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN, 
        PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN, 
        LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN, 
        LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN, 
        LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN, 
        LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN, 
        LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN, 
        LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN, 
        UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN, 
        UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN, 
        UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN, 
        UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN, 
        UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN, 
        EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN, 
        EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN, 
        EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN, 
        EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN, 
        EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN, 
        EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN, 
        EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN, 
        EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN, 
        EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN, 
        EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN, 
        EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN, 
        EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN, 
        EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN, 
        EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN, 
        EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN, 
        EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN, 
        EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN, 
        EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN, 
        EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN, 
        EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN, 
        EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN, 
        REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN, 
        REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN, 
        REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN, 
        REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN, 
        REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, keyinput_f0, keyinput_f1, 
        keyinput_f2, keyinput_f3, keyinput_f4, keyinput_f5, keyinput_f6, 
        keyinput_f7, keyinput_f8, keyinput_f9, keyinput_f10, keyinput_f11, 
        keyinput_f12, keyinput_f13, keyinput_f14, keyinput_f15, keyinput_f16, 
        keyinput_f17, keyinput_f18, keyinput_f19, keyinput_f20, keyinput_f21, 
        keyinput_f22, keyinput_f23, keyinput_f24, keyinput_f25, keyinput_f26, 
        keyinput_f27, keyinput_f28, keyinput_f29, keyinput_f30, keyinput_f31, 
        keyinput_f32, keyinput_f33, keyinput_f34, keyinput_f35, keyinput_f36, 
        keyinput_f37, keyinput_f38, keyinput_f39, keyinput_f40, keyinput_f41, 
        keyinput_f42, keyinput_f43, keyinput_f44, keyinput_f45, keyinput_f46, 
        keyinput_f47, keyinput_f48, keyinput_f49, keyinput_f50, keyinput_f51, 
        keyinput_f52, keyinput_f53, keyinput_f54, keyinput_f55, keyinput_f56, 
        keyinput_f57, keyinput_f58, keyinput_f59, keyinput_f60, keyinput_f61, 
        keyinput_f62, keyinput_f63, keyinput_g0, keyinput_g1, keyinput_g2, 
        keyinput_g3, keyinput_g4, keyinput_g5, keyinput_g6, keyinput_g7, 
        keyinput_g8, keyinput_g9, keyinput_g10, keyinput_g11, keyinput_g12, 
        keyinput_g13, keyinput_g14, keyinput_g15, keyinput_g16, keyinput_g17, 
        keyinput_g18, keyinput_g19, keyinput_g20, keyinput_g21, keyinput_g22, 
        keyinput_g23, keyinput_g24, keyinput_g25, keyinput_g26, keyinput_g27, 
        keyinput_g28, keyinput_g29, keyinput_g30, keyinput_g31, keyinput_g32, 
        keyinput_g33, keyinput_g34, keyinput_g35, keyinput_g36, keyinput_g37, 
        keyinput_g38, keyinput_g39, keyinput_g40, keyinput_g41, keyinput_g42, 
        keyinput_g43, keyinput_g44, keyinput_g45, keyinput_g46, keyinput_g47, 
        keyinput_g48, keyinput_g49, keyinput_g50, keyinput_g51, keyinput_g52, 
        keyinput_g53, keyinput_g54, keyinput_g55, keyinput_g56, keyinput_g57, 
        keyinput_g58, keyinput_g59, keyinput_g60, keyinput_g61, keyinput_g62, 
        keyinput_g63, U3445, U3446, U3447, U3448, U3213, U3212, U3211, U3210, 
        U3209, U3208, U3207, U3206, U3205, U3204, U3203, U3202, U3201, U3200, 
        U3199, U3198, U3197, U3196, U3195, U3194, U3193, U3192, U3191, U3190, 
        U3189, U3188, U3187, U3186, U3185, U3184, U3183, U3182, U3181, U3451, 
        U3452, U3180, U3179, U3178, U3177, U3176, U3175, U3174, U3173, U3172, 
        U3171, U3170, U3169, U3168, U3167, U3166, U3165, U3164, U3163, U3162, 
        U3161, U3160, U3159, U3158, U3157, U3156, U3155, U3154, U3153, U3152, 
        U3151, U3453, U3150, U3149, U3148, U3147, U3146, U3145, U3144, U3143, 
        U3142, U3141, U3140, U3139, U3138, U3137, U3136, U3135, U3134, U3133, 
        U3132, U3131, U3130, U3129, U3128, U3127, U3126, U3125, U3124, U3123, 
        U3122, U3121, U3120, U3119, U3118, U3117, U3116, U3115, U3114, U3113, 
        U3112, U3111, U3110, U3109, U3108, U3107, U3106, U3105, U3104, U3103, 
        U3102, U3101, U3100, U3099, U3098, U3097, U3096, U3095, U3094, U3093, 
        U3092, U3091, U3090, U3089, U3088, U3087, U3086, U3085, U3084, U3083, 
        U3082, U3081, U3080, U3079, U3078, U3077, U3076, U3075, U3074, U3073, 
        U3072, U3071, U3070, U3069, U3068, U3067, U3066, U3065, U3064, U3063, 
        U3062, U3061, U3060, U3059, U3058, U3057, U3056, U3055, U3054, U3053, 
        U3052, U3051, U3050, U3049, U3048, U3047, U3046, U3045, U3044, U3043, 
        U3042, U3041, U3040, U3039, U3038, U3037, U3036, U3035, U3034, U3033, 
        U3032, U3031, U3030, U3029, U3028, U3027, U3026, U3025, U3024, U3023, 
        U3022, U3021, U3020, U3455, U3456, U3459, U3460, U3461, U3019, U3462, 
        U3463, U3464, U3465, U3018, U3017, U3016, U3015, U3014, U3013, U3012, 
        U3011, U3010, U3009, U3008, U3007, U3006, U3005, U3004, U3003, U3002, 
        U3001, U3000, U2999, U2998, U2997, U2996, U2995, U2994, U2993, U2992, 
        U2991, U2990, U2989, U2988, U2987, U2986, U2985, U2984, U2983, U2982, 
        U2981, U2980, U2979, U2978, U2977, U2976, U2975, U2974, U2973, U2972, 
        U2971, U2970, U2969, U2968, U2967, U2966, U2965, U2964, U2963, U2962, 
        U2961, U2960, U2959, U2958, U2957, U2956, U2955, U2954, U2953, U2952, 
        U2951, U2950, U2949, U2948, U2947, U2946, U2945, U2944, U2943, U2942, 
        U2941, U2940, U2939, U2938, U2937, U2936, U2935, U2934, U2933, U2932, 
        U2931, U2930, U2929, U2928, U2927, U2926, U2925, U2924, U2923, U2922, 
        U2921, U2920, U2919, U2918, U2917, U2916, U2915, U2914, U2913, U2912, 
        U2911, U2910, U2909, U2908, U2907, U2906, U2905, U2904, U2903, U2902, 
        U2901, U2900, U2899, U2898, U2897, U2896, U2895, U2894, U2893, U2892, 
        U2891, U2890, U2889, U2888, U2887, U2886, U2885, U2884, U2883, U2882, 
        U2881, U2880, U2879, U2878, U2877, U2876, U2875, U2874, U2873, U2872, 
        U2871, U2870, U2869, U2868, U2867, U2866, U2865, U2864, U2863, U2862, 
        U2861, U2860, U2859, U2858, U2857, U2856, U2855, U2854, U2853, U2852, 
        U2851, U2850, U2849, U2848, U2847, U2846, U2845, U2844, U2843, U2842, 
        U2841, U2840, U2839, U2838, U2837, U2836, U2835, U2834, U2833, U2832, 
        U2831, U2830, U2829, U2828, U2827, U2826, U2825, U2824, U2823, U2822, 
        U2821, U2820, U2819, U2818, U2817, U2816, U2815, U2814, U2813, U2812, 
        U2811, U2810, U2809, U2808, U2807, U2806, U2805, U2804, U2803, U2802, 
        U2801, U2800, U2799, U2798, U2797, U2796, U2795, U3468, U2794, U3469, 
        U3470, U2793, U3471, U2792, U3472, U2791, U3473, U2790, U2789, U3474, 
        U2788 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, READY_N, HOLD,
         READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, CODEFETCH_REG_SCAN_IN,
         M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, REQUESTPENDING_REG_SCAN_IN,
         STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, FLUSH_REG_SCAN_IN,
         W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN,
         BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN,
         BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN,
         REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN,
         REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN,
         REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN,
         REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN,
         REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN,
         BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN,
         ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN,
         ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN,
         ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN,
         ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN,
         ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN,
         ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN,
         ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN,
         ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN,
         ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN,
         ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN,
         ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN,
         ADDRESS_REG_7__SCAN_IN, ADDRESS_REG_6__SCAN_IN,
         ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN,
         ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN,
         ADDRESS_REG_1__SCAN_IN, ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN,
         STATE_REG_1__SCAN_IN, STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN,
         DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN,
         DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN,
         DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN,
         DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN,
         DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN,
         DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN,
         DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN,
         DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN,
         DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN,
         DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN,
         DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN,
         DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN,
         DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN,
         DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN,
         DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN,
         DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN,
         STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN,
         INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN,
         INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN,
         INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN,
         INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN,
         INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN,
         INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN,
         INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN,
         INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN,
         INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN,
         INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN,
         INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN,
         INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN,
         INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN,
         INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN,
         INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN,
         INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN,
         INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN,
         INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN,
         INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN,
         INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN,
         INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN,
         INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN,
         INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN,
         INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN,
         INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN,
         INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN,
         INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN,
         INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN,
         INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN,
         INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN,
         INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN,
         INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN,
         INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN,
         INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN,
         INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN,
         INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN,
         INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN,
         INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN,
         INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN,
         INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN,
         INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN,
         INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN,
         INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN,
         INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN,
         INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN,
         INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN,
         INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN,
         INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN,
         INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN,
         INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN,
         INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN,
         INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN,
         INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN,
         INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN,
         INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN,
         INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN,
         INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN,
         INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN,
         INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN,
         INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN,
         INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN,
         INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN,
         INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN,
         INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN,
         INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN,
         INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN,
         INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN,
         INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN,
         INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN,
         INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN,
         INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN,
         INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN,
         INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN,
         INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN,
         INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN,
         INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN,
         INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN,
         INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN,
         INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN,
         INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN,
         PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN,
         PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN,
         PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN,
         PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN,
         PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN,
         PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN,
         PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN,
         PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN,
         PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN,
         PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN,
         PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN,
         PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN,
         PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN,
         PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN,
         PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN,
         PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN,
         LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN,
         LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN,
         LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN,
         LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN,
         LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN,
         LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN,
         UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN,
         UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN,
         UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN,
         UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN,
         UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN,
         DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN,
         DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN,
         DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN,
         DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN,
         DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN,
         DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN,
         DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN,
         DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN,
         DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN,
         DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN,
         EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN,
         EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN,
         EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN,
         EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN,
         EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN,
         EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN,
         EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN,
         EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN,
         EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN,
         EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN,
         EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN,
         EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN,
         EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN,
         EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN,
         EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN,
         EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN,
         EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN,
         EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN,
         EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN,
         EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN,
         EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN,
         EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN,
         REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN,
         REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN,
         REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN,
         REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN,
         REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, keyinput_f0, keyinput_f1,
         keyinput_f2, keyinput_f3, keyinput_f4, keyinput_f5, keyinput_f6,
         keyinput_f7, keyinput_f8, keyinput_f9, keyinput_f10, keyinput_f11,
         keyinput_f12, keyinput_f13, keyinput_f14, keyinput_f15, keyinput_f16,
         keyinput_f17, keyinput_f18, keyinput_f19, keyinput_f20, keyinput_f21,
         keyinput_f22, keyinput_f23, keyinput_f24, keyinput_f25, keyinput_f26,
         keyinput_f27, keyinput_f28, keyinput_f29, keyinput_f30, keyinput_f31,
         keyinput_f32, keyinput_f33, keyinput_f34, keyinput_f35, keyinput_f36,
         keyinput_f37, keyinput_f38, keyinput_f39, keyinput_f40, keyinput_f41,
         keyinput_f42, keyinput_f43, keyinput_f44, keyinput_f45, keyinput_f46,
         keyinput_f47, keyinput_f48, keyinput_f49, keyinput_f50, keyinput_f51,
         keyinput_f52, keyinput_f53, keyinput_f54, keyinput_f55, keyinput_f56,
         keyinput_f57, keyinput_f58, keyinput_f59, keyinput_f60, keyinput_f61,
         keyinput_f62, keyinput_f63, keyinput_g0, keyinput_g1, keyinput_g2,
         keyinput_g3, keyinput_g4, keyinput_g5, keyinput_g6, keyinput_g7,
         keyinput_g8, keyinput_g9, keyinput_g10, keyinput_g11, keyinput_g12,
         keyinput_g13, keyinput_g14, keyinput_g15, keyinput_g16, keyinput_g17,
         keyinput_g18, keyinput_g19, keyinput_g20, keyinput_g21, keyinput_g22,
         keyinput_g23, keyinput_g24, keyinput_g25, keyinput_g26, keyinput_g27,
         keyinput_g28, keyinput_g29, keyinput_g30, keyinput_g31, keyinput_g32,
         keyinput_g33, keyinput_g34, keyinput_g35, keyinput_g36, keyinput_g37,
         keyinput_g38, keyinput_g39, keyinput_g40, keyinput_g41, keyinput_g42,
         keyinput_g43, keyinput_g44, keyinput_g45, keyinput_g46, keyinput_g47,
         keyinput_g48, keyinput_g49, keyinput_g50, keyinput_g51, keyinput_g52,
         keyinput_g53, keyinput_g54, keyinput_g55, keyinput_g56, keyinput_g57,
         keyinput_g58, keyinput_g59, keyinput_g60, keyinput_g61, keyinput_g62,
         keyinput_g63;
  output U3445, U3446, U3447, U3448, U3213, U3212, U3211, U3210, U3209, U3208,
         U3207, U3206, U3205, U3204, U3203, U3202, U3201, U3200, U3199, U3198,
         U3197, U3196, U3195, U3194, U3193, U3192, U3191, U3190, U3189, U3188,
         U3187, U3186, U3185, U3184, U3183, U3182, U3181, U3451, U3452, U3180,
         U3179, U3178, U3177, U3176, U3175, U3174, U3173, U3172, U3171, U3170,
         U3169, U3168, U3167, U3166, U3165, U3164, U3163, U3162, U3161, U3160,
         U3159, U3158, U3157, U3156, U3155, U3154, U3153, U3152, U3151, U3453,
         U3150, U3149, U3148, U3147, U3146, U3145, U3144, U3143, U3142, U3141,
         U3140, U3139, U3138, U3137, U3136, U3135, U3134, U3133, U3132, U3131,
         U3130, U3129, U3128, U3127, U3126, U3125, U3124, U3123, U3122, U3121,
         U3120, U3119, U3118, U3117, U3116, U3115, U3114, U3113, U3112, U3111,
         U3110, U3109, U3108, U3107, U3106, U3105, U3104, U3103, U3102, U3101,
         U3100, U3099, U3098, U3097, U3096, U3095, U3094, U3093, U3092, U3091,
         U3090, U3089, U3088, U3087, U3086, U3085, U3084, U3083, U3082, U3081,
         U3080, U3079, U3078, U3077, U3076, U3075, U3074, U3073, U3072, U3071,
         U3070, U3069, U3068, U3067, U3066, U3065, U3064, U3063, U3062, U3061,
         U3060, U3059, U3058, U3057, U3056, U3055, U3054, U3053, U3052, U3051,
         U3050, U3049, U3048, U3047, U3046, U3045, U3044, U3043, U3042, U3041,
         U3040, U3039, U3038, U3037, U3036, U3035, U3034, U3033, U3032, U3031,
         U3030, U3029, U3028, U3027, U3026, U3025, U3024, U3023, U3022, U3021,
         U3020, U3455, U3456, U3459, U3460, U3461, U3019, U3462, U3463, U3464,
         U3465, U3018, U3017, U3016, U3015, U3014, U3013, U3012, U3011, U3010,
         U3009, U3008, U3007, U3006, U3005, U3004, U3003, U3002, U3001, U3000,
         U2999, U2998, U2997, U2996, U2995, U2994, U2993, U2992, U2991, U2990,
         U2989, U2988, U2987, U2986, U2985, U2984, U2983, U2982, U2981, U2980,
         U2979, U2978, U2977, U2976, U2975, U2974, U2973, U2972, U2971, U2970,
         U2969, U2968, U2967, U2966, U2965, U2964, U2963, U2962, U2961, U2960,
         U2959, U2958, U2957, U2956, U2955, U2954, U2953, U2952, U2951, U2950,
         U2949, U2948, U2947, U2946, U2945, U2944, U2943, U2942, U2941, U2940,
         U2939, U2938, U2937, U2936, U2935, U2934, U2933, U2932, U2931, U2930,
         U2929, U2928, U2927, U2926, U2925, U2924, U2923, U2922, U2921, U2920,
         U2919, U2918, U2917, U2916, U2915, U2914, U2913, U2912, U2911, U2910,
         U2909, U2908, U2907, U2906, U2905, U2904, U2903, U2902, U2901, U2900,
         U2899, U2898, U2897, U2896, U2895, U2894, U2893, U2892, U2891, U2890,
         U2889, U2888, U2887, U2886, U2885, U2884, U2883, U2882, U2881, U2880,
         U2879, U2878, U2877, U2876, U2875, U2874, U2873, U2872, U2871, U2870,
         U2869, U2868, U2867, U2866, U2865, U2864, U2863, U2862, U2861, U2860,
         U2859, U2858, U2857, U2856, U2855, U2854, U2853, U2852, U2851, U2850,
         U2849, U2848, U2847, U2846, U2845, U2844, U2843, U2842, U2841, U2840,
         U2839, U2838, U2837, U2836, U2835, U2834, U2833, U2832, U2831, U2830,
         U2829, U2828, U2827, U2826, U2825, U2824, U2823, U2822, U2821, U2820,
         U2819, U2818, U2817, U2816, U2815, U2814, U2813, U2812, U2811, U2810,
         U2809, U2808, U2807, U2806, U2805, U2804, U2803, U2802, U2801, U2800,
         U2799, U2798, U2797, U2796, U2795, U3468, U2794, U3469, U3470, U2793,
         U3471, U2792, U3472, U2791, U3473, U2790, U2789, U3474, U2788;
  wire   n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994,
         n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004,
         n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014,
         n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024,
         n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034,
         n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044,
         n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054,
         n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064,
         n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074,
         n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084,
         n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094,
         n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104,
         n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114,
         n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124,
         n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134,
         n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144,
         n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154,
         n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164,
         n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174,
         n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184,
         n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194,
         n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204,
         n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214,
         n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224,
         n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234,
         n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244,
         n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254,
         n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264,
         n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274,
         n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284,
         n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294,
         n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304,
         n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314,
         n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324,
         n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334,
         n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344,
         n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354,
         n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364,
         n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374,
         n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384,
         n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394,
         n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404,
         n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414,
         n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424,
         n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434,
         n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444,
         n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454,
         n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464,
         n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474,
         n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484,
         n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494,
         n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504,
         n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514,
         n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524,
         n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534,
         n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544,
         n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554,
         n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564,
         n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574,
         n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584,
         n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594,
         n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604,
         n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614,
         n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624,
         n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634,
         n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644,
         n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654,
         n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664,
         n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674,
         n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684,
         n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694,
         n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704,
         n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714,
         n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724,
         n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734,
         n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744,
         n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754,
         n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764,
         n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774,
         n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784,
         n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794,
         n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804,
         n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814,
         n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824,
         n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834,
         n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844,
         n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854,
         n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864,
         n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874,
         n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884,
         n3885, n3886, n3887, n3888, n3890, n3891, n3892, n3893, n3894, n3895,
         n3896, n3897, n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906,
         n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916,
         n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926,
         n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936,
         n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946,
         n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956,
         n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966,
         n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976,
         n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986,
         n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996,
         n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4007,
         n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017,
         n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027,
         n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037,
         n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047,
         n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057,
         n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067,
         n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077,
         n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087,
         n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097,
         n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107,
         n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117,
         n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127,
         n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137,
         n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147,
         n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157,
         n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167,
         n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177,
         n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187,
         n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197,
         n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207,
         n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217,
         n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227,
         n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237,
         n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247,
         n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257,
         n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267,
         n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277,
         n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287,
         n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297,
         n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307,
         n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317,
         n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327,
         n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337,
         n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347,
         n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357,
         n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367,
         n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377,
         n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387,
         n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397,
         n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407,
         n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417,
         n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427,
         n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437,
         n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447,
         n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457,
         n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467,
         n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477,
         n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487,
         n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497,
         n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507,
         n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517,
         n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527,
         n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537,
         n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547,
         n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557,
         n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567,
         n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577,
         n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587,
         n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597,
         n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607,
         n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617,
         n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627,
         n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637,
         n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647,
         n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657,
         n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667,
         n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677,
         n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687,
         n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697,
         n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707,
         n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717,
         n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727,
         n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737,
         n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747,
         n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757,
         n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767,
         n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777,
         n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787,
         n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797,
         n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807,
         n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817,
         n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827,
         n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837,
         n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847,
         n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857,
         n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867,
         n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877,
         n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887,
         n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897,
         n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907,
         n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917,
         n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927,
         n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937,
         n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947,
         n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957,
         n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967,
         n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977,
         n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987,
         n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997,
         n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007,
         n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017,
         n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027,
         n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037,
         n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047,
         n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057,
         n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067,
         n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077,
         n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087,
         n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097,
         n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107,
         n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117,
         n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127,
         n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137,
         n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147,
         n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157,
         n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167,
         n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177,
         n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187,
         n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197,
         n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207,
         n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217,
         n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227,
         n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237,
         n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247,
         n5248, n5249, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258,
         n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268,
         n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278,
         n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288,
         n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298,
         n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308,
         n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5317, n5318, n5319,
         n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329,
         n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339,
         n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349,
         n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359,
         n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369,
         n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379,
         n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389,
         n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399,
         n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409,
         n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419,
         n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429,
         n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439,
         n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449,
         n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459,
         n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469,
         n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479,
         n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489,
         n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499,
         n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509,
         n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519,
         n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529,
         n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539,
         n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549,
         n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559,
         n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569,
         n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579,
         n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589,
         n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599,
         n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609,
         n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619,
         n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629,
         n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639,
         n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649,
         n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659,
         n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669,
         n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679,
         n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689,
         n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699,
         n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709,
         n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719,
         n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729,
         n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739,
         n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749,
         n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759,
         n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769,
         n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779,
         n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789,
         n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799,
         n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809,
         n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819,
         n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829,
         n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839,
         n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849,
         n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859,
         n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869,
         n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879,
         n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889,
         n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899,
         n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909,
         n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919,
         n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929,
         n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939,
         n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949,
         n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959,
         n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969,
         n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979,
         n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989,
         n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999,
         n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009,
         n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019,
         n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029,
         n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039,
         n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049,
         n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059,
         n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069,
         n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079,
         n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089,
         n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099,
         n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109,
         n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119,
         n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129,
         n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139,
         n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149,
         n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159,
         n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169,
         n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179,
         n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189,
         n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199,
         n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209,
         n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219,
         n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229,
         n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239,
         n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249,
         n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259,
         n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269,
         n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279,
         n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289,
         n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299,
         n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309,
         n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319,
         n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329,
         n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339,
         n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349,
         n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359,
         n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369,
         n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379,
         n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389,
         n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399,
         n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409,
         n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419,
         n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429,
         n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439,
         n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449,
         n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459,
         n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469,
         n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479,
         n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489,
         n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499,
         n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509,
         n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519,
         n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529,
         n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539,
         n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549,
         n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559,
         n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569,
         n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579,
         n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589,
         n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599,
         n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609,
         n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619,
         n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629,
         n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639,
         n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649,
         n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659,
         n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669,
         n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679,
         n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689,
         n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699,
         n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709,
         n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719,
         n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729,
         n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739,
         n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749,
         n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759,
         n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769,
         n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779,
         n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789,
         n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799,
         n6800, n6801, n6802, n6803, n6804, n6805, n6806;

  BUF_X1 U3433 ( .A(n4288), .Z(n5615) );
  INV_X2 U3434 ( .A(n3437), .ZN(n5683) );
  OAI21_X1 U3435 ( .B1(n4861), .B2(n3425), .A(n3288), .ZN(n4352) );
  AND2_X1 U3436 ( .A1(n3895), .A2(n3894), .ZN(n4355) );
  INV_X2 U3437 ( .A(n3888), .ZN(n5374) );
  CLKBUF_X2 U3439 ( .A(n3191), .Z(n4063) );
  CLKBUF_X2 U3440 ( .A(n3106), .Z(n4116) );
  CLKBUF_X2 U3441 ( .A(n3608), .Z(n3853) );
  CLKBUF_X2 U3442 ( .A(n3231), .Z(n4125) );
  CLKBUF_X2 U3443 ( .A(n3253), .Z(n4117) );
  CLKBUF_X2 U3444 ( .A(n3225), .Z(n2994) );
  CLKBUF_X2 U34450 ( .A(n3190), .Z(n4021) );
  CLKBUF_X2 U34460 ( .A(n3107), .Z(n4022) );
  CLKBUF_X2 U34470 ( .A(n3197), .Z(n4027) );
  AND2_X1 U3449 ( .A1(n4513), .A2(n4518), .ZN(n3461) );
  CLKBUF_X1 U3450 ( .A(n3136), .Z(n4509) );
  INV_X2 U34510 ( .A(n4181), .ZN(n4513) );
  INV_X1 U34520 ( .A(n3144), .ZN(n3121) );
  OR2_X1 U34530 ( .A1(n3059), .A2(n3058), .ZN(n3164) );
  INV_X1 U3454 ( .A(n3133), .ZN(n4518) );
  INV_X1 U34560 ( .A(n3135), .ZN(n4493) );
  NAND4_X1 U3457 ( .A1(n3100), .A2(n3099), .A3(n3098), .A4(n3097), .ZN(n3133)
         );
  AND4_X1 U3458 ( .A1(n3018), .A2(n3017), .A3(n3016), .A4(n3015), .ZN(n3019)
         );
  AND2_X2 U34590 ( .A1(n3014), .A2(n4463), .ZN(n3832) );
  AND2_X2 U34600 ( .A1(n5839), .A2(n4430), .ZN(n3198) );
  AND2_X2 U34610 ( .A1(n5839), .A2(n3014), .ZN(n3106) );
  CLKBUF_X1 U34620 ( .A(n6572), .Z(n2985) );
  NOR2_X1 U34630 ( .A1(STATE_REG_2__SCAN_IN), .A2(n6803), .ZN(n6572) );
  NAND2_X1 U34640 ( .A1(n5186), .A2(n2989), .ZN(n2986) );
  AND2_X2 U34650 ( .A1(n2986), .A2(n2987), .ZN(n6213) );
  OR2_X1 U3466 ( .A1(n2988), .A2(n3435), .ZN(n2987) );
  INV_X1 U3467 ( .A(n5248), .ZN(n2988) );
  AND2_X1 U34680 ( .A1(n3434), .A2(n5248), .ZN(n2989) );
  AND2_X1 U34690 ( .A1(n3128), .A2(STATE2_REG_0__SCAN_IN), .ZN(n2990) );
  INV_X1 U34700 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n2991) );
  OAI211_X2 U34710 ( .C1(n4247), .C2(n3127), .A(n4236), .B(n4238), .ZN(n3128)
         );
  AOI21_X1 U34730 ( .B1(n3268), .B2(n3281), .A(n3424), .ZN(n3294) );
  NAND2_X1 U34740 ( .A1(n3990), .A2(n5562), .ZN(n4353) );
  AND2_X2 U3475 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4429) );
  INV_X1 U3476 ( .A(n5971), .ZN(n6036) );
  INV_X2 U3477 ( .A(n6335), .ZN(n2993) );
  NAND2_X2 U3478 ( .A1(n3285), .A2(n3284), .ZN(n4861) );
  INV_X1 U3479 ( .A(n5194), .ZN(n6071) );
  NAND2_X2 U3480 ( .A1(n3274), .A2(n3273), .ZN(n3362) );
  AND2_X1 U3482 ( .A1(n3709), .A2(n3697), .ZN(n5241) );
  CLKBUF_X1 U3483 ( .A(n3559), .Z(n5412) );
  NOR2_X1 U3484 ( .A1(n3263), .A2(n6498), .ZN(n3424) );
  BUF_X2 U3485 ( .A(n3162), .Z(n6130) );
  CLKBUF_X2 U3486 ( .A(n3912), .Z(n4380) );
  INV_X1 U3487 ( .A(n4182), .ZN(n3298) );
  CLKBUF_X2 U3488 ( .A(n3196), .Z(n4119) );
  AND2_X2 U3489 ( .A1(n4451), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n5839)
         );
  AOI211_X1 U3490 ( .C1(n6217), .C2(n5612), .A(n5611), .B(n5610), .ZN(n5613)
         );
  NOR2_X1 U3491 ( .A1(n4326), .A2(n4272), .ZN(n4275) );
  XNOR2_X1 U3492 ( .A(n4326), .B(n4148), .ZN(n5577) );
  CLKBUF_X1 U3493 ( .A(n4230), .Z(n5621) );
  CLKBUF_X1 U3494 ( .A(n5431), .Z(n5446) );
  CLKBUF_X1 U3495 ( .A(n5444), .Z(n5445) );
  CLKBUF_X1 U3496 ( .A(n5459), .Z(n5472) );
  CLKBUF_X1 U3497 ( .A(n4020), .Z(n5549) );
  CLKBUF_X1 U3498 ( .A(n5370), .Z(n5568) );
  CLKBUF_X1 U3499 ( .A(n5266), .Z(n5270) );
  CLKBUF_X1 U3500 ( .A(n5284), .Z(n5570) );
  CLKBUF_X1 U3501 ( .A(n5298), .Z(n5311) );
  AOI21_X1 U3502 ( .B1(n3607), .B2(n3733), .A(n3606), .ZN(n4851) );
  NAND2_X1 U3503 ( .A1(n3423), .A2(n3427), .ZN(n3437) );
  AOI21_X1 U3504 ( .B1(n3600), .B2(n3733), .A(n3599), .ZN(n4789) );
  NAND2_X1 U3505 ( .A1(n3569), .A2(n3692), .ZN(n4573) );
  OR2_X1 U3506 ( .A1(n4482), .A2(n3622), .ZN(n3569) );
  CLKBUF_X1 U3507 ( .A(n4482), .Z(n5831) );
  NOR2_X1 U3508 ( .A1(n5905), .A2(n5260), .ZN(n3945) );
  AND2_X2 U3509 ( .A1(n3332), .A2(n3331), .ZN(n4533) );
  CLKBUF_X1 U3510 ( .A(n4421), .Z(n4799) );
  NAND2_X1 U3511 ( .A1(n3206), .A2(n3205), .ZN(n3209) );
  NAND2_X1 U3512 ( .A1(n4421), .A2(n6498), .ZN(n3332) );
  XNOR2_X1 U3513 ( .A(n4465), .B(n4864), .ZN(n4421) );
  OR2_X1 U3514 ( .A1(n3312), .A2(n3311), .ZN(n4465) );
  NAND2_X1 U3515 ( .A1(n3224), .A2(n3223), .ZN(n3292) );
  NAND2_X1 U3516 ( .A1(n3920), .A2(n3003), .ZN(n4852) );
  CLKBUF_X1 U3517 ( .A(n4484), .Z(n6074) );
  CLKBUF_X1 U3518 ( .A(n3178), .Z(n2996) );
  OAI21_X1 U3519 ( .B1(n3180), .B2(n3153), .A(n3154), .ZN(n3246) );
  INV_X1 U3520 ( .A(n3262), .ZN(n3283) );
  AND2_X1 U3521 ( .A1(n3124), .A2(n3123), .ZN(n4002) );
  NAND2_X1 U3522 ( .A1(n3893), .A2(n3892), .ZN(n3896) );
  OAI21_X1 U3524 ( .B1(n3517), .B2(n3207), .A(n3143), .ZN(n3170) );
  INV_X1 U3525 ( .A(n3912), .ZN(n4012) );
  NAND2_X1 U3526 ( .A1(n3156), .A2(n4493), .ZN(n3517) );
  CLKBUF_X1 U3527 ( .A(n3156), .Z(n3157) );
  AND2_X1 U3528 ( .A1(n4513), .A2(n4360), .ZN(n3162) );
  NAND2_X1 U3529 ( .A1(n3156), .A2(n3136), .ZN(n3140) );
  CLKBUF_X1 U3530 ( .A(n3137), .Z(n3138) );
  NAND2_X1 U3532 ( .A1(n3029), .A2(n3028), .ZN(n3135) );
  AND4_X1 U3533 ( .A1(n3084), .A2(n3083), .A3(n3082), .A4(n3081), .ZN(n3100)
         );
  AND4_X1 U3534 ( .A1(n3096), .A2(n3095), .A3(n3094), .A4(n3093), .ZN(n3097)
         );
  AND4_X1 U3535 ( .A1(n3092), .A2(n3091), .A3(n3090), .A4(n3089), .ZN(n3098)
         );
  AND4_X1 U3536 ( .A1(n3037), .A2(n3036), .A3(n3035), .A4(n3034), .ZN(n3048)
         );
  AND4_X1 U3537 ( .A1(n3027), .A2(n3026), .A3(n3025), .A4(n3024), .ZN(n3028)
         );
  AND4_X1 U3538 ( .A1(n3033), .A2(n3032), .A3(n3031), .A4(n3030), .ZN(n3049)
         );
  AND4_X1 U3539 ( .A1(n3023), .A2(n3022), .A3(n3021), .A4(n3020), .ZN(n3029)
         );
  AND4_X1 U3540 ( .A1(n3088), .A2(n3087), .A3(n3086), .A4(n3085), .ZN(n3099)
         );
  AND4_X1 U3541 ( .A1(n3041), .A2(n3040), .A3(n3039), .A4(n3038), .ZN(n3047)
         );
  BUF_X2 U3542 ( .A(n3832), .Z(n4120) );
  BUF_X2 U3543 ( .A(n3198), .Z(n4126) );
  BUF_X2 U3544 ( .A(n3226), .Z(n4118) );
  AND2_X2 U3545 ( .A1(n3013), .A2(n5839), .ZN(n3608) );
  AND2_X2 U3546 ( .A1(n3013), .A2(n4463), .ZN(n3196) );
  AND2_X2 U3547 ( .A1(n4463), .A2(n4430), .ZN(n3107) );
  AND2_X2 U3548 ( .A1(n4463), .A2(n4420), .ZN(n3197) );
  INV_X1 U3549 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4451) );
  NAND2_X1 U3550 ( .A1(n3354), .A2(n3335), .ZN(n2995) );
  OAI211_X1 U3551 ( .C1(n3180), .C2(n2991), .A(n3151), .B(n3150), .ZN(n3178)
         );
  AND2_X1 U3552 ( .A1(n3157), .A2(n4181), .ZN(n3464) );
  AND2_X1 U3554 ( .A1(n4222), .A2(n3453), .ZN(n5665) );
  INV_X1 U3555 ( .A(n3115), .ZN(n3136) );
  AND2_X1 U3557 ( .A1(n4463), .A2(n4420), .ZN(n2997) );
  XNOR2_X2 U3558 ( .A(n3896), .B(n4355), .ZN(n6086) );
  NOR2_X2 U3559 ( .A1(n4230), .A2(n4228), .ZN(n4288) );
  NOR2_X2 U3560 ( .A1(n5596), .A2(n5622), .ZN(n4230) );
  NAND2_X1 U3561 ( .A1(n2990), .A2(n3001), .ZN(n3152) );
  NAND2_X1 U3562 ( .A1(n3246), .A2(n3245), .ZN(n3210) );
  NOR2_X1 U3563 ( .A1(n3170), .A2(n4182), .ZN(n4189) );
  NAND2_X1 U3564 ( .A1(n5511), .A2(n5512), .ZN(n4020) );
  XNOR2_X1 U3565 ( .A(n3423), .B(n3414), .ZN(n3607) );
  NOR2_X1 U3566 ( .A1(STATE2_REG_2__SCAN_IN), .A2(STATEBS16_REG_SCAN_IN), .ZN(
        n3811) );
  AND2_X1 U3567 ( .A1(n5321), .A2(n3446), .ZN(n5670) );
  AND2_X1 U3568 ( .A1(n3458), .A2(n3207), .ZN(n3499) );
  OR2_X1 U3569 ( .A1(n6595), .A2(n4260), .ZN(n6046) );
  INV_X1 U3570 ( .A(n6500), .ZN(n4394) );
  NAND2_X1 U3571 ( .A1(n4324), .A2(n4327), .ZN(n4326) );
  NOR2_X1 U3572 ( .A1(n5629), .A2(n4231), .ZN(n4289) );
  NOR2_X2 U3573 ( .A1(n4852), .A2(n4853), .ZN(n5026) );
  OR2_X1 U3574 ( .A1(n4244), .A2(n4428), .ZN(n5336) );
  NAND2_X1 U3575 ( .A1(n4335), .A2(n4336), .ZN(n6595) );
  INV_X1 U3576 ( .A(n3139), .ZN(n3127) );
  OR2_X1 U3577 ( .A1(n3397), .A2(n3396), .ZN(n3416) );
  AND2_X1 U3578 ( .A1(n3498), .A2(n3497), .ZN(n4160) );
  AND3_X1 U3579 ( .A1(n3174), .A2(n3173), .A3(n3172), .ZN(n3175) );
  NAND2_X1 U3580 ( .A1(n3796), .A2(n3795), .ZN(n5370) );
  INV_X1 U3581 ( .A(n5284), .ZN(n3796) );
  INV_X1 U3582 ( .A(n3409), .ZN(n3411) );
  NAND2_X1 U3583 ( .A1(n4012), .A2(n3988), .ZN(n3984) );
  AND3_X1 U3584 ( .A1(n3243), .A2(n3248), .A3(n3242), .ZN(n3291) );
  NAND2_X1 U3585 ( .A1(n4484), .A2(n6498), .ZN(n3224) );
  AND2_X1 U3586 ( .A1(n3506), .A2(n3505), .ZN(n4165) );
  OR2_X1 U3587 ( .A1(n3504), .A2(n3503), .ZN(n3506) );
  NAND2_X1 U3588 ( .A1(n3499), .A2(n3464), .ZN(n3511) );
  NAND2_X1 U3589 ( .A1(n3149), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3180) );
  AND2_X1 U3590 ( .A1(n3129), .A2(n3184), .ZN(n4866) );
  AOI22_X1 U3591 ( .A1(n3198), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n3226), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3024) );
  NOR2_X1 U3592 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n4492), .ZN(n4757) );
  OR2_X1 U3593 ( .A1(n4448), .A2(n4447), .ZN(n4469) );
  OR2_X1 U3594 ( .A1(n6126), .A2(n4248), .ZN(n4335) );
  OR3_X1 U3595 ( .A1(n6126), .A2(READY_N), .A3(n4441), .ZN(n6131) );
  CLKBUF_X1 U3596 ( .A(n4324), .Z(n4325) );
  NOR2_X2 U3597 ( .A1(n4020), .A2(n4019), .ZN(n5474) );
  OR2_X1 U3598 ( .A1(n4018), .A2(n5548), .ZN(n4019) );
  AND2_X1 U3599 ( .A1(PHYADDRPOINTER_REG_16__SCAN_IN), .A2(n3752), .ZN(n3772)
         );
  AND2_X1 U3600 ( .A1(n5215), .A2(n5214), .ZN(n5280) );
  OR2_X1 U3601 ( .A1(n5223), .A2(n5224), .ZN(n5278) );
  OR2_X1 U3602 ( .A1(n5213), .A2(n5212), .ZN(n5223) );
  NAND2_X1 U3603 ( .A1(n4475), .A2(n4394), .ZN(n6126) );
  INV_X1 U3604 ( .A(n5657), .ZN(n3454) );
  AND2_X1 U3605 ( .A1(n5674), .A2(n5345), .ZN(n3448) );
  NOR2_X1 U3606 ( .A1(n5629), .A2(n6254), .ZN(n5267) );
  AND2_X1 U3607 ( .A1(n6212), .A2(n3439), .ZN(n3440) );
  OR2_X1 U3608 ( .A1(n5629), .A2(n3928), .ZN(n6212) );
  OR2_X1 U3609 ( .A1(n3987), .A2(EBX_REG_6__SCAN_IN), .ZN(n3919) );
  AND2_X1 U3610 ( .A1(n3164), .A2(n3554), .ZN(n4398) );
  NAND2_X1 U3611 ( .A1(n4178), .A2(n4394), .ZN(n4244) );
  NOR2_X1 U3612 ( .A1(n5831), .A2(n3333), .ZN(n4668) );
  AND2_X1 U3613 ( .A1(n4313), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4314) );
  OR2_X1 U3614 ( .A1(n5193), .A2(n4252), .ZN(n6065) );
  INV_X1 U3615 ( .A(n5397), .ZN(n6102) );
  AND2_X1 U3616 ( .A1(n5397), .A2(n4398), .ZN(n6099) );
  AND2_X1 U3617 ( .A1(n5397), .A2(n4399), .ZN(n6103) );
  INV_X1 U3618 ( .A(n4272), .ZN(n4148) );
  OAI21_X1 U3619 ( .B1(n4325), .B2(n4327), .A(n4326), .ZN(n5420) );
  INV_X1 U3620 ( .A(n6249), .ZN(n6217) );
  INV_X1 U3621 ( .A(n5691), .ZN(n6239) );
  OR2_X1 U3622 ( .A1(n6508), .A2(n5835), .ZN(n5697) );
  XNOR2_X1 U3623 ( .A(n4292), .B(n4299), .ZN(n4323) );
  OR2_X1 U3624 ( .A1(n3283), .A2(n3282), .ZN(n3284) );
  AND2_X1 U3625 ( .A1(n3131), .A2(n3130), .ZN(n3150) );
  NAND2_X1 U3626 ( .A1(n3114), .A2(n4159), .ZN(n3139) );
  INV_X1 U3627 ( .A(n4181), .ZN(n3114) );
  AND2_X2 U3628 ( .A1(n3181), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3013)
         );
  OR2_X1 U3629 ( .A1(n4360), .A2(n6498), .ZN(n3318) );
  OR2_X1 U3630 ( .A1(n3207), .A2(n6498), .ZN(n3319) );
  NOR2_X1 U3631 ( .A1(n3362), .A2(n4533), .ZN(n3364) );
  NAND2_X1 U3632 ( .A1(n3387), .A2(n3386), .ZN(n3409) );
  INV_X1 U3633 ( .A(n3385), .ZN(n3387) );
  OR2_X1 U3634 ( .A1(n3374), .A2(n3373), .ZN(n3400) );
  INV_X1 U3635 ( .A(n3461), .ZN(n4240) );
  OR2_X1 U3636 ( .A1(n3517), .A2(n6599), .ZN(n4007) );
  AND2_X1 U3637 ( .A1(n4360), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3458) );
  INV_X1 U3638 ( .A(n3319), .ZN(n3240) );
  INV_X1 U3639 ( .A(n3291), .ZN(n3244) );
  NAND2_X1 U3640 ( .A1(n3121), .A2(n4518), .ZN(n3122) );
  NAND2_X1 U3641 ( .A1(n3189), .A2(n3188), .ZN(n3310) );
  OR2_X1 U3642 ( .A1(n3180), .A2(n3182), .ZN(n3189) );
  AOI22_X1 U3643 ( .A1(n3832), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n3197), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3105) );
  AOI22_X1 U3644 ( .A1(n3608), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3106), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3020) );
  AOI22_X1 U3645 ( .A1(n4127), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3324), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3026) );
  NAND2_X1 U3646 ( .A1(n3319), .A2(n3318), .ZN(n3507) );
  OR2_X2 U3647 ( .A1(n3080), .A2(n3079), .ZN(n4182) );
  NOR2_X1 U3648 ( .A1(n5459), .A2(n5460), .ZN(n5444) );
  NAND2_X1 U3649 ( .A1(n5474), .A2(n5473), .ZN(n5459) );
  NOR2_X1 U3650 ( .A1(n5842), .A2(n6498), .ZN(n4111) );
  INV_X1 U3651 ( .A(n4789), .ZN(n3601) );
  AND2_X1 U3652 ( .A1(n5629), .A2(n5750), .ZN(n4228) );
  NAND2_X1 U3653 ( .A1(n5476), .A2(n5475), .ZN(n5462) );
  NAND2_X1 U3654 ( .A1(n5319), .A2(n3443), .ZN(n3450) );
  AND2_X1 U3655 ( .A1(n5320), .A2(n3442), .ZN(n3443) );
  NOR2_X1 U3656 ( .A1(n5227), .A2(n5226), .ZN(n5225) );
  NAND2_X1 U3657 ( .A1(n3607), .A2(n3464), .ZN(n3420) );
  INV_X1 U3658 ( .A(n3897), .ZN(n3987) );
  NOR2_X1 U3659 ( .A1(n4182), .A2(n3156), .ZN(n3125) );
  INV_X1 U3660 ( .A(n3296), .ZN(n3264) );
  CLKBUF_X1 U3661 ( .A(n4002), .Z(n4003) );
  INV_X1 U3662 ( .A(n3210), .ZN(n3211) );
  AOI21_X1 U3663 ( .B1(n6507), .B2(n4478), .A(n5415), .ZN(n4492) );
  INV_X1 U3664 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6464) );
  INV_X1 U3665 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n6468) );
  CLKBUF_X1 U3666 ( .A(n4167), .Z(n4168) );
  INV_X1 U3667 ( .A(n3162), .ZN(n6599) );
  NOR2_X1 U3669 ( .A1(n3724), .A2(n5967), .ZN(n3752) );
  XNOR2_X1 U3670 ( .A(n3247), .B(n3246), .ZN(n3559) );
  AND2_X1 U3671 ( .A1(n3941), .A2(n3940), .ZN(n5903) );
  INV_X1 U3672 ( .A(n6125), .ZN(n4361) );
  NOR2_X1 U3673 ( .A1(n4041), .A2(n5623), .ZN(n4042) );
  NAND2_X1 U3674 ( .A1(n4042), .A2(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n4078)
         );
  OR2_X1 U3675 ( .A1(n4038), .A2(n5490), .ZN(n4041) );
  AND2_X1 U3676 ( .A1(n3848), .A2(n3847), .ZN(n5512) );
  AND2_X1 U3677 ( .A1(n3831), .A2(n3830), .ZN(n5557) );
  OR2_X1 U3678 ( .A1(n5866), .A2(n4139), .ZN(n3830) );
  CLKBUF_X1 U3679 ( .A(n5372), .Z(n5558) );
  NAND2_X1 U3680 ( .A1(n3772), .A2(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n3790)
         );
  AND2_X1 U3681 ( .A1(n3774), .A2(n3773), .ZN(n5285) );
  CLKBUF_X1 U3682 ( .A(n5282), .Z(n5283) );
  NAND2_X1 U3683 ( .A1(n5246), .A2(n3709), .ZN(n5258) );
  INV_X1 U3684 ( .A(n3689), .ZN(n3710) );
  AND2_X1 U3685 ( .A1(n3619), .A2(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n3690)
         );
  NAND2_X1 U3686 ( .A1(n3690), .A2(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n3689)
         );
  NAND2_X1 U3687 ( .A1(n5241), .A2(n5242), .ZN(n5246) );
  NAND2_X1 U3688 ( .A1(n3640), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n3624)
         );
  INV_X1 U3689 ( .A(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n6002) );
  NOR2_X1 U3690 ( .A1(n3655), .A2(n6011), .ZN(n3640) );
  CLKBUF_X1 U3691 ( .A(n4910), .Z(n4911) );
  NOR2_X1 U3692 ( .A1(n3591), .A2(n4846), .ZN(n3595) );
  AND2_X1 U3693 ( .A1(n3595), .A2(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n3603)
         );
  CLKBUF_X1 U3694 ( .A(n4788), .Z(n4850) );
  INV_X1 U3695 ( .A(n3563), .ZN(n3574) );
  AND2_X1 U3696 ( .A1(PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n3574), .ZN(n3585)
         );
  AOI21_X1 U3697 ( .B1(n4861), .B2(n4493), .A(n6497), .ZN(n4370) );
  OR2_X1 U3698 ( .A1(n5596), .A2(n5597), .ZN(n5605) );
  CLKBUF_X1 U3699 ( .A(n5504), .Z(n5505) );
  INV_X1 U3700 ( .A(n5376), .ZN(n3956) );
  NAND2_X1 U3701 ( .A1(n5629), .A2(n5799), .ZN(n3453) );
  AND2_X1 U3703 ( .A1(n5670), .A2(n3447), .ZN(n5345) );
  CLKBUF_X1 U3704 ( .A(n5301), .Z(n5314) );
  OR2_X1 U3705 ( .A1(n3445), .A2(n5892), .ZN(n5321) );
  OR2_X1 U3706 ( .A1(n4244), .A2(n4193), .ZN(n5326) );
  INV_X1 U3707 ( .A(n4588), .ZN(n3920) );
  NAND2_X1 U3708 ( .A1(n3903), .A2(n3902), .ZN(n4578) );
  INV_X1 U3709 ( .A(n4575), .ZN(n3902) );
  INV_X1 U3710 ( .A(n4576), .ZN(n3903) );
  NOR2_X2 U3711 ( .A1(n4578), .A2(n4529), .ZN(n4567) );
  CLKBUF_X1 U3712 ( .A(n4236), .Z(n4237) );
  NAND2_X1 U3713 ( .A1(n3559), .A2(n6498), .ZN(n3279) );
  XNOR2_X1 U3714 ( .A(n3292), .B(n3291), .ZN(n3293) );
  CLKBUF_X1 U3715 ( .A(n4449), .Z(n5833) );
  AND2_X2 U3716 ( .A1(n3007), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n5838)
         );
  INV_X1 U3717 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3007) );
  OR2_X1 U3718 ( .A1(n3517), .A2(n3516), .ZN(n5842) );
  INV_X1 U3719 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3181) );
  OR2_X1 U3720 ( .A1(n3510), .A2(n3509), .ZN(n3514) );
  INV_X1 U3721 ( .A(n4469), .ZN(n6459) );
  NOR2_X1 U3722 ( .A1(n4799), .A2(n5835), .ZN(n6348) );
  NOR2_X1 U3723 ( .A1(n2995), .A2(n4640), .ZN(n4620) );
  NOR2_X1 U3724 ( .A1(n2995), .A2(n4915), .ZN(n4601) );
  AND2_X1 U3725 ( .A1(n5833), .A2(n5829), .ZN(n5033) );
  NOR2_X1 U3726 ( .A1(n4532), .A2(n5827), .ZN(n4862) );
  INV_X1 U3727 ( .A(n4861), .ZN(n4711) );
  OR3_X1 U3728 ( .A1(n6581), .A2(STATE2_REG_0__SCAN_IN), .A3(n4492), .ZN(n4519) );
  INV_X1 U3729 ( .A(n4757), .ZN(n4867) );
  AND2_X1 U3730 ( .A1(n5413), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3515) );
  INV_X1 U3731 ( .A(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n6011) );
  AND2_X1 U3732 ( .A1(n4267), .A2(n4250), .ZN(n6047) );
  AND2_X1 U3733 ( .A1(n6046), .A2(STATE2_REG_3__SCAN_IN), .ZN(n6059) );
  INV_X1 U3734 ( .A(n6065), .ZN(n6083) );
  INV_X1 U3735 ( .A(n6047), .ZN(n6087) );
  AND2_X1 U3736 ( .A1(n5191), .A2(n5971), .ZN(n6058) );
  OR2_X1 U3737 ( .A1(n4293), .A2(n4298), .ZN(n5430) );
  INV_X1 U3738 ( .A(n5555), .ZN(n6092) );
  NAND2_X1 U3739 ( .A1(n4396), .A2(n6131), .ZN(n5397) );
  BUF_X1 U3740 ( .A(n6123), .Z(n6118) );
  INV_X1 U3741 ( .A(n6486), .ZN(n6597) );
  CLKBUF_X2 U3742 ( .A(n6208), .Z(n6201) );
  INV_X1 U3743 ( .A(n6131), .ZN(n6207) );
  XNOR2_X1 U3744 ( .A(n4278), .B(n4277), .ZN(n4313) );
  OR2_X1 U3745 ( .A1(n4276), .A2(n5408), .ZN(n4278) );
  XNOR2_X1 U3746 ( .A(n4275), .B(n4274), .ZN(n5399) );
  AND2_X1 U3747 ( .A1(n5278), .A2(n5277), .ZN(n5279) );
  INV_X1 U3749 ( .A(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n4846) );
  NAND2_X1 U3750 ( .A1(n6221), .A2(n3878), .ZN(n5691) );
  OAI21_X1 U3751 ( .B1(INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n5404), .A(n5403), 
        .ZN(n5405) );
  OR2_X1 U3752 ( .A1(n5430), .A2(n6337), .ZN(n4304) );
  AND2_X1 U3753 ( .A1(n5767), .A2(n4211), .ZN(n5751) );
  AND2_X1 U3754 ( .A1(n5778), .A2(n5630), .ZN(n5756) );
  AND2_X1 U3755 ( .A1(n5817), .A2(n5338), .ZN(n6324) );
  OR2_X1 U3756 ( .A1(n4244), .A2(n6462), .ZN(n5909) );
  INV_X1 U3757 ( .A(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n5031) );
  CLKBUF_X1 U3758 ( .A(n4483), .Z(n5827) );
  INV_X1 U3759 ( .A(STATE2_REG_1__SCAN_IN), .ZN(n5413) );
  CLKBUF_X1 U3760 ( .A(n3181), .Z(n3182) );
  AND2_X1 U3761 ( .A1(n4475), .A2(STATE2_REG_3__SCAN_IN), .ZN(n5415) );
  INV_X1 U3762 ( .A(n5137), .ZN(n5173) );
  OAI211_X1 U3763 ( .C1(n6389), .C2(n6581), .A(n6359), .B(n6474), .ZN(n6393)
         );
  NAND2_X1 U3764 ( .A1(n4601), .A2(n4795), .ZN(n6457) );
  NOR2_X1 U3765 ( .A1(n4532), .A2(n4749), .ZN(n5137) );
  INV_X1 U3766 ( .A(STATE2_REG_0__SCAN_IN), .ZN(n6498) );
  NAND2_X1 U3767 ( .A1(n5577), .A2(n6036), .ZN(n4321) );
  NAND2_X1 U3768 ( .A1(n5577), .A2(n4149), .ZN(n4152) );
  INV_X1 U3769 ( .A(n5577), .ZN(n5580) );
  INV_X1 U3770 ( .A(n4332), .ZN(n4333) );
  OAI21_X1 U3771 ( .B1(n5420), .B2(n5697), .A(n4331), .ZN(n4332) );
  INV_X4 U3772 ( .A(n5683), .ZN(n5629) );
  OR2_X2 U3773 ( .A1(n3070), .A2(n3069), .ZN(n3144) );
  INV_X1 U3774 ( .A(n3164), .ZN(n5396) );
  INV_X1 U3775 ( .A(n2995), .ZN(n4750) );
  AND2_X1 U3776 ( .A1(n5999), .A2(n5218), .ZN(n5217) );
  NAND2_X1 U3777 ( .A1(n5629), .A2(n5790), .ZN(n2998) );
  OR2_X1 U3778 ( .A1(n4295), .A2(n4153), .ZN(n2999) );
  NAND2_X1 U3779 ( .A1(n5629), .A2(n5674), .ZN(n3000) );
  OR2_X1 U3780 ( .A1(n3132), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3001)
         );
  AND4_X1 U3781 ( .A1(n3012), .A2(n3011), .A3(n3010), .A4(n3009), .ZN(n3002)
         );
  NAND2_X1 U3782 ( .A1(n3919), .A2(n3918), .ZN(n3003) );
  INV_X1 U3783 ( .A(n3560), .ZN(n3756) );
  INV_X1 U3784 ( .A(n5576), .ZN(n4149) );
  INV_X1 U3785 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3153) );
  NAND4_X1 U3786 ( .A1(n3049), .A2(n3048), .A3(n3047), .A4(n3046), .ZN(n3115)
         );
  INV_X1 U3787 ( .A(n6095), .ZN(n4150) );
  AND3_X1 U3788 ( .A1(n4220), .A2(n5630), .A3(n4219), .ZN(n3004) );
  AND2_X1 U3789 ( .A1(n5683), .A2(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n3005)
         );
  OR2_X1 U3790 ( .A1(n6126), .A2(n6479), .ZN(n6221) );
  INV_X1 U3791 ( .A(n6221), .ZN(n6243) );
  INV_X1 U3792 ( .A(n3908), .ZN(n3990) );
  OR2_X1 U3793 ( .A1(n3274), .A2(n3273), .ZN(n3006) );
  AND2_X1 U3794 ( .A1(n3156), .A2(n3135), .ZN(n3117) );
  OR2_X1 U3795 ( .A1(n3140), .A2(n3888), .ZN(n3167) );
  OR2_X1 U3796 ( .A1(n3204), .A2(n3203), .ZN(n3275) );
  NAND2_X1 U3797 ( .A1(n3137), .A2(n3135), .ZN(n4010) );
  OR2_X1 U3798 ( .A1(n3351), .A2(n3350), .ZN(n3401) );
  AND2_X1 U3799 ( .A1(n4518), .A2(n3144), .ZN(n3276) );
  NOR2_X1 U3800 ( .A1(n3140), .A2(n3122), .ZN(n3123) );
  AOI22_X1 U3801 ( .A1(n3106), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n3190), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3074) );
  AND2_X2 U3802 ( .A1(n4420), .A2(n4429), .ZN(n3226) );
  OR3_X1 U3803 ( .A1(n3504), .A2(n6346), .A3(INSTQUEUERD_ADDR_REG_4__SCAN_IN), 
        .ZN(n3498) );
  INV_X1 U3804 ( .A(n5300), .ZN(n3740) );
  OR2_X1 U3805 ( .A1(n3238), .A2(n3237), .ZN(n3429) );
  NAND2_X1 U3806 ( .A1(n3144), .A2(n4181), .ZN(n3888) );
  OR2_X1 U3807 ( .A1(n3437), .A2(n3438), .ZN(n3439) );
  OR2_X1 U3808 ( .A1(n3222), .A2(n3221), .ZN(n3295) );
  INV_X1 U3809 ( .A(n4533), .ZN(n3333) );
  AND2_X1 U3810 ( .A1(n3272), .A2(n3271), .ZN(n3273) );
  AOI22_X1 U3811 ( .A1(n3253), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n3190), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3111) );
  AND4_X1 U3812 ( .A1(n3045), .A2(n3044), .A3(n3043), .A4(n3042), .ZN(n3046)
         );
  OR2_X1 U3813 ( .A1(n3330), .A2(n3329), .ZN(n3355) );
  INV_X1 U3814 ( .A(n5571), .ZN(n3795) );
  OR2_X1 U3815 ( .A1(n3696), .A2(n3695), .ZN(n3709) );
  NAND2_X1 U3816 ( .A1(n3411), .A2(n3410), .ZN(n3423) );
  XNOR2_X1 U3817 ( .A(n3409), .B(n3410), .ZN(n3600) );
  AND2_X1 U3818 ( .A1(n3125), .A2(n3121), .ZN(n3126) );
  AND2_X1 U3819 ( .A1(n3931), .A2(n3930), .ZN(n5226) );
  AND2_X1 U3820 ( .A1(n3901), .A2(n3900), .ZN(n4575) );
  OR2_X1 U3821 ( .A1(n3260), .A2(n3259), .ZN(n3296) );
  AND2_X2 U3822 ( .A1(n3008), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3014)
         );
  OR2_X1 U3823 ( .A1(n4165), .A2(n4164), .ZN(n4249) );
  INV_X1 U3825 ( .A(n5374), .ZN(n3988) );
  OR2_X1 U3826 ( .A1(n4080), .A2(n5436), .ZN(n4144) );
  NOR2_X1 U3827 ( .A1(n3846), .A2(n5650), .ZN(n3864) );
  INV_X1 U3828 ( .A(n4111), .ZN(n4142) );
  INV_X1 U3829 ( .A(n3756), .ZN(n4094) );
  NOR2_X1 U3830 ( .A1(n3164), .A2(n6497), .ZN(n3560) );
  AND2_X1 U3831 ( .A1(n5629), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n4229)
         );
  AND2_X1 U3832 ( .A1(n3126), .A2(n3461), .ZN(n4423) );
  AND2_X1 U3833 ( .A1(n5891), .A2(n3444), .ZN(n5320) );
  INV_X1 U3834 ( .A(n5996), .ZN(n3935) );
  AND2_X1 U3835 ( .A1(n3915), .A2(n3914), .ZN(n4586) );
  INV_X1 U3836 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4434) );
  NAND2_X1 U3837 ( .A1(n3362), .A2(n3006), .ZN(n4482) );
  INV_X1 U3838 ( .A(n5096), .ZN(n5139) );
  OR2_X1 U3839 ( .A1(n3180), .A2(n4434), .ZN(n3317) );
  XNOR2_X1 U3840 ( .A(n3294), .B(n3293), .ZN(n4483) );
  INV_X1 U3841 ( .A(n3811), .ZN(n4139) );
  NAND2_X1 U3842 ( .A1(n3512), .A2(n4165), .ZN(n3513) );
  NAND2_X1 U3843 ( .A1(n3875), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n4038)
         );
  NAND2_X1 U3844 ( .A1(n3810), .A2(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n3828)
         );
  NAND2_X1 U3845 ( .A1(n3710), .A2(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n3724)
         );
  NAND2_X1 U3846 ( .A1(n3682), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n3655)
         );
  AND2_X1 U3847 ( .A1(n4567), .A2(n4566), .ZN(n4565) );
  INV_X1 U3848 ( .A(n6059), .ZN(n6078) );
  INV_X1 U3849 ( .A(n3997), .ZN(n3998) );
  NOR2_X1 U3850 ( .A1(n5431), .A2(n5432), .ZN(n4324) );
  NOR2_X1 U3851 ( .A1(n4562), .A2(n4561), .ZN(n4563) );
  AND2_X1 U3852 ( .A1(n3864), .A2(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n3875)
         );
  AND2_X1 U3853 ( .A1(n5671), .A2(n5670), .ZN(n5673) );
  NOR2_X1 U3854 ( .A1(n3624), .A2(n6002), .ZN(n3619) );
  AND2_X1 U3855 ( .A1(n3603), .A2(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n3682)
         );
  INV_X1 U3856 ( .A(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n4234) );
  NAND2_X1 U3857 ( .A1(n5404), .A2(n4291), .ZN(n4292) );
  NOR2_X2 U3858 ( .A1(n5506), .A2(n5381), .ZN(n5476) );
  INV_X1 U3859 ( .A(n5641), .ZN(n5642) );
  INV_X1 U3860 ( .A(n5286), .ZN(n5575) );
  NAND2_X1 U3861 ( .A1(n5217), .A2(n5903), .ZN(n5905) );
  AND2_X1 U3862 ( .A1(n5225), .A2(n3935), .ZN(n5999) );
  OAI21_X1 U3863 ( .B1(n6330), .B2(n5337), .A(n5336), .ZN(n5817) );
  NAND2_X1 U3864 ( .A1(n4796), .A2(n2995), .ZN(n4961) );
  INV_X1 U3865 ( .A(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6474) );
  AND2_X1 U3866 ( .A1(n5827), .A2(n4711), .ZN(n4600) );
  INV_X1 U3867 ( .A(n6418), .ZN(n5121) );
  INV_X1 U3868 ( .A(n5831), .ZN(n4915) );
  NAND2_X1 U3869 ( .A1(n4601), .A2(n4600), .ZN(n6450) );
  NAND2_X1 U3870 ( .A1(n3317), .A2(n3316), .ZN(n4864) );
  INV_X1 U3871 ( .A(n4600), .ZN(n4749) );
  INV_X1 U3872 ( .A(n4139), .ZN(n4256) );
  NAND2_X1 U3873 ( .A1(n3514), .A2(n3513), .ZN(n4475) );
  OR2_X1 U3874 ( .A1(n3828), .A2(n3827), .ZN(n3846) );
  NOR2_X1 U3875 ( .A1(n3790), .A2(n3789), .ZN(n3810) );
  INV_X1 U3876 ( .A(n6030), .ZN(n6072) );
  AND2_X1 U3877 ( .A1(n6046), .A2(n4314), .ZN(n5194) );
  NAND2_X1 U3878 ( .A1(n5181), .A2(n5180), .ZN(n5227) );
  OR2_X1 U3879 ( .A1(n5551), .A2(n5497), .ZN(n5499) );
  CLKBUF_X1 U3880 ( .A(n4583), .Z(n4790) );
  CLKBUF_X2 U3881 ( .A(n3133), .Z(n4360) );
  NOR2_X1 U3882 ( .A1(n6597), .A2(n4361), .ZN(n6123) );
  OR2_X1 U3883 ( .A1(n5549), .A2(n5548), .ZN(n5551) );
  NOR2_X1 U3884 ( .A1(n5673), .A2(n5672), .ZN(n5701) );
  NOR2_X1 U3885 ( .A1(n5280), .A2(n5279), .ZN(n6218) );
  NAND2_X1 U3886 ( .A1(n3585), .A2(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n3591)
         );
  NAND2_X1 U3887 ( .A1(PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n3563) );
  OAI22_X1 U3888 ( .A1(n5632), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .B1(n5643), .B2(n3456), .ZN(n3457) );
  INV_X1 U3889 ( .A(n6324), .ZN(n6314) );
  INV_X1 U3890 ( .A(n6300), .ZN(n6340) );
  INV_X1 U3891 ( .A(n6337), .ZN(n6323) );
  INV_X1 U3892 ( .A(n5826), .ZN(n5835) );
  OAI21_X1 U3893 ( .B1(n5136), .B2(n5135), .A(n5134), .ZN(n5170) );
  AND2_X1 U3894 ( .A1(n4641), .A2(n2995), .ZN(n4647) );
  AND2_X1 U3895 ( .A1(n4647), .A2(n4711), .ZN(n4838) );
  INV_X1 U3896 ( .A(n5041), .ZN(n4921) );
  AND2_X1 U3897 ( .A1(n4668), .A2(n4600), .ZN(n6418) );
  AND2_X1 U3898 ( .A1(n4620), .A2(n4711), .ZN(n5017) );
  AND2_X1 U3899 ( .A1(n5827), .A2(n4861), .ZN(n4795) );
  INV_X1 U3900 ( .A(n4870), .ZN(n5074) );
  INV_X1 U3901 ( .A(n4744), .ZN(n4521) );
  INV_X1 U3902 ( .A(n6595), .ZN(n5193) );
  NAND2_X1 U3903 ( .A1(n5399), .A2(n6036), .ZN(n4280) );
  NAND2_X1 U3904 ( .A1(n6046), .A2(n4279), .ZN(n5971) );
  OR2_X1 U3905 ( .A1(n5193), .A2(n4312), .ZN(n6030) );
  NAND2_X1 U3906 ( .A1(n5399), .A2(n5398), .ZN(n5401) );
  OR3_X1 U3907 ( .A1(n6126), .A2(n4359), .A3(n6519), .ZN(n6125) );
  AND2_X1 U3908 ( .A1(n3886), .A2(n3885), .ZN(n3887) );
  NAND2_X1 U3909 ( .A1(n5691), .A2(n3881), .ZN(n6249) );
  AND2_X1 U3910 ( .A1(n4304), .A2(n4303), .ZN(n4305) );
  OR2_X1 U3911 ( .A1(n4244), .A2(n4180), .ZN(n6337) );
  OR2_X1 U3912 ( .A1(n4244), .A2(n4243), .ZN(n6300) );
  NAND2_X1 U3913 ( .A1(n4647), .A2(n4861), .ZN(n5178) );
  INV_X1 U3914 ( .A(n4803), .ZN(n4841) );
  NAND2_X1 U3915 ( .A1(n4674), .A2(n4861), .ZN(n4787) );
  NAND2_X1 U3916 ( .A1(n4668), .A2(n4795), .ZN(n6424) );
  NAND2_X1 U3917 ( .A1(n4620), .A2(n4861), .ZN(n5127) );
  INV_X1 U3918 ( .A(n4983), .ZN(n5023) );
  NOR2_X1 U3919 ( .A1(n4869), .A2(n4868), .ZN(n4908) );
  NAND2_X1 U3920 ( .A1(n4862), .A2(n4711), .ZN(n5076) );
  INV_X1 U3921 ( .A(n4488), .ZN(n4525) );
  INV_X1 U3922 ( .A(n6578), .ZN(n6511) );
  INV_X1 U3923 ( .A(n6565), .ZN(n6804) );
  AND2_X2 U3924 ( .A1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4420) );
  AND2_X2 U3925 ( .A1(n5838), .A2(n4420), .ZN(n3190) );
  AND2_X2 U3926 ( .A1(n5839), .A2(n4420), .ZN(n3231) );
  AOI22_X1 U3927 ( .A1(n3190), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n3231), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3012) );
  NOR2_X4 U3928 ( .A1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4430) );
  AND2_X2 U3929 ( .A1(n5838), .A2(n4430), .ZN(n3225) );
  NOR2_X4 U3930 ( .A1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4463) );
  AOI22_X1 U3931 ( .A1(n3225), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n3196), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3011) );
  INV_X1 U3932 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3008) );
  AND2_X4 U3933 ( .A1(n3014), .A2(n4429), .ZN(n3254) );
  AOI22_X1 U3934 ( .A1(n3254), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n3107), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3010) );
  AND2_X4 U3935 ( .A1(n4430), .A2(n4429), .ZN(n3324) );
  AOI22_X1 U3936 ( .A1(n3324), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .B1(n2997), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3009) );
  AND2_X4 U3937 ( .A1(n3013), .A2(n5838), .ZN(n4127) );
  AOI22_X1 U3938 ( .A1(n4127), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3832), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3018) );
  AND2_X2 U3939 ( .A1(n5838), .A2(n3014), .ZN(n3253) );
  AND2_X2 U3940 ( .A1(n3013), .A2(n4429), .ZN(n3191) );
  AOI22_X1 U3941 ( .A1(n3253), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n3191), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n3017) );
  AOI22_X1 U3942 ( .A1(n3198), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n3226), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3016) );
  AOI22_X1 U3943 ( .A1(n3608), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3106), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3015) );
  AND2_X2 U3944 ( .A1(n3002), .A2(n3019), .ZN(n3137) );
  AOI22_X1 U3945 ( .A1(n3253), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3190), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3023) );
  AOI22_X1 U3946 ( .A1(n3231), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3107), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3022) );
  AOI22_X1 U3947 ( .A1(n3191), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3254), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3021) );
  AOI22_X1 U3948 ( .A1(n3225), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n3196), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3027) );
  AOI22_X1 U3949 ( .A1(n3197), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n3832), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3025) );
  NAND2_X1 U3950 ( .A1(n3106), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3033) );
  NAND2_X1 U3951 ( .A1(n3608), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3032) );
  NAND2_X1 U3952 ( .A1(n3253), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3031) );
  NAND2_X1 U3953 ( .A1(n3190), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3030)
         );
  NAND2_X1 U3954 ( .A1(n3832), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3037) );
  NAND2_X1 U3955 ( .A1(n4127), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n3036)
         );
  NAND2_X1 U3956 ( .A1(n3324), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3035) );
  NAND2_X1 U3957 ( .A1(n3197), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3034)
         );
  NAND2_X1 U3958 ( .A1(n3225), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3041) );
  NAND2_X1 U3959 ( .A1(n3196), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3040) );
  NAND2_X1 U3960 ( .A1(n3198), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3039) );
  NAND2_X1 U3961 ( .A1(n3226), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3038)
         );
  NAND2_X1 U3962 ( .A1(n3231), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3045)
         );
  NAND2_X1 U3963 ( .A1(n3191), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n3044)
         );
  NAND2_X1 U3964 ( .A1(n3254), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3043) );
  NAND2_X1 U3965 ( .A1(n3107), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3042) );
  NAND2_X1 U3966 ( .A1(n4010), .A2(n3136), .ZN(n3169) );
  INV_X1 U3967 ( .A(n3169), .ZN(n3060) );
  AOI22_X1 U3968 ( .A1(n3608), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3106), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3053) );
  AOI22_X1 U3969 ( .A1(n3253), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n3190), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3052) );
  AOI22_X1 U3970 ( .A1(n3191), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3254), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n3051) );
  AOI22_X1 U3971 ( .A1(n3231), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3107), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3050) );
  NAND4_X1 U3972 ( .A1(n3053), .A2(n3052), .A3(n3051), .A4(n3050), .ZN(n3059)
         );
  AOI22_X1 U3973 ( .A1(n3832), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n3197), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n3057) );
  AOI22_X1 U3974 ( .A1(n4127), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3324), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3056) );
  AOI22_X1 U3975 ( .A1(n3225), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n3196), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3055) );
  AOI22_X1 U3976 ( .A1(n3198), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n3226), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3054) );
  NAND4_X1 U3977 ( .A1(n3057), .A2(n3056), .A3(n3055), .A4(n3054), .ZN(n3058)
         );
  NAND2_X1 U3978 ( .A1(n3060), .A2(n3164), .ZN(n3134) );
  AOI22_X1 U3979 ( .A1(n3191), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3254), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3064) );
  AOI22_X1 U3980 ( .A1(n3608), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3106), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3063) );
  AOI22_X1 U3981 ( .A1(n3253), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3190), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3062) );
  AOI22_X1 U3982 ( .A1(n3231), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3107), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3061) );
  NAND4_X1 U3983 ( .A1(n3064), .A2(n3063), .A3(n3062), .A4(n3061), .ZN(n3070)
         );
  AOI22_X1 U3984 ( .A1(n3832), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n3197), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3068) );
  AOI22_X1 U3985 ( .A1(n4127), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3324), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3067) );
  AOI22_X1 U3986 ( .A1(n3225), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n3196), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3066) );
  AOI22_X1 U3987 ( .A1(n3198), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n3226), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3065) );
  NAND4_X1 U3988 ( .A1(n3068), .A2(n3067), .A3(n3066), .A4(n3065), .ZN(n3069)
         );
  NOR2_X2 U3989 ( .A1(n3134), .A2(n3121), .ZN(n3161) );
  AOI22_X1 U3990 ( .A1(n3253), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n3191), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n3073) );
  AOI22_X1 U3991 ( .A1(n4127), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3198), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3072) );
  AOI22_X1 U3992 ( .A1(n3225), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n3254), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3071) );
  NAND4_X1 U3993 ( .A1(n3074), .A2(n3073), .A3(n3072), .A4(n3071), .ZN(n3080)
         );
  AOI22_X1 U3994 ( .A1(n3608), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3231), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3078) );
  AOI22_X1 U3995 ( .A1(n3196), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3107), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3077) );
  AOI22_X1 U3996 ( .A1(n3832), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n3197), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3076) );
  AOI22_X1 U3997 ( .A1(n3324), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .B1(n3226), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3075) );
  NAND4_X1 U3998 ( .A1(n3078), .A2(n3077), .A3(n3076), .A4(n3075), .ZN(n3079)
         );
  INV_X2 U3999 ( .A(n3137), .ZN(n3156) );
  NAND2_X1 U4000 ( .A1(n3161), .A2(n3125), .ZN(n4167) );
  INV_X1 U4001 ( .A(n4167), .ZN(n3101) );
  NAND2_X1 U4002 ( .A1(n4127), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3084)
         );
  NAND2_X1 U4003 ( .A1(n3191), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3083)
         );
  NAND2_X1 U4004 ( .A1(n3226), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3082)
         );
  NAND2_X1 U4005 ( .A1(n3197), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3081)
         );
  NAND2_X1 U4006 ( .A1(n3106), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3088) );
  NAND2_X1 U4007 ( .A1(n3608), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3087) );
  NAND2_X1 U4008 ( .A1(n3196), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3086) );
  NAND2_X1 U4009 ( .A1(n3254), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3085) );
  NAND2_X1 U4010 ( .A1(n3253), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3092) );
  NAND2_X1 U4011 ( .A1(n3190), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3091)
         );
  NAND2_X1 U4012 ( .A1(n3231), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3090)
         );
  NAND2_X1 U4013 ( .A1(n3107), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3089) );
  NAND2_X1 U4014 ( .A1(n3198), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3096) );
  NAND2_X1 U4015 ( .A1(n3225), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3095) );
  NAND2_X1 U4016 ( .A1(n3832), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3094) );
  NAND2_X1 U4017 ( .A1(n3324), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3093) );
  NAND2_X1 U4018 ( .A1(n3101), .A2(n4360), .ZN(n4247) );
  AOI22_X1 U4019 ( .A1(n4127), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n3324), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3104) );
  AOI22_X1 U4020 ( .A1(n3225), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n3196), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3103) );
  AOI22_X1 U4021 ( .A1(n3198), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n3226), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3102) );
  NAND4_X1 U4022 ( .A1(n3105), .A2(n3104), .A3(n3103), .A4(n3102), .ZN(n3113)
         );
  AOI22_X1 U4023 ( .A1(n3608), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n3106), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3110) );
  AOI22_X1 U4024 ( .A1(n3191), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n3254), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3109) );
  AOI22_X1 U4025 ( .A1(n3231), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n3107), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3108) );
  NAND4_X1 U4026 ( .A1(n3111), .A2(n3110), .A3(n3109), .A4(n3108), .ZN(n3112)
         );
  NAND2_X1 U4027 ( .A1(STATE_REG_1__SCAN_IN), .A2(STATE_REG_2__SCAN_IN), .ZN(
        n6514) );
  OAI21_X1 U4028 ( .B1(STATE_REG_1__SCAN_IN), .B2(STATE_REG_2__SCAN_IN), .A(
        n6514), .ZN(n4159) );
  OAI21_X1 U4029 ( .B1(n3554), .B2(n3115), .A(n3164), .ZN(n3116) );
  INV_X1 U4030 ( .A(n3116), .ZN(n3120) );
  NAND2_X1 U4031 ( .A1(n3140), .A2(n4182), .ZN(n3119) );
  NAND2_X1 U4032 ( .A1(n3117), .A2(n3298), .ZN(n3118) );
  NAND3_X1 U4033 ( .A1(n3120), .A2(n3119), .A3(n3118), .ZN(n3147) );
  INV_X1 U4034 ( .A(n3147), .ZN(n3124) );
  NAND2_X1 U4035 ( .A1(n4002), .A2(n4513), .ZN(n4236) );
  NAND2_X1 U4036 ( .A1(n4423), .A2(n4398), .ZN(n4238) );
  NAND2_X1 U4037 ( .A1(n3128), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3151) );
  NOR2_X1 U4038 ( .A1(STATE2_REG_1__SCAN_IN), .A2(STATE2_REG_3__SCAN_IN), .ZN(
        n5840) );
  NAND2_X1 U4039 ( .A1(n5840), .A2(n6498), .ZN(n3882) );
  INV_X1 U4040 ( .A(n3882), .ZN(n3187) );
  NAND2_X1 U4041 ( .A1(n6464), .A2(n5031), .ZN(n3129) );
  NAND2_X1 U4042 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3184) );
  NAND2_X1 U4043 ( .A1(n3187), .A2(n4866), .ZN(n3131) );
  INV_X1 U4044 ( .A(n3515), .ZN(n3186) );
  NAND2_X1 U4045 ( .A1(n3186), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3130) );
  INV_X1 U4046 ( .A(n3150), .ZN(n3132) );
  NAND2_X1 U4047 ( .A1(n3517), .A2(n4360), .ZN(n4004) );
  NAND2_X1 U4048 ( .A1(n3139), .A2(n3138), .ZN(n3141) );
  OAI211_X1 U4049 ( .C1(n4004), .C2(n4509), .A(n3141), .B(n3167), .ZN(n3142)
         );
  AOI21_X1 U4050 ( .B1(n3162), .B2(n3134), .A(n3142), .ZN(n3148) );
  AND2_X1 U4051 ( .A1(n3144), .A2(n3164), .ZN(n3143) );
  NAND2_X1 U4052 ( .A1(n3276), .A2(n3517), .ZN(n3145) );
  NAND2_X1 U4053 ( .A1(n4518), .A2(n4181), .ZN(n5192) );
  NAND2_X1 U4054 ( .A1(n3145), .A2(n5192), .ZN(n3146) );
  AOI21_X1 U4055 ( .B1(n3147), .B2(n4518), .A(n3146), .ZN(n3155) );
  NAND3_X1 U4056 ( .A1(n3148), .A2(n4189), .A3(n3155), .ZN(n3149) );
  NAND2_X1 U4057 ( .A1(n3152), .A2(n3178), .ZN(n3212) );
  INV_X1 U4058 ( .A(n3212), .ZN(n3177) );
  MUX2_X1 U4059 ( .A(n3515), .B(n3882), .S(n5031), .Z(n3154) );
  INV_X1 U4060 ( .A(n3155), .ZN(n3159) );
  NAND2_X1 U4061 ( .A1(n3464), .A2(n4509), .ZN(n3158) );
  NAND2_X1 U4062 ( .A1(n3159), .A2(n3158), .ZN(n3160) );
  NAND2_X1 U4063 ( .A1(n3160), .A2(n4007), .ZN(n4191) );
  INV_X1 U4064 ( .A(n4191), .ZN(n3176) );
  INV_X1 U4065 ( .A(n3161), .ZN(n3163) );
  NAND2_X1 U4066 ( .A1(n3163), .A2(n6130), .ZN(n3174) );
  NAND2_X1 U4067 ( .A1(n3207), .A2(n3164), .ZN(n3516) );
  INV_X1 U4068 ( .A(n3516), .ZN(n3166) );
  NOR2_X1 U4069 ( .A1(n4182), .A2(n3554), .ZN(n3165) );
  NAND3_X1 U4070 ( .A1(n3166), .A2(n3121), .A3(n3165), .ZN(n4456) );
  NAND2_X1 U4071 ( .A1(n5840), .A2(STATE2_REG_0__SCAN_IN), .ZN(n6501) );
  AOI21_X1 U4072 ( .B1(n4182), .B2(n4360), .A(n6501), .ZN(n3168) );
  AND3_X1 U4073 ( .A1(n4456), .A2(n3168), .A3(n3167), .ZN(n3173) );
  AND2_X1 U4074 ( .A1(n3169), .A2(n3517), .ZN(n3171) );
  OAI21_X1 U4075 ( .B1(n3171), .B2(n3170), .A(n4181), .ZN(n3172) );
  NAND2_X1 U4076 ( .A1(n3176), .A2(n3175), .ZN(n3245) );
  NAND2_X1 U4077 ( .A1(n3177), .A2(n3210), .ZN(n3179) );
  NAND2_X1 U4078 ( .A1(n3179), .A2(n2996), .ZN(n3312) );
  INV_X1 U4079 ( .A(n3184), .ZN(n3183) );
  NAND2_X1 U4080 ( .A1(n3183), .A2(n6468), .ZN(n4918) );
  NAND2_X1 U4081 ( .A1(n3184), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3185) );
  NAND2_X1 U4082 ( .A1(n4918), .A2(n3185), .ZN(n4718) );
  AOI22_X1 U4083 ( .A1(n3187), .A2(n4718), .B1(n3186), .B2(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3188) );
  XNOR2_X1 U4084 ( .A(n3312), .B(n3310), .ZN(n4449) );
  NAND2_X1 U4085 ( .A1(n4449), .A2(n6498), .ZN(n3206) );
  AOI22_X1 U4086 ( .A1(n3853), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n4116), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3195) );
  AOI22_X1 U4087 ( .A1(n4117), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n4021), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3194) );
  AOI22_X1 U4088 ( .A1(n4063), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n2992), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3193) );
  AOI22_X1 U4089 ( .A1(n4125), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n4022), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3192) );
  NAND4_X1 U4090 ( .A1(n3195), .A2(n3194), .A3(n3193), .A4(n3192), .ZN(n3204)
         );
  AOI22_X1 U4091 ( .A1(n2994), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .B1(n4119), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3202) );
  BUF_X1 U4092 ( .A(n4127), .Z(n3675) );
  AOI22_X1 U4093 ( .A1(n3675), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3324), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3201) );
  AOI22_X1 U4094 ( .A1(n4120), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n4027), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3200) );
  AOI22_X1 U4095 ( .A1(n4126), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n4118), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3199) );
  NAND4_X1 U4096 ( .A1(n3202), .A2(n3201), .A3(n3200), .A4(n3199), .ZN(n3203)
         );
  NAND2_X1 U4097 ( .A1(n3240), .A2(n3275), .ZN(n3205) );
  INV_X1 U4098 ( .A(n3318), .ZN(n3241) );
  AOI22_X1 U4099 ( .A1(n3499), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n3241), 
        .B2(n3275), .ZN(n3208) );
  XNOR2_X1 U4100 ( .A(n3212), .B(n3211), .ZN(n4484) );
  AOI22_X1 U4101 ( .A1(n4117), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n4125), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3216) );
  AOI22_X1 U4102 ( .A1(INSTQUEUE_REG_9__1__SCAN_IN), .A2(n4119), .B1(n2994), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3215) );
  AOI22_X1 U4103 ( .A1(n4063), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n4022), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3214) );
  AOI22_X1 U4104 ( .A1(n4127), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n4118), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3213) );
  NAND4_X1 U4105 ( .A1(n3216), .A2(n3215), .A3(n3214), .A4(n3213), .ZN(n3222)
         );
  AOI22_X1 U4106 ( .A1(n3853), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n4116), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3220) );
  AOI22_X1 U4107 ( .A1(n4021), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n2992), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3219) );
  AOI22_X1 U4108 ( .A1(INSTQUEUE_REG_2__1__SCAN_IN), .A2(n4126), .B1(n3324), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3218) );
  AOI22_X1 U4109 ( .A1(INSTQUEUE_REG_5__1__SCAN_IN), .A2(n4120), .B1(n4027), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3217) );
  NAND4_X1 U4110 ( .A1(n3220), .A2(n3219), .A3(n3218), .A4(n3217), .ZN(n3221)
         );
  NAND2_X1 U4111 ( .A1(n3240), .A2(n3295), .ZN(n3223) );
  NAND2_X1 U4112 ( .A1(n3499), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3243) );
  AOI22_X1 U4113 ( .A1(n4116), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n4117), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n3230) );
  AOI22_X1 U4114 ( .A1(n3675), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3198), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3229) );
  AOI22_X1 U4115 ( .A1(n4063), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n2992), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3228) );
  AOI22_X1 U4116 ( .A1(n2994), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n4118), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3227) );
  NAND4_X1 U4117 ( .A1(n3230), .A2(n3229), .A3(n3228), .A4(n3227), .ZN(n3238)
         );
  AOI22_X1 U4118 ( .A1(n3853), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n4021), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3236) );
  AOI22_X1 U4119 ( .A1(n4125), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n4022), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3235) );
  AOI22_X1 U4120 ( .A1(n3196), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3232), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3234) );
  AOI22_X1 U4121 ( .A1(n4120), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n4027), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3233) );
  NAND4_X1 U4122 ( .A1(n3236), .A2(n3235), .A3(n3234), .A4(n3233), .ZN(n3237)
         );
  INV_X1 U4123 ( .A(n3429), .ZN(n3239) );
  NAND2_X1 U4124 ( .A1(n3240), .A2(n3239), .ZN(n3248) );
  NAND2_X1 U4125 ( .A1(n3241), .A2(n3295), .ZN(n3242) );
  NAND2_X1 U4126 ( .A1(n3292), .A2(n3244), .ZN(n3269) );
  INV_X1 U4127 ( .A(n3245), .ZN(n3247) );
  INV_X1 U4128 ( .A(n3248), .ZN(n3261) );
  NAND2_X1 U4129 ( .A1(n4509), .A2(n3429), .ZN(n3263) );
  AOI22_X1 U4130 ( .A1(n3853), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n4116), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3252) );
  AOI22_X1 U4131 ( .A1(n2994), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .B1(n3198), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3251) );
  AOI22_X1 U4132 ( .A1(n3196), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n4022), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3250) );
  AOI22_X1 U4133 ( .A1(n4127), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n4027), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3249) );
  NAND4_X1 U4134 ( .A1(n3252), .A2(n3251), .A3(n3250), .A4(n3249), .ZN(n3260)
         );
  AOI22_X1 U4135 ( .A1(n4117), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n4021), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3258) );
  AOI22_X1 U4136 ( .A1(n4125), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n4063), 
        .B2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3257) );
  AOI22_X1 U4137 ( .A1(n2992), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n4118), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3256) );
  AOI22_X1 U4138 ( .A1(n4120), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n3324), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3255) );
  NAND4_X1 U4139 ( .A1(n3258), .A2(n3257), .A3(n3256), .A4(n3255), .ZN(n3259)
         );
  MUX2_X1 U4140 ( .A(n3261), .B(n3424), .S(n3264), .Z(n3262) );
  NAND2_X1 U4141 ( .A1(n3279), .A2(n3283), .ZN(n3268) );
  NAND2_X1 U4142 ( .A1(n3499), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3267) );
  OAI211_X1 U4143 ( .C1(n3264), .C2(n4360), .A(n3263), .B(
        STATE2_REG_0__SCAN_IN), .ZN(n3265) );
  INV_X1 U4144 ( .A(n3265), .ZN(n3266) );
  NAND2_X1 U4145 ( .A1(n3267), .A2(n3266), .ZN(n3281) );
  NAND2_X1 U4146 ( .A1(n3269), .A2(n3294), .ZN(n3272) );
  INV_X1 U4147 ( .A(n3292), .ZN(n3270) );
  NAND2_X1 U4148 ( .A1(n3270), .A2(n3291), .ZN(n3271) );
  INV_X1 U4149 ( .A(n3464), .ZN(n3425) );
  NAND2_X1 U4150 ( .A1(n3296), .A2(n3295), .ZN(n3337) );
  INV_X1 U4151 ( .A(n3275), .ZN(n3336) );
  XNOR2_X1 U4152 ( .A(n3337), .B(n3336), .ZN(n3277) );
  AOI21_X1 U4153 ( .B1(n3277), .B2(n6130), .A(n3276), .ZN(n3278) );
  OAI21_X2 U4154 ( .B1(n4482), .B2(n3425), .A(n3278), .ZN(n6240) );
  NAND2_X1 U4155 ( .A1(n6240), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n3305)
         );
  NAND2_X1 U4156 ( .A1(n3279), .A2(n3281), .ZN(n3280) );
  NAND2_X1 U4157 ( .A1(n3280), .A2(n3283), .ZN(n3285) );
  INV_X1 U4158 ( .A(n3281), .ZN(n3282) );
  INV_X1 U4159 ( .A(n3276), .ZN(n3286) );
  OAI21_X1 U4160 ( .B1(n6599), .B2(n3296), .A(n3286), .ZN(n3287) );
  INV_X1 U4161 ( .A(n3287), .ZN(n3288) );
  NAND2_X1 U4162 ( .A1(n4352), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n3289)
         );
  INV_X1 U4163 ( .A(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n6331) );
  NAND2_X1 U4164 ( .A1(n3289), .A2(n6331), .ZN(n3290) );
  AND2_X1 U4165 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n6333) );
  NAND2_X1 U4166 ( .A1(n4352), .A2(n6333), .ZN(n3303) );
  AND2_X1 U4167 ( .A1(n3290), .A2(n3303), .ZN(n4378) );
  NAND2_X1 U4168 ( .A1(n4483), .A2(n3464), .ZN(n3302) );
  OAI21_X1 U4169 ( .B1(n3296), .B2(n3295), .A(n3337), .ZN(n3297) );
  INV_X1 U4170 ( .A(n3297), .ZN(n3300) );
  NAND3_X1 U4171 ( .A1(n3298), .A2(n3157), .A3(n3144), .ZN(n3299) );
  AOI21_X1 U4172 ( .B1(n3300), .B2(n6130), .A(n3299), .ZN(n3301) );
  NAND2_X1 U4173 ( .A1(n3302), .A2(n3301), .ZN(n4379) );
  INV_X1 U4174 ( .A(n3303), .ZN(n3304) );
  AOI21_X1 U4175 ( .B1(n4378), .B2(n4379), .A(n3304), .ZN(n6241) );
  NAND2_X1 U4176 ( .A1(n3305), .A2(n6241), .ZN(n3309) );
  INV_X1 U4177 ( .A(n6240), .ZN(n3307) );
  INV_X1 U4178 ( .A(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n3306) );
  NAND2_X1 U4179 ( .A1(n3307), .A2(n3306), .ZN(n3308) );
  AND2_X1 U4180 ( .A1(n3309), .A2(n3308), .ZN(n4540) );
  INV_X1 U4181 ( .A(n3362), .ZN(n3334) );
  INV_X1 U4182 ( .A(n3310), .ZN(n3311) );
  NAND3_X1 U4183 ( .A1(n6474), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6347) );
  INV_X1 U4184 ( .A(n6347), .ZN(n3313) );
  NAND2_X1 U4185 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n3313), .ZN(n4554) );
  NAND2_X1 U4186 ( .A1(n6474), .A2(n4554), .ZN(n3314) );
  NOR3_X1 U4187 ( .A1(n6474), .A2(n6468), .A3(n6464), .ZN(n4489) );
  NAND2_X1 U4188 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4489), .ZN(n4485) );
  NAND2_X1 U4189 ( .A1(n3314), .A2(n4485), .ZN(n4865) );
  OAI22_X1 U4190 ( .A1(n3882), .A2(n4865), .B1(n3515), .B2(n6474), .ZN(n3315)
         );
  INV_X1 U4191 ( .A(n3315), .ZN(n3316) );
  AOI22_X1 U4192 ( .A1(n4117), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n4021), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3323) );
  AOI22_X1 U4193 ( .A1(n4125), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n4119), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n3322) );
  AOI22_X1 U4194 ( .A1(n4126), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n4120), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3321) );
  AOI22_X1 U4195 ( .A1(n2994), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .B1(n4118), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3320) );
  NAND4_X1 U4196 ( .A1(n3323), .A2(n3322), .A3(n3321), .A4(n3320), .ZN(n3330)
         );
  AOI22_X1 U4197 ( .A1(n3853), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n4116), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3328) );
  AOI22_X1 U4198 ( .A1(n3675), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n2992), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3327) );
  AOI22_X1 U4199 ( .A1(n4063), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n4022), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3326) );
  AOI22_X1 U4200 ( .A1(n3324), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n4027), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3325) );
  NAND4_X1 U4201 ( .A1(n3328), .A2(n3327), .A3(n3326), .A4(n3325), .ZN(n3329)
         );
  AOI22_X1 U4202 ( .A1(n3499), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n3507), 
        .B2(n3355), .ZN(n3331) );
  NAND2_X1 U4203 ( .A1(n3334), .A2(n3333), .ZN(n3354) );
  NAND2_X1 U4204 ( .A1(n3362), .A2(n4533), .ZN(n3335) );
  NAND2_X1 U4205 ( .A1(n3354), .A2(n3335), .ZN(n3573) );
  NAND2_X1 U4206 ( .A1(n3337), .A2(n3336), .ZN(n3356) );
  XNOR2_X1 U4207 ( .A(n3356), .B(n3355), .ZN(n3338) );
  OR2_X1 U4208 ( .A1(n3338), .A2(n6599), .ZN(n3339) );
  OAI21_X2 U4209 ( .B1(n3573), .B2(n3425), .A(n3339), .ZN(n3340) );
  INV_X1 U4210 ( .A(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n6328) );
  XNOR2_X1 U4211 ( .A(n3340), .B(n6328), .ZN(n4541) );
  NAND2_X1 U4212 ( .A1(n4540), .A2(n4541), .ZN(n4539) );
  NAND2_X1 U4213 ( .A1(n3340), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n3341)
         );
  NAND2_X1 U4214 ( .A1(n4539), .A2(n3341), .ZN(n6232) );
  NAND2_X1 U4215 ( .A1(n3499), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3353) );
  AOI22_X1 U4216 ( .A1(n3853), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n4116), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3345) );
  AOI22_X1 U4217 ( .A1(n4117), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n4021), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3344) );
  AOI22_X1 U4218 ( .A1(n4063), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n2992), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3343) );
  AOI22_X1 U4219 ( .A1(n4125), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n4022), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3342) );
  NAND4_X1 U4220 ( .A1(n3345), .A2(n3344), .A3(n3343), .A4(n3342), .ZN(n3351)
         );
  AOI22_X1 U4221 ( .A1(n2994), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .B1(n4119), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3349) );
  AOI22_X1 U4222 ( .A1(n3675), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n3232), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3348) );
  AOI22_X1 U4223 ( .A1(n4120), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n4027), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3347) );
  AOI22_X1 U4224 ( .A1(n4126), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .B1(n4118), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3346) );
  NAND4_X1 U4225 ( .A1(n3349), .A2(n3348), .A3(n3347), .A4(n3346), .ZN(n3350)
         );
  NAND2_X1 U4226 ( .A1(n3507), .A2(n3401), .ZN(n3352) );
  NAND2_X1 U4227 ( .A1(n3353), .A2(n3352), .ZN(n3363) );
  XNOR2_X1 U4228 ( .A(n3354), .B(n3363), .ZN(n3589) );
  NAND2_X1 U4229 ( .A1(n3589), .A2(n3464), .ZN(n3359) );
  NAND2_X1 U4230 ( .A1(n3356), .A2(n3355), .ZN(n3403) );
  XNOR2_X1 U4231 ( .A(n3403), .B(n3401), .ZN(n3357) );
  NAND2_X1 U4232 ( .A1(n3357), .A2(n6130), .ZN(n3358) );
  NAND2_X1 U4233 ( .A1(n3359), .A2(n3358), .ZN(n3360) );
  INV_X1 U4234 ( .A(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n6320) );
  XNOR2_X1 U4235 ( .A(n3360), .B(n6320), .ZN(n6231) );
  NAND2_X1 U4236 ( .A1(n6232), .A2(n6231), .ZN(n6230) );
  NAND2_X1 U4237 ( .A1(n3360), .A2(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n3361)
         );
  NAND2_X1 U4238 ( .A1(n6230), .A2(n3361), .ZN(n4844) );
  NAND2_X1 U4239 ( .A1(n3364), .A2(n3363), .ZN(n3385) );
  NAND2_X1 U4240 ( .A1(n3499), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3376) );
  AOI22_X1 U4241 ( .A1(n4116), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n4021), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3368) );
  AOI22_X1 U4242 ( .A1(n4119), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n4126), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3367) );
  AOI22_X1 U4243 ( .A1(n4117), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n2992), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3366) );
  AOI22_X1 U4244 ( .A1(n3675), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n4027), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3365) );
  NAND4_X1 U4245 ( .A1(n3368), .A2(n3367), .A3(n3366), .A4(n3365), .ZN(n3374)
         );
  AOI22_X1 U4246 ( .A1(n3853), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n4125), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3372) );
  AOI22_X1 U4247 ( .A1(n4063), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n4022), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3371) );
  AOI22_X1 U4248 ( .A1(n4120), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n3232), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3370) );
  AOI22_X1 U4249 ( .A1(n2994), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .B1(n4118), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3369) );
  NAND4_X1 U4250 ( .A1(n3372), .A2(n3371), .A3(n3370), .A4(n3369), .ZN(n3373)
         );
  NAND2_X1 U4251 ( .A1(n3507), .A2(n3400), .ZN(n3375) );
  NAND2_X1 U4252 ( .A1(n3376), .A2(n3375), .ZN(n3386) );
  XNOR2_X1 U4253 ( .A(n3385), .B(n3386), .ZN(n3590) );
  NAND2_X1 U4254 ( .A1(n3590), .A2(n3464), .ZN(n3381) );
  INV_X1 U4255 ( .A(n3401), .ZN(n3377) );
  OR2_X1 U4256 ( .A1(n3403), .A2(n3377), .ZN(n3378) );
  XNOR2_X1 U4257 ( .A(n3378), .B(n3400), .ZN(n3379) );
  NAND2_X1 U4258 ( .A1(n3379), .A2(n6130), .ZN(n3380) );
  NAND2_X1 U4259 ( .A1(n3381), .A2(n3380), .ZN(n3383) );
  INV_X1 U4260 ( .A(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n3382) );
  XNOR2_X1 U4261 ( .A(n3383), .B(n3382), .ZN(n4843) );
  NAND2_X1 U4262 ( .A1(n4844), .A2(n4843), .ZN(n4842) );
  NAND2_X1 U4263 ( .A1(n3383), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n3384)
         );
  NAND2_X1 U4264 ( .A1(n4842), .A2(n3384), .ZN(n6224) );
  NAND2_X1 U4265 ( .A1(n3499), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3399) );
  AOI22_X1 U4266 ( .A1(n3853), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n4116), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3391) );
  AOI22_X1 U4267 ( .A1(n4117), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n4021), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3390) );
  AOI22_X1 U4268 ( .A1(n4063), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n2992), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3389) );
  AOI22_X1 U4269 ( .A1(n4125), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n4022), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3388) );
  NAND4_X1 U4270 ( .A1(n3391), .A2(n3390), .A3(n3389), .A4(n3388), .ZN(n3397)
         );
  AOI22_X1 U4271 ( .A1(n2994), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n4119), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n3395) );
  AOI22_X1 U4272 ( .A1(n3675), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3232), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3394) );
  AOI22_X1 U4273 ( .A1(n4120), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n4027), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3393) );
  AOI22_X1 U4274 ( .A1(n4126), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n4118), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3392) );
  NAND4_X1 U4275 ( .A1(n3395), .A2(n3394), .A3(n3393), .A4(n3392), .ZN(n3396)
         );
  NAND2_X1 U4276 ( .A1(n3507), .A2(n3416), .ZN(n3398) );
  NAND2_X1 U4277 ( .A1(n3399), .A2(n3398), .ZN(n3410) );
  NAND2_X1 U4278 ( .A1(n3600), .A2(n3464), .ZN(n3406) );
  NAND2_X1 U4279 ( .A1(n3401), .A2(n3400), .ZN(n3402) );
  OR2_X1 U4280 ( .A1(n3403), .A2(n3402), .ZN(n3415) );
  XNOR2_X1 U4281 ( .A(n3415), .B(n3416), .ZN(n3404) );
  NAND2_X1 U4282 ( .A1(n3404), .A2(n6130), .ZN(n3405) );
  NAND2_X1 U4283 ( .A1(n3406), .A2(n3405), .ZN(n3407) );
  INV_X1 U4284 ( .A(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n6304) );
  XNOR2_X1 U4285 ( .A(n3407), .B(n6304), .ZN(n6223) );
  NAND2_X1 U4286 ( .A1(n6224), .A2(n6223), .ZN(n6222) );
  NAND2_X1 U4287 ( .A1(n3407), .A2(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n3408)
         );
  NAND2_X1 U4288 ( .A1(n6222), .A2(n3408), .ZN(n4857) );
  NAND2_X1 U4289 ( .A1(n3499), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3413) );
  NAND2_X1 U4290 ( .A1(n3507), .A2(n3429), .ZN(n3412) );
  NAND2_X1 U4291 ( .A1(n3413), .A2(n3412), .ZN(n3414) );
  INV_X1 U4292 ( .A(n3415), .ZN(n3417) );
  NAND2_X1 U4293 ( .A1(n3417), .A2(n3416), .ZN(n3428) );
  XNOR2_X1 U4294 ( .A(n3428), .B(n3429), .ZN(n3418) );
  NAND2_X1 U4295 ( .A1(n3418), .A2(n6130), .ZN(n3419) );
  NAND2_X1 U4296 ( .A1(n3420), .A2(n3419), .ZN(n3421) );
  INV_X1 U4297 ( .A(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n6295) );
  XNOR2_X1 U4298 ( .A(n3421), .B(n6295), .ZN(n4856) );
  NAND2_X1 U4299 ( .A1(n4857), .A2(n4856), .ZN(n4855) );
  NAND2_X1 U4300 ( .A1(n3421), .A2(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n3422)
         );
  NAND2_X1 U4301 ( .A1(n4855), .A2(n3422), .ZN(n4969) );
  INV_X1 U4302 ( .A(n3424), .ZN(n3426) );
  NOR2_X1 U4303 ( .A1(n3426), .A2(n3425), .ZN(n3427) );
  INV_X1 U4304 ( .A(n3428), .ZN(n3430) );
  NAND3_X1 U4305 ( .A1(n3430), .A2(n6130), .A3(n3429), .ZN(n3431) );
  NAND2_X1 U4306 ( .A1(n3437), .A2(n3431), .ZN(n3432) );
  INV_X1 U4307 ( .A(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n3922) );
  XNOR2_X1 U4308 ( .A(n3432), .B(n3922), .ZN(n4968) );
  NAND2_X1 U4309 ( .A1(n4969), .A2(n4968), .ZN(n4967) );
  NAND2_X1 U4310 ( .A1(n3432), .A2(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n3433)
         );
  NAND2_X1 U4311 ( .A1(n4967), .A2(n3433), .ZN(n5186) );
  INV_X1 U4312 ( .A(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n5184) );
  NAND2_X1 U4313 ( .A1(n5629), .A2(n5184), .ZN(n3434) );
  NAND2_X1 U4314 ( .A1(n5186), .A2(n3434), .ZN(n3436) );
  OR2_X1 U4315 ( .A1(n5629), .A2(n5184), .ZN(n3435) );
  NAND2_X1 U4316 ( .A1(n3436), .A2(n3435), .ZN(n5249) );
  INV_X1 U4317 ( .A(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n3928) );
  NAND2_X1 U4318 ( .A1(n5629), .A2(n3928), .ZN(n5248) );
  INV_X1 U4319 ( .A(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n3438) );
  AND2_X1 U4320 ( .A1(n5629), .A2(n3438), .ZN(n3441) );
  OAI21_X2 U4321 ( .B1(n6213), .B2(n3441), .A(n3440), .ZN(n5266) );
  INV_X1 U4322 ( .A(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n6254) );
  OR2_X2 U4323 ( .A1(n5266), .A2(n5267), .ZN(n5319) );
  NAND2_X1 U4324 ( .A1(n5629), .A2(n6254), .ZN(n5891) );
  NAND2_X1 U4325 ( .A1(n5629), .A2(n4196), .ZN(n3444) );
  INV_X1 U4326 ( .A(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n5322) );
  AND2_X1 U4327 ( .A1(n5629), .A2(n5322), .ZN(n5672) );
  INV_X1 U4328 ( .A(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n5675) );
  AND2_X1 U4329 ( .A1(n5629), .A2(n5675), .ZN(n5698) );
  NOR2_X1 U4330 ( .A1(n5672), .A2(n5698), .ZN(n5346) );
  INV_X1 U4331 ( .A(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5674) );
  AND2_X1 U4332 ( .A1(n5346), .A2(n3000), .ZN(n3442) );
  INV_X1 U4333 ( .A(n3444), .ZN(n3445) );
  XNOR2_X1 U4334 ( .A(n5629), .B(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n5892)
         );
  OR2_X1 U4335 ( .A1(n5629), .A2(n5322), .ZN(n3446) );
  NOR2_X1 U4336 ( .A1(n5629), .A2(n5675), .ZN(n5699) );
  INV_X1 U4337 ( .A(n5699), .ZN(n3447) );
  NAND2_X1 U4338 ( .A1(n3450), .A2(n3448), .ZN(n5682) );
  INV_X1 U4339 ( .A(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5820) );
  INV_X1 U4340 ( .A(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n5786) );
  NAND2_X1 U4341 ( .A1(n5820), .A2(n5786), .ZN(n3449) );
  OAI21_X1 U4342 ( .B1(n5682), .B2(n3449), .A(n5683), .ZN(n3452) );
  INV_X1 U4343 ( .A(n3450), .ZN(n5669) );
  AND2_X1 U4344 ( .A1(INSTADDRPOINTER_REG_17__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n4201) );
  NAND2_X1 U4345 ( .A1(n5669), .A2(n4201), .ZN(n3451) );
  NAND2_X1 U4346 ( .A1(n3452), .A2(n3451), .ZN(n4222) );
  INV_X1 U4347 ( .A(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5799) );
  NOR2_X1 U4348 ( .A1(n5629), .A2(n5799), .ZN(n5661) );
  NOR2_X2 U4349 ( .A1(n5665), .A2(n5661), .ZN(n5657) );
  INV_X1 U4350 ( .A(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5790) );
  AOI21_X2 U4351 ( .B1(n3454), .B2(n2998), .A(n3005), .ZN(n5649) );
  XNOR2_X1 U4352 ( .A(n5629), .B(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5648)
         );
  NAND2_X1 U4353 ( .A1(n5649), .A2(n5648), .ZN(n5647) );
  INV_X1 U4354 ( .A(n5647), .ZN(n3455) );
  NOR2_X1 U4355 ( .A1(n3437), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5640)
         );
  NAND2_X1 U4356 ( .A1(n3455), .A2(n5640), .ZN(n5632) );
  OAI21_X1 U4357 ( .B1(n5683), .B2(INSTADDRPOINTER_REG_21__SCAN_IN), .A(n5647), 
        .ZN(n5643) );
  NAND3_X1 U4358 ( .A1(n5629), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n3456) );
  XNOR2_X1 U4359 ( .A(n3457), .B(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5386)
         );
  NAND2_X1 U4360 ( .A1(n5031), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3463) );
  OAI21_X1 U4361 ( .B1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n5031), .A(n3463), 
        .ZN(n3465) );
  INV_X1 U4362 ( .A(n3465), .ZN(n3460) );
  INV_X1 U4363 ( .A(n3458), .ZN(n3459) );
  AOI21_X1 U4364 ( .B1(n3140), .B2(n3460), .A(n3459), .ZN(n3469) );
  NAND2_X1 U4365 ( .A1(n4513), .A2(n3157), .ZN(n3462) );
  NAND2_X1 U4366 ( .A1(n4240), .A2(n3462), .ZN(n3483) );
  AOI21_X1 U4367 ( .B1(n3507), .B2(n4181), .A(n3138), .ZN(n3470) );
  INV_X1 U4368 ( .A(n3463), .ZN(n3478) );
  XNOR2_X1 U4369 ( .A(n6464), .B(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3477)
         );
  XNOR2_X1 U4370 ( .A(n3478), .B(n3477), .ZN(n4161) );
  NAND2_X1 U4371 ( .A1(n4161), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3471) );
  NAND2_X1 U4372 ( .A1(n3470), .A2(n3471), .ZN(n3468) );
  INV_X1 U4373 ( .A(n3507), .ZN(n3466) );
  OAI21_X1 U4374 ( .B1(n3466), .B2(n3465), .A(n3511), .ZN(n3467) );
  OAI211_X1 U4375 ( .C1(n3469), .C2(n3483), .A(n3468), .B(n3467), .ZN(n3476)
         );
  INV_X1 U4376 ( .A(n3470), .ZN(n3474) );
  INV_X1 U4377 ( .A(n4161), .ZN(n3473) );
  NAND2_X1 U4378 ( .A1(n3511), .A2(n3471), .ZN(n3472) );
  OAI21_X1 U4379 ( .B1(n3474), .B2(n3473), .A(n3472), .ZN(n3475) );
  NAND2_X1 U4380 ( .A1(n3476), .A2(n3475), .ZN(n3487) );
  INV_X1 U4381 ( .A(n3477), .ZN(n3479) );
  NAND2_X1 U4382 ( .A1(n3479), .A2(n3478), .ZN(n3481) );
  NAND2_X1 U4383 ( .A1(n6464), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3480) );
  NAND2_X1 U4384 ( .A1(n3481), .A2(n3480), .ZN(n3489) );
  XNOR2_X1 U4385 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3488) );
  INV_X1 U4386 ( .A(n3488), .ZN(n3482) );
  XNOR2_X1 U4387 ( .A(n3489), .B(n3482), .ZN(n4163) );
  OAI211_X1 U4388 ( .C1(n3487), .C2(n3483), .A(n4163), .B(n3507), .ZN(n3502)
         );
  INV_X1 U4389 ( .A(n3499), .ZN(n3485) );
  INV_X1 U4390 ( .A(n3483), .ZN(n3484) );
  OAI21_X1 U4391 ( .B1(n4163), .B2(n3485), .A(n3484), .ZN(n3486) );
  NAND2_X1 U4392 ( .A1(n3487), .A2(n3486), .ZN(n3501) );
  NAND2_X1 U4393 ( .A1(n3489), .A2(n3488), .ZN(n3491) );
  NAND2_X1 U4394 ( .A1(n6468), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3490) );
  NAND2_X1 U4395 ( .A1(n3491), .A2(n3490), .ZN(n3496) );
  XNOR2_X1 U4396 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n3494) );
  NAND2_X1 U4397 ( .A1(n3496), .A2(n3494), .ZN(n3493) );
  NAND2_X1 U4398 ( .A1(n6474), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3492) );
  NAND2_X1 U4399 ( .A1(n3493), .A2(n3492), .ZN(n3504) );
  INV_X1 U4400 ( .A(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n6346) );
  INV_X1 U4401 ( .A(n3494), .ZN(n3495) );
  XNOR2_X1 U4402 ( .A(n3496), .B(n3495), .ZN(n3497) );
  NOR2_X1 U4403 ( .A1(n4160), .A2(n3499), .ZN(n3500) );
  AOI21_X1 U4404 ( .B1(n3502), .B2(n3501), .A(n3500), .ZN(n3510) );
  AND2_X1 U4405 ( .A1(n6346), .A2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n3503)
         );
  INV_X1 U4406 ( .A(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n3582) );
  NAND2_X1 U4407 ( .A1(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n3582), .ZN(n3505) );
  AOI22_X1 U4408 ( .A1(n4165), .A2(n3507), .B1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n6498), .ZN(n3508) );
  OAI21_X1 U4409 ( .B1(n3511), .B2(n4160), .A(n3508), .ZN(n3509) );
  INV_X1 U4410 ( .A(n3511), .ZN(n3512) );
  NAND2_X1 U4411 ( .A1(n3515), .A2(STATE2_REG_0__SCAN_IN), .ZN(n6500) );
  NAND2_X1 U4412 ( .A1(n5842), .A2(n4518), .ZN(n3518) );
  NAND2_X1 U4413 ( .A1(n4189), .A2(n3518), .ZN(n4241) );
  OR2_X1 U4414 ( .A1(n4241), .A2(n3140), .ZN(n6479) );
  AOI22_X1 U4415 ( .A1(n3853), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n4116), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3522) );
  AOI22_X1 U4416 ( .A1(n4021), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n4063), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3521) );
  AOI22_X1 U4417 ( .A1(n2994), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n4118), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3520) );
  AOI22_X1 U4418 ( .A1(n4127), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n3232), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3519) );
  NAND4_X1 U4419 ( .A1(n3522), .A2(n3521), .A3(n3520), .A4(n3519), .ZN(n3528)
         );
  AOI22_X1 U4420 ( .A1(n4117), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n4125), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3526) );
  AOI22_X1 U4421 ( .A1(n4119), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n4126), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3525) );
  AOI22_X1 U4422 ( .A1(n2992), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n4022), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3524) );
  AOI22_X1 U4423 ( .A1(n4120), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n4027), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3523) );
  NAND4_X1 U4424 ( .A1(n3526), .A2(n3525), .A3(n3524), .A4(n3523), .ZN(n3527)
         );
  NOR2_X1 U4425 ( .A1(n3528), .A2(n3527), .ZN(n3870) );
  AOI22_X1 U4426 ( .A1(n4116), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n4117), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n3532) );
  AOI22_X1 U4427 ( .A1(n2994), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n4119), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n3531) );
  AOI22_X1 U4428 ( .A1(n4125), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .B1(n4022), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3530) );
  AOI22_X1 U4429 ( .A1(n4120), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n4027), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3529) );
  NAND4_X1 U4430 ( .A1(n3532), .A2(n3531), .A3(n3530), .A4(n3529), .ZN(n3538)
         );
  AOI22_X1 U4431 ( .A1(n3853), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n4021), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3536) );
  AOI22_X1 U4432 ( .A1(n4063), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n2992), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n3535) );
  AOI22_X1 U4433 ( .A1(n4126), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n4118), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3534) );
  AOI22_X1 U4434 ( .A1(n4127), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3232), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3533) );
  NAND4_X1 U4435 ( .A1(n3536), .A2(n3535), .A3(n3534), .A4(n3533), .ZN(n3537)
         );
  NOR2_X1 U4436 ( .A1(n3538), .A2(n3537), .ZN(n3869) );
  NOR2_X1 U4437 ( .A1(n3870), .A2(n3869), .ZN(n4035) );
  AOI22_X1 U4438 ( .A1(n3853), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n4116), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3542) );
  AOI22_X1 U4439 ( .A1(n4117), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n4021), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3541) );
  AOI22_X1 U4440 ( .A1(n4063), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n3254), 
        .B2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3540) );
  AOI22_X1 U4441 ( .A1(n4125), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n4022), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3539) );
  NAND4_X1 U4442 ( .A1(n3542), .A2(n3541), .A3(n3540), .A4(n3539), .ZN(n3548)
         );
  AOI22_X1 U4443 ( .A1(INSTQUEUE_REG_6__1__SCAN_IN), .A2(n2994), .B1(n4119), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3546) );
  AOI22_X1 U4444 ( .A1(n4127), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n3232), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3545) );
  AOI22_X1 U4445 ( .A1(INSTQUEUE_REG_8__1__SCAN_IN), .A2(n4120), .B1(n4027), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3544) );
  AOI22_X1 U4446 ( .A1(n4126), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n4118), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3543) );
  NAND4_X1 U4447 ( .A1(n3546), .A2(n3545), .A3(n3544), .A4(n3543), .ZN(n3547)
         );
  OR2_X1 U4448 ( .A1(n3548), .A2(n3547), .ZN(n4034) );
  INV_X1 U4449 ( .A(n4034), .ZN(n3549) );
  XNOR2_X1 U4450 ( .A(n4035), .B(n3549), .ZN(n3553) );
  INV_X1 U4451 ( .A(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n5967) );
  INV_X1 U4452 ( .A(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n3789) );
  INV_X1 U4453 ( .A(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n3827) );
  INV_X1 U4454 ( .A(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n5650) );
  XNOR2_X1 U4455 ( .A(n4038), .B(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n5494)
         );
  INV_X2 U4456 ( .A(STATE2_REG_2__SCAN_IN), .ZN(n6497) );
  NAND2_X1 U4457 ( .A1(n6497), .A2(STATEBS16_REG_SCAN_IN), .ZN(n3692) );
  INV_X1 U4458 ( .A(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n5490) );
  NOR2_X1 U4459 ( .A1(n3692), .A2(n5490), .ZN(n3550) );
  AOI21_X1 U4460 ( .B1(n4094), .B2(EAX_REG_24__SCAN_IN), .A(n3550), .ZN(n3551)
         );
  OAI21_X1 U4461 ( .B1(n5494), .B2(n4139), .A(n3551), .ZN(n3552) );
  AOI21_X1 U4462 ( .B1(n3553), .B2(n4111), .A(n3552), .ZN(n4017) );
  NOR2_X2 U4463 ( .A1(n3554), .A2(n6497), .ZN(n3733) );
  NAND2_X1 U4464 ( .A1(n4483), .A2(n3733), .ZN(n3558) );
  AOI22_X1 U4465 ( .A1(n3560), .A2(EAX_REG_1__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n6497), .ZN(n3556) );
  AND2_X1 U4466 ( .A1(n4398), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3577) );
  NAND2_X1 U4467 ( .A1(n3577), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3555) );
  AND2_X1 U4468 ( .A1(n3556), .A2(n3555), .ZN(n3557) );
  NAND2_X1 U4469 ( .A1(n3558), .A2(n3557), .ZN(n4401) );
  INV_X1 U4470 ( .A(n3577), .ZN(n3583) );
  NAND2_X1 U4471 ( .A1(n5412), .A2(n3733), .ZN(n3562) );
  AOI22_X1 U4472 ( .A1(n3560), .A2(EAX_REG_0__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n6497), .ZN(n3561) );
  OAI211_X1 U4473 ( .C1(n3583), .C2(n3153), .A(n3562), .B(n3561), .ZN(n4369)
         );
  MUX2_X1 U4474 ( .A(n4256), .B(n4370), .S(n4369), .Z(n4402) );
  NAND2_X1 U4475 ( .A1(n4401), .A2(n4402), .ZN(n4400) );
  NAND2_X1 U4476 ( .A1(n3577), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3568) );
  INV_X1 U4477 ( .A(PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n3565) );
  OAI21_X1 U4478 ( .B1(PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .A(n3563), .ZN(n6248) );
  NAND2_X1 U4479 ( .A1(n4256), .A2(n6248), .ZN(n3564) );
  OAI21_X1 U4480 ( .B1(n3565), .B2(n3692), .A(n3564), .ZN(n3566) );
  AOI21_X1 U4481 ( .B1(n3560), .B2(EAX_REG_2__SCAN_IN), .A(n3566), .ZN(n3567)
         );
  AND2_X1 U4482 ( .A1(n3568), .A2(n3567), .ZN(n4571) );
  NOR2_X1 U4483 ( .A1(n4400), .A2(n4571), .ZN(n3571) );
  INV_X1 U4484 ( .A(n3733), .ZN(n3622) );
  NAND2_X1 U4485 ( .A1(n4400), .A2(n4571), .ZN(n3570) );
  OAI21_X1 U4486 ( .B1(n3571), .B2(n4573), .A(n3570), .ZN(n3572) );
  INV_X1 U4487 ( .A(n3572), .ZN(n4526) );
  NOR2_X1 U4488 ( .A1(PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n3574), .ZN(n3575)
         );
  NOR2_X1 U4489 ( .A1(n3585), .A2(n3575), .ZN(n6055) );
  INV_X1 U4490 ( .A(PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n4544) );
  OAI22_X1 U4491 ( .A1(n6055), .A2(n4139), .B1(n3692), .B2(n4544), .ZN(n3576)
         );
  AOI21_X1 U4492 ( .B1(n4094), .B2(EAX_REG_3__SCAN_IN), .A(n3576), .ZN(n3579)
         );
  NAND2_X1 U4493 ( .A1(n3577), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3578) );
  OAI211_X1 U4494 ( .C1(n2995), .C2(n3622), .A(n3579), .B(n3578), .ZN(n4528)
         );
  NAND2_X1 U4495 ( .A1(n4526), .A2(n4528), .ZN(n4562) );
  NAND2_X1 U4496 ( .A1(n6497), .A2(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n3581)
         );
  NAND2_X1 U4497 ( .A1(n4094), .A2(EAX_REG_4__SCAN_IN), .ZN(n3580) );
  OAI211_X1 U4498 ( .C1(n3583), .C2(n3582), .A(n3581), .B(n3580), .ZN(n3584)
         );
  NAND2_X1 U4499 ( .A1(n3584), .A2(n4139), .ZN(n3587) );
  OAI21_X1 U4500 ( .B1(n3585), .B2(PHYADDRPOINTER_REG_4__SCAN_IN), .A(n3591), 
        .ZN(n6238) );
  NAND2_X1 U4501 ( .A1(n6238), .A2(n4256), .ZN(n3586) );
  NAND2_X1 U4502 ( .A1(n3587), .A2(n3586), .ZN(n3588) );
  AOI21_X1 U4503 ( .B1(n3589), .B2(n3733), .A(n3588), .ZN(n4561) );
  NAND2_X1 U4504 ( .A1(n3590), .A2(n3733), .ZN(n3594) );
  XNOR2_X1 U4505 ( .A(n3591), .B(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n5209) );
  OAI22_X1 U4506 ( .A1(n5209), .A2(n4139), .B1(n3692), .B2(n4846), .ZN(n3592)
         );
  AOI21_X1 U4507 ( .B1(n4094), .B2(EAX_REG_5__SCAN_IN), .A(n3592), .ZN(n3593)
         );
  NAND2_X1 U4508 ( .A1(n3594), .A2(n3593), .ZN(n4584) );
  NAND2_X1 U4509 ( .A1(n4563), .A2(n4584), .ZN(n4583) );
  INV_X1 U4510 ( .A(n4583), .ZN(n3602) );
  NOR2_X1 U4511 ( .A1(n3595), .A2(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n3596)
         );
  OR2_X1 U4512 ( .A1(n3603), .A2(n3596), .ZN(n6229) );
  INV_X1 U4513 ( .A(EAX_REG_6__SCAN_IN), .ZN(n6181) );
  INV_X1 U4514 ( .A(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n3597) );
  OAI22_X1 U4515 ( .A1(n3756), .A2(n6181), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n3597), .ZN(n3598) );
  MUX2_X1 U4516 ( .A(n6229), .B(n3598), .S(n4139), .Z(n3599) );
  NAND2_X1 U4517 ( .A1(n3602), .A2(n3601), .ZN(n4788) );
  INV_X1 U4518 ( .A(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n5078) );
  NAND2_X1 U4519 ( .A1(n4094), .A2(EAX_REG_7__SCAN_IN), .ZN(n3605) );
  XNOR2_X1 U4520 ( .A(n3603), .B(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n5084) );
  NAND2_X1 U4521 ( .A1(n5084), .A2(n3811), .ZN(n3604) );
  OAI211_X1 U4522 ( .C1(n5078), .C2(n3692), .A(n3605), .B(n3604), .ZN(n3606)
         );
  NOR2_X2 U4523 ( .A1(n4788), .A2(n4851), .ZN(n4910) );
  AOI22_X1 U4524 ( .A1(n3853), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n4116), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3612) );
  AOI22_X1 U4525 ( .A1(n4117), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n4021), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3611) );
  AOI22_X1 U4526 ( .A1(n4119), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n3254), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3610) );
  AOI22_X1 U4527 ( .A1(n3232), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n4118), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3609) );
  NAND4_X1 U4528 ( .A1(n3612), .A2(n3611), .A3(n3610), .A4(n3609), .ZN(n3618)
         );
  AOI22_X1 U4529 ( .A1(n4063), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n2994), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3616) );
  AOI22_X1 U4530 ( .A1(n3675), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n4126), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3615) );
  AOI22_X1 U4531 ( .A1(n4125), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n4022), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3614) );
  AOI22_X1 U4532 ( .A1(n4120), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n4027), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3613) );
  NAND4_X1 U4533 ( .A1(n3616), .A2(n3615), .A3(n3614), .A4(n3613), .ZN(n3617)
         );
  NOR2_X1 U4534 ( .A1(n3618), .A2(n3617), .ZN(n3623) );
  XNOR2_X1 U4535 ( .A(n3619), .B(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n5272)
         );
  NAND2_X1 U4536 ( .A1(n5272), .A2(n3811), .ZN(n3621) );
  INV_X1 U4537 ( .A(n3692), .ZN(n4273) );
  AOI22_X1 U4538 ( .A1(n3560), .A2(EAX_REG_12__SCAN_IN), .B1(n4273), .B2(
        PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n3620) );
  OAI211_X1 U4539 ( .C1(n3623), .C2(n3622), .A(n3621), .B(n3620), .ZN(n5216)
         );
  XOR2_X1 U4540 ( .A(n6002), .B(n3624), .Z(n6216) );
  INV_X1 U4541 ( .A(n6216), .ZN(n3639) );
  AOI22_X1 U4542 ( .A1(n3853), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n4021), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3628) );
  AOI22_X1 U4543 ( .A1(n3675), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n4119), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n3627) );
  AOI22_X1 U4544 ( .A1(n4063), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n2992), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n3626) );
  AOI22_X1 U4545 ( .A1(n4120), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3232), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3625) );
  NAND4_X1 U4546 ( .A1(n3628), .A2(n3627), .A3(n3626), .A4(n3625), .ZN(n3634)
         );
  AOI22_X1 U4547 ( .A1(n4116), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n4117), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3632) );
  AOI22_X1 U4548 ( .A1(n4125), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n4022), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3631) );
  AOI22_X1 U4549 ( .A1(n4126), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .B1(n4027), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3630) );
  AOI22_X1 U4550 ( .A1(n2994), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n4118), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3629) );
  NAND4_X1 U4551 ( .A1(n3632), .A2(n3631), .A3(n3630), .A4(n3629), .ZN(n3633)
         );
  OAI21_X1 U4552 ( .B1(n3634), .B2(n3633), .A(n3733), .ZN(n3637) );
  NAND2_X1 U4553 ( .A1(n4094), .A2(EAX_REG_11__SCAN_IN), .ZN(n3636) );
  NAND2_X1 U4554 ( .A1(n4273), .A2(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n3635)
         );
  NAND3_X1 U4555 ( .A1(n3637), .A2(n3636), .A3(n3635), .ZN(n3638) );
  AOI21_X1 U4556 ( .B1(n3639), .B2(n3811), .A(n3638), .ZN(n5277) );
  XNOR2_X1 U4557 ( .A(n3640), .B(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n5528)
         );
  AOI22_X1 U4558 ( .A1(n4116), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n4117), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3644) );
  AOI22_X1 U4559 ( .A1(n4063), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n2992), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3643) );
  AOI22_X1 U4560 ( .A1(n2994), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n4119), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n3642) );
  AOI22_X1 U4561 ( .A1(n4126), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .B1(n4120), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3641) );
  NAND4_X1 U4562 ( .A1(n3644), .A2(n3643), .A3(n3642), .A4(n3641), .ZN(n3650)
         );
  AOI22_X1 U4563 ( .A1(n3853), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n4021), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3648) );
  AOI22_X1 U4564 ( .A1(n4125), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n4022), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3647) );
  AOI22_X1 U4565 ( .A1(n3232), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n4027), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3646) );
  AOI22_X1 U4566 ( .A1(n3675), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n4118), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3645) );
  NAND4_X1 U4567 ( .A1(n3648), .A2(n3647), .A3(n3646), .A4(n3645), .ZN(n3649)
         );
  OAI21_X1 U4568 ( .B1(n3650), .B2(n3649), .A(n3733), .ZN(n3653) );
  NAND2_X1 U4569 ( .A1(n4094), .A2(EAX_REG_10__SCAN_IN), .ZN(n3652) );
  NAND2_X1 U4570 ( .A1(n4273), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n3651)
         );
  NAND3_X1 U4571 ( .A1(n3653), .A2(n3652), .A3(n3651), .ZN(n3654) );
  AOI21_X1 U4572 ( .B1(n5528), .B2(n3811), .A(n3654), .ZN(n5224) );
  NOR2_X1 U4573 ( .A1(n5277), .A2(n5224), .ZN(n5214) );
  NAND2_X1 U4574 ( .A1(n5216), .A2(n5214), .ZN(n3670) );
  XOR2_X1 U4575 ( .A(n6011), .B(n3655), .Z(n6015) );
  INV_X1 U4576 ( .A(n6015), .ZN(n5187) );
  AOI22_X1 U4577 ( .A1(n3853), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n4021), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3659) );
  AOI22_X1 U4578 ( .A1(n3675), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n4126), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3658) );
  AOI22_X1 U4579 ( .A1(n4125), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n4022), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3657) );
  AOI22_X1 U4580 ( .A1(INSTQUEUE_REG_6__1__SCAN_IN), .A2(n4120), .B1(n4027), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3656) );
  NAND4_X1 U4581 ( .A1(n3659), .A2(n3658), .A3(n3657), .A4(n3656), .ZN(n3665)
         );
  AOI22_X1 U4582 ( .A1(n4116), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n4117), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3663) );
  AOI22_X1 U4583 ( .A1(n2994), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n4119), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3662) );
  AOI22_X1 U4584 ( .A1(INSTQUEUE_REG_13__1__SCAN_IN), .A2(n4063), .B1(n2992), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3661) );
  AOI22_X1 U4585 ( .A1(n3232), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n4118), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3660) );
  NAND4_X1 U4586 ( .A1(n3663), .A2(n3662), .A3(n3661), .A4(n3660), .ZN(n3664)
         );
  OAI21_X1 U4587 ( .B1(n3665), .B2(n3664), .A(n3733), .ZN(n3668) );
  NAND2_X1 U4588 ( .A1(n4094), .A2(EAX_REG_9__SCAN_IN), .ZN(n3667) );
  NAND2_X1 U4589 ( .A1(n4273), .A2(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n3666)
         );
  NAND3_X1 U4590 ( .A1(n3668), .A2(n3667), .A3(n3666), .ZN(n3669) );
  AOI21_X1 U4591 ( .B1(n5187), .B2(n3811), .A(n3669), .ZN(n5212) );
  NOR2_X1 U4592 ( .A1(n3670), .A2(n5212), .ZN(n3687) );
  AOI22_X1 U4593 ( .A1(n3853), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n4117), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3674) );
  AOI22_X1 U4594 ( .A1(n2994), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n4119), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3673) );
  AOI22_X1 U4595 ( .A1(n4125), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n2992), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3672) );
  AOI22_X1 U4596 ( .A1(n4027), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n4118), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3671) );
  NAND4_X1 U4597 ( .A1(n3674), .A2(n3673), .A3(n3672), .A4(n3671), .ZN(n3681)
         );
  AOI22_X1 U4598 ( .A1(n4116), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n4021), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3679) );
  AOI22_X1 U4599 ( .A1(n3675), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n4126), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3678) );
  AOI22_X1 U4600 ( .A1(n4063), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n4022), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3677) );
  AOI22_X1 U4601 ( .A1(n4120), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n3232), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3676) );
  NAND4_X1 U4602 ( .A1(n3679), .A2(n3678), .A3(n3677), .A4(n3676), .ZN(n3680)
         );
  OAI21_X1 U4603 ( .B1(n3681), .B2(n3680), .A(n3733), .ZN(n3686) );
  NAND2_X1 U4604 ( .A1(n4094), .A2(EAX_REG_8__SCAN_IN), .ZN(n3685) );
  INV_X1 U4605 ( .A(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n4972) );
  XNOR2_X1 U4606 ( .A(n3682), .B(n4972), .ZN(n6027) );
  OR2_X1 U4607 ( .A1(n6027), .A2(n4139), .ZN(n3684) );
  NAND2_X1 U4608 ( .A1(n4273), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n3683)
         );
  NAND4_X1 U4609 ( .A1(n3686), .A2(n3685), .A3(n3684), .A4(n3683), .ZN(n4912)
         );
  AND2_X1 U4610 ( .A1(n3687), .A2(n4912), .ZN(n3688) );
  NAND2_X1 U4611 ( .A1(n4910), .A2(n3688), .ZN(n3696) );
  INV_X1 U4612 ( .A(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n3693) );
  OAI21_X1 U4613 ( .B1(PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n3690), .A(n3689), 
        .ZN(n5995) );
  NAND2_X1 U4614 ( .A1(n5995), .A2(n3811), .ZN(n3691) );
  OAI21_X1 U4615 ( .B1(n3693), .B2(n3692), .A(n3691), .ZN(n3694) );
  AOI21_X1 U4616 ( .B1(n4094), .B2(EAX_REG_13__SCAN_IN), .A(n3694), .ZN(n3695)
         );
  NAND2_X1 U4617 ( .A1(n3696), .A2(n3695), .ZN(n3697) );
  AOI22_X1 U4618 ( .A1(n4116), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n4117), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3701) );
  AOI22_X1 U4619 ( .A1(n4063), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n2994), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3700) );
  AOI22_X1 U4620 ( .A1(n3675), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n4126), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3699) );
  AOI22_X1 U4621 ( .A1(n3232), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n4027), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3698) );
  NAND4_X1 U4622 ( .A1(n3701), .A2(n3700), .A3(n3699), .A4(n3698), .ZN(n3707)
         );
  AOI22_X1 U4623 ( .A1(n3853), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n4021), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3705) );
  AOI22_X1 U4624 ( .A1(n4119), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3254), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3704) );
  AOI22_X1 U4625 ( .A1(n4125), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n4022), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3703) );
  AOI22_X1 U4626 ( .A1(n4120), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n4118), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3702) );
  NAND4_X1 U4627 ( .A1(n3705), .A2(n3704), .A3(n3703), .A4(n3702), .ZN(n3706)
         );
  OR2_X1 U4628 ( .A1(n3707), .A2(n3706), .ZN(n3708) );
  AND2_X1 U4629 ( .A1(n3733), .A2(n3708), .ZN(n5242) );
  XOR2_X1 U4630 ( .A(PHYADDRPOINTER_REG_14__SCAN_IN), .B(n3710), .Z(n5983) );
  AOI22_X1 U4631 ( .A1(n3853), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n4116), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3714) );
  AOI22_X1 U4632 ( .A1(n4021), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n4125), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3713) );
  AOI22_X1 U4633 ( .A1(n4063), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n4022), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3712) );
  AOI22_X1 U4634 ( .A1(n2994), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n3232), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3711) );
  NAND4_X1 U4635 ( .A1(n3714), .A2(n3713), .A3(n3712), .A4(n3711), .ZN(n3720)
         );
  AOI22_X1 U4636 ( .A1(n3675), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n4126), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3718) );
  AOI22_X1 U4637 ( .A1(n4117), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n2992), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n3717) );
  AOI22_X1 U4638 ( .A1(n4119), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n4118), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3716) );
  AOI22_X1 U4639 ( .A1(n4120), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n4027), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3715) );
  NAND4_X1 U4640 ( .A1(n3718), .A2(n3717), .A3(n3716), .A4(n3715), .ZN(n3719)
         );
  OR2_X1 U4641 ( .A1(n3720), .A2(n3719), .ZN(n3721) );
  AOI22_X1 U4642 ( .A1(n3733), .A2(n3721), .B1(n4273), .B2(
        PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n3723) );
  NAND2_X1 U4643 ( .A1(n3560), .A2(EAX_REG_14__SCAN_IN), .ZN(n3722) );
  OAI211_X1 U4644 ( .C1(n5983), .C2(n4139), .A(n3723), .B(n3722), .ZN(n5257)
         );
  NAND2_X1 U4645 ( .A1(n5258), .A2(n5257), .ZN(n5256) );
  INV_X1 U4646 ( .A(n5256), .ZN(n3741) );
  XNOR2_X1 U4647 ( .A(n3724), .B(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n5974)
         );
  INV_X1 U4648 ( .A(n5974), .ZN(n5703) );
  AOI22_X1 U4649 ( .A1(n3853), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n4117), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3728) );
  AOI22_X1 U4650 ( .A1(n4119), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n2992), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n3727) );
  AOI22_X1 U4651 ( .A1(n4125), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n4022), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3726) );
  AOI22_X1 U4652 ( .A1(n4126), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n3232), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3725) );
  NAND4_X1 U4653 ( .A1(n3728), .A2(n3727), .A3(n3726), .A4(n3725), .ZN(n3735)
         );
  AOI22_X1 U4654 ( .A1(n4116), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n4021), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3732) );
  AOI22_X1 U4655 ( .A1(n4063), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n2994), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3731) );
  AOI22_X1 U4656 ( .A1(n3675), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n4118), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3730) );
  AOI22_X1 U4657 ( .A1(n4120), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n4027), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3729) );
  NAND4_X1 U4658 ( .A1(n3732), .A2(n3731), .A3(n3730), .A4(n3729), .ZN(n3734)
         );
  OAI21_X1 U4659 ( .B1(n3735), .B2(n3734), .A(n3733), .ZN(n3738) );
  NAND2_X1 U4660 ( .A1(n4094), .A2(EAX_REG_15__SCAN_IN), .ZN(n3737) );
  NAND2_X1 U4661 ( .A1(n4273), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n3736)
         );
  NAND3_X1 U4662 ( .A1(n3738), .A2(n3737), .A3(n3736), .ZN(n3739) );
  AOI21_X1 U4663 ( .B1(n5703), .B2(n3811), .A(n3739), .ZN(n5300) );
  NAND2_X1 U4664 ( .A1(n3741), .A2(n3740), .ZN(n5298) );
  AOI22_X1 U4665 ( .A1(n4116), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n4021), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3745) );
  AOI22_X1 U4666 ( .A1(n4063), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n2992), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3744) );
  AOI22_X1 U4667 ( .A1(n4119), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n4120), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3743) );
  AOI22_X1 U4668 ( .A1(n4125), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .B1(n4022), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3742) );
  NAND4_X1 U4669 ( .A1(n3745), .A2(n3744), .A3(n3743), .A4(n3742), .ZN(n3751)
         );
  AOI22_X1 U4670 ( .A1(n3853), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n4117), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3749) );
  AOI22_X1 U4671 ( .A1(n3675), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n4126), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3748) );
  AOI22_X1 U4672 ( .A1(n2994), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n4118), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3747) );
  AOI22_X1 U4673 ( .A1(n3232), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n4027), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3746) );
  NAND4_X1 U4674 ( .A1(n3749), .A2(n3748), .A3(n3747), .A4(n3746), .ZN(n3750)
         );
  OR2_X1 U4675 ( .A1(n3751), .A2(n3750), .ZN(n3758) );
  INV_X1 U4676 ( .A(EAX_REG_16__SCAN_IN), .ZN(n3755) );
  XOR2_X1 U4677 ( .A(PHYADDRPOINTER_REG_16__SCAN_IN), .B(n3752), .Z(n5962) );
  INV_X1 U4678 ( .A(n5962), .ZN(n3753) );
  AOI22_X1 U4679 ( .A1(PHYADDRPOINTER_REG_16__SCAN_IN), .A2(n4273), .B1(n4256), 
        .B2(n3753), .ZN(n3754) );
  OAI21_X1 U4680 ( .B1(n3756), .B2(n3755), .A(n3754), .ZN(n3757) );
  AOI21_X1 U4681 ( .B1(n4111), .B2(n3758), .A(n3757), .ZN(n5310) );
  NOR2_X2 U4682 ( .A1(n5298), .A2(n5310), .ZN(n5282) );
  AOI22_X1 U4683 ( .A1(n3853), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n4116), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3762) );
  AOI22_X1 U4684 ( .A1(INSTQUEUE_REG_14__1__SCAN_IN), .A2(n4063), .B1(n2992), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3761) );
  AOI22_X1 U4685 ( .A1(n4126), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n3832), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3760) );
  AOI22_X1 U4686 ( .A1(n2994), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n4118), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3759) );
  NAND4_X1 U4687 ( .A1(n3762), .A2(n3761), .A3(n3760), .A4(n3759), .ZN(n3768)
         );
  AOI22_X1 U4688 ( .A1(INSTQUEUE_REG_9__1__SCAN_IN), .A2(n4117), .B1(n4021), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3766) );
  AOI22_X1 U4689 ( .A1(INSTQUEUE_REG_13__1__SCAN_IN), .A2(n3675), .B1(n4119), 
        .B2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3765) );
  AOI22_X1 U4690 ( .A1(INSTQUEUE_REG_0__1__SCAN_IN), .A2(n4125), .B1(n4022), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3764) );
  AOI22_X1 U4691 ( .A1(INSTQUEUE_REG_6__1__SCAN_IN), .A2(n3232), .B1(n4027), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3763) );
  NAND4_X1 U4692 ( .A1(n3766), .A2(n3765), .A3(n3764), .A4(n3763), .ZN(n3767)
         );
  NOR2_X1 U4693 ( .A1(n3768), .A2(n3767), .ZN(n3771) );
  INV_X1 U4694 ( .A(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n5690) );
  OAI21_X1 U4695 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n5690), .A(n4139), .ZN(
        n3769) );
  AOI21_X1 U4696 ( .B1(n4094), .B2(EAX_REG_17__SCAN_IN), .A(n3769), .ZN(n3770)
         );
  OAI21_X1 U4697 ( .B1(n4142), .B2(n3771), .A(n3770), .ZN(n3774) );
  XNOR2_X1 U4698 ( .A(n3772), .B(n5690), .ZN(n5693) );
  NAND2_X1 U4699 ( .A1(n5693), .A2(n3811), .ZN(n3773) );
  NAND2_X1 U4700 ( .A1(n5282), .A2(n5285), .ZN(n5284) );
  AOI22_X1 U4701 ( .A1(n4116), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n4117), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3778) );
  AOI22_X1 U4702 ( .A1(n4063), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n4119), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n3777) );
  AOI22_X1 U4703 ( .A1(n2994), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n4126), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3776) );
  AOI22_X1 U4704 ( .A1(n3232), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n4027), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3775) );
  NAND4_X1 U4705 ( .A1(n3778), .A2(n3777), .A3(n3776), .A4(n3775), .ZN(n3784)
         );
  AOI22_X1 U4706 ( .A1(n3853), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n4021), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3782) );
  AOI22_X1 U4707 ( .A1(n3675), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n3832), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3781) );
  AOI22_X1 U4708 ( .A1(n4125), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n4022), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3780) );
  AOI22_X1 U4709 ( .A1(n2992), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n4118), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3779) );
  NAND4_X1 U4710 ( .A1(n3782), .A2(n3781), .A3(n3780), .A4(n3779), .ZN(n3783)
         );
  NOR2_X1 U4711 ( .A1(n3784), .A2(n3783), .ZN(n3788) );
  INV_X1 U4712 ( .A(STATEBS16_REG_SCAN_IN), .ZN(n6657) );
  OAI21_X1 U4713 ( .B1(PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n6657), .A(n6497), 
        .ZN(n3785) );
  INV_X1 U4714 ( .A(n3785), .ZN(n3786) );
  AOI21_X1 U4715 ( .B1(n4094), .B2(EAX_REG_18__SCAN_IN), .A(n3786), .ZN(n3787)
         );
  OAI21_X1 U4716 ( .B1(n4142), .B2(n3788), .A(n3787), .ZN(n3794) );
  AND2_X1 U4717 ( .A1(n3790), .A2(n3789), .ZN(n3791) );
  OR2_X1 U4718 ( .A1(n3791), .A2(n3810), .ZN(n5952) );
  INV_X1 U4719 ( .A(n5952), .ZN(n3792) );
  NAND2_X1 U4720 ( .A1(n3792), .A2(n3811), .ZN(n3793) );
  NAND2_X1 U4721 ( .A1(n3794), .A2(n3793), .ZN(n5571) );
  AOI22_X1 U4722 ( .A1(n3853), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n4116), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3800) );
  AOI22_X1 U4723 ( .A1(n4117), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n4021), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3799) );
  AOI22_X1 U4724 ( .A1(n4063), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n2992), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n3798) );
  AOI22_X1 U4725 ( .A1(n4125), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n4022), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3797) );
  NAND4_X1 U4726 ( .A1(n3800), .A2(n3799), .A3(n3798), .A4(n3797), .ZN(n3806)
         );
  AOI22_X1 U4727 ( .A1(n2994), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n4119), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n3804) );
  AOI22_X1 U4728 ( .A1(n3675), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3232), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3803) );
  AOI22_X1 U4729 ( .A1(n4120), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n4027), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3802) );
  AOI22_X1 U4730 ( .A1(n4126), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n4118), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3801) );
  NAND4_X1 U4731 ( .A1(n3804), .A2(n3803), .A3(n3802), .A4(n3801), .ZN(n3805)
         );
  NOR2_X1 U4732 ( .A1(n3806), .A2(n3805), .ZN(n3809) );
  INV_X1 U4733 ( .A(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n5869) );
  AOI21_X1 U4734 ( .B1(n5869), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n3807) );
  AOI21_X1 U4735 ( .B1(n4094), .B2(EAX_REG_19__SCAN_IN), .A(n3807), .ZN(n3808)
         );
  OAI21_X1 U4736 ( .B1(n4142), .B2(n3809), .A(n3808), .ZN(n3813) );
  XNOR2_X1 U4737 ( .A(n3810), .B(n5869), .ZN(n5873) );
  NAND2_X1 U4738 ( .A1(n5873), .A2(n3811), .ZN(n3812) );
  NAND2_X1 U4739 ( .A1(n3813), .A2(n3812), .ZN(n5371) );
  NOR2_X2 U4740 ( .A1(n5370), .A2(n5371), .ZN(n5372) );
  AOI22_X1 U4741 ( .A1(n4117), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n4021), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3817) );
  AOI22_X1 U4742 ( .A1(n4119), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n4126), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3816) );
  AOI22_X1 U4743 ( .A1(n2992), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n4022), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3815) );
  AOI22_X1 U4744 ( .A1(n4120), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n4027), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3814) );
  NAND4_X1 U4745 ( .A1(n3817), .A2(n3816), .A3(n3815), .A4(n3814), .ZN(n3823)
         );
  AOI22_X1 U4746 ( .A1(n3853), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n4116), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3821) );
  AOI22_X1 U4747 ( .A1(n4125), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .B1(n4063), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3820) );
  AOI22_X1 U4748 ( .A1(n2994), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n4118), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3819) );
  AOI22_X1 U4749 ( .A1(n3675), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n3232), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3818) );
  NAND4_X1 U4750 ( .A1(n3821), .A2(n3820), .A3(n3819), .A4(n3818), .ZN(n3822)
         );
  NOR2_X1 U4751 ( .A1(n3823), .A2(n3822), .ZN(n3826) );
  OAI21_X1 U4752 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n3827), .A(n4139), .ZN(
        n3824) );
  AOI21_X1 U4753 ( .B1(n4094), .B2(EAX_REG_20__SCAN_IN), .A(n3824), .ZN(n3825)
         );
  OAI21_X1 U4754 ( .B1(n4142), .B2(n3826), .A(n3825), .ZN(n3831) );
  NAND2_X1 U4755 ( .A1(n3828), .A2(n3827), .ZN(n3829) );
  NAND2_X1 U4756 ( .A1(n3846), .A2(n3829), .ZN(n5866) );
  AND2_X2 U4757 ( .A1(n5372), .A2(n5557), .ZN(n5511) );
  AOI22_X1 U4758 ( .A1(n3853), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n4117), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3836) );
  AOI22_X1 U4759 ( .A1(n4125), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .B1(n4063), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3835) );
  AOI22_X1 U4760 ( .A1(n3675), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n3832), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3834) );
  AOI22_X1 U4761 ( .A1(n3254), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n4118), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3833) );
  NAND4_X1 U4762 ( .A1(n3836), .A2(n3835), .A3(n3834), .A4(n3833), .ZN(n3842)
         );
  AOI22_X1 U4763 ( .A1(n4116), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n4021), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3840) );
  AOI22_X1 U4764 ( .A1(n2994), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n4126), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3839) );
  AOI22_X1 U4765 ( .A1(n4119), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n4022), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3838) );
  AOI22_X1 U4766 ( .A1(n3324), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n4027), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3837) );
  NAND4_X1 U4767 ( .A1(n3840), .A2(n3839), .A3(n3838), .A4(n3837), .ZN(n3841)
         );
  NOR2_X1 U4768 ( .A1(n3842), .A2(n3841), .ZN(n3845) );
  OAI21_X1 U4769 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n5650), .A(n4139), .ZN(
        n3843) );
  AOI21_X1 U4770 ( .B1(n4094), .B2(EAX_REG_21__SCAN_IN), .A(n3843), .ZN(n3844)
         );
  OAI21_X1 U4771 ( .B1(n4142), .B2(n3845), .A(n3844), .ZN(n3848) );
  XNOR2_X1 U4772 ( .A(n3846), .B(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n5652)
         );
  NAND2_X1 U4773 ( .A1(n5652), .A2(n4256), .ZN(n3847) );
  AOI22_X1 U4774 ( .A1(n4116), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n4117), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n3852) );
  AOI22_X1 U4775 ( .A1(n3191), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n2994), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3851) );
  AOI22_X1 U4776 ( .A1(n4125), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n4022), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3850) );
  AOI22_X1 U4777 ( .A1(n4120), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n3232), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3849) );
  NAND4_X1 U4778 ( .A1(n3852), .A2(n3851), .A3(n3850), .A4(n3849), .ZN(n3859)
         );
  AOI22_X1 U4779 ( .A1(n3853), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n4021), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3857) );
  AOI22_X1 U4780 ( .A1(n4119), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3254), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n3856) );
  AOI22_X1 U4781 ( .A1(n4126), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n4118), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3855) );
  AOI22_X1 U4782 ( .A1(n4127), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n4027), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3854) );
  NAND4_X1 U4783 ( .A1(n3857), .A2(n3856), .A3(n3855), .A4(n3854), .ZN(n3858)
         );
  NOR2_X1 U4784 ( .A1(n3859), .A2(n3858), .ZN(n3863) );
  NAND2_X1 U4785 ( .A1(n6497), .A2(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n3860)
         );
  NAND2_X1 U4786 ( .A1(n4139), .A2(n3860), .ZN(n3861) );
  AOI21_X1 U4787 ( .B1(n4094), .B2(EAX_REG_22__SCAN_IN), .A(n3861), .ZN(n3862)
         );
  OAI21_X1 U4788 ( .B1(n4142), .B2(n3863), .A(n3862), .ZN(n3868) );
  NOR2_X1 U4789 ( .A1(n3864), .A2(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n3865)
         );
  OR2_X1 U4790 ( .A1(n3875), .A2(n3865), .ZN(n5854) );
  INV_X1 U4791 ( .A(n5854), .ZN(n3866) );
  NAND2_X1 U4792 ( .A1(n3866), .A2(n4256), .ZN(n3867) );
  NAND2_X1 U4793 ( .A1(n3868), .A2(n3867), .ZN(n5548) );
  XOR2_X1 U4794 ( .A(n3870), .B(n3869), .Z(n3871) );
  NAND2_X1 U4795 ( .A1(n3871), .A2(n4111), .ZN(n3874) );
  INV_X1 U4796 ( .A(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n5634) );
  AOI21_X1 U4797 ( .B1(n5634), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n3872) );
  AOI21_X1 U4798 ( .B1(n4094), .B2(EAX_REG_23__SCAN_IN), .A(n3872), .ZN(n3873)
         );
  NAND2_X1 U4799 ( .A1(n3874), .A2(n3873), .ZN(n3877) );
  XNOR2_X1 U4800 ( .A(n3875), .B(n5634), .ZN(n5638) );
  NAND2_X1 U4801 ( .A1(n5638), .A2(n4256), .ZN(n3876) );
  NAND2_X1 U4802 ( .A1(n3877), .A2(n3876), .ZN(n5497) );
  XOR2_X1 U4803 ( .A(n4017), .B(n5499), .Z(n5486) );
  AND2_X1 U4804 ( .A1(n6498), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4257) );
  NAND2_X1 U4805 ( .A1(n4257), .A2(STATEBS16_REG_SCAN_IN), .ZN(n6508) );
  NOR2_X2 U4806 ( .A1(STATE2_REG_2__SCAN_IN), .A2(STATE2_REG_3__SCAN_IN), .ZN(
        n5826) );
  INV_X2 U4807 ( .A(n5697), .ZN(n6244) );
  NAND2_X1 U4808 ( .A1(n5486), .A2(n6244), .ZN(n3886) );
  NAND2_X1 U4809 ( .A1(n5835), .A2(n3882), .ZN(n6596) );
  NAND2_X1 U4810 ( .A1(n6596), .A2(n6498), .ZN(n3878) );
  NAND2_X1 U4811 ( .A1(n6498), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3880) );
  NAND2_X1 U4812 ( .A1(n6657), .A2(STATE2_REG_1__SCAN_IN), .ZN(n3879) );
  AND2_X1 U4813 ( .A1(n3880), .A2(n3879), .ZN(n4372) );
  INV_X1 U4814 ( .A(n4372), .ZN(n3881) );
  OR2_X2 U4815 ( .A1(n3882), .A2(STATE2_REG_2__SCAN_IN), .ZN(n6335) );
  INV_X1 U4816 ( .A(REIP_REG_24__SCAN_IN), .ZN(n3883) );
  NOR2_X1 U4817 ( .A1(n6335), .A2(n3883), .ZN(n5384) );
  NOR2_X1 U4818 ( .A1(n5691), .A2(n5490), .ZN(n3884) );
  AOI211_X1 U4819 ( .C1(n6217), .C2(n5494), .A(n5384), .B(n3884), .ZN(n3885)
         );
  OAI21_X1 U4820 ( .B1(n5386), .B2(n6221), .A(n3887), .ZN(U2962) );
  NAND2_X1 U4821 ( .A1(n4181), .A2(n3133), .ZN(n3912) );
  AND2_X4 U4822 ( .A1(n5374), .A2(n4012), .ZN(n3897) );
  INV_X1 U4823 ( .A(EBX_REG_1__SCAN_IN), .ZN(n3890) );
  NAND2_X1 U4824 ( .A1(n3897), .A2(n3890), .ZN(n3893) );
  NAND2_X1 U4825 ( .A1(n3121), .A2(n4360), .ZN(n3907) );
  NAND2_X1 U4826 ( .A1(n3907), .A2(n6331), .ZN(n3891) );
  OAI211_X1 U4827 ( .C1(n3912), .C2(EBX_REG_1__SCAN_IN), .A(n3891), .B(n3888), 
        .ZN(n3892) );
  NAND2_X1 U4828 ( .A1(n3907), .A2(EBX_REG_0__SCAN_IN), .ZN(n3895) );
  OR2_X1 U4829 ( .A1(n5374), .A2(EBX_REG_0__SCAN_IN), .ZN(n3894) );
  OAI21_X1 U4830 ( .B1(n6086), .B2(n4380), .A(n3896), .ZN(n4576) );
  INV_X1 U4831 ( .A(EBX_REG_2__SCAN_IN), .ZN(n4579) );
  NAND2_X1 U4832 ( .A1(n3897), .A2(n4579), .ZN(n3901) );
  NAND2_X1 U4833 ( .A1(n3990), .A2(n3306), .ZN(n3899) );
  OAI211_X1 U4834 ( .C1(n4380), .C2(EBX_REG_2__SCAN_IN), .A(n3899), .B(n5562), 
        .ZN(n3900) );
  MUX2_X1 U4835 ( .A(n3984), .B(n3988), .S(EBX_REG_3__SCAN_IN), .Z(n3905) );
  INV_X1 U4836 ( .A(n5374), .ZN(n5562) );
  OR2_X1 U4837 ( .A1(n4353), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n3904)
         );
  NAND2_X1 U4838 ( .A1(n3905), .A2(n3904), .ZN(n4529) );
  INV_X1 U4839 ( .A(EBX_REG_4__SCAN_IN), .ZN(n3906) );
  NAND2_X1 U4840 ( .A1(n3897), .A2(n3906), .ZN(n3911) );
  INV_X1 U4841 ( .A(n3907), .ZN(n3908) );
  NAND2_X1 U4842 ( .A1(n3990), .A2(n6320), .ZN(n3909) );
  OAI211_X1 U4843 ( .C1(n4380), .C2(EBX_REG_4__SCAN_IN), .A(n3909), .B(n5562), 
        .ZN(n3910) );
  NAND2_X1 U4844 ( .A1(n3911), .A2(n3910), .ZN(n4566) );
  OR2_X1 U4845 ( .A1(n3984), .A2(EBX_REG_5__SCAN_IN), .ZN(n3915) );
  NAND2_X1 U4846 ( .A1(n3988), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n3913)
         );
  OAI211_X1 U4847 ( .C1(n4380), .C2(EBX_REG_5__SCAN_IN), .A(n3990), .B(n3913), 
        .ZN(n3914) );
  NAND2_X1 U4848 ( .A1(n4565), .A2(n4586), .ZN(n4588) );
  NAND2_X1 U4849 ( .A1(n5562), .A2(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n3916)
         );
  NAND2_X1 U4850 ( .A1(n3990), .A2(n3916), .ZN(n3917) );
  OAI21_X1 U4851 ( .B1(EBX_REG_6__SCAN_IN), .B2(n4380), .A(n3917), .ZN(n3918)
         );
  MUX2_X1 U4852 ( .A(n3984), .B(n3988), .S(EBX_REG_7__SCAN_IN), .Z(n3921) );
  OAI21_X1 U4853 ( .B1(INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n4353), .A(n3921), 
        .ZN(n4853) );
  INV_X1 U4854 ( .A(EBX_REG_8__SCAN_IN), .ZN(n6031) );
  NAND2_X1 U4855 ( .A1(n3897), .A2(n6031), .ZN(n3925) );
  NAND2_X1 U4856 ( .A1(n3990), .A2(n3922), .ZN(n3923) );
  OAI211_X1 U4857 ( .C1(n4380), .C2(EBX_REG_8__SCAN_IN), .A(n3923), .B(n3988), 
        .ZN(n3924) );
  NAND2_X1 U4858 ( .A1(n3925), .A2(n3924), .ZN(n5025) );
  AND2_X2 U4859 ( .A1(n5026), .A2(n5025), .ZN(n5181) );
  OR2_X1 U4860 ( .A1(n4353), .A2(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n3927)
         );
  MUX2_X1 U4861 ( .A(n3984), .B(n3988), .S(EBX_REG_9__SCAN_IN), .Z(n3926) );
  AND2_X1 U4862 ( .A1(n3927), .A2(n3926), .ZN(n5180) );
  INV_X1 U4863 ( .A(EBX_REG_10__SCAN_IN), .ZN(n5525) );
  NAND2_X1 U4864 ( .A1(n3897), .A2(n5525), .ZN(n3931) );
  NAND2_X1 U4865 ( .A1(n3990), .A2(n3928), .ZN(n3929) );
  OAI211_X1 U4866 ( .C1(n4380), .C2(EBX_REG_10__SCAN_IN), .A(n3929), .B(n3988), 
        .ZN(n3930) );
  OR2_X1 U4867 ( .A1(n3984), .A2(EBX_REG_11__SCAN_IN), .ZN(n3934) );
  NAND2_X1 U4868 ( .A1(n5562), .A2(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n3932) );
  OAI211_X1 U4869 ( .C1(n4380), .C2(EBX_REG_11__SCAN_IN), .A(n3990), .B(n3932), 
        .ZN(n3933) );
  NAND2_X1 U4870 ( .A1(n3934), .A2(n3933), .ZN(n5996) );
  INV_X1 U4871 ( .A(EBX_REG_12__SCAN_IN), .ZN(n5237) );
  NAND2_X1 U4872 ( .A1(n3897), .A2(n5237), .ZN(n3938) );
  NAND2_X1 U4873 ( .A1(n3990), .A2(n6254), .ZN(n3936) );
  OAI211_X1 U4874 ( .C1(n4380), .C2(EBX_REG_12__SCAN_IN), .A(n3936), .B(n5562), 
        .ZN(n3937) );
  NAND2_X1 U4875 ( .A1(n3938), .A2(n3937), .ZN(n5218) );
  OR2_X1 U4876 ( .A1(n3984), .A2(EBX_REG_13__SCAN_IN), .ZN(n3941) );
  NAND2_X1 U4877 ( .A1(n3988), .A2(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n3939) );
  OAI211_X1 U4878 ( .C1(n4380), .C2(EBX_REG_13__SCAN_IN), .A(n3990), .B(n3939), 
        .ZN(n3940) );
  INV_X1 U4879 ( .A(EBX_REG_14__SCAN_IN), .ZN(n5979) );
  NAND2_X1 U4880 ( .A1(n3897), .A2(n5979), .ZN(n3944) );
  NAND2_X1 U4881 ( .A1(n3990), .A2(n5322), .ZN(n3942) );
  OAI211_X1 U4882 ( .C1(n4380), .C2(EBX_REG_14__SCAN_IN), .A(n3942), .B(n3988), 
        .ZN(n3943) );
  AND2_X1 U4883 ( .A1(n3944), .A2(n3943), .ZN(n5260) );
  INV_X1 U4884 ( .A(n3945), .ZN(n5302) );
  MUX2_X1 U4885 ( .A(n3984), .B(n3988), .S(EBX_REG_15__SCAN_IN), .Z(n3946) );
  OAI21_X1 U4886 ( .B1(n4353), .B2(INSTADDRPOINTER_REG_15__SCAN_IN), .A(n3946), 
        .ZN(n5303) );
  NOR2_X2 U4887 ( .A1(n5302), .A2(n5303), .ZN(n5301) );
  INV_X1 U4888 ( .A(EBX_REG_16__SCAN_IN), .ZN(n5960) );
  NAND2_X1 U4889 ( .A1(n3897), .A2(n5960), .ZN(n3949) );
  NAND2_X1 U4890 ( .A1(n3990), .A2(n5674), .ZN(n3947) );
  OAI211_X1 U4891 ( .C1(n4380), .C2(EBX_REG_16__SCAN_IN), .A(n3947), .B(n3988), 
        .ZN(n3948) );
  NAND2_X1 U4892 ( .A1(n3949), .A2(n3948), .ZN(n5313) );
  NAND2_X1 U4893 ( .A1(n5301), .A2(n5313), .ZN(n5287) );
  MUX2_X1 U4894 ( .A(n3984), .B(n5562), .S(EBX_REG_17__SCAN_IN), .Z(n3951) );
  OR2_X1 U4895 ( .A1(n4353), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n3950)
         );
  NAND2_X1 U4896 ( .A1(n3951), .A2(n3950), .ZN(n5288) );
  NOR2_X2 U4897 ( .A1(n5287), .A2(n5288), .ZN(n5286) );
  OR2_X1 U4898 ( .A1(n3987), .A2(EBX_REG_19__SCAN_IN), .ZN(n3955) );
  NAND2_X1 U4899 ( .A1(n3988), .A2(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n3952) );
  NAND2_X1 U4900 ( .A1(n3990), .A2(n3952), .ZN(n3953) );
  OAI21_X1 U4901 ( .B1(EBX_REG_19__SCAN_IN), .B2(n4380), .A(n3953), .ZN(n3954)
         );
  AND2_X1 U4902 ( .A1(n3955), .A2(n3954), .ZN(n5376) );
  NAND2_X1 U4903 ( .A1(n5286), .A2(n3956), .ZN(n5561) );
  OR2_X1 U4904 ( .A1(n4353), .A2(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n3959)
         );
  INV_X1 U4905 ( .A(EBX_REG_20__SCAN_IN), .ZN(n3957) );
  NAND2_X1 U4906 ( .A1(n4012), .A2(n3957), .ZN(n3958) );
  AND2_X1 U4907 ( .A1(n3959), .A2(n3958), .ZN(n5564) );
  OR2_X1 U4908 ( .A1(n4353), .A2(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n3961)
         );
  INV_X1 U4909 ( .A(EBX_REG_18__SCAN_IN), .ZN(n3960) );
  NAND2_X1 U4910 ( .A1(n4012), .A2(n3960), .ZN(n5375) );
  NAND2_X1 U4911 ( .A1(n3961), .A2(n5375), .ZN(n5563) );
  NAND2_X1 U4912 ( .A1(n5374), .A2(EBX_REG_20__SCAN_IN), .ZN(n3963) );
  NAND2_X1 U4913 ( .A1(n5563), .A2(n5562), .ZN(n3962) );
  OAI211_X1 U4914 ( .C1(n5564), .C2(n5563), .A(n3963), .B(n3962), .ZN(n3964)
         );
  NOR2_X2 U4915 ( .A1(n5561), .A2(n3964), .ZN(n5517) );
  MUX2_X1 U4916 ( .A(n3984), .B(n3988), .S(EBX_REG_21__SCAN_IN), .Z(n3966) );
  OR2_X1 U4917 ( .A1(n4353), .A2(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n3965)
         );
  AND2_X1 U4918 ( .A1(n3966), .A2(n3965), .ZN(n5516) );
  AND2_X2 U4919 ( .A1(n5517), .A2(n5516), .ZN(n5515) );
  OR2_X1 U4920 ( .A1(n3987), .A2(EBX_REG_22__SCAN_IN), .ZN(n3970) );
  NAND2_X1 U4921 ( .A1(n3988), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n3967) );
  NAND2_X1 U4922 ( .A1(n3990), .A2(n3967), .ZN(n3968) );
  OAI21_X1 U4923 ( .B1(EBX_REG_22__SCAN_IN), .B2(n4380), .A(n3968), .ZN(n3969)
         );
  NAND2_X1 U4924 ( .A1(n3970), .A2(n3969), .ZN(n5552) );
  NAND2_X1 U4925 ( .A1(n5515), .A2(n5552), .ZN(n5504) );
  OR2_X1 U4926 ( .A1(n3984), .A2(EBX_REG_23__SCAN_IN), .ZN(n3973) );
  NAND2_X1 U4927 ( .A1(n3988), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n3971) );
  OAI211_X1 U4928 ( .C1(n4380), .C2(EBX_REG_23__SCAN_IN), .A(n3990), .B(n3971), 
        .ZN(n3972) );
  NAND2_X1 U4929 ( .A1(n3973), .A2(n3972), .ZN(n5508) );
  OR2_X2 U4930 ( .A1(n5504), .A2(n5508), .ZN(n5506) );
  INV_X1 U4931 ( .A(EBX_REG_24__SCAN_IN), .ZN(n5491) );
  NAND2_X1 U4932 ( .A1(n3897), .A2(n5491), .ZN(n3977) );
  INV_X1 U4933 ( .A(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n3974) );
  NAND2_X1 U4934 ( .A1(n3990), .A2(n3974), .ZN(n3975) );
  OAI211_X1 U4935 ( .C1(n4380), .C2(EBX_REG_24__SCAN_IN), .A(n3975), .B(n3988), 
        .ZN(n3976) );
  AND2_X1 U4936 ( .A1(n3977), .A2(n3976), .ZN(n5381) );
  MUX2_X1 U4937 ( .A(n3984), .B(n3988), .S(EBX_REG_25__SCAN_IN), .Z(n3979) );
  OR2_X1 U4938 ( .A1(n4353), .A2(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n3978)
         );
  AND2_X1 U4939 ( .A1(n3979), .A2(n3978), .ZN(n5475) );
  OR2_X1 U4940 ( .A1(n3987), .A2(EBX_REG_26__SCAN_IN), .ZN(n3983) );
  NAND2_X1 U4941 ( .A1(n5562), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n3980) );
  NAND2_X1 U4942 ( .A1(n3990), .A2(n3980), .ZN(n3981) );
  OAI21_X1 U4943 ( .B1(EBX_REG_26__SCAN_IN), .B2(n4380), .A(n3981), .ZN(n3982)
         );
  AND2_X1 U4944 ( .A1(n3983), .A2(n3982), .ZN(n5463) );
  OR2_X2 U4945 ( .A1(n5462), .A2(n5463), .ZN(n5464) );
  MUX2_X1 U4946 ( .A(n3984), .B(n3988), .S(EBX_REG_27__SCAN_IN), .Z(n3986) );
  OR2_X1 U4947 ( .A1(n4353), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n3985)
         );
  NAND2_X1 U4948 ( .A1(n3986), .A2(n3985), .ZN(n5448) );
  OR2_X4 U4949 ( .A1(n5464), .A2(n5448), .ZN(n5450) );
  OR2_X1 U4950 ( .A1(n3987), .A2(EBX_REG_28__SCAN_IN), .ZN(n3993) );
  NAND2_X1 U4951 ( .A1(n3988), .A2(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n3989) );
  NAND2_X1 U4952 ( .A1(n3990), .A2(n3989), .ZN(n3991) );
  OAI21_X1 U4953 ( .B1(EBX_REG_28__SCAN_IN), .B2(n4380), .A(n3991), .ZN(n3992)
         );
  AND2_X1 U4954 ( .A1(n3993), .A2(n3992), .ZN(n5433) );
  NOR2_X4 U4955 ( .A1(n5450), .A2(n5433), .ZN(n5434) );
  INV_X1 U4956 ( .A(n4353), .ZN(n4188) );
  INV_X1 U4957 ( .A(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n4299) );
  NOR2_X1 U4958 ( .A1(n4380), .A2(EBX_REG_29__SCAN_IN), .ZN(n3994) );
  AOI21_X1 U4959 ( .B1(n4188), .B2(n4299), .A(n3994), .ZN(n4294) );
  AND2_X2 U4960 ( .A1(n5434), .A2(n4294), .ZN(n3999) );
  INV_X1 U4961 ( .A(n3999), .ZN(n4154) );
  AND2_X1 U4962 ( .A1(n4380), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n3995)
         );
  AOI21_X1 U4963 ( .B1(n4353), .B2(EBX_REG_30__SCAN_IN), .A(n3995), .ZN(n4156)
         );
  INV_X1 U4964 ( .A(n4156), .ZN(n3996) );
  NOR2_X1 U4965 ( .A1(n3999), .A2(n5374), .ZN(n4155) );
  AOI211_X1 U4966 ( .C1(n5434), .C2(n4154), .A(n3996), .B(n4155), .ZN(n4001)
         );
  INV_X1 U4967 ( .A(n5434), .ZN(n4153) );
  AOI21_X1 U4968 ( .B1(n4153), .B2(n5374), .A(n4156), .ZN(n3997) );
  NOR2_X1 U4969 ( .A1(n3999), .A2(n3998), .ZN(n4000) );
  NOR2_X1 U4970 ( .A1(n4001), .A2(n4000), .ZN(n5707) );
  INV_X1 U4971 ( .A(n4003), .ZN(n4343) );
  INV_X1 U4972 ( .A(n4004), .ZN(n4005) );
  NAND2_X1 U4973 ( .A1(n3134), .A2(n4005), .ZN(n4186) );
  NAND2_X1 U4974 ( .A1(n4186), .A2(n4007), .ZN(n4008) );
  OR2_X1 U4975 ( .A1(n4241), .A2(n4008), .ZN(n4009) );
  NAND2_X1 U4976 ( .A1(n4343), .A2(n4009), .ZN(n4176) );
  OR2_X1 U4977 ( .A1(n5192), .A2(n4182), .ZN(n4184) );
  AND2_X1 U4978 ( .A1(n4176), .A2(n4184), .ZN(n4444) );
  NOR2_X1 U4979 ( .A1(n5842), .A2(n4513), .ZN(n4174) );
  NAND2_X1 U4980 ( .A1(n4444), .A2(n4174), .ZN(n4428) );
  INV_X1 U4981 ( .A(n4010), .ZN(n4014) );
  NAND2_X1 U4982 ( .A1(n5396), .A2(n4509), .ZN(n4392) );
  INV_X1 U4983 ( .A(n4392), .ZN(n4013) );
  NOR2_X1 U4984 ( .A1(n4182), .A2(n3144), .ZN(n4011) );
  NAND4_X1 U4985 ( .A1(n4014), .A2(n4013), .A3(n4012), .A4(n4011), .ZN(n4015)
         );
  OAI21_X1 U4986 ( .B1(n4475), .B2(n4428), .A(n4015), .ZN(n4016) );
  AND2_X2 U4987 ( .A1(n4016), .A2(n4394), .ZN(n6095) );
  NAND2_X1 U4988 ( .A1(n6095), .A2(n5396), .ZN(n5555) );
  OR2_X1 U4989 ( .A1(n4017), .A2(n5497), .ZN(n4018) );
  AOI22_X1 U4990 ( .A1(n3853), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n4116), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n4026) );
  AOI22_X1 U4991 ( .A1(n4117), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n4021), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n4025) );
  AOI22_X1 U4992 ( .A1(n4063), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n2992), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n4024) );
  AOI22_X1 U4993 ( .A1(n4125), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n4022), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n4023) );
  NAND4_X1 U4994 ( .A1(n4026), .A2(n4025), .A3(n4024), .A4(n4023), .ZN(n4033)
         );
  AOI22_X1 U4995 ( .A1(n2994), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n4119), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n4031) );
  AOI22_X1 U4996 ( .A1(n3675), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n3232), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n4030) );
  AOI22_X1 U4997 ( .A1(n4120), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n4027), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n4029) );
  AOI22_X1 U4998 ( .A1(n4126), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n4118), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n4028) );
  NAND4_X1 U4999 ( .A1(n4031), .A2(n4030), .A3(n4029), .A4(n4028), .ZN(n4032)
         );
  NOR2_X1 U5000 ( .A1(n4033), .A2(n4032), .ZN(n4046) );
  NAND2_X1 U5001 ( .A1(n4035), .A2(n4034), .ZN(n4045) );
  XOR2_X1 U5002 ( .A(n4046), .B(n4045), .Z(n4036) );
  NAND2_X1 U5003 ( .A1(n4036), .A2(n4111), .ZN(n4040) );
  INV_X1 U5004 ( .A(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n5623) );
  NOR2_X1 U5005 ( .A1(n5623), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4037) );
  AOI211_X1 U5006 ( .C1(n3560), .C2(EAX_REG_25__SCAN_IN), .A(n4256), .B(n4037), 
        .ZN(n4039) );
  XNOR2_X1 U5007 ( .A(n4041), .B(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n5627)
         );
  AOI22_X1 U5008 ( .A1(n4040), .A2(n4039), .B1(n4256), .B2(n5627), .ZN(n5473)
         );
  INV_X1 U5009 ( .A(n4042), .ZN(n4043) );
  INV_X1 U5010 ( .A(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n5461) );
  NAND2_X1 U5011 ( .A1(n4043), .A2(n5461), .ZN(n4044) );
  NAND2_X1 U5012 ( .A1(n4078), .A2(n4044), .ZN(n5617) );
  NOR2_X1 U5013 ( .A1(n4046), .A2(n4045), .ZN(n4062) );
  AOI22_X1 U5014 ( .A1(n3853), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n4116), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n4050) );
  AOI22_X1 U5015 ( .A1(n4117), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n4021), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n4049) );
  AOI22_X1 U5016 ( .A1(n4063), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n2992), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n4048) );
  AOI22_X1 U5017 ( .A1(n4125), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n4022), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n4047) );
  NAND4_X1 U5018 ( .A1(n4050), .A2(n4049), .A3(n4048), .A4(n4047), .ZN(n4056)
         );
  AOI22_X1 U5019 ( .A1(n2994), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n4119), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n4054) );
  AOI22_X1 U5020 ( .A1(n3675), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3232), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n4053) );
  AOI22_X1 U5021 ( .A1(n4120), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n4027), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n4052) );
  AOI22_X1 U5022 ( .A1(n4126), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n4118), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n4051) );
  NAND4_X1 U5023 ( .A1(n4054), .A2(n4053), .A3(n4052), .A4(n4051), .ZN(n4055)
         );
  OR2_X1 U5024 ( .A1(n4056), .A2(n4055), .ZN(n4061) );
  XNOR2_X1 U5025 ( .A(n4062), .B(n4061), .ZN(n4059) );
  AOI21_X1 U5026 ( .B1(PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n6497), .A(n4256), 
        .ZN(n4058) );
  NAND2_X1 U5027 ( .A1(n3560), .A2(EAX_REG_26__SCAN_IN), .ZN(n4057) );
  OAI211_X1 U5028 ( .C1(n4059), .C2(n4142), .A(n4058), .B(n4057), .ZN(n4060)
         );
  OAI21_X1 U5029 ( .B1(n4139), .B2(n5617), .A(n4060), .ZN(n5460) );
  NAND2_X1 U5030 ( .A1(n4062), .A2(n4061), .ZN(n4082) );
  AOI22_X1 U5031 ( .A1(n4125), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n4063), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n4067) );
  AOI22_X1 U5032 ( .A1(n4119), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n3254), 
        .B2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n4066) );
  AOI22_X1 U5033 ( .A1(n2994), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n4118), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n4065) );
  AOI22_X1 U5034 ( .A1(n4120), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n3197), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4064) );
  NAND4_X1 U5035 ( .A1(n4067), .A2(n4066), .A3(n4065), .A4(n4064), .ZN(n4073)
         );
  AOI22_X1 U5036 ( .A1(n3853), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n4116), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n4071) );
  AOI22_X1 U5037 ( .A1(n4117), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n4021), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n4070) );
  AOI22_X1 U5038 ( .A1(n4126), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n4022), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n4069) );
  AOI22_X1 U5039 ( .A1(n4127), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n3232), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n4068) );
  NAND4_X1 U5040 ( .A1(n4071), .A2(n4070), .A3(n4069), .A4(n4068), .ZN(n4072)
         );
  NOR2_X1 U5041 ( .A1(n4073), .A2(n4072), .ZN(n4083) );
  XOR2_X1 U5042 ( .A(n4082), .B(n4083), .Z(n4074) );
  NAND2_X1 U5043 ( .A1(n4074), .A2(n4111), .ZN(n4077) );
  INV_X1 U5044 ( .A(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n5608) );
  AOI21_X1 U5045 ( .B1(n5608), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n4075) );
  AOI21_X1 U5046 ( .B1(n3560), .B2(EAX_REG_27__SCAN_IN), .A(n4075), .ZN(n4076)
         );
  XNOR2_X1 U5047 ( .A(n4078), .B(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n5612)
         );
  AOI22_X1 U5048 ( .A1(n4077), .A2(n4076), .B1(n4256), .B2(n5612), .ZN(n5447)
         );
  NAND2_X1 U5049 ( .A1(n5444), .A2(n5447), .ZN(n5431) );
  INV_X1 U5050 ( .A(n4078), .ZN(n4079) );
  NAND2_X1 U5051 ( .A1(n4079), .A2(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n4080)
         );
  INV_X1 U5052 ( .A(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n5436) );
  NAND2_X1 U5053 ( .A1(n4080), .A2(n5436), .ZN(n4081) );
  NAND2_X1 U5054 ( .A1(n4144), .A2(n4081), .ZN(n5601) );
  NOR2_X1 U5055 ( .A1(n4083), .A2(n4082), .ZN(n4100) );
  AOI22_X1 U5056 ( .A1(n3853), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n4116), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n4087) );
  AOI22_X1 U5057 ( .A1(n4117), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n4021), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n4086) );
  AOI22_X1 U5058 ( .A1(n4063), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n2992), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n4085) );
  AOI22_X1 U5059 ( .A1(n4125), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n4022), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n4084) );
  NAND4_X1 U5060 ( .A1(n4087), .A2(n4086), .A3(n4085), .A4(n4084), .ZN(n4093)
         );
  AOI22_X1 U5061 ( .A1(n2994), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n4119), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n4091) );
  AOI22_X1 U5062 ( .A1(n4127), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n3324), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n4090) );
  AOI22_X1 U5063 ( .A1(n4120), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3197), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4089) );
  AOI22_X1 U5064 ( .A1(n4126), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n4118), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n4088) );
  NAND4_X1 U5065 ( .A1(n4091), .A2(n4090), .A3(n4089), .A4(n4088), .ZN(n4092)
         );
  OR2_X1 U5066 ( .A1(n4093), .A2(n4092), .ZN(n4099) );
  XNOR2_X1 U5067 ( .A(n4100), .B(n4099), .ZN(n4097) );
  AOI21_X1 U5068 ( .B1(PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n6497), .A(n4256), 
        .ZN(n4096) );
  NAND2_X1 U5069 ( .A1(n4094), .A2(EAX_REG_28__SCAN_IN), .ZN(n4095) );
  OAI211_X1 U5070 ( .C1(n4097), .C2(n4142), .A(n4096), .B(n4095), .ZN(n4098)
         );
  OAI21_X1 U5071 ( .B1(n4139), .B2(n5601), .A(n4098), .ZN(n5432) );
  NAND2_X1 U5072 ( .A1(n4100), .A2(n4099), .ZN(n4134) );
  AOI22_X1 U5073 ( .A1(n3853), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3106), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n4104) );
  AOI22_X1 U5074 ( .A1(n4063), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n4022), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n4103) );
  AOI22_X1 U5075 ( .A1(n4127), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n3324), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n4102) );
  AOI22_X1 U5076 ( .A1(n4126), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n4118), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n4101) );
  NAND4_X1 U5077 ( .A1(n4104), .A2(n4103), .A3(n4102), .A4(n4101), .ZN(n4110)
         );
  AOI22_X1 U5078 ( .A1(n4117), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n4021), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n4108) );
  AOI22_X1 U5079 ( .A1(n2994), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n4119), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n4107) );
  AOI22_X1 U5080 ( .A1(n4125), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n2992), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n4106) );
  AOI22_X1 U5081 ( .A1(n4120), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n2997), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4105) );
  NAND4_X1 U5082 ( .A1(n4108), .A2(n4107), .A3(n4106), .A4(n4105), .ZN(n4109)
         );
  NOR2_X1 U5083 ( .A1(n4110), .A2(n4109), .ZN(n4135) );
  XOR2_X1 U5084 ( .A(n4134), .B(n4135), .Z(n4112) );
  NAND2_X1 U5085 ( .A1(n4112), .A2(n4111), .ZN(n4115) );
  INV_X1 U5086 ( .A(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n4328) );
  NOR2_X1 U5087 ( .A1(n4328), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4113) );
  AOI211_X1 U5088 ( .C1(n3560), .C2(EAX_REG_29__SCAN_IN), .A(n4256), .B(n4113), 
        .ZN(n4114) );
  XNOR2_X1 U5089 ( .A(n4144), .B(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n5423)
         );
  AOI22_X1 U5090 ( .A1(n4115), .A2(n4114), .B1(n4256), .B2(n5423), .ZN(n4327)
         );
  AOI22_X1 U5091 ( .A1(n4116), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n4021), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n4124) );
  AOI22_X1 U5092 ( .A1(n4117), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3254), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n4123) );
  AOI22_X1 U5093 ( .A1(n4119), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n4118), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n4122) );
  AOI22_X1 U5094 ( .A1(n4120), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3324), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n4121) );
  NAND4_X1 U5095 ( .A1(n4124), .A2(n4123), .A3(n4122), .A4(n4121), .ZN(n4133)
         );
  AOI22_X1 U5096 ( .A1(n3853), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n4125), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n4131) );
  AOI22_X1 U5097 ( .A1(n2994), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n4126), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n4130) );
  AOI22_X1 U5098 ( .A1(n4063), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n4022), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n4129) );
  AOI22_X1 U5099 ( .A1(n4127), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3197), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4128) );
  NAND4_X1 U5100 ( .A1(n4131), .A2(n4130), .A3(n4129), .A4(n4128), .ZN(n4132)
         );
  NOR2_X1 U5101 ( .A1(n4133), .A2(n4132), .ZN(n4137) );
  NOR2_X1 U5102 ( .A1(n4135), .A2(n4134), .ZN(n4136) );
  XOR2_X1 U5103 ( .A(n4137), .B(n4136), .Z(n4143) );
  NAND2_X1 U5104 ( .A1(n6497), .A2(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n4138)
         );
  NAND2_X1 U5105 ( .A1(n4139), .A2(n4138), .ZN(n4140) );
  AOI21_X1 U5106 ( .B1(n3560), .B2(EAX_REG_30__SCAN_IN), .A(n4140), .ZN(n4141)
         );
  OAI21_X1 U5107 ( .B1(n4143), .B2(n4142), .A(n4141), .ZN(n4147) );
  INV_X1 U5108 ( .A(n4144), .ZN(n4145) );
  NAND2_X1 U5109 ( .A1(n4145), .A2(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n4276)
         );
  XNOR2_X1 U5110 ( .A(n4276), .B(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n5406)
         );
  NAND2_X1 U5111 ( .A1(n5406), .A2(n4256), .ZN(n4146) );
  NAND2_X1 U5112 ( .A1(n4147), .A2(n4146), .ZN(n4272) );
  NAND2_X1 U5113 ( .A1(n6095), .A2(n3164), .ZN(n5576) );
  INV_X1 U5114 ( .A(EBX_REG_30__SCAN_IN), .ZN(n4316) );
  NAND2_X1 U5115 ( .A1(n4150), .A2(EBX_REG_30__SCAN_IN), .ZN(n4151) );
  OAI211_X1 U5116 ( .C1(n5707), .C2(n5555), .A(n4152), .B(n4151), .ZN(U2829)
         );
  INV_X1 U5117 ( .A(EBX_REG_29__SCAN_IN), .ZN(n5380) );
  NAND2_X1 U5118 ( .A1(n3897), .A2(n5380), .ZN(n4295) );
  OAI21_X1 U5119 ( .B1(n4154), .B2(n5374), .A(n2999), .ZN(n4293) );
  AOI21_X1 U5120 ( .B1(n4156), .B2(n4293), .A(n4155), .ZN(n4158) );
  OAI22_X1 U5121 ( .A1(n4353), .A2(INSTADDRPOINTER_REG_31__SCAN_IN), .B1(
        EBX_REG_31__SCAN_IN), .B2(n4380), .ZN(n4157) );
  OR2_X1 U5122 ( .A1(n4159), .A2(STATE_REG_0__SCAN_IN), .ZN(n6519) );
  NAND2_X1 U5123 ( .A1(n4181), .A2(n6519), .ZN(n4166) );
  AND2_X1 U5124 ( .A1(n4161), .A2(n4160), .ZN(n4162) );
  AND2_X1 U5125 ( .A1(n4163), .A2(n4162), .ZN(n4164) );
  NOR2_X1 U5126 ( .A1(READY_N), .A2(n4249), .ZN(n4389) );
  NAND2_X1 U5127 ( .A1(n4166), .A2(n4389), .ZN(n4173) );
  NAND2_X1 U5128 ( .A1(n4513), .A2(n6519), .ZN(n4251) );
  NAND2_X1 U5129 ( .A1(n4251), .A2(n6487), .ZN(n4170) );
  INV_X1 U5130 ( .A(n4398), .ZN(n4169) );
  OAI211_X1 U5131 ( .C1(n4168), .C2(n4170), .A(n4360), .B(n4169), .ZN(n4171)
         );
  NAND2_X1 U5132 ( .A1(n4475), .A2(n4171), .ZN(n4172) );
  MUX2_X1 U5133 ( .A(n4173), .B(n4172), .S(n3298), .Z(n4177) );
  INV_X1 U5134 ( .A(n4174), .ZN(n4175) );
  OR2_X1 U5135 ( .A1(n4475), .A2(n4175), .ZN(n4446) );
  NAND3_X1 U5136 ( .A1(n4177), .A2(n4176), .A3(n4446), .ZN(n4178) );
  OR2_X1 U5137 ( .A1(n4168), .A2(n6599), .ZN(n6490) );
  NAND3_X1 U5138 ( .A1(n4423), .A2(n4509), .A3(n4398), .ZN(n4179) );
  AND2_X1 U5139 ( .A1(n6490), .A2(n4179), .ZN(n4180) );
  NAND2_X1 U5140 ( .A1(n4003), .A2(n4181), .ZN(n6462) );
  NAND2_X1 U5141 ( .A1(n4398), .A2(n4518), .ZN(n4183) );
  NAND2_X1 U5142 ( .A1(n4183), .A2(n4182), .ZN(n4185) );
  AND3_X1 U5143 ( .A1(n4186), .A2(n4185), .A3(n4184), .ZN(n4187) );
  OAI21_X1 U5144 ( .B1(n4189), .B2(n4188), .A(n4187), .ZN(n4190) );
  OR2_X1 U5145 ( .A1(n4191), .A2(n4190), .ZN(n4422) );
  INV_X1 U5146 ( .A(n4456), .ZN(n4192) );
  NOR2_X1 U5147 ( .A1(n4422), .A2(n4192), .ZN(n4193) );
  NAND2_X1 U5148 ( .A1(n5909), .A2(n5326), .ZN(n5784) );
  INV_X1 U5149 ( .A(n5784), .ZN(n4194) );
  NAND2_X1 U5150 ( .A1(n4194), .A2(n5336), .ZN(n6297) );
  NAND2_X1 U5151 ( .A1(INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n4300) );
  INV_X1 U5152 ( .A(n4300), .ZN(n5719) );
  AND2_X1 U5153 ( .A1(INSTADDRPOINTER_REG_30__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n4195) );
  NAND2_X1 U5154 ( .A1(n5719), .A2(n4195), .ZN(n4214) );
  INV_X1 U5155 ( .A(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n5387) );
  NAND2_X1 U5156 ( .A1(n5909), .A2(n5387), .ZN(n4385) );
  NAND2_X1 U5157 ( .A1(n5784), .A2(n4385), .ZN(n6330) );
  INV_X1 U5158 ( .A(n6330), .ZN(n4198) );
  NAND2_X1 U5159 ( .A1(INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n5337) );
  NAND3_X1 U5160 ( .A1(INSTADDRPOINTER_REG_3__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_4__SCAN_IN), .A3(INSTADDRPOINTER_REG_5__SCAN_IN), 
        .ZN(n6296) );
  NOR2_X1 U5161 ( .A1(n6304), .A2(n6296), .ZN(n6263) );
  NAND2_X1 U5162 ( .A1(INSTADDRPOINTER_REG_7__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n6282) );
  INV_X1 U5163 ( .A(n6282), .ZN(n6265) );
  NAND4_X1 U5164 ( .A1(INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_10__SCAN_IN), .A3(n6263), .A4(n6265), .ZN(n5339)
         );
  NOR2_X1 U5165 ( .A1(n5337), .A2(n5339), .ZN(n5911) );
  INV_X1 U5166 ( .A(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n4196) );
  NAND2_X1 U5167 ( .A1(INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n5334) );
  NOR2_X1 U5168 ( .A1(n4196), .A2(n5334), .ZN(n5350) );
  NAND2_X1 U5169 ( .A1(INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n5350), .ZN(n5351) );
  NAND2_X1 U5170 ( .A1(INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5355) );
  NOR2_X1 U5171 ( .A1(n5351), .A2(n5355), .ZN(n4199) );
  NAND2_X1 U5172 ( .A1(n5911), .A2(n4199), .ZN(n4203) );
  INV_X1 U5173 ( .A(n4203), .ZN(n4197) );
  NAND2_X1 U5174 ( .A1(n4198), .A2(n4197), .ZN(n5805) );
  INV_X1 U5175 ( .A(n5336), .ZN(n6334) );
  NOR2_X1 U5176 ( .A1(INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n6333), .ZN(n6298)
         );
  NOR2_X1 U5177 ( .A1(n5339), .A2(n6298), .ZN(n5327) );
  AND2_X1 U5178 ( .A1(n5327), .A2(n4199), .ZN(n5816) );
  NAND2_X1 U5179 ( .A1(n6334), .A2(n5816), .ZN(n4200) );
  NAND2_X1 U5180 ( .A1(n5805), .A2(n4200), .ZN(n4202) );
  AND2_X1 U5181 ( .A1(INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n4219) );
  AND2_X1 U5182 ( .A1(n4201), .A2(n4219), .ZN(n4205) );
  NAND2_X1 U5183 ( .A1(n4202), .A2(n4205), .ZN(n4213) );
  AND2_X1 U5184 ( .A1(INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5630) );
  OR2_X1 U5185 ( .A1(n4213), .A2(n5630), .ZN(n5765) );
  NAND2_X1 U5186 ( .A1(n4244), .A2(n6335), .ZN(n4382) );
  OAI21_X1 U5187 ( .B1(n5326), .B2(INSTADDRPOINTER_REG_0__SCAN_IN), .A(n4382), 
        .ZN(n5331) );
  AND2_X1 U5188 ( .A1(n5784), .A2(n4203), .ZN(n4204) );
  NOR2_X1 U5189 ( .A1(n5331), .A2(n4204), .ZN(n5783) );
  INV_X1 U5190 ( .A(n5816), .ZN(n4207) );
  INV_X1 U5191 ( .A(n4205), .ZN(n4206) );
  OAI21_X1 U5192 ( .B1(n4207), .B2(n4206), .A(n6297), .ZN(n4208) );
  AND2_X1 U5193 ( .A1(n5783), .A2(n4208), .ZN(n5775) );
  AND2_X1 U5194 ( .A1(n5765), .A2(n5775), .ZN(n5767) );
  NAND2_X1 U5195 ( .A1(n6330), .A2(n5336), .ZN(n4210) );
  AND2_X1 U5196 ( .A1(INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n4220) );
  INV_X1 U5197 ( .A(n4220), .ZN(n4209) );
  NAND2_X1 U5198 ( .A1(n4210), .A2(n4209), .ZN(n4211) );
  NAND2_X1 U5199 ( .A1(INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5739) );
  NAND2_X1 U5200 ( .A1(n6297), .A2(n5739), .ZN(n4212) );
  NAND2_X1 U5201 ( .A1(n5751), .A2(n4212), .ZN(n5733) );
  AOI21_X1 U5202 ( .B1(n6297), .B2(n4214), .A(n5733), .ZN(n4217) );
  NAND2_X1 U5203 ( .A1(n2993), .A2(REIP_REG_31__SCAN_IN), .ZN(n4283) );
  INV_X1 U5204 ( .A(n4213), .ZN(n5778) );
  NAND2_X1 U5205 ( .A1(n5756), .A2(n4220), .ZN(n5737) );
  NOR2_X1 U5206 ( .A1(n5737), .A2(n5739), .ZN(n5711) );
  INV_X1 U5207 ( .A(n4214), .ZN(n4215) );
  NAND3_X1 U5208 ( .A1(n5711), .A2(n4215), .A3(n4234), .ZN(n4216) );
  OAI211_X1 U5209 ( .C1(n4217), .C2(n4234), .A(n4283), .B(n4216), .ZN(n4218)
         );
  AOI21_X1 U5210 ( .B1(n5538), .B2(n6323), .A(n4218), .ZN(n4246) );
  NAND2_X1 U5211 ( .A1(n4222), .A2(n3004), .ZN(n4221) );
  NAND2_X1 U5212 ( .A1(n4221), .A2(n5629), .ZN(n4227) );
  INV_X1 U5213 ( .A(n4222), .ZN(n5662) );
  NOR2_X1 U5214 ( .A1(INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n4224) );
  NOR2_X1 U5215 ( .A1(INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n4223) );
  INV_X1 U5216 ( .A(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5777) );
  AND4_X1 U5217 ( .A1(n4224), .A2(n4223), .A3(n5777), .A4(n5799), .ZN(n4225)
         );
  NAND2_X1 U5218 ( .A1(n5662), .A2(n4225), .ZN(n4226) );
  AND2_X2 U5219 ( .A1(n4227), .A2(n4226), .ZN(n5596) );
  XOR2_X1 U5220 ( .A(INSTADDRPOINTER_REG_25__SCAN_IN), .B(n5629), .Z(n5622) );
  INV_X1 U5221 ( .A(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5750) );
  NAND2_X1 U5222 ( .A1(n4288), .A2(n4229), .ZN(n5606) );
  NOR2_X2 U5223 ( .A1(n5606), .A2(n4300), .ZN(n5402) );
  NAND2_X1 U5224 ( .A1(n5402), .A2(n4195), .ZN(n4233) );
  NOR2_X1 U5225 ( .A1(INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5720) );
  INV_X1 U5226 ( .A(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5742) );
  NAND2_X1 U5227 ( .A1(n5720), .A2(n5742), .ZN(n4231) );
  INV_X1 U5228 ( .A(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n5710) );
  NAND4_X1 U5229 ( .A1(n5621), .A2(n4289), .A3(n5710), .A4(n4299), .ZN(n4232)
         );
  NAND2_X1 U5230 ( .A1(n4233), .A2(n4232), .ZN(n4235) );
  XNOR2_X1 U5231 ( .A(n4235), .B(n4234), .ZN(n4285) );
  OR2_X1 U5232 ( .A1(n4238), .A2(n4509), .ZN(n4239) );
  AND2_X1 U5233 ( .A1(n6479), .A2(n4239), .ZN(n4242) );
  NOR2_X1 U5234 ( .A1(n4241), .A2(n4240), .ZN(n4388) );
  INV_X1 U5235 ( .A(n4388), .ZN(n4427) );
  OR2_X1 U5236 ( .A1(n4168), .A2(n4380), .ZN(n4441) );
  AND4_X1 U5237 ( .A1(n4237), .A2(n4242), .A3(n4427), .A4(n4441), .ZN(n4243)
         );
  NAND2_X1 U5238 ( .A1(n4285), .A2(n6340), .ZN(n4245) );
  NAND2_X1 U5239 ( .A1(n4246), .A2(n4245), .ZN(U2987) );
  INV_X1 U5240 ( .A(n4249), .ZN(n4344) );
  AND2_X1 U5241 ( .A1(n4003), .A2(n4344), .ZN(n4338) );
  NAND2_X1 U5242 ( .A1(n4338), .A2(n4394), .ZN(n4336) );
  INV_X1 U5243 ( .A(EBX_REG_31__SCAN_IN), .ZN(n5539) );
  NOR2_X1 U5244 ( .A1(n5193), .A2(n5539), .ZN(n4267) );
  NOR2_X1 U5245 ( .A1(STATEBS16_REG_SCAN_IN), .A2(READY_N), .ZN(n4308) );
  NOR2_X1 U5246 ( .A1(n4380), .A2(n4308), .ZN(n4250) );
  INV_X1 U5247 ( .A(REIP_REG_22__SCAN_IN), .ZN(n6560) );
  NAND3_X1 U5248 ( .A1(n4251), .A2(n4308), .A3(n4360), .ZN(n4252) );
  INV_X1 U5249 ( .A(REIP_REG_19__SCAN_IN), .ZN(n6706) );
  INV_X1 U5250 ( .A(REIP_REG_17__SCAN_IN), .ZN(n6555) );
  INV_X1 U5251 ( .A(REIP_REG_15__SCAN_IN), .ZN(n6552) );
  INV_X1 U5252 ( .A(REIP_REG_13__SCAN_IN), .ZN(n6549) );
  INV_X1 U5253 ( .A(REIP_REG_12__SCAN_IN), .ZN(n6547) );
  INV_X1 U5254 ( .A(REIP_REG_10__SCAN_IN), .ZN(n6544) );
  INV_X1 U5255 ( .A(REIP_REG_7__SCAN_IN), .ZN(n4253) );
  INV_X1 U5256 ( .A(REIP_REG_4__SCAN_IN), .ZN(n6536) );
  NAND3_X1 U5257 ( .A1(REIP_REG_1__SCAN_IN), .A2(REIP_REG_3__SCAN_IN), .A3(
        REIP_REG_2__SCAN_IN), .ZN(n6040) );
  NOR2_X1 U5258 ( .A1(n6536), .A2(n6040), .ZN(n5202) );
  NAND2_X1 U5259 ( .A1(REIP_REG_5__SCAN_IN), .A2(n5202), .ZN(n5079) );
  INV_X1 U5260 ( .A(n5079), .ZN(n5080) );
  NAND2_X1 U5261 ( .A1(REIP_REG_6__SCAN_IN), .A2(n5080), .ZN(n5081) );
  NOR2_X1 U5262 ( .A1(n4253), .A2(n5081), .ZN(n6022) );
  NAND2_X1 U5263 ( .A1(REIP_REG_8__SCAN_IN), .A2(n6022), .ZN(n6021) );
  INV_X1 U5264 ( .A(n6021), .ZN(n5531) );
  NAND2_X1 U5265 ( .A1(REIP_REG_9__SCAN_IN), .A2(n5531), .ZN(n5527) );
  NOR2_X1 U5266 ( .A1(n6544), .A2(n5527), .ZN(n6001) );
  NAND2_X1 U5267 ( .A1(REIP_REG_11__SCAN_IN), .A2(n6001), .ZN(n5988) );
  NOR3_X1 U5268 ( .A1(n6549), .A2(n6547), .A3(n5988), .ZN(n5978) );
  NAND2_X1 U5269 ( .A1(REIP_REG_14__SCAN_IN), .A2(n5978), .ZN(n5953) );
  NOR2_X1 U5270 ( .A1(n6552), .A2(n5953), .ZN(n5956) );
  NAND2_X1 U5271 ( .A1(REIP_REG_16__SCAN_IN), .A2(n5956), .ZN(n5295) );
  NOR2_X1 U5272 ( .A1(n6555), .A2(n5295), .ZN(n5944) );
  NAND2_X1 U5273 ( .A1(REIP_REG_18__SCAN_IN), .A2(n5944), .ZN(n5867) );
  NOR2_X1 U5274 ( .A1(n6706), .A2(n5867), .ZN(n5859) );
  NAND2_X1 U5275 ( .A1(REIP_REG_20__SCAN_IN), .A2(n5859), .ZN(n4261) );
  NOR2_X1 U5276 ( .A1(n6065), .A2(n4261), .ZN(n5519) );
  NAND2_X1 U5277 ( .A1(REIP_REG_21__SCAN_IN), .A2(n5519), .ZN(n5851) );
  NOR2_X1 U5278 ( .A1(n6560), .A2(n5851), .ZN(n5502) );
  NAND2_X1 U5279 ( .A1(REIP_REG_23__SCAN_IN), .A2(n5502), .ZN(n5489) );
  NAND3_X1 U5280 ( .A1(REIP_REG_24__SCAN_IN), .A2(REIP_REG_26__SCAN_IN), .A3(
        REIP_REG_25__SCAN_IN), .ZN(n5452) );
  INV_X1 U5281 ( .A(n5452), .ZN(n4262) );
  NAND2_X1 U5282 ( .A1(REIP_REG_27__SCAN_IN), .A2(n4262), .ZN(n4254) );
  NOR2_X1 U5283 ( .A1(n5489), .A2(n4254), .ZN(n5438) );
  NAND2_X1 U5284 ( .A1(n5438), .A2(REIP_REG_28__SCAN_IN), .ZN(n5426) );
  INV_X1 U5285 ( .A(REIP_REG_31__SCAN_IN), .ZN(n4255) );
  NAND3_X1 U5286 ( .A1(n4255), .A2(REIP_REG_30__SCAN_IN), .A3(
        REIP_REG_29__SCAN_IN), .ZN(n4270) );
  INV_X1 U5287 ( .A(REIP_REG_23__SCAN_IN), .ZN(n6666) );
  INV_X1 U5288 ( .A(REIP_REG_21__SCAN_IN), .ZN(n6703) );
  INV_X1 U5289 ( .A(STATE2_REG_3__SCAN_IN), .ZN(n6581) );
  NOR2_X1 U5290 ( .A1(STATE2_REG_1__SCAN_IN), .A2(STATE2_REG_2__SCAN_IN), .ZN(
        n6600) );
  INV_X1 U5291 ( .A(n6600), .ZN(n6507) );
  NOR3_X1 U5292 ( .A1(n6498), .A2(n6581), .A3(n6507), .ZN(n6492) );
  AND2_X1 U5293 ( .A1(n4257), .A2(n4256), .ZN(n6502) );
  INV_X1 U5294 ( .A(n6502), .ZN(n4258) );
  NAND2_X1 U5295 ( .A1(n4258), .A2(n6335), .ZN(n4259) );
  OR2_X1 U5296 ( .A1(n6492), .A2(n4259), .ZN(n4260) );
  INV_X1 U5297 ( .A(n6046), .ZN(n6075) );
  OR2_X1 U5298 ( .A1(n4261), .A2(n6075), .ZN(n5514) );
  NOR4_X1 U5299 ( .A1(n6666), .A2(n6560), .A3(n6703), .A4(n5514), .ZN(n5487)
         );
  AND2_X1 U5300 ( .A1(n5487), .A2(n4262), .ZN(n4263) );
  NAND2_X1 U5301 ( .A1(n6065), .A2(n6046), .ZN(n6067) );
  INV_X1 U5302 ( .A(n6067), .ZN(n5488) );
  OR2_X1 U5303 ( .A1(n4263), .A2(n5488), .ZN(n5470) );
  NAND2_X1 U5304 ( .A1(REIP_REG_28__SCAN_IN), .A2(REIP_REG_27__SCAN_IN), .ZN(
        n4264) );
  NAND2_X1 U5305 ( .A1(n6083), .A2(n4264), .ZN(n4265) );
  AND2_X1 U5306 ( .A1(n5470), .A2(n4265), .ZN(n5422) );
  OAI211_X1 U5307 ( .C1(REIP_REG_29__SCAN_IN), .C2(n6065), .A(n5422), .B(
        REIP_REG_30__SCAN_IN), .ZN(n4320) );
  NAND3_X1 U5308 ( .A1(n4320), .A2(REIP_REG_31__SCAN_IN), .A3(n6067), .ZN(
        n4269) );
  INV_X1 U5309 ( .A(n6519), .ZN(n4266) );
  NAND2_X1 U5310 ( .A1(n4266), .A2(n4308), .ZN(n6491) );
  AND2_X1 U5311 ( .A1(n6130), .A2(n6491), .ZN(n4311) );
  AOI22_X1 U5312 ( .A1(n4267), .A2(n4311), .B1(PHYADDRPOINTER_REG_31__SCAN_IN), 
        .B2(n6059), .ZN(n4268) );
  OAI211_X1 U5313 ( .C1(n5426), .C2(n4270), .A(n4269), .B(n4268), .ZN(n4271)
         );
  AOI21_X1 U5314 ( .B1(n5538), .B2(n6047), .A(n4271), .ZN(n4281) );
  AOI22_X1 U5315 ( .A1(n4094), .A2(EAX_REG_31__SCAN_IN), .B1(n4273), .B2(
        PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n4274) );
  INV_X1 U5316 ( .A(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n5408) );
  INV_X1 U5317 ( .A(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n4277) );
  NOR2_X1 U5318 ( .A1(n4313), .A2(n5413), .ZN(n4279) );
  NAND2_X1 U5319 ( .A1(n4281), .A2(n4280), .ZN(U2796) );
  NAND2_X1 U5320 ( .A1(n6239), .A2(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n4282)
         );
  OAI211_X1 U5321 ( .C1(n6249), .C2(n4313), .A(n4283), .B(n4282), .ZN(n4284)
         );
  AOI21_X1 U5322 ( .B1(n5399), .B2(n6244), .A(n4284), .ZN(n4287) );
  NAND2_X1 U5323 ( .A1(n4285), .A2(n6243), .ZN(n4286) );
  NAND2_X1 U5324 ( .A1(n4287), .A2(n4286), .ZN(U2955) );
  INV_X1 U5325 ( .A(n5615), .ZN(n4290) );
  NAND2_X1 U5326 ( .A1(n4290), .A2(n4289), .ZN(n5404) );
  INV_X1 U5327 ( .A(n5402), .ZN(n4291) );
  NAND2_X1 U5328 ( .A1(n4323), .A2(n6340), .ZN(n4306) );
  NAND2_X1 U5329 ( .A1(n4294), .A2(n5562), .ZN(n4296) );
  NAND2_X1 U5330 ( .A1(n4296), .A2(n4295), .ZN(n4297) );
  NOR2_X1 U5331 ( .A1(n5434), .A2(n4297), .ZN(n4298) );
  AOI211_X1 U5332 ( .C1(n4300), .C2(n6297), .A(n4299), .B(n5733), .ZN(n5708)
         );
  INV_X1 U5333 ( .A(n5708), .ZN(n4302) );
  INV_X1 U5334 ( .A(n5711), .ZN(n5729) );
  OAI21_X1 U5335 ( .B1(n5729), .B2(n4300), .A(n4299), .ZN(n4301) );
  INV_X1 U5336 ( .A(REIP_REG_29__SCAN_IN), .ZN(n6702) );
  NOR2_X1 U5337 ( .A1(n6335), .A2(n6702), .ZN(n4330) );
  AOI21_X1 U5338 ( .B1(n4302), .B2(n4301), .A(n4330), .ZN(n4303) );
  NAND2_X1 U5339 ( .A1(n4306), .A2(n4305), .ZN(U2989) );
  INV_X1 U5340 ( .A(REIP_REG_30__SCAN_IN), .ZN(n4307) );
  OAI21_X1 U5341 ( .B1(n5426), .B2(n6702), .A(n4307), .ZN(n4319) );
  NOR2_X1 U5342 ( .A1(n4308), .A2(EBX_REG_31__SCAN_IN), .ZN(n4309) );
  AND2_X1 U5343 ( .A1(n4360), .A2(n4309), .ZN(n4310) );
  NOR2_X1 U5344 ( .A1(n4311), .A2(n4310), .ZN(n4312) );
  AOI22_X1 U5345 ( .A1(PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n6059), .B1(n5194), 
        .B2(n5406), .ZN(n4315) );
  OAI21_X1 U5346 ( .B1(n4316), .B2(n6030), .A(n4315), .ZN(n4318) );
  NOR2_X1 U5347 ( .A1(n5707), .A2(n6087), .ZN(n4317) );
  AOI211_X1 U5348 ( .C1(n4320), .C2(n4319), .A(n4318), .B(n4317), .ZN(n4322)
         );
  NAND2_X1 U5349 ( .A1(n4322), .A2(n4321), .ZN(U2797) );
  NAND2_X1 U5350 ( .A1(n4323), .A2(n6243), .ZN(n4334) );
  NOR2_X1 U5351 ( .A1(n5691), .A2(n4328), .ZN(n4329) );
  AOI211_X1 U5352 ( .C1(n6217), .C2(n5423), .A(n4330), .B(n4329), .ZN(n4331)
         );
  NAND2_X1 U5353 ( .A1(n4334), .A2(n4333), .ZN(U2957) );
  AND2_X1 U5354 ( .A1(n5826), .A2(n5413), .ZN(n4349) );
  INV_X1 U5355 ( .A(n4335), .ZN(n6129) );
  AOI211_X1 U5356 ( .C1(MEMORYFETCH_REG_SCAN_IN), .C2(n4336), .A(n4349), .B(
        n6129), .ZN(n4337) );
  INV_X1 U5357 ( .A(n4337), .ZN(U2788) );
  OR2_X1 U5358 ( .A1(n4475), .A2(n3461), .ZN(n4341) );
  INV_X1 U5359 ( .A(n4338), .ZN(n4339) );
  NAND2_X1 U5360 ( .A1(n4339), .A2(n4248), .ZN(n4340) );
  NAND2_X1 U5361 ( .A1(n4341), .A2(n4340), .ZN(n5923) );
  INV_X1 U5362 ( .A(n5192), .ZN(n4342) );
  OR2_X1 U5363 ( .A1(n6130), .A2(n4342), .ZN(n4351) );
  AOI21_X1 U5364 ( .B1(n4351), .B2(n6519), .A(READY_N), .ZN(n6598) );
  NOR2_X1 U5365 ( .A1(n5923), .A2(n6598), .ZN(n6478) );
  OR2_X1 U5366 ( .A1(n6478), .A2(n6500), .ZN(n5927) );
  INV_X1 U5367 ( .A(n4428), .ZN(n4347) );
  AND3_X1 U5368 ( .A1(n4427), .A2(n6479), .A3(n4248), .ZN(n4345) );
  OAI22_X1 U5369 ( .A1(n4475), .A2(n4345), .B1(n4344), .B2(n4343), .ZN(n4346)
         );
  AOI21_X1 U5370 ( .B1(n4347), .B2(n4475), .A(n4346), .ZN(n6480) );
  NAND2_X1 U5371 ( .A1(n5927), .A2(MORE_REG_SCAN_IN), .ZN(n4348) );
  OAI21_X1 U5372 ( .B1(n5927), .B2(n6480), .A(n4348), .ZN(U3471) );
  OAI21_X1 U5373 ( .B1(n4349), .B2(READREQUEST_REG_SCAN_IN), .A(n5193), .ZN(
        n4350) );
  OAI21_X1 U5374 ( .B1(n5193), .B2(n4351), .A(n4350), .ZN(U3474) );
  XNOR2_X1 U5375 ( .A(n4352), .B(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4373)
         );
  NOR2_X1 U5376 ( .A1(n4353), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4354)
         );
  OR2_X1 U5377 ( .A1(n4355), .A2(n4354), .ZN(n5197) );
  INV_X1 U5378 ( .A(n5197), .ZN(n4357) );
  AND2_X1 U5379 ( .A1(n2993), .A2(REIP_REG_0__SCAN_IN), .ZN(n4375) );
  AOI21_X1 U5380 ( .B1(n5909), .B2(n4382), .A(n5387), .ZN(n4356) );
  AOI211_X1 U5381 ( .C1(n6323), .C2(n4357), .A(n4375), .B(n4356), .ZN(n4358)
         );
  NAND2_X1 U5382 ( .A1(n5336), .A2(n5326), .ZN(n5333) );
  NAND2_X1 U5383 ( .A1(n5333), .A2(n5387), .ZN(n4381) );
  OAI211_X1 U5384 ( .C1(n4373), .C2(n6300), .A(n4358), .B(n4381), .ZN(U3018)
         );
  INV_X1 U5385 ( .A(EAX_REG_25__SCAN_IN), .ZN(n6150) );
  AND2_X1 U5386 ( .A1(n6490), .A2(n6462), .ZN(n4359) );
  NAND2_X1 U5387 ( .A1(n4361), .A2(n4360), .ZN(n4419) );
  NAND2_X1 U5388 ( .A1(STATE2_REG_1__SCAN_IN), .A2(STATE2_REG_2__SCAN_IN), 
        .ZN(n4478) );
  NOR2_X1 U5389 ( .A1(n4478), .A2(STATE2_REG_0__SCAN_IN), .ZN(n6112) );
  INV_X1 U5390 ( .A(n6112), .ZN(n6486) );
  AOI22_X1 U5391 ( .A1(n6597), .A2(UWORD_REG_9__SCAN_IN), .B1(n6123), .B2(
        DATAO_REG_25__SCAN_IN), .ZN(n4362) );
  OAI21_X1 U5392 ( .B1(n6150), .B2(n4419), .A(n4362), .ZN(U2898) );
  INV_X1 U5393 ( .A(EAX_REG_26__SCAN_IN), .ZN(n6152) );
  AOI22_X1 U5394 ( .A1(n6597), .A2(UWORD_REG_10__SCAN_IN), .B1(n6123), .B2(
        DATAO_REG_26__SCAN_IN), .ZN(n4363) );
  OAI21_X1 U5395 ( .B1(n6152), .B2(n4419), .A(n4363), .ZN(U2897) );
  INV_X1 U5396 ( .A(EAX_REG_27__SCAN_IN), .ZN(n6154) );
  AOI22_X1 U5397 ( .A1(n6597), .A2(UWORD_REG_11__SCAN_IN), .B1(n6123), .B2(
        DATAO_REG_27__SCAN_IN), .ZN(n4364) );
  OAI21_X1 U5398 ( .B1(n6154), .B2(n4419), .A(n4364), .ZN(U2896) );
  INV_X1 U5399 ( .A(EAX_REG_28__SCAN_IN), .ZN(n6156) );
  AOI22_X1 U5400 ( .A1(n6597), .A2(UWORD_REG_12__SCAN_IN), .B1(n6123), .B2(
        DATAO_REG_28__SCAN_IN), .ZN(n4365) );
  OAI21_X1 U5401 ( .B1(n6156), .B2(n4419), .A(n4365), .ZN(U2895) );
  INV_X1 U5402 ( .A(EAX_REG_29__SCAN_IN), .ZN(n6158) );
  AOI22_X1 U5403 ( .A1(n6597), .A2(UWORD_REG_13__SCAN_IN), .B1(n6123), .B2(
        DATAO_REG_29__SCAN_IN), .ZN(n4366) );
  OAI21_X1 U5404 ( .B1(n6158), .B2(n4419), .A(n4366), .ZN(U2894) );
  INV_X1 U5405 ( .A(EAX_REG_24__SCAN_IN), .ZN(n6148) );
  AOI22_X1 U5406 ( .A1(n6597), .A2(UWORD_REG_8__SCAN_IN), .B1(n6123), .B2(
        DATAO_REG_24__SCAN_IN), .ZN(n4367) );
  OAI21_X1 U5407 ( .B1(n6148), .B2(n4419), .A(n4367), .ZN(U2899) );
  INV_X1 U5408 ( .A(EAX_REG_30__SCAN_IN), .ZN(n6160) );
  AOI22_X1 U5409 ( .A1(n6597), .A2(UWORD_REG_14__SCAN_IN), .B1(n6123), .B2(
        DATAO_REG_30__SCAN_IN), .ZN(n4368) );
  OAI21_X1 U5410 ( .B1(n6160), .B2(n4419), .A(n4368), .ZN(U2893) );
  INV_X1 U5411 ( .A(EBX_REG_0__SCAN_IN), .ZN(n4371) );
  XNOR2_X1 U5412 ( .A(n4370), .B(n4369), .ZN(n5201) );
  OAI222_X1 U5413 ( .A1(n5197), .A2(n5555), .B1(n4371), .B2(n6095), .C1(n5576), 
        .C2(n5201), .ZN(U2859) );
  NAND2_X1 U5414 ( .A1(n4372), .A2(n5691), .ZN(n4376) );
  NOR2_X1 U5415 ( .A1(n4373), .A2(n6221), .ZN(n4374) );
  AOI211_X1 U5416 ( .C1(PHYADDRPOINTER_REG_0__SCAN_IN), .C2(n4376), .A(n4375), 
        .B(n4374), .ZN(n4377) );
  OAI21_X1 U5417 ( .B1(n5201), .B2(n5697), .A(n4377), .ZN(U2986) );
  XNOR2_X1 U5418 ( .A(n4379), .B(n4378), .ZN(n4409) );
  XNOR2_X1 U5419 ( .A(n6086), .B(n4380), .ZN(n4404) );
  AOI21_X1 U5420 ( .B1(n4382), .B2(n4381), .A(n6331), .ZN(n4384) );
  INV_X1 U5421 ( .A(REIP_REG_1__SCAN_IN), .ZN(n6531) );
  NOR2_X1 U5422 ( .A1(n6335), .A2(n6531), .ZN(n4383) );
  AOI211_X1 U5423 ( .C1(n6323), .C2(n4404), .A(n4384), .B(n4383), .ZN(n4387)
         );
  NAND3_X1 U5424 ( .A1(n6297), .A2(n6331), .A3(n4385), .ZN(n4386) );
  OAI211_X1 U5425 ( .C1(n4409), .C2(n6300), .A(n4387), .B(n4386), .ZN(U3017)
         );
  NAND2_X1 U5426 ( .A1(n4475), .A2(n4388), .ZN(n4391) );
  INV_X1 U5427 ( .A(n4237), .ZN(n4467) );
  NAND2_X1 U5428 ( .A1(n4467), .A2(n4389), .ZN(n4390) );
  NAND2_X1 U5429 ( .A1(n4391), .A2(n4390), .ZN(n4447) );
  NOR2_X1 U5430 ( .A1(n4392), .A2(n4493), .ZN(n4393) );
  AND2_X1 U5431 ( .A1(n4423), .A2(n4393), .ZN(n4395) );
  OAI21_X1 U5432 ( .B1(n4447), .B2(n4395), .A(n4394), .ZN(n4396) );
  AND2_X1 U5433 ( .A1(n3138), .A2(n3164), .ZN(n4399) );
  NOR2_X1 U5434 ( .A1(n4399), .A2(n4398), .ZN(n4397) );
  NAND2_X2 U5435 ( .A1(n5397), .A2(n4397), .ZN(n5878) );
  INV_X1 U5436 ( .A(EAX_REG_0__SCAN_IN), .ZN(n6163) );
  INV_X1 U5437 ( .A(DATAI_0_), .ZN(n6732) );
  NOR2_X2 U5438 ( .A1(n6099), .A2(n6103), .ZN(n5305) );
  OAI222_X1 U5439 ( .A1(n5878), .A2(n5201), .B1(n5397), .B2(n6163), .C1(n6732), 
        .C2(n5305), .ZN(U2891) );
  OR2_X1 U5440 ( .A1(n4402), .A2(n4401), .ZN(n4403) );
  AND2_X1 U5441 ( .A1(n4400), .A2(n4403), .ZN(n6082) );
  INV_X1 U5442 ( .A(n6082), .ZN(n4410) );
  AOI22_X1 U5443 ( .A1(n6092), .A2(n4404), .B1(EBX_REG_1__SCAN_IN), .B2(n4150), 
        .ZN(n4405) );
  OAI21_X1 U5444 ( .B1(n4410), .B2(n5576), .A(n4405), .ZN(U2858) );
  AOI22_X1 U5445 ( .A1(n6239), .A2(PHYADDRPOINTER_REG_1__SCAN_IN), .B1(n2993), 
        .B2(REIP_REG_1__SCAN_IN), .ZN(n4406) );
  OAI21_X1 U5446 ( .B1(PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n6249), .A(n4406), 
        .ZN(n4407) );
  AOI21_X1 U5447 ( .B1(n6082), .B2(n6244), .A(n4407), .ZN(n4408) );
  OAI21_X1 U5448 ( .B1(n4409), .B2(n6221), .A(n4408), .ZN(U2985) );
  INV_X1 U5449 ( .A(DATAI_1_), .ZN(n6737) );
  INV_X1 U5450 ( .A(EAX_REG_1__SCAN_IN), .ZN(n6166) );
  OAI222_X1 U5451 ( .A1(n4410), .A2(n5878), .B1(n5305), .B2(n6737), .C1(n5397), 
        .C2(n6166), .ZN(U2890) );
  INV_X1 U5452 ( .A(EAX_REG_20__SCAN_IN), .ZN(n6140) );
  AOI22_X1 U5453 ( .A1(n6112), .A2(UWORD_REG_4__SCAN_IN), .B1(n6118), .B2(
        DATAO_REG_20__SCAN_IN), .ZN(n4411) );
  OAI21_X1 U5454 ( .B1(n6140), .B2(n4419), .A(n4411), .ZN(U2903) );
  INV_X1 U5455 ( .A(EAX_REG_17__SCAN_IN), .ZN(n6134) );
  AOI22_X1 U5456 ( .A1(n6112), .A2(UWORD_REG_1__SCAN_IN), .B1(n6118), .B2(
        DATAO_REG_17__SCAN_IN), .ZN(n4412) );
  OAI21_X1 U5457 ( .B1(n6134), .B2(n4419), .A(n4412), .ZN(U2906) );
  AOI22_X1 U5458 ( .A1(n6112), .A2(UWORD_REG_0__SCAN_IN), .B1(n6118), .B2(
        DATAO_REG_16__SCAN_IN), .ZN(n4413) );
  OAI21_X1 U5459 ( .B1(n3755), .B2(n4419), .A(n4413), .ZN(U2907) );
  INV_X1 U5460 ( .A(EAX_REG_21__SCAN_IN), .ZN(n6142) );
  AOI22_X1 U5461 ( .A1(n6112), .A2(UWORD_REG_5__SCAN_IN), .B1(n6118), .B2(
        DATAO_REG_21__SCAN_IN), .ZN(n4414) );
  OAI21_X1 U5462 ( .B1(n6142), .B2(n4419), .A(n4414), .ZN(U2902) );
  INV_X1 U5463 ( .A(EAX_REG_18__SCAN_IN), .ZN(n6136) );
  AOI22_X1 U5464 ( .A1(n6112), .A2(UWORD_REG_2__SCAN_IN), .B1(n6118), .B2(
        DATAO_REG_18__SCAN_IN), .ZN(n4415) );
  OAI21_X1 U5465 ( .B1(n6136), .B2(n4419), .A(n4415), .ZN(U2905) );
  INV_X1 U5466 ( .A(EAX_REG_19__SCAN_IN), .ZN(n6138) );
  AOI22_X1 U5467 ( .A1(n6112), .A2(UWORD_REG_3__SCAN_IN), .B1(n6118), .B2(
        DATAO_REG_19__SCAN_IN), .ZN(n4416) );
  OAI21_X1 U5468 ( .B1(n6138), .B2(n4419), .A(n4416), .ZN(U2904) );
  INV_X1 U5469 ( .A(EAX_REG_23__SCAN_IN), .ZN(n6146) );
  AOI22_X1 U5470 ( .A1(n6597), .A2(UWORD_REG_7__SCAN_IN), .B1(n6118), .B2(
        DATAO_REG_23__SCAN_IN), .ZN(n4417) );
  OAI21_X1 U5471 ( .B1(n6146), .B2(n4419), .A(n4417), .ZN(U2900) );
  INV_X1 U5472 ( .A(EAX_REG_22__SCAN_IN), .ZN(n6144) );
  AOI22_X1 U5473 ( .A1(n6597), .A2(UWORD_REG_6__SCAN_IN), .B1(n6118), .B2(
        DATAO_REG_22__SCAN_IN), .ZN(n4418) );
  OAI21_X1 U5474 ( .B1(n6144), .B2(n4419), .A(n4418), .ZN(U2901) );
  INV_X1 U5475 ( .A(FLUSH_REG_SCAN_IN), .ZN(n6696) );
  NAND2_X1 U5476 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n6696), .ZN(n4462) );
  INV_X1 U5477 ( .A(n4420), .ZN(n4461) );
  INV_X1 U5478 ( .A(n4422), .ZN(n4426) );
  INV_X1 U5479 ( .A(n4423), .ZN(n4424) );
  AND3_X1 U5480 ( .A1(n4237), .A2(n4168), .A3(n4424), .ZN(n4425) );
  NAND2_X1 U5481 ( .A1(n4426), .A2(n4425), .ZN(n5844) );
  NAND2_X1 U5482 ( .A1(n4799), .A2(n5844), .ZN(n4440) );
  NAND2_X1 U5483 ( .A1(n4428), .A2(n4427), .ZN(n4450) );
  CLKBUF_X1 U5484 ( .A(n4429), .Z(n5392) );
  MUX2_X1 U5485 ( .A(n4430), .B(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(n5392), 
        .Z(n4431) );
  NOR2_X1 U5486 ( .A1(n4431), .A2(n4420), .ZN(n4438) );
  NAND2_X1 U5487 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4433) );
  INV_X1 U5488 ( .A(n4433), .ZN(n4432) );
  MUX2_X1 U5489 ( .A(n4433), .B(n4432), .S(INSTQUEUERD_ADDR_REG_3__SCAN_IN), 
        .Z(n4436) );
  AOI21_X1 U5490 ( .B1(n5392), .B2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(n4434), 
        .ZN(n4435) );
  NOR2_X1 U5491 ( .A1(n3254), .A2(n4435), .ZN(n6584) );
  OAI22_X1 U5492 ( .A1(n6462), .A2(n4436), .B1(n6584), .B2(n4456), .ZN(n4437)
         );
  AOI21_X1 U5493 ( .B1(n4450), .B2(n4438), .A(n4437), .ZN(n4439) );
  NAND2_X1 U5494 ( .A1(n4440), .A2(n4439), .ZN(n6582) );
  INV_X1 U5495 ( .A(n4441), .ZN(n4443) );
  AOI21_X1 U5496 ( .B1(n6462), .B2(n4168), .A(n6519), .ZN(n4442) );
  INV_X1 U5497 ( .A(READY_N), .ZN(n6487) );
  OAI211_X1 U5498 ( .C1(n4443), .C2(n4442), .A(n4475), .B(n6487), .ZN(n4445)
         );
  NAND3_X1 U5499 ( .A1(n4446), .A2(n4445), .A3(n4444), .ZN(n4448) );
  MUX2_X1 U5500 ( .A(n6582), .B(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(n6459), 
        .Z(n6475) );
  XNOR2_X1 U5501 ( .A(n5392), .B(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4455)
         );
  NAND2_X1 U5502 ( .A1(n4450), .A2(n4455), .ZN(n4454) );
  INV_X1 U5503 ( .A(n6462), .ZN(n5417) );
  NAND2_X1 U5504 ( .A1(n5417), .A2(n4451), .ZN(n5841) );
  NAND2_X1 U5505 ( .A1(n5417), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4452) );
  MUX2_X1 U5506 ( .A(n5841), .B(n4452), .S(n3182), .Z(n4453) );
  OAI211_X1 U5507 ( .C1(n4456), .C2(n4455), .A(n4454), .B(n4453), .ZN(n4457)
         );
  AOI21_X1 U5508 ( .B1(n5833), .B2(n5844), .A(n4457), .ZN(n5389) );
  MUX2_X1 U5509 ( .A(n3182), .B(n5389), .S(n4469), .Z(n6470) );
  INV_X1 U5510 ( .A(n6470), .ZN(n4458) );
  AND2_X1 U5511 ( .A1(n4458), .A2(n5413), .ZN(n4459) );
  NAND2_X1 U5512 ( .A1(n6475), .A2(n4459), .ZN(n4460) );
  OAI21_X1 U5513 ( .B1(n4462), .B2(n4461), .A(n4460), .ZN(n6484) );
  INV_X1 U5514 ( .A(n4463), .ZN(n4464) );
  NAND2_X1 U5515 ( .A1(n6484), .A2(n4464), .ZN(n4477) );
  INV_X1 U5516 ( .A(n4864), .ZN(n4669) );
  NOR2_X1 U5517 ( .A1(n4465), .A2(n4669), .ZN(n4466) );
  XNOR2_X1 U5518 ( .A(n4466), .B(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n6041)
         );
  NAND2_X1 U5519 ( .A1(n4467), .A2(n5413), .ZN(n4468) );
  OR2_X1 U5520 ( .A1(n6041), .A2(n4468), .ZN(n5918) );
  MUX2_X1 U5521 ( .A(n4469), .B(FLUSH_REG_SCAN_IN), .S(STATE2_REG_1__SCAN_IN), 
        .Z(n4470) );
  OR2_X1 U5522 ( .A1(n4470), .A2(n3582), .ZN(n4471) );
  NAND2_X1 U5523 ( .A1(n5918), .A2(n4471), .ZN(n6483) );
  INV_X1 U5524 ( .A(n6483), .ZN(n4472) );
  NAND3_X1 U5525 ( .A1(n4477), .A2(n4472), .A3(n6696), .ZN(n4474) );
  OR2_X1 U5526 ( .A1(n6498), .A2(n4478), .ZN(n6579) );
  INV_X1 U5527 ( .A(n6579), .ZN(n4473) );
  NAND2_X1 U5528 ( .A1(n4474), .A2(n4473), .ZN(n4476) );
  NAND2_X1 U5529 ( .A1(n4476), .A2(n4867), .ZN(n6345) );
  INV_X1 U5530 ( .A(n4477), .ZN(n4479) );
  NOR3_X1 U5531 ( .A1(n4479), .A2(n4478), .A3(n6483), .ZN(n6493) );
  INV_X1 U5532 ( .A(n5412), .ZN(n4594) );
  NAND2_X1 U5533 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n6581), .ZN(n4535) );
  INV_X1 U5534 ( .A(n4535), .ZN(n5834) );
  OAI22_X1 U5535 ( .A1(n4861), .A2(n5835), .B1(n4594), .B2(n5834), .ZN(n4480)
         );
  OAI21_X1 U5536 ( .B1(n6493), .B2(n4480), .A(n6345), .ZN(n4481) );
  OAI21_X1 U5537 ( .B1(n6345), .B2(n5031), .A(n4481), .ZN(U3465) );
  OR2_X1 U5538 ( .A1(n5831), .A2(n4533), .ZN(n4532) );
  INV_X1 U5539 ( .A(n4532), .ZN(n4491) );
  AOI21_X1 U5540 ( .B1(n4491), .B2(n5827), .A(n5697), .ZN(n4486) );
  AND2_X1 U5541 ( .A1(n5826), .A2(n6657), .ZN(n5128) );
  AND2_X1 U5542 ( .A1(n4799), .A2(n5412), .ZN(n5034) );
  NAND2_X1 U5543 ( .A1(n5833), .A2(n6074), .ZN(n6352) );
  INV_X1 U5544 ( .A(n6352), .ZN(n4720) );
  INV_X1 U5545 ( .A(n4485), .ZN(n4520) );
  AOI21_X1 U5546 ( .B1(n5034), .B2(n4720), .A(n4520), .ZN(n4490) );
  OAI21_X1 U5547 ( .B1(n4486), .B2(n5128), .A(n4490), .ZN(n4487) );
  AOI21_X1 U5548 ( .B1(n5031), .B2(STATE2_REG_3__SCAN_IN), .A(n4867), .ZN(
        n5041) );
  OAI211_X1 U5549 ( .C1(n4489), .C2(n5826), .A(n4487), .B(n5041), .ZN(n4488)
         );
  INV_X1 U5550 ( .A(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n4496) );
  NAND2_X1 U5551 ( .A1(n6244), .A2(DATAI_22_), .ZN(n6386) );
  INV_X1 U5552 ( .A(n6386), .ZN(n6417) );
  INV_X1 U5553 ( .A(DATAI_6_), .ZN(n6715) );
  NOR2_X1 U5554 ( .A1(n6715), .A2(n4867), .ZN(n6420) );
  INV_X1 U5555 ( .A(n4489), .ZN(n4712) );
  OAI22_X1 U5556 ( .A1(n4490), .A2(n5835), .B1(n6497), .B2(n4712), .ZN(n4517)
         );
  AOI22_X1 U5557 ( .A1(n5137), .A2(n6417), .B1(n6420), .B2(n4517), .ZN(n4495)
         );
  NAND2_X1 U5558 ( .A1(n4491), .A2(n4795), .ZN(n4744) );
  NAND2_X1 U5559 ( .A1(n6244), .A2(DATAI_30_), .ZN(n6425) );
  INV_X1 U5560 ( .A(n6425), .ZN(n6383) );
  NOR2_X2 U5561 ( .A1(n4519), .A2(n4493), .ZN(n6415) );
  AOI22_X1 U5562 ( .A1(n4521), .A2(n6383), .B1(n4520), .B2(n6415), .ZN(n4494)
         );
  OAI211_X1 U5563 ( .C1(n4525), .C2(n4496), .A(n4495), .B(n4494), .ZN(U3146)
         );
  INV_X1 U5564 ( .A(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n4499) );
  NAND2_X1 U5565 ( .A1(n6244), .A2(DATAI_21_), .ZN(n6449) );
  INV_X1 U5566 ( .A(n6449), .ZN(n6412) );
  INV_X1 U5567 ( .A(DATAI_5_), .ZN(n6719) );
  NOR2_X2 U5568 ( .A1(n6719), .A2(n4867), .ZN(n6453) );
  AOI22_X1 U5569 ( .A1(n5137), .A2(n6412), .B1(n6453), .B2(n4517), .ZN(n4498)
         );
  NAND2_X1 U5570 ( .A1(n6244), .A2(DATAI_29_), .ZN(n6458) );
  INV_X1 U5571 ( .A(n6458), .ZN(n6380) );
  NOR2_X2 U5572 ( .A1(n4519), .A2(n3138), .ZN(n6411) );
  AOI22_X1 U5573 ( .A1(n4521), .A2(n6380), .B1(n4520), .B2(n6411), .ZN(n4497)
         );
  OAI211_X1 U5574 ( .C1(n4525), .C2(n4499), .A(n4498), .B(n4497), .ZN(U3145)
         );
  INV_X1 U5575 ( .A(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n4502) );
  NAND2_X1 U5576 ( .A1(n6244), .A2(DATAI_18_), .ZN(n6371) );
  INV_X1 U5577 ( .A(n6371), .ZN(n4947) );
  INV_X1 U5578 ( .A(DATAI_2_), .ZN(n6729) );
  NOR2_X1 U5579 ( .A1(n6729), .A2(n4867), .ZN(n6366) );
  AOI22_X1 U5580 ( .A1(n5137), .A2(n4947), .B1(n6366), .B2(n4517), .ZN(n4501)
         );
  INV_X1 U5581 ( .A(DATAI_26_), .ZN(n6769) );
  NOR2_X1 U5582 ( .A1(n5697), .A2(n6769), .ZN(n6368) );
  NOR2_X2 U5583 ( .A1(n4519), .A2(n3298), .ZN(n6367) );
  AOI22_X1 U5584 ( .A1(n4521), .A2(n6368), .B1(n4520), .B2(n6367), .ZN(n4500)
         );
  OAI211_X1 U5585 ( .C1(n4525), .C2(n4502), .A(n4501), .B(n4500), .ZN(U3142)
         );
  INV_X1 U5586 ( .A(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n4505) );
  NAND2_X1 U5587 ( .A1(n6244), .A2(DATAI_23_), .ZN(n6396) );
  INV_X1 U5588 ( .A(n6396), .ZN(n4952) );
  INV_X1 U5589 ( .A(DATAI_7_), .ZN(n6713) );
  NOR2_X1 U5590 ( .A1(n6713), .A2(n4867), .ZN(n6388) );
  AOI22_X1 U5591 ( .A1(n5137), .A2(n4952), .B1(n6388), .B2(n4517), .ZN(n4504)
         );
  INV_X1 U5592 ( .A(DATAI_31_), .ZN(n6744) );
  NOR2_X1 U5593 ( .A1(n5697), .A2(n6744), .ZN(n6392) );
  NOR2_X2 U5594 ( .A1(n4519), .A2(n5396), .ZN(n6390) );
  AOI22_X1 U5595 ( .A1(n4521), .A2(n6392), .B1(n4520), .B2(n6390), .ZN(n4503)
         );
  OAI211_X1 U5596 ( .C1(n4525), .C2(n4505), .A(n4504), .B(n4503), .ZN(U3147)
         );
  INV_X1 U5597 ( .A(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n4508) );
  NAND2_X1 U5598 ( .A1(n6244), .A2(DATAI_19_), .ZN(n6375) );
  INV_X1 U5599 ( .A(n6375), .ZN(n6406) );
  INV_X1 U5600 ( .A(DATAI_3_), .ZN(n6802) );
  NOR2_X1 U5601 ( .A1(n6802), .A2(n4867), .ZN(n6407) );
  AOI22_X1 U5602 ( .A1(n5137), .A2(n6406), .B1(n6407), .B2(n4517), .ZN(n4507)
         );
  NAND2_X1 U5603 ( .A1(n6244), .A2(DATAI_27_), .ZN(n6410) );
  INV_X1 U5604 ( .A(n6410), .ZN(n6372) );
  NOR2_X2 U5605 ( .A1(n4519), .A2(n3121), .ZN(n6405) );
  AOI22_X1 U5606 ( .A1(n4521), .A2(n6372), .B1(n4520), .B2(n6405), .ZN(n4506)
         );
  OAI211_X1 U5607 ( .C1(n4525), .C2(n4508), .A(n4507), .B(n4506), .ZN(U3143)
         );
  INV_X1 U5608 ( .A(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n4512) );
  NAND2_X1 U5609 ( .A1(n6244), .A2(DATAI_20_), .ZN(n6441) );
  INV_X1 U5610 ( .A(n6441), .ZN(n4958) );
  INV_X1 U5611 ( .A(DATAI_4_), .ZN(n6721) );
  NOR2_X2 U5612 ( .A1(n6721), .A2(n4867), .ZN(n6443) );
  AOI22_X1 U5613 ( .A1(n5137), .A2(n4958), .B1(n6443), .B2(n4517), .ZN(n4511)
         );
  NAND2_X1 U5614 ( .A1(n6244), .A2(DATAI_28_), .ZN(n6446) );
  INV_X1 U5615 ( .A(n6446), .ZN(n6377) );
  NOR2_X2 U5616 ( .A1(n4519), .A2(n4509), .ZN(n6376) );
  AOI22_X1 U5617 ( .A1(n4521), .A2(n6377), .B1(n4520), .B2(n6376), .ZN(n4510)
         );
  OAI211_X1 U5618 ( .C1(n4525), .C2(n4512), .A(n4511), .B(n4510), .ZN(U3144)
         );
  INV_X1 U5619 ( .A(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n4516) );
  NAND2_X1 U5620 ( .A1(n6244), .A2(DATAI_17_), .ZN(n6434) );
  INV_X1 U5621 ( .A(n6434), .ZN(n6402) );
  NOR2_X2 U5622 ( .A1(n6737), .A2(n4867), .ZN(n6436) );
  AOI22_X1 U5623 ( .A1(n5137), .A2(n6402), .B1(n6436), .B2(n4517), .ZN(n4515)
         );
  NAND2_X1 U5624 ( .A1(n6244), .A2(DATAI_25_), .ZN(n6439) );
  INV_X1 U5625 ( .A(n6439), .ZN(n6363) );
  NOR2_X2 U5626 ( .A1(n4519), .A2(n4513), .ZN(n6401) );
  AOI22_X1 U5627 ( .A1(n4521), .A2(n6363), .B1(n4520), .B2(n6401), .ZN(n4514)
         );
  OAI211_X1 U5628 ( .C1(n4525), .C2(n4516), .A(n4515), .B(n4514), .ZN(U3141)
         );
  INV_X1 U5629 ( .A(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n4524) );
  NAND2_X1 U5630 ( .A1(n6244), .A2(DATAI_16_), .ZN(n6427) );
  INV_X1 U5631 ( .A(n6427), .ZN(n6398) );
  NOR2_X2 U5632 ( .A1(n6732), .A2(n4867), .ZN(n6429) );
  AOI22_X1 U5633 ( .A1(n5137), .A2(n6398), .B1(n6429), .B2(n4517), .ZN(n4523)
         );
  NAND2_X1 U5634 ( .A1(n6244), .A2(DATAI_24_), .ZN(n6432) );
  INV_X1 U5635 ( .A(n6432), .ZN(n6360) );
  NOR2_X2 U5636 ( .A1(n4519), .A2(n4518), .ZN(n6397) );
  AOI22_X1 U5637 ( .A1(n4521), .A2(n6360), .B1(n4520), .B2(n6397), .ZN(n4522)
         );
  OAI211_X1 U5638 ( .C1(n4525), .C2(n4524), .A(n4523), .B(n4522), .ZN(U3140)
         );
  CLKBUF_X1 U5639 ( .A(n4526), .Z(n4527) );
  OAI21_X1 U5640 ( .B1(n4527), .B2(n4528), .A(n4562), .ZN(n6053) );
  AND2_X1 U5641 ( .A1(n4578), .A2(n4529), .ZN(n4530) );
  NOR2_X1 U5642 ( .A1(n4567), .A2(n4530), .ZN(n6322) );
  AOI22_X1 U5643 ( .A1(n6092), .A2(n6322), .B1(EBX_REG_3__SCAN_IN), .B2(n4150), 
        .ZN(n4531) );
  OAI21_X1 U5644 ( .B1(n6053), .B2(n5576), .A(n4531), .ZN(U2856) );
  NAND2_X1 U5645 ( .A1(n4862), .A2(STATEBS16_REG_SCAN_IN), .ZN(n5038) );
  INV_X1 U5646 ( .A(n4601), .ZN(n4534) );
  AND2_X1 U5647 ( .A1(n5827), .A2(STATEBS16_REG_SCAN_IN), .ZN(n4914) );
  NAND2_X1 U5648 ( .A1(n4668), .A2(n4914), .ZN(n4549) );
  NAND3_X1 U5649 ( .A1(n5038), .A2(n4534), .A3(n4549), .ZN(n4916) );
  AOI222_X1 U5650 ( .A1(n4916), .A2(n5826), .B1(n4750), .B2(n5128), .C1(n4799), 
        .C2(n4535), .ZN(n4538) );
  INV_X1 U5651 ( .A(n6345), .ZN(n4537) );
  NAND2_X1 U5652 ( .A1(n4537), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n4536) );
  OAI21_X1 U5653 ( .B1(n4538), .B2(n4537), .A(n4536), .ZN(U3462) );
  OAI21_X1 U5654 ( .B1(n4541), .B2(n4540), .A(n4539), .ZN(n4542) );
  INV_X1 U5655 ( .A(n4542), .ZN(n6325) );
  NAND2_X1 U5656 ( .A1(n6325), .A2(n6243), .ZN(n4547) );
  INV_X1 U5657 ( .A(REIP_REG_3__SCAN_IN), .ZN(n4543) );
  NOR2_X1 U5658 ( .A1(n6335), .A2(n4543), .ZN(n6321) );
  NOR2_X1 U5659 ( .A1(n5691), .A2(n4544), .ZN(n4545) );
  AOI211_X1 U5660 ( .C1(n6217), .C2(n6055), .A(n6321), .B(n4545), .ZN(n4546)
         );
  OAI211_X1 U5661 ( .C1(n5697), .C2(n6053), .A(n4547), .B(n4546), .ZN(U2983)
         );
  INV_X1 U5662 ( .A(n4799), .ZN(n6050) );
  NAND3_X1 U5663 ( .A1(n6050), .A2(n4720), .A3(n5412), .ZN(n4548) );
  AND2_X1 U5664 ( .A1(n4548), .A2(n4554), .ZN(n4553) );
  INV_X1 U5665 ( .A(n4553), .ZN(n4551) );
  NAND2_X1 U5666 ( .A1(n5826), .A2(n4549), .ZN(n4552) );
  AOI21_X1 U5667 ( .B1(n6347), .B2(n5835), .A(n4921), .ZN(n4550) );
  OAI21_X1 U5668 ( .B1(n4551), .B2(n4552), .A(n4550), .ZN(n6421) );
  OAI22_X1 U5669 ( .A1(n4553), .A2(n4552), .B1(n6497), .B2(n6347), .ZN(n6419)
         );
  AOI22_X1 U5670 ( .A1(INSTQUEUE_REG_7__4__SCAN_IN), .A2(n6421), .B1(n6443), 
        .B2(n6419), .ZN(n4556) );
  INV_X1 U5671 ( .A(n4554), .ZN(n6416) );
  AOI22_X1 U5672 ( .A1(n6418), .A2(n4958), .B1(n6416), .B2(n6376), .ZN(n4555)
         );
  OAI211_X1 U5673 ( .C1(n6446), .C2(n6424), .A(n4556), .B(n4555), .ZN(U3080)
         );
  INV_X1 U5674 ( .A(n6368), .ZN(n5158) );
  AOI22_X1 U5675 ( .A1(INSTQUEUE_REG_7__2__SCAN_IN), .A2(n6421), .B1(n6366), 
        .B2(n6419), .ZN(n4558) );
  AOI22_X1 U5676 ( .A1(n6418), .A2(n4947), .B1(n6416), .B2(n6367), .ZN(n4557)
         );
  OAI211_X1 U5677 ( .C1(n5158), .C2(n6424), .A(n4558), .B(n4557), .ZN(U3078)
         );
  INV_X1 U5678 ( .A(n6392), .ZN(n5153) );
  AOI22_X1 U5679 ( .A1(INSTQUEUE_REG_7__7__SCAN_IN), .A2(n6421), .B1(n6388), 
        .B2(n6419), .ZN(n4560) );
  AOI22_X1 U5680 ( .A1(n6418), .A2(n4952), .B1(n6416), .B2(n6390), .ZN(n4559)
         );
  OAI211_X1 U5681 ( .C1(n5153), .C2(n6424), .A(n4560), .B(n4559), .ZN(U3083)
         );
  INV_X1 U5682 ( .A(EAX_REG_3__SCAN_IN), .ZN(n6172) );
  OAI222_X1 U5683 ( .A1(n6053), .A2(n5878), .B1(n5305), .B2(n6802), .C1(n5397), 
        .C2(n6172), .ZN(U2888) );
  AND2_X1 U5684 ( .A1(n4562), .A2(n4561), .ZN(n4564) );
  CLKBUF_X1 U5685 ( .A(n4563), .Z(n4585) );
  OR2_X1 U5686 ( .A1(n4564), .A2(n4585), .ZN(n6234) );
  CLKBUF_X1 U5687 ( .A(n4565), .Z(n4587) );
  NOR2_X1 U5688 ( .A1(n4567), .A2(n4566), .ZN(n4568) );
  OR2_X1 U5689 ( .A1(n4587), .A2(n4568), .ZN(n6313) );
  INV_X1 U5690 ( .A(n6313), .ZN(n4569) );
  AOI22_X1 U5691 ( .A1(n6092), .A2(n4569), .B1(EBX_REG_4__SCAN_IN), .B2(n4150), 
        .ZN(n4570) );
  OAI21_X1 U5692 ( .B1(n6234), .B2(n5576), .A(n4570), .ZN(U2855) );
  INV_X1 U5693 ( .A(n4571), .ZN(n4572) );
  NOR2_X1 U5694 ( .A1(n4573), .A2(n4572), .ZN(n4574) );
  AOI21_X1 U5695 ( .B1(n4574), .B2(n4400), .A(n4527), .ZN(n6245) );
  NAND2_X1 U5696 ( .A1(n4576), .A2(n4575), .ZN(n4577) );
  NAND2_X1 U5697 ( .A1(n4578), .A2(n4577), .ZN(n6336) );
  OAI22_X1 U5698 ( .A1(n5555), .A2(n6336), .B1(n4579), .B2(n6095), .ZN(n4580)
         );
  AOI21_X1 U5699 ( .B1(n6245), .B2(n4149), .A(n4580), .ZN(n4581) );
  INV_X1 U5700 ( .A(n4581), .ZN(U2857) );
  INV_X1 U5701 ( .A(EAX_REG_4__SCAN_IN), .ZN(n6175) );
  OAI222_X1 U5702 ( .A1(n6234), .A2(n5878), .B1(n5305), .B2(n6721), .C1(n5397), 
        .C2(n6175), .ZN(U2887) );
  INV_X1 U5703 ( .A(n6245), .ZN(n4582) );
  INV_X1 U5704 ( .A(EAX_REG_2__SCAN_IN), .ZN(n6169) );
  OAI222_X1 U5705 ( .A1(n4582), .A2(n5878), .B1(n5305), .B2(n6729), .C1(n5397), 
        .C2(n6169), .ZN(U2889) );
  OAI21_X1 U5706 ( .B1(n4585), .B2(n4584), .A(n4790), .ZN(n5211) );
  INV_X1 U5707 ( .A(n4586), .ZN(n4590) );
  INV_X1 U5708 ( .A(n4587), .ZN(n4589) );
  INV_X1 U5709 ( .A(n4588), .ZN(n4792) );
  AOI21_X1 U5710 ( .B1(n4590), .B2(n4589), .A(n4792), .ZN(n6307) );
  AOI22_X1 U5711 ( .A1(n6307), .A2(n6092), .B1(EBX_REG_5__SCAN_IN), .B2(n4150), 
        .ZN(n4591) );
  OAI21_X1 U5712 ( .B1(n5211), .B2(n5576), .A(n4591), .ZN(U2854) );
  INV_X1 U5713 ( .A(EAX_REG_5__SCAN_IN), .ZN(n6178) );
  OAI222_X1 U5714 ( .A1(n5211), .A2(n5878), .B1(n5305), .B2(n6719), .C1(n5397), 
        .C2(n6178), .ZN(U2886) );
  NAND3_X1 U5715 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(n6468), .ZN(n4978) );
  AOI21_X1 U5716 ( .B1(n4601), .B2(n4914), .A(n5835), .ZN(n4596) );
  INV_X1 U5717 ( .A(n6074), .ZN(n5829) );
  OR2_X1 U5718 ( .A1(n5833), .A2(n5829), .ZN(n4798) );
  INV_X1 U5719 ( .A(n4798), .ZN(n4592) );
  NAND2_X1 U5720 ( .A1(n4592), .A2(n4799), .ZN(n4986) );
  INV_X1 U5721 ( .A(n4918), .ZN(n4593) );
  NAND2_X1 U5722 ( .A1(n4593), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6447) );
  OAI21_X1 U5723 ( .B1(n4986), .B2(n4594), .A(n6447), .ZN(n4598) );
  NAND2_X1 U5724 ( .A1(n4596), .A2(n4598), .ZN(n4595) );
  OAI21_X1 U5725 ( .B1(n4978), .B2(n6497), .A(n4595), .ZN(n6452) );
  INV_X1 U5726 ( .A(n6452), .ZN(n4614) );
  INV_X1 U5727 ( .A(n6407), .ZN(n5140) );
  INV_X1 U5728 ( .A(n4596), .ZN(n4599) );
  AOI21_X1 U5729 ( .B1(n5835), .B2(n4978), .A(n4921), .ZN(n4597) );
  OAI21_X1 U5730 ( .B1(n4599), .B2(n4598), .A(n4597), .ZN(n6454) );
  NOR2_X1 U5731 ( .A1(n6457), .A2(n6410), .ZN(n4603) );
  INV_X1 U5732 ( .A(n6405), .ZN(n5055) );
  OAI22_X1 U5733 ( .A1(n6450), .A2(n6375), .B1(n5055), .B2(n6447), .ZN(n4602)
         );
  AOI211_X1 U5734 ( .C1(n6454), .C2(INSTQUEUE_REG_11__3__SCAN_IN), .A(n4603), 
        .B(n4602), .ZN(n4604) );
  OAI21_X1 U5735 ( .B1(n4614), .B2(n5140), .A(n4604), .ZN(U3111) );
  INV_X1 U5736 ( .A(n6366), .ZN(n5157) );
  NOR2_X1 U5737 ( .A1(n6457), .A2(n5158), .ZN(n4606) );
  INV_X1 U5738 ( .A(n6367), .ZN(n5051) );
  OAI22_X1 U5739 ( .A1(n6450), .A2(n6371), .B1(n5051), .B2(n6447), .ZN(n4605)
         );
  AOI211_X1 U5740 ( .C1(n6454), .C2(INSTQUEUE_REG_11__2__SCAN_IN), .A(n4606), 
        .B(n4605), .ZN(n4607) );
  OAI21_X1 U5741 ( .B1(n4614), .B2(n5157), .A(n4607), .ZN(U3110) );
  INV_X1 U5742 ( .A(n6388), .ZN(n5152) );
  NOR2_X1 U5743 ( .A1(n6457), .A2(n5153), .ZN(n4609) );
  INV_X1 U5744 ( .A(n6390), .ZN(n5072) );
  OAI22_X1 U5745 ( .A1(n6450), .A2(n6396), .B1(n5072), .B2(n6447), .ZN(n4608)
         );
  AOI211_X1 U5746 ( .C1(n6454), .C2(INSTQUEUE_REG_11__7__SCAN_IN), .A(n4609), 
        .B(n4608), .ZN(n4610) );
  OAI21_X1 U5747 ( .B1(n4614), .B2(n5152), .A(n4610), .ZN(U3115) );
  INV_X1 U5748 ( .A(n6420), .ZN(n5148) );
  NOR2_X1 U5749 ( .A1(n6457), .A2(n6425), .ZN(n4612) );
  INV_X1 U5750 ( .A(n6415), .ZN(n5065) );
  OAI22_X1 U5751 ( .A1(n6450), .A2(n6386), .B1(n5065), .B2(n6447), .ZN(n4611)
         );
  AOI211_X1 U5752 ( .C1(n6454), .C2(INSTQUEUE_REG_11__6__SCAN_IN), .A(n4612), 
        .B(n4611), .ZN(n4613) );
  OAI21_X1 U5753 ( .B1(n4614), .B2(n5148), .A(n4613), .ZN(U3114) );
  INV_X1 U5754 ( .A(n5827), .ZN(n4667) );
  NAND2_X1 U5755 ( .A1(n5831), .A2(n4667), .ZN(n4640) );
  OR2_X1 U5756 ( .A1(n5833), .A2(n6074), .ZN(n5096) );
  NAND3_X1 U5757 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n6468), .A3(n6464), .ZN(n5089) );
  NOR2_X1 U5758 ( .A1(n5031), .A2(n5089), .ZN(n4637) );
  AOI21_X1 U5759 ( .B1(n5034), .B2(n5139), .A(n4637), .ZN(n4619) );
  INV_X1 U5760 ( .A(n4619), .ZN(n4617) );
  INV_X1 U5761 ( .A(n4620), .ZN(n4615) );
  OAI21_X1 U5762 ( .B1(n4615), .B2(n6657), .A(n5826), .ZN(n4618) );
  AOI21_X1 U5763 ( .B1(n5835), .B2(n5089), .A(n4921), .ZN(n4616) );
  OAI21_X1 U5764 ( .B1(n4617), .B2(n4618), .A(n4616), .ZN(n4636) );
  OAI22_X1 U5765 ( .A1(n4619), .A2(n4618), .B1(n6497), .B2(n5089), .ZN(n4635)
         );
  AOI22_X1 U5766 ( .A1(INSTQUEUE_REG_9__2__SCAN_IN), .A2(n4636), .B1(n6366), 
        .B2(n4635), .ZN(n4622) );
  AOI22_X1 U5767 ( .A1(n5017), .A2(n4947), .B1(n6367), .B2(n4637), .ZN(n4621)
         );
  OAI211_X1 U5768 ( .C1(n5158), .C2(n5127), .A(n4622), .B(n4621), .ZN(U3094)
         );
  AOI22_X1 U5769 ( .A1(INSTQUEUE_REG_9__4__SCAN_IN), .A2(n4636), .B1(n6443), 
        .B2(n4635), .ZN(n4624) );
  AOI22_X1 U5770 ( .A1(n5017), .A2(n4958), .B1(n6376), .B2(n4637), .ZN(n4623)
         );
  OAI211_X1 U5771 ( .C1(n6446), .C2(n5127), .A(n4624), .B(n4623), .ZN(U3096)
         );
  AOI22_X1 U5772 ( .A1(INSTQUEUE_REG_9__5__SCAN_IN), .A2(n4636), .B1(n6453), 
        .B2(n4635), .ZN(n4626) );
  AOI22_X1 U5773 ( .A1(n5017), .A2(n6412), .B1(n6411), .B2(n4637), .ZN(n4625)
         );
  OAI211_X1 U5774 ( .C1(n6458), .C2(n5127), .A(n4626), .B(n4625), .ZN(U3097)
         );
  AOI22_X1 U5775 ( .A1(INSTQUEUE_REG_9__7__SCAN_IN), .A2(n4636), .B1(n6388), 
        .B2(n4635), .ZN(n4628) );
  AOI22_X1 U5776 ( .A1(n5017), .A2(n4952), .B1(n6390), .B2(n4637), .ZN(n4627)
         );
  OAI211_X1 U5777 ( .C1(n5153), .C2(n5127), .A(n4628), .B(n4627), .ZN(U3099)
         );
  AOI22_X1 U5778 ( .A1(INSTQUEUE_REG_9__6__SCAN_IN), .A2(n4636), .B1(n6420), 
        .B2(n4635), .ZN(n4630) );
  AOI22_X1 U5779 ( .A1(n5017), .A2(n6417), .B1(n6415), .B2(n4637), .ZN(n4629)
         );
  OAI211_X1 U5780 ( .C1(n6425), .C2(n5127), .A(n4630), .B(n4629), .ZN(U3098)
         );
  AOI22_X1 U5781 ( .A1(INSTQUEUE_REG_9__3__SCAN_IN), .A2(n4636), .B1(n6407), 
        .B2(n4635), .ZN(n4632) );
  AOI22_X1 U5782 ( .A1(n5017), .A2(n6406), .B1(n6405), .B2(n4637), .ZN(n4631)
         );
  OAI211_X1 U5783 ( .C1(n6410), .C2(n5127), .A(n4632), .B(n4631), .ZN(U3095)
         );
  AOI22_X1 U5784 ( .A1(INSTQUEUE_REG_9__0__SCAN_IN), .A2(n4636), .B1(n6429), 
        .B2(n4635), .ZN(n4634) );
  AOI22_X1 U5785 ( .A1(n5017), .A2(n6398), .B1(n6397), .B2(n4637), .ZN(n4633)
         );
  OAI211_X1 U5786 ( .C1(n6432), .C2(n5127), .A(n4634), .B(n4633), .ZN(U3092)
         );
  AOI22_X1 U5787 ( .A1(INSTQUEUE_REG_9__1__SCAN_IN), .A2(n4636), .B1(n6436), 
        .B2(n4635), .ZN(n4639) );
  AOI22_X1 U5788 ( .A1(n5017), .A2(n6402), .B1(n6401), .B2(n4637), .ZN(n4638)
         );
  OAI211_X1 U5789 ( .C1(n6439), .C2(n5127), .A(n4639), .B(n4638), .ZN(U3093)
         );
  INV_X1 U5790 ( .A(n4640), .ZN(n4641) );
  INV_X1 U5791 ( .A(n4647), .ZN(n4642) );
  OAI21_X1 U5792 ( .B1(n4642), .B2(n6657), .A(n5826), .ZN(n4645) );
  NOR2_X1 U5793 ( .A1(n4799), .A2(n5096), .ZN(n5135) );
  NAND3_X1 U5794 ( .A1(n6474), .A2(n6468), .A3(n6464), .ZN(n5130) );
  NOR2_X1 U5795 ( .A1(n5031), .A2(n5130), .ZN(n4664) );
  AOI21_X1 U5796 ( .B1(n5135), .B2(n5412), .A(n4664), .ZN(n4646) );
  INV_X1 U5797 ( .A(n4646), .ZN(n4644) );
  AOI21_X1 U5798 ( .B1(n5835), .B2(n5130), .A(n4921), .ZN(n4643) );
  OAI21_X1 U5799 ( .B1(n4645), .B2(n4644), .A(n4643), .ZN(n4663) );
  OAI22_X1 U5800 ( .A1(n4646), .A2(n4645), .B1(n6497), .B2(n5130), .ZN(n4662)
         );
  AOI22_X1 U5801 ( .A1(INSTQUEUE_REG_1__3__SCAN_IN), .A2(n4663), .B1(n6407), 
        .B2(n4662), .ZN(n4649) );
  AOI22_X1 U5802 ( .A1(n4838), .A2(n6406), .B1(n6405), .B2(n4664), .ZN(n4648)
         );
  OAI211_X1 U5803 ( .C1(n6410), .C2(n5178), .A(n4649), .B(n4648), .ZN(U3031)
         );
  AOI22_X1 U5804 ( .A1(INSTQUEUE_REG_1__1__SCAN_IN), .A2(n4663), .B1(n6436), 
        .B2(n4662), .ZN(n4651) );
  AOI22_X1 U5805 ( .A1(n4838), .A2(n6402), .B1(n6401), .B2(n4664), .ZN(n4650)
         );
  OAI211_X1 U5806 ( .C1(n6439), .C2(n5178), .A(n4651), .B(n4650), .ZN(U3029)
         );
  AOI22_X1 U5807 ( .A1(INSTQUEUE_REG_1__7__SCAN_IN), .A2(n4663), .B1(n6388), 
        .B2(n4662), .ZN(n4653) );
  AOI22_X1 U5808 ( .A1(n4838), .A2(n4952), .B1(n6390), .B2(n4664), .ZN(n4652)
         );
  OAI211_X1 U5809 ( .C1(n5153), .C2(n5178), .A(n4653), .B(n4652), .ZN(U3035)
         );
  AOI22_X1 U5810 ( .A1(INSTQUEUE_REG_1__5__SCAN_IN), .A2(n4663), .B1(n6453), 
        .B2(n4662), .ZN(n4655) );
  AOI22_X1 U5811 ( .A1(n4838), .A2(n6412), .B1(n6411), .B2(n4664), .ZN(n4654)
         );
  OAI211_X1 U5812 ( .C1(n6458), .C2(n5178), .A(n4655), .B(n4654), .ZN(U3033)
         );
  AOI22_X1 U5813 ( .A1(INSTQUEUE_REG_1__4__SCAN_IN), .A2(n4663), .B1(n6443), 
        .B2(n4662), .ZN(n4657) );
  AOI22_X1 U5814 ( .A1(n4838), .A2(n4958), .B1(n6376), .B2(n4664), .ZN(n4656)
         );
  OAI211_X1 U5815 ( .C1(n6446), .C2(n5178), .A(n4657), .B(n4656), .ZN(U3032)
         );
  AOI22_X1 U5816 ( .A1(INSTQUEUE_REG_1__6__SCAN_IN), .A2(n4663), .B1(n6420), 
        .B2(n4662), .ZN(n4659) );
  AOI22_X1 U5817 ( .A1(n4838), .A2(n6417), .B1(n6415), .B2(n4664), .ZN(n4658)
         );
  OAI211_X1 U5818 ( .C1(n6425), .C2(n5178), .A(n4659), .B(n4658), .ZN(U3034)
         );
  AOI22_X1 U5819 ( .A1(INSTQUEUE_REG_1__2__SCAN_IN), .A2(n4663), .B1(n6366), 
        .B2(n4662), .ZN(n4661) );
  AOI22_X1 U5820 ( .A1(n4838), .A2(n4947), .B1(n6367), .B2(n4664), .ZN(n4660)
         );
  OAI211_X1 U5821 ( .C1(n5158), .C2(n5178), .A(n4661), .B(n4660), .ZN(U3030)
         );
  AOI22_X1 U5822 ( .A1(INSTQUEUE_REG_1__0__SCAN_IN), .A2(n4663), .B1(n6429), 
        .B2(n4662), .ZN(n4666) );
  AOI22_X1 U5823 ( .A1(n4838), .A2(n6398), .B1(n6397), .B2(n4664), .ZN(n4665)
         );
  OAI211_X1 U5824 ( .C1(n6432), .C2(n5178), .A(n4666), .B(n4665), .ZN(U3028)
         );
  NAND2_X1 U5825 ( .A1(n4668), .A2(n4667), .ZN(n4675) );
  OAI21_X1 U5826 ( .B1(n4675), .B2(n6657), .A(n5826), .ZN(n4673) );
  INV_X1 U5827 ( .A(n4673), .ZN(n4753) );
  AND2_X1 U5828 ( .A1(n5033), .A2(n4669), .ZN(n4751) );
  NAND3_X1 U5829 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n6474), .A3(n6464), .ZN(n4755) );
  NOR2_X1 U5830 ( .A1(n5031), .A2(n4755), .ZN(n4704) );
  AOI21_X1 U5831 ( .B1(n4751), .B2(n5412), .A(n4704), .ZN(n4672) );
  INV_X1 U5832 ( .A(n4755), .ZN(n4670) );
  NOR2_X1 U5833 ( .A1(n5826), .A2(n4670), .ZN(n4671) );
  AOI211_X2 U5834 ( .C1(n4753), .C2(n4672), .A(n4921), .B(n4671), .ZN(n4710)
         );
  INV_X1 U5835 ( .A(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n4679) );
  OAI22_X1 U5836 ( .A1(n4673), .A2(n4672), .B1(n4755), .B2(n6497), .ZN(n4707)
         );
  INV_X1 U5837 ( .A(n4675), .ZN(n4674) );
  NOR2_X2 U5838 ( .A1(n4675), .A2(n4861), .ZN(n6391) );
  AOI22_X1 U5839 ( .A1(n6391), .A2(n6402), .B1(n6401), .B2(n4704), .ZN(n4676)
         );
  OAI21_X1 U5840 ( .B1(n6439), .B2(n4787), .A(n4676), .ZN(n4677) );
  AOI21_X1 U5841 ( .B1(n6436), .B2(n4707), .A(n4677), .ZN(n4678) );
  OAI21_X1 U5842 ( .B1(n4710), .B2(n4679), .A(n4678), .ZN(U3061) );
  INV_X1 U5843 ( .A(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n4683) );
  AOI22_X1 U5844 ( .A1(n6391), .A2(n6412), .B1(n6411), .B2(n4704), .ZN(n4680)
         );
  OAI21_X1 U5845 ( .B1(n6458), .B2(n4787), .A(n4680), .ZN(n4681) );
  AOI21_X1 U5846 ( .B1(n6453), .B2(n4707), .A(n4681), .ZN(n4682) );
  OAI21_X1 U5847 ( .B1(n4710), .B2(n4683), .A(n4682), .ZN(U3065) );
  INV_X1 U5848 ( .A(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n4687) );
  AOI22_X1 U5849 ( .A1(n6391), .A2(n6398), .B1(n6397), .B2(n4704), .ZN(n4684)
         );
  OAI21_X1 U5850 ( .B1(n6432), .B2(n4787), .A(n4684), .ZN(n4685) );
  AOI21_X1 U5851 ( .B1(n6429), .B2(n4707), .A(n4685), .ZN(n4686) );
  OAI21_X1 U5852 ( .B1(n4710), .B2(n4687), .A(n4686), .ZN(U3060) );
  INV_X1 U5853 ( .A(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n4691) );
  AOI22_X1 U5854 ( .A1(n6391), .A2(n6406), .B1(n6405), .B2(n4704), .ZN(n4688)
         );
  OAI21_X1 U5855 ( .B1(n6410), .B2(n4787), .A(n4688), .ZN(n4689) );
  AOI21_X1 U5856 ( .B1(n6407), .B2(n4707), .A(n4689), .ZN(n4690) );
  OAI21_X1 U5857 ( .B1(n4710), .B2(n4691), .A(n4690), .ZN(U3063) );
  INV_X1 U5858 ( .A(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n4695) );
  AOI22_X1 U5859 ( .A1(n6391), .A2(n4947), .B1(n6367), .B2(n4704), .ZN(n4692)
         );
  OAI21_X1 U5860 ( .B1(n5158), .B2(n4787), .A(n4692), .ZN(n4693) );
  AOI21_X1 U5861 ( .B1(n6366), .B2(n4707), .A(n4693), .ZN(n4694) );
  OAI21_X1 U5862 ( .B1(n4710), .B2(n4695), .A(n4694), .ZN(U3062) );
  INV_X1 U5863 ( .A(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n4699) );
  AOI22_X1 U5864 ( .A1(n6391), .A2(n4958), .B1(n6376), .B2(n4704), .ZN(n4696)
         );
  OAI21_X1 U5865 ( .B1(n6446), .B2(n4787), .A(n4696), .ZN(n4697) );
  AOI21_X1 U5866 ( .B1(n6443), .B2(n4707), .A(n4697), .ZN(n4698) );
  OAI21_X1 U5867 ( .B1(n4710), .B2(n4699), .A(n4698), .ZN(U3064) );
  INV_X1 U5868 ( .A(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n4703) );
  AOI22_X1 U5869 ( .A1(n6391), .A2(n6417), .B1(n6415), .B2(n4704), .ZN(n4700)
         );
  OAI21_X1 U5870 ( .B1(n6425), .B2(n4787), .A(n4700), .ZN(n4701) );
  AOI21_X1 U5871 ( .B1(n6420), .B2(n4707), .A(n4701), .ZN(n4702) );
  OAI21_X1 U5872 ( .B1(n4710), .B2(n4703), .A(n4702), .ZN(U3066) );
  INV_X1 U5873 ( .A(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n4709) );
  AOI22_X1 U5874 ( .A1(n6391), .A2(n4952), .B1(n6390), .B2(n4704), .ZN(n4705)
         );
  OAI21_X1 U5875 ( .B1(n5153), .B2(n4787), .A(n4705), .ZN(n4706) );
  AOI21_X1 U5876 ( .B1(n6388), .B2(n4707), .A(n4706), .ZN(n4708) );
  OAI21_X1 U5877 ( .B1(n4710), .B2(n4709), .A(n4708), .ZN(U3067) );
  AOI21_X1 U5878 ( .B1(n5076), .B2(n4744), .A(n6657), .ZN(n4717) );
  AND2_X1 U5879 ( .A1(n6352), .A2(n5826), .ZN(n6358) );
  INV_X1 U5880 ( .A(n6358), .ZN(n4716) );
  NOR2_X1 U5881 ( .A1(n4718), .A2(n6497), .ZN(n6356) );
  OAI21_X1 U5882 ( .B1(n4866), .B2(n6497), .A(n4757), .ZN(n6355) );
  NOR2_X1 U5883 ( .A1(n6356), .A2(n6355), .ZN(n4715) );
  NOR2_X1 U5884 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4712), .ZN(n4746)
         );
  INV_X1 U5885 ( .A(n4746), .ZN(n4713) );
  AOI21_X1 U5886 ( .B1(STATE2_REG_3__SCAN_IN), .B2(n4713), .A(n6474), .ZN(
        n4714) );
  OAI211_X1 U5887 ( .C1(n4717), .C2(n4716), .A(n4715), .B(n4714), .ZN(n4742)
         );
  NAND2_X1 U5888 ( .A1(n4742), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n4723)
         );
  AND2_X1 U5889 ( .A1(n4799), .A2(n5826), .ZN(n5091) );
  NAND2_X1 U5890 ( .A1(n4866), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n4984) );
  INV_X1 U5891 ( .A(n4984), .ZN(n4719) );
  AND2_X1 U5892 ( .A1(n4718), .A2(STATE2_REG_2__SCAN_IN), .ZN(n5132) );
  AOI22_X1 U5893 ( .A1(n5091), .A2(n4720), .B1(n4719), .B2(n5132), .ZN(n4743)
         );
  OAI22_X1 U5894 ( .A1(n4744), .A2(n6375), .B1(n4743), .B2(n5140), .ZN(n4721)
         );
  AOI21_X1 U5895 ( .B1(n6405), .B2(n4746), .A(n4721), .ZN(n4722) );
  OAI211_X1 U5896 ( .C1(n5076), .C2(n6410), .A(n4723), .B(n4722), .ZN(U3135)
         );
  NAND2_X1 U5897 ( .A1(n4742), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n4726)
         );
  OAI22_X1 U5898 ( .A1(n4744), .A2(n6396), .B1(n4743), .B2(n5152), .ZN(n4724)
         );
  AOI21_X1 U5899 ( .B1(n6390), .B2(n4746), .A(n4724), .ZN(n4725) );
  OAI211_X1 U5900 ( .C1(n5076), .C2(n5153), .A(n4726), .B(n4725), .ZN(U3139)
         );
  NAND2_X1 U5901 ( .A1(n4742), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n4729)
         );
  INV_X1 U5902 ( .A(n6453), .ZN(n5171) );
  OAI22_X1 U5903 ( .A1(n4744), .A2(n6449), .B1(n4743), .B2(n5171), .ZN(n4727)
         );
  AOI21_X1 U5904 ( .B1(n6411), .B2(n4746), .A(n4727), .ZN(n4728) );
  OAI211_X1 U5905 ( .C1(n5076), .C2(n6458), .A(n4729), .B(n4728), .ZN(U3137)
         );
  NAND2_X1 U5906 ( .A1(n4742), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n4732)
         );
  OAI22_X1 U5907 ( .A1(n4744), .A2(n6371), .B1(n4743), .B2(n5157), .ZN(n4730)
         );
  AOI21_X1 U5908 ( .B1(n6367), .B2(n4746), .A(n4730), .ZN(n4731) );
  OAI211_X1 U5909 ( .C1(n5076), .C2(n5158), .A(n4732), .B(n4731), .ZN(U3134)
         );
  NAND2_X1 U5910 ( .A1(n4742), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n4735)
         );
  INV_X1 U5911 ( .A(n6429), .ZN(n5166) );
  OAI22_X1 U5912 ( .A1(n4744), .A2(n6427), .B1(n4743), .B2(n5166), .ZN(n4733)
         );
  AOI21_X1 U5913 ( .B1(n6397), .B2(n4746), .A(n4733), .ZN(n4734) );
  OAI211_X1 U5914 ( .C1(n5076), .C2(n6432), .A(n4735), .B(n4734), .ZN(U3132)
         );
  NAND2_X1 U5915 ( .A1(n4742), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n4738)
         );
  INV_X1 U5916 ( .A(n6443), .ZN(n5144) );
  OAI22_X1 U5917 ( .A1(n4744), .A2(n6441), .B1(n4743), .B2(n5144), .ZN(n4736)
         );
  AOI21_X1 U5918 ( .B1(n6376), .B2(n4746), .A(n4736), .ZN(n4737) );
  OAI211_X1 U5919 ( .C1(n5076), .C2(n6446), .A(n4738), .B(n4737), .ZN(U3136)
         );
  NAND2_X1 U5920 ( .A1(n4742), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n4741)
         );
  OAI22_X1 U5921 ( .A1(n4744), .A2(n6386), .B1(n4743), .B2(n5148), .ZN(n4739)
         );
  AOI21_X1 U5922 ( .B1(n6415), .B2(n4746), .A(n4739), .ZN(n4740) );
  OAI211_X1 U5923 ( .C1(n5076), .C2(n6425), .A(n4741), .B(n4740), .ZN(U3138)
         );
  NAND2_X1 U5924 ( .A1(n4742), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n4748)
         );
  INV_X1 U5925 ( .A(n6436), .ZN(n5162) );
  OAI22_X1 U5926 ( .A1(n4744), .A2(n6434), .B1(n4743), .B2(n5162), .ZN(n4745)
         );
  AOI21_X1 U5927 ( .B1(n6401), .B2(n4746), .A(n4745), .ZN(n4747) );
  OAI211_X1 U5928 ( .C1(n5076), .C2(n6439), .A(n4748), .B(n4747), .ZN(U3133)
         );
  NOR3_X4 U5929 ( .A1(n4750), .A2(n4915), .A3(n4749), .ZN(n4959) );
  INV_X1 U5930 ( .A(n4959), .ZN(n4754) );
  INV_X1 U5931 ( .A(n4751), .ZN(n4752) );
  OAI211_X1 U5932 ( .C1(n4754), .C2(n5128), .A(n4753), .B(n4752), .ZN(n4759)
         );
  OR2_X1 U5933 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4755), .ZN(n4783)
         );
  INV_X1 U5934 ( .A(n4865), .ZN(n4756) );
  NOR2_X1 U5935 ( .A1(n4756), .A2(n4866), .ZN(n5138) );
  OAI21_X1 U5936 ( .B1(n5138), .B2(n6497), .A(n4757), .ZN(n5131) );
  AOI211_X1 U5937 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n4783), .A(n6356), .B(
        n5131), .ZN(n4758) );
  NAND2_X1 U5938 ( .A1(n4759), .A2(n4758), .ZN(n4781) );
  NAND2_X1 U5939 ( .A1(n4781), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n4762) );
  INV_X1 U5940 ( .A(n6401), .ZN(n6433) );
  AOI22_X1 U5941 ( .A1(n6348), .A2(n5033), .B1(n5132), .B2(n5138), .ZN(n4782)
         );
  OAI22_X1 U5942 ( .A1(n6433), .A2(n4783), .B1(n4782), .B2(n5162), .ZN(n4760)
         );
  AOI21_X1 U5943 ( .B1(n4959), .B2(n6363), .A(n4760), .ZN(n4761) );
  OAI211_X1 U5944 ( .C1(n4787), .C2(n6434), .A(n4762), .B(n4761), .ZN(U3053)
         );
  NAND2_X1 U5945 ( .A1(n4781), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n4765) );
  OAI22_X1 U5946 ( .A1(n5055), .A2(n4783), .B1(n4782), .B2(n5140), .ZN(n4763)
         );
  AOI21_X1 U5947 ( .B1(n4959), .B2(n6372), .A(n4763), .ZN(n4764) );
  OAI211_X1 U5948 ( .C1(n4787), .C2(n6375), .A(n4765), .B(n4764), .ZN(U3055)
         );
  NAND2_X1 U5949 ( .A1(n4781), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n4768) );
  INV_X1 U5950 ( .A(n6397), .ZN(n6426) );
  OAI22_X1 U5951 ( .A1(n6426), .A2(n4783), .B1(n4782), .B2(n5166), .ZN(n4766)
         );
  AOI21_X1 U5952 ( .B1(n4959), .B2(n6360), .A(n4766), .ZN(n4767) );
  OAI211_X1 U5953 ( .C1(n4787), .C2(n6427), .A(n4768), .B(n4767), .ZN(U3052)
         );
  NAND2_X1 U5954 ( .A1(n4781), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n4771) );
  INV_X1 U5955 ( .A(n6411), .ZN(n6448) );
  OAI22_X1 U5956 ( .A1(n6448), .A2(n4783), .B1(n4782), .B2(n5171), .ZN(n4769)
         );
  AOI21_X1 U5957 ( .B1(n4959), .B2(n6380), .A(n4769), .ZN(n4770) );
  OAI211_X1 U5958 ( .C1(n4787), .C2(n6449), .A(n4771), .B(n4770), .ZN(U3057)
         );
  NAND2_X1 U5959 ( .A1(n4781), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n4774) );
  OAI22_X1 U5960 ( .A1(n5065), .A2(n4783), .B1(n4782), .B2(n5148), .ZN(n4772)
         );
  AOI21_X1 U5961 ( .B1(n4959), .B2(n6383), .A(n4772), .ZN(n4773) );
  OAI211_X1 U5962 ( .C1(n4787), .C2(n6386), .A(n4774), .B(n4773), .ZN(U3058)
         );
  NAND2_X1 U5963 ( .A1(n4781), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n4777) );
  OAI22_X1 U5964 ( .A1(n5051), .A2(n4783), .B1(n4782), .B2(n5157), .ZN(n4775)
         );
  AOI21_X1 U5965 ( .B1(n4959), .B2(n6368), .A(n4775), .ZN(n4776) );
  OAI211_X1 U5966 ( .C1(n4787), .C2(n6371), .A(n4777), .B(n4776), .ZN(U3054)
         );
  NAND2_X1 U5967 ( .A1(n4781), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n4780) );
  OAI22_X1 U5968 ( .A1(n5072), .A2(n4783), .B1(n4782), .B2(n5152), .ZN(n4778)
         );
  AOI21_X1 U5969 ( .B1(n4959), .B2(n6392), .A(n4778), .ZN(n4779) );
  OAI211_X1 U5970 ( .C1(n4787), .C2(n6396), .A(n4780), .B(n4779), .ZN(U3059)
         );
  NAND2_X1 U5971 ( .A1(n4781), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n4786) );
  INV_X1 U5972 ( .A(n6376), .ZN(n6440) );
  OAI22_X1 U5973 ( .A1(n6440), .A2(n4783), .B1(n4782), .B2(n5144), .ZN(n4784)
         );
  AOI21_X1 U5974 ( .B1(n4959), .B2(n6377), .A(n4784), .ZN(n4785) );
  OAI211_X1 U5975 ( .C1(n4787), .C2(n6441), .A(n4786), .B(n4785), .ZN(U3056)
         );
  NAND2_X1 U5976 ( .A1(n4790), .A2(n4789), .ZN(n4791) );
  AND2_X1 U5977 ( .A1(n4850), .A2(n4791), .ZN(n6225) );
  INV_X1 U5978 ( .A(n6225), .ZN(n4794) );
  INV_X1 U5979 ( .A(EBX_REG_6__SCAN_IN), .ZN(n4793) );
  OAI21_X1 U5980 ( .B1(n4792), .B2(n3003), .A(n4852), .ZN(n6301) );
  OAI222_X1 U5981 ( .A1(n4794), .A2(n5576), .B1(n4793), .B2(n6095), .C1(n5555), 
        .C2(n6301), .ZN(U2853) );
  OAI222_X1 U5982 ( .A1(n4794), .A2(n5878), .B1(n5305), .B2(n6715), .C1(n6181), 
        .C2(n5397), .ZN(U2885) );
  NAND3_X1 U5983 ( .A1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n6474), .A3(n6468), .ZN(n4924) );
  NOR2_X1 U5984 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4924), .ZN(n4835)
         );
  AND2_X1 U5985 ( .A1(n5831), .A2(n4795), .ZN(n4796) );
  INV_X1 U5986 ( .A(n4961), .ZN(n4797) );
  NOR2_X1 U5987 ( .A1(n4838), .A2(n4797), .ZN(n4801) );
  NOR2_X1 U5988 ( .A1(n4799), .A2(n4798), .ZN(n4919) );
  INV_X1 U5989 ( .A(n4919), .ZN(n4800) );
  OAI21_X1 U5990 ( .B1(n4801), .B2(n5128), .A(n4800), .ZN(n4802) );
  NOR2_X1 U5991 ( .A1(n5132), .A2(n6355), .ZN(n4982) );
  OAI221_X1 U5992 ( .B1(n4835), .B2(n6581), .C1(n4835), .C2(n4802), .A(n4982), 
        .ZN(n4803) );
  INV_X1 U5993 ( .A(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n4809) );
  NAND2_X1 U5994 ( .A1(n4919), .A2(n5826), .ZN(n4805) );
  AND2_X1 U5995 ( .A1(n4866), .A2(n6474), .ZN(n6349) );
  NAND2_X1 U5996 ( .A1(n6356), .A2(n6349), .ZN(n4804) );
  NAND2_X1 U5997 ( .A1(n4805), .A2(n4804), .ZN(n4834) );
  AOI22_X1 U5998 ( .A1(n6401), .A2(n4835), .B1(n6436), .B2(n4834), .ZN(n4806)
         );
  OAI21_X1 U5999 ( .B1(n6434), .B2(n4961), .A(n4806), .ZN(n4807) );
  AOI21_X1 U6000 ( .B1(n6363), .B2(n4838), .A(n4807), .ZN(n4808) );
  OAI21_X1 U6001 ( .B1(n4841), .B2(n4809), .A(n4808), .ZN(U3037) );
  INV_X1 U6002 ( .A(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n4813) );
  AOI22_X1 U6003 ( .A1(n6415), .A2(n4835), .B1(n6420), .B2(n4834), .ZN(n4810)
         );
  OAI21_X1 U6004 ( .B1(n6386), .B2(n4961), .A(n4810), .ZN(n4811) );
  AOI21_X1 U6005 ( .B1(n6383), .B2(n4838), .A(n4811), .ZN(n4812) );
  OAI21_X1 U6006 ( .B1(n4841), .B2(n4813), .A(n4812), .ZN(U3042) );
  INV_X1 U6007 ( .A(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n4817) );
  AOI22_X1 U6008 ( .A1(n6376), .A2(n4835), .B1(n6443), .B2(n4834), .ZN(n4814)
         );
  OAI21_X1 U6009 ( .B1(n6441), .B2(n4961), .A(n4814), .ZN(n4815) );
  AOI21_X1 U6010 ( .B1(n6377), .B2(n4838), .A(n4815), .ZN(n4816) );
  OAI21_X1 U6011 ( .B1(n4841), .B2(n4817), .A(n4816), .ZN(U3040) );
  INV_X1 U6012 ( .A(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n4821) );
  AOI22_X1 U6013 ( .A1(n6405), .A2(n4835), .B1(n6407), .B2(n4834), .ZN(n4818)
         );
  OAI21_X1 U6014 ( .B1(n6375), .B2(n4961), .A(n4818), .ZN(n4819) );
  AOI21_X1 U6015 ( .B1(n6372), .B2(n4838), .A(n4819), .ZN(n4820) );
  OAI21_X1 U6016 ( .B1(n4841), .B2(n4821), .A(n4820), .ZN(U3039) );
  INV_X1 U6017 ( .A(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n4825) );
  AOI22_X1 U6018 ( .A1(n6397), .A2(n4835), .B1(n6429), .B2(n4834), .ZN(n4822)
         );
  OAI21_X1 U6019 ( .B1(n6427), .B2(n4961), .A(n4822), .ZN(n4823) );
  AOI21_X1 U6020 ( .B1(n6360), .B2(n4838), .A(n4823), .ZN(n4824) );
  OAI21_X1 U6021 ( .B1(n4841), .B2(n4825), .A(n4824), .ZN(U3036) );
  INV_X1 U6022 ( .A(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n4829) );
  AOI22_X1 U6023 ( .A1(n6390), .A2(n4835), .B1(n6388), .B2(n4834), .ZN(n4826)
         );
  OAI21_X1 U6024 ( .B1(n6396), .B2(n4961), .A(n4826), .ZN(n4827) );
  AOI21_X1 U6025 ( .B1(n6392), .B2(n4838), .A(n4827), .ZN(n4828) );
  OAI21_X1 U6026 ( .B1(n4841), .B2(n4829), .A(n4828), .ZN(U3043) );
  INV_X1 U6027 ( .A(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n4833) );
  AOI22_X1 U6028 ( .A1(n6367), .A2(n4835), .B1(n6366), .B2(n4834), .ZN(n4830)
         );
  OAI21_X1 U6029 ( .B1(n6371), .B2(n4961), .A(n4830), .ZN(n4831) );
  AOI21_X1 U6030 ( .B1(n6368), .B2(n4838), .A(n4831), .ZN(n4832) );
  OAI21_X1 U6031 ( .B1(n4841), .B2(n4833), .A(n4832), .ZN(U3038) );
  INV_X1 U6032 ( .A(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n4840) );
  AOI22_X1 U6033 ( .A1(n6411), .A2(n4835), .B1(n6453), .B2(n4834), .ZN(n4836)
         );
  OAI21_X1 U6034 ( .B1(n6449), .B2(n4961), .A(n4836), .ZN(n4837) );
  AOI21_X1 U6035 ( .B1(n6380), .B2(n4838), .A(n4837), .ZN(n4839) );
  OAI21_X1 U6036 ( .B1(n4841), .B2(n4840), .A(n4839), .ZN(U3041) );
  OAI21_X1 U6037 ( .B1(n4844), .B2(n4843), .A(n4842), .ZN(n6306) );
  INV_X1 U6038 ( .A(REIP_REG_5__SCAN_IN), .ZN(n4845) );
  OAI22_X1 U6039 ( .A1(n5691), .A2(n4846), .B1(n6335), .B2(n4845), .ZN(n4848)
         );
  NOR2_X1 U6040 ( .A1(n5211), .A2(n5697), .ZN(n4847) );
  AOI211_X1 U6041 ( .C1(n6217), .C2(n5209), .A(n4848), .B(n4847), .ZN(n4849)
         );
  OAI21_X1 U6042 ( .B1(n6221), .B2(n6306), .A(n4849), .ZN(U2981) );
  XOR2_X1 U6043 ( .A(n4851), .B(n4850), .Z(n5087) );
  INV_X1 U6044 ( .A(n5087), .ZN(n4909) );
  AOI21_X1 U6045 ( .B1(n4853), .B2(n4852), .A(n5026), .ZN(n6288) );
  AOI22_X1 U6046 ( .A1(n6288), .A2(n6092), .B1(EBX_REG_7__SCAN_IN), .B2(n4150), 
        .ZN(n4854) );
  OAI21_X1 U6047 ( .B1(n4909), .B2(n5576), .A(n4854), .ZN(U2852) );
  OAI21_X1 U6048 ( .B1(n4857), .B2(n4856), .A(n4855), .ZN(n6289) );
  NOR2_X1 U6049 ( .A1(n6335), .A2(n4253), .ZN(n6287) );
  AOI21_X1 U6050 ( .B1(n6239), .B2(PHYADDRPOINTER_REG_7__SCAN_IN), .A(n6287), 
        .ZN(n4858) );
  OAI21_X1 U6051 ( .B1(n5084), .B2(n6249), .A(n4858), .ZN(n4859) );
  AOI21_X1 U6052 ( .B1(n5087), .B2(n6244), .A(n4859), .ZN(n4860) );
  OAI21_X1 U6053 ( .B1(n6289), .B2(n6221), .A(n4860), .ZN(U2979) );
  NAND2_X1 U6054 ( .A1(n4862), .A2(n4861), .ZN(n4870) );
  AOI21_X1 U6055 ( .B1(n6450), .B2(n4870), .A(n6657), .ZN(n4863) );
  AOI211_X1 U6056 ( .C1(n5033), .C2(n4864), .A(n5835), .B(n4863), .ZN(n4869)
         );
  NOR3_X1 U6057 ( .A1(n6468), .A2(n6474), .A3(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), 
        .ZN(n5037) );
  INV_X1 U6058 ( .A(n5037), .ZN(n5030) );
  NOR2_X1 U6059 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5030), .ZN(n4903)
         );
  INV_X1 U6060 ( .A(n6356), .ZN(n4985) );
  OR2_X1 U6061 ( .A1(n4866), .A2(n4865), .ZN(n4871) );
  AOI21_X1 U6062 ( .B1(n4871), .B2(STATE2_REG_2__SCAN_IN), .A(n4867), .ZN(
        n5093) );
  OAI211_X1 U6063 ( .C1(n6581), .C2(n4903), .A(n4985), .B(n5093), .ZN(n4868)
         );
  INV_X1 U6064 ( .A(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n4877) );
  NAND2_X1 U6065 ( .A1(n5091), .A2(n5033), .ZN(n4873) );
  INV_X1 U6066 ( .A(n4871), .ZN(n5090) );
  NAND2_X1 U6067 ( .A1(n5090), .A2(n5132), .ZN(n4872) );
  NAND2_X1 U6068 ( .A1(n4873), .A2(n4872), .ZN(n4902) );
  AOI22_X1 U6069 ( .A1(n6401), .A2(n4903), .B1(n6436), .B2(n4902), .ZN(n4874)
         );
  OAI21_X1 U6070 ( .B1(n6450), .B2(n6439), .A(n4874), .ZN(n4875) );
  AOI21_X1 U6071 ( .B1(n6402), .B2(n5074), .A(n4875), .ZN(n4876) );
  OAI21_X1 U6072 ( .B1(n4908), .B2(n4877), .A(n4876), .ZN(U3117) );
  INV_X1 U6073 ( .A(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n4881) );
  AOI22_X1 U6074 ( .A1(n6397), .A2(n4903), .B1(n6429), .B2(n4902), .ZN(n4878)
         );
  OAI21_X1 U6075 ( .B1(n6450), .B2(n6432), .A(n4878), .ZN(n4879) );
  AOI21_X1 U6076 ( .B1(n6398), .B2(n5074), .A(n4879), .ZN(n4880) );
  OAI21_X1 U6077 ( .B1(n4908), .B2(n4881), .A(n4880), .ZN(U3116) );
  INV_X1 U6078 ( .A(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n4885) );
  AOI22_X1 U6079 ( .A1(n6411), .A2(n4903), .B1(n6453), .B2(n4902), .ZN(n4882)
         );
  OAI21_X1 U6080 ( .B1(n6450), .B2(n6458), .A(n4882), .ZN(n4883) );
  AOI21_X1 U6081 ( .B1(n6412), .B2(n5074), .A(n4883), .ZN(n4884) );
  OAI21_X1 U6082 ( .B1(n4908), .B2(n4885), .A(n4884), .ZN(U3121) );
  INV_X1 U6083 ( .A(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n4889) );
  AOI22_X1 U6084 ( .A1(n6367), .A2(n4903), .B1(n6366), .B2(n4902), .ZN(n4886)
         );
  OAI21_X1 U6085 ( .B1(n6450), .B2(n5158), .A(n4886), .ZN(n4887) );
  AOI21_X1 U6086 ( .B1(n4947), .B2(n5074), .A(n4887), .ZN(n4888) );
  OAI21_X1 U6087 ( .B1(n4908), .B2(n4889), .A(n4888), .ZN(U3118) );
  INV_X1 U6088 ( .A(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n4893) );
  AOI22_X1 U6089 ( .A1(n6405), .A2(n4903), .B1(n6407), .B2(n4902), .ZN(n4890)
         );
  OAI21_X1 U6090 ( .B1(n6450), .B2(n6410), .A(n4890), .ZN(n4891) );
  AOI21_X1 U6091 ( .B1(n6406), .B2(n5074), .A(n4891), .ZN(n4892) );
  OAI21_X1 U6092 ( .B1(n4908), .B2(n4893), .A(n4892), .ZN(U3119) );
  INV_X1 U6093 ( .A(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n4897) );
  AOI22_X1 U6094 ( .A1(n6415), .A2(n4903), .B1(n6420), .B2(n4902), .ZN(n4894)
         );
  OAI21_X1 U6095 ( .B1(n6450), .B2(n6425), .A(n4894), .ZN(n4895) );
  AOI21_X1 U6096 ( .B1(n6417), .B2(n5074), .A(n4895), .ZN(n4896) );
  OAI21_X1 U6097 ( .B1(n4908), .B2(n4897), .A(n4896), .ZN(U3122) );
  INV_X1 U6098 ( .A(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n4901) );
  AOI22_X1 U6099 ( .A1(n6390), .A2(n4903), .B1(n6388), .B2(n4902), .ZN(n4898)
         );
  OAI21_X1 U6100 ( .B1(n6450), .B2(n5153), .A(n4898), .ZN(n4899) );
  AOI21_X1 U6101 ( .B1(n4952), .B2(n5074), .A(n4899), .ZN(n4900) );
  OAI21_X1 U6102 ( .B1(n4908), .B2(n4901), .A(n4900), .ZN(U3123) );
  INV_X1 U6103 ( .A(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n4907) );
  AOI22_X1 U6104 ( .A1(n6376), .A2(n4903), .B1(n6443), .B2(n4902), .ZN(n4904)
         );
  OAI21_X1 U6105 ( .B1(n6450), .B2(n6446), .A(n4904), .ZN(n4905) );
  AOI21_X1 U6106 ( .B1(n4958), .B2(n5074), .A(n4905), .ZN(n4906) );
  OAI21_X1 U6107 ( .B1(n4908), .B2(n4907), .A(n4906), .ZN(U3120) );
  INV_X1 U6108 ( .A(EAX_REG_7__SCAN_IN), .ZN(n6184) );
  OAI222_X1 U6109 ( .A1(n5878), .A2(n4909), .B1(n5397), .B2(n6184), .C1(n6713), 
        .C2(n5305), .ZN(U2884) );
  NAND2_X1 U6110 ( .A1(n4911), .A2(n4912), .ZN(n5213) );
  OAI21_X1 U6111 ( .B1(n4911), .B2(n4912), .A(n5213), .ZN(n5024) );
  INV_X1 U6112 ( .A(DATAI_8_), .ZN(n4913) );
  INV_X1 U6113 ( .A(EAX_REG_8__SCAN_IN), .ZN(n6187) );
  OAI222_X1 U6114 ( .A1(n5024), .A2(n5878), .B1(n5305), .B2(n4913), .C1(n5397), 
        .C2(n6187), .ZN(U2883) );
  INV_X1 U6115 ( .A(n4914), .ZN(n5832) );
  NOR3_X1 U6116 ( .A1(n4916), .A2(n4915), .A3(n5832), .ZN(n4917) );
  NOR2_X1 U6117 ( .A1(n4917), .A2(n5835), .ZN(n4923) );
  NOR2_X1 U6118 ( .A1(n4918), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n4957)
         );
  AOI21_X1 U6119 ( .B1(n4919), .B2(n5412), .A(n4957), .ZN(n4925) );
  INV_X1 U6120 ( .A(n4924), .ZN(n4920) );
  NOR2_X1 U6121 ( .A1(n5826), .A2(n4920), .ZN(n4922) );
  AOI211_X2 U6122 ( .C1(n4923), .C2(n4925), .A(n4922), .B(n4921), .ZN(n4966)
         );
  INV_X1 U6123 ( .A(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n4930) );
  INV_X1 U6124 ( .A(n4923), .ZN(n4926) );
  OAI22_X1 U6125 ( .A1(n4926), .A2(n4925), .B1(n4924), .B2(n6497), .ZN(n4963)
         );
  AOI22_X1 U6126 ( .A1(n4959), .A2(n6398), .B1(n6397), .B2(n4957), .ZN(n4927)
         );
  OAI21_X1 U6127 ( .B1(n6432), .B2(n4961), .A(n4927), .ZN(n4928) );
  AOI21_X1 U6128 ( .B1(n4963), .B2(n6429), .A(n4928), .ZN(n4929) );
  OAI21_X1 U6129 ( .B1(n4966), .B2(n4930), .A(n4929), .ZN(U3044) );
  INV_X1 U6130 ( .A(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n4934) );
  AOI22_X1 U6131 ( .A1(n4959), .A2(n6406), .B1(n6405), .B2(n4957), .ZN(n4931)
         );
  OAI21_X1 U6132 ( .B1(n6410), .B2(n4961), .A(n4931), .ZN(n4932) );
  AOI21_X1 U6133 ( .B1(n4963), .B2(n6407), .A(n4932), .ZN(n4933) );
  OAI21_X1 U6134 ( .B1(n4966), .B2(n4934), .A(n4933), .ZN(U3047) );
  INV_X1 U6135 ( .A(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n4938) );
  AOI22_X1 U6136 ( .A1(n4959), .A2(n6402), .B1(n6401), .B2(n4957), .ZN(n4935)
         );
  OAI21_X1 U6137 ( .B1(n6439), .B2(n4961), .A(n4935), .ZN(n4936) );
  AOI21_X1 U6138 ( .B1(n4963), .B2(n6436), .A(n4936), .ZN(n4937) );
  OAI21_X1 U6139 ( .B1(n4966), .B2(n4938), .A(n4937), .ZN(U3045) );
  INV_X1 U6140 ( .A(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n4942) );
  AOI22_X1 U6141 ( .A1(n4959), .A2(n6412), .B1(n6411), .B2(n4957), .ZN(n4939)
         );
  OAI21_X1 U6142 ( .B1(n6458), .B2(n4961), .A(n4939), .ZN(n4940) );
  AOI21_X1 U6143 ( .B1(n4963), .B2(n6453), .A(n4940), .ZN(n4941) );
  OAI21_X1 U6144 ( .B1(n4966), .B2(n4942), .A(n4941), .ZN(U3049) );
  INV_X1 U6145 ( .A(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n4946) );
  AOI22_X1 U6146 ( .A1(n4959), .A2(n6417), .B1(n6415), .B2(n4957), .ZN(n4943)
         );
  OAI21_X1 U6147 ( .B1(n6425), .B2(n4961), .A(n4943), .ZN(n4944) );
  AOI21_X1 U6148 ( .B1(n4963), .B2(n6420), .A(n4944), .ZN(n4945) );
  OAI21_X1 U6149 ( .B1(n4966), .B2(n4946), .A(n4945), .ZN(U3050) );
  INV_X1 U6150 ( .A(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n4951) );
  AOI22_X1 U6151 ( .A1(n4959), .A2(n4947), .B1(n6367), .B2(n4957), .ZN(n4948)
         );
  OAI21_X1 U6152 ( .B1(n5158), .B2(n4961), .A(n4948), .ZN(n4949) );
  AOI21_X1 U6153 ( .B1(n4963), .B2(n6366), .A(n4949), .ZN(n4950) );
  OAI21_X1 U6154 ( .B1(n4966), .B2(n4951), .A(n4950), .ZN(U3046) );
  INV_X1 U6155 ( .A(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n4956) );
  AOI22_X1 U6156 ( .A1(n4959), .A2(n4952), .B1(n6390), .B2(n4957), .ZN(n4953)
         );
  OAI21_X1 U6157 ( .B1(n5153), .B2(n4961), .A(n4953), .ZN(n4954) );
  AOI21_X1 U6158 ( .B1(n4963), .B2(n6388), .A(n4954), .ZN(n4955) );
  OAI21_X1 U6159 ( .B1(n4966), .B2(n4956), .A(n4955), .ZN(U3051) );
  INV_X1 U6160 ( .A(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n4965) );
  AOI22_X1 U6161 ( .A1(n4959), .A2(n4958), .B1(n6376), .B2(n4957), .ZN(n4960)
         );
  OAI21_X1 U6162 ( .B1(n6446), .B2(n4961), .A(n4960), .ZN(n4962) );
  AOI21_X1 U6163 ( .B1(n4963), .B2(n6443), .A(n4962), .ZN(n4964) );
  OAI21_X1 U6164 ( .B1(n4966), .B2(n4965), .A(n4964), .ZN(U3048) );
  OAI21_X1 U6165 ( .B1(n4969), .B2(n4968), .A(n4967), .ZN(n4970) );
  INV_X1 U6166 ( .A(n4970), .ZN(n6281) );
  NAND2_X1 U6167 ( .A1(n6281), .A2(n6243), .ZN(n4975) );
  INV_X1 U6168 ( .A(REIP_REG_8__SCAN_IN), .ZN(n4971) );
  NOR2_X1 U6169 ( .A1(n6335), .A2(n4971), .ZN(n6279) );
  NOR2_X1 U6170 ( .A1(n5691), .A2(n4972), .ZN(n4973) );
  AOI211_X1 U6171 ( .C1(n6217), .C2(n6027), .A(n6279), .B(n4973), .ZN(n4974)
         );
  OAI211_X1 U6172 ( .C1(n5697), .C2(n5024), .A(n4975), .B(n4974), .ZN(U2978)
         );
  INV_X1 U6173 ( .A(n6457), .ZN(n4976) );
  OAI21_X1 U6174 ( .B1(n4976), .B2(n5017), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n4977) );
  NAND2_X1 U6175 ( .A1(n4977), .A2(n5826), .ZN(n4987) );
  INV_X1 U6176 ( .A(n4987), .ZN(n4980) );
  NOR2_X1 U6177 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4978), .ZN(n5016)
         );
  INV_X1 U6178 ( .A(n5016), .ZN(n4979) );
  AOI22_X1 U6179 ( .A1(n4980), .A2(n4986), .B1(STATE2_REG_3__SCAN_IN), .B2(
        n4979), .ZN(n4981) );
  OAI211_X1 U6180 ( .C1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .C2(n6497), .A(n4982), .B(n4981), .ZN(n4983) );
  INV_X1 U6181 ( .A(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n4991) );
  OAI22_X1 U6182 ( .A1(n4987), .A2(n4986), .B1(n4985), .B2(n4984), .ZN(n5020)
         );
  AOI22_X1 U6183 ( .A1(n5017), .A2(n6360), .B1(n6397), .B2(n5016), .ZN(n4988)
         );
  OAI21_X1 U6184 ( .B1(n6457), .B2(n6427), .A(n4988), .ZN(n4989) );
  AOI21_X1 U6185 ( .B1(n5020), .B2(n6429), .A(n4989), .ZN(n4990) );
  OAI21_X1 U6186 ( .B1(n5023), .B2(n4991), .A(n4990), .ZN(U3100) );
  INV_X1 U6187 ( .A(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n4995) );
  AOI22_X1 U6188 ( .A1(n5017), .A2(n6372), .B1(n5016), .B2(n6405), .ZN(n4992)
         );
  OAI21_X1 U6189 ( .B1(n6457), .B2(n6375), .A(n4992), .ZN(n4993) );
  AOI21_X1 U6190 ( .B1(n5020), .B2(n6407), .A(n4993), .ZN(n4994) );
  OAI21_X1 U6191 ( .B1(n5023), .B2(n4995), .A(n4994), .ZN(U3103) );
  INV_X1 U6192 ( .A(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n4999) );
  AOI22_X1 U6193 ( .A1(n5017), .A2(n6392), .B1(n5016), .B2(n6390), .ZN(n4996)
         );
  OAI21_X1 U6194 ( .B1(n6457), .B2(n6396), .A(n4996), .ZN(n4997) );
  AOI21_X1 U6195 ( .B1(n5020), .B2(n6388), .A(n4997), .ZN(n4998) );
  OAI21_X1 U6196 ( .B1(n5023), .B2(n4999), .A(n4998), .ZN(U3107) );
  INV_X1 U6197 ( .A(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n5003) );
  AOI22_X1 U6198 ( .A1(n5017), .A2(n6383), .B1(n5016), .B2(n6415), .ZN(n5000)
         );
  OAI21_X1 U6199 ( .B1(n6457), .B2(n6386), .A(n5000), .ZN(n5001) );
  AOI21_X1 U6200 ( .B1(n5020), .B2(n6420), .A(n5001), .ZN(n5002) );
  OAI21_X1 U6201 ( .B1(n5023), .B2(n5003), .A(n5002), .ZN(U3106) );
  INV_X1 U6202 ( .A(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n5007) );
  AOI22_X1 U6203 ( .A1(n5017), .A2(n6368), .B1(n5016), .B2(n6367), .ZN(n5004)
         );
  OAI21_X1 U6204 ( .B1(n6457), .B2(n6371), .A(n5004), .ZN(n5005) );
  AOI21_X1 U6205 ( .B1(n5020), .B2(n6366), .A(n5005), .ZN(n5006) );
  OAI21_X1 U6206 ( .B1(n5023), .B2(n5007), .A(n5006), .ZN(U3102) );
  INV_X1 U6207 ( .A(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n5011) );
  AOI22_X1 U6208 ( .A1(n5017), .A2(n6363), .B1(n5016), .B2(n6401), .ZN(n5008)
         );
  OAI21_X1 U6209 ( .B1(n6457), .B2(n6434), .A(n5008), .ZN(n5009) );
  AOI21_X1 U6210 ( .B1(n5020), .B2(n6436), .A(n5009), .ZN(n5010) );
  OAI21_X1 U6211 ( .B1(n5023), .B2(n5011), .A(n5010), .ZN(U3101) );
  INV_X1 U6212 ( .A(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n5015) );
  AOI22_X1 U6213 ( .A1(n5017), .A2(n6377), .B1(n5016), .B2(n6376), .ZN(n5012)
         );
  OAI21_X1 U6214 ( .B1(n6457), .B2(n6441), .A(n5012), .ZN(n5013) );
  AOI21_X1 U6215 ( .B1(n5020), .B2(n6443), .A(n5013), .ZN(n5014) );
  OAI21_X1 U6216 ( .B1(n5023), .B2(n5015), .A(n5014), .ZN(U3104) );
  INV_X1 U6217 ( .A(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n5022) );
  AOI22_X1 U6218 ( .A1(n5017), .A2(n6380), .B1(n5016), .B2(n6411), .ZN(n5018)
         );
  OAI21_X1 U6219 ( .B1(n6457), .B2(n6449), .A(n5018), .ZN(n5019) );
  AOI21_X1 U6220 ( .B1(n5020), .B2(n6453), .A(n5019), .ZN(n5021) );
  OAI21_X1 U6221 ( .B1(n5023), .B2(n5022), .A(n5021), .ZN(U3105) );
  INV_X1 U6222 ( .A(n5024), .ZN(n6020) );
  NOR2_X1 U6223 ( .A1(n5026), .A2(n5025), .ZN(n5027) );
  OR2_X1 U6224 ( .A1(n5181), .A2(n5027), .ZN(n6018) );
  OAI22_X1 U6225 ( .A1(n6018), .A2(n5555), .B1(n6031), .B2(n6095), .ZN(n5028)
         );
  AOI21_X1 U6226 ( .B1(n6020), .B2(n4149), .A(n5028), .ZN(n5029) );
  INV_X1 U6227 ( .A(n5029), .ZN(U2851) );
  NOR2_X1 U6228 ( .A1(n5031), .A2(n5030), .ZN(n5032) );
  INV_X1 U6229 ( .A(n5032), .ZN(n5071) );
  AOI21_X1 U6230 ( .B1(n5034), .B2(n5033), .A(n5032), .ZN(n5039) );
  OR2_X1 U6231 ( .A1(n5039), .A2(n5835), .ZN(n5036) );
  NAND2_X1 U6232 ( .A1(STATE2_REG_2__SCAN_IN), .A2(n5037), .ZN(n5035) );
  NAND2_X1 U6233 ( .A1(n5036), .A2(n5035), .ZN(n5069) );
  OR2_X1 U6234 ( .A1(n5826), .A2(n5037), .ZN(n5043) );
  AND2_X1 U6235 ( .A1(n5039), .A2(n5038), .ZN(n5040) );
  NAND2_X1 U6236 ( .A1(n5826), .A2(n5040), .ZN(n5042) );
  NAND3_X1 U6237 ( .A1(n5043), .A2(n5042), .A3(n5041), .ZN(n5068) );
  AOI22_X1 U6238 ( .A1(n5069), .A2(n6429), .B1(INSTQUEUE_REG_13__0__SCAN_IN), 
        .B2(n5068), .ZN(n5044) );
  OAI21_X1 U6239 ( .B1(n6426), .B2(n5071), .A(n5044), .ZN(n5045) );
  AOI21_X1 U6240 ( .B1(n5074), .B2(n6360), .A(n5045), .ZN(n5046) );
  OAI21_X1 U6241 ( .B1(n6427), .B2(n5076), .A(n5046), .ZN(U3124) );
  AOI22_X1 U6242 ( .A1(n5069), .A2(n6436), .B1(INSTQUEUE_REG_13__1__SCAN_IN), 
        .B2(n5068), .ZN(n5047) );
  OAI21_X1 U6243 ( .B1(n6433), .B2(n5071), .A(n5047), .ZN(n5048) );
  AOI21_X1 U6244 ( .B1(n5074), .B2(n6363), .A(n5048), .ZN(n5049) );
  OAI21_X1 U6245 ( .B1(n6434), .B2(n5076), .A(n5049), .ZN(U3125) );
  AOI22_X1 U6246 ( .A1(n5069), .A2(n6366), .B1(INSTQUEUE_REG_13__2__SCAN_IN), 
        .B2(n5068), .ZN(n5050) );
  OAI21_X1 U6247 ( .B1(n5051), .B2(n5071), .A(n5050), .ZN(n5052) );
  AOI21_X1 U6248 ( .B1(n5074), .B2(n6368), .A(n5052), .ZN(n5053) );
  OAI21_X1 U6249 ( .B1(n6371), .B2(n5076), .A(n5053), .ZN(U3126) );
  AOI22_X1 U6250 ( .A1(n5069), .A2(n6407), .B1(INSTQUEUE_REG_13__3__SCAN_IN), 
        .B2(n5068), .ZN(n5054) );
  OAI21_X1 U6251 ( .B1(n5055), .B2(n5071), .A(n5054), .ZN(n5056) );
  AOI21_X1 U6252 ( .B1(n5074), .B2(n6372), .A(n5056), .ZN(n5057) );
  OAI21_X1 U6253 ( .B1(n6375), .B2(n5076), .A(n5057), .ZN(U3127) );
  AOI22_X1 U6254 ( .A1(n5069), .A2(n6443), .B1(INSTQUEUE_REG_13__4__SCAN_IN), 
        .B2(n5068), .ZN(n5058) );
  OAI21_X1 U6255 ( .B1(n6440), .B2(n5071), .A(n5058), .ZN(n5059) );
  AOI21_X1 U6256 ( .B1(n5074), .B2(n6377), .A(n5059), .ZN(n5060) );
  OAI21_X1 U6257 ( .B1(n6441), .B2(n5076), .A(n5060), .ZN(U3128) );
  AOI22_X1 U6258 ( .A1(n5069), .A2(n6453), .B1(INSTQUEUE_REG_13__5__SCAN_IN), 
        .B2(n5068), .ZN(n5061) );
  OAI21_X1 U6259 ( .B1(n6448), .B2(n5071), .A(n5061), .ZN(n5062) );
  AOI21_X1 U6260 ( .B1(n5074), .B2(n6380), .A(n5062), .ZN(n5063) );
  OAI21_X1 U6261 ( .B1(n6449), .B2(n5076), .A(n5063), .ZN(U3129) );
  AOI22_X1 U6262 ( .A1(n5069), .A2(n6420), .B1(INSTQUEUE_REG_13__6__SCAN_IN), 
        .B2(n5068), .ZN(n5064) );
  OAI21_X1 U6263 ( .B1(n5065), .B2(n5071), .A(n5064), .ZN(n5066) );
  AOI21_X1 U6264 ( .B1(n5074), .B2(n6383), .A(n5066), .ZN(n5067) );
  OAI21_X1 U6265 ( .B1(n6386), .B2(n5076), .A(n5067), .ZN(U3130) );
  AOI22_X1 U6266 ( .A1(n5069), .A2(n6388), .B1(INSTQUEUE_REG_13__7__SCAN_IN), 
        .B2(n5068), .ZN(n5070) );
  OAI21_X1 U6267 ( .B1(n5072), .B2(n5071), .A(n5070), .ZN(n5073) );
  AOI21_X1 U6268 ( .B1(n5074), .B2(n6392), .A(n5073), .ZN(n5075) );
  OAI21_X1 U6269 ( .B1(n6396), .B2(n5076), .A(n5075), .ZN(U3131) );
  AOI22_X1 U6270 ( .A1(EBX_REG_7__SCAN_IN), .A2(n6072), .B1(n6047), .B2(n6288), 
        .ZN(n5077) );
  OAI211_X1 U6271 ( .C1(n6078), .C2(n5078), .A(n5077), .B(n6335), .ZN(n5086)
         );
  NOR3_X1 U6272 ( .A1(n6065), .A2(REIP_REG_6__SCAN_IN), .A3(n5079), .ZN(n6032)
         );
  OAI21_X1 U6273 ( .B1(n6065), .B2(n5080), .A(n6046), .ZN(n6035) );
  OAI21_X1 U6274 ( .B1(n6032), .B2(n6035), .A(REIP_REG_7__SCAN_IN), .ZN(n5083)
         );
  OR3_X1 U6275 ( .A1(n6065), .A2(REIP_REG_7__SCAN_IN), .A3(n5081), .ZN(n5082)
         );
  OAI211_X1 U6276 ( .C1(n6071), .C2(n5084), .A(n5083), .B(n5082), .ZN(n5085)
         );
  AOI211_X1 U6277 ( .C1(n5087), .C2(n6036), .A(n5086), .B(n5085), .ZN(n5088)
         );
  INV_X1 U6278 ( .A(n5088), .ZN(U2820) );
  NOR2_X1 U6279 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5089), .ZN(n5123)
         );
  AOI22_X1 U6280 ( .A1(n5091), .A2(n5139), .B1(n6356), .B2(n5090), .ZN(n5120)
         );
  OAI22_X1 U6281 ( .A1(n5121), .A2(n6425), .B1(n5120), .B2(n5148), .ZN(n5092)
         );
  AOI21_X1 U6282 ( .B1(n6415), .B2(n5123), .A(n5092), .ZN(n5101) );
  INV_X1 U6283 ( .A(n5132), .ZN(n6350) );
  OAI211_X1 U6284 ( .C1(n6581), .C2(n5123), .A(n6350), .B(n5093), .ZN(n5094)
         );
  INV_X1 U6285 ( .A(n5094), .ZN(n5099) );
  NOR2_X1 U6286 ( .A1(n5139), .A2(n5835), .ZN(n5095) );
  OAI211_X1 U6287 ( .C1(n6348), .C2(n5095), .A(n5121), .B(n5127), .ZN(n5098)
         );
  NAND2_X1 U6288 ( .A1(n5096), .A2(n5128), .ZN(n5097) );
  NAND3_X1 U6289 ( .A1(n5099), .A2(n5098), .A3(n5097), .ZN(n5124) );
  NAND2_X1 U6290 ( .A1(n5124), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n5100) );
  OAI211_X1 U6291 ( .C1(n5127), .C2(n6386), .A(n5101), .B(n5100), .ZN(U3090)
         );
  OAI22_X1 U6292 ( .A1(n5121), .A2(n6458), .B1(n5120), .B2(n5171), .ZN(n5102)
         );
  AOI21_X1 U6293 ( .B1(n6411), .B2(n5123), .A(n5102), .ZN(n5104) );
  NAND2_X1 U6294 ( .A1(n5124), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n5103) );
  OAI211_X1 U6295 ( .C1(n5127), .C2(n6449), .A(n5104), .B(n5103), .ZN(U3089)
         );
  OAI22_X1 U6296 ( .A1(n5121), .A2(n6446), .B1(n5120), .B2(n5144), .ZN(n5105)
         );
  AOI21_X1 U6297 ( .B1(n6376), .B2(n5123), .A(n5105), .ZN(n5107) );
  NAND2_X1 U6298 ( .A1(n5124), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n5106) );
  OAI211_X1 U6299 ( .C1(n5127), .C2(n6441), .A(n5107), .B(n5106), .ZN(U3088)
         );
  OAI22_X1 U6300 ( .A1(n5121), .A2(n5158), .B1(n5120), .B2(n5157), .ZN(n5108)
         );
  AOI21_X1 U6301 ( .B1(n6367), .B2(n5123), .A(n5108), .ZN(n5110) );
  NAND2_X1 U6302 ( .A1(n5124), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n5109) );
  OAI211_X1 U6303 ( .C1(n5127), .C2(n6371), .A(n5110), .B(n5109), .ZN(U3086)
         );
  OAI22_X1 U6304 ( .A1(n5121), .A2(n6410), .B1(n5120), .B2(n5140), .ZN(n5111)
         );
  AOI21_X1 U6305 ( .B1(n6405), .B2(n5123), .A(n5111), .ZN(n5113) );
  NAND2_X1 U6306 ( .A1(n5124), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n5112) );
  OAI211_X1 U6307 ( .C1(n5127), .C2(n6375), .A(n5113), .B(n5112), .ZN(U3087)
         );
  OAI22_X1 U6308 ( .A1(n5121), .A2(n6432), .B1(n5120), .B2(n5166), .ZN(n5114)
         );
  AOI21_X1 U6309 ( .B1(n6397), .B2(n5123), .A(n5114), .ZN(n5116) );
  NAND2_X1 U6310 ( .A1(n5124), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n5115) );
  OAI211_X1 U6311 ( .C1(n5127), .C2(n6427), .A(n5116), .B(n5115), .ZN(U3084)
         );
  OAI22_X1 U6312 ( .A1(n5121), .A2(n6439), .B1(n5120), .B2(n5162), .ZN(n5117)
         );
  AOI21_X1 U6313 ( .B1(n6401), .B2(n5123), .A(n5117), .ZN(n5119) );
  NAND2_X1 U6314 ( .A1(n5124), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n5118) );
  OAI211_X1 U6315 ( .C1(n5127), .C2(n6434), .A(n5119), .B(n5118), .ZN(U3085)
         );
  OAI22_X1 U6316 ( .A1(n5121), .A2(n5153), .B1(n5120), .B2(n5152), .ZN(n5122)
         );
  AOI21_X1 U6317 ( .B1(n6390), .B2(n5123), .A(n5122), .ZN(n5126) );
  NAND2_X1 U6318 ( .A1(n5124), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n5125) );
  OAI211_X1 U6319 ( .C1(n5127), .C2(n6396), .A(n5126), .B(n5125), .ZN(U3091)
         );
  NOR2_X1 U6320 ( .A1(n5137), .A2(n5835), .ZN(n5129) );
  AOI21_X1 U6321 ( .B1(n5129), .B2(n5178), .A(n5128), .ZN(n5136) );
  NOR2_X1 U6322 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5130), .ZN(n5175)
         );
  INV_X1 U6323 ( .A(n5175), .ZN(n5133) );
  AOI211_X1 U6324 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n5133), .A(n5132), .B(
        n5131), .ZN(n5134) );
  NAND2_X1 U6325 ( .A1(n5170), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n5143) );
  AOI22_X1 U6326 ( .A1(n6348), .A2(n5139), .B1(n6356), .B2(n5138), .ZN(n5172)
         );
  OAI22_X1 U6327 ( .A1(n5173), .A2(n6410), .B1(n5172), .B2(n5140), .ZN(n5141)
         );
  AOI21_X1 U6328 ( .B1(n6405), .B2(n5175), .A(n5141), .ZN(n5142) );
  OAI211_X1 U6329 ( .C1(n5178), .C2(n6375), .A(n5143), .B(n5142), .ZN(U3023)
         );
  NAND2_X1 U6330 ( .A1(n5170), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n5147) );
  OAI22_X1 U6331 ( .A1(n5173), .A2(n6446), .B1(n5172), .B2(n5144), .ZN(n5145)
         );
  AOI21_X1 U6332 ( .B1(n6376), .B2(n5175), .A(n5145), .ZN(n5146) );
  OAI211_X1 U6333 ( .C1(n5178), .C2(n6441), .A(n5147), .B(n5146), .ZN(U3024)
         );
  NAND2_X1 U6334 ( .A1(n5170), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n5151) );
  OAI22_X1 U6335 ( .A1(n5173), .A2(n6425), .B1(n5172), .B2(n5148), .ZN(n5149)
         );
  AOI21_X1 U6336 ( .B1(n6415), .B2(n5175), .A(n5149), .ZN(n5150) );
  OAI211_X1 U6337 ( .C1(n5178), .C2(n6386), .A(n5151), .B(n5150), .ZN(U3026)
         );
  NAND2_X1 U6338 ( .A1(n5170), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n5156) );
  OAI22_X1 U6339 ( .A1(n5173), .A2(n5153), .B1(n5172), .B2(n5152), .ZN(n5154)
         );
  AOI21_X1 U6340 ( .B1(n6390), .B2(n5175), .A(n5154), .ZN(n5155) );
  OAI211_X1 U6341 ( .C1(n5178), .C2(n6396), .A(n5156), .B(n5155), .ZN(U3027)
         );
  NAND2_X1 U6342 ( .A1(n5170), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n5161) );
  OAI22_X1 U6343 ( .A1(n5173), .A2(n5158), .B1(n5172), .B2(n5157), .ZN(n5159)
         );
  AOI21_X1 U6344 ( .B1(n6367), .B2(n5175), .A(n5159), .ZN(n5160) );
  OAI211_X1 U6345 ( .C1(n5178), .C2(n6371), .A(n5161), .B(n5160), .ZN(U3022)
         );
  NAND2_X1 U6346 ( .A1(n5170), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n5165) );
  OAI22_X1 U6347 ( .A1(n5173), .A2(n6439), .B1(n5172), .B2(n5162), .ZN(n5163)
         );
  AOI21_X1 U6348 ( .B1(n6401), .B2(n5175), .A(n5163), .ZN(n5164) );
  OAI211_X1 U6349 ( .C1(n5178), .C2(n6434), .A(n5165), .B(n5164), .ZN(U3021)
         );
  NAND2_X1 U6350 ( .A1(n5170), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n5169) );
  OAI22_X1 U6351 ( .A1(n5173), .A2(n6432), .B1(n5172), .B2(n5166), .ZN(n5167)
         );
  AOI21_X1 U6352 ( .B1(n6397), .B2(n5175), .A(n5167), .ZN(n5168) );
  OAI211_X1 U6353 ( .C1(n5178), .C2(n6427), .A(n5169), .B(n5168), .ZN(U3020)
         );
  NAND2_X1 U6354 ( .A1(n5170), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n5177) );
  OAI22_X1 U6355 ( .A1(n5173), .A2(n6458), .B1(n5172), .B2(n5171), .ZN(n5174)
         );
  AOI21_X1 U6356 ( .B1(n6411), .B2(n5175), .A(n5174), .ZN(n5176) );
  OAI211_X1 U6357 ( .C1(n5178), .C2(n6449), .A(n5177), .B(n5176), .ZN(U3025)
         );
  NAND2_X1 U6358 ( .A1(n5213), .A2(n5212), .ZN(n5179) );
  NAND2_X1 U6359 ( .A1(n5223), .A2(n5179), .ZN(n6008) );
  INV_X1 U6360 ( .A(EBX_REG_9__SCAN_IN), .ZN(n5182) );
  OAI21_X1 U6361 ( .B1(n5181), .B2(n5180), .A(n5227), .ZN(n6009) );
  OAI222_X1 U6362 ( .A1(n6008), .A2(n5576), .B1(n5182), .B2(n6095), .C1(n5555), 
        .C2(n6009), .ZN(U2850) );
  INV_X1 U6363 ( .A(DATAI_9_), .ZN(n5183) );
  INV_X1 U6364 ( .A(EAX_REG_9__SCAN_IN), .ZN(n6190) );
  OAI222_X1 U6365 ( .A1(n6008), .A2(n5878), .B1(n5305), .B2(n5183), .C1(n5397), 
        .C2(n6190), .ZN(U2882) );
  XNOR2_X1 U6366 ( .A(n3437), .B(n5184), .ZN(n5185) );
  XNOR2_X1 U6367 ( .A(n5186), .B(n5185), .ZN(n6276) );
  NAND2_X1 U6368 ( .A1(n6276), .A2(n6243), .ZN(n5190) );
  INV_X1 U6369 ( .A(REIP_REG_9__SCAN_IN), .ZN(n5532) );
  NOR2_X1 U6370 ( .A1(n6335), .A2(n5532), .ZN(n6271) );
  NOR2_X1 U6371 ( .A1(n6249), .A2(n5187), .ZN(n5188) );
  AOI211_X1 U6372 ( .C1(n6239), .C2(PHYADDRPOINTER_REG_9__SCAN_IN), .A(n6271), 
        .B(n5188), .ZN(n5189) );
  OAI211_X1 U6373 ( .C1(n5697), .C2(n6008), .A(n5190), .B(n5189), .ZN(U2977)
         );
  NAND2_X1 U6374 ( .A1(n6595), .A2(n3461), .ZN(n5191) );
  OR2_X1 U6375 ( .A1(n5193), .A2(n5192), .ZN(n6061) );
  INV_X1 U6376 ( .A(n6061), .ZN(n6073) );
  OAI21_X1 U6377 ( .B1(n6059), .B2(n5194), .A(PHYADDRPOINTER_REG_0__SCAN_IN), 
        .ZN(n5195) );
  OAI21_X1 U6378 ( .B1(n6030), .B2(n4371), .A(n5195), .ZN(n5199) );
  INV_X1 U6379 ( .A(REIP_REG_0__SCAN_IN), .ZN(n5196) );
  OAI22_X1 U6380 ( .A1(n6087), .A2(n5197), .B1(n5488), .B2(n5196), .ZN(n5198)
         );
  AOI211_X1 U6381 ( .C1(n5412), .C2(n6073), .A(n5199), .B(n5198), .ZN(n5200)
         );
  OAI21_X1 U6382 ( .B1(n6058), .B2(n5201), .A(n5200), .ZN(U2827) );
  INV_X1 U6383 ( .A(n6035), .ZN(n5204) );
  AOI21_X1 U6384 ( .B1(n6083), .B2(n5202), .A(REIP_REG_5__SCAN_IN), .ZN(n5203)
         );
  NOR2_X1 U6385 ( .A1(n5204), .A2(n5203), .ZN(n5208) );
  INV_X1 U6386 ( .A(EBX_REG_5__SCAN_IN), .ZN(n5206) );
  AOI22_X1 U6387 ( .A1(PHYADDRPOINTER_REG_5__SCAN_IN), .A2(n6059), .B1(n6047), 
        .B2(n6307), .ZN(n5205) );
  OAI211_X1 U6388 ( .C1(n6030), .C2(n5206), .A(n5205), .B(n6335), .ZN(n5207)
         );
  AOI211_X1 U6389 ( .C1(n5194), .C2(n5209), .A(n5208), .B(n5207), .ZN(n5210)
         );
  OAI21_X1 U6390 ( .B1(n6058), .B2(n5211), .A(n5210), .ZN(U2822) );
  NOR2_X1 U6391 ( .A1(n5213), .A2(n5212), .ZN(n5215) );
  XOR2_X1 U6392 ( .A(n5216), .B(n5280), .Z(n5274) );
  NOR2_X1 U6393 ( .A1(n5999), .A2(n5218), .ZN(n5219) );
  OR2_X1 U6394 ( .A1(n5217), .A2(n5219), .ZN(n5232) );
  OAI22_X1 U6395 ( .A1(n5232), .A2(n5555), .B1(n5237), .B2(n6095), .ZN(n5220)
         );
  AOI21_X1 U6396 ( .B1(n5274), .B2(n4149), .A(n5220), .ZN(n5221) );
  INV_X1 U6397 ( .A(n5221), .ZN(U2847) );
  INV_X1 U6398 ( .A(n5278), .ZN(n5222) );
  AOI21_X1 U6399 ( .B1(n5224), .B2(n5223), .A(n5222), .ZN(n5524) );
  INV_X1 U6400 ( .A(n5225), .ZN(n5997) );
  NAND2_X1 U6401 ( .A1(n5227), .A2(n5226), .ZN(n5228) );
  NAND2_X1 U6402 ( .A1(n5997), .A2(n5228), .ZN(n6266) );
  OAI22_X1 U6403 ( .A1(n6266), .A2(n5555), .B1(n5525), .B2(n6095), .ZN(n5229)
         );
  AOI21_X1 U6404 ( .B1(n5524), .B2(n4149), .A(n5229), .ZN(n5230) );
  INV_X1 U6405 ( .A(n5230), .ZN(U2849) );
  INV_X1 U6406 ( .A(n5524), .ZN(n5231) );
  INV_X1 U6407 ( .A(DATAI_10_), .ZN(n6734) );
  INV_X1 U6408 ( .A(EAX_REG_10__SCAN_IN), .ZN(n6193) );
  OAI222_X1 U6409 ( .A1(n5231), .A2(n5878), .B1(n5305), .B2(n6734), .C1(n5397), 
        .C2(n6193), .ZN(U2881) );
  INV_X1 U6410 ( .A(n5274), .ZN(n5255) );
  INV_X1 U6411 ( .A(n5272), .ZN(n5239) );
  INV_X1 U6412 ( .A(n5232), .ZN(n6250) );
  INV_X1 U6413 ( .A(n5988), .ZN(n5233) );
  NOR2_X1 U6414 ( .A1(n6065), .A2(n5233), .ZN(n6000) );
  INV_X1 U6415 ( .A(n6000), .ZN(n5234) );
  NAND2_X1 U6416 ( .A1(n6046), .A2(n5234), .ZN(n6004) );
  AOI22_X1 U6417 ( .A1(n6047), .A2(n6250), .B1(REIP_REG_12__SCAN_IN), .B2(
        n6004), .ZN(n5236) );
  NOR3_X1 U6418 ( .A1(n6065), .A2(REIP_REG_12__SCAN_IN), .A3(n5988), .ZN(n5989) );
  AOI211_X1 U6419 ( .C1(n6059), .C2(PHYADDRPOINTER_REG_12__SCAN_IN), .A(n2993), 
        .B(n5989), .ZN(n5235) );
  OAI211_X1 U6420 ( .C1(n5237), .C2(n6030), .A(n5236), .B(n5235), .ZN(n5238)
         );
  AOI21_X1 U6421 ( .B1(n5194), .B2(n5239), .A(n5238), .ZN(n5240) );
  OAI21_X1 U6422 ( .B1(n5255), .B2(n5971), .A(n5240), .ZN(U2815) );
  INV_X1 U6423 ( .A(n5241), .ZN(n5244) );
  INV_X1 U6424 ( .A(n5242), .ZN(n5243) );
  NAND2_X1 U6425 ( .A1(n5244), .A2(n5243), .ZN(n5245) );
  AND2_X1 U6426 ( .A1(n5246), .A2(n5245), .ZN(n6089) );
  INV_X1 U6427 ( .A(n6089), .ZN(n5247) );
  INV_X1 U6428 ( .A(DATAI_13_), .ZN(n6700) );
  INV_X1 U6429 ( .A(EAX_REG_13__SCAN_IN), .ZN(n6203) );
  OAI222_X1 U6430 ( .A1(n5247), .A2(n5878), .B1(n5305), .B2(n6700), .C1(n5397), 
        .C2(n6203), .ZN(U2878) );
  NAND2_X1 U6431 ( .A1(n6212), .A2(n5248), .ZN(n5251) );
  XOR2_X1 U6432 ( .A(n5251), .B(n5249), .Z(n6264) );
  AOI22_X1 U6433 ( .A1(n6239), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .B1(n2993), 
        .B2(REIP_REG_10__SCAN_IN), .ZN(n5252) );
  OAI21_X1 U6434 ( .B1(n5528), .B2(n6249), .A(n5252), .ZN(n5253) );
  AOI21_X1 U6435 ( .B1(n5524), .B2(n6244), .A(n5253), .ZN(n5254) );
  OAI21_X1 U6436 ( .B1(n6264), .B2(n6221), .A(n5254), .ZN(U2976) );
  INV_X1 U6437 ( .A(EAX_REG_12__SCAN_IN), .ZN(n6199) );
  INV_X1 U6438 ( .A(DATAI_12_), .ZN(n6697) );
  OAI222_X1 U6439 ( .A1(n5878), .A2(n5255), .B1(n5397), .B2(n6199), .C1(n6697), 
        .C2(n5305), .ZN(U2879) );
  OR2_X1 U6440 ( .A1(n5258), .A2(n5257), .ZN(n5259) );
  AND2_X1 U6441 ( .A1(n5256), .A2(n5259), .ZN(n5984) );
  NAND2_X1 U6442 ( .A1(n5905), .A2(n5260), .ZN(n5261) );
  NAND2_X1 U6443 ( .A1(n5302), .A2(n5261), .ZN(n5987) );
  OAI22_X1 U6444 ( .A1(n5987), .A2(n5555), .B1(n5979), .B2(n6095), .ZN(n5262)
         );
  AOI21_X1 U6445 ( .B1(n5984), .B2(n4149), .A(n5262), .ZN(n5263) );
  INV_X1 U6446 ( .A(n5263), .ZN(U2845) );
  INV_X1 U6447 ( .A(n5984), .ZN(n5265) );
  INV_X1 U6448 ( .A(DATAI_14_), .ZN(n5264) );
  INV_X1 U6449 ( .A(EAX_REG_14__SCAN_IN), .ZN(n6206) );
  OAI222_X1 U6450 ( .A1(n5265), .A2(n5878), .B1(n5305), .B2(n5264), .C1(n5397), 
        .C2(n6206), .ZN(U2877) );
  INV_X1 U6451 ( .A(n5267), .ZN(n5268) );
  NAND2_X1 U6452 ( .A1(n5268), .A2(n5891), .ZN(n5269) );
  XNOR2_X1 U6453 ( .A(n5270), .B(n5269), .ZN(n6251) );
  INV_X1 U6454 ( .A(n6251), .ZN(n5276) );
  AOI22_X1 U6455 ( .A1(n6239), .A2(PHYADDRPOINTER_REG_12__SCAN_IN), .B1(n2993), 
        .B2(REIP_REG_12__SCAN_IN), .ZN(n5271) );
  OAI21_X1 U6456 ( .B1(n5272), .B2(n6249), .A(n5271), .ZN(n5273) );
  AOI21_X1 U6457 ( .B1(n5274), .B2(n6244), .A(n5273), .ZN(n5275) );
  OAI21_X1 U6458 ( .B1(n5276), .B2(n6221), .A(n5275), .ZN(U2974) );
  INV_X1 U6459 ( .A(n6218), .ZN(n5281) );
  INV_X1 U6460 ( .A(DATAI_11_), .ZN(n6699) );
  INV_X1 U6461 ( .A(EAX_REG_11__SCAN_IN), .ZN(n6196) );
  OAI222_X1 U6462 ( .A1(n5281), .A2(n5878), .B1(n5305), .B2(n6699), .C1(n5397), 
        .C2(n6196), .ZN(U2880) );
  OAI21_X1 U6463 ( .B1(n5283), .B2(n5285), .A(n5570), .ZN(n5696) );
  NAND2_X1 U6464 ( .A1(n5287), .A2(n5288), .ZN(n5289) );
  AND2_X1 U6465 ( .A1(n5575), .A2(n5289), .ZN(n5823) );
  INV_X1 U6466 ( .A(n5944), .ZN(n5290) );
  NAND2_X1 U6467 ( .A1(n6083), .A2(n5290), .ZN(n5294) );
  INV_X1 U6468 ( .A(EBX_REG_17__SCAN_IN), .ZN(n5309) );
  OAI22_X1 U6469 ( .A1(n5309), .A2(n6030), .B1(n5690), .B2(n6078), .ZN(n5291)
         );
  AOI211_X1 U6470 ( .C1(n5194), .C2(n5693), .A(n5291), .B(n2993), .ZN(n5293)
         );
  NAND2_X1 U6471 ( .A1(n5294), .A2(n6046), .ZN(n5945) );
  NAND2_X1 U6472 ( .A1(n5945), .A2(REIP_REG_17__SCAN_IN), .ZN(n5292) );
  OAI211_X1 U6473 ( .C1(n5295), .C2(n5294), .A(n5293), .B(n5292), .ZN(n5296)
         );
  AOI21_X1 U6474 ( .B1(n5823), .B2(n6047), .A(n5296), .ZN(n5297) );
  OAI21_X1 U6475 ( .B1(n5696), .B2(n5971), .A(n5297), .ZN(U2810) );
  INV_X1 U6476 ( .A(n5311), .ZN(n5299) );
  AOI21_X1 U6477 ( .B1(n5300), .B2(n5256), .A(n5299), .ZN(n5705) );
  INV_X1 U6478 ( .A(n5705), .ZN(n5972) );
  INV_X1 U6479 ( .A(EBX_REG_15__SCAN_IN), .ZN(n5304) );
  AOI21_X1 U6480 ( .B1(n5303), .B2(n5302), .A(n5314), .ZN(n5898) );
  INV_X1 U6481 ( .A(n5898), .ZN(n5976) );
  OAI222_X1 U6482 ( .A1(n5972), .A2(n5576), .B1(n6095), .B2(n5304), .C1(n5976), 
        .C2(n5555), .ZN(U2844) );
  INV_X1 U6483 ( .A(DATAI_15_), .ZN(n6705) );
  INV_X1 U6484 ( .A(EAX_REG_15__SCAN_IN), .ZN(n6211) );
  OAI222_X1 U6485 ( .A1(n5972), .A2(n5878), .B1(n6705), .B2(n5305), .C1(n5397), 
        .C2(n6211), .ZN(U2876) );
  AOI22_X1 U6486 ( .A1(n6099), .A2(DATAI_17_), .B1(n6102), .B2(
        EAX_REG_17__SCAN_IN), .ZN(n5307) );
  NAND2_X1 U6487 ( .A1(n6103), .A2(DATAI_1_), .ZN(n5306) );
  OAI211_X1 U6488 ( .C1(n5696), .C2(n5878), .A(n5307), .B(n5306), .ZN(U2874)
         );
  INV_X1 U6489 ( .A(n5823), .ZN(n5308) );
  OAI222_X1 U6490 ( .A1(n5696), .A2(n5576), .B1(n6095), .B2(n5309), .C1(n5308), 
        .C2(n5555), .ZN(U2842) );
  AND2_X1 U6491 ( .A1(n5311), .A2(n5310), .ZN(n5312) );
  NOR2_X1 U6492 ( .A1(n5283), .A2(n5312), .ZN(n6101) );
  OR2_X1 U6493 ( .A1(n5314), .A2(n5313), .ZN(n5315) );
  NAND2_X1 U6494 ( .A1(n5287), .A2(n5315), .ZN(n5965) );
  OAI22_X1 U6495 ( .A1(n5965), .A2(n5555), .B1(n5960), .B2(n6095), .ZN(n5317)
         );
  AOI21_X1 U6496 ( .B1(n6101), .B2(n4149), .A(n5317), .ZN(n5318) );
  INV_X1 U6497 ( .A(n5318), .ZN(U2843) );
  NAND2_X1 U6498 ( .A1(n5319), .A2(n5320), .ZN(n5671) );
  AND2_X1 U6499 ( .A1(n5671), .A2(n5321), .ZN(n5324) );
  XNOR2_X1 U6500 ( .A(n3437), .B(n5322), .ZN(n5323) );
  XNOR2_X1 U6501 ( .A(n5324), .B(n5323), .ZN(n5369) );
  INV_X1 U6502 ( .A(n5911), .ZN(n5325) );
  NOR3_X1 U6503 ( .A1(n5326), .A2(n5387), .A3(n5325), .ZN(n5328) );
  NOR2_X1 U6504 ( .A1(n5334), .A2(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n5910)
         );
  OAI211_X1 U6505 ( .C1(n6334), .C2(n5328), .A(n5327), .B(n5910), .ZN(n5329)
         );
  INV_X1 U6506 ( .A(n5329), .ZN(n5908) );
  INV_X1 U6507 ( .A(n5339), .ZN(n5332) );
  INV_X1 U6508 ( .A(n6298), .ZN(n5338) );
  NOR2_X1 U6509 ( .A1(n5336), .A2(n5338), .ZN(n6339) );
  AOI21_X1 U6510 ( .B1(n5784), .B2(n5337), .A(n5331), .ZN(n5330) );
  INV_X1 U6511 ( .A(n5330), .ZN(n6332) );
  NOR2_X1 U6512 ( .A1(n6339), .A2(n6332), .ZN(n6329) );
  NOR2_X1 U6513 ( .A1(n5331), .A2(n6297), .ZN(n6262) );
  AOI21_X1 U6514 ( .B1(n5332), .B2(n6329), .A(n6262), .ZN(n6258) );
  AOI211_X1 U6515 ( .C1(n5334), .C2(n5333), .A(n5908), .B(n6258), .ZN(n5335)
         );
  OAI21_X1 U6516 ( .B1(n5350), .B2(n5909), .A(n5335), .ZN(n5907) );
  NOR2_X1 U6517 ( .A1(n5339), .A2(n6314), .ZN(n6257) );
  NAND2_X1 U6518 ( .A1(n5350), .A2(n6257), .ZN(n5340) );
  NOR2_X1 U6519 ( .A1(n5340), .A2(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n5343)
         );
  INV_X1 U6520 ( .A(REIP_REG_14__SCAN_IN), .ZN(n5341) );
  OR2_X1 U6521 ( .A1(n6335), .A2(n5341), .ZN(n5364) );
  OAI21_X1 U6522 ( .B1(n5987), .B2(n6337), .A(n5364), .ZN(n5342) );
  AOI211_X1 U6523 ( .C1(n5907), .C2(INSTADDRPOINTER_REG_14__SCAN_IN), .A(n5343), .B(n5342), .ZN(n5344) );
  OAI21_X1 U6524 ( .B1(n5369), .B2(n6300), .A(n5344), .ZN(U3004) );
  NAND2_X1 U6525 ( .A1(n5671), .A2(n5345), .ZN(n5347) );
  NAND2_X1 U6526 ( .A1(n5347), .A2(n5346), .ZN(n5349) );
  XNOR2_X1 U6527 ( .A(n3437), .B(n5674), .ZN(n5348) );
  XNOR2_X1 U6528 ( .A(n5349), .B(n5348), .ZN(n5363) );
  NAND3_X1 U6529 ( .A1(INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n5350), .A3(n6257), .ZN(n5902) );
  AOI21_X1 U6530 ( .B1(n5675), .B2(n5674), .A(n5902), .ZN(n5356) );
  AND2_X1 U6531 ( .A1(n6297), .A2(n5351), .ZN(n5352) );
  OR2_X1 U6532 ( .A1(n6258), .A2(n5352), .ZN(n5896) );
  NAND2_X1 U6533 ( .A1(n5896), .A2(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5353) );
  NAND2_X1 U6534 ( .A1(n2993), .A2(REIP_REG_16__SCAN_IN), .ZN(n5358) );
  OAI211_X1 U6535 ( .C1(n6337), .C2(n5965), .A(n5353), .B(n5358), .ZN(n5354)
         );
  AOI21_X1 U6536 ( .B1(n5356), .B2(n5355), .A(n5354), .ZN(n5357) );
  OAI21_X1 U6537 ( .B1(n5363), .B2(n6300), .A(n5357), .ZN(U3002) );
  INV_X1 U6538 ( .A(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n5360) );
  NAND2_X1 U6539 ( .A1(n6217), .A2(n5962), .ZN(n5359) );
  OAI211_X1 U6540 ( .C1(n5691), .C2(n5360), .A(n5359), .B(n5358), .ZN(n5361)
         );
  AOI21_X1 U6541 ( .B1(n6101), .B2(n6244), .A(n5361), .ZN(n5362) );
  OAI21_X1 U6542 ( .B1(n5363), .B2(n6221), .A(n5362), .ZN(U2970) );
  INV_X1 U6543 ( .A(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n5365) );
  OAI21_X1 U6544 ( .B1(n5691), .B2(n5365), .A(n5364), .ZN(n5366) );
  AOI21_X1 U6545 ( .B1(n6217), .B2(n5983), .A(n5366), .ZN(n5368) );
  NAND2_X1 U6546 ( .A1(n5984), .A2(n6244), .ZN(n5367) );
  OAI211_X1 U6547 ( .C1(n5369), .C2(n6221), .A(n5368), .B(n5367), .ZN(U2972)
         );
  AND2_X1 U6548 ( .A1(n5568), .A2(n5371), .ZN(n5373) );
  OR2_X1 U6549 ( .A1(n5373), .A2(n5558), .ZN(n5872) );
  INV_X1 U6550 ( .A(EBX_REG_19__SCAN_IN), .ZN(n5377) );
  MUX2_X1 U6551 ( .A(n5563), .B(n5375), .S(n5374), .Z(n5574) );
  OR2_X1 U6552 ( .A1(n5575), .A2(n5574), .ZN(n5572) );
  XNOR2_X1 U6553 ( .A(n5572), .B(n5376), .ZN(n5876) );
  OAI222_X1 U6554 ( .A1(n5872), .A2(n5576), .B1(n6095), .B2(n5377), .C1(n5555), 
        .C2(n5876), .ZN(U2840) );
  AOI22_X1 U6555 ( .A1(n6099), .A2(DATAI_29_), .B1(n6102), .B2(
        EAX_REG_29__SCAN_IN), .ZN(n5379) );
  NAND2_X1 U6556 ( .A1(n6103), .A2(DATAI_13_), .ZN(n5378) );
  OAI211_X1 U6557 ( .C1(n5420), .C2(n5878), .A(n5379), .B(n5378), .ZN(U2862)
         );
  OAI222_X1 U6558 ( .A1(n5576), .A2(n5420), .B1(n5380), .B2(n6095), .C1(n5430), 
        .C2(n5555), .ZN(U2830) );
  AOI21_X1 U6559 ( .B1(n5381), .B2(n5506), .A(n5476), .ZN(n5545) );
  AOI21_X1 U6560 ( .B1(n5756), .B2(INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5382) );
  NOR2_X1 U6561 ( .A1(n5751), .A2(n5382), .ZN(n5383) );
  AOI211_X1 U6562 ( .C1(n5545), .C2(n6323), .A(n5384), .B(n5383), .ZN(n5385)
         );
  OAI21_X1 U6563 ( .B1(n5386), .B2(n6300), .A(n5385), .ZN(U2994) );
  NOR2_X1 U6564 ( .A1(n5413), .A2(n5387), .ZN(n5414) );
  AOI22_X1 U6565 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n4234), .B1(
        INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n6331), .ZN(n5388) );
  INV_X1 U6566 ( .A(n5388), .ZN(n5846) );
  INV_X1 U6567 ( .A(n5415), .ZN(n6583) );
  NOR2_X1 U6568 ( .A1(n6583), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n5391)
         );
  INV_X1 U6569 ( .A(n5389), .ZN(n5390) );
  AOI222_X1 U6570 ( .A1(n5414), .A2(n5846), .B1(n5392), .B2(n5391), .C1(n5390), 
        .C2(n5840), .ZN(n5395) );
  OAI22_X1 U6571 ( .A1(n6459), .A2(n6500), .B1(n6579), .B2(n6696), .ZN(n5919)
         );
  AOI21_X1 U6572 ( .B1(STATE2_REG_3__SCAN_IN), .B2(n6498), .A(n5919), .ZN(
        n5917) );
  INV_X1 U6573 ( .A(n5392), .ZN(n5393) );
  AOI21_X1 U6574 ( .B1(n5415), .B2(n5393), .A(n5917), .ZN(n5394) );
  OAI22_X1 U6575 ( .A1(n5395), .A2(n5917), .B1(n5394), .B2(n3182), .ZN(U3459)
         );
  AND2_X1 U6576 ( .A1(n5397), .A2(n5396), .ZN(n5398) );
  AOI22_X1 U6577 ( .A1(n6099), .A2(DATAI_31_), .B1(EAX_REG_31__SCAN_IN), .B2(
        n6102), .ZN(n5400) );
  NAND2_X1 U6578 ( .A1(n5401), .A2(n5400), .ZN(U2860) );
  NAND2_X1 U6579 ( .A1(n5402), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5403) );
  XNOR2_X1 U6580 ( .A(n5405), .B(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n5718)
         );
  NAND2_X1 U6581 ( .A1(n6217), .A2(n5406), .ZN(n5407) );
  NAND2_X1 U6582 ( .A1(n2993), .A2(REIP_REG_30__SCAN_IN), .ZN(n5712) );
  OAI211_X1 U6583 ( .C1(n5408), .C2(n5691), .A(n5407), .B(n5712), .ZN(n5409)
         );
  AOI21_X1 U6584 ( .B1(n5577), .B2(n6244), .A(n5409), .ZN(n5410) );
  OAI21_X1 U6585 ( .B1(n5718), .B2(n6221), .A(n5410), .ZN(U2956) );
  INV_X1 U6586 ( .A(n5842), .ZN(n5411) );
  AOI22_X1 U6587 ( .A1(n5412), .A2(n5844), .B1(n5411), .B2(n3153), .ZN(n6461)
         );
  OAI21_X1 U6588 ( .B1(n6461), .B2(STATE2_REG_3__SCAN_IN), .A(n5413), .ZN(
        n5416) );
  INV_X1 U6589 ( .A(n5414), .ZN(n5847) );
  AOI22_X1 U6590 ( .A1(n5416), .A2(n5847), .B1(n5415), .B2(n3153), .ZN(n5419)
         );
  AOI21_X1 U6591 ( .B1(n5417), .B2(n5840), .A(n5917), .ZN(n5418) );
  OAI22_X1 U6592 ( .A1(n5419), .A2(n5917), .B1(n5418), .B2(n3153), .ZN(U3461)
         );
  INV_X1 U6593 ( .A(n5420), .ZN(n5421) );
  NAND2_X1 U6594 ( .A1(n5421), .A2(n6036), .ZN(n5429) );
  INV_X1 U6595 ( .A(n5422), .ZN(n5442) );
  AOI22_X1 U6596 ( .A1(PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n6059), .B1(n5194), 
        .B2(n5423), .ZN(n5425) );
  NAND2_X1 U6597 ( .A1(n6072), .A2(EBX_REG_29__SCAN_IN), .ZN(n5424) );
  OAI211_X1 U6598 ( .C1(n5426), .C2(REIP_REG_29__SCAN_IN), .A(n5425), .B(n5424), .ZN(n5427) );
  AOI21_X1 U6599 ( .B1(n5442), .B2(REIP_REG_29__SCAN_IN), .A(n5427), .ZN(n5428) );
  OAI211_X1 U6600 ( .C1(n6087), .C2(n5430), .A(n5429), .B(n5428), .ZN(U2798)
         );
  AOI21_X1 U6601 ( .B1(n5432), .B2(n5446), .A(n4325), .ZN(n5603) );
  INV_X1 U6602 ( .A(n5603), .ZN(n5583) );
  AND2_X1 U6603 ( .A1(n5450), .A2(n5433), .ZN(n5435) );
  OR2_X1 U6604 ( .A1(n5435), .A2(n5434), .ZN(n5723) );
  OAI22_X1 U6605 ( .A1(n5436), .A2(n6078), .B1(n6071), .B2(n5601), .ZN(n5437)
         );
  AOI21_X1 U6606 ( .B1(n6072), .B2(EBX_REG_28__SCAN_IN), .A(n5437), .ZN(n5440)
         );
  INV_X1 U6607 ( .A(REIP_REG_28__SCAN_IN), .ZN(n6771) );
  NAND2_X1 U6608 ( .A1(n5438), .A2(n6771), .ZN(n5439) );
  OAI211_X1 U6609 ( .C1(n5723), .C2(n6087), .A(n5440), .B(n5439), .ZN(n5441)
         );
  AOI21_X1 U6610 ( .B1(REIP_REG_28__SCAN_IN), .B2(n5442), .A(n5441), .ZN(n5443) );
  OAI21_X1 U6611 ( .B1(n5583), .B2(n5971), .A(n5443), .ZN(U2799) );
  OAI21_X1 U6612 ( .B1(n5445), .B2(n5447), .A(n5446), .ZN(n5609) );
  INV_X1 U6613 ( .A(n5470), .ZN(n5457) );
  NAND2_X1 U6614 ( .A1(n5464), .A2(n5448), .ZN(n5449) );
  NAND2_X1 U6615 ( .A1(n5450), .A2(n5449), .ZN(n5730) );
  INV_X1 U6616 ( .A(n5612), .ZN(n5451) );
  OAI22_X1 U6617 ( .A1(n5608), .A2(n6078), .B1(n6071), .B2(n5451), .ZN(n5454)
         );
  NOR3_X1 U6618 ( .A1(n5489), .A2(REIP_REG_27__SCAN_IN), .A3(n5452), .ZN(n5453) );
  AOI211_X1 U6619 ( .C1(EBX_REG_27__SCAN_IN), .C2(n6072), .A(n5454), .B(n5453), 
        .ZN(n5455) );
  OAI21_X1 U6620 ( .B1(n5730), .B2(n6087), .A(n5455), .ZN(n5456) );
  AOI21_X1 U6621 ( .B1(REIP_REG_27__SCAN_IN), .B2(n5457), .A(n5456), .ZN(n5458) );
  OAI21_X1 U6622 ( .B1(n5609), .B2(n5971), .A(n5458), .ZN(U2800) );
  NOR2_X1 U6623 ( .A1(n3883), .A2(n5489), .ZN(n5481) );
  AOI21_X1 U6624 ( .B1(n5481), .B2(REIP_REG_25__SCAN_IN), .A(
        REIP_REG_26__SCAN_IN), .ZN(n5471) );
  AOI21_X1 U6625 ( .B1(n5460), .B2(n5472), .A(n5445), .ZN(n5619) );
  NAND2_X1 U6626 ( .A1(n5619), .A2(n6036), .ZN(n5469) );
  OAI22_X1 U6627 ( .A1(n5461), .A2(n6078), .B1(n6071), .B2(n5617), .ZN(n5467)
         );
  INV_X1 U6628 ( .A(n5462), .ZN(n5477) );
  INV_X1 U6629 ( .A(n5463), .ZN(n5465) );
  OAI21_X1 U6630 ( .B1(n5477), .B2(n5465), .A(n5464), .ZN(n5736) );
  NOR2_X1 U6631 ( .A1(n5736), .A2(n6087), .ZN(n5466) );
  AOI211_X1 U6632 ( .C1(n6072), .C2(EBX_REG_26__SCAN_IN), .A(n5467), .B(n5466), 
        .ZN(n5468) );
  OAI211_X1 U6633 ( .C1(n5471), .C2(n5470), .A(n5469), .B(n5468), .ZN(U2801)
         );
  OAI21_X1 U6634 ( .B1(n5474), .B2(n5473), .A(n5472), .ZN(n5624) );
  INV_X1 U6635 ( .A(n5475), .ZN(n5479) );
  INV_X1 U6636 ( .A(n5476), .ZN(n5478) );
  AOI21_X1 U6637 ( .B1(n5479), .B2(n5478), .A(n5477), .ZN(n5753) );
  OAI22_X1 U6638 ( .A1(n5488), .A2(n5487), .B1(REIP_REG_24__SCAN_IN), .B2(
        n5489), .ZN(n5480) );
  AOI22_X1 U6639 ( .A1(n5627), .A2(n5194), .B1(REIP_REG_25__SCAN_IN), .B2(
        n5480), .ZN(n5483) );
  INV_X1 U6640 ( .A(REIP_REG_25__SCAN_IN), .ZN(n6749) );
  AOI22_X1 U6641 ( .A1(EBX_REG_25__SCAN_IN), .A2(n6072), .B1(n5481), .B2(n6749), .ZN(n5482) );
  OAI211_X1 U6642 ( .C1(n5623), .C2(n6078), .A(n5483), .B(n5482), .ZN(n5484)
         );
  AOI21_X1 U6643 ( .B1(n5753), .B2(n6047), .A(n5484), .ZN(n5485) );
  OAI21_X1 U6644 ( .B1(n5624), .B2(n5971), .A(n5485), .ZN(U2802) );
  INV_X1 U6645 ( .A(n5486), .ZN(n5593) );
  NOR2_X1 U6646 ( .A1(n5488), .A2(n5487), .ZN(n5503) );
  NOR2_X1 U6647 ( .A1(REIP_REG_24__SCAN_IN), .A2(n5489), .ZN(n5493) );
  OAI22_X1 U6648 ( .A1(n5491), .A2(n6030), .B1(n5490), .B2(n6078), .ZN(n5492)
         );
  AOI211_X1 U6649 ( .C1(n5503), .C2(REIP_REG_24__SCAN_IN), .A(n5493), .B(n5492), .ZN(n5496) );
  AOI22_X1 U6650 ( .A1(n5545), .A2(n6047), .B1(n5494), .B2(n5194), .ZN(n5495)
         );
  OAI211_X1 U6651 ( .C1(n5593), .C2(n5971), .A(n5496), .B(n5495), .ZN(U2803)
         );
  NAND2_X1 U6652 ( .A1(n5551), .A2(n5497), .ZN(n5498) );
  NAND2_X1 U6653 ( .A1(n5499), .A2(n5498), .ZN(n5635) );
  INV_X1 U6654 ( .A(EBX_REG_23__SCAN_IN), .ZN(n5500) );
  OAI22_X1 U6655 ( .A1(n5500), .A2(n6030), .B1(n5634), .B2(n6078), .ZN(n5501)
         );
  AOI221_X1 U6656 ( .B1(REIP_REG_23__SCAN_IN), .B2(n5503), .C1(n5502), .C2(
        n5503), .A(n5501), .ZN(n5510) );
  INV_X1 U6657 ( .A(n5506), .ZN(n5507) );
  AOI21_X1 U6658 ( .B1(n5508), .B2(n5505), .A(n5507), .ZN(n5761) );
  AOI22_X1 U6659 ( .A1(n5761), .A2(n6047), .B1(n5638), .B2(n5194), .ZN(n5509)
         );
  OAI211_X1 U6660 ( .C1(n5635), .C2(n5971), .A(n5510), .B(n5509), .ZN(U2804)
         );
  OR2_X1 U6661 ( .A1(n5511), .A2(n5512), .ZN(n5513) );
  NAND2_X1 U6662 ( .A1(n5549), .A2(n5513), .ZN(n5655) );
  INV_X1 U6663 ( .A(n5655), .ZN(n5882) );
  NAND2_X1 U6664 ( .A1(n6067), .A2(n5514), .ZN(n5860) );
  OAI22_X1 U6665 ( .A1(n5650), .A2(n6078), .B1(n6703), .B2(n5860), .ZN(n5522)
         );
  NOR2_X1 U6666 ( .A1(n5517), .A2(n5516), .ZN(n5518) );
  OR2_X1 U6667 ( .A1(n5515), .A2(n5518), .ZN(n5781) );
  NAND2_X1 U6668 ( .A1(n5519), .A2(n6703), .ZN(n5849) );
  AOI22_X1 U6669 ( .A1(n6072), .A2(EBX_REG_21__SCAN_IN), .B1(n5652), .B2(n5194), .ZN(n5520) );
  OAI211_X1 U6670 ( .C1(n5781), .C2(n6087), .A(n5849), .B(n5520), .ZN(n5521)
         );
  AOI211_X1 U6671 ( .C1(n5882), .C2(n6036), .A(n5522), .B(n5521), .ZN(n5523)
         );
  INV_X1 U6672 ( .A(n5523), .ZN(U2806) );
  NAND2_X1 U6673 ( .A1(n5524), .A2(n6036), .ZN(n5537) );
  OAI22_X1 U6674 ( .A1(n5525), .A2(n6030), .B1(n6087), .B2(n6266), .ZN(n5526)
         );
  AOI211_X1 U6675 ( .C1(n6059), .C2(PHYADDRPOINTER_REG_10__SCAN_IN), .A(n5526), 
        .B(n2993), .ZN(n5536) );
  NOR2_X1 U6676 ( .A1(REIP_REG_10__SCAN_IN), .A2(n5527), .ZN(n5530) );
  INV_X1 U6677 ( .A(n5528), .ZN(n5529) );
  AOI22_X1 U6678 ( .A1(n6083), .A2(n5530), .B1(n5529), .B2(n5194), .ZN(n5535)
         );
  OAI21_X1 U6679 ( .B1(n6065), .B2(n5531), .A(n6046), .ZN(n6019) );
  NAND2_X1 U6680 ( .A1(n5532), .A2(n5531), .ZN(n5533) );
  NOR2_X1 U6681 ( .A1(n6065), .A2(n5533), .ZN(n6013) );
  OAI21_X1 U6682 ( .B1(n6019), .B2(n6013), .A(REIP_REG_10__SCAN_IN), .ZN(n5534) );
  NAND4_X1 U6683 ( .A1(n5537), .A2(n5536), .A3(n5535), .A4(n5534), .ZN(U2817)
         );
  INV_X1 U6684 ( .A(n5538), .ZN(n5540) );
  OAI22_X1 U6685 ( .A1(n5540), .A2(n5555), .B1(n6095), .B2(n5539), .ZN(U2828)
         );
  INV_X1 U6686 ( .A(EBX_REG_28__SCAN_IN), .ZN(n5541) );
  OAI222_X1 U6687 ( .A1(n5576), .A2(n5583), .B1(n5541), .B2(n6095), .C1(n5723), 
        .C2(n5555), .ZN(U2831) );
  INV_X1 U6688 ( .A(EBX_REG_27__SCAN_IN), .ZN(n5542) );
  OAI222_X1 U6689 ( .A1(n5576), .A2(n5609), .B1(n5542), .B2(n6095), .C1(n5730), 
        .C2(n5555), .ZN(U2832) );
  INV_X1 U6690 ( .A(n5619), .ZN(n5588) );
  INV_X1 U6691 ( .A(EBX_REG_26__SCAN_IN), .ZN(n5543) );
  OAI222_X1 U6692 ( .A1(n5576), .A2(n5588), .B1(n5543), .B2(n6095), .C1(n5736), 
        .C2(n5555), .ZN(U2833) );
  AOI22_X1 U6693 ( .A1(n5753), .A2(n6092), .B1(EBX_REG_25__SCAN_IN), .B2(n4150), .ZN(n5544) );
  OAI21_X1 U6694 ( .B1(n5624), .B2(n5576), .A(n5544), .ZN(U2834) );
  AOI22_X1 U6695 ( .A1(n5545), .A2(n6092), .B1(EBX_REG_24__SCAN_IN), .B2(n4150), .ZN(n5546) );
  OAI21_X1 U6696 ( .B1(n5593), .B2(n5576), .A(n5546), .ZN(U2835) );
  AOI22_X1 U6697 ( .A1(n5761), .A2(n6092), .B1(EBX_REG_23__SCAN_IN), .B2(n4150), .ZN(n5547) );
  OAI21_X1 U6698 ( .B1(n5635), .B2(n5576), .A(n5547), .ZN(U2836) );
  NAND2_X1 U6699 ( .A1(n5549), .A2(n5548), .ZN(n5550) );
  NAND2_X1 U6700 ( .A1(n5551), .A2(n5550), .ZN(n5877) );
  INV_X1 U6701 ( .A(EBX_REG_22__SCAN_IN), .ZN(n5554) );
  OR2_X1 U6702 ( .A1(n5515), .A2(n5552), .ZN(n5553) );
  NAND2_X1 U6703 ( .A1(n5505), .A2(n5553), .ZN(n5858) );
  OAI222_X1 U6704 ( .A1(n5576), .A2(n5877), .B1(n5554), .B2(n6095), .C1(n5858), 
        .C2(n5555), .ZN(U2837) );
  INV_X1 U6705 ( .A(EBX_REG_21__SCAN_IN), .ZN(n5556) );
  OAI222_X1 U6706 ( .A1(n5576), .A2(n5655), .B1(n5556), .B2(n6095), .C1(n5781), 
        .C2(n5555), .ZN(U2838) );
  INV_X1 U6707 ( .A(n5557), .ZN(n5560) );
  INV_X1 U6708 ( .A(n5558), .ZN(n5559) );
  AOI21_X1 U6709 ( .B1(n5560), .B2(n5559), .A(n5511), .ZN(n5885) );
  INV_X1 U6710 ( .A(n5885), .ZN(n5567) );
  MUX2_X1 U6711 ( .A(n5563), .B(n5562), .S(n5561), .Z(n5565) );
  XNOR2_X1 U6712 ( .A(n5565), .B(n5564), .ZN(n5863) );
  AOI22_X1 U6713 ( .A1(n5863), .A2(n6092), .B1(EBX_REG_20__SCAN_IN), .B2(n4150), .ZN(n5566) );
  OAI21_X1 U6714 ( .B1(n5567), .B2(n5576), .A(n5566), .ZN(U2839) );
  INV_X1 U6715 ( .A(n5568), .ZN(n5569) );
  AOI21_X1 U6716 ( .B1(n5571), .B2(n5570), .A(n5569), .ZN(n6096) );
  INV_X1 U6717 ( .A(n6096), .ZN(n5948) );
  INV_X1 U6718 ( .A(n5572), .ZN(n5573) );
  AOI21_X1 U6719 ( .B1(n5575), .B2(n5574), .A(n5573), .ZN(n5811) );
  INV_X1 U6720 ( .A(n5811), .ZN(n5947) );
  OAI222_X1 U6721 ( .A1(n5948), .A2(n5576), .B1(n6095), .B2(n3960), .C1(n5947), 
        .C2(n5555), .ZN(U2841) );
  AOI22_X1 U6722 ( .A1(n6099), .A2(DATAI_30_), .B1(n6102), .B2(
        EAX_REG_30__SCAN_IN), .ZN(n5579) );
  NAND2_X1 U6723 ( .A1(n6103), .A2(DATAI_14_), .ZN(n5578) );
  OAI211_X1 U6724 ( .C1(n5580), .C2(n5878), .A(n5579), .B(n5578), .ZN(U2861)
         );
  AOI22_X1 U6725 ( .A1(n6099), .A2(DATAI_28_), .B1(n6102), .B2(
        EAX_REG_28__SCAN_IN), .ZN(n5582) );
  NAND2_X1 U6726 ( .A1(n6103), .A2(DATAI_12_), .ZN(n5581) );
  OAI211_X1 U6727 ( .C1(n5583), .C2(n5878), .A(n5582), .B(n5581), .ZN(U2863)
         );
  AOI22_X1 U6728 ( .A1(n6099), .A2(DATAI_27_), .B1(n6102), .B2(
        EAX_REG_27__SCAN_IN), .ZN(n5585) );
  NAND2_X1 U6729 ( .A1(n6103), .A2(DATAI_11_), .ZN(n5584) );
  OAI211_X1 U6730 ( .C1(n5609), .C2(n5878), .A(n5585), .B(n5584), .ZN(U2864)
         );
  AOI22_X1 U6731 ( .A1(n6099), .A2(DATAI_26_), .B1(n6102), .B2(
        EAX_REG_26__SCAN_IN), .ZN(n5587) );
  NAND2_X1 U6732 ( .A1(n6103), .A2(DATAI_10_), .ZN(n5586) );
  OAI211_X1 U6733 ( .C1(n5588), .C2(n5878), .A(n5587), .B(n5586), .ZN(U2865)
         );
  AOI22_X1 U6734 ( .A1(n6099), .A2(DATAI_25_), .B1(n6102), .B2(
        EAX_REG_25__SCAN_IN), .ZN(n5590) );
  NAND2_X1 U6735 ( .A1(n6103), .A2(DATAI_9_), .ZN(n5589) );
  OAI211_X1 U6736 ( .C1(n5624), .C2(n5878), .A(n5590), .B(n5589), .ZN(U2866)
         );
  AOI22_X1 U6737 ( .A1(n6099), .A2(DATAI_24_), .B1(n6102), .B2(
        EAX_REG_24__SCAN_IN), .ZN(n5592) );
  NAND2_X1 U6738 ( .A1(n6103), .A2(DATAI_8_), .ZN(n5591) );
  OAI211_X1 U6739 ( .C1(n5593), .C2(n5878), .A(n5592), .B(n5591), .ZN(U2867)
         );
  AOI22_X1 U6740 ( .A1(n6099), .A2(DATAI_23_), .B1(n6102), .B2(
        EAX_REG_23__SCAN_IN), .ZN(n5595) );
  NAND2_X1 U6741 ( .A1(n6103), .A2(DATAI_7_), .ZN(n5594) );
  OAI211_X1 U6742 ( .C1(n5635), .C2(n5878), .A(n5595), .B(n5594), .ZN(U2868)
         );
  NAND3_X1 U6743 ( .A1(n5615), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .A3(n5629), .ZN(n5598) );
  NAND2_X1 U6744 ( .A1(n5750), .A2(n5742), .ZN(n5738) );
  OR2_X1 U6745 ( .A1(n5629), .A2(n5738), .ZN(n5597) );
  AOI22_X1 U6746 ( .A1(n5598), .A2(n5605), .B1(INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n5742), .ZN(n5599) );
  XNOR2_X1 U6747 ( .A(n5599), .B(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5727)
         );
  NOR2_X1 U6748 ( .A1(n6335), .A2(n6771), .ZN(n5722) );
  AOI21_X1 U6749 ( .B1(n6239), .B2(PHYADDRPOINTER_REG_28__SCAN_IN), .A(n5722), 
        .ZN(n5600) );
  OAI21_X1 U6750 ( .B1(n5601), .B2(n6249), .A(n5600), .ZN(n5602) );
  AOI21_X1 U6751 ( .B1(n5603), .B2(n6244), .A(n5602), .ZN(n5604) );
  OAI21_X1 U6752 ( .B1(n6221), .B2(n5727), .A(n5604), .ZN(U2958) );
  NAND2_X1 U6753 ( .A1(n5606), .A2(n5605), .ZN(n5607) );
  XNOR2_X1 U6754 ( .A(n5607), .B(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5735)
         );
  NAND2_X1 U6755 ( .A1(n2993), .A2(REIP_REG_27__SCAN_IN), .ZN(n5728) );
  OAI21_X1 U6756 ( .B1(n5691), .B2(n5608), .A(n5728), .ZN(n5611) );
  NOR2_X1 U6757 ( .A1(n5609), .A2(n5697), .ZN(n5610) );
  OAI21_X1 U6758 ( .B1(n5735), .B2(n6221), .A(n5613), .ZN(U2959) );
  XNOR2_X1 U6759 ( .A(n3437), .B(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5614)
         );
  XNOR2_X1 U6760 ( .A(n5615), .B(n5614), .ZN(n5746) );
  NAND2_X1 U6761 ( .A1(n2993), .A2(REIP_REG_26__SCAN_IN), .ZN(n5741) );
  NAND2_X1 U6762 ( .A1(n6239), .A2(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n5616)
         );
  OAI211_X1 U6763 ( .C1(n6249), .C2(n5617), .A(n5741), .B(n5616), .ZN(n5618)
         );
  AOI21_X1 U6764 ( .B1(n5619), .B2(n6244), .A(n5618), .ZN(n5620) );
  OAI21_X1 U6765 ( .B1(n5746), .B2(n6221), .A(n5620), .ZN(U2960) );
  AOI21_X1 U6766 ( .B1(n5596), .B2(n5622), .A(n5621), .ZN(n5755) );
  NAND2_X1 U6767 ( .A1(n2993), .A2(REIP_REG_25__SCAN_IN), .ZN(n5749) );
  OAI21_X1 U6768 ( .B1(n5691), .B2(n5623), .A(n5749), .ZN(n5626) );
  NOR2_X1 U6769 ( .A1(n5624), .A2(n5697), .ZN(n5625) );
  AOI211_X1 U6770 ( .C1(n6217), .C2(n5627), .A(n5626), .B(n5625), .ZN(n5628)
         );
  OAI21_X1 U6771 ( .B1(n5755), .B2(n6221), .A(n5628), .ZN(U2961) );
  NAND4_X1 U6772 ( .A1(n5665), .A2(n5630), .A3(INSTADDRPOINTER_REG_20__SCAN_IN), .A4(n5629), .ZN(n5631) );
  NAND2_X1 U6773 ( .A1(n5632), .A2(n5631), .ZN(n5633) );
  XNOR2_X1 U6774 ( .A(n5633), .B(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5763)
         );
  NAND2_X1 U6775 ( .A1(n2993), .A2(REIP_REG_23__SCAN_IN), .ZN(n5758) );
  OAI21_X1 U6776 ( .B1(n5691), .B2(n5634), .A(n5758), .ZN(n5637) );
  NOR2_X1 U6777 ( .A1(n5635), .A2(n5697), .ZN(n5636) );
  AOI211_X1 U6778 ( .C1(n6217), .C2(n5638), .A(n5637), .B(n5636), .ZN(n5639)
         );
  OAI21_X1 U6779 ( .B1(n5763), .B2(n6221), .A(n5639), .ZN(U2963) );
  AOI21_X1 U6780 ( .B1(INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n3437), .A(n5640), 
        .ZN(n5641) );
  XNOR2_X1 U6781 ( .A(n5643), .B(n5642), .ZN(n5764) );
  NAND2_X1 U6782 ( .A1(n5764), .A2(n6243), .ZN(n5646) );
  NOR2_X1 U6783 ( .A1(n6335), .A2(n6560), .ZN(n5769) );
  NOR2_X1 U6784 ( .A1(n6249), .A2(n5854), .ZN(n5644) );
  AOI211_X1 U6785 ( .C1(n6239), .C2(PHYADDRPOINTER_REG_22__SCAN_IN), .A(n5769), 
        .B(n5644), .ZN(n5645) );
  OAI211_X1 U6786 ( .C1(n5697), .C2(n5877), .A(n5646), .B(n5645), .ZN(U2964)
         );
  OAI21_X1 U6787 ( .B1(n5649), .B2(n5648), .A(n5647), .ZN(n5773) );
  NAND2_X1 U6788 ( .A1(n5773), .A2(n6243), .ZN(n5654) );
  NAND2_X1 U6789 ( .A1(n2993), .A2(REIP_REG_21__SCAN_IN), .ZN(n5774) );
  OAI21_X1 U6790 ( .B1(n5691), .B2(n5650), .A(n5774), .ZN(n5651) );
  AOI21_X1 U6791 ( .B1(n6217), .B2(n5652), .A(n5651), .ZN(n5653) );
  OAI211_X1 U6792 ( .C1(n5697), .C2(n5655), .A(n5654), .B(n5653), .ZN(U2965)
         );
  XNOR2_X1 U6793 ( .A(n3437), .B(n5790), .ZN(n5656) );
  XNOR2_X1 U6794 ( .A(n5657), .B(n5656), .ZN(n5793) );
  NAND2_X1 U6795 ( .A1(n2993), .A2(REIP_REG_20__SCAN_IN), .ZN(n5789) );
  NAND2_X1 U6796 ( .A1(n6239), .A2(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n5658)
         );
  OAI211_X1 U6797 ( .C1(n6249), .C2(n5866), .A(n5789), .B(n5658), .ZN(n5659)
         );
  AOI21_X1 U6798 ( .B1(n5885), .B2(n6244), .A(n5659), .ZN(n5660) );
  OAI21_X1 U6799 ( .B1(n5793), .B2(n6221), .A(n5660), .ZN(U2966) );
  INV_X1 U6800 ( .A(n5661), .ZN(n5664) );
  XNOR2_X1 U6801 ( .A(n5629), .B(n5799), .ZN(n5663) );
  AOI22_X1 U6802 ( .A1(n5665), .A2(n5664), .B1(n5662), .B2(n5663), .ZN(n5794)
         );
  NAND2_X1 U6803 ( .A1(n5794), .A2(n6243), .ZN(n5668) );
  NOR2_X1 U6804 ( .A1(n6335), .A2(n6706), .ZN(n5795) );
  NOR2_X1 U6805 ( .A1(n5691), .A2(n5869), .ZN(n5666) );
  AOI211_X1 U6806 ( .C1(n6217), .C2(n5873), .A(n5795), .B(n5666), .ZN(n5667)
         );
  OAI211_X1 U6807 ( .C1(n5697), .C2(n5872), .A(n5668), .B(n5667), .ZN(U2967)
         );
  INV_X1 U6808 ( .A(n5669), .ZN(n5684) );
  NOR3_X1 U6809 ( .A1(n5684), .A2(n5683), .A3(n5820), .ZN(n5688) );
  NAND4_X1 U6810 ( .A1(n5683), .A2(n5675), .A3(n5674), .A4(n5820), .ZN(n5676)
         );
  NOR2_X1 U6811 ( .A1(n5701), .A2(n5676), .ZN(n5686) );
  NOR2_X1 U6812 ( .A1(n5688), .A2(n5686), .ZN(n5677) );
  XNOR2_X1 U6813 ( .A(n5677), .B(n5786), .ZN(n5814) );
  INV_X1 U6814 ( .A(REIP_REG_18__SCAN_IN), .ZN(n5678) );
  NOR2_X1 U6815 ( .A1(n6335), .A2(n5678), .ZN(n5809) );
  AOI21_X1 U6816 ( .B1(n6239), .B2(PHYADDRPOINTER_REG_18__SCAN_IN), .A(n5809), 
        .ZN(n5679) );
  OAI21_X1 U6817 ( .B1(n5952), .B2(n6249), .A(n5679), .ZN(n5680) );
  AOI21_X1 U6818 ( .B1(n6096), .B2(n6244), .A(n5680), .ZN(n5681) );
  OAI21_X1 U6819 ( .B1(n5814), .B2(n6221), .A(n5681), .ZN(U2968) );
  AOI21_X1 U6820 ( .B1(n5684), .B2(n5820), .A(n5683), .ZN(n5685) );
  AOI21_X1 U6821 ( .B1(INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n5682), .A(n5685), 
        .ZN(n5689) );
  INV_X1 U6822 ( .A(n5686), .ZN(n5687) );
  OAI21_X1 U6823 ( .B1(n5689), .B2(n5688), .A(n5687), .ZN(n5815) );
  NAND2_X1 U6824 ( .A1(n5815), .A2(n6243), .ZN(n5695) );
  NAND2_X1 U6825 ( .A1(n2993), .A2(REIP_REG_17__SCAN_IN), .ZN(n5818) );
  OAI21_X1 U6826 ( .B1(n5691), .B2(n5690), .A(n5818), .ZN(n5692) );
  AOI21_X1 U6827 ( .B1(n6217), .B2(n5693), .A(n5692), .ZN(n5694) );
  OAI211_X1 U6828 ( .C1(n5697), .C2(n5696), .A(n5695), .B(n5694), .ZN(U2969)
         );
  NOR2_X1 U6829 ( .A1(n5699), .A2(n5698), .ZN(n5700) );
  XNOR2_X1 U6830 ( .A(n5701), .B(n5700), .ZN(n5897) );
  AOI22_X1 U6831 ( .A1(n6239), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .B1(n2993), 
        .B2(REIP_REG_15__SCAN_IN), .ZN(n5702) );
  OAI21_X1 U6832 ( .B1(n5703), .B2(n6249), .A(n5702), .ZN(n5704) );
  AOI21_X1 U6833 ( .B1(n5705), .B2(n6244), .A(n5704), .ZN(n5706) );
  OAI21_X1 U6834 ( .B1(n5897), .B2(n6221), .A(n5706), .ZN(U2971) );
  INV_X1 U6835 ( .A(n5707), .ZN(n5716) );
  INV_X1 U6836 ( .A(n6297), .ZN(n5709) );
  AOI211_X1 U6837 ( .C1(n5709), .C2(n5751), .A(n5710), .B(n5708), .ZN(n5715)
         );
  NAND4_X1 U6838 ( .A1(n5711), .A2(n5719), .A3(INSTADDRPOINTER_REG_29__SCAN_IN), .A4(n5710), .ZN(n5713) );
  NAND2_X1 U6839 ( .A1(n5713), .A2(n5712), .ZN(n5714) );
  AOI211_X1 U6840 ( .C1(n5716), .C2(n6323), .A(n5715), .B(n5714), .ZN(n5717)
         );
  OAI21_X1 U6841 ( .B1(n5718), .B2(n6300), .A(n5717), .ZN(U2988) );
  NOR3_X1 U6842 ( .A1(n5729), .A2(n5720), .A3(n5719), .ZN(n5721) );
  AOI211_X1 U6843 ( .C1(INSTADDRPOINTER_REG_28__SCAN_IN), .C2(n5733), .A(n5722), .B(n5721), .ZN(n5726) );
  INV_X1 U6844 ( .A(n5723), .ZN(n5724) );
  NAND2_X1 U6845 ( .A1(n5724), .A2(n6323), .ZN(n5725) );
  OAI211_X1 U6846 ( .C1(n5727), .C2(n6300), .A(n5726), .B(n5725), .ZN(U2990)
         );
  OAI21_X1 U6847 ( .B1(n5729), .B2(INSTADDRPOINTER_REG_27__SCAN_IN), .A(n5728), 
        .ZN(n5732) );
  NOR2_X1 U6848 ( .A1(n5730), .A2(n6337), .ZN(n5731) );
  AOI211_X1 U6849 ( .C1(INSTADDRPOINTER_REG_27__SCAN_IN), .C2(n5733), .A(n5732), .B(n5731), .ZN(n5734) );
  OAI21_X1 U6850 ( .B1(n5735), .B2(n6300), .A(n5734), .ZN(U2991) );
  INV_X1 U6851 ( .A(n5736), .ZN(n5744) );
  INV_X1 U6852 ( .A(n5737), .ZN(n5747) );
  NAND3_X1 U6853 ( .A1(n5747), .A2(n5739), .A3(n5738), .ZN(n5740) );
  OAI211_X1 U6854 ( .C1(n5751), .C2(n5742), .A(n5741), .B(n5740), .ZN(n5743)
         );
  AOI21_X1 U6855 ( .B1(n5744), .B2(n6323), .A(n5743), .ZN(n5745) );
  OAI21_X1 U6856 ( .B1(n5746), .B2(n6300), .A(n5745), .ZN(U2992) );
  NAND2_X1 U6857 ( .A1(n5747), .A2(n5750), .ZN(n5748) );
  OAI211_X1 U6858 ( .C1(n5751), .C2(n5750), .A(n5749), .B(n5748), .ZN(n5752)
         );
  AOI21_X1 U6859 ( .B1(n5753), .B2(n6323), .A(n5752), .ZN(n5754) );
  OAI21_X1 U6860 ( .B1(n5755), .B2(n6300), .A(n5754), .ZN(U2993) );
  INV_X1 U6861 ( .A(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5759) );
  NAND2_X1 U6862 ( .A1(n5756), .A2(n5759), .ZN(n5757) );
  OAI211_X1 U6863 ( .C1(n5767), .C2(n5759), .A(n5758), .B(n5757), .ZN(n5760)
         );
  AOI21_X1 U6864 ( .B1(n5761), .B2(n6323), .A(n5760), .ZN(n5762) );
  OAI21_X1 U6865 ( .B1(n5763), .B2(n6300), .A(n5762), .ZN(U2995) );
  NAND2_X1 U6866 ( .A1(n5764), .A2(n6340), .ZN(n5772) );
  INV_X1 U6867 ( .A(n5765), .ZN(n5770) );
  INV_X1 U6868 ( .A(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5766) );
  NOR2_X1 U6869 ( .A1(n5767), .A2(n5766), .ZN(n5768) );
  AOI211_X1 U6870 ( .C1(n5770), .C2(INSTADDRPOINTER_REG_21__SCAN_IN), .A(n5769), .B(n5768), .ZN(n5771) );
  OAI211_X1 U6871 ( .C1(n6337), .C2(n5858), .A(n5772), .B(n5771), .ZN(U2996)
         );
  NAND2_X1 U6872 ( .A1(n5773), .A2(n6340), .ZN(n5780) );
  OAI21_X1 U6873 ( .B1(n5775), .B2(n5777), .A(n5774), .ZN(n5776) );
  AOI21_X1 U6874 ( .B1(n5778), .B2(n5777), .A(n5776), .ZN(n5779) );
  OAI211_X1 U6875 ( .C1(n6337), .C2(n5781), .A(n5780), .B(n5779), .ZN(U2997)
         );
  NAND2_X1 U6876 ( .A1(n5816), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5806) );
  NAND2_X1 U6877 ( .A1(n6334), .A2(n5806), .ZN(n5782) );
  AND2_X1 U6878 ( .A1(n5783), .A2(n5782), .ZN(n5821) );
  AOI22_X1 U6879 ( .A1(n6297), .A2(n5786), .B1(n5820), .B2(n5784), .ZN(n5785)
         );
  AND2_X1 U6880 ( .A1(n5821), .A2(n5785), .ZN(n5800) );
  NOR2_X1 U6881 ( .A1(n5806), .A2(n5786), .ZN(n5796) );
  XNOR2_X1 U6882 ( .A(n5799), .B(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5787)
         );
  NAND3_X1 U6883 ( .A1(n5817), .A2(n5796), .A3(n5787), .ZN(n5788) );
  OAI211_X1 U6884 ( .C1(n5800), .C2(n5790), .A(n5789), .B(n5788), .ZN(n5791)
         );
  AOI21_X1 U6885 ( .B1(n5863), .B2(n6323), .A(n5791), .ZN(n5792) );
  OAI21_X1 U6886 ( .B1(n5793), .B2(n6300), .A(n5792), .ZN(U2998) );
  INV_X1 U6887 ( .A(n5794), .ZN(n5804) );
  INV_X1 U6888 ( .A(n5876), .ZN(n5802) );
  INV_X1 U6889 ( .A(n5795), .ZN(n5798) );
  NAND3_X1 U6890 ( .A1(n5817), .A2(n5796), .A3(n5799), .ZN(n5797) );
  OAI211_X1 U6891 ( .C1(n5800), .C2(n5799), .A(n5798), .B(n5797), .ZN(n5801)
         );
  AOI21_X1 U6892 ( .B1(n5802), .B2(n6323), .A(n5801), .ZN(n5803) );
  OAI21_X1 U6893 ( .B1(n5804), .B2(n6300), .A(n5803), .ZN(U2999) );
  OAI21_X1 U6894 ( .B1(INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n5805), .A(n5821), 
        .ZN(n5810) );
  INV_X1 U6895 ( .A(n5817), .ZN(n5807) );
  NOR3_X1 U6896 ( .A1(n5807), .A2(INSTADDRPOINTER_REG_18__SCAN_IN), .A3(n5806), 
        .ZN(n5808) );
  AOI211_X1 U6897 ( .C1(INSTADDRPOINTER_REG_18__SCAN_IN), .C2(n5810), .A(n5809), .B(n5808), .ZN(n5813) );
  NAND2_X1 U6898 ( .A1(n5811), .A2(n6323), .ZN(n5812) );
  OAI211_X1 U6899 ( .C1(n5814), .C2(n6300), .A(n5813), .B(n5812), .ZN(U3000)
         );
  INV_X1 U6900 ( .A(n5815), .ZN(n5825) );
  NAND3_X1 U6901 ( .A1(n5817), .A2(n5816), .A3(n5820), .ZN(n5819) );
  OAI211_X1 U6902 ( .C1(n5821), .C2(n5820), .A(n5819), .B(n5818), .ZN(n5822)
         );
  AOI21_X1 U6903 ( .B1(n5823), .B2(n6323), .A(n5822), .ZN(n5824) );
  OAI21_X1 U6904 ( .B1(n5825), .B2(n6300), .A(n5824), .ZN(U3001) );
  OAI211_X1 U6905 ( .C1(STATEBS16_REG_SCAN_IN), .C2(n5827), .A(n5832), .B(
        n5826), .ZN(n5828) );
  OAI21_X1 U6906 ( .B1(n5834), .B2(n5829), .A(n5828), .ZN(n5830) );
  MUX2_X1 U6907 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(n5830), .S(n6345), 
        .Z(U3464) );
  XNOR2_X1 U6908 ( .A(n5832), .B(n5831), .ZN(n5836) );
  INV_X1 U6909 ( .A(n5833), .ZN(n6062) );
  OAI22_X1 U6910 ( .A1(n5836), .A2(n5835), .B1(n6062), .B2(n5834), .ZN(n5837)
         );
  MUX2_X1 U6911 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B(n5837), .S(n6345), 
        .Z(U3463) );
  NOR2_X1 U6912 ( .A1(n5839), .A2(n5838), .ZN(n5845) );
  INV_X1 U6913 ( .A(n5840), .ZN(n6585) );
  OAI21_X1 U6914 ( .B1(n5845), .B2(n5842), .A(n5841), .ZN(n5843) );
  AOI21_X1 U6915 ( .B1(n6074), .B2(n5844), .A(n5843), .ZN(n6460) );
  OAI222_X1 U6916 ( .A1(n5847), .A2(n5846), .B1(n6583), .B2(n5845), .C1(n6585), 
        .C2(n6460), .ZN(n5848) );
  MUX2_X1 U6917 ( .A(n5848), .B(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .S(n5917), 
        .Z(U3460) );
  AND2_X1 U6918 ( .A1(n6118), .A2(DATAO_REG_31__SCAN_IN), .ZN(U2892) );
  AOI21_X1 U6919 ( .B1(n5860), .B2(n5849), .A(n6560), .ZN(n5853) );
  INV_X1 U6920 ( .A(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n5850) );
  OAI22_X1 U6921 ( .A1(REIP_REG_22__SCAN_IN), .A2(n5851), .B1(n5850), .B2(
        n6078), .ZN(n5852) );
  AOI211_X1 U6922 ( .C1(n6072), .C2(EBX_REG_22__SCAN_IN), .A(n5853), .B(n5852), 
        .ZN(n5857) );
  OAI22_X1 U6923 ( .A1(n5877), .A2(n5971), .B1(n5854), .B2(n6071), .ZN(n5855)
         );
  INV_X1 U6924 ( .A(n5855), .ZN(n5856) );
  OAI211_X1 U6925 ( .C1(n5858), .C2(n6087), .A(n5857), .B(n5856), .ZN(U2805)
         );
  AOI21_X1 U6926 ( .B1(n6083), .B2(n5859), .A(REIP_REG_20__SCAN_IN), .ZN(n5861) );
  OAI22_X1 U6927 ( .A1(n5861), .A2(n5860), .B1(n3827), .B2(n6078), .ZN(n5862)
         );
  AOI21_X1 U6928 ( .B1(EBX_REG_20__SCAN_IN), .B2(n6072), .A(n5862), .ZN(n5865)
         );
  AOI22_X1 U6929 ( .A1(n5885), .A2(n6036), .B1(n5863), .B2(n6047), .ZN(n5864)
         );
  OAI211_X1 U6930 ( .C1(n5866), .C2(n6071), .A(n5865), .B(n5864), .ZN(U2807)
         );
  NOR3_X1 U6931 ( .A1(n6065), .A2(REIP_REG_19__SCAN_IN), .A3(n5867), .ZN(n5871) );
  NOR2_X1 U6932 ( .A1(n6065), .A2(REIP_REG_18__SCAN_IN), .ZN(n5943) );
  OAI21_X1 U6933 ( .B1(n5945), .B2(n5943), .A(REIP_REG_19__SCAN_IN), .ZN(n5868) );
  OAI211_X1 U6934 ( .C1(n6078), .C2(n5869), .A(n5868), .B(n6335), .ZN(n5870)
         );
  AOI211_X1 U6935 ( .C1(n6072), .C2(EBX_REG_19__SCAN_IN), .A(n5871), .B(n5870), 
        .ZN(n5875) );
  INV_X1 U6936 ( .A(n5872), .ZN(n5888) );
  AOI22_X1 U6937 ( .A1(n5888), .A2(n6036), .B1(n5873), .B2(n5194), .ZN(n5874)
         );
  OAI211_X1 U6938 ( .C1(n5876), .C2(n6087), .A(n5875), .B(n5874), .ZN(U2808)
         );
  INV_X1 U6939 ( .A(n5877), .ZN(n5879) );
  INV_X1 U6940 ( .A(n5878), .ZN(n6100) );
  AOI22_X1 U6941 ( .A1(n5879), .A2(n6100), .B1(n6099), .B2(DATAI_22_), .ZN(
        n5881) );
  AOI22_X1 U6942 ( .A1(n6103), .A2(DATAI_6_), .B1(n6102), .B2(
        EAX_REG_22__SCAN_IN), .ZN(n5880) );
  NAND2_X1 U6943 ( .A1(n5881), .A2(n5880), .ZN(U2869) );
  AOI22_X1 U6944 ( .A1(n5882), .A2(n6100), .B1(n6099), .B2(DATAI_21_), .ZN(
        n5884) );
  AOI22_X1 U6945 ( .A1(n6103), .A2(DATAI_5_), .B1(n6102), .B2(
        EAX_REG_21__SCAN_IN), .ZN(n5883) );
  NAND2_X1 U6946 ( .A1(n5884), .A2(n5883), .ZN(U2870) );
  AOI22_X1 U6947 ( .A1(n5885), .A2(n6100), .B1(n6099), .B2(DATAI_20_), .ZN(
        n5887) );
  AOI22_X1 U6948 ( .A1(n6103), .A2(DATAI_4_), .B1(n6102), .B2(
        EAX_REG_20__SCAN_IN), .ZN(n5886) );
  NAND2_X1 U6949 ( .A1(n5887), .A2(n5886), .ZN(U2871) );
  AOI22_X1 U6950 ( .A1(n5888), .A2(n6100), .B1(n6099), .B2(DATAI_19_), .ZN(
        n5890) );
  AOI22_X1 U6951 ( .A1(n6103), .A2(DATAI_3_), .B1(n6102), .B2(
        EAX_REG_19__SCAN_IN), .ZN(n5889) );
  NAND2_X1 U6952 ( .A1(n5890), .A2(n5889), .ZN(U2872) );
  AOI22_X1 U6953 ( .A1(n2993), .A2(REIP_REG_13__SCAN_IN), .B1(n6239), .B2(
        PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n5895) );
  NAND2_X1 U6954 ( .A1(n5319), .A2(n5891), .ZN(n5893) );
  XNOR2_X1 U6955 ( .A(n5893), .B(n5892), .ZN(n5906) );
  AOI22_X1 U6956 ( .A1(n5906), .A2(n6243), .B1(n6244), .B2(n6089), .ZN(n5894)
         );
  OAI211_X1 U6957 ( .C1(n6249), .C2(n5995), .A(n5895), .B(n5894), .ZN(U2973)
         );
  INV_X1 U6958 ( .A(n5896), .ZN(n5901) );
  INV_X1 U6959 ( .A(n5897), .ZN(n5899) );
  AOI222_X1 U6960 ( .A1(n5899), .A2(n6340), .B1(n6323), .B2(n5898), .C1(
        REIP_REG_15__SCAN_IN), .C2(n2993), .ZN(n5900) );
  OAI221_X1 U6961 ( .B1(INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n5902), .C1(
        n5675), .C2(n5901), .A(n5900), .ZN(U3003) );
  OR2_X1 U6962 ( .A1(n5217), .A2(n5903), .ZN(n5904) );
  AND2_X1 U6963 ( .A1(n5905), .A2(n5904), .ZN(n6088) );
  AOI22_X1 U6964 ( .A1(n5906), .A2(n6340), .B1(n6323), .B2(n6088), .ZN(n5916)
         );
  NAND2_X1 U6965 ( .A1(n2993), .A2(REIP_REG_13__SCAN_IN), .ZN(n5915) );
  OAI21_X1 U6966 ( .B1(INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n5908), .A(n5907), 
        .ZN(n5914) );
  INV_X1 U6967 ( .A(n5909), .ZN(n5912) );
  NAND3_X1 U6968 ( .A1(n5912), .A2(n5911), .A3(n5910), .ZN(n5913) );
  NAND4_X1 U6969 ( .A1(n5916), .A2(n5915), .A3(n5914), .A4(n5913), .ZN(U3005)
         );
  INV_X1 U6970 ( .A(n5917), .ZN(n6587) );
  INV_X1 U6971 ( .A(n5918), .ZN(n5920) );
  NAND3_X1 U6972 ( .A1(n5920), .A2(n6581), .A3(n5919), .ZN(n5921) );
  OAI21_X1 U6973 ( .B1(n6587), .B2(n3582), .A(n5921), .ZN(U3455) );
  INV_X1 U6974 ( .A(ADS_N_REG_SCAN_IN), .ZN(n6751) );
  INV_X1 U6975 ( .A(STATE_REG_0__SCAN_IN), .ZN(n6522) );
  INV_X1 U6976 ( .A(STATE_REG_1__SCAN_IN), .ZN(n5922) );
  NAND2_X1 U6977 ( .A1(n6522), .A2(STATE_REG_1__SCAN_IN), .ZN(n6565) );
  AOI221_X1 U6978 ( .B1(STATE_REG_2__SCAN_IN), .B2(STATE_REG_0__SCAN_IN), .C1(
        n5922), .C2(STATE_REG_0__SCAN_IN), .A(n6804), .ZN(n6578) );
  OAI21_X1 U6979 ( .B1(n6751), .B2(n6522), .A(n6511), .ZN(U2789) );
  OAI21_X1 U6980 ( .B1(n5923), .B2(n6500), .A(CODEFETCH_REG_SCAN_IN), .ZN(
        n5924) );
  OAI21_X1 U6981 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n6501), .A(n5924), .ZN(
        U2790) );
  INV_X1 U6982 ( .A(D_C_N_REG_SCAN_IN), .ZN(n6671) );
  NOR2_X1 U6983 ( .A1(STATE_REG_0__SCAN_IN), .A2(STATE_REG_2__SCAN_IN), .ZN(
        n5926) );
  NOR2_X1 U6984 ( .A1(n6804), .A2(n5926), .ZN(n5925) );
  AOI22_X1 U6985 ( .A1(CODEFETCH_REG_SCAN_IN), .A2(n6804), .B1(n6671), .B2(
        n5925), .ZN(U2791) );
  OAI21_X1 U6986 ( .B1(BS16_N), .B2(n5926), .A(n6578), .ZN(n6576) );
  OAI21_X1 U6987 ( .B1(n6578), .B2(n6657), .A(n6576), .ZN(U2792) );
  INV_X1 U6988 ( .A(n5927), .ZN(n5928) );
  OAI21_X1 U6989 ( .B1(n5928), .B2(n6696), .A(n6221), .ZN(U2793) );
  NOR4_X1 U6990 ( .A1(DATAWIDTH_REG_20__SCAN_IN), .A2(
        DATAWIDTH_REG_21__SCAN_IN), .A3(DATAWIDTH_REG_22__SCAN_IN), .A4(
        DATAWIDTH_REG_23__SCAN_IN), .ZN(n5932) );
  NOR4_X1 U6991 ( .A1(DATAWIDTH_REG_16__SCAN_IN), .A2(
        DATAWIDTH_REG_17__SCAN_IN), .A3(DATAWIDTH_REG_18__SCAN_IN), .A4(
        DATAWIDTH_REG_19__SCAN_IN), .ZN(n5931) );
  NOR4_X1 U6992 ( .A1(DATAWIDTH_REG_28__SCAN_IN), .A2(
        DATAWIDTH_REG_29__SCAN_IN), .A3(DATAWIDTH_REG_30__SCAN_IN), .A4(
        DATAWIDTH_REG_31__SCAN_IN), .ZN(n5930) );
  NOR4_X1 U6993 ( .A1(DATAWIDTH_REG_24__SCAN_IN), .A2(
        DATAWIDTH_REG_25__SCAN_IN), .A3(DATAWIDTH_REG_26__SCAN_IN), .A4(
        DATAWIDTH_REG_27__SCAN_IN), .ZN(n5929) );
  NAND4_X1 U6994 ( .A1(n5932), .A2(n5931), .A3(n5930), .A4(n5929), .ZN(n5938)
         );
  NOR4_X1 U6995 ( .A1(DATAWIDTH_REG_4__SCAN_IN), .A2(DATAWIDTH_REG_5__SCAN_IN), 
        .A3(DATAWIDTH_REG_6__SCAN_IN), .A4(DATAWIDTH_REG_7__SCAN_IN), .ZN(
        n5936) );
  AOI211_X1 U6996 ( .C1(DATAWIDTH_REG_0__SCAN_IN), .C2(
        DATAWIDTH_REG_1__SCAN_IN), .A(DATAWIDTH_REG_2__SCAN_IN), .B(
        DATAWIDTH_REG_3__SCAN_IN), .ZN(n5935) );
  NOR4_X1 U6997 ( .A1(DATAWIDTH_REG_12__SCAN_IN), .A2(
        DATAWIDTH_REG_13__SCAN_IN), .A3(DATAWIDTH_REG_14__SCAN_IN), .A4(
        DATAWIDTH_REG_15__SCAN_IN), .ZN(n5934) );
  NOR4_X1 U6998 ( .A1(DATAWIDTH_REG_8__SCAN_IN), .A2(DATAWIDTH_REG_9__SCAN_IN), 
        .A3(DATAWIDTH_REG_10__SCAN_IN), .A4(DATAWIDTH_REG_11__SCAN_IN), .ZN(
        n5933) );
  NAND4_X1 U6999 ( .A1(n5936), .A2(n5935), .A3(n5934), .A4(n5933), .ZN(n5937)
         );
  NOR2_X1 U7000 ( .A1(n5938), .A2(n5937), .ZN(n6593) );
  INV_X1 U7001 ( .A(BYTEENABLE_REG_1__SCAN_IN), .ZN(n6748) );
  NOR3_X1 U7002 ( .A1(REIP_REG_0__SCAN_IN), .A2(DATAWIDTH_REG_1__SCAN_IN), 
        .A3(DATAWIDTH_REG_0__SCAN_IN), .ZN(n5940) );
  OAI21_X1 U7003 ( .B1(REIP_REG_1__SCAN_IN), .B2(n5940), .A(n6593), .ZN(n5939)
         );
  OAI21_X1 U7004 ( .B1(n6593), .B2(n6748), .A(n5939), .ZN(U2794) );
  INV_X1 U7005 ( .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6577) );
  AOI21_X1 U7006 ( .B1(n6531), .B2(n6577), .A(n5940), .ZN(n5942) );
  INV_X1 U7007 ( .A(BYTEENABLE_REG_3__SCAN_IN), .ZN(n5941) );
  INV_X1 U7008 ( .A(n6593), .ZN(n6591) );
  AOI22_X1 U7009 ( .A1(n6593), .A2(n5942), .B1(n5941), .B2(n6591), .ZN(U2795)
         );
  AOI22_X1 U7010 ( .A1(REIP_REG_18__SCAN_IN), .A2(n5945), .B1(n5944), .B2(
        n5943), .ZN(n5946) );
  OAI211_X1 U7011 ( .C1(n6078), .C2(n3789), .A(n5946), .B(n6335), .ZN(n5950)
         );
  OAI22_X1 U7012 ( .A1(n5948), .A2(n5971), .B1(n6087), .B2(n5947), .ZN(n5949)
         );
  AOI211_X1 U7013 ( .C1(EBX_REG_18__SCAN_IN), .C2(n6072), .A(n5950), .B(n5949), 
        .ZN(n5951) );
  OAI21_X1 U7014 ( .B1(n5952), .B2(n6071), .A(n5951), .ZN(U2809) );
  NOR3_X1 U7015 ( .A1(n6065), .A2(REIP_REG_15__SCAN_IN), .A3(n5953), .ZN(n5968) );
  INV_X1 U7016 ( .A(n5953), .ZN(n5954) );
  NAND2_X1 U7017 ( .A1(n6046), .A2(n5954), .ZN(n5955) );
  AND2_X1 U7018 ( .A1(n6067), .A2(n5955), .ZN(n5977) );
  OAI21_X1 U7019 ( .B1(n5968), .B2(n5977), .A(REIP_REG_16__SCAN_IN), .ZN(n5959) );
  INV_X1 U7020 ( .A(REIP_REG_16__SCAN_IN), .ZN(n5957) );
  NAND3_X1 U7021 ( .A1(n6083), .A2(n5957), .A3(n5956), .ZN(n5958) );
  OAI211_X1 U7022 ( .C1(n6030), .C2(n5960), .A(n5959), .B(n5958), .ZN(n5961)
         );
  AOI211_X1 U7023 ( .C1(n6059), .C2(PHYADDRPOINTER_REG_16__SCAN_IN), .A(n2993), 
        .B(n5961), .ZN(n5964) );
  AOI22_X1 U7024 ( .A1(n6101), .A2(n6036), .B1(n5194), .B2(n5962), .ZN(n5963)
         );
  OAI211_X1 U7025 ( .C1(n6087), .C2(n5965), .A(n5964), .B(n5963), .ZN(U2811)
         );
  NAND2_X1 U7026 ( .A1(n6072), .A2(EBX_REG_15__SCAN_IN), .ZN(n5966) );
  OAI211_X1 U7027 ( .C1(n6078), .C2(n5967), .A(n5966), .B(n6335), .ZN(n5969)
         );
  AOI211_X1 U7028 ( .C1(n5977), .C2(REIP_REG_15__SCAN_IN), .A(n5969), .B(n5968), .ZN(n5970) );
  OAI21_X1 U7029 ( .B1(n5972), .B2(n5971), .A(n5970), .ZN(n5973) );
  AOI21_X1 U7030 ( .B1(n5974), .B2(n5194), .A(n5973), .ZN(n5975) );
  OAI21_X1 U7031 ( .B1(n6087), .B2(n5976), .A(n5975), .ZN(U2812) );
  INV_X1 U7032 ( .A(n5977), .ZN(n5981) );
  AOI21_X1 U7033 ( .B1(n6083), .B2(n5978), .A(REIP_REG_14__SCAN_IN), .ZN(n5980) );
  OAI22_X1 U7034 ( .A1(n5981), .A2(n5980), .B1(n5979), .B2(n6030), .ZN(n5982)
         );
  AOI211_X1 U7035 ( .C1(n6059), .C2(PHYADDRPOINTER_REG_14__SCAN_IN), .A(n2993), 
        .B(n5982), .ZN(n5986) );
  AOI22_X1 U7036 ( .A1(n5984), .A2(n6036), .B1(n5194), .B2(n5983), .ZN(n5985)
         );
  OAI211_X1 U7037 ( .C1(n6087), .C2(n5987), .A(n5986), .B(n5985), .ZN(U2813)
         );
  NOR4_X1 U7038 ( .A1(n6065), .A2(n5988), .A3(n6547), .A4(REIP_REG_13__SCAN_IN), .ZN(n5992) );
  OAI21_X1 U7039 ( .B1(n5989), .B2(n6004), .A(REIP_REG_13__SCAN_IN), .ZN(n5990) );
  OAI211_X1 U7040 ( .C1(n6078), .C2(n3693), .A(n6335), .B(n5990), .ZN(n5991)
         );
  AOI211_X1 U7041 ( .C1(n6072), .C2(EBX_REG_13__SCAN_IN), .A(n5992), .B(n5991), 
        .ZN(n5994) );
  AOI22_X1 U7042 ( .A1(n6089), .A2(n6036), .B1(n6047), .B2(n6088), .ZN(n5993)
         );
  OAI211_X1 U7043 ( .C1(n5995), .C2(n6071), .A(n5994), .B(n5993), .ZN(U2814)
         );
  AND2_X1 U7044 ( .A1(n5997), .A2(n5996), .ZN(n5998) );
  NOR2_X1 U7045 ( .A1(n5999), .A2(n5998), .ZN(n6256) );
  AOI22_X1 U7046 ( .A1(n6047), .A2(n6256), .B1(n6001), .B2(n6000), .ZN(n6007)
         );
  INV_X1 U7047 ( .A(EBX_REG_11__SCAN_IN), .ZN(n6094) );
  OAI22_X1 U7048 ( .A1(n6094), .A2(n6030), .B1(n6002), .B2(n6078), .ZN(n6003)
         );
  AOI211_X1 U7049 ( .C1(REIP_REG_11__SCAN_IN), .C2(n6004), .A(n2993), .B(n6003), .ZN(n6006) );
  AOI22_X1 U7050 ( .A1(n6218), .A2(n6036), .B1(n5194), .B2(n6216), .ZN(n6005)
         );
  NAND3_X1 U7051 ( .A1(n6007), .A2(n6006), .A3(n6005), .ZN(U2816) );
  INV_X1 U7052 ( .A(n6008), .ZN(n6014) );
  INV_X1 U7053 ( .A(n6009), .ZN(n6272) );
  AOI22_X1 U7054 ( .A1(EBX_REG_9__SCAN_IN), .A2(n6072), .B1(n6047), .B2(n6272), 
        .ZN(n6010) );
  OAI211_X1 U7055 ( .C1(n6078), .C2(n6011), .A(n6010), .B(n6335), .ZN(n6012)
         );
  AOI211_X1 U7056 ( .C1(n6014), .C2(n6036), .A(n6013), .B(n6012), .ZN(n6017)
         );
  AOI22_X1 U7057 ( .A1(n6015), .A2(n5194), .B1(REIP_REG_9__SCAN_IN), .B2(n6019), .ZN(n6016) );
  NAND2_X1 U7058 ( .A1(n6017), .A2(n6016), .ZN(U2818) );
  INV_X1 U7059 ( .A(n6018), .ZN(n6280) );
  AOI22_X1 U7060 ( .A1(n6047), .A2(n6280), .B1(REIP_REG_8__SCAN_IN), .B2(n6019), .ZN(n6029) );
  NAND2_X1 U7061 ( .A1(n6020), .A2(n6036), .ZN(n6025) );
  NAND3_X1 U7062 ( .A1(n6083), .A2(n6022), .A3(n6021), .ZN(n6024) );
  NAND2_X1 U7063 ( .A1(n6059), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n6023)
         );
  NAND4_X1 U7064 ( .A1(n6025), .A2(n6335), .A3(n6024), .A4(n6023), .ZN(n6026)
         );
  AOI21_X1 U7065 ( .B1(n6027), .B2(n5194), .A(n6026), .ZN(n6028) );
  OAI211_X1 U7066 ( .C1(n6031), .C2(n6030), .A(n6029), .B(n6028), .ZN(U2819)
         );
  AOI211_X1 U7067 ( .C1(n6059), .C2(PHYADDRPOINTER_REG_6__SCAN_IN), .A(n2993), 
        .B(n6032), .ZN(n6033) );
  OAI21_X1 U7068 ( .B1(n6087), .B2(n6301), .A(n6033), .ZN(n6034) );
  AOI21_X1 U7069 ( .B1(EBX_REG_6__SCAN_IN), .B2(n6072), .A(n6034), .ZN(n6038)
         );
  AOI22_X1 U7070 ( .A1(n6225), .A2(n6036), .B1(REIP_REG_6__SCAN_IN), .B2(n6035), .ZN(n6037) );
  OAI211_X1 U7071 ( .C1(n6229), .C2(n6071), .A(n6038), .B(n6037), .ZN(U2821)
         );
  NOR3_X1 U7072 ( .A1(n6065), .A2(n6040), .A3(REIP_REG_4__SCAN_IN), .ZN(n6039)
         );
  AOI211_X1 U7073 ( .C1(n6059), .C2(PHYADDRPOINTER_REG_4__SCAN_IN), .A(n2993), 
        .B(n6039), .ZN(n6045) );
  OAI21_X1 U7074 ( .B1(n6075), .B2(n6040), .A(n6067), .ZN(n6057) );
  OAI22_X1 U7075 ( .A1(n6057), .A2(n6536), .B1(n6041), .B2(n6061), .ZN(n6043)
         );
  OAI22_X1 U7076 ( .A1(n6234), .A2(n6058), .B1(n6238), .B2(n6071), .ZN(n6042)
         );
  AOI211_X1 U7077 ( .C1(EBX_REG_4__SCAN_IN), .C2(n6072), .A(n6043), .B(n6042), 
        .ZN(n6044) );
  OAI211_X1 U7078 ( .C1(n6087), .C2(n6313), .A(n6045), .B(n6044), .ZN(U2823)
         );
  NAND3_X1 U7079 ( .A1(REIP_REG_1__SCAN_IN), .A2(n6046), .A3(
        REIP_REG_2__SCAN_IN), .ZN(n6066) );
  NAND2_X1 U7080 ( .A1(n6047), .A2(n6322), .ZN(n6049) );
  AOI22_X1 U7081 ( .A1(n6072), .A2(EBX_REG_3__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n6059), .ZN(n6048) );
  OAI211_X1 U7082 ( .C1(n6050), .C2(n6061), .A(n6049), .B(n6048), .ZN(n6051)
         );
  INV_X1 U7083 ( .A(n6051), .ZN(n6052) );
  OAI21_X1 U7084 ( .B1(n6053), .B2(n6058), .A(n6052), .ZN(n6054) );
  AOI21_X1 U7085 ( .B1(n6055), .B2(n5194), .A(n6054), .ZN(n6056) );
  OAI221_X1 U7086 ( .B1(n6057), .B2(n4543), .C1(n6057), .C2(n6066), .A(n6056), 
        .ZN(U2824) );
  INV_X1 U7087 ( .A(n6058), .ZN(n6081) );
  NOR2_X1 U7088 ( .A1(n6087), .A2(n6336), .ZN(n6064) );
  AOI22_X1 U7089 ( .A1(n6072), .A2(EBX_REG_2__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n6059), .ZN(n6060) );
  OAI21_X1 U7090 ( .B1(n6062), .B2(n6061), .A(n6060), .ZN(n6063) );
  AOI211_X1 U7091 ( .C1(n6245), .C2(n6081), .A(n6064), .B(n6063), .ZN(n6070)
         );
  NOR2_X1 U7092 ( .A1(n6065), .A2(n6531), .ZN(n6068) );
  OAI211_X1 U7093 ( .C1(n6068), .C2(REIP_REG_2__SCAN_IN), .A(n6067), .B(n6066), 
        .ZN(n6069) );
  OAI211_X1 U7094 ( .C1(n6071), .C2(n6248), .A(n6070), .B(n6069), .ZN(U2825)
         );
  INV_X1 U7095 ( .A(PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n6079) );
  AOI22_X1 U7096 ( .A1(n6074), .A2(n6073), .B1(n6072), .B2(EBX_REG_1__SCAN_IN), 
        .ZN(n6077) );
  AOI22_X1 U7097 ( .A1(n5194), .A2(n6079), .B1(n6075), .B2(REIP_REG_1__SCAN_IN), .ZN(n6076) );
  OAI211_X1 U7098 ( .C1(n6079), .C2(n6078), .A(n6077), .B(n6076), .ZN(n6080)
         );
  AOI21_X1 U7099 ( .B1(n6082), .B2(n6081), .A(n6080), .ZN(n6085) );
  NAND2_X1 U7100 ( .A1(n6083), .A2(n6531), .ZN(n6084) );
  OAI211_X1 U7101 ( .C1(n6087), .C2(n6086), .A(n6085), .B(n6084), .ZN(U2826)
         );
  INV_X1 U7102 ( .A(EBX_REG_13__SCAN_IN), .ZN(n6091) );
  AOI22_X1 U7103 ( .A1(n6089), .A2(n4149), .B1(n6092), .B2(n6088), .ZN(n6090)
         );
  OAI21_X1 U7104 ( .B1(n6095), .B2(n6091), .A(n6090), .ZN(U2846) );
  AOI22_X1 U7105 ( .A1(n6218), .A2(n4149), .B1(n6092), .B2(n6256), .ZN(n6093)
         );
  OAI21_X1 U7106 ( .B1(n6095), .B2(n6094), .A(n6093), .ZN(U2848) );
  AOI22_X1 U7107 ( .A1(n6096), .A2(n6100), .B1(n6099), .B2(DATAI_18_), .ZN(
        n6098) );
  AOI22_X1 U7108 ( .A1(n6103), .A2(DATAI_2_), .B1(n6102), .B2(
        EAX_REG_18__SCAN_IN), .ZN(n6097) );
  NAND2_X1 U7109 ( .A1(n6098), .A2(n6097), .ZN(U2873) );
  AOI22_X1 U7110 ( .A1(n6101), .A2(n6100), .B1(n6099), .B2(DATAI_16_), .ZN(
        n6105) );
  AOI22_X1 U7111 ( .A1(n6103), .A2(DATAI_0_), .B1(n6102), .B2(
        EAX_REG_16__SCAN_IN), .ZN(n6104) );
  NAND2_X1 U7112 ( .A1(n6105), .A2(n6104), .ZN(U2875) );
  AOI22_X1 U7113 ( .A1(n6597), .A2(LWORD_REG_15__SCAN_IN), .B1(n6118), .B2(
        DATAO_REG_15__SCAN_IN), .ZN(n6106) );
  OAI21_X1 U7114 ( .B1(n6211), .B2(n6125), .A(n6106), .ZN(U2908) );
  AOI22_X1 U7115 ( .A1(n6597), .A2(LWORD_REG_14__SCAN_IN), .B1(n6118), .B2(
        DATAO_REG_14__SCAN_IN), .ZN(n6107) );
  OAI21_X1 U7116 ( .B1(n6206), .B2(n6125), .A(n6107), .ZN(U2909) );
  AOI22_X1 U7117 ( .A1(n6597), .A2(LWORD_REG_13__SCAN_IN), .B1(n6118), .B2(
        DATAO_REG_13__SCAN_IN), .ZN(n6108) );
  OAI21_X1 U7118 ( .B1(n6203), .B2(n6125), .A(n6108), .ZN(U2910) );
  AOI22_X1 U7119 ( .A1(n6112), .A2(LWORD_REG_12__SCAN_IN), .B1(n6118), .B2(
        DATAO_REG_12__SCAN_IN), .ZN(n6109) );
  OAI21_X1 U7120 ( .B1(n6199), .B2(n6125), .A(n6109), .ZN(U2911) );
  AOI22_X1 U7121 ( .A1(n6112), .A2(LWORD_REG_11__SCAN_IN), .B1(n6118), .B2(
        DATAO_REG_11__SCAN_IN), .ZN(n6110) );
  OAI21_X1 U7122 ( .B1(n6196), .B2(n6125), .A(n6110), .ZN(U2912) );
  AOI22_X1 U7123 ( .A1(n6112), .A2(LWORD_REG_10__SCAN_IN), .B1(n6118), .B2(
        DATAO_REG_10__SCAN_IN), .ZN(n6111) );
  OAI21_X1 U7124 ( .B1(n6193), .B2(n6125), .A(n6111), .ZN(U2913) );
  AOI22_X1 U7125 ( .A1(n6112), .A2(LWORD_REG_9__SCAN_IN), .B1(n6118), .B2(
        DATAO_REG_9__SCAN_IN), .ZN(n6113) );
  OAI21_X1 U7126 ( .B1(n6190), .B2(n6125), .A(n6113), .ZN(U2914) );
  AOI22_X1 U7127 ( .A1(n6597), .A2(LWORD_REG_8__SCAN_IN), .B1(n6118), .B2(
        DATAO_REG_8__SCAN_IN), .ZN(n6114) );
  OAI21_X1 U7128 ( .B1(n6187), .B2(n6125), .A(n6114), .ZN(U2915) );
  AOI22_X1 U7129 ( .A1(n6597), .A2(LWORD_REG_7__SCAN_IN), .B1(n6118), .B2(
        DATAO_REG_7__SCAN_IN), .ZN(n6115) );
  OAI21_X1 U7130 ( .B1(n6184), .B2(n6125), .A(n6115), .ZN(U2916) );
  AOI22_X1 U7131 ( .A1(n6597), .A2(LWORD_REG_6__SCAN_IN), .B1(n6118), .B2(
        DATAO_REG_6__SCAN_IN), .ZN(n6116) );
  OAI21_X1 U7132 ( .B1(n6181), .B2(n6125), .A(n6116), .ZN(U2917) );
  AOI22_X1 U7133 ( .A1(n6597), .A2(LWORD_REG_5__SCAN_IN), .B1(n6118), .B2(
        DATAO_REG_5__SCAN_IN), .ZN(n6117) );
  OAI21_X1 U7134 ( .B1(n6178), .B2(n6125), .A(n6117), .ZN(U2918) );
  AOI22_X1 U7135 ( .A1(n6597), .A2(LWORD_REG_4__SCAN_IN), .B1(n6118), .B2(
        DATAO_REG_4__SCAN_IN), .ZN(n6119) );
  OAI21_X1 U7136 ( .B1(n6175), .B2(n6125), .A(n6119), .ZN(U2919) );
  AOI22_X1 U7137 ( .A1(n6597), .A2(LWORD_REG_3__SCAN_IN), .B1(n6123), .B2(
        DATAO_REG_3__SCAN_IN), .ZN(n6120) );
  OAI21_X1 U7138 ( .B1(n6172), .B2(n6125), .A(n6120), .ZN(U2920) );
  AOI22_X1 U7139 ( .A1(n6597), .A2(LWORD_REG_2__SCAN_IN), .B1(n6123), .B2(
        DATAO_REG_2__SCAN_IN), .ZN(n6121) );
  OAI21_X1 U7140 ( .B1(n6169), .B2(n6125), .A(n6121), .ZN(U2921) );
  AOI22_X1 U7141 ( .A1(n6597), .A2(LWORD_REG_1__SCAN_IN), .B1(n6123), .B2(
        DATAO_REG_1__SCAN_IN), .ZN(n6122) );
  OAI21_X1 U7142 ( .B1(n6166), .B2(n6125), .A(n6122), .ZN(U2922) );
  AOI22_X1 U7143 ( .A1(n6597), .A2(LWORD_REG_0__SCAN_IN), .B1(n6123), .B2(
        DATAO_REG_0__SCAN_IN), .ZN(n6124) );
  OAI21_X1 U7144 ( .B1(n6163), .B2(n6125), .A(n6124), .ZN(U2923) );
  INV_X1 U7145 ( .A(n6126), .ZN(n6128) );
  INV_X1 U7146 ( .A(n6490), .ZN(n6127) );
  NAND2_X2 U7147 ( .A1(n6128), .A2(n6127), .ZN(n6210) );
  OAI21_X1 U7148 ( .B1(n6487), .B2(n6130), .A(n6129), .ZN(n6208) );
  AND2_X1 U7149 ( .A1(n6207), .A2(DATAI_0_), .ZN(n6161) );
  AOI21_X1 U7150 ( .B1(UWORD_REG_0__SCAN_IN), .B2(n6208), .A(n6161), .ZN(n6132) );
  OAI21_X1 U7151 ( .B1(n3755), .B2(n6210), .A(n6132), .ZN(U2924) );
  AND2_X1 U7152 ( .A1(n6207), .A2(DATAI_1_), .ZN(n6164) );
  AOI21_X1 U7153 ( .B1(UWORD_REG_1__SCAN_IN), .B2(n6208), .A(n6164), .ZN(n6133) );
  OAI21_X1 U7154 ( .B1(n6134), .B2(n6210), .A(n6133), .ZN(U2925) );
  AND2_X1 U7155 ( .A1(n6207), .A2(DATAI_2_), .ZN(n6167) );
  AOI21_X1 U7156 ( .B1(UWORD_REG_2__SCAN_IN), .B2(n6208), .A(n6167), .ZN(n6135) );
  OAI21_X1 U7157 ( .B1(n6136), .B2(n6210), .A(n6135), .ZN(U2926) );
  AND2_X1 U7158 ( .A1(n6207), .A2(DATAI_3_), .ZN(n6170) );
  AOI21_X1 U7159 ( .B1(UWORD_REG_3__SCAN_IN), .B2(n6201), .A(n6170), .ZN(n6137) );
  OAI21_X1 U7160 ( .B1(n6138), .B2(n6210), .A(n6137), .ZN(U2927) );
  AND2_X1 U7161 ( .A1(n6207), .A2(DATAI_4_), .ZN(n6173) );
  AOI21_X1 U7162 ( .B1(UWORD_REG_4__SCAN_IN), .B2(n6201), .A(n6173), .ZN(n6139) );
  OAI21_X1 U7163 ( .B1(n6140), .B2(n6210), .A(n6139), .ZN(U2928) );
  AND2_X1 U7164 ( .A1(n6207), .A2(DATAI_5_), .ZN(n6176) );
  AOI21_X1 U7165 ( .B1(UWORD_REG_5__SCAN_IN), .B2(n6201), .A(n6176), .ZN(n6141) );
  OAI21_X1 U7166 ( .B1(n6142), .B2(n6210), .A(n6141), .ZN(U2929) );
  AND2_X1 U7167 ( .A1(n6207), .A2(DATAI_6_), .ZN(n6179) );
  AOI21_X1 U7168 ( .B1(UWORD_REG_6__SCAN_IN), .B2(n6201), .A(n6179), .ZN(n6143) );
  OAI21_X1 U7169 ( .B1(n6144), .B2(n6210), .A(n6143), .ZN(U2930) );
  AND2_X1 U7170 ( .A1(n6207), .A2(DATAI_7_), .ZN(n6182) );
  AOI21_X1 U7171 ( .B1(UWORD_REG_7__SCAN_IN), .B2(n6201), .A(n6182), .ZN(n6145) );
  OAI21_X1 U7172 ( .B1(n6146), .B2(n6210), .A(n6145), .ZN(U2931) );
  AND2_X1 U7173 ( .A1(n6207), .A2(DATAI_8_), .ZN(n6185) );
  AOI21_X1 U7174 ( .B1(UWORD_REG_8__SCAN_IN), .B2(n6201), .A(n6185), .ZN(n6147) );
  OAI21_X1 U7175 ( .B1(n6148), .B2(n6210), .A(n6147), .ZN(U2932) );
  AND2_X1 U7176 ( .A1(n6207), .A2(DATAI_9_), .ZN(n6188) );
  AOI21_X1 U7177 ( .B1(UWORD_REG_9__SCAN_IN), .B2(n6201), .A(n6188), .ZN(n6149) );
  OAI21_X1 U7178 ( .B1(n6150), .B2(n6210), .A(n6149), .ZN(U2933) );
  AND2_X1 U7179 ( .A1(n6207), .A2(DATAI_10_), .ZN(n6191) );
  AOI21_X1 U7180 ( .B1(UWORD_REG_10__SCAN_IN), .B2(n6201), .A(n6191), .ZN(
        n6151) );
  OAI21_X1 U7181 ( .B1(n6152), .B2(n6210), .A(n6151), .ZN(U2934) );
  AND2_X1 U7182 ( .A1(n6207), .A2(DATAI_11_), .ZN(n6194) );
  AOI21_X1 U7183 ( .B1(UWORD_REG_11__SCAN_IN), .B2(n6201), .A(n6194), .ZN(
        n6153) );
  OAI21_X1 U7184 ( .B1(n6154), .B2(n6210), .A(n6153), .ZN(U2935) );
  AND2_X1 U7185 ( .A1(n6207), .A2(DATAI_12_), .ZN(n6197) );
  AOI21_X1 U7186 ( .B1(UWORD_REG_12__SCAN_IN), .B2(n6201), .A(n6197), .ZN(
        n6155) );
  OAI21_X1 U7187 ( .B1(n6156), .B2(n6210), .A(n6155), .ZN(U2936) );
  AND2_X1 U7188 ( .A1(n6207), .A2(DATAI_13_), .ZN(n6200) );
  AOI21_X1 U7189 ( .B1(UWORD_REG_13__SCAN_IN), .B2(n6201), .A(n6200), .ZN(
        n6157) );
  OAI21_X1 U7190 ( .B1(n6158), .B2(n6210), .A(n6157), .ZN(U2937) );
  AND2_X1 U7191 ( .A1(n6207), .A2(DATAI_14_), .ZN(n6204) );
  AOI21_X1 U7192 ( .B1(UWORD_REG_14__SCAN_IN), .B2(n6201), .A(n6204), .ZN(
        n6159) );
  OAI21_X1 U7193 ( .B1(n6160), .B2(n6210), .A(n6159), .ZN(U2938) );
  AOI21_X1 U7194 ( .B1(LWORD_REG_0__SCAN_IN), .B2(n6201), .A(n6161), .ZN(n6162) );
  OAI21_X1 U7195 ( .B1(n6163), .B2(n6210), .A(n6162), .ZN(U2939) );
  AOI21_X1 U7196 ( .B1(LWORD_REG_1__SCAN_IN), .B2(n6201), .A(n6164), .ZN(n6165) );
  OAI21_X1 U7197 ( .B1(n6166), .B2(n6210), .A(n6165), .ZN(U2940) );
  AOI21_X1 U7198 ( .B1(LWORD_REG_2__SCAN_IN), .B2(n6201), .A(n6167), .ZN(n6168) );
  OAI21_X1 U7199 ( .B1(n6169), .B2(n6210), .A(n6168), .ZN(U2941) );
  AOI21_X1 U7200 ( .B1(LWORD_REG_3__SCAN_IN), .B2(n6201), .A(n6170), .ZN(n6171) );
  OAI21_X1 U7201 ( .B1(n6172), .B2(n6210), .A(n6171), .ZN(U2942) );
  AOI21_X1 U7202 ( .B1(LWORD_REG_4__SCAN_IN), .B2(n6201), .A(n6173), .ZN(n6174) );
  OAI21_X1 U7203 ( .B1(n6175), .B2(n6210), .A(n6174), .ZN(U2943) );
  AOI21_X1 U7204 ( .B1(LWORD_REG_5__SCAN_IN), .B2(n6201), .A(n6176), .ZN(n6177) );
  OAI21_X1 U7205 ( .B1(n6178), .B2(n6210), .A(n6177), .ZN(U2944) );
  AOI21_X1 U7206 ( .B1(LWORD_REG_6__SCAN_IN), .B2(n6201), .A(n6179), .ZN(n6180) );
  OAI21_X1 U7207 ( .B1(n6181), .B2(n6210), .A(n6180), .ZN(U2945) );
  AOI21_X1 U7208 ( .B1(LWORD_REG_7__SCAN_IN), .B2(n6201), .A(n6182), .ZN(n6183) );
  OAI21_X1 U7209 ( .B1(n6184), .B2(n6210), .A(n6183), .ZN(U2946) );
  AOI21_X1 U7210 ( .B1(LWORD_REG_8__SCAN_IN), .B2(n6201), .A(n6185), .ZN(n6186) );
  OAI21_X1 U7211 ( .B1(n6187), .B2(n6210), .A(n6186), .ZN(U2947) );
  AOI21_X1 U7212 ( .B1(LWORD_REG_9__SCAN_IN), .B2(n6201), .A(n6188), .ZN(n6189) );
  OAI21_X1 U7213 ( .B1(n6190), .B2(n6210), .A(n6189), .ZN(U2948) );
  AOI21_X1 U7214 ( .B1(LWORD_REG_10__SCAN_IN), .B2(n6201), .A(n6191), .ZN(
        n6192) );
  OAI21_X1 U7215 ( .B1(n6193), .B2(n6210), .A(n6192), .ZN(U2949) );
  AOI21_X1 U7216 ( .B1(LWORD_REG_11__SCAN_IN), .B2(n6201), .A(n6194), .ZN(
        n6195) );
  OAI21_X1 U7217 ( .B1(n6196), .B2(n6210), .A(n6195), .ZN(U2950) );
  AOI21_X1 U7218 ( .B1(LWORD_REG_12__SCAN_IN), .B2(n6201), .A(n6197), .ZN(
        n6198) );
  OAI21_X1 U7219 ( .B1(n6199), .B2(n6210), .A(n6198), .ZN(U2951) );
  AOI21_X1 U7220 ( .B1(LWORD_REG_13__SCAN_IN), .B2(n6201), .A(n6200), .ZN(
        n6202) );
  OAI21_X1 U7221 ( .B1(n6203), .B2(n6210), .A(n6202), .ZN(U2952) );
  AOI21_X1 U7222 ( .B1(LWORD_REG_14__SCAN_IN), .B2(n6208), .A(n6204), .ZN(
        n6205) );
  OAI21_X1 U7223 ( .B1(n6206), .B2(n6210), .A(n6205), .ZN(U2953) );
  AOI22_X1 U7224 ( .A1(n6208), .A2(LWORD_REG_15__SCAN_IN), .B1(n6207), .B2(
        DATAI_15_), .ZN(n6209) );
  OAI21_X1 U7225 ( .B1(n6211), .B2(n6210), .A(n6209), .ZN(U2954) );
  NAND2_X1 U7226 ( .A1(n6213), .A2(n6212), .ZN(n6215) );
  XNOR2_X1 U7227 ( .A(n3437), .B(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n6214)
         );
  XNOR2_X1 U7228 ( .A(n6215), .B(n6214), .ZN(n6261) );
  AOI22_X1 U7229 ( .A1(n2993), .A2(REIP_REG_11__SCAN_IN), .B1(n6239), .B2(
        PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n6220) );
  AOI22_X1 U7230 ( .A1(n6218), .A2(n6244), .B1(n6217), .B2(n6216), .ZN(n6219)
         );
  OAI211_X1 U7231 ( .C1(n6261), .C2(n6221), .A(n6220), .B(n6219), .ZN(U2975)
         );
  AOI22_X1 U7232 ( .A1(n2993), .A2(REIP_REG_6__SCAN_IN), .B1(n6239), .B2(
        PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n6228) );
  OAI21_X1 U7233 ( .B1(n6224), .B2(n6223), .A(n6222), .ZN(n6299) );
  INV_X1 U7234 ( .A(n6299), .ZN(n6226) );
  AOI22_X1 U7235 ( .A1(n6226), .A2(n6243), .B1(n6244), .B2(n6225), .ZN(n6227)
         );
  OAI211_X1 U7236 ( .C1(n6249), .C2(n6229), .A(n6228), .B(n6227), .ZN(U2980)
         );
  AOI22_X1 U7237 ( .A1(n2993), .A2(REIP_REG_4__SCAN_IN), .B1(n6239), .B2(
        PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n6237) );
  OAI21_X1 U7238 ( .B1(n6232), .B2(n6231), .A(n6230), .ZN(n6233) );
  INV_X1 U7239 ( .A(n6233), .ZN(n6318) );
  INV_X1 U7240 ( .A(n6234), .ZN(n6235) );
  AOI22_X1 U7241 ( .A1(n6318), .A2(n6243), .B1(n6244), .B2(n6235), .ZN(n6236)
         );
  OAI211_X1 U7242 ( .C1(n6249), .C2(n6238), .A(n6237), .B(n6236), .ZN(U2982)
         );
  AOI22_X1 U7243 ( .A1(n2993), .A2(REIP_REG_2__SCAN_IN), .B1(n6239), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n6247) );
  XNOR2_X1 U7244 ( .A(n6240), .B(n3306), .ZN(n6242) );
  XNOR2_X1 U7245 ( .A(n6242), .B(n6241), .ZN(n6341) );
  AOI22_X1 U7246 ( .A1(n6245), .A2(n6244), .B1(n6243), .B2(n6341), .ZN(n6246)
         );
  OAI211_X1 U7247 ( .C1(n6249), .C2(n6248), .A(n6247), .B(n6246), .ZN(U2984)
         );
  NAND2_X1 U7248 ( .A1(INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n6257), .ZN(n6255) );
  AOI21_X1 U7249 ( .B1(n6257), .B2(n3438), .A(n6258), .ZN(n6253) );
  AOI222_X1 U7250 ( .A1(n6251), .A2(n6340), .B1(n6323), .B2(n6250), .C1(
        REIP_REG_12__SCAN_IN), .C2(n2993), .ZN(n6252) );
  OAI221_X1 U7251 ( .B1(INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n6255), .C1(
        n6254), .C2(n6253), .A(n6252), .ZN(U3006) );
  AOI22_X1 U7252 ( .A1(n6256), .A2(n6323), .B1(n2993), .B2(
        REIP_REG_11__SCAN_IN), .ZN(n6260) );
  AOI22_X1 U7253 ( .A1(INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n6258), .B1(n6257), .B2(n3438), .ZN(n6259) );
  OAI211_X1 U7254 ( .C1(n6261), .C2(n6300), .A(n6260), .B(n6259), .ZN(U3007)
         );
  AOI21_X1 U7255 ( .B1(n6263), .B2(n6329), .A(n6262), .ZN(n6286) );
  AOI21_X1 U7256 ( .B1(n6282), .B2(n6297), .A(n6286), .ZN(n6278) );
  INV_X1 U7257 ( .A(n6264), .ZN(n6269) );
  NOR3_X1 U7258 ( .A1(n6304), .A2(n6296), .A3(n6314), .ZN(n6290) );
  NAND2_X1 U7259 ( .A1(n6265), .A2(n6290), .ZN(n6274) );
  AOI221_X1 U7260 ( .B1(INSTADDRPOINTER_REG_9__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_10__SCAN_IN), .C1(n5184), .C2(n3928), .A(n6274), 
        .ZN(n6268) );
  OAI22_X1 U7261 ( .A1(n6266), .A2(n6337), .B1(n6544), .B2(n6335), .ZN(n6267)
         );
  AOI211_X1 U7262 ( .C1(n6269), .C2(n6340), .A(n6268), .B(n6267), .ZN(n6270)
         );
  OAI21_X1 U7263 ( .B1(n6278), .B2(n3928), .A(n6270), .ZN(U3008) );
  AOI21_X1 U7264 ( .B1(n6272), .B2(n6323), .A(n6271), .ZN(n6273) );
  OAI21_X1 U7265 ( .B1(n6274), .B2(INSTADDRPOINTER_REG_9__SCAN_IN), .A(n6273), 
        .ZN(n6275) );
  AOI21_X1 U7266 ( .B1(n6276), .B2(n6340), .A(n6275), .ZN(n6277) );
  OAI21_X1 U7267 ( .B1(n6278), .B2(n5184), .A(n6277), .ZN(U3009) );
  AOI21_X1 U7268 ( .B1(n6280), .B2(n6323), .A(n6279), .ZN(n6285) );
  AOI22_X1 U7269 ( .A1(n6281), .A2(n6340), .B1(INSTADDRPOINTER_REG_8__SCAN_IN), 
        .B2(n6286), .ZN(n6284) );
  OAI211_X1 U7270 ( .C1(INSTADDRPOINTER_REG_7__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_8__SCAN_IN), .A(n6290), .B(n6282), .ZN(n6283) );
  NAND3_X1 U7271 ( .A1(n6285), .A2(n6284), .A3(n6283), .ZN(U3010) );
  INV_X1 U7272 ( .A(n6286), .ZN(n6294) );
  AOI21_X1 U7273 ( .B1(n6288), .B2(n6323), .A(n6287), .ZN(n6293) );
  INV_X1 U7274 ( .A(n6289), .ZN(n6291) );
  AOI22_X1 U7275 ( .A1(n6291), .A2(n6340), .B1(n6290), .B2(n6295), .ZN(n6292)
         );
  OAI211_X1 U7276 ( .C1(n6295), .C2(n6294), .A(n6293), .B(n6292), .ZN(U3011)
         );
  OR2_X1 U7277 ( .A1(n6296), .A2(n6314), .ZN(n6305) );
  AOI221_X1 U7278 ( .B1(n6298), .B2(n6297), .C1(n6296), .C2(n6297), .A(n6332), 
        .ZN(n6312) );
  INV_X1 U7279 ( .A(REIP_REG_6__SCAN_IN), .ZN(n6539) );
  OAI222_X1 U7280 ( .A1(n6301), .A2(n6337), .B1(n6335), .B2(n6539), .C1(n6300), 
        .C2(n6299), .ZN(n6302) );
  INV_X1 U7281 ( .A(n6302), .ZN(n6303) );
  OAI221_X1 U7282 ( .B1(INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n6305), .C1(n6304), .C2(n6312), .A(n6303), .ZN(U3012) );
  NOR2_X1 U7283 ( .A1(n6328), .A2(n6320), .ZN(n6315) );
  AOI21_X1 U7284 ( .B1(n6315), .B2(n6324), .A(INSTADDRPOINTER_REG_5__SCAN_IN), 
        .ZN(n6311) );
  INV_X1 U7285 ( .A(n6306), .ZN(n6308) );
  AOI22_X1 U7286 ( .A1(n6308), .A2(n6340), .B1(n6323), .B2(n6307), .ZN(n6310)
         );
  NAND2_X1 U7287 ( .A1(n2993), .A2(REIP_REG_5__SCAN_IN), .ZN(n6309) );
  OAI211_X1 U7288 ( .C1(n6312), .C2(n6311), .A(n6310), .B(n6309), .ZN(U3013)
         );
  OAI22_X1 U7289 ( .A1(n6337), .A2(n6313), .B1(n6536), .B2(n6335), .ZN(n6317)
         );
  AOI211_X1 U7290 ( .C1(n6328), .C2(n6320), .A(n6315), .B(n6314), .ZN(n6316)
         );
  AOI211_X1 U7291 ( .C1(n6318), .C2(n6340), .A(n6317), .B(n6316), .ZN(n6319)
         );
  OAI21_X1 U7292 ( .B1(n6329), .B2(n6320), .A(n6319), .ZN(U3014) );
  AOI21_X1 U7293 ( .B1(n6323), .B2(n6322), .A(n6321), .ZN(n6327) );
  AOI22_X1 U7294 ( .A1(n6325), .A2(n6340), .B1(n6324), .B2(n6328), .ZN(n6326)
         );
  OAI211_X1 U7295 ( .C1(n6329), .C2(n6328), .A(n6327), .B(n6326), .ZN(U3015)
         );
  OR2_X1 U7296 ( .A1(n6331), .A2(n6330), .ZN(n6344) );
  AOI21_X1 U7297 ( .B1(n6334), .B2(n6333), .A(n6332), .ZN(n6343) );
  INV_X1 U7298 ( .A(REIP_REG_2__SCAN_IN), .ZN(n6533) );
  OAI22_X1 U7299 ( .A1(n6337), .A2(n6336), .B1(n6533), .B2(n6335), .ZN(n6338)
         );
  AOI211_X1 U7300 ( .C1(n6341), .C2(n6340), .A(n6339), .B(n6338), .ZN(n6342)
         );
  OAI221_X1 U7301 ( .B1(INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n6344), .C1(n3306), .C2(n6343), .A(n6342), .ZN(U3016) );
  NOR2_X1 U7302 ( .A1(n6346), .A2(n6345), .ZN(U3019) );
  NOR2_X1 U7303 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6347), .ZN(n6389)
         );
  INV_X1 U7304 ( .A(n6348), .ZN(n6353) );
  INV_X1 U7305 ( .A(n6349), .ZN(n6351) );
  OAI22_X1 U7306 ( .A1(n6353), .A2(n6352), .B1(n6351), .B2(n6350), .ZN(n6387)
         );
  AOI22_X1 U7307 ( .A1(n6397), .A2(n6389), .B1(n6429), .B2(n6387), .ZN(n6362)
         );
  INV_X1 U7308 ( .A(n6424), .ZN(n6354) );
  OAI21_X1 U7309 ( .B1(n6391), .B2(n6354), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n6357) );
  AOI211_X1 U7310 ( .C1(n6358), .C2(n6357), .A(n6356), .B(n6355), .ZN(n6359)
         );
  AOI22_X1 U7311 ( .A1(n6393), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n6360), 
        .B2(n6391), .ZN(n6361) );
  OAI211_X1 U7312 ( .C1(n6427), .C2(n6424), .A(n6362), .B(n6361), .ZN(U3068)
         );
  AOI22_X1 U7313 ( .A1(n6401), .A2(n6389), .B1(n6436), .B2(n6387), .ZN(n6365)
         );
  AOI22_X1 U7314 ( .A1(n6393), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n6363), 
        .B2(n6391), .ZN(n6364) );
  OAI211_X1 U7315 ( .C1(n6434), .C2(n6424), .A(n6365), .B(n6364), .ZN(U3069)
         );
  AOI22_X1 U7316 ( .A1(n6367), .A2(n6389), .B1(n6366), .B2(n6387), .ZN(n6370)
         );
  AOI22_X1 U7317 ( .A1(n6393), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n6368), 
        .B2(n6391), .ZN(n6369) );
  OAI211_X1 U7318 ( .C1(n6371), .C2(n6424), .A(n6370), .B(n6369), .ZN(U3070)
         );
  AOI22_X1 U7319 ( .A1(n6405), .A2(n6389), .B1(n6407), .B2(n6387), .ZN(n6374)
         );
  AOI22_X1 U7320 ( .A1(n6393), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n6372), 
        .B2(n6391), .ZN(n6373) );
  OAI211_X1 U7321 ( .C1(n6375), .C2(n6424), .A(n6374), .B(n6373), .ZN(U3071)
         );
  AOI22_X1 U7322 ( .A1(n6376), .A2(n6389), .B1(n6443), .B2(n6387), .ZN(n6379)
         );
  AOI22_X1 U7323 ( .A1(n6393), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n6377), 
        .B2(n6391), .ZN(n6378) );
  OAI211_X1 U7324 ( .C1(n6441), .C2(n6424), .A(n6379), .B(n6378), .ZN(U3072)
         );
  AOI22_X1 U7325 ( .A1(n6411), .A2(n6389), .B1(n6453), .B2(n6387), .ZN(n6382)
         );
  AOI22_X1 U7326 ( .A1(n6393), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n6380), 
        .B2(n6391), .ZN(n6381) );
  OAI211_X1 U7327 ( .C1(n6449), .C2(n6424), .A(n6382), .B(n6381), .ZN(U3073)
         );
  AOI22_X1 U7328 ( .A1(n6415), .A2(n6389), .B1(n6420), .B2(n6387), .ZN(n6385)
         );
  AOI22_X1 U7329 ( .A1(n6393), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n6383), 
        .B2(n6391), .ZN(n6384) );
  OAI211_X1 U7330 ( .C1(n6386), .C2(n6424), .A(n6385), .B(n6384), .ZN(U3074)
         );
  AOI22_X1 U7331 ( .A1(n6390), .A2(n6389), .B1(n6388), .B2(n6387), .ZN(n6395)
         );
  AOI22_X1 U7332 ( .A1(n6393), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n6392), 
        .B2(n6391), .ZN(n6394) );
  OAI211_X1 U7333 ( .C1(n6396), .C2(n6424), .A(n6395), .B(n6394), .ZN(U3075)
         );
  AOI22_X1 U7334 ( .A1(n6418), .A2(n6398), .B1(n6416), .B2(n6397), .ZN(n6400)
         );
  AOI22_X1 U7335 ( .A1(INSTQUEUE_REG_7__0__SCAN_IN), .A2(n6421), .B1(n6429), 
        .B2(n6419), .ZN(n6399) );
  OAI211_X1 U7336 ( .C1(n6432), .C2(n6424), .A(n6400), .B(n6399), .ZN(U3076)
         );
  AOI22_X1 U7337 ( .A1(n6418), .A2(n6402), .B1(n6416), .B2(n6401), .ZN(n6404)
         );
  AOI22_X1 U7338 ( .A1(INSTQUEUE_REG_7__1__SCAN_IN), .A2(n6421), .B1(n6436), 
        .B2(n6419), .ZN(n6403) );
  OAI211_X1 U7339 ( .C1(n6439), .C2(n6424), .A(n6404), .B(n6403), .ZN(U3077)
         );
  AOI22_X1 U7340 ( .A1(n6418), .A2(n6406), .B1(n6416), .B2(n6405), .ZN(n6409)
         );
  AOI22_X1 U7341 ( .A1(INSTQUEUE_REG_7__3__SCAN_IN), .A2(n6421), .B1(n6407), 
        .B2(n6419), .ZN(n6408) );
  OAI211_X1 U7342 ( .C1(n6410), .C2(n6424), .A(n6409), .B(n6408), .ZN(U3079)
         );
  AOI22_X1 U7343 ( .A1(n6418), .A2(n6412), .B1(n6416), .B2(n6411), .ZN(n6414)
         );
  AOI22_X1 U7344 ( .A1(INSTQUEUE_REG_7__5__SCAN_IN), .A2(n6421), .B1(n6453), 
        .B2(n6419), .ZN(n6413) );
  OAI211_X1 U7345 ( .C1(n6458), .C2(n6424), .A(n6414), .B(n6413), .ZN(U3081)
         );
  AOI22_X1 U7346 ( .A1(n6418), .A2(n6417), .B1(n6416), .B2(n6415), .ZN(n6423)
         );
  AOI22_X1 U7347 ( .A1(INSTQUEUE_REG_7__6__SCAN_IN), .A2(n6421), .B1(n6420), 
        .B2(n6419), .ZN(n6422) );
  OAI211_X1 U7348 ( .C1(n6425), .C2(n6424), .A(n6423), .B(n6422), .ZN(U3082)
         );
  OAI22_X1 U7349 ( .A1(n6450), .A2(n6427), .B1(n6426), .B2(n6447), .ZN(n6428)
         );
  INV_X1 U7350 ( .A(n6428), .ZN(n6431) );
  AOI22_X1 U7351 ( .A1(INSTQUEUE_REG_11__0__SCAN_IN), .A2(n6454), .B1(n6429), 
        .B2(n6452), .ZN(n6430) );
  OAI211_X1 U7352 ( .C1(n6432), .C2(n6457), .A(n6431), .B(n6430), .ZN(U3108)
         );
  OAI22_X1 U7353 ( .A1(n6450), .A2(n6434), .B1(n6433), .B2(n6447), .ZN(n6435)
         );
  INV_X1 U7354 ( .A(n6435), .ZN(n6438) );
  AOI22_X1 U7355 ( .A1(INSTQUEUE_REG_11__1__SCAN_IN), .A2(n6454), .B1(n6436), 
        .B2(n6452), .ZN(n6437) );
  OAI211_X1 U7356 ( .C1(n6439), .C2(n6457), .A(n6438), .B(n6437), .ZN(U3109)
         );
  OAI22_X1 U7357 ( .A1(n6450), .A2(n6441), .B1(n6440), .B2(n6447), .ZN(n6442)
         );
  INV_X1 U7358 ( .A(n6442), .ZN(n6445) );
  AOI22_X1 U7359 ( .A1(INSTQUEUE_REG_11__4__SCAN_IN), .A2(n6454), .B1(n6443), 
        .B2(n6452), .ZN(n6444) );
  OAI211_X1 U7360 ( .C1(n6446), .C2(n6457), .A(n6445), .B(n6444), .ZN(U3112)
         );
  OAI22_X1 U7361 ( .A1(n6450), .A2(n6449), .B1(n6448), .B2(n6447), .ZN(n6451)
         );
  INV_X1 U7362 ( .A(n6451), .ZN(n6456) );
  AOI22_X1 U7363 ( .A1(INSTQUEUE_REG_11__5__SCAN_IN), .A2(n6454), .B1(n6453), 
        .B2(n6452), .ZN(n6455) );
  OAI211_X1 U7364 ( .C1(n6458), .C2(n6457), .A(n6456), .B(n6455), .ZN(U3113)
         );
  INV_X1 U7365 ( .A(n6475), .ZN(n6477) );
  NOR2_X1 U7366 ( .A1(n6460), .A2(n6459), .ZN(n6465) );
  NAND2_X1 U7367 ( .A1(n6465), .A2(n6464), .ZN(n6467) );
  OAI211_X1 U7368 ( .C1(n3153), .C2(n6462), .A(n6461), .B(
        INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n6463) );
  OAI21_X1 U7369 ( .B1(n6465), .B2(n6464), .A(n6463), .ZN(n6466) );
  NAND2_X1 U7370 ( .A1(n6467), .A2(n6466), .ZN(n6469) );
  INV_X1 U7371 ( .A(n6469), .ZN(n6472) );
  NAND2_X1 U7372 ( .A1(n6469), .A2(n6468), .ZN(n6471) );
  AOI22_X1 U7373 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n6472), .B1(n6471), .B2(n6470), .ZN(n6473) );
  AOI21_X1 U7374 ( .B1(n6475), .B2(n6474), .A(n6473), .ZN(n6476) );
  AOI211_X1 U7375 ( .C1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .C2(n6477), .A(
        INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B(n6476), .ZN(n6485) );
  OAI21_X1 U7376 ( .B1(FLUSH_REG_SCAN_IN), .B2(MORE_REG_SCAN_IN), .A(n6478), 
        .ZN(n6481) );
  NAND3_X1 U7377 ( .A1(n6481), .A2(n6480), .A3(n6479), .ZN(n6482) );
  NOR4_X1 U7378 ( .A1(n6485), .A2(n6484), .A3(n6483), .A4(n6482), .ZN(n6496)
         );
  INV_X1 U7379 ( .A(n6496), .ZN(n6488) );
  OAI22_X1 U7380 ( .A1(n6488), .A2(n6500), .B1(n6487), .B2(n6486), .ZN(n6489)
         );
  OAI21_X1 U7381 ( .B1(n6491), .B2(n6490), .A(n6489), .ZN(n6580) );
  OAI21_X1 U7382 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n6487), .A(n6580), .ZN(
        n6499) );
  AOI221_X1 U7383 ( .B1(n6493), .B2(STATE2_REG_0__SCAN_IN), .C1(n6499), .C2(
        STATE2_REG_0__SCAN_IN), .A(n6492), .ZN(n6495) );
  OAI211_X1 U7384 ( .C1(n6507), .C2(n6583), .A(n6498), .B(n6580), .ZN(n6494)
         );
  OAI211_X1 U7385 ( .C1(n6496), .C2(n6500), .A(n6495), .B(n6494), .ZN(U3148)
         );
  NAND2_X1 U7386 ( .A1(n6498), .A2(n6497), .ZN(n6506) );
  NAND3_X1 U7387 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n6506), .A3(n6499), .ZN(
        n6505) );
  OAI21_X1 U7388 ( .B1(READY_N), .B2(n6501), .A(n6500), .ZN(n6503) );
  AOI21_X1 U7389 ( .B1(n6503), .B2(n6580), .A(n6502), .ZN(n6504) );
  NAND2_X1 U7390 ( .A1(n6505), .A2(n6504), .ZN(U3149) );
  INV_X1 U7391 ( .A(n6506), .ZN(n6510) );
  OAI211_X1 U7392 ( .C1(STATE2_REG_2__SCAN_IN), .C2(n6487), .A(n6579), .B(
        n6507), .ZN(n6509) );
  OAI21_X1 U7393 ( .B1(n6510), .B2(n6509), .A(n6508), .ZN(U3150) );
  AND2_X1 U7394 ( .A1(DATAWIDTH_REG_31__SCAN_IN), .A2(n6511), .ZN(U3151) );
  AND2_X1 U7395 ( .A1(DATAWIDTH_REG_30__SCAN_IN), .A2(n6511), .ZN(U3152) );
  AND2_X1 U7396 ( .A1(DATAWIDTH_REG_29__SCAN_IN), .A2(n6511), .ZN(U3153) );
  AND2_X1 U7397 ( .A1(DATAWIDTH_REG_28__SCAN_IN), .A2(n6511), .ZN(U3154) );
  AND2_X1 U7398 ( .A1(DATAWIDTH_REG_27__SCAN_IN), .A2(n6511), .ZN(U3155) );
  AND2_X1 U7399 ( .A1(DATAWIDTH_REG_26__SCAN_IN), .A2(n6511), .ZN(U3156) );
  AND2_X1 U7400 ( .A1(DATAWIDTH_REG_25__SCAN_IN), .A2(n6511), .ZN(U3157) );
  AND2_X1 U7401 ( .A1(DATAWIDTH_REG_24__SCAN_IN), .A2(n6511), .ZN(U3158) );
  AND2_X1 U7402 ( .A1(DATAWIDTH_REG_23__SCAN_IN), .A2(n6511), .ZN(U3159) );
  AND2_X1 U7403 ( .A1(DATAWIDTH_REG_22__SCAN_IN), .A2(n6511), .ZN(U3160) );
  AND2_X1 U7404 ( .A1(DATAWIDTH_REG_21__SCAN_IN), .A2(n6511), .ZN(U3161) );
  AND2_X1 U7405 ( .A1(DATAWIDTH_REG_20__SCAN_IN), .A2(n6511), .ZN(U3162) );
  AND2_X1 U7406 ( .A1(DATAWIDTH_REG_19__SCAN_IN), .A2(n6511), .ZN(U3163) );
  AND2_X1 U7407 ( .A1(DATAWIDTH_REG_18__SCAN_IN), .A2(n6511), .ZN(U3164) );
  AND2_X1 U7408 ( .A1(DATAWIDTH_REG_17__SCAN_IN), .A2(n6511), .ZN(U3165) );
  AND2_X1 U7409 ( .A1(DATAWIDTH_REG_16__SCAN_IN), .A2(n6511), .ZN(U3166) );
  AND2_X1 U7410 ( .A1(DATAWIDTH_REG_15__SCAN_IN), .A2(n6511), .ZN(U3167) );
  AND2_X1 U7411 ( .A1(DATAWIDTH_REG_14__SCAN_IN), .A2(n6511), .ZN(U3168) );
  AND2_X1 U7412 ( .A1(DATAWIDTH_REG_13__SCAN_IN), .A2(n6511), .ZN(U3169) );
  AND2_X1 U7413 ( .A1(DATAWIDTH_REG_12__SCAN_IN), .A2(n6511), .ZN(U3170) );
  AND2_X1 U7414 ( .A1(DATAWIDTH_REG_11__SCAN_IN), .A2(n6511), .ZN(U3171) );
  AND2_X1 U7415 ( .A1(DATAWIDTH_REG_10__SCAN_IN), .A2(n6511), .ZN(U3172) );
  AND2_X1 U7416 ( .A1(DATAWIDTH_REG_9__SCAN_IN), .A2(n6511), .ZN(U3173) );
  AND2_X1 U7417 ( .A1(DATAWIDTH_REG_8__SCAN_IN), .A2(n6511), .ZN(U3174) );
  AND2_X1 U7418 ( .A1(DATAWIDTH_REG_7__SCAN_IN), .A2(n6511), .ZN(U3175) );
  AND2_X1 U7419 ( .A1(DATAWIDTH_REG_6__SCAN_IN), .A2(n6511), .ZN(U3176) );
  AND2_X1 U7420 ( .A1(DATAWIDTH_REG_5__SCAN_IN), .A2(n6511), .ZN(U3177) );
  AND2_X1 U7421 ( .A1(DATAWIDTH_REG_4__SCAN_IN), .A2(n6511), .ZN(U3178) );
  AND2_X1 U7422 ( .A1(DATAWIDTH_REG_3__SCAN_IN), .A2(n6511), .ZN(U3179) );
  AND2_X1 U7423 ( .A1(DATAWIDTH_REG_2__SCAN_IN), .A2(n6511), .ZN(U3180) );
  NAND2_X1 U7424 ( .A1(STATE_REG_1__SCAN_IN), .A2(HOLD), .ZN(n6517) );
  NAND2_X1 U7425 ( .A1(STATE_REG_2__SCAN_IN), .A2(HOLD), .ZN(n6516) );
  NAND2_X1 U7426 ( .A1(READY_N), .A2(STATE_REG_1__SCAN_IN), .ZN(n6524) );
  NAND2_X1 U7427 ( .A1(n6516), .A2(n6524), .ZN(n6513) );
  INV_X1 U7428 ( .A(NA_N), .ZN(n6633) );
  INV_X1 U7429 ( .A(n6514), .ZN(n6512) );
  AOI211_X1 U7430 ( .C1(STATE_REG_2__SCAN_IN), .C2(n6633), .A(
        STATE_REG_0__SCAN_IN), .B(n6512), .ZN(n6529) );
  AOI21_X1 U7431 ( .B1(n6514), .B2(n6513), .A(n6529), .ZN(n6515) );
  OAI221_X1 U7432 ( .B1(n6804), .B2(REQUESTPENDING_REG_SCAN_IN), .C1(n6804), 
        .C2(n6517), .A(n6515), .ZN(U3181) );
  INV_X1 U7433 ( .A(n6516), .ZN(n6521) );
  INV_X1 U7434 ( .A(n6517), .ZN(n6518) );
  AOI21_X1 U7435 ( .B1(REQUESTPENDING_REG_SCAN_IN), .B2(STATE_REG_0__SCAN_IN), 
        .A(n6518), .ZN(n6520) );
  OAI211_X1 U7436 ( .C1(n6521), .C2(n6520), .A(n6519), .B(n6524), .ZN(U3182)
         );
  AOI221_X1 U7437 ( .B1(NA_N), .B2(STATE_REG_1__SCAN_IN), .C1(n6487), .C2(
        STATE_REG_1__SCAN_IN), .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n6523) );
  AOI221_X1 U7438 ( .B1(STATE_REG_2__SCAN_IN), .B2(HOLD), .C1(n6523), .C2(HOLD), .A(n6522), .ZN(n6528) );
  INV_X1 U7439 ( .A(n6524), .ZN(n6525) );
  NAND4_X1 U7440 ( .A1(REQUESTPENDING_REG_SCAN_IN), .A2(STATE_REG_0__SCAN_IN), 
        .A3(n6525), .A4(n6633), .ZN(n6527) );
  NAND3_X1 U7441 ( .A1(READY_N), .A2(STATE_REG_2__SCAN_IN), .A3(
        STATE_REG_1__SCAN_IN), .ZN(n6526) );
  OAI211_X1 U7442 ( .C1(n6529), .C2(n6528), .A(n6527), .B(n6526), .ZN(U3183)
         );
  NAND2_X1 U7443 ( .A1(STATE_REG_2__SCAN_IN), .A2(n6804), .ZN(n6574) );
  INV_X1 U7444 ( .A(n6804), .ZN(n6803) );
  AOI22_X1 U7445 ( .A1(REIP_REG_2__SCAN_IN), .A2(n2985), .B1(
        ADDRESS_REG_0__SCAN_IN), .B2(n6803), .ZN(n6530) );
  OAI21_X1 U7446 ( .B1(n6531), .B2(n6574), .A(n6530), .ZN(U3184) );
  AOI22_X1 U7447 ( .A1(REIP_REG_3__SCAN_IN), .A2(n2985), .B1(
        ADDRESS_REG_1__SCAN_IN), .B2(n6803), .ZN(n6532) );
  OAI21_X1 U7448 ( .B1(n6533), .B2(n6574), .A(n6532), .ZN(U3185) );
  AOI22_X1 U7449 ( .A1(REIP_REG_4__SCAN_IN), .A2(n2985), .B1(
        ADDRESS_REG_2__SCAN_IN), .B2(n6565), .ZN(n6534) );
  OAI21_X1 U7450 ( .B1(n4543), .B2(n6574), .A(n6534), .ZN(U3186) );
  AOI22_X1 U7451 ( .A1(REIP_REG_5__SCAN_IN), .A2(n2985), .B1(
        ADDRESS_REG_3__SCAN_IN), .B2(n6565), .ZN(n6535) );
  OAI21_X1 U7452 ( .B1(n6536), .B2(n6574), .A(n6535), .ZN(U3187) );
  INV_X1 U7453 ( .A(n2985), .ZN(n6564) );
  INV_X1 U7454 ( .A(n6574), .ZN(n6562) );
  AOI22_X1 U7455 ( .A1(REIP_REG_5__SCAN_IN), .A2(n6562), .B1(
        ADDRESS_REG_4__SCAN_IN), .B2(n6565), .ZN(n6537) );
  OAI21_X1 U7456 ( .B1(n6539), .B2(n6564), .A(n6537), .ZN(U3188) );
  AOI22_X1 U7457 ( .A1(REIP_REG_7__SCAN_IN), .A2(n2985), .B1(
        ADDRESS_REG_5__SCAN_IN), .B2(n6565), .ZN(n6538) );
  OAI21_X1 U7458 ( .B1(n6539), .B2(n6574), .A(n6538), .ZN(U3189) );
  AOI22_X1 U7459 ( .A1(REIP_REG_7__SCAN_IN), .A2(n6562), .B1(
        ADDRESS_REG_6__SCAN_IN), .B2(n6565), .ZN(n6540) );
  OAI21_X1 U7460 ( .B1(n4971), .B2(n6564), .A(n6540), .ZN(U3190) );
  AOI22_X1 U7461 ( .A1(REIP_REG_9__SCAN_IN), .A2(n2985), .B1(
        ADDRESS_REG_7__SCAN_IN), .B2(n6565), .ZN(n6541) );
  OAI21_X1 U7462 ( .B1(n4971), .B2(n6574), .A(n6541), .ZN(U3191) );
  AOI22_X1 U7463 ( .A1(REIP_REG_9__SCAN_IN), .A2(n6562), .B1(
        ADDRESS_REG_8__SCAN_IN), .B2(n6565), .ZN(n6542) );
  OAI21_X1 U7464 ( .B1(n6544), .B2(n6564), .A(n6542), .ZN(U3192) );
  AOI22_X1 U7465 ( .A1(REIP_REG_11__SCAN_IN), .A2(n2985), .B1(
        ADDRESS_REG_9__SCAN_IN), .B2(n6565), .ZN(n6543) );
  OAI21_X1 U7466 ( .B1(n6544), .B2(n6574), .A(n6543), .ZN(U3193) );
  AOI22_X1 U7467 ( .A1(REIP_REG_11__SCAN_IN), .A2(n6562), .B1(
        ADDRESS_REG_10__SCAN_IN), .B2(n6565), .ZN(n6545) );
  OAI21_X1 U7468 ( .B1(n6547), .B2(n6564), .A(n6545), .ZN(U3194) );
  AOI22_X1 U7469 ( .A1(REIP_REG_13__SCAN_IN), .A2(n2985), .B1(
        ADDRESS_REG_11__SCAN_IN), .B2(n6565), .ZN(n6546) );
  OAI21_X1 U7470 ( .B1(n6547), .B2(n6574), .A(n6546), .ZN(U3195) );
  AOI22_X1 U7471 ( .A1(REIP_REG_14__SCAN_IN), .A2(n2985), .B1(
        ADDRESS_REG_12__SCAN_IN), .B2(n6565), .ZN(n6548) );
  OAI21_X1 U7472 ( .B1(n6549), .B2(n6574), .A(n6548), .ZN(U3196) );
  AOI22_X1 U7473 ( .A1(REIP_REG_14__SCAN_IN), .A2(n6562), .B1(
        ADDRESS_REG_13__SCAN_IN), .B2(n6565), .ZN(n6550) );
  OAI21_X1 U7474 ( .B1(n6552), .B2(n6564), .A(n6550), .ZN(U3197) );
  AOI22_X1 U7475 ( .A1(REIP_REG_16__SCAN_IN), .A2(n2985), .B1(
        ADDRESS_REG_14__SCAN_IN), .B2(n6565), .ZN(n6551) );
  OAI21_X1 U7476 ( .B1(n6552), .B2(n6574), .A(n6551), .ZN(U3198) );
  AOI22_X1 U7477 ( .A1(REIP_REG_16__SCAN_IN), .A2(n6562), .B1(
        ADDRESS_REG_15__SCAN_IN), .B2(n6565), .ZN(n6553) );
  OAI21_X1 U7478 ( .B1(n6555), .B2(n6564), .A(n6553), .ZN(U3199) );
  AOI22_X1 U7479 ( .A1(REIP_REG_18__SCAN_IN), .A2(n2985), .B1(
        ADDRESS_REG_16__SCAN_IN), .B2(n6565), .ZN(n6554) );
  OAI21_X1 U7480 ( .B1(n6555), .B2(n6574), .A(n6554), .ZN(U3200) );
  AOI22_X1 U7481 ( .A1(REIP_REG_18__SCAN_IN), .A2(n6562), .B1(
        ADDRESS_REG_17__SCAN_IN), .B2(n6565), .ZN(n6556) );
  OAI21_X1 U7482 ( .B1(n6706), .B2(n6564), .A(n6556), .ZN(U3201) );
  AOI22_X1 U7483 ( .A1(REIP_REG_20__SCAN_IN), .A2(n2985), .B1(
        ADDRESS_REG_18__SCAN_IN), .B2(n6565), .ZN(n6557) );
  OAI21_X1 U7484 ( .B1(n6706), .B2(n6574), .A(n6557), .ZN(U3202) );
  INV_X1 U7485 ( .A(REIP_REG_20__SCAN_IN), .ZN(n6640) );
  AOI22_X1 U7486 ( .A1(REIP_REG_21__SCAN_IN), .A2(n2985), .B1(
        ADDRESS_REG_19__SCAN_IN), .B2(n6565), .ZN(n6558) );
  OAI21_X1 U7487 ( .B1(n6640), .B2(n6574), .A(n6558), .ZN(U3203) );
  AOI22_X1 U7488 ( .A1(REIP_REG_21__SCAN_IN), .A2(n6562), .B1(
        ADDRESS_REG_20__SCAN_IN), .B2(n6565), .ZN(n6559) );
  OAI21_X1 U7489 ( .B1(n6560), .B2(n6564), .A(n6559), .ZN(U3204) );
  AOI22_X1 U7490 ( .A1(REIP_REG_22__SCAN_IN), .A2(n6562), .B1(
        ADDRESS_REG_21__SCAN_IN), .B2(n6565), .ZN(n6561) );
  OAI21_X1 U7491 ( .B1(n6666), .B2(n6564), .A(n6561), .ZN(U3205) );
  AOI22_X1 U7492 ( .A1(REIP_REG_23__SCAN_IN), .A2(n6562), .B1(
        ADDRESS_REG_22__SCAN_IN), .B2(n6565), .ZN(n6563) );
  OAI21_X1 U7493 ( .B1(n3883), .B2(n6564), .A(n6563), .ZN(U3206) );
  AOI22_X1 U7494 ( .A1(REIP_REG_25__SCAN_IN), .A2(n2985), .B1(
        ADDRESS_REG_23__SCAN_IN), .B2(n6565), .ZN(n6566) );
  OAI21_X1 U7495 ( .B1(n3883), .B2(n6574), .A(n6566), .ZN(U3207) );
  AOI22_X1 U7496 ( .A1(REIP_REG_26__SCAN_IN), .A2(n2985), .B1(
        ADDRESS_REG_24__SCAN_IN), .B2(n6803), .ZN(n6567) );
  OAI21_X1 U7497 ( .B1(n6749), .B2(n6574), .A(n6567), .ZN(U3208) );
  INV_X1 U7498 ( .A(REIP_REG_26__SCAN_IN), .ZN(n6731) );
  AOI22_X1 U7499 ( .A1(REIP_REG_27__SCAN_IN), .A2(n2985), .B1(
        ADDRESS_REG_25__SCAN_IN), .B2(n6803), .ZN(n6568) );
  OAI21_X1 U7500 ( .B1(n6731), .B2(n6574), .A(n6568), .ZN(U3209) );
  INV_X1 U7501 ( .A(REIP_REG_27__SCAN_IN), .ZN(n6611) );
  AOI22_X1 U7502 ( .A1(REIP_REG_28__SCAN_IN), .A2(n2985), .B1(
        ADDRESS_REG_26__SCAN_IN), .B2(n6803), .ZN(n6569) );
  OAI21_X1 U7503 ( .B1(n6611), .B2(n6574), .A(n6569), .ZN(U3210) );
  AOI22_X1 U7504 ( .A1(REIP_REG_29__SCAN_IN), .A2(n2985), .B1(
        ADDRESS_REG_27__SCAN_IN), .B2(n6803), .ZN(n6570) );
  OAI21_X1 U7505 ( .B1(n6771), .B2(n6574), .A(n6570), .ZN(U3211) );
  AOI22_X1 U7506 ( .A1(REIP_REG_30__SCAN_IN), .A2(n2985), .B1(
        ADDRESS_REG_28__SCAN_IN), .B2(n6803), .ZN(n6571) );
  OAI21_X1 U7507 ( .B1(n6702), .B2(n6574), .A(n6571), .ZN(U3212) );
  AOI22_X1 U7508 ( .A1(REIP_REG_31__SCAN_IN), .A2(n2985), .B1(
        ADDRESS_REG_29__SCAN_IN), .B2(n6803), .ZN(n6573) );
  OAI21_X1 U7509 ( .B1(n4307), .B2(n6574), .A(n6573), .ZN(U3213) );
  MUX2_X1 U7510 ( .A(BYTEENABLE_REG_2__SCAN_IN), .B(BE_N_REG_2__SCAN_IN), .S(
        n6803), .Z(U3446) );
  MUX2_X1 U7511 ( .A(BYTEENABLE_REG_1__SCAN_IN), .B(BE_N_REG_1__SCAN_IN), .S(
        n6803), .Z(U3447) );
  MUX2_X1 U7512 ( .A(BYTEENABLE_REG_0__SCAN_IN), .B(BE_N_REG_0__SCAN_IN), .S(
        n6803), .Z(U3448) );
  OAI21_X1 U7513 ( .B1(DATAWIDTH_REG_0__SCAN_IN), .B2(n6578), .A(n6576), .ZN(
        n6575) );
  INV_X1 U7514 ( .A(n6575), .ZN(U3451) );
  OAI21_X1 U7515 ( .B1(n6578), .B2(n6577), .A(n6576), .ZN(U3452) );
  OAI221_X1 U7516 ( .B1(n6581), .B2(STATE2_REG_0__SCAN_IN), .C1(n6581), .C2(
        n6580), .A(n6579), .ZN(U3453) );
  INV_X1 U7517 ( .A(n6582), .ZN(n6586) );
  OAI22_X1 U7518 ( .A1(n6586), .A2(n6585), .B1(n6584), .B2(n6583), .ZN(n6588)
         );
  MUX2_X1 U7519 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n6588), .S(n6587), 
        .Z(U3456) );
  AOI211_X1 U7520 ( .C1(REIP_REG_0__SCAN_IN), .C2(DATAWIDTH_REG_0__SCAN_IN), 
        .A(REIP_REG_1__SCAN_IN), .B(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6589) );
  AOI21_X1 U7521 ( .B1(REIP_REG_1__SCAN_IN), .B2(REIP_REG_0__SCAN_IN), .A(
        n6589), .ZN(n6590) );
  INV_X1 U7522 ( .A(BYTEENABLE_REG_2__SCAN_IN), .ZN(n6609) );
  AOI22_X1 U7523 ( .A1(n6593), .A2(n6590), .B1(n6609), .B2(n6591), .ZN(U3468)
         );
  NOR2_X1 U7524 ( .A1(REIP_REG_1__SCAN_IN), .A2(REIP_REG_0__SCAN_IN), .ZN(
        n6592) );
  INV_X1 U7525 ( .A(BYTEENABLE_REG_0__SCAN_IN), .ZN(n6627) );
  AOI22_X1 U7526 ( .A1(n6593), .A2(n6592), .B1(n6627), .B2(n6591), .ZN(U3469)
         );
  INV_X1 U7527 ( .A(READREQUEST_REG_SCAN_IN), .ZN(n6735) );
  OAI22_X1 U7528 ( .A1(n6803), .A2(n6735), .B1(W_R_N_REG_SCAN_IN), .B2(n6804), 
        .ZN(n6594) );
  INV_X1 U7529 ( .A(n6594), .ZN(U3470) );
  AOI211_X1 U7530 ( .C1(n6597), .C2(n6487), .A(n6596), .B(n6595), .ZN(n6604)
         );
  OAI211_X1 U7531 ( .C1(STATEBS16_REG_SCAN_IN), .C2(n6599), .A(n6598), .B(
        STATE2_REG_2__SCAN_IN), .ZN(n6601) );
  AOI21_X1 U7532 ( .B1(n6601), .B2(STATE2_REG_0__SCAN_IN), .A(n6600), .ZN(
        n6603) );
  NAND2_X1 U7533 ( .A1(n6604), .A2(REQUESTPENDING_REG_SCAN_IN), .ZN(n6602) );
  OAI21_X1 U7534 ( .B1(n6604), .B2(n6603), .A(n6602), .ZN(U3472) );
  OAI22_X1 U7535 ( .A1(n6803), .A2(MEMORYFETCH_REG_SCAN_IN), .B1(
        M_IO_N_REG_SCAN_IN), .B2(n6804), .ZN(n6605) );
  INV_X1 U7536 ( .A(n6605), .ZN(U3473) );
  INV_X1 U7537 ( .A(keyinput_f28), .ZN(n6694) );
  OAI22_X1 U7538 ( .A1(DATAI_14_), .A2(keyinput_f17), .B1(keyinput_f12), .B2(
        DATAI_19_), .ZN(n6606) );
  AOI221_X1 U7539 ( .B1(DATAI_14_), .B2(keyinput_f17), .C1(DATAI_19_), .C2(
        keyinput_f12), .A(n6606), .ZN(n6615) );
  OAI22_X1 U7540 ( .A1(REIP_REG_31__SCAN_IN), .A2(keyinput_f51), .B1(BS16_N), 
        .B2(keyinput_f34), .ZN(n6607) );
  AOI221_X1 U7541 ( .B1(REIP_REG_31__SCAN_IN), .B2(keyinput_f51), .C1(
        keyinput_f34), .C2(BS16_N), .A(n6607), .ZN(n6614) );
  OAI22_X1 U7542 ( .A1(keyinput_f49), .A2(n6609), .B1(n6751), .B2(keyinput_f38), .ZN(n6608) );
  AOI221_X1 U7543 ( .B1(n6609), .B2(keyinput_f49), .C1(n6751), .C2(
        keyinput_f38), .A(n6608), .ZN(n6613) );
  OAI22_X1 U7544 ( .A1(n6611), .A2(keyinput_f55), .B1(M_IO_N_REG_SCAN_IN), 
        .B2(keyinput_f40), .ZN(n6610) );
  AOI221_X1 U7545 ( .B1(n6611), .B2(keyinput_f55), .C1(keyinput_f40), .C2(
        M_IO_N_REG_SCAN_IN), .A(n6610), .ZN(n6612) );
  NAND4_X1 U7546 ( .A1(n6615), .A2(n6614), .A3(n6613), .A4(n6612), .ZN(n6692)
         );
  OAI22_X1 U7547 ( .A1(REIP_REG_19__SCAN_IN), .A2(keyinput_f63), .B1(DATAI_4_), 
        .B2(keyinput_f27), .ZN(n6616) );
  AOI221_X1 U7548 ( .B1(REIP_REG_19__SCAN_IN), .B2(keyinput_f63), .C1(
        keyinput_f27), .C2(DATAI_4_), .A(n6616), .ZN(n6623) );
  OAI22_X1 U7549 ( .A1(DATAI_1_), .A2(keyinput_f30), .B1(DATAI_17_), .B2(
        keyinput_f14), .ZN(n6617) );
  AOI221_X1 U7550 ( .B1(DATAI_1_), .B2(keyinput_f30), .C1(keyinput_f14), .C2(
        DATAI_17_), .A(n6617), .ZN(n6622) );
  OAI22_X1 U7551 ( .A1(keyinput_f36), .A2(HOLD), .B1(keyinput_f50), .B2(
        BYTEENABLE_REG_3__SCAN_IN), .ZN(n6618) );
  AOI221_X1 U7552 ( .B1(keyinput_f36), .B2(HOLD), .C1(
        BYTEENABLE_REG_3__SCAN_IN), .C2(keyinput_f50), .A(n6618), .ZN(n6621)
         );
  OAI22_X1 U7553 ( .A1(REIP_REG_22__SCAN_IN), .A2(keyinput_f60), .B1(DATAI_8_), 
        .B2(keyinput_f23), .ZN(n6619) );
  AOI221_X1 U7554 ( .B1(REIP_REG_22__SCAN_IN), .B2(keyinput_f60), .C1(
        keyinput_f23), .C2(DATAI_8_), .A(n6619), .ZN(n6620) );
  NAND4_X1 U7555 ( .A1(n6623), .A2(n6622), .A3(n6621), .A4(n6620), .ZN(n6691)
         );
  INV_X1 U7556 ( .A(DATAI_24_), .ZN(n6738) );
  INV_X1 U7557 ( .A(MORE_REG_SCAN_IN), .ZN(n6625) );
  OAI22_X1 U7558 ( .A1(n6738), .A2(keyinput_f7), .B1(n6625), .B2(keyinput_f44), 
        .ZN(n6624) );
  AOI221_X1 U7559 ( .B1(n6738), .B2(keyinput_f7), .C1(keyinput_f44), .C2(n6625), .A(n6624), .ZN(n6648) );
  OAI22_X1 U7560 ( .A1(n6702), .A2(keyinput_f53), .B1(n6627), .B2(keyinput_f47), .ZN(n6626) );
  AOI221_X1 U7561 ( .B1(n6702), .B2(keyinput_f53), .C1(keyinput_f47), .C2(
        n6627), .A(n6626), .ZN(n6647) );
  INV_X1 U7562 ( .A(DATAI_16_), .ZN(n6629) );
  OAI22_X1 U7563 ( .A1(n6629), .A2(keyinput_f15), .B1(n6748), .B2(keyinput_f48), .ZN(n6628) );
  AOI221_X1 U7564 ( .B1(n6629), .B2(keyinput_f15), .C1(keyinput_f48), .C2(
        n6748), .A(n6628), .ZN(n6631) );
  INV_X1 U7565 ( .A(DATAI_28_), .ZN(n6722) );
  XOR2_X1 U7566 ( .A(n6722), .B(keyinput_f3), .Z(n6630) );
  OAI211_X1 U7567 ( .C1(n6633), .C2(keyinput_f33), .A(n6631), .B(n6630), .ZN(
        n6632) );
  AOI21_X1 U7568 ( .B1(n6633), .B2(keyinput_f33), .A(n6632), .ZN(n6646) );
  AOI22_X1 U7569 ( .A1(n6699), .A2(keyinput_f20), .B1(keyinput_f16), .B2(n6705), .ZN(n6634) );
  OAI221_X1 U7570 ( .B1(n6699), .B2(keyinput_f20), .C1(n6705), .C2(
        keyinput_f16), .A(n6634), .ZN(n6644) );
  INV_X1 U7571 ( .A(MEMORYFETCH_REG_SCAN_IN), .ZN(n6636) );
  AOI22_X1 U7572 ( .A1(n6636), .A2(keyinput_f32), .B1(n6732), .B2(keyinput_f31), .ZN(n6635) );
  OAI221_X1 U7573 ( .B1(n6636), .B2(keyinput_f32), .C1(n6732), .C2(
        keyinput_f31), .A(n6635), .ZN(n6643) );
  INV_X1 U7574 ( .A(DATAI_29_), .ZN(n6638) );
  AOI22_X1 U7575 ( .A1(n6697), .A2(keyinput_f19), .B1(n6638), .B2(keyinput_f2), 
        .ZN(n6637) );
  OAI221_X1 U7576 ( .B1(n6697), .B2(keyinput_f19), .C1(n6638), .C2(keyinput_f2), .A(n6637), .ZN(n6642) );
  INV_X1 U7577 ( .A(CODEFETCH_REG_SCAN_IN), .ZN(n6728) );
  AOI22_X1 U7578 ( .A1(n6728), .A2(keyinput_f39), .B1(n6640), .B2(keyinput_f62), .ZN(n6639) );
  OAI221_X1 U7579 ( .B1(n6728), .B2(keyinput_f39), .C1(n6640), .C2(
        keyinput_f62), .A(n6639), .ZN(n6641) );
  NOR4_X1 U7580 ( .A1(n6644), .A2(n6643), .A3(n6642), .A4(n6641), .ZN(n6645)
         );
  NAND4_X1 U7581 ( .A1(n6648), .A2(n6647), .A3(n6646), .A4(n6645), .ZN(n6690)
         );
  AOI22_X1 U7582 ( .A1(keyinput_f46), .A2(W_R_N_REG_SCAN_IN), .B1(
        REIP_REG_21__SCAN_IN), .B2(keyinput_f61), .ZN(n6649) );
  OAI221_X1 U7583 ( .B1(keyinput_f46), .B2(W_R_N_REG_SCAN_IN), .C1(
        REIP_REG_21__SCAN_IN), .C2(keyinput_f61), .A(n6649), .ZN(n6656) );
  AOI22_X1 U7584 ( .A1(DATAI_2_), .A2(keyinput_f29), .B1(REIP_REG_28__SCAN_IN), 
        .B2(keyinput_f54), .ZN(n6650) );
  OAI221_X1 U7585 ( .B1(DATAI_2_), .B2(keyinput_f29), .C1(REIP_REG_28__SCAN_IN), .C2(keyinput_f54), .A(n6650), .ZN(n6655) );
  AOI22_X1 U7586 ( .A1(REQUESTPENDING_REG_SCAN_IN), .A2(keyinput_f42), .B1(
        DATAI_9_), .B2(keyinput_f22), .ZN(n6651) );
  OAI221_X1 U7587 ( .B1(REQUESTPENDING_REG_SCAN_IN), .B2(keyinput_f42), .C1(
        DATAI_9_), .C2(keyinput_f22), .A(n6651), .ZN(n6654) );
  AOI22_X1 U7588 ( .A1(DATAI_20_), .A2(keyinput_f11), .B1(REIP_REG_30__SCAN_IN), .B2(keyinput_f52), .ZN(n6652) );
  OAI221_X1 U7589 ( .B1(DATAI_20_), .B2(keyinput_f11), .C1(
        REIP_REG_30__SCAN_IN), .C2(keyinput_f52), .A(n6652), .ZN(n6653) );
  NOR4_X1 U7590 ( .A1(n6656), .A2(n6655), .A3(n6654), .A4(n6653), .ZN(n6688)
         );
  XOR2_X1 U7591 ( .A(n6657), .B(keyinput_f43), .Z(n6664) );
  AOI22_X1 U7592 ( .A1(DATAI_31_), .A2(keyinput_f0), .B1(n6735), .B2(
        keyinput_f37), .ZN(n6658) );
  OAI221_X1 U7593 ( .B1(DATAI_31_), .B2(keyinput_f0), .C1(n6735), .C2(
        keyinput_f37), .A(n6658), .ZN(n6663) );
  AOI22_X1 U7594 ( .A1(DATAI_6_), .A2(keyinput_f25), .B1(REIP_REG_24__SCAN_IN), 
        .B2(keyinput_f58), .ZN(n6659) );
  OAI221_X1 U7595 ( .B1(DATAI_6_), .B2(keyinput_f25), .C1(REIP_REG_24__SCAN_IN), .C2(keyinput_f58), .A(n6659), .ZN(n6662) );
  AOI22_X1 U7596 ( .A1(DATAI_21_), .A2(keyinput_f10), .B1(DATAI_5_), .B2(
        keyinput_f26), .ZN(n6660) );
  OAI221_X1 U7597 ( .B1(DATAI_21_), .B2(keyinput_f10), .C1(DATAI_5_), .C2(
        keyinput_f26), .A(n6660), .ZN(n6661) );
  NOR4_X1 U7598 ( .A1(n6664), .A2(n6663), .A3(n6662), .A4(n6661), .ZN(n6687)
         );
  AOI22_X1 U7599 ( .A1(n6769), .A2(keyinput_f5), .B1(n6666), .B2(keyinput_f59), 
        .ZN(n6665) );
  OAI221_X1 U7600 ( .B1(n6769), .B2(keyinput_f5), .C1(n6666), .C2(keyinput_f59), .A(n6665), .ZN(n6675) );
  INV_X1 U7601 ( .A(DATAI_30_), .ZN(n6668) );
  INV_X1 U7602 ( .A(DATAI_18_), .ZN(n6716) );
  AOI22_X1 U7603 ( .A1(n6668), .A2(keyinput_f1), .B1(keyinput_f13), .B2(n6716), 
        .ZN(n6667) );
  OAI221_X1 U7604 ( .B1(n6668), .B2(keyinput_f1), .C1(n6716), .C2(keyinput_f13), .A(n6667), .ZN(n6674) );
  INV_X1 U7605 ( .A(DATAI_22_), .ZN(n6718) );
  AOI22_X1 U7606 ( .A1(n6696), .A2(keyinput_f45), .B1(n6718), .B2(keyinput_f9), 
        .ZN(n6669) );
  OAI221_X1 U7607 ( .B1(n6696), .B2(keyinput_f45), .C1(n6718), .C2(keyinput_f9), .A(n6669), .ZN(n6673) );
  INV_X1 U7608 ( .A(DATAI_25_), .ZN(n6746) );
  AOI22_X1 U7609 ( .A1(n6746), .A2(keyinput_f6), .B1(keyinput_f41), .B2(n6671), 
        .ZN(n6670) );
  OAI221_X1 U7610 ( .B1(n6746), .B2(keyinput_f6), .C1(n6671), .C2(keyinput_f41), .A(n6670), .ZN(n6672) );
  NOR4_X1 U7611 ( .A1(n6675), .A2(n6674), .A3(n6673), .A4(n6672), .ZN(n6686)
         );
  AOI22_X1 U7612 ( .A1(n6731), .A2(keyinput_f56), .B1(keyinput_f18), .B2(n6700), .ZN(n6676) );
  OAI221_X1 U7613 ( .B1(n6731), .B2(keyinput_f56), .C1(n6700), .C2(
        keyinput_f18), .A(n6676), .ZN(n6684) );
  INV_X1 U7614 ( .A(DATAI_27_), .ZN(n6678) );
  AOI22_X1 U7615 ( .A1(n6734), .A2(keyinput_f21), .B1(n6678), .B2(keyinput_f4), 
        .ZN(n6677) );
  OAI221_X1 U7616 ( .B1(n6734), .B2(keyinput_f21), .C1(n6678), .C2(keyinput_f4), .A(n6677), .ZN(n6683) );
  AOI22_X1 U7617 ( .A1(n6713), .A2(keyinput_f24), .B1(n6749), .B2(keyinput_f57), .ZN(n6679) );
  OAI221_X1 U7618 ( .B1(n6713), .B2(keyinput_f24), .C1(n6749), .C2(
        keyinput_f57), .A(n6679), .ZN(n6682) );
  INV_X1 U7619 ( .A(DATAI_23_), .ZN(n6712) );
  AOI22_X1 U7620 ( .A1(n6712), .A2(keyinput_f8), .B1(n6487), .B2(keyinput_f35), 
        .ZN(n6680) );
  OAI221_X1 U7621 ( .B1(n6712), .B2(keyinput_f8), .C1(n6487), .C2(keyinput_f35), .A(n6680), .ZN(n6681) );
  NOR4_X1 U7622 ( .A1(n6684), .A2(n6683), .A3(n6682), .A4(n6681), .ZN(n6685)
         );
  NAND4_X1 U7623 ( .A1(n6688), .A2(n6687), .A3(n6686), .A4(n6685), .ZN(n6689)
         );
  NOR4_X1 U7624 ( .A1(n6692), .A2(n6691), .A3(n6690), .A4(n6689), .ZN(n6693)
         );
  AOI221_X1 U7625 ( .B1(DATAI_3_), .B2(keyinput_f28), .C1(n6802), .C2(n6694), 
        .A(n6693), .ZN(n6801) );
  AOI22_X1 U7626 ( .A1(n6697), .A2(keyinput_g19), .B1(keyinput_g45), .B2(n6696), .ZN(n6695) );
  OAI221_X1 U7627 ( .B1(n6697), .B2(keyinput_g19), .C1(n6696), .C2(
        keyinput_g45), .A(n6695), .ZN(n6710) );
  AOI22_X1 U7628 ( .A1(n6700), .A2(keyinput_g18), .B1(keyinput_g20), .B2(n6699), .ZN(n6698) );
  OAI221_X1 U7629 ( .B1(n6700), .B2(keyinput_g18), .C1(n6699), .C2(
        keyinput_g20), .A(n6698), .ZN(n6709) );
  AOI22_X1 U7630 ( .A1(n6703), .A2(keyinput_g61), .B1(n6702), .B2(keyinput_g53), .ZN(n6701) );
  OAI221_X1 U7631 ( .B1(n6703), .B2(keyinput_g61), .C1(n6702), .C2(
        keyinput_g53), .A(n6701), .ZN(n6708) );
  AOI22_X1 U7632 ( .A1(n6706), .A2(keyinput_g63), .B1(keyinput_g16), .B2(n6705), .ZN(n6704) );
  OAI221_X1 U7633 ( .B1(n6706), .B2(keyinput_g63), .C1(n6705), .C2(
        keyinput_g16), .A(n6704), .ZN(n6707) );
  NOR4_X1 U7634 ( .A1(n6710), .A2(n6709), .A3(n6708), .A4(n6707), .ZN(n6760)
         );
  AOI22_X1 U7635 ( .A1(n6713), .A2(keyinput_g24), .B1(keyinput_g8), .B2(n6712), 
        .ZN(n6711) );
  OAI221_X1 U7636 ( .B1(n6713), .B2(keyinput_g24), .C1(n6712), .C2(keyinput_g8), .A(n6711), .ZN(n6726) );
  AOI22_X1 U7637 ( .A1(n6716), .A2(keyinput_g13), .B1(n6715), .B2(keyinput_g25), .ZN(n6714) );
  OAI221_X1 U7638 ( .B1(n6716), .B2(keyinput_g13), .C1(n6715), .C2(
        keyinput_g25), .A(n6714), .ZN(n6725) );
  AOI22_X1 U7639 ( .A1(n6719), .A2(keyinput_g26), .B1(n6718), .B2(keyinput_g9), 
        .ZN(n6717) );
  OAI221_X1 U7640 ( .B1(n6719), .B2(keyinput_g26), .C1(n6718), .C2(keyinput_g9), .A(n6717), .ZN(n6724) );
  AOI22_X1 U7641 ( .A1(n6722), .A2(keyinput_g3), .B1(keyinput_g27), .B2(n6721), 
        .ZN(n6720) );
  OAI221_X1 U7642 ( .B1(n6722), .B2(keyinput_g3), .C1(n6721), .C2(keyinput_g27), .A(n6720), .ZN(n6723) );
  NOR4_X1 U7643 ( .A1(n6726), .A2(n6725), .A3(n6724), .A4(n6723), .ZN(n6759)
         );
  AOI22_X1 U7644 ( .A1(n6729), .A2(keyinput_g29), .B1(keyinput_g39), .B2(n6728), .ZN(n6727) );
  OAI221_X1 U7645 ( .B1(n6729), .B2(keyinput_g29), .C1(n6728), .C2(
        keyinput_g39), .A(n6727), .ZN(n6742) );
  AOI22_X1 U7646 ( .A1(n6732), .A2(keyinput_g31), .B1(n6731), .B2(keyinput_g56), .ZN(n6730) );
  OAI221_X1 U7647 ( .B1(n6732), .B2(keyinput_g31), .C1(n6731), .C2(
        keyinput_g56), .A(n6730), .ZN(n6741) );
  AOI22_X1 U7648 ( .A1(n6735), .A2(keyinput_g37), .B1(n6734), .B2(keyinput_g21), .ZN(n6733) );
  OAI221_X1 U7649 ( .B1(n6735), .B2(keyinput_g37), .C1(n6734), .C2(
        keyinput_g21), .A(n6733), .ZN(n6740) );
  AOI22_X1 U7650 ( .A1(n6738), .A2(keyinput_g7), .B1(keyinput_g30), .B2(n6737), 
        .ZN(n6736) );
  OAI221_X1 U7651 ( .B1(n6738), .B2(keyinput_g7), .C1(n6737), .C2(keyinput_g30), .A(n6736), .ZN(n6739) );
  NOR4_X1 U7652 ( .A1(n6742), .A2(n6741), .A3(n6740), .A4(n6739), .ZN(n6758)
         );
  AOI22_X1 U7653 ( .A1(n6744), .A2(keyinput_g0), .B1(n6487), .B2(keyinput_g35), 
        .ZN(n6743) );
  OAI221_X1 U7654 ( .B1(n6744), .B2(keyinput_g0), .C1(n6487), .C2(keyinput_g35), .A(n6743), .ZN(n6756) );
  AOI22_X1 U7655 ( .A1(n4307), .A2(keyinput_g52), .B1(keyinput_g6), .B2(n6746), 
        .ZN(n6745) );
  OAI221_X1 U7656 ( .B1(n4307), .B2(keyinput_g52), .C1(n6746), .C2(keyinput_g6), .A(n6745), .ZN(n6755) );
  AOI22_X1 U7657 ( .A1(n6749), .A2(keyinput_g57), .B1(keyinput_g48), .B2(n6748), .ZN(n6747) );
  OAI221_X1 U7658 ( .B1(n6749), .B2(keyinput_g57), .C1(n6748), .C2(
        keyinput_g48), .A(n6747), .ZN(n6754) );
  INV_X1 U7659 ( .A(DATAI_21_), .ZN(n6752) );
  AOI22_X1 U7660 ( .A1(n6752), .A2(keyinput_g10), .B1(keyinput_g38), .B2(n6751), .ZN(n6750) );
  OAI221_X1 U7661 ( .B1(n6752), .B2(keyinput_g10), .C1(n6751), .C2(
        keyinput_g38), .A(n6750), .ZN(n6753) );
  NOR4_X1 U7662 ( .A1(n6756), .A2(n6755), .A3(n6754), .A4(n6753), .ZN(n6757)
         );
  NAND4_X1 U7663 ( .A1(n6760), .A2(n6759), .A3(n6758), .A4(n6757), .ZN(n6799)
         );
  AOI22_X1 U7664 ( .A1(DATAI_20_), .A2(keyinput_g11), .B1(DATAI_8_), .B2(
        keyinput_g23), .ZN(n6761) );
  OAI221_X1 U7665 ( .B1(DATAI_20_), .B2(keyinput_g11), .C1(DATAI_8_), .C2(
        keyinput_g23), .A(n6761), .ZN(n6768) );
  AOI22_X1 U7666 ( .A1(REQUESTPENDING_REG_SCAN_IN), .A2(keyinput_g42), .B1(
        REIP_REG_31__SCAN_IN), .B2(keyinput_g51), .ZN(n6762) );
  OAI221_X1 U7667 ( .B1(REQUESTPENDING_REG_SCAN_IN), .B2(keyinput_g42), .C1(
        REIP_REG_31__SCAN_IN), .C2(keyinput_g51), .A(n6762), .ZN(n6767) );
  AOI22_X1 U7668 ( .A1(BS16_N), .A2(keyinput_g34), .B1(DATAI_19_), .B2(
        keyinput_g12), .ZN(n6763) );
  OAI221_X1 U7669 ( .B1(BS16_N), .B2(keyinput_g34), .C1(DATAI_19_), .C2(
        keyinput_g12), .A(n6763), .ZN(n6766) );
  AOI22_X1 U7670 ( .A1(W_R_N_REG_SCAN_IN), .A2(keyinput_g46), .B1(
        REIP_REG_27__SCAN_IN), .B2(keyinput_g55), .ZN(n6764) );
  OAI221_X1 U7671 ( .B1(W_R_N_REG_SCAN_IN), .B2(keyinput_g46), .C1(
        REIP_REG_27__SCAN_IN), .C2(keyinput_g55), .A(n6764), .ZN(n6765) );
  NOR4_X1 U7672 ( .A1(n6768), .A2(n6767), .A3(n6766), .A4(n6765), .ZN(n6797)
         );
  XOR2_X1 U7673 ( .A(n6769), .B(keyinput_g5), .Z(n6777) );
  AOI22_X1 U7674 ( .A1(HOLD), .A2(keyinput_g36), .B1(n6771), .B2(keyinput_g54), 
        .ZN(n6770) );
  OAI221_X1 U7675 ( .B1(HOLD), .B2(keyinput_g36), .C1(n6771), .C2(keyinput_g54), .A(n6770), .ZN(n6776) );
  AOI22_X1 U7676 ( .A1(D_C_N_REG_SCAN_IN), .A2(keyinput_g41), .B1(DATAI_16_), 
        .B2(keyinput_g15), .ZN(n6772) );
  OAI221_X1 U7677 ( .B1(D_C_N_REG_SCAN_IN), .B2(keyinput_g41), .C1(DATAI_16_), 
        .C2(keyinput_g15), .A(n6772), .ZN(n6775) );
  AOI22_X1 U7678 ( .A1(BYTEENABLE_REG_3__SCAN_IN), .A2(keyinput_g50), .B1(
        DATAI_27_), .B2(keyinput_g4), .ZN(n6773) );
  OAI221_X1 U7679 ( .B1(BYTEENABLE_REG_3__SCAN_IN), .B2(keyinput_g50), .C1(
        DATAI_27_), .C2(keyinput_g4), .A(n6773), .ZN(n6774) );
  NOR4_X1 U7680 ( .A1(n6777), .A2(n6776), .A3(n6775), .A4(n6774), .ZN(n6796)
         );
  AOI22_X1 U7681 ( .A1(DATAI_9_), .A2(keyinput_g22), .B1(STATEBS16_REG_SCAN_IN), .B2(keyinput_g43), .ZN(n6778) );
  OAI221_X1 U7682 ( .B1(DATAI_9_), .B2(keyinput_g22), .C1(
        STATEBS16_REG_SCAN_IN), .C2(keyinput_g43), .A(n6778), .ZN(n6785) );
  AOI22_X1 U7683 ( .A1(BYTEENABLE_REG_0__SCAN_IN), .A2(keyinput_g47), .B1(
        REIP_REG_24__SCAN_IN), .B2(keyinput_g58), .ZN(n6779) );
  OAI221_X1 U7684 ( .B1(BYTEENABLE_REG_0__SCAN_IN), .B2(keyinput_g47), .C1(
        REIP_REG_24__SCAN_IN), .C2(keyinput_g58), .A(n6779), .ZN(n6784) );
  AOI22_X1 U7685 ( .A1(NA_N), .A2(keyinput_g33), .B1(M_IO_N_REG_SCAN_IN), .B2(
        keyinput_g40), .ZN(n6780) );
  OAI221_X1 U7686 ( .B1(NA_N), .B2(keyinput_g33), .C1(M_IO_N_REG_SCAN_IN), 
        .C2(keyinput_g40), .A(n6780), .ZN(n6783) );
  AOI22_X1 U7687 ( .A1(BYTEENABLE_REG_2__SCAN_IN), .A2(keyinput_g49), .B1(
        DATAI_14_), .B2(keyinput_g17), .ZN(n6781) );
  OAI221_X1 U7688 ( .B1(BYTEENABLE_REG_2__SCAN_IN), .B2(keyinput_g49), .C1(
        DATAI_14_), .C2(keyinput_g17), .A(n6781), .ZN(n6782) );
  NOR4_X1 U7689 ( .A1(n6785), .A2(n6784), .A3(n6783), .A4(n6782), .ZN(n6795)
         );
  AOI22_X1 U7690 ( .A1(DATAI_17_), .A2(keyinput_g14), .B1(REIP_REG_22__SCAN_IN), .B2(keyinput_g60), .ZN(n6786) );
  OAI221_X1 U7691 ( .B1(DATAI_17_), .B2(keyinput_g14), .C1(
        REIP_REG_22__SCAN_IN), .C2(keyinput_g60), .A(n6786), .ZN(n6793) );
  AOI22_X1 U7692 ( .A1(DATAI_29_), .A2(keyinput_g2), .B1(DATAI_30_), .B2(
        keyinput_g1), .ZN(n6787) );
  OAI221_X1 U7693 ( .B1(DATAI_29_), .B2(keyinput_g2), .C1(DATAI_30_), .C2(
        keyinput_g1), .A(n6787), .ZN(n6792) );
  AOI22_X1 U7694 ( .A1(REIP_REG_20__SCAN_IN), .A2(keyinput_g62), .B1(
        REIP_REG_23__SCAN_IN), .B2(keyinput_g59), .ZN(n6788) );
  OAI221_X1 U7695 ( .B1(REIP_REG_20__SCAN_IN), .B2(keyinput_g62), .C1(
        REIP_REG_23__SCAN_IN), .C2(keyinput_g59), .A(n6788), .ZN(n6791) );
  AOI22_X1 U7696 ( .A1(MEMORYFETCH_REG_SCAN_IN), .A2(keyinput_g32), .B1(
        MORE_REG_SCAN_IN), .B2(keyinput_g44), .ZN(n6789) );
  OAI221_X1 U7697 ( .B1(MEMORYFETCH_REG_SCAN_IN), .B2(keyinput_g32), .C1(
        MORE_REG_SCAN_IN), .C2(keyinput_g44), .A(n6789), .ZN(n6790) );
  NOR4_X1 U7698 ( .A1(n6793), .A2(n6792), .A3(n6791), .A4(n6790), .ZN(n6794)
         );
  NAND4_X1 U7699 ( .A1(n6797), .A2(n6796), .A3(n6795), .A4(n6794), .ZN(n6798)
         );
  OAI22_X1 U7700 ( .A1(keyinput_g28), .A2(n6802), .B1(n6799), .B2(n6798), .ZN(
        n6800) );
  AOI211_X1 U7701 ( .C1(keyinput_g28), .C2(n6802), .A(n6801), .B(n6800), .ZN(
        n6806) );
  AOI22_X1 U7702 ( .A1(n6804), .A2(BYTEENABLE_REG_3__SCAN_IN), .B1(
        BE_N_REG_3__SCAN_IN), .B2(n6803), .ZN(n6805) );
  XNOR2_X1 U7703 ( .A(n6806), .B(n6805), .ZN(U3445) );
  CLKBUF_X1 U34480 ( .A(n3254), .Z(n2992) );
  CLKBUF_X1 U3438 ( .A(n3324), .Z(n3232) );
  CLKBUF_X1 U34550 ( .A(n3115), .Z(n3207) );
  XNOR2_X1 U34720 ( .A(n3209), .B(n3208), .ZN(n3274) );
  CLKBUF_X1 U3481 ( .A(n4247), .Z(n4248) );
  CLKBUF_X1 U3523 ( .A(n3135), .Z(n3554) );
  OR2_X2 U3531 ( .A1(n3113), .A2(n3112), .ZN(n4181) );
  XNOR2_X1 U3553 ( .A(n4158), .B(n4157), .ZN(n5538) );
endmodule

