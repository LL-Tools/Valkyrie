

module b14_C_lock ( keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, 
        keyinput_5, keyinput_6, keyinput_7, keyinput_8, keyinput_9, 
        keyinput_10, keyinput_11, keyinput_12, keyinput_13, keyinput_14, 
        keyinput_15, keyinput_16, keyinput_17, keyinput_18, keyinput_19, 
        keyinput_20, keyinput_21, keyinput_22, keyinput_23, keyinput_24, 
        keyinput_25, keyinput_26, keyinput_27, keyinput_28, keyinput_29, 
        keyinput_30, keyinput_31, keyinput_32, keyinput_33, keyinput_34, 
        keyinput_35, keyinput_36, keyinput_37, keyinput_38, keyinput_39, 
        keyinput_40, keyinput_41, keyinput_42, keyinput_43, keyinput_44, 
        keyinput_45, keyinput_46, keyinput_47, keyinput_48, keyinput_49, 
        keyinput_50, keyinput_51, keyinput_52, keyinput_53, keyinput_54, 
        keyinput_55, keyinput_56, keyinput_57, keyinput_58, keyinput_59, 
        keyinput_60, keyinput_61, keyinput_62, keyinput_63, keyinput_64, 
        keyinput_65, keyinput_66, keyinput_67, keyinput_68, keyinput_69, 
        keyinput_70, keyinput_71, keyinput_72, keyinput_73, keyinput_74, 
        keyinput_75, keyinput_76, keyinput_77, keyinput_78, keyinput_79, 
        keyinput_80, keyinput_81, keyinput_82, keyinput_83, keyinput_84, 
        keyinput_85, keyinput_86, keyinput_87, keyinput_88, keyinput_89, 
        keyinput_90, keyinput_91, keyinput_92, keyinput_93, keyinput_94, 
        keyinput_95, keyinput_96, keyinput_97, keyinput_98, keyinput_99, 
        keyinput_100, keyinput_101, keyinput_102, keyinput_103, keyinput_104, 
        keyinput_105, keyinput_106, keyinput_107, keyinput_108, keyinput_109, 
        keyinput_110, keyinput_111, keyinput_112, keyinput_113, keyinput_114, 
        keyinput_115, keyinput_116, keyinput_117, keyinput_118, keyinput_119, 
        keyinput_120, keyinput_121, keyinput_122, keyinput_123, keyinput_124, 
        keyinput_125, keyinput_126, keyinput_127, keyinput_128, keyinput_129, 
        keyinput_130, keyinput_131, keyinput_132, keyinput_133, keyinput_134, 
        keyinput_135, keyinput_136, keyinput_137, keyinput_138, keyinput_139, 
        keyinput_140, keyinput_141, keyinput_142, keyinput_143, keyinput_144, 
        keyinput_145, keyinput_146, keyinput_147, keyinput_148, keyinput_149, 
        keyinput_150, keyinput_151, keyinput_152, keyinput_153, keyinput_154, 
        keyinput_155, keyinput_156, keyinput_157, keyinput_158, keyinput_159, 
        keyinput_160, keyinput_161, keyinput_162, keyinput_163, keyinput_164, 
        keyinput_165, keyinput_166, keyinput_167, keyinput_168, keyinput_169, 
        keyinput_170, keyinput_171, keyinput_172, keyinput_173, keyinput_174, 
        keyinput_175, keyinput_176, keyinput_177, keyinput_178, keyinput_179, 
        keyinput_180, keyinput_181, keyinput_182, keyinput_183, keyinput_184, 
        keyinput_185, keyinput_186, keyinput_187, keyinput_188, keyinput_189, 
        keyinput_190, keyinput_191, keyinput_192, keyinput_193, keyinput_194, 
        keyinput_195, keyinput_196, keyinput_197, keyinput_198, keyinput_199, 
        keyinput_200, keyinput_201, keyinput_202, keyinput_203, keyinput_204, 
        keyinput_205, keyinput_206, keyinput_207, keyinput_208, keyinput_209, 
        keyinput_210, keyinput_211, keyinput_212, keyinput_213, keyinput_214, 
        keyinput_215, keyinput_216, keyinput_217, keyinput_218, keyinput_219, 
        keyinput_220, keyinput_221, keyinput_222, keyinput_223, keyinput_224, 
        keyinput_225, keyinput_226, keyinput_227, keyinput_228, keyinput_229, 
        keyinput_230, keyinput_231, keyinput_232, keyinput_233, keyinput_234, 
        keyinput_235, keyinput_236, keyinput_237, keyinput_238, keyinput_239, 
        keyinput_240, keyinput_241, keyinput_242, keyinput_243, keyinput_244, 
        keyinput_245, keyinput_246, keyinput_247, keyinput_248, keyinput_249, 
        keyinput_250, keyinput_251, keyinput_252, keyinput_253, keyinput_254, 
        keyinput_255, DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, 
        DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, 
        DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, 
        DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, 
        DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, 
        DATAI_1_, DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN, 
        REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN, 
        REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN, 
        REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN, 
        REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN, 
        REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN, 
        REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN, 
        REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN, 
        IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN, 
        IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN, 
        IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN, 
        IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN, 
        IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN, 
        IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN, 
        IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN, 
        IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN, 
        IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN, 
        IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN, 
        IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN, 
        D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN, D_REG_4__SCAN_IN, 
        D_REG_5__SCAN_IN, D_REG_6__SCAN_IN, D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, 
        D_REG_9__SCAN_IN, D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, 
        D_REG_12__SCAN_IN, D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, 
        D_REG_15__SCAN_IN, D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, 
        D_REG_18__SCAN_IN, D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, 
        D_REG_21__SCAN_IN, D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, 
        D_REG_24__SCAN_IN, D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, 
        D_REG_27__SCAN_IN, D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, 
        D_REG_30__SCAN_IN, D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, 
        REG0_REG_1__SCAN_IN, REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, 
        REG0_REG_4__SCAN_IN, REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, 
        REG0_REG_7__SCAN_IN, REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, 
        REG0_REG_10__SCAN_IN, REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, 
        REG0_REG_13__SCAN_IN, REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, 
        REG0_REG_16__SCAN_IN, REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, 
        REG0_REG_19__SCAN_IN, REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, 
        REG0_REG_22__SCAN_IN, REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, 
        REG0_REG_25__SCAN_IN, REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, 
        REG0_REG_28__SCAN_IN, REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, 
        REG0_REG_31__SCAN_IN, REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, 
        REG1_REG_2__SCAN_IN, REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, 
        REG1_REG_5__SCAN_IN, REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, 
        REG1_REG_8__SCAN_IN, REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, 
        REG1_REG_11__SCAN_IN, REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, 
        REG1_REG_14__SCAN_IN, REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, 
        REG1_REG_17__SCAN_IN, REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, 
        REG1_REG_20__SCAN_IN, REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, 
        REG1_REG_23__SCAN_IN, REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, 
        REG1_REG_26__SCAN_IN, REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, 
        REG1_REG_29__SCAN_IN, REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, 
        REG2_REG_0__SCAN_IN, REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, 
        REG2_REG_3__SCAN_IN, REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, 
        REG2_REG_6__SCAN_IN, REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, 
        REG2_REG_9__SCAN_IN, REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, 
        REG2_REG_12__SCAN_IN, REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, 
        REG2_REG_15__SCAN_IN, REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, 
        REG2_REG_18__SCAN_IN, REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, 
        REG2_REG_21__SCAN_IN, REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, 
        REG2_REG_24__SCAN_IN, REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, 
        REG2_REG_27__SCAN_IN, REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, 
        REG2_REG_30__SCAN_IN, REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, 
        ADDR_REG_18__SCAN_IN, ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, 
        ADDR_REG_15__SCAN_IN, ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, 
        ADDR_REG_12__SCAN_IN, ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, 
        ADDR_REG_9__SCAN_IN, ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, 
        ADDR_REG_6__SCAN_IN, ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, 
        ADDR_REG_3__SCAN_IN, ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, 
        ADDR_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        B_REG_SCAN_IN, REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, 
        REG3_REG_6__SCAN_IN, REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, 
        REG3_REG_11__SCAN_IN, REG3_REG_22__SCAN_IN, U3352, U3351, U3350, U3349, 
        U3348, U3347, U3346, U3345, U3344, U3343, U3342, U3341, U3340, U3339, 
        U3338, U3337, U3336, U3335, U3334, U3333, U3332, U3331, U3330, U3329, 
        U3328, U3327, U3326, U3325, U3324, U3323, U3322, U3321, U3458, U3459, 
        U3320, U3319, U3318, U3317, U3316, U3315, U3314, U3313, U3312, U3311, 
        U3310, U3309, U3308, U3307, U3306, U3305, U3304, U3303, U3302, U3301, 
        U3300, U3299, U3298, U3297, U3296, U3295, U3294, U3293, U3292, U3291, 
        U3467, U3469, U3471, U3473, U3475, U3477, U3479, U3481, U3483, U3485, 
        U3487, U3489, U3491, U3493, U3495, U3497, U3499, U3501, U3503, U3505, 
        U3506, U3507, U3508, U3509, U3510, U3511, U3512, U3513, U3514, U3515, 
        U3516, U3517, U3518, U3519, U3520, U3521, U3522, U3523, U3524, U3525, 
        U3526, U3527, U3528, U3529, U3530, U3531, U3532, U3533, U3534, U3535, 
        U3536, U3537, U3538, U3539, U3540, U3541, U3542, U3543, U3544, U3545, 
        U3546, U3547, U3548, U3549, U3290, U3289, U3288, U3287, U3286, U3285, 
        U3284, U3283, U3282, U3281, U3280, U3279, U3278, U3277, U3276, U3275, 
        U3274, U3273, U3272, U3271, U3270, U3269, U3268, U3267, U3266, U3265, 
        U3264, U3263, U3262, U3354, U3261, U3260, U3259, U3258, U3257, U3256, 
        U3255, U3254, U3253, U3252, U3251, U3250, U3249, U3248, U3247, U3246, 
        U3245, U3244, U3243, U3242, U3241, U3240, U3550, U3551, U3552, U3553, 
        U3554, U3555, U3556, U3557, U3558, U3559, U3560, U3561, U3562, U3563, 
        U3564, U3565, U3566, U3567, U3568, U3569, U3570, U3571, U3572, U3573, 
        U3574, U3575, U3576, U3577, U3578, U3579, U3580, U3581, U3239, U3238, 
        U3237, U3236, U3235, U3234, U3233, U3232, U3231, U3230, U3229, U3228, 
        U3227, U3226, U3225, U3224, U3223, U3222, U3221, U3220, U3219, U3218, 
        U3217, U3216, U3215, U3214, U3213, U3212, U3211, U3210, U3149, U3148, 
        U4043 );
  input keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, keyinput_5,
         keyinput_6, keyinput_7, keyinput_8, keyinput_9, keyinput_10,
         keyinput_11, keyinput_12, keyinput_13, keyinput_14, keyinput_15,
         keyinput_16, keyinput_17, keyinput_18, keyinput_19, keyinput_20,
         keyinput_21, keyinput_22, keyinput_23, keyinput_24, keyinput_25,
         keyinput_26, keyinput_27, keyinput_28, keyinput_29, keyinput_30,
         keyinput_31, keyinput_32, keyinput_33, keyinput_34, keyinput_35,
         keyinput_36, keyinput_37, keyinput_38, keyinput_39, keyinput_40,
         keyinput_41, keyinput_42, keyinput_43, keyinput_44, keyinput_45,
         keyinput_46, keyinput_47, keyinput_48, keyinput_49, keyinput_50,
         keyinput_51, keyinput_52, keyinput_53, keyinput_54, keyinput_55,
         keyinput_56, keyinput_57, keyinput_58, keyinput_59, keyinput_60,
         keyinput_61, keyinput_62, keyinput_63, keyinput_64, keyinput_65,
         keyinput_66, keyinput_67, keyinput_68, keyinput_69, keyinput_70,
         keyinput_71, keyinput_72, keyinput_73, keyinput_74, keyinput_75,
         keyinput_76, keyinput_77, keyinput_78, keyinput_79, keyinput_80,
         keyinput_81, keyinput_82, keyinput_83, keyinput_84, keyinput_85,
         keyinput_86, keyinput_87, keyinput_88, keyinput_89, keyinput_90,
         keyinput_91, keyinput_92, keyinput_93, keyinput_94, keyinput_95,
         keyinput_96, keyinput_97, keyinput_98, keyinput_99, keyinput_100,
         keyinput_101, keyinput_102, keyinput_103, keyinput_104, keyinput_105,
         keyinput_106, keyinput_107, keyinput_108, keyinput_109, keyinput_110,
         keyinput_111, keyinput_112, keyinput_113, keyinput_114, keyinput_115,
         keyinput_116, keyinput_117, keyinput_118, keyinput_119, keyinput_120,
         keyinput_121, keyinput_122, keyinput_123, keyinput_124, keyinput_125,
         keyinput_126, keyinput_127, keyinput_128, keyinput_129, keyinput_130,
         keyinput_131, keyinput_132, keyinput_133, keyinput_134, keyinput_135,
         keyinput_136, keyinput_137, keyinput_138, keyinput_139, keyinput_140,
         keyinput_141, keyinput_142, keyinput_143, keyinput_144, keyinput_145,
         keyinput_146, keyinput_147, keyinput_148, keyinput_149, keyinput_150,
         keyinput_151, keyinput_152, keyinput_153, keyinput_154, keyinput_155,
         keyinput_156, keyinput_157, keyinput_158, keyinput_159, keyinput_160,
         keyinput_161, keyinput_162, keyinput_163, keyinput_164, keyinput_165,
         keyinput_166, keyinput_167, keyinput_168, keyinput_169, keyinput_170,
         keyinput_171, keyinput_172, keyinput_173, keyinput_174, keyinput_175,
         keyinput_176, keyinput_177, keyinput_178, keyinput_179, keyinput_180,
         keyinput_181, keyinput_182, keyinput_183, keyinput_184, keyinput_185,
         keyinput_186, keyinput_187, keyinput_188, keyinput_189, keyinput_190,
         keyinput_191, keyinput_192, keyinput_193, keyinput_194, keyinput_195,
         keyinput_196, keyinput_197, keyinput_198, keyinput_199, keyinput_200,
         keyinput_201, keyinput_202, keyinput_203, keyinput_204, keyinput_205,
         keyinput_206, keyinput_207, keyinput_208, keyinput_209, keyinput_210,
         keyinput_211, keyinput_212, keyinput_213, keyinput_214, keyinput_215,
         keyinput_216, keyinput_217, keyinput_218, keyinput_219, keyinput_220,
         keyinput_221, keyinput_222, keyinput_223, keyinput_224, keyinput_225,
         keyinput_226, keyinput_227, keyinput_228, keyinput_229, keyinput_230,
         keyinput_231, keyinput_232, keyinput_233, keyinput_234, keyinput_235,
         keyinput_236, keyinput_237, keyinput_238, keyinput_239, keyinput_240,
         keyinput_241, keyinput_242, keyinput_243, keyinput_244, keyinput_245,
         keyinput_246, keyinput_247, keyinput_248, keyinput_249, keyinput_250,
         keyinput_251, keyinput_252, keyinput_253, keyinput_254, keyinput_255,
         DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN,
         REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN,
         REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN,
         REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN,
         REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN,
         REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN,
         REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN,
         REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN,
         IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN,
         IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN,
         IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN,
         IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN,
         IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN,
         IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN,
         IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN,
         IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN,
         IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN,
         IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN,
         IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN,
         D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN,
         D_REG_4__SCAN_IN, D_REG_5__SCAN_IN, D_REG_6__SCAN_IN,
         D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, D_REG_9__SCAN_IN,
         D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, D_REG_12__SCAN_IN,
         D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, D_REG_15__SCAN_IN,
         D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, D_REG_18__SCAN_IN,
         D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, D_REG_21__SCAN_IN,
         D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, D_REG_24__SCAN_IN,
         D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, D_REG_27__SCAN_IN,
         D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, D_REG_30__SCAN_IN,
         D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, REG0_REG_1__SCAN_IN,
         REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, REG0_REG_4__SCAN_IN,
         REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, REG0_REG_7__SCAN_IN,
         REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, REG0_REG_10__SCAN_IN,
         REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, REG0_REG_13__SCAN_IN,
         REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, REG0_REG_16__SCAN_IN,
         REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, REG0_REG_19__SCAN_IN,
         REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, REG0_REG_22__SCAN_IN,
         REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, REG0_REG_25__SCAN_IN,
         REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, REG0_REG_28__SCAN_IN,
         REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, REG0_REG_31__SCAN_IN,
         REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, REG1_REG_2__SCAN_IN,
         REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, REG1_REG_5__SCAN_IN,
         REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, REG1_REG_8__SCAN_IN,
         REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, REG1_REG_11__SCAN_IN,
         REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, REG1_REG_14__SCAN_IN,
         REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, REG1_REG_17__SCAN_IN,
         REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, REG1_REG_20__SCAN_IN,
         REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, REG1_REG_23__SCAN_IN,
         REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, REG1_REG_26__SCAN_IN,
         REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, REG1_REG_29__SCAN_IN,
         REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, REG2_REG_0__SCAN_IN,
         REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, REG2_REG_3__SCAN_IN,
         REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, REG2_REG_6__SCAN_IN,
         REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, REG2_REG_9__SCAN_IN,
         REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, REG2_REG_12__SCAN_IN,
         REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, REG2_REG_15__SCAN_IN,
         REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, REG2_REG_18__SCAN_IN,
         REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, REG2_REG_21__SCAN_IN,
         REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, REG2_REG_24__SCAN_IN,
         REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, REG2_REG_27__SCAN_IN,
         REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, REG2_REG_30__SCAN_IN,
         REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, ADDR_REG_18__SCAN_IN,
         ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, ADDR_REG_15__SCAN_IN,
         ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, ADDR_REG_12__SCAN_IN,
         ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, ADDR_REG_9__SCAN_IN,
         ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, ADDR_REG_6__SCAN_IN,
         ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, ADDR_REG_3__SCAN_IN,
         ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, ADDR_REG_0__SCAN_IN,
         DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, DATAO_REG_2__SCAN_IN,
         DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, DATAO_REG_5__SCAN_IN,
         DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, DATAO_REG_8__SCAN_IN,
         DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, DATAO_REG_11__SCAN_IN,
         DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, DATAO_REG_14__SCAN_IN,
         DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, DATAO_REG_17__SCAN_IN,
         DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, DATAO_REG_20__SCAN_IN,
         DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, DATAO_REG_23__SCAN_IN,
         DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, DATAO_REG_26__SCAN_IN,
         DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, DATAO_REG_29__SCAN_IN,
         DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, B_REG_SCAN_IN,
         REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, REG3_REG_6__SCAN_IN,
         REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, REG3_REG_11__SCAN_IN,
         REG3_REG_22__SCAN_IN;
  output U3352, U3351, U3350, U3349, U3348, U3347, U3346, U3345, U3344, U3343,
         U3342, U3341, U3340, U3339, U3338, U3337, U3336, U3335, U3334, U3333,
         U3332, U3331, U3330, U3329, U3328, U3327, U3326, U3325, U3324, U3323,
         U3322, U3321, U3458, U3459, U3320, U3319, U3318, U3317, U3316, U3315,
         U3314, U3313, U3312, U3311, U3310, U3309, U3308, U3307, U3306, U3305,
         U3304, U3303, U3302, U3301, U3300, U3299, U3298, U3297, U3296, U3295,
         U3294, U3293, U3292, U3291, U3467, U3469, U3471, U3473, U3475, U3477,
         U3479, U3481, U3483, U3485, U3487, U3489, U3491, U3493, U3495, U3497,
         U3499, U3501, U3503, U3505, U3506, U3507, U3508, U3509, U3510, U3511,
         U3512, U3513, U3514, U3515, U3516, U3517, U3518, U3519, U3520, U3521,
         U3522, U3523, U3524, U3525, U3526, U3527, U3528, U3529, U3530, U3531,
         U3532, U3533, U3534, U3535, U3536, U3537, U3538, U3539, U3540, U3541,
         U3542, U3543, U3544, U3545, U3546, U3547, U3548, U3549, U3290, U3289,
         U3288, U3287, U3286, U3285, U3284, U3283, U3282, U3281, U3280, U3279,
         U3278, U3277, U3276, U3275, U3274, U3273, U3272, U3271, U3270, U3269,
         U3268, U3267, U3266, U3265, U3264, U3263, U3262, U3354, U3261, U3260,
         U3259, U3258, U3257, U3256, U3255, U3254, U3253, U3252, U3251, U3250,
         U3249, U3248, U3247, U3246, U3245, U3244, U3243, U3242, U3241, U3240,
         U3550, U3551, U3552, U3553, U3554, U3555, U3556, U3557, U3558, U3559,
         U3560, U3561, U3562, U3563, U3564, U3565, U3566, U3567, U3568, U3569,
         U3570, U3571, U3572, U3573, U3574, U3575, U3576, U3577, U3578, U3579,
         U3580, U3581, U3239, U3238, U3237, U3236, U3235, U3234, U3233, U3232,
         U3231, U3230, U3229, U3228, U3227, U3226, U3225, U3224, U3223, U3222,
         U3221, U3220, U3219, U3218, U3217, U3216, U3215, U3214, U3213, U3212,
         U3211, U3210, U3149, U3148, U4043;
  wire   n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519,
         n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529,
         n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539,
         n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549,
         n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559,
         n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569,
         n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579,
         n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589,
         n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599,
         n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609,
         n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619,
         n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629,
         n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639,
         n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649,
         n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659,
         n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669,
         n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679,
         n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689,
         n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699,
         n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709,
         n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719,
         n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729,
         n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739,
         n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749,
         n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759,
         n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769,
         n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779,
         n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789,
         n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799,
         n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809,
         n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819,
         n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829,
         n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839,
         n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849,
         n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859,
         n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869,
         n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879,
         n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889,
         n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899,
         n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909,
         n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919,
         n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929,
         n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939,
         n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949,
         n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959,
         n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969,
         n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979,
         n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989,
         n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999,
         n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009,
         n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019,
         n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029,
         n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039,
         n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049,
         n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059,
         n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069,
         n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079,
         n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089,
         n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099,
         n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109,
         n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119,
         n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129,
         n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139,
         n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149,
         n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159,
         n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169,
         n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179,
         n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189,
         n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199,
         n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209,
         n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219,
         n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229,
         n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239,
         n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249,
         n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259,
         n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269,
         n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279,
         n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289,
         n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299,
         n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309,
         n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319,
         n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329,
         n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339,
         n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349,
         n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359,
         n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369,
         n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379,
         n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389,
         n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399,
         n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409,
         n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419,
         n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429,
         n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439,
         n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449,
         n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459,
         n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469,
         n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479,
         n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489,
         n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499,
         n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509,
         n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519,
         n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529,
         n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539,
         n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549,
         n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559,
         n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569,
         n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579,
         n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589,
         n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599,
         n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609,
         n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619,
         n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629,
         n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639,
         n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649,
         n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659,
         n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669,
         n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679,
         n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689,
         n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699,
         n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709,
         n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719,
         n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729,
         n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739,
         n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749,
         n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759,
         n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769,
         n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779,
         n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789,
         n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799,
         n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809,
         n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819,
         n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829,
         n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839,
         n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849,
         n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859,
         n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869,
         n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879,
         n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889,
         n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899,
         n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909,
         n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919,
         n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929,
         n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939,
         n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949,
         n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959,
         n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969,
         n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979,
         n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989,
         n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999,
         n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009,
         n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019,
         n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029,
         n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039,
         n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049,
         n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059,
         n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069,
         n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079,
         n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089,
         n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099,
         n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109,
         n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119,
         n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129,
         n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139,
         n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149,
         n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159,
         n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169,
         n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179,
         n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189,
         n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199,
         n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209,
         n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219,
         n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229,
         n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239,
         n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249,
         n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259,
         n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269,
         n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279,
         n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289,
         n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299,
         n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309,
         n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319,
         n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329,
         n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339,
         n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349,
         n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359,
         n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369,
         n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379,
         n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389,
         n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399,
         n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409,
         n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419,
         n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429,
         n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439,
         n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449,
         n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459,
         n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469,
         n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479,
         n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489,
         n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499,
         n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509,
         n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519,
         n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529,
         n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539,
         n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549,
         n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559,
         n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569,
         n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579,
         n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589,
         n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599,
         n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609,
         n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619,
         n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629,
         n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639,
         n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649,
         n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659,
         n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669,
         n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679,
         n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689,
         n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699,
         n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709,
         n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719,
         n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729,
         n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739,
         n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749,
         n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759,
         n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769,
         n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779,
         n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789,
         n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799,
         n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809,
         n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819,
         n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829,
         n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839,
         n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849,
         n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859,
         n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869,
         n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879,
         n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889,
         n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899,
         n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909,
         n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919,
         n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929,
         n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939,
         n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949,
         n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959,
         n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969,
         n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979,
         n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989,
         n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999,
         n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009,
         n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019,
         n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029,
         n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039,
         n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049,
         n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059,
         n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069,
         n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079,
         n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089,
         n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099,
         n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109,
         n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119,
         n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129,
         n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139,
         n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149,
         n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159,
         n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169,
         n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179,
         n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189,
         n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199,
         n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209,
         n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219,
         n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229,
         n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239,
         n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249,
         n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259,
         n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269,
         n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279,
         n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289,
         n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299,
         n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309,
         n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319,
         n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329,
         n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339,
         n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349,
         n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359,
         n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369,
         n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379,
         n5380, n5381;

  INV_X1 U2545 ( .A(n3829), .ZN(n3782) );
  CLKBUF_X2 U2546 ( .A(n3054), .Z(n3835) );
  INV_X1 U2547 ( .A(n3740), .ZN(n3798) );
  INV_X1 U2548 ( .A(n3814), .ZN(n3740) );
  NOR2_X1 U2549 ( .A1(n3069), .A2(n2782), .ZN(n2785) );
  NAND2_X1 U2550 ( .A1(n3912), .A2(n3654), .ZN(n3913) );
  AOI21_X1 U2552 ( .B1(n3913), .B2(n3663), .A(n2753), .ZN(n5346) );
  CLKBUF_X3 U2553 ( .A(n3107), .Z(n4064) );
  NAND2_X1 U2554 ( .A1(n3866), .A2(n3758), .ZN(n3869) );
  AND4_X1 U2555 ( .A1(n3059), .A2(n3058), .A3(n3057), .A4(n3056), .ZN(n5133)
         );
  NAND2_X1 U2556 ( .A1(n3023), .A2(n2999), .ZN(n5333) );
  INV_X2 U2557 ( .A(IR_REG_31__SCAN_IN), .ZN(n2871) );
  NAND2_X1 U2558 ( .A1(n3023), .A2(n4921), .ZN(n3209) );
  OR2_X1 U2559 ( .A1(n3023), .A2(n5106), .ZN(n5266) );
  NAND2_X2 U2560 ( .A1(n2525), .A2(n2690), .ZN(n3023) );
  BUF_X1 U2561 ( .A(n4470), .Z(n2510) );
  AND2_X1 U2562 ( .A1(n3003), .A2(n3002), .ZN(n3051) );
  NAND2_X1 U2563 ( .A1(n2998), .A2(n3129), .ZN(n3814) );
  AOI21_X2 U2564 ( .B1(n5047), .B2(n5046), .A(n2839), .ZN(n2938) );
  INV_X1 U2565 ( .A(n3110), .ZN(n3752) );
  INV_X1 U2566 ( .A(n4163), .ZN(n3251) );
  XNOR2_X1 U2567 ( .A(n2785), .B(n5154), .ZN(n5090) );
  XNOR2_X1 U2568 ( .A(n2987), .B(n4843), .ZN(n2989) );
  NOR2_X1 U2569 ( .A1(n2968), .A2(n2967), .ZN(n2986) );
  NAND2_X1 U2570 ( .A1(n2564), .A2(n2514), .ZN(n4260) );
  NAND2_X1 U2571 ( .A1(n3742), .A2(n3741), .ZN(n3866) );
  NAND2_X1 U2572 ( .A1(n2582), .A2(n2516), .ZN(n4326) );
  NOR2_X1 U2573 ( .A1(n5024), .A2(n2610), .ZN(n2822) );
  NAND2_X1 U2574 ( .A1(n3234), .A2(n3997), .ZN(n3274) );
  OR2_X1 U2575 ( .A1(n5006), .A2(n2803), .ZN(n2807) );
  AND2_X1 U2576 ( .A1(n2750), .A2(n3263), .ZN(n3166) );
  OR2_X1 U2577 ( .A1(n3161), .A2(n3160), .ZN(n3167) );
  INV_X1 U2578 ( .A(n3200), .ZN(n4084) );
  NOR2_X1 U2579 ( .A1(n3114), .A2(n3113), .ZN(n3345) );
  INV_X2 U2580 ( .A(n5380), .ZN(n2512) );
  CLKBUF_X1 U2581 ( .A(n3183), .Z(n5103) );
  BUF_X2 U2582 ( .A(n3110), .Z(n3800) );
  NAND2_X1 U2583 ( .A1(n3000), .A2(n5333), .ZN(n3110) );
  NAND4_X1 U2584 ( .A1(n3098), .A2(n3097), .A3(n3096), .A4(n3095), .ZN(n4163)
         );
  INV_X1 U2585 ( .A(n3108), .ZN(n3815) );
  NAND4_X1 U2586 ( .A1(n2996), .A2(n2995), .A3(n2994), .A4(n2993), .ZN(n4165)
         );
  INV_X2 U2587 ( .A(n3026), .ZN(n4052) );
  NAND2_X2 U2588 ( .A1(n3209), .A2(n3047), .ZN(n3829) );
  NAND2_X1 U2589 ( .A1(n2990), .A2(n4918), .ZN(n3054) );
  CLKBUF_X3 U2590 ( .A(n3094), .Z(n2513) );
  NAND2_X1 U2591 ( .A1(n5071), .A2(n2926), .ZN(n3107) );
  NAND2_X1 U2592 ( .A1(n2992), .A2(n2989), .ZN(n3094) );
  XNOR2_X1 U2593 ( .A(n2970), .B(n2969), .ZN(n2992) );
  NAND2_X1 U2594 ( .A1(n4916), .A2(IR_REG_31__SCAN_IN), .ZN(n2970) );
  NAND2_X1 U2595 ( .A1(n2865), .A2(IR_REG_31__SCAN_IN), .ZN(n2866) );
  OR2_X1 U2596 ( .A1(n2986), .A2(n2871), .ZN(n2987) );
  AND2_X1 U2597 ( .A1(n5030), .A2(REG1_REG_13__SCAN_IN), .ZN(n2610) );
  OR2_X1 U2598 ( .A1(n2966), .A2(IR_REG_28__SCAN_IN), .ZN(n2967) );
  AND2_X1 U2599 ( .A1(n2853), .A2(n2792), .ZN(n2747) );
  AND3_X1 U2600 ( .A1(n2765), .A2(n2768), .A3(n2767), .ZN(n4926) );
  AND2_X1 U2601 ( .A1(n2748), .A2(n2591), .ZN(n2590) );
  AND2_X1 U2602 ( .A1(n2799), .A2(n2756), .ZN(n2804) );
  NOR2_X2 U2603 ( .A1(IR_REG_0__SCAN_IN), .A2(IR_REG_1__SCAN_IN), .ZN(n2769)
         );
  INV_X1 U2604 ( .A(IR_REG_30__SCAN_IN), .ZN(n2969) );
  INV_X1 U2605 ( .A(IR_REG_2__SCAN_IN), .ZN(n4800) );
  INV_X1 U2606 ( .A(IR_REG_3__SCAN_IN), .ZN(n2778) );
  INV_X1 U2607 ( .A(IR_REG_4__SCAN_IN), .ZN(n4607) );
  INV_X1 U2608 ( .A(IR_REG_18__SCAN_IN), .ZN(n4628) );
  INV_X1 U2609 ( .A(IR_REG_17__SCAN_IN), .ZN(n4822) );
  NOR2_X1 U2610 ( .A1(IR_REG_12__SCAN_IN), .A2(IR_REG_11__SCAN_IN), .ZN(n2758)
         );
  NOR2_X1 U2611 ( .A1(IR_REG_8__SCAN_IN), .A2(IR_REG_7__SCAN_IN), .ZN(n2799)
         );
  INV_X1 U2612 ( .A(IR_REG_16__SCAN_IN), .ZN(n4623) );
  NAND2_X4 U2613 ( .A1(n3209), .A2(n3129), .ZN(n3108) );
  AND2_X1 U2614 ( .A1(n3846), .A2(n2671), .ZN(n2670) );
  NAND2_X1 U2615 ( .A1(n2537), .A2(n3803), .ZN(n2671) );
  NAND2_X1 U2616 ( .A1(n3517), .A2(n3516), .ZN(n2681) );
  NOR2_X1 U2617 ( .A1(n4172), .A2(n2916), .ZN(n2917) );
  AND2_X1 U2618 ( .A1(n4924), .A2(REG2_REG_15__SCAN_IN), .ZN(n2916) );
  INV_X1 U2619 ( .A(n2714), .ZN(n2713) );
  AOI21_X1 U2620 ( .B1(n2707), .B2(n2701), .A(n2706), .ZN(n2700) );
  AOI21_X1 U2621 ( .B1(n2707), .B2(n2704), .A(n3592), .ZN(n2703) );
  NOR2_X1 U2622 ( .A1(n2751), .A2(n5308), .ZN(n2704) );
  OAI21_X1 U2623 ( .B1(n3833), .B2(n2667), .A(n2664), .ZN(n2663) );
  NAND2_X1 U2624 ( .A1(n2667), .A2(n2665), .ZN(n2664) );
  NAND2_X1 U2625 ( .A1(n2669), .A2(n2666), .ZN(n2665) );
  INV_X1 U2626 ( .A(n5241), .ZN(n2682) );
  INV_X1 U2627 ( .A(n3209), .ZN(n2998) );
  AND4_X1 U2628 ( .A1(n3797), .A2(n3796), .A3(n3795), .A4(n3794), .ZN(n4214)
         );
  OR2_X1 U2629 ( .A1(n5029), .A2(n3629), .ZN(n2624) );
  AND2_X1 U2630 ( .A1(n2912), .A2(n5042), .ZN(n2915) );
  NAND2_X1 U2631 ( .A1(n2918), .A2(n2632), .ZN(n2628) );
  INV_X1 U2632 ( .A(n5051), .ZN(n2632) );
  NAND2_X1 U2633 ( .A1(n4178), .A2(n2833), .ZN(n5047) );
  AOI21_X1 U2634 ( .B1(n2734), .B2(n2739), .A(n4241), .ZN(n2733) );
  NOR2_X1 U2635 ( .A1(n2735), .A2(n2731), .ZN(n2730) );
  NAND2_X1 U2636 ( .A1(n3499), .A2(n5265), .ZN(n2727) );
  NAND2_X1 U2637 ( .A1(n5178), .A2(n5174), .ZN(n2578) );
  AND2_X1 U2638 ( .A1(n4165), .A2(n3227), .ZN(n3217) );
  AND2_X1 U2639 ( .A1(n3129), .A2(n2984), .ZN(n3037) );
  AND2_X1 U2640 ( .A1(n2747), .A2(n2588), .ZN(n2861) );
  AND4_X1 U2641 ( .A1(n2590), .A2(n2531), .A3(n2755), .A4(n2804), .ZN(n2588)
         );
  AND2_X1 U2642 ( .A1(n2804), .A2(n2528), .ZN(n2759) );
  AND2_X1 U2643 ( .A1(n2791), .A2(n2792), .ZN(n2811) );
  AND2_X1 U2644 ( .A1(n2580), .A2(n4104), .ZN(n2579) );
  OR2_X1 U2645 ( .A1(n5174), .A2(n2581), .ZN(n2580) );
  INV_X1 U2646 ( .A(n4009), .ZN(n2581) );
  XNOR2_X1 U2647 ( .A(n3157), .B(n3829), .ZN(n3161) );
  NAND2_X1 U2648 ( .A1(n3027), .A2(REG0_REG_2__SCAN_IN), .ZN(n3057) );
  INV_X1 U2649 ( .A(n4983), .ZN(n2639) );
  AOI21_X1 U2650 ( .B1(REG1_REG_7__SCAN_IN), .B2(n5171), .A(n4986), .ZN(n2797)
         );
  NOR2_X1 U2651 ( .A1(n5003), .A2(n2906), .ZN(n2907) );
  AND2_X1 U2652 ( .A1(n5010), .A2(REG2_REG_9__SCAN_IN), .ZN(n2906) );
  AOI21_X1 U2653 ( .B1(REG2_REG_11__SCAN_IN), .B2(n5021), .A(n5014), .ZN(n2910) );
  OR2_X1 U2654 ( .A1(n2822), .A2(n2956), .ZN(n2824) );
  OR2_X1 U2655 ( .A1(n4220), .A2(n2737), .ZN(n2736) );
  NAND2_X1 U2656 ( .A1(n4216), .A2(n4215), .ZN(n2737) );
  INV_X1 U2657 ( .A(n2571), .ZN(n2570) );
  NAND2_X1 U2658 ( .A1(n2569), .A2(n2571), .ZN(n2568) );
  INV_X1 U2659 ( .A(n4131), .ZN(n2569) );
  NOR2_X1 U2660 ( .A1(n2572), .A2(n4130), .ZN(n2571) );
  OR2_X1 U2661 ( .A1(n4228), .A2(n4292), .ZN(n2599) );
  INV_X1 U2662 ( .A(n4211), .ZN(n2745) );
  INV_X1 U2663 ( .A(n4327), .ZN(n2742) );
  OR2_X1 U2664 ( .A1(n3835), .A2(n4293), .ZN(n3779) );
  INV_X1 U2665 ( .A(n2712), .ZN(n2711) );
  OAI21_X1 U2666 ( .B1(n2534), .B2(n2713), .A(n4207), .ZN(n2712) );
  AND2_X1 U2667 ( .A1(n4403), .A2(n4428), .ZN(n2600) );
  NOR2_X1 U2668 ( .A1(n4119), .A2(n4118), .ZN(n4439) );
  NAND2_X1 U2669 ( .A1(n5304), .A2(n2596), .ZN(n2595) );
  INV_X1 U2670 ( .A(n4077), .ZN(n2724) );
  NOR2_X1 U2671 ( .A1(n5261), .A2(n2726), .ZN(n2725) );
  INV_X1 U2672 ( .A(n3497), .ZN(n2726) );
  NAND2_X1 U2673 ( .A1(n5257), .A2(n5265), .ZN(n3500) );
  NOR2_X1 U2674 ( .A1(n5174), .A2(n2535), .ZN(n2720) );
  NAND2_X1 U2675 ( .A1(n2547), .A2(n2719), .ZN(n2718) );
  OR2_X1 U2676 ( .A1(n3395), .A2(n2535), .ZN(n2719) );
  INV_X1 U2677 ( .A(n5179), .ZN(n5187) );
  NAND2_X1 U2678 ( .A1(n2856), .A2(n2855), .ZN(n2883) );
  NOR2_X1 U2679 ( .A1(IR_REG_24__SCAN_IN), .A2(IR_REG_23__SCAN_IN), .ZN(n2855)
         );
  INV_X1 U2680 ( .A(n2872), .ZN(n2856) );
  OAI21_X1 U2681 ( .B1(n2968), .B2(n2872), .A(IR_REG_31__SCAN_IN), .ZN(n2873)
         );
  NOR2_X1 U2682 ( .A1(n2852), .A2(n2851), .ZN(n2853) );
  INV_X1 U2683 ( .A(IR_REG_19__SCAN_IN), .ZN(n2849) );
  XNOR2_X1 U2684 ( .A(n3102), .B(n3829), .ZN(n3105) );
  INV_X1 U2685 ( .A(n2688), .ZN(n2687) );
  OAI21_X1 U2686 ( .B1(n3879), .B2(n2689), .A(n3943), .ZN(n2688) );
  NAND2_X1 U2687 ( .A1(n2683), .A2(n5239), .ZN(n2679) );
  NAND2_X1 U2688 ( .A1(n3122), .A2(n3347), .ZN(n3264) );
  AND2_X1 U2689 ( .A1(n3123), .A2(n3124), .ZN(n3122) );
  NAND2_X1 U2690 ( .A1(n2527), .A2(n2681), .ZN(n2675) );
  NAND2_X1 U2691 ( .A1(n2677), .A2(n2681), .ZN(n2676) );
  INV_X1 U2692 ( .A(n2679), .ZN(n2677) );
  NOR2_X1 U2693 ( .A1(n3345), .A2(n3115), .ZN(n3968) );
  NOR2_X1 U2694 ( .A1(IR_REG_27__SCAN_IN), .A2(IR_REG_31__SCAN_IN), .ZN(n2859)
         );
  NOR2_X1 U2695 ( .A1(n5056), .A2(n2893), .ZN(n2894) );
  OAI21_X1 U2696 ( .B1(n5090), .B2(n2612), .A(n2611), .ZN(n4972) );
  NAND2_X1 U2697 ( .A1(n2615), .A2(REG1_REG_4__SCAN_IN), .ZN(n2612) );
  INV_X1 U2698 ( .A(n4973), .ZN(n2615) );
  NOR2_X1 U2699 ( .A1(n4972), .A2(n2790), .ZN(n2794) );
  AND2_X1 U2700 ( .A1(n4979), .A2(REG1_REG_5__SCAN_IN), .ZN(n2790) );
  AND3_X1 U2701 ( .A1(n2648), .A2(n2646), .A3(n2551), .ZN(n2899) );
  OR2_X1 U2702 ( .A1(n3076), .A2(n3287), .ZN(n2638) );
  XNOR2_X1 U2703 ( .A(n2797), .B(n3315), .ZN(n4993) );
  XNOR2_X1 U2704 ( .A(n2907), .B(n3483), .ZN(n3485) );
  NOR2_X1 U2705 ( .A1(n3480), .A2(n2809), .ZN(n5018) );
  OR2_X1 U2706 ( .A1(n5018), .A2(n5017), .ZN(n2601) );
  NOR2_X1 U2707 ( .A1(n5026), .A2(n5025), .ZN(n5024) );
  NOR2_X1 U2708 ( .A1(n5039), .A2(n5300), .ZN(n5038) );
  NAND2_X1 U2709 ( .A1(n2629), .A2(n2627), .ZN(n2939) );
  NAND2_X1 U2710 ( .A1(n2628), .A2(n2919), .ZN(n2627) );
  AND2_X1 U2711 ( .A1(n2919), .A2(n4181), .ZN(n2630) );
  NOR2_X1 U2712 ( .A1(n2939), .A2(n2940), .ZN(n2941) );
  OR2_X1 U2713 ( .A1(n2520), .A2(n4229), .ZN(n5370) );
  OR2_X1 U2714 ( .A1(n3822), .A2(n4579), .ZN(n4231) );
  INV_X1 U2715 ( .A(n4221), .ZN(n4246) );
  INV_X1 U2716 ( .A(n4215), .ZN(n2740) );
  AND4_X1 U2717 ( .A1(n3828), .A2(n3827), .A3(n3826), .A4(n3825), .ZN(n4255)
         );
  AND2_X1 U2718 ( .A1(n4191), .A2(n4085), .ZN(n4256) );
  AND2_X1 U2719 ( .A1(n2573), .A2(n4075), .ZN(n4275) );
  AOI21_X1 U2720 ( .B1(n4326), .B2(n4127), .A(n4126), .ZN(n4311) );
  AND2_X1 U2721 ( .A1(n4360), .A2(n4351), .ZN(n4343) );
  NAND2_X1 U2722 ( .A1(n2515), .A2(n2543), .ZN(n2714) );
  NAND2_X1 U2723 ( .A1(n4444), .A2(n4428), .ZN(n4203) );
  NOR2_X1 U2724 ( .A1(n2519), .A2(n4442), .ZN(n4434) );
  NAND2_X1 U2725 ( .A1(n2698), .A2(n2697), .ZN(n4436) );
  AOI22_X1 U2726 ( .A1(n2703), .A2(n2705), .B1(n2700), .B2(n2702), .ZN(n2697)
         );
  NAND2_X1 U2727 ( .A1(n2707), .A2(n2706), .ZN(n2705) );
  OR2_X1 U2728 ( .A1(n3522), .A2(n4572), .ZN(n3562) );
  AND2_X1 U2729 ( .A1(n3533), .A2(n3558), .ZN(n4077) );
  NAND2_X1 U2730 ( .A1(n3498), .A2(n2725), .ZN(n2728) );
  NAND2_X1 U2731 ( .A1(n3470), .A2(n4158), .ZN(n3497) );
  AND2_X1 U2732 ( .A1(n4019), .A2(n4022), .ZN(n5261) );
  OAI21_X1 U2733 ( .B1(n5173), .B2(n2716), .A(n2715), .ZN(n3474) );
  OAI21_X1 U2734 ( .B1(n2718), .B2(n2552), .A(n2717), .ZN(n2715) );
  NAND2_X1 U2735 ( .A1(n2720), .A2(n2717), .ZN(n2716) );
  INV_X1 U2736 ( .A(n4093), .ZN(n2717) );
  AND4_X1 U2737 ( .A1(n3419), .A2(n3418), .A3(n3417), .A4(n3416), .ZN(n3499)
         );
  AND2_X1 U2738 ( .A1(n3171), .A2(REG3_REG_7__SCAN_IN), .ZN(n3333) );
  NAND2_X1 U2739 ( .A1(n3380), .A2(n4082), .ZN(n3381) );
  NAND2_X1 U2740 ( .A1(n3394), .A2(n3393), .ZN(n5176) );
  OAI21_X1 U2741 ( .B1(n5128), .B2(n3207), .A(n3206), .ZN(n3242) );
  AND2_X1 U2742 ( .A1(n4140), .A2(n3190), .ZN(n5138) );
  OR2_X1 U2743 ( .A1(n2968), .A2(n2966), .ZN(n2865) );
  INV_X1 U2744 ( .A(n2968), .ZN(n2885) );
  AOI22_X1 U2745 ( .A1(n2997), .A2(n2694), .B1(n2692), .B2(n2691), .ZN(n2690)
         );
  NAND2_X1 U2746 ( .A1(IR_REG_20__SCAN_IN), .A2(n2693), .ZN(n2692) );
  AND2_X1 U2747 ( .A1(n2804), .A2(n2757), .ZN(n2810) );
  NAND2_X1 U2748 ( .A1(n2975), .A2(n2521), .ZN(n3129) );
  NOR2_X1 U2749 ( .A1(n2661), .A2(n5344), .ZN(n2659) );
  AND2_X1 U2750 ( .A1(n2663), .A2(n2532), .ZN(n2661) );
  NAND2_X1 U2751 ( .A1(n2663), .A2(n2545), .ZN(n2662) );
  INV_X1 U2752 ( .A(n4014), .ZN(n3472) );
  NAND2_X1 U2753 ( .A1(n3041), .A2(n2891), .ZN(n3043) );
  INV_X1 U2754 ( .A(n3382), .ZN(n4161) );
  OR2_X1 U2755 ( .A1(n3026), .A2(n2991), .ZN(n2994) );
  NAND2_X1 U2756 ( .A1(n2914), .A2(n2913), .ZN(n5037) );
  INV_X1 U2757 ( .A(n5069), .ZN(n5098) );
  XNOR2_X1 U2758 ( .A(n2574), .B(n5366), .ZN(n5378) );
  NOR2_X1 U2759 ( .A1(n5370), .A2(n5369), .ZN(n2574) );
  NAND2_X1 U2760 ( .A1(n2811), .A2(n2759), .ZN(n2760) );
  NAND2_X1 U2761 ( .A1(n2867), .A2(n2854), .ZN(n2872) );
  INV_X1 U2762 ( .A(n3169), .ZN(n2657) );
  AND2_X1 U2763 ( .A1(n2655), .A2(n3300), .ZN(n2654) );
  INV_X1 U2764 ( .A(n3167), .ZN(n2656) );
  NAND2_X1 U2765 ( .A1(n3300), .A2(n2657), .ZN(n2652) );
  OR2_X1 U2766 ( .A1(n3640), .A2(n3639), .ZN(n3652) );
  INV_X1 U2767 ( .A(n4213), .ZN(n2731) );
  AND2_X1 U2768 ( .A1(REG3_REG_17__SCAN_IN), .A2(n3584), .ZN(n3666) );
  AND2_X1 U2769 ( .A1(n3438), .A2(n3437), .ZN(n3449) );
  INV_X1 U2770 ( .A(n3436), .ZN(n3438) );
  NOR2_X1 U2771 ( .A1(n5186), .A2(n3472), .ZN(n2586) );
  NAND2_X1 U2772 ( .A1(n5135), .A2(n3191), .ZN(n3999) );
  AOI21_X1 U2773 ( .B1(n2579), .B2(n2581), .A(n2577), .ZN(n2576) );
  INV_X1 U2774 ( .A(n4008), .ZN(n2577) );
  OR2_X1 U2775 ( .A1(n3018), .A2(n3014), .ZN(n4462) );
  AND2_X1 U2776 ( .A1(n2589), .A2(n2757), .ZN(n2587) );
  NAND2_X1 U2777 ( .A1(IR_REG_19__SCAN_IN), .A2(IR_REG_31__SCAN_IN), .ZN(n2693) );
  NOR2_X1 U2778 ( .A1(n4633), .A2(n2871), .ZN(n2694) );
  NAND2_X1 U2779 ( .A1(n4633), .A2(IR_REG_31__SCAN_IN), .ZN(n2691) );
  INV_X1 U2780 ( .A(IR_REG_14__SCAN_IN), .ZN(n2835) );
  INV_X1 U2781 ( .A(IR_REG_5__SCAN_IN), .ZN(n2591) );
  AOI21_X1 U2782 ( .B1(n2670), .B2(n2668), .A(n2541), .ZN(n2667) );
  INV_X1 U2783 ( .A(n3803), .ZN(n2668) );
  INV_X1 U2784 ( .A(n2670), .ZN(n2669) );
  INV_X1 U2785 ( .A(n3833), .ZN(n2666) );
  AND2_X1 U2786 ( .A1(n3446), .A2(n3445), .ZN(n3515) );
  AOI21_X1 U2787 ( .B1(n3001), .B2(REG1_REG_0__SCAN_IN), .A(n3050), .ZN(n3052)
         );
  NAND2_X1 U2788 ( .A1(n2674), .A2(n2672), .ZN(n3636) );
  AOI21_X1 U2789 ( .B1(n2676), .B2(n2675), .A(n2673), .ZN(n2672) );
  INV_X1 U2790 ( .A(n3520), .ZN(n2673) );
  INV_X1 U2791 ( .A(n3958), .ZN(n3741) );
  INV_X1 U2792 ( .A(REG3_REG_6__SCAN_IN), .ZN(n3146) );
  NOR2_X1 U2793 ( .A1(n3147), .A2(n3146), .ZN(n3171) );
  OR2_X1 U2794 ( .A1(n3375), .A2(n5072), .ZN(n3982) );
  INV_X1 U2795 ( .A(n3210), .ZN(n3060) );
  OR2_X1 U2796 ( .A1(n3835), .A2(n4267), .ZN(n3811) );
  OR2_X1 U2797 ( .A1(n3835), .A2(n4320), .ZN(n3766) );
  AND4_X1 U2798 ( .A1(n3591), .A2(n3590), .A3(n3589), .A4(n3588), .ZN(n4418)
         );
  AND4_X1 U2799 ( .A1(n3090), .A2(n3089), .A3(n3088), .A4(n3087), .ZN(n3189)
         );
  OR2_X1 U2800 ( .A1(n3054), .A2(n3257), .ZN(n3058) );
  NAND2_X1 U2801 ( .A1(n2773), .A2(n2772), .ZN(n2774) );
  INV_X1 U2802 ( .A(IR_REG_1__SCAN_IN), .ZN(n2771) );
  OAI22_X1 U2803 ( .A1(n2891), .A2(REG2_REG_1__SCAN_IN), .B1(n2889), .B2(n2890), .ZN(n4961) );
  NOR2_X1 U2804 ( .A1(n5062), .A2(n5063), .ZN(n5061) );
  XNOR2_X1 U2805 ( .A(n2781), .B(n3099), .ZN(n3070) );
  NOR2_X1 U2806 ( .A1(n3070), .A2(n5144), .ZN(n3069) );
  NOR2_X1 U2807 ( .A1(n3067), .A2(n2895), .ZN(n2896) );
  OR2_X1 U2808 ( .A1(n5093), .A2(n2649), .ZN(n2648) );
  OR2_X1 U2809 ( .A1(n4977), .A2(n5094), .ZN(n2649) );
  NAND2_X1 U2810 ( .A1(n2897), .A2(n2647), .ZN(n2646) );
  INV_X1 U2811 ( .A(n4977), .ZN(n2647) );
  OR2_X1 U2812 ( .A1(n5093), .A2(n5094), .ZN(n2651) );
  OR2_X1 U2813 ( .A1(n5090), .A2(n5158), .ZN(n2614) );
  NAND2_X1 U2814 ( .A1(n2636), .A2(n2517), .ZN(n2635) );
  NAND2_X1 U2815 ( .A1(n2635), .A2(n2633), .ZN(n2903) );
  AND2_X1 U2816 ( .A1(n2634), .A2(n2901), .ZN(n2633) );
  NAND2_X1 U2817 ( .A1(n2619), .A2(REG1_REG_8__SCAN_IN), .ZN(n2618) );
  NAND2_X1 U2818 ( .A1(n2798), .A2(n2619), .ZN(n2617) );
  INV_X1 U2819 ( .A(n5007), .ZN(n2619) );
  NOR2_X1 U2820 ( .A1(n4993), .A2(n5205), .ZN(n4992) );
  NOR2_X1 U2821 ( .A1(n3485), .A2(n3486), .ZN(n3484) );
  NAND2_X1 U2822 ( .A1(n2601), .A2(n2813), .ZN(n2819) );
  OR2_X1 U2823 ( .A1(n3628), .A2(n3629), .ZN(n2626) );
  INV_X1 U2824 ( .A(n2824), .ZN(n2825) );
  NOR2_X1 U2825 ( .A1(n4166), .A2(n2827), .ZN(n2832) );
  AND2_X1 U2826 ( .A1(n4924), .A2(REG1_REG_15__SCAN_IN), .ZN(n2827) );
  INV_X1 U2827 ( .A(n2843), .ZN(n2609) );
  AND2_X1 U2828 ( .A1(n4923), .A2(REG2_REG_18__SCAN_IN), .ZN(n2921) );
  NAND2_X1 U2829 ( .A1(n2567), .A2(n2565), .ZN(n4240) );
  AOI21_X1 U2830 ( .B1(n2514), .B2(n2570), .A(n2566), .ZN(n2565) );
  INV_X1 U2831 ( .A(n4191), .ZN(n2566) );
  AND4_X1 U2832 ( .A1(n3840), .A2(n3839), .A3(n3838), .A4(n3837), .ZN(n4242)
         );
  INV_X1 U2833 ( .A(n2599), .ZN(n2598) );
  OR2_X1 U2834 ( .A1(n4298), .A2(n2570), .ZN(n2564) );
  NAND2_X1 U2835 ( .A1(n2573), .A2(n2571), .ZN(n4258) );
  NOR3_X1 U2836 ( .A1(n4308), .A2(n2599), .A3(n4217), .ZN(n4264) );
  INV_X1 U2837 ( .A(n4218), .ZN(n4276) );
  NOR2_X1 U2838 ( .A1(n4308), .A2(n2599), .ZN(n4280) );
  INV_X1 U2839 ( .A(n2744), .ZN(n2743) );
  AOI21_X1 U2840 ( .B1(n2744), .B2(n2742), .A(n2544), .ZN(n2741) );
  NOR2_X1 U2841 ( .A1(n4312), .A2(n2745), .ZN(n2744) );
  AND2_X1 U2842 ( .A1(n4075), .A2(n4074), .ZN(n4299) );
  AND4_X1 U2843 ( .A1(n3781), .A2(n3780), .A3(n3779), .A4(n3778), .ZN(n4313)
         );
  NAND2_X1 U2844 ( .A1(n4335), .A2(n4314), .ZN(n4308) );
  OR2_X1 U2845 ( .A1(n3744), .A2(n4762), .ZN(n3762) );
  AOI21_X1 U2846 ( .B1(n4367), .B2(n4107), .A(n4123), .ZN(n2583) );
  INV_X1 U2847 ( .A(n4152), .ZN(n4330) );
  AND2_X1 U2848 ( .A1(n4343), .A2(n4333), .ZN(n4335) );
  OR2_X1 U2849 ( .A1(n3732), .A2(n3959), .ZN(n3744) );
  NAND2_X1 U2850 ( .A1(n2585), .A2(n4107), .ZN(n4349) );
  AOI21_X1 U2851 ( .B1(n2711), .B2(n2713), .A(n2538), .ZN(n2709) );
  OR2_X1 U2852 ( .A1(n4124), .A2(n4123), .ZN(n4350) );
  AND4_X1 U2853 ( .A1(n3704), .A2(n3703), .A3(n3702), .A4(n3701), .ZN(n4365)
         );
  OR2_X1 U2854 ( .A1(n4368), .A2(n4367), .ZN(n2585) );
  NAND2_X1 U2855 ( .A1(n3713), .A2(REG3_REG_21__SCAN_IN), .ZN(n3732) );
  NOR2_X1 U2856 ( .A1(n3698), .A2(n3949), .ZN(n3713) );
  AND2_X1 U2857 ( .A1(n4434), .A2(n2555), .ZN(n4360) );
  NAND2_X1 U2858 ( .A1(n4434), .A2(n2518), .ZN(n4391) );
  NAND2_X1 U2859 ( .A1(n4434), .A2(n2600), .ZN(n4412) );
  NAND2_X1 U2860 ( .A1(n3683), .A2(REG3_REG_19__SCAN_IN), .ZN(n3698) );
  NAND2_X1 U2861 ( .A1(n4434), .A2(n4428), .ZN(n4427) );
  OAI22_X1 U2862 ( .A1(n4436), .A2(n4440), .B1(n4442), .B2(n4201), .ZN(n4426)
         );
  AOI21_X1 U2863 ( .B1(n3601), .B2(n2751), .A(n2546), .ZN(n2707) );
  NAND2_X1 U2864 ( .A1(n4073), .A2(n3598), .ZN(n3601) );
  NAND2_X1 U2865 ( .A1(n2594), .A2(n2593), .ZN(n2592) );
  NOR2_X1 U2866 ( .A1(n3859), .A2(n4200), .ZN(n2593) );
  INV_X1 U2867 ( .A(n2595), .ZN(n2594) );
  INV_X1 U2868 ( .A(REG3_REG_15__SCAN_IN), .ZN(n4169) );
  NOR2_X1 U2869 ( .A1(n3562), .A2(n4169), .ZN(n3578) );
  INV_X1 U2870 ( .A(REG3_REG_14__SCAN_IN), .ZN(n4572) );
  NOR3_X1 U2871 ( .A1(n3543), .A2(n3859), .A3(n3559), .ZN(n3616) );
  NOR2_X1 U2872 ( .A1(n3543), .A2(n3559), .ZN(n3555) );
  INV_X1 U2873 ( .A(n2722), .ZN(n2721) );
  OAI22_X1 U2874 ( .A1(n4077), .A2(n2727), .B1(n4156), .B2(n3540), .ZN(n2722)
         );
  OR2_X1 U2875 ( .A1(n3500), .A2(n3540), .ZN(n3543) );
  NOR2_X1 U2876 ( .A1(n5211), .A2(n3470), .ZN(n5257) );
  NAND2_X1 U2877 ( .A1(n2586), .A2(n5215), .ZN(n5211) );
  NAND2_X1 U2878 ( .A1(n5188), .A2(n5187), .ZN(n5186) );
  INV_X1 U2879 ( .A(n2586), .ZN(n5209) );
  AND4_X1 U2880 ( .A1(n3309), .A2(n3308), .A3(n3307), .A4(n3306), .ZN(n5183)
         );
  INV_X1 U2881 ( .A(n5246), .ZN(n5180) );
  AND2_X1 U2882 ( .A1(n3285), .A2(n3389), .ZN(n5188) );
  AND4_X1 U2883 ( .A1(n3176), .A2(n3175), .A3(n3174), .A4(n3173), .ZN(n3382)
         );
  AND4_X1 U2884 ( .A1(n3141), .A2(n3140), .A3(n3139), .A4(n3138), .ZN(n3281)
         );
  AND2_X1 U2885 ( .A1(n4006), .A2(n4002), .ZN(n4082) );
  NOR2_X1 U2886 ( .A1(n3237), .A2(n3270), .ZN(n3285) );
  OR2_X1 U2887 ( .A1(n2926), .A2(n3210), .ZN(n5246) );
  NAND2_X1 U2888 ( .A1(n2562), .A2(n3191), .ZN(n3237) );
  INV_X1 U2889 ( .A(n2563), .ZN(n2562) );
  INV_X1 U2890 ( .A(n3350), .ZN(n5132) );
  AND2_X1 U2891 ( .A1(n3996), .A2(n3993), .ZN(n5131) );
  NAND2_X1 U2892 ( .A1(n4084), .A2(n2560), .ZN(n3221) );
  INV_X1 U2893 ( .A(n3184), .ZN(n3222) );
  INV_X1 U2894 ( .A(n3227), .ZN(n5105) );
  AND2_X1 U2895 ( .A1(n3037), .A2(n3127), .ZN(n4463) );
  OR2_X1 U2896 ( .A1(n3018), .A2(D_REG_0__SCAN_IN), .ZN(n3020) );
  NAND2_X1 U2897 ( .A1(n4325), .A2(n4327), .ZN(n2746) );
  AOI21_X1 U2898 ( .B1(n3394), .B2(n2720), .A(n2718), .ZN(n5207) );
  INV_X1 U2899 ( .A(n5335), .ZN(n5296) );
  NAND2_X1 U2900 ( .A1(n5102), .A2(n5122), .ZN(n5335) );
  INV_X1 U2901 ( .A(n4465), .ZN(n4504) );
  INV_X1 U2902 ( .A(IR_REG_29__SCAN_IN), .ZN(n4843) );
  INV_X1 U2903 ( .A(IR_REG_28__SCAN_IN), .ZN(n4839) );
  XNOR2_X1 U2904 ( .A(n2887), .B(n4834), .ZN(n2978) );
  NAND2_X1 U2905 ( .A1(n2886), .A2(IR_REG_31__SCAN_IN), .ZN(n2887) );
  INV_X1 U2906 ( .A(n2883), .ZN(n2884) );
  INV_X1 U2907 ( .A(IR_REG_15__SCAN_IN), .ZN(n2834) );
  INV_X1 U2908 ( .A(IR_REG_9__SCAN_IN), .ZN(n2756) );
  AND2_X1 U2909 ( .A1(n3349), .A2(n3968), .ZN(n3121) );
  NAND2_X1 U2910 ( .A1(n2686), .A2(n2684), .ZN(n3893) );
  AOI21_X1 U2911 ( .B1(n2687), .B2(n2689), .A(n2685), .ZN(n2684) );
  INV_X1 U2912 ( .A(n3944), .ZN(n2685) );
  OR2_X1 U2913 ( .A1(n3426), .A2(n2679), .ZN(n2678) );
  OAI21_X1 U2914 ( .B1(n3933), .B2(n3935), .A(n3932), .ZN(n3905) );
  OR2_X1 U2915 ( .A1(n3035), .A2(n4146), .ZN(n3375) );
  NAND2_X1 U2916 ( .A1(n3877), .A2(n3696), .ZN(n3945) );
  NOR2_X1 U2917 ( .A1(n3426), .A2(n2680), .ZN(n5243) );
  INV_X1 U2918 ( .A(n5302), .ZN(n3980) );
  OAI21_X1 U2919 ( .B1(n3038), .B2(n5266), .A(n5231), .ZN(n3972) );
  INV_X1 U2920 ( .A(n5305), .ZN(n5339) );
  NAND2_X1 U2921 ( .A1(n3262), .A2(n3167), .ZN(n3168) );
  INV_X1 U2922 ( .A(n3599), .ZN(n5304) );
  INV_X1 U2923 ( .A(n3972), .ZN(n5305) );
  AND4_X1 U2924 ( .A1(n3528), .A2(n3527), .A3(n3526), .A4(n3525), .ZN(n5303)
         );
  INV_X1 U2925 ( .A(n3982), .ZN(n5309) );
  INV_X1 U2926 ( .A(n4214), .ZN(n4303) );
  INV_X1 U2927 ( .A(n4313), .ZN(n4212) );
  INV_X1 U2928 ( .A(n4418), .ZN(n4201) );
  INV_X1 U2929 ( .A(n3499), .ZN(n4157) );
  INV_X1 U2930 ( .A(n3281), .ZN(n4162) );
  INV_X1 U2931 ( .A(n3189), .ZN(n5135) );
  INV_X1 U2932 ( .A(n5133), .ZN(n4164) );
  NAND2_X1 U2933 ( .A1(n2864), .A2(n2863), .ZN(n5071) );
  NAND2_X1 U2934 ( .A1(n2881), .A2(n2862), .ZN(n2863) );
  NOR2_X1 U2935 ( .A1(n2857), .A2(n2871), .ZN(n2862) );
  NOR2_X1 U2936 ( .A1(n3066), .A2(n3068), .ZN(n3067) );
  INV_X1 U2937 ( .A(n2614), .ZN(n5089) );
  NAND2_X1 U2938 ( .A1(n2646), .A2(n2648), .ZN(n4976) );
  INV_X1 U2939 ( .A(n2786), .ZN(n2613) );
  INV_X1 U2940 ( .A(n2638), .ZN(n3075) );
  NAND2_X1 U2941 ( .A1(n2635), .A2(n2634), .ZN(n4982) );
  INV_X1 U2942 ( .A(n2900), .ZN(n2637) );
  XNOR2_X1 U2943 ( .A(n2903), .B(n4999), .ZN(n4996) );
  NOR2_X1 U2944 ( .A1(n4995), .A2(n4996), .ZN(n4994) );
  OAI21_X1 U2945 ( .B1(n3485), .B2(n2641), .A(n2640), .ZN(n5014) );
  NAND2_X1 U2946 ( .A1(n2642), .A2(REG2_REG_10__SCAN_IN), .ZN(n2641) );
  INV_X1 U2947 ( .A(n2601), .ZN(n5016) );
  XNOR2_X1 U2948 ( .A(n2819), .B(n2818), .ZN(n3623) );
  OAI21_X1 U2949 ( .B1(n5037), .B2(n2644), .A(n2643), .ZN(n4172) );
  NAND2_X1 U2950 ( .A1(n2645), .A2(REG2_REG_14__SCAN_IN), .ZN(n2644) );
  INV_X1 U2951 ( .A(n4173), .ZN(n2645) );
  XNOR2_X1 U2952 ( .A(n2832), .B(n2831), .ZN(n4179) );
  NAND2_X1 U2953 ( .A1(n4179), .A2(n5329), .ZN(n4178) );
  OR2_X1 U2954 ( .A1(n4958), .A2(n5072), .ZN(n5069) );
  INV_X1 U2955 ( .A(n2628), .ZN(n2631) );
  NAND2_X1 U2956 ( .A1(n4180), .A2(n2918), .ZN(n5050) );
  OR2_X1 U2957 ( .A1(n4958), .A2(n5074), .ZN(n5091) );
  NAND2_X1 U2958 ( .A1(n2938), .A2(n2556), .ZN(n2603) );
  OR2_X1 U2959 ( .A1(n2609), .A2(n2847), .ZN(n2608) );
  INV_X1 U2960 ( .A(n2606), .ZN(n2605) );
  OAI21_X1 U2961 ( .B1(n2608), .B2(n2937), .A(n2607), .ZN(n2606) );
  NAND2_X1 U2962 ( .A1(n2847), .A2(n2609), .ZN(n2607) );
  NOR2_X1 U2963 ( .A1(n2941), .A2(n2921), .ZN(n2925) );
  INV_X1 U2964 ( .A(n4225), .ZN(n4226) );
  NAND2_X1 U2965 ( .A1(n4222), .A2(n4221), .ZN(n4223) );
  NAND2_X1 U2966 ( .A1(n2732), .A2(n2734), .ZN(n4238) );
  NAND2_X1 U2967 ( .A1(n4273), .A2(n2738), .ZN(n2732) );
  OAI21_X1 U2968 ( .B1(n4273), .B2(n4216), .A(n4215), .ZN(n4254) );
  NAND2_X1 U2969 ( .A1(n2710), .A2(n2714), .ZN(n4359) );
  NAND2_X1 U2970 ( .A1(n4407), .A2(n2534), .ZN(n2710) );
  NAND2_X1 U2971 ( .A1(n4407), .A2(n4205), .ZN(n4375) );
  AND2_X1 U2972 ( .A1(n2728), .A2(n2727), .ZN(n3541) );
  NAND2_X1 U2973 ( .A1(n3498), .A2(n3497), .ZN(n5255) );
  NAND2_X1 U2974 ( .A1(n2578), .A2(n4009), .ZN(n3462) );
  NAND2_X1 U2975 ( .A1(n5176), .A2(n3395), .ZN(n3473) );
  AND2_X1 U2976 ( .A1(n5226), .A2(n5177), .ZN(n4437) );
  INV_X1 U2977 ( .A(n4461), .ZN(n3036) );
  NAND2_X1 U2978 ( .A1(n4084), .A2(n2561), .ZN(n3218) );
  INV_X1 U2979 ( .A(n3217), .ZN(n2561) );
  AND2_X1 U2980 ( .A1(n5226), .A2(n4138), .ZN(n4247) );
  AOI21_X1 U2981 ( .B1(n5378), .B2(n5377), .A(n5376), .ZN(n5381) );
  INV_X1 U2982 ( .A(n2989), .ZN(n4918) );
  AND2_X1 U2983 ( .A1(n2882), .A2(n2881), .ZN(n4919) );
  MUX2_X1 U2984 ( .A(IR_REG_31__SCAN_IN), .B(n2880), .S(IR_REG_26__SCAN_IN), 
        .Z(n2882) );
  XNOR2_X1 U2985 ( .A(n2877), .B(IR_REG_24__SCAN_IN), .ZN(n2975) );
  AND2_X1 U2986 ( .A1(n3128), .A2(STATE_REG_SCAN_IN), .ZN(n2984) );
  XNOR2_X1 U2987 ( .A(n2869), .B(n2854), .ZN(n3208) );
  XNOR2_X1 U2988 ( .A(n2870), .B(IR_REG_21__SCAN_IN), .ZN(n4921) );
  AND2_X1 U2989 ( .A1(n2840), .A2(n2838), .ZN(n5048) );
  XNOR2_X1 U2990 ( .A(n2815), .B(IR_REG_11__SCAN_IN), .ZN(n5021) );
  XNOR2_X1 U2991 ( .A(n2801), .B(IR_REG_9__SCAN_IN), .ZN(n5010) );
  XNOR2_X1 U2992 ( .A(n2764), .B(IR_REG_7__SCAN_IN), .ZN(n5171) );
  XNOR2_X1 U2993 ( .A(n2788), .B(IR_REG_5__SCAN_IN), .ZN(n4979) );
  NAND2_X1 U2994 ( .A1(n2871), .A2(n4800), .ZN(n2767) );
  NAND2_X1 U2995 ( .A1(n2766), .A2(IR_REG_2__SCAN_IN), .ZN(n2768) );
  NAND2_X1 U2996 ( .A1(n2662), .A2(n5314), .ZN(n2660) );
  NAND2_X1 U2997 ( .A1(n2621), .A2(n2620), .ZN(n5031) );
  OAI21_X1 U2998 ( .B1(n2602), .B2(n2604), .A(n2935), .ZN(U3259) );
  AND2_X1 U2999 ( .A1(n2934), .A2(n2933), .ZN(n2935) );
  OAI21_X1 U3000 ( .B1(n2938), .B2(n2608), .A(n2605), .ZN(n2604) );
  NAND2_X1 U3001 ( .A1(n2603), .A2(n5065), .ZN(n2602) );
  AOI22_X1 U3002 ( .A1(n5381), .A2(n5363), .B1(n5379), .B2(n4056), .ZN(U3549)
         );
  AND2_X1 U3003 ( .A1(n2526), .A2(n2568), .ZN(n2514) );
  NAND2_X1 U3004 ( .A1(n2774), .A2(n2775), .ZN(n2889) );
  AND2_X1 U3005 ( .A1(n4007), .A2(n4009), .ZN(n5174) );
  INV_X1 U3006 ( .A(n5174), .ZN(n3393) );
  OR2_X1 U3007 ( .A1(n4206), .A2(n4390), .ZN(n2515) );
  INV_X1 U3008 ( .A(n4132), .ZN(n2572) );
  OR2_X1 U3009 ( .A1(n2583), .A2(n4124), .ZN(n2516) );
  AND2_X1 U3010 ( .A1(n2639), .A2(REG2_REG_6__SCAN_IN), .ZN(n2517) );
  INV_X1 U3011 ( .A(n5338), .ZN(n4428) );
  AND2_X1 U3012 ( .A1(n2600), .A2(n4386), .ZN(n2518) );
  OR2_X1 U3013 ( .A1(n3543), .A2(n2592), .ZN(n2519) );
  OR2_X1 U3014 ( .A1(n4308), .A2(n2597), .ZN(n2520) );
  AND2_X1 U3015 ( .A1(n4919), .A2(n4920), .ZN(n2521) );
  INV_X1 U3016 ( .A(IR_REG_20__SCAN_IN), .ZN(n4633) );
  AND4_X1 U3017 ( .A1(n3032), .A2(n3031), .A3(n3030), .A4(n3029), .ZN(n3185)
         );
  OR2_X1 U3018 ( .A1(n2910), .A2(n3626), .ZN(n2522) );
  NAND2_X1 U3019 ( .A1(n3043), .A2(n3042), .ZN(n3184) );
  NAND2_X1 U3020 ( .A1(n2746), .A2(n4211), .ZN(n4309) );
  NAND2_X1 U3021 ( .A1(n2992), .A2(n4918), .ZN(n3136) );
  INV_X1 U3022 ( .A(n2889), .ZN(n2891) );
  OR2_X1 U3023 ( .A1(n4289), .A2(n4299), .ZN(n2749) );
  NAND2_X1 U3024 ( .A1(n2755), .A2(n2748), .ZN(n2787) );
  INV_X1 U3025 ( .A(IR_REG_21__SCAN_IN), .ZN(n2867) );
  AND2_X1 U3026 ( .A1(n2891), .A2(REG2_REG_1__SCAN_IN), .ZN(n2523) );
  AND2_X1 U3027 ( .A1(n2631), .A2(n4180), .ZN(n2524) );
  OR3_X1 U3028 ( .A1(n2997), .A2(IR_REG_20__SCAN_IN), .A3(IR_REG_19__SCAN_IN), 
        .ZN(n2525) );
  AND2_X1 U3029 ( .A1(n4256), .A2(n4257), .ZN(n2526) );
  INV_X1 U3030 ( .A(n2683), .ZN(n2680) );
  NAND2_X1 U3031 ( .A1(n3427), .A2(n3428), .ZN(n2683) );
  NAND2_X1 U3032 ( .A1(n2682), .A2(n3518), .ZN(n2527) );
  AND2_X1 U3033 ( .A1(n2758), .A2(n2757), .ZN(n2528) );
  AND2_X1 U3034 ( .A1(n4926), .A2(REG1_REG_2__SCAN_IN), .ZN(n2529) );
  AND2_X1 U3035 ( .A1(n3324), .A2(n2652), .ZN(n2530) );
  AND2_X1 U3036 ( .A1(n2587), .A2(n2758), .ZN(n2531) );
  NAND2_X1 U3037 ( .A1(n2667), .A2(n2666), .ZN(n2532) );
  INV_X1 U3038 ( .A(IR_REG_13__SCAN_IN), .ZN(n2696) );
  INV_X1 U3039 ( .A(IR_REG_26__SCAN_IN), .ZN(n2589) );
  INV_X1 U3040 ( .A(IR_REG_22__SCAN_IN), .ZN(n2854) );
  NAND2_X1 U3041 ( .A1(n2723), .A2(n2721), .ZN(n3597) );
  INV_X1 U3042 ( .A(IR_REG_10__SCAN_IN), .ZN(n2757) );
  INV_X1 U3043 ( .A(n4109), .ZN(n2560) );
  NOR2_X1 U3044 ( .A1(n4308), .A2(n4292), .ZN(n2533) );
  AND2_X1 U3045 ( .A1(n2515), .A2(n4205), .ZN(n2534) );
  INV_X1 U3046 ( .A(n4444), .ZN(n4202) );
  AND2_X1 U3047 ( .A1(n5183), .A2(n4014), .ZN(n2535) );
  AND2_X1 U3048 ( .A1(n2699), .A2(n2707), .ZN(n2536) );
  NOR2_X1 U3049 ( .A1(n3976), .A2(n3977), .ZN(n2537) );
  AND2_X1 U3050 ( .A1(n4208), .A2(n4361), .ZN(n2538) );
  AND2_X1 U3051 ( .A1(n2626), .A2(n2522), .ZN(n2539) );
  OR3_X1 U3052 ( .A1(n3543), .A2(n2595), .A3(n3859), .ZN(n2540) );
  NOR2_X1 U3053 ( .A1(n5037), .A2(n5036), .ZN(n5035) );
  AND2_X1 U3054 ( .A1(n3819), .A2(n3820), .ZN(n2541) );
  NOR2_X1 U3055 ( .A1(n5035), .A2(n2915), .ZN(n2542) );
  AND2_X1 U3056 ( .A1(n4206), .A2(n4390), .ZN(n2543) );
  AND2_X1 U3057 ( .A1(n4330), .A2(n4314), .ZN(n2544) );
  INV_X1 U3058 ( .A(n2739), .ZN(n2738) );
  OR2_X1 U3059 ( .A1(n4220), .A2(n2740), .ZN(n2739) );
  OR2_X1 U3060 ( .A1(n2669), .A2(n2666), .ZN(n2545) );
  INV_X1 U3061 ( .A(IR_REG_27__SCAN_IN), .ZN(n2857) );
  INV_X1 U3062 ( .A(n2735), .ZN(n2734) );
  NAND2_X1 U3063 ( .A1(n2736), .A2(n4219), .ZN(n2735) );
  INV_X1 U3064 ( .A(n4124), .ZN(n2584) );
  NOR2_X1 U3065 ( .A1(n3643), .A2(n5304), .ZN(n2546) );
  NAND4_X1 U3066 ( .A1(n3582), .A2(n3581), .A3(n3580), .A4(n3579), .ZN(n5308)
         );
  INV_X1 U3067 ( .A(n5308), .ZN(n2706) );
  NAND2_X1 U3068 ( .A1(n4160), .A2(n3472), .ZN(n2547) );
  AND2_X1 U3069 ( .A1(n2678), .A2(n2682), .ZN(n2548) );
  OR2_X1 U3070 ( .A1(n2703), .A2(n2700), .ZN(n2549) );
  AND2_X1 U3071 ( .A1(n2724), .A2(n2725), .ZN(n2550) );
  NAND2_X1 U3072 ( .A1(n4979), .A2(REG2_REG_5__SCAN_IN), .ZN(n2551) );
  INV_X1 U3073 ( .A(n5344), .ZN(n5314) );
  NAND2_X1 U3074 ( .A1(n3168), .A2(n3169), .ZN(n3301) );
  INV_X1 U3075 ( .A(IR_REG_6__SCAN_IN), .ZN(n2792) );
  AND2_X1 U3076 ( .A1(n4159), .A2(n5208), .ZN(n2552) );
  INV_X1 U3077 ( .A(n4364), .ZN(n4361) );
  NOR2_X1 U3078 ( .A1(n4992), .A2(n2798), .ZN(n2553) );
  NOR2_X1 U3079 ( .A1(n3484), .A2(n2908), .ZN(n2554) );
  AND2_X1 U3080 ( .A1(n4064), .A2(DATAI_20_), .ZN(n4390) );
  AND2_X1 U3081 ( .A1(n2518), .A2(n4364), .ZN(n2555) );
  INV_X1 U3082 ( .A(n5029), .ZN(n2625) );
  XNOR2_X1 U3083 ( .A(n2866), .B(n4839), .ZN(n2926) );
  INV_X1 U3084 ( .A(n3559), .ZN(n2596) );
  OR2_X1 U3085 ( .A1(n4958), .A2(n4954), .ZN(n5088) );
  AND2_X1 U3086 ( .A1(n2937), .A2(n2847), .ZN(n2556) );
  AND2_X1 U3087 ( .A1(n2638), .A2(n2637), .ZN(n2557) );
  AND2_X1 U3088 ( .A1(n2614), .A2(n2613), .ZN(n2558) );
  AND2_X1 U3089 ( .A1(n2651), .A2(n2650), .ZN(n2559) );
  INV_X1 U3090 ( .A(n4217), .ZN(n4266) );
  NAND2_X1 U3091 ( .A1(n4114), .A2(n3208), .ZN(n5106) );
  OAI21_X1 U3092 ( .B1(n5132), .B2(n5129), .A(n2563), .ZN(n5147) );
  AOI21_X1 U3093 ( .B1(n2563), .B2(n3240), .A(n5333), .ZN(n3197) );
  NAND2_X1 U3094 ( .A1(n5132), .A2(n5129), .ZN(n2563) );
  NAND2_X1 U3095 ( .A1(n4298), .A2(n4131), .ZN(n2573) );
  NAND2_X1 U3096 ( .A1(n4298), .A2(n2514), .ZN(n2567) );
  NAND2_X1 U3097 ( .A1(n5178), .A2(n2579), .ZN(n2575) );
  NAND2_X1 U3098 ( .A1(n2575), .A2(n2576), .ZN(n5213) );
  OAI21_X2 U3099 ( .B1(n3274), .B2(n4080), .A(n4000), .ZN(n3380) );
  NAND3_X1 U3100 ( .A1(n4368), .A2(n4107), .A3(n2584), .ZN(n2582) );
  INV_X1 U3101 ( .A(n2585), .ZN(n4366) );
  AND2_X1 U3102 ( .A1(n2590), .A2(n2755), .ZN(n2791) );
  NAND3_X1 U3103 ( .A1(n2747), .A2(n2759), .A3(n2791), .ZN(n2968) );
  NAND3_X1 U3104 ( .A1(n2598), .A2(n4266), .A3(n4246), .ZN(n2597) );
  NOR2_X1 U3105 ( .A1(n5061), .A2(n2529), .ZN(n2781) );
  NAND2_X1 U3106 ( .A1(n2938), .A2(n2937), .ZN(n2936) );
  NAND2_X1 U3107 ( .A1(n2786), .A2(n2615), .ZN(n2611) );
  NAND3_X1 U3108 ( .A1(n2775), .A2(n2774), .A3(REG1_REG_1__SCAN_IN), .ZN(n2616) );
  NAND2_X1 U3109 ( .A1(n2777), .A2(n2616), .ZN(n4965) );
  OAI21_X1 U3110 ( .B1(n4993), .B2(n2618), .A(n2617), .ZN(n5006) );
  NOR2_X1 U3111 ( .A1(n3623), .A2(n5288), .ZN(n3622) );
  NAND2_X1 U3112 ( .A1(n3628), .A2(n2522), .ZN(n2620) );
  AOI21_X1 U3113 ( .B1(n2522), .B2(n3629), .A(n5029), .ZN(n2621) );
  OAI211_X1 U3114 ( .C1(n3628), .C2(n2624), .A(n2622), .B(n2911), .ZN(n2912)
         );
  NAND2_X1 U3115 ( .A1(n2623), .A2(n2625), .ZN(n2622) );
  INV_X1 U3116 ( .A(n2522), .ZN(n2623) );
  INV_X1 U3117 ( .A(n2626), .ZN(n3627) );
  NAND2_X1 U3118 ( .A1(n4182), .A2(n2630), .ZN(n2629) );
  NAND2_X1 U3119 ( .A1(n4182), .A2(n4181), .ZN(n4180) );
  INV_X1 U3120 ( .A(n3076), .ZN(n2636) );
  NAND2_X1 U3121 ( .A1(n2900), .A2(n2639), .ZN(n2634) );
  NAND2_X1 U3122 ( .A1(n2908), .A2(n2642), .ZN(n2640) );
  INV_X1 U3123 ( .A(n5015), .ZN(n2642) );
  NAND2_X1 U3124 ( .A1(n2915), .A2(n2645), .ZN(n2643) );
  INV_X1 U3125 ( .A(n2651), .ZN(n5092) );
  INV_X1 U3126 ( .A(n2897), .ZN(n2650) );
  NAND2_X1 U3127 ( .A1(n2656), .A2(n3169), .ZN(n2655) );
  NAND2_X1 U3128 ( .A1(n3262), .A2(n2654), .ZN(n2653) );
  NAND2_X1 U3129 ( .A1(n2653), .A2(n2530), .ZN(n3362) );
  OAI21_X1 U3130 ( .B1(n3262), .B2(n2657), .A(n2654), .ZN(n3325) );
  NAND2_X1 U3131 ( .A1(n3804), .A2(n2659), .ZN(n2658) );
  OAI211_X1 U3132 ( .C1(n3804), .C2(n2660), .A(n2658), .B(n3845), .ZN(U3217)
         );
  OAI21_X1 U3133 ( .B1(n3804), .B2(n2537), .A(n3803), .ZN(n3847) );
  NAND2_X1 U3134 ( .A1(n3426), .A2(n2675), .ZN(n2674) );
  OAI21_X1 U3135 ( .B1(n3426), .B2(n2676), .A(n2675), .ZN(n3519) );
  NAND2_X1 U3136 ( .A1(n3878), .A2(n2687), .ZN(n2686) );
  INV_X1 U3137 ( .A(n3696), .ZN(n2689) );
  NAND2_X1 U3138 ( .A1(n3878), .A2(n3879), .ZN(n3877) );
  AOI21_X2 U3139 ( .B1(n3869), .B2(n3772), .A(n3773), .ZN(n3933) );
  NAND2_X1 U3140 ( .A1(n2695), .A2(IR_REG_31__SCAN_IN), .ZN(n2837) );
  NAND4_X1 U3141 ( .A1(n2759), .A2(n2791), .A3(n2696), .A4(n2792), .ZN(n2695)
         );
  NAND2_X1 U3142 ( .A1(n3602), .A2(n2549), .ZN(n2698) );
  NAND2_X1 U3143 ( .A1(n3602), .A2(n2751), .ZN(n2699) );
  INV_X1 U3144 ( .A(n2751), .ZN(n2701) );
  INV_X1 U3145 ( .A(n2707), .ZN(n2702) );
  NAND2_X1 U3146 ( .A1(n4407), .A2(n2711), .ZN(n2708) );
  NAND2_X1 U3147 ( .A1(n2708), .A2(n2709), .ZN(n4342) );
  NAND2_X1 U31480 ( .A1(n3498), .A2(n2550), .ZN(n2723) );
  INV_X1 U31490 ( .A(n2728), .ZN(n5254) );
  NAND2_X1 U3150 ( .A1(n2749), .A2(n4213), .ZN(n4273) );
  NAND2_X1 U3151 ( .A1(n2729), .A2(n2733), .ZN(n4224) );
  NAND2_X1 U3152 ( .A1(n2749), .A2(n2730), .ZN(n2729) );
  OAI21_X1 U3153 ( .B1(n4325), .B2(n2743), .A(n2741), .ZN(n4289) );
  NAND2_X1 U3154 ( .A1(n3107), .A2(DATAI_1_), .ZN(n3042) );
  INV_X1 U3155 ( .A(n3107), .ZN(n3041) );
  NAND2_X1 U3156 ( .A1(n3264), .A2(n3166), .ZN(n3262) );
  OR2_X1 U3157 ( .A1(n3026), .A2(n4321), .ZN(n3767) );
  NAND2_X1 U3158 ( .A1(n2837), .A2(n2836), .ZN(n2845) );
  INV_X1 U3159 ( .A(n3185), .ZN(n3183) );
  NAND2_X1 U3160 ( .A1(n3854), .A2(n2754), .ZN(n5311) );
  XNOR2_X1 U3161 ( .A(n3049), .B(n3116), .ZN(n3119) );
  XNOR2_X1 U3162 ( .A(n3048), .B(n3829), .ZN(n3116) );
  XNOR2_X1 U3163 ( .A(n3106), .B(n3105), .ZN(n3349) );
  INV_X1 U3164 ( .A(n2992), .ZN(n2990) );
  AND2_X1 U3165 ( .A1(n4607), .A2(n2778), .ZN(n2748) );
  AND4_X1 U3166 ( .A1(n3371), .A2(n3370), .A3(n3369), .A4(n3368), .ZN(n5247)
         );
  INV_X1 U3167 ( .A(n4403), .ZN(n4410) );
  AND2_X1 U3168 ( .A1(n3167), .A2(n3162), .ZN(n2750) );
  AND2_X1 U3169 ( .A1(n3608), .A2(n3600), .ZN(n2751) );
  AND2_X1 U3170 ( .A1(n3001), .A2(IR_REG_0__SCAN_IN), .ZN(n2752) );
  NOR2_X1 U3171 ( .A1(n3662), .A2(n3925), .ZN(n2753) );
  AND2_X1 U3172 ( .A1(n3653), .A2(n3652), .ZN(n2754) );
  INV_X1 U3173 ( .A(n2846), .ZN(n4138) );
  INV_X1 U3174 ( .A(n3046), .ZN(n2846) );
  OR2_X1 U3175 ( .A1(n4153), .A2(n3599), .ZN(n3600) );
  INV_X1 U3176 ( .A(n3651), .ZN(n3653) );
  AND2_X1 U3177 ( .A1(n2857), .A2(n2589), .ZN(n2858) );
  NAND2_X1 U3178 ( .A1(n2889), .A2(n2776), .ZN(n2777) );
  OR2_X1 U3179 ( .A1(n4208), .A2(n4361), .ZN(n4207) );
  AND2_X1 U3180 ( .A1(n3302), .A2(n3303), .ZN(n3300) );
  NAND2_X1 U3181 ( .A1(n3161), .A2(n3160), .ZN(n3162) );
  AND2_X1 U3182 ( .A1(n3915), .A2(n5311), .ZN(n3654) );
  NAND2_X1 U3183 ( .A1(n3185), .A2(n3184), .ZN(n3990) );
  AND2_X1 U3184 ( .A1(n3326), .A2(n3327), .ZN(n3324) );
  AOI21_X1 U3185 ( .B1(n3740), .B2(n3227), .A(n2752), .ZN(n3002) );
  AND2_X1 U3186 ( .A1(REG3_REG_12__SCAN_IN), .A2(REG3_REG_11__SCAN_IN), .ZN(
        n3437) );
  AND2_X1 U3187 ( .A1(n3114), .A2(n3113), .ZN(n3115) );
  OR2_X1 U3188 ( .A1(n3791), .A2(n3981), .ZN(n3807) );
  INV_X1 U3189 ( .A(n4153), .ZN(n3643) );
  NAND2_X1 U3190 ( .A1(n3028), .A2(REG1_REG_1__SCAN_IN), .ZN(n3029) );
  INV_X1 U3191 ( .A(n3626), .ZN(n2818) );
  INV_X1 U3192 ( .A(n4187), .ZN(n2831) );
  INV_X1 U3193 ( .A(n2923), .ZN(n2924) );
  NAND2_X1 U3194 ( .A1(n3774), .A2(REG3_REG_25__SCAN_IN), .ZN(n3791) );
  OR2_X1 U3195 ( .A1(n3762), .A2(n4781), .ZN(n3775) );
  INV_X1 U3196 ( .A(n4419), .ZN(n4204) );
  INV_X1 U3197 ( .A(n3859), .ZN(n3637) );
  INV_X1 U3198 ( .A(n4999), .ZN(n3315) );
  INV_X1 U3199 ( .A(n4282), .ZN(n4228) );
  INV_X1 U3200 ( .A(n5260), .ZN(n5265) );
  INV_X1 U3201 ( .A(n3386), .ZN(n3389) );
  INV_X1 U3202 ( .A(n3202), .ZN(n4083) );
  INV_X1 U3203 ( .A(n4921), .ZN(n4114) );
  INV_X1 U3204 ( .A(IR_REG_23__SCAN_IN), .ZN(n4830) );
  AND2_X1 U3205 ( .A1(n3410), .A2(n3411), .ZN(n3409) );
  AND2_X1 U3206 ( .A1(n3666), .A2(REG3_REG_18__SCAN_IN), .ZN(n3683) );
  OR2_X1 U3207 ( .A1(n3375), .A2(n2926), .ZN(n5302) );
  OR2_X1 U3208 ( .A1(n3835), .A2(n4248), .ZN(n3826) );
  OR2_X1 U3209 ( .A1(n3835), .A2(n4283), .ZN(n3795) );
  INV_X1 U32100 ( .A(n5266), .ZN(n5365) );
  AND2_X1 U32110 ( .A1(n4064), .A2(DATAI_25_), .ZN(n4292) );
  NAND2_X1 U32120 ( .A1(n4403), .A2(n4204), .ZN(n4205) );
  NAND2_X1 U32130 ( .A1(n4426), .A2(n4425), .ZN(n4424) );
  AND2_X1 U32140 ( .A1(REG3_REG_9__SCAN_IN), .A2(REG3_REG_8__SCAN_IN), .ZN(
        n3332) );
  AND2_X1 U32150 ( .A1(n2926), .A2(n3060), .ZN(n5136) );
  AND2_X1 U32160 ( .A1(n4376), .A2(n4076), .ZN(n4440) );
  INV_X1 U32170 ( .A(n5136), .ZN(n5244) );
  OR2_X1 U32180 ( .A1(n5112), .A2(n5106), .ZN(n4461) );
  INV_X1 U32190 ( .A(IR_REG_25__SCAN_IN), .ZN(n4834) );
  OR2_X1 U32200 ( .A1(n2811), .A2(n2871), .ZN(n2764) );
  AND2_X1 U32210 ( .A1(REG3_REG_3__SCAN_IN), .A2(REG3_REG_4__SCAN_IN), .ZN(
        n3135) );
  NAND2_X1 U32220 ( .A1(n3449), .A2(REG3_REG_13__SCAN_IN), .ZN(n3522) );
  NAND2_X1 U32230 ( .A1(n3366), .A2(REG3_REG_10__SCAN_IN), .ZN(n3436) );
  OR2_X1 U32240 ( .A1(n3035), .A2(n3021), .ZN(n3038) );
  INV_X1 U32250 ( .A(n3208), .ZN(n4455) );
  INV_X2 U32260 ( .A(n3028), .ZN(n4061) );
  OR2_X1 U32270 ( .A1(n3835), .A2(n4346), .ZN(n3736) );
  AND4_X1 U32280 ( .A1(n3674), .A2(n3673), .A3(n3672), .A4(n3671), .ZN(n4444)
         );
  AND4_X1 U32290 ( .A1(n3443), .A2(n3442), .A3(n3441), .A4(n3440), .ZN(n5245)
         );
  INV_X1 U32300 ( .A(n5088), .ZN(n5065) );
  INV_X1 U32310 ( .A(n5374), .ZN(n4450) );
  AND2_X1 U32320 ( .A1(n3333), .A2(n3332), .ZN(n3366) );
  INV_X1 U32330 ( .A(n5138), .ZN(n5268) );
  AND2_X1 U32340 ( .A1(n4247), .A2(n5377), .ZN(n5372) );
  NAND2_X1 U32350 ( .A1(n3020), .A2(n3019), .ZN(n4465) );
  INV_X1 U32360 ( .A(n5333), .ZN(n5377) );
  NAND2_X1 U32370 ( .A1(n2977), .A2(n4919), .ZN(n3018) );
  OR2_X1 U32380 ( .A1(n2812), .A2(n2871), .ZN(n2815) );
  OR2_X1 U32390 ( .A1(n3038), .A2(n3025), .ZN(n5344) );
  NAND4_X1 U32400 ( .A1(n3813), .A2(n3812), .A3(n3811), .A4(n3810), .ZN(n4218)
         );
  INV_X1 U32410 ( .A(n4365), .ZN(n4206) );
  INV_X1 U32420 ( .A(n5245), .ZN(n4156) );
  INV_X1 U32430 ( .A(n5183), .ZN(n4160) );
  CLKBUF_X2 U32440 ( .A(U4043), .Z(n5082) );
  NOR2_X1 U32450 ( .A1(n2947), .A2(n2946), .ZN(n2948) );
  INV_X1 U32460 ( .A(n4437), .ZN(n4399) );
  NAND2_X1 U32470 ( .A1(n3196), .A2(n5231), .ZN(n5226) );
  OR2_X1 U32480 ( .A1(n4505), .A2(n4465), .ZN(n5379) );
  AND2_X1 U32490 ( .A1(n5270), .A2(n5272), .ZN(n5271) );
  OR2_X1 U32500 ( .A1(n4505), .A2(n4504), .ZN(n5380) );
  NOR2_X1 U32510 ( .A1(n3129), .A2(n2951), .ZN(U4043) );
  INV_X2 U32520 ( .A(STATE_REG_SCAN_IN), .ZN(U3149) );
  NAND2_X1 U32530 ( .A1(n2769), .A2(n4800), .ZN(n2765) );
  INV_X1 U32540 ( .A(n2765), .ZN(n2755) );
  NAND2_X1 U32550 ( .A1(n2760), .A2(IR_REG_31__SCAN_IN), .ZN(n2761) );
  XNOR2_X1 U32560 ( .A(n2761), .B(IR_REG_13__SCAN_IN), .ZN(n5030) );
  INV_X1 U32570 ( .A(REG1_REG_8__SCAN_IN), .ZN(n5205) );
  INV_X1 U32580 ( .A(IR_REG_7__SCAN_IN), .ZN(n4806) );
  NAND2_X1 U32590 ( .A1(n2764), .A2(n4806), .ZN(n2762) );
  NAND2_X1 U32600 ( .A1(n2762), .A2(IR_REG_31__SCAN_IN), .ZN(n2763) );
  XNOR2_X1 U32610 ( .A(n2763), .B(IR_REG_8__SCAN_IN), .ZN(n4999) );
  NOR2_X1 U32620 ( .A1(n2769), .A2(n2871), .ZN(n2766) );
  INV_X1 U32630 ( .A(n2769), .ZN(n2775) );
  NAND2_X1 U32640 ( .A1(IR_REG_0__SCAN_IN), .A2(IR_REG_31__SCAN_IN), .ZN(n2770) );
  NAND2_X1 U32650 ( .A1(n2770), .A2(IR_REG_1__SCAN_IN), .ZN(n2773) );
  NAND2_X1 U32660 ( .A1(n2771), .A2(IR_REG_31__SCAN_IN), .ZN(n2772) );
  INV_X1 U32670 ( .A(IR_REG_0__SCAN_IN), .ZN(n5078) );
  INV_X1 U32680 ( .A(REG1_REG_0__SCAN_IN), .ZN(n5107) );
  INV_X1 U32690 ( .A(REG1_REG_1__SCAN_IN), .ZN(n2776) );
  NOR3_X1 U32700 ( .A1(n5078), .A2(n5107), .A3(n4965), .ZN(n4963) );
  AOI21_X1 U32710 ( .B1(n2891), .B2(REG1_REG_1__SCAN_IN), .A(n4963), .ZN(n5062) );
  INV_X1 U32720 ( .A(REG1_REG_2__SCAN_IN), .ZN(n3055) );
  MUX2_X1 U32730 ( .A(n3055), .B(REG1_REG_2__SCAN_IN), .S(n4926), .Z(n5063) );
  NAND2_X1 U32740 ( .A1(n2765), .A2(IR_REG_31__SCAN_IN), .ZN(n2779) );
  NAND2_X1 U32750 ( .A1(n2779), .A2(n2778), .ZN(n2783) );
  OR2_X1 U32760 ( .A1(n2779), .A2(n2778), .ZN(n2780) );
  NAND2_X1 U32770 ( .A1(n2783), .A2(n2780), .ZN(n3099) );
  INV_X1 U32780 ( .A(REG1_REG_3__SCAN_IN), .ZN(n5144) );
  NOR2_X1 U32790 ( .A1(n2781), .A2(n3099), .ZN(n2782) );
  NAND2_X1 U32800 ( .A1(n2783), .A2(IR_REG_31__SCAN_IN), .ZN(n2784) );
  XNOR2_X1 U32810 ( .A(n2784), .B(n4607), .ZN(n5154) );
  NOR2_X1 U32820 ( .A1(n2785), .A2(n5154), .ZN(n2786) );
  INV_X1 U32830 ( .A(REG1_REG_4__SCAN_IN), .ZN(n5158) );
  NAND2_X1 U32840 ( .A1(n2787), .A2(IR_REG_31__SCAN_IN), .ZN(n2788) );
  NAND2_X1 U32850 ( .A1(REG1_REG_5__SCAN_IN), .A2(n4979), .ZN(n2789) );
  OAI21_X1 U32860 ( .B1(n4979), .B2(REG1_REG_5__SCAN_IN), .A(n2789), .ZN(n4973) );
  OR2_X1 U32870 ( .A1(n2791), .A2(n2871), .ZN(n2793) );
  XNOR2_X1 U32880 ( .A(n2793), .B(n2792), .ZN(n5163) );
  NOR2_X1 U32890 ( .A1(n2794), .A2(n5163), .ZN(n2795) );
  INV_X1 U32900 ( .A(REG1_REG_6__SCAN_IN), .ZN(n5168) );
  XNOR2_X1 U32910 ( .A(n2794), .B(n5163), .ZN(n3079) );
  NOR2_X1 U32920 ( .A1(n5168), .A2(n3079), .ZN(n3078) );
  NOR2_X1 U32930 ( .A1(n2795), .A2(n3078), .ZN(n4988) );
  NAND2_X1 U32940 ( .A1(n5171), .A2(REG1_REG_7__SCAN_IN), .ZN(n2796) );
  OAI21_X1 U32950 ( .B1(n5171), .B2(REG1_REG_7__SCAN_IN), .A(n2796), .ZN(n4987) );
  NOR2_X1 U32960 ( .A1(n4988), .A2(n4987), .ZN(n4986) );
  NOR2_X1 U32970 ( .A1(n2797), .A2(n3315), .ZN(n2798) );
  NAND2_X1 U32980 ( .A1(n2811), .A2(n2799), .ZN(n2800) );
  NAND2_X1 U32990 ( .A1(n2800), .A2(IR_REG_31__SCAN_IN), .ZN(n2801) );
  NAND2_X1 U33000 ( .A1(n5010), .A2(REG1_REG_9__SCAN_IN), .ZN(n2802) );
  OAI21_X1 U33010 ( .B1(n5010), .B2(REG1_REG_9__SCAN_IN), .A(n2802), .ZN(n5007) );
  AND2_X1 U33020 ( .A1(n5010), .A2(REG1_REG_9__SCAN_IN), .ZN(n2803) );
  NAND2_X1 U33030 ( .A1(n2811), .A2(n2804), .ZN(n2805) );
  NAND2_X1 U33040 ( .A1(n2805), .A2(IR_REG_31__SCAN_IN), .ZN(n2806) );
  XNOR2_X1 U33050 ( .A(n2806), .B(n2757), .ZN(n3483) );
  XNOR2_X1 U33060 ( .A(n2807), .B(n3401), .ZN(n3479) );
  INV_X1 U33070 ( .A(REG1_REG_10__SCAN_IN), .ZN(n5237) );
  NOR2_X1 U33080 ( .A1(n3479), .A2(n5237), .ZN(n3480) );
  INV_X1 U33090 ( .A(n2807), .ZN(n2808) );
  NOR2_X1 U33100 ( .A1(n2808), .A2(n3483), .ZN(n2809) );
  AND2_X1 U33110 ( .A1(n2811), .A2(n2810), .ZN(n2812) );
  NAND2_X1 U33120 ( .A1(n5021), .A2(REG1_REG_11__SCAN_IN), .ZN(n2813) );
  OAI21_X1 U33130 ( .B1(n5021), .B2(REG1_REG_11__SCAN_IN), .A(n2813), .ZN(
        n5017) );
  INV_X1 U33140 ( .A(IR_REG_11__SCAN_IN), .ZN(n2814) );
  NAND2_X1 U33150 ( .A1(n2815), .A2(n2814), .ZN(n2816) );
  NAND2_X1 U33160 ( .A1(n2816), .A2(IR_REG_31__SCAN_IN), .ZN(n2817) );
  INV_X1 U33170 ( .A(IR_REG_12__SCAN_IN), .ZN(n4813) );
  XNOR2_X1 U33180 ( .A(n2817), .B(n4813), .ZN(n3626) );
  INV_X1 U33190 ( .A(REG1_REG_12__SCAN_IN), .ZN(n5288) );
  INV_X1 U33200 ( .A(n2819), .ZN(n2820) );
  NOR2_X1 U33210 ( .A1(n2820), .A2(n3626), .ZN(n2821) );
  NOR2_X1 U33220 ( .A1(n3622), .A2(n2821), .ZN(n5026) );
  XNOR2_X1 U33230 ( .A(n5030), .B(REG1_REG_13__SCAN_IN), .ZN(n5025) );
  XNOR2_X1 U33240 ( .A(n2837), .B(IR_REG_14__SCAN_IN), .ZN(n5042) );
  INV_X1 U33250 ( .A(n5042), .ZN(n2956) );
  NAND2_X1 U33260 ( .A1(n2822), .A2(n2956), .ZN(n2823) );
  NAND2_X1 U33270 ( .A1(n2824), .A2(n2823), .ZN(n5039) );
  INV_X1 U33280 ( .A(REG1_REG_14__SCAN_IN), .ZN(n5300) );
  NOR2_X1 U33290 ( .A1(n5038), .A2(n2825), .ZN(n4167) );
  NAND2_X1 U33300 ( .A1(n2837), .A2(n2835), .ZN(n2826) );
  NAND2_X1 U33310 ( .A1(n2826), .A2(IR_REG_31__SCAN_IN), .ZN(n2828) );
  XNOR2_X1 U33320 ( .A(n2828), .B(IR_REG_15__SCAN_IN), .ZN(n4924) );
  INV_X1 U33330 ( .A(n4924), .ZN(n4171) );
  INV_X1 U33340 ( .A(REG1_REG_15__SCAN_IN), .ZN(n5324) );
  AOI22_X1 U33350 ( .A1(REG1_REG_15__SCAN_IN), .A2(n4171), .B1(n4924), .B2(
        n5324), .ZN(n4168) );
  NOR2_X1 U33360 ( .A1(n4167), .A2(n4168), .ZN(n4166) );
  NAND2_X1 U33370 ( .A1(n2828), .A2(n2834), .ZN(n2829) );
  NAND2_X1 U33380 ( .A1(n2829), .A2(IR_REG_31__SCAN_IN), .ZN(n2830) );
  XNOR2_X1 U33390 ( .A(n2830), .B(n4623), .ZN(n4187) );
  INV_X1 U33400 ( .A(REG1_REG_16__SCAN_IN), .ZN(n5329) );
  NAND2_X1 U33410 ( .A1(n2832), .A2(n4187), .ZN(n2833) );
  NAND3_X1 U33420 ( .A1(n2835), .A2(n4623), .A3(n2834), .ZN(n2851) );
  NAND2_X1 U33430 ( .A1(n2851), .A2(IR_REG_31__SCAN_IN), .ZN(n2836) );
  OR2_X1 U33440 ( .A1(n2845), .A2(IR_REG_17__SCAN_IN), .ZN(n2840) );
  NAND2_X1 U33450 ( .A1(n2845), .A2(IR_REG_17__SCAN_IN), .ZN(n2838) );
  INV_X1 U33460 ( .A(REG1_REG_17__SCAN_IN), .ZN(n3587) );
  XNOR2_X1 U33470 ( .A(n5048), .B(n3587), .ZN(n5046) );
  NOR2_X1 U33480 ( .A1(n5048), .A2(REG1_REG_17__SCAN_IN), .ZN(n2839) );
  NAND2_X1 U33490 ( .A1(n2840), .A2(IR_REG_31__SCAN_IN), .ZN(n2841) );
  XNOR2_X1 U33500 ( .A(n2841), .B(IR_REG_18__SCAN_IN), .ZN(n4923) );
  OR2_X1 U33510 ( .A1(n4923), .A2(REG1_REG_18__SCAN_IN), .ZN(n2842) );
  NAND2_X1 U33520 ( .A1(n4923), .A2(REG1_REG_18__SCAN_IN), .ZN(n2843) );
  AND2_X1 U3353 ( .A1(n2842), .A2(n2843), .ZN(n2937) );
  NAND2_X1 U33540 ( .A1(n4628), .A2(n4822), .ZN(n2848) );
  AND2_X1 U3355 ( .A1(n2848), .A2(IR_REG_31__SCAN_IN), .ZN(n2844) );
  OR2_X2 U3356 ( .A1(n2845), .A2(n2844), .ZN(n2997) );
  XNOR2_X1 U3357 ( .A(n2997), .B(IR_REG_19__SCAN_IN), .ZN(n3046) );
  XNOR2_X1 U3358 ( .A(n4138), .B(REG1_REG_19__SCAN_IN), .ZN(n2847) );
  INV_X1 U3359 ( .A(n2848), .ZN(n2850) );
  NAND4_X1 U3360 ( .A1(n2850), .A2(n4633), .A3(n2696), .A4(n2849), .ZN(n2852)
         );
  NOR2_X2 U3361 ( .A1(n2883), .A2(IR_REG_25__SCAN_IN), .ZN(n2878) );
  NAND2_X1 U3362 ( .A1(n2878), .A2(n2858), .ZN(n2966) );
  INV_X1 U3363 ( .A(n2865), .ZN(n2860) );
  NOR2_X1 U3364 ( .A1(n2860), .A2(n2859), .ZN(n2864) );
  NAND2_X1 U3365 ( .A1(n2861), .A2(n2878), .ZN(n2881) );
  NAND2_X1 U3366 ( .A1(n2885), .A2(n2867), .ZN(n2868) );
  NAND2_X1 U3367 ( .A1(n2868), .A2(IR_REG_31__SCAN_IN), .ZN(n2869) );
  NAND2_X1 U3368 ( .A1(n2968), .A2(IR_REG_31__SCAN_IN), .ZN(n2870) );
  NAND2_X1 U3369 ( .A1(n4455), .A2(n4921), .ZN(n3210) );
  OR2_X1 U3370 ( .A1(n2873), .A2(n4830), .ZN(n2874) );
  NAND2_X1 U3371 ( .A1(n2873), .A2(n4830), .ZN(n2876) );
  NAND2_X1 U3372 ( .A1(n2874), .A2(n2876), .ZN(n3128) );
  NAND2_X1 U3373 ( .A1(n3060), .A2(n3128), .ZN(n2875) );
  AND2_X1 U3374 ( .A1(n4064), .A2(n2875), .ZN(n2929) );
  NAND2_X1 U3375 ( .A1(n2876), .A2(IR_REG_31__SCAN_IN), .ZN(n2877) );
  NAND2_X1 U3376 ( .A1(n2878), .A2(n2885), .ZN(n2879) );
  NAND2_X1 U3377 ( .A1(n2879), .A2(IR_REG_31__SCAN_IN), .ZN(n2880) );
  NAND2_X1 U3378 ( .A1(n2885), .A2(n2884), .ZN(n2886) );
  INV_X1 U3379 ( .A(n2978), .ZN(n4920) );
  INV_X1 U3380 ( .A(n3037), .ZN(n3021) );
  INV_X1 U3381 ( .A(n3128), .ZN(n2888) );
  NAND2_X1 U3382 ( .A1(n2888), .A2(STATE_REG_SCAN_IN), .ZN(n4149) );
  NAND2_X1 U3383 ( .A1(n3021), .A2(n4149), .ZN(n2928) );
  NAND2_X1 U3384 ( .A1(n2929), .A2(n2928), .ZN(n4958) );
  INV_X1 U3385 ( .A(n5071), .ZN(n4954) );
  NAND2_X1 U3386 ( .A1(IR_REG_0__SCAN_IN), .A2(REG2_REG_0__SCAN_IN), .ZN(n5075) );
  INV_X1 U3387 ( .A(REG2_REG_1__SCAN_IN), .ZN(n2890) );
  NOR2_X1 U3388 ( .A1(n5075), .A2(n4961), .ZN(n4960) );
  NOR2_X1 U3389 ( .A1(n4960), .A2(n2523), .ZN(n5057) );
  INV_X1 U3390 ( .A(n4926), .ZN(n5068) );
  INV_X1 U3391 ( .A(REG2_REG_2__SCAN_IN), .ZN(n2892) );
  AOI22_X1 U3392 ( .A1(REG2_REG_2__SCAN_IN), .A2(n5068), .B1(n4926), .B2(n2892), .ZN(n5058) );
  NOR2_X1 U3393 ( .A1(n5057), .A2(n5058), .ZN(n5056) );
  AND2_X1 U3394 ( .A1(n4926), .A2(REG2_REG_2__SCAN_IN), .ZN(n2893) );
  XNOR2_X1 U3395 ( .A(n2894), .B(n3099), .ZN(n3066) );
  INV_X1 U3396 ( .A(REG2_REG_3__SCAN_IN), .ZN(n3068) );
  NOR2_X1 U3397 ( .A1(n2894), .A2(n3099), .ZN(n2895) );
  NOR2_X1 U3398 ( .A1(n2896), .A2(n5154), .ZN(n2897) );
  INV_X1 U3399 ( .A(REG2_REG_4__SCAN_IN), .ZN(n5094) );
  XNOR2_X1 U3400 ( .A(n2896), .B(n5154), .ZN(n5093) );
  NAND2_X1 U3401 ( .A1(REG2_REG_5__SCAN_IN), .A2(n4979), .ZN(n2898) );
  OAI21_X1 U3402 ( .B1(REG2_REG_5__SCAN_IN), .B2(n4979), .A(n2898), .ZN(n4977)
         );
  NOR2_X1 U3403 ( .A1(n2899), .A2(n5163), .ZN(n2900) );
  INV_X1 U3404 ( .A(REG2_REG_6__SCAN_IN), .ZN(n3287) );
  XNOR2_X1 U3405 ( .A(n5163), .B(n2899), .ZN(n3076) );
  NAND2_X1 U3406 ( .A1(n5171), .A2(REG2_REG_7__SCAN_IN), .ZN(n2901) );
  OAI21_X1 U3407 ( .B1(n5171), .B2(REG2_REG_7__SCAN_IN), .A(n2901), .ZN(n4983)
         );
  INV_X1 U3408 ( .A(n2903), .ZN(n2902) );
  NOR2_X1 U3409 ( .A1(n2902), .A2(n3315), .ZN(n2904) );
  INV_X1 U3410 ( .A(REG2_REG_8__SCAN_IN), .ZN(n4995) );
  NOR2_X1 U3411 ( .A1(n2904), .A2(n4994), .ZN(n5005) );
  NAND2_X1 U3412 ( .A1(n5010), .A2(REG2_REG_9__SCAN_IN), .ZN(n2905) );
  OAI21_X1 U3413 ( .B1(n5010), .B2(REG2_REG_9__SCAN_IN), .A(n2905), .ZN(n5004)
         );
  NOR2_X1 U3414 ( .A1(n5005), .A2(n5004), .ZN(n5003) );
  INV_X1 U3415 ( .A(REG2_REG_10__SCAN_IN), .ZN(n3486) );
  NOR2_X1 U3416 ( .A1(n2907), .A2(n3483), .ZN(n2908) );
  NAND2_X1 U3417 ( .A1(n5021), .A2(REG2_REG_11__SCAN_IN), .ZN(n2909) );
  OAI21_X1 U3418 ( .B1(n5021), .B2(REG2_REG_11__SCAN_IN), .A(n2909), .ZN(n5015) );
  XNOR2_X1 U3419 ( .A(n2910), .B(n3626), .ZN(n3628) );
  INV_X1 U3420 ( .A(REG2_REG_12__SCAN_IN), .ZN(n3629) );
  XNOR2_X1 U3421 ( .A(n5030), .B(REG2_REG_13__SCAN_IN), .ZN(n5029) );
  NAND2_X1 U3422 ( .A1(n5030), .A2(REG2_REG_13__SCAN_IN), .ZN(n2911) );
  INV_X1 U3423 ( .A(n2915), .ZN(n2914) );
  OR2_X1 U3424 ( .A1(n2912), .A2(n5042), .ZN(n2913) );
  INV_X1 U3425 ( .A(REG2_REG_14__SCAN_IN), .ZN(n5036) );
  AOI22_X1 U3426 ( .A1(REG2_REG_15__SCAN_IN), .A2(n4171), .B1(n4924), .B2(
        n3617), .ZN(n4173) );
  XNOR2_X1 U3427 ( .A(n2917), .B(n2831), .ZN(n4182) );
  INV_X1 U3428 ( .A(REG2_REG_16__SCAN_IN), .ZN(n4181) );
  NAND2_X1 U3429 ( .A1(n2917), .A2(n4187), .ZN(n2918) );
  NAND2_X1 U3430 ( .A1(n5048), .A2(REG2_REG_17__SCAN_IN), .ZN(n2919) );
  OAI21_X1 U3431 ( .B1(n5048), .B2(REG2_REG_17__SCAN_IN), .A(n2919), .ZN(n5051) );
  NAND2_X1 U3432 ( .A1(REG2_REG_18__SCAN_IN), .A2(n4923), .ZN(n2920) );
  OAI21_X1 U3433 ( .B1(REG2_REG_18__SCAN_IN), .B2(n4923), .A(n2920), .ZN(n2940) );
  INV_X1 U3434 ( .A(REG2_REG_19__SCAN_IN), .ZN(n2922) );
  MUX2_X1 U3435 ( .A(REG2_REG_19__SCAN_IN), .B(n2922), .S(n4138), .Z(n2923) );
  XNOR2_X1 U3436 ( .A(n2925), .B(n2924), .ZN(n2927) );
  INV_X1 U3437 ( .A(n2926), .ZN(n5072) );
  NAND2_X1 U3438 ( .A1(n5072), .A2(n4954), .ZN(n5074) );
  INV_X1 U3439 ( .A(n5091), .ZN(n5060) );
  NAND2_X1 U3440 ( .A1(n2927), .A2(n5060), .ZN(n2934) );
  INV_X1 U3441 ( .A(n2928), .ZN(n2930) );
  NOR2_X2 U3442 ( .A1(n2930), .A2(n2929), .ZN(n5087) );
  NAND2_X1 U3443 ( .A1(n5087), .A2(ADDR_REG_19__SCAN_IN), .ZN(n2931) );
  NAND2_X1 U3444 ( .A1(U3149), .A2(REG3_REG_19__SCAN_IN), .ZN(n3882) );
  OAI211_X1 U3445 ( .C1(n4138), .C2(n5069), .A(n2931), .B(n3882), .ZN(n2932)
         );
  INV_X1 U3446 ( .A(n2932), .ZN(n2933) );
  OAI211_X1 U3447 ( .C1(n2938), .C2(n2937), .A(n2936), .B(n5065), .ZN(n2950)
         );
  NAND2_X1 U3448 ( .A1(n2939), .A2(n2940), .ZN(n2943) );
  NOR2_X1 U3449 ( .A1(n5091), .A2(n2941), .ZN(n2942) );
  NAND2_X1 U3450 ( .A1(n2943), .A2(n2942), .ZN(n2949) );
  AOI22_X1 U3451 ( .A1(REG3_REG_18__SCAN_IN), .A2(U3149), .B1(n5087), .B2(
        ADDR_REG_18__SCAN_IN), .ZN(n2944) );
  INV_X1 U3452 ( .A(n2944), .ZN(n2947) );
  INV_X1 U3453 ( .A(n4923), .ZN(n2945) );
  NOR2_X1 U3454 ( .A1(n5069), .A2(n2945), .ZN(n2946) );
  NAND3_X1 U3455 ( .A1(n2950), .A2(n2949), .A3(n2948), .ZN(U3258) );
  INV_X1 U3456 ( .A(n2984), .ZN(n2951) );
  INV_X1 U3457 ( .A(DATAI_10_), .ZN(n2952) );
  MUX2_X1 U34580 ( .A(n3483), .B(n2952), .S(U3149), .Z(n2953) );
  INV_X1 U34590 ( .A(n2953), .ZN(U3342) );
  INV_X1 U3460 ( .A(DATAI_12_), .ZN(n2954) );
  MUX2_X1 U3461 ( .A(n3626), .B(n2954), .S(U3149), .Z(n2955) );
  INV_X1 U3462 ( .A(n2955), .ZN(U3340) );
  INV_X1 U3463 ( .A(DATAI_14_), .ZN(n2957) );
  MUX2_X1 U3464 ( .A(n2957), .B(n2956), .S(STATE_REG_SCAN_IN), .Z(n2958) );
  INV_X1 U3465 ( .A(n2958), .ZN(U3338) );
  INV_X1 U3466 ( .A(DATAI_23_), .ZN(n2959) );
  AOI21_X1 U34670 ( .B1(U3149), .B2(n2959), .A(n2984), .ZN(U3329) );
  INV_X1 U3468 ( .A(DATAI_22_), .ZN(n2960) );
  MUX2_X1 U34690 ( .A(n3208), .B(n2960), .S(U3149), .Z(n2961) );
  INV_X1 U3470 ( .A(n2961), .ZN(U3330) );
  INV_X1 U34710 ( .A(DATAI_28_), .ZN(n2962) );
  MUX2_X1 U3472 ( .A(n2962), .B(n2926), .S(STATE_REG_SCAN_IN), .Z(n2963) );
  INV_X1 U34730 ( .A(n2963), .ZN(U3324) );
  INV_X1 U3474 ( .A(DATAI_16_), .ZN(n2964) );
  MUX2_X1 U34750 ( .A(n2964), .B(n4187), .S(STATE_REG_SCAN_IN), .Z(n2965) );
  INV_X1 U3476 ( .A(n2965), .ZN(U3336) );
  INV_X1 U34770 ( .A(DATAI_30_), .ZN(n2971) );
  NAND2_X1 U3478 ( .A1(n2986), .A2(n4843), .ZN(n4916) );
  MUX2_X1 U34790 ( .A(n2971), .B(n2992), .S(STATE_REG_SCAN_IN), .Z(n2972) );
  INV_X1 U3480 ( .A(n2972), .ZN(U3322) );
  INV_X1 U34810 ( .A(DATAI_19_), .ZN(n2973) );
  MUX2_X1 U3482 ( .A(n4138), .B(n2973), .S(U3149), .Z(n2974) );
  INV_X1 U34830 ( .A(n2974), .ZN(U3333) );
  NAND2_X1 U3484 ( .A1(n2978), .A2(B_REG_SCAN_IN), .ZN(n2976) );
  MUX2_X1 U34850 ( .A(n2976), .B(B_REG_SCAN_IN), .S(n2975), .Z(n2977) );
  NAND2_X1 U3486 ( .A1(n3037), .A2(n3018), .ZN(n4951) );
  INV_X1 U34870 ( .A(D_REG_1__SCAN_IN), .ZN(n2980) );
  INV_X1 U3488 ( .A(n4919), .ZN(n2982) );
  NAND2_X1 U34890 ( .A1(n2982), .A2(n2978), .ZN(n3015) );
  INV_X1 U3490 ( .A(n3015), .ZN(n2979) );
  AOI22_X1 U34910 ( .A1(n4951), .A2(n2980), .B1(n2984), .B2(n2979), .ZN(U3459)
         );
  INV_X1 U3492 ( .A(D_REG_0__SCAN_IN), .ZN(n2985) );
  INV_X1 U34930 ( .A(n2975), .ZN(n2981) );
  NAND2_X1 U3494 ( .A1(n2982), .A2(n2981), .ZN(n3019) );
  INV_X1 U34950 ( .A(n3019), .ZN(n2983) );
  AOI22_X1 U3496 ( .A1(n4951), .A2(n2985), .B1(n2984), .B2(n2983), .ZN(U3458)
         );
  NOR2_X1 U34970 ( .A1(n5087), .A2(n5082), .ZN(U3148) );
  INV_X1 U3498 ( .A(n3129), .ZN(n3001) );
  INV_X1 U34990 ( .A(REG0_REG_0__SCAN_IN), .ZN(n5108) );
  OR2_X1 U3500 ( .A1(n3094), .A2(n5108), .ZN(n2996) );
  INV_X1 U35010 ( .A(REG3_REG_0__SCAN_IN), .ZN(n2988) );
  OR2_X1 U3502 ( .A1(n3054), .A2(n2988), .ZN(n2995) );
  NAND2_X2 U35030 ( .A1(n2990), .A2(n2989), .ZN(n3026) );
  INV_X1 U3504 ( .A(REG2_REG_0__SCAN_IN), .ZN(n2991) );
  OR2_X1 U35050 ( .A1(n3136), .A2(n5107), .ZN(n2993) );
  INV_X1 U35060 ( .A(n4165), .ZN(n3186) );
  MUX2_X1 U35070 ( .A(IR_REG_0__SCAN_IN), .B(DATAI_0_), .S(n3107), .Z(n3227)
         );
  OAI22_X1 U35080 ( .A1(n3186), .A2(n2511), .B1(n3108), .B2(n5105), .ZN(n3050)
         );
  INV_X1 U35090 ( .A(n3108), .ZN(n3000) );
  INV_X1 U35100 ( .A(n5106), .ZN(n2999) );
  NAND2_X1 U35110 ( .A1(n3752), .A2(n4165), .ZN(n3003) );
  XNOR2_X1 U35120 ( .A(n3052), .B(n3051), .ZN(n5073) );
  NOR4_X1 U35130 ( .A1(D_REG_13__SCAN_IN), .A2(D_REG_15__SCAN_IN), .A3(
        D_REG_16__SCAN_IN), .A4(D_REG_18__SCAN_IN), .ZN(n3004) );
  INV_X1 U35140 ( .A(D_REG_7__SCAN_IN), .ZN(n4932) );
  INV_X1 U35150 ( .A(D_REG_5__SCAN_IN), .ZN(n4930) );
  NAND3_X1 U35160 ( .A1(n3004), .A2(n4932), .A3(n4930), .ZN(n3010) );
  NOR4_X1 U35170 ( .A1(D_REG_12__SCAN_IN), .A2(D_REG_11__SCAN_IN), .A3(
        D_REG_8__SCAN_IN), .A4(D_REG_2__SCAN_IN), .ZN(n3008) );
  NOR4_X1 U35180 ( .A1(D_REG_21__SCAN_IN), .A2(D_REG_27__SCAN_IN), .A3(
        D_REG_25__SCAN_IN), .A4(D_REG_19__SCAN_IN), .ZN(n3007) );
  NOR4_X1 U35190 ( .A1(D_REG_31__SCAN_IN), .A2(D_REG_30__SCAN_IN), .A3(
        D_REG_29__SCAN_IN), .A4(D_REG_14__SCAN_IN), .ZN(n3006) );
  NOR4_X1 U35200 ( .A1(D_REG_20__SCAN_IN), .A2(D_REG_23__SCAN_IN), .A3(
        D_REG_28__SCAN_IN), .A4(D_REG_26__SCAN_IN), .ZN(n3005) );
  NAND4_X1 U35210 ( .A1(n3008), .A2(n3007), .A3(n3006), .A4(n3005), .ZN(n3009)
         );
  NOR4_X1 U35220 ( .A1(D_REG_6__SCAN_IN), .A2(D_REG_10__SCAN_IN), .A3(n3010), 
        .A4(n3009), .ZN(n3013) );
  INV_X1 U35230 ( .A(D_REG_3__SCAN_IN), .ZN(n4928) );
  INV_X1 U35240 ( .A(D_REG_4__SCAN_IN), .ZN(n4929) );
  INV_X1 U35250 ( .A(D_REG_17__SCAN_IN), .ZN(n4941) );
  INV_X1 U35260 ( .A(D_REG_9__SCAN_IN), .ZN(n4934) );
  NAND4_X1 U35270 ( .A1(n4928), .A2(n4929), .A3(n4941), .A4(n4934), .ZN(n3011)
         );
  NOR3_X1 U35280 ( .A1(D_REG_24__SCAN_IN), .A2(D_REG_22__SCAN_IN), .A3(n3011), 
        .ZN(n3012) );
  AND2_X1 U35290 ( .A1(n3013), .A2(n3012), .ZN(n3014) );
  INV_X1 U35300 ( .A(n4462), .ZN(n3017) );
  OR2_X1 U35310 ( .A1(n3018), .A2(D_REG_1__SCAN_IN), .ZN(n3016) );
  NAND2_X1 U35320 ( .A1(n3016), .A2(n3015), .ZN(n4464) );
  NOR2_X1 U35330 ( .A1(n3017), .A2(n4464), .ZN(n3195) );
  NAND2_X1 U35340 ( .A1(n3195), .A2(n4504), .ZN(n3035) );
  OAI21_X1 U35350 ( .B1(n5106), .B2(n4138), .A(n3210), .ZN(n3022) );
  INV_X1 U35360 ( .A(n3022), .ZN(n3024) );
  AND2_X1 U35370 ( .A1(n3024), .A2(n5266), .ZN(n3033) );
  INV_X1 U35380 ( .A(n3033), .ZN(n3025) );
  NAND2_X1 U35390 ( .A1(n3023), .A2(n4138), .ZN(n4117) );
  NAND2_X1 U35400 ( .A1(n4117), .A2(n3060), .ZN(n3127) );
  NAND2_X1 U35410 ( .A1(n4463), .A2(n3060), .ZN(n4146) );
  INV_X1 U35420 ( .A(n3026), .ZN(n3053) );
  NAND2_X1 U35430 ( .A1(n3053), .A2(REG2_REG_1__SCAN_IN), .ZN(n3032) );
  INV_X1 U35440 ( .A(REG3_REG_1__SCAN_IN), .ZN(n3229) );
  OR2_X1 U35450 ( .A1(n3054), .A2(n3229), .ZN(n3031) );
  INV_X1 U35460 ( .A(n3094), .ZN(n3027) );
  NAND2_X1 U35470 ( .A1(n3027), .A2(REG0_REG_1__SCAN_IN), .ZN(n3030) );
  INV_X1 U35480 ( .A(n3136), .ZN(n3028) );
  NAND2_X1 U35490 ( .A1(n3035), .A2(n3033), .ZN(n3130) );
  OAI21_X1 U35500 ( .B1(n5266), .B2(U3149), .A(n4146), .ZN(n3034) );
  NAND2_X1 U35510 ( .A1(n3035), .A2(n3034), .ZN(n3132) );
  NAND3_X1 U35520 ( .A1(n3130), .A2(n3132), .A3(n4463), .ZN(n3970) );
  AOI22_X1 U35530 ( .A1(n5309), .A2(n5103), .B1(n3970), .B2(
        REG3_REG_0__SCAN_IN), .ZN(n3040) );
  NAND2_X1 U35540 ( .A1(n3023), .A2(n2846), .ZN(n5112) );
  NAND2_X2 U35550 ( .A1(n3037), .A2(n3036), .ZN(n5231) );
  NAND2_X1 U35560 ( .A1(n3972), .A2(n3227), .ZN(n3039) );
  OAI211_X1 U35570 ( .C1(n5073), .C2(n5344), .A(n3040), .B(n3039), .ZN(U3229)
         );
  OR2_X1 U35580 ( .A1(n3185), .A2(n3110), .ZN(n3045) );
  NAND2_X1 U35590 ( .A1(n3184), .A2(n3740), .ZN(n3044) );
  NAND2_X1 U35600 ( .A1(n3045), .A2(n3044), .ZN(n3117) );
  INV_X1 U35610 ( .A(n3117), .ZN(n3049) );
  OAI22_X1 U35620 ( .A1(n3185), .A2(n2511), .B1(n3108), .B2(n3222), .ZN(n3048)
         );
  NAND2_X1 U35630 ( .A1(n4455), .A2(n3046), .ZN(n3047) );
  OAI22_X1 U35640 ( .A1(n3052), .A2(n3051), .B1(n3829), .B2(n3050), .ZN(n3118)
         );
  XNOR2_X1 U35650 ( .A(n3119), .B(n3118), .ZN(n3065) );
  NAND2_X1 U35660 ( .A1(n3053), .A2(REG2_REG_2__SCAN_IN), .ZN(n3059) );
  INV_X1 U35670 ( .A(REG3_REG_2__SCAN_IN), .ZN(n3257) );
  OR2_X1 U35680 ( .A1(n3136), .A2(n3055), .ZN(n3056) );
  OR2_X1 U35690 ( .A1(n5133), .A2(n5244), .ZN(n3062) );
  NAND2_X1 U35700 ( .A1(n4165), .A2(n5180), .ZN(n3061) );
  NAND2_X1 U35710 ( .A1(n3062), .A2(n3061), .ZN(n3223) );
  INV_X1 U35720 ( .A(n3375), .ZN(n5348) );
  AOI22_X1 U35730 ( .A1(n3223), .A2(n5348), .B1(REG3_REG_1__SCAN_IN), .B2(
        n3970), .ZN(n3064) );
  NAND2_X1 U35740 ( .A1(n3972), .A2(n3184), .ZN(n3063) );
  OAI211_X1 U35750 ( .C1(n3065), .C2(n5344), .A(n3064), .B(n3063), .ZN(U3219)
         );
  AOI21_X1 U35760 ( .B1(n3068), .B2(n3066), .A(n3067), .ZN(n3072) );
  AOI211_X1 U35770 ( .C1(n3070), .C2(n5144), .A(n3069), .B(n5088), .ZN(n3071)
         );
  AOI21_X1 U35780 ( .B1(n5060), .B2(n3072), .A(n3071), .ZN(n3074) );
  INV_X1 U35790 ( .A(REG3_REG_3__SCAN_IN), .ZN(n5146) );
  NOR2_X1 U35800 ( .A1(STATE_REG_SCAN_IN), .A2(n5146), .ZN(n3351) );
  AOI21_X1 U35810 ( .B1(n5087), .B2(ADDR_REG_3__SCAN_IN), .A(n3351), .ZN(n3073) );
  OAI211_X1 U3582 ( .C1(n3099), .C2(n5069), .A(n3074), .B(n3073), .ZN(U3243)
         );
  AOI21_X1 U3583 ( .B1(n3287), .B2(n3076), .A(n3075), .ZN(n3082) );
  AND2_X1 U3584 ( .A1(U3149), .A2(REG3_REG_6__SCAN_IN), .ZN(n3177) );
  AOI21_X1 U3585 ( .B1(n5087), .B2(ADDR_REG_6__SCAN_IN), .A(n3177), .ZN(n3077)
         );
  OAI21_X1 U3586 ( .B1(n5163), .B2(n5069), .A(n3077), .ZN(n3081) );
  AOI211_X1 U3587 ( .C1(n3079), .C2(n5168), .A(n3078), .B(n5088), .ZN(n3080)
         );
  AOI211_X1 U3588 ( .C1(n3082), .C2(n5060), .A(n3081), .B(n3080), .ZN(n3083)
         );
  INV_X1 U3589 ( .A(n3083), .ZN(U3246) );
  NAND2_X1 U3590 ( .A1(n4052), .A2(REG2_REG_4__SCAN_IN), .ZN(n3090) );
  OR2_X1 U3591 ( .A1(n3136), .A2(n5158), .ZN(n3089) );
  INV_X1 U3592 ( .A(n3135), .ZN(n3086) );
  INV_X1 U3593 ( .A(REG3_REG_4__SCAN_IN), .ZN(n3084) );
  NAND2_X1 U3594 ( .A1(n5146), .A2(n3084), .ZN(n3085) );
  NAND2_X1 U3595 ( .A1(n3086), .A2(n3085), .ZN(n3198) );
  OR2_X1 U3596 ( .A1(n3835), .A2(n3198), .ZN(n3088) );
  INV_X1 U3597 ( .A(REG0_REG_4__SCAN_IN), .ZN(n4898) );
  OR2_X1 U3598 ( .A1(n2513), .A2(n4898), .ZN(n3087) );
  INV_X1 U3599 ( .A(n5154), .ZN(n5097) );
  MUX2_X1 U3600 ( .A(n5097), .B(DATAI_4_), .S(n4064), .Z(n3240) );
  INV_X1 U3601 ( .A(n3240), .ZN(n3191) );
  OAI22_X1 U3602 ( .A1(n3189), .A2(n3798), .B1(n3108), .B2(n3191), .ZN(n3091)
         );
  XNOR2_X1 U3603 ( .A(n3091), .B(n3782), .ZN(n3163) );
  OR2_X1 U3604 ( .A1(n3189), .A2(n3800), .ZN(n3093) );
  INV_X2 U3605 ( .A(n2511), .ZN(n3293) );
  NAND2_X1 U3606 ( .A1(n3240), .A2(n3293), .ZN(n3092) );
  NAND2_X1 U3607 ( .A1(n3093), .A2(n3092), .ZN(n3164) );
  XNOR2_X1 U3608 ( .A(n3163), .B(n3164), .ZN(n3123) );
  NAND2_X1 U3609 ( .A1(n4052), .A2(REG2_REG_3__SCAN_IN), .ZN(n3098) );
  OR2_X1 U3610 ( .A1(n3136), .A2(n5144), .ZN(n3097) );
  INV_X1 U3611 ( .A(REG0_REG_3__SCAN_IN), .ZN(n4899) );
  OR2_X1 U3612 ( .A1(n2513), .A2(n4899), .ZN(n3096) );
  OR2_X1 U3613 ( .A1(n3054), .A2(REG3_REG_3__SCAN_IN), .ZN(n3095) );
  NAND2_X1 U3614 ( .A1(n4163), .A2(n3740), .ZN(n3101) );
  INV_X1 U3615 ( .A(n3099), .ZN(n4925) );
  MUX2_X1 U3616 ( .A(n4925), .B(DATAI_3_), .S(n4064), .Z(n3350) );
  NAND2_X1 U3617 ( .A1(n3350), .A2(n3815), .ZN(n3100) );
  NAND2_X1 U3618 ( .A1(n3101), .A2(n3100), .ZN(n3102) );
  INV_X1 U3619 ( .A(n3105), .ZN(n3104) );
  OAI22_X1 U3620 ( .A1(n3251), .A2(n3110), .B1(n2511), .B2(n5132), .ZN(n3103)
         );
  INV_X1 U3621 ( .A(n3103), .ZN(n3106) );
  NAND2_X1 U3622 ( .A1(n3104), .A2(n3106), .ZN(n3124) );
  MUX2_X1 U3623 ( .A(n4926), .B(DATAI_2_), .S(n3107), .Z(n3971) );
  INV_X1 U3624 ( .A(n3971), .ZN(n3204) );
  OAI22_X1 U3625 ( .A1(n3204), .A2(n3108), .B1(n5133), .B2(n2511), .ZN(n3109)
         );
  XNOR2_X1 U3626 ( .A(n3109), .B(n3829), .ZN(n3114) );
  OR2_X1 U3627 ( .A1(n5133), .A2(n3110), .ZN(n3112) );
  NAND2_X1 U3628 ( .A1(n3971), .A2(n3740), .ZN(n3111) );
  NAND2_X1 U3629 ( .A1(n3112), .A2(n3111), .ZN(n3113) );
  AOI22_X1 U3630 ( .A1(n3119), .A2(n3118), .B1(n3117), .B2(n3116), .ZN(n3967)
         );
  AND2_X1 U3631 ( .A1(n3349), .A2(n3345), .ZN(n3120) );
  AOI21_X2 U3632 ( .B1(n3121), .B2(n3967), .A(n3120), .ZN(n3347) );
  INV_X1 U3633 ( .A(n3264), .ZN(n3126) );
  AOI21_X1 U3634 ( .B1(n3347), .B2(n3124), .A(n3123), .ZN(n3125) );
  NOR3_X1 U3635 ( .A1(n3126), .A2(n3125), .A3(n5344), .ZN(n3145) );
  NAND4_X1 U3636 ( .A1(n3130), .A2(n3129), .A3(n3128), .A4(n3127), .ZN(n3131)
         );
  NAND2_X1 U3637 ( .A1(n3131), .A2(STATE_REG_SCAN_IN), .ZN(n3133) );
  AND2_X2 U3638 ( .A1(n3133), .A2(n3132), .ZN(n5354) );
  AOI22_X1 U3639 ( .A1(n3240), .A2(n3972), .B1(n3980), .B2(n4163), .ZN(n3143)
         );
  NAND2_X1 U3640 ( .A1(n4052), .A2(REG2_REG_5__SCAN_IN), .ZN(n3141) );
  INV_X1 U3641 ( .A(REG0_REG_5__SCAN_IN), .ZN(n3134) );
  OR2_X1 U3642 ( .A1(n2513), .A2(n3134), .ZN(n3140) );
  NAND2_X1 U3643 ( .A1(n3135), .A2(REG3_REG_5__SCAN_IN), .ZN(n3147) );
  OAI21_X1 U3644 ( .B1(n3135), .B2(REG3_REG_5__SCAN_IN), .A(n3147), .ZN(n3273)
         );
  OR2_X1 U3645 ( .A1(n3835), .A2(n3273), .ZN(n3139) );
  INV_X1 U3646 ( .A(REG1_REG_5__SCAN_IN), .ZN(n3137) );
  OR2_X1 U3647 ( .A1(n4061), .A2(n3137), .ZN(n3138) );
  AND2_X1 U3648 ( .A1(U3149), .A2(REG3_REG_4__SCAN_IN), .ZN(n5086) );
  AOI21_X1 U3649 ( .B1(n5309), .B2(n4162), .A(n5086), .ZN(n3142) );
  OAI211_X1 U3650 ( .C1(n5354), .C2(n3198), .A(n3143), .B(n3142), .ZN(n3144)
         );
  OR2_X1 U3651 ( .A1(n3145), .A2(n3144), .ZN(U3227) );
  NAND2_X1 U3652 ( .A1(n4052), .A2(REG2_REG_6__SCAN_IN), .ZN(n3152) );
  OR2_X1 U3653 ( .A1(n4061), .A2(n5168), .ZN(n3151) );
  AND2_X1 U3654 ( .A1(n3147), .A2(n3146), .ZN(n3148) );
  OR2_X1 U3655 ( .A1(n3148), .A2(n3171), .ZN(n3286) );
  OR2_X1 U3656 ( .A1(n3835), .A2(n3286), .ZN(n3150) );
  INV_X1 U3657 ( .A(REG0_REG_6__SCAN_IN), .ZN(n5169) );
  OR2_X1 U3658 ( .A1(n2513), .A2(n5169), .ZN(n3149) );
  NAND4_X1 U3659 ( .A1(n3152), .A2(n3151), .A3(n3150), .A4(n3149), .ZN(n5181)
         );
  INV_X1 U3660 ( .A(n5181), .ZN(n3390) );
  INV_X1 U3661 ( .A(n5163), .ZN(n3153) );
  MUX2_X1 U3662 ( .A(n3153), .B(DATAI_6_), .S(n4064), .Z(n3386) );
  OAI22_X1 U3663 ( .A1(n3390), .A2(n3800), .B1(n2511), .B2(n3389), .ZN(n3297)
         );
  NAND2_X1 U3664 ( .A1(n5181), .A2(n3293), .ZN(n3155) );
  NAND2_X1 U3665 ( .A1(n3386), .A2(n3815), .ZN(n3154) );
  NAND2_X1 U3666 ( .A1(n3155), .A2(n3154), .ZN(n3156) );
  XNOR2_X1 U3667 ( .A(n3156), .B(n3829), .ZN(n3296) );
  XOR2_X1 U3668 ( .A(n3297), .B(n3296), .Z(n3169) );
  MUX2_X1 U3669 ( .A(n4979), .B(DATAI_5_), .S(n4064), .Z(n3270) );
  INV_X1 U3670 ( .A(n3270), .ZN(n3280) );
  OAI22_X1 U3671 ( .A1(n3281), .A2(n3798), .B1(n3108), .B2(n3280), .ZN(n3157)
         );
  OR2_X1 U3672 ( .A1(n3281), .A2(n3800), .ZN(n3159) );
  NAND2_X1 U3673 ( .A1(n3270), .A2(n3293), .ZN(n3158) );
  NAND2_X1 U3674 ( .A1(n3159), .A2(n3158), .ZN(n3160) );
  INV_X1 U3675 ( .A(n3163), .ZN(n3165) );
  NAND2_X1 U3676 ( .A1(n3165), .A2(n3164), .ZN(n3263) );
  OAI21_X1 U3677 ( .B1(n3169), .B2(n3168), .A(n3301), .ZN(n3181) );
  AOI22_X1 U3678 ( .A1(n3386), .A2(n3972), .B1(n3980), .B2(n4162), .ZN(n3179)
         );
  NAND2_X1 U3679 ( .A1(n4052), .A2(REG2_REG_7__SCAN_IN), .ZN(n3176) );
  INV_X1 U3680 ( .A(REG1_REG_7__SCAN_IN), .ZN(n3170) );
  OR2_X1 U3681 ( .A1(n4061), .A2(n3170), .ZN(n3175) );
  NOR2_X1 U3682 ( .A1(n3171), .A2(REG3_REG_7__SCAN_IN), .ZN(n3172) );
  OR2_X1 U3683 ( .A1(n3333), .A2(n3172), .ZN(n5189) );
  OR2_X1 U3684 ( .A1(n3835), .A2(n5189), .ZN(n3174) );
  INV_X1 U3685 ( .A(REG0_REG_7__SCAN_IN), .ZN(n5199) );
  OR2_X1 U3686 ( .A1(n2513), .A2(n5199), .ZN(n3173) );
  AOI21_X1 U3687 ( .B1(n5309), .B2(n4161), .A(n3177), .ZN(n3178) );
  OAI211_X1 U3688 ( .C1(n5354), .C2(n3286), .A(n3179), .B(n3178), .ZN(n3180)
         );
  AOI21_X1 U3689 ( .B1(n3181), .B2(n5314), .A(n3180), .ZN(n3182) );
  INV_X1 U3690 ( .A(n3182), .ZN(U3236) );
  NAND2_X1 U3691 ( .A1(n3183), .A2(n3222), .ZN(n3989) );
  NAND2_X1 U3692 ( .A1(n3989), .A2(n3990), .ZN(n3200) );
  NAND2_X1 U3693 ( .A1(n3186), .A2(n3227), .ZN(n4109) );
  NAND2_X1 U3694 ( .A1(n3221), .A2(n3990), .ZN(n3249) );
  NAND2_X1 U3695 ( .A1(n4164), .A2(n3204), .ZN(n3994) );
  NAND2_X1 U3696 ( .A1(n5133), .A2(n3971), .ZN(n3991) );
  NAND2_X1 U3697 ( .A1(n3994), .A2(n3991), .ZN(n3202) );
  NAND2_X1 U3698 ( .A1(n3249), .A2(n4083), .ZN(n3187) );
  NAND2_X1 U3699 ( .A1(n3187), .A2(n3991), .ZN(n5130) );
  NAND2_X1 U3700 ( .A1(n3251), .A2(n3350), .ZN(n3996) );
  NAND2_X1 U3701 ( .A1(n4163), .A2(n5132), .ZN(n3993) );
  NAND2_X1 U3702 ( .A1(n5130), .A2(n5131), .ZN(n3188) );
  NAND2_X1 U3703 ( .A1(n3188), .A2(n3996), .ZN(n3233) );
  NAND2_X1 U3704 ( .A1(n3189), .A2(n3240), .ZN(n3997) );
  NAND2_X1 U3705 ( .A1(n3997), .A2(n3999), .ZN(n4079) );
  XNOR2_X1 U3706 ( .A(n3233), .B(n4079), .ZN(n3194) );
  OR2_X1 U3707 ( .A1(n3023), .A2(n4114), .ZN(n4140) );
  OR2_X1 U3708 ( .A1(n4138), .A2(n3208), .ZN(n3190) );
  OAI22_X1 U3709 ( .A1(n3251), .A2(n5246), .B1(n5266), .B2(n3191), .ZN(n3192)
         );
  AOI21_X1 U3710 ( .B1(n5136), .B2(n4162), .A(n3192), .ZN(n3193) );
  OAI21_X1 U3711 ( .B1(n3194), .B2(n5138), .A(n3193), .ZN(n5155) );
  INV_X1 U3712 ( .A(n5155), .ZN(n3215) );
  NAND3_X1 U3713 ( .A1(n3195), .A2(n4463), .A3(n4465), .ZN(n3196) );
  NAND2_X1 U3714 ( .A1(n5105), .A2(n3222), .ZN(n3256) );
  NOR2_X1 U3715 ( .A1(n3256), .A2(n3971), .ZN(n5129) );
  AND2_X1 U3716 ( .A1(n3197), .A2(n3237), .ZN(n5156) );
  INV_X2 U3717 ( .A(n5226), .ZN(n5374) );
  OAI22_X1 U3718 ( .A1(n5226), .A2(n5094), .B1(n3198), .B2(n5231), .ZN(n3199)
         );
  AOI21_X1 U3719 ( .B1(n5156), .B2(n4247), .A(n3199), .ZN(n3214) );
  NAND2_X1 U3720 ( .A1(n3200), .A2(n3217), .ZN(n3216) );
  NAND2_X1 U3721 ( .A1(n5103), .A2(n3184), .ZN(n3201) );
  NAND2_X1 U3722 ( .A1(n3216), .A2(n3201), .ZN(n3247) );
  INV_X1 U3723 ( .A(n3247), .ZN(n3203) );
  NAND2_X1 U3724 ( .A1(n3203), .A2(n3202), .ZN(n3246) );
  NAND2_X1 U3725 ( .A1(n5133), .A2(n3204), .ZN(n3205) );
  NAND2_X1 U3726 ( .A1(n3246), .A2(n3205), .ZN(n5128) );
  NOR2_X1 U3727 ( .A1(n4163), .A2(n3350), .ZN(n3207) );
  NAND2_X1 U3728 ( .A1(n4163), .A2(n3350), .ZN(n3206) );
  XOR2_X1 U3729 ( .A(n3242), .B(n4079), .Z(n5157) );
  NAND2_X1 U3730 ( .A1(n3209), .A2(n3208), .ZN(n3212) );
  AND2_X1 U3731 ( .A1(n3210), .A2(n4138), .ZN(n3211) );
  NAND2_X1 U3732 ( .A1(n3212), .A2(n3211), .ZN(n5102) );
  OR2_X1 U3733 ( .A1(n5112), .A2(n4114), .ZN(n3219) );
  NAND2_X1 U3734 ( .A1(n5102), .A2(n3219), .ZN(n5177) );
  NAND2_X1 U3735 ( .A1(n5157), .A2(n4437), .ZN(n3213) );
  OAI211_X1 U3736 ( .C1(n3215), .C2(n5374), .A(n3214), .B(n3213), .ZN(U3286)
         );
  NAND2_X1 U3737 ( .A1(n3216), .A2(n3218), .ZN(n5117) );
  INV_X1 U3738 ( .A(n3219), .ZN(n3220) );
  AND2_X1 U3739 ( .A1(n5226), .A2(n3220), .ZN(n5279) );
  INV_X1 U3740 ( .A(n5279), .ZN(n3261) );
  OAI21_X1 U3741 ( .B1(n4084), .B2(n2560), .A(n3221), .ZN(n3225) );
  NOR2_X1 U3742 ( .A1(n3222), .A2(n5266), .ZN(n3224) );
  AOI211_X1 U3743 ( .C1(n3225), .C2(n5268), .A(n3224), .B(n3223), .ZN(n3226)
         );
  OAI21_X1 U3744 ( .B1(n5102), .B2(n5117), .A(n3226), .ZN(n5118) );
  NAND2_X1 U3745 ( .A1(n5118), .A2(n4450), .ZN(n3232) );
  NAND2_X1 U3746 ( .A1(n3227), .A2(n3184), .ZN(n3228) );
  AND3_X1 U3747 ( .A1(n3256), .A2(n5377), .A3(n3228), .ZN(n5119) );
  OAI22_X1 U3748 ( .A1(n4450), .A2(n2890), .B1(n3229), .B2(n5231), .ZN(n3230)
         );
  AOI21_X1 U3749 ( .B1(n4247), .B2(n5119), .A(n3230), .ZN(n3231) );
  OAI211_X1 U3750 ( .C1(n5117), .C2(n3261), .A(n3232), .B(n3231), .ZN(U3289)
         );
  NAND2_X1 U3751 ( .A1(n3281), .A2(n3270), .ZN(n4004) );
  NAND2_X1 U3752 ( .A1(n4162), .A2(n3280), .ZN(n4000) );
  NAND2_X1 U3753 ( .A1(n4004), .A2(n4000), .ZN(n4080) );
  NAND2_X1 U3754 ( .A1(n3233), .A2(n3999), .ZN(n3234) );
  XOR2_X1 U3755 ( .A(n4080), .B(n3274), .Z(n3236) );
  AOI22_X1 U3756 ( .A1(n5135), .A2(n5180), .B1(n5136), .B2(n5181), .ZN(n3268)
         );
  OAI21_X1 U3757 ( .B1(n5266), .B2(n3280), .A(n3268), .ZN(n3235) );
  AOI21_X1 U3758 ( .B1(n3236), .B2(n5268), .A(n3235), .ZN(n4520) );
  AOI21_X1 U3759 ( .B1(n3270), .B2(n3237), .A(n3285), .ZN(n4518) );
  INV_X1 U3760 ( .A(REG2_REG_5__SCAN_IN), .ZN(n3238) );
  OAI22_X1 U3761 ( .A1(n4450), .A2(n3238), .B1(n3273), .B2(n5231), .ZN(n3239)
         );
  AOI21_X1 U3762 ( .B1(n4518), .B2(n5372), .A(n3239), .ZN(n3245) );
  AND2_X1 U3763 ( .A1(n5135), .A2(n3240), .ZN(n3241) );
  AOI21_X1 U3764 ( .B1(n3242), .B2(n4079), .A(n3241), .ZN(n3243) );
  NAND2_X1 U3765 ( .A1(n3243), .A2(n4080), .ZN(n3283) );
  OAI21_X1 U3766 ( .B1(n3243), .B2(n4080), .A(n3283), .ZN(n4519) );
  NAND2_X1 U3767 ( .A1(n4519), .A2(n4437), .ZN(n3244) );
  OAI211_X1 U3768 ( .C1(n4520), .C2(n5374), .A(n3245), .B(n3244), .ZN(U3285)
         );
  NAND2_X1 U3769 ( .A1(n3247), .A2(n4083), .ZN(n3248) );
  NAND2_X1 U3770 ( .A1(n3246), .A2(n3248), .ZN(n3253) );
  INV_X1 U3771 ( .A(n3253), .ZN(n5123) );
  XOR2_X1 U3772 ( .A(n4083), .B(n3249), .Z(n3255) );
  INV_X1 U3773 ( .A(n5102), .ZN(n5274) );
  AOI22_X1 U3774 ( .A1(n5103), .A2(n5180), .B1(n5365), .B2(n3971), .ZN(n3250)
         );
  OAI21_X1 U3775 ( .B1(n3251), .B2(n5244), .A(n3250), .ZN(n3252) );
  AOI21_X1 U3776 ( .B1(n3253), .B2(n5274), .A(n3252), .ZN(n3254) );
  OAI21_X1 U3777 ( .B1(n3255), .B2(n5138), .A(n3254), .ZN(n5124) );
  NAND2_X1 U3778 ( .A1(n5124), .A2(n5226), .ZN(n3260) );
  AOI21_X1 U3779 ( .B1(n3971), .B2(n3256), .A(n5129), .ZN(n5126) );
  OAI22_X1 U3780 ( .A1(n4450), .A2(n2892), .B1(n3257), .B2(n5231), .ZN(n3258)
         );
  AOI21_X1 U3781 ( .B1(n5126), .B2(n5372), .A(n3258), .ZN(n3259) );
  OAI211_X1 U3782 ( .C1(n5123), .C2(n3261), .A(n3260), .B(n3259), .ZN(U3288)
         );
  INV_X1 U3783 ( .A(n3262), .ZN(n3266) );
  AOI21_X1 U3784 ( .B1(n3264), .B2(n3263), .A(n2750), .ZN(n3265) );
  OAI21_X1 U3785 ( .B1(n3266), .B2(n3265), .A(n5314), .ZN(n3272) );
  INV_X1 U3786 ( .A(REG3_REG_5__SCAN_IN), .ZN(n3267) );
  NOR2_X1 U3787 ( .A1(STATE_REG_SCAN_IN), .A2(n3267), .ZN(n4974) );
  NOR2_X1 U3788 ( .A1(n3268), .A2(n3375), .ZN(n3269) );
  AOI211_X1 U3789 ( .C1(n3270), .C2(n5339), .A(n4974), .B(n3269), .ZN(n3271)
         );
  OAI211_X1 U3790 ( .C1(n5354), .C2(n3273), .A(n3272), .B(n3271), .ZN(U3224)
         );
  NAND2_X1 U3791 ( .A1(n3390), .A2(n3386), .ZN(n4006) );
  NAND2_X1 U3792 ( .A1(n5181), .A2(n3389), .ZN(n4002) );
  INV_X1 U3793 ( .A(n4082), .ZN(n3275) );
  XNOR2_X1 U3794 ( .A(n3380), .B(n3275), .ZN(n3276) );
  NAND2_X1 U3795 ( .A1(n3276), .A2(n5268), .ZN(n3279) );
  OAI22_X1 U3796 ( .A1(n3281), .A2(n5246), .B1(n5266), .B2(n3389), .ZN(n3277)
         );
  INV_X1 U3797 ( .A(n3277), .ZN(n3278) );
  OAI211_X1 U3798 ( .C1(n3382), .C2(n5244), .A(n3279), .B(n3278), .ZN(n5165)
         );
  INV_X1 U3799 ( .A(n5165), .ZN(n3291) );
  NAND2_X1 U3800 ( .A1(n3281), .A2(n3280), .ZN(n3282) );
  NAND2_X1 U3801 ( .A1(n3283), .A2(n3282), .ZN(n3388) );
  XOR2_X1 U3802 ( .A(n3388), .B(n4082), .Z(n5167) );
  INV_X1 U3803 ( .A(n5188), .ZN(n3284) );
  OAI21_X1 U3804 ( .B1(n3285), .B2(n3389), .A(n3284), .ZN(n5164) );
  INV_X1 U3805 ( .A(n5372), .ZN(n4454) );
  NOR2_X1 U3806 ( .A1(n5164), .A2(n4454), .ZN(n3289) );
  OAI22_X1 U3807 ( .A1(n4450), .A2(n3287), .B1(n3286), .B2(n5231), .ZN(n3288)
         );
  AOI211_X1 U3808 ( .C1(n5167), .C2(n4437), .A(n3289), .B(n3288), .ZN(n3290)
         );
  OAI21_X1 U3809 ( .B1(n5374), .B2(n3291), .A(n3290), .ZN(U3284) );
  MUX2_X1 U3810 ( .A(n5171), .B(DATAI_7_), .S(n4064), .Z(n5179) );
  OAI22_X1 U3811 ( .A1(n3382), .A2(n3798), .B1(n3108), .B2(n5187), .ZN(n3292)
         );
  XNOR2_X1 U3812 ( .A(n3292), .B(n3782), .ZN(n3321) );
  OR2_X1 U3813 ( .A1(n3382), .A2(n3800), .ZN(n3295) );
  NAND2_X1 U3814 ( .A1(n5179), .A2(n3293), .ZN(n3294) );
  NAND2_X1 U3815 ( .A1(n3295), .A2(n3294), .ZN(n3322) );
  XNOR2_X1 U3816 ( .A(n3321), .B(n3322), .ZN(n3302) );
  INV_X1 U3817 ( .A(n3296), .ZN(n3299) );
  INV_X1 U3818 ( .A(n3297), .ZN(n3298) );
  NAND2_X1 U3819 ( .A1(n3299), .A2(n3298), .ZN(n3303) );
  INV_X1 U3820 ( .A(n3325), .ZN(n3305) );
  AOI21_X1 U3821 ( .B1(n3301), .B2(n3303), .A(n3302), .ZN(n3304) );
  NOR3_X1 U3822 ( .A1(n3305), .A2(n3304), .A3(n5344), .ZN(n3314) );
  AOI22_X1 U3823 ( .A1(n5179), .A2(n5339), .B1(n3980), .B2(n5181), .ZN(n3312)
         );
  NAND2_X1 U3824 ( .A1(n4052), .A2(REG2_REG_8__SCAN_IN), .ZN(n3309) );
  OR2_X1 U3825 ( .A1(n4061), .A2(n5205), .ZN(n3308) );
  XNOR2_X1 U3826 ( .A(n3333), .B(REG3_REG_8__SCAN_IN), .ZN(n3397) );
  OR2_X1 U3827 ( .A1(n3835), .A2(n3397), .ZN(n3307) );
  INV_X1 U3828 ( .A(REG0_REG_8__SCAN_IN), .ZN(n4709) );
  OR2_X1 U3829 ( .A1(n2513), .A2(n4709), .ZN(n3306) );
  INV_X1 U3830 ( .A(REG3_REG_7__SCAN_IN), .ZN(n3310) );
  NOR2_X1 U3831 ( .A1(STATE_REG_SCAN_IN), .A2(n3310), .ZN(n4984) );
  AOI21_X1 U3832 ( .B1(n5309), .B2(n4160), .A(n4984), .ZN(n3311) );
  OAI211_X1 U3833 ( .C1(n5354), .C2(n5189), .A(n3312), .B(n3311), .ZN(n3313)
         );
  OR2_X1 U3834 ( .A1(n3314), .A2(n3313), .ZN(U3210) );
  INV_X1 U3835 ( .A(DATAI_8_), .ZN(n4739) );
  MUX2_X1 U3836 ( .A(n3315), .B(n4739), .S(n4064), .Z(n4014) );
  OAI22_X1 U3837 ( .A1(n5183), .A2(n3798), .B1(n3108), .B2(n4014), .ZN(n3316)
         );
  XNOR2_X1 U3838 ( .A(n3316), .B(n3829), .ZN(n3320) );
  OR2_X1 U3839 ( .A1(n5183), .A2(n3800), .ZN(n3318) );
  NAND2_X1 U3840 ( .A1(n3472), .A2(n3293), .ZN(n3317) );
  NAND2_X1 U3841 ( .A1(n3318), .A2(n3317), .ZN(n3319) );
  NOR2_X1 U3842 ( .A1(n3320), .A2(n3319), .ZN(n3360) );
  AOI21_X1 U3843 ( .B1(n3320), .B2(n3319), .A(n3360), .ZN(n3326) );
  INV_X1 U3844 ( .A(n3321), .ZN(n3323) );
  NAND2_X1 U3845 ( .A1(n3323), .A2(n3322), .ZN(n3327) );
  INV_X1 U3846 ( .A(n3362), .ZN(n3329) );
  AOI21_X1 U3847 ( .B1(n3325), .B2(n3327), .A(n3326), .ZN(n3328) );
  OAI21_X1 U3848 ( .B1(n3329), .B2(n3328), .A(n5314), .ZN(n3344) );
  OR2_X1 U3849 ( .A1(n3382), .A2(n5246), .ZN(n3340) );
  NAND2_X1 U3850 ( .A1(n4052), .A2(REG2_REG_9__SCAN_IN), .ZN(n3338) );
  INV_X1 U3851 ( .A(REG1_REG_9__SCAN_IN), .ZN(n3330) );
  OR2_X1 U3852 ( .A1(n4061), .A2(n3330), .ZN(n3337) );
  INV_X1 U3853 ( .A(REG0_REG_9__SCAN_IN), .ZN(n3331) );
  OR2_X1 U3854 ( .A1(n2513), .A2(n3331), .ZN(n3336) );
  AOI21_X1 U3855 ( .B1(n3333), .B2(REG3_REG_8__SCAN_IN), .A(
        REG3_REG_9__SCAN_IN), .ZN(n3334) );
  OR2_X1 U3856 ( .A1(n3366), .A2(n3334), .ZN(n5230) );
  OR2_X1 U3857 ( .A1(n3835), .A2(n5230), .ZN(n3335) );
  NAND4_X1 U3858 ( .A1(n3338), .A2(n3337), .A3(n3336), .A4(n3335), .ZN(n4159)
         );
  NAND2_X1 U3859 ( .A1(n4159), .A2(n5136), .ZN(n3339) );
  NAND2_X1 U3860 ( .A1(n3340), .A2(n3339), .ZN(n3383) );
  INV_X1 U3861 ( .A(n3383), .ZN(n3341) );
  NAND2_X1 U3862 ( .A1(REG3_REG_8__SCAN_IN), .A2(U3149), .ZN(n5000) );
  OAI21_X1 U3863 ( .B1(n3341), .B2(n3375), .A(n5000), .ZN(n3342) );
  AOI21_X1 U3864 ( .B1(n3472), .B2(n5339), .A(n3342), .ZN(n3343) );
  OAI211_X1 U3865 ( .C1(n5354), .C2(n3397), .A(n3344), .B(n3343), .ZN(U3218)
         );
  NAND2_X1 U3866 ( .A1(n3967), .A2(n3968), .ZN(n3966) );
  INV_X1 U3867 ( .A(n3345), .ZN(n3346) );
  NAND2_X1 U3868 ( .A1(n3966), .A2(n3346), .ZN(n3348) );
  OAI21_X1 U3869 ( .B1(n3349), .B2(n3348), .A(n3347), .ZN(n3355) );
  AOI22_X1 U3870 ( .A1(n3350), .A2(n5339), .B1(n3980), .B2(n4164), .ZN(n3353)
         );
  AOI21_X1 U3871 ( .B1(n5309), .B2(n5135), .A(n3351), .ZN(n3352) );
  OAI211_X1 U3872 ( .C1(REG3_REG_3__SCAN_IN), .C2(n5354), .A(n3353), .B(n3352), 
        .ZN(n3354) );
  AOI21_X1 U3873 ( .B1(n3355), .B2(n5314), .A(n3354), .ZN(n3356) );
  INV_X1 U3874 ( .A(n3356), .ZN(U3215) );
  INV_X1 U3875 ( .A(n4159), .ZN(n3463) );
  MUX2_X1 U3876 ( .A(n5010), .B(DATAI_9_), .S(n4064), .Z(n5208) );
  INV_X1 U3877 ( .A(n5208), .ZN(n5215) );
  OAI22_X1 U3878 ( .A1(n3463), .A2(n3800), .B1(n3798), .B2(n5215), .ZN(n3406)
         );
  NAND2_X1 U3879 ( .A1(n4159), .A2(n3293), .ZN(n3358) );
  NAND2_X1 U3880 ( .A1(n5208), .A2(n3815), .ZN(n3357) );
  NAND2_X1 U3881 ( .A1(n3358), .A2(n3357), .ZN(n3359) );
  XNOR2_X1 U3882 ( .A(n3359), .B(n3829), .ZN(n3405) );
  XOR2_X1 U3883 ( .A(n3406), .B(n3405), .Z(n3364) );
  INV_X1 U3884 ( .A(n3360), .ZN(n3361) );
  NAND2_X1 U3885 ( .A1(n3362), .A2(n3361), .ZN(n3363) );
  NAND2_X1 U3886 ( .A1(n3363), .A2(n3364), .ZN(n3412) );
  OAI21_X1 U3887 ( .B1(n3364), .B2(n3363), .A(n3412), .ZN(n3378) );
  NOR2_X1 U3888 ( .A1(n5354), .A2(n5230), .ZN(n3377) );
  NAND2_X1 U3889 ( .A1(n4052), .A2(REG2_REG_10__SCAN_IN), .ZN(n3371) );
  INV_X1 U3890 ( .A(REG0_REG_10__SCAN_IN), .ZN(n3365) );
  OR2_X1 U3891 ( .A1(n2513), .A2(n3365), .ZN(n3370) );
  OR2_X1 U3892 ( .A1(n3366), .A2(REG3_REG_10__SCAN_IN), .ZN(n3367) );
  NAND2_X1 U3893 ( .A1(n3436), .A2(n3367), .ZN(n3471) );
  OR2_X1 U3894 ( .A1(n3835), .A2(n3471), .ZN(n3369) );
  OR2_X1 U3895 ( .A1(n4061), .A2(n5237), .ZN(n3368) );
  OR2_X1 U3896 ( .A1(n5247), .A2(n5244), .ZN(n3373) );
  OR2_X1 U3897 ( .A1(n5183), .A2(n5246), .ZN(n3372) );
  AND2_X1 U3898 ( .A1(n3373), .A2(n3372), .ZN(n5214) );
  NAND2_X1 U3899 ( .A1(REG3_REG_9__SCAN_IN), .A2(U3149), .ZN(n5011) );
  NAND2_X1 U3900 ( .A1(n3972), .A2(n5208), .ZN(n3374) );
  OAI211_X1 U3901 ( .C1(n5214), .C2(n3375), .A(n5011), .B(n3374), .ZN(n3376)
         );
  AOI211_X1 U3902 ( .C1(n3378), .C2(n5314), .A(n3377), .B(n3376), .ZN(n3379)
         );
  INV_X1 U3903 ( .A(n3379), .ZN(U3228) );
  XNOR2_X1 U3904 ( .A(n4160), .B(n3472), .ZN(n4104) );
  NAND2_X1 U3905 ( .A1(n3381), .A2(n4002), .ZN(n5178) );
  NAND2_X1 U3906 ( .A1(n3382), .A2(n5179), .ZN(n4007) );
  NAND2_X1 U3907 ( .A1(n4161), .A2(n5187), .ZN(n4009) );
  XOR2_X1 U3908 ( .A(n4104), .B(n3462), .Z(n3385) );
  NOR2_X1 U3909 ( .A1(n4014), .A2(n5266), .ZN(n3384) );
  AOI211_X1 U3910 ( .C1(n3385), .C2(n5268), .A(n3384), .B(n3383), .ZN(n5201)
         );
  NAND2_X1 U3911 ( .A1(n5181), .A2(n3386), .ZN(n3387) );
  NAND2_X1 U3912 ( .A1(n3388), .A2(n3387), .ZN(n3392) );
  NAND2_X1 U3913 ( .A1(n3390), .A2(n3389), .ZN(n3391) );
  NAND2_X1 U3914 ( .A1(n3392), .A2(n3391), .ZN(n5173) );
  INV_X1 U3915 ( .A(n5173), .ZN(n3394) );
  NAND2_X1 U3916 ( .A1(n4161), .A2(n5179), .ZN(n3395) );
  XNOR2_X1 U3917 ( .A(n3473), .B(n4104), .ZN(n5204) );
  INV_X1 U3918 ( .A(n5186), .ZN(n3396) );
  OAI21_X1 U3919 ( .B1(n3396), .B2(n4014), .A(n5209), .ZN(n5202) );
  NOR2_X1 U3920 ( .A1(n5202), .A2(n4454), .ZN(n3399) );
  OAI22_X1 U3921 ( .A1(n4450), .A2(n4995), .B1(n3397), .B2(n5231), .ZN(n3398)
         );
  AOI211_X1 U3922 ( .C1(n5204), .C2(n4437), .A(n3399), .B(n3398), .ZN(n3400)
         );
  OAI21_X1 U3923 ( .B1(n5201), .B2(n5374), .A(n3400), .ZN(U3282) );
  INV_X1 U3924 ( .A(n3483), .ZN(n3401) );
  MUX2_X1 U3925 ( .A(n3401), .B(DATAI_10_), .S(n4064), .Z(n3470) );
  INV_X1 U3926 ( .A(n3470), .ZN(n3496) );
  OAI22_X1 U3927 ( .A1(n5247), .A2(n3798), .B1(n3108), .B2(n3496), .ZN(n3402)
         );
  XNOR2_X1 U3928 ( .A(n3402), .B(n3782), .ZN(n3425) );
  OR2_X1 U3929 ( .A1(n5247), .A2(n3110), .ZN(n3404) );
  NAND2_X1 U3930 ( .A1(n3470), .A2(n3740), .ZN(n3403) );
  NAND2_X1 U3931 ( .A1(n3404), .A2(n3403), .ZN(n3428) );
  XNOR2_X1 U3932 ( .A(n3425), .B(n3428), .ZN(n3410) );
  INV_X1 U3933 ( .A(n3405), .ZN(n3408) );
  INV_X1 U3934 ( .A(n3406), .ZN(n3407) );
  NAND2_X1 U3935 ( .A1(n3408), .A2(n3407), .ZN(n3411) );
  AND2_X2 U3936 ( .A1(n3412), .A2(n3409), .ZN(n3426) );
  AOI21_X1 U3937 ( .B1(n3412), .B2(n3411), .A(n3410), .ZN(n3413) );
  NOR3_X1 U3938 ( .A1(n3426), .A2(n3413), .A3(n5344), .ZN(n3424) );
  AOI22_X1 U3939 ( .A1(n3470), .A2(n5339), .B1(n3980), .B2(n4159), .ZN(n3422)
         );
  NAND2_X1 U3940 ( .A1(n4052), .A2(REG2_REG_11__SCAN_IN), .ZN(n3419) );
  INV_X1 U3941 ( .A(REG0_REG_11__SCAN_IN), .ZN(n3414) );
  OR2_X1 U3942 ( .A1(n2513), .A2(n3414), .ZN(n3418) );
  INV_X1 U3943 ( .A(REG1_REG_11__SCAN_IN), .ZN(n3415) );
  OR2_X1 U3944 ( .A1(n4061), .A2(n3415), .ZN(n3417) );
  INV_X1 U3945 ( .A(REG3_REG_11__SCAN_IN), .ZN(n3435) );
  XNOR2_X1 U3946 ( .A(n3436), .B(n3435), .ZN(n5275) );
  OR2_X1 U3947 ( .A1(n3835), .A2(n5275), .ZN(n3416) );
  INV_X1 U3948 ( .A(REG3_REG_10__SCAN_IN), .ZN(n3420) );
  NOR2_X1 U3949 ( .A1(STATE_REG_SCAN_IN), .A2(n3420), .ZN(n3481) );
  AOI21_X1 U3950 ( .B1(n5309), .B2(n4157), .A(n3481), .ZN(n3421) );
  OAI211_X1 U3951 ( .C1(n5354), .C2(n3471), .A(n3422), .B(n3421), .ZN(n3423)
         );
  OR2_X1 U3952 ( .A1(n3424), .A2(n3423), .ZN(U3214) );
  INV_X1 U3953 ( .A(n3425), .ZN(n3427) );
  MUX2_X1 U3954 ( .A(n5021), .B(DATAI_11_), .S(n4064), .Z(n5260) );
  OAI22_X1 U3955 ( .A1(n3499), .A2(n3798), .B1(n3108), .B2(n5265), .ZN(n3429)
         );
  XNOR2_X1 U3956 ( .A(n3429), .B(n3829), .ZN(n3433) );
  OR2_X1 U3957 ( .A1(n3499), .A2(n3800), .ZN(n3431) );
  NAND2_X1 U3958 ( .A1(n5260), .A2(n3293), .ZN(n3430) );
  NAND2_X1 U3959 ( .A1(n3431), .A2(n3430), .ZN(n3432) );
  NAND2_X1 U3960 ( .A1(n3433), .A2(n3432), .ZN(n5239) );
  NOR2_X1 U3961 ( .A1(n3433), .A2(n3432), .ZN(n5241) );
  NAND2_X1 U3962 ( .A1(n4052), .A2(REG2_REG_12__SCAN_IN), .ZN(n3443) );
  INV_X1 U3963 ( .A(REG0_REG_12__SCAN_IN), .ZN(n3434) );
  OR2_X1 U3964 ( .A1(n2513), .A2(n3434), .ZN(n3442) );
  INV_X1 U3965 ( .A(REG3_REG_12__SCAN_IN), .ZN(n4776) );
  OAI21_X1 U3966 ( .B1(n3436), .B2(n3435), .A(n4776), .ZN(n3439) );
  INV_X1 U3967 ( .A(n3449), .ZN(n3450) );
  NAND2_X1 U3968 ( .A1(n3439), .A2(n3450), .ZN(n3502) );
  OR2_X1 U3969 ( .A1(n3835), .A2(n3502), .ZN(n3441) );
  OR2_X1 U3970 ( .A1(n4061), .A2(n5288), .ZN(n3440) );
  MUX2_X1 U3971 ( .A(n2818), .B(DATAI_12_), .S(n4064), .Z(n3540) );
  INV_X1 U3972 ( .A(n3540), .ZN(n3501) );
  OAI22_X1 U3973 ( .A1(n5245), .A2(n3798), .B1(n3108), .B2(n3501), .ZN(n3444)
         );
  XNOR2_X1 U3974 ( .A(n3444), .B(n3782), .ZN(n3514) );
  OR2_X1 U3975 ( .A1(n5245), .A2(n3800), .ZN(n3446) );
  NAND2_X1 U3976 ( .A1(n3540), .A2(n3293), .ZN(n3445) );
  XNOR2_X1 U3977 ( .A(n3514), .B(n3515), .ZN(n3447) );
  XNOR2_X1 U3978 ( .A(n2548), .B(n3447), .ZN(n3460) );
  AOI22_X1 U3979 ( .A1(n3540), .A2(n5339), .B1(n3980), .B2(n4157), .ZN(n3458)
         );
  NAND2_X1 U3980 ( .A1(n4052), .A2(REG2_REG_13__SCAN_IN), .ZN(n3456) );
  INV_X1 U3981 ( .A(REG1_REG_13__SCAN_IN), .ZN(n3448) );
  OR2_X1 U3982 ( .A1(n4061), .A2(n3448), .ZN(n3455) );
  INV_X1 U3983 ( .A(REG3_REG_13__SCAN_IN), .ZN(n3529) );
  NAND2_X1 U3984 ( .A1(n3450), .A2(n3529), .ZN(n3451) );
  NAND2_X1 U3985 ( .A1(n3522), .A2(n3451), .ZN(n3544) );
  OR2_X1 U3986 ( .A1(n3835), .A2(n3544), .ZN(n3454) );
  INV_X1 U3987 ( .A(REG0_REG_13__SCAN_IN), .ZN(n3452) );
  OR2_X1 U3988 ( .A1(n2513), .A2(n3452), .ZN(n3453) );
  NAND4_X1 U3989 ( .A1(n3456), .A2(n3455), .A3(n3454), .A4(n3453), .ZN(n4155)
         );
  NOR2_X1 U3990 ( .A1(STATE_REG_SCAN_IN), .A2(n4776), .ZN(n3624) );
  AOI21_X1 U3991 ( .B1(n5309), .B2(n4155), .A(n3624), .ZN(n3457) );
  OAI211_X1 U3992 ( .C1(n5354), .C2(n3502), .A(n3458), .B(n3457), .ZN(n3459)
         );
  AOI21_X1 U3993 ( .B1(n3460), .B2(n5314), .A(n3459), .ZN(n3461) );
  INV_X1 U3994 ( .A(n3461), .ZN(U3221) );
  NAND2_X1 U3995 ( .A1(n4160), .A2(n4014), .ZN(n4008) );
  NAND2_X1 U3996 ( .A1(n3463), .A2(n5208), .ZN(n4012) );
  AND2_X1 U3997 ( .A1(n4159), .A2(n5215), .ZN(n4016) );
  AOI21_X1 U3998 ( .B1(n5213), .B2(n4012), .A(n4016), .ZN(n3492) );
  NAND2_X1 U3999 ( .A1(n5247), .A2(n3470), .ZN(n3491) );
  INV_X1 U4000 ( .A(n5247), .ZN(n4158) );
  NAND2_X1 U4001 ( .A1(n4158), .A2(n3496), .ZN(n4015) );
  NAND2_X1 U4002 ( .A1(n3491), .A2(n4015), .ZN(n4081) );
  INV_X1 U4003 ( .A(n4081), .ZN(n3464) );
  XNOR2_X1 U4004 ( .A(n3492), .B(n3464), .ZN(n3465) );
  NAND2_X1 U4005 ( .A1(n3465), .A2(n5268), .ZN(n3469) );
  AOI22_X1 U4006 ( .A1(n4159), .A2(n5180), .B1(n5365), .B2(n3470), .ZN(n3466)
         );
  OAI21_X1 U4007 ( .B1(n3499), .B2(n5244), .A(n3466), .ZN(n3467) );
  INV_X1 U4008 ( .A(n3467), .ZN(n3468) );
  NAND2_X1 U4009 ( .A1(n3469), .A2(n3468), .ZN(n5235) );
  INV_X1 U4010 ( .A(n5235), .ZN(n3478) );
  AOI21_X1 U4011 ( .B1(n3470), .B2(n5211), .A(n5257), .ZN(n5236) );
  OAI22_X1 U4012 ( .A1(n4450), .A2(n3486), .B1(n3471), .B2(n5231), .ZN(n3476)
         );
  NOR2_X1 U4013 ( .A1(n4159), .A2(n5208), .ZN(n4093) );
  NOR2_X1 U4014 ( .A1(n3474), .A2(n4081), .ZN(n5233) );
  NAND2_X1 U4015 ( .A1(n3474), .A2(n4081), .ZN(n3498) );
  INV_X1 U4016 ( .A(n3498), .ZN(n5232) );
  NOR3_X1 U4017 ( .A1(n5233), .A2(n5232), .A3(n4399), .ZN(n3475) );
  AOI211_X1 U4018 ( .C1(n5372), .C2(n5236), .A(n3476), .B(n3475), .ZN(n3477)
         );
  OAI21_X1 U4019 ( .B1(n5374), .B2(n3478), .A(n3477), .ZN(U3280) );
  AOI21_X1 U4020 ( .B1(n5237), .B2(n3479), .A(n3480), .ZN(n3489) );
  AOI21_X1 U4021 ( .B1(n5087), .B2(ADDR_REG_10__SCAN_IN), .A(n3481), .ZN(n3482) );
  OAI21_X1 U4022 ( .B1(n3483), .B2(n5069), .A(n3482), .ZN(n3488) );
  AOI211_X1 U4023 ( .C1(n3486), .C2(n3485), .A(n3484), .B(n5091), .ZN(n3487)
         );
  AOI211_X1 U4024 ( .C1(n5065), .C2(n3489), .A(n3488), .B(n3487), .ZN(n3490)
         );
  INV_X1 U4025 ( .A(n3490), .ZN(U3250) );
  INV_X1 U4026 ( .A(n3491), .ZN(n4023) );
  AOI21_X1 U4027 ( .B1(n3492), .B2(n4015), .A(n4023), .ZN(n5263) );
  NAND2_X1 U4028 ( .A1(n3499), .A2(n5260), .ZN(n4019) );
  NAND2_X1 U4029 ( .A1(n4157), .A2(n5265), .ZN(n4022) );
  INV_X1 U4030 ( .A(n4022), .ZN(n4018) );
  AOI21_X1 U4031 ( .B1(n5263), .B2(n5261), .A(n4018), .ZN(n3534) );
  NAND2_X1 U4032 ( .A1(n5245), .A2(n3540), .ZN(n3533) );
  NAND2_X1 U4033 ( .A1(n4156), .A2(n3501), .ZN(n3558) );
  XNOR2_X1 U4034 ( .A(n3534), .B(n4077), .ZN(n3495) );
  INV_X1 U4035 ( .A(n4155), .ZN(n3560) );
  AOI22_X1 U4036 ( .A1(n4157), .A2(n5180), .B1(n5365), .B2(n3540), .ZN(n3493)
         );
  OAI21_X1 U4037 ( .B1(n3560), .B2(n5244), .A(n3493), .ZN(n3494) );
  AOI21_X1 U4038 ( .B1(n3495), .B2(n5268), .A(n3494), .ZN(n5284) );
  XNOR2_X1 U4039 ( .A(n3541), .B(n4077), .ZN(n5287) );
  NAND2_X1 U4040 ( .A1(n5287), .A2(n4437), .ZN(n3506) );
  INV_X1 U4041 ( .A(n3500), .ZN(n5258) );
  OAI21_X1 U4042 ( .B1(n5258), .B2(n3501), .A(n3543), .ZN(n5285) );
  INV_X1 U40430 ( .A(n5285), .ZN(n3504) );
  OAI22_X1 U4044 ( .A1(n4450), .A2(n3629), .B1(n3502), .B2(n5231), .ZN(n3503)
         );
  AOI21_X1 U4045 ( .B1(n3504), .B2(n5372), .A(n3503), .ZN(n3505) );
  OAI211_X1 U4046 ( .C1(n5374), .C2(n5284), .A(n3506), .B(n3505), .ZN(U3278)
         );
  NAND2_X1 U4047 ( .A1(n4155), .A2(n3293), .ZN(n3508) );
  MUX2_X1 U4048 ( .A(n5030), .B(DATAI_13_), .S(n4064), .Z(n3559) );
  NAND2_X1 U4049 ( .A1(n3559), .A2(n3815), .ZN(n3507) );
  NAND2_X1 U4050 ( .A1(n3508), .A2(n3507), .ZN(n3509) );
  XNOR2_X1 U4051 ( .A(n3509), .B(n3829), .ZN(n3513) );
  NAND2_X1 U4052 ( .A1(n4155), .A2(n3752), .ZN(n3511) );
  NAND2_X1 U4053 ( .A1(n3559), .A2(n3293), .ZN(n3510) );
  NAND2_X1 U4054 ( .A1(n3511), .A2(n3510), .ZN(n3512) );
  NOR2_X1 U4055 ( .A1(n3513), .A2(n3512), .ZN(n3634) );
  AOI21_X1 U4056 ( .B1(n3513), .B2(n3512), .A(n3634), .ZN(n3520) );
  NAND2_X1 U4057 ( .A1(n3514), .A2(n3515), .ZN(n3518) );
  INV_X1 U4058 ( .A(n3514), .ZN(n3517) );
  INV_X1 U4059 ( .A(n3515), .ZN(n3516) );
  OAI21_X1 U4060 ( .B1(n3520), .B2(n3519), .A(n3636), .ZN(n3521) );
  NAND2_X1 U4061 ( .A1(n3521), .A2(n5314), .ZN(n3532) );
  NAND2_X1 U4062 ( .A1(n4052), .A2(REG2_REG_14__SCAN_IN), .ZN(n3528) );
  OR2_X1 U4063 ( .A1(n4061), .A2(n5300), .ZN(n3527) );
  NAND2_X1 U4064 ( .A1(n3522), .A2(n4572), .ZN(n3523) );
  NAND2_X1 U4065 ( .A1(n3562), .A2(n3523), .ZN(n3862) );
  OR2_X1 U4066 ( .A1(n3835), .A2(n3862), .ZN(n3526) );
  INV_X1 U4067 ( .A(REG0_REG_14__SCAN_IN), .ZN(n3524) );
  OR2_X1 U4068 ( .A1(n2513), .A2(n3524), .ZN(n3525) );
  INV_X1 U4069 ( .A(n5303), .ZN(n4154) );
  NOR2_X1 U4070 ( .A1(STATE_REG_SCAN_IN), .A2(n3529), .ZN(n5027) );
  OAI22_X1 U4071 ( .A1(n5305), .A2(n2596), .B1(n5245), .B2(n5302), .ZN(n3530)
         );
  AOI211_X1 U4072 ( .C1(n5309), .C2(n4154), .A(n5027), .B(n3530), .ZN(n3531)
         );
  OAI211_X1 U4073 ( .C1(n5354), .C2(n3544), .A(n3532), .B(n3531), .ZN(U3231)
         );
  INV_X1 U4074 ( .A(n3533), .ZN(n4020) );
  NOR2_X1 U4075 ( .A1(n3534), .A2(n4020), .ZN(n3561) );
  INV_X1 U4076 ( .A(n3558), .ZN(n3535) );
  NOR2_X1 U4077 ( .A1(n3561), .A2(n3535), .ZN(n3536) );
  NAND2_X1 U4078 ( .A1(n4155), .A2(n3559), .ZN(n3598) );
  INV_X1 U4079 ( .A(n3598), .ZN(n3551) );
  NOR2_X1 U4080 ( .A1(n4155), .A2(n3559), .ZN(n3596) );
  OR2_X1 U4081 ( .A1(n3551), .A2(n3596), .ZN(n3542) );
  XNOR2_X1 U4082 ( .A(n3536), .B(n3542), .ZN(n3537) );
  NAND2_X1 U4083 ( .A1(n3537), .A2(n5268), .ZN(n3539) );
  AOI22_X1 U4084 ( .A1(n4156), .A2(n5180), .B1(n5365), .B2(n3559), .ZN(n3538)
         );
  OAI211_X1 U4085 ( .C1(n5303), .C2(n5244), .A(n3539), .B(n3538), .ZN(n5290)
         );
  INV_X1 U4086 ( .A(n5290), .ZN(n3549) );
  INV_X1 U4087 ( .A(n3542), .ZN(n4101) );
  XNOR2_X1 U4088 ( .A(n3597), .B(n4101), .ZN(n5292) );
  NAND2_X1 U4089 ( .A1(n5292), .A2(n4437), .ZN(n3548) );
  AOI211_X1 U4090 ( .C1(n3559), .C2(n3543), .A(n5333), .B(n3555), .ZN(n5291)
         );
  INV_X1 U4091 ( .A(REG2_REG_13__SCAN_IN), .ZN(n3545) );
  OAI22_X1 U4092 ( .A1(n4450), .A2(n3545), .B1(n3544), .B2(n5231), .ZN(n3546)
         );
  AOI21_X1 U4093 ( .B1(n5291), .B2(n4247), .A(n3546), .ZN(n3547) );
  OAI211_X1 U4094 ( .C1(n5374), .C2(n3549), .A(n3548), .B(n3547), .ZN(U3277)
         );
  INV_X1 U4095 ( .A(n3597), .ZN(n3552) );
  INV_X1 U4096 ( .A(n3596), .ZN(n3550) );
  OAI21_X1 U4097 ( .B1(n3552), .B2(n3551), .A(n3550), .ZN(n3553) );
  MUX2_X1 U4098 ( .A(n5042), .B(DATAI_14_), .S(n4064), .Z(n3859) );
  NAND2_X1 U4099 ( .A1(n5303), .A2(n3859), .ZN(n4025) );
  NAND2_X1 U4100 ( .A1(n4154), .A2(n3637), .ZN(n4031) );
  NAND2_X1 U4101 ( .A1(n4025), .A2(n4031), .ZN(n4073) );
  NAND2_X1 U4102 ( .A1(n3553), .A2(n4073), .ZN(n3609) );
  OAI21_X1 U4103 ( .B1(n3553), .B2(n4073), .A(n3609), .ZN(n3554) );
  INV_X1 U4104 ( .A(n3554), .ZN(n5297) );
  INV_X1 U4105 ( .A(n3555), .ZN(n3556) );
  AOI21_X1 U4106 ( .B1(n3859), .B2(n3556), .A(n3616), .ZN(n5294) );
  OAI22_X1 U4107 ( .A1(n5226), .A2(n5036), .B1(n3862), .B2(n5231), .ZN(n3557)
         );
  AOI21_X1 U4108 ( .B1(n5294), .B2(n5372), .A(n3557), .ZN(n3574) );
  OAI21_X1 U4109 ( .B1(n3560), .B2(n3559), .A(n3558), .ZN(n4026) );
  NAND2_X1 U4110 ( .A1(n3560), .A2(n3559), .ZN(n4024) );
  OAI21_X1 U4111 ( .B1(n3561), .B2(n4026), .A(n4024), .ZN(n3576) );
  XNOR2_X1 U4112 ( .A(n3576), .B(n4073), .ZN(n3572) );
  NAND2_X1 U4113 ( .A1(n4052), .A2(REG2_REG_15__SCAN_IN), .ZN(n3568) );
  OR2_X1 U4114 ( .A1(n4061), .A2(n5324), .ZN(n3567) );
  AND2_X1 U4115 ( .A1(n3562), .A2(n4169), .ZN(n3563) );
  OR2_X1 U4116 ( .A1(n3578), .A2(n3563), .ZN(n5318) );
  OR2_X1 U4117 ( .A1(n3835), .A2(n5318), .ZN(n3566) );
  INV_X1 U4118 ( .A(REG0_REG_15__SCAN_IN), .ZN(n3564) );
  OR2_X1 U4119 ( .A1(n2513), .A2(n3564), .ZN(n3565) );
  NAND4_X1 U4120 ( .A1(n3568), .A2(n3567), .A3(n3566), .A4(n3565), .ZN(n4153)
         );
  NAND2_X1 U4121 ( .A1(n4153), .A2(n5136), .ZN(n3570) );
  NAND2_X1 U4122 ( .A1(n4155), .A2(n5180), .ZN(n3569) );
  NAND2_X1 U4123 ( .A1(n3570), .A2(n3569), .ZN(n3858) );
  AOI21_X1 U4124 ( .B1(n5365), .B2(n3859), .A(n3858), .ZN(n3571) );
  OAI21_X1 U4125 ( .B1(n3572), .B2(n5138), .A(n3571), .ZN(n5299) );
  NAND2_X1 U4126 ( .A1(n5299), .A2(n5226), .ZN(n3573) );
  OAI211_X1 U4127 ( .C1(n5297), .C2(n4399), .A(n3574), .B(n3573), .ZN(U3276)
         );
  INV_X1 U4128 ( .A(n4025), .ZN(n3575) );
  OAI21_X1 U4129 ( .B1(n3576), .B2(n3575), .A(n4031), .ZN(n3612) );
  MUX2_X1 U4130 ( .A(n4924), .B(DATAI_15_), .S(n4064), .Z(n3599) );
  AND2_X1 U4131 ( .A1(n4153), .A2(n5304), .ZN(n3610) );
  NAND2_X1 U4132 ( .A1(n3643), .A2(n3599), .ZN(n4033) );
  OAI21_X1 U4133 ( .B1(n3612), .B2(n3610), .A(n4033), .ZN(n4119) );
  NAND2_X1 U4134 ( .A1(n4052), .A2(REG2_REG_16__SCAN_IN), .ZN(n3582) );
  INV_X1 U4135 ( .A(REG0_REG_16__SCAN_IN), .ZN(n3577) );
  OR2_X1 U4136 ( .A1(n2513), .A2(n3577), .ZN(n3581) );
  OR2_X1 U4137 ( .A1(n4061), .A2(n5329), .ZN(n3580) );
  NAND2_X1 U4138 ( .A1(n3578), .A2(REG3_REG_16__SCAN_IN), .ZN(n3585) );
  OAI21_X1 U4139 ( .B1(n3578), .B2(REG3_REG_16__SCAN_IN), .A(n3585), .ZN(n3918) );
  OR2_X1 U4140 ( .A1(n3835), .A2(n3918), .ZN(n3579) );
  MUX2_X1 U4141 ( .A(n2831), .B(DATAI_16_), .S(n4064), .Z(n4200) );
  INV_X1 U4142 ( .A(n4200), .ZN(n3592) );
  AND2_X1 U4143 ( .A1(n5308), .A2(n3592), .ZN(n4438) );
  NOR2_X1 U4144 ( .A1(n5308), .A2(n3592), .ZN(n4118) );
  OR2_X1 U4145 ( .A1(n4438), .A2(n4118), .ZN(n4099) );
  XNOR2_X1 U4146 ( .A(n4119), .B(n4099), .ZN(n3595) );
  NAND2_X1 U4147 ( .A1(n4052), .A2(REG2_REG_17__SCAN_IN), .ZN(n3591) );
  INV_X1 U4148 ( .A(REG0_REG_17__SCAN_IN), .ZN(n3583) );
  OR2_X1 U4149 ( .A1(n2513), .A2(n3583), .ZN(n3590) );
  INV_X1 U4150 ( .A(n3585), .ZN(n3584) );
  INV_X1 U4151 ( .A(n3666), .ZN(n3668) );
  INV_X1 U4152 ( .A(REG3_REG_17__SCAN_IN), .ZN(n3926) );
  NAND2_X1 U4153 ( .A1(n3926), .A2(n3585), .ZN(n3586) );
  NAND2_X1 U4154 ( .A1(n3668), .A2(n3586), .ZN(n4447) );
  OR2_X1 U4155 ( .A1(n3835), .A2(n4447), .ZN(n3589) );
  OR2_X1 U4156 ( .A1(n4061), .A2(n3587), .ZN(n3588) );
  OAI22_X1 U4157 ( .A1(n3643), .A2(n5246), .B1(n5266), .B2(n3592), .ZN(n3593)
         );
  AOI21_X1 U4158 ( .B1(n5136), .B2(n4201), .A(n3593), .ZN(n3594) );
  OAI21_X1 U4159 ( .B1(n3595), .B2(n5138), .A(n3594), .ZN(n5326) );
  INV_X1 U4160 ( .A(n5326), .ZN(n3607) );
  NOR2_X1 U4161 ( .A1(n3597), .A2(n3596), .ZN(n3602) );
  NAND2_X1 U4162 ( .A1(n5303), .A2(n3637), .ZN(n3608) );
  XNOR2_X1 U4163 ( .A(n2536), .B(n4099), .ZN(n5328) );
  NAND2_X1 U4164 ( .A1(n5328), .A2(n4437), .ZN(n3606) );
  AOI21_X1 U4165 ( .B1(n2540), .B2(n4200), .A(n5333), .ZN(n3603) );
  AND2_X1 U4166 ( .A1(n3603), .A2(n2519), .ZN(n5327) );
  OAI22_X1 U4167 ( .A1(n5226), .A2(n4181), .B1(n3918), .B2(n5231), .ZN(n3604)
         );
  AOI21_X1 U4168 ( .B1(n5327), .B2(n4247), .A(n3604), .ZN(n3605) );
  OAI211_X1 U4169 ( .C1(n5374), .C2(n3607), .A(n3606), .B(n3605), .ZN(U3274)
         );
  NAND2_X1 U4170 ( .A1(n3609), .A2(n3608), .ZN(n3611) );
  INV_X1 U4171 ( .A(n3610), .ZN(n4032) );
  NAND2_X1 U4172 ( .A1(n4032), .A2(n4033), .ZN(n4100) );
  XNOR2_X1 U4173 ( .A(n3611), .B(n4100), .ZN(n5323) );
  INV_X1 U4174 ( .A(n5323), .ZN(n3621) );
  XOR2_X1 U4175 ( .A(n4100), .B(n3612), .Z(n3615) );
  OAI22_X1 U4176 ( .A1(n2706), .A2(n5244), .B1(n5266), .B2(n5304), .ZN(n3613)
         );
  AOI21_X1 U4177 ( .B1(n5180), .B2(n4154), .A(n3613), .ZN(n3614) );
  OAI21_X1 U4178 ( .B1(n3615), .B2(n5138), .A(n3614), .ZN(n5321) );
  NOR2_X1 U4179 ( .A1(n3616), .A2(n5304), .ZN(n5320) );
  INV_X1 U4180 ( .A(n2540), .ZN(n5319) );
  NOR3_X1 U4181 ( .A1(n5320), .A2(n5319), .A3(n4454), .ZN(n3619) );
  INV_X1 U4182 ( .A(REG2_REG_15__SCAN_IN), .ZN(n3617) );
  OAI22_X1 U4183 ( .A1(n4450), .A2(n3617), .B1(n5318), .B2(n5231), .ZN(n3618)
         );
  AOI211_X1 U4184 ( .C1(n5321), .C2(n4450), .A(n3619), .B(n3618), .ZN(n3620)
         );
  OAI21_X1 U4185 ( .B1(n3621), .B2(n4399), .A(n3620), .ZN(U3275) );
  AOI21_X1 U4186 ( .B1(n5288), .B2(n3623), .A(n3622), .ZN(n3632) );
  AOI21_X1 U4187 ( .B1(n5087), .B2(ADDR_REG_12__SCAN_IN), .A(n3624), .ZN(n3625) );
  OAI21_X1 U4188 ( .B1(n3626), .B2(n5069), .A(n3625), .ZN(n3631) );
  AOI211_X1 U4189 ( .C1(n3629), .C2(n3628), .A(n3627), .B(n5091), .ZN(n3630)
         );
  AOI211_X1 U4190 ( .C1(n5065), .C2(n3632), .A(n3631), .B(n3630), .ZN(n3633)
         );
  INV_X1 U4191 ( .A(n3633), .ZN(U3252) );
  INV_X1 U4192 ( .A(n3634), .ZN(n3635) );
  NAND2_X1 U4193 ( .A1(n3636), .A2(n3635), .ZN(n3855) );
  OAI22_X1 U4194 ( .A1(n5303), .A2(n3800), .B1(n3798), .B2(n3637), .ZN(n3639)
         );
  OAI22_X1 U4195 ( .A1(n5303), .A2(n3798), .B1(n3108), .B2(n3637), .ZN(n3638)
         );
  XNOR2_X1 U4196 ( .A(n3638), .B(n3829), .ZN(n3640) );
  XOR2_X1 U4197 ( .A(n3639), .B(n3640), .Z(n3856) );
  NAND2_X1 U4198 ( .A1(n3855), .A2(n3856), .ZN(n3854) );
  NAND2_X1 U4199 ( .A1(n3854), .A2(n3652), .ZN(n3642) );
  OAI22_X1 U4200 ( .A1(n3643), .A2(n3798), .B1(n3108), .B2(n5304), .ZN(n3641)
         );
  XOR2_X1 U4201 ( .A(n3829), .B(n3641), .Z(n3651) );
  NAND2_X1 U4202 ( .A1(n3642), .A2(n3651), .ZN(n5310) );
  OAI22_X1 U4203 ( .A1(n3643), .A2(n3800), .B1(n2511), .B2(n5304), .ZN(n5312)
         );
  NAND2_X1 U4204 ( .A1(n5310), .A2(n5312), .ZN(n3912) );
  NAND2_X1 U4205 ( .A1(n5308), .A2(n3293), .ZN(n3645) );
  NAND2_X1 U4206 ( .A1(n4200), .A2(n3815), .ZN(n3644) );
  NAND2_X1 U4207 ( .A1(n3645), .A2(n3644), .ZN(n3646) );
  XNOR2_X1 U4208 ( .A(n3646), .B(n3829), .ZN(n3650) );
  NAND2_X1 U4209 ( .A1(n5308), .A2(n3752), .ZN(n3648) );
  NAND2_X1 U4210 ( .A1(n4200), .A2(n3293), .ZN(n3647) );
  NAND2_X1 U4211 ( .A1(n3648), .A2(n3647), .ZN(n3649) );
  NOR2_X1 U4212 ( .A1(n3650), .A2(n3649), .ZN(n3655) );
  AOI21_X1 U4213 ( .B1(n3650), .B2(n3649), .A(n3655), .ZN(n3915) );
  INV_X1 U4214 ( .A(n3655), .ZN(n3922) );
  MUX2_X1 U4215 ( .A(n5048), .B(DATAI_17_), .S(n4064), .Z(n4442) );
  INV_X1 U4216 ( .A(n4442), .ZN(n4037) );
  OAI22_X1 U4217 ( .A1(n4418), .A2(n3798), .B1(n3108), .B2(n4037), .ZN(n3656)
         );
  XNOR2_X1 U4218 ( .A(n3656), .B(n3829), .ZN(n3660) );
  INV_X1 U4219 ( .A(n3660), .ZN(n3658) );
  OAI22_X1 U4220 ( .A1(n4418), .A2(n3800), .B1(n2511), .B2(n4037), .ZN(n3661)
         );
  INV_X1 U4221 ( .A(n3661), .ZN(n3657) );
  NAND2_X1 U4222 ( .A1(n3658), .A2(n3657), .ZN(n3659) );
  AND2_X1 U4223 ( .A1(n3922), .A2(n3659), .ZN(n3663) );
  INV_X1 U4224 ( .A(n3659), .ZN(n3662) );
  XOR2_X1 U4225 ( .A(n3661), .B(n3660), .Z(n3925) );
  NAND2_X1 U4226 ( .A1(n4052), .A2(REG2_REG_18__SCAN_IN), .ZN(n3674) );
  INV_X1 U4227 ( .A(REG0_REG_18__SCAN_IN), .ZN(n3664) );
  OR2_X1 U4228 ( .A1(n2513), .A2(n3664), .ZN(n3673) );
  INV_X1 U4229 ( .A(REG1_REG_18__SCAN_IN), .ZN(n3665) );
  OR2_X1 U4230 ( .A1(n4061), .A2(n3665), .ZN(n3672) );
  INV_X1 U4231 ( .A(n3683), .ZN(n3670) );
  INV_X1 U4232 ( .A(REG3_REG_18__SCAN_IN), .ZN(n3667) );
  NAND2_X1 U4233 ( .A1(n3668), .A2(n3667), .ZN(n3669) );
  NAND2_X1 U4234 ( .A1(n3670), .A2(n3669), .ZN(n5353) );
  OR2_X1 U4235 ( .A1(n3835), .A2(n5353), .ZN(n3671) );
  MUX2_X1 U4236 ( .A(n4923), .B(DATAI_18_), .S(n4064), .Z(n5338) );
  OAI22_X1 U4237 ( .A1(n4444), .A2(n3798), .B1(n3108), .B2(n4428), .ZN(n3675)
         );
  XNOR2_X1 U4238 ( .A(n3675), .B(n3829), .ZN(n3678) );
  OR2_X1 U4239 ( .A1(n4444), .A2(n3800), .ZN(n3677) );
  NAND2_X1 U4240 ( .A1(n5338), .A2(n3293), .ZN(n3676) );
  NAND2_X1 U4241 ( .A1(n3677), .A2(n3676), .ZN(n3679) );
  NAND2_X1 U4242 ( .A1(n3678), .A2(n3679), .ZN(n5340) );
  NAND2_X1 U4243 ( .A1(n5346), .A2(n5340), .ZN(n5341) );
  INV_X1 U4244 ( .A(n3678), .ZN(n3681) );
  INV_X1 U4245 ( .A(n3679), .ZN(n3680) );
  NAND2_X1 U4246 ( .A1(n3681), .A2(n3680), .ZN(n5343) );
  NAND2_X1 U4247 ( .A1(n5341), .A2(n5343), .ZN(n3878) );
  NAND2_X1 U4248 ( .A1(n4052), .A2(REG2_REG_19__SCAN_IN), .ZN(n3688) );
  INV_X1 U4249 ( .A(REG0_REG_19__SCAN_IN), .ZN(n3682) );
  OR2_X1 U4250 ( .A1(n2513), .A2(n3682), .ZN(n3687) );
  OAI21_X1 U4251 ( .B1(n3683), .B2(REG3_REG_19__SCAN_IN), .A(n3698), .ZN(n4413) );
  OR2_X1 U4252 ( .A1(n3835), .A2(n4413), .ZN(n3686) );
  INV_X1 U4253 ( .A(REG1_REG_19__SCAN_IN), .ZN(n3684) );
  OR2_X1 U4254 ( .A1(n4061), .A2(n3684), .ZN(n3685) );
  NAND4_X1 U4255 ( .A1(n3688), .A2(n3687), .A3(n3686), .A4(n3685), .ZN(n4419)
         );
  MUX2_X1 U4256 ( .A(n4138), .B(n2973), .S(n4064), .Z(n4403) );
  OAI22_X1 U4257 ( .A1(n4204), .A2(n3800), .B1(n2511), .B2(n4403), .ZN(n3693)
         );
  NAND2_X1 U4258 ( .A1(n4419), .A2(n3293), .ZN(n3690) );
  NAND2_X1 U4259 ( .A1(n4410), .A2(n3815), .ZN(n3689) );
  NAND2_X1 U4260 ( .A1(n3690), .A2(n3689), .ZN(n3691) );
  XNOR2_X1 U4261 ( .A(n3691), .B(n3829), .ZN(n3692) );
  XOR2_X1 U4262 ( .A(n3693), .B(n3692), .Z(n3879) );
  INV_X1 U4263 ( .A(n3692), .ZN(n3695) );
  INV_X1 U4264 ( .A(n3693), .ZN(n3694) );
  NAND2_X1 U4265 ( .A1(n3695), .A2(n3694), .ZN(n3696) );
  NAND2_X1 U4266 ( .A1(n4052), .A2(REG2_REG_20__SCAN_IN), .ZN(n3704) );
  INV_X1 U4267 ( .A(REG1_REG_20__SCAN_IN), .ZN(n3697) );
  OR2_X1 U4268 ( .A1(n4061), .A2(n3697), .ZN(n3703) );
  INV_X1 U4269 ( .A(REG3_REG_20__SCAN_IN), .ZN(n3949) );
  AND2_X1 U4270 ( .A1(n3698), .A2(n3949), .ZN(n3699) );
  OR2_X1 U4271 ( .A1(n3699), .A2(n3713), .ZN(n4393) );
  OR2_X1 U4272 ( .A1(n3835), .A2(n4393), .ZN(n3702) );
  INV_X1 U4273 ( .A(REG0_REG_20__SCAN_IN), .ZN(n3700) );
  OR2_X1 U4274 ( .A1(n2513), .A2(n3700), .ZN(n3701) );
  INV_X1 U4275 ( .A(n4390), .ZN(n4386) );
  OAI22_X1 U4276 ( .A1(n4365), .A2(n3798), .B1(n3108), .B2(n4386), .ZN(n3705)
         );
  XNOR2_X1 U4277 ( .A(n3705), .B(n3829), .ZN(n3708) );
  OR2_X1 U4278 ( .A1(n4365), .A2(n3800), .ZN(n3707) );
  NAND2_X1 U4279 ( .A1(n4390), .A2(n3293), .ZN(n3706) );
  NAND2_X1 U4280 ( .A1(n3707), .A2(n3706), .ZN(n3709) );
  NAND2_X1 U4281 ( .A1(n3708), .A2(n3709), .ZN(n3943) );
  INV_X1 U4282 ( .A(n3708), .ZN(n3711) );
  INV_X1 U4283 ( .A(n3709), .ZN(n3710) );
  NAND2_X1 U4284 ( .A1(n3711), .A2(n3710), .ZN(n3944) );
  INV_X1 U4285 ( .A(n3893), .ZN(n3725) );
  NAND2_X1 U4286 ( .A1(n4052), .A2(REG2_REG_21__SCAN_IN), .ZN(n3719) );
  INV_X1 U4287 ( .A(REG1_REG_21__SCAN_IN), .ZN(n3712) );
  OR2_X1 U4288 ( .A1(n4061), .A2(n3712), .ZN(n3718) );
  OR2_X1 U4289 ( .A1(n3713), .A2(REG3_REG_21__SCAN_IN), .ZN(n3714) );
  NAND2_X1 U4290 ( .A1(n3732), .A2(n3714), .ZN(n4362) );
  OR2_X1 U4291 ( .A1(n3835), .A2(n4362), .ZN(n3717) );
  INV_X1 U4292 ( .A(REG0_REG_21__SCAN_IN), .ZN(n3715) );
  OR2_X1 U4293 ( .A1(n2513), .A2(n3715), .ZN(n3716) );
  NAND4_X1 U4294 ( .A1(n3719), .A2(n3718), .A3(n3717), .A4(n3716), .ZN(n4208)
         );
  NAND2_X1 U4295 ( .A1(n4208), .A2(n3293), .ZN(n3721) );
  NAND2_X1 U4296 ( .A1(n4064), .A2(DATAI_21_), .ZN(n4364) );
  NAND2_X1 U4297 ( .A1(n4361), .A2(n3815), .ZN(n3720) );
  NAND2_X1 U4298 ( .A1(n3721), .A2(n3720), .ZN(n3722) );
  XNOR2_X1 U4299 ( .A(n3722), .B(n3782), .ZN(n3726) );
  NOR2_X1 U4300 ( .A1(n4364), .A2(n3798), .ZN(n3723) );
  AOI21_X1 U4301 ( .B1(n4208), .B2(n3752), .A(n3723), .ZN(n3727) );
  AND2_X1 U4302 ( .A1(n3726), .A2(n3727), .ZN(n3890) );
  INV_X1 U4303 ( .A(n3890), .ZN(n3724) );
  NAND2_X1 U4304 ( .A1(n3725), .A2(n3724), .ZN(n3730) );
  INV_X1 U4305 ( .A(n3726), .ZN(n3729) );
  INV_X1 U4306 ( .A(n3727), .ZN(n3728) );
  NAND2_X1 U4307 ( .A1(n3729), .A2(n3728), .ZN(n3889) );
  NAND2_X1 U4308 ( .A1(n3730), .A2(n3889), .ZN(n3957) );
  INV_X1 U4309 ( .A(n3957), .ZN(n3742) );
  NAND2_X1 U4310 ( .A1(n4052), .A2(REG2_REG_22__SCAN_IN), .ZN(n3738) );
  INV_X1 U4311 ( .A(REG1_REG_22__SCAN_IN), .ZN(n3731) );
  OR2_X1 U4312 ( .A1(n4061), .A2(n3731), .ZN(n3737) );
  INV_X1 U4313 ( .A(REG3_REG_22__SCAN_IN), .ZN(n3959) );
  NAND2_X1 U4314 ( .A1(n3732), .A2(n3959), .ZN(n3733) );
  NAND2_X1 U4315 ( .A1(n3744), .A2(n3733), .ZN(n4346) );
  INV_X1 U4316 ( .A(REG0_REG_22__SCAN_IN), .ZN(n3734) );
  OR2_X1 U4317 ( .A1(n2513), .A2(n3734), .ZN(n3735) );
  NAND4_X1 U4318 ( .A1(n3738), .A2(n3737), .A3(n3736), .A4(n3735), .ZN(n4371)
         );
  NAND2_X1 U4319 ( .A1(n4064), .A2(DATAI_22_), .ZN(n4351) );
  INV_X1 U4320 ( .A(n4351), .ZN(n4345) );
  AOI22_X1 U4321 ( .A1(n4371), .A2(n3740), .B1(n3815), .B2(n4345), .ZN(n3739)
         );
  XNOR2_X1 U4322 ( .A(n3739), .B(n3829), .ZN(n3754) );
  AOI22_X1 U4323 ( .A1(n4371), .A2(n3752), .B1(n3740), .B2(n4345), .ZN(n3755)
         );
  XNOR2_X1 U4324 ( .A(n3754), .B(n3755), .ZN(n3958) );
  NAND2_X1 U4325 ( .A1(n4052), .A2(REG2_REG_23__SCAN_IN), .ZN(n3750) );
  INV_X1 U4326 ( .A(REG1_REG_23__SCAN_IN), .ZN(n3743) );
  OR2_X1 U4327 ( .A1(n4061), .A2(n3743), .ZN(n3749) );
  INV_X1 U4328 ( .A(REG3_REG_23__SCAN_IN), .ZN(n4762) );
  NAND2_X1 U4329 ( .A1(n3744), .A2(n4762), .ZN(n3745) );
  NAND2_X1 U4330 ( .A1(n3762), .A2(n3745), .ZN(n4336) );
  OR2_X1 U4331 ( .A1(n3835), .A2(n4336), .ZN(n3748) );
  INV_X1 U4332 ( .A(REG0_REG_23__SCAN_IN), .ZN(n3746) );
  OR2_X1 U4333 ( .A1(n2513), .A2(n3746), .ZN(n3747) );
  NAND4_X1 U4334 ( .A1(n3750), .A2(n3749), .A3(n3748), .A4(n3747), .ZN(n4354)
         );
  NAND2_X1 U4335 ( .A1(n4064), .A2(DATAI_23_), .ZN(n4333) );
  NOR2_X1 U4336 ( .A1(n4333), .A2(n2511), .ZN(n3751) );
  AOI21_X1 U4337 ( .B1(n4354), .B2(n3752), .A(n3751), .ZN(n3760) );
  INV_X1 U4338 ( .A(n4354), .ZN(n4315) );
  OAI22_X1 U4339 ( .A1(n4315), .A2(n3798), .B1(n3108), .B2(n4333), .ZN(n3753)
         );
  XNOR2_X1 U4340 ( .A(n3753), .B(n3829), .ZN(n3759) );
  XOR2_X1 U4341 ( .A(n3760), .B(n3759), .Z(n3867) );
  INV_X1 U4342 ( .A(n3754), .ZN(n3757) );
  INV_X1 U4343 ( .A(n3755), .ZN(n3756) );
  NOR2_X1 U4344 ( .A1(n3757), .A2(n3756), .ZN(n3868) );
  NOR2_X1 U4345 ( .A1(n3867), .A2(n3868), .ZN(n3758) );
  INV_X1 U4346 ( .A(n3759), .ZN(n3761) );
  OR2_X1 U4347 ( .A1(n3761), .A2(n3760), .ZN(n3772) );
  NAND2_X1 U4348 ( .A1(n3028), .A2(REG1_REG_24__SCAN_IN), .ZN(n3768) );
  INV_X1 U4349 ( .A(REG2_REG_24__SCAN_IN), .ZN(n4321) );
  INV_X1 U4350 ( .A(REG3_REG_24__SCAN_IN), .ZN(n4781) );
  NAND2_X1 U4351 ( .A1(n3762), .A2(n4781), .ZN(n3763) );
  NAND2_X1 U4352 ( .A1(n3775), .A2(n3763), .ZN(n4320) );
  INV_X1 U4353 ( .A(REG0_REG_24__SCAN_IN), .ZN(n3764) );
  OR2_X1 U4354 ( .A1(n2513), .A2(n3764), .ZN(n3765) );
  NAND4_X1 U4355 ( .A1(n3768), .A2(n3767), .A3(n3766), .A4(n3765), .ZN(n4152)
         );
  NAND2_X1 U4356 ( .A1(n4152), .A2(n3293), .ZN(n3770) );
  NAND2_X1 U4357 ( .A1(n4064), .A2(DATAI_24_), .ZN(n4314) );
  INV_X1 U4358 ( .A(n4314), .ZN(n4049) );
  NAND2_X1 U4359 ( .A1(n4049), .A2(n3815), .ZN(n3769) );
  NAND2_X1 U4360 ( .A1(n3770), .A2(n3769), .ZN(n3771) );
  XNOR2_X1 U4361 ( .A(n3771), .B(n3782), .ZN(n3773) );
  OAI22_X1 U4362 ( .A1(n4330), .A2(n3800), .B1(n2511), .B2(n4314), .ZN(n3935)
         );
  NAND3_X1 U4363 ( .A1(n3869), .A2(n3773), .A3(n3772), .ZN(n3932) );
  NAND2_X1 U4364 ( .A1(n3028), .A2(REG1_REG_25__SCAN_IN), .ZN(n3781) );
  INV_X1 U4365 ( .A(REG2_REG_25__SCAN_IN), .ZN(n4294) );
  OR2_X1 U4366 ( .A1(n3026), .A2(n4294), .ZN(n3780) );
  INV_X1 U4367 ( .A(n3775), .ZN(n3774) );
  INV_X1 U4368 ( .A(REG3_REG_25__SCAN_IN), .ZN(n4777) );
  NAND2_X1 U4369 ( .A1(n3775), .A2(n4777), .ZN(n3776) );
  NAND2_X1 U4370 ( .A1(n3791), .A2(n3776), .ZN(n4293) );
  INV_X1 U4371 ( .A(REG0_REG_25__SCAN_IN), .ZN(n3777) );
  OR2_X1 U4372 ( .A1(n2513), .A2(n3777), .ZN(n3778) );
  INV_X1 U4373 ( .A(n4292), .ZN(n4301) );
  OAI22_X1 U4374 ( .A1(n4313), .A2(n2511), .B1(n4301), .B2(n3108), .ZN(n3783)
         );
  XNOR2_X1 U4375 ( .A(n3783), .B(n3782), .ZN(n3786) );
  OR2_X1 U4376 ( .A1(n4313), .A2(n3800), .ZN(n3785) );
  NAND2_X1 U4377 ( .A1(n4292), .A2(n3293), .ZN(n3784) );
  AND2_X1 U4378 ( .A1(n3785), .A2(n3784), .ZN(n3787) );
  AND2_X1 U4379 ( .A1(n3786), .A2(n3787), .ZN(n3901) );
  INV_X1 U4380 ( .A(n3786), .ZN(n3789) );
  INV_X1 U4381 ( .A(n3787), .ZN(n3788) );
  NAND2_X1 U4382 ( .A1(n3789), .A2(n3788), .ZN(n3902) );
  OAI21_X1 U4383 ( .B1(n3905), .B2(n3901), .A(n3902), .ZN(n3979) );
  INV_X1 U4384 ( .A(n3979), .ZN(n3804) );
  NAND2_X1 U4385 ( .A1(n4052), .A2(REG2_REG_26__SCAN_IN), .ZN(n3797) );
  INV_X1 U4386 ( .A(REG1_REG_26__SCAN_IN), .ZN(n3790) );
  OR2_X1 U4387 ( .A1(n4061), .A2(n3790), .ZN(n3796) );
  INV_X1 U4388 ( .A(REG3_REG_26__SCAN_IN), .ZN(n3981) );
  NAND2_X1 U4389 ( .A1(n3791), .A2(n3981), .ZN(n3792) );
  NAND2_X1 U4390 ( .A1(n3807), .A2(n3792), .ZN(n4283) );
  INV_X1 U4391 ( .A(REG0_REG_26__SCAN_IN), .ZN(n3793) );
  OR2_X1 U4392 ( .A1(n2513), .A2(n3793), .ZN(n3794) );
  NAND2_X1 U4393 ( .A1(n4064), .A2(DATAI_26_), .ZN(n4282) );
  OAI22_X1 U4394 ( .A1(n4214), .A2(n3798), .B1(n3108), .B2(n4282), .ZN(n3799)
         );
  XNOR2_X1 U4395 ( .A(n3799), .B(n3829), .ZN(n3976) );
  OR2_X1 U4396 ( .A1(n4214), .A2(n3800), .ZN(n3802) );
  NAND2_X1 U4397 ( .A1(n4228), .A2(n3293), .ZN(n3801) );
  NAND2_X1 U4398 ( .A1(n3802), .A2(n3801), .ZN(n3977) );
  NAND2_X1 U4399 ( .A1(n3976), .A2(n3977), .ZN(n3803) );
  NAND2_X1 U4400 ( .A1(n4052), .A2(REG2_REG_27__SCAN_IN), .ZN(n3813) );
  INV_X1 U4401 ( .A(REG1_REG_27__SCAN_IN), .ZN(n3805) );
  OR2_X1 U4402 ( .A1(n4061), .A2(n3805), .ZN(n3812) );
  INV_X1 U4403 ( .A(n3807), .ZN(n3806) );
  NAND2_X1 U4404 ( .A1(n3806), .A2(REG3_REG_27__SCAN_IN), .ZN(n3822) );
  INV_X1 U4405 ( .A(REG3_REG_27__SCAN_IN), .ZN(n4755) );
  NAND2_X1 U4406 ( .A1(n3807), .A2(n4755), .ZN(n3808) );
  NAND2_X1 U4407 ( .A1(n3822), .A2(n3808), .ZN(n4267) );
  INV_X1 U4408 ( .A(REG0_REG_27__SCAN_IN), .ZN(n3809) );
  OR2_X1 U4409 ( .A1(n2513), .A2(n3809), .ZN(n3810) );
  AND2_X1 U4410 ( .A1(n4064), .A2(DATAI_27_), .ZN(n4217) );
  OAI22_X1 U4411 ( .A1(n4276), .A2(n3110), .B1(n2511), .B2(n4266), .ZN(n3820)
         );
  NAND2_X1 U4412 ( .A1(n4218), .A2(n3293), .ZN(n3817) );
  NAND2_X1 U4413 ( .A1(n4217), .A2(n3815), .ZN(n3816) );
  NAND2_X1 U4414 ( .A1(n3817), .A2(n3816), .ZN(n3818) );
  XNOR2_X1 U4415 ( .A(n3818), .B(n3829), .ZN(n3819) );
  XOR2_X1 U4416 ( .A(n3820), .B(n3819), .Z(n3846) );
  NAND2_X1 U4417 ( .A1(n4052), .A2(REG2_REG_28__SCAN_IN), .ZN(n3828) );
  INV_X1 U4418 ( .A(REG1_REG_28__SCAN_IN), .ZN(n3821) );
  OR2_X1 U4419 ( .A1(n4061), .A2(n3821), .ZN(n3827) );
  INV_X1 U4420 ( .A(REG3_REG_28__SCAN_IN), .ZN(n4579) );
  NAND2_X1 U4421 ( .A1(n3822), .A2(n4579), .ZN(n3823) );
  NAND2_X1 U4422 ( .A1(n4231), .A2(n3823), .ZN(n4248) );
  INV_X1 U4423 ( .A(REG0_REG_28__SCAN_IN), .ZN(n3824) );
  OR2_X1 U4424 ( .A1(n2513), .A2(n3824), .ZN(n3825) );
  AND2_X1 U4425 ( .A1(n4064), .A2(DATAI_28_), .ZN(n4221) );
  OAI22_X1 U4426 ( .A1(n4255), .A2(n2511), .B1(n3108), .B2(n4246), .ZN(n3830)
         );
  XNOR2_X1 U4427 ( .A(n3830), .B(n3829), .ZN(n3832) );
  OAI22_X1 U4428 ( .A1(n4255), .A2(n3800), .B1(n2511), .B2(n4246), .ZN(n3831)
         );
  XNOR2_X1 U4429 ( .A(n3832), .B(n3831), .ZN(n3833) );
  AOI22_X1 U4430 ( .A1(n4221), .A2(n3972), .B1(n3980), .B2(n4218), .ZN(n3843)
         );
  NAND2_X1 U4431 ( .A1(n4052), .A2(REG2_REG_29__SCAN_IN), .ZN(n3840) );
  INV_X1 U4432 ( .A(REG1_REG_29__SCAN_IN), .ZN(n3834) );
  OR2_X1 U4433 ( .A1(n4061), .A2(n3834), .ZN(n3839) );
  OR2_X1 U4434 ( .A1(n3835), .A2(n4231), .ZN(n3838) );
  INV_X1 U4435 ( .A(REG0_REG_29__SCAN_IN), .ZN(n3836) );
  OR2_X1 U4436 ( .A1(n2513), .A2(n3836), .ZN(n3837) );
  OAI22_X1 U4437 ( .A1(n3982), .A2(n4242), .B1(STATE_REG_SCAN_IN), .B2(n4579), 
        .ZN(n3841) );
  INV_X1 U4438 ( .A(n3841), .ZN(n3842) );
  OAI211_X1 U4439 ( .C1(n5354), .C2(n4248), .A(n3843), .B(n3842), .ZN(n3844)
         );
  INV_X1 U4440 ( .A(n3844), .ZN(n3845) );
  XNOR2_X1 U4441 ( .A(n3847), .B(n3846), .ZN(n3853) );
  AOI22_X1 U4442 ( .A1(n4217), .A2(n5339), .B1(n3980), .B2(n4303), .ZN(n3850)
         );
  OAI22_X1 U4443 ( .A1(n3982), .A2(n4255), .B1(STATE_REG_SCAN_IN), .B2(n4755), 
        .ZN(n3848) );
  INV_X1 U4444 ( .A(n3848), .ZN(n3849) );
  OAI211_X1 U4445 ( .C1(n5354), .C2(n4267), .A(n3850), .B(n3849), .ZN(n3851)
         );
  INV_X1 U4446 ( .A(n3851), .ZN(n3852) );
  OAI21_X1 U4447 ( .B1(n3853), .B2(n5344), .A(n3852), .ZN(U3211) );
  OAI21_X1 U4448 ( .B1(n3856), .B2(n3855), .A(n3854), .ZN(n3864) );
  NAND2_X1 U4449 ( .A1(REG3_REG_14__SCAN_IN), .A2(U3149), .ZN(n5043) );
  INV_X1 U4450 ( .A(n5043), .ZN(n3857) );
  AOI21_X1 U4451 ( .B1(n3858), .B2(n5348), .A(n3857), .ZN(n3861) );
  NAND2_X1 U4452 ( .A1(n5339), .A2(n3859), .ZN(n3860) );
  OAI211_X1 U4453 ( .C1(n5354), .C2(n3862), .A(n3861), .B(n3860), .ZN(n3863)
         );
  AOI21_X1 U4454 ( .B1(n3864), .B2(n5314), .A(n3863), .ZN(n3865) );
  INV_X1 U4455 ( .A(n3865), .ZN(U3212) );
  INV_X1 U4456 ( .A(n3866), .ZN(n3956) );
  OAI21_X1 U4457 ( .B1(n3956), .B2(n3868), .A(n3867), .ZN(n3870) );
  NAND3_X1 U4458 ( .A1(n3870), .A2(n5314), .A3(n3869), .ZN(n3876) );
  INV_X1 U4459 ( .A(n4371), .ZN(n3871) );
  OAI22_X1 U4460 ( .A1(n5302), .A2(n3871), .B1(STATE_REG_SCAN_IN), .B2(n4762), 
        .ZN(n3872) );
  INV_X1 U4461 ( .A(n3872), .ZN(n3875) );
  INV_X1 U4462 ( .A(n4333), .ZN(n4328) );
  AOI22_X1 U4463 ( .A1(n4328), .A2(n5339), .B1(n5309), .B2(n4152), .ZN(n3874)
         );
  OR2_X1 U4464 ( .A1(n5354), .A2(n4336), .ZN(n3873) );
  NAND4_X1 U4465 ( .A1(n3876), .A2(n3875), .A3(n3874), .A4(n3873), .ZN(U3213)
         );
  OAI21_X1 U4466 ( .B1(n3879), .B2(n3878), .A(n3877), .ZN(n3887) );
  OR2_X1 U4467 ( .A1(n4365), .A2(n5244), .ZN(n3881) );
  OR2_X1 U4468 ( .A1(n4444), .A2(n5246), .ZN(n3880) );
  NAND2_X1 U4469 ( .A1(n3881), .A2(n3880), .ZN(n4404) );
  INV_X1 U4470 ( .A(n3882), .ZN(n3883) );
  AOI21_X1 U4471 ( .B1(n4404), .B2(n5348), .A(n3883), .ZN(n3885) );
  NAND2_X1 U4472 ( .A1(n5339), .A2(n4410), .ZN(n3884) );
  OAI211_X1 U4473 ( .C1(n5354), .C2(n4413), .A(n3885), .B(n3884), .ZN(n3886)
         );
  AOI21_X1 U4474 ( .B1(n3887), .B2(n5314), .A(n3886), .ZN(n3888) );
  INV_X1 U4475 ( .A(n3888), .ZN(U3216) );
  INV_X1 U4476 ( .A(n3889), .ZN(n3891) );
  NOR2_X1 U4477 ( .A1(n3891), .A2(n3890), .ZN(n3892) );
  XNOR2_X1 U4478 ( .A(n3893), .B(n3892), .ZN(n3899) );
  AOI22_X1 U4479 ( .A1(n4361), .A2(n3972), .B1(n5309), .B2(n4371), .ZN(n3897)
         );
  INV_X1 U4480 ( .A(REG3_REG_21__SCAN_IN), .ZN(n3894) );
  OAI22_X1 U4481 ( .A1(n5302), .A2(n4365), .B1(STATE_REG_SCAN_IN), .B2(n3894), 
        .ZN(n3895) );
  INV_X1 U4482 ( .A(n3895), .ZN(n3896) );
  OAI211_X1 U4483 ( .C1(n5354), .C2(n4362), .A(n3897), .B(n3896), .ZN(n3898)
         );
  AOI21_X1 U4484 ( .B1(n3899), .B2(n5314), .A(n3898), .ZN(n3900) );
  INV_X1 U4485 ( .A(n3900), .ZN(U3220) );
  INV_X1 U4486 ( .A(n3901), .ZN(n3903) );
  NAND2_X1 U4487 ( .A1(n3903), .A2(n3902), .ZN(n3904) );
  XNOR2_X1 U4488 ( .A(n3905), .B(n3904), .ZN(n3911) );
  AOI22_X1 U4489 ( .A1(n4292), .A2(n5339), .B1(n5309), .B2(n4303), .ZN(n3908)
         );
  OAI22_X1 U4490 ( .A1(n5302), .A2(n4330), .B1(STATE_REG_SCAN_IN), .B2(n4777), 
        .ZN(n3906) );
  INV_X1 U4491 ( .A(n3906), .ZN(n3907) );
  OAI211_X1 U4492 ( .C1(n5354), .C2(n4293), .A(n3908), .B(n3907), .ZN(n3909)
         );
  INV_X1 U4493 ( .A(n3909), .ZN(n3910) );
  OAI21_X1 U4494 ( .B1(n3911), .B2(n5344), .A(n3910), .ZN(U3222) );
  AND2_X1 U4495 ( .A1(n3912), .A2(n5311), .ZN(n3914) );
  OAI21_X1 U4496 ( .B1(n3915), .B2(n3914), .A(n3913), .ZN(n3920) );
  AOI22_X1 U4497 ( .A1(n4200), .A2(n3972), .B1(n5309), .B2(n4201), .ZN(n3917)
         );
  INV_X1 U4498 ( .A(REG3_REG_16__SCAN_IN), .ZN(n4590) );
  NOR2_X1 U4499 ( .A1(STATE_REG_SCAN_IN), .A2(n4590), .ZN(n4184) );
  AOI21_X1 U4500 ( .B1(n3980), .B2(n4153), .A(n4184), .ZN(n3916) );
  OAI211_X1 U4501 ( .C1(n3918), .C2(n5354), .A(n3917), .B(n3916), .ZN(n3919)
         );
  AOI21_X1 U4502 ( .B1(n3920), .B2(n5314), .A(n3919), .ZN(n3921) );
  INV_X1 U4503 ( .A(n3921), .ZN(U3223) );
  NAND2_X1 U4504 ( .A1(n3913), .A2(n3922), .ZN(n3924) );
  NAND2_X1 U4505 ( .A1(n3924), .A2(n3925), .ZN(n3923) );
  OAI21_X1 U4506 ( .B1(n3925), .B2(n3924), .A(n3923), .ZN(n3930) );
  AOI22_X1 U4507 ( .A1(n4442), .A2(n3972), .B1(n5309), .B2(n4202), .ZN(n3928)
         );
  NOR2_X1 U4508 ( .A1(STATE_REG_SCAN_IN), .A2(n3926), .ZN(n5053) );
  AOI21_X1 U4509 ( .B1(n3980), .B2(n5308), .A(n5053), .ZN(n3927) );
  OAI211_X1 U4510 ( .C1(n5354), .C2(n4447), .A(n3928), .B(n3927), .ZN(n3929)
         );
  AOI21_X1 U4511 ( .B1(n3930), .B2(n5314), .A(n3929), .ZN(n3931) );
  INV_X1 U4512 ( .A(n3931), .ZN(U3225) );
  INV_X1 U4513 ( .A(n3932), .ZN(n3934) );
  NOR2_X1 U4514 ( .A1(n3934), .A2(n3933), .ZN(n3936) );
  XNOR2_X1 U4515 ( .A(n3936), .B(n3935), .ZN(n3942) );
  AOI22_X1 U4516 ( .A1(n4049), .A2(n5339), .B1(n5309), .B2(n4212), .ZN(n3939)
         );
  OAI22_X1 U4517 ( .A1(n5302), .A2(n4315), .B1(STATE_REG_SCAN_IN), .B2(n4781), 
        .ZN(n3937) );
  INV_X1 U4518 ( .A(n3937), .ZN(n3938) );
  OAI211_X1 U4519 ( .C1(n5354), .C2(n4320), .A(n3939), .B(n3938), .ZN(n3940)
         );
  INV_X1 U4520 ( .A(n3940), .ZN(n3941) );
  OAI21_X1 U4521 ( .B1(n3942), .B2(n5344), .A(n3941), .ZN(U3226) );
  NAND2_X1 U4522 ( .A1(n3944), .A2(n3943), .ZN(n3946) );
  XOR2_X1 U4523 ( .A(n3946), .B(n3945), .Z(n3954) );
  NAND2_X1 U4524 ( .A1(n4208), .A2(n5136), .ZN(n3948) );
  NAND2_X1 U4525 ( .A1(n4419), .A2(n5180), .ZN(n3947) );
  NAND2_X1 U4526 ( .A1(n3948), .A2(n3947), .ZN(n4387) );
  NOR2_X1 U4527 ( .A1(n3949), .A2(STATE_REG_SCAN_IN), .ZN(n3950) );
  AOI21_X1 U4528 ( .B1(n4387), .B2(n5348), .A(n3950), .ZN(n3952) );
  NAND2_X1 U4529 ( .A1(n5339), .A2(n4390), .ZN(n3951) );
  OAI211_X1 U4530 ( .C1(n5354), .C2(n4393), .A(n3952), .B(n3951), .ZN(n3953)
         );
  AOI21_X1 U4531 ( .B1(n3954), .B2(n5314), .A(n3953), .ZN(n3955) );
  INV_X1 U4532 ( .A(n3955), .ZN(U3230) );
  AOI21_X1 U4533 ( .B1(n3958), .B2(n3957), .A(n3956), .ZN(n3965) );
  INV_X1 U4534 ( .A(n4346), .ZN(n3963) );
  INV_X1 U4535 ( .A(n5354), .ZN(n3962) );
  INV_X1 U4536 ( .A(n4208), .ZN(n4352) );
  OAI22_X1 U4537 ( .A1(n5302), .A2(n4352), .B1(STATE_REG_SCAN_IN), .B2(n3959), 
        .ZN(n3961) );
  OAI22_X1 U4538 ( .A1(n5305), .A2(n4351), .B1(n4315), .B2(n3982), .ZN(n3960)
         );
  AOI211_X1 U4539 ( .C1(n3963), .C2(n3962), .A(n3961), .B(n3960), .ZN(n3964)
         );
  OAI21_X1 U4540 ( .B1(n3965), .B2(n5344), .A(n3964), .ZN(U3232) );
  OAI21_X1 U4541 ( .B1(n3968), .B2(n3967), .A(n3966), .ZN(n3969) );
  NAND2_X1 U4542 ( .A1(n3969), .A2(n5314), .ZN(n3975) );
  AOI22_X1 U4543 ( .A1(n5309), .A2(n4163), .B1(n3980), .B2(n5103), .ZN(n3974)
         );
  AOI22_X1 U4544 ( .A1(n3972), .A2(n3971), .B1(REG3_REG_2__SCAN_IN), .B2(n3970), .ZN(n3973) );
  NAND3_X1 U4545 ( .A1(n3975), .A2(n3974), .A3(n3973), .ZN(U3234) );
  XOR2_X1 U4546 ( .A(n3977), .B(n3976), .Z(n3978) );
  XNOR2_X1 U4547 ( .A(n3979), .B(n3978), .ZN(n3988) );
  AOI22_X1 U4548 ( .A1(n4228), .A2(n5339), .B1(n3980), .B2(n4212), .ZN(n3985)
         );
  OAI22_X1 U4549 ( .A1(n3982), .A2(n4276), .B1(STATE_REG_SCAN_IN), .B2(n3981), 
        .ZN(n3983) );
  INV_X1 U4550 ( .A(n3983), .ZN(n3984) );
  OAI211_X1 U4551 ( .C1(n5354), .C2(n4283), .A(n3985), .B(n3984), .ZN(n3986)
         );
  INV_X1 U4552 ( .A(n3986), .ZN(n3987) );
  OAI21_X1 U4553 ( .B1(n3988), .B2(n5344), .A(n3987), .ZN(U3237) );
  INV_X1 U4554 ( .A(n5112), .ZN(n4145) );
  NOR2_X1 U4555 ( .A1(n4371), .A2(n4351), .ZN(n4123) );
  NAND2_X1 U4556 ( .A1(n4354), .A2(n4333), .ZN(n4127) );
  NAND2_X1 U4557 ( .A1(n4165), .A2(n5105), .ZN(n4108) );
  OAI211_X1 U4558 ( .C1(n2560), .C2(n4921), .A(n4108), .B(n3989), .ZN(n3992)
         );
  NAND3_X1 U4559 ( .A1(n3992), .A2(n3991), .A3(n3990), .ZN(n3995) );
  NAND3_X1 U4560 ( .A1(n3995), .A2(n3994), .A3(n3993), .ZN(n3998) );
  NAND3_X1 U4561 ( .A1(n3998), .A2(n3997), .A3(n3996), .ZN(n4001) );
  NAND3_X1 U4562 ( .A1(n4001), .A2(n4000), .A3(n3999), .ZN(n4005) );
  INV_X1 U4563 ( .A(n4002), .ZN(n4003) );
  AOI21_X1 U4564 ( .B1(n4005), .B2(n4004), .A(n4003), .ZN(n4011) );
  NAND2_X1 U4565 ( .A1(n4007), .A2(n4006), .ZN(n4010) );
  OAI211_X1 U4566 ( .C1(n4011), .C2(n4010), .A(n4009), .B(n4008), .ZN(n4013)
         );
  OAI211_X1 U4567 ( .C1(n4160), .C2(n4014), .A(n4013), .B(n4012), .ZN(n4030)
         );
  INV_X1 U4568 ( .A(n4015), .ZN(n4017) );
  NOR4_X1 U4569 ( .A1(n4026), .A2(n4018), .A3(n4017), .A4(n4016), .ZN(n4029)
         );
  INV_X1 U4570 ( .A(n4019), .ZN(n4021) );
  AOI211_X1 U4571 ( .C1(n4023), .C2(n4022), .A(n4021), .B(n4020), .ZN(n4027)
         );
  OAI211_X1 U4572 ( .C1(n4027), .C2(n4026), .A(n4025), .B(n4024), .ZN(n4028)
         );
  AOI21_X1 U4573 ( .B1(n4030), .B2(n4029), .A(n4028), .ZN(n4036) );
  NAND2_X1 U4574 ( .A1(n4032), .A2(n4031), .ZN(n4035) );
  INV_X1 U4575 ( .A(n4118), .ZN(n4034) );
  OAI211_X1 U4576 ( .C1(n4036), .C2(n4035), .A(n4034), .B(n4033), .ZN(n4042)
         );
  NAND2_X1 U4577 ( .A1(n4201), .A2(n4037), .ZN(n4076) );
  INV_X1 U4578 ( .A(n4076), .ZN(n4038) );
  NOR2_X1 U4579 ( .A1(n4438), .A2(n4038), .ZN(n4378) );
  NAND2_X1 U4580 ( .A1(n4202), .A2(n4428), .ZN(n4400) );
  NAND2_X1 U4581 ( .A1(n4419), .A2(n4403), .ZN(n4039) );
  AND2_X1 U4582 ( .A1(n4400), .A2(n4039), .ZN(n4383) );
  NAND2_X1 U4583 ( .A1(n4206), .A2(n4386), .ZN(n4086) );
  NAND3_X1 U4584 ( .A1(n4378), .A2(n4383), .A3(n4086), .ZN(n4121) );
  INV_X1 U4585 ( .A(n4121), .ZN(n4041) );
  NAND2_X1 U4586 ( .A1(n4352), .A2(n4361), .ZN(n4106) );
  INV_X1 U4587 ( .A(n4106), .ZN(n4040) );
  AOI21_X1 U4588 ( .B1(n4042), .B2(n4041), .A(n4040), .ZN(n4046) );
  NAND2_X1 U4589 ( .A1(n4418), .A2(n4442), .ZN(n4376) );
  NAND2_X1 U4590 ( .A1(n4444), .A2(n5338), .ZN(n4380) );
  NAND2_X1 U4591 ( .A1(n4376), .A2(n4380), .ZN(n4043) );
  NAND2_X1 U4592 ( .A1(n4043), .A2(n4383), .ZN(n4044) );
  NAND2_X1 U4593 ( .A1(n4365), .A2(n4390), .ZN(n4087) );
  NAND2_X1 U4594 ( .A1(n4204), .A2(n4410), .ZN(n4381) );
  NAND3_X1 U4595 ( .A1(n4044), .A2(n4087), .A3(n4381), .ZN(n4045) );
  NAND2_X1 U4596 ( .A1(n4045), .A2(n4086), .ZN(n4120) );
  AND2_X1 U4597 ( .A1(n4371), .A2(n4351), .ZN(n4124) );
  AND2_X1 U4598 ( .A1(n4208), .A2(n4364), .ZN(n4122) );
  AOI211_X1 U4599 ( .C1(n4046), .C2(n4120), .A(n4124), .B(n4122), .ZN(n4047)
         );
  NOR2_X1 U4600 ( .A1(n4152), .A2(n4314), .ZN(n4128) );
  AOI221_X1 U4601 ( .B1(n4123), .B2(n4127), .C1(n4047), .C2(n4127), .A(n4128), 
        .ZN(n4048) );
  NAND2_X1 U4602 ( .A1(n4315), .A2(n4328), .ZN(n4125) );
  NAND2_X1 U4603 ( .A1(n4048), .A2(n4125), .ZN(n4051) );
  NOR2_X1 U4604 ( .A1(n4330), .A2(n4049), .ZN(n4296) );
  NAND2_X1 U4605 ( .A1(n4212), .A2(n4301), .ZN(n4074) );
  INV_X1 U4606 ( .A(n4074), .ZN(n4050) );
  NOR2_X1 U4607 ( .A1(n4296), .A2(n4050), .ZN(n4131) );
  NAND2_X1 U4608 ( .A1(n4313), .A2(n4292), .ZN(n4075) );
  INV_X1 U4609 ( .A(n4075), .ZN(n4130) );
  NAND2_X1 U4610 ( .A1(n4214), .A2(n4228), .ZN(n4132) );
  AOI211_X1 U4611 ( .C1(n4051), .C2(n4131), .A(n4130), .B(n2572), .ZN(n4066)
         );
  INV_X1 U4612 ( .A(REG1_REG_31__SCAN_IN), .ZN(n4056) );
  NAND2_X1 U4613 ( .A1(n4052), .A2(REG2_REG_31__SCAN_IN), .ZN(n4055) );
  INV_X1 U4614 ( .A(REG0_REG_31__SCAN_IN), .ZN(n4053) );
  OR2_X1 U4615 ( .A1(n2513), .A2(n4053), .ZN(n4054) );
  OAI211_X1 U4616 ( .C1(n4061), .C2(n4056), .A(n4055), .B(n4054), .ZN(n5356)
         );
  NAND2_X1 U4617 ( .A1(n4064), .A2(DATAI_31_), .ZN(n5371) );
  OR2_X1 U4618 ( .A1(n5356), .A2(n5371), .ZN(n4063) );
  INV_X1 U4619 ( .A(REG1_REG_30__SCAN_IN), .ZN(n4060) );
  NAND2_X1 U4620 ( .A1(n4052), .A2(REG2_REG_30__SCAN_IN), .ZN(n4059) );
  INV_X1 U4621 ( .A(REG0_REG_30__SCAN_IN), .ZN(n4057) );
  OR2_X1 U4622 ( .A1(n2513), .A2(n4057), .ZN(n4058) );
  OAI211_X1 U4623 ( .C1(n4061), .C2(n4060), .A(n4059), .B(n4058), .ZN(n4197)
         );
  NAND2_X1 U4624 ( .A1(n4064), .A2(DATAI_30_), .ZN(n5358) );
  NAND2_X1 U4625 ( .A1(n4197), .A2(n5358), .ZN(n4062) );
  AND2_X1 U4626 ( .A1(n4063), .A2(n4062), .ZN(n4135) );
  INV_X1 U4627 ( .A(n4135), .ZN(n4096) );
  INV_X1 U4628 ( .A(n4242), .ZN(n4151) );
  AND2_X1 U4629 ( .A1(n4064), .A2(DATAI_29_), .ZN(n4229) );
  INV_X1 U4630 ( .A(n4229), .ZN(n4195) );
  NAND2_X1 U4631 ( .A1(n4151), .A2(n4195), .ZN(n4094) );
  INV_X1 U4632 ( .A(n4255), .ZN(n4222) );
  NAND2_X1 U4633 ( .A1(n4222), .A2(n4246), .ZN(n4098) );
  NAND2_X1 U4634 ( .A1(n4094), .A2(n4098), .ZN(n4133) );
  NAND2_X1 U4635 ( .A1(n4303), .A2(n4282), .ZN(n4257) );
  NAND2_X1 U4636 ( .A1(n4218), .A2(n4266), .ZN(n4085) );
  NAND2_X1 U4637 ( .A1(n4257), .A2(n4085), .ZN(n4065) );
  NOR4_X1 U4638 ( .A1(n4066), .A2(n4096), .A3(n4133), .A4(n4065), .ZN(n4072)
         );
  NAND2_X1 U4639 ( .A1(n5356), .A2(n5371), .ZN(n4070) );
  NAND2_X1 U4640 ( .A1(n4255), .A2(n4221), .ZN(n4192) );
  NAND2_X1 U4641 ( .A1(n4276), .A2(n4217), .ZN(n4191) );
  AOI21_X1 U4642 ( .B1(n4192), .B2(n4191), .A(n4133), .ZN(n4069) );
  NAND2_X1 U4643 ( .A1(n4242), .A2(n4229), .ZN(n4095) );
  INV_X1 U4644 ( .A(n4095), .ZN(n4068) );
  OR2_X1 U4645 ( .A1(n4197), .A2(n5358), .ZN(n4067) );
  NAND2_X1 U4646 ( .A1(n4070), .A2(n4067), .ZN(n4097) );
  NOR3_X1 U4647 ( .A1(n4069), .A2(n4068), .A3(n4097), .ZN(n4134) );
  AOI21_X1 U4648 ( .B1(n4070), .B2(n4096), .A(n4134), .ZN(n4071) );
  NOR2_X1 U4649 ( .A1(n4072), .A2(n4071), .ZN(n4144) );
  INV_X1 U4650 ( .A(n4073), .ZN(n4078) );
  NAND4_X1 U4651 ( .A1(n4078), .A2(n4299), .A3(n4440), .A4(n4077), .ZN(n4092)
         );
  OR4_X1 U4652 ( .A1(n3393), .A2(n4081), .A3(n4080), .A4(n4079), .ZN(n4091) );
  NAND4_X1 U4653 ( .A1(n4084), .A2(n4083), .A3(n5131), .A4(n4082), .ZN(n4090)
         );
  NAND2_X1 U4654 ( .A1(n4132), .A2(n4257), .ZN(n4274) );
  INV_X1 U4655 ( .A(n4274), .ZN(n4088) );
  AND2_X1 U4656 ( .A1(n4087), .A2(n4086), .ZN(n4385) );
  NAND4_X1 U4657 ( .A1(n4088), .A2(n5261), .A3(n4256), .A4(n4385), .ZN(n4089)
         );
  NOR4_X1 U4658 ( .A1(n4092), .A2(n4091), .A3(n4090), .A4(n4089), .ZN(n4105)
         );
  NOR2_X1 U4659 ( .A1(n2552), .A2(n4093), .ZN(n5212) );
  NAND2_X1 U4660 ( .A1(n4095), .A2(n4094), .ZN(n4225) );
  NOR4_X1 U4661 ( .A1(n5212), .A2(n4225), .A3(n4097), .A4(n4096), .ZN(n4103)
         );
  NAND2_X1 U4662 ( .A1(n4192), .A2(n4098), .ZN(n4237) );
  NOR4_X1 U4663 ( .A1(n4101), .A2(n4100), .A3(n4099), .A4(n4237), .ZN(n4102)
         );
  NAND4_X1 U4664 ( .A1(n4105), .A2(n4104), .A3(n4103), .A4(n4102), .ZN(n4112)
         );
  XNOR2_X1 U4665 ( .A(n4202), .B(n4428), .ZN(n4425) );
  INV_X1 U4666 ( .A(n4122), .ZN(n4107) );
  NAND2_X1 U4667 ( .A1(n4107), .A2(n4106), .ZN(n4367) );
  NAND2_X1 U4668 ( .A1(n4109), .A2(n4108), .ZN(n5114) );
  NAND2_X1 U4669 ( .A1(n4125), .A2(n4127), .ZN(n4327) );
  NOR4_X1 U4670 ( .A1(n4350), .A2(n4367), .A3(n5114), .A4(n4327), .ZN(n4110)
         );
  XOR2_X1 U4671 ( .A(n4152), .B(n4314), .Z(n4312) );
  NAND2_X1 U4672 ( .A1(n4110), .A2(n4312), .ZN(n4111) );
  XNOR2_X1 U4673 ( .A(n4419), .B(n4403), .ZN(n4408) );
  NOR4_X1 U4674 ( .A1(n4112), .A2(n4425), .A3(n4111), .A4(n4408), .ZN(n4113)
         );
  XNOR2_X1 U4675 ( .A(n4113), .B(n4138), .ZN(n4115) );
  INV_X1 U4676 ( .A(n3023), .ZN(n4922) );
  NAND3_X1 U4677 ( .A1(n4115), .A2(n4922), .A3(n4114), .ZN(n4116) );
  OAI21_X1 U4678 ( .B1(n4144), .B2(n4117), .A(n4116), .ZN(n4143) );
  OAI21_X1 U4679 ( .B1(n4439), .B2(n4121), .A(n4120), .ZN(n4368) );
  INV_X1 U4680 ( .A(n4125), .ZN(n4126) );
  INV_X1 U4681 ( .A(n4128), .ZN(n4129) );
  NAND2_X1 U4682 ( .A1(n4311), .A2(n4129), .ZN(n4298) );
  NOR2_X1 U4683 ( .A1(n4260), .A2(n4133), .ZN(n4137) );
  OAI21_X1 U4684 ( .B1(n5356), .B2(n5358), .A(n4134), .ZN(n4136) );
  OAI22_X1 U4685 ( .A1(n4137), .A2(n4136), .B1(n4135), .B2(n5371), .ZN(n4139)
         );
  XNOR2_X1 U4686 ( .A(n4139), .B(n4138), .ZN(n4141) );
  NOR2_X1 U4687 ( .A1(n4141), .A2(n4140), .ZN(n4142) );
  AOI211_X1 U4688 ( .C1(n4145), .C2(n4144), .A(n4143), .B(n4142), .ZN(n4150)
         );
  NOR2_X1 U4689 ( .A1(n4146), .A2(n5074), .ZN(n4148) );
  OAI21_X1 U4690 ( .B1(n4149), .B2(n4455), .A(B_REG_SCAN_IN), .ZN(n4147) );
  OAI22_X1 U4691 ( .A1(n4150), .A2(n4149), .B1(n4148), .B2(n4147), .ZN(U3239)
         );
  MUX2_X1 U4692 ( .A(DATAO_REG_31__SCAN_IN), .B(n5356), .S(n5082), .Z(U3581)
         );
  MUX2_X1 U4693 ( .A(DATAO_REG_30__SCAN_IN), .B(n4197), .S(n5082), .Z(U3580)
         );
  MUX2_X1 U4694 ( .A(DATAO_REG_29__SCAN_IN), .B(n4151), .S(n5082), .Z(U3579)
         );
  MUX2_X1 U4695 ( .A(DATAO_REG_28__SCAN_IN), .B(n4222), .S(U4043), .Z(U3578)
         );
  MUX2_X1 U4696 ( .A(DATAO_REG_27__SCAN_IN), .B(n4218), .S(U4043), .Z(U3577)
         );
  MUX2_X1 U4697 ( .A(DATAO_REG_26__SCAN_IN), .B(n4303), .S(U4043), .Z(U3576)
         );
  MUX2_X1 U4698 ( .A(DATAO_REG_25__SCAN_IN), .B(n4212), .S(n5082), .Z(U3575)
         );
  MUX2_X1 U4699 ( .A(DATAO_REG_24__SCAN_IN), .B(n4152), .S(n5082), .Z(U3574)
         );
  MUX2_X1 U4700 ( .A(DATAO_REG_23__SCAN_IN), .B(n4354), .S(n5082), .Z(U3573)
         );
  MUX2_X1 U4701 ( .A(DATAO_REG_22__SCAN_IN), .B(n4371), .S(n5082), .Z(U3572)
         );
  MUX2_X1 U4702 ( .A(DATAO_REG_21__SCAN_IN), .B(n4208), .S(n5082), .Z(U3571)
         );
  MUX2_X1 U4703 ( .A(DATAO_REG_20__SCAN_IN), .B(n4206), .S(n5082), .Z(U3570)
         );
  MUX2_X1 U4704 ( .A(DATAO_REG_19__SCAN_IN), .B(n4419), .S(n5082), .Z(U3569)
         );
  MUX2_X1 U4705 ( .A(DATAO_REG_18__SCAN_IN), .B(n4202), .S(n5082), .Z(U3568)
         );
  MUX2_X1 U4706 ( .A(DATAO_REG_17__SCAN_IN), .B(n4201), .S(n5082), .Z(U3567)
         );
  MUX2_X1 U4707 ( .A(DATAO_REG_16__SCAN_IN), .B(n5308), .S(n5082), .Z(U3566)
         );
  MUX2_X1 U4708 ( .A(DATAO_REG_15__SCAN_IN), .B(n4153), .S(n5082), .Z(U3565)
         );
  MUX2_X1 U4709 ( .A(DATAO_REG_14__SCAN_IN), .B(n4154), .S(n5082), .Z(U3564)
         );
  MUX2_X1 U4710 ( .A(DATAO_REG_13__SCAN_IN), .B(n4155), .S(n5082), .Z(U3563)
         );
  MUX2_X1 U4711 ( .A(DATAO_REG_12__SCAN_IN), .B(n4156), .S(n5082), .Z(U3562)
         );
  MUX2_X1 U4712 ( .A(DATAO_REG_11__SCAN_IN), .B(n4157), .S(n5082), .Z(U3561)
         );
  MUX2_X1 U4713 ( .A(DATAO_REG_10__SCAN_IN), .B(n4158), .S(n5082), .Z(U3560)
         );
  MUX2_X1 U4714 ( .A(DATAO_REG_9__SCAN_IN), .B(n4159), .S(n5082), .Z(U3559) );
  MUX2_X1 U4715 ( .A(DATAO_REG_8__SCAN_IN), .B(n4160), .S(n5082), .Z(U3558) );
  MUX2_X1 U4716 ( .A(DATAO_REG_7__SCAN_IN), .B(n4161), .S(n5082), .Z(U3557) );
  MUX2_X1 U4717 ( .A(DATAO_REG_6__SCAN_IN), .B(n5181), .S(n5082), .Z(U3556) );
  MUX2_X1 U4718 ( .A(DATAO_REG_5__SCAN_IN), .B(n4162), .S(n5082), .Z(U3555) );
  MUX2_X1 U4719 ( .A(DATAO_REG_4__SCAN_IN), .B(n5135), .S(n5082), .Z(U3554) );
  MUX2_X1 U4720 ( .A(DATAO_REG_3__SCAN_IN), .B(n4163), .S(n5082), .Z(U3553) );
  MUX2_X1 U4721 ( .A(DATAO_REG_2__SCAN_IN), .B(n4164), .S(n5082), .Z(U3552) );
  MUX2_X1 U4722 ( .A(DATAO_REG_1__SCAN_IN), .B(n5103), .S(n5082), .Z(U3551) );
  MUX2_X1 U4723 ( .A(DATAO_REG_0__SCAN_IN), .B(n4165), .S(n5082), .Z(U3550) );
  AOI21_X1 U4724 ( .B1(n4168), .B2(n4167), .A(n4166), .ZN(n4176) );
  NOR2_X1 U4725 ( .A1(STATE_REG_SCAN_IN), .A2(n4169), .ZN(n5307) );
  AOI21_X1 U4726 ( .B1(n5087), .B2(ADDR_REG_15__SCAN_IN), .A(n5307), .ZN(n4170) );
  OAI21_X1 U4727 ( .B1(n4171), .B2(n5069), .A(n4170), .ZN(n4175) );
  AOI211_X1 U4728 ( .C1(n2542), .C2(n4173), .A(n4172), .B(n5091), .ZN(n4174)
         );
  AOI211_X1 U4729 ( .C1(n5065), .C2(n4176), .A(n4175), .B(n4174), .ZN(n4177)
         );
  INV_X1 U4730 ( .A(n4177), .ZN(U3255) );
  OAI21_X1 U4731 ( .B1(n4179), .B2(n5329), .A(n4178), .ZN(n4189) );
  OAI21_X1 U4732 ( .B1(n4182), .B2(n4181), .A(n4180), .ZN(n4183) );
  NAND2_X1 U4733 ( .A1(n4183), .A2(n5060), .ZN(n4186) );
  AOI21_X1 U4734 ( .B1(n5087), .B2(ADDR_REG_16__SCAN_IN), .A(n4184), .ZN(n4185) );
  OAI211_X1 U4735 ( .C1(n5069), .C2(n4187), .A(n4186), .B(n4185), .ZN(n4188)
         );
  AOI21_X1 U4736 ( .B1(n5065), .B2(n4189), .A(n4188), .ZN(n4190) );
  INV_X1 U4737 ( .A(n4190), .ZN(U3256) );
  INV_X1 U4738 ( .A(n4237), .ZN(n4241) );
  NAND2_X1 U4739 ( .A1(n4240), .A2(n4241), .ZN(n4239) );
  NAND2_X1 U4740 ( .A1(n4239), .A2(n4192), .ZN(n4193) );
  XNOR2_X1 U4741 ( .A(n4193), .B(n4225), .ZN(n4199) );
  NAND2_X1 U4742 ( .A1(n4954), .A2(B_REG_SCAN_IN), .ZN(n4194) );
  AND2_X1 U4743 ( .A1(n5136), .A2(n4194), .ZN(n5355) );
  OAI22_X1 U4744 ( .A1(n4255), .A2(n5246), .B1(n5266), .B2(n4195), .ZN(n4196)
         );
  AOI21_X1 U4745 ( .B1(n5355), .B2(n4197), .A(n4196), .ZN(n4198) );
  OAI21_X1 U4746 ( .B1(n4199), .B2(n5138), .A(n4198), .ZN(n4458) );
  INV_X1 U4747 ( .A(n4458), .ZN(n4236) );
  NAND2_X1 U4748 ( .A1(n4424), .A2(n4203), .ZN(n4409) );
  NAND2_X1 U4749 ( .A1(n4409), .A2(n4408), .ZN(n4407) );
  NAND2_X1 U4750 ( .A1(n4342), .A2(n4350), .ZN(n4210) );
  NAND2_X1 U4751 ( .A1(n4371), .A2(n4345), .ZN(n4209) );
  NAND2_X1 U4752 ( .A1(n4210), .A2(n4209), .ZN(n4325) );
  NAND2_X1 U4753 ( .A1(n4354), .A2(n4328), .ZN(n4211) );
  NAND2_X1 U4754 ( .A1(n4212), .A2(n4292), .ZN(n4213) );
  NOR2_X1 U4755 ( .A1(n4214), .A2(n4282), .ZN(n4216) );
  NAND2_X1 U4756 ( .A1(n4214), .A2(n4282), .ZN(n4215) );
  NOR2_X1 U4757 ( .A1(n4218), .A2(n4217), .ZN(n4220) );
  NAND2_X1 U4758 ( .A1(n4218), .A2(n4217), .ZN(n4219) );
  NAND2_X1 U4759 ( .A1(n4224), .A2(n4223), .ZN(n4227) );
  XNOR2_X1 U4760 ( .A(n4227), .B(n4226), .ZN(n4456) );
  NAND2_X1 U4761 ( .A1(n4456), .A2(n4437), .ZN(n4235) );
  AOI21_X1 U4762 ( .B1(n2520), .B2(n4229), .A(n5333), .ZN(n4230) );
  AND2_X1 U4763 ( .A1(n4230), .A2(n5370), .ZN(n4457) );
  INV_X1 U4764 ( .A(REG2_REG_29__SCAN_IN), .ZN(n4232) );
  OAI22_X1 U4765 ( .A1(n5226), .A2(n4232), .B1(n4231), .B2(n5231), .ZN(n4233)
         );
  AOI21_X1 U4766 ( .B1(n4457), .B2(n4247), .A(n4233), .ZN(n4234) );
  OAI211_X1 U4767 ( .C1(n4236), .C2(n5374), .A(n4235), .B(n4234), .ZN(U3354)
         );
  XNOR2_X1 U4768 ( .A(n4238), .B(n4237), .ZN(n4468) );
  OAI21_X1 U4769 ( .B1(n4241), .B2(n4240), .A(n4239), .ZN(n4245) );
  NOR2_X1 U4770 ( .A1(n4242), .A2(n5244), .ZN(n4244) );
  OAI22_X1 U4771 ( .A1(n4276), .A2(n5246), .B1(n5266), .B2(n4246), .ZN(n4243)
         );
  AOI211_X1 U4772 ( .C1(n4245), .C2(n5268), .A(n4244), .B(n4243), .ZN(n4467)
         );
  INV_X1 U4773 ( .A(n4467), .ZN(n4252) );
  OAI211_X1 U4774 ( .C1(n4264), .C2(n4246), .A(n5377), .B(n2520), .ZN(n4466)
         );
  INV_X1 U4775 ( .A(n4247), .ZN(n4429) );
  INV_X1 U4776 ( .A(n4248), .ZN(n4249) );
  INV_X1 U4777 ( .A(n5231), .ZN(n5276) );
  AOI22_X1 U4778 ( .A1(n5374), .A2(REG2_REG_28__SCAN_IN), .B1(n4249), .B2(
        n5276), .ZN(n4250) );
  OAI21_X1 U4779 ( .B1(n4466), .B2(n4429), .A(n4250), .ZN(n4251) );
  AOI21_X1 U4780 ( .B1(n4252), .B2(n5226), .A(n4251), .ZN(n4253) );
  OAI21_X1 U4781 ( .B1(n4468), .B2(n4399), .A(n4253), .ZN(U3262) );
  XNOR2_X1 U4782 ( .A(n4254), .B(n4256), .ZN(n4471) );
  OAI22_X1 U4783 ( .A1(n4255), .A2(n5244), .B1(n5266), .B2(n4266), .ZN(n4263)
         );
  AOI21_X1 U4784 ( .B1(n4258), .B2(n4257), .A(n4256), .ZN(n4259) );
  INV_X1 U4785 ( .A(n4259), .ZN(n4261) );
  AOI21_X1 U4786 ( .B1(n4261), .B2(n4260), .A(n5138), .ZN(n4262) );
  AOI211_X1 U4787 ( .C1(n5180), .C2(n4303), .A(n4263), .B(n4262), .ZN(n4470)
         );
  INV_X1 U4788 ( .A(n2510), .ZN(n4271) );
  INV_X1 U4789 ( .A(n4264), .ZN(n4265) );
  OAI211_X1 U4790 ( .C1(n4280), .C2(n4266), .A(n4265), .B(n5377), .ZN(n4469)
         );
  INV_X1 U4791 ( .A(n4267), .ZN(n4268) );
  AOI22_X1 U4792 ( .A1(n5374), .A2(REG2_REG_27__SCAN_IN), .B1(n4268), .B2(
        n5276), .ZN(n4269) );
  OAI21_X1 U4793 ( .B1(n4469), .B2(n4429), .A(n4269), .ZN(n4270) );
  AOI21_X1 U4794 ( .B1(n4271), .B2(n5226), .A(n4270), .ZN(n4272) );
  OAI21_X1 U4795 ( .B1(n4471), .B2(n4399), .A(n4272), .ZN(U3263) );
  XNOR2_X1 U4796 ( .A(n4273), .B(n4274), .ZN(n4474) );
  XNOR2_X1 U4797 ( .A(n4275), .B(n4274), .ZN(n4279) );
  NOR2_X1 U4798 ( .A1(n4313), .A2(n5246), .ZN(n4278) );
  OAI22_X1 U4799 ( .A1(n4276), .A2(n5244), .B1(n5266), .B2(n4282), .ZN(n4277)
         );
  AOI211_X1 U4800 ( .C1(n4279), .C2(n5268), .A(n4278), .B(n4277), .ZN(n4473)
         );
  INV_X1 U4801 ( .A(n4473), .ZN(n4287) );
  INV_X1 U4802 ( .A(n4280), .ZN(n4281) );
  OAI211_X1 U4803 ( .C1(n2533), .C2(n4282), .A(n4281), .B(n5377), .ZN(n4472)
         );
  INV_X1 U4804 ( .A(n4283), .ZN(n4284) );
  AOI22_X1 U4805 ( .A1(n5374), .A2(REG2_REG_26__SCAN_IN), .B1(n4284), .B2(
        n5276), .ZN(n4285) );
  OAI21_X1 U4806 ( .B1(n4472), .B2(n4429), .A(n4285), .ZN(n4286) );
  AOI21_X1 U4807 ( .B1(n4287), .B2(n5226), .A(n4286), .ZN(n4288) );
  OAI21_X1 U4808 ( .B1(n4474), .B2(n4399), .A(n4288), .ZN(U3264) );
  INV_X1 U4809 ( .A(n4289), .ZN(n4291) );
  INV_X1 U4810 ( .A(n4299), .ZN(n4290) );
  OAI21_X1 U4811 ( .B1(n4291), .B2(n4290), .A(n2749), .ZN(n4478) );
  AOI21_X1 U4812 ( .B1(n4292), .B2(n4308), .A(n2533), .ZN(n4476) );
  OAI22_X1 U4813 ( .A1(n5226), .A2(n4294), .B1(n4293), .B2(n5231), .ZN(n4295)
         );
  AOI21_X1 U4814 ( .B1(n4476), .B2(n5372), .A(n4295), .ZN(n4307) );
  INV_X1 U4815 ( .A(n4296), .ZN(n4297) );
  NAND2_X1 U4816 ( .A1(n4298), .A2(n4297), .ZN(n4300) );
  XNOR2_X1 U4817 ( .A(n4300), .B(n4299), .ZN(n4305) );
  OAI22_X1 U4818 ( .A1(n4330), .A2(n5246), .B1(n5266), .B2(n4301), .ZN(n4302)
         );
  AOI21_X1 U4819 ( .B1(n5136), .B2(n4303), .A(n4302), .ZN(n4304) );
  OAI21_X1 U4820 ( .B1(n4305), .B2(n5138), .A(n4304), .ZN(n4475) );
  NAND2_X1 U4821 ( .A1(n4475), .A2(n4450), .ZN(n4306) );
  OAI211_X1 U4822 ( .C1(n4478), .C2(n4399), .A(n4307), .B(n4306), .ZN(U3265)
         );
  OAI211_X1 U4823 ( .C1(n4335), .C2(n4314), .A(n5377), .B(n4308), .ZN(n4479)
         );
  XOR2_X1 U4824 ( .A(n4312), .B(n4309), .Z(n4481) );
  INV_X1 U4825 ( .A(n4481), .ZN(n4310) );
  NAND2_X1 U4826 ( .A1(n4310), .A2(n5177), .ZN(n4319) );
  XOR2_X1 U4827 ( .A(n4312), .B(n4311), .Z(n4318) );
  NOR2_X1 U4828 ( .A1(n4313), .A2(n5244), .ZN(n4317) );
  OAI22_X1 U4829 ( .A1(n4315), .A2(n5246), .B1(n5266), .B2(n4314), .ZN(n4316)
         );
  AOI211_X1 U4830 ( .C1(n4318), .C2(n5268), .A(n4317), .B(n4316), .ZN(n4480)
         );
  OAI211_X1 U4831 ( .C1(n4479), .C2(n2846), .A(n4319), .B(n4480), .ZN(n4323)
         );
  OAI22_X1 U4832 ( .A1(n5226), .A2(n4321), .B1(n4320), .B2(n5231), .ZN(n4322)
         );
  AOI21_X1 U4833 ( .B1(n4323), .B2(n4450), .A(n4322), .ZN(n4324) );
  INV_X1 U4834 ( .A(n4324), .ZN(U3266) );
  XNOR2_X1 U4835 ( .A(n4325), .B(n4327), .ZN(n4484) );
  XOR2_X1 U4836 ( .A(n4327), .B(n4326), .Z(n4332) );
  AOI22_X1 U4837 ( .A1(n4371), .A2(n5180), .B1(n5365), .B2(n4328), .ZN(n4329)
         );
  OAI21_X1 U4838 ( .B1(n4330), .B2(n5244), .A(n4329), .ZN(n4331) );
  AOI21_X1 U4839 ( .B1(n4332), .B2(n5268), .A(n4331), .ZN(n4483) );
  INV_X1 U4840 ( .A(n4483), .ZN(n4340) );
  OAI21_X1 U4841 ( .B1(n4343), .B2(n4333), .A(n5377), .ZN(n4334) );
  OR2_X1 U4842 ( .A1(n4335), .A2(n4334), .ZN(n4482) );
  INV_X1 U4843 ( .A(n4336), .ZN(n4337) );
  AOI22_X1 U4844 ( .A1(n5374), .A2(REG2_REG_23__SCAN_IN), .B1(n4337), .B2(
        n5276), .ZN(n4338) );
  OAI21_X1 U4845 ( .B1(n4482), .B2(n4429), .A(n4338), .ZN(n4339) );
  AOI21_X1 U4846 ( .B1(n4340), .B2(n5226), .A(n4339), .ZN(n4341) );
  OAI21_X1 U4847 ( .B1(n4484), .B2(n4399), .A(n4341), .ZN(U3267) );
  XNOR2_X1 U4848 ( .A(n4342), .B(n4350), .ZN(n4488) );
  INV_X1 U4849 ( .A(n4360), .ZN(n4344) );
  AOI21_X1 U4850 ( .B1(n4345), .B2(n4344), .A(n4343), .ZN(n4486) );
  INV_X1 U4851 ( .A(REG2_REG_22__SCAN_IN), .ZN(n4347) );
  OAI22_X1 U4852 ( .A1(n5226), .A2(n4347), .B1(n4346), .B2(n5231), .ZN(n4348)
         );
  AOI21_X1 U4853 ( .B1(n4486), .B2(n5372), .A(n4348), .ZN(n4358) );
  XOR2_X1 U4854 ( .A(n4350), .B(n4349), .Z(n4356) );
  OAI22_X1 U4855 ( .A1(n4352), .A2(n5246), .B1(n5266), .B2(n4351), .ZN(n4353)
         );
  AOI21_X1 U4856 ( .B1(n5136), .B2(n4354), .A(n4353), .ZN(n4355) );
  OAI21_X1 U4857 ( .B1(n4356), .B2(n5138), .A(n4355), .ZN(n4485) );
  NAND2_X1 U4858 ( .A1(n4485), .A2(n5226), .ZN(n4357) );
  OAI211_X1 U4859 ( .C1(n4488), .C2(n4399), .A(n4358), .B(n4357), .ZN(U3268)
         );
  XNOR2_X1 U4860 ( .A(n4359), .B(n4367), .ZN(n4492) );
  AOI21_X1 U4861 ( .B1(n4361), .B2(n4391), .A(n4360), .ZN(n4489) );
  INV_X1 U4862 ( .A(REG2_REG_21__SCAN_IN), .ZN(n4363) );
  OAI22_X1 U4863 ( .A1(n5226), .A2(n4363), .B1(n4362), .B2(n5231), .ZN(n4373)
         );
  OAI22_X1 U4864 ( .A1(n4365), .A2(n5246), .B1(n5266), .B2(n4364), .ZN(n4370)
         );
  AOI211_X1 U4865 ( .C1(n4368), .C2(n4367), .A(n5138), .B(n4366), .ZN(n4369)
         );
  AOI211_X1 U4866 ( .C1(n5136), .C2(n4371), .A(n4370), .B(n4369), .ZN(n4491)
         );
  NOR2_X1 U4867 ( .A1(n4491), .A2(n5374), .ZN(n4372) );
  AOI211_X1 U4868 ( .C1(n4489), .C2(n5372), .A(n4373), .B(n4372), .ZN(n4374)
         );
  OAI21_X1 U4869 ( .B1(n4492), .B2(n4399), .A(n4374), .ZN(U3269) );
  XNOR2_X1 U4870 ( .A(n4375), .B(n4385), .ZN(n4495) );
  INV_X1 U4871 ( .A(n4439), .ZN(n4379) );
  INV_X1 U4872 ( .A(n4376), .ZN(n4377) );
  AOI21_X1 U4873 ( .B1(n4379), .B2(n4378), .A(n4377), .ZN(n4417) );
  NAND2_X1 U4874 ( .A1(n4417), .A2(n4380), .ZN(n4401) );
  INV_X1 U4875 ( .A(n4381), .ZN(n4382) );
  AOI21_X1 U4876 ( .B1(n4401), .B2(n4383), .A(n4382), .ZN(n4384) );
  XOR2_X1 U4877 ( .A(n4385), .B(n4384), .Z(n4389) );
  NOR2_X1 U4878 ( .A1(n4386), .A2(n5266), .ZN(n4388) );
  AOI211_X1 U4879 ( .C1(n4389), .C2(n5268), .A(n4388), .B(n4387), .ZN(n4494)
         );
  INV_X1 U4880 ( .A(n4494), .ZN(n4397) );
  AOI21_X1 U4881 ( .B1(n4412), .B2(n4390), .A(n5333), .ZN(n4392) );
  NAND2_X1 U4882 ( .A1(n4392), .A2(n4391), .ZN(n4493) );
  INV_X1 U4883 ( .A(n4393), .ZN(n4394) );
  AOI22_X1 U4884 ( .A1(n5374), .A2(REG2_REG_20__SCAN_IN), .B1(n4394), .B2(
        n5276), .ZN(n4395) );
  OAI21_X1 U4885 ( .B1(n4493), .B2(n4429), .A(n4395), .ZN(n4396) );
  AOI21_X1 U4886 ( .B1(n4397), .B2(n4450), .A(n4396), .ZN(n4398) );
  OAI21_X1 U4887 ( .B1(n4495), .B2(n4399), .A(n4398), .ZN(U3270) );
  NAND2_X1 U4888 ( .A1(n4401), .A2(n4400), .ZN(n4402) );
  XNOR2_X1 U4889 ( .A(n4402), .B(n4408), .ZN(n4406) );
  NOR2_X1 U4890 ( .A1(n4403), .A2(n5266), .ZN(n4405) );
  AOI211_X1 U4891 ( .C1(n4406), .C2(n5268), .A(n4405), .B(n4404), .ZN(n4497)
         );
  OAI21_X1 U4892 ( .B1(n4409), .B2(n4408), .A(n4407), .ZN(n4496) );
  NAND2_X1 U4893 ( .A1(n4427), .A2(n4410), .ZN(n4411) );
  NAND2_X1 U4894 ( .A1(n4412), .A2(n4411), .ZN(n4499) );
  NOR2_X1 U4895 ( .A1(n4499), .A2(n4454), .ZN(n4415) );
  OAI22_X1 U4896 ( .A1(n4450), .A2(n2922), .B1(n4413), .B2(n5231), .ZN(n4414)
         );
  AOI211_X1 U4897 ( .C1(n4496), .C2(n4437), .A(n4415), .B(n4414), .ZN(n4416)
         );
  OAI21_X1 U4898 ( .B1(n5374), .B2(n4497), .A(n4416), .ZN(U3271) );
  XNOR2_X1 U4899 ( .A(n4417), .B(n4425), .ZN(n4423) );
  NOR2_X1 U4900 ( .A1(n4428), .A2(n5266), .ZN(n4422) );
  OR2_X1 U4901 ( .A1(n4418), .A2(n5246), .ZN(n4421) );
  NAND2_X1 U4902 ( .A1(n4419), .A2(n5136), .ZN(n4420) );
  NAND2_X1 U4903 ( .A1(n4421), .A2(n4420), .ZN(n5347) );
  AOI211_X1 U4904 ( .C1(n4423), .C2(n5268), .A(n4422), .B(n5347), .ZN(n4502)
         );
  OAI21_X1 U4905 ( .B1(n4426), .B2(n4425), .A(n4424), .ZN(n4500) );
  OAI211_X1 U4906 ( .C1(n4434), .C2(n4428), .A(n4427), .B(n5377), .ZN(n4501)
         );
  NOR2_X1 U4907 ( .A1(n4501), .A2(n4429), .ZN(n4432) );
  INV_X1 U4908 ( .A(REG2_REG_18__SCAN_IN), .ZN(n4430) );
  OAI22_X1 U4909 ( .A1(n4450), .A2(n4430), .B1(n5353), .B2(n5231), .ZN(n4431)
         );
  AOI211_X1 U4910 ( .C1(n4500), .C2(n4437), .A(n4432), .B(n4431), .ZN(n4433)
         );
  OAI21_X1 U4911 ( .B1(n5374), .B2(n4502), .A(n4433), .ZN(U3272) );
  AND2_X1 U4912 ( .A1(n2519), .A2(n4442), .ZN(n4435) );
  OR2_X1 U4913 ( .A1(n4435), .A2(n4434), .ZN(n5332) );
  XNOR2_X1 U4914 ( .A(n4436), .B(n4440), .ZN(n5336) );
  NAND2_X1 U4915 ( .A1(n5336), .A2(n4437), .ZN(n4453) );
  NOR2_X1 U4916 ( .A1(n4439), .A2(n4438), .ZN(n4441) );
  XNOR2_X1 U4917 ( .A(n4441), .B(n4440), .ZN(n4446) );
  AOI22_X1 U4918 ( .A1(n5308), .A2(n5180), .B1(n5365), .B2(n4442), .ZN(n4443)
         );
  OAI21_X1 U4919 ( .B1(n4444), .B2(n5244), .A(n4443), .ZN(n4445) );
  AOI21_X1 U4920 ( .B1(n4446), .B2(n5268), .A(n4445), .ZN(n5331) );
  OAI21_X1 U4921 ( .B1(n4447), .B2(n5231), .A(n5331), .ZN(n4451) );
  INV_X1 U4922 ( .A(REG2_REG_17__SCAN_IN), .ZN(n4448) );
  NOR2_X1 U4923 ( .A1(n4450), .A2(n4448), .ZN(n4449) );
  AOI21_X1 U4924 ( .B1(n4451), .B2(n4450), .A(n4449), .ZN(n4452) );
  OAI211_X1 U4925 ( .C1(n5332), .C2(n4454), .A(n4453), .B(n4452), .ZN(U3273)
         );
  OR2_X1 U4926 ( .A1(n5112), .A2(n4455), .ZN(n5122) );
  NAND2_X1 U4927 ( .A1(n4456), .A2(n5335), .ZN(n4460) );
  NOR2_X1 U4928 ( .A1(n4458), .A2(n4457), .ZN(n4459) );
  NAND2_X1 U4929 ( .A1(n4460), .A2(n4459), .ZN(n4506) );
  NAND4_X1 U4930 ( .A1(n4464), .A2(n4463), .A3(n4462), .A4(n4461), .ZN(n4505)
         );
  MUX2_X1 U4931 ( .A(REG1_REG_29__SCAN_IN), .B(n4506), .S(n5363), .Z(U3547) );
  OAI211_X1 U4932 ( .C1(n4468), .C2(n5296), .A(n4467), .B(n4466), .ZN(n4507)
         );
  MUX2_X1 U4933 ( .A(REG1_REG_28__SCAN_IN), .B(n4507), .S(n5363), .Z(U3546) );
  OAI211_X1 U4934 ( .C1(n4471), .C2(n5296), .A(n2510), .B(n4469), .ZN(n4508)
         );
  MUX2_X1 U4935 ( .A(REG1_REG_27__SCAN_IN), .B(n4508), .S(n5363), .Z(U3545) );
  OAI211_X1 U4936 ( .C1(n4474), .C2(n5296), .A(n4473), .B(n4472), .ZN(n4509)
         );
  MUX2_X1 U4937 ( .A(REG1_REG_26__SCAN_IN), .B(n4509), .S(n5363), .Z(U3544) );
  AOI21_X1 U4938 ( .B1(n5377), .B2(n4476), .A(n4475), .ZN(n4477) );
  OAI21_X1 U4939 ( .B1(n4478), .B2(n5296), .A(n4477), .ZN(n4510) );
  MUX2_X1 U4940 ( .A(REG1_REG_25__SCAN_IN), .B(n4510), .S(n5363), .Z(U3543) );
  OAI211_X1 U4941 ( .C1(n4481), .C2(n5296), .A(n4480), .B(n4479), .ZN(n4511)
         );
  MUX2_X1 U4942 ( .A(REG1_REG_24__SCAN_IN), .B(n4511), .S(n5363), .Z(U3542) );
  OAI211_X1 U4943 ( .C1(n4484), .C2(n5296), .A(n4483), .B(n4482), .ZN(n4512)
         );
  MUX2_X1 U4944 ( .A(REG1_REG_23__SCAN_IN), .B(n4512), .S(n5363), .Z(U3541) );
  AOI21_X1 U4945 ( .B1(n5377), .B2(n4486), .A(n4485), .ZN(n4487) );
  OAI21_X1 U4946 ( .B1(n4488), .B2(n5296), .A(n4487), .ZN(n4513) );
  MUX2_X1 U4947 ( .A(REG1_REG_22__SCAN_IN), .B(n4513), .S(n5363), .Z(U3540) );
  NAND2_X1 U4948 ( .A1(n4489), .A2(n5377), .ZN(n4490) );
  OAI211_X1 U4949 ( .C1(n4492), .C2(n5296), .A(n4491), .B(n4490), .ZN(n4514)
         );
  MUX2_X1 U4950 ( .A(REG1_REG_21__SCAN_IN), .B(n4514), .S(n5363), .Z(U3539) );
  OAI211_X1 U4951 ( .C1(n4495), .C2(n5296), .A(n4494), .B(n4493), .ZN(n4515)
         );
  MUX2_X1 U4952 ( .A(REG1_REG_20__SCAN_IN), .B(n4515), .S(n5363), .Z(U3538) );
  NAND2_X1 U4953 ( .A1(n4496), .A2(n5335), .ZN(n4498) );
  OAI211_X1 U4954 ( .C1(n5333), .C2(n4499), .A(n4498), .B(n4497), .ZN(n4516)
         );
  MUX2_X1 U4955 ( .A(REG1_REG_19__SCAN_IN), .B(n4516), .S(n5363), .Z(U3537) );
  INV_X1 U4956 ( .A(n4500), .ZN(n4503) );
  OAI211_X1 U4957 ( .C1(n4503), .C2(n5296), .A(n4502), .B(n4501), .ZN(n4517)
         );
  MUX2_X1 U4958 ( .A(REG1_REG_18__SCAN_IN), .B(n4517), .S(n5363), .Z(U3536) );
  MUX2_X1 U4959 ( .A(REG0_REG_29__SCAN_IN), .B(n4506), .S(n2512), .Z(U3515) );
  MUX2_X1 U4960 ( .A(REG0_REG_28__SCAN_IN), .B(n4507), .S(n2512), .Z(U3514) );
  MUX2_X1 U4961 ( .A(REG0_REG_27__SCAN_IN), .B(n4508), .S(n2512), .Z(U3513) );
  MUX2_X1 U4962 ( .A(REG0_REG_26__SCAN_IN), .B(n4509), .S(n2512), .Z(U3512) );
  MUX2_X1 U4963 ( .A(REG0_REG_25__SCAN_IN), .B(n4510), .S(n2512), .Z(U3511) );
  MUX2_X1 U4964 ( .A(REG0_REG_24__SCAN_IN), .B(n4511), .S(n2512), .Z(U3510) );
  MUX2_X1 U4965 ( .A(REG0_REG_23__SCAN_IN), .B(n4512), .S(n2512), .Z(U3509) );
  MUX2_X1 U4966 ( .A(REG0_REG_22__SCAN_IN), .B(n4513), .S(n2512), .Z(U3508) );
  MUX2_X1 U4967 ( .A(REG0_REG_21__SCAN_IN), .B(n4514), .S(n2512), .Z(U3507) );
  MUX2_X1 U4968 ( .A(REG0_REG_20__SCAN_IN), .B(n4515), .S(n2512), .Z(U3506) );
  MUX2_X1 U4969 ( .A(REG0_REG_19__SCAN_IN), .B(n4516), .S(n2512), .Z(U3505) );
  MUX2_X1 U4970 ( .A(REG0_REG_18__SCAN_IN), .B(n4517), .S(n2512), .Z(U3503) );
  AOI22_X1 U4971 ( .A1(n4519), .A2(n5335), .B1(n5377), .B2(n4518), .ZN(n4521)
         );
  NAND2_X1 U4972 ( .A1(n4521), .A2(n4520), .ZN(n5160) );
  MUX2_X1 U4973 ( .A(REG0_REG_5__SCAN_IN), .B(n5160), .S(n2512), .Z(n4915) );
  XOR2_X1 U4974 ( .A(DATAI_30_), .B(keyinput_129), .Z(n4525) );
  XOR2_X1 U4975 ( .A(DATAI_31_), .B(keyinput_128), .Z(n4524) );
  XOR2_X1 U4976 ( .A(DATAI_28_), .B(keyinput_131), .Z(n4523) );
  XOR2_X1 U4977 ( .A(DATAI_29_), .B(keyinput_130), .Z(n4522) );
  AOI211_X1 U4978 ( .C1(n4525), .C2(n4524), .A(n4523), .B(n4522), .ZN(n4528)
         );
  XOR2_X1 U4979 ( .A(DATAI_27_), .B(keyinput_132), .Z(n4527) );
  XNOR2_X1 U4980 ( .A(DATAI_26_), .B(keyinput_133), .ZN(n4526) );
  OAI21_X1 U4981 ( .B1(n4528), .B2(n4527), .A(n4526), .ZN(n4531) );
  XNOR2_X1 U4982 ( .A(DATAI_25_), .B(keyinput_134), .ZN(n4530) );
  XNOR2_X1 U4983 ( .A(DATAI_24_), .B(keyinput_135), .ZN(n4529) );
  AOI21_X1 U4984 ( .B1(n4531), .B2(n4530), .A(n4529), .ZN(n4534) );
  XOR2_X1 U4985 ( .A(DATAI_23_), .B(keyinput_136), .Z(n4533) );
  XNOR2_X1 U4986 ( .A(DATAI_22_), .B(keyinput_137), .ZN(n4532) );
  OAI21_X1 U4987 ( .B1(n4534), .B2(n4533), .A(n4532), .ZN(n4537) );
  XOR2_X1 U4988 ( .A(DATAI_21_), .B(keyinput_138), .Z(n4536) );
  XNOR2_X1 U4989 ( .A(DATAI_20_), .B(keyinput_139), .ZN(n4535) );
  AOI21_X1 U4990 ( .B1(n4537), .B2(n4536), .A(n4535), .ZN(n4540) );
  XNOR2_X1 U4991 ( .A(DATAI_18_), .B(keyinput_141), .ZN(n4539) );
  XNOR2_X1 U4992 ( .A(DATAI_19_), .B(keyinput_140), .ZN(n4538) );
  NOR3_X1 U4993 ( .A1(n4540), .A2(n4539), .A3(n4538), .ZN(n4550) );
  XNOR2_X1 U4994 ( .A(DATAI_17_), .B(keyinput_142), .ZN(n4549) );
  XOR2_X1 U4995 ( .A(DATAI_13_), .B(keyinput_146), .Z(n4544) );
  XNOR2_X1 U4996 ( .A(DATAI_15_), .B(keyinput_144), .ZN(n4543) );
  XNOR2_X1 U4997 ( .A(DATAI_11_), .B(keyinput_148), .ZN(n4542) );
  XNOR2_X1 U4998 ( .A(DATAI_12_), .B(keyinput_147), .ZN(n4541) );
  NAND4_X1 U4999 ( .A1(n4544), .A2(n4543), .A3(n4542), .A4(n4541), .ZN(n4547)
         );
  XNOR2_X1 U5000 ( .A(DATAI_16_), .B(keyinput_143), .ZN(n4546) );
  XNOR2_X1 U5001 ( .A(DATAI_14_), .B(keyinput_145), .ZN(n4545) );
  NOR3_X1 U5002 ( .A1(n4547), .A2(n4546), .A3(n4545), .ZN(n4548) );
  OAI21_X1 U5003 ( .B1(n4550), .B2(n4549), .A(n4548), .ZN(n4556) );
  XNOR2_X1 U5004 ( .A(DATAI_10_), .B(keyinput_149), .ZN(n4555) );
  XOR2_X1 U5005 ( .A(DATAI_9_), .B(keyinput_150), .Z(n4553) );
  XOR2_X1 U5006 ( .A(DATAI_7_), .B(keyinput_152), .Z(n4552) );
  XNOR2_X1 U5007 ( .A(DATAI_8_), .B(keyinput_151), .ZN(n4551) );
  NAND3_X1 U5008 ( .A1(n4553), .A2(n4552), .A3(n4551), .ZN(n4554) );
  AOI21_X1 U5009 ( .B1(n4556), .B2(n4555), .A(n4554), .ZN(n4559) );
  INV_X1 U5010 ( .A(DATAI_6_), .ZN(n5162) );
  XNOR2_X1 U5011 ( .A(n5162), .B(keyinput_153), .ZN(n4558) );
  XOR2_X1 U5012 ( .A(DATAI_5_), .B(keyinput_154), .Z(n4557) );
  NOR3_X1 U5013 ( .A1(n4559), .A2(n4558), .A3(n4557), .ZN(n4562) );
  INV_X1 U5014 ( .A(DATAI_4_), .ZN(n5153) );
  XNOR2_X1 U5015 ( .A(n5153), .B(keyinput_155), .ZN(n4561) );
  XOR2_X1 U5016 ( .A(DATAI_3_), .B(keyinput_156), .Z(n4560) );
  NOR3_X1 U5017 ( .A1(n4562), .A2(n4561), .A3(n4560), .ZN(n4565) );
  XOR2_X1 U5018 ( .A(DATAI_2_), .B(keyinput_157), .Z(n4564) );
  XOR2_X1 U5019 ( .A(DATAI_1_), .B(keyinput_158), .Z(n4563) );
  OAI21_X1 U5020 ( .B1(n4565), .B2(n4564), .A(n4563), .ZN(n4571) );
  XOR2_X1 U5021 ( .A(DATAI_0_), .B(keyinput_159), .Z(n4570) );
  XOR2_X1 U5022 ( .A(REG3_REG_7__SCAN_IN), .B(keyinput_161), .Z(n4568) );
  XNOR2_X1 U5023 ( .A(U3149), .B(keyinput_160), .ZN(n4567) );
  XNOR2_X1 U5024 ( .A(REG3_REG_27__SCAN_IN), .B(keyinput_162), .ZN(n4566) );
  NAND3_X1 U5025 ( .A1(n4568), .A2(n4567), .A3(n4566), .ZN(n4569) );
  AOI21_X1 U5026 ( .B1(n4571), .B2(n4570), .A(n4569), .ZN(n4578) );
  XNOR2_X1 U5027 ( .A(n4572), .B(keyinput_163), .ZN(n4577) );
  XOR2_X1 U5028 ( .A(REG3_REG_10__SCAN_IN), .B(keyinput_165), .Z(n4575) );
  XNOR2_X1 U5029 ( .A(REG3_REG_23__SCAN_IN), .B(keyinput_164), .ZN(n4574) );
  XNOR2_X1 U5030 ( .A(REG3_REG_3__SCAN_IN), .B(keyinput_166), .ZN(n4573) );
  NOR3_X1 U5031 ( .A1(n4575), .A2(n4574), .A3(n4573), .ZN(n4576) );
  OAI21_X1 U5032 ( .B1(n4578), .B2(n4577), .A(n4576), .ZN(n4582) );
  XNOR2_X1 U5033 ( .A(REG3_REG_19__SCAN_IN), .B(keyinput_167), .ZN(n4581) );
  XNOR2_X1 U5034 ( .A(n4579), .B(keyinput_168), .ZN(n4580) );
  AOI21_X1 U5035 ( .B1(n4582), .B2(n4581), .A(n4580), .ZN(n4586) );
  XNOR2_X1 U5036 ( .A(REG3_REG_8__SCAN_IN), .B(keyinput_169), .ZN(n4585) );
  XOR2_X1 U5037 ( .A(REG3_REG_21__SCAN_IN), .B(keyinput_171), .Z(n4584) );
  XNOR2_X1 U5038 ( .A(REG3_REG_1__SCAN_IN), .B(keyinput_170), .ZN(n4583) );
  OAI211_X1 U5039 ( .C1(n4586), .C2(n4585), .A(n4584), .B(n4583), .ZN(n4589)
         );
  XNOR2_X1 U5040 ( .A(REG3_REG_12__SCAN_IN), .B(keyinput_172), .ZN(n4588) );
  XNOR2_X1 U5041 ( .A(REG3_REG_25__SCAN_IN), .B(keyinput_173), .ZN(n4587) );
  AOI21_X1 U5042 ( .B1(n4589), .B2(n4588), .A(n4587), .ZN(n4597) );
  XNOR2_X1 U5043 ( .A(n4590), .B(keyinput_174), .ZN(n4596) );
  XOR2_X1 U5044 ( .A(REG3_REG_5__SCAN_IN), .B(keyinput_175), .Z(n4594) );
  XNOR2_X1 U5045 ( .A(REG3_REG_4__SCAN_IN), .B(keyinput_178), .ZN(n4593) );
  XNOR2_X1 U5046 ( .A(REG3_REG_24__SCAN_IN), .B(keyinput_177), .ZN(n4592) );
  XNOR2_X1 U5047 ( .A(REG3_REG_17__SCAN_IN), .B(keyinput_176), .ZN(n4591) );
  NOR4_X1 U5048 ( .A1(n4594), .A2(n4593), .A3(n4592), .A4(n4591), .ZN(n4595)
         );
  OAI21_X1 U5049 ( .B1(n4597), .B2(n4596), .A(n4595), .ZN(n4601) );
  XNOR2_X1 U5050 ( .A(REG3_REG_20__SCAN_IN), .B(keyinput_181), .ZN(n4600) );
  XNOR2_X1 U5051 ( .A(REG3_REG_9__SCAN_IN), .B(keyinput_179), .ZN(n4599) );
  XNOR2_X1 U5052 ( .A(REG3_REG_0__SCAN_IN), .B(keyinput_180), .ZN(n4598) );
  NAND4_X1 U5053 ( .A1(n4601), .A2(n4600), .A3(n4599), .A4(n4598), .ZN(n4605)
         );
  XOR2_X1 U5054 ( .A(IR_REG_0__SCAN_IN), .B(keyinput_183), .Z(n4604) );
  XNOR2_X1 U5055 ( .A(IR_REG_1__SCAN_IN), .B(keyinput_184), .ZN(n4603) );
  XNOR2_X1 U5056 ( .A(REG3_REG_13__SCAN_IN), .B(keyinput_182), .ZN(n4602) );
  NAND4_X1 U5057 ( .A1(n4605), .A2(n4604), .A3(n4603), .A4(n4602), .ZN(n4614)
         );
  AOI22_X1 U5058 ( .A1(n2792), .A2(keyinput_189), .B1(n4800), .B2(keyinput_185), .ZN(n4606) );
  OAI221_X1 U5059 ( .B1(n2792), .B2(keyinput_189), .C1(n4800), .C2(
        keyinput_185), .A(n4606), .ZN(n4611) );
  XNOR2_X1 U5060 ( .A(n2778), .B(keyinput_186), .ZN(n4610) );
  XNOR2_X1 U5061 ( .A(n4607), .B(keyinput_187), .ZN(n4609) );
  XNOR2_X1 U5062 ( .A(IR_REG_5__SCAN_IN), .B(keyinput_188), .ZN(n4608) );
  NOR4_X1 U5063 ( .A1(n4611), .A2(n4610), .A3(n4609), .A4(n4608), .ZN(n4613)
         );
  XNOR2_X1 U5064 ( .A(IR_REG_7__SCAN_IN), .B(keyinput_190), .ZN(n4612) );
  AOI21_X1 U5065 ( .B1(n4614), .B2(n4613), .A(n4612), .ZN(n4618) );
  XNOR2_X1 U5066 ( .A(IR_REG_8__SCAN_IN), .B(keyinput_191), .ZN(n4617) );
  XNOR2_X1 U5067 ( .A(n2757), .B(keyinput_193), .ZN(n4616) );
  XNOR2_X1 U5068 ( .A(IR_REG_9__SCAN_IN), .B(keyinput_192), .ZN(n4615) );
  OAI211_X1 U5069 ( .C1(n4618), .C2(n4617), .A(n4616), .B(n4615), .ZN(n4622)
         );
  XNOR2_X1 U5070 ( .A(IR_REG_11__SCAN_IN), .B(keyinput_194), .ZN(n4621) );
  XNOR2_X1 U5071 ( .A(IR_REG_12__SCAN_IN), .B(keyinput_195), .ZN(n4620) );
  XNOR2_X1 U5072 ( .A(IR_REG_13__SCAN_IN), .B(keyinput_196), .ZN(n4619) );
  AOI211_X1 U5073 ( .C1(n4622), .C2(n4621), .A(n4620), .B(n4619), .ZN(n4627)
         );
  XNOR2_X1 U5074 ( .A(IR_REG_14__SCAN_IN), .B(keyinput_197), .ZN(n4626) );
  XNOR2_X1 U5075 ( .A(n4623), .B(keyinput_199), .ZN(n4625) );
  XNOR2_X1 U5076 ( .A(IR_REG_15__SCAN_IN), .B(keyinput_198), .ZN(n4624) );
  OAI211_X1 U5077 ( .C1(n4627), .C2(n4626), .A(n4625), .B(n4624), .ZN(n4632)
         );
  XNOR2_X1 U5078 ( .A(n4628), .B(keyinput_201), .ZN(n4631) );
  XNOR2_X1 U5079 ( .A(IR_REG_17__SCAN_IN), .B(keyinput_200), .ZN(n4630) );
  XNOR2_X1 U5080 ( .A(IR_REG_19__SCAN_IN), .B(keyinput_202), .ZN(n4629) );
  NAND4_X1 U5081 ( .A1(n4632), .A2(n4631), .A3(n4630), .A4(n4629), .ZN(n4636)
         );
  XNOR2_X1 U5082 ( .A(n4633), .B(keyinput_203), .ZN(n4635) );
  XNOR2_X1 U5083 ( .A(IR_REG_21__SCAN_IN), .B(keyinput_204), .ZN(n4634) );
  AOI21_X1 U5084 ( .B1(n4636), .B2(n4635), .A(n4634), .ZN(n4639) );
  XNOR2_X1 U5085 ( .A(IR_REG_22__SCAN_IN), .B(keyinput_205), .ZN(n4638) );
  XNOR2_X1 U5086 ( .A(n4830), .B(keyinput_206), .ZN(n4637) );
  OAI21_X1 U5087 ( .B1(n4639), .B2(n4638), .A(n4637), .ZN(n4643) );
  XNOR2_X1 U5088 ( .A(IR_REG_24__SCAN_IN), .B(keyinput_207), .ZN(n4642) );
  XNOR2_X1 U5089 ( .A(n4834), .B(keyinput_208), .ZN(n4641) );
  XNOR2_X1 U5090 ( .A(IR_REG_26__SCAN_IN), .B(keyinput_209), .ZN(n4640) );
  AOI211_X1 U5091 ( .C1(n4643), .C2(n4642), .A(n4641), .B(n4640), .ZN(n4649)
         );
  XOR2_X1 U5092 ( .A(IR_REG_27__SCAN_IN), .B(keyinput_210), .Z(n4645) );
  XNOR2_X1 U5093 ( .A(IR_REG_28__SCAN_IN), .B(keyinput_211), .ZN(n4644) );
  NAND2_X1 U5094 ( .A1(n4645), .A2(n4644), .ZN(n4648) );
  XOR2_X1 U5095 ( .A(IR_REG_30__SCAN_IN), .B(keyinput_213), .Z(n4647) );
  XNOR2_X1 U5096 ( .A(IR_REG_29__SCAN_IN), .B(keyinput_212), .ZN(n4646) );
  OAI211_X1 U5097 ( .C1(n4649), .C2(n4648), .A(n4647), .B(n4646), .ZN(n4652)
         );
  XNOR2_X1 U5098 ( .A(IR_REG_31__SCAN_IN), .B(keyinput_214), .ZN(n4651) );
  XOR2_X1 U5099 ( .A(D_REG_0__SCAN_IN), .B(keyinput_215), .Z(n4650) );
  AOI21_X1 U5100 ( .B1(n4652), .B2(n4651), .A(n4650), .ZN(n4658) );
  XNOR2_X1 U5101 ( .A(D_REG_1__SCAN_IN), .B(keyinput_216), .ZN(n4657) );
  XOR2_X1 U5102 ( .A(D_REG_4__SCAN_IN), .B(keyinput_219), .Z(n4655) );
  XOR2_X1 U5103 ( .A(D_REG_3__SCAN_IN), .B(keyinput_218), .Z(n4654) );
  INV_X1 U5104 ( .A(D_REG_2__SCAN_IN), .ZN(n4927) );
  XNOR2_X1 U5105 ( .A(n4927), .B(keyinput_217), .ZN(n4653) );
  NOR3_X1 U5106 ( .A1(n4655), .A2(n4654), .A3(n4653), .ZN(n4656) );
  OAI21_X1 U5107 ( .B1(n4658), .B2(n4657), .A(n4656), .ZN(n4661) );
  XNOR2_X1 U5108 ( .A(D_REG_5__SCAN_IN), .B(keyinput_220), .ZN(n4660) );
  INV_X1 U5109 ( .A(D_REG_6__SCAN_IN), .ZN(n4931) );
  XNOR2_X1 U5110 ( .A(n4931), .B(keyinput_221), .ZN(n4659) );
  AOI21_X1 U5111 ( .B1(n4661), .B2(n4660), .A(n4659), .ZN(n4667) );
  XNOR2_X1 U5112 ( .A(D_REG_7__SCAN_IN), .B(keyinput_222), .ZN(n4666) );
  XOR2_X1 U5113 ( .A(D_REG_9__SCAN_IN), .B(keyinput_224), .Z(n4664) );
  INV_X1 U5114 ( .A(D_REG_10__SCAN_IN), .ZN(n4935) );
  XNOR2_X1 U5115 ( .A(n4935), .B(keyinput_225), .ZN(n4663) );
  XNOR2_X1 U5116 ( .A(D_REG_8__SCAN_IN), .B(keyinput_223), .ZN(n4662) );
  NOR3_X1 U5117 ( .A1(n4664), .A2(n4663), .A3(n4662), .ZN(n4665) );
  OAI21_X1 U5118 ( .B1(n4667), .B2(n4666), .A(n4665), .ZN(n4670) );
  XNOR2_X1 U5119 ( .A(D_REG_11__SCAN_IN), .B(keyinput_226), .ZN(n4669) );
  XNOR2_X1 U5120 ( .A(D_REG_12__SCAN_IN), .B(keyinput_227), .ZN(n4668) );
  NAND3_X1 U5121 ( .A1(n4670), .A2(n4669), .A3(n4668), .ZN(n4673) );
  XOR2_X1 U5122 ( .A(D_REG_14__SCAN_IN), .B(keyinput_229), .Z(n4672) );
  XNOR2_X1 U5123 ( .A(D_REG_13__SCAN_IN), .B(keyinput_228), .ZN(n4671) );
  NAND3_X1 U5124 ( .A1(n4673), .A2(n4672), .A3(n4671), .ZN(n4676) );
  INV_X1 U5125 ( .A(D_REG_15__SCAN_IN), .ZN(n4939) );
  XNOR2_X1 U5126 ( .A(n4939), .B(keyinput_230), .ZN(n4675) );
  INV_X1 U5127 ( .A(D_REG_16__SCAN_IN), .ZN(n4940) );
  XNOR2_X1 U5128 ( .A(n4940), .B(keyinput_231), .ZN(n4674) );
  AOI21_X1 U5129 ( .B1(n4676), .B2(n4675), .A(n4674), .ZN(n4680) );
  XOR2_X1 U5130 ( .A(D_REG_17__SCAN_IN), .B(keyinput_232), .Z(n4679) );
  INV_X1 U5131 ( .A(D_REG_18__SCAN_IN), .ZN(n4942) );
  XNOR2_X1 U5132 ( .A(n4942), .B(keyinput_233), .ZN(n4678) );
  XNOR2_X1 U5133 ( .A(D_REG_19__SCAN_IN), .B(keyinput_234), .ZN(n4677) );
  NOR4_X1 U5134 ( .A1(n4680), .A2(n4679), .A3(n4678), .A4(n4677), .ZN(n4686)
         );
  INV_X1 U5135 ( .A(D_REG_20__SCAN_IN), .ZN(n4944) );
  XNOR2_X1 U5136 ( .A(n4944), .B(keyinput_235), .ZN(n4685) );
  INV_X1 U5137 ( .A(D_REG_23__SCAN_IN), .ZN(n4946) );
  XNOR2_X1 U5138 ( .A(n4946), .B(keyinput_238), .ZN(n4683) );
  INV_X1 U5139 ( .A(D_REG_21__SCAN_IN), .ZN(n4945) );
  XNOR2_X1 U5140 ( .A(n4945), .B(keyinput_236), .ZN(n4682) );
  XNOR2_X1 U5141 ( .A(D_REG_22__SCAN_IN), .B(keyinput_237), .ZN(n4681) );
  NOR3_X1 U5142 ( .A1(n4683), .A2(n4682), .A3(n4681), .ZN(n4684) );
  OAI21_X1 U5143 ( .B1(n4686), .B2(n4685), .A(n4684), .ZN(n4693) );
  XOR2_X1 U5144 ( .A(D_REG_28__SCAN_IN), .B(keyinput_243), .Z(n4692) );
  XOR2_X1 U5145 ( .A(keyinput_240), .B(D_REG_25__SCAN_IN), .Z(n4689) );
  XOR2_X1 U5146 ( .A(keyinput_242), .B(D_REG_27__SCAN_IN), .Z(n4688) );
  XNOR2_X1 U5147 ( .A(D_REG_24__SCAN_IN), .B(keyinput_239), .ZN(n4687) );
  NOR3_X1 U5148 ( .A1(n4689), .A2(n4688), .A3(n4687), .ZN(n4691) );
  XNOR2_X1 U5149 ( .A(D_REG_26__SCAN_IN), .B(keyinput_241), .ZN(n4690) );
  NAND4_X1 U5150 ( .A1(n4693), .A2(n4692), .A3(n4691), .A4(n4690), .ZN(n4697)
         );
  XOR2_X1 U5151 ( .A(D_REG_30__SCAN_IN), .B(keyinput_245), .Z(n4696) );
  XOR2_X1 U5152 ( .A(D_REG_29__SCAN_IN), .B(keyinput_244), .Z(n4695) );
  INV_X1 U5153 ( .A(D_REG_31__SCAN_IN), .ZN(n4952) );
  XNOR2_X1 U5154 ( .A(n4952), .B(keyinput_246), .ZN(n4694) );
  NAND4_X1 U5155 ( .A1(n4697), .A2(n4696), .A3(n4695), .A4(n4694), .ZN(n4700)
         );
  XOR2_X1 U5156 ( .A(REG0_REG_0__SCAN_IN), .B(keyinput_247), .Z(n4699) );
  INV_X1 U5157 ( .A(REG0_REG_1__SCAN_IN), .ZN(n4894) );
  XNOR2_X1 U5158 ( .A(n4894), .B(keyinput_248), .ZN(n4698) );
  NAND3_X1 U5159 ( .A1(n4700), .A2(n4699), .A3(n4698), .ZN(n4705) );
  XNOR2_X1 U5160 ( .A(n4899), .B(keyinput_250), .ZN(n4704) );
  INV_X1 U5161 ( .A(REG0_REG_2__SCAN_IN), .ZN(n4701) );
  XNOR2_X1 U5162 ( .A(n4701), .B(keyinput_249), .ZN(n4703) );
  XNOR2_X1 U5163 ( .A(REG0_REG_4__SCAN_IN), .B(keyinput_251), .ZN(n4702) );
  NAND4_X1 U5164 ( .A1(n4705), .A2(n4704), .A3(n4703), .A4(n4702), .ZN(n4708)
         );
  XOR2_X1 U5165 ( .A(REG0_REG_5__SCAN_IN), .B(keyinput_252), .Z(n4707) );
  XNOR2_X1 U5166 ( .A(REG0_REG_6__SCAN_IN), .B(keyinput_253), .ZN(n4706) );
  NAND3_X1 U5167 ( .A1(n4708), .A2(n4707), .A3(n4706), .ZN(n4913) );
  XNOR2_X1 U5168 ( .A(REG0_REG_7__SCAN_IN), .B(keyinput_254), .ZN(n4912) );
  XNOR2_X1 U5169 ( .A(n4709), .B(keyinput_255), .ZN(n4911) );
  XOR2_X1 U5170 ( .A(DATAI_31_), .B(keyinput_0), .Z(n4713) );
  XOR2_X1 U5171 ( .A(DATAI_30_), .B(keyinput_1), .Z(n4712) );
  XOR2_X1 U5172 ( .A(DATAI_29_), .B(keyinput_2), .Z(n4711) );
  XOR2_X1 U5173 ( .A(DATAI_28_), .B(keyinput_3), .Z(n4710) );
  AOI211_X1 U5174 ( .C1(n4713), .C2(n4712), .A(n4711), .B(n4710), .ZN(n4716)
         );
  XNOR2_X1 U5175 ( .A(DATAI_27_), .B(keyinput_4), .ZN(n4715) );
  XNOR2_X1 U5176 ( .A(DATAI_26_), .B(keyinput_5), .ZN(n4714) );
  OAI21_X1 U5177 ( .B1(n4716), .B2(n4715), .A(n4714), .ZN(n4719) );
  XOR2_X1 U5178 ( .A(DATAI_25_), .B(keyinput_6), .Z(n4718) );
  XOR2_X1 U5179 ( .A(DATAI_24_), .B(keyinput_7), .Z(n4717) );
  AOI21_X1 U5180 ( .B1(n4719), .B2(n4718), .A(n4717), .ZN(n4722) );
  XNOR2_X1 U5181 ( .A(DATAI_23_), .B(keyinput_8), .ZN(n4721) );
  XOR2_X1 U5182 ( .A(DATAI_22_), .B(keyinput_9), .Z(n4720) );
  OAI21_X1 U5183 ( .B1(n4722), .B2(n4721), .A(n4720), .ZN(n4725) );
  XNOR2_X1 U5184 ( .A(DATAI_21_), .B(keyinput_10), .ZN(n4724) );
  XOR2_X1 U5185 ( .A(DATAI_20_), .B(keyinput_11), .Z(n4723) );
  AOI21_X1 U5186 ( .B1(n4725), .B2(n4724), .A(n4723), .ZN(n4728) );
  XOR2_X1 U5187 ( .A(DATAI_18_), .B(keyinput_13), .Z(n4727) );
  XNOR2_X1 U5188 ( .A(DATAI_19_), .B(keyinput_12), .ZN(n4726) );
  NOR3_X1 U5189 ( .A1(n4728), .A2(n4727), .A3(n4726), .ZN(n4738) );
  XOR2_X1 U5190 ( .A(DATAI_17_), .B(keyinput_14), .Z(n4737) );
  XNOR2_X1 U5191 ( .A(DATAI_13_), .B(keyinput_18), .ZN(n4732) );
  XNOR2_X1 U5192 ( .A(DATAI_16_), .B(keyinput_15), .ZN(n4731) );
  XNOR2_X1 U5193 ( .A(DATAI_11_), .B(keyinput_20), .ZN(n4730) );
  XNOR2_X1 U5194 ( .A(DATAI_12_), .B(keyinput_19), .ZN(n4729) );
  NAND4_X1 U5195 ( .A1(n4732), .A2(n4731), .A3(n4730), .A4(n4729), .ZN(n4735)
         );
  XNOR2_X1 U5196 ( .A(DATAI_15_), .B(keyinput_16), .ZN(n4734) );
  XNOR2_X1 U5197 ( .A(DATAI_14_), .B(keyinput_17), .ZN(n4733) );
  NOR3_X1 U5198 ( .A1(n4735), .A2(n4734), .A3(n4733), .ZN(n4736) );
  OAI21_X1 U5199 ( .B1(n4738), .B2(n4737), .A(n4736), .ZN(n4745) );
  XNOR2_X1 U5200 ( .A(DATAI_10_), .B(keyinput_21), .ZN(n4744) );
  XOR2_X1 U5201 ( .A(DATAI_7_), .B(keyinput_24), .Z(n4742) );
  XNOR2_X1 U5202 ( .A(n4739), .B(keyinput_23), .ZN(n4741) );
  XNOR2_X1 U5203 ( .A(DATAI_9_), .B(keyinput_22), .ZN(n4740) );
  NAND3_X1 U5204 ( .A1(n4742), .A2(n4741), .A3(n4740), .ZN(n4743) );
  AOI21_X1 U5205 ( .B1(n4745), .B2(n4744), .A(n4743), .ZN(n4748) );
  XOR2_X1 U5206 ( .A(DATAI_5_), .B(keyinput_26), .Z(n4747) );
  XNOR2_X1 U5207 ( .A(DATAI_6_), .B(keyinput_25), .ZN(n4746) );
  NOR3_X1 U5208 ( .A1(n4748), .A2(n4747), .A3(n4746), .ZN(n4751) );
  XOR2_X1 U5209 ( .A(DATAI_3_), .B(keyinput_28), .Z(n4750) );
  XNOR2_X1 U5210 ( .A(DATAI_4_), .B(keyinput_27), .ZN(n4749) );
  NOR3_X1 U5211 ( .A1(n4751), .A2(n4750), .A3(n4749), .ZN(n4754) );
  XOR2_X1 U5212 ( .A(DATAI_2_), .B(keyinput_29), .Z(n4753) );
  XNOR2_X1 U5213 ( .A(DATAI_1_), .B(keyinput_30), .ZN(n4752) );
  OAI21_X1 U5214 ( .B1(n4754), .B2(n4753), .A(n4752), .ZN(n4761) );
  XNOR2_X1 U5215 ( .A(DATAI_0_), .B(keyinput_31), .ZN(n4760) );
  XOR2_X1 U5216 ( .A(REG3_REG_7__SCAN_IN), .B(keyinput_33), .Z(n4758) );
  XNOR2_X1 U5217 ( .A(n4755), .B(keyinput_34), .ZN(n4757) );
  XNOR2_X1 U5218 ( .A(STATE_REG_SCAN_IN), .B(keyinput_32), .ZN(n4756) );
  NAND3_X1 U5219 ( .A1(n4758), .A2(n4757), .A3(n4756), .ZN(n4759) );
  AOI21_X1 U5220 ( .B1(n4761), .B2(n4760), .A(n4759), .ZN(n4768) );
  XNOR2_X1 U5221 ( .A(REG3_REG_14__SCAN_IN), .B(keyinput_35), .ZN(n4767) );
  XNOR2_X1 U5222 ( .A(n4762), .B(keyinput_36), .ZN(n4765) );
  XNOR2_X1 U5223 ( .A(REG3_REG_3__SCAN_IN), .B(keyinput_38), .ZN(n4764) );
  XNOR2_X1 U5224 ( .A(REG3_REG_10__SCAN_IN), .B(keyinput_37), .ZN(n4763) );
  NOR3_X1 U5225 ( .A1(n4765), .A2(n4764), .A3(n4763), .ZN(n4766) );
  OAI21_X1 U5226 ( .B1(n4768), .B2(n4767), .A(n4766), .ZN(n4771) );
  XNOR2_X1 U5227 ( .A(REG3_REG_19__SCAN_IN), .B(keyinput_39), .ZN(n4770) );
  XNOR2_X1 U5228 ( .A(REG3_REG_28__SCAN_IN), .B(keyinput_40), .ZN(n4769) );
  AOI21_X1 U5229 ( .B1(n4771), .B2(n4770), .A(n4769), .ZN(n4775) );
  XOR2_X1 U5230 ( .A(REG3_REG_8__SCAN_IN), .B(keyinput_41), .Z(n4774) );
  XNOR2_X1 U5231 ( .A(REG3_REG_21__SCAN_IN), .B(keyinput_43), .ZN(n4773) );
  XNOR2_X1 U5232 ( .A(REG3_REG_1__SCAN_IN), .B(keyinput_42), .ZN(n4772) );
  OAI211_X1 U5233 ( .C1(n4775), .C2(n4774), .A(n4773), .B(n4772), .ZN(n4780)
         );
  XNOR2_X1 U5234 ( .A(n4776), .B(keyinput_44), .ZN(n4779) );
  XNOR2_X1 U5235 ( .A(n4777), .B(keyinput_45), .ZN(n4778) );
  AOI21_X1 U5236 ( .B1(n4780), .B2(n4779), .A(n4778), .ZN(n4788) );
  XNOR2_X1 U5237 ( .A(keyinput_46), .B(REG3_REG_16__SCAN_IN), .ZN(n4787) );
  XOR2_X1 U5238 ( .A(REG3_REG_5__SCAN_IN), .B(keyinput_47), .Z(n4785) );
  XNOR2_X1 U5239 ( .A(n4781), .B(keyinput_49), .ZN(n4784) );
  XNOR2_X1 U5240 ( .A(REG3_REG_17__SCAN_IN), .B(keyinput_48), .ZN(n4783) );
  XNOR2_X1 U5241 ( .A(REG3_REG_4__SCAN_IN), .B(keyinput_50), .ZN(n4782) );
  NOR4_X1 U5242 ( .A1(n4785), .A2(n4784), .A3(n4783), .A4(n4782), .ZN(n4786)
         );
  OAI21_X1 U5243 ( .B1(n4788), .B2(n4787), .A(n4786), .ZN(n4794) );
  INV_X1 U5244 ( .A(REG3_REG_9__SCAN_IN), .ZN(n4790) );
  OAI22_X1 U5245 ( .A1(n4790), .A2(keyinput_51), .B1(REG3_REG_20__SCAN_IN), 
        .B2(keyinput_53), .ZN(n4789) );
  AOI21_X1 U5246 ( .B1(n4790), .B2(keyinput_51), .A(n4789), .ZN(n4793) );
  XNOR2_X1 U5247 ( .A(REG3_REG_0__SCAN_IN), .B(keyinput_52), .ZN(n4792) );
  NAND2_X1 U5248 ( .A1(REG3_REG_20__SCAN_IN), .A2(keyinput_53), .ZN(n4791) );
  NAND4_X1 U5249 ( .A1(n4794), .A2(n4793), .A3(n4792), .A4(n4791), .ZN(n4798)
         );
  XNOR2_X1 U5250 ( .A(IR_REG_1__SCAN_IN), .B(keyinput_56), .ZN(n4797) );
  XNOR2_X1 U5251 ( .A(IR_REG_0__SCAN_IN), .B(keyinput_55), .ZN(n4796) );
  XNOR2_X1 U5252 ( .A(REG3_REG_13__SCAN_IN), .B(keyinput_54), .ZN(n4795) );
  NAND4_X1 U5253 ( .A1(n4798), .A2(n4797), .A3(n4796), .A4(n4795), .ZN(n4805)
         );
  OAI22_X1 U5254 ( .A1(IR_REG_3__SCAN_IN), .A2(keyinput_58), .B1(keyinput_61), 
        .B2(IR_REG_6__SCAN_IN), .ZN(n4799) );
  AOI221_X1 U5255 ( .B1(IR_REG_3__SCAN_IN), .B2(keyinput_58), .C1(
        IR_REG_6__SCAN_IN), .C2(keyinput_61), .A(n4799), .ZN(n4804) );
  XNOR2_X1 U5256 ( .A(n4800), .B(keyinput_57), .ZN(n4803) );
  OAI22_X1 U5257 ( .A1(IR_REG_4__SCAN_IN), .A2(keyinput_59), .B1(keyinput_60), 
        .B2(IR_REG_5__SCAN_IN), .ZN(n4801) );
  AOI221_X1 U5258 ( .B1(IR_REG_4__SCAN_IN), .B2(keyinput_59), .C1(
        IR_REG_5__SCAN_IN), .C2(keyinput_60), .A(n4801), .ZN(n4802) );
  NAND4_X1 U5259 ( .A1(n4805), .A2(n4804), .A3(n4803), .A4(n4802), .ZN(n4809)
         );
  XNOR2_X1 U5260 ( .A(n4806), .B(keyinput_62), .ZN(n4808) );
  XOR2_X1 U5261 ( .A(IR_REG_8__SCAN_IN), .B(keyinput_63), .Z(n4807) );
  AOI21_X1 U5262 ( .B1(n4809), .B2(n4808), .A(n4807), .ZN(n4812) );
  XNOR2_X1 U5263 ( .A(n2757), .B(keyinput_65), .ZN(n4811) );
  XOR2_X1 U5264 ( .A(IR_REG_9__SCAN_IN), .B(keyinput_64), .Z(n4810) );
  NOR3_X1 U5265 ( .A1(n4812), .A2(n4811), .A3(n4810), .ZN(n4817) );
  XNOR2_X1 U5266 ( .A(IR_REG_11__SCAN_IN), .B(keyinput_66), .ZN(n4816) );
  XNOR2_X1 U5267 ( .A(n4813), .B(keyinput_67), .ZN(n4815) );
  XNOR2_X1 U5268 ( .A(IR_REG_13__SCAN_IN), .B(keyinput_68), .ZN(n4814) );
  OAI211_X1 U5269 ( .C1(n4817), .C2(n4816), .A(n4815), .B(n4814), .ZN(n4821)
         );
  XNOR2_X1 U5270 ( .A(IR_REG_14__SCAN_IN), .B(keyinput_69), .ZN(n4820) );
  XNOR2_X1 U5271 ( .A(IR_REG_16__SCAN_IN), .B(keyinput_71), .ZN(n4819) );
  XNOR2_X1 U5272 ( .A(IR_REG_15__SCAN_IN), .B(keyinput_70), .ZN(n4818) );
  AOI211_X1 U5273 ( .C1(n4821), .C2(n4820), .A(n4819), .B(n4818), .ZN(n4826)
         );
  XNOR2_X1 U5274 ( .A(n4822), .B(keyinput_72), .ZN(n4825) );
  XNOR2_X1 U5275 ( .A(IR_REG_19__SCAN_IN), .B(keyinput_74), .ZN(n4824) );
  XNOR2_X1 U5276 ( .A(IR_REG_18__SCAN_IN), .B(keyinput_73), .ZN(n4823) );
  NOR4_X1 U5277 ( .A1(n4826), .A2(n4825), .A3(n4824), .A4(n4823), .ZN(n4829)
         );
  XNOR2_X1 U5278 ( .A(IR_REG_20__SCAN_IN), .B(keyinput_75), .ZN(n4828) );
  XNOR2_X1 U5279 ( .A(n2867), .B(keyinput_76), .ZN(n4827) );
  OAI21_X1 U5280 ( .B1(n4829), .B2(n4828), .A(n4827), .ZN(n4833) );
  XNOR2_X1 U5281 ( .A(IR_REG_22__SCAN_IN), .B(keyinput_77), .ZN(n4832) );
  XNOR2_X1 U5282 ( .A(n4830), .B(keyinput_78), .ZN(n4831) );
  AOI21_X1 U5283 ( .B1(n4833), .B2(n4832), .A(n4831), .ZN(n4838) );
  XNOR2_X1 U5284 ( .A(IR_REG_24__SCAN_IN), .B(keyinput_79), .ZN(n4837) );
  XNOR2_X1 U5285 ( .A(n4834), .B(keyinput_80), .ZN(n4836) );
  XOR2_X1 U5286 ( .A(IR_REG_26__SCAN_IN), .B(keyinput_81), .Z(n4835) );
  OAI211_X1 U5287 ( .C1(n4838), .C2(n4837), .A(n4836), .B(n4835), .ZN(n4842)
         );
  XOR2_X1 U5288 ( .A(IR_REG_27__SCAN_IN), .B(keyinput_82), .Z(n4841) );
  XNOR2_X1 U5289 ( .A(n4839), .B(keyinput_83), .ZN(n4840) );
  NAND3_X1 U5290 ( .A1(n4842), .A2(n4841), .A3(n4840), .ZN(n4846) );
  XOR2_X1 U5291 ( .A(IR_REG_30__SCAN_IN), .B(keyinput_85), .Z(n4845) );
  XNOR2_X1 U5292 ( .A(n4843), .B(keyinput_84), .ZN(n4844) );
  NAND3_X1 U5293 ( .A1(n4846), .A2(n4845), .A3(n4844), .ZN(n4849) );
  XOR2_X1 U5294 ( .A(IR_REG_31__SCAN_IN), .B(keyinput_86), .Z(n4848) );
  XNOR2_X1 U5295 ( .A(D_REG_0__SCAN_IN), .B(keyinput_87), .ZN(n4847) );
  AOI21_X1 U5296 ( .B1(n4849), .B2(n4848), .A(n4847), .ZN(n4855) );
  XOR2_X1 U5297 ( .A(D_REG_1__SCAN_IN), .B(keyinput_88), .Z(n4854) );
  XOR2_X1 U5298 ( .A(keyinput_91), .B(D_REG_4__SCAN_IN), .Z(n4852) );
  XOR2_X1 U5299 ( .A(keyinput_90), .B(D_REG_3__SCAN_IN), .Z(n4851) );
  XNOR2_X1 U5300 ( .A(keyinput_89), .B(D_REG_2__SCAN_IN), .ZN(n4850) );
  NOR3_X1 U5301 ( .A1(n4852), .A2(n4851), .A3(n4850), .ZN(n4853) );
  OAI21_X1 U5302 ( .B1(n4855), .B2(n4854), .A(n4853), .ZN(n4858) );
  XNOR2_X1 U5303 ( .A(keyinput_92), .B(D_REG_5__SCAN_IN), .ZN(n4857) );
  XNOR2_X1 U5304 ( .A(keyinput_93), .B(D_REG_6__SCAN_IN), .ZN(n4856) );
  AOI21_X1 U5305 ( .B1(n4858), .B2(n4857), .A(n4856), .ZN(n4864) );
  XNOR2_X1 U5306 ( .A(keyinput_94), .B(D_REG_7__SCAN_IN), .ZN(n4863) );
  XOR2_X1 U5307 ( .A(keyinput_96), .B(D_REG_9__SCAN_IN), .Z(n4861) );
  INV_X1 U5308 ( .A(D_REG_8__SCAN_IN), .ZN(n4933) );
  XNOR2_X1 U5309 ( .A(n4933), .B(keyinput_95), .ZN(n4860) );
  XNOR2_X1 U5310 ( .A(keyinput_97), .B(D_REG_10__SCAN_IN), .ZN(n4859) );
  NOR3_X1 U5311 ( .A1(n4861), .A2(n4860), .A3(n4859), .ZN(n4862) );
  OAI21_X1 U5312 ( .B1(n4864), .B2(n4863), .A(n4862), .ZN(n4867) );
  INV_X1 U5313 ( .A(D_REG_11__SCAN_IN), .ZN(n4936) );
  XNOR2_X1 U5314 ( .A(n4936), .B(keyinput_98), .ZN(n4866) );
  INV_X1 U5315 ( .A(D_REG_12__SCAN_IN), .ZN(n4937) );
  XNOR2_X1 U5316 ( .A(n4937), .B(keyinput_99), .ZN(n4865) );
  NAND3_X1 U5317 ( .A1(n4867), .A2(n4866), .A3(n4865), .ZN(n4870) );
  INV_X1 U5318 ( .A(D_REG_13__SCAN_IN), .ZN(n4938) );
  XNOR2_X1 U5319 ( .A(n4938), .B(keyinput_100), .ZN(n4869) );
  XOR2_X1 U5320 ( .A(D_REG_14__SCAN_IN), .B(keyinput_101), .Z(n4868) );
  NAND3_X1 U5321 ( .A1(n4870), .A2(n4869), .A3(n4868), .ZN(n4873) );
  XNOR2_X1 U5322 ( .A(keyinput_102), .B(D_REG_15__SCAN_IN), .ZN(n4872) );
  XNOR2_X1 U5323 ( .A(n4940), .B(keyinput_103), .ZN(n4871) );
  AOI21_X1 U5324 ( .B1(n4873), .B2(n4872), .A(n4871), .ZN(n4877) );
  INV_X1 U5325 ( .A(D_REG_19__SCAN_IN), .ZN(n4943) );
  XNOR2_X1 U5326 ( .A(n4943), .B(keyinput_106), .ZN(n4876) );
  XOR2_X1 U5327 ( .A(keyinput_104), .B(D_REG_17__SCAN_IN), .Z(n4875) );
  XNOR2_X1 U5328 ( .A(keyinput_105), .B(D_REG_18__SCAN_IN), .ZN(n4874) );
  NOR4_X1 U5329 ( .A1(n4877), .A2(n4876), .A3(n4875), .A4(n4874), .ZN(n4883)
         );
  XNOR2_X1 U5330 ( .A(n4944), .B(keyinput_107), .ZN(n4882) );
  XNOR2_X1 U5331 ( .A(n4945), .B(keyinput_108), .ZN(n4880) );
  XNOR2_X1 U5332 ( .A(keyinput_110), .B(D_REG_23__SCAN_IN), .ZN(n4879) );
  XNOR2_X1 U5333 ( .A(D_REG_22__SCAN_IN), .B(keyinput_109), .ZN(n4878) );
  NOR3_X1 U5334 ( .A1(n4880), .A2(n4879), .A3(n4878), .ZN(n4881) );
  OAI21_X1 U5335 ( .B1(n4883), .B2(n4882), .A(n4881), .ZN(n4889) );
  INV_X1 U5336 ( .A(D_REG_28__SCAN_IN), .ZN(n4950) );
  OAI22_X1 U5337 ( .A1(n4950), .A2(keyinput_115), .B1(D_REG_24__SCAN_IN), .B2(
        keyinput_111), .ZN(n4884) );
  AOI221_X1 U5338 ( .B1(n4950), .B2(keyinput_115), .C1(keyinput_111), .C2(
        D_REG_24__SCAN_IN), .A(n4884), .ZN(n4888) );
  INV_X1 U5339 ( .A(D_REG_26__SCAN_IN), .ZN(n4948) );
  XNOR2_X1 U5340 ( .A(n4948), .B(keyinput_113), .ZN(n4887) );
  INV_X1 U5341 ( .A(D_REG_27__SCAN_IN), .ZN(n4949) );
  INV_X1 U5342 ( .A(D_REG_25__SCAN_IN), .ZN(n4947) );
  OAI22_X1 U5343 ( .A1(n4949), .A2(keyinput_114), .B1(n4947), .B2(keyinput_112), .ZN(n4885) );
  AOI221_X1 U5344 ( .B1(n4949), .B2(keyinput_114), .C1(keyinput_112), .C2(
        n4947), .A(n4885), .ZN(n4886) );
  NAND4_X1 U5345 ( .A1(n4889), .A2(n4888), .A3(n4887), .A4(n4886), .ZN(n4893)
         );
  XOR2_X1 U5346 ( .A(D_REG_29__SCAN_IN), .B(keyinput_116), .Z(n4892) );
  XNOR2_X1 U5347 ( .A(keyinput_118), .B(D_REG_31__SCAN_IN), .ZN(n4891) );
  XNOR2_X1 U5348 ( .A(D_REG_30__SCAN_IN), .B(keyinput_117), .ZN(n4890) );
  NAND4_X1 U5349 ( .A1(n4893), .A2(n4892), .A3(n4891), .A4(n4890), .ZN(n4897)
         );
  XNOR2_X1 U5350 ( .A(n4894), .B(keyinput_120), .ZN(n4896) );
  XNOR2_X1 U5351 ( .A(REG0_REG_0__SCAN_IN), .B(keyinput_119), .ZN(n4895) );
  NAND3_X1 U5352 ( .A1(n4897), .A2(n4896), .A3(n4895), .ZN(n4903) );
  XNOR2_X1 U5353 ( .A(n4898), .B(keyinput_123), .ZN(n4902) );
  XNOR2_X1 U5354 ( .A(n4899), .B(keyinput_122), .ZN(n4901) );
  XNOR2_X1 U5355 ( .A(REG0_REG_2__SCAN_IN), .B(keyinput_121), .ZN(n4900) );
  NAND4_X1 U5356 ( .A1(n4903), .A2(n4902), .A3(n4901), .A4(n4900), .ZN(n4906)
         );
  XOR2_X1 U5357 ( .A(REG0_REG_5__SCAN_IN), .B(keyinput_124), .Z(n4905) );
  XNOR2_X1 U5358 ( .A(REG0_REG_6__SCAN_IN), .B(keyinput_125), .ZN(n4904) );
  NAND3_X1 U5359 ( .A1(n4906), .A2(n4905), .A3(n4904), .ZN(n4909) );
  XNOR2_X1 U5360 ( .A(REG0_REG_7__SCAN_IN), .B(keyinput_126), .ZN(n4908) );
  XOR2_X1 U5361 ( .A(keyinput_255), .B(keyinput_127), .Z(n4907) );
  AOI21_X1 U5362 ( .B1(n4909), .B2(n4908), .A(n4907), .ZN(n4910) );
  AOI211_X1 U5363 ( .C1(n4913), .C2(n4912), .A(n4911), .B(n4910), .ZN(n4914)
         );
  XOR2_X1 U5364 ( .A(n4915), .B(n4914), .Z(U3477) );
  NOR3_X1 U5365 ( .A1(n4916), .A2(IR_REG_30__SCAN_IN), .A3(n2871), .ZN(n4917)
         );
  MUX2_X1 U5366 ( .A(DATAI_31_), .B(n4917), .S(STATE_REG_SCAN_IN), .Z(U3321)
         );
  MUX2_X1 U5367 ( .A(n4918), .B(DATAI_29_), .S(U3149), .Z(U3323) );
  MUX2_X1 U5368 ( .A(n4954), .B(DATAI_27_), .S(U3149), .Z(U3325) );
  MUX2_X1 U5369 ( .A(n4919), .B(DATAI_26_), .S(U3149), .Z(U3326) );
  MUX2_X1 U5370 ( .A(DATAI_25_), .B(n4920), .S(STATE_REG_SCAN_IN), .Z(U3327)
         );
  MUX2_X1 U5371 ( .A(DATAI_24_), .B(n2975), .S(STATE_REG_SCAN_IN), .Z(U3328)
         );
  MUX2_X1 U5372 ( .A(n4921), .B(DATAI_21_), .S(U3149), .Z(U3331) );
  MUX2_X1 U5373 ( .A(DATAI_20_), .B(n4922), .S(STATE_REG_SCAN_IN), .Z(U3332)
         );
  MUX2_X1 U5374 ( .A(n4923), .B(DATAI_18_), .S(U3149), .Z(U3334) );
  MUX2_X1 U5375 ( .A(n5048), .B(DATAI_17_), .S(U3149), .Z(U3335) );
  MUX2_X1 U5376 ( .A(DATAI_15_), .B(n4924), .S(STATE_REG_SCAN_IN), .Z(U3337)
         );
  MUX2_X1 U5377 ( .A(DATAI_13_), .B(n5030), .S(STATE_REG_SCAN_IN), .Z(U3339)
         );
  MUX2_X1 U5378 ( .A(n5021), .B(DATAI_11_), .S(U3149), .Z(U3341) );
  MUX2_X1 U5379 ( .A(DATAI_9_), .B(n5010), .S(STATE_REG_SCAN_IN), .Z(U3343) );
  MUX2_X1 U5380 ( .A(n4999), .B(DATAI_8_), .S(U3149), .Z(U3344) );
  MUX2_X1 U5381 ( .A(n4979), .B(DATAI_5_), .S(U3149), .Z(U3347) );
  MUX2_X1 U5382 ( .A(DATAI_3_), .B(n4925), .S(STATE_REG_SCAN_IN), .Z(U3349) );
  MUX2_X1 U5383 ( .A(n4926), .B(DATAI_2_), .S(U3149), .Z(U3350) );
  MUX2_X1 U5384 ( .A(n2891), .B(DATAI_1_), .S(U3149), .Z(U3351) );
  MUX2_X1 U5385 ( .A(DATAI_0_), .B(IR_REG_0__SCAN_IN), .S(STATE_REG_SCAN_IN), 
        .Z(U3352) );
  INV_X2 U5386 ( .A(n4951), .ZN(n4953) );
  NOR2_X1 U5387 ( .A1(n4953), .A2(n4927), .ZN(U3320) );
  NOR2_X1 U5388 ( .A1(n4953), .A2(n4928), .ZN(U3319) );
  NOR2_X1 U5389 ( .A1(n4953), .A2(n4929), .ZN(U3318) );
  NOR2_X1 U5390 ( .A1(n4953), .A2(n4930), .ZN(U3317) );
  NOR2_X1 U5391 ( .A1(n4953), .A2(n4931), .ZN(U3316) );
  NOR2_X1 U5392 ( .A1(n4953), .A2(n4932), .ZN(U3315) );
  NOR2_X1 U5393 ( .A1(n4953), .A2(n4933), .ZN(U3314) );
  NOR2_X1 U5394 ( .A1(n4953), .A2(n4934), .ZN(U3313) );
  NOR2_X1 U5395 ( .A1(n4953), .A2(n4935), .ZN(U3312) );
  NOR2_X1 U5396 ( .A1(n4953), .A2(n4936), .ZN(U3311) );
  NOR2_X1 U5397 ( .A1(n4953), .A2(n4937), .ZN(U3310) );
  NOR2_X1 U5398 ( .A1(n4953), .A2(n4938), .ZN(U3309) );
  AND2_X1 U5399 ( .A1(n4951), .A2(D_REG_14__SCAN_IN), .ZN(U3308) );
  NOR2_X1 U5400 ( .A1(n4953), .A2(n4939), .ZN(U3307) );
  NOR2_X1 U5401 ( .A1(n4953), .A2(n4940), .ZN(U3306) );
  NOR2_X1 U5402 ( .A1(n4953), .A2(n4941), .ZN(U3305) );
  NOR2_X1 U5403 ( .A1(n4953), .A2(n4942), .ZN(U3304) );
  NOR2_X1 U5404 ( .A1(n4953), .A2(n4943), .ZN(U3303) );
  NOR2_X1 U5405 ( .A1(n4953), .A2(n4944), .ZN(U3302) );
  NOR2_X1 U5406 ( .A1(n4953), .A2(n4945), .ZN(U3301) );
  AND2_X1 U5407 ( .A1(n4951), .A2(D_REG_22__SCAN_IN), .ZN(U3300) );
  NOR2_X1 U5408 ( .A1(n4953), .A2(n4946), .ZN(U3299) );
  AND2_X1 U5409 ( .A1(n4951), .A2(D_REG_24__SCAN_IN), .ZN(U3298) );
  NOR2_X1 U5410 ( .A1(n4953), .A2(n4947), .ZN(U3297) );
  NOR2_X1 U5411 ( .A1(n4953), .A2(n4948), .ZN(U3296) );
  NOR2_X1 U5412 ( .A1(n4953), .A2(n4949), .ZN(U3295) );
  NOR2_X1 U5413 ( .A1(n4953), .A2(n4950), .ZN(U3294) );
  AND2_X1 U5414 ( .A1(n4951), .A2(D_REG_29__SCAN_IN), .ZN(U3293) );
  AND2_X1 U5415 ( .A1(n4951), .A2(D_REG_30__SCAN_IN), .ZN(U3292) );
  NOR2_X1 U5416 ( .A1(n4953), .A2(n4952), .ZN(U3291) );
  NAND2_X1 U5417 ( .A1(n4954), .A2(n2991), .ZN(n4955) );
  NAND2_X1 U5418 ( .A1(n5072), .A2(n4955), .ZN(n5079) );
  AOI21_X1 U5419 ( .B1(n5071), .B2(n5107), .A(n5079), .ZN(n4956) );
  XNOR2_X1 U5420 ( .A(n4956), .B(IR_REG_0__SCAN_IN), .ZN(n4959) );
  AOI22_X1 U5421 ( .A1(ADDR_REG_0__SCAN_IN), .A2(n5087), .B1(
        REG3_REG_0__SCAN_IN), .B2(U3149), .ZN(n4957) );
  OAI21_X1 U5422 ( .B1(n4959), .B2(n4958), .A(n4957), .ZN(U3240) );
  AOI22_X1 U5423 ( .A1(ADDR_REG_1__SCAN_IN), .A2(n5087), .B1(
        REG3_REG_1__SCAN_IN), .B2(U3149), .ZN(n4971) );
  AOI21_X1 U5424 ( .B1(n4961), .B2(n5075), .A(n4960), .ZN(n4962) );
  NAND2_X1 U5425 ( .A1(n5060), .A2(n4962), .ZN(n4968) );
  NAND2_X1 U5426 ( .A1(IR_REG_0__SCAN_IN), .A2(REG1_REG_0__SCAN_IN), .ZN(n4964) );
  AOI21_X1 U5427 ( .B1(n4965), .B2(n4964), .A(n4963), .ZN(n4966) );
  NAND2_X1 U5428 ( .A1(n5065), .A2(n4966), .ZN(n4967) );
  OAI211_X1 U5429 ( .C1(n5069), .C2(n2889), .A(n4968), .B(n4967), .ZN(n4969)
         );
  INV_X1 U5430 ( .A(n4969), .ZN(n4970) );
  NAND2_X1 U5431 ( .A1(n4971), .A2(n4970), .ZN(U3241) );
  AOI211_X1 U5432 ( .C1(n2558), .C2(n4973), .A(n4972), .B(n5088), .ZN(n4975)
         );
  AOI211_X1 U5433 ( .C1(n5087), .C2(ADDR_REG_5__SCAN_IN), .A(n4975), .B(n4974), 
        .ZN(n4981) );
  AOI211_X1 U5434 ( .C1(n2559), .C2(n4977), .A(n4976), .B(n5091), .ZN(n4978)
         );
  AOI21_X1 U5435 ( .B1(n5098), .B2(n4979), .A(n4978), .ZN(n4980) );
  NAND2_X1 U5436 ( .A1(n4981), .A2(n4980), .ZN(U3245) );
  AOI211_X1 U5437 ( .C1(n2557), .C2(n4983), .A(n4982), .B(n5091), .ZN(n4985)
         );
  AOI211_X1 U5438 ( .C1(n5087), .C2(ADDR_REG_7__SCAN_IN), .A(n4985), .B(n4984), 
        .ZN(n4991) );
  AOI211_X1 U5439 ( .C1(n4988), .C2(n4987), .A(n4986), .B(n5088), .ZN(n4989)
         );
  AOI21_X1 U5440 ( .B1(n5098), .B2(n5171), .A(n4989), .ZN(n4990) );
  NAND2_X1 U5441 ( .A1(n4991), .A2(n4990), .ZN(U3247) );
  NAND2_X1 U5442 ( .A1(ADDR_REG_8__SCAN_IN), .A2(n5087), .ZN(n5002) );
  AOI211_X1 U5443 ( .C1(n4993), .C2(n5205), .A(n4992), .B(n5088), .ZN(n4998)
         );
  AOI211_X1 U5444 ( .C1(n4996), .C2(n4995), .A(n4994), .B(n5091), .ZN(n4997)
         );
  AOI211_X1 U5445 ( .C1(n5098), .C2(n4999), .A(n4998), .B(n4997), .ZN(n5001)
         );
  NAND3_X1 U5446 ( .A1(n5002), .A2(n5001), .A3(n5000), .ZN(U3248) );
  NAND2_X1 U5447 ( .A1(ADDR_REG_9__SCAN_IN), .A2(n5087), .ZN(n5013) );
  AOI211_X1 U5448 ( .C1(n5005), .C2(n5004), .A(n5003), .B(n5091), .ZN(n5009)
         );
  AOI211_X1 U5449 ( .C1(n2553), .C2(n5007), .A(n5006), .B(n5088), .ZN(n5008)
         );
  AOI211_X1 U5450 ( .C1(n5098), .C2(n5010), .A(n5009), .B(n5008), .ZN(n5012)
         );
  NAND3_X1 U5451 ( .A1(n5013), .A2(n5012), .A3(n5011), .ZN(U3249) );
  AOI22_X1 U5452 ( .A1(REG3_REG_11__SCAN_IN), .A2(U3149), .B1(n5087), .B2(
        ADDR_REG_11__SCAN_IN), .ZN(n5023) );
  AOI211_X1 U5453 ( .C1(n2554), .C2(n5015), .A(n5014), .B(n5091), .ZN(n5020)
         );
  AOI211_X1 U5454 ( .C1(n5018), .C2(n5017), .A(n5016), .B(n5088), .ZN(n5019)
         );
  AOI211_X1 U5455 ( .C1(n5098), .C2(n5021), .A(n5020), .B(n5019), .ZN(n5022)
         );
  NAND2_X1 U5456 ( .A1(n5023), .A2(n5022), .ZN(U3251) );
  AOI211_X1 U5457 ( .C1(n5026), .C2(n5025), .A(n5088), .B(n5024), .ZN(n5028)
         );
  AOI211_X1 U5458 ( .C1(n5087), .C2(ADDR_REG_13__SCAN_IN), .A(n5028), .B(n5027), .ZN(n5034) );
  AOI21_X1 U5459 ( .B1(n2539), .B2(n5029), .A(n5091), .ZN(n5032) );
  AOI22_X1 U5460 ( .A1(n5032), .A2(n5031), .B1(n5030), .B2(n5098), .ZN(n5033)
         );
  NAND2_X1 U5461 ( .A1(n5034), .A2(n5033), .ZN(U3253) );
  NAND2_X1 U5462 ( .A1(ADDR_REG_14__SCAN_IN), .A2(n5087), .ZN(n5045) );
  AOI211_X1 U5463 ( .C1(n5037), .C2(n5036), .A(n5035), .B(n5091), .ZN(n5041)
         );
  AOI211_X1 U5464 ( .C1(n5300), .C2(n5039), .A(n5088), .B(n5038), .ZN(n5040)
         );
  AOI211_X1 U5465 ( .C1(n5098), .C2(n5042), .A(n5041), .B(n5040), .ZN(n5044)
         );
  NAND3_X1 U5466 ( .A1(n5045), .A2(n5044), .A3(n5043), .ZN(U3254) );
  XNOR2_X1 U5467 ( .A(n5047), .B(n5046), .ZN(n5049) );
  AOI22_X1 U5468 ( .A1(n5049), .A2(n5065), .B1(n5048), .B2(n5098), .ZN(n5055)
         );
  AOI211_X1 U5469 ( .C1(n5051), .C2(n5050), .A(n2524), .B(n5091), .ZN(n5052)
         );
  AOI211_X1 U5470 ( .C1(n5087), .C2(ADDR_REG_17__SCAN_IN), .A(n5053), .B(n5052), .ZN(n5054) );
  NAND2_X1 U5471 ( .A1(n5055), .A2(n5054), .ZN(U3257) );
  AOI22_X1 U5472 ( .A1(ADDR_REG_2__SCAN_IN), .A2(n5087), .B1(
        REG3_REG_2__SCAN_IN), .B2(U3149), .ZN(n5085) );
  AOI21_X1 U5473 ( .B1(n5058), .B2(n5057), .A(n5056), .ZN(n5059) );
  NAND2_X1 U5474 ( .A1(n5060), .A2(n5059), .ZN(n5067) );
  AOI21_X1 U5475 ( .B1(n5063), .B2(n5062), .A(n5061), .ZN(n5064) );
  NAND2_X1 U5476 ( .A1(n5065), .A2(n5064), .ZN(n5066) );
  OAI211_X1 U5477 ( .C1(n5069), .C2(n5068), .A(n5067), .B(n5066), .ZN(n5070)
         );
  INV_X1 U5478 ( .A(n5070), .ZN(n5084) );
  NAND3_X1 U5479 ( .A1(n5073), .A2(n5072), .A3(n5071), .ZN(n5083) );
  INV_X1 U5480 ( .A(n5074), .ZN(n5077) );
  INV_X1 U5481 ( .A(n5075), .ZN(n5076) );
  NAND2_X1 U5482 ( .A1(n5077), .A2(n5076), .ZN(n5081) );
  NAND2_X1 U5483 ( .A1(n5079), .A2(n5078), .ZN(n5080) );
  NAND4_X1 U5484 ( .A1(n5083), .A2(n5082), .A3(n5081), .A4(n5080), .ZN(n5099)
         );
  NAND3_X1 U5485 ( .A1(n5085), .A2(n5084), .A3(n5099), .ZN(U3242) );
  AOI21_X1 U5486 ( .B1(n5087), .B2(ADDR_REG_4__SCAN_IN), .A(n5086), .ZN(n5101)
         );
  AOI211_X1 U5487 ( .C1(n5090), .C2(n5158), .A(n5089), .B(n5088), .ZN(n5096)
         );
  AOI211_X1 U5488 ( .C1(n5094), .C2(n5093), .A(n5092), .B(n5091), .ZN(n5095)
         );
  AOI211_X1 U5489 ( .C1(n5098), .C2(n5097), .A(n5096), .B(n5095), .ZN(n5100)
         );
  NAND3_X1 U5490 ( .A1(n5101), .A2(n5100), .A3(n5099), .ZN(U3244) );
  INV_X2 U5491 ( .A(n5379), .ZN(n5363) );
  INV_X1 U5492 ( .A(n5122), .ZN(n5143) );
  NAND2_X1 U5493 ( .A1(n5102), .A2(n5138), .ZN(n5104) );
  AOI22_X1 U5494 ( .A1(n5114), .A2(n5104), .B1(n5136), .B2(n5103), .ZN(n5110)
         );
  OAI21_X1 U5495 ( .B1(n5106), .B2(n5105), .A(n5110), .ZN(n5111) );
  AOI21_X1 U5496 ( .B1(n5143), .B2(n5114), .A(n5111), .ZN(n5109) );
  AOI22_X1 U5497 ( .A1(n5363), .A2(n5109), .B1(n5107), .B2(n5379), .ZN(U3518)
         );
  AOI22_X1 U5498 ( .A1(n2512), .A2(n5109), .B1(n5108), .B2(n5380), .ZN(U3467)
         );
  INV_X1 U5499 ( .A(n5110), .ZN(n5113) );
  OAI21_X1 U5500 ( .B1(n5113), .B2(n5112), .A(n5111), .ZN(n5116) );
  AOI22_X1 U5501 ( .A1(n5114), .A2(n5279), .B1(REG3_REG_0__SCAN_IN), .B2(n5276), .ZN(n5115) );
  OAI221_X1 U5502 ( .B1(n5374), .B2(n5116), .C1(n5226), .C2(n2991), .A(n5115), 
        .ZN(U3290) );
  INV_X1 U5503 ( .A(n5117), .ZN(n5120) );
  AOI211_X1 U5504 ( .C1(n5120), .C2(n5143), .A(n5119), .B(n5118), .ZN(n5121)
         );
  AOI22_X1 U5505 ( .A1(n5363), .A2(n5121), .B1(n2776), .B2(n5379), .ZN(U3519)
         );
  AOI22_X1 U5506 ( .A1(n2512), .A2(n5121), .B1(n4894), .B2(n5380), .ZN(U3469)
         );
  NOR2_X1 U5507 ( .A1(n5123), .A2(n5122), .ZN(n5125) );
  AOI211_X1 U5508 ( .C1(n5377), .C2(n5126), .A(n5125), .B(n5124), .ZN(n5127)
         );
  AOI22_X1 U5509 ( .A1(n5363), .A2(n5127), .B1(n3055), .B2(n5379), .ZN(U3520)
         );
  AOI22_X1 U5510 ( .A1(n2512), .A2(n5127), .B1(n4701), .B2(n5380), .ZN(U3471)
         );
  XOR2_X1 U5511 ( .A(n5128), .B(n5131), .Z(n5149) );
  NOR2_X1 U5512 ( .A1(n5147), .A2(n5333), .ZN(n5142) );
  XOR2_X1 U5513 ( .A(n5131), .B(n5130), .Z(n5139) );
  OAI22_X1 U5514 ( .A1(n5133), .A2(n5246), .B1(n5266), .B2(n5132), .ZN(n5134)
         );
  AOI21_X1 U5515 ( .B1(n5136), .B2(n5135), .A(n5134), .ZN(n5137) );
  OAI21_X1 U5516 ( .B1(n5139), .B2(n5138), .A(n5137), .ZN(n5140) );
  AOI21_X1 U5517 ( .B1(n5274), .B2(n5149), .A(n5140), .ZN(n5152) );
  INV_X1 U5518 ( .A(n5152), .ZN(n5141) );
  AOI211_X1 U5519 ( .C1(n5143), .C2(n5149), .A(n5142), .B(n5141), .ZN(n5145)
         );
  AOI22_X1 U5520 ( .A1(n5363), .A2(n5145), .B1(n5144), .B2(n5379), .ZN(U3521)
         );
  AOI22_X1 U5521 ( .A1(n2512), .A2(n5145), .B1(n4899), .B2(n5380), .ZN(U3473)
         );
  AOI22_X1 U5522 ( .A1(n5374), .A2(REG2_REG_3__SCAN_IN), .B1(n5276), .B2(n5146), .ZN(n5151) );
  INV_X1 U5523 ( .A(n5147), .ZN(n5148) );
  AOI22_X1 U5524 ( .A1(n5149), .A2(n5279), .B1(n5372), .B2(n5148), .ZN(n5150)
         );
  OAI211_X1 U5525 ( .C1(n5374), .C2(n5152), .A(n5151), .B(n5150), .ZN(U3287)
         );
  AOI22_X1 U5526 ( .A1(STATE_REG_SCAN_IN), .A2(n5154), .B1(n5153), .B2(U3149), 
        .ZN(U3348) );
  AOI211_X1 U5527 ( .C1(n5157), .C2(n5335), .A(n5156), .B(n5155), .ZN(n5159)
         );
  AOI22_X1 U5528 ( .A1(n5363), .A2(n5159), .B1(n5158), .B2(n5379), .ZN(U3522)
         );
  AOI22_X1 U5529 ( .A1(n2512), .A2(n5159), .B1(n4898), .B2(n5380), .ZN(U3475)
         );
  OAI22_X1 U5530 ( .A1(n5379), .A2(n5160), .B1(REG1_REG_5__SCAN_IN), .B2(n5363), .ZN(n5161) );
  INV_X1 U5531 ( .A(n5161), .ZN(U3523) );
  AOI22_X1 U5532 ( .A1(STATE_REG_SCAN_IN), .A2(n5163), .B1(n5162), .B2(U3149), 
        .ZN(U3346) );
  NOR2_X1 U5533 ( .A1(n5164), .A2(n5333), .ZN(n5166) );
  AOI211_X1 U5534 ( .C1(n5167), .C2(n5335), .A(n5166), .B(n5165), .ZN(n5170)
         );
  AOI22_X1 U5535 ( .A1(n5363), .A2(n5170), .B1(n5168), .B2(n5379), .ZN(U3524)
         );
  AOI22_X1 U5536 ( .A1(n2512), .A2(n5170), .B1(n5169), .B2(n5380), .ZN(U3479)
         );
  OAI22_X1 U5537 ( .A1(U3149), .A2(n5171), .B1(DATAI_7_), .B2(
        STATE_REG_SCAN_IN), .ZN(n5172) );
  INV_X1 U5538 ( .A(n5172), .ZN(U3345) );
  INV_X1 U5539 ( .A(REG2_REG_7__SCAN_IN), .ZN(n5194) );
  NAND2_X1 U5540 ( .A1(n5173), .A2(n5174), .ZN(n5175) );
  NAND2_X1 U5541 ( .A1(n5176), .A2(n5175), .ZN(n5197) );
  INV_X1 U5542 ( .A(n5177), .ZN(n5224) );
  XNOR2_X1 U5543 ( .A(n5178), .B(n3393), .ZN(n5185) );
  AOI22_X1 U5544 ( .A1(n5181), .A2(n5180), .B1(n5365), .B2(n5179), .ZN(n5182)
         );
  OAI21_X1 U5545 ( .B1(n5183), .B2(n5244), .A(n5182), .ZN(n5184) );
  AOI21_X1 U5546 ( .B1(n5185), .B2(n5268), .A(n5184), .ZN(n5196) );
  OAI211_X1 U5547 ( .C1(n5188), .C2(n5187), .A(n5377), .B(n5186), .ZN(n5195)
         );
  OAI22_X1 U5548 ( .A1(n5195), .A2(n2846), .B1(n5189), .B2(n5231), .ZN(n5190)
         );
  INV_X1 U5549 ( .A(n5190), .ZN(n5191) );
  OAI211_X1 U5550 ( .C1(n5197), .C2(n5224), .A(n5196), .B(n5191), .ZN(n5192)
         );
  INV_X1 U5551 ( .A(n5192), .ZN(n5193) );
  AOI22_X1 U5552 ( .A1(n5374), .A2(n5194), .B1(n5193), .B2(n5226), .ZN(U3283)
         );
  OAI211_X1 U5553 ( .C1(n5197), .C2(n5296), .A(n5196), .B(n5195), .ZN(n5198)
         );
  INV_X1 U5554 ( .A(n5198), .ZN(n5200) );
  AOI22_X1 U5555 ( .A1(n5363), .A2(n5200), .B1(n3170), .B2(n5379), .ZN(U3525)
         );
  AOI22_X1 U5556 ( .A1(n2512), .A2(n5200), .B1(n5199), .B2(n5380), .ZN(U3481)
         );
  OAI21_X1 U5557 ( .B1(n5333), .B2(n5202), .A(n5201), .ZN(n5203) );
  AOI21_X1 U5558 ( .B1(n5204), .B2(n5335), .A(n5203), .ZN(n5206) );
  AOI22_X1 U5559 ( .A1(n5363), .A2(n5206), .B1(n5205), .B2(n5379), .ZN(U3526)
         );
  AOI22_X1 U5560 ( .A1(n2512), .A2(n5206), .B1(n4709), .B2(n5380), .ZN(U3483)
         );
  XNOR2_X1 U5561 ( .A(n5207), .B(n5212), .ZN(n5222) );
  NAND2_X1 U5562 ( .A1(n5209), .A2(n5208), .ZN(n5210) );
  NAND2_X1 U5563 ( .A1(n5211), .A2(n5210), .ZN(n5220) );
  XNOR2_X1 U5564 ( .A(n5213), .B(n5212), .ZN(n5217) );
  OAI21_X1 U5565 ( .B1(n5266), .B2(n5215), .A(n5214), .ZN(n5216) );
  AOI21_X1 U5566 ( .B1(n5217), .B2(n5268), .A(n5216), .ZN(n5223) );
  OAI21_X1 U5567 ( .B1(n5333), .B2(n5220), .A(n5223), .ZN(n5218) );
  AOI21_X1 U5568 ( .B1(n5335), .B2(n5222), .A(n5218), .ZN(n5219) );
  AOI22_X1 U5569 ( .A1(n5363), .A2(n5219), .B1(n3330), .B2(n5379), .ZN(U3527)
         );
  AOI22_X1 U5570 ( .A1(n2512), .A2(n5219), .B1(n3331), .B2(n5380), .ZN(U3485)
         );
  INV_X1 U5571 ( .A(n5220), .ZN(n5221) );
  AOI22_X1 U5572 ( .A1(n5221), .A2(n5372), .B1(REG2_REG_9__SCAN_IN), .B2(n5374), .ZN(n5229) );
  INV_X1 U5573 ( .A(n5222), .ZN(n5225) );
  OAI21_X1 U5574 ( .B1(n5225), .B2(n5224), .A(n5223), .ZN(n5227) );
  NAND2_X1 U5575 ( .A1(n5227), .A2(n5226), .ZN(n5228) );
  OAI211_X1 U5576 ( .C1(n5231), .C2(n5230), .A(n5229), .B(n5228), .ZN(U3281)
         );
  NOR3_X1 U5577 ( .A1(n5233), .A2(n5232), .A3(n5296), .ZN(n5234) );
  AOI211_X1 U5578 ( .C1(n5377), .C2(n5236), .A(n5235), .B(n5234), .ZN(n5238)
         );
  AOI22_X1 U5579 ( .A1(n5363), .A2(n5238), .B1(n5237), .B2(n5379), .ZN(U3528)
         );
  AOI22_X1 U5580 ( .A1(n2512), .A2(n5238), .B1(n3365), .B2(n5380), .ZN(U3487)
         );
  AOI22_X1 U5581 ( .A1(n5339), .A2(n5260), .B1(REG3_REG_11__SCAN_IN), .B2(
        U3149), .ZN(n5253) );
  INV_X1 U5582 ( .A(n5239), .ZN(n5240) );
  NOR2_X1 U5583 ( .A1(n5241), .A2(n5240), .ZN(n5242) );
  XNOR2_X1 U5584 ( .A(n5243), .B(n5242), .ZN(n5251) );
  OR2_X1 U5585 ( .A1(n5245), .A2(n5244), .ZN(n5249) );
  OR2_X1 U5586 ( .A1(n5247), .A2(n5246), .ZN(n5248) );
  AND2_X1 U5587 ( .A1(n5249), .A2(n5248), .ZN(n5264) );
  INV_X1 U5588 ( .A(n5264), .ZN(n5250) );
  AOI22_X1 U5589 ( .A1(n5251), .A2(n5314), .B1(n5348), .B2(n5250), .ZN(n5252)
         );
  OAI211_X1 U5590 ( .C1(n5354), .C2(n5275), .A(n5253), .B(n5252), .ZN(U3233)
         );
  AOI21_X1 U5591 ( .B1(n5261), .B2(n5255), .A(n5254), .ZN(n5256) );
  INV_X1 U5592 ( .A(n5256), .ZN(n5280) );
  INV_X1 U5593 ( .A(n5257), .ZN(n5259) );
  AOI21_X1 U5594 ( .B1(n5260), .B2(n5259), .A(n5258), .ZN(n5278) );
  AOI22_X1 U5595 ( .A1(n5280), .A2(n5335), .B1(n5377), .B2(n5278), .ZN(n5270)
         );
  INV_X1 U5596 ( .A(n5261), .ZN(n5262) );
  XNOR2_X1 U5597 ( .A(n5263), .B(n5262), .ZN(n5269) );
  OAI21_X1 U5598 ( .B1(n5266), .B2(n5265), .A(n5264), .ZN(n5267) );
  AOI21_X1 U5599 ( .B1(n5269), .B2(n5268), .A(n5267), .ZN(n5272) );
  AOI22_X1 U5600 ( .A1(n5363), .A2(n5271), .B1(n3415), .B2(n5379), .ZN(U3529)
         );
  AOI22_X1 U5601 ( .A1(n2512), .A2(n5271), .B1(n3414), .B2(n5380), .ZN(U3489)
         );
  INV_X1 U5602 ( .A(n5272), .ZN(n5273) );
  AOI21_X1 U5603 ( .B1(n5280), .B2(n5274), .A(n5273), .ZN(n5283) );
  INV_X1 U5604 ( .A(n5275), .ZN(n5277) );
  AOI22_X1 U5605 ( .A1(n5277), .A2(n5276), .B1(REG2_REG_11__SCAN_IN), .B2(
        n5374), .ZN(n5282) );
  AOI22_X1 U5606 ( .A1(n5280), .A2(n5279), .B1(n5372), .B2(n5278), .ZN(n5281)
         );
  OAI211_X1 U5607 ( .C1(n5374), .C2(n5283), .A(n5282), .B(n5281), .ZN(U3279)
         );
  OAI21_X1 U5608 ( .B1(n5333), .B2(n5285), .A(n5284), .ZN(n5286) );
  AOI21_X1 U5609 ( .B1(n5287), .B2(n5335), .A(n5286), .ZN(n5289) );
  AOI22_X1 U5610 ( .A1(n5363), .A2(n5289), .B1(n5288), .B2(n5379), .ZN(U3530)
         );
  AOI22_X1 U5611 ( .A1(n2512), .A2(n5289), .B1(n3434), .B2(n5380), .ZN(U3491)
         );
  AOI211_X1 U5612 ( .C1(n5292), .C2(n5335), .A(n5291), .B(n5290), .ZN(n5293)
         );
  AOI22_X1 U5613 ( .A1(n5363), .A2(n5293), .B1(n3448), .B2(n5379), .ZN(U3531)
         );
  AOI22_X1 U5614 ( .A1(n2512), .A2(n5293), .B1(n3452), .B2(n5380), .ZN(U3493)
         );
  INV_X1 U5615 ( .A(n5294), .ZN(n5295) );
  OAI22_X1 U5616 ( .A1(n5297), .A2(n5296), .B1(n5333), .B2(n5295), .ZN(n5298)
         );
  NOR2_X1 U5617 ( .A1(n5299), .A2(n5298), .ZN(n5301) );
  AOI22_X1 U5618 ( .A1(n5363), .A2(n5301), .B1(n5300), .B2(n5379), .ZN(U3532)
         );
  AOI22_X1 U5619 ( .A1(n2512), .A2(n5301), .B1(n3524), .B2(n5380), .ZN(U3495)
         );
  OAI22_X1 U5620 ( .A1(n5305), .A2(n5304), .B1(n5303), .B2(n5302), .ZN(n5306)
         );
  AOI211_X1 U5621 ( .C1(n5309), .C2(n5308), .A(n5307), .B(n5306), .ZN(n5317)
         );
  NAND2_X1 U5622 ( .A1(n5311), .A2(n5310), .ZN(n5313) );
  XNOR2_X1 U5623 ( .A(n5313), .B(n5312), .ZN(n5315) );
  NAND2_X1 U5624 ( .A1(n5315), .A2(n5314), .ZN(n5316) );
  OAI211_X1 U5625 ( .C1(n5354), .C2(n5318), .A(n5317), .B(n5316), .ZN(U3238)
         );
  NOR3_X1 U5626 ( .A1(n5320), .A2(n5319), .A3(n5333), .ZN(n5322) );
  AOI211_X1 U5627 ( .C1(n5323), .C2(n5335), .A(n5322), .B(n5321), .ZN(n5325)
         );
  AOI22_X1 U5628 ( .A1(n5363), .A2(n5325), .B1(n5324), .B2(n5379), .ZN(U3533)
         );
  AOI22_X1 U5629 ( .A1(n2512), .A2(n5325), .B1(n3564), .B2(n5380), .ZN(U3497)
         );
  AOI211_X1 U5630 ( .C1(n5328), .C2(n5335), .A(n5327), .B(n5326), .ZN(n5330)
         );
  AOI22_X1 U5631 ( .A1(n5363), .A2(n5330), .B1(n5329), .B2(n5379), .ZN(U3534)
         );
  AOI22_X1 U5632 ( .A1(n2512), .A2(n5330), .B1(n3577), .B2(n5380), .ZN(U3499)
         );
  OAI21_X1 U5633 ( .B1(n5333), .B2(n5332), .A(n5331), .ZN(n5334) );
  AOI21_X1 U5634 ( .B1(n5336), .B2(n5335), .A(n5334), .ZN(n5337) );
  AOI22_X1 U5635 ( .A1(n5363), .A2(n5337), .B1(n3587), .B2(n5379), .ZN(U3535)
         );
  AOI22_X1 U5636 ( .A1(n2512), .A2(n5337), .B1(n3583), .B2(n5380), .ZN(U3501)
         );
  AOI22_X1 U5637 ( .A1(n5339), .A2(n5338), .B1(REG3_REG_18__SCAN_IN), .B2(
        U3149), .ZN(n5352) );
  AND2_X1 U5638 ( .A1(n5343), .A2(n5340), .ZN(n5342) );
  OAI21_X1 U5639 ( .B1(n5342), .B2(n5346), .A(n5341), .ZN(n5350) );
  INV_X1 U5640 ( .A(n5343), .ZN(n5345) );
  AOI21_X1 U5641 ( .B1(n5346), .B2(n5345), .A(n5344), .ZN(n5349) );
  AOI22_X1 U5642 ( .A1(n5350), .A2(n5349), .B1(n5348), .B2(n5347), .ZN(n5351)
         );
  OAI211_X1 U5643 ( .C1(n5354), .C2(n5353), .A(n5352), .B(n5351), .ZN(U3235)
         );
  NAND2_X1 U5644 ( .A1(n5356), .A2(n5355), .ZN(n5368) );
  INV_X1 U5645 ( .A(n5358), .ZN(n5369) );
  NAND2_X1 U5646 ( .A1(n5369), .A2(n5365), .ZN(n5357) );
  AND2_X1 U5647 ( .A1(n5368), .A2(n5357), .ZN(n5360) );
  XNOR2_X1 U5648 ( .A(n5370), .B(n5358), .ZN(n5362) );
  AOI22_X1 U5649 ( .A1(n5362), .A2(n5372), .B1(REG2_REG_30__SCAN_IN), .B2(
        n5374), .ZN(n5359) );
  OAI21_X1 U5650 ( .B1(n5374), .B2(n5360), .A(n5359), .ZN(U3261) );
  INV_X1 U5651 ( .A(n5360), .ZN(n5361) );
  AOI21_X1 U5652 ( .B1(n5362), .B2(n5377), .A(n5361), .ZN(n5364) );
  AOI22_X1 U5653 ( .A1(n5363), .A2(n5364), .B1(n4060), .B2(n5379), .ZN(U3548)
         );
  AOI22_X1 U5654 ( .A1(n2512), .A2(n5364), .B1(n4057), .B2(n5380), .ZN(U3516)
         );
  INV_X1 U5655 ( .A(n5371), .ZN(n5366) );
  NAND2_X1 U5656 ( .A1(n5366), .A2(n5365), .ZN(n5367) );
  AND2_X1 U5657 ( .A1(n5368), .A2(n5367), .ZN(n5375) );
  AOI22_X1 U5658 ( .A1(n5378), .A2(n5372), .B1(n5374), .B2(
        REG2_REG_31__SCAN_IN), .ZN(n5373) );
  OAI21_X1 U5659 ( .B1(n5374), .B2(n5375), .A(n5373), .ZN(U3260) );
  INV_X1 U5660 ( .A(n5375), .ZN(n5376) );
  AOI22_X1 U5661 ( .A1(n2512), .A2(n5381), .B1(n4053), .B2(n5380), .ZN(U3517)
         );
  CLKBUF_X3 U2551 ( .A(n3814), .Z(n2511) );
endmodule

