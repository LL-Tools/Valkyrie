

module b22_C_gen_AntiSAT_k_256_7 ( P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN, 
        P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN, 
        P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN, 
        P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN, 
        P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN, 
        P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN, 
        P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN, 
        P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN, 
        P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN, 
        P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN, P3_REG3_REG_0__SCAN_IN, 
        P3_REG3_REG_20__SCAN_IN, P3_REG3_REG_13__SCAN_IN, 
        P3_REG3_REG_22__SCAN_IN, P3_REG3_REG_11__SCAN_IN, 
        P3_REG3_REG_2__SCAN_IN, P3_REG3_REG_18__SCAN_IN, 
        P3_REG3_REG_6__SCAN_IN, P3_REG3_REG_26__SCAN_IN, 
        P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_ADDR_REG_0__SCAN_IN, 
        P3_ADDR_REG_1__SCAN_IN, P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN, 
        P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN, P3_ADDR_REG_6__SCAN_IN, 
        P3_ADDR_REG_7__SCAN_IN, P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, 
        P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, 
        P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, 
        P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, 
        P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, 
        P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, 
        P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, 
        P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, 
        P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, 
        P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, 
        P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, 
        P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, 
        P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, 
        P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, 
        P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, 
        P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, 
        P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, 
        P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, 
        P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, 
        P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, 
        P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, 
        P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, 
        P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, 
        P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, 
        P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, 
        P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, 
        P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN, 
        P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN, 
        P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN, 
        P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN, 
        P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN, 
        P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN, 
        P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN, 
        P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN, 
        P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN, 
        P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN, 
        P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN, 
        P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN, 
        P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN, 
        P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN, 
        P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN, 
        P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN, 
        P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN, 
        P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_4__SCAN_IN, 
        P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_17__SCAN_IN, 
        P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_16__SCAN_IN, 
        P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_12__SCAN_IN, 
        P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_1__SCAN_IN, 
        P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_28__SCAN_IN, 
        P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_3__SCAN_IN, 
        P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_23__SCAN_IN, 
        P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_27__SCAN_IN, 
        P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN, P2_RD_REG_SCAN_IN, 
        P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN, P3_IR_REG_1__SCAN_IN, 
        P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN, P3_IR_REG_4__SCAN_IN, 
        P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN, P3_IR_REG_7__SCAN_IN, 
        P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN, P3_IR_REG_10__SCAN_IN, 
        P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN, P3_IR_REG_13__SCAN_IN, 
        P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN, P3_IR_REG_16__SCAN_IN, 
        P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN, P3_IR_REG_19__SCAN_IN, 
        P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN, P3_IR_REG_22__SCAN_IN, 
        P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN, P3_IR_REG_25__SCAN_IN, 
        P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN, P3_IR_REG_28__SCAN_IN, 
        P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN, P3_IR_REG_31__SCAN_IN, 
        P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN, P3_D_REG_2__SCAN_IN, 
        P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN, P3_D_REG_5__SCAN_IN, 
        P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN, P3_D_REG_8__SCAN_IN, 
        P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN, P3_D_REG_11__SCAN_IN, 
        P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN, P3_D_REG_14__SCAN_IN, 
        P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN, P3_D_REG_17__SCAN_IN, 
        P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN, P3_D_REG_20__SCAN_IN, 
        P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN, P3_D_REG_23__SCAN_IN, 
        P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN, P3_D_REG_26__SCAN_IN, 
        P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN, P3_D_REG_29__SCAN_IN, 
        P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN, P3_REG0_REG_0__SCAN_IN, 
        P3_REG0_REG_1__SCAN_IN, P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN, 
        P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN, P3_REG0_REG_6__SCAN_IN, 
        P3_REG0_REG_7__SCAN_IN, P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN, 
        P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN, 
        P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN, 
        P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN, 
        P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN, 
        P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN, 
        P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN, 
        P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN, 
        P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN, 
        P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN, 
        P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN, 
        P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN, 
        P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN, P3_REG1_REG_2__SCAN_IN, 
        P3_REG1_REG_3__SCAN_IN, P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN, 
        P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN, P3_REG1_REG_8__SCAN_IN, 
        P3_REG1_REG_9__SCAN_IN, P3_REG1_REG_10__SCAN_IN, 
        P3_REG1_REG_11__SCAN_IN, P3_REG1_REG_12__SCAN_IN, 
        P3_REG1_REG_13__SCAN_IN, P3_REG1_REG_14__SCAN_IN, 
        P3_REG1_REG_15__SCAN_IN, P3_REG1_REG_16__SCAN_IN, 
        P3_REG1_REG_17__SCAN_IN, P3_REG1_REG_18__SCAN_IN, 
        P3_REG1_REG_19__SCAN_IN, P3_REG1_REG_20__SCAN_IN, 
        P3_REG1_REG_21__SCAN_IN, P3_REG1_REG_22__SCAN_IN, 
        P3_REG1_REG_23__SCAN_IN, P3_REG1_REG_24__SCAN_IN, 
        P3_REG1_REG_25__SCAN_IN, P3_REG1_REG_26__SCAN_IN, 
        P3_REG1_REG_27__SCAN_IN, P3_REG1_REG_28__SCAN_IN, 
        P3_REG1_REG_29__SCAN_IN, P3_REG1_REG_30__SCAN_IN, 
        P3_REG1_REG_31__SCAN_IN, P3_REG2_REG_0__SCAN_IN, 
        P3_REG2_REG_1__SCAN_IN, P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN, 
        P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN, P3_REG2_REG_6__SCAN_IN, 
        P3_REG2_REG_7__SCAN_IN, P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN, 
        P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN, 
        P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN, 
        P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN, 
        P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN, 
        P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN, 
        P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN, 
        P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN, 
        P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN, 
        P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN, 
        P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN, 
        P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN, 
        P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN, 
        P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN, 
        P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN, 
        P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN, 
        P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, keyinput_f0, 
        keyinput_f1, keyinput_f2, keyinput_f3, keyinput_f4, keyinput_f5, 
        keyinput_f6, keyinput_f7, keyinput_f8, keyinput_f9, keyinput_f10, 
        keyinput_f11, keyinput_f12, keyinput_f13, keyinput_f14, keyinput_f15, 
        keyinput_f16, keyinput_f17, keyinput_f18, keyinput_f19, keyinput_f20, 
        keyinput_f21, keyinput_f22, keyinput_f23, keyinput_f24, keyinput_f25, 
        keyinput_f26, keyinput_f27, keyinput_f28, keyinput_f29, keyinput_f30, 
        keyinput_f31, keyinput_f32, keyinput_f33, keyinput_f34, keyinput_f35, 
        keyinput_f36, keyinput_f37, keyinput_f38, keyinput_f39, keyinput_f40, 
        keyinput_f41, keyinput_f42, keyinput_f43, keyinput_f44, keyinput_f45, 
        keyinput_f46, keyinput_f47, keyinput_f48, keyinput_f49, keyinput_f50, 
        keyinput_f51, keyinput_f52, keyinput_f53, keyinput_f54, keyinput_f55, 
        keyinput_f56, keyinput_f57, keyinput_f58, keyinput_f59, keyinput_f60, 
        keyinput_f61, keyinput_f62, keyinput_f63, keyinput_f64, keyinput_f65, 
        keyinput_f66, keyinput_f67, keyinput_f68, keyinput_f69, keyinput_f70, 
        keyinput_f71, keyinput_f72, keyinput_f73, keyinput_f74, keyinput_f75, 
        keyinput_f76, keyinput_f77, keyinput_f78, keyinput_f79, keyinput_f80, 
        keyinput_f81, keyinput_f82, keyinput_f83, keyinput_f84, keyinput_f85, 
        keyinput_f86, keyinput_f87, keyinput_f88, keyinput_f89, keyinput_f90, 
        keyinput_f91, keyinput_f92, keyinput_f93, keyinput_f94, keyinput_f95, 
        keyinput_f96, keyinput_f97, keyinput_f98, keyinput_f99, keyinput_f100, 
        keyinput_f101, keyinput_f102, keyinput_f103, keyinput_f104, 
        keyinput_f105, keyinput_f106, keyinput_f107, keyinput_f108, 
        keyinput_f109, keyinput_f110, keyinput_f111, keyinput_f112, 
        keyinput_f113, keyinput_f114, keyinput_f115, keyinput_f116, 
        keyinput_f117, keyinput_f118, keyinput_f119, keyinput_f120, 
        keyinput_f121, keyinput_f122, keyinput_f123, keyinput_f124, 
        keyinput_f125, keyinput_f126, keyinput_f127, keyinput_g0, keyinput_g1, 
        keyinput_g2, keyinput_g3, keyinput_g4, keyinput_g5, keyinput_g6, 
        keyinput_g7, keyinput_g8, keyinput_g9, keyinput_g10, keyinput_g11, 
        keyinput_g12, keyinput_g13, keyinput_g14, keyinput_g15, keyinput_g16, 
        keyinput_g17, keyinput_g18, keyinput_g19, keyinput_g20, keyinput_g21, 
        keyinput_g22, keyinput_g23, keyinput_g24, keyinput_g25, keyinput_g26, 
        keyinput_g27, keyinput_g28, keyinput_g29, keyinput_g30, keyinput_g31, 
        keyinput_g32, keyinput_g33, keyinput_g34, keyinput_g35, keyinput_g36, 
        keyinput_g37, keyinput_g38, keyinput_g39, keyinput_g40, keyinput_g41, 
        keyinput_g42, keyinput_g43, keyinput_g44, keyinput_g45, keyinput_g46, 
        keyinput_g47, keyinput_g48, keyinput_g49, keyinput_g50, keyinput_g51, 
        keyinput_g52, keyinput_g53, keyinput_g54, keyinput_g55, keyinput_g56, 
        keyinput_g57, keyinput_g58, keyinput_g59, keyinput_g60, keyinput_g61, 
        keyinput_g62, keyinput_g63, keyinput_g64, keyinput_g65, keyinput_g66, 
        keyinput_g67, keyinput_g68, keyinput_g69, keyinput_g70, keyinput_g71, 
        keyinput_g72, keyinput_g73, keyinput_g74, keyinput_g75, keyinput_g76, 
        keyinput_g77, keyinput_g78, keyinput_g79, keyinput_g80, keyinput_g81, 
        keyinput_g82, keyinput_g83, keyinput_g84, keyinput_g85, keyinput_g86, 
        keyinput_g87, keyinput_g88, keyinput_g89, keyinput_g90, keyinput_g91, 
        keyinput_g92, keyinput_g93, keyinput_g94, keyinput_g95, keyinput_g96, 
        keyinput_g97, keyinput_g98, keyinput_g99, keyinput_g100, keyinput_g101, 
        keyinput_g102, keyinput_g103, keyinput_g104, keyinput_g105, 
        keyinput_g106, keyinput_g107, keyinput_g108, keyinput_g109, 
        keyinput_g110, keyinput_g111, keyinput_g112, keyinput_g113, 
        keyinput_g114, keyinput_g115, keyinput_g116, keyinput_g117, 
        keyinput_g118, keyinput_g119, keyinput_g120, keyinput_g121, 
        keyinput_g122, keyinput_g123, keyinput_g124, keyinput_g125, 
        keyinput_g126, keyinput_g127, SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, 
        SUB_1596_U64, SUB_1596_U65, SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, 
        SUB_1596_U69, SUB_1596_U70, SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, 
        SUB_1596_U57, SUB_1596_U58, SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, 
        SUB_1596_U5, SUB_1596_U53, U29, U28, P1_U3355, P1_U3354, P1_U3353, 
        P1_U3352, P1_U3351, P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, 
        P1_U3345, P1_U3344, P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, 
        P1_U3338, P1_U3337, P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, 
        P1_U3331, P1_U3330, P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, 
        P1_U3324, P1_U3445, P1_U3446, P1_U3323, P1_U3322, P1_U3321, P1_U3320, 
        P1_U3319, P1_U3318, P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, 
        P1_U3312, P1_U3311, P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, 
        P1_U3305, P1_U3304, P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, 
        P1_U3298, P1_U3297, P1_U3296, P1_U3295, P1_U3294, P1_U3459, P1_U3462, 
        P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483, 
        P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504, 
        P1_U3507, P1_U3510, P1_U3513, P1_U3515, P1_U3516, P1_U3517, P1_U3518, 
        P1_U3519, P1_U3520, P1_U3521, P1_U3522, P1_U3523, P1_U3524, P1_U3525, 
        P1_U3526, P1_U3527, P1_U3528, P1_U3529, P1_U3530, P1_U3531, P1_U3532, 
        P1_U3533, P1_U3534, P1_U3535, P1_U3536, P1_U3537, P1_U3538, P1_U3539, 
        P1_U3540, P1_U3541, P1_U3542, P1_U3543, P1_U3544, P1_U3545, P1_U3546, 
        P1_U3547, P1_U3548, P1_U3549, P1_U3550, P1_U3551, P1_U3552, P1_U3553, 
        P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3293, 
        P1_U3292, P1_U3291, P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, 
        P1_U3285, P1_U3284, P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, 
        P1_U3278, P1_U3277, P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, 
        P1_U3271, P1_U3270, P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, 
        P1_U3356, P1_U3264, P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, 
        P1_U3258, P1_U3257, P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, 
        P1_U3251, P1_U3250, P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, 
        P1_U3244, P1_U3243, P1_U3560, P1_U3561, P1_U3562, P1_U3563, P1_U3564, 
        P1_U3565, P1_U3566, P1_U3567, P1_U3568, P1_U3569, P1_U3570, P1_U3571, 
        P1_U3572, P1_U3573, P1_U3574, P1_U3575, P1_U3576, P1_U3577, P1_U3578, 
        P1_U3579, P1_U3580, P1_U3581, P1_U3582, P1_U3583, P1_U3584, P1_U3585, 
        P1_U3586, P1_U3587, P1_U3588, P1_U3589, P1_U3590, P1_U3591, P1_U3242, 
        P1_U3241, P1_U3240, P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, 
        P1_U3234, P1_U3233, P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, 
        P1_U3227, P1_U3226, P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, 
        P1_U3220, P1_U3219, P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, 
        P1_U3213, P1_U3086, P1_U3085, P1_U4016, P2_U3327, P2_U3326, P2_U3325, 
        P2_U3324, P2_U3323, P2_U3322, P2_U3321, P2_U3320, P2_U3319, P2_U3318, 
        P2_U3317, P2_U3316, P2_U3315, P2_U3314, P2_U3313, P2_U3312, P2_U3311, 
        P2_U3310, P2_U3309, P2_U3308, P2_U3307, P2_U3306, P2_U3305, P2_U3304, 
        P2_U3303, P2_U3302, P2_U3301, P2_U3300, P2_U3299, P2_U3298, P2_U3297, 
        P2_U3296, P2_U3416, P2_U3417, P2_U3295, P2_U3294, P2_U3293, P2_U3292, 
        P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, 
        P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, 
        P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, 
        P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3430, P2_U3433, 
        P2_U3436, P2_U3439, P2_U3442, P2_U3445, P2_U3448, P2_U3451, P2_U3454, 
        P2_U3457, P2_U3460, P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, 
        P2_U3478, P2_U3481, P2_U3484, P2_U3486, P2_U3487, P2_U3488, P2_U3489, 
        P2_U3490, P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, 
        P2_U3497, P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, 
        P2_U3504, P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, 
        P2_U3511, P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, 
        P2_U3518, P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, 
        P2_U3525, P2_U3526, P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3265, 
        P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258, 
        P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251, 
        P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244, 
        P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, 
        P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, 
        P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, 
        P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, 
        P2_U3215, P2_U3214, P2_U3531, P2_U3532, P2_U3533, P2_U3534, P2_U3535, 
        P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540, P2_U3541, P2_U3542, 
        P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547, P2_U3548, P2_U3549, 
        P2_U3550, P2_U3551, P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, 
        P2_U3557, P2_U3558, P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3328, 
        P2_U3213, P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3208, P2_U3207, 
        P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, 
        P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, 
        P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, 
        P2_U3185, P2_U3088, P2_U3087, P2_U3947, P3_U3295, P3_U3294, P3_U3293, 
        P3_U3292, P3_U3291, P3_U3290, P3_U3289, P3_U3288, P3_U3287, P3_U3286, 
        P3_U3285, P3_U3284, P3_U3283, P3_U3282, P3_U3281, P3_U3280, P3_U3279, 
        P3_U3278, P3_U3277, P3_U3276, P3_U3275, P3_U3274, P3_U3273, P3_U3272, 
        P3_U3271, P3_U3270, P3_U3269, P3_U3268, P3_U3267, P3_U3266, P3_U3265, 
        P3_U3264, P3_U3376, P3_U3377, P3_U3263, P3_U3262, P3_U3261, P3_U3260, 
        P3_U3259, P3_U3258, P3_U3257, P3_U3256, P3_U3255, P3_U3254, P3_U3253, 
        P3_U3252, P3_U3251, P3_U3250, P3_U3249, P3_U3248, P3_U3247, P3_U3246, 
        P3_U3245, P3_U3244, P3_U3243, P3_U3242, P3_U3241, P3_U3240, P3_U3239, 
        P3_U3238, P3_U3237, P3_U3236, P3_U3235, P3_U3234, P3_U3390, P3_U3393, 
        P3_U3396, P3_U3399, P3_U3402, P3_U3405, P3_U3408, P3_U3411, P3_U3414, 
        P3_U3417, P3_U3420, P3_U3423, P3_U3426, P3_U3429, P3_U3432, P3_U3435, 
        P3_U3438, P3_U3441, P3_U3444, P3_U3446, P3_U3447, P3_U3448, P3_U3449, 
        P3_U3450, P3_U3451, P3_U3452, P3_U3453, P3_U3454, P3_U3455, P3_U3456, 
        P3_U3457, P3_U3458, P3_U3459, P3_U3460, P3_U3461, P3_U3462, P3_U3463, 
        P3_U3464, P3_U3465, P3_U3466, P3_U3467, P3_U3468, P3_U3469, P3_U3470, 
        P3_U3471, P3_U3472, P3_U3473, P3_U3474, P3_U3475, P3_U3476, P3_U3477, 
        P3_U3478, P3_U3479, P3_U3480, P3_U3481, P3_U3482, P3_U3483, P3_U3484, 
        P3_U3485, P3_U3486, P3_U3487, P3_U3488, P3_U3489, P3_U3490, P3_U3233, 
        P3_U3232, P3_U3231, P3_U3230, P3_U3229, P3_U3228, P3_U3227, P3_U3226, 
        P3_U3225, P3_U3224, P3_U3223, P3_U3222, P3_U3221, P3_U3220, P3_U3219, 
        P3_U3218, P3_U3217, P3_U3216, P3_U3215, P3_U3214, P3_U3213, P3_U3212, 
        P3_U3211, P3_U3210, P3_U3209, P3_U3208, P3_U3207, P3_U3206, P3_U3205, 
        P3_U3204, P3_U3203, P3_U3202, P3_U3201, P3_U3200, P3_U3199, P3_U3198, 
        P3_U3197, P3_U3196, P3_U3195, P3_U3194, P3_U3193, P3_U3192, P3_U3191, 
        P3_U3190, P3_U3189, P3_U3188, P3_U3187, P3_U3186, P3_U3185, P3_U3184, 
        P3_U3183, P3_U3182, P3_U3491, P3_U3492, P3_U3493, P3_U3494, P3_U3495, 
        P3_U3496, P3_U3497, P3_U3498, P3_U3499, P3_U3500, P3_U3501, P3_U3502, 
        P3_U3503, P3_U3504, P3_U3505, P3_U3506, P3_U3507, P3_U3508, P3_U3509, 
        P3_U3510, P3_U3511, P3_U3512, P3_U3513, P3_U3514, P3_U3515, P3_U3516, 
        P3_U3517, P3_U3518, P3_U3519, P3_U3520, P3_U3521, P3_U3522, P3_U3296, 
        P3_U3181, P3_U3180, P3_U3179, P3_U3178, P3_U3177, P3_U3176, P3_U3175, 
        P3_U3174, P3_U3173, P3_U3172, P3_U3171, P3_U3170, P3_U3169, P3_U3168, 
        P3_U3167, P3_U3166, P3_U3165, P3_U3164, P3_U3163, P3_U3162, P3_U3161, 
        P3_U3160, P3_U3159, P3_U3158, P3_U3157, P3_U3156, P3_U3155, P3_U3154, 
        P3_U3153, P3_U3151, P3_U3150, P3_U3897 );
  input P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN,
         P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN,
         P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN,
         P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN,
         P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN,
         P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN,
         P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN,
         P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN,
         P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN,
         P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN,
         P3_REG3_REG_0__SCAN_IN, P3_REG3_REG_20__SCAN_IN,
         P3_REG3_REG_13__SCAN_IN, P3_REG3_REG_22__SCAN_IN,
         P3_REG3_REG_11__SCAN_IN, P3_REG3_REG_2__SCAN_IN,
         P3_REG3_REG_18__SCAN_IN, P3_REG3_REG_6__SCAN_IN,
         P3_REG3_REG_26__SCAN_IN, P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN,
         P3_DATAO_REG_31__SCAN_IN, P3_DATAO_REG_30__SCAN_IN,
         P3_DATAO_REG_29__SCAN_IN, P3_DATAO_REG_28__SCAN_IN,
         P3_DATAO_REG_27__SCAN_IN, P3_DATAO_REG_26__SCAN_IN,
         P3_DATAO_REG_25__SCAN_IN, P3_DATAO_REG_24__SCAN_IN,
         P3_DATAO_REG_23__SCAN_IN, P3_DATAO_REG_22__SCAN_IN,
         P3_DATAO_REG_21__SCAN_IN, P3_DATAO_REG_20__SCAN_IN,
         P3_DATAO_REG_19__SCAN_IN, P3_DATAO_REG_18__SCAN_IN,
         P3_DATAO_REG_17__SCAN_IN, P3_DATAO_REG_16__SCAN_IN,
         P3_DATAO_REG_15__SCAN_IN, P3_DATAO_REG_14__SCAN_IN,
         P3_DATAO_REG_13__SCAN_IN, P3_DATAO_REG_12__SCAN_IN,
         P3_DATAO_REG_11__SCAN_IN, P3_DATAO_REG_10__SCAN_IN,
         P3_DATAO_REG_9__SCAN_IN, P3_DATAO_REG_8__SCAN_IN,
         P3_DATAO_REG_7__SCAN_IN, P3_DATAO_REG_6__SCAN_IN,
         P3_DATAO_REG_5__SCAN_IN, P3_DATAO_REG_4__SCAN_IN,
         P3_DATAO_REG_3__SCAN_IN, P3_DATAO_REG_2__SCAN_IN,
         P3_DATAO_REG_1__SCAN_IN, P3_DATAO_REG_0__SCAN_IN,
         P3_ADDR_REG_0__SCAN_IN, P3_ADDR_REG_1__SCAN_IN,
         P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN,
         P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN,
         P3_ADDR_REG_6__SCAN_IN, P3_ADDR_REG_7__SCAN_IN,
         P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, P1_IR_REG_0__SCAN_IN,
         P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN,
         P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN,
         P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN,
         P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN,
         P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN,
         P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN,
         P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN,
         P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN,
         P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN,
         P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN,
         P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN,
         P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN,
         P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN,
         P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN,
         P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN,
         P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN,
         P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN,
         P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN,
         P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN,
         P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN,
         P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN,
         P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN,
         P2_RD_REG_SCAN_IN, P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN,
         P3_IR_REG_1__SCAN_IN, P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN,
         P3_IR_REG_4__SCAN_IN, P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN,
         P3_IR_REG_7__SCAN_IN, P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN,
         P3_IR_REG_10__SCAN_IN, P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN,
         P3_IR_REG_13__SCAN_IN, P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN,
         P3_IR_REG_16__SCAN_IN, P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN,
         P3_IR_REG_19__SCAN_IN, P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN,
         P3_IR_REG_22__SCAN_IN, P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN,
         P3_IR_REG_25__SCAN_IN, P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN,
         P3_IR_REG_28__SCAN_IN, P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN,
         P3_IR_REG_31__SCAN_IN, P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN,
         P3_D_REG_2__SCAN_IN, P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN,
         P3_D_REG_5__SCAN_IN, P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN,
         P3_D_REG_8__SCAN_IN, P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN,
         P3_D_REG_11__SCAN_IN, P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN,
         P3_D_REG_14__SCAN_IN, P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN,
         P3_D_REG_17__SCAN_IN, P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN,
         P3_D_REG_20__SCAN_IN, P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN,
         P3_D_REG_23__SCAN_IN, P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN,
         P3_D_REG_26__SCAN_IN, P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN,
         P3_D_REG_29__SCAN_IN, P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN,
         P3_REG0_REG_0__SCAN_IN, P3_REG0_REG_1__SCAN_IN,
         P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN,
         P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN,
         P3_REG0_REG_6__SCAN_IN, P3_REG0_REG_7__SCAN_IN,
         P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN,
         P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN,
         P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN,
         P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN,
         P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN,
         P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN,
         P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN,
         P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN,
         P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN,
         P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN,
         P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN,
         P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN,
         P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN,
         P3_REG1_REG_2__SCAN_IN, P3_REG1_REG_3__SCAN_IN,
         P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN,
         P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN,
         P3_REG1_REG_8__SCAN_IN, P3_REG1_REG_9__SCAN_IN,
         P3_REG1_REG_10__SCAN_IN, P3_REG1_REG_11__SCAN_IN,
         P3_REG1_REG_12__SCAN_IN, P3_REG1_REG_13__SCAN_IN,
         P3_REG1_REG_14__SCAN_IN, P3_REG1_REG_15__SCAN_IN,
         P3_REG1_REG_16__SCAN_IN, P3_REG1_REG_17__SCAN_IN,
         P3_REG1_REG_18__SCAN_IN, P3_REG1_REG_19__SCAN_IN,
         P3_REG1_REG_20__SCAN_IN, P3_REG1_REG_21__SCAN_IN,
         P3_REG1_REG_22__SCAN_IN, P3_REG1_REG_23__SCAN_IN,
         P3_REG1_REG_24__SCAN_IN, P3_REG1_REG_25__SCAN_IN,
         P3_REG1_REG_26__SCAN_IN, P3_REG1_REG_27__SCAN_IN,
         P3_REG1_REG_28__SCAN_IN, P3_REG1_REG_29__SCAN_IN,
         P3_REG1_REG_30__SCAN_IN, P3_REG1_REG_31__SCAN_IN,
         P3_REG2_REG_0__SCAN_IN, P3_REG2_REG_1__SCAN_IN,
         P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN,
         P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN,
         P3_REG2_REG_6__SCAN_IN, P3_REG2_REG_7__SCAN_IN,
         P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN,
         P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN,
         P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN,
         P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN,
         P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN,
         P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN,
         P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN,
         P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN,
         P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN,
         P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN,
         P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN,
         P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN,
         P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN,
         P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN,
         P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN,
         P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN,
         P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, keyinput_f0,
         keyinput_f1, keyinput_f2, keyinput_f3, keyinput_f4, keyinput_f5,
         keyinput_f6, keyinput_f7, keyinput_f8, keyinput_f9, keyinput_f10,
         keyinput_f11, keyinput_f12, keyinput_f13, keyinput_f14, keyinput_f15,
         keyinput_f16, keyinput_f17, keyinput_f18, keyinput_f19, keyinput_f20,
         keyinput_f21, keyinput_f22, keyinput_f23, keyinput_f24, keyinput_f25,
         keyinput_f26, keyinput_f27, keyinput_f28, keyinput_f29, keyinput_f30,
         keyinput_f31, keyinput_f32, keyinput_f33, keyinput_f34, keyinput_f35,
         keyinput_f36, keyinput_f37, keyinput_f38, keyinput_f39, keyinput_f40,
         keyinput_f41, keyinput_f42, keyinput_f43, keyinput_f44, keyinput_f45,
         keyinput_f46, keyinput_f47, keyinput_f48, keyinput_f49, keyinput_f50,
         keyinput_f51, keyinput_f52, keyinput_f53, keyinput_f54, keyinput_f55,
         keyinput_f56, keyinput_f57, keyinput_f58, keyinput_f59, keyinput_f60,
         keyinput_f61, keyinput_f62, keyinput_f63, keyinput_f64, keyinput_f65,
         keyinput_f66, keyinput_f67, keyinput_f68, keyinput_f69, keyinput_f70,
         keyinput_f71, keyinput_f72, keyinput_f73, keyinput_f74, keyinput_f75,
         keyinput_f76, keyinput_f77, keyinput_f78, keyinput_f79, keyinput_f80,
         keyinput_f81, keyinput_f82, keyinput_f83, keyinput_f84, keyinput_f85,
         keyinput_f86, keyinput_f87, keyinput_f88, keyinput_f89, keyinput_f90,
         keyinput_f91, keyinput_f92, keyinput_f93, keyinput_f94, keyinput_f95,
         keyinput_f96, keyinput_f97, keyinput_f98, keyinput_f99, keyinput_f100,
         keyinput_f101, keyinput_f102, keyinput_f103, keyinput_f104,
         keyinput_f105, keyinput_f106, keyinput_f107, keyinput_f108,
         keyinput_f109, keyinput_f110, keyinput_f111, keyinput_f112,
         keyinput_f113, keyinput_f114, keyinput_f115, keyinput_f116,
         keyinput_f117, keyinput_f118, keyinput_f119, keyinput_f120,
         keyinput_f121, keyinput_f122, keyinput_f123, keyinput_f124,
         keyinput_f125, keyinput_f126, keyinput_f127, keyinput_g0, keyinput_g1,
         keyinput_g2, keyinput_g3, keyinput_g4, keyinput_g5, keyinput_g6,
         keyinput_g7, keyinput_g8, keyinput_g9, keyinput_g10, keyinput_g11,
         keyinput_g12, keyinput_g13, keyinput_g14, keyinput_g15, keyinput_g16,
         keyinput_g17, keyinput_g18, keyinput_g19, keyinput_g20, keyinput_g21,
         keyinput_g22, keyinput_g23, keyinput_g24, keyinput_g25, keyinput_g26,
         keyinput_g27, keyinput_g28, keyinput_g29, keyinput_g30, keyinput_g31,
         keyinput_g32, keyinput_g33, keyinput_g34, keyinput_g35, keyinput_g36,
         keyinput_g37, keyinput_g38, keyinput_g39, keyinput_g40, keyinput_g41,
         keyinput_g42, keyinput_g43, keyinput_g44, keyinput_g45, keyinput_g46,
         keyinput_g47, keyinput_g48, keyinput_g49, keyinput_g50, keyinput_g51,
         keyinput_g52, keyinput_g53, keyinput_g54, keyinput_g55, keyinput_g56,
         keyinput_g57, keyinput_g58, keyinput_g59, keyinput_g60, keyinput_g61,
         keyinput_g62, keyinput_g63, keyinput_g64, keyinput_g65, keyinput_g66,
         keyinput_g67, keyinput_g68, keyinput_g69, keyinput_g70, keyinput_g71,
         keyinput_g72, keyinput_g73, keyinput_g74, keyinput_g75, keyinput_g76,
         keyinput_g77, keyinput_g78, keyinput_g79, keyinput_g80, keyinput_g81,
         keyinput_g82, keyinput_g83, keyinput_g84, keyinput_g85, keyinput_g86,
         keyinput_g87, keyinput_g88, keyinput_g89, keyinput_g90, keyinput_g91,
         keyinput_g92, keyinput_g93, keyinput_g94, keyinput_g95, keyinput_g96,
         keyinput_g97, keyinput_g98, keyinput_g99, keyinput_g100,
         keyinput_g101, keyinput_g102, keyinput_g103, keyinput_g104,
         keyinput_g105, keyinput_g106, keyinput_g107, keyinput_g108,
         keyinput_g109, keyinput_g110, keyinput_g111, keyinput_g112,
         keyinput_g113, keyinput_g114, keyinput_g115, keyinput_g116,
         keyinput_g117, keyinput_g118, keyinput_g119, keyinput_g120,
         keyinput_g121, keyinput_g122, keyinput_g123, keyinput_g124,
         keyinput_g125, keyinput_g126, keyinput_g127;
  output SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65,
         SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70,
         SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58,
         SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53,
         U29, U28, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350,
         P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343,
         P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336,
         P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329,
         P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446,
         P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317,
         P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310,
         P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303,
         P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296,
         P1_U3295, P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471,
         P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492,
         P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556,
         P1_U3557, P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290,
         P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283,
         P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276,
         P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269,
         P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263,
         P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256,
         P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249,
         P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588,
         P1_U3589, P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239,
         P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232,
         P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085,
         P1_U4016, P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322,
         P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315,
         P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308,
         P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301,
         P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417,
         P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289,
         P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282,
         P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275,
         P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268,
         P2_U3267, P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442,
         P2_U3445, P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463,
         P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484,
         P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492,
         P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499,
         P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506,
         P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513,
         P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520,
         P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527,
         P2_U3528, P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262,
         P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255,
         P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248,
         P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241,
         P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234,
         P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227,
         P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220,
         P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531,
         P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538,
         P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545,
         P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552,
         P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559,
         P2_U3560, P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204,
         P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197,
         P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190,
         P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087,
         P2_U3947, P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290,
         P3_U3289, P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283,
         P3_U3282, P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276,
         P3_U3275, P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269,
         P3_U3268, P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377,
         P3_U3263, P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257,
         P3_U3256, P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250,
         P3_U3249, P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243,
         P3_U3242, P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236,
         P3_U3235, P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402,
         P3_U3405, P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423,
         P3_U3426, P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444,
         P3_U3446, P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452,
         P3_U3453, P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459,
         P3_U3460, P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466,
         P3_U3467, P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473,
         P3_U3474, P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480,
         P3_U3481, P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487,
         P3_U3488, P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230,
         P3_U3229, P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223,
         P3_U3222, P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216,
         P3_U3215, P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209,
         P3_U3208, P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202,
         P3_U3201, P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195,
         P3_U3194, P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188,
         P3_U3187, P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491,
         P3_U3492, P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498,
         P3_U3499, P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505,
         P3_U3506, P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512,
         P3_U3513, P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519,
         P3_U3520, P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179,
         P3_U3178, P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172,
         P3_U3171, P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165,
         P3_U3164, P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158,
         P3_U3157, P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150,
         P3_U3897;
  wire   n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6674, n6675,
         n6676, n6677, n6678, n6679, n6680, n6681, n6683, n6684, n6685, n6686,
         n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696,
         n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706,
         n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716,
         n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726,
         n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736,
         n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746,
         n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756,
         n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766,
         n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776,
         n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786,
         n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796,
         n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806,
         n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816,
         n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826,
         n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836,
         n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846,
         n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856,
         n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866,
         n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876,
         n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886,
         n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896,
         n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906,
         n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916,
         n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926,
         n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936,
         n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946,
         n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956,
         n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966,
         n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976,
         n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986,
         n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996,
         n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006,
         n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016,
         n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026,
         n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036,
         n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046,
         n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056,
         n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066,
         n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076,
         n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086,
         n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096,
         n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106,
         n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116,
         n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126,
         n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136,
         n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146,
         n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156,
         n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166,
         n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176,
         n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186,
         n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196,
         n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206,
         n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216,
         n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226,
         n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236,
         n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246,
         n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256,
         n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266,
         n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276,
         n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286,
         n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296,
         n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306,
         n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316,
         n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326,
         n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336,
         n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346,
         n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356,
         n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366,
         n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376,
         n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386,
         n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396,
         n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406,
         n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416,
         n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426,
         n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436,
         n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446,
         n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456,
         n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466,
         n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476,
         n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486,
         n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496,
         n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506,
         n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516,
         n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526,
         n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536,
         n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546,
         n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556,
         n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566,
         n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576,
         n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586,
         n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596,
         n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606,
         n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616,
         n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626,
         n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636,
         n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646,
         n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656,
         n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666,
         n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676,
         n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686,
         n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696,
         n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706,
         n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716,
         n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726,
         n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736,
         n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746,
         n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756,
         n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766,
         n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776,
         n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786,
         n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796,
         n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806,
         n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816,
         n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826,
         n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836,
         n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846,
         n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856,
         n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866,
         n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876,
         n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886,
         n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896,
         n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906,
         n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916,
         n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926,
         n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936,
         n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946,
         n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956,
         n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966,
         n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976,
         n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986,
         n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996,
         n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006,
         n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016,
         n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026,
         n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036,
         n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046,
         n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056,
         n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066,
         n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076,
         n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086,
         n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096,
         n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106,
         n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116,
         n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126,
         n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136,
         n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146,
         n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156,
         n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166,
         n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176,
         n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186,
         n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196,
         n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206,
         n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216,
         n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226,
         n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236,
         n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246,
         n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256,
         n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266,
         n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276,
         n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286,
         n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296,
         n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306,
         n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316,
         n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326,
         n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336,
         n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346,
         n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356,
         n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366,
         n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376,
         n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386,
         n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396,
         n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406,
         n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416,
         n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426,
         n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436,
         n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446,
         n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456,
         n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466,
         n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476,
         n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486,
         n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496,
         n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506,
         n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516,
         n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526,
         n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536,
         n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546,
         n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556,
         n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566,
         n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576,
         n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586,
         n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596,
         n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606,
         n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616,
         n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626,
         n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636,
         n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646,
         n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656,
         n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666,
         n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676,
         n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686,
         n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696,
         n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706,
         n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716,
         n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726,
         n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736,
         n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746,
         n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756,
         n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766,
         n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776,
         n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786,
         n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796,
         n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806,
         n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816,
         n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826,
         n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836,
         n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846,
         n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856,
         n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866,
         n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876,
         n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886,
         n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896,
         n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906,
         n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916,
         n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926,
         n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936,
         n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946,
         n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956,
         n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966,
         n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976,
         n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986,
         n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996,
         n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006,
         n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9017,
         n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027,
         n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037,
         n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047,
         n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057,
         n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067,
         n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077,
         n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087,
         n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097,
         n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107,
         n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117,
         n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127,
         n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137,
         n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147,
         n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157,
         n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167,
         n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177,
         n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187,
         n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197,
         n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207,
         n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217,
         n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227,
         n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237,
         n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247,
         n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257,
         n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267,
         n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277,
         n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287,
         n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297,
         n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307,
         n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317,
         n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327,
         n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337,
         n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347,
         n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357,
         n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367,
         n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377,
         n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387,
         n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397,
         n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407,
         n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417,
         n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427,
         n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437,
         n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447,
         n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457,
         n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467,
         n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477,
         n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487,
         n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497,
         n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507,
         n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517,
         n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527,
         n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537,
         n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547,
         n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557,
         n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567,
         n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577,
         n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587,
         n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597,
         n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607,
         n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617,
         n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627,
         n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637,
         n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647,
         n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657,
         n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667,
         n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677,
         n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687,
         n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697,
         n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707,
         n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717,
         n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727,
         n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737,
         n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747,
         n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757,
         n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767,
         n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777,
         n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787,
         n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797,
         n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807,
         n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817,
         n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827,
         n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837,
         n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847,
         n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857,
         n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867,
         n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877,
         n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887,
         n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897,
         n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907,
         n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917,
         n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927,
         n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937,
         n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947,
         n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957,
         n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967,
         n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977,
         n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987,
         n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997,
         n9998, n9999, n10000, n10001, n10002, n10003, n10004, n10005, n10006,
         n10007, n10008, n10009, n10010, n10011, n10012, n10013, n10014,
         n10015, n10016, n10017, n10018, n10019, n10020, n10021, n10022,
         n10023, n10024, n10025, n10026, n10027, n10028, n10029, n10030,
         n10031, n10032, n10033, n10034, n10035, n10036, n10037, n10038,
         n10039, n10040, n10041, n10042, n10043, n10044, n10045, n10046,
         n10047, n10048, n10049, n10050, n10051, n10052, n10053, n10054,
         n10055, n10056, n10057, n10058, n10059, n10060, n10061, n10062,
         n10063, n10064, n10065, n10066, n10067, n10068, n10069, n10070,
         n10071, n10072, n10073, n10074, n10075, n10076, n10077, n10078,
         n10079, n10080, n10081, n10082, n10083, n10084, n10085, n10086,
         n10087, n10088, n10089, n10090, n10091, n10092, n10093, n10094,
         n10095, n10096, n10097, n10098, n10099, n10100, n10101, n10102,
         n10103, n10104, n10105, n10106, n10107, n10108, n10109, n10110,
         n10111, n10112, n10113, n10114, n10115, n10116, n10117, n10118,
         n10119, n10120, n10121, n10122, n10123, n10124, n10125, n10126,
         n10127, n10128, n10129, n10130, n10131, n10132, n10133, n10134,
         n10135, n10136, n10137, n10138, n10139, n10140, n10141, n10142,
         n10143, n10144, n10145, n10146, n10147, n10148, n10149, n10150,
         n10151, n10152, n10153, n10154, n10155, n10156, n10157, n10158,
         n10159, n10160, n10161, n10162, n10163, n10164, n10165, n10166,
         n10167, n10168, n10169, n10170, n10171, n10172, n10173, n10174,
         n10175, n10176, n10177, n10178, n10179, n10180, n10181, n10182,
         n10183, n10184, n10185, n10186, n10187, n10188, n10189, n10190,
         n10191, n10192, n10193, n10194, n10195, n10196, n10197, n10198,
         n10199, n10200, n10201, n10202, n10203, n10204, n10205, n10206,
         n10207, n10208, n10209, n10210, n10211, n10212, n10213, n10214,
         n10215, n10216, n10217, n10218, n10219, n10220, n10221, n10222,
         n10223, n10224, n10225, n10226, n10227, n10228, n10229, n10230,
         n10231, n10232, n10233, n10234, n10235, n10236, n10237, n10238,
         n10239, n10240, n10241, n10242, n10243, n10244, n10245, n10246,
         n10247, n10248, n10249, n10250, n10251, n10252, n10253, n10254,
         n10255, n10256, n10257, n10258, n10259, n10260, n10261, n10262,
         n10263, n10264, n10265, n10266, n10267, n10268, n10269, n10270,
         n10271, n10272, n10273, n10274, n10275, n10276, n10277, n10278,
         n10279, n10280, n10281, n10282, n10283, n10284, n10285, n10286,
         n10287, n10288, n10289, n10290, n10291, n10292, n10293, n10294,
         n10295, n10296, n10297, n10298, n10299, n10300, n10301, n10302,
         n10303, n10304, n10305, n10306, n10307, n10308, n10309, n10310,
         n10311, n10312, n10313, n10314, n10315, n10316, n10317, n10318,
         n10319, n10320, n10321, n10322, n10323, n10324, n10325, n10326,
         n10327, n10328, n10329, n10330, n10331, n10332, n10333, n10334,
         n10335, n10336, n10337, n10338, n10339, n10340, n10341, n10342,
         n10343, n10344, n10345, n10346, n10347, n10348, n10349, n10350,
         n10351, n10352, n10353, n10354, n10355, n10356, n10357, n10358,
         n10359, n10360, n10361, n10362, n10363, n10364, n10365, n10366,
         n10367, n10368, n10369, n10370, n10371, n10372, n10373, n10374,
         n10375, n10376, n10377, n10378, n10379, n10380, n10381, n10382,
         n10383, n10384, n10385, n10386, n10387, n10388, n10389, n10390,
         n10391, n10392, n10393, n10394, n10395, n10396, n10397, n10398,
         n10399, n10400, n10401, n10402, n10403, n10404, n10405, n10406,
         n10407, n10408, n10409, n10410, n10411, n10412, n10413, n10414,
         n10415, n10416, n10417, n10418, n10419, n10420, n10421, n10422,
         n10423, n10424, n10425, n10426, n10427, n10428, n10429, n10430,
         n10431, n10432, n10433, n10434, n10435, n10436, n10437, n10438,
         n10439, n10440, n10441, n10442, n10443, n10444, n10445, n10446,
         n10447, n10448, n10449, n10450, n10451, n10452, n10453, n10454,
         n10455, n10456, n10457, n10458, n10459, n10460, n10461, n10462,
         n10463, n10464, n10465, n10466, n10467, n10468, n10469, n10470,
         n10471, n10472, n10473, n10474, n10475, n10476, n10477, n10478,
         n10479, n10480, n10481, n10482, n10483, n10484, n10485, n10486,
         n10487, n10488, n10489, n10490, n10491, n10492, n10493, n10494,
         n10495, n10496, n10497, n10498, n10499, n10500, n10501, n10502,
         n10503, n10504, n10505, n10506, n10507, n10508, n10509, n10510,
         n10511, n10512, n10513, n10514, n10515, n10516, n10517, n10518,
         n10519, n10520, n10521, n10522, n10523, n10524, n10525, n10526,
         n10527, n10528, n10529, n10530, n10531, n10532, n10533, n10534,
         n10535, n10536, n10537, n10538, n10539, n10540, n10541, n10542,
         n10543, n10544, n10545, n10546, n10547, n10548, n10549, n10550,
         n10551, n10552, n10553, n10554, n10555, n10556, n10557, n10558,
         n10559, n10560, n10561, n10562, n10563, n10564, n10565, n10566,
         n10567, n10568, n10569, n10570, n10571, n10572, n10573, n10574,
         n10575, n10576, n10577, n10578, n10579, n10580, n10581, n10582,
         n10583, n10584, n10585, n10586, n10587, n10588, n10589, n10590,
         n10591, n10592, n10593, n10594, n10595, n10596, n10597, n10598,
         n10599, n10600, n10601, n10602, n10603, n10604, n10605, n10606,
         n10607, n10608, n10609, n10610, n10611, n10612, n10613, n10614,
         n10615, n10616, n10617, n10618, n10619, n10620, n10621, n10622,
         n10623, n10624, n10625, n10626, n10627, n10628, n10629, n10630,
         n10631, n10632, n10633, n10634, n10635, n10636, n10637, n10638,
         n10639, n10640, n10641, n10642, n10643, n10644, n10645, n10646,
         n10647, n10648, n10649, n10650, n10651, n10652, n10653, n10654,
         n10655, n10656, n10657, n10658, n10659, n10660, n10661, n10662,
         n10663, n10664, n10665, n10666, n10667, n10668, n10669, n10670,
         n10671, n10672, n10673, n10674, n10675, n10676, n10677, n10678,
         n10679, n10680, n10681, n10682, n10683, n10684, n10685, n10686,
         n10687, n10688, n10689, n10690, n10691, n10692, n10693, n10694,
         n10695, n10696, n10697, n10698, n10699, n10700, n10701, n10702,
         n10703, n10704, n10705, n10706, n10707, n10708, n10709, n10710,
         n10711, n10712, n10713, n10714, n10715, n10716, n10717, n10718,
         n10719, n10720, n10721, n10722, n10723, n10724, n10725, n10726,
         n10727, n10728, n10729, n10730, n10731, n10732, n10733, n10734,
         n10735, n10736, n10737, n10738, n10739, n10740, n10741, n10742,
         n10743, n10744, n10745, n10746, n10747, n10748, n10749, n10750,
         n10751, n10752, n10753, n10754, n10755, n10756, n10757, n10758,
         n10759, n10760, n10761, n10762, n10763, n10764, n10765, n10766,
         n10767, n10768, n10769, n10770, n10771, n10772, n10773, n10774,
         n10775, n10776, n10777, n10778, n10779, n10780, n10781, n10782,
         n10783, n10784, n10785, n10786, n10787, n10788, n10789, n10790,
         n10791, n10792, n10793, n10794, n10795, n10796, n10797, n10798,
         n10799, n10800, n10801, n10802, n10803, n10804, n10805, n10806,
         n10807, n10808, n10809, n10810, n10811, n10812, n10813, n10814,
         n10815, n10816, n10817, n10818, n10819, n10820, n10821, n10822,
         n10823, n10824, n10825, n10826, n10827, n10828, n10829, n10830,
         n10831, n10832, n10833, n10834, n10835, n10836, n10837, n10838,
         n10839, n10840, n10841, n10842, n10843, n10844, n10845, n10846,
         n10847, n10848, n10849, n10850, n10851, n10852, n10853, n10854,
         n10855, n10856, n10857, n10858, n10859, n10860, n10861, n10862,
         n10863, n10864, n10865, n10866, n10867, n10868, n10869, n10870,
         n10871, n10872, n10873, n10874, n10875, n10876, n10877, n10878,
         n10879, n10880, n10881, n10882, n10883, n10884, n10885, n10886,
         n10887, n10888, n10889, n10890, n10891, n10892, n10893, n10894,
         n10895, n10896, n10897, n10898, n10899, n10900, n10901, n10902,
         n10903, n10904, n10905, n10906, n10907, n10908, n10909, n10910,
         n10911, n10912, n10913, n10914, n10915, n10916, n10917, n10918,
         n10919, n10920, n10921, n10922, n10923, n10924, n10925, n10926,
         n10927, n10928, n10929, n10930, n10931, n10932, n10933, n10934,
         n10935, n10936, n10937, n10938, n10939, n10940, n10941, n10942,
         n10943, n10944, n10945, n10946, n10947, n10948, n10949, n10950,
         n10951, n10952, n10953, n10954, n10955, n10956, n10957, n10958,
         n10959, n10960, n10961, n10962, n10963, n10964, n10965, n10966,
         n10967, n10968, n10969, n10970, n10971, n10972, n10973, n10974,
         n10975, n10976, n10977, n10978, n10979, n10980, n10981, n10982,
         n10983, n10984, n10985, n10986, n10987, n10988, n10989, n10990,
         n10991, n10992, n10993, n10994, n10995, n10996, n10997, n10998,
         n10999, n11000, n11001, n11002, n11003, n11004, n11005, n11006,
         n11007, n11008, n11009, n11010, n11011, n11012, n11013, n11014,
         n11015, n11016, n11017, n11018, n11019, n11020, n11021, n11022,
         n11023, n11024, n11025, n11026, n11027, n11028, n11029, n11030,
         n11031, n11032, n11033, n11034, n11035, n11036, n11037, n11038,
         n11039, n11040, n11041, n11042, n11043, n11044, n11045, n11046,
         n11047, n11048, n11049, n11050, n11051, n11052, n11053, n11054,
         n11055, n11056, n11057, n11058, n11059, n11060, n11061, n11062,
         n11063, n11064, n11065, n11066, n11067, n11068, n11069, n11070,
         n11071, n11072, n11073, n11074, n11075, n11076, n11077, n11078,
         n11079, n11080, n11081, n11082, n11083, n11084, n11085, n11086,
         n11087, n11088, n11089, n11090, n11091, n11092, n11093, n11094,
         n11095, n11096, n11097, n11098, n11099, n11100, n11101, n11102,
         n11103, n11104, n11105, n11106, n11107, n11108, n11109, n11110,
         n11111, n11112, n11113, n11114, n11115, n11116, n11117, n11118,
         n11119, n11120, n11121, n11122, n11123, n11124, n11125, n11126,
         n11127, n11128, n11129, n11130, n11131, n11132, n11133, n11134,
         n11135, n11136, n11137, n11138, n11139, n11140, n11141, n11142,
         n11143, n11144, n11145, n11146, n11147, n11148, n11149, n11150,
         n11151, n11152, n11153, n11154, n11155, n11156, n11157, n11158,
         n11159, n11160, n11161, n11162, n11163, n11164, n11165, n11166,
         n11167, n11168, n11169, n11170, n11171, n11172, n11173, n11174,
         n11175, n11176, n11177, n11178, n11179, n11180, n11181, n11182,
         n11183, n11184, n11185, n11186, n11187, n11188, n11189, n11190,
         n11191, n11192, n11193, n11194, n11195, n11196, n11197, n11198,
         n11199, n11200, n11201, n11202, n11203, n11204, n11205, n11206,
         n11207, n11208, n11209, n11210, n11211, n11212, n11213, n11214,
         n11215, n11216, n11217, n11218, n11219, n11220, n11221, n11222,
         n11223, n11224, n11225, n11226, n11227, n11228, n11229, n11230,
         n11231, n11232, n11233, n11234, n11235, n11236, n11237, n11238,
         n11239, n11240, n11241, n11242, n11243, n11244, n11245, n11246,
         n11247, n11248, n11249, n11250, n11251, n11252, n11253, n11254,
         n11255, n11256, n11257, n11258, n11259, n11260, n11261, n11262,
         n11263, n11264, n11265, n11266, n11267, n11268, n11269, n11270,
         n11271, n11272, n11273, n11274, n11275, n11276, n11277, n11278,
         n11279, n11280, n11281, n11282, n11283, n11284, n11285, n11286,
         n11287, n11288, n11289, n11290, n11291, n11292, n11293, n11294,
         n11295, n11296, n11297, n11298, n11299, n11300, n11301, n11302,
         n11303, n11304, n11305, n11306, n11307, n11308, n11309, n11310,
         n11311, n11312, n11313, n11314, n11315, n11316, n11317, n11318,
         n11319, n11320, n11321, n11322, n11323, n11324, n11325, n11326,
         n11327, n11328, n11329, n11330, n11331, n11332, n11333, n11334,
         n11335, n11336, n11337, n11338, n11339, n11340, n11341, n11342,
         n11343, n11344, n11345, n11346, n11347, n11348, n11349, n11350,
         n11351, n11352, n11353, n11354, n11355, n11356, n11357, n11358,
         n11359, n11360, n11361, n11362, n11363, n11364, n11365, n11366,
         n11367, n11368, n11369, n11370, n11371, n11372, n11373, n11374,
         n11375, n11376, n11377, n11378, n11379, n11380, n11381, n11382,
         n11383, n11384, n11385, n11386, n11387, n11388, n11389, n11390,
         n11391, n11392, n11393, n11394, n11395, n11396, n11397, n11398,
         n11399, n11400, n11401, n11402, n11403, n11404, n11405, n11406,
         n11407, n11408, n11409, n11410, n11411, n11412, n11413, n11414,
         n11415, n11416, n11417, n11418, n11419, n11420, n11421, n11422,
         n11423, n11424, n11425, n11426, n11427, n11428, n11429, n11430,
         n11431, n11432, n11433, n11434, n11435, n11436, n11437, n11438,
         n11439, n11440, n11441, n11442, n11443, n11444, n11445, n11446,
         n11447, n11448, n11449, n11450, n11451, n11452, n11453, n11454,
         n11455, n11456, n11457, n11458, n11459, n11460, n11461, n11462,
         n11463, n11464, n11465, n11466, n11467, n11468, n11469, n11470,
         n11471, n11472, n11473, n11474, n11475, n11476, n11477, n11478,
         n11479, n11480, n11481, n11482, n11483, n11484, n11485, n11486,
         n11487, n11488, n11489, n11490, n11491, n11492, n11493, n11494,
         n11495, n11496, n11497, n11498, n11499, n11500, n11501, n11502,
         n11503, n11504, n11505, n11506, n11507, n11508, n11509, n11510,
         n11511, n11512, n11513, n11514, n11515, n11516, n11517, n11518,
         n11519, n11520, n11521, n11522, n11523, n11524, n11525, n11526,
         n11527, n11528, n11529, n11530, n11531, n11532, n11533, n11534,
         n11535, n11536, n11537, n11538, n11539, n11540, n11541, n11542,
         n11543, n11544, n11545, n11546, n11547, n11548, n11549, n11550,
         n11551, n11552, n11553, n11554, n11555, n11556, n11557, n11558,
         n11559, n11560, n11561, n11562, n11563, n11564, n11565, n11566,
         n11567, n11568, n11569, n11570, n11571, n11572, n11573, n11574,
         n11575, n11576, n11577, n11578, n11579, n11580, n11581, n11582,
         n11583, n11584, n11585, n11586, n11587, n11588, n11589, n11590,
         n11591, n11592, n11593, n11594, n11595, n11596, n11597, n11598,
         n11599, n11600, n11601, n11602, n11603, n11604, n11605, n11606,
         n11607, n11608, n11609, n11610, n11611, n11612, n11613, n11614,
         n11615, n11616, n11617, n11618, n11619, n11620, n11621, n11622,
         n11623, n11624, n11625, n11626, n11627, n11628, n11629, n11630,
         n11631, n11632, n11633, n11634, n11635, n11636, n11637, n11638,
         n11639, n11640, n11641, n11642, n11643, n11644, n11645, n11646,
         n11647, n11648, n11649, n11650, n11651, n11652, n11653, n11654,
         n11655, n11656, n11657, n11658, n11659, n11660, n11661, n11662,
         n11663, n11664, n11665, n11666, n11667, n11668, n11669, n11670,
         n11671, n11672, n11673, n11674, n11675, n11676, n11677, n11678,
         n11679, n11680, n11681, n11682, n11683, n11684, n11685, n11686,
         n11687, n11688, n11689, n11690, n11691, n11692, n11693, n11694,
         n11695, n11696, n11697, n11698, n11699, n11700, n11701, n11702,
         n11703, n11704, n11705, n11706, n11707, n11708, n11709, n11710,
         n11711, n11712, n11713, n11714, n11715, n11716, n11717, n11718,
         n11719, n11720, n11721, n11722, n11723, n11724, n11725, n11726,
         n11727, n11728, n11729, n11730, n11731, n11732, n11733, n11734,
         n11735, n11736, n11737, n11738, n11739, n11740, n11741, n11742,
         n11743, n11744, n11745, n11746, n11747, n11748, n11749, n11750,
         n11751, n11752, n11753, n11754, n11755, n11756, n11757, n11758,
         n11759, n11760, n11761, n11762, n11763, n11764, n11765, n11766,
         n11767, n11768, n11769, n11770, n11771, n11772, n11773, n11774,
         n11775, n11776, n11777, n11778, n11779, n11780, n11781, n11782,
         n11783, n11784, n11785, n11786, n11787, n11788, n11789, n11790,
         n11791, n11792, n11793, n11794, n11795, n11796, n11797, n11798,
         n11799, n11800, n11801, n11802, n11803, n11804, n11805, n11806,
         n11807, n11808, n11809, n11810, n11811, n11812, n11813, n11814,
         n11815, n11816, n11817, n11818, n11819, n11820, n11821, n11822,
         n11823, n11824, n11825, n11826, n11827, n11828, n11829, n11830,
         n11831, n11832, n11833, n11834, n11835, n11836, n11837, n11838,
         n11839, n11840, n11841, n11842, n11843, n11844, n11845, n11846,
         n11847, n11848, n11849, n11850, n11851, n11852, n11853, n11854,
         n11855, n11856, n11857, n11858, n11859, n11860, n11861, n11862,
         n11863, n11864, n11865, n11866, n11867, n11868, n11869, n11870,
         n11871, n11872, n11873, n11874, n11875, n11876, n11877, n11878,
         n11879, n11880, n11881, n11882, n11883, n11884, n11885, n11886,
         n11887, n11888, n11889, n11890, n11891, n11892, n11893, n11894,
         n11895, n11896, n11897, n11898, n11899, n11900, n11901, n11902,
         n11903, n11904, n11905, n11906, n11907, n11908, n11909, n11910,
         n11911, n11912, n11913, n11914, n11915, n11916, n11917, n11918,
         n11919, n11920, n11921, n11922, n11923, n11924, n11925, n11926,
         n11927, n11928, n11929, n11930, n11931, n11932, n11933, n11934,
         n11935, n11936, n11937, n11938, n11939, n11940, n11941, n11942,
         n11943, n11944, n11945, n11946, n11947, n11948, n11949, n11950,
         n11951, n11952, n11953, n11954, n11955, n11956, n11957, n11958,
         n11959, n11960, n11961, n11962, n11963, n11964, n11965, n11966,
         n11967, n11968, n11969, n11970, n11971, n11972, n11973, n11974,
         n11975, n11976, n11977, n11978, n11979, n11980, n11981, n11982,
         n11983, n11984, n11985, n11986, n11987, n11988, n11989, n11990,
         n11991, n11992, n11993, n11994, n11995, n11996, n11997, n11998,
         n11999, n12000, n12001, n12002, n12003, n12004, n12005, n12006,
         n12007, n12008, n12009, n12010, n12011, n12012, n12013, n12014,
         n12015, n12016, n12017, n12018, n12019, n12020, n12021, n12022,
         n12023, n12024, n12025, n12026, n12027, n12028, n12029, n12030,
         n12031, n12032, n12033, n12034, n12035, n12036, n12037, n12038,
         n12039, n12040, n12041, n12042, n12043, n12044, n12045, n12046,
         n12047, n12048, n12049, n12050, n12051, n12052, n12053, n12054,
         n12055, n12056, n12057, n12058, n12059, n12060, n12061, n12062,
         n12063, n12064, n12065, n12066, n12067, n12068, n12069, n12070,
         n12071, n12072, n12073, n12074, n12075, n12076, n12077, n12078,
         n12079, n12080, n12081, n12082, n12083, n12084, n12085, n12086,
         n12087, n12088, n12089, n12090, n12091, n12092, n12093, n12094,
         n12095, n12096, n12097, n12098, n12099, n12100, n12101, n12102,
         n12103, n12104, n12105, n12106, n12107, n12108, n12109, n12110,
         n12111, n12112, n12113, n12114, n12115, n12116, n12117, n12118,
         n12119, n12120, n12121, n12122, n12123, n12124, n12125, n12126,
         n12127, n12128, n12129, n12130, n12131, n12132, n12133, n12134,
         n12135, n12136, n12137, n12138, n12139, n12140, n12141, n12142,
         n12143, n12144, n12145, n12146, n12147, n12148, n12149, n12150,
         n12151, n12152, n12153, n12154, n12155, n12156, n12157, n12158,
         n12159, n12160, n12161, n12162, n12163, n12164, n12165, n12166,
         n12167, n12168, n12169, n12170, n12171, n12172, n12173, n12174,
         n12175, n12176, n12177, n12178, n12179, n12180, n12181, n12182,
         n12183, n12184, n12185, n12186, n12187, n12188, n12189, n12190,
         n12191, n12192, n12193, n12194, n12195, n12196, n12197, n12198,
         n12199, n12200, n12201, n12202, n12203, n12204, n12205, n12206,
         n12207, n12208, n12209, n12210, n12211, n12212, n12213, n12214,
         n12215, n12216, n12217, n12218, n12219, n12220, n12221, n12222,
         n12223, n12224, n12225, n12226, n12227, n12228, n12229, n12230,
         n12231, n12232, n12233, n12234, n12235, n12236, n12237, n12238,
         n12239, n12240, n12241, n12242, n12243, n12244, n12245, n12246,
         n12247, n12248, n12249, n12250, n12251, n12252, n12253, n12254,
         n12255, n12256, n12257, n12258, n12259, n12260, n12261, n12262,
         n12263, n12264, n12265, n12266, n12267, n12268, n12269, n12270,
         n12271, n12272, n12273, n12274, n12275, n12276, n12277, n12278,
         n12279, n12280, n12281, n12282, n12283, n12284, n12285, n12286,
         n12287, n12288, n12289, n12290, n12291, n12292, n12293, n12294,
         n12295, n12296, n12297, n12298, n12299, n12300, n12301, n12302,
         n12303, n12304, n12305, n12306, n12307, n12308, n12309, n12310,
         n12311, n12312, n12313, n12314, n12315, n12316, n12317, n12318,
         n12319, n12320, n12321, n12322, n12323, n12324, n12325, n12326,
         n12327, n12328, n12329, n12330, n12331, n12332, n12333, n12334,
         n12335, n12336, n12337, n12338, n12339, n12340, n12341, n12342,
         n12343, n12344, n12345, n12346, n12347, n12348, n12349, n12350,
         n12351, n12352, n12353, n12354, n12355, n12356, n12357, n12358,
         n12359, n12360, n12361, n12362, n12363, n12364, n12365, n12366,
         n12367, n12368, n12369, n12370, n12371, n12372, n12373, n12374,
         n12375, n12376, n12377, n12378, n12379, n12380, n12381, n12382,
         n12383, n12384, n12385, n12386, n12387, n12388, n12389, n12390,
         n12391, n12392, n12393, n12394, n12395, n12396, n12397, n12398,
         n12399, n12400, n12401, n12402, n12403, n12404, n12405, n12406,
         n12407, n12408, n12409, n12410, n12411, n12412, n12413, n12414,
         n12415, n12416, n12417, n12418, n12419, n12420, n12421, n12422,
         n12423, n12424, n12425, n12426, n12427, n12428, n12429, n12430,
         n12431, n12432, n12433, n12434, n12435, n12436, n12437, n12438,
         n12439, n12440, n12441, n12442, n12443, n12444, n12445, n12446,
         n12447, n12448, n12449, n12450, n12451, n12452, n12453, n12454,
         n12455, n12456, n12457, n12458, n12459, n12460, n12461, n12462,
         n12463, n12464, n12465, n12466, n12467, n12468, n12469, n12470,
         n12471, n12472, n12473, n12474, n12475, n12476, n12477, n12478,
         n12479, n12480, n12481, n12482, n12483, n12484, n12485, n12486,
         n12487, n12488, n12489, n12490, n12491, n12492, n12493, n12494,
         n12495, n12496, n12497, n12498, n12499, n12500, n12501, n12502,
         n12503, n12504, n12505, n12506, n12507, n12508, n12509, n12510,
         n12511, n12512, n12513, n12514, n12515, n12516, n12517, n12518,
         n12519, n12520, n12521, n12522, n12523, n12524, n12525, n12526,
         n12527, n12528, n12529, n12530, n12531, n12532, n12533, n12534,
         n12535, n12536, n12537, n12538, n12539, n12540, n12541, n12542,
         n12543, n12544, n12545, n12546, n12547, n12548, n12549, n12550,
         n12551, n12552, n12553, n12554, n12555, n12556, n12557, n12558,
         n12559, n12560, n12561, n12562, n12563, n12564, n12565, n12566,
         n12567, n12568, n12569, n12570, n12571, n12572, n12573, n12574,
         n12575, n12576, n12577, n12578, n12579, n12580, n12581, n12582,
         n12583, n12584, n12585, n12586, n12587, n12588, n12589, n12590,
         n12591, n12592, n12593, n12594, n12595, n12596, n12597, n12598,
         n12599, n12600, n12601, n12602, n12603, n12604, n12605, n12606,
         n12607, n12608, n12609, n12610, n12611, n12612, n12613, n12614,
         n12615, n12616, n12617, n12618, n12619, n12620, n12621, n12622,
         n12623, n12624, n12625, n12626, n12627, n12628, n12629, n12630,
         n12631, n12632, n12633, n12634, n12635, n12636, n12637, n12638,
         n12639, n12640, n12641, n12642, n12643, n12644, n12645, n12646,
         n12647, n12648, n12649, n12650, n12651, n12652, n12653, n12654,
         n12655, n12656, n12657, n12658, n12659, n12660, n12661, n12662,
         n12663, n12664, n12665, n12666, n12667, n12668, n12669, n12670,
         n12671, n12672, n12673, n12674, n12675, n12676, n12677, n12678,
         n12679, n12680, n12681, n12682, n12683, n12684, n12685, n12686,
         n12687, n12688, n12689, n12690, n12691, n12692, n12693, n12694,
         n12695, n12696, n12697, n12698, n12699, n12700, n12701, n12702,
         n12703, n12704, n12705, n12706, n12707, n12708, n12709, n12710,
         n12711, n12712, n12713, n12714, n12715, n12716, n12717, n12718,
         n12719, n12720, n12721, n12722, n12723, n12724, n12725, n12726,
         n12727, n12728, n12729, n12730, n12731, n12732, n12733, n12734,
         n12735, n12736, n12737, n12738, n12739, n12740, n12741, n12742,
         n12743, n12744, n12745, n12746, n12747, n12748, n12749, n12750,
         n12751, n12752, n12753, n12754, n12755, n12756, n12757, n12758,
         n12759, n12760, n12761, n12762, n12763, n12764, n12765, n12766,
         n12767, n12768, n12769, n12770, n12771, n12772, n12773, n12774,
         n12775, n12776, n12777, n12778, n12779, n12780, n12781, n12782,
         n12783, n12784, n12785, n12786, n12787, n12788, n12789, n12790,
         n12791, n12792, n12793, n12794, n12795, n12796, n12797, n12798,
         n12799, n12800, n12801, n12802, n12803, n12804, n12805, n12806,
         n12807, n12808, n12809, n12810, n12811, n12812, n12813, n12814,
         n12815, n12816, n12817, n12818, n12819, n12820, n12821, n12822,
         n12823, n12824, n12825, n12826, n12827, n12828, n12829, n12830,
         n12831, n12832, n12833, n12834, n12835, n12836, n12837, n12838,
         n12839, n12840, n12841, n12842, n12843, n12844, n12845, n12846,
         n12847, n12848, n12849, n12850, n12851, n12852, n12853, n12854,
         n12855, n12856, n12857, n12858, n12859, n12860, n12861, n12862,
         n12863, n12864, n12865, n12866, n12867, n12868, n12869, n12870,
         n12871, n12872, n12873, n12874, n12875, n12876, n12877, n12878,
         n12879, n12880, n12881, n12882, n12883, n12884, n12885, n12886,
         n12887, n12888, n12889, n12890, n12891, n12892, n12893, n12894,
         n12895, n12896, n12897, n12898, n12899, n12900, n12901, n12902,
         n12903, n12904, n12905, n12906, n12907, n12908, n12909, n12910,
         n12911, n12912, n12913, n12914, n12915, n12916, n12917, n12918,
         n12919, n12920, n12921, n12922, n12923, n12924, n12925, n12926,
         n12927, n12928, n12929, n12930, n12931, n12932, n12933, n12934,
         n12935, n12936, n12937, n12938, n12939, n12940, n12941, n12942,
         n12943, n12944, n12945, n12946, n12947, n12948, n12949, n12950,
         n12951, n12952, n12953, n12954, n12955, n12956, n12957, n12958,
         n12959, n12960, n12961, n12962, n12963, n12964, n12965, n12966,
         n12967, n12968, n12969, n12970, n12971, n12972, n12973, n12974,
         n12975, n12976, n12977, n12978, n12979, n12980, n12981, n12982,
         n12983, n12984, n12985, n12986, n12987, n12988, n12989, n12990,
         n12991, n12992, n12993, n12994, n12995, n12996, n12997, n12998,
         n12999, n13000, n13001, n13002, n13003, n13004, n13005, n13006,
         n13007, n13008, n13009, n13010, n13011, n13012, n13013, n13014,
         n13015, n13016, n13017, n13018, n13019, n13020, n13021, n13022,
         n13023, n13024, n13025, n13026, n13027, n13028, n13029, n13030,
         n13031, n13032, n13033, n13034, n13035, n13036, n13037, n13038,
         n13039, n13040, n13041, n13042, n13043, n13044, n13045, n13046,
         n13047, n13048, n13049, n13050, n13051, n13052, n13053, n13054,
         n13055, n13056, n13057, n13058, n13059, n13060, n13061, n13062,
         n13063, n13064, n13065, n13066, n13067, n13068, n13069, n13070,
         n13071, n13072, n13073, n13074, n13075, n13076, n13077, n13078,
         n13079, n13080, n13081, n13082, n13083, n13084, n13085, n13086,
         n13087, n13088, n13089, n13090, n13091, n13092, n13093, n13094,
         n13095, n13096, n13097, n13098, n13099, n13100, n13101, n13102,
         n13103, n13104, n13105, n13106, n13107, n13108, n13109, n13110,
         n13111, n13112, n13113, n13114, n13115, n13116, n13117, n13118,
         n13119, n13120, n13121, n13122, n13123, n13124, n13125, n13126,
         n13127, n13128, n13129, n13130, n13131, n13132, n13133, n13134,
         n13135, n13136, n13137, n13138, n13139, n13140, n13141, n13142,
         n13143, n13144, n13145, n13146, n13147, n13148, n13149, n13150,
         n13151, n13152, n13153, n13154, n13155, n13156, n13157, n13158,
         n13159, n13160, n13161, n13162, n13163, n13164, n13165, n13166,
         n13167, n13168, n13169, n13170, n13171, n13172, n13173, n13174,
         n13175, n13176, n13177, n13178, n13179, n13180, n13181, n13182,
         n13183, n13184, n13185, n13186, n13187, n13188, n13189, n13190,
         n13191, n13192, n13193, n13194, n13195, n13196, n13197, n13198,
         n13199, n13200, n13201, n13202, n13203, n13204, n13205, n13206,
         n13207, n13208, n13209, n13210, n13211, n13212, n13213, n13214,
         n13215, n13216, n13217, n13218, n13219, n13220, n13221, n13222,
         n13223, n13224, n13225, n13226, n13227, n13228, n13229, n13230,
         n13231, n13232, n13233, n13234, n13235, n13236, n13237, n13238,
         n13239, n13240, n13241, n13242, n13243, n13244, n13245, n13246,
         n13247, n13248, n13249, n13250, n13251, n13252, n13253, n13254,
         n13255, n13256, n13257, n13258, n13259, n13260, n13261, n13262,
         n13263, n13264, n13265, n13266, n13267, n13268, n13269, n13270,
         n13271, n13272, n13273, n13274, n13275, n13276, n13277, n13278,
         n13279, n13280, n13281, n13282, n13283, n13284, n13285, n13286,
         n13287, n13288, n13289, n13290, n13291, n13292, n13293, n13294,
         n13295, n13296, n13297, n13298, n13299, n13300, n13301, n13302,
         n13303, n13304, n13305, n13306, n13307, n13308, n13309, n13310,
         n13311, n13312, n13313, n13314, n13315, n13316, n13317, n13318,
         n13319, n13320, n13321, n13322, n13323, n13324, n13325, n13326,
         n13327, n13328, n13329, n13330, n13331, n13332, n13333, n13334,
         n13335, n13336, n13337, n13338, n13339, n13340, n13341, n13342,
         n13343, n13344, n13345, n13346, n13347, n13348, n13349, n13350,
         n13351, n13352, n13353, n13354, n13355, n13356, n13357, n13358,
         n13359, n13360, n13361, n13362, n13363, n13364, n13365, n13366,
         n13367, n13368, n13369, n13370, n13371, n13372, n13373, n13374,
         n13375, n13376, n13377, n13378, n13379, n13380, n13381, n13382,
         n13383, n13384, n13385, n13386, n13387, n13388, n13389, n13390,
         n13391, n13392, n13393, n13394, n13395, n13396, n13397, n13398,
         n13399, n13400, n13401, n13402, n13403, n13404, n13405, n13406,
         n13407, n13408, n13409, n13410, n13411, n13412, n13413, n13414,
         n13415, n13416, n13417, n13418, n13419, n13420, n13421, n13422,
         n13423, n13424, n13425, n13426, n13427, n13428, n13429, n13430,
         n13431, n13432, n13433, n13434, n13435, n13436, n13437, n13438,
         n13439, n13440, n13441, n13442, n13443, n13444, n13445, n13446,
         n13447, n13448, n13449, n13450, n13451, n13452, n13453, n13454,
         n13455, n13456, n13457, n13458, n13459, n13460, n13461, n13462,
         n13463, n13464, n13465, n13466, n13467, n13468, n13469, n13470,
         n13471, n13472, n13473, n13474, n13475, n13476, n13477, n13478,
         n13479, n13480, n13481, n13482, n13483, n13484, n13485, n13486,
         n13487, n13488, n13489, n13490, n13491, n13492, n13493, n13494,
         n13495, n13496, n13497, n13498, n13499, n13500, n13501, n13502,
         n13503, n13504, n13505, n13506, n13507, n13508, n13509, n13510,
         n13511, n13512, n13513, n13514, n13515, n13516, n13517, n13518,
         n13519, n13520, n13521, n13522, n13523, n13524, n13525, n13526,
         n13527, n13528, n13529, n13530, n13531, n13532, n13533, n13534,
         n13535, n13536, n13537, n13538, n13539, n13540, n13541, n13542,
         n13543, n13544, n13545, n13546, n13547, n13548, n13549, n13550,
         n13551, n13552, n13553, n13554, n13555, n13556, n13557, n13558,
         n13559, n13560, n13561, n13562, n13563, n13564, n13565, n13566,
         n13567, n13568, n13569, n13570, n13571, n13572, n13573, n13574,
         n13575, n13576, n13577, n13578, n13579, n13580, n13581, n13582,
         n13583, n13584, n13585, n13586, n13587, n13588, n13589, n13590,
         n13591, n13592, n13593, n13594, n13595, n13596, n13597, n13598,
         n13599, n13600, n13601, n13602, n13603, n13604, n13605, n13606,
         n13607, n13608, n13609, n13610, n13611, n13612, n13613, n13614,
         n13615, n13616, n13617, n13618, n13619, n13620, n13621, n13622,
         n13623, n13624, n13625, n13626, n13627, n13628, n13629, n13630,
         n13631, n13632, n13633, n13634, n13635, n13636, n13637, n13638,
         n13639, n13640, n13641, n13642, n13643, n13644, n13645, n13646,
         n13647, n13648, n13649, n13650, n13651, n13652, n13653, n13654,
         n13655, n13656, n13657, n13658, n13659, n13660, n13661, n13662,
         n13663, n13664, n13665, n13666, n13667, n13668, n13669, n13670,
         n13671, n13672, n13673, n13674, n13675, n13676, n13677, n13678,
         n13679, n13680, n13681, n13682, n13683, n13684, n13685, n13686,
         n13687, n13688, n13689, n13690, n13691, n13692, n13693, n13694,
         n13695, n13696, n13697, n13698, n13699, n13700, n13701, n13702,
         n13703, n13704, n13705, n13706, n13707, n13708, n13709, n13710,
         n13711, n13712, n13713, n13714, n13715, n13716, n13717, n13718,
         n13719, n13720, n13721, n13722, n13723, n13724, n13725, n13726,
         n13727, n13728, n13729, n13730, n13731, n13732, n13733, n13734,
         n13735, n13736, n13737, n13738, n13739, n13740, n13741, n13742,
         n13743, n13744, n13745, n13746, n13747, n13748, n13749, n13750,
         n13751, n13752, n13753, n13754, n13755, n13756, n13757, n13758,
         n13759, n13760, n13761, n13762, n13763, n13764, n13765, n13766,
         n13767, n13768, n13769, n13770, n13771, n13772, n13773, n13774,
         n13775, n13776, n13777, n13778, n13779, n13780, n13781, n13782,
         n13783, n13784, n13785, n13786, n13787, n13788, n13789, n13790,
         n13791, n13792, n13793, n13794, n13795, n13796, n13797, n13798,
         n13799, n13800, n13801, n13802, n13803, n13804, n13805, n13806,
         n13807, n13808, n13809, n13810, n13811, n13812, n13813, n13814,
         n13815, n13816, n13817, n13818, n13819, n13820, n13821, n13822,
         n13823, n13824, n13825, n13826, n13827, n13828, n13829, n13830,
         n13831, n13832, n13833, n13834, n13835, n13836, n13837, n13839,
         n13840, n13841, n13842, n13843, n13844, n13845, n13846, n13847,
         n13848, n13849, n13850, n13851, n13852, n13853, n13854, n13855,
         n13856, n13857, n13858, n13859, n13860, n13861, n13862, n13863,
         n13864, n13865, n13866, n13867, n13868, n13869, n13870, n13871,
         n13872, n13873, n13874, n13875, n13876, n13877, n13878, n13879,
         n13880, n13881, n13882, n13883, n13884, n13885, n13886, n13887,
         n13888, n13889, n13890, n13891, n13892, n13893, n13894, n13895,
         n13896, n13897, n13898, n13899, n13900, n13901, n13902, n13903,
         n13904, n13905, n13906, n13907, n13908, n13909, n13910, n13911,
         n13912, n13913, n13914, n13915, n13916, n13917, n13918, n13919,
         n13920, n13921, n13922, n13923, n13924, n13925, n13926, n13927,
         n13928, n13929, n13930, n13931, n13932, n13933, n13934, n13935,
         n13936, n13937, n13938, n13939, n13940, n13941, n13942, n13943,
         n13944, n13945, n13946, n13947, n13948, n13949, n13950, n13951,
         n13952, n13953, n13954, n13955, n13956, n13957, n13958, n13959,
         n13960, n13961, n13962, n13963, n13964, n13965, n13966, n13967,
         n13968, n13969, n13970, n13971, n13972, n13973, n13974, n13975,
         n13976, n13977, n13978, n13979, n13980, n13981, n13982, n13983,
         n13984, n13985, n13986, n13987, n13988, n13989, n13990, n13991,
         n13992, n13993, n13994, n13995, n13996, n13997, n13998, n13999,
         n14000, n14001, n14002, n14003, n14004, n14005, n14006, n14007,
         n14008, n14009, n14010, n14011, n14012, n14013, n14014, n14015,
         n14016, n14017, n14018, n14019, n14020, n14021, n14022, n14023,
         n14024, n14025, n14026, n14027, n14028, n14029, n14030, n14031,
         n14032, n14033, n14034, n14035, n14036, n14037, n14038, n14039,
         n14040, n14041, n14042, n14043, n14044, n14045, n14046, n14047,
         n14048, n14049, n14050, n14051, n14052, n14053, n14054, n14055,
         n14056, n14057, n14058, n14059, n14060, n14061, n14062, n14063,
         n14064, n14065, n14066, n14067, n14068, n14069, n14070, n14071,
         n14072, n14073, n14074, n14075, n14076, n14077, n14078, n14079,
         n14080, n14081, n14082, n14083, n14084, n14085, n14086, n14087,
         n14088, n14089, n14090, n14091, n14092, n14093, n14094, n14095,
         n14096, n14097, n14098, n14099, n14100, n14101, n14102, n14103,
         n14104, n14105, n14106, n14107, n14108, n14109, n14110, n14111,
         n14112, n14113, n14114, n14115, n14116, n14117, n14118, n14119,
         n14120, n14121, n14122, n14123, n14124, n14125, n14126, n14127,
         n14128, n14129, n14130, n14131, n14132, n14133, n14134, n14135,
         n14136, n14137, n14138, n14139, n14140, n14141, n14142, n14143,
         n14144, n14145, n14146, n14147, n14148, n14149, n14150, n14151,
         n14152, n14153, n14154, n14155, n14156, n14157, n14158, n14159,
         n14160, n14161, n14162, n14163, n14164, n14165, n14166, n14167,
         n14168, n14169, n14170, n14171, n14172, n14173, n14174, n14175,
         n14176, n14177, n14178, n14179, n14180, n14181, n14182, n14183,
         n14184, n14185, n14186, n14187, n14188, n14189, n14190, n14191,
         n14192, n14193, n14194, n14195, n14196, n14197, n14198, n14199,
         n14200, n14201, n14202, n14203, n14204, n14205, n14206, n14207,
         n14208, n14209, n14210, n14211, n14212, n14213, n14214, n14215,
         n14216, n14217, n14218, n14219, n14220, n14221, n14222, n14223,
         n14224, n14225, n14226, n14227, n14228, n14229, n14230, n14231,
         n14232, n14233, n14234, n14235, n14236, n14237, n14238, n14239,
         n14240, n14241, n14242, n14243, n14244, n14245, n14246, n14247,
         n14248, n14249, n14250, n14251, n14252, n14253, n14254, n14255,
         n14256, n14257, n14258, n14259, n14260, n14261, n14262, n14263,
         n14264, n14265, n14266, n14267, n14268, n14269, n14270, n14271,
         n14272, n14273, n14274, n14275, n14276, n14277, n14278, n14279,
         n14280, n14281, n14282, n14283, n14284, n14285, n14286, n14287,
         n14288, n14289, n14290, n14291, n14292, n14293, n14294, n14295,
         n14296, n14297, n14298, n14299, n14300, n14301, n14302, n14303,
         n14304, n14305, n14306, n14307, n14308, n14309, n14310, n14311,
         n14312, n14313, n14314, n14315, n14316, n14317, n14318, n14319,
         n14320, n14321, n14322, n14323, n14324, n14325, n14326, n14327,
         n14328, n14329, n14330, n14331, n14332, n14333, n14334, n14335,
         n14336, n14337, n14338, n14339, n14340, n14341, n14342, n14343,
         n14344, n14345, n14346, n14347, n14348, n14349, n14350, n14351,
         n14352, n14353, n14354, n14355, n14356, n14357, n14358, n14359,
         n14360, n14361, n14362, n14363, n14364, n14365, n14366, n14367,
         n14368, n14369, n14370, n14371, n14372, n14373, n14374, n14375,
         n14376, n14377, n14378, n14379, n14380, n14381, n14382, n14383,
         n14384, n14385, n14386, n14387, n14388, n14389, n14390, n14391,
         n14392, n14393, n14394, n14395, n14396, n14397, n14398, n14399,
         n14400, n14401, n14402, n14403, n14404, n14405, n14406, n14407,
         n14408, n14409, n14410, n14411, n14412, n14413, n14414, n14415,
         n14416, n14417, n14418, n14419, n14420, n14421, n14422, n14423,
         n14424, n14425, n14426, n14427, n14428, n14429, n14430, n14431,
         n14432, n14433, n14434, n14435, n14436, n14437, n14438, n14439,
         n14440, n14441, n14442, n14443, n14444, n14445, n14446, n14447,
         n14448, n14449, n14450, n14451, n14452, n14453, n14454, n14455,
         n14456, n14457, n14458, n14459, n14460, n14461, n14462, n14463,
         n14464, n14465, n14466, n14467, n14468, n14469, n14470, n14471,
         n14472, n14473, n14474, n14475, n14476, n14477, n14478, n14479,
         n14480, n14481, n14482, n14483, n14484, n14485, n14486, n14487,
         n14488, n14489, n14490, n14491, n14492, n14493, n14494, n14495,
         n14496, n14497, n14498, n14499, n14500, n14501, n14502, n14503,
         n14504, n14505, n14506, n14507, n14508, n14509, n14510, n14511,
         n14512, n14513, n14514, n14515, n14516, n14517, n14518, n14519,
         n14520, n14521, n14522, n14523, n14524, n14525, n14526, n14527,
         n14528, n14529, n14530, n14531, n14532, n14533, n14534, n14535,
         n14536, n14537, n14538, n14539, n14540, n14541, n14542, n14543,
         n14544, n14545, n14546, n14547, n14548, n14549, n14550, n14551,
         n14552, n14553, n14554, n14555, n14556, n14557, n14558, n14559,
         n14560, n14561, n14562, n14563, n14564, n14565, n14566, n14567,
         n14568, n14569, n14570, n14571, n14572, n14573, n14574, n14575,
         n14576, n14577, n14578, n14579, n14580, n14581, n14582, n14583,
         n14584, n14585, n14586, n14587, n14588, n14589, n14590, n14591,
         n14592, n14593, n14594, n14595, n14596, n14597, n14598, n14599,
         n14600, n14601, n14602, n14603, n14604, n14605, n14606, n14607,
         n14608, n14609, n14610, n14611, n14612, n14613, n14614, n14615,
         n14616, n14617, n14618, n14619, n14620, n14621, n14622, n14623,
         n14624, n14625, n14626, n14627, n14628, n14629, n14630, n14631,
         n14632, n14633, n14634, n14635, n14636, n14637, n14638, n14639,
         n14640, n14641, n14642, n14643, n14644, n14645, n14646, n14647,
         n14648, n14649, n14650, n14651, n14652, n14653, n14654, n14655,
         n14656, n14657, n14658, n14659, n14660, n14661, n14662, n14663,
         n14664, n14665, n14666, n14667, n14668, n14669, n14670, n14671,
         n14672, n14673, n14674, n14675, n14676, n14677, n14678, n14679,
         n14680, n14681, n14682, n14683, n14684, n14685, n14686, n14687,
         n14688, n14689, n14690, n14691, n14692, n14693, n14694, n14695,
         n14696, n14697, n14698, n14699, n14700, n14701, n14702, n14703,
         n14704, n14705, n14706, n14707, n14708, n14709, n14710, n14711,
         n14712, n14713, n14714, n14715, n14716, n14717, n14718, n14719,
         n14720, n14721, n14722, n14723, n14724, n14725, n14726, n14727,
         n14728, n14729, n14730, n14731, n14732, n14733, n14734, n14735,
         n14736, n14737, n14738, n14739, n14740, n14741, n14742, n14743,
         n14744, n14745, n14746, n14747, n14748, n14749, n14750, n14751,
         n14752, n14753, n14754, n14755, n14756, n14757, n14758, n14759,
         n14760, n14761, n14762, n14763, n14764, n14765, n14766, n14767,
         n14768, n14769, n14770, n14771, n14772, n14773, n14774, n14775,
         n14776, n14777, n14778, n14779, n14780, n14781, n14782, n14783,
         n14784, n14785, n14786, n14787, n14788, n14789, n14790, n14791,
         n14792, n14793, n14794, n14795, n14796, n14797, n14798, n14799,
         n14800, n14801, n14802, n14803, n14804, n14805, n14806, n14807,
         n14808, n14809, n14810, n14811, n14812, n14813, n14814, n14815,
         n14816, n14817, n14818, n14819, n14820, n14821, n14822, n14823,
         n14824, n14825, n14826, n14827, n14828, n14829, n14830, n14831,
         n14832, n14833, n14834, n14835, n14836, n14837, n14838, n14839,
         n14840, n14841, n14842, n14843, n14844, n14845, n14846, n14847,
         n14848, n14849, n14850, n14851, n14852, n14853, n14854, n14855,
         n14856, n14857, n14858, n14859, n14860, n14861, n14862, n14863,
         n14864, n14865, n14866, n14867, n14868, n14869, n14870, n14871,
         n14872, n14873, n14874, n14875, n14876, n14877, n14878, n14879,
         n14880, n14881, n14882, n14883, n14884, n14885, n14886, n14887,
         n14888, n14889, n14890, n14891, n14892, n14893, n14894, n14895,
         n14896, n14897, n14898, n14899, n14900, n14901, n14902, n14903,
         n14904, n14905, n14906, n14907, n14908, n14909, n14910, n14911,
         n14912, n14913, n14914, n14915, n14916, n14917, n14918, n14919,
         n14920, n14921, n14922, n14923, n14924, n14925, n14926, n14927,
         n14928, n14929, n14930, n14931, n14932, n14933, n14934, n14935,
         n14936, n14937, n14938, n14939, n14940, n14941, n14942, n14943,
         n14944, n14945, n14946, n14947, n14948, n14949, n14950, n14951,
         n14952, n14953, n14954, n14955, n14956, n14957, n14958, n14959,
         n14960, n14961, n14962, n14963, n14964, n14965, n14966, n14967,
         n14968, n14969, n14970, n14971, n14972, n14973, n14974, n14975,
         n14976, n14977, n14978, n14979, n14980, n14981, n14982, n14983,
         n14984, n14985, n14986, n14987, n14988, n14989, n14990, n14991,
         n14992, n14993, n14994, n14995, n14996, n14997, n14998, n14999,
         n15000, n15001, n15002, n15003, n15004, n15005, n15006, n15007,
         n15008, n15009, n15010, n15011, n15012, n15013, n15014, n15015,
         n15016, n15017, n15018, n15019, n15020, n15021, n15022, n15023,
         n15024, n15025, n15026, n15027, n15028, n15029, n15030, n15031,
         n15032, n15033, n15034, n15035, n15036, n15037, n15038, n15039,
         n15040, n15041, n15042, n15043, n15044, n15045, n15046, n15047,
         n15048, n15049, n15050, n15051, n15052, n15053, n15054, n15055,
         n15056, n15057, n15058, n15059, n15060, n15061, n15062, n15063,
         n15064, n15065, n15066, n15067, n15068, n15069, n15070, n15071,
         n15072, n15073, n15074, n15075, n15076, n15077, n15078, n15079,
         n15080, n15081, n15082, n15083, n15084, n15085, n15086, n15087,
         n15088, n15089, n15090, n15091, n15092, n15093, n15094, n15095,
         n15096, n15097, n15098, n15099, n15100, n15101, n15102, n15103,
         n15104, n15105, n15106, n15107, n15108, n15109, n15110, n15111,
         n15112, n15113, n15114, n15115, n15116, n15117, n15118, n15119,
         n15120, n15121, n15122, n15123, n15124, n15125, n15126, n15127,
         n15128, n15129, n15130, n15131, n15132, n15133, n15134, n15135,
         n15136, n15137, n15138, n15139, n15140, n15141, n15142, n15143,
         n15144, n15145, n15146, n15147, n15148, n15149, n15150, n15151,
         n15152, n15153, n15154, n15155, n15156, n15157, n15158, n15159,
         n15160, n15161, n15162, n15163, n15164, n15165, n15166, n15167,
         n15168, n15169, n15170, n15171, n15172, n15173, n15174, n15175,
         n15176, n15177, n15178, n15179, n15180, n15181, n15182, n15183,
         n15184, n15185, n15186, n15187, n15188, n15189, n15190, n15191,
         n15192, n15193, n15194, n15195, n15196, n15197, n15198, n15199,
         n15200, n15201, n15202, n15203, n15204, n15205, n15206, n15207,
         n15208, n15209, n15210, n15211, n15212, n15213, n15214, n15215,
         n15216, n15217, n15218, n15219, n15220, n15221, n15222, n15223,
         n15224, n15225, n15226, n15227, n15228, n15229, n15230, n15231,
         n15232, n15233, n15234, n15235, n15236, n15237, n15238, n15239,
         n15240, n15241, n15242, n15243, n15244, n15245, n15246, n15247,
         n15248, n15249, n15250, n15251, n15252, n15253, n15254, n15255,
         n15256, n15257, n15258, n15259, n15260, n15261, n15262, n15263,
         n15264, n15265, n15266, n15267, n15268, n15269, n15270, n15271,
         n15272, n15273, n15274, n15275, n15276, n15277, n15278, n15279,
         n15280, n15281, n15282, n15283, n15284, n15285, n15286, n15287,
         n15288, n15289, n15290, n15291, n15292, n15293, n15294, n15295,
         n15296, n15297, n15298, n15299, n15300, n15301, n15302, n15303,
         n15304, n15305, n15306, n15307, n15308, n15309, n15310, n15311,
         n15312, n15313, n15314, n15315, n15316, n15317, n15318, n15319,
         n15320, n15321, n15322, n15323, n15324, n15325, n15326, n15327,
         n15328, n15329, n15330, n15331, n15332, n15333, n15334, n15335,
         n15336, n15337, n15338, n15339, n15340, n15341, n15342, n15343,
         n15344, n15345, n15346, n15347, n15348, n15349, n15350, n15351,
         n15352, n15353, n15354, n15355, n15356, n15357, n15358, n15359,
         n15360, n15361, n15362, n15363, n15364, n15365, n15366, n15367,
         n15368, n15369, n15370, n15371, n15372, n15373, n15374, n15375,
         n15376, n15377, n15378, n15379, n15380, n15381, n15382, n15383,
         n15384, n15385, n15386, n15387, n15388, n15389, n15390, n15391,
         n15392, n15393, n15394, n15395, n15396, n15397, n15398, n15399,
         n15400, n15401, n15402, n15403, n15404, n15405, n15406, n15407,
         n15408, n15409, n15410, n15411, n15412, n15413, n15414, n15415,
         n15416, n15417, n15418, n15419, n15420, n15421, n15422, n15423,
         n15424, n15425, n15426, n15427, n15428, n15429, n15430, n15431,
         n15432, n15433, n15434, n15435, n15436, n15437, n15438, n15439,
         n15440, n15441, n15442, n15443, n15444, n15445, n15446, n15447,
         n15448, n15449, n15450, n15451, n15452, n15453, n15454, n15455,
         n15456, n15457, n15458, n15459, n15460, n15461, n15462, n15463,
         n15464, n15465, n15466, n15467, n15468, n15469, n15470, n15471,
         n15472, n15473, n15474, n15475, n15476, n15477, n15478, n15479,
         n15480, n15481, n15482, n15483, n15484, n15485, n15486, n15487,
         n15488, n15489, n15490, n15491, n15492, n15493, n15494, n15495,
         n15496, n15497, n15498, n15499, n15500, n15501, n15502, n15503,
         n15504, n15505, n15506, n15507, n15508, n15509, n15510, n15511,
         n15512, n15513, n15514, n15515, n15516, n15517, n15518, n15519,
         n15520, n15521, n15522, n15523, n15524, n15525, n15526, n15527,
         n15528, n15529, n15530, n15531, n15532, n15533, n15534, n15535,
         n15536, n15537, n15538, n15539, n15540, n15541, n15542, n15543,
         n15544, n15545, n15546, n15547, n15548, n15549, n15550, n15551,
         n15552, n15553, n15554, n15555, n15556, n15557, n15558, n15559,
         n15560, n15561, n15562, n15563, n15564, n15565, n15566, n15567,
         n15568, n15569, n15570, n15571, n15572, n15573, n15574, n15575,
         n15576, n15577, n15578, n15579, n15580, n15581, n15582, n15583,
         n15584, n15585, n15586, n15587, n15588, n15589, n15590, n15591,
         n15592, n15593, n15594, n15595, n15596, n15597, n15598, n15599,
         n15600, n15601, n15602, n15603, n15604, n15605, n15606, n15607,
         n15608, n15609, n15610, n15611, n15612, n15613, n15614, n15615,
         n15616, n15617, n15618, n15619, n15620, n15621, n15622, n15623,
         n15624, n15625, n15626, n15627, n15628, n15629, n15630, n15631,
         n15632, n15633, n15634, n15635, n15636, n15637, n15638, n15639,
         n15640, n15641, n15642, n15643, n15644, n15645, n15646, n15647,
         n15648, n15649, n15650, n15651, n15652, n15653, n15654, n15655,
         n15656, n15657, n15658, n15659, n15660, n15661, n15662, n15663,
         n15664, n15665, n15666, n15667, n15668, n15669, n15670, n15671,
         n15672, n15673, n15674, n15675, n15676, n15677, n15678, n15679,
         n15680, n15681, n15682, n15683, n15684, n15685, n15686, n15687,
         n15688, n15689, n15690, n15691, n15692, n15693, n15694, n15695,
         n15696, n15697, n15698, n15699, n15700, n15701, n15702, n15703,
         n15704, n15705, n15706, n15707, n15708, n15709, n15710, n15711,
         n15712, n15713, n15714, n15715, n15716, n15717, n15718, n15719,
         n15720, n15721, n15722, n15723, n15724, n15725, n15726, n15727,
         n15728, n15729, n15730, n15731, n15732, n15733, n15734, n15735,
         n15736, n15737, n15738, n15739, n15740, n15741, n15742, n15743,
         n15744, n15745, n15746, n15747, n15748, n15749, n15750, n15751,
         n15752, n15753, n15754, n15755, n15756, n15757, n15758, n15759,
         n15760, n15761, n15762, n15763, n15764, n15765, n15766, n15767,
         n15768, n15769, n15770, n15771, n15772, n15773, n15774, n15775,
         n15776, n15777, n15778, n15779, n15780, n15781, n15782, n15783,
         n15784, n15785, n15786, n15787, n15788, n15789, n15790, n15791,
         n15792, n15793, n15794, n15795, n15796, n15797, n15798, n15799,
         n15800, n15801;

  INV_X2 U7413 ( .A(n14206), .ZN(n6670) );
  AND2_X1 U7414 ( .A1(n11285), .A2(n10999), .ZN(n10746) );
  INV_X2 U7415 ( .A(n9851), .ZN(n6921) );
  NAND2_X2 U7416 ( .A1(n8441), .A2(n8440), .ZN(n15671) );
  INV_X2 U7418 ( .A(n9388), .ZN(n9479) );
  INV_X1 U7419 ( .A(n9695), .ZN(n11053) );
  AND4_X1 U7420 ( .A1(n9056), .A2(n9055), .A3(n9054), .A4(n9053), .ZN(n11224)
         );
  BUF_X1 U7421 ( .A(n8322), .Z(n8508) );
  AND2_X1 U7422 ( .A1(n9018), .A2(n13842), .ZN(n9089) );
  NAND2_X2 U7423 ( .A1(n9033), .A2(n9032), .ZN(n10826) );
  AND2_X2 U7424 ( .A1(n13837), .A2(n13842), .ZN(n9138) );
  NAND2_X1 U7425 ( .A1(n15092), .A2(n15085), .ZN(n12597) );
  INV_X1 U7426 ( .A(n10746), .ZN(n9771) );
  AND2_X1 U7428 ( .A1(n9290), .A2(n9289), .ZN(n9294) );
  INV_X2 U7429 ( .A(n8369), .ZN(n8382) );
  AND2_X1 U7430 ( .A1(n11022), .A2(n11021), .ZN(n11081) );
  CLKBUF_X2 U7433 ( .A(n10829), .Z(n13254) );
  NAND2_X1 U7434 ( .A1(n9656), .A2(n9657), .ZN(n13567) );
  NAND2_X1 U7435 ( .A1(n9015), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9017) );
  OAI21_X1 U7436 ( .B1(n8558), .B2(n7025), .A(n7023), .ZN(n12128) );
  NAND2_X1 U7437 ( .A1(n6726), .A2(n6730), .ZN(n7012) );
  NOR2_X1 U7438 ( .A1(n13878), .A2(n8784), .ZN(n13949) );
  INV_X1 U7439 ( .A(n12448), .ZN(n12415) );
  INV_X1 U7440 ( .A(n6666), .ZN(n6680) );
  NAND2_X2 U7441 ( .A1(n10187), .A2(n9941), .ZN(n12448) );
  INV_X1 U7442 ( .A(n12609), .ZN(n11544) );
  OAI21_X1 U7443 ( .B1(n8660), .B2(n7677), .A(n8285), .ZN(n8678) );
  XNOR2_X1 U7444 ( .A(n8257), .B(SI_8_), .ZN(n8468) );
  NAND2_X1 U7445 ( .A1(n13949), .A2(n13948), .ZN(n13947) );
  NAND2_X1 U7446 ( .A1(n8398), .A2(n8397), .ZN(n15659) );
  NAND3_X1 U7447 ( .A1(n8368), .A2(n8367), .A3(n8366), .ZN(n12882) );
  NAND2_X1 U7448 ( .A1(n12257), .A2(n12256), .ZN(n12255) );
  OAI211_X2 U7449 ( .C1(n10076), .C2(n10261), .A(n8348), .B(n8347), .ZN(n8886)
         );
  NAND2_X1 U7450 ( .A1(n14960), .A2(n12545), .ZN(n14937) );
  AOI21_X1 U7451 ( .B1(n9737), .B2(n15722), .A(n9736), .ZN(n13174) );
  NAND2_X1 U7452 ( .A1(n13947), .A2(n7036), .ZN(n12847) );
  OAI21_X1 U7453 ( .B1(n7064), .B2(n7063), .A(n9848), .ZN(n12593) );
  NAND2_X1 U7454 ( .A1(n9844), .A2(n9850), .ZN(n14553) );
  XOR2_X1 U7455 ( .A(n13155), .B(n8859), .Z(n6665) );
  INV_X1 U7456 ( .A(n9138), .ZN(n9070) );
  NAND2_X1 U7457 ( .A1(n9821), .A2(n15234), .ZN(n6666) );
  INV_X2 U7458 ( .A(n12888), .ZN(n12891) );
  AOI21_X2 U7459 ( .B1(n8346), .B2(n8345), .A(n8238), .ZN(n8239) );
  NAND2_X2 U7460 ( .A1(n13419), .A2(n13418), .ZN(n13438) );
  NOR2_X4 U7461 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n8342) );
  NAND2_X2 U7462 ( .A1(n10947), .A2(n6763), .ZN(n12620) );
  NAND2_X1 U7463 ( .A1(n12866), .A2(n12863), .ZN(n13120) );
  OAI222_X1 U7464 ( .A1(n12861), .A2(n10531), .B1(n14396), .B2(n9980), .C1(
        P2_U3088), .C2(n10166), .ZN(P2_U3324) );
  OAI222_X1 U7465 ( .A1(n14750), .A2(P1_U3086), .B1(n15238), .B2(n9980), .C1(
        n9963), .C2(n15239), .ZN(P1_U3352) );
  OR2_X1 U7466 ( .A1(n9980), .A2(n9889), .ZN(n9842) );
  OAI21_X2 U7467 ( .B1(n12575), .B2(n12574), .A(n12573), .ZN(n12576) );
  OAI222_X1 U7468 ( .A1(P1_U3086), .A2(n9941), .B1(n15238), .B2(n15237), .C1(
        n15236), .C2(n15239), .ZN(P1_U3327) );
  AOI21_X2 U7469 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(n7839), .A(n15297), .ZN(
        n15247) );
  NAND2_X2 U7470 ( .A1(n11322), .A2(n11323), .ZN(n11458) );
  OAI22_X2 U7471 ( .A1(n11319), .A2(n11318), .B1(n11317), .B2(n11331), .ZN(
        n11322) );
  XNOR2_X2 U7472 ( .A(n9243), .B(P2_DATAO_REG_13__SCAN_IN), .ZN(n9242) );
  AOI22_X1 U7473 ( .A1(n8680), .A2(P1_DATAO_REG_4__SCAN_IN), .B1(n8679), .B2(
        n10309), .ZN(n8397) );
  NAND2_X2 U7474 ( .A1(n9816), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9818) );
  NAND4_X2 U7475 ( .A1(n9038), .A2(n9037), .A3(n9036), .A4(n9035), .ZN(n9512)
         );
  NAND2_X2 U7476 ( .A1(n9835), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9832) );
  INV_X1 U7477 ( .A(n14557), .ZN(n6676) );
  NOR2_X2 U7478 ( .A1(n9081), .A2(P3_IR_REG_4__SCAN_IN), .ZN(n9080) );
  BUF_X4 U7479 ( .A(n14553), .Z(n6667) );
  INV_X1 U7480 ( .A(n9474), .ZN(n6668) );
  INV_X2 U7481 ( .A(n9474), .ZN(n9184) );
  OAI222_X1 U7482 ( .A1(P1_U3086), .A2(n15234), .B1(n15238), .B2(n15233), .C1(
        n15232), .C2(n15239), .ZN(P1_U3326) );
  AND2_X1 U7483 ( .A1(n9820), .A2(n15234), .ZN(n6878) );
  NOR2_X4 U7484 ( .A1(n9820), .A2(n15234), .ZN(n9865) );
  INV_X2 U7485 ( .A(n9821), .ZN(n9820) );
  OAI21_X2 U7486 ( .B1(n14120), .B2(n7429), .A(n7427), .ZN(n14085) );
  NAND2_X2 U7487 ( .A1(n14139), .A2(n8929), .ZN(n14120) );
  NOR2_X2 U7488 ( .A1(n8859), .A2(n13156), .ZN(n12871) );
  NOR4_X1 U7489 ( .A1(n13602), .A2(n13567), .A3(n13615), .A4(n9521), .ZN(n9522) );
  BUF_X4 U7490 ( .A(n9435), .Z(n6678) );
  AOI21_X2 U7491 ( .B1(n8454), .B2(n8256), .A(n8468), .ZN(n7685) );
  XNOR2_X2 U7492 ( .A(n8255), .B(SI_7_), .ZN(n8454) );
  OAI211_X1 U7494 ( .C1(n12448), .C2(n14734), .A(n9891), .B(n9890), .ZN(n12609) );
  NAND2_X4 U7495 ( .A1(n8992), .A2(n8326), .ZN(n8369) );
  MUX2_X2 U7496 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9030), .S(
        P3_IR_REG_1__SCAN_IN), .Z(n9033) );
  AOI21_X1 U7497 ( .B1(n13313), .B2(n13630), .A(n13206), .ZN(n13210) );
  NAND2_X1 U7498 ( .A1(n7243), .A2(n7242), .ZN(n15024) );
  OR2_X1 U7499 ( .A1(n9420), .A2(n7116), .ZN(n7115) );
  NAND2_X1 U7500 ( .A1(n14634), .A2(n7394), .ZN(n15377) );
  BUF_X1 U7501 ( .A(n13549), .Z(n6675) );
  NAND2_X1 U7502 ( .A1(n11398), .A2(n11397), .ZN(n12641) );
  NAND2_X1 U7503 ( .A1(n10936), .A2(n15727), .ZN(n15733) );
  NAND2_X1 U7504 ( .A1(n8422), .A2(n8421), .ZN(n12907) );
  CLKBUF_X2 U7505 ( .A(P2_U3947), .Z(n6672) );
  NAND2_X1 U7506 ( .A1(n10625), .A2(n15747), .ZN(n9554) );
  INV_X2 U7507 ( .A(n10829), .ZN(n13207) );
  CLKBUF_X1 U7508 ( .A(n9844), .Z(n9928) );
  INV_X4 U7509 ( .A(n6674), .ZN(n12789) );
  INV_X2 U7510 ( .A(n12891), .ZN(n13088) );
  INV_X2 U7511 ( .A(n12891), .ZN(n13096) );
  INV_X2 U7512 ( .A(n12891), .ZN(n12984) );
  OR2_X2 U7513 ( .A1(n9901), .A2(n9809), .ZN(n9844) );
  CLKBUF_X3 U7514 ( .A(n12603), .Z(n6674) );
  NAND4_X1 U7515 ( .A1(n11043), .A2(n11042), .A3(n11041), .A4(n11040), .ZN(
        n14703) );
  AND2_X1 U7516 ( .A1(n7340), .A2(n7200), .ZN(n10686) );
  NAND4_X1 U7517 ( .A1(n10959), .A2(n10958), .A3(n10957), .A4(n10956), .ZN(
        n14704) );
  OR2_X1 U7518 ( .A1(n9888), .A2(n9962), .ZN(n9891) );
  INV_X2 U7519 ( .A(n9888), .ZN(n7282) );
  INV_X1 U7520 ( .A(n12871), .ZN(n12888) );
  CLKBUF_X1 U7521 ( .A(n6878), .Z(n6683) );
  AND2_X1 U7522 ( .A1(n6941), .A2(n9748), .ZN(n9752) );
  AOI21_X1 U7523 ( .B1(n7685), .B2(n7686), .A(n6775), .ZN(n7683) );
  INV_X1 U7525 ( .A(n9975), .ZN(n8253) );
  NAND2_X4 U7526 ( .A1(n7420), .A2(n7421), .ZN(n9975) );
  XNOR2_X1 U7527 ( .A(n8936), .B(n6990), .ZN(n7442) );
  XNOR2_X1 U7528 ( .A(n13553), .B(n13552), .ZN(n13721) );
  XNOR2_X1 U7529 ( .A(n12572), .B(n12793), .ZN(n15110) );
  AOI21_X1 U7530 ( .B1(n12856), .B2(n12855), .A(n12854), .ZN(n12857) );
  NAND2_X1 U7531 ( .A1(n14862), .A2(n6762), .ZN(n12570) );
  OR2_X1 U7532 ( .A1(n13064), .A2(n13063), .ZN(n6858) );
  NAND2_X1 U7533 ( .A1(n14875), .A2(n6755), .ZN(n14862) );
  AOI21_X1 U7534 ( .B1(n12529), .B2(n15280), .A(n12528), .ZN(n15115) );
  NAND2_X1 U7535 ( .A1(n13547), .A2(n13546), .ZN(n13545) );
  NAND2_X1 U7536 ( .A1(n7296), .A2(n7295), .ZN(n13253) );
  NOR2_X1 U7537 ( .A1(n9523), .A2(n7459), .ZN(n7458) );
  OR2_X1 U7538 ( .A1(n14904), .A2(n12547), .ZN(n14905) );
  NAND2_X1 U7539 ( .A1(n7612), .A2(n6767), .ZN(n13055) );
  AND2_X1 U7540 ( .A1(n7566), .A2(n7562), .ZN(n7561) );
  NAND2_X1 U7541 ( .A1(n7565), .A2(n7564), .ZN(n7563) );
  NAND2_X1 U7542 ( .A1(n7558), .A2(n7557), .ZN(n7566) );
  OR3_X1 U7543 ( .A1(n13041), .A2(n13044), .A3(n7614), .ZN(n7612) );
  OAI211_X1 U7544 ( .C1(n6906), .C2(n13211), .A(n6904), .B(n13214), .ZN(n13270) );
  INV_X1 U7545 ( .A(n7436), .ZN(n6671) );
  NAND2_X1 U7546 ( .A1(n9352), .A2(n9636), .ZN(n13639) );
  INV_X1 U7547 ( .A(n7148), .ZN(n14027) );
  AND2_X1 U7548 ( .A1(n9720), .A2(n9719), .ZN(n7747) );
  XNOR2_X1 U7549 ( .A(n13205), .B(n13203), .ZN(n13313) );
  NAND2_X1 U7550 ( .A1(n14224), .A2(n14223), .ZN(n14222) );
  AOI21_X1 U7551 ( .B1(n13627), .B2(n9718), .A(n7624), .ZN(n7623) );
  AND2_X1 U7552 ( .A1(n9652), .A2(n9651), .ZN(n13574) );
  AND2_X1 U7553 ( .A1(n9532), .A2(n9533), .ZN(n13592) );
  NAND2_X1 U7554 ( .A1(n15024), .A2(n12410), .ZN(n14998) );
  NAND2_X1 U7555 ( .A1(n13243), .A2(n13198), .ZN(n13307) );
  AND2_X1 U7556 ( .A1(n13938), .A2(n8676), .ZN(n13861) );
  NAND2_X1 U7557 ( .A1(n9375), .A2(n9374), .ZN(n13318) );
  NAND2_X1 U7558 ( .A1(n14673), .A2(n14674), .ZN(n14672) );
  NAND2_X1 U7559 ( .A1(n8759), .A2(n8758), .ZN(n14343) );
  XNOR2_X1 U7560 ( .A(n14426), .B(n14424), .ZN(n14673) );
  NAND2_X1 U7561 ( .A1(n7303), .A2(n7301), .ZN(n13289) );
  OAI21_X1 U7562 ( .B1(n9405), .B2(P2_DATAO_REG_24__SCAN_IN), .A(n9406), .ZN(
        n9418) );
  NAND2_X1 U7563 ( .A1(n15377), .A2(n14420), .ZN(n14426) );
  OAI21_X1 U7564 ( .B1(n13183), .B2(n6911), .A(n6908), .ZN(n13191) );
  NAND2_X1 U7565 ( .A1(n8306), .A2(n8305), .ZN(n8772) );
  AND2_X1 U7566 ( .A1(n15007), .A2(n15173), .ZN(n14986) );
  NAND2_X1 U7567 ( .A1(n12460), .A2(n12459), .ZN(n15148) );
  NAND2_X1 U7568 ( .A1(n8717), .A2(n8716), .ZN(n14285) );
  OAI21_X1 U7569 ( .B1(n11620), .B2(n8971), .A(n8972), .ZN(n11712) );
  NAND2_X1 U7570 ( .A1(n12437), .A2(n12436), .ZN(n15158) );
  NAND2_X1 U7571 ( .A1(n6929), .A2(n9355), .ZN(n9369) );
  XNOR2_X1 U7572 ( .A(n6902), .B(n6901), .ZN(n12224) );
  NOR2_X1 U7573 ( .A1(n13359), .A2(n6826), .ZN(n13383) );
  AOI21_X1 U7574 ( .B1(n6910), .B2(n7288), .A(n6909), .ZN(n6908) );
  NAND2_X1 U7575 ( .A1(n8299), .A2(n8298), .ZN(n8743) );
  NAND2_X1 U7576 ( .A1(n15426), .A2(n15424), .ZN(n15429) );
  NAND2_X1 U7577 ( .A1(n11943), .A2(n11942), .ZN(n11944) );
  NAND2_X1 U7578 ( .A1(n11400), .A2(n12804), .ZN(n11823) );
  NAND2_X1 U7579 ( .A1(n9325), .A2(n9324), .ZN(n9339) );
  NAND2_X1 U7580 ( .A1(n8586), .A2(n8585), .ZN(n12988) );
  NAND2_X1 U7581 ( .A1(n12335), .A2(n12334), .ZN(n15380) );
  NAND2_X1 U7582 ( .A1(n11713), .A2(n15363), .ZN(n11811) );
  NAND2_X1 U7583 ( .A1(n9700), .A2(n9513), .ZN(n11794) );
  XNOR2_X1 U7584 ( .A(n8284), .B(SI_18_), .ZN(n8660) );
  NAND2_X1 U7585 ( .A1(n6848), .A2(n8282), .ZN(n8284) );
  NAND2_X1 U7586 ( .A1(n10910), .A2(n8900), .ZN(n11106) );
  NAND2_X1 U7587 ( .A1(n6926), .A2(n6924), .ZN(n9307) );
  NAND2_X1 U7588 ( .A1(n12397), .A2(n12396), .ZN(n15192) );
  NAND2_X1 U7589 ( .A1(n8627), .A2(n8626), .ZN(n14376) );
  NAND2_X1 U7590 ( .A1(n11482), .A2(n11413), .ZN(n11577) );
  NAND2_X1 U7591 ( .A1(n8527), .A2(n8526), .ZN(n15349) );
  NOR2_X1 U7592 ( .A1(n11326), .A2(n7496), .ZN(n11438) );
  NAND2_X1 U7593 ( .A1(n10832), .A2(n6976), .ZN(n11008) );
  NAND2_X1 U7594 ( .A1(n6968), .A2(n6731), .ZN(n6995) );
  AND2_X1 U7595 ( .A1(n10412), .A2(n8375), .ZN(n8393) );
  NAND2_X1 U7596 ( .A1(n7682), .A2(n8271), .ZN(n8561) );
  NAND2_X1 U7597 ( .A1(n11820), .A2(n11819), .ZN(n12650) );
  NAND2_X1 U7598 ( .A1(n8473), .A2(n8472), .ZN(n12935) );
  NAND2_X1 U7599 ( .A1(n8511), .A2(n8510), .ZN(n12947) );
  INV_X2 U7600 ( .A(n15093), .ZN(n15067) );
  AND2_X1 U7601 ( .A1(n10833), .A2(n10831), .ZN(n6976) );
  AND2_X1 U7602 ( .A1(n8374), .A2(n8375), .ZN(n10414) );
  NOR2_X1 U7603 ( .A1(n10868), .A2(n6869), .ZN(n10985) );
  XNOR2_X1 U7604 ( .A(n8455), .B(n8454), .ZN(n11343) );
  NAND2_X1 U7605 ( .A1(n8252), .A2(n8251), .ZN(n8455) );
  OR2_X1 U7606 ( .A1(n10888), .A2(n11434), .ZN(n6870) );
  AND3_X1 U7607 ( .A1(n9134), .A2(n9133), .A3(n9132), .ZN(n11896) );
  AND3_X1 U7608 ( .A1(n9153), .A2(n9152), .A3(n9151), .ZN(n12173) );
  NAND2_X1 U7609 ( .A1(n9157), .A2(n6758), .ZN(n12018) );
  BUF_X1 U7610 ( .A(n12874), .Z(n13988) );
  XNOR2_X1 U7611 ( .A(n8438), .B(n8437), .ZN(n11232) );
  NAND3_X1 U7612 ( .A1(n9052), .A2(n7482), .A3(n7481), .ZN(n10674) );
  AOI21_X1 U7613 ( .B1(n7208), .B2(n7210), .A(n7205), .ZN(n7204) );
  AND3_X1 U7614 ( .A1(n9067), .A2(n9066), .A3(n9065), .ZN(n10830) );
  NAND4_X1 U7615 ( .A1(n8403), .A2(n8402), .A3(n8401), .A4(n8400), .ZN(n13985)
         );
  NAND2_X1 U7616 ( .A1(n14706), .A2(n10686), .ZN(n12602) );
  NAND4_X1 U7617 ( .A1(n8388), .A2(n8387), .A3(n8386), .A4(n8385), .ZN(n13986)
         );
  NAND2_X1 U7618 ( .A1(n7663), .A2(n8248), .ZN(n8438) );
  INV_X1 U7619 ( .A(n14702), .ZN(n11582) );
  OAI21_X1 U7620 ( .B1(n8395), .B2(n7662), .A(n7661), .ZN(n7663) );
  INV_X1 U7621 ( .A(n15092), .ZN(n14706) );
  NAND3_X1 U7622 ( .A1(n9843), .A2(n7732), .A3(n9842), .ZN(n15496) );
  INV_X2 U7623 ( .A(n9070), .ZN(n9476) );
  INV_X2 U7624 ( .A(n13358), .ZN(P3_U3897) );
  NOR2_X1 U7625 ( .A1(n10786), .A2(n10785), .ZN(n10787) );
  NAND2_X1 U7626 ( .A1(n7406), .A2(n7405), .ZN(n7404) );
  AND2_X2 U7627 ( .A1(n8216), .A2(n12564), .ZN(n8384) );
  NAND4_X1 U7628 ( .A1(n9945), .A2(n9944), .A3(n9943), .A4(n9942), .ZN(n14705)
         );
  INV_X2 U7629 ( .A(n12888), .ZN(n13097) );
  BUF_X4 U7630 ( .A(n9089), .Z(n9475) );
  AND2_X1 U7631 ( .A1(n8218), .A2(n14388), .ZN(n8336) );
  NAND2_X1 U7632 ( .A1(n9733), .A2(n8253), .ZN(n9474) );
  NAND2_X1 U7633 ( .A1(n12448), .A2(n8253), .ZN(n9889) );
  NAND2_X1 U7634 ( .A1(n9688), .A2(n9689), .ZN(n9733) );
  BUF_X1 U7635 ( .A(n8217), .Z(n12564) );
  INV_X1 U7636 ( .A(n6666), .ZN(n6681) );
  CLKBUF_X3 U7637 ( .A(n9688), .Z(n6945) );
  XNOR2_X1 U7638 ( .A(n8209), .B(n8208), .ZN(n8217) );
  AND2_X2 U7639 ( .A1(n12594), .A2(n12770), .ZN(n12592) );
  NAND2_X1 U7640 ( .A1(n8325), .A2(n13099), .ZN(n13156) );
  OAI21_X1 U7641 ( .B1(n9799), .B2(P1_IR_REG_24__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n9798) );
  XNOR2_X1 U7642 ( .A(n9827), .B(P1_IR_REG_21__SCAN_IN), .ZN(n12594) );
  XNOR2_X1 U7643 ( .A(n9830), .B(n9829), .ZN(n12770) );
  OR2_X1 U7644 ( .A1(n13830), .A2(n9682), .ZN(n9014) );
  NAND2_X1 U7645 ( .A1(n9839), .A2(n9838), .ZN(n10187) );
  XNOR2_X1 U7646 ( .A(n9150), .B(n9149), .ZN(n11331) );
  OAI21_X1 U7647 ( .B1(n8645), .B2(P2_IR_REG_18__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n7031) );
  XNOR2_X1 U7648 ( .A(n9681), .B(P3_IR_REG_26__SCAN_IN), .ZN(n9748) );
  NAND2_X1 U7649 ( .A1(n9503), .A2(n9674), .ZN(n11171) );
  OAI211_X1 U7650 ( .C1(n6896), .C2(n9679), .A(n6894), .B(n6892), .ZN(n9688)
         );
  OR2_X1 U7651 ( .A1(n9834), .A2(n9813), .ZN(n9839) );
  NOR2_X1 U7652 ( .A1(n9826), .A2(n7382), .ZN(n7381) );
  XNOR2_X1 U7653 ( .A(n9507), .B(n9506), .ZN(n10926) );
  NAND2_X1 U7654 ( .A1(n9826), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9827) );
  XNOR2_X1 U7655 ( .A(n9131), .B(P3_IR_REG_7__SCAN_IN), .ZN(n10986) );
  OAI21_X1 U7656 ( .B1(n9326), .B2(P3_IR_REG_18__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n7287) );
  OR2_X1 U7657 ( .A1(n9679), .A2(n9682), .ZN(n9681) );
  MUX2_X1 U7658 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8316), .S(
        P2_IR_REG_28__SCAN_IN), .Z(n8318) );
  XNOR2_X1 U7659 ( .A(n8228), .B(P2_IR_REG_21__SCAN_IN), .ZN(n8321) );
  XNOR2_X1 U7660 ( .A(n8226), .B(n8225), .ZN(n13099) );
  NAND2_X1 U7661 ( .A1(n7722), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6876) );
  NAND2_X1 U7662 ( .A1(n9795), .A2(n9829), .ZN(n9826) );
  XNOR2_X1 U7663 ( .A(n9685), .B(n9684), .ZN(n12124) );
  NAND2_X1 U7664 ( .A1(n9294), .A2(n9293), .ZN(n9326) );
  XNOR2_X1 U7665 ( .A(n8231), .B(n8230), .ZN(n11849) );
  NAND2_X1 U7666 ( .A1(n8227), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8228) );
  NAND2_X2 U7667 ( .A1(n9950), .A2(P1_U3086), .ZN(n15239) );
  OR2_X1 U7668 ( .A1(n8229), .A2(n14381), .ZN(n8231) );
  NAND2_X2 U7669 ( .A1(n9084), .A2(n9083), .ZN(n10801) );
  NOR2_X1 U7670 ( .A1(n8470), .A2(n7616), .ZN(n7615) );
  AND2_X1 U7671 ( .A1(n8322), .A2(n8202), .ZN(n8229) );
  NAND2_X1 U7672 ( .A1(n7383), .A2(n9810), .ZN(n7382) );
  NAND2_X1 U7673 ( .A1(n8195), .A2(n8194), .ZN(n8470) );
  INV_X1 U7674 ( .A(n8361), .ZN(n8194) );
  NAND2_X1 U7675 ( .A1(n6799), .A2(n8224), .ZN(n7616) );
  NAND2_X1 U7676 ( .A1(n7284), .A2(P1_ADDR_REG_19__SCAN_IN), .ZN(n7420) );
  INV_X1 U7677 ( .A(n7384), .ZN(n7383) );
  AND4_X1 U7678 ( .A1(n8192), .A2(n8191), .A3(n8190), .A4(n8418), .ZN(n8195)
         );
  AND3_X1 U7679 ( .A1(n9007), .A2(n9006), .A3(n9005), .ZN(n9499) );
  NAND4_X1 U7680 ( .A1(n9886), .A2(n9789), .A3(n9859), .A4(n7704), .ZN(n9986)
         );
  AND3_X1 U7681 ( .A1(n7285), .A2(n7008), .A3(n7286), .ZN(n9004) );
  NOR2_X1 U7682 ( .A1(P3_IR_REG_11__SCAN_IN), .A2(P3_IR_REG_6__SCAN_IN), .ZN(
        n7285) );
  NOR2_X1 U7683 ( .A1(P3_IR_REG_8__SCAN_IN), .A2(P3_IR_REG_9__SCAN_IN), .ZN(
        n7286) );
  INV_X1 U7684 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n9789) );
  NOR2_X1 U7685 ( .A1(P3_IR_REG_20__SCAN_IN), .A2(P3_IR_REG_23__SCAN_IN), .ZN(
        n9010) );
  NOR2_X1 U7686 ( .A1(P3_IR_REG_10__SCAN_IN), .A2(P3_IR_REG_7__SCAN_IN), .ZN(
        n7008) );
  NOR2_X1 U7687 ( .A1(P2_IR_REG_21__SCAN_IN), .A2(P2_IR_REG_20__SCAN_IN), .ZN(
        n8224) );
  INV_X1 U7688 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n8643) );
  INV_X1 U7689 ( .A(P3_ADDR_REG_2__SCAN_IN), .ZN(n8106) );
  NOR2_X1 U7690 ( .A1(P3_IR_REG_16__SCAN_IN), .A2(P3_IR_REG_15__SCAN_IN), .ZN(
        n9006) );
  NOR2_X1 U7691 ( .A1(P3_IR_REG_19__SCAN_IN), .A2(P3_IR_REG_17__SCAN_IN), .ZN(
        n9005) );
  NOR2_X1 U7692 ( .A1(P2_IR_REG_13__SCAN_IN), .A2(P2_IR_REG_15__SCAN_IN), .ZN(
        n8198) );
  INV_X1 U7693 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n8624) );
  NOR2_X1 U7694 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(P1_IR_REG_8__SCAN_IN), .ZN(
        n10241) );
  INV_X1 U7695 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n10240) );
  INV_X1 U7696 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n10244) );
  NOR2_X1 U7697 ( .A1(P2_IR_REG_7__SCAN_IN), .A2(P2_IR_REG_4__SCAN_IN), .ZN(
        n8192) );
  INV_X1 U7698 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n10239) );
  INV_X1 U7699 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n9886) );
  INV_X1 U7700 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n8418) );
  INV_X4 U7701 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  INV_X1 U7702 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n10453) );
  INV_X1 U7703 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n9846) );
  INV_X1 U7704 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n9810) );
  INV_X1 U7705 ( .A(P3_ADDR_REG_0__SCAN_IN), .ZN(n8141) );
  INV_X1 U7706 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n9794) );
  INV_X1 U7707 ( .A(P3_IR_REG_8__SCAN_IN), .ZN(n9149) );
  INV_X1 U7708 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n9829) );
  NOR2_X1 U7709 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P1_IR_REG_16__SCAN_IN), .ZN(
        n7364) );
  INV_X1 U7710 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n10456) );
  INV_X4 U7711 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3088) );
  AND3_X2 U7712 ( .A1(n7718), .A2(n9793), .A3(n9990), .ZN(n9807) );
  NAND2_X2 U7713 ( .A1(n12602), .A2(n12597), .ZN(n12794) );
  OAI222_X1 U7714 ( .A1(P1_U3086), .A2(n9821), .B1(n15238), .B2(n13093), .C1(
        n12862), .C2(n15239), .ZN(P1_U3325) );
  INV_X1 U7715 ( .A(n8886), .ZN(n8887) );
  INV_X1 U7716 ( .A(n9346), .ZN(n9388) );
  NAND4_X2 U7717 ( .A1(n9884), .A2(n9883), .A3(n9882), .A4(n9881), .ZN(n10689)
         );
  INV_X2 U7718 ( .A(n14557), .ZN(n9893) );
  AOI21_X2 U7719 ( .B1(n15287), .B2(n15288), .A(n6724), .ZN(n15059) );
  XNOR2_X2 U7720 ( .A(n8314), .B(n8313), .ZN(n8938) );
  BUF_X4 U7721 ( .A(n9880), .Z(n6677) );
  AND2_X2 U7722 ( .A1(n9820), .A2(n9819), .ZN(n9880) );
  NOR2_X2 U7724 ( .A1(n9063), .A2(n7451), .ZN(n7450) );
  INV_X2 U7725 ( .A(n10585), .ZN(n6957) );
  NAND4_X1 U7726 ( .A1(n9023), .A2(n9022), .A3(n9024), .A4(n9021), .ZN(n10585)
         );
  NAND2_X1 U7727 ( .A1(n9733), .A2(n9975), .ZN(n9435) );
  AND2_X1 U7728 ( .A1(n9018), .A2(n13842), .ZN(n6679) );
  NOR2_X2 U7729 ( .A1(n9986), .A2(P1_IR_REG_4__SCAN_IN), .ZN(n9990) );
  NAND2_X1 U7730 ( .A1(n7342), .A2(n7341), .ZN(n7340) );
  AND2_X1 U7731 ( .A1(n9821), .A2(n15234), .ZN(n9864) );
  XNOR2_X2 U7732 ( .A(n6876), .B(n9815), .ZN(n9821) );
  INV_X1 U7733 ( .A(n6683), .ZN(n6684) );
  AND2_X1 U7734 ( .A1(n9727), .A2(n9726), .ZN(n13547) );
  OR2_X1 U7735 ( .A1(n7263), .A2(n6722), .ZN(n6687) );
  INV_X1 U7736 ( .A(n7264), .ZN(n7263) );
  OAI21_X1 U7737 ( .B1(n7266), .B2(n7265), .A(n12501), .ZN(n7264) );
  AND2_X1 U7738 ( .A1(n14936), .A2(n6737), .ZN(n7255) );
  OR2_X1 U7739 ( .A1(n15158), .A2(n14969), .ZN(n12545) );
  OR2_X1 U7740 ( .A1(n15380), .A2(n14637), .ZN(n12678) );
  NAND2_X1 U7741 ( .A1(n7309), .A2(n7308), .ZN(n6903) );
  NOR2_X1 U7742 ( .A1(n11866), .A2(n11863), .ZN(n7308) );
  NOR2_X1 U7743 ( .A1(n13468), .A2(n13469), .ZN(n13502) );
  OR2_X1 U7744 ( .A1(n12658), .A2(n15385), .ZN(n15278) );
  NOR2_X1 U7745 ( .A1(n15260), .A2(n15259), .ZN(n15258) );
  OR2_X1 U7746 ( .A1(n12887), .A2(n12886), .ZN(n12896) );
  INV_X1 U7747 ( .A(n12761), .ZN(n7076) );
  INV_X1 U7748 ( .A(n7225), .ZN(n7224) );
  AND2_X1 U7749 ( .A1(n10604), .A2(n9693), .ZN(n15716) );
  INV_X1 U7750 ( .A(n10591), .ZN(n6959) );
  INV_X1 U7751 ( .A(n10772), .ZN(n7495) );
  NAND2_X1 U7752 ( .A1(n7408), .A2(n7407), .ZN(n7406) );
  INV_X1 U7753 ( .A(n10758), .ZN(n7407) );
  NOR2_X1 U7754 ( .A1(n10809), .A2(n15713), .ZN(n6869) );
  OR2_X1 U7755 ( .A1(n13540), .A2(n6675), .ZN(n9666) );
  OR2_X1 U7756 ( .A1(n13318), .A2(n13630), .ZN(n9536) );
  OR2_X1 U7757 ( .A1(n9707), .A2(n11749), .ZN(n9708) );
  OR2_X1 U7758 ( .A1(n9705), .A2(n12002), .ZN(n9709) );
  INV_X1 U7759 ( .A(n7470), .ZN(n7469) );
  OAI21_X1 U7760 ( .B1(n12023), .B2(n7471), .A(n9171), .ZN(n7470) );
  NAND2_X1 U7761 ( .A1(n15716), .A2(n9545), .ZN(n10596) );
  NAND2_X1 U7762 ( .A1(n7453), .A2(n7452), .ZN(n7451) );
  INV_X1 U7763 ( .A(P3_IR_REG_13__SCAN_IN), .ZN(n7453) );
  INV_X1 U7764 ( .A(P3_IR_REG_4__SCAN_IN), .ZN(n7452) );
  NOR2_X1 U7765 ( .A1(P3_IR_REG_5__SCAN_IN), .A2(P3_IR_REG_12__SCAN_IN), .ZN(
        n7625) );
  NAND2_X1 U7766 ( .A1(n9031), .A2(n9002), .ZN(n9063) );
  NOR2_X1 U7767 ( .A1(P3_IR_REG_3__SCAN_IN), .A2(P3_IR_REG_2__SCAN_IN), .ZN(
        n9002) );
  INV_X1 U7768 ( .A(n14388), .ZN(n8216) );
  AND2_X1 U7769 ( .A1(n12181), .A2(n8916), .ZN(n7446) );
  NAND2_X1 U7770 ( .A1(n11708), .A2(n13136), .ZN(n8913) );
  AND2_X1 U7771 ( .A1(n8894), .A2(n7531), .ZN(n13123) );
  INV_X1 U7772 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n8200) );
  NAND2_X1 U7773 ( .A1(n7283), .A2(n8233), .ZN(n7421) );
  INV_X1 U7774 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n7139) );
  NOR2_X1 U7775 ( .A1(n7719), .A2(n9803), .ZN(n7718) );
  INV_X1 U7776 ( .A(n8661), .ZN(n7677) );
  NOR2_X1 U7777 ( .A1(n10667), .A2(P1_IR_REG_17__SCAN_IN), .ZN(n11257) );
  OR2_X1 U7778 ( .A1(n7683), .A2(n8488), .ZN(n6849) );
  NAND2_X1 U7779 ( .A1(n13191), .A2(n6819), .ZN(n7303) );
  NAND2_X1 U7780 ( .A1(n6903), .A2(n6721), .ZN(n6902) );
  NAND2_X1 U7781 ( .A1(n7489), .A2(n10764), .ZN(n7488) );
  XNOR2_X1 U7782 ( .A(n10769), .B(n10768), .ZN(n10846) );
  NOR2_X1 U7783 ( .A1(n13503), .A2(n13502), .ZN(n13507) );
  NAND2_X1 U7784 ( .A1(n7635), .A2(n7634), .ZN(n13563) );
  AOI21_X1 U7785 ( .B1(n6688), .B2(n13592), .A(n6773), .ZN(n7634) );
  AOI21_X1 U7786 ( .B1(n7643), .B2(n7646), .A(n7642), .ZN(n7641) );
  NOR2_X1 U7787 ( .A1(n13772), .A2(n13693), .ZN(n7642) );
  NOR2_X1 U7788 ( .A1(n13710), .A2(n6720), .ZN(n7643) );
  OAI21_X1 U7789 ( .B1(n12197), .B2(n9601), .A(n9603), .ZN(n12267) );
  XNOR2_X1 U7790 ( .A(n12018), .B(n15759), .ZN(n12034) );
  NAND2_X1 U7791 ( .A1(n10600), .A2(n10746), .ZN(n13696) );
  OR2_X1 U7792 ( .A1(n10600), .A2(n9771), .ZN(n13694) );
  NAND2_X1 U7793 ( .A1(n9777), .A2(n9732), .ZN(n15722) );
  NAND2_X1 U7794 ( .A1(n10933), .A2(n10932), .ZN(n10936) );
  INV_X1 U7795 ( .A(n9671), .ZN(n9769) );
  NOR2_X1 U7796 ( .A1(n9781), .A2(n13827), .ZN(n10602) );
  NOR2_X1 U7797 ( .A1(n6897), .A2(P3_IR_REG_28__SCAN_IN), .ZN(n6891) );
  NAND2_X1 U7798 ( .A1(n7114), .A2(n7113), .ZN(n9445) );
  NAND2_X1 U7799 ( .A1(P2_DATAO_REG_26__SCAN_IN), .A2(n14394), .ZN(n7113) );
  INV_X1 U7800 ( .A(P3_IR_REG_17__SCAN_IN), .ZN(n9293) );
  NAND2_X1 U7801 ( .A1(n7027), .A2(n8582), .ZN(n7026) );
  INV_X1 U7802 ( .A(n11963), .ZN(n7027) );
  AOI21_X1 U7803 ( .B1(n7574), .B2(n12846), .A(n7573), .ZN(n7572) );
  AND2_X1 U7804 ( .A1(n8805), .A2(n8826), .ZN(n7573) );
  NOR2_X1 U7805 ( .A1(n7580), .A2(n7579), .ZN(n7578) );
  INV_X1 U7806 ( .A(n7733), .ZN(n7580) );
  INV_X1 U7807 ( .A(n8540), .ZN(n7579) );
  NAND2_X1 U7808 ( .A1(n8885), .A2(n8884), .ZN(n14031) );
  NAND2_X1 U7809 ( .A1(n8814), .A2(n8813), .ZN(n14247) );
  NAND2_X1 U7810 ( .A1(n7166), .A2(n6745), .ZN(n14124) );
  INV_X1 U7811 ( .A(n7162), .ZN(n7161) );
  OAI22_X1 U7812 ( .A1(n6690), .A2(n7163), .B1(n13868), .B2(n13914), .ZN(n7162) );
  OR2_X1 U7813 ( .A1(n12980), .A2(n8917), .ZN(n12211) );
  AOI21_X1 U7814 ( .B1(n7175), .B2(n7532), .A(n14057), .ZN(n7174) );
  INV_X1 U7815 ( .A(n7533), .ZN(n7175) );
  INV_X1 U7816 ( .A(n13149), .ZN(n14057) );
  NAND2_X1 U7817 ( .A1(n8320), .A2(n8319), .ZN(n14256) );
  NAND2_X1 U7818 ( .A1(n14151), .A2(n14161), .ZN(n8986) );
  NAND2_X1 U7819 ( .A1(n14222), .A2(n6690), .ZN(n14201) );
  NAND2_X1 U7820 ( .A1(n13156), .A2(n7033), .ZN(n7032) );
  OR2_X1 U7821 ( .A1(n8325), .A2(n13099), .ZN(n7033) );
  AND2_X1 U7822 ( .A1(n9787), .A2(n12058), .ZN(n8868) );
  XNOR2_X1 U7823 ( .A(n12064), .B(n14445), .ZN(n12241) );
  XNOR2_X1 U7824 ( .A(n12241), .B(n6944), .ZN(n12070) );
  NAND2_X1 U7825 ( .A1(n11768), .A2(n11767), .ZN(n12068) );
  INV_X1 U7826 ( .A(n11770), .ZN(n11768) );
  NAND2_X1 U7827 ( .A1(n6687), .A2(n14859), .ZN(n7261) );
  AOI21_X1 U7828 ( .B1(n6687), .B2(n7260), .A(n7259), .ZN(n7258) );
  NOR2_X1 U7829 ( .A1(n15121), .A2(n14688), .ZN(n7259) );
  AOI21_X1 U7830 ( .B1(n7255), .B2(n7254), .A(n6770), .ZN(n7253) );
  INV_X1 U7831 ( .A(n14963), .ZN(n7254) );
  INV_X1 U7832 ( .A(n7255), .ZN(n7252) );
  NAND2_X1 U7833 ( .A1(n15163), .A2(n7353), .ZN(n14960) );
  NOR2_X1 U7834 ( .A1(n14963), .A2(n7354), .ZN(n7353) );
  INV_X1 U7835 ( .A(n12544), .ZN(n7354) );
  NAND2_X1 U7836 ( .A1(n7245), .A2(n7244), .ZN(n7243) );
  INV_X1 U7837 ( .A(n7249), .ZN(n7244) );
  INV_X1 U7838 ( .A(n15184), .ZN(n15032) );
  OR2_X1 U7839 ( .A1(n15196), .A2(n15372), .ZN(n12681) );
  NAND2_X1 U7840 ( .A1(n12355), .A2(n12810), .ZN(n6874) );
  AND2_X2 U7841 ( .A1(n9807), .A2(n9806), .ZN(n9814) );
  INV_X1 U7842 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n9806) );
  NAND2_X1 U7843 ( .A1(n15788), .A2(n7821), .ZN(n7825) );
  OAI21_X1 U7844 ( .B1(P1_ADDR_REG_8__SCAN_IN), .B2(n8104), .A(n7765), .ZN(
        n7800) );
  OAI21_X1 U7845 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(n7771), .A(n7770), .ZN(
        n7794) );
  OR2_X1 U7846 ( .A1(n9474), .A2(n9029), .ZN(n6983) );
  OR2_X1 U7847 ( .A1(n9435), .A2(n9955), .ZN(n6982) );
  XNOR2_X1 U7848 ( .A(n13485), .B(n13501), .ZN(n13464) );
  AND2_X1 U7849 ( .A1(n10860), .A2(n9689), .ZN(n13529) );
  NAND2_X1 U7850 ( .A1(n7035), .A2(n7034), .ZN(n12855) );
  INV_X1 U7851 ( .A(n12846), .ZN(n7034) );
  INV_X1 U7852 ( .A(n12847), .ZN(n7035) );
  INV_X1 U7853 ( .A(n13099), .ZN(n13169) );
  NAND2_X1 U7854 ( .A1(n14875), .A2(n12549), .ZN(n14860) );
  NOR2_X1 U7855 ( .A1(n15258), .A2(n7833), .ZN(n15262) );
  INV_X1 U7856 ( .A(n6802), .ZN(n7588) );
  NAND2_X1 U7857 ( .A1(n12630), .A2(n12632), .ZN(n7711) );
  AND2_X1 U7858 ( .A1(n6801), .A2(n7059), .ZN(n7058) );
  NAND2_X1 U7859 ( .A1(n12634), .A2(n7060), .ZN(n7059) );
  INV_X1 U7860 ( .A(n12634), .ZN(n7061) );
  INV_X1 U7861 ( .A(n12937), .ZN(n7552) );
  NAND2_X1 U7862 ( .A1(n12932), .A2(n6743), .ZN(n7550) );
  NOR2_X1 U7863 ( .A1(n6766), .A2(n7084), .ZN(n7083) );
  AND2_X1 U7864 ( .A1(n12651), .A2(n7085), .ZN(n7084) );
  INV_X1 U7865 ( .A(n12655), .ZN(n7708) );
  NAND2_X1 U7866 ( .A1(n12950), .A2(n6748), .ZN(n7599) );
  OAI21_X1 U7867 ( .B1(n12943), .B2(n12942), .A(n6754), .ZN(n7600) );
  OAI21_X1 U7868 ( .B1(n12684), .B2(n7092), .A(n12683), .ZN(n7091) );
  INV_X1 U7869 ( .A(n12671), .ZN(n7092) );
  INV_X1 U7870 ( .A(n12702), .ZN(n12703) );
  OAI21_X1 U7871 ( .B1(n12720), .B2(n12719), .A(n12718), .ZN(n12722) );
  NAND2_X1 U7872 ( .A1(n12723), .A2(n12725), .ZN(n7724) );
  INV_X1 U7873 ( .A(n12726), .ZN(n7070) );
  AND2_X1 U7874 ( .A1(n7705), .A2(n7068), .ZN(n7067) );
  NAND2_X1 U7875 ( .A1(n7069), .A2(n12726), .ZN(n7068) );
  MUX2_X1 U7876 ( .A(n14690), .B(n15133), .S(n12789), .Z(n12741) );
  INV_X1 U7877 ( .A(n12748), .ZN(n7080) );
  MUX2_X1 U7878 ( .A(n14689), .B(n14516), .S(n12789), .Z(n12748) );
  NOR2_X1 U7879 ( .A1(n8713), .A2(SI_21_), .ZN(n8292) );
  INV_X1 U7880 ( .A(n8638), .ZN(n8281) );
  INV_X1 U7881 ( .A(n8279), .ZN(n6847) );
  INV_X1 U7882 ( .A(n9393), .ZN(n7111) );
  OR2_X1 U7883 ( .A1(n13057), .A2(n13056), .ZN(n13062) );
  NAND2_X1 U7884 ( .A1(n6860), .A2(n7593), .ZN(n7592) );
  NAND2_X1 U7885 ( .A1(n6694), .A2(n6772), .ZN(n7593) );
  MUX2_X1 U7886 ( .A(n15113), .B(n14687), .S(n6674), .Z(n12757) );
  AOI21_X1 U7887 ( .B1(n12756), .B2(n12755), .A(n7075), .ZN(n7073) );
  NOR2_X1 U7888 ( .A1(n7076), .A2(n12760), .ZN(n7075) );
  XNOR2_X1 U7889 ( .A(n12593), .B(n15244), .ZN(n12767) );
  INV_X1 U7890 ( .A(n12491), .ZN(n7265) );
  INV_X1 U7891 ( .A(n12592), .ZN(n9850) );
  AOI21_X1 U7892 ( .B1(n8771), .B2(n7675), .A(n7674), .ZN(n7673) );
  AOI21_X1 U7893 ( .B1(n8771), .B2(n8310), .A(SI_26_), .ZN(n7676) );
  NAND2_X1 U7894 ( .A1(n8743), .A2(n8300), .ZN(n8303) );
  NAND2_X1 U7895 ( .A1(n8677), .A2(n8289), .ZN(n7214) );
  NOR2_X1 U7896 ( .A1(n6813), .A2(n7217), .ZN(n7216) );
  INV_X1 U7897 ( .A(n8289), .ZN(n7217) );
  NAND2_X1 U7898 ( .A1(n8286), .A2(n10544), .ZN(n8289) );
  INV_X1 U7899 ( .A(n9957), .ZN(n7483) );
  AND2_X1 U7900 ( .A1(n15309), .A2(n15303), .ZN(n9668) );
  INV_X1 U7901 ( .A(n9508), .ZN(n9669) );
  AND2_X1 U7902 ( .A1(n9665), .A2(n9666), .ZN(n7119) );
  NAND2_X1 U7903 ( .A1(n11177), .A2(n10754), .ZN(n10755) );
  NAND2_X1 U7904 ( .A1(n10801), .A2(P3_REG2_REG_4__SCAN_IN), .ZN(n7405) );
  NAND2_X1 U7905 ( .A1(n7413), .A2(n7412), .ZN(n6954) );
  NAND2_X1 U7906 ( .A1(n11331), .A2(P3_REG2_REG_8__SCAN_IN), .ZN(n7412) );
  NAND2_X1 U7907 ( .A1(n13377), .A2(P3_REG1_REG_12__SCAN_IN), .ZN(n6981) );
  NOR2_X1 U7908 ( .A1(n13523), .A2(n13525), .ZN(n7526) );
  AOI21_X1 U7909 ( .B1(n13506), .B2(n7526), .A(n6838), .ZN(n7525) );
  INV_X1 U7910 ( .A(n7461), .ZN(n7459) );
  OR2_X1 U7911 ( .A1(n13267), .A2(n13638), .ZN(n9538) );
  OR2_X1 U7912 ( .A1(n13813), .A2(n13664), .ZN(n9716) );
  INV_X1 U7913 ( .A(n7653), .ZN(n7652) );
  NAND2_X1 U7914 ( .A1(n13650), .A2(n7654), .ZN(n7653) );
  INV_X1 U7915 ( .A(n7655), .ZN(n7654) );
  OR2_X1 U7916 ( .A1(n7641), .A2(n7639), .ZN(n7638) );
  AND2_X1 U7917 ( .A1(n9711), .A2(n7627), .ZN(n7626) );
  INV_X1 U7918 ( .A(n9154), .ZN(n7471) );
  INV_X1 U7919 ( .A(n11285), .ZN(n9768) );
  AND2_X1 U7920 ( .A1(n9013), .A2(n9026), .ZN(n7659) );
  NOR2_X1 U7921 ( .A1(n7322), .A2(n7107), .ZN(n7105) );
  INV_X1 U7922 ( .A(n9257), .ZN(n7323) );
  NOR2_X1 U7923 ( .A1(n9128), .A2(n7325), .ZN(n7324) );
  INV_X1 U7924 ( .A(n9116), .ZN(n7325) );
  NAND2_X1 U7925 ( .A1(n7317), .A2(n9057), .ZN(n7315) );
  INV_X1 U7926 ( .A(n9046), .ZN(n7317) );
  INV_X1 U7927 ( .A(n8467), .ZN(n7015) );
  INV_X1 U7928 ( .A(n13853), .ZN(n7564) );
  AND2_X1 U7929 ( .A1(n13918), .A2(n8731), .ZN(n7052) );
  NAND2_X1 U7930 ( .A1(n7051), .A2(n8731), .ZN(n7050) );
  INV_X1 U7931 ( .A(n7598), .ZN(n7051) );
  INV_X1 U7932 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n8562) );
  NAND2_X1 U7933 ( .A1(n14104), .A2(n14116), .ZN(n7429) );
  OR2_X1 U7934 ( .A1(n14274), .A2(n13048), .ZN(n14116) );
  NOR2_X1 U7935 ( .A1(n13135), .A2(n7426), .ZN(n7425) );
  INV_X1 U7936 ( .A(n8909), .ZN(n7426) );
  NAND2_X1 U7937 ( .A1(n10384), .A2(n12882), .ZN(n8894) );
  INV_X1 U7938 ( .A(n8983), .ZN(n7538) );
  INV_X1 U7939 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n8830) );
  OR2_X2 U7940 ( .A1(n14553), .A2(n15291), .ZN(n14555) );
  NAND2_X1 U7941 ( .A1(n13083), .A2(n11026), .ZN(n7689) );
  NOR2_X1 U7942 ( .A1(n7265), .A2(n6722), .ZN(n7262) );
  AND2_X1 U7943 ( .A1(n12818), .A2(n12548), .ZN(n7367) );
  NOR2_X1 U7944 ( .A1(n15154), .A2(n7195), .ZN(n7194) );
  INV_X1 U7945 ( .A(n7196), .ZN(n7195) );
  NOR2_X1 U7946 ( .A1(n12710), .A2(n7360), .ZN(n7359) );
  INV_X1 U7947 ( .A(n12540), .ZN(n7360) );
  INV_X1 U7948 ( .A(n12709), .ZN(n7356) );
  NOR2_X1 U7949 ( .A1(n15196), .A2(n7190), .ZN(n7189) );
  INV_X1 U7950 ( .A(n7191), .ZN(n7190) );
  NAND2_X1 U7951 ( .A1(n11581), .A2(n11414), .ZN(n7344) );
  INV_X1 U7952 ( .A(n7701), .ZN(n7700) );
  AOI21_X1 U7953 ( .B1(n7701), .B2(n7699), .A(n7698), .ZN(n7697) );
  INV_X1 U7954 ( .A(n12778), .ZN(n7698) );
  INV_X1 U7955 ( .A(n12556), .ZN(n7699) );
  OAI21_X1 U7956 ( .B1(n8883), .B2(n8882), .A(n8881), .ZN(n12557) );
  INV_X1 U7957 ( .A(n7668), .ZN(n7667) );
  INV_X1 U7958 ( .A(n9835), .ZN(n9837) );
  AND2_X1 U7959 ( .A1(n7671), .A2(n7669), .ZN(n7668) );
  NAND2_X1 U7960 ( .A1(n7676), .A2(n7672), .ZN(n7671) );
  NAND2_X1 U7961 ( .A1(n7673), .A2(n7670), .ZN(n7669) );
  INV_X1 U7962 ( .A(n8310), .ZN(n7672) );
  OAI21_X1 U7963 ( .B1(n8678), .B2(n8677), .A(n8289), .ZN(n8710) );
  MUX2_X1 U7964 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(P1_DATAO_REG_20__SCAN_IN), 
        .S(n9950), .Z(n8708) );
  AOI21_X1 U7965 ( .B1(n7222), .B2(n7224), .A(n7220), .ZN(n7219) );
  INV_X1 U7966 ( .A(n8277), .ZN(n7220) );
  OR2_X1 U7967 ( .A1(n10358), .A2(P1_IR_REG_11__SCAN_IN), .ZN(n10359) );
  NAND2_X1 U7968 ( .A1(n6862), .A2(n8243), .ZN(n8395) );
  NAND2_X1 U7969 ( .A1(n6863), .A2(n8241), .ZN(n6861) );
  AND2_X1 U7970 ( .A1(n8237), .A2(SI_1_), .ZN(n8238) );
  XNOR2_X1 U7971 ( .A(P3_ADDR_REG_1__SCAN_IN), .B(P1_ADDR_REG_1__SCAN_IN), 
        .ZN(n7808) );
  OAI21_X1 U7972 ( .B1(P1_ADDR_REG_2__SCAN_IN), .B2(n8106), .A(n7751), .ZN(
        n7752) );
  XNOR2_X1 U7973 ( .A(n7755), .B(n7138), .ZN(n7803) );
  XNOR2_X1 U7974 ( .A(n7757), .B(n7136), .ZN(n7817) );
  INV_X1 U7975 ( .A(P3_ADDR_REG_5__SCAN_IN), .ZN(n7136) );
  INV_X1 U7976 ( .A(P3_ADDR_REG_9__SCAN_IN), .ZN(n8083) );
  INV_X1 U7977 ( .A(n13216), .ZN(n7300) );
  AND2_X1 U7978 ( .A1(n13332), .A2(n7299), .ZN(n7298) );
  OR2_X1 U7979 ( .A1(n13271), .A2(n7300), .ZN(n7299) );
  XNOR2_X1 U7980 ( .A(n13250), .B(n13565), .ZN(n13252) );
  OR2_X1 U7981 ( .A1(n9346), .A2(n9123), .ZN(n9124) );
  NOR2_X1 U7982 ( .A1(n9121), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n9136) );
  NAND2_X1 U7983 ( .A1(n6915), .A2(n11297), .ZN(n6918) );
  AND2_X1 U7984 ( .A1(n9136), .A2(n10983), .ZN(n9155) );
  AOI21_X1 U7985 ( .B1(n12224), .B2(n12223), .A(n6900), .ZN(n12382) );
  OAI21_X1 U7986 ( .B1(n13307), .B2(n7305), .A(n6898), .ZN(n13205) );
  AOI21_X1 U7987 ( .B1(n7304), .B2(n6899), .A(n6744), .ZN(n6898) );
  INV_X1 U7988 ( .A(n13306), .ZN(n6899) );
  OR2_X1 U7989 ( .A1(n9376), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n9386) );
  NAND2_X1 U7990 ( .A1(n6882), .A2(n6884), .ZN(n6881) );
  NAND2_X1 U7991 ( .A1(n6883), .A2(n10596), .ZN(n6882) );
  AND2_X1 U7992 ( .A1(n13225), .A2(n7291), .ZN(n7290) );
  NAND2_X1 U7993 ( .A1(n7292), .A2(n13185), .ZN(n7291) );
  INV_X1 U7994 ( .A(n13182), .ZN(n7292) );
  NAND2_X1 U7995 ( .A1(n9089), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n9035) );
  NAND2_X1 U7996 ( .A1(n7488), .A2(n7487), .ZN(n10818) );
  XNOR2_X1 U7997 ( .A(n10755), .B(n10768), .ZN(n10848) );
  NAND2_X1 U7998 ( .A1(n7494), .A2(n7492), .ZN(n10786) );
  NAND2_X1 U7999 ( .A1(n7495), .A2(n7493), .ZN(n7492) );
  INV_X1 U8000 ( .A(n10770), .ZN(n7493) );
  NAND2_X1 U8001 ( .A1(n6872), .A2(P3_REG2_REG_7__SCAN_IN), .ZN(n6968) );
  INV_X1 U8002 ( .A(n7511), .ZN(n7503) );
  OAI21_X1 U8003 ( .B1(n10790), .B2(n7508), .A(n7505), .ZN(n7504) );
  OR2_X1 U8004 ( .A1(n10789), .A2(n10986), .ZN(n7508) );
  INV_X1 U8005 ( .A(n7506), .ZN(n7505) );
  OAI21_X1 U8006 ( .B1(n7511), .B2(n7507), .A(n7509), .ZN(n7506) );
  NAND2_X1 U8007 ( .A1(n6995), .A2(n6994), .ZN(n7413) );
  INV_X1 U8008 ( .A(n10989), .ZN(n6994) );
  XNOR2_X1 U8009 ( .A(n6954), .B(n11332), .ZN(n11333) );
  AND2_X1 U8010 ( .A1(n11331), .A2(P3_REG1_REG_8__SCAN_IN), .ZN(n7496) );
  NOR2_X1 U8011 ( .A1(n11327), .A2(n15780), .ZN(n11439) );
  NOR2_X1 U8012 ( .A1(n11450), .A2(n11449), .ZN(n11900) );
  NOR2_X1 U8013 ( .A1(n11900), .A2(n7414), .ZN(n11971) );
  AND2_X1 U8014 ( .A1(n11914), .A2(P3_REG2_REG_10__SCAN_IN), .ZN(n7414) );
  OR2_X1 U8015 ( .A1(n13378), .A2(n9234), .ZN(n7491) );
  NOR2_X1 U8016 ( .A1(n13450), .A2(n13451), .ZN(n13454) );
  INV_X1 U8017 ( .A(n6953), .ZN(n13448) );
  XNOR2_X1 U8018 ( .A(n13434), .B(n13449), .ZN(n13428) );
  AOI21_X1 U8019 ( .B1(n13440), .B2(n13449), .A(n13439), .ZN(n13478) );
  NAND2_X1 U8020 ( .A1(n7636), .A2(n6688), .ZN(n13575) );
  INV_X1 U8021 ( .A(n13603), .ZN(n13580) );
  OR2_X1 U8022 ( .A1(n13588), .A2(n13592), .ZN(n7636) );
  OR2_X1 U8023 ( .A1(n13626), .A2(n13627), .ZN(n13624) );
  INV_X1 U8024 ( .A(n7476), .ZN(n7475) );
  OAI21_X1 U8025 ( .B1(n13662), .B2(n7477), .A(n9634), .ZN(n7476) );
  OR2_X1 U8026 ( .A1(n13670), .A2(n13681), .ZN(n9623) );
  NOR2_X1 U8027 ( .A1(n7656), .A2(n13670), .ZN(n7655) );
  OR2_X1 U8028 ( .A1(n13660), .A2(n7653), .ZN(n13649) );
  NOR2_X1 U8029 ( .A1(n13661), .A2(n13662), .ZN(n13660) );
  AND4_X1 U8030 ( .A1(n9285), .A2(n9284), .A3(n9283), .A4(n9282), .ZN(n13680)
         );
  INV_X1 U8031 ( .A(n13326), .ZN(n13695) );
  NAND2_X1 U8032 ( .A1(n7646), .A2(n7645), .ZN(n7644) );
  INV_X1 U8033 ( .A(n9606), .ZN(n7484) );
  NAND2_X1 U8034 ( .A1(n7647), .A2(n6695), .ZN(n7646) );
  NAND2_X1 U8035 ( .A1(n12088), .A2(n9712), .ZN(n12193) );
  OR2_X1 U8036 ( .A1(n9192), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n9209) );
  NAND2_X1 U8037 ( .A1(n12043), .A2(n9588), .ZN(n12087) );
  NAND2_X1 U8038 ( .A1(n11997), .A2(n7472), .ZN(n12043) );
  NOR2_X1 U8039 ( .A1(n7627), .A2(n7473), .ZN(n7472) );
  AND4_X1 U8040 ( .A1(n9178), .A2(n9177), .A3(n9176), .A4(n9175), .ZN(n12050)
         );
  NAND2_X1 U8041 ( .A1(n7632), .A2(n7631), .ZN(n7630) );
  NAND2_X1 U8042 ( .A1(n11794), .A2(n9711), .ZN(n7631) );
  NAND2_X1 U8043 ( .A1(n7630), .A2(n7627), .ZN(n12091) );
  XNOR2_X1 U8044 ( .A(n13357), .B(n12173), .ZN(n12016) );
  INV_X1 U8045 ( .A(n12016), .ZN(n12023) );
  NAND2_X1 U8046 ( .A1(n12024), .A2(n12023), .ZN(n12022) );
  OR2_X1 U8047 ( .A1(n10748), .A2(n10768), .ZN(n9065) );
  AND2_X1 U8048 ( .A1(n13826), .A2(n10500), .ZN(n10934) );
  AND2_X1 U8049 ( .A1(n9472), .A2(n9471), .ZN(n9486) );
  NOR2_X1 U8050 ( .A1(n7333), .A2(n9469), .ZN(n7331) );
  NAND2_X1 U8051 ( .A1(n9445), .A2(n7336), .ZN(n7332) );
  AOI21_X1 U8052 ( .B1(n6893), .B2(P3_IR_REG_26__SCAN_IN), .A(n6779), .ZN(
        n6892) );
  NAND2_X1 U8053 ( .A1(n9679), .A2(n6895), .ZN(n6894) );
  INV_X1 U8054 ( .A(n6896), .ZN(n6893) );
  AND2_X1 U8055 ( .A1(n12390), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n7116) );
  NAND2_X1 U8056 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(P3_IR_REG_25__SCAN_IN), 
        .ZN(n6949) );
  INV_X1 U8057 ( .A(P3_IR_REG_21__SCAN_IN), .ZN(n9009) );
  INV_X1 U8058 ( .A(P3_IR_REG_24__SCAN_IN), .ZN(n9684) );
  XNOR2_X1 U8059 ( .A(n9404), .B(P1_DATAO_REG_24__SCAN_IN), .ZN(n9405) );
  NAND2_X1 U8060 ( .A1(n6830), .A2(n6713), .ZN(n7327) );
  INV_X1 U8061 ( .A(n9371), .ZN(n7328) );
  NAND2_X1 U8062 ( .A1(P1_DATAO_REG_21__SCAN_IN), .A2(n9370), .ZN(n9371) );
  OR2_X1 U8063 ( .A1(n9502), .A2(P3_IR_REG_21__SCAN_IN), .ZN(n9674) );
  NAND2_X1 U8064 ( .A1(n9354), .A2(n12426), .ZN(n6929) );
  XNOR2_X1 U8065 ( .A(n9353), .B(n11848), .ZN(n9354) );
  NAND2_X1 U8066 ( .A1(P1_DATAO_REG_16__SCAN_IN), .A2(n6925), .ZN(n6924) );
  NAND2_X1 U8067 ( .A1(n9288), .A2(n9287), .ZN(n6926) );
  NAND2_X1 U8068 ( .A1(n7106), .A2(n9244), .ZN(n9256) );
  NAND2_X1 U8069 ( .A1(n9242), .A2(P1_DATAO_REG_13__SCAN_IN), .ZN(n7106) );
  INV_X1 U8070 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n9181) );
  OR2_X1 U8071 ( .A1(n9148), .A2(P3_IR_REG_7__SCAN_IN), .ZN(n9164) );
  NAND2_X1 U8072 ( .A1(n9100), .A2(n9099), .ZN(n9115) );
  CLKBUF_X1 U8073 ( .A(n9063), .Z(n9081) );
  OR2_X1 U8074 ( .A1(n10566), .A2(n7020), .ZN(n7019) );
  INV_X1 U8075 ( .A(n7026), .ZN(n7025) );
  AND2_X1 U8076 ( .A1(n12129), .A2(n7024), .ZN(n7023) );
  NAND2_X1 U8077 ( .A1(n7026), .A2(n7029), .ZN(n7024) );
  INV_X1 U8078 ( .A(n8453), .ZN(n7017) );
  OR2_X1 U8079 ( .A1(n8520), .A2(n8519), .ZN(n8521) );
  NAND2_X1 U8080 ( .A1(n11264), .A2(n6752), .ZN(n7039) );
  INV_X1 U8081 ( .A(n8505), .ZN(n7040) );
  AND2_X1 U8082 ( .A1(n8620), .A2(n7582), .ZN(n7581) );
  INV_X1 U8083 ( .A(n13888), .ZN(n7582) );
  AND2_X1 U8084 ( .A1(n8675), .A2(n8659), .ZN(n7601) );
  NAND2_X1 U8085 ( .A1(n7042), .A2(n13896), .ZN(n13898) );
  NAND2_X1 U8086 ( .A1(n13887), .A2(n13895), .ZN(n7042) );
  NAND4_X1 U8087 ( .A1(n8340), .A2(n8339), .A3(n8338), .A4(n8337), .ZN(n12874)
         );
  AND2_X1 U8088 ( .A1(n7150), .A2(n7148), .ZN(n14037) );
  OAI21_X1 U8089 ( .B1(n14062), .B2(n7146), .A(n7145), .ZN(n7150) );
  NOR2_X1 U8090 ( .A1(n14062), .A2(n14247), .ZN(n14048) );
  NAND2_X1 U8091 ( .A1(n14058), .A2(n14057), .ZN(n14056) );
  AND2_X1 U8092 ( .A1(n14343), .A2(n13965), .ZN(n7537) );
  NAND2_X1 U8093 ( .A1(n14089), .A2(n7183), .ZN(n7182) );
  INV_X1 U8094 ( .A(n7537), .ZN(n7183) );
  INV_X1 U8095 ( .A(n7429), .ZN(n7430) );
  AND2_X1 U8096 ( .A1(n14118), .A2(n14116), .ZN(n14100) );
  NAND2_X1 U8097 ( .A1(n14120), .A2(n8987), .ZN(n14118) );
  AND2_X1 U8098 ( .A1(n8926), .A2(n8925), .ZN(n14170) );
  INV_X1 U8099 ( .A(n14222), .ZN(n7160) );
  AND2_X1 U8100 ( .A1(n12211), .A2(n8918), .ZN(n12181) );
  NAND2_X1 U8101 ( .A1(n6967), .A2(n6966), .ZN(n12102) );
  INV_X1 U8102 ( .A(n11712), .ZN(n8974) );
  NAND2_X1 U8103 ( .A1(n11106), .A2(n13128), .ZN(n11105) );
  NAND2_X1 U8104 ( .A1(n13124), .A2(n11156), .ZN(n7155) );
  NAND2_X1 U8105 ( .A1(n13086), .A2(n13085), .ZN(n14020) );
  NAND2_X1 U8106 ( .A1(n6866), .A2(n13094), .ZN(n14019) );
  OR2_X1 U8107 ( .A1(n13093), .A2(n8358), .ZN(n6866) );
  NOR2_X1 U8108 ( .A1(n14246), .A2(n6993), .ZN(n6992) );
  AND2_X1 U8109 ( .A1(n14247), .A2(n15672), .ZN(n6993) );
  NAND2_X1 U8110 ( .A1(n8792), .A2(n8791), .ZN(n14329) );
  AND2_X1 U8111 ( .A1(n13118), .A2(n13117), .ZN(n14080) );
  NAND2_X1 U8112 ( .A1(n14124), .A2(n8988), .ZN(n14105) );
  XNOR2_X1 U8113 ( .A(n14343), .B(n13965), .ZN(n14104) );
  NOR2_X1 U8114 ( .A1(n14105), .A2(n14104), .ZN(n14107) );
  NOR2_X1 U8115 ( .A1(n6986), .A2(n7165), .ZN(n7164) );
  INV_X1 U8116 ( .A(n8985), .ZN(n7165) );
  NAND2_X1 U8117 ( .A1(n12435), .A2(n8412), .ZN(n8717) );
  AOI21_X1 U8118 ( .B1(n6685), .B2(n7163), .A(n6769), .ZN(n7157) );
  OAI21_X1 U8119 ( .B1(n12101), .B2(n6777), .A(n7541), .ZN(n12204) );
  NAND2_X1 U8120 ( .A1(n7543), .A2(n8980), .ZN(n7541) );
  INV_X1 U8121 ( .A(n12181), .ZN(n13142) );
  NAND2_X1 U8122 ( .A1(n8978), .A2(n13141), .ZN(n12099) );
  INV_X1 U8123 ( .A(n12101), .ZN(n8978) );
  AND2_X1 U8124 ( .A1(n8840), .A2(n8839), .ZN(n15628) );
  NAND2_X1 U8125 ( .A1(n8229), .A2(n7184), .ZN(n8317) );
  AND2_X1 U8126 ( .A1(n8206), .A2(n7185), .ZN(n7184) );
  INV_X1 U8127 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n7185) );
  NOR2_X1 U8128 ( .A1(P2_IR_REG_29__SCAN_IN), .A2(P2_IR_REG_31__SCAN_IN), .ZN(
        n8212) );
  INV_X1 U8129 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n8833) );
  AND2_X1 U8130 ( .A1(n8855), .A2(n8857), .ZN(n8831) );
  NAND2_X1 U8131 ( .A1(n8831), .A2(n8830), .ZN(n8836) );
  XNOR2_X1 U8132 ( .A(n8858), .B(n8857), .ZN(n12058) );
  NOR2_X1 U8133 ( .A1(n8470), .A2(P2_IR_REG_8__SCAN_IN), .ZN(n8490) );
  NAND2_X1 U8134 ( .A1(n12417), .A2(n12416), .ZN(n14448) );
  NAND2_X1 U8135 ( .A1(n6879), .A2(n9820), .ZN(n9855) );
  AND2_X1 U8136 ( .A1(n15234), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n6879) );
  AOI21_X1 U8137 ( .B1(n7379), .B2(n14570), .A(n7378), .ZN(n7377) );
  INV_X1 U8138 ( .A(n14645), .ZN(n7378) );
  NOR2_X1 U8139 ( .A1(n9862), .A2(n9861), .ZN(n9878) );
  NOR2_X1 U8140 ( .A1(n14656), .A2(n7387), .ZN(n7386) );
  INV_X1 U8141 ( .A(n14440), .ZN(n7387) );
  OR2_X1 U8142 ( .A1(n7696), .A2(n12832), .ZN(n7695) );
  AND2_X1 U8143 ( .A1(n12834), .A2(n12833), .ZN(n7696) );
  AND4_X1 U8144 ( .A1(n12823), .A2(n7729), .A3(n12822), .A4(n7744), .ZN(n12824) );
  OAI21_X1 U8145 ( .B1(n12777), .B2(n12776), .A(n12775), .ZN(n12792) );
  OAI21_X1 U8146 ( .B1(n12774), .B2(n12773), .A(n12772), .ZN(n12775) );
  NAND2_X1 U8147 ( .A1(n7689), .A2(n7687), .ZN(n7690) );
  NOR2_X1 U8148 ( .A1(n12789), .A2(n7688), .ZN(n7687) );
  INV_X1 U8149 ( .A(n12782), .ZN(n7688) );
  INV_X1 U8150 ( .A(n12770), .ZN(n12787) );
  AND4_X1 U8151 ( .A1(n12343), .A2(n12342), .A3(n12341), .A4(n12340), .ZN(
        n14637) );
  NAND2_X1 U8152 ( .A1(n7689), .A2(n12782), .ZN(n14844) );
  NAND2_X1 U8153 ( .A1(n14899), .A2(n7199), .ZN(n14867) );
  NAND2_X1 U8154 ( .A1(n12503), .A2(n12502), .ZN(n14866) );
  INV_X1 U8155 ( .A(n12819), .ZN(n14876) );
  NAND2_X1 U8156 ( .A1(n7267), .A2(n7266), .ZN(n14889) );
  NAND2_X1 U8157 ( .A1(n14905), .A2(n12548), .ZN(n14897) );
  NAND2_X1 U8158 ( .A1(n7251), .A2(n7250), .ZN(n14925) );
  AOI21_X1 U8159 ( .B1(n7252), .B2(n7253), .A(n14921), .ZN(n7251) );
  INV_X1 U8160 ( .A(n14692), .ZN(n14942) );
  AND2_X1 U8161 ( .A1(n15027), .A2(n15014), .ZN(n15007) );
  AND2_X1 U8162 ( .A1(n14985), .A2(n6735), .ZN(n7278) );
  NOR2_X1 U8163 ( .A1(n12539), .A2(n7363), .ZN(n7362) );
  INV_X1 U8164 ( .A(n12536), .ZN(n7363) );
  INV_X1 U8165 ( .A(n12814), .ZN(n14999) );
  NOR2_X1 U8166 ( .A1(n7248), .A2(n15019), .ZN(n7242) );
  NAND2_X1 U8167 ( .A1(n15278), .A2(n7269), .ZN(n7268) );
  AOI21_X1 U8168 ( .B1(n6696), .B2(n15278), .A(n15288), .ZN(n7270) );
  INV_X1 U8169 ( .A(n12285), .ZN(n7269) );
  INV_X1 U8170 ( .A(n15271), .ZN(n12658) );
  AOI21_X1 U8171 ( .B1(n6729), .B2(n7352), .A(n7349), .ZN(n7348) );
  INV_X1 U8172 ( .A(n12274), .ZN(n7349) );
  NAND2_X1 U8173 ( .A1(n11944), .A2(n12809), .ZN(n12161) );
  NAND2_X1 U8174 ( .A1(n11834), .A2(n11833), .ZN(n11836) );
  NAND2_X1 U8175 ( .A1(n11577), .A2(n12803), .ZN(n11576) );
  AND2_X1 U8176 ( .A1(n12401), .A2(n12400), .ZN(n15184) );
  INV_X1 U8177 ( .A(n15398), .ZN(n15409) );
  INV_X1 U8178 ( .A(n15495), .ZN(n15518) );
  INV_X1 U8179 ( .A(n15280), .ZN(n15481) );
  AND2_X1 U8180 ( .A1(n7702), .A2(n12560), .ZN(n7701) );
  INV_X1 U8181 ( .A(n12562), .ZN(n7702) );
  NAND2_X1 U8182 ( .A1(n9814), .A2(n9813), .ZN(n9835) );
  INV_X1 U8183 ( .A(n7719), .ZN(n7402) );
  NOR2_X1 U8184 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), .ZN(
        n9847) );
  NAND2_X1 U8185 ( .A1(n7207), .A2(n8263), .ZN(n8522) );
  NAND2_X1 U8186 ( .A1(n8506), .A2(n8261), .ZN(n7207) );
  XNOR2_X1 U8187 ( .A(n8489), .B(n8488), .ZN(n11818) );
  XNOR2_X1 U8188 ( .A(n8242), .B(n9960), .ZN(n7203) );
  XNOR2_X1 U8189 ( .A(n7817), .B(P1_ADDR_REG_5__SCAN_IN), .ZN(n7818) );
  AND2_X1 U8190 ( .A1(n7230), .A2(n6787), .ZN(n7829) );
  NOR2_X1 U8191 ( .A1(n7835), .A2(n7768), .ZN(n7798) );
  NOR2_X1 U8192 ( .A1(P3_ADDR_REG_10__SCAN_IN), .A2(n7834), .ZN(n7768) );
  AOI22_X1 U8193 ( .A1(P3_ADDR_REG_13__SCAN_IN), .A2(n7792), .B1(n7794), .B2(
        n7772), .ZN(n7790) );
  INV_X1 U8194 ( .A(P3_ADDR_REG_19__SCAN_IN), .ZN(n8232) );
  INV_X1 U8195 ( .A(n13357), .ZN(n11640) );
  OAI21_X1 U8196 ( .B1(n13289), .B2(n6914), .A(n6912), .ZN(n13245) );
  AOI21_X1 U8197 ( .B1(n13324), .B2(n6913), .A(n6778), .ZN(n6912) );
  INV_X1 U8198 ( .A(n13324), .ZN(n6914) );
  INV_X1 U8199 ( .A(n13194), .ZN(n6913) );
  NAND2_X1 U8200 ( .A1(n13245), .A2(n13244), .ZN(n13243) );
  OR2_X1 U8201 ( .A1(n6678), .A2(n8127), .ZN(n9449) );
  AND4_X1 U8202 ( .A1(n9270), .A2(n9269), .A3(n9268), .A4(n9267), .ZN(n13693)
         );
  AND4_X1 U8203 ( .A1(n9215), .A2(n9214), .A3(n9213), .A4(n9212), .ZN(n12230)
         );
  AOI21_X1 U8204 ( .B1(n10017), .B2(n6668), .A(n9233), .ZN(n15318) );
  OR2_X1 U8205 ( .A1(n6678), .A2(n9373), .ZN(n9374) );
  OR2_X1 U8206 ( .A1(n6678), .A2(n13849), .ZN(n9423) );
  INV_X1 U8207 ( .A(n13680), .ZN(n13707) );
  INV_X1 U8208 ( .A(n12050), .ZN(n12145) );
  AOI21_X1 U8209 ( .B1(n9388), .B2(P3_REG1_REG_9__SCAN_IN), .A(n6703), .ZN(
        n7633) );
  NAND2_X1 U8210 ( .A1(n10822), .A2(n15697), .ZN(n11189) );
  XNOR2_X1 U8211 ( .A(n11971), .B(n11977), .ZN(n11901) );
  NOR2_X1 U8212 ( .A1(n11901), .A2(n12052), .ZN(n11972) );
  NAND2_X1 U8213 ( .A1(n13513), .A2(P3_REG2_REG_18__SCAN_IN), .ZN(n6997) );
  INV_X1 U8214 ( .A(n13512), .ZN(n6873) );
  NOR2_X1 U8215 ( .A1(n6836), .A2(n7530), .ZN(n7529) );
  NAND2_X1 U8216 ( .A1(n13471), .A2(n7524), .ZN(n7522) );
  OR2_X1 U8217 ( .A1(n10773), .A2(n10760), .ZN(n15694) );
  NAND2_X1 U8218 ( .A1(n13545), .A2(n9728), .ZN(n13532) );
  AOI21_X1 U8219 ( .B1(n13721), .B2(n13554), .A(n7009), .ZN(n13722) );
  INV_X1 U8220 ( .A(n13555), .ZN(n7009) );
  INV_X1 U8221 ( .A(n13714), .ZN(n15707) );
  AND2_X1 U8222 ( .A1(n9769), .A2(n10926), .ZN(n15715) );
  NAND2_X1 U8223 ( .A1(n13556), .A2(n6989), .ZN(n6988) );
  INV_X1 U8224 ( .A(n13825), .ZN(n6989) );
  AND2_X1 U8225 ( .A1(n9385), .A2(n9384), .ZN(n13797) );
  AND2_X1 U8226 ( .A1(n9750), .A2(n9749), .ZN(n13827) );
  NAND2_X1 U8227 ( .A1(n6897), .A2(n6888), .ZN(n6887) );
  NOR2_X1 U8228 ( .A1(n6891), .A2(n6890), .ZN(n6889) );
  NOR2_X1 U8229 ( .A1(n9682), .A2(n9025), .ZN(n6888) );
  INV_X1 U8230 ( .A(P3_IR_REG_19__SCAN_IN), .ZN(n9327) );
  NAND2_X1 U8231 ( .A1(n14329), .A2(n15350), .ZN(n12853) );
  NOR2_X1 U8232 ( .A1(n6699), .A2(n13935), .ZN(n7569) );
  NAND2_X1 U8233 ( .A1(n7572), .A2(n7576), .ZN(n7571) );
  OR2_X1 U8234 ( .A1(n12846), .A2(n7577), .ZN(n7576) );
  INV_X1 U8235 ( .A(n8826), .ZN(n7577) );
  OR2_X1 U8236 ( .A1(n8786), .A2(n8787), .ZN(n7036) );
  NAND2_X1 U8237 ( .A1(n8546), .A2(n8545), .ZN(n12959) );
  AND2_X1 U8238 ( .A1(n10075), .A2(n10081), .ZN(n13951) );
  OR2_X1 U8239 ( .A1(n13165), .A2(n13164), .ZN(n6856) );
  NAND2_X1 U8240 ( .A1(n8817), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n7545) );
  AND3_X1 U8241 ( .A1(n8353), .A2(n8354), .A3(n8355), .ZN(n7544) );
  AND2_X1 U8242 ( .A1(n14032), .A2(n8816), .ZN(n14049) );
  NAND2_X1 U8243 ( .A1(n7169), .A2(n7173), .ZN(n14042) );
  NAND2_X1 U8244 ( .A1(n8682), .A2(n8681), .ZN(n14295) );
  NAND2_X1 U8245 ( .A1(n7424), .A2(n8922), .ZN(n14197) );
  AND2_X1 U8246 ( .A1(n7174), .A2(n14041), .ZN(n7172) );
  OAI21_X1 U8247 ( .B1(n7173), .B2(n7171), .A(n6774), .ZN(n7170) );
  AOI21_X1 U8248 ( .B1(n7534), .B2(n7533), .A(n7176), .ZN(n14055) );
  AND2_X1 U8249 ( .A1(n8868), .A2(P2_STATE_REG_SCAN_IN), .ZN(n15635) );
  INV_X1 U8250 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n8225) );
  AND2_X1 U8251 ( .A1(n14417), .A2(n14415), .ZN(n7394) );
  AND4_X1 U8252 ( .A1(n12354), .A2(n12353), .A3(n12352), .A4(n12351), .ZN(
        n15372) );
  NAND2_X1 U8253 ( .A1(n11770), .A2(n7392), .ZN(n6998) );
  NAND2_X1 U8254 ( .A1(n11937), .A2(n11936), .ZN(n12654) );
  NAND2_X1 U8255 ( .A1(n10657), .A2(n9899), .ZN(n9924) );
  AND4_X1 U8256 ( .A1(n12525), .A2(n12524), .A3(n12523), .A4(n12522), .ZN(
        n14562) );
  NOR2_X1 U8257 ( .A1(n9863), .A2(n9878), .ZN(n10578) );
  AND2_X1 U8258 ( .A1(n9862), .A2(n9861), .ZN(n9863) );
  NAND2_X1 U8259 ( .A1(n6923), .A2(n6920), .ZN(n10577) );
  NAND2_X1 U8260 ( .A1(n10438), .A2(n10437), .ZN(n6923) );
  NAND2_X1 U8261 ( .A1(n6922), .A2(n6921), .ZN(n6920) );
  NAND2_X1 U8262 ( .A1(n11082), .A2(n11081), .ZN(n7400) );
  NAND2_X1 U8263 ( .A1(n12067), .A2(n12068), .ZN(n12069) );
  INV_X1 U8264 ( .A(n15014), .ZN(n15180) );
  AND2_X1 U8265 ( .A1(n9936), .A2(n15058), .ZN(n14683) );
  INV_X1 U8266 ( .A(n15392), .ZN(n14675) );
  AND2_X1 U8267 ( .A1(n12763), .A2(n12762), .ZN(n15103) );
  OR2_X1 U8268 ( .A1(n13093), .A2(n9889), .ZN(n12763) );
  INV_X1 U8269 ( .A(n14866), .ZN(n15121) );
  AOI21_X1 U8270 ( .B1(n15118), .B2(n15080), .A(n14863), .ZN(n14864) );
  NAND2_X1 U8271 ( .A1(n15163), .A2(n12544), .ZN(n14962) );
  INV_X1 U8272 ( .A(n12593), .ZN(n15048) );
  OR2_X1 U8273 ( .A1(n9935), .A2(n10684), .ZN(n15058) );
  AND2_X1 U8274 ( .A1(n6736), .A2(n9817), .ZN(n7721) );
  XNOR2_X1 U8275 ( .A(n7825), .B(n7822), .ZN(n15256) );
  OR2_X1 U8276 ( .A1(n15256), .A2(n15257), .ZN(n7230) );
  OR2_X1 U8277 ( .A1(n15263), .A2(n7135), .ZN(n7132) );
  AND2_X1 U8278 ( .A1(n15263), .A2(n7135), .ZN(n7133) );
  INV_X1 U8279 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n7135) );
  NAND2_X1 U8280 ( .A1(n15429), .A2(n15430), .ZN(n15428) );
  NAND2_X1 U8281 ( .A1(n7121), .A2(n15428), .ZN(n15433) );
  OAI21_X1 U8282 ( .B1(n15429), .B2(n15430), .A(n7122), .ZN(n7121) );
  INV_X1 U8283 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n7122) );
  NAND2_X1 U8284 ( .A1(n7129), .A2(n7128), .ZN(n7237) );
  INV_X1 U8285 ( .A(n15248), .ZN(n7128) );
  INV_X1 U8286 ( .A(n15247), .ZN(n7129) );
  AND2_X1 U8287 ( .A1(n10689), .A2(n6669), .ZN(n12608) );
  NAND2_X1 U8288 ( .A1(n7589), .A2(n6802), .ZN(n7585) );
  INV_X1 U8289 ( .A(n12921), .ZN(n7603) );
  INV_X1 U8290 ( .A(n12920), .ZN(n7604) );
  MUX2_X1 U8291 ( .A(n14705), .B(n12620), .S(n12789), .Z(n12621) );
  MUX2_X1 U8292 ( .A(n14703), .B(n12633), .S(n12789), .Z(n12634) );
  AOI21_X1 U8293 ( .B1(n7058), .B2(n6756), .A(n6686), .ZN(n7056) );
  MUX2_X1 U8294 ( .A(n14701), .B(n12641), .S(n12789), .Z(n12642) );
  NAND2_X1 U8295 ( .A1(n7549), .A2(n7546), .ZN(n12943) );
  INV_X1 U8296 ( .A(n12936), .ZN(n7553) );
  AOI21_X1 U8297 ( .B1(n7083), .B2(n7086), .A(n7707), .ZN(n7082) );
  NOR2_X1 U8298 ( .A1(n7085), .A2(n12651), .ZN(n7086) );
  OAI22_X1 U8299 ( .A1(n7605), .A2(n12956), .B1(n7606), .B2(n12963), .ZN(
        n12970) );
  INV_X1 U8300 ( .A(n12962), .ZN(n7606) );
  OAI21_X1 U8301 ( .B1(n12955), .B2(n12954), .A(n6753), .ZN(n7605) );
  INV_X1 U8302 ( .A(n13011), .ZN(n7611) );
  NAND2_X1 U8303 ( .A1(n12707), .A2(n12706), .ZN(n12711) );
  AND2_X1 U8304 ( .A1(n12705), .A2(n12704), .ZN(n12706) );
  NAND2_X1 U8305 ( .A1(n12703), .A2(n15032), .ZN(n12704) );
  AOI21_X1 U8306 ( .B1(n7610), .B2(n7609), .A(n6771), .ZN(n7608) );
  NOR2_X1 U8307 ( .A1(n6723), .A2(n7611), .ZN(n7610) );
  NAND2_X1 U8308 ( .A1(n6723), .A2(n7611), .ZN(n7609) );
  INV_X1 U8309 ( .A(n13026), .ZN(n7584) );
  AOI21_X1 U8310 ( .B1(n7067), .B2(n6702), .A(n6781), .ZN(n7066) );
  NOR2_X1 U8311 ( .A1(n13049), .A2(n13050), .ZN(n7614) );
  INV_X1 U8312 ( .A(n13049), .ZN(n7613) );
  NAND2_X1 U8313 ( .A1(n12749), .A2(n7080), .ZN(n7078) );
  NAND2_X1 U8314 ( .A1(n12750), .A2(n12748), .ZN(n7079) );
  INV_X1 U8315 ( .A(n12751), .ZN(n7713) );
  NAND2_X1 U8316 ( .A1(n7745), .A2(n7596), .ZN(n7595) );
  OAI22_X1 U8317 ( .A1(n13071), .A2(n13070), .B1(n13075), .B2(n13076), .ZN(
        n7596) );
  AND2_X1 U8318 ( .A1(n8310), .A2(SI_26_), .ZN(n7675) );
  INV_X1 U8319 ( .A(P3_ADDR_REG_1__SCAN_IN), .ZN(n8102) );
  NAND2_X1 U8320 ( .A1(n9723), .A2(n13548), .ZN(n9724) );
  AND2_X1 U8321 ( .A1(n9701), .A2(n11998), .ZN(n9706) );
  NAND2_X1 U8322 ( .A1(n8770), .A2(n7564), .ZN(n7559) );
  NAND2_X1 U8323 ( .A1(n13102), .A2(n13101), .ZN(n13109) );
  INV_X1 U8324 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n8191) );
  INV_X1 U8325 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n8190) );
  INV_X1 U8326 ( .A(n7675), .ZN(n7670) );
  NAND2_X1 U8327 ( .A1(n8280), .A2(n6846), .ZN(n6848) );
  NOR2_X1 U8328 ( .A1(n6847), .A2(n8283), .ZN(n6846) );
  INV_X1 U8329 ( .A(n7223), .ZN(n7222) );
  OAI21_X1 U8330 ( .B1(n7226), .B2(n7224), .A(n7227), .ZN(n7223) );
  AND2_X1 U8331 ( .A1(n8273), .A2(n8275), .ZN(n7227) );
  NOR2_X1 U8332 ( .A1(n10715), .A2(P1_IR_REG_15__SCAN_IN), .ZN(n9845) );
  OR2_X1 U8333 ( .A1(n8272), .A2(n10016), .ZN(n7226) );
  NAND2_X1 U8334 ( .A1(n8272), .A2(n10016), .ZN(n7225) );
  INV_X1 U8335 ( .A(n7735), .ZN(n7205) );
  NAND2_X1 U8336 ( .A1(n8268), .A2(n9999), .ZN(n8271) );
  AOI21_X1 U8337 ( .B1(n8394), .B2(n8246), .A(n8410), .ZN(n7661) );
  INV_X1 U8338 ( .A(n13341), .ZN(n6909) );
  NAND2_X1 U8339 ( .A1(n7485), .A2(n10767), .ZN(n10769) );
  NAND2_X1 U8340 ( .A1(n10771), .A2(n6956), .ZN(n10772) );
  OR2_X1 U8341 ( .A1(n10801), .A2(P3_REG1_REG_4__SCAN_IN), .ZN(n6956) );
  NAND2_X1 U8342 ( .A1(n10847), .A2(n10756), .ZN(n7408) );
  INV_X1 U8343 ( .A(n10789), .ZN(n7507) );
  NAND2_X1 U8344 ( .A1(n7512), .A2(n10986), .ZN(n7511) );
  INV_X1 U8345 ( .A(n7513), .ZN(n7512) );
  NAND2_X1 U8346 ( .A1(n7513), .A2(n7510), .ZN(n7509) );
  NOR2_X1 U8347 ( .A1(n13467), .A2(n13466), .ZN(n13500) );
  AND2_X1 U8348 ( .A1(n9483), .A2(n13533), .ZN(n9509) );
  NOR2_X1 U8349 ( .A1(n9396), .A2(P3_REG3_REG_24__SCAN_IN), .ZN(n9410) );
  INV_X1 U8350 ( .A(n9623), .ZN(n7479) );
  NAND2_X1 U8351 ( .A1(n9236), .A2(n9235), .ZN(n9249) );
  OR2_X1 U8352 ( .A1(n9173), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n9192) );
  AND2_X1 U8353 ( .A1(n12016), .A2(n9703), .ZN(n12000) );
  OR2_X1 U8354 ( .A1(n9704), .A2(n12031), .ZN(n12001) );
  NAND2_X1 U8355 ( .A1(n12017), .A2(n11893), .ZN(n9573) );
  NAND2_X1 U8356 ( .A1(n7619), .A2(n11221), .ZN(n11422) );
  INV_X1 U8357 ( .A(n9698), .ZN(n7620) );
  INV_X1 U8358 ( .A(n11171), .ZN(n10999) );
  AND2_X1 U8359 ( .A1(n7659), .A2(n7658), .ZN(n7657) );
  NOR2_X1 U8360 ( .A1(P3_IR_REG_28__SCAN_IN), .A2(P3_IR_REG_25__SCAN_IN), .ZN(
        n7658) );
  NAND2_X1 U8361 ( .A1(n15236), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n7337) );
  AND2_X1 U8362 ( .A1(n7338), .A2(n7337), .ZN(n7336) );
  NAND2_X1 U8363 ( .A1(P3_IR_REG_27__SCAN_IN), .A2(P3_IR_REG_31__SCAN_IN), 
        .ZN(n6896) );
  AND2_X1 U8364 ( .A1(n9013), .A2(n9026), .ZN(n6895) );
  INV_X1 U8365 ( .A(P3_IR_REG_22__SCAN_IN), .ZN(n9008) );
  NAND2_X1 U8366 ( .A1(n7109), .A2(n7108), .ZN(n9404) );
  NAND2_X1 U8367 ( .A1(n7110), .A2(n6712), .ZN(n7108) );
  NAND2_X1 U8368 ( .A1(n7310), .A2(n9340), .ZN(n9353) );
  NAND2_X1 U8369 ( .A1(P1_DATAO_REG_19__SCAN_IN), .A2(n11316), .ZN(n9340) );
  NOR2_X1 U8370 ( .A1(n7559), .A2(n8755), .ZN(n7555) );
  INV_X1 U8371 ( .A(n8770), .ZN(n7560) );
  OR2_X1 U8372 ( .A1(n7559), .A2(n7557), .ZN(n7556) );
  NAND2_X1 U8373 ( .A1(n6859), .A2(n6858), .ZN(n7590) );
  INV_X1 U8374 ( .A(n7592), .ZN(n6859) );
  OR2_X1 U8375 ( .A1(n7592), .A2(n7594), .ZN(n7591) );
  AND2_X1 U8376 ( .A1(n6694), .A2(n6796), .ZN(n7594) );
  NAND2_X1 U8377 ( .A1(n13071), .A2(n13070), .ZN(n7597) );
  NAND2_X1 U8378 ( .A1(n8817), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n8340) );
  NAND2_X1 U8379 ( .A1(n8817), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n8332) );
  NAND2_X1 U8380 ( .A1(n14074), .A2(n7147), .ZN(n7148) );
  NOR2_X1 U8381 ( .A1(n7149), .A2(n14329), .ZN(n7147) );
  OR2_X1 U8382 ( .A1(n14031), .A2(n14247), .ZN(n7149) );
  AND2_X1 U8383 ( .A1(n14152), .A2(n6707), .ZN(n14090) );
  AND2_X1 U8384 ( .A1(n14132), .A2(n6704), .ZN(n7143) );
  NOR2_X1 U8385 ( .A1(n14192), .A2(n14289), .ZN(n14152) );
  NOR2_X1 U8386 ( .A1(n12980), .A2(n14376), .ZN(n7152) );
  NOR2_X1 U8387 ( .A1(n8611), .A2(n12258), .ZN(n8610) );
  CLKBUF_X1 U8388 ( .A(n10384), .Z(n6962) );
  INV_X1 U8389 ( .A(n14104), .ZN(n7179) );
  NAND2_X1 U8390 ( .A1(n8889), .A2(n7536), .ZN(n7535) );
  INV_X1 U8391 ( .A(n7182), .ZN(n7181) );
  OR2_X1 U8392 ( .A1(n14207), .A2(n14295), .ZN(n14192) );
  NAND3_X1 U8393 ( .A1(n12109), .A2(n7151), .A3(n6689), .ZN(n14207) );
  NAND2_X1 U8394 ( .A1(n12109), .A2(n6689), .ZN(n14231) );
  INV_X1 U8395 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n8857) );
  INV_X1 U8396 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n7617) );
  INV_X1 U8397 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n8197) );
  INV_X1 U8398 ( .A(n7380), .ZN(n7379) );
  OAI21_X1 U8399 ( .B1(n14462), .B2(n14570), .A(n14644), .ZN(n7380) );
  NAND2_X1 U8400 ( .A1(n7071), .A2(n7074), .ZN(n12774) );
  NAND2_X1 U8401 ( .A1(n12760), .A2(n7076), .ZN(n7074) );
  NAND2_X1 U8402 ( .A1(n7073), .A2(n7072), .ZN(n7071) );
  NOR2_X1 U8403 ( .A1(n7262), .A2(n14857), .ZN(n7260) );
  NOR2_X1 U8404 ( .A1(n14516), .A2(n14866), .ZN(n7199) );
  NOR2_X1 U8405 ( .A1(n15158), .A2(n14977), .ZN(n7196) );
  NAND2_X1 U8406 ( .A1(n15040), .A2(n12681), .ZN(n7249) );
  NOR2_X1 U8407 ( .A1(n15380), .A2(n15286), .ZN(n7191) );
  OR2_X1 U8408 ( .A1(n12809), .A2(n7352), .ZN(n7351) );
  INV_X1 U8409 ( .A(n12160), .ZN(n7352) );
  NAND2_X1 U8410 ( .A1(n7187), .A2(n7186), .ZN(n11840) );
  INV_X1 U8411 ( .A(n11569), .ZN(n7187) );
  AND2_X1 U8412 ( .A1(n7194), .A2(n7193), .ZN(n7192) );
  AND2_X1 U8413 ( .A1(n12678), .A2(n12677), .ZN(n15060) );
  NAND2_X1 U8414 ( .A1(n7282), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n7281) );
  OR2_X1 U8415 ( .A1(n8302), .A2(n8147), .ZN(n7679) );
  AND2_X1 U8416 ( .A1(n8302), .A2(n8147), .ZN(n7681) );
  NAND2_X1 U8417 ( .A1(n8743), .A2(n6715), .ZN(n7678) );
  NAND2_X1 U8418 ( .A1(n7215), .A2(n7212), .ZN(n8297) );
  INV_X1 U8419 ( .A(n7213), .ZN(n7212) );
  OAI21_X1 U8420 ( .B1(n6813), .B2(n7214), .A(n8295), .ZN(n7213) );
  NAND2_X1 U8421 ( .A1(n9796), .A2(n7385), .ZN(n7384) );
  INV_X1 U8422 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n7385) );
  XNOR2_X1 U8423 ( .A(n8297), .B(n9373), .ZN(n8296) );
  INV_X1 U8424 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n7720) );
  NAND2_X1 U8425 ( .A1(n9845), .A2(n7094), .ZN(n10667) );
  INV_X1 U8426 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n7094) );
  INV_X1 U8427 ( .A(n9845), .ZN(n10717) );
  NAND2_X1 U8428 ( .A1(n7211), .A2(n8263), .ZN(n7210) );
  INV_X1 U8429 ( .A(n8523), .ZN(n7211) );
  INV_X1 U8430 ( .A(n7209), .ZN(n7208) );
  OAI21_X1 U8431 ( .B1(n8261), .B2(n7210), .A(n8267), .ZN(n7209) );
  INV_X1 U8432 ( .A(n8256), .ZN(n7686) );
  OAI211_X1 U8433 ( .C1(n7421), .C2(n9982), .A(n6865), .B(n6864), .ZN(n8237)
         );
  OR2_X1 U8434 ( .A1(n7420), .A2(n9982), .ZN(n6865) );
  NAND2_X1 U8435 ( .A1(n7137), .A2(n7756), .ZN(n7757) );
  NAND2_X1 U8436 ( .A1(n7803), .A2(n15462), .ZN(n7137) );
  OAI21_X1 U8437 ( .B1(P1_ADDR_REG_6__SCAN_IN), .B2(n7761), .A(n7760), .ZN(
        n7762) );
  OAI21_X1 U8438 ( .B1(P1_ADDR_REG_9__SCAN_IN), .B2(n8083), .A(n7766), .ZN(
        n7767) );
  OAI21_X1 U8439 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(n11904), .A(n7769), .ZN(
        n7796) );
  INV_X1 U8440 ( .A(P3_REG3_REG_8__SCAN_IN), .ZN(n10983) );
  NAND2_X1 U8441 ( .A1(n6973), .A2(n9041), .ZN(n6884) );
  INV_X1 U8442 ( .A(P3_REG3_REG_5__SCAN_IN), .ZN(n10889) );
  INV_X1 U8443 ( .A(P3_REG3_REG_17__SCAN_IN), .ZN(n9297) );
  INV_X1 U8444 ( .A(n11299), .ZN(n6917) );
  INV_X1 U8445 ( .A(n11614), .ZN(n6974) );
  CLKBUF_X1 U8446 ( .A(n15716), .Z(n6935) );
  INV_X1 U8447 ( .A(n15718), .ZN(n10836) );
  OR2_X1 U8448 ( .A1(n9474), .A2(n7483), .ZN(n7482) );
  OR2_X1 U8449 ( .A1(n9435), .A2(SI_2_), .ZN(n7481) );
  OR2_X1 U8450 ( .A1(n9316), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n9331) );
  AOI21_X1 U8451 ( .B1(n7290), .B2(n7293), .A(n6739), .ZN(n7288) );
  INV_X1 U8452 ( .A(n13185), .ZN(n7293) );
  INV_X1 U8453 ( .A(n13315), .ZN(n13343) );
  INV_X1 U8454 ( .A(n9732), .ZN(n7311) );
  NOR2_X1 U8455 ( .A1(n9672), .A2(n10591), .ZN(n7101) );
  NAND2_X1 U8456 ( .A1(n9667), .A2(n7117), .ZN(n9670) );
  AND4_X1 U8457 ( .A1(n9113), .A2(n9112), .A3(n9111), .A4(n9110), .ZN(n11602)
         );
  NAND2_X1 U8458 ( .A1(n6952), .A2(P3_REG2_REG_1__SCAN_IN), .ZN(n10815) );
  NAND2_X1 U8459 ( .A1(n11194), .A2(P3_REG1_REG_2__SCAN_IN), .ZN(n10761) );
  OR2_X1 U8460 ( .A1(n11194), .A2(P3_REG1_REG_2__SCAN_IN), .ZN(n10762) );
  INV_X1 U8461 ( .A(P3_ADDR_REG_3__SCAN_IN), .ZN(n8121) );
  NAND2_X1 U8462 ( .A1(n10848), .A2(P3_REG2_REG_3__SCAN_IN), .ZN(n10847) );
  NAND2_X1 U8463 ( .A1(n10846), .A2(P3_REG1_REG_3__SCAN_IN), .ZN(n10845) );
  INV_X1 U8464 ( .A(n7406), .ZN(n10800) );
  INV_X1 U8465 ( .A(n7408), .ZN(n10759) );
  AND2_X1 U8466 ( .A1(n6870), .A2(n6738), .ZN(n10805) );
  INV_X1 U8467 ( .A(n7404), .ZN(n10803) );
  NOR2_X1 U8468 ( .A1(n10805), .A2(n10804), .ZN(n10868) );
  AND2_X1 U8469 ( .A1(n10979), .A2(n10986), .ZN(n7003) );
  NOR2_X1 U8470 ( .A1(n10809), .A2(n9109), .ZN(n7513) );
  INV_X1 U8471 ( .A(n6954), .ZN(n11444) );
  INV_X1 U8472 ( .A(P3_ADDR_REG_11__SCAN_IN), .ZN(n11904) );
  OAI21_X1 U8473 ( .B1(n11913), .B2(n7519), .A(n7514), .ZN(n11915) );
  NOR2_X1 U8474 ( .A1(n11909), .A2(n11908), .ZN(n11985) );
  NOR2_X1 U8475 ( .A1(n13370), .A2(n7004), .ZN(n13400) );
  NAND2_X1 U8476 ( .A1(n7006), .A2(n7005), .ZN(n7004) );
  INV_X1 U8477 ( .A(n13369), .ZN(n7005) );
  INV_X1 U8478 ( .A(n13368), .ZN(n7006) );
  AND2_X1 U8479 ( .A1(n7491), .A2(n6786), .ZN(n13392) );
  NOR2_X1 U8480 ( .A1(n13392), .A2(n13396), .ZN(n13426) );
  OR2_X1 U8481 ( .A1(n13410), .A2(n13411), .ZN(n6953) );
  NOR2_X1 U8482 ( .A1(n13421), .A2(n13420), .ZN(n13439) );
  NOR2_X1 U8483 ( .A1(n13426), .A2(n13425), .ZN(n13434) );
  INV_X1 U8484 ( .A(n7526), .ZN(n7523) );
  NAND2_X1 U8485 ( .A1(n7525), .A2(n7527), .ZN(n7524) );
  NAND2_X1 U8486 ( .A1(n7528), .A2(n13525), .ZN(n7527) );
  INV_X1 U8487 ( .A(n13506), .ZN(n7528) );
  INV_X1 U8488 ( .A(n13526), .ZN(n7530) );
  NAND2_X1 U8489 ( .A1(n7455), .A2(n7457), .ZN(n9738) );
  AOI21_X1 U8490 ( .B1(n7458), .B2(n7462), .A(n7456), .ZN(n7455) );
  INV_X1 U8491 ( .A(n9663), .ZN(n7456) );
  NOR2_X1 U8492 ( .A1(n9510), .A2(n9509), .ZN(n9739) );
  NAND2_X1 U8493 ( .A1(n7464), .A2(n9662), .ZN(n7461) );
  NAND2_X1 U8494 ( .A1(n13552), .A2(n7465), .ZN(n7464) );
  NAND2_X1 U8495 ( .A1(n7466), .A2(n9657), .ZN(n7465) );
  INV_X1 U8496 ( .A(n9656), .ZN(n7466) );
  NAND2_X1 U8497 ( .A1(n9662), .A2(n9657), .ZN(n7462) );
  AND2_X1 U8498 ( .A1(n9523), .A2(n9728), .ZN(n7621) );
  AND2_X1 U8499 ( .A1(n9666), .A2(n9663), .ZN(n13537) );
  OR2_X1 U8500 ( .A1(n13338), .A2(n13548), .ZN(n9656) );
  AND2_X1 U8501 ( .A1(n9660), .A2(n9662), .ZN(n13552) );
  NAND2_X1 U8502 ( .A1(n13591), .A2(n9533), .ZN(n13573) );
  INV_X1 U8503 ( .A(n7650), .ZN(n7649) );
  OAI21_X1 U8504 ( .B1(n7653), .B2(n7651), .A(n9716), .ZN(n7650) );
  AOI21_X1 U8505 ( .B1(n7637), .B2(n6698), .A(n6783), .ZN(n13678) );
  NOR2_X1 U8506 ( .A1(n9264), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n9280) );
  NAND2_X1 U8507 ( .A1(n9227), .A2(n9598), .ZN(n12197) );
  NOR2_X1 U8508 ( .A1(n9209), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n9236) );
  NAND2_X1 U8509 ( .A1(n7629), .A2(n7628), .ZN(n12088) );
  AOI21_X1 U8510 ( .B1(n7469), .B2(n7471), .A(n6776), .ZN(n7468) );
  AND2_X1 U8511 ( .A1(n12005), .A2(n12001), .ZN(n12002) );
  AND2_X1 U8512 ( .A1(n12034), .A2(n12030), .ZN(n12031) );
  OAI21_X1 U8513 ( .B1(n7447), .B2(n7448), .A(n9562), .ZN(n11789) );
  NOR2_X1 U8514 ( .A1(n11219), .A2(n7449), .ZN(n7447) );
  INV_X1 U8515 ( .A(n9088), .ZN(n7449) );
  AND2_X1 U8516 ( .A1(n9570), .A2(n9568), .ZN(n11790) );
  OR2_X1 U8517 ( .A1(n9107), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n9121) );
  NAND2_X1 U8518 ( .A1(n11221), .A2(n9698), .ZN(n11424) );
  NAND2_X1 U8519 ( .A1(n11223), .A2(n11222), .ZN(n11221) );
  INV_X1 U8520 ( .A(n11218), .ZN(n11222) );
  NAND2_X1 U8521 ( .A1(n15721), .A2(n15720), .ZN(n7618) );
  NAND2_X1 U8522 ( .A1(n9744), .A2(n9772), .ZN(n13554) );
  NAND2_X1 U8523 ( .A1(n11050), .A2(n11053), .ZN(n11049) );
  AND2_X1 U8524 ( .A1(n9766), .A2(n9765), .ZN(n10933) );
  INV_X1 U8525 ( .A(n11432), .ZN(n15753) );
  INV_X1 U8526 ( .A(n15316), .ZN(n15327) );
  INV_X1 U8527 ( .A(n15745), .ZN(n15769) );
  OR2_X1 U8528 ( .A1(n9474), .A2(n7734), .ZN(n6972) );
  OR2_X1 U8529 ( .A1(n9435), .A2(n9953), .ZN(n6971) );
  NAND2_X1 U8530 ( .A1(n9754), .A2(n9753), .ZN(n10592) );
  NAND2_X1 U8531 ( .A1(n13848), .A2(n12124), .ZN(n9753) );
  NAND2_X1 U8532 ( .A1(n9752), .A2(n9751), .ZN(n9754) );
  NAND2_X1 U8533 ( .A1(n7335), .A2(n7334), .ZN(n7333) );
  NAND2_X1 U8534 ( .A1(n6840), .A2(n7337), .ZN(n7334) );
  NAND2_X1 U8535 ( .A1(n7336), .A2(n9446), .ZN(n7335) );
  NOR2_X1 U8536 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(P3_IR_REG_28__SCAN_IN), .ZN(
        n6890) );
  NAND2_X1 U8537 ( .A1(n9678), .A2(n6764), .ZN(n6897) );
  NAND2_X1 U8538 ( .A1(P1_DATAO_REG_27__SCAN_IN), .A2(n7339), .ZN(n7338) );
  XNOR2_X1 U8539 ( .A(n9676), .B(n9675), .ZN(n10745) );
  INV_X1 U8540 ( .A(P3_IR_REG_23__SCAN_IN), .ZN(n9675) );
  OAI21_X1 U8541 ( .B1(n9674), .B2(P3_IR_REG_22__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n9676) );
  INV_X1 U8542 ( .A(P3_IR_REG_20__SCAN_IN), .ZN(n9506) );
  NAND2_X1 U8543 ( .A1(n9309), .A2(n9308), .ZN(n9322) );
  NAND2_X1 U8544 ( .A1(P1_DATAO_REG_17__SCAN_IN), .A2(n10671), .ZN(n9308) );
  NAND2_X1 U8545 ( .A1(n9307), .A2(n9306), .ZN(n9309) );
  NAND2_X1 U8546 ( .A1(n9275), .A2(n7307), .ZN(n7306) );
  INV_X1 U8547 ( .A(P3_IR_REG_15__SCAN_IN), .ZN(n9275) );
  INV_X1 U8548 ( .A(P3_IR_REG_16__SCAN_IN), .ZN(n9289) );
  AOI21_X1 U8549 ( .B1(n7321), .B2(n7323), .A(n6824), .ZN(n7319) );
  OR2_X1 U8550 ( .A1(n9244), .A2(n7322), .ZN(n7103) );
  INV_X1 U8551 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n9161) );
  XNOR2_X1 U8552 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(P2_DATAO_REG_8__SCAN_IN), 
        .ZN(n9159) );
  AOI211_X1 U8553 ( .C1(n9100), .C2(n6742), .A(n7095), .B(n6691), .ZN(n7097)
         );
  AND2_X1 U8554 ( .A1(n7324), .A2(n7096), .ZN(n7095) );
  XNOR2_X1 U8555 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .ZN(n9143) );
  INV_X1 U8556 ( .A(P3_IR_REG_6__SCAN_IN), .ZN(n9130) );
  XNOR2_X1 U8557 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(P2_DATAO_REG_4__SCAN_IN), 
        .ZN(n9097) );
  OAI211_X1 U8558 ( .C1(n7316), .C2(n7318), .A(n9059), .B(n7315), .ZN(n9076)
         );
  XNOR2_X1 U8559 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(P2_DATAO_REG_3__SCAN_IN), 
        .ZN(n9075) );
  AND2_X1 U8560 ( .A1(n9064), .A2(n9081), .ZN(n10768) );
  XNOR2_X1 U8561 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(P2_DATAO_REG_2__SCAN_IN), 
        .ZN(n9057) );
  XNOR2_X1 U8562 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .ZN(n9028) );
  OR2_X1 U8563 ( .A1(n8746), .A2(n8184), .ZN(n8761) );
  INV_X1 U8564 ( .A(n11121), .ZN(n7021) );
  AOI21_X1 U8565 ( .B1(n10721), .B2(n7017), .A(n7015), .ZN(n7014) );
  AND2_X1 U8566 ( .A1(n8730), .A2(n8706), .ZN(n7598) );
  INV_X1 U8567 ( .A(n13909), .ZN(n7562) );
  INV_X1 U8568 ( .A(n8754), .ZN(n7558) );
  INV_X1 U8569 ( .A(n13852), .ZN(n7565) );
  AOI21_X1 U8570 ( .B1(n7050), .B2(n7048), .A(n6730), .ZN(n7047) );
  INV_X1 U8571 ( .A(n7050), .ZN(n7049) );
  INV_X1 U8572 ( .A(n7052), .ZN(n7048) );
  OR2_X1 U8573 ( .A1(n8718), .A2(n13874), .ZN(n8746) );
  OR2_X1 U8574 ( .A1(n8513), .A2(n8512), .ZN(n8529) );
  OR2_X1 U8575 ( .A1(n8529), .A2(n8528), .ZN(n8548) );
  AND2_X1 U8576 ( .A1(n13169), .A2(n8321), .ZN(n10075) );
  AOI21_X1 U8577 ( .B1(n7430), .B2(n7428), .A(n6734), .ZN(n7427) );
  INV_X1 U8578 ( .A(n8987), .ZN(n7428) );
  NAND2_X1 U8579 ( .A1(n14152), .A2(n7143), .ZN(n14127) );
  NOR2_X1 U8580 ( .A1(n6692), .A2(n6746), .ZN(n14140) );
  NAND2_X1 U8581 ( .A1(n14152), .A2(n14158), .ZN(n14153) );
  AND2_X1 U8582 ( .A1(n7739), .A2(n8922), .ZN(n7423) );
  INV_X1 U8583 ( .A(n12211), .ZN(n7445) );
  OR2_X1 U8584 ( .A1(n8587), .A2(n12132), .ZN(n8611) );
  NAND2_X1 U8585 ( .A1(n12109), .A2(n8888), .ZN(n12205) );
  NAND2_X1 U8586 ( .A1(n7446), .A2(n12102), .ZN(n12213) );
  NAND2_X1 U8587 ( .A1(n7141), .A2(n15357), .ZN(n12110) );
  INV_X1 U8588 ( .A(n11811), .ZN(n7141) );
  AND2_X1 U8589 ( .A1(n13137), .A2(n8912), .ZN(n7422) );
  NAND2_X1 U8590 ( .A1(n8913), .A2(n8912), .ZN(n11805) );
  NAND2_X1 U8591 ( .A1(n8970), .A2(n8969), .ZN(n11620) );
  XNOR2_X1 U8592 ( .A(n12935), .B(n13981), .ZN(n13130) );
  OAI21_X1 U8593 ( .B1(n7155), .B2(n11515), .A(n7153), .ZN(n10908) );
  AOI21_X1 U8594 ( .B1(n13126), .B2(n7154), .A(n6768), .ZN(n7153) );
  INV_X1 U8595 ( .A(n8958), .ZN(n7154) );
  CLKBUF_X1 U8596 ( .A(n13123), .Z(n6961) );
  INV_X1 U8597 ( .A(n6961), .ZN(n10476) );
  AOI21_X1 U8598 ( .B1(n7174), .B2(n7176), .A(n6782), .ZN(n7173) );
  AND2_X1 U8599 ( .A1(n7439), .A2(n8949), .ZN(n7436) );
  NOR2_X1 U8600 ( .A1(n14037), .A2(n7440), .ZN(n7439) );
  AND2_X1 U8601 ( .A1(n14031), .A2(n15672), .ZN(n7440) );
  NAND2_X1 U8602 ( .A1(n14078), .A2(n8989), .ZN(n7533) );
  INV_X1 U8603 ( .A(n14071), .ZN(n7534) );
  NAND2_X1 U8604 ( .A1(n7180), .A2(n7177), .ZN(n14071) );
  INV_X1 U8605 ( .A(n7178), .ZN(n7177) );
  NAND2_X1 U8606 ( .A1(n14105), .A2(n7181), .ZN(n7180) );
  OAI21_X1 U8607 ( .B1(n7182), .B2(n7179), .A(n7535), .ZN(n7178) );
  NAND2_X1 U8608 ( .A1(n12204), .A2(n12212), .ZN(n12203) );
  INV_X1 U8609 ( .A(n13139), .ZN(n12212) );
  OR2_X1 U8610 ( .A1(n12967), .A2(n13976), .ZN(n7540) );
  NAND2_X1 U8611 ( .A1(n8992), .A2(n15675), .ZN(n15366) );
  NAND2_X1 U8612 ( .A1(n8365), .A2(n8364), .ZN(n8366) );
  OR2_X1 U8613 ( .A1(n8379), .A2(n9977), .ZN(n8368) );
  OR2_X1 U8614 ( .A1(n9976), .A2(n8358), .ZN(n8367) );
  INV_X1 U8615 ( .A(n15644), .ZN(n15672) );
  INV_X1 U8616 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n8208) );
  NAND2_X1 U8617 ( .A1(n14382), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8209) );
  INV_X1 U8618 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n8313) );
  INV_X1 U8619 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n8837) );
  INV_X1 U8620 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n8230) );
  CLKBUF_X1 U8621 ( .A(n8361), .Z(n8362) );
  INV_X1 U8622 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n9039) );
  AOI21_X1 U8623 ( .B1(n14525), .B2(n14522), .A(n14552), .ZN(n7374) );
  INV_X1 U8624 ( .A(n7374), .ZN(n7372) );
  NAND2_X1 U8625 ( .A1(n14463), .A2(n14462), .ZN(n14569) );
  AND2_X1 U8626 ( .A1(n14510), .A2(n14508), .ZN(n14581) );
  INV_X1 U8627 ( .A(n7398), .ZN(n7399) );
  INV_X1 U8628 ( .A(n12067), .ZN(n7393) );
  AOI21_X1 U8629 ( .B1(n14517), .B2(n14707), .A(n9877), .ZN(n10438) );
  OR2_X1 U8630 ( .A1(n12429), .A2(n14628), .ZN(n12439) );
  NOR2_X1 U8631 ( .A1(n11947), .A2(n11946), .ZN(n11948) );
  XNOR2_X1 U8632 ( .A(n9892), .B(n14445), .ZN(n9898) );
  OR2_X1 U8633 ( .A1(n12403), .A2(n12402), .ZN(n12405) );
  NOR2_X1 U8634 ( .A1(n12405), .A2(n10523), .ZN(n12418) );
  NAND2_X1 U8635 ( .A1(n14583), .A2(n14510), .ZN(n14664) );
  AND2_X1 U8636 ( .A1(n12349), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n12362) );
  NAND2_X1 U8637 ( .A1(n6677), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n9867) );
  NAND2_X1 U8638 ( .A1(n14899), .A2(n7198), .ZN(n14851) );
  AND2_X1 U8639 ( .A1(n6697), .A2(n12759), .ZN(n7198) );
  AND2_X1 U8640 ( .A1(n14899), .A2(n6697), .ZN(n12577) );
  NAND2_X1 U8641 ( .A1(n7257), .A2(n6687), .ZN(n14856) );
  AOI21_X1 U8642 ( .B1(n7367), .B2(n12547), .A(n6741), .ZN(n7365) );
  NAND2_X1 U8643 ( .A1(n14905), .A2(n7367), .ZN(n14896) );
  AOI21_X1 U8644 ( .B1(n14937), .B2(n14938), .A(n6725), .ZN(n14922) );
  NOR2_X1 U8645 ( .A1(n12439), .A2(n12438), .ZN(n12449) );
  NAND2_X1 U8646 ( .A1(n14986), .A2(n7194), .ZN(n14944) );
  NAND2_X1 U8647 ( .A1(n14986), .A2(n15166), .ZN(n14974) );
  OR2_X1 U8648 ( .A1(n7278), .A2(n7277), .ZN(n7276) );
  INV_X1 U8649 ( .A(n12424), .ZN(n7277) );
  AOI21_X1 U8650 ( .B1(n7359), .B2(n7357), .A(n7356), .ZN(n7355) );
  INV_X1 U8651 ( .A(n7359), .ZN(n7358) );
  INV_X1 U8652 ( .A(n7362), .ZN(n7357) );
  INV_X1 U8653 ( .A(n15192), .ZN(n7188) );
  NAND2_X1 U8654 ( .A1(n12360), .A2(n7189), .ZN(n15045) );
  AND2_X1 U8655 ( .A1(n15061), .A2(n12357), .ZN(n12358) );
  NAND2_X1 U8656 ( .A1(n12358), .A2(n12813), .ZN(n12534) );
  NOR2_X1 U8657 ( .A1(n12337), .A2(n12336), .ZN(n12349) );
  NAND2_X1 U8658 ( .A1(n12360), .A2(n12359), .ZN(n15290) );
  OR2_X1 U8659 ( .A1(n12289), .A2(n12288), .ZN(n12337) );
  AND2_X1 U8660 ( .A1(n11945), .A2(n12243), .ZN(n12162) );
  OR2_X1 U8661 ( .A1(n11402), .A2(n11401), .ZN(n11827) );
  OR2_X1 U8662 ( .A1(n11827), .A2(n11826), .ZN(n11947) );
  NOR2_X1 U8663 ( .A1(n11840), .A2(n12650), .ZN(n11945) );
  NAND2_X1 U8664 ( .A1(n11836), .A2(n11835), .ZN(n11943) );
  NAND2_X1 U8665 ( .A1(n11823), .A2(n11822), .ZN(n11825) );
  INV_X1 U8666 ( .A(n15069), .ZN(n15001) );
  AND2_X1 U8667 ( .A1(n10184), .A2(n9941), .ZN(n15002) );
  NAND2_X1 U8668 ( .A1(n7346), .A2(n7347), .ZN(n7345) );
  NAND2_X1 U8669 ( .A1(n11417), .A2(n11416), .ZN(n11834) );
  NAND2_X1 U8670 ( .A1(n11589), .A2(n15511), .ZN(n11569) );
  NOR2_X1 U8671 ( .A1(n11590), .A2(n12633), .ZN(n11589) );
  AND3_X1 U8672 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .A3(P1_REG3_REG_5__SCAN_IN), .ZN(n11039) );
  INV_X1 U8673 ( .A(n11584), .ZN(n15080) );
  OR2_X1 U8674 ( .A1(n11483), .A2(n12629), .ZN(n11590) );
  NAND2_X1 U8675 ( .A1(n11412), .A2(n11411), .ZN(n11480) );
  NAND2_X1 U8676 ( .A1(n11480), .A2(n12800), .ZN(n11482) );
  NAND2_X1 U8677 ( .A1(n11387), .A2(n7280), .ZN(n10950) );
  NAND2_X1 U8678 ( .A1(n14705), .A2(n11410), .ZN(n7280) );
  NAND2_X1 U8679 ( .A1(n10949), .A2(n10950), .ZN(n11412) );
  NAND2_X1 U8680 ( .A1(n11525), .A2(n7055), .ZN(n11524) );
  NAND2_X1 U8681 ( .A1(n12794), .A2(n15077), .ZN(n15079) );
  OR3_X1 U8682 ( .A1(n11201), .A2(n11200), .A3(n11199), .ZN(n12584) );
  NAND2_X1 U8683 ( .A1(n12471), .A2(n12470), .ZN(n15141) );
  INV_X1 U8684 ( .A(n15291), .ZN(n15488) );
  INV_X1 U8685 ( .A(n15413), .ZN(n15482) );
  NAND2_X1 U8686 ( .A1(n9904), .A2(n9903), .ZN(n10018) );
  XNOR2_X1 U8687 ( .A(n12781), .B(n12780), .ZN(n13083) );
  OAI21_X1 U8688 ( .B1(n12557), .B2(n7700), .A(n7697), .ZN(n12781) );
  XNOR2_X1 U8689 ( .A(n12557), .B(n12556), .ZN(n14386) );
  AOI21_X1 U8690 ( .B1(n6714), .B2(n7666), .A(n6831), .ZN(n7665) );
  INV_X1 U8691 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n9831) );
  NOR2_X1 U8692 ( .A1(n9837), .A2(n9836), .ZN(n9838) );
  OAI21_X1 U8693 ( .B1(n8772), .B2(n6714), .A(n7668), .ZN(n8809) );
  AND2_X1 U8694 ( .A1(n9808), .A2(n9833), .ZN(n9905) );
  OAI21_X1 U8695 ( .B1(n8772), .B2(n8771), .A(n8310), .ZN(n8789) );
  INV_X1 U8696 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n9797) );
  INV_X1 U8697 ( .A(n8296), .ZN(n8732) );
  XNOR2_X1 U8698 ( .A(n8715), .B(n8714), .ZN(n12435) );
  NAND2_X1 U8699 ( .A1(n8280), .A2(n8279), .ZN(n8640) );
  OR2_X1 U8700 ( .A1(n10243), .A2(n10242), .ZN(n10358) );
  NAND2_X1 U8701 ( .A1(n7660), .A2(n8246), .ZN(n8411) );
  NAND2_X1 U8702 ( .A1(n8395), .A2(n8244), .ZN(n7660) );
  INV_X1 U8703 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n7704) );
  NOR2_X1 U8704 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n9885) );
  XNOR2_X1 U8705 ( .A(n8237), .B(n9955), .ZN(n8346) );
  NAND2_X1 U8706 ( .A1(n7750), .A2(n7749), .ZN(n7807) );
  NAND2_X1 U8707 ( .A1(P3_ADDR_REG_1__SCAN_IN), .A2(n7748), .ZN(n7749) );
  INV_X1 U8708 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n7804) );
  NAND2_X1 U8709 ( .A1(n15792), .A2(n7830), .ZN(n7832) );
  AND2_X1 U8710 ( .A1(n7767), .A2(n10465), .ZN(n7834) );
  NOR2_X1 U8711 ( .A1(n7767), .A2(n10465), .ZN(n7835) );
  OAI21_X1 U8712 ( .B1(n15422), .B2(n15421), .A(n7232), .ZN(n7231) );
  INV_X1 U8713 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n7232) );
  OAI21_X1 U8714 ( .B1(P3_ADDR_REG_14__SCAN_IN), .B2(n10613), .A(n7773), .ZN(
        n7788) );
  AOI21_X1 U8715 ( .B1(n7298), .B2(n7300), .A(n6749), .ZN(n7295) );
  NAND2_X1 U8716 ( .A1(n13183), .A2(n13182), .ZN(n7289) );
  AND3_X1 U8717 ( .A1(n9189), .A2(n9188), .A3(n9187), .ZN(n15766) );
  INV_X1 U8718 ( .A(n6903), .ZN(n12140) );
  XNOR2_X1 U8719 ( .A(n11007), .B(n11224), .ZN(n10833) );
  INV_X1 U8720 ( .A(n13652), .ZN(n13629) );
  AND4_X1 U8721 ( .A1(n9127), .A2(n9126), .A3(n9125), .A4(n9124), .ZN(n11858)
         );
  NAND2_X1 U8722 ( .A1(n6880), .A2(n6885), .ZN(n10675) );
  INV_X1 U8723 ( .A(n6881), .ZN(n6880) );
  NAND2_X1 U8724 ( .A1(n13305), .A2(n13200), .ZN(n13262) );
  NAND2_X1 U8725 ( .A1(n9358), .A2(n9357), .ZN(n13267) );
  NAND2_X1 U8726 ( .A1(n9408), .A2(n9407), .ZN(n13581) );
  OR2_X1 U8727 ( .A1(n6678), .A2(n12178), .ZN(n9407) );
  AOI21_X1 U8728 ( .B1(n10434), .B2(n6668), .A(n9296), .ZN(n13295) );
  NOR2_X1 U8729 ( .A1(n13287), .A2(n7302), .ZN(n7301) );
  INV_X1 U8730 ( .A(n13192), .ZN(n7302) );
  NAND2_X1 U8731 ( .A1(n7303), .A2(n13192), .ZN(n13288) );
  AND2_X1 U8732 ( .A1(n9416), .A2(n9415), .ZN(n13590) );
  NAND2_X1 U8733 ( .A1(n11007), .A2(n10625), .ZN(n7294) );
  INV_X1 U8734 ( .A(n7309), .ZN(n11864) );
  NAND2_X1 U8735 ( .A1(n13307), .A2(n13306), .ZN(n13305) );
  AND4_X1 U8736 ( .A1(n9198), .A2(n9197), .A3(n9196), .A4(n9195), .ZN(n12377)
         );
  NAND2_X1 U8737 ( .A1(n10676), .A2(n10677), .ZN(n10832) );
  NAND2_X1 U8738 ( .A1(n6881), .A2(n6885), .ZN(n10676) );
  INV_X1 U8739 ( .A(n13308), .ZN(n13664) );
  NAND2_X1 U8740 ( .A1(n13325), .A2(n13324), .ZN(n13323) );
  NAND2_X1 U8741 ( .A1(n13289), .A2(n13194), .ZN(n13325) );
  NAND2_X1 U8742 ( .A1(n7297), .A2(n13216), .ZN(n13331) );
  NAND2_X1 U8743 ( .A1(n13270), .A2(n13271), .ZN(n7297) );
  NAND2_X1 U8744 ( .A1(n10512), .A2(n10934), .ZN(n13352) );
  NAND2_X1 U8745 ( .A1(n6907), .A2(n7288), .ZN(n13342) );
  NAND2_X1 U8746 ( .A1(n13183), .A2(n7290), .ZN(n6907) );
  AOI21_X1 U8747 ( .B1(n13557), .B2(n9300), .A(n9444), .ZN(n13565) );
  INV_X1 U8748 ( .A(n13590), .ZN(n13333) );
  AND3_X1 U8749 ( .A1(n9380), .A2(n9379), .A3(n9378), .ZN(n13630) );
  INV_X1 U8750 ( .A(n12230), .ZN(n13356) );
  INV_X1 U8751 ( .A(n12377), .ZN(n12223) );
  NAND4_X1 U8752 ( .A1(n9142), .A2(n9141), .A3(n9140), .A4(n9139), .ZN(n13357)
         );
  INV_X1 U8753 ( .A(n11858), .ZN(n12017) );
  INV_X1 U8754 ( .A(n11602), .ZN(n11751) );
  OR2_X1 U8755 ( .A1(n9346), .A2(n15689), .ZN(n9037) );
  NAND2_X1 U8756 ( .A1(n9138), .A2(P3_REG0_REG_0__SCAN_IN), .ZN(n9036) );
  OAI21_X1 U8757 ( .B1(n6945), .B2(n15690), .A(n7007), .ZN(n10728) );
  NAND2_X1 U8758 ( .A1(n6945), .A2(P3_REG1_REG_0__SCAN_IN), .ZN(n7007) );
  NAND2_X1 U8759 ( .A1(n7488), .A2(n10765), .ZN(n7490) );
  AND3_X2 U8760 ( .A1(n9051), .A2(n9061), .A3(n9050), .ZN(n11194) );
  OR2_X1 U8761 ( .A1(n9031), .A2(n6871), .ZN(n9051) );
  NAND2_X1 U8762 ( .A1(n9682), .A2(n9049), .ZN(n9050) );
  NAND2_X1 U8763 ( .A1(P3_IR_REG_2__SCAN_IN), .A2(P3_IR_REG_31__SCAN_IN), .ZN(
        n6871) );
  AOI21_X1 U8764 ( .B1(n11189), .B2(n11188), .A(n11187), .ZN(n11186) );
  NOR2_X1 U8765 ( .A1(n10788), .A2(n10883), .ZN(n10790) );
  INV_X1 U8766 ( .A(n6968), .ZN(n10987) );
  INV_X1 U8767 ( .A(n6995), .ZN(n10990) );
  INV_X1 U8768 ( .A(n7413), .ZN(n11330) );
  NOR2_X1 U8769 ( .A1(n11440), .A2(n11439), .ZN(n11443) );
  NOR2_X1 U8770 ( .A1(n11443), .A2(n11442), .ZN(n11913) );
  NOR2_X1 U8771 ( .A1(n11972), .A2(n11973), .ZN(n11976) );
  INV_X1 U8772 ( .A(n7491), .ZN(n13389) );
  NOR2_X1 U8773 ( .A1(n13384), .A2(n13385), .ZN(n13386) );
  NOR2_X1 U8774 ( .A1(n13386), .A2(n13397), .ZN(n13410) );
  NOR2_X1 U8775 ( .A1(n13412), .A2(n13413), .ZN(n13450) );
  XNOR2_X1 U8776 ( .A(n6953), .B(n13427), .ZN(n13412) );
  NAND2_X1 U8777 ( .A1(n6817), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9260) );
  NOR2_X1 U8778 ( .A1(n13449), .A2(n13434), .ZN(n13436) );
  NOR2_X1 U8779 ( .A1(n13428), .A2(n13429), .ZN(n13435) );
  OAI21_X1 U8780 ( .B1(n13428), .B2(n7498), .A(n7497), .ZN(n13467) );
  NAND2_X1 U8781 ( .A1(n7499), .A2(P3_REG1_REG_15__SCAN_IN), .ZN(n7498) );
  NAND2_X1 U8782 ( .A1(n13436), .A2(n7499), .ZN(n7497) );
  INV_X1 U8783 ( .A(n13437), .ZN(n7499) );
  OAI21_X1 U8784 ( .B1(n13478), .B2(n13477), .A(n13476), .ZN(n13479) );
  NOR2_X1 U8785 ( .A1(n13464), .A2(n13684), .ZN(n13486) );
  AOI21_X1 U8786 ( .B1(n7002), .B2(n7001), .A(n15692), .ZN(n13498) );
  NAND2_X1 U8787 ( .A1(n13496), .A2(n13497), .ZN(n7001) );
  INV_X1 U8788 ( .A(n13514), .ZN(n7002) );
  NOR2_X1 U8789 ( .A1(n13507), .A2(n13506), .ZN(n13522) );
  OAI21_X1 U8790 ( .B1(n13464), .B2(n7410), .A(n7409), .ZN(n13512) );
  NAND2_X1 U8791 ( .A1(n7411), .A2(P3_REG2_REG_17__SCAN_IN), .ZN(n7410) );
  INV_X1 U8792 ( .A(n13489), .ZN(n7411) );
  AND2_X1 U8793 ( .A1(n7636), .A2(n6716), .ZN(n13576) );
  CLKBUF_X1 U8794 ( .A(n13599), .Z(n13600) );
  NAND2_X1 U8795 ( .A1(n13624), .A2(n9718), .ZN(n13611) );
  CLKBUF_X1 U8796 ( .A(n13614), .Z(n13616) );
  CLKBUF_X1 U8797 ( .A(n13622), .Z(n13623) );
  NAND2_X1 U8798 ( .A1(n13757), .A2(n9623), .ZN(n13648) );
  NOR2_X1 U8799 ( .A1(n13660), .A2(n7655), .ZN(n13651) );
  NAND2_X1 U8800 ( .A1(n7480), .A2(n13662), .ZN(n13757) );
  INV_X1 U8801 ( .A(n13672), .ZN(n7480) );
  CLKBUF_X1 U8802 ( .A(n13675), .Z(n13676) );
  OAI21_X1 U8803 ( .B1(n9714), .B2(n7644), .A(n7641), .ZN(n13690) );
  CLKBUF_X1 U8804 ( .A(n13697), .Z(n13698) );
  NAND2_X1 U8805 ( .A1(n7640), .A2(n7646), .ZN(n13705) );
  NAND2_X1 U8806 ( .A1(n9714), .A2(n6720), .ZN(n7640) );
  NAND2_X1 U8807 ( .A1(n9714), .A2(n9713), .ZN(n12264) );
  NAND2_X1 U8808 ( .A1(n11997), .A2(n9593), .ZN(n12045) );
  INV_X1 U8809 ( .A(n7630), .ZN(n12047) );
  NAND2_X1 U8810 ( .A1(n12022), .A2(n9154), .ZN(n12029) );
  AND2_X1 U8811 ( .A1(n15733), .A2(n15703), .ZN(n13716) );
  NAND2_X1 U8812 ( .A1(n10938), .A2(n10937), .ZN(n13714) );
  INV_X1 U8813 ( .A(n15709), .ZN(n15727) );
  AND2_X1 U8814 ( .A1(n15311), .A2(n15310), .ZN(n15332) );
  INV_X1 U8815 ( .A(P3_REG0_REG_27__SCAN_IN), .ZN(n6969) );
  AOI21_X1 U8816 ( .B1(n12126), .B2(n9184), .A(n9395), .ZN(n13793) );
  INV_X1 U8817 ( .A(n13318), .ZN(n13801) );
  INV_X1 U8818 ( .A(n13267), .ZN(n13805) );
  AND2_X1 U8819 ( .A1(n9342), .A2(n9341), .ZN(n13809) );
  NAND2_X1 U8820 ( .A1(n9330), .A2(n9329), .ZN(n13813) );
  NAND2_X1 U8821 ( .A1(n9248), .A2(n9247), .ZN(n13824) );
  INV_X1 U8822 ( .A(n9693), .ZN(n10939) );
  XNOR2_X1 U8823 ( .A(n9492), .B(n9491), .ZN(n13829) );
  CLKBUF_X1 U8824 ( .A(n13830), .Z(n13831) );
  INV_X1 U8825 ( .A(SI_29_), .ZN(n13841) );
  INV_X1 U8826 ( .A(n9020), .ZN(n13842) );
  INV_X1 U8827 ( .A(n7333), .ZN(n7330) );
  OAI21_X1 U8828 ( .B1(n9445), .B2(n9446), .A(n7338), .ZN(n9457) );
  INV_X1 U8829 ( .A(n7115), .ZN(n9432) );
  OR2_X1 U8830 ( .A1(n9678), .A2(n6949), .ZN(n6948) );
  NAND2_X1 U8831 ( .A1(n7112), .A2(n7327), .ZN(n9394) );
  NAND2_X1 U8832 ( .A1(n9369), .A2(n6825), .ZN(n7112) );
  NAND2_X1 U8833 ( .A1(n7329), .A2(n9371), .ZN(n9383) );
  NAND2_X1 U8834 ( .A1(n9369), .A2(n9368), .ZN(n7329) );
  XNOR2_X1 U8835 ( .A(n9530), .B(P3_IR_REG_22__SCAN_IN), .ZN(n11285) );
  INV_X1 U8836 ( .A(SI_20_), .ZN(n10924) );
  INV_X1 U8837 ( .A(SI_19_), .ZN(n10544) );
  INV_X1 U8838 ( .A(SI_15_), .ZN(n10130) );
  NAND2_X1 U8839 ( .A1(n7320), .A2(n9257), .ZN(n9273) );
  NAND2_X1 U8840 ( .A1(n9256), .A2(n9255), .ZN(n7320) );
  INV_X1 U8841 ( .A(SI_13_), .ZN(n10016) );
  INV_X1 U8842 ( .A(SI_12_), .ZN(n9999) );
  XNOR2_X1 U8843 ( .A(n9186), .B(n9185), .ZN(n11914) );
  NAND2_X1 U8844 ( .A1(n7326), .A2(n9116), .ZN(n9129) );
  NAND2_X1 U8845 ( .A1(n9115), .A2(n9114), .ZN(n7326) );
  INV_X1 U8846 ( .A(P3_IR_REG_0__SCAN_IN), .ZN(n10763) );
  NAND2_X1 U8847 ( .A1(n7022), .A2(n7026), .ZN(n12130) );
  NAND2_X1 U8848 ( .A1(n8558), .A2(n7028), .ZN(n7022) );
  NAND2_X1 U8849 ( .A1(n11264), .A2(n8505), .ZN(n11308) );
  OR2_X1 U8850 ( .A1(n9980), .A2(n8358), .ZN(n7433) );
  OAI21_X1 U8851 ( .B1(n10076), .B2(n10166), .A(n8380), .ZN(n7432) );
  NAND2_X1 U8852 ( .A1(n7567), .A2(n8467), .ZN(n11122) );
  OAI211_X1 U8853 ( .C1(n7018), .C2(n7017), .A(n6829), .B(n10721), .ZN(n7567)
         );
  NAND2_X1 U8854 ( .A1(n8335), .A2(n7730), .ZN(n10404) );
  NAND2_X1 U8855 ( .A1(n13922), .A2(n8706), .ZN(n13870) );
  NAND2_X1 U8856 ( .A1(n13922), .A2(n7598), .ZN(n13871) );
  NAND2_X1 U8857 ( .A1(n12255), .A2(n8620), .ZN(n13886) );
  NAND2_X1 U8858 ( .A1(n7563), .A2(n7566), .ZN(n13908) );
  NAND2_X1 U8859 ( .A1(n8702), .A2(n13918), .ZN(n13922) );
  NAND2_X1 U8860 ( .A1(n8558), .A2(n11699), .ZN(n11964) );
  NAND2_X1 U8861 ( .A1(n11964), .A2(n11963), .ZN(n11962) );
  NAND2_X1 U8862 ( .A1(n13926), .A2(n7012), .ZN(n13927) );
  NAND2_X1 U8863 ( .A1(n7039), .A2(n8521), .ZN(n15343) );
  NOR2_X1 U8864 ( .A1(n15342), .A2(n7038), .ZN(n7037) );
  INV_X1 U8865 ( .A(n8521), .ZN(n7038) );
  NAND2_X1 U8866 ( .A1(n7041), .A2(n7043), .ZN(n13938) );
  AND2_X1 U8867 ( .A1(n7601), .A2(n7044), .ZN(n7043) );
  NAND2_X1 U8868 ( .A1(n13896), .A2(n7045), .ZN(n7044) );
  NAND2_X1 U8869 ( .A1(n13898), .A2(n8659), .ZN(n13937) );
  INV_X1 U8870 ( .A(n15354), .ZN(n13944) );
  INV_X1 U8871 ( .A(n15350), .ZN(n13958) );
  INV_X1 U8872 ( .A(n13171), .ZN(n6853) );
  NAND2_X1 U8873 ( .A1(n6933), .A2(n14082), .ZN(n14254) );
  NAND2_X1 U8874 ( .A1(n6934), .A2(n15617), .ZN(n6933) );
  OR2_X1 U8875 ( .A1(n14107), .A2(n7182), .ZN(n14088) );
  NAND2_X1 U8876 ( .A1(n14118), .A2(n7430), .ZN(n14099) );
  AND2_X1 U8877 ( .A1(n7166), .A2(n6727), .ZN(n14126) );
  NAND2_X1 U8878 ( .A1(n7158), .A2(n7161), .ZN(n14167) );
  NAND2_X1 U8879 ( .A1(n7160), .A2(n7159), .ZN(n7158) );
  NAND2_X1 U8880 ( .A1(n14222), .A2(n8983), .ZN(n14199) );
  NAND2_X1 U8881 ( .A1(n8976), .A2(n8975), .ZN(n11803) );
  NAND2_X1 U8882 ( .A1(n11369), .A2(n8909), .ZN(n11623) );
  NAND2_X1 U8883 ( .A1(n11105), .A2(n8901), .ZN(n10900) );
  NAND2_X1 U8884 ( .A1(n7155), .A2(n8958), .ZN(n11508) );
  INV_X1 U8885 ( .A(n14234), .ZN(n14134) );
  INV_X1 U8886 ( .A(n14157), .ZN(n14228) );
  OR2_X1 U8887 ( .A1(n15688), .A2(n8954), .ZN(n7437) );
  INV_X1 U8888 ( .A(n13152), .ZN(n6990) );
  AOI21_X1 U8889 ( .B1(n7436), .B2(n14220), .A(n7435), .ZN(n7434) );
  NAND2_X1 U8890 ( .A1(n8493), .A2(n8492), .ZN(n12940) );
  INV_X1 U8891 ( .A(n14020), .ZN(n14320) );
  INV_X1 U8892 ( .A(n14019), .ZN(n14325) );
  NAND2_X1 U8893 ( .A1(n7441), .A2(n6985), .ZN(n7229) );
  NOR2_X1 U8894 ( .A1(n6671), .A2(n15678), .ZN(n6985) );
  OR2_X1 U8895 ( .A1(n15680), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n7228) );
  NAND2_X1 U8896 ( .A1(n6931), .A2(n6930), .ZN(n14326) );
  INV_X1 U8897 ( .A(n6991), .ZN(n6930) );
  INV_X1 U8898 ( .A(n14245), .ZN(n6931) );
  NAND2_X1 U8899 ( .A1(n8986), .A2(n8985), .ZN(n14138) );
  NAND2_X1 U8900 ( .A1(n14201), .A2(n8984), .ZN(n14187) );
  NAND2_X1 U8901 ( .A1(n12099), .A2(n7542), .ZN(n12189) );
  AND2_X1 U8902 ( .A1(n12099), .A2(n8979), .ZN(n7738) );
  AND2_X1 U8903 ( .A1(n15680), .A2(n15672), .ZN(n14375) );
  OR2_X1 U8904 ( .A1(n8211), .A2(n8207), .ZN(n8215) );
  XNOR2_X1 U8905 ( .A(n8838), .B(n8837), .ZN(n14395) );
  OAI21_X1 U8906 ( .B1(n8836), .B2(P2_IR_REG_25__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n8838) );
  XNOR2_X1 U8907 ( .A(n8834), .B(n8833), .ZN(n12388) );
  INV_X1 U8908 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n12390) );
  NAND2_X1 U8909 ( .A1(n8832), .A2(n8836), .ZN(n12322) );
  INV_X1 U8910 ( .A(n8829), .ZN(n8832) );
  INV_X1 U8911 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n11848) );
  INV_X1 U8912 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n10238) );
  INV_X1 U8913 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n10002) );
  INV_X1 U8914 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n9996) );
  INV_X1 U8915 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n9985) );
  INV_X1 U8916 ( .A(n12637), .ZN(n15511) );
  NAND2_X1 U8917 ( .A1(n14634), .A2(n14415), .ZN(n15375) );
  INV_X1 U8918 ( .A(n14697), .ZN(n15373) );
  INV_X1 U8919 ( .A(n14705), .ZN(n11529) );
  NAND2_X1 U8920 ( .A1(n14543), .A2(n14451), .ZN(n14546) );
  NAND2_X1 U8921 ( .A1(n11764), .A2(n7000), .ZN(n6999) );
  INV_X1 U8922 ( .A(n11766), .ZN(n7000) );
  AND2_X1 U8923 ( .A1(n12278), .A2(n12277), .ZN(n15271) );
  NAND2_X1 U8924 ( .A1(n14672), .A2(n14427), .ZN(n14594) );
  INV_X1 U8925 ( .A(n14699), .ZN(n15386) );
  NAND2_X1 U8926 ( .A1(n12158), .A2(n12157), .ZN(n15398) );
  NAND2_X1 U8927 ( .A1(n10576), .A2(n9879), .ZN(n10658) );
  NAND2_X1 U8928 ( .A1(n10658), .A2(n10659), .ZN(n10657) );
  AND2_X1 U8929 ( .A1(n9932), .A2(n12844), .ZN(n15402) );
  NAND2_X1 U8930 ( .A1(n9934), .A2(n9923), .ZN(n15392) );
  NAND2_X1 U8931 ( .A1(n7388), .A2(n14440), .ZN(n14655) );
  NAND2_X1 U8932 ( .A1(n14574), .A2(n15002), .ZN(n15384) );
  INV_X1 U8933 ( .A(n15402), .ZN(n14680) );
  AND2_X1 U8934 ( .A1(n7694), .A2(n7693), .ZN(n7692) );
  NOR2_X1 U8935 ( .A1(n12831), .A2(n7695), .ZN(n7694) );
  AOI211_X1 U8936 ( .C1(n12827), .C2(n14848), .A(n12825), .B(n12790), .ZN(
        n12838) );
  AND4_X1 U8937 ( .A1(n10322), .A2(n10321), .A3(n10320), .A4(n10319), .ZN(
        n15385) );
  INV_X1 U8938 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n10531) );
  INV_X1 U8939 ( .A(n14844), .ZN(n15100) );
  NAND2_X1 U8940 ( .A1(n12570), .A2(n12569), .ZN(n12572) );
  NAND2_X1 U8941 ( .A1(n14862), .A2(n12550), .ZN(n12552) );
  NAND2_X1 U8942 ( .A1(n14889), .A2(n12491), .ZN(n14874) );
  OAI21_X1 U8943 ( .B1(n14953), .B2(n7252), .A(n7253), .ZN(n14927) );
  AND2_X1 U8944 ( .A1(n7256), .A2(n6737), .ZN(n14939) );
  NAND2_X1 U8945 ( .A1(n14953), .A2(n14963), .ZN(n7256) );
  INV_X1 U8946 ( .A(n14979), .ZN(n12543) );
  INV_X1 U8947 ( .A(n14978), .ZN(n6877) );
  NAND2_X1 U8948 ( .A1(n7279), .A2(n7278), .ZN(n14984) );
  AND2_X1 U8949 ( .A1(n7279), .A2(n6735), .ZN(n7740) );
  NAND2_X1 U8950 ( .A1(n14998), .A2(n14999), .ZN(n7279) );
  AND2_X1 U8951 ( .A1(n12413), .A2(n12412), .ZN(n15014) );
  NAND2_X1 U8952 ( .A1(n7361), .A2(n12540), .ZN(n14997) );
  NAND2_X1 U8953 ( .A1(n12537), .A2(n7362), .ZN(n7361) );
  NAND2_X1 U8954 ( .A1(n7243), .A2(n7247), .ZN(n15020) );
  NAND2_X1 U8955 ( .A1(n12393), .A2(n12392), .ZN(n7246) );
  NAND2_X1 U8956 ( .A1(n12161), .A2(n12160), .ZN(n12273) );
  NAND2_X1 U8957 ( .A1(n11576), .A2(n11414), .ZN(n11559) );
  INV_X1 U8958 ( .A(n15063), .ZN(n15294) );
  NAND2_X1 U8959 ( .A1(n15093), .A2(n11203), .ZN(n15013) );
  NOR2_X1 U8960 ( .A1(n15067), .A2(n12785), .ZN(n15086) );
  INV_X1 U8961 ( .A(n15013), .ZN(n15285) );
  NAND2_X1 U8962 ( .A1(n6955), .A2(n6740), .ZN(n15211) );
  INV_X1 U8963 ( .A(n15122), .ZN(n6955) );
  INV_X2 U8964 ( .A(n15524), .ZN(n15526) );
  NAND2_X1 U8965 ( .A1(n6868), .A2(n6867), .ZN(n13093) );
  NAND2_X1 U8966 ( .A1(n7703), .A2(n7701), .ZN(n6867) );
  INV_X1 U8967 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n9815) );
  XNOR2_X1 U8968 ( .A(n8883), .B(n8882), .ZN(n15235) );
  INV_X1 U8969 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n15236) );
  CLKBUF_X1 U8970 ( .A(n10187), .Z(n14718) );
  INV_X1 U8971 ( .A(n9905), .ZN(n15242) );
  CLKBUF_X1 U8972 ( .A(n9901), .Z(n12387) );
  INV_X1 U8973 ( .A(n9795), .ZN(n9828) );
  NAND2_X1 U8974 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_19__SCAN_IN), 
        .ZN(n7063) );
  INV_X1 U8975 ( .A(n11260), .ZN(n7064) );
  INV_X1 U8976 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n10719) );
  INV_X1 U8977 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n10458) );
  INV_X1 U8978 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n10360) );
  INV_X1 U8979 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n10246) );
  INV_X1 U8980 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n10073) );
  INV_X1 U8981 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n10013) );
  INV_X1 U8982 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n10008) );
  OR2_X1 U8983 ( .A1(n10007), .A2(n10006), .ZN(n14782) );
  OR2_X1 U8984 ( .A1(n15800), .A2(n15801), .ZN(n7240) );
  XNOR2_X1 U8985 ( .A(n7819), .B(n7820), .ZN(n15790) );
  NAND2_X1 U8986 ( .A1(n15790), .A2(n15789), .ZN(n15788) );
  XNOR2_X1 U8987 ( .A(n7829), .B(P2_ADDR_REG_7__SCAN_IN), .ZN(n15793) );
  XNOR2_X1 U8988 ( .A(n7832), .B(n7831), .ZN(n15260) );
  OAI21_X1 U8989 ( .B1(n7134), .B2(n7131), .A(n7130), .ZN(n15422) );
  NAND2_X1 U8990 ( .A1(n15267), .A2(n7233), .ZN(n7130) );
  NOR2_X1 U8991 ( .A1(n15267), .A2(n7233), .ZN(n7131) );
  INV_X1 U8992 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n7233) );
  NAND2_X1 U8993 ( .A1(n15422), .A2(n15421), .ZN(n15420) );
  NOR2_X1 U8994 ( .A1(n7837), .A2(n6718), .ZN(n15425) );
  INV_X1 U8995 ( .A(n15425), .ZN(n15426) );
  NAND2_X1 U8996 ( .A1(n15427), .A2(n15567), .ZN(n15424) );
  OAI21_X1 U8997 ( .B1(n7838), .B2(P2_ADDR_REG_14__SCAN_IN), .A(n15432), .ZN(
        n15438) );
  NAND2_X1 U8998 ( .A1(n15438), .A2(n15437), .ZN(n15436) );
  NAND2_X1 U8999 ( .A1(n7125), .A2(n15436), .ZN(n15441) );
  OAI21_X1 U9000 ( .B1(n15438), .B2(n15437), .A(n7234), .ZN(n7125) );
  INV_X1 U9001 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n7234) );
  NAND2_X1 U9002 ( .A1(n15441), .A2(n15442), .ZN(n15440) );
  NAND2_X1 U9003 ( .A1(n7123), .A2(n15440), .ZN(n15298) );
  OAI21_X1 U9004 ( .B1(n15441), .B2(n15442), .A(n7124), .ZN(n7123) );
  INV_X1 U9005 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n7124) );
  NOR2_X1 U9006 ( .A1(n13527), .A2(n13528), .ZN(n6947) );
  NAND2_X1 U9007 ( .A1(n6928), .A2(n6820), .ZN(P3_U3488) );
  NAND2_X1 U9008 ( .A1(n15782), .A2(P3_REG1_REG_29__SCAN_IN), .ZN(n6927) );
  OR2_X1 U9009 ( .A1(n15784), .A2(P3_REG1_REG_28__SCAN_IN), .ZN(n6951) );
  INV_X1 U9010 ( .A(n6978), .ZN(n6977) );
  NAND2_X1 U9011 ( .A1(n6970), .A2(n6711), .ZN(P3_U3454) );
  NAND2_X1 U9012 ( .A1(n12853), .A2(n12852), .ZN(n12854) );
  NAND2_X1 U9013 ( .A1(n7571), .A2(n15345), .ZN(n7570) );
  NAND2_X1 U9014 ( .A1(n6854), .A2(n6853), .ZN(n6852) );
  INV_X1 U9015 ( .A(n6964), .ZN(n6963) );
  OAI21_X1 U9016 ( .B1(n14040), .B2(n14234), .A(n14039), .ZN(n6964) );
  NAND2_X1 U9017 ( .A1(n7438), .A2(n7167), .ZN(P2_U3528) );
  INV_X1 U9018 ( .A(n7168), .ZN(n7167) );
  OAI21_X1 U9019 ( .B1(n7442), .B2(n6671), .A(n7434), .ZN(n7438) );
  OAI21_X1 U9020 ( .B1(n14040), .B2(n14316), .A(n7437), .ZN(n7168) );
  INV_X1 U9021 ( .A(n6937), .ZN(n6936) );
  OAI21_X1 U9022 ( .B1(n14332), .B2(n14316), .A(n14252), .ZN(n6937) );
  INV_X1 U9023 ( .A(n6939), .ZN(n6938) );
  OAI21_X1 U9024 ( .B1(n14332), .B2(n14379), .A(n14330), .ZN(n6939) );
  XNOR2_X1 U9025 ( .A(n14524), .B(n14525), .ZN(n14531) );
  INV_X1 U9026 ( .A(n7230), .ZN(n15255) );
  NOR2_X1 U9027 ( .A1(n15262), .A2(n15263), .ZN(n15261) );
  NAND2_X1 U9028 ( .A1(n15266), .A2(n15267), .ZN(n15265) );
  INV_X1 U9029 ( .A(n7134), .ZN(n15266) );
  XNOR2_X1 U9030 ( .A(n7126), .B(P2_ADDR_REG_18__SCAN_IN), .ZN(SUB_1596_U62)
         );
  NAND2_X1 U9031 ( .A1(n7237), .A2(n7127), .ZN(n7126) );
  NAND2_X1 U9032 ( .A1(n15247), .A2(n15248), .ZN(n7127) );
  XNOR2_X1 U9033 ( .A(n7236), .B(n7235), .ZN(SUB_1596_U4) );
  XNOR2_X1 U9034 ( .A(n8178), .B(n6845), .ZN(n7235) );
  NAND2_X1 U9035 ( .A1(n7238), .A2(n7237), .ZN(n7236) );
  AND2_X1 U9036 ( .A1(n7161), .A2(n6759), .ZN(n6685) );
  AND2_X1 U9037 ( .A1(n12638), .A2(n12640), .ZN(n6686) );
  INV_X2 U9038 ( .A(P3_IR_REG_31__SCAN_IN), .ZN(n9682) );
  INV_X2 U9039 ( .A(n14445), .ZN(n9851) );
  INV_X1 U9040 ( .A(n6677), .ZN(n12451) );
  INV_X1 U9041 ( .A(n8755), .ZN(n7557) );
  AND2_X1 U9042 ( .A1(n9722), .A2(n6716), .ZN(n6688) );
  NAND2_X1 U9043 ( .A1(n8986), .A2(n7164), .ZN(n7166) );
  AND2_X1 U9044 ( .A1(n7152), .A2(n14229), .ZN(n6689) );
  NOR2_X1 U9045 ( .A1(n14198), .A2(n7538), .ZN(n6690) );
  AND2_X1 U9046 ( .A1(n10008), .A2(P1_DATAO_REG_6__SCAN_IN), .ZN(n6691) );
  AND2_X1 U9047 ( .A1(n14162), .A2(n8927), .ZN(n6692) );
  AND2_X1 U9048 ( .A1(n6788), .A2(n7240), .ZN(n6693) );
  NOR2_X1 U9049 ( .A1(n13151), .A2(n13091), .ZN(n6694) );
  OR2_X1 U9050 ( .A1(n13824), .A2(n9715), .ZN(n6695) );
  INV_X1 U9051 ( .A(n14041), .ZN(n7171) );
  OR2_X1 U9052 ( .A1(n12810), .A2(n7274), .ZN(n6696) );
  INV_X1 U9053 ( .A(n13615), .ZN(n7624) );
  NAND2_X1 U9054 ( .A1(n8774), .A2(n8773), .ZN(n14262) );
  AND2_X1 U9055 ( .A1(n7199), .A2(n14563), .ZN(n6697) );
  NOR2_X1 U9056 ( .A1(n7644), .A2(n7639), .ZN(n6698) );
  AND2_X1 U9057 ( .A1(n7572), .A2(n7575), .ZN(n6699) );
  AND2_X1 U9058 ( .A1(n12616), .A2(n12610), .ZN(n6700) );
  AND2_X1 U9059 ( .A1(n6665), .A2(n13158), .ZN(n6701) );
  AND2_X1 U9060 ( .A1(n12728), .A2(n7070), .ZN(n6702) );
  INV_X1 U9061 ( .A(n7163), .ZN(n7159) );
  NAND2_X1 U9062 ( .A1(n6728), .A2(n8984), .ZN(n7163) );
  AND2_X1 U9063 ( .A1(n9300), .A2(n12038), .ZN(n6703) );
  AND2_X1 U9064 ( .A1(n14158), .A2(n7144), .ZN(n6704) );
  INV_X1 U9065 ( .A(P3_IR_REG_28__SCAN_IN), .ZN(n9025) );
  MUX2_X1 U9066 ( .A(n14702), .B(n12637), .S(n12789), .Z(n12639) );
  AND2_X1 U9067 ( .A1(n11822), .A2(n12805), .ZN(n6705) );
  OR2_X1 U9068 ( .A1(n9673), .A2(n10594), .ZN(n6706) );
  XNOR2_X1 U9069 ( .A(n13212), .B(n13580), .ZN(n13297) );
  AND2_X1 U9070 ( .A1(n7143), .A2(n7142), .ZN(n6707) );
  NAND2_X1 U9071 ( .A1(n12967), .A2(n13976), .ZN(n6708) );
  OR2_X1 U9072 ( .A1(n14295), .A2(n13914), .ZN(n6709) );
  OR2_X1 U9073 ( .A1(n7560), .A2(n7562), .ZN(n6710) );
  AND2_X1 U9074 ( .A1(n6988), .A2(n6828), .ZN(n6711) );
  INV_X1 U9075 ( .A(n13141), .ZN(n6966) );
  NAND2_X1 U9076 ( .A1(n12060), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n6712) );
  NAND2_X1 U9077 ( .A1(n12860), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n6713) );
  INV_X2 U9078 ( .A(n15773), .ZN(n15775) );
  NOR2_X1 U9079 ( .A1(n7676), .A2(n7673), .ZN(n6714) );
  AND2_X1 U9080 ( .A1(n8300), .A2(SI_24_), .ZN(n6715) );
  INV_X1 U9081 ( .A(n13935), .ZN(n15345) );
  CLKBUF_X3 U9082 ( .A(n8336), .Z(n8941) );
  NAND2_X2 U9083 ( .A1(n8381), .A2(n8253), .ZN(n8379) );
  NAND2_X1 U9084 ( .A1(n13793), .A2(n13580), .ZN(n6716) );
  AND2_X1 U9085 ( .A1(n6998), .A2(n7391), .ZN(n6717) );
  AND2_X1 U9086 ( .A1(n7231), .A2(n15420), .ZN(n6718) );
  AND2_X1 U9087 ( .A1(n9080), .A2(n9003), .ZN(n9102) );
  AND2_X1 U9088 ( .A1(n14569), .A2(n14470), .ZN(n6719) );
  AND2_X1 U9089 ( .A1(n6695), .A2(n9713), .ZN(n6720) );
  NAND2_X1 U9090 ( .A1(n12141), .A2(n12145), .ZN(n6721) );
  INV_X1 U9091 ( .A(n9636), .ZN(n13641) );
  AND2_X1 U9092 ( .A1(n9639), .A2(n9638), .ZN(n9636) );
  AND2_X1 U9093 ( .A1(n14516), .A2(n12500), .ZN(n6722) );
  AND2_X1 U9094 ( .A1(n13010), .A2(n13009), .ZN(n6723) );
  OAI21_X1 U9095 ( .B1(n8702), .B2(n7049), .A(n7047), .ZN(n13926) );
  NOR2_X1 U9096 ( .A1(n15286), .A2(n14697), .ZN(n6724) );
  NOR2_X1 U9097 ( .A1(n15154), .A2(n14693), .ZN(n6725) );
  INV_X1 U9098 ( .A(n12240), .ZN(n6944) );
  AND2_X1 U9099 ( .A1(n7046), .A2(n7050), .ZN(n6726) );
  INV_X1 U9100 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n15227) );
  INV_X1 U9101 ( .A(n13145), .ZN(n6986) );
  INV_X1 U9102 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n14381) );
  XNOR2_X1 U9103 ( .A(n8754), .B(n8755), .ZN(n13852) );
  NAND2_X1 U9104 ( .A1(n14351), .A2(n13967), .ZN(n6727) );
  OR2_X1 U9105 ( .A1(n14295), .A2(n13970), .ZN(n6728) );
  AND2_X1 U9106 ( .A1(n7351), .A2(n12272), .ZN(n6729) );
  XOR2_X1 U9107 ( .A(n14351), .B(n8382), .Z(n6730) );
  NAND2_X1 U9108 ( .A1(n6942), .A2(n10595), .ZN(n10829) );
  OR2_X1 U9109 ( .A1(n10986), .A2(n10985), .ZN(n6731) );
  INV_X1 U9110 ( .A(n13689), .ZN(n7639) );
  INV_X1 U9111 ( .A(n12266), .ZN(n7647) );
  NAND2_X1 U9112 ( .A1(n12493), .A2(n12492), .ZN(n14516) );
  NAND2_X1 U9113 ( .A1(n12513), .A2(n12512), .ZN(n15113) );
  INV_X1 U9114 ( .A(n15113), .ZN(n14563) );
  AND4_X1 U9115 ( .A1(n11850), .A2(n11852), .A3(n11604), .A4(n11603), .ZN(
        n6732) );
  AND2_X1 U9116 ( .A1(n12428), .A2(n12427), .ZN(n15166) );
  INV_X1 U9117 ( .A(n15166), .ZN(n14977) );
  INV_X1 U9118 ( .A(n14888), .ZN(n7267) );
  AND2_X1 U9119 ( .A1(n9673), .A2(n15715), .ZN(n6733) );
  AND2_X1 U9120 ( .A1(n14343), .A2(n8930), .ZN(n6734) );
  NAND2_X1 U9121 ( .A1(n15014), .A2(n14988), .ZN(n6735) );
  AND2_X1 U9122 ( .A1(n9813), .A2(n9831), .ZN(n6736) );
  OR2_X1 U9123 ( .A1(n15158), .A2(n14941), .ZN(n6737) );
  INV_X1 U9124 ( .A(n12636), .ZN(n7060) );
  INV_X1 U9125 ( .A(n14859), .ZN(n14857) );
  XNOR2_X1 U9126 ( .A(n14866), .B(n14688), .ZN(n14859) );
  OR2_X1 U9127 ( .A1(n10802), .A2(n10803), .ZN(n6738) );
  AND2_X1 U9128 ( .A1(n13186), .A2(n13706), .ZN(n6739) );
  NAND2_X1 U9129 ( .A1(n8898), .A2(n8897), .ZN(n13126) );
  MUX2_X1 U9130 ( .A(n14704), .B(n12629), .S(n12789), .Z(n12631) );
  MUX2_X1 U9131 ( .A(n14692), .B(n15148), .S(n12789), .Z(n12730) );
  AND2_X1 U9132 ( .A1(n14865), .A2(n14864), .ZN(n6740) );
  INV_X1 U9133 ( .A(n14525), .ZN(n7375) );
  INV_X1 U9134 ( .A(n10986), .ZN(n7510) );
  AND2_X1 U9135 ( .A1(n15133), .A2(n14690), .ZN(n6741) );
  AND2_X1 U9136 ( .A1(n7324), .A2(n9099), .ZN(n6742) );
  AND2_X1 U9137 ( .A1(n12937), .A2(n12931), .ZN(n6743) );
  AND2_X1 U9138 ( .A1(n15243), .A2(n12448), .ZN(n15154) );
  NAND2_X1 U9139 ( .A1(n9885), .A2(n9886), .ZN(n9840) );
  AND2_X1 U9140 ( .A1(n13202), .A2(n13638), .ZN(n6744) );
  AND2_X1 U9141 ( .A1(n14125), .A2(n6727), .ZN(n6745) );
  INV_X1 U9142 ( .A(n12863), .ZN(n15616) );
  AND2_X1 U9143 ( .A1(n14285), .A2(n13916), .ZN(n6746) );
  AND2_X1 U9144 ( .A1(n6932), .A2(n7743), .ZN(n6747) );
  AND2_X1 U9145 ( .A1(n12946), .A2(n12945), .ZN(n6748) );
  AND2_X1 U9146 ( .A1(n13217), .A2(n13548), .ZN(n6749) );
  NOR2_X1 U9147 ( .A1(n13486), .A2(n13487), .ZN(n6750) );
  NOR2_X1 U9148 ( .A1(n13435), .A2(n13436), .ZN(n6751) );
  NAND2_X1 U9149 ( .A1(n12348), .A2(n12347), .ZN(n15196) );
  INV_X1 U9150 ( .A(n13338), .ZN(n9723) );
  NAND2_X1 U9151 ( .A1(n9424), .A2(n9423), .ZN(n13338) );
  NOR2_X1 U9152 ( .A1(n11307), .A2(n7040), .ZN(n6752) );
  INV_X1 U9153 ( .A(n15286), .ZN(n12359) );
  NAND2_X1 U9154 ( .A1(n12330), .A2(n12329), .ZN(n15286) );
  OR2_X1 U9155 ( .A1(n12962), .A2(n12964), .ZN(n6753) );
  OR2_X1 U9156 ( .A1(n12950), .A2(n6748), .ZN(n6754) );
  INV_X1 U9157 ( .A(n7532), .ZN(n7176) );
  NAND2_X1 U9158 ( .A1(n14256), .A2(n13963), .ZN(n7532) );
  AND2_X1 U9159 ( .A1(n14857), .A2(n12549), .ZN(n6755) );
  AND2_X1 U9160 ( .A1(n7061), .A2(n12636), .ZN(n6756) );
  INV_X1 U9161 ( .A(n11414), .ZN(n7347) );
  AND2_X1 U9162 ( .A1(n7563), .A2(n7561), .ZN(n6757) );
  INV_X1 U9163 ( .A(n12728), .ZN(n7069) );
  AND2_X1 U9164 ( .A1(n9158), .A2(n7633), .ZN(n6758) );
  NAND2_X1 U9165 ( .A1(n14289), .A2(n13969), .ZN(n6759) );
  AND2_X1 U9166 ( .A1(n12940), .A2(n8907), .ZN(n6760) );
  NAND2_X1 U9167 ( .A1(n13699), .A2(n13707), .ZN(n6761) );
  INV_X1 U9168 ( .A(n7248), .ZN(n7247) );
  OAI21_X1 U9169 ( .B1(n12392), .B2(n7249), .A(n12398), .ZN(n7248) );
  AND2_X1 U9170 ( .A1(n12551), .A2(n12550), .ZN(n6762) );
  AND2_X1 U9171 ( .A1(n10946), .A2(n7281), .ZN(n6763) );
  INV_X1 U9172 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n7030) );
  INV_X1 U9173 ( .A(n7274), .ZN(n7273) );
  AND2_X1 U9174 ( .A1(n7659), .A2(n9012), .ZN(n6764) );
  AND2_X1 U9175 ( .A1(n7518), .A2(n7517), .ZN(n6765) );
  MUX2_X1 U9176 ( .A(n14969), .B(n15158), .S(n12789), .Z(n12724) );
  NOR2_X1 U9177 ( .A1(n12655), .A2(n12657), .ZN(n6766) );
  OR2_X1 U9178 ( .A1(n13046), .A2(n7613), .ZN(n6767) );
  NOR2_X1 U9179 ( .A1(n13985), .A2(n15659), .ZN(n6768) );
  NOR2_X1 U9180 ( .A1(n14289), .A2(n13969), .ZN(n6769) );
  INV_X1 U9181 ( .A(n7029), .ZN(n7028) );
  NAND2_X1 U9182 ( .A1(n8582), .A2(n11699), .ZN(n7029) );
  AND2_X1 U9183 ( .A1(n15154), .A2(n14573), .ZN(n6770) );
  AND2_X1 U9184 ( .A1(n9623), .A2(n9628), .ZN(n13662) );
  INV_X1 U9185 ( .A(n13662), .ZN(n7651) );
  INV_X1 U9186 ( .A(n7575), .ZN(n7574) );
  OR2_X1 U9187 ( .A1(n8805), .A2(n8826), .ZN(n7575) );
  AND2_X1 U9188 ( .A1(n13014), .A2(n13013), .ZN(n6771) );
  NAND2_X1 U9189 ( .A1(n7595), .A2(n13092), .ZN(n6772) );
  AND2_X1 U9190 ( .A1(n13581), .A2(n13333), .ZN(n6773) );
  NAND2_X1 U9191 ( .A1(n14247), .A2(n13961), .ZN(n6774) );
  AND2_X1 U9192 ( .A1(n8257), .A2(SI_8_), .ZN(n6775) );
  AND2_X1 U9193 ( .A1(n9172), .A2(n9582), .ZN(n6776) );
  NAND2_X1 U9194 ( .A1(n13141), .A2(n8980), .ZN(n6777) );
  AND2_X1 U9195 ( .A1(n13196), .A2(n7656), .ZN(n6778) );
  INV_X1 U9196 ( .A(n7305), .ZN(n7304) );
  NAND2_X1 U9197 ( .A1(n13201), .A2(n13200), .ZN(n7305) );
  XNOR2_X1 U9198 ( .A(n13207), .B(n10830), .ZN(n11007) );
  AND2_X1 U9199 ( .A1(n9026), .A2(n9682), .ZN(n6779) );
  INV_X1 U9200 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n9796) );
  NOR2_X1 U9201 ( .A1(n7708), .A2(n12656), .ZN(n7707) );
  OR2_X1 U9202 ( .A1(n10864), .A2(n10869), .ZN(n6780) );
  AND2_X1 U9203 ( .A1(n12729), .A2(n12731), .ZN(n6781) );
  NOR2_X1 U9204 ( .A1(n14068), .A2(n8990), .ZN(n6782) );
  NAND2_X1 U9205 ( .A1(n7638), .A2(n6761), .ZN(n6783) );
  INV_X1 U9206 ( .A(n7543), .ZN(n7542) );
  NAND2_X1 U9207 ( .A1(n13142), .A2(n8979), .ZN(n7543) );
  OR2_X1 U9208 ( .A1(n7560), .A2(n8755), .ZN(n6784) );
  INV_X1 U9209 ( .A(n12729), .ZN(n7706) );
  INV_X1 U9210 ( .A(n12630), .ZN(n7710) );
  INV_X1 U9211 ( .A(n9688), .ZN(n13517) );
  OR2_X1 U9212 ( .A1(n12920), .A2(n12921), .ZN(n6785) );
  INV_X1 U9213 ( .A(n9975), .ZN(n7202) );
  OR2_X1 U9214 ( .A1(n13388), .A2(n13387), .ZN(n6786) );
  OR2_X1 U9215 ( .A1(n7825), .A2(n7822), .ZN(n6787) );
  MUX2_X1 U9216 ( .A(n14700), .B(n12650), .S(n12789), .Z(n12653) );
  INV_X1 U9217 ( .A(n12653), .ZN(n7085) );
  OR2_X1 U9218 ( .A1(n7812), .A2(n7809), .ZN(n6788) );
  AOI21_X1 U9219 ( .B1(n14386), .B2(n11026), .A(n12571), .ZN(n12759) );
  OR2_X1 U9220 ( .A1(n13109), .A2(n13110), .ZN(n6789) );
  AND2_X1 U9221 ( .A1(n12241), .A2(n6944), .ZN(n6790) );
  AND2_X1 U9222 ( .A1(n12937), .A2(n12927), .ZN(n6791) );
  AND2_X1 U9223 ( .A1(n13251), .A2(n13565), .ZN(n6792) );
  NOR2_X1 U9224 ( .A1(n14107), .A2(n7537), .ZN(n6793) );
  AND2_X1 U9225 ( .A1(n7189), .A2(n7188), .ZN(n6794) );
  AND2_X1 U9226 ( .A1(n10836), .A2(n10674), .ZN(n6795) );
  AND2_X1 U9227 ( .A1(n7745), .A2(n7597), .ZN(n6796) );
  AND2_X1 U9228 ( .A1(n12616), .A2(n12614), .ZN(n6797) );
  AND2_X1 U9229 ( .A1(n14999), .A2(n12424), .ZN(n6798) );
  AND2_X1 U9230 ( .A1(n7617), .A2(n8196), .ZN(n6799) );
  NAND2_X1 U9231 ( .A1(n8745), .A2(n8744), .ZN(n14274) );
  OR2_X1 U9232 ( .A1(n13025), .A2(n13026), .ZN(n6800) );
  OR2_X1 U9233 ( .A1(n12640), .A2(n12638), .ZN(n6801) );
  AND2_X1 U9234 ( .A1(n12617), .A2(n12618), .ZN(n12616) );
  AND2_X1 U9235 ( .A1(n12903), .A2(n12902), .ZN(n6802) );
  NAND2_X1 U9236 ( .A1(n12089), .A2(n12090), .ZN(n6803) );
  INV_X1 U9237 ( .A(n7478), .ZN(n7477) );
  NOR2_X1 U9238 ( .A1(n9337), .A2(n7479), .ZN(n7478) );
  AND2_X1 U9239 ( .A1(n7715), .A2(n7079), .ZN(n6804) );
  OR2_X1 U9240 ( .A1(n7583), .A2(n7584), .ZN(n6805) );
  NAND2_X1 U9241 ( .A1(n9682), .A2(n9012), .ZN(n6806) );
  INV_X1 U9242 ( .A(P3_IR_REG_27__SCAN_IN), .ZN(n9026) );
  INV_X1 U9243 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n9817) );
  OR2_X1 U9244 ( .A1(n7604), .A2(n7603), .ZN(n6807) );
  AND2_X1 U9245 ( .A1(n6784), .A2(n7556), .ZN(n6808) );
  AND2_X1 U9246 ( .A1(n9538), .A2(n9537), .ZN(n13627) );
  AND2_X1 U9247 ( .A1(n14295), .A2(n13914), .ZN(n6809) );
  OR2_X1 U9248 ( .A1(n7375), .A2(n7373), .ZN(n6810) );
  NAND2_X1 U9249 ( .A1(n9508), .A2(n15305), .ZN(n6811) );
  INV_X2 U9250 ( .A(n15733), .ZN(n15735) );
  AND2_X1 U9251 ( .A1(n14226), .A2(n8859), .ZN(n14160) );
  XNOR2_X1 U9252 ( .A(n7287), .B(n9327), .ZN(n9671) );
  OAI21_X1 U9253 ( .B1(n12382), .B2(n12378), .A(n12379), .ZN(n13183) );
  NOR2_X1 U9254 ( .A1(n12362), .A2(n12350), .ZN(n6812) );
  NOR2_X1 U9255 ( .A1(n12286), .A2(n12285), .ZN(n7272) );
  OR2_X1 U9256 ( .A1(n7272), .A2(n6696), .ZN(n12325) );
  NAND2_X1 U9257 ( .A1(n7581), .A2(n12255), .ZN(n13887) );
  NAND2_X1 U9258 ( .A1(n8641), .A2(n8643), .ZN(n8645) );
  NAND2_X1 U9259 ( .A1(n7454), .A2(n9080), .ZN(n9223) );
  INV_X1 U9260 ( .A(n13964), .ZN(n7536) );
  AND4_X1 U9261 ( .A1(n9321), .A2(n9320), .A3(n9319), .A4(n9318), .ZN(n13681)
         );
  OR2_X1 U9262 ( .A1(n8290), .A2(n8292), .ZN(n6813) );
  INV_X1 U9263 ( .A(n13710), .ZN(n7645) );
  AND2_X1 U9264 ( .A1(n14152), .A2(n6704), .ZN(n6814) );
  AND2_X1 U9265 ( .A1(n12360), .A2(n7191), .ZN(n6815) );
  AND2_X1 U9266 ( .A1(n12109), .A2(n7152), .ZN(n6816) );
  OR2_X1 U9267 ( .A1(n9259), .A2(P3_IR_REG_14__SCAN_IN), .ZN(n6817) );
  INV_X1 U9268 ( .A(n7322), .ZN(n7321) );
  OAI21_X1 U9269 ( .B1(n9255), .B2(n7323), .A(n9272), .ZN(n7322) );
  NAND2_X1 U9270 ( .A1(n7289), .A2(n13185), .ZN(n13224) );
  NAND2_X1 U9271 ( .A1(n7246), .A2(n12681), .ZN(n15039) );
  XNOR2_X1 U9272 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(P2_DATAO_REG_5__SCAN_IN), 
        .ZN(n9114) );
  INV_X1 U9273 ( .A(n9114), .ZN(n7096) );
  INV_X1 U9274 ( .A(n14343), .ZN(n7142) );
  INV_X1 U9275 ( .A(P3_IR_REG_14__SCAN_IN), .ZN(n7307) );
  INV_X1 U9276 ( .A(n13556), .ZN(n13782) );
  NAND2_X1 U9277 ( .A1(n9437), .A2(n9436), .ZN(n13556) );
  NAND2_X1 U9278 ( .A1(n8570), .A2(n8569), .ZN(n12967) );
  NAND2_X1 U9279 ( .A1(n8735), .A2(n8734), .ZN(n14351) );
  INV_X1 U9280 ( .A(n14351), .ZN(n7144) );
  INV_X1 U9281 ( .A(n15148), .ZN(n7193) );
  INV_X1 U9282 ( .A(n9593), .ZN(n7473) );
  NOR2_X1 U9283 ( .A1(n12110), .A2(n12988), .ZN(n12109) );
  AND2_X1 U9284 ( .A1(n11914), .A2(P3_REG1_REG_10__SCAN_IN), .ZN(n7520) );
  INV_X1 U9285 ( .A(n7520), .ZN(n7517) );
  OAI21_X1 U9286 ( .B1(n12286), .B2(n7268), .A(n7270), .ZN(n15277) );
  OR2_X1 U9287 ( .A1(n13277), .A2(n13680), .ZN(n6818) );
  NAND2_X1 U9288 ( .A1(n14986), .A2(n7196), .ZN(n7197) );
  AND2_X1 U9289 ( .A1(n6818), .A2(n13190), .ZN(n6819) );
  AND2_X1 U9290 ( .A1(n7726), .A2(n6927), .ZN(n6820) );
  AND2_X1 U9291 ( .A1(n12102), .A2(n8916), .ZN(n6821) );
  AND2_X1 U9292 ( .A1(n13305), .A2(n7304), .ZN(n6822) );
  OR2_X1 U9293 ( .A1(n9826), .A2(n7384), .ZN(n6823) );
  NOR2_X1 U9294 ( .A1(n8623), .A2(P2_IR_REG_16__SCAN_IN), .ZN(n8641) );
  AND2_X1 U9295 ( .A1(n10719), .A2(P1_DATAO_REG_15__SCAN_IN), .ZN(n6824) );
  INV_X1 U9296 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n6925) );
  NOR2_X1 U9297 ( .A1(n7667), .A2(n8808), .ZN(n7666) );
  INV_X1 U9298 ( .A(n13298), .ZN(n13613) );
  INV_X1 U9299 ( .A(n12222), .ZN(n6901) );
  INV_X1 U9300 ( .A(P3_IR_REG_25__SCAN_IN), .ZN(n9012) );
  AND2_X2 U9301 ( .A1(n8997), .A2(n8953), .ZN(n15688) );
  NAND2_X1 U9302 ( .A1(n9671), .A2(n10926), .ZN(n10594) );
  NAND2_X1 U9303 ( .A1(n8664), .A2(n8663), .ZN(n14210) );
  INV_X1 U9304 ( .A(n14210), .ZN(n7151) );
  INV_X1 U9305 ( .A(n12048), .ZN(n7627) );
  AND2_X1 U9306 ( .A1(n9368), .A2(n6713), .ZN(n6825) );
  INV_X2 U9307 ( .A(n15534), .ZN(n15537) );
  NAND2_X1 U9308 ( .A1(n6874), .A2(n12356), .ZN(n15287) );
  NAND2_X1 U9309 ( .A1(n15341), .A2(n8540), .ZN(n11698) );
  INV_X1 U9310 ( .A(n13895), .ZN(n7045) );
  AND2_X1 U9311 ( .A1(n13377), .A2(P3_REG2_REG_12__SCAN_IN), .ZN(n6826) );
  NAND2_X1 U9312 ( .A1(n7039), .A2(n7037), .ZN(n15341) );
  AND2_X1 U9313 ( .A1(n12068), .A2(n7392), .ZN(n6827) );
  NOR2_X1 U9314 ( .A1(n12280), .A2(n12658), .ZN(n12360) );
  OR2_X1 U9315 ( .A1(n15775), .A2(n6969), .ZN(n6828) );
  INV_X1 U9316 ( .A(n8788), .ZN(n7674) );
  OR2_X1 U9317 ( .A1(n10533), .A2(n7017), .ZN(n6829) );
  OR2_X1 U9318 ( .A1(n9382), .A2(n7328), .ZN(n6830) );
  AND2_X1 U9319 ( .A1(n8807), .A2(SI_27_), .ZN(n6831) );
  INV_X1 U9320 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n10656) );
  NAND2_X1 U9321 ( .A1(n7327), .A2(n7111), .ZN(n7110) );
  OR2_X1 U9322 ( .A1(P3_REG0_REG_28__SCAN_IN), .A2(n15775), .ZN(n6832) );
  NOR2_X1 U9323 ( .A1(n13399), .A2(n13398), .ZN(n6833) );
  AND2_X1 U9324 ( .A1(n6825), .A2(n6712), .ZN(n6834) );
  AND2_X1 U9325 ( .A1(n7679), .A2(n8757), .ZN(n6835) );
  OR2_X1 U9326 ( .A1(n8860), .A2(n13122), .ZN(n8753) );
  INV_X1 U9327 ( .A(n8753), .ZN(n14206) );
  NAND2_X1 U9328 ( .A1(n6889), .A2(n6887), .ZN(n9689) );
  INV_X1 U9329 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n7339) );
  AND2_X2 U9330 ( .A1(n10933), .A2(n9776), .ZN(n15784) );
  AND2_X2 U9331 ( .A1(n8997), .A2(n11064), .ZN(n15680) );
  INV_X1 U9332 ( .A(n15680), .ZN(n15678) );
  INV_X1 U9333 ( .A(n10437), .ZN(n6922) );
  NAND2_X1 U9334 ( .A1(n7618), .A2(n9694), .ZN(n11052) );
  AND2_X1 U9335 ( .A1(n15698), .A2(P3_ADDR_REG_19__SCAN_IN), .ZN(n6836) );
  XOR2_X1 U9336 ( .A(n8389), .B(n8390), .Z(n6837) );
  INV_X1 U9337 ( .A(n9512), .ZN(n10604) );
  INV_X1 U9338 ( .A(n12641), .ZN(n7186) );
  NAND2_X1 U9339 ( .A1(n8876), .A2(n8863), .ZN(n13935) );
  AND2_X1 U9340 ( .A1(n13525), .A2(n13523), .ZN(n6838) );
  NAND2_X1 U9341 ( .A1(n7525), .A2(n7523), .ZN(n6839) );
  AND2_X1 U9342 ( .A1(P2_DATAO_REG_28__SCAN_IN), .A2(n14392), .ZN(n6840) );
  INV_X1 U9343 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n15240) );
  INV_X1 U9344 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n12567) );
  OR2_X1 U9345 ( .A1(P2_DATAO_REG_26__SCAN_IN), .A2(n14394), .ZN(n6841) );
  AND2_X1 U9346 ( .A1(n6885), .A2(n6884), .ZN(n6842) );
  AND2_X1 U9347 ( .A1(n13471), .A2(n6839), .ZN(n6843) );
  INV_X1 U9348 ( .A(SI_26_), .ZN(n13849) );
  AND2_X1 U9349 ( .A1(n10845), .A2(n10770), .ZN(n6844) );
  INV_X1 U9350 ( .A(P3_ADDR_REG_4__SCAN_IN), .ZN(n7138) );
  INV_X1 U9351 ( .A(n8321), .ZN(n13158) );
  NAND2_X1 U9352 ( .A1(n9814), .A2(n7721), .ZN(n7722) );
  INV_X1 U9353 ( .A(n14710), .ZN(n7341) );
  XOR2_X1 U9354 ( .A(n7840), .B(P1_ADDR_REG_19__SCAN_IN), .Z(n6845) );
  INV_X1 U9355 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n7107) );
  INV_X1 U9356 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n7748) );
  INV_X1 U9357 ( .A(P1_RD_REG_SCAN_IN), .ZN(n7140) );
  NAND2_X1 U9358 ( .A1(n10911), .A2(n10912), .ZN(n10910) );
  INV_X1 U9359 ( .A(n13987), .ZN(n10384) );
  NAND2_X1 U9360 ( .A1(n12215), .A2(n8920), .ZN(n14218) );
  NAND2_X1 U9361 ( .A1(n7442), .A2(n15617), .ZN(n7441) );
  AND2_X1 U9362 ( .A1(n9928), .A2(n10024), .ZN(n10182) );
  NOR2_X1 U9363 ( .A1(n14021), .A2(n6670), .ZN(n14238) );
  OR2_X1 U9364 ( .A1(n14031), .A2(n6670), .ZN(n7145) );
  OR2_X1 U9365 ( .A1(n14247), .A2(n6670), .ZN(n7146) );
  AND2_X2 U9366 ( .A1(n11129), .A2(n15621), .ZN(n15627) );
  NAND3_X1 U9367 ( .A1(n6850), .A2(n6849), .A3(n8260), .ZN(n8506) );
  NAND3_X1 U9368 ( .A1(n8455), .A2(n8258), .A3(n7685), .ZN(n6850) );
  NAND2_X1 U9369 ( .A1(n6851), .A2(n7683), .ZN(n8489) );
  NAND2_X1 U9370 ( .A1(n8455), .A2(n7685), .ZN(n6851) );
  NAND2_X1 U9371 ( .A1(n6852), .A2(n13170), .ZN(P2_U3328) );
  NAND3_X1 U9372 ( .A1(n6857), .A2(n6856), .A3(n6855), .ZN(n6854) );
  NAND2_X1 U9373 ( .A1(n13165), .A2(n13163), .ZN(n6855) );
  OAI21_X1 U9374 ( .B1(n13165), .B2(n15620), .A(n6701), .ZN(n6857) );
  INV_X1 U9375 ( .A(n13111), .ZN(n6860) );
  NAND2_X1 U9376 ( .A1(n6861), .A2(n7203), .ZN(n6862) );
  NAND2_X1 U9377 ( .A1(n8357), .A2(n8356), .ZN(n6863) );
  NAND2_X1 U9378 ( .A1(n6863), .A2(n8241), .ZN(n8378) );
  NAND3_X1 U9379 ( .A1(n7421), .A2(P2_DATAO_REG_1__SCAN_IN), .A3(n7420), .ZN(
        n6864) );
  NAND2_X1 U9380 ( .A1(n12563), .A2(n12562), .ZN(n6868) );
  INV_X1 U9381 ( .A(n6870), .ZN(n10887) );
  NOR2_X4 U9382 ( .A1(P3_IR_REG_0__SCAN_IN), .A2(P3_IR_REG_1__SCAN_IN), .ZN(
        n9031) );
  INV_X1 U9383 ( .A(n10870), .ZN(n6872) );
  NAND2_X1 U9384 ( .A1(n6873), .A2(n6997), .ZN(n6996) );
  NAND4_X1 U9385 ( .A1(n10456), .A2(n10453), .A3(n10239), .A4(n10240), .ZN(
        n9791) );
  NAND2_X1 U9386 ( .A1(n7350), .A2(n7348), .ZN(n12355) );
  MUX2_X1 U9387 ( .A(n6875), .B(P1_REG1_REG_29__SCAN_IN), .S(n15534), .Z(
        P1_U3557) );
  MUX2_X1 U9388 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n6875), .S(n15526), .Z(
        P1_U3525) );
  OAI21_X1 U9389 ( .B1(n15110), .B2(n15482), .A(n6747), .ZN(n6875) );
  NAND2_X2 U9390 ( .A1(n15038), .A2(n12535), .ZN(n12537) );
  NAND2_X2 U9391 ( .A1(n12534), .A2(n12533), .ZN(n15038) );
  NAND2_X2 U9392 ( .A1(n6877), .A2(n12543), .ZN(n15163) );
  NAND2_X1 U9393 ( .A1(n12542), .A2(n12541), .ZN(n14978) );
  NAND2_X1 U9394 ( .A1(n6878), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n9866) );
  NAND2_X1 U9395 ( .A1(n13207), .A2(n15720), .ZN(n6883) );
  NAND2_X1 U9396 ( .A1(n6958), .A2(n6957), .ZN(n6885) );
  INV_X1 U9397 ( .A(n9011), .ZN(n6886) );
  NAND2_X2 U9398 ( .A1(n7450), .A2(n7454), .ZN(n9259) );
  AND3_X2 U9399 ( .A1(n7450), .A2(n7454), .A3(n6886), .ZN(n9683) );
  AND2_X1 U9400 ( .A1(n6902), .A2(n12222), .ZN(n6900) );
  NAND3_X1 U9401 ( .A1(n13235), .A2(n13297), .A3(n13613), .ZN(n6904) );
  NAND2_X1 U9402 ( .A1(n6905), .A2(n13211), .ZN(n13296) );
  NAND2_X1 U9403 ( .A1(n13235), .A2(n13613), .ZN(n6905) );
  INV_X1 U9404 ( .A(n13297), .ZN(n6906) );
  INV_X1 U9405 ( .A(n7290), .ZN(n6910) );
  INV_X1 U9406 ( .A(n7288), .ZN(n6911) );
  NAND2_X1 U9407 ( .A1(n6918), .A2(n6917), .ZN(n6919) );
  INV_X1 U9408 ( .A(n11298), .ZN(n6915) );
  NAND2_X1 U9409 ( .A1(n6919), .A2(n6732), .ZN(n6916) );
  NAND2_X1 U9410 ( .A1(n6916), .A2(n11611), .ZN(n11613) );
  INV_X1 U9411 ( .A(n6918), .ZN(n11300) );
  INV_X1 U9412 ( .A(n11613), .ZN(n6975) );
  INV_X1 U9413 ( .A(n6919), .ZN(n11612) );
  XNOR2_X1 U9414 ( .A(n15714), .B(n13207), .ZN(n6958) );
  OAI21_X1 U9415 ( .B1(n11237), .B2(n11236), .A(n11235), .ZN(n11242) );
  NOR2_X2 U9416 ( .A1(n6717), .A2(n12245), .ZN(n15391) );
  XNOR2_X1 U9417 ( .A(n9738), .B(n9739), .ZN(n13178) );
  XNOR2_X1 U9418 ( .A(n9798), .B(n9797), .ZN(n9901) );
  NAND2_X1 U9420 ( .A1(n9498), .A2(n9497), .ZN(n7314) );
  NAND2_X1 U9421 ( .A1(n9784), .A2(n15784), .ZN(n6928) );
  NAND2_X1 U9422 ( .A1(n9322), .A2(n9323), .ZN(n9325) );
  NAND2_X1 U9423 ( .A1(n7115), .A2(n6841), .ZN(n7114) );
  INV_X1 U9424 ( .A(n10715), .ZN(n7403) );
  OAI21_X1 U9425 ( .B1(P2_DATAO_REG_12__SCAN_IN), .B2(n10352), .A(n9230), .ZN(
        n9243) );
  NAND2_X1 U9426 ( .A1(n9146), .A2(n9145), .ZN(n9160) );
  NAND2_X1 U9427 ( .A1(n9202), .A2(n9201), .ZN(n9217) );
  NAND3_X1 U9428 ( .A1(n7395), .A2(n6943), .A3(n7400), .ZN(n11237) );
  NOR2_X1 U9429 ( .A1(n15388), .A2(n12311), .ZN(n12314) );
  AOI21_X2 U9430 ( .B1(n11145), .B2(n11144), .A(n6760), .ZN(n7725) );
  NAND2_X1 U9431 ( .A1(n15109), .A2(n15280), .ZN(n6932) );
  INV_X1 U9432 ( .A(n12818), .ZN(n7266) );
  XNOR2_X1 U9433 ( .A(n14081), .B(n14080), .ZN(n6934) );
  OAI21_X2 U9434 ( .B1(n12102), .B2(n7445), .A(n7443), .ZN(n12215) );
  NAND2_X1 U9435 ( .A1(n10479), .A2(n13123), .ZN(n10478) );
  NAND2_X1 U9436 ( .A1(n11516), .A2(n11515), .ZN(n11518) );
  XNOR2_X1 U9437 ( .A(n8239), .B(SI_2_), .ZN(n8357) );
  INV_X1 U9438 ( .A(n8217), .ZN(n8218) );
  NAND2_X1 U9439 ( .A1(n8913), .A2(n7422), .ZN(n11807) );
  NAND2_X1 U9440 ( .A1(n11621), .A2(n8911), .ZN(n11708) );
  NOR2_X2 U9441 ( .A1(n14256), .A2(n14091), .ZN(n14074) );
  OAI21_X1 U9442 ( .B1(n14248), .B2(n15656), .A(n6992), .ZN(n6991) );
  NAND3_X1 U9443 ( .A1(n6948), .A2(n9680), .A3(n6806), .ZN(n12180) );
  INV_X1 U9444 ( .A(n11425), .ZN(n11301) );
  OAI21_X1 U9445 ( .B1(n7449), .B2(n11218), .A(n11426), .ZN(n7448) );
  NAND2_X1 U9446 ( .A1(n13781), .A2(n15775), .ZN(n6970) );
  NAND2_X1 U9447 ( .A1(n11807), .A2(n8914), .ZN(n12104) );
  NAND2_X1 U9448 ( .A1(n11160), .A2(n8896), .ZN(n11516) );
  INV_X1 U9449 ( .A(n12882), .ZN(n11501) );
  NAND2_X1 U9450 ( .A1(n7725), .A2(n8908), .ZN(n11369) );
  NAND2_X1 U9451 ( .A1(n14169), .A2(n14170), .ZN(n14168) );
  OAI21_X1 U9452 ( .B1(n14182), .B2(n6809), .A(n6709), .ZN(n6984) );
  NAND2_X1 U9453 ( .A1(n14253), .A2(n6936), .ZN(P2_U3526) );
  NAND2_X1 U9454 ( .A1(n14331), .A2(n6938), .ZN(P2_U3494) );
  INV_X1 U9455 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n8193) );
  NAND2_X1 U9456 ( .A1(n7441), .A2(n8949), .ZN(n14038) );
  NAND2_X1 U9457 ( .A1(n8893), .A2(n8892), .ZN(n10479) );
  NAND2_X1 U9458 ( .A1(n8214), .A2(n8215), .ZN(n14388) );
  NAND2_X1 U9459 ( .A1(n8924), .A2(n8923), .ZN(n14182) );
  AND4_X2 U9460 ( .A1(n8332), .A2(n8330), .A3(n8331), .A4(n8333), .ZN(n12866)
         );
  AND2_X2 U9461 ( .A1(n7403), .A2(n7402), .ZN(n9795) );
  NAND2_X1 U9462 ( .A1(n11242), .A2(n11241), .ZN(n11351) );
  NOR2_X1 U9463 ( .A1(n6957), .A2(n10829), .ZN(n6973) );
  AND2_X1 U9464 ( .A1(n7416), .A2(n8903), .ZN(n6940) );
  NAND4_X2 U9465 ( .A1(n8448), .A2(n8447), .A3(n8446), .A4(n8445), .ZN(n13983)
         );
  INV_X1 U9466 ( .A(n8901), .ZN(n7419) );
  XNOR2_X1 U9467 ( .A(n15671), .B(n13983), .ZN(n13128) );
  NAND2_X1 U9468 ( .A1(n7425), .A2(n11369), .ZN(n11621) );
  NAND2_X2 U9469 ( .A1(n8938), .A2(n8875), .ZN(n8381) );
  NAND2_X1 U9470 ( .A1(n11094), .A2(n13130), .ZN(n8906) );
  NAND2_X1 U9471 ( .A1(n7415), .A2(n6940), .ZN(n11094) );
  NAND2_X1 U9472 ( .A1(n7417), .A2(n7419), .ZN(n7416) );
  OR2_X1 U9473 ( .A1(n13128), .A2(n7419), .ZN(n7418) );
  NAND2_X1 U9474 ( .A1(n9746), .A2(n12180), .ZN(n6941) );
  NAND2_X1 U9475 ( .A1(n6960), .A2(n6959), .ZN(n6942) );
  NAND2_X1 U9476 ( .A1(n7398), .A2(n7396), .ZN(n6943) );
  INV_X2 U9477 ( .A(n15496), .ZN(n11538) );
  XNOR2_X1 U9478 ( .A(n8378), .B(n7203), .ZN(n9980) );
  AOI21_X1 U9479 ( .B1(n11771), .B2(n7392), .A(n6790), .ZN(n7391) );
  NOR2_X1 U9480 ( .A1(n12070), .A2(n7393), .ZN(n7392) );
  OAI21_X1 U9481 ( .B1(n7446), .B2(n7445), .A(n13139), .ZN(n7444) );
  NOR2_X1 U9482 ( .A1(n8213), .A2(n8212), .ZN(n8214) );
  OAI211_X1 U9483 ( .C1(n13531), .C2(n15694), .A(n6947), .B(n6946), .ZN(
        P3_U3201) );
  NAND2_X1 U9484 ( .A1(n13530), .A2(n13529), .ZN(n6946) );
  NOR2_X1 U9485 ( .A1(n11907), .A2(n11906), .ZN(n11909) );
  AOI21_X1 U9486 ( .B1(n10981), .B2(n10980), .A(n7003), .ZN(n11319) );
  XNOR2_X1 U9487 ( .A(n13210), .B(n13208), .ZN(n13235) );
  NAND3_X1 U9488 ( .A1(n6972), .A2(n6971), .A3(n9040), .ZN(n9693) );
  NOR2_X1 U9489 ( .A1(n11011), .A2(n11010), .ZN(n11298) );
  NAND2_X1 U9490 ( .A1(n6975), .A2(n6974), .ZN(n7309) );
  NAND2_X1 U9491 ( .A1(n7397), .A2(n9899), .ZN(n7398) );
  NAND2_X1 U9492 ( .A1(n9793), .A2(n9990), .ZN(n10715) );
  NAND2_X1 U9493 ( .A1(n7460), .A2(n7461), .ZN(n13538) );
  OAI21_X1 U9494 ( .B1(n13778), .B2(n15782), .A(n6951), .ZN(n13720) );
  OAI21_X1 U9495 ( .B1(n13778), .B2(n15773), .A(n6832), .ZN(n13779) );
  OAI21_X2 U9496 ( .B1(n12537), .B2(n7358), .A(n7355), .ZN(n14983) );
  XNOR2_X1 U9497 ( .A(n6996), .B(n13518), .ZN(n13531) );
  INV_X1 U9498 ( .A(n10813), .ZN(n6952) );
  NOR2_X1 U9499 ( .A1(n11334), .A2(n11333), .ZN(n11446) );
  XNOR2_X1 U9500 ( .A(n7404), .B(n10886), .ZN(n10888) );
  NOR2_X1 U9501 ( .A1(n13463), .A2(n13462), .ZN(n13485) );
  NOR2_X1 U9502 ( .A1(n11447), .A2(n11446), .ZN(n11450) );
  NAND2_X1 U9503 ( .A1(n7206), .A2(n7204), .ZN(n7682) );
  XNOR2_X1 U9504 ( .A(n13387), .B(n13388), .ZN(n13378) );
  NAND3_X1 U9505 ( .A1(n7495), .A2(n10846), .A3(P3_REG1_REG_3__SCAN_IN), .ZN(
        n7494) );
  NOR2_X1 U9506 ( .A1(n10977), .A2(n10976), .ZN(n11326) );
  OAI21_X1 U9507 ( .B1(n13376), .B2(n13375), .A(n6981), .ZN(n6980) );
  INV_X1 U9508 ( .A(n9041), .ZN(n15714) );
  NAND3_X1 U9509 ( .A1(n6983), .A2(n6982), .A3(n9034), .ZN(n9041) );
  NAND2_X1 U9510 ( .A1(n11008), .A2(n7294), .ZN(n11011) );
  AOI21_X1 U9511 ( .B1(n13253), .B2(n13252), .A(n6792), .ZN(n13256) );
  INV_X1 U9512 ( .A(n12104), .ZN(n6967) );
  NAND2_X1 U9513 ( .A1(n14168), .A2(n8926), .ZN(n14162) );
  INV_X1 U9514 ( .A(n10592), .ZN(n6960) );
  NAND2_X1 U9515 ( .A1(n14038), .A2(n14226), .ZN(n6965) );
  NAND2_X1 U9516 ( .A1(n15714), .A2(n10585), .ZN(n9545) );
  NAND2_X1 U9517 ( .A1(n6965), .A2(n6963), .ZN(P2_U3236) );
  NAND2_X1 U9518 ( .A1(n10478), .A2(n8894), .ZN(n11161) );
  NAND2_X1 U9519 ( .A1(n11106), .A2(n7417), .ZN(n7415) );
  AND3_X2 U9520 ( .A1(n8194), .A2(n8195), .A3(n6799), .ZN(n8322) );
  INV_X1 U9521 ( .A(n8317), .ZN(n8210) );
  NAND3_X1 U9522 ( .A1(n7343), .A2(n7345), .A3(n11415), .ZN(n11417) );
  AND3_X4 U9523 ( .A1(n9857), .A2(n9853), .A3(n9854), .ZN(n15092) );
  OR2_X1 U9524 ( .A1(n12879), .A2(n12878), .ZN(n12885) );
  NAND2_X1 U9525 ( .A1(n13116), .A2(n13115), .ZN(n13165) );
  NAND2_X1 U9526 ( .A1(n7586), .A2(n7585), .ZN(n12912) );
  NAND2_X1 U9527 ( .A1(n7602), .A2(n6785), .ZN(n12929) );
  NAND2_X1 U9528 ( .A1(n7366), .A2(n7365), .ZN(n14877) );
  NAND2_X1 U9529 ( .A1(n12932), .A2(n12931), .ZN(n7547) );
  NAND2_X1 U9530 ( .A1(n6987), .A2(n6800), .ZN(n13032) );
  NAND2_X1 U9531 ( .A1(n13032), .A2(n13033), .ZN(n13031) );
  OAI21_X1 U9532 ( .B1(n12992), .B2(n12991), .A(n7741), .ZN(n13008) );
  NOR2_X1 U9533 ( .A1(n13360), .A2(n13361), .ZN(n13384) );
  NAND2_X1 U9534 ( .A1(n7463), .A2(n9657), .ZN(n13553) );
  XNOR2_X1 U9535 ( .A(n10985), .B(n10986), .ZN(n10870) );
  XNOR2_X1 U9536 ( .A(n13383), .B(n13388), .ZN(n13360) );
  NAND2_X1 U9537 ( .A1(n10818), .A2(n10765), .ZN(n11174) );
  NAND2_X1 U9538 ( .A1(n14218), .A2(n8921), .ZN(n7424) );
  INV_X1 U9539 ( .A(n6980), .ZN(n13387) );
  NOR2_X1 U9540 ( .A1(n10861), .A2(n7513), .ZN(n10972) );
  NOR2_X1 U9541 ( .A1(n10974), .A2(n10973), .ZN(n10977) );
  INV_X1 U9542 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n8233) );
  XNOR2_X1 U9543 ( .A(n11749), .B(n13207), .ZN(n11850) );
  NAND2_X2 U9544 ( .A1(n9573), .A2(n9574), .ZN(n11749) );
  NAND3_X1 U9545 ( .A1(n7590), .A2(n6789), .A3(n7591), .ZN(n13116) );
  NAND2_X1 U9546 ( .A1(n8772), .A2(n7666), .ZN(n7664) );
  NAND2_X1 U9547 ( .A1(n7703), .A2(n12560), .ZN(n12563) );
  NAND2_X1 U9548 ( .A1(n14435), .A2(n7389), .ZN(n7388) );
  NAND2_X1 U9549 ( .A1(n7684), .A2(n8256), .ZN(n8469) );
  NAND2_X1 U9550 ( .A1(n13372), .A2(n6833), .ZN(n13419) );
  NAND2_X1 U9551 ( .A1(n10863), .A2(n6780), .ZN(n10981) );
  AOI21_X1 U9552 ( .B1(n13495), .B2(n13494), .A(n13493), .ZN(n13516) );
  NAND2_X1 U9553 ( .A1(n14140), .A2(n6986), .ZN(n14139) );
  INV_X1 U9554 ( .A(n6984), .ZN(n14169) );
  NAND2_X1 U9555 ( .A1(n11355), .A2(n11354), .ZN(n11765) );
  NAND2_X1 U9556 ( .A1(n14546), .A2(n14457), .ZN(n14463) );
  INV_X1 U9557 ( .A(n9925), .ZN(n7397) );
  XNOR2_X1 U9558 ( .A(n9852), .B(n14445), .ZN(n11024) );
  NAND2_X1 U9559 ( .A1(n6979), .A2(n6977), .ZN(P3_U3486) );
  OAI22_X1 U9560 ( .A1(n13782), .A2(n13777), .B1(n15784), .B2(n9443), .ZN(
        n6978) );
  NAND2_X1 U9561 ( .A1(n13781), .A2(n15784), .ZN(n6979) );
  XNOR2_X1 U9562 ( .A(n11438), .B(n11445), .ZN(n11327) );
  AND2_X2 U9563 ( .A1(n9004), .A2(n7625), .ZN(n7454) );
  INV_X1 U9564 ( .A(n13124), .ZN(n11162) );
  INV_X1 U9565 ( .A(n7432), .ZN(n7431) );
  NAND2_X1 U9566 ( .A1(n8932), .A2(n8931), .ZN(n14081) );
  NAND2_X1 U9567 ( .A1(n7229), .A2(n7228), .ZN(n9001) );
  NAND3_X1 U9568 ( .A1(n7587), .A2(n12901), .A3(n12900), .ZN(n7586) );
  NAND3_X1 U9569 ( .A1(n13021), .A2(n13022), .A3(n6805), .ZN(n6987) );
  OAI21_X1 U9570 ( .B1(n15769), .B2(n13723), .A(n13722), .ZN(n13781) );
  NAND3_X1 U9571 ( .A1(n7139), .A2(n7140), .A3(P3_ADDR_REG_19__SCAN_IN), .ZN(
        n7283) );
  NAND2_X1 U9572 ( .A1(n13270), .A2(n7298), .ZN(n7296) );
  NAND2_X1 U9573 ( .A1(n7424), .A2(n7423), .ZN(n8924) );
  NAND2_X1 U9574 ( .A1(n7221), .A2(n7225), .ZN(n8600) );
  INV_X1 U9575 ( .A(n7444), .ZN(n7443) );
  INV_X1 U9576 ( .A(n11025), .ZN(n7396) );
  NAND2_X2 U9577 ( .A1(n14664), .A2(n14665), .ZN(n14663) );
  NAND2_X2 U9578 ( .A1(n11765), .A2(n6999), .ZN(n11770) );
  NOR2_X1 U9579 ( .A1(n9259), .A2(n9500), .ZN(n9504) );
  NAND2_X2 U9580 ( .A1(n11754), .A2(n9574), .ZN(n12024) );
  XNOR2_X2 U9581 ( .A(n9087), .B(n11425), .ZN(n11218) );
  NAND2_X2 U9582 ( .A1(n9191), .A2(n9190), .ZN(n11997) );
  NAND2_X1 U9583 ( .A1(n7011), .A2(n8409), .ZN(n10534) );
  NAND2_X1 U9584 ( .A1(n7011), .A2(n7010), .ZN(n10445) );
  OR2_X1 U9585 ( .A1(n10444), .A2(n10443), .ZN(n7010) );
  NAND2_X1 U9586 ( .A1(n10444), .A2(n10443), .ZN(n7011) );
  XNOR2_X1 U9587 ( .A(n8393), .B(n6837), .ZN(n10390) );
  NAND2_X2 U9588 ( .A1(n7012), .A2(n8741), .ZN(n8754) );
  NAND3_X1 U9589 ( .A1(n7021), .A2(n7014), .A3(n7013), .ZN(n11119) );
  NAND3_X1 U9590 ( .A1(n10533), .A2(n7018), .A3(n10721), .ZN(n7013) );
  NAND2_X1 U9591 ( .A1(n10533), .A2(n8436), .ZN(n10567) );
  OAI21_X1 U9592 ( .B1(n7016), .B2(n7019), .A(n8453), .ZN(n10722) );
  INV_X1 U9593 ( .A(n10533), .ZN(n7016) );
  INV_X1 U9594 ( .A(n7019), .ZN(n7018) );
  INV_X1 U9595 ( .A(n8436), .ZN(n7020) );
  NAND2_X1 U9596 ( .A1(n8486), .A2(n8487), .ZN(n11121) );
  NAND2_X2 U9597 ( .A1(n7032), .A2(n8859), .ZN(n8992) );
  XNOR2_X2 U9598 ( .A(n7031), .B(n7030), .ZN(n8859) );
  NAND3_X1 U9599 ( .A1(n12255), .A2(n7581), .A3(n13896), .ZN(n7041) );
  NAND2_X1 U9600 ( .A1(n8702), .A2(n7052), .ZN(n7046) );
  NAND3_X1 U9601 ( .A1(n7054), .A2(n12619), .A3(n7053), .ZN(n12623) );
  NAND2_X1 U9602 ( .A1(n12615), .A2(n6797), .ZN(n7053) );
  NAND2_X1 U9603 ( .A1(n6700), .A2(n12611), .ZN(n7054) );
  INV_X1 U9604 ( .A(n12616), .ZN(n7055) );
  NAND2_X1 U9605 ( .A1(n12635), .A2(n7058), .ZN(n7057) );
  NAND2_X1 U9606 ( .A1(n7057), .A2(n7056), .ZN(n12644) );
  XNOR2_X2 U9607 ( .A(n7062), .B(P1_IR_REG_22__SCAN_IN), .ZN(n15244) );
  OAI21_X2 U9608 ( .B1(n9826), .B2(P1_IR_REG_21__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n7062) );
  NAND2_X1 U9609 ( .A1(n12727), .A2(n7067), .ZN(n7065) );
  NAND2_X1 U9610 ( .A1(n7065), .A2(n7066), .ZN(n12734) );
  NAND2_X1 U9611 ( .A1(n12758), .A2(n12757), .ZN(n7072) );
  NAND2_X1 U9612 ( .A1(n7077), .A2(n6804), .ZN(n7714) );
  NAND3_X1 U9613 ( .A1(n12747), .A2(n7078), .A3(n12746), .ZN(n7077) );
  NAND2_X1 U9614 ( .A1(n12652), .A2(n7083), .ZN(n7081) );
  NAND2_X1 U9615 ( .A1(n7081), .A2(n7082), .ZN(n12664) );
  NAND2_X1 U9616 ( .A1(n7089), .A2(n7087), .ZN(n12707) );
  NAND2_X1 U9617 ( .A1(n7088), .A2(n7090), .ZN(n7087) );
  NAND3_X1 U9618 ( .A1(n7093), .A2(n12672), .A3(n12691), .ZN(n7088) );
  NAND3_X1 U9619 ( .A1(n12667), .A2(n12666), .A3(n7090), .ZN(n7089) );
  NAND2_X1 U9620 ( .A1(n7091), .A2(n12691), .ZN(n7090) );
  INV_X1 U9621 ( .A(n12684), .ZN(n7093) );
  INV_X1 U9622 ( .A(n7097), .ZN(n9144) );
  NAND2_X1 U9623 ( .A1(n7098), .A2(n9692), .ZN(P3_U3296) );
  NAND2_X1 U9624 ( .A1(n7099), .A2(n9677), .ZN(n7098) );
  NAND3_X1 U9625 ( .A1(n7102), .A2(n6706), .A3(n7100), .ZN(n7099) );
  NOR2_X1 U9626 ( .A1(n7101), .A2(n6733), .ZN(n7100) );
  NAND2_X1 U9627 ( .A1(n7312), .A2(n7311), .ZN(n7102) );
  NAND2_X1 U9628 ( .A1(n9242), .A2(n7105), .ZN(n7104) );
  NAND3_X1 U9629 ( .A1(n7104), .A2(n7319), .A3(n7103), .ZN(n9288) );
  NAND2_X1 U9630 ( .A1(n9369), .A2(n6834), .ZN(n7109) );
  NAND3_X1 U9631 ( .A1(n7120), .A2(n7119), .A3(n7118), .ZN(n7117) );
  NAND4_X1 U9632 ( .A1(n9664), .A2(n10746), .A3(n9663), .A4(n9662), .ZN(n7118)
         );
  NAND3_X1 U9633 ( .A1(n13537), .A2(n9661), .A3(n9771), .ZN(n7120) );
  OAI21_X1 U9634 ( .B1(n15262), .B2(n7133), .A(n7132), .ZN(n7134) );
  AND2_X2 U9635 ( .A1(n11628), .A2(n11783), .ZN(n11713) );
  NOR2_X2 U9636 ( .A1(n11368), .A2(n12947), .ZN(n11628) );
  NAND2_X1 U9637 ( .A1(n14074), .A2(n14068), .ZN(n14062) );
  NAND2_X1 U9638 ( .A1(n14222), .A2(n6685), .ZN(n7156) );
  NAND2_X1 U9639 ( .A1(n7157), .A2(n7156), .ZN(n14151) );
  INV_X1 U9640 ( .A(n7166), .ZN(n14137) );
  NAND2_X1 U9641 ( .A1(n7534), .A2(n7174), .ZN(n7169) );
  AOI21_X1 U9642 ( .B1(n7534), .B2(n7172), .A(n7170), .ZN(n8991) );
  NAND2_X1 U9643 ( .A1(n8817), .A2(n8383), .ZN(n8388) );
  AND2_X4 U9644 ( .A1(n8218), .A2(n8216), .ZN(n8817) );
  NAND2_X1 U9645 ( .A1(n8229), .A2(n8206), .ZN(n8315) );
  NAND2_X1 U9646 ( .A1(n8317), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8211) );
  NAND2_X1 U9647 ( .A1(n6794), .A2(n12360), .ZN(n15043) );
  NAND2_X1 U9648 ( .A1(n14986), .A2(n7192), .ZN(n14923) );
  INV_X1 U9649 ( .A(n7197), .ZN(n14943) );
  NAND2_X1 U9650 ( .A1(n14899), .A2(n15125), .ZN(n14879) );
  NAND2_X1 U9651 ( .A1(n12448), .A2(n7201), .ZN(n7200) );
  NAND2_X2 U9652 ( .A1(n12448), .A2(n9975), .ZN(n9888) );
  OAI22_X1 U9653 ( .A1(n9981), .A2(n9950), .B1(n8234), .B2(n8253), .ZN(n7201)
         );
  NAND3_X1 U9654 ( .A1(n7680), .A2(n7678), .A3(n7679), .ZN(n8756) );
  NAND2_X1 U9655 ( .A1(n8506), .A2(n7208), .ZN(n7206) );
  OAI21_X1 U9656 ( .B1(n8506), .B2(n7210), .A(n7208), .ZN(n8541) );
  NAND2_X1 U9657 ( .A1(n8678), .A2(n7216), .ZN(n7215) );
  NAND2_X1 U9658 ( .A1(n8561), .A2(n7222), .ZN(n7218) );
  NAND2_X1 U9659 ( .A1(n7218), .A2(n7219), .ZN(n8622) );
  NAND2_X1 U9660 ( .A1(n8561), .A2(n7226), .ZN(n7221) );
  NAND2_X1 U9661 ( .A1(n7239), .A2(P2_ADDR_REG_18__SCAN_IN), .ZN(n7238) );
  NAND2_X1 U9662 ( .A1(n15247), .A2(n15248), .ZN(n7239) );
  INV_X1 U9663 ( .A(n7240), .ZN(n15799) );
  XNOR2_X1 U9664 ( .A(n7812), .B(n7809), .ZN(n15800) );
  XNOR2_X1 U9665 ( .A(n7808), .B(n7241), .ZN(n7812) );
  INV_X1 U9666 ( .A(n7810), .ZN(n7241) );
  INV_X1 U9667 ( .A(n12393), .ZN(n7245) );
  NAND2_X1 U9668 ( .A1(n14953), .A2(n7253), .ZN(n7250) );
  NAND2_X1 U9669 ( .A1(n14888), .A2(n7262), .ZN(n7257) );
  OAI21_X2 U9670 ( .B1(n14888), .B2(n7261), .A(n7258), .ZN(n12575) );
  INV_X1 U9671 ( .A(n7272), .ZN(n7271) );
  NAND2_X1 U9672 ( .A1(n7271), .A2(n7273), .ZN(n12287) );
  NOR2_X1 U9673 ( .A1(n15409), .A2(n14698), .ZN(n7274) );
  NAND2_X1 U9674 ( .A1(n14998), .A2(n6798), .ZN(n7275) );
  NAND2_X1 U9675 ( .A1(n7275), .A2(n7276), .ZN(n14968) );
  INV_X1 U9676 ( .A(n12620), .ZN(n11410) );
  NAND3_X1 U9677 ( .A1(n8232), .A2(P2_ADDR_REG_19__SCAN_IN), .A3(n15251), .ZN(
        n7284) );
  NAND2_X1 U9678 ( .A1(n11823), .A2(n6705), .ZN(n11933) );
  NAND2_X1 U9679 ( .A1(n13191), .A2(n13190), .ZN(n13279) );
  NOR2_X2 U9680 ( .A1(n9259), .A2(n7306), .ZN(n9290) );
  NAND2_X1 U9681 ( .A1(n9339), .A2(n9338), .ZN(n7310) );
  XNOR2_X1 U9682 ( .A(n7313), .B(n9769), .ZN(n7312) );
  NAND2_X1 U9683 ( .A1(n7314), .A2(n6811), .ZN(n7313) );
  NAND2_X1 U9684 ( .A1(n9028), .A2(n9057), .ZN(n7316) );
  INV_X1 U9685 ( .A(n9027), .ZN(n7318) );
  NAND2_X1 U9686 ( .A1(n9047), .A2(n9046), .ZN(n9058) );
  NAND2_X1 U9687 ( .A1(n9028), .A2(n9027), .ZN(n9047) );
  NAND2_X1 U9688 ( .A1(n7332), .A2(n7330), .ZN(n9470) );
  NAND2_X1 U9689 ( .A1(n7332), .A2(n7331), .ZN(n9472) );
  INV_X1 U9690 ( .A(n10686), .ZN(n15085) );
  INV_X1 U9691 ( .A(n12448), .ZN(n7342) );
  NAND2_X1 U9692 ( .A1(n7346), .A2(n11577), .ZN(n7343) );
  AND2_X1 U9693 ( .A1(n7344), .A2(n12801), .ZN(n7346) );
  NAND2_X1 U9694 ( .A1(n11944), .A2(n6729), .ZN(n7350) );
  NAND2_X1 U9695 ( .A1(n12537), .A2(n12536), .ZN(n15017) );
  NAND4_X1 U9696 ( .A1(n7364), .A2(n7720), .A3(n9846), .A4(n9794), .ZN(n7719)
         );
  NAND2_X1 U9697 ( .A1(n14904), .A2(n7367), .ZN(n7366) );
  NAND2_X1 U9698 ( .A1(n14663), .A2(n14523), .ZN(n14524) );
  OAI211_X1 U9699 ( .C1(n14663), .C2(n6810), .A(n7370), .B(n7368), .ZN(n14568)
         );
  NAND2_X1 U9700 ( .A1(n14663), .A2(n7369), .ZN(n7368) );
  NOR2_X1 U9701 ( .A1(n7372), .A2(n14560), .ZN(n7369) );
  OAI22_X1 U9702 ( .A1(n7372), .A2(n7371), .B1(n14560), .B2(n7374), .ZN(n7370)
         );
  NOR2_X1 U9703 ( .A1(n14525), .A2(n14560), .ZN(n7371) );
  INV_X1 U9704 ( .A(n14560), .ZN(n7373) );
  NAND2_X1 U9705 ( .A1(n7376), .A2(n7377), .ZN(n14533) );
  NAND2_X1 U9706 ( .A1(n14463), .A2(n7379), .ZN(n7376) );
  INV_X1 U9707 ( .A(n7381), .ZN(n9799) );
  NAND2_X1 U9708 ( .A1(n7388), .A2(n7386), .ZN(n14543) );
  NAND2_X1 U9709 ( .A1(n14435), .A2(n14434), .ZN(n14602) );
  NOR2_X1 U9710 ( .A1(n14441), .A2(n7390), .ZN(n7389) );
  INV_X1 U9711 ( .A(n14434), .ZN(n7390) );
  NAND2_X2 U9712 ( .A1(n14636), .A2(n14635), .ZN(n14634) );
  NAND3_X1 U9713 ( .A1(n7396), .A2(n10658), .A3(n10659), .ZN(n7395) );
  NAND2_X1 U9714 ( .A1(n10657), .A2(n7399), .ZN(n7401) );
  INV_X1 U9715 ( .A(n7401), .ZN(n11079) );
  NOR2_X2 U9716 ( .A1(n9792), .A2(n9791), .ZN(n9793) );
  NAND2_X1 U9717 ( .A1(n13487), .A2(n7411), .ZN(n7409) );
  AND2_X1 U9718 ( .A1(n7418), .A2(n8902), .ZN(n7417) );
  INV_X1 U9719 ( .A(n15652), .ZN(n11158) );
  NAND2_X2 U9720 ( .A1(n7433), .A2(n7431), .ZN(n15652) );
  INV_X2 U9721 ( .A(n15688), .ZN(n7435) );
  NAND2_X1 U9722 ( .A1(n11217), .A2(n9088), .ZN(n11427) );
  NAND2_X1 U9723 ( .A1(n11219), .A2(n11218), .ZN(n11217) );
  OR2_X1 U9724 ( .A1(n13566), .A2(n7462), .ZN(n7460) );
  NAND2_X1 U9725 ( .A1(n13566), .A2(n7458), .ZN(n7457) );
  NAND2_X1 U9726 ( .A1(n13566), .A2(n9656), .ZN(n7463) );
  NAND2_X1 U9727 ( .A1(n12024), .A2(n7469), .ZN(n7467) );
  NAND2_X1 U9728 ( .A1(n7467), .A2(n7468), .ZN(n11995) );
  NAND2_X1 U9729 ( .A1(n13671), .A2(n7478), .ZN(n7474) );
  NAND2_X1 U9730 ( .A1(n7474), .A2(n7475), .ZN(n13642) );
  XNOR2_X2 U9731 ( .A(n10674), .B(n15718), .ZN(n9695) );
  OAI21_X2 U9732 ( .B1(n12267), .B2(n7484), .A(n9607), .ZN(n13709) );
  AND2_X2 U9733 ( .A1(n9678), .A2(n9012), .ZN(n9679) );
  AND2_X2 U9734 ( .A1(n9683), .A2(n9684), .ZN(n9678) );
  NAND2_X1 U9735 ( .A1(n11174), .A2(n11175), .ZN(n7485) );
  OAI21_X1 U9736 ( .B1(n11175), .B2(n11174), .A(n7485), .ZN(n11176) );
  INV_X1 U9737 ( .A(n10765), .ZN(n7486) );
  INV_X1 U9738 ( .A(n10826), .ZN(n7489) );
  NOR2_X1 U9739 ( .A1(n7486), .A2(n9019), .ZN(n7487) );
  NAND2_X1 U9740 ( .A1(n7490), .A2(n9019), .ZN(n10817) );
  NAND2_X1 U9741 ( .A1(n7500), .A2(n7502), .ZN(n10862) );
  INV_X1 U9742 ( .A(n7504), .ZN(n7500) );
  NOR2_X1 U9743 ( .A1(n7504), .A2(n7501), .ZN(n10973) );
  NAND2_X1 U9744 ( .A1(n7502), .A2(P3_REG1_REG_7__SCAN_IN), .ZN(n7501) );
  NAND2_X1 U9745 ( .A1(n10790), .A2(n7503), .ZN(n7502) );
  NOR2_X1 U9746 ( .A1(n10790), .A2(n10789), .ZN(n10861) );
  NAND2_X1 U9747 ( .A1(n7515), .A2(n7516), .ZN(n7514) );
  NAND2_X1 U9748 ( .A1(n11443), .A2(n7517), .ZN(n7515) );
  AOI21_X1 U9749 ( .B1(n11442), .B2(n7517), .A(n11977), .ZN(n7516) );
  INV_X1 U9750 ( .A(n11913), .ZN(n7518) );
  NOR2_X1 U9751 ( .A1(n11915), .A2(n9194), .ZN(n11978) );
  OR2_X1 U9752 ( .A1(n7520), .A2(n11981), .ZN(n7519) );
  NAND2_X1 U9753 ( .A1(n13507), .A2(n6843), .ZN(n7521) );
  OAI211_X1 U9754 ( .C1(n13507), .C2(n7522), .A(n7521), .B(n7529), .ZN(n13527)
         );
  NAND2_X2 U9755 ( .A1(n7544), .A2(n7545), .ZN(n13987) );
  NAND2_X1 U9756 ( .A1(n11501), .A2(n13987), .ZN(n7531) );
  NAND3_X1 U9757 ( .A1(n8976), .A2(n6708), .A3(n8975), .ZN(n7539) );
  NAND2_X1 U9758 ( .A1(n7539), .A2(n7540), .ZN(n12101) );
  NAND2_X1 U9759 ( .A1(n13987), .A2(n8753), .ZN(n8372) );
  INV_X1 U9760 ( .A(n8372), .ZN(n8371) );
  NAND3_X1 U9761 ( .A1(n7548), .A2(n7547), .A3(n7552), .ZN(n7546) );
  NAND2_X1 U9762 ( .A1(n12928), .A2(n12927), .ZN(n7548) );
  NAND3_X1 U9763 ( .A1(n7551), .A2(n7550), .A3(n7553), .ZN(n7549) );
  NAND2_X1 U9764 ( .A1(n12928), .A2(n6791), .ZN(n7551) );
  NAND2_X1 U9765 ( .A1(n8754), .A2(n7555), .ZN(n7554) );
  OAI211_X1 U9766 ( .C1(n8754), .C2(n6808), .A(n6710), .B(n7554), .ZN(n13880)
         );
  NAND2_X1 U9767 ( .A1(n12847), .A2(n7569), .ZN(n7568) );
  OAI211_X1 U9768 ( .C1(n12847), .C2(n7570), .A(n7568), .B(n7746), .ZN(
        P2_U3192) );
  NAND2_X1 U9769 ( .A1(n15341), .A2(n7578), .ZN(n8558) );
  INV_X1 U9770 ( .A(n13025), .ZN(n7583) );
  NAND2_X1 U9771 ( .A1(n12912), .A2(n12913), .ZN(n12911) );
  INV_X1 U9772 ( .A(n12904), .ZN(n7589) );
  NAND2_X1 U9773 ( .A1(n12904), .A2(n7588), .ZN(n7587) );
  OAI21_X1 U9774 ( .B1(n7600), .B2(n12944), .A(n7599), .ZN(n12955) );
  NAND3_X1 U9775 ( .A1(n12917), .A2(n12916), .A3(n6807), .ZN(n7602) );
  OAI21_X1 U9776 ( .B1(n13012), .B2(n7610), .A(n7609), .ZN(n13019) );
  NAND2_X1 U9777 ( .A1(n7607), .A2(n7608), .ZN(n13018) );
  NAND2_X1 U9778 ( .A1(n13012), .A2(n7609), .ZN(n7607) );
  NAND2_X1 U9779 ( .A1(n8202), .A2(n7615), .ZN(n8827) );
  AOI21_X1 U9780 ( .B1(n11052), .B2(n9695), .A(n6795), .ZN(n7742) );
  NOR2_X1 U9781 ( .A1(n11426), .A2(n7620), .ZN(n7619) );
  NAND2_X1 U9782 ( .A1(n13545), .A2(n7621), .ZN(n13535) );
  NAND2_X1 U9783 ( .A1(n7622), .A2(n7623), .ZN(n9720) );
  NAND2_X1 U9784 ( .A1(n13626), .A2(n9718), .ZN(n7622) );
  NAND3_X1 U9785 ( .A1(n9080), .A2(n9004), .A3(n9003), .ZN(n9221) );
  AOI21_X1 U9786 ( .B1(n11794), .B2(n7626), .A(n6803), .ZN(n7628) );
  NAND2_X1 U9787 ( .A1(n9710), .A2(n7627), .ZN(n7629) );
  INV_X1 U9788 ( .A(n9710), .ZN(n7632) );
  NAND2_X1 U9789 ( .A1(n13588), .A2(n6688), .ZN(n7635) );
  INV_X1 U9790 ( .A(n7636), .ZN(n13587) );
  INV_X1 U9791 ( .A(n9714), .ZN(n7637) );
  NAND2_X1 U9792 ( .A1(n7648), .A2(n7649), .ZN(n13636) );
  NAND2_X1 U9793 ( .A1(n13661), .A2(n7652), .ZN(n7648) );
  INV_X1 U9794 ( .A(n13681), .ZN(n7656) );
  NAND2_X1 U9795 ( .A1(n9678), .A2(n7657), .ZN(n9015) );
  INV_X1 U9796 ( .A(n8246), .ZN(n7662) );
  NAND2_X1 U9797 ( .A1(n7664), .A2(n7665), .ZN(n8883) );
  NAND3_X1 U9798 ( .A1(n7680), .A2(n6835), .A3(n7678), .ZN(n8306) );
  NAND2_X1 U9799 ( .A1(n8303), .A2(n8302), .ZN(n8304) );
  NAND2_X1 U9800 ( .A1(n8303), .A2(n7681), .ZN(n7680) );
  NAND2_X1 U9801 ( .A1(n8455), .A2(n8254), .ZN(n7684) );
  XNOR2_X1 U9802 ( .A(n7690), .B(n12791), .ZN(n12830) );
  INV_X1 U9803 ( .A(n7690), .ZN(n12827) );
  NAND2_X1 U9804 ( .A1(n7691), .A2(n12828), .ZN(n7693) );
  XNOR2_X1 U9805 ( .A(n12824), .B(n12593), .ZN(n7691) );
  NAND2_X1 U9806 ( .A1(n7692), .A2(n12836), .ZN(n12837) );
  NAND2_X1 U9807 ( .A1(n12557), .A2(n12556), .ZN(n7703) );
  NAND2_X1 U9808 ( .A1(n12730), .A2(n7706), .ZN(n7705) );
  NAND3_X1 U9809 ( .A1(n12628), .A2(n12627), .A3(n7709), .ZN(n7712) );
  NAND2_X1 U9810 ( .A1(n12631), .A2(n7710), .ZN(n7709) );
  NAND2_X1 U9811 ( .A1(n7712), .A2(n7711), .ZN(n12635) );
  NAND2_X1 U9812 ( .A1(n12752), .A2(n7713), .ZN(n7715) );
  NAND2_X1 U9813 ( .A1(n7714), .A2(n7716), .ZN(n12753) );
  NAND2_X1 U9814 ( .A1(n7717), .A2(n12751), .ZN(n7716) );
  INV_X1 U9815 ( .A(n12752), .ZN(n7717) );
  NAND2_X1 U9816 ( .A1(n9814), .A2(n6736), .ZN(n9816) );
  NAND2_X1 U9817 ( .A1(n7723), .A2(n7724), .ZN(n12727) );
  OAI211_X1 U9818 ( .C1(n12723), .C2(n12725), .A(n12722), .B(n12721), .ZN(
        n7723) );
  NAND2_X1 U9819 ( .A1(n10696), .A2(n10695), .ZN(n10952) );
  INV_X1 U9820 ( .A(n12797), .ZN(n10696) );
  NAND2_X1 U9821 ( .A1(n14968), .A2(n14979), .ZN(n14967) );
  MUX2_X1 U9822 ( .A(n15211), .B(P1_REG1_REG_27__SCAN_IN), .S(n15534), .Z(
        P1_U3555) );
  MUX2_X1 U9823 ( .A(n15211), .B(P1_REG0_REG_27__SCAN_IN), .S(n15524), .Z(
        P1_U3523) );
  XNOR2_X1 U9824 ( .A(n9800), .B(P1_IR_REG_24__SCAN_IN), .ZN(n9900) );
  INV_X1 U9825 ( .A(n14569), .ZN(n14571) );
  CLKBUF_X1 U9826 ( .A(n9900), .Z(n9906) );
  NAND2_X1 U9827 ( .A1(n10578), .A2(n10577), .ZN(n10576) );
  AND2_X1 U9828 ( .A1(n13205), .A2(n13204), .ZN(n13206) );
  CLKBUF_X1 U9829 ( .A(n13709), .Z(n13711) );
  NAND2_X1 U9830 ( .A1(n8999), .A2(n8998), .ZN(n9000) );
  INV_X1 U9831 ( .A(n10830), .ZN(n15747) );
  XNOR2_X1 U9832 ( .A(n12575), .B(n12821), .ZN(n12529) );
  CLKBUF_X1 U9833 ( .A(n13671), .Z(n13672) );
  NAND2_X1 U9834 ( .A1(n8318), .A2(n8317), .ZN(n8875) );
  NAND2_X1 U9835 ( .A1(n12737), .A2(n12736), .ZN(n12743) );
  MUX2_X2 U9836 ( .A(P3_REG0_REG_29__SCAN_IN), .B(n9784), .S(n15775), .Z(n9785) );
  INV_X1 U9837 ( .A(n12570), .ZN(n15117) );
  NAND2_X1 U9838 ( .A1(n12733), .A2(n12732), .ZN(n12744) );
  NAND3_X1 U9839 ( .A1(n12607), .A2(n12606), .A3(n12605), .ZN(n12612) );
  BUF_X2 U9840 ( .A(n8381), .Z(n10076) );
  INV_X1 U9841 ( .A(n12613), .ZN(n12614) );
  NOR2_X1 U9842 ( .A1(n8827), .A2(P2_IR_REG_22__SCAN_IN), .ZN(n8855) );
  OAI21_X2 U9843 ( .B1(n8827), .B2(n8312), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n8314) );
  NOR2_X1 U9844 ( .A1(n9795), .A2(n9847), .ZN(n9848) );
  OAI21_X1 U9845 ( .B1(n12711), .B2(n12709), .A(n12708), .ZN(n12713) );
  OR2_X1 U9846 ( .A1(n15244), .A2(n12594), .ZN(n9920) );
  NAND2_X1 U9847 ( .A1(n9388), .A2(P3_REG1_REG_4__SCAN_IN), .ZN(n9074) );
  AOI21_X1 U9848 ( .B1(n13829), .B2(n9184), .A(n9493), .ZN(n15309) );
  INV_X1 U9849 ( .A(n12866), .ZN(n13989) );
  NAND2_X1 U9850 ( .A1(n12018), .A2(n15759), .ZN(n9171) );
  AND2_X4 U9851 ( .A1(n9018), .A2(n9020), .ZN(n9300) );
  INV_X1 U9852 ( .A(n9018), .ZN(n13837) );
  NAND2_X1 U9853 ( .A1(n9709), .A2(n9708), .ZN(n9710) );
  INV_X1 U9854 ( .A(n8817), .ZN(n8874) );
  AOI21_X1 U9855 ( .B1(n12839), .B2(n12838), .A(n12837), .ZN(n12845) );
  INV_X1 U9856 ( .A(n14382), .ZN(n8213) );
  INV_X1 U9857 ( .A(n14040), .ZN(n8999) );
  AOI21_X1 U9858 ( .B1(n12847), .B2(n12846), .A(n13935), .ZN(n12856) );
  NAND4_X2 U9859 ( .A1(n9869), .A2(n9868), .A3(n9867), .A4(n9866), .ZN(n14707)
         );
  NAND2_X1 U9860 ( .A1(n9865), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n9868) );
  INV_X1 U9861 ( .A(n12805), .ZN(n11835) );
  INV_X1 U9862 ( .A(n14921), .ZN(n14926) );
  AND2_X1 U9863 ( .A1(n9812), .A2(n13826), .ZN(n10860) );
  OR2_X1 U9864 ( .A1(n13176), .A2(n13777), .ZN(n7726) );
  OR2_X1 U9865 ( .A1(n13176), .A2(n13825), .ZN(n7727) );
  INV_X1 U9866 ( .A(n13540), .ZN(n13780) );
  OR2_X1 U9867 ( .A1(n13809), .A2(n13629), .ZN(n7728) );
  XNOR2_X1 U9868 ( .A(n14843), .B(n14685), .ZN(n7729) );
  NAND2_X1 U9869 ( .A1(n15616), .A2(n8369), .ZN(n7730) );
  AND2_X1 U9870 ( .A1(n8392), .A2(n8391), .ZN(n7731) );
  INV_X1 U9871 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n11262) );
  OR2_X1 U9872 ( .A1(n12448), .A2(n14750), .ZN(n7732) );
  NAND2_X1 U9873 ( .A1(n8554), .A2(n8555), .ZN(n7733) );
  INV_X1 U9874 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n9813) );
  XOR2_X1 U9875 ( .A(n9039), .B(P2_DATAO_REG_0__SCAN_IN), .Z(n7734) );
  INV_X1 U9876 ( .A(P3_ADDR_REG_8__SCAN_IN), .ZN(n8104) );
  AND2_X1 U9877 ( .A1(n8271), .A2(n8270), .ZN(n7735) );
  AND2_X1 U9878 ( .A1(n7202), .A2(P1_U3086), .ZN(n12056) );
  INV_X1 U9879 ( .A(n13501), .ZN(n13494) );
  INV_X1 U9880 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n10671) );
  INV_X1 U9881 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n10652) );
  INV_X1 U9882 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n12566) );
  INV_X1 U9883 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n11960) );
  NOR2_X1 U9884 ( .A1(n9601), .A2(n9511), .ZN(n7736) );
  AND2_X1 U9885 ( .A1(n12986), .A2(n12985), .ZN(n7737) );
  INV_X1 U9886 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n11256) );
  OR2_X1 U9887 ( .A1(n14210), .A2(n13863), .ZN(n7739) );
  INV_X1 U9888 ( .A(P3_IR_REG_2__SCAN_IN), .ZN(n9049) );
  INV_X1 U9889 ( .A(n12813), .ZN(n12392) );
  INV_X1 U9890 ( .A(n12980), .ZN(n8888) );
  INV_X1 U9891 ( .A(n12804), .ZN(n11416) );
  AND2_X1 U9892 ( .A1(n12993), .A2(n12990), .ZN(n7741) );
  AND4_X1 U9893 ( .A1(n15108), .A2(n15107), .A3(n15106), .A4(n15105), .ZN(
        n7743) );
  AND4_X1 U9894 ( .A1(n12821), .A2(n12820), .A3(n14859), .A4(n12819), .ZN(
        n7744) );
  AND2_X1 U9895 ( .A1(n13078), .A2(n13077), .ZN(n7745) );
  AND2_X1 U9896 ( .A1(n8880), .A2(n8879), .ZN(n7746) );
  INV_X1 U9897 ( .A(n13548), .ZN(n13577) );
  AOI21_X1 U9898 ( .B1(n13539), .B2(n9300), .A(n9456), .ZN(n13549) );
  INV_X1 U9899 ( .A(n6675), .ZN(n9729) );
  INV_X1 U9900 ( .A(n14379), .ZN(n8998) );
  NAND2_X1 U9901 ( .A1(n12863), .A2(n12871), .ZN(n12868) );
  NAND2_X1 U9902 ( .A1(n12873), .A2(n12872), .ZN(n12876) );
  INV_X1 U9903 ( .A(n12897), .ZN(n12898) );
  INV_X1 U9904 ( .A(n12913), .ZN(n12914) );
  INV_X1 U9905 ( .A(n12930), .ZN(n12931) );
  INV_X1 U9906 ( .A(n12994), .ZN(n12989) );
  NAND2_X1 U9907 ( .A1(n7737), .A2(n12989), .ZN(n12990) );
  INV_X1 U9908 ( .A(n13033), .ZN(n13034) );
  MUX2_X1 U9909 ( .A(n14688), .B(n14866), .S(n12789), .Z(n12752) );
  INV_X1 U9910 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n8204) );
  INV_X1 U9911 ( .A(n13355), .ZN(n13180) );
  NAND2_X1 U9912 ( .A1(n11194), .A2(P3_REG2_REG_2__SCAN_IN), .ZN(n10753) );
  INV_X1 U9913 ( .A(P3_IR_REG_26__SCAN_IN), .ZN(n9013) );
  INV_X1 U9914 ( .A(n13990), .ZN(n8364) );
  OAI22_X1 U9915 ( .A1(n15092), .A2(n14557), .B1(n10686), .B2(n6667), .ZN(
        n9860) );
  AND2_X1 U9916 ( .A1(n10594), .A2(n10593), .ZN(n10595) );
  INV_X1 U9917 ( .A(P3_REG3_REG_13__SCAN_IN), .ZN(n9235) );
  OAI21_X1 U9918 ( .B1(n11194), .B2(P3_REG2_REG_2__SCAN_IN), .A(n10753), .ZN(
        n11179) );
  AND2_X1 U9919 ( .A1(n10801), .A2(P3_REG1_REG_4__SCAN_IN), .ZN(n10785) );
  INV_X1 U9920 ( .A(P3_REG3_REG_16__SCAN_IN), .ZN(n13280) );
  NAND2_X1 U9921 ( .A1(n13540), .A2(n9729), .ZN(n9730) );
  INV_X1 U9922 ( .A(n13574), .ZN(n9722) );
  INV_X1 U9923 ( .A(n13706), .ZN(n9715) );
  INV_X1 U9924 ( .A(n11000), .ZN(n9696) );
  INV_X1 U9925 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n9487) );
  INV_X1 U9926 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n9370) );
  INV_X1 U9927 ( .A(P3_IR_REG_5__SCAN_IN), .ZN(n9003) );
  AND2_X1 U9928 ( .A1(n8610), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n8628) );
  INV_X1 U9929 ( .A(n14262), .ZN(n8889) );
  INV_X1 U9930 ( .A(n13134), .ZN(n8908) );
  INV_X1 U9931 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n8196) );
  NOR2_X1 U9932 ( .A1(n14923), .A2(n15141), .ZN(n12530) );
  INV_X1 U9933 ( .A(n8806), .ZN(n8807) );
  NAND2_X1 U9934 ( .A1(n13184), .A2(n13355), .ZN(n13185) );
  AND2_X1 U9935 ( .A1(n9280), .A2(n13280), .ZN(n9298) );
  OR2_X1 U9936 ( .A1(n9249), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n9264) );
  NAND2_X1 U9937 ( .A1(n9362), .A2(n9361), .ZN(n9376) );
  OR2_X1 U9938 ( .A1(n9425), .A2(P3_REG3_REG_26__SCAN_IN), .ZN(n9438) );
  OR2_X1 U9939 ( .A1(n15304), .A2(n9452), .ZN(n13539) );
  NAND2_X1 U9940 ( .A1(P2_DATAO_REG_30__SCAN_IN), .A2(n9487), .ZN(n9488) );
  AND2_X1 U9941 ( .A1(n10002), .A2(P2_DATAO_REG_6__SCAN_IN), .ZN(n9128) );
  AND2_X1 U9942 ( .A1(n8188), .A2(n8187), .ZN(n8793) );
  OAI22_X1 U9943 ( .A1(n8947), .A2(n13913), .B1(n14022), .B2(n8946), .ZN(n8948) );
  NAND2_X1 U9944 ( .A1(n8974), .A2(n13977), .ZN(n8975) );
  AND2_X1 U9945 ( .A1(n10075), .A2(n8875), .ZN(n13952) );
  OR2_X1 U9946 ( .A1(n15620), .A2(n8860), .ZN(n8865) );
  NAND2_X1 U9947 ( .A1(n14090), .A2(n8889), .ZN(n14091) );
  XNOR2_X1 U9948 ( .A(n12874), .B(n8886), .ZN(n11654) );
  INV_X1 U9949 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n8207) );
  INV_X1 U9950 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n11243) );
  INV_X1 U9951 ( .A(n11771), .ZN(n11767) );
  INV_X1 U9952 ( .A(n9897), .ZN(n9896) );
  OR2_X1 U9953 ( .A1(n15113), .A2(n14556), .ZN(n12573) );
  INV_X1 U9954 ( .A(n12530), .ZN(n14913) );
  NOR2_X1 U9955 ( .A1(n15043), .A2(n15032), .ZN(n15027) );
  OR2_X1 U9956 ( .A1(n11535), .A2(n12620), .ZN(n11483) );
  NOR2_X1 U9957 ( .A1(P1_IR_REG_27__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), .ZN(
        n9836) );
  NAND2_X1 U9958 ( .A1(n9799), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9800) );
  INV_X1 U9959 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n10004) );
  INV_X1 U9960 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n8234) );
  OR2_X1 U9961 ( .A1(n9386), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n9396) );
  NOR2_X1 U9962 ( .A1(n9331), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n9344) );
  NAND2_X1 U9963 ( .A1(n9298), .A2(n9297), .ZN(n9316) );
  NAND2_X1 U9964 ( .A1(n9155), .A2(n11335), .ZN(n9173) );
  AND2_X1 U9965 ( .A1(n9344), .A2(n9343), .ZN(n9362) );
  AND2_X1 U9966 ( .A1(n9431), .A2(n9430), .ZN(n13548) );
  INV_X1 U9967 ( .A(n11332), .ZN(n11445) );
  NOR2_X1 U9968 ( .A1(n11979), .A2(n11978), .ZN(n13376) );
  NOR2_X1 U9969 ( .A1(n9438), .A2(P3_REG3_REG_27__SCAN_IN), .ZN(n9451) );
  AND2_X1 U9970 ( .A1(n9610), .A2(n9615), .ZN(n13710) );
  AND2_X2 U9971 ( .A1(n9562), .A2(n9566), .ZN(n11426) );
  AND2_X1 U9972 ( .A1(n10931), .A2(n10930), .ZN(n10932) );
  OR2_X1 U9973 ( .A1(n6678), .A2(n13845), .ZN(n9436) );
  INV_X1 U9974 ( .A(n15722), .ZN(n13691) );
  NAND2_X1 U9975 ( .A1(n15232), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n9471) );
  NAND2_X1 U9976 ( .A1(P1_DATAO_REG_18__SCAN_IN), .A2(n11262), .ZN(n9324) );
  INV_X1 U9977 ( .A(P3_IR_REG_9__SCAN_IN), .ZN(n9166) );
  NAND2_X1 U9978 ( .A1(n9031), .A2(n9049), .ZN(n9061) );
  INV_X1 U9979 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n12132) );
  XNOR2_X1 U9980 ( .A(n8350), .B(n8349), .ZN(n10405) );
  NAND2_X1 U9981 ( .A1(n8185), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n8775) );
  INV_X1 U9982 ( .A(n13936), .ZN(n8675) );
  AND3_X1 U9983 ( .A1(n10134), .A2(n10133), .A3(n10132), .ZN(n14023) );
  OR2_X1 U9984 ( .A1(n8665), .A2(n13942), .ZN(n8684) );
  OR2_X1 U9985 ( .A1(n10102), .A2(n13167), .ZN(n14009) );
  INV_X1 U9986 ( .A(n8948), .ZN(n8949) );
  INV_X1 U9987 ( .A(n14152), .ZN(n14176) );
  CLKBUF_X1 U9988 ( .A(n11654), .Z(n13121) );
  INV_X1 U9989 ( .A(n8951), .ZN(n8993) );
  OR2_X1 U9990 ( .A1(n8995), .A2(n8994), .ZN(n8952) );
  INV_X1 U9991 ( .A(n13146), .ZN(n14089) );
  INV_X1 U9992 ( .A(n13968), .ZN(n13916) );
  INV_X1 U9993 ( .A(n12109), .ZN(n12186) );
  AND2_X1 U9994 ( .A1(n8937), .A2(n13162), .ZN(n14220) );
  OR3_X1 U9995 ( .A1(n12322), .A2(n14395), .A3(n12388), .ZN(n9787) );
  NAND2_X1 U9996 ( .A1(n11347), .A2(n11349), .ZN(n11350) );
  INV_X1 U9997 ( .A(n12473), .ZN(n12472) );
  AND2_X1 U9998 ( .A1(n12310), .A2(n12309), .ZN(n12311) );
  NOR3_X1 U9999 ( .A1(n15391), .A2(n15390), .A3(n15389), .ZN(n15388) );
  XNOR2_X1 U10000 ( .A(n9896), .B(n9898), .ZN(n10659) );
  AND2_X1 U10001 ( .A1(n12507), .A2(n12521), .ZN(n14869) );
  INV_X1 U10002 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n14759) );
  INV_X1 U10003 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n10190) );
  NAND2_X1 U10004 ( .A1(n10189), .A2(n10186), .ZN(n10193) );
  OR3_X1 U10005 ( .A1(n14987), .A2(n14986), .A3(n15488), .ZN(n15172) );
  NAND2_X1 U10006 ( .A1(n9933), .A2(n9921), .ZN(n15495) );
  OR2_X1 U10007 ( .A1(n11210), .A2(n15048), .ZN(n11584) );
  INV_X1 U10008 ( .A(n15002), .ZN(n15091) );
  INV_X1 U10009 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n9992) );
  INV_X1 U10010 ( .A(P3_ADDR_REG_6__SCAN_IN), .ZN(n7761) );
  INV_X1 U10011 ( .A(n13346), .ZN(n13281) );
  AND2_X1 U10012 ( .A1(n10515), .A2(n10514), .ZN(n13337) );
  NAND2_X1 U10013 ( .A1(n9403), .A2(n9402), .ZN(n13603) );
  INV_X1 U10014 ( .A(n9689), .ZN(n10750) );
  INV_X1 U10015 ( .A(n13521), .ZN(n15699) );
  AND2_X1 U10016 ( .A1(n9451), .A2(n8142), .ZN(n15304) );
  AND2_X1 U10017 ( .A1(n9621), .A2(n9620), .ZN(n13677) );
  INV_X1 U10018 ( .A(n13694), .ZN(n15717) );
  AND3_X1 U10019 ( .A1(n15715), .A2(n10934), .A3(n15765), .ZN(n15709) );
  AND2_X1 U10020 ( .A1(n15733), .A2(n11216), .ZN(n13561) );
  AND2_X1 U10021 ( .A1(n15303), .A2(n15302), .ZN(n15313) );
  NAND2_X1 U10022 ( .A1(n9768), .A2(n11171), .ZN(n15758) );
  INV_X1 U10023 ( .A(n15758), .ZN(n15765) );
  OR2_X1 U10024 ( .A1(n13554), .A2(n15745), .ZN(n15316) );
  AND2_X1 U10025 ( .A1(n15715), .A2(n9768), .ZN(n15745) );
  OR2_X1 U10026 ( .A1(n8815), .A2(n8877), .ZN(n14032) );
  INV_X1 U10027 ( .A(n10131), .ZN(n8945) );
  INV_X1 U10028 ( .A(n14009), .ZN(n15609) );
  OAI21_X1 U10029 ( .B1(n10908), .B2(n8960), .A(n8959), .ZN(n11104) );
  INV_X1 U10030 ( .A(n14220), .ZN(n15617) );
  NAND2_X1 U10031 ( .A1(n15635), .A2(n8866), .ZN(n15621) );
  AND2_X1 U10032 ( .A1(n15688), .A2(n15672), .ZN(n14313) );
  AND2_X1 U10033 ( .A1(n8996), .A2(n8995), .ZN(n11064) );
  AND2_X1 U10034 ( .A1(n8420), .A2(n8456), .ZN(n10296) );
  XNOR2_X1 U10035 ( .A(n9811), .B(n9810), .ZN(n10183) );
  INV_X1 U10036 ( .A(n14683), .ZN(n15397) );
  NAND2_X1 U10037 ( .A1(n10184), .A2(n14721), .ZN(n15069) );
  AND3_X1 U10038 ( .A1(n12433), .A2(n12432), .A3(n12431), .ZN(n14572) );
  NOR2_X1 U10039 ( .A1(n10529), .A2(n10528), .ZN(n15022) );
  INV_X1 U10040 ( .A(n15468), .ZN(n14833) );
  INV_X1 U10041 ( .A(n15476), .ZN(n14819) );
  NAND2_X1 U10042 ( .A1(n12527), .A2(n12526), .ZN(n12528) );
  NAND2_X1 U10043 ( .A1(n10698), .A2(n10697), .ZN(n15280) );
  INV_X1 U10044 ( .A(n14994), .ZN(n15293) );
  NAND2_X1 U10045 ( .A1(n12584), .A2(n15058), .ZN(n15093) );
  NAND2_X1 U10046 ( .A1(n9907), .A2(n10019), .ZN(n10711) );
  OR2_X1 U10047 ( .A1(n12593), .A2(n12783), .ZN(n15499) );
  NAND2_X1 U10048 ( .A1(n11584), .A2(n15499), .ZN(n15413) );
  INV_X1 U10049 ( .A(n10711), .ZN(n11201) );
  OR2_X1 U10050 ( .A1(n9906), .A2(n9905), .ZN(n10019) );
  INV_X1 U10051 ( .A(n7818), .ZN(n7819) );
  AND2_X1 U10052 ( .A1(n10776), .A2(n10775), .ZN(n15698) );
  INV_X1 U10053 ( .A(n13337), .ZN(n13347) );
  AND2_X1 U10054 ( .A1(n9482), .A2(n9481), .ZN(n11102) );
  AND3_X1 U10055 ( .A1(n9366), .A2(n9365), .A3(n9364), .ZN(n13638) );
  INV_X1 U10056 ( .A(n10860), .ZN(n13358) );
  INV_X1 U10057 ( .A(n13529), .ZN(n15692) );
  OR2_X1 U10058 ( .A1(n10773), .A2(n13517), .ZN(n15693) );
  INV_X1 U10059 ( .A(n13716), .ZN(n13688) );
  NAND2_X1 U10060 ( .A1(n15784), .A2(n15765), .ZN(n13777) );
  INV_X1 U10061 ( .A(n15784), .ZN(n15782) );
  AND2_X1 U10062 ( .A1(n9783), .A2(n9782), .ZN(n15773) );
  AND2_X1 U10063 ( .A1(n10745), .A2(P3_STATE_REG_SCAN_IN), .ZN(n13826) );
  INV_X1 U10064 ( .A(n9748), .ZN(n13848) );
  INV_X1 U10065 ( .A(SI_16_), .ZN(n10250) );
  INV_X1 U10066 ( .A(SI_11_), .ZN(n9984) );
  INV_X1 U10067 ( .A(n10809), .ZN(n10869) );
  NAND2_X1 U10068 ( .A1(n8876), .A2(n13166), .ZN(n13953) );
  OR2_X1 U10069 ( .A1(n8655), .A2(n8654), .ZN(n13972) );
  INV_X1 U10070 ( .A(n15603), .ZN(n10350) );
  NAND2_X1 U10071 ( .A1(n14226), .A2(n11070), .ZN(n14157) );
  AND2_X1 U10072 ( .A1(n15623), .A2(n11130), .ZN(n14234) );
  INV_X1 U10073 ( .A(n14160), .ZN(n14213) );
  AND4_X1 U10074 ( .A1(n15668), .A2(n15667), .A3(n15666), .A4(n15665), .ZN(
        n15686) );
  OR2_X1 U10075 ( .A1(n15629), .A2(n15628), .ZN(n15630) );
  INV_X1 U10076 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n14394) );
  INV_X1 U10077 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n10352) );
  NAND2_X1 U10078 ( .A1(n10183), .A2(P1_STATE_REG_SCAN_IN), .ZN(n12840) );
  INV_X1 U10079 ( .A(n14448), .ZN(n15173) );
  INV_X1 U10080 ( .A(n15154), .ZN(n14946) );
  INV_X1 U10081 ( .A(n14516), .ZN(n15125) );
  NAND4_X1 U10082 ( .A1(n12511), .A2(n12510), .A3(n12509), .A4(n12508), .ZN(
        n14688) );
  OAI21_X1 U10083 ( .B1(n14956), .B2(n12451), .A(n12445), .ZN(n14969) );
  INV_X1 U10084 ( .A(n14637), .ZN(n14696) );
  INV_X1 U10085 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n15462) );
  INV_X1 U10086 ( .A(n15457), .ZN(n15472) );
  NAND2_X1 U10087 ( .A1(n11202), .A2(n12593), .ZN(n14994) );
  NAND2_X1 U10088 ( .A1(n15093), .A2(n11211), .ZN(n15063) );
  OR2_X1 U10089 ( .A1(n10712), .A2(n10711), .ZN(n15534) );
  AND2_X1 U10090 ( .A1(n15515), .A2(n15514), .ZN(n15533) );
  OR2_X1 U10091 ( .A1(n10712), .A2(n11201), .ZN(n15524) );
  INV_X1 U10092 ( .A(n12840), .ZN(n10024) );
  INV_X1 U10093 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n11316) );
  INV_X1 U10094 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n10650) );
  XNOR2_X1 U10095 ( .A(n8177), .B(n8176), .ZN(n8178) );
  NOR2_X1 U10096 ( .A1(n10079), .A2(P2_U3088), .ZN(P2_U3947) );
  NOR2_X2 U10097 ( .A1(n9928), .A2(n12840), .ZN(P1_U4016) );
  INV_X1 U10098 ( .A(P3_ADDR_REG_15__SCAN_IN), .ZN(n13415) );
  INV_X1 U10099 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n15477) );
  NOR2_X1 U10100 ( .A1(P3_ADDR_REG_15__SCAN_IN), .A2(n15477), .ZN(n7774) );
  INV_X1 U10101 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n10613) );
  XOR2_X1 U10102 ( .A(P3_ADDR_REG_14__SCAN_IN), .B(n10613), .Z(n7791) );
  INV_X1 U10103 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n7792) );
  INV_X1 U10104 ( .A(P3_ADDR_REG_12__SCAN_IN), .ZN(n7771) );
  XOR2_X1 U10105 ( .A(P1_ADDR_REG_12__SCAN_IN), .B(n7771), .Z(n7795) );
  INV_X1 U10106 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n14792) );
  XNOR2_X1 U10107 ( .A(n14792), .B(n8083), .ZN(n7799) );
  XOR2_X1 U10108 ( .A(n10190), .B(P3_ADDR_REG_8__SCAN_IN), .Z(n7801) );
  XOR2_X1 U10109 ( .A(P1_ADDR_REG_6__SCAN_IN), .B(n7761), .Z(n7823) );
  XOR2_X1 U10110 ( .A(P1_ADDR_REG_2__SCAN_IN), .B(n8106), .Z(n7806) );
  NOR2_X1 U10111 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(n8141), .ZN(n7810) );
  NAND2_X1 U10112 ( .A1(n7808), .A2(n7810), .ZN(n7750) );
  NAND2_X1 U10113 ( .A1(n7806), .A2(n7807), .ZN(n7751) );
  NAND2_X1 U10114 ( .A1(P3_ADDR_REG_3__SCAN_IN), .A2(n7752), .ZN(n7754) );
  XNOR2_X1 U10115 ( .A(n8121), .B(n7752), .ZN(n7805) );
  NAND2_X1 U10116 ( .A1(n7805), .A2(n7804), .ZN(n7753) );
  NAND2_X1 U10117 ( .A1(n7754), .A2(n7753), .ZN(n7755) );
  NAND2_X1 U10118 ( .A1(P3_ADDR_REG_4__SCAN_IN), .A2(n7755), .ZN(n7756) );
  NAND2_X1 U10119 ( .A1(P3_ADDR_REG_5__SCAN_IN), .A2(n7757), .ZN(n7759) );
  NAND2_X1 U10120 ( .A1(n7817), .A2(n14759), .ZN(n7758) );
  NAND2_X1 U10121 ( .A1(n7759), .A2(n7758), .ZN(n7824) );
  NAND2_X1 U10122 ( .A1(n7823), .A2(n7824), .ZN(n7760) );
  NAND2_X1 U10123 ( .A1(P3_ADDR_REG_7__SCAN_IN), .A2(n7762), .ZN(n7764) );
  XOR2_X1 U10124 ( .A(P3_ADDR_REG_7__SCAN_IN), .B(n7762), .Z(n7828) );
  INV_X1 U10125 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n7827) );
  NAND2_X1 U10126 ( .A1(n7828), .A2(n7827), .ZN(n7763) );
  NAND2_X1 U10127 ( .A1(n7764), .A2(n7763), .ZN(n7802) );
  NAND2_X1 U10128 ( .A1(n7801), .A2(n7802), .ZN(n7765) );
  NAND2_X1 U10129 ( .A1(n7799), .A2(n7800), .ZN(n7766) );
  INV_X1 U10130 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n10465) );
  INV_X1 U10131 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n10425) );
  XNOR2_X1 U10132 ( .A(n10425), .B(n11904), .ZN(n7797) );
  NAND2_X1 U10133 ( .A1(n7798), .A2(n7797), .ZN(n7769) );
  NAND2_X1 U10134 ( .A1(n7795), .A2(n7796), .ZN(n7770) );
  INV_X1 U10135 ( .A(P3_ADDR_REG_13__SCAN_IN), .ZN(n13364) );
  NAND2_X1 U10136 ( .A1(P1_ADDR_REG_13__SCAN_IN), .A2(n13364), .ZN(n7772) );
  NAND2_X1 U10137 ( .A1(n7791), .A2(n7790), .ZN(n7773) );
  OAI22_X1 U10138 ( .A1(P1_ADDR_REG_15__SCAN_IN), .A2(n13415), .B1(n7774), 
        .B2(n7788), .ZN(n7775) );
  INV_X1 U10139 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n7776) );
  NOR2_X1 U10140 ( .A1(n7775), .A2(n7776), .ZN(n7778) );
  XNOR2_X1 U10141 ( .A(n7776), .B(n7775), .ZN(n7785) );
  NOR2_X1 U10142 ( .A1(P3_ADDR_REG_16__SCAN_IN), .A2(n7785), .ZN(n7777) );
  NOR2_X1 U10143 ( .A1(n7778), .A2(n7777), .ZN(n7780) );
  INV_X1 U10144 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n7779) );
  NAND2_X1 U10145 ( .A1(n7780), .A2(n7779), .ZN(n7782) );
  INV_X1 U10146 ( .A(P3_ADDR_REG_17__SCAN_IN), .ZN(n13475) );
  XOR2_X1 U10147 ( .A(P1_ADDR_REG_17__SCAN_IN), .B(n7780), .Z(n7784) );
  OR2_X1 U10148 ( .A1(n13475), .A2(n7784), .ZN(n7781) );
  NAND2_X1 U10149 ( .A1(n7782), .A2(n7781), .ZN(n7841) );
  INV_X1 U10150 ( .A(P3_ADDR_REG_18__SCAN_IN), .ZN(n13491) );
  NOR2_X1 U10151 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(n13491), .ZN(n7783) );
  AOI21_X1 U10152 ( .B1(P1_ADDR_REG_18__SCAN_IN), .B2(n13491), .A(n7783), .ZN(
        n7842) );
  XOR2_X1 U10153 ( .A(n7841), .B(n7842), .Z(n15248) );
  XOR2_X1 U10154 ( .A(n13475), .B(n7784), .Z(n15299) );
  INV_X1 U10155 ( .A(P3_ADDR_REG_16__SCAN_IN), .ZN(n7786) );
  XOR2_X1 U10156 ( .A(n7786), .B(n7785), .Z(n15442) );
  NOR2_X1 U10157 ( .A1(P1_ADDR_REG_15__SCAN_IN), .A2(n13415), .ZN(n7787) );
  AOI21_X1 U10158 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(n13415), .A(n7787), .ZN(
        n7789) );
  XNOR2_X1 U10159 ( .A(n7789), .B(n7788), .ZN(n15437) );
  XNOR2_X1 U10160 ( .A(n7791), .B(n7790), .ZN(n15434) );
  XNOR2_X1 U10161 ( .A(n7792), .B(P3_ADDR_REG_13__SCAN_IN), .ZN(n7793) );
  XNOR2_X1 U10162 ( .A(n7794), .B(n7793), .ZN(n15430) );
  XNOR2_X1 U10163 ( .A(n7796), .B(n7795), .ZN(n7837) );
  XOR2_X1 U10164 ( .A(n7798), .B(n7797), .Z(n15421) );
  XOR2_X1 U10165 ( .A(n7800), .B(n7799), .Z(n15263) );
  XOR2_X1 U10166 ( .A(n7802), .B(n7801), .Z(n7831) );
  XNOR2_X1 U10167 ( .A(n15462), .B(n7803), .ZN(n7815) );
  AND2_X1 U10168 ( .A1(n7815), .A2(P2_ADDR_REG_4__SCAN_IN), .ZN(n7816) );
  XOR2_X1 U10169 ( .A(n7805), .B(n7804), .Z(n15797) );
  XOR2_X1 U10170 ( .A(n7807), .B(n7806), .Z(n15253) );
  INV_X1 U10171 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n7809) );
  AOI21_X1 U10172 ( .B1(n8141), .B2(P1_ADDR_REG_0__SCAN_IN), .A(n7810), .ZN(
        n7811) );
  INV_X1 U10173 ( .A(n7811), .ZN(n15791) );
  NAND2_X1 U10174 ( .A1(P2_ADDR_REG_0__SCAN_IN), .A2(n15791), .ZN(n15801) );
  NOR2_X1 U10175 ( .A1(n15253), .A2(n6693), .ZN(n7813) );
  NAND2_X1 U10176 ( .A1(n15253), .A2(n6693), .ZN(n15252) );
  OAI21_X1 U10177 ( .B1(P2_ADDR_REG_2__SCAN_IN), .B2(n7813), .A(n15252), .ZN(
        n15796) );
  NAND2_X1 U10178 ( .A1(n15797), .A2(n15796), .ZN(n7814) );
  NOR2_X1 U10179 ( .A1(n15797), .A2(n15796), .ZN(n15795) );
  AOI21_X1 U10180 ( .B1(P2_ADDR_REG_3__SCAN_IN), .B2(n7814), .A(n15795), .ZN(
        n15787) );
  XNOR2_X1 U10181 ( .A(P2_ADDR_REG_4__SCAN_IN), .B(n7815), .ZN(n15786) );
  NOR2_X1 U10182 ( .A1(n15787), .A2(n15786), .ZN(n15785) );
  NOR2_X1 U10183 ( .A1(n7816), .A2(n15785), .ZN(n7820) );
  NAND2_X1 U10184 ( .A1(n7820), .A2(n7818), .ZN(n7821) );
  INV_X1 U10185 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n15789) );
  INV_X1 U10186 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n7822) );
  XOR2_X1 U10187 ( .A(n7824), .B(n7823), .Z(n15257) );
  INV_X1 U10188 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n7826) );
  NAND2_X1 U10189 ( .A1(n7829), .A2(n7826), .ZN(n7830) );
  XOR2_X1 U10190 ( .A(n7828), .B(n7827), .Z(n15794) );
  NAND2_X1 U10191 ( .A1(n15794), .A2(n15793), .ZN(n15792) );
  NOR2_X1 U10192 ( .A1(n7831), .A2(n7832), .ZN(n7833) );
  INV_X1 U10193 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n15259) );
  INV_X1 U10194 ( .A(P3_ADDR_REG_10__SCAN_IN), .ZN(n11461) );
  NOR2_X1 U10195 ( .A1(n7835), .A2(n7834), .ZN(n7836) );
  XNOR2_X1 U10196 ( .A(n11461), .B(n7836), .ZN(n15267) );
  INV_X1 U10197 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n15567) );
  NAND2_X1 U10198 ( .A1(n6718), .A2(n7837), .ZN(n15427) );
  NOR2_X1 U10199 ( .A1(n15434), .A2(n15433), .ZN(n7838) );
  NAND2_X1 U10200 ( .A1(n15434), .A2(n15433), .ZN(n15432) );
  NAND2_X1 U10201 ( .A1(n15299), .A2(n15298), .ZN(n7839) );
  NOR2_X1 U10202 ( .A1(n15299), .A2(n15298), .ZN(n15297) );
  XNOR2_X1 U10203 ( .A(n8232), .B(P2_ADDR_REG_19__SCAN_IN), .ZN(n7840) );
  NAND2_X1 U10204 ( .A1(n7842), .A2(n7841), .ZN(n7843) );
  OAI21_X1 U10205 ( .B1(n13491), .B2(P1_ADDR_REG_18__SCAN_IN), .A(n7843), .ZN(
        n8177) );
  OAI22_X1 U10206 ( .A1(SI_24_), .A2(keyinput_g8), .B1(SI_21_), .B2(
        keyinput_g11), .ZN(n7844) );
  AOI221_X1 U10207 ( .B1(SI_24_), .B2(keyinput_g8), .C1(keyinput_g11), .C2(
        SI_21_), .A(n7844), .ZN(n7851) );
  OAI22_X1 U10208 ( .A1(SI_3_), .A2(keyinput_g29), .B1(P3_REG3_REG_0__SCAN_IN), 
        .B2(keyinput_g54), .ZN(n7845) );
  AOI221_X1 U10209 ( .B1(SI_3_), .B2(keyinput_g29), .C1(keyinput_g54), .C2(
        P3_REG3_REG_0__SCAN_IN), .A(n7845), .ZN(n7850) );
  OAI22_X1 U10210 ( .A1(P3_REG3_REG_1__SCAN_IN), .A2(keyinput_g44), .B1(
        P3_ADDR_REG_7__SCAN_IN), .B2(keyinput_g104), .ZN(n7846) );
  AOI221_X1 U10211 ( .B1(P3_REG3_REG_1__SCAN_IN), .B2(keyinput_g44), .C1(
        keyinput_g104), .C2(P3_ADDR_REG_7__SCAN_IN), .A(n7846), .ZN(n7849) );
  OAI22_X1 U10212 ( .A1(P3_REG3_REG_16__SCAN_IN), .A2(keyinput_g48), .B1(
        P3_DATAO_REG_12__SCAN_IN), .B2(keyinput_g84), .ZN(n7847) );
  AOI221_X1 U10213 ( .B1(P3_REG3_REG_16__SCAN_IN), .B2(keyinput_g48), .C1(
        keyinput_g84), .C2(P3_DATAO_REG_12__SCAN_IN), .A(n7847), .ZN(n7848) );
  NAND4_X1 U10214 ( .A1(n7851), .A2(n7850), .A3(n7849), .A4(n7848), .ZN(n7879)
         );
  OAI22_X1 U10215 ( .A1(P3_REG3_REG_13__SCAN_IN), .A2(keyinput_g56), .B1(
        keyinput_g0), .B2(P3_WR_REG_SCAN_IN), .ZN(n7852) );
  AOI221_X1 U10216 ( .B1(P3_REG3_REG_13__SCAN_IN), .B2(keyinput_g56), .C1(
        P3_WR_REG_SCAN_IN), .C2(keyinput_g0), .A(n7852), .ZN(n7859) );
  OAI22_X1 U10217 ( .A1(SI_19_), .A2(keyinput_g13), .B1(keyinput_g116), .B2(
        P1_IR_REG_9__SCAN_IN), .ZN(n7853) );
  AOI221_X1 U10218 ( .B1(SI_19_), .B2(keyinput_g13), .C1(P1_IR_REG_9__SCAN_IN), 
        .C2(keyinput_g116), .A(n7853), .ZN(n7858) );
  OAI22_X1 U10219 ( .A1(P3_REG3_REG_18__SCAN_IN), .A2(keyinput_g60), .B1(
        SI_26_), .B2(keyinput_g6), .ZN(n7854) );
  AOI221_X1 U10220 ( .B1(P3_REG3_REG_18__SCAN_IN), .B2(keyinput_g60), .C1(
        keyinput_g6), .C2(SI_26_), .A(n7854), .ZN(n7857) );
  OAI22_X1 U10221 ( .A1(SI_30_), .A2(keyinput_g2), .B1(SI_25_), .B2(
        keyinput_g7), .ZN(n7855) );
  AOI221_X1 U10222 ( .B1(SI_30_), .B2(keyinput_g2), .C1(keyinput_g7), .C2(
        SI_25_), .A(n7855), .ZN(n7856) );
  NAND4_X1 U10223 ( .A1(n7859), .A2(n7858), .A3(n7857), .A4(n7856), .ZN(n7878)
         );
  OAI22_X1 U10224 ( .A1(P1_IR_REG_18__SCAN_IN), .A2(keyinput_g125), .B1(
        keyinput_g75), .B2(P3_DATAO_REG_21__SCAN_IN), .ZN(n7860) );
  AOI221_X1 U10225 ( .B1(P1_IR_REG_18__SCAN_IN), .B2(keyinput_g125), .C1(
        P3_DATAO_REG_21__SCAN_IN), .C2(keyinput_g75), .A(n7860), .ZN(n7867) );
  OAI22_X1 U10226 ( .A1(P3_REG3_REG_26__SCAN_IN), .A2(keyinput_g62), .B1(
        keyinput_g4), .B2(SI_28_), .ZN(n7861) );
  AOI221_X1 U10227 ( .B1(P3_REG3_REG_26__SCAN_IN), .B2(keyinput_g62), .C1(
        SI_28_), .C2(keyinput_g4), .A(n7861), .ZN(n7866) );
  OAI22_X1 U10228 ( .A1(SI_29_), .A2(keyinput_g3), .B1(keyinput_g114), .B2(
        P1_IR_REG_7__SCAN_IN), .ZN(n7862) );
  AOI221_X1 U10229 ( .B1(SI_29_), .B2(keyinput_g3), .C1(P1_IR_REG_7__SCAN_IN), 
        .C2(keyinput_g114), .A(n7862), .ZN(n7865) );
  OAI22_X1 U10230 ( .A1(P1_IR_REG_2__SCAN_IN), .A2(keyinput_g109), .B1(
        keyinput_g81), .B2(P3_DATAO_REG_15__SCAN_IN), .ZN(n7863) );
  AOI221_X1 U10231 ( .B1(P1_IR_REG_2__SCAN_IN), .B2(keyinput_g109), .C1(
        P3_DATAO_REG_15__SCAN_IN), .C2(keyinput_g81), .A(n7863), .ZN(n7864) );
  NAND4_X1 U10232 ( .A1(n7867), .A2(n7866), .A3(n7865), .A4(n7864), .ZN(n7877)
         );
  OAI22_X1 U10233 ( .A1(SI_2_), .A2(keyinput_g30), .B1(keyinput_g90), .B2(
        P3_DATAO_REG_6__SCAN_IN), .ZN(n7868) );
  AOI221_X1 U10234 ( .B1(SI_2_), .B2(keyinput_g30), .C1(
        P3_DATAO_REG_6__SCAN_IN), .C2(keyinput_g90), .A(n7868), .ZN(n7875) );
  OAI22_X1 U10235 ( .A1(SI_27_), .A2(keyinput_g5), .B1(SI_15_), .B2(
        keyinput_g17), .ZN(n7869) );
  AOI221_X1 U10236 ( .B1(SI_27_), .B2(keyinput_g5), .C1(keyinput_g17), .C2(
        SI_15_), .A(n7869), .ZN(n7874) );
  OAI22_X1 U10237 ( .A1(SI_20_), .A2(keyinput_g12), .B1(keyinput_g86), .B2(
        P3_DATAO_REG_10__SCAN_IN), .ZN(n7870) );
  AOI221_X1 U10238 ( .B1(SI_20_), .B2(keyinput_g12), .C1(
        P3_DATAO_REG_10__SCAN_IN), .C2(keyinput_g86), .A(n7870), .ZN(n7873) );
  OAI22_X1 U10239 ( .A1(P3_STATE_REG_SCAN_IN), .A2(keyinput_g34), .B1(
        keyinput_g15), .B2(SI_17_), .ZN(n7871) );
  AOI221_X1 U10240 ( .B1(P3_STATE_REG_SCAN_IN), .B2(keyinput_g34), .C1(SI_17_), 
        .C2(keyinput_g15), .A(n7871), .ZN(n7872) );
  NAND4_X1 U10241 ( .A1(n7875), .A2(n7874), .A3(n7873), .A4(n7872), .ZN(n7876)
         );
  NOR4_X1 U10242 ( .A1(n7879), .A2(n7878), .A3(n7877), .A4(n7876), .ZN(n8174)
         );
  OAI22_X1 U10243 ( .A1(P1_IR_REG_14__SCAN_IN), .A2(keyinput_g121), .B1(
        keyinput_g85), .B2(P3_DATAO_REG_11__SCAN_IN), .ZN(n7880) );
  AOI221_X1 U10244 ( .B1(P1_IR_REG_14__SCAN_IN), .B2(keyinput_g121), .C1(
        P3_DATAO_REG_11__SCAN_IN), .C2(keyinput_g85), .A(n7880), .ZN(n7887) );
  OAI22_X1 U10245 ( .A1(P3_REG3_REG_14__SCAN_IN), .A2(keyinput_g37), .B1(
        P1_IR_REG_12__SCAN_IN), .B2(keyinput_g119), .ZN(n7881) );
  AOI221_X1 U10246 ( .B1(P3_REG3_REG_14__SCAN_IN), .B2(keyinput_g37), .C1(
        keyinput_g119), .C2(P1_IR_REG_12__SCAN_IN), .A(n7881), .ZN(n7886) );
  OAI22_X1 U10247 ( .A1(P3_DATAO_REG_29__SCAN_IN), .A2(keyinput_g67), .B1(
        keyinput_g95), .B2(P3_DATAO_REG_1__SCAN_IN), .ZN(n7882) );
  AOI221_X1 U10248 ( .B1(P3_DATAO_REG_29__SCAN_IN), .B2(keyinput_g67), .C1(
        P3_DATAO_REG_1__SCAN_IN), .C2(keyinput_g95), .A(n7882), .ZN(n7885) );
  OAI22_X1 U10249 ( .A1(SI_0_), .A2(keyinput_g32), .B1(P1_IR_REG_1__SCAN_IN), 
        .B2(keyinput_g108), .ZN(n7883) );
  AOI221_X1 U10250 ( .B1(SI_0_), .B2(keyinput_g32), .C1(keyinput_g108), .C2(
        P1_IR_REG_1__SCAN_IN), .A(n7883), .ZN(n7884) );
  NAND4_X1 U10251 ( .A1(n7887), .A2(n7886), .A3(n7885), .A4(n7884), .ZN(n8000)
         );
  OAI22_X1 U10252 ( .A1(P3_REG3_REG_21__SCAN_IN), .A2(keyinput_g45), .B1(
        keyinput_g83), .B2(P3_DATAO_REG_13__SCAN_IN), .ZN(n7888) );
  AOI221_X1 U10253 ( .B1(P3_REG3_REG_21__SCAN_IN), .B2(keyinput_g45), .C1(
        P3_DATAO_REG_13__SCAN_IN), .C2(keyinput_g83), .A(n7888), .ZN(n7913) );
  INV_X1 U10254 ( .A(P3_DATAO_REG_16__SCAN_IN), .ZN(n10563) );
  OAI22_X1 U10255 ( .A1(P1_IR_REG_6__SCAN_IN), .A2(keyinput_g113), .B1(
        keyinput_g103), .B2(P3_ADDR_REG_6__SCAN_IN), .ZN(n7889) );
  AOI221_X1 U10256 ( .B1(P1_IR_REG_6__SCAN_IN), .B2(keyinput_g113), .C1(
        P3_ADDR_REG_6__SCAN_IN), .C2(keyinput_g103), .A(n7889), .ZN(n7892) );
  OAI22_X1 U10257 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(keyinput_g126), .B1(
        P3_ADDR_REG_5__SCAN_IN), .B2(keyinput_g102), .ZN(n7890) );
  AOI221_X1 U10258 ( .B1(P1_IR_REG_19__SCAN_IN), .B2(keyinput_g126), .C1(
        keyinput_g102), .C2(P3_ADDR_REG_5__SCAN_IN), .A(n7890), .ZN(n7891) );
  OAI211_X1 U10259 ( .C1(n10563), .C2(keyinput_g80), .A(n7892), .B(n7891), 
        .ZN(n7893) );
  AOI21_X1 U10260 ( .B1(n10563), .B2(keyinput_g80), .A(n7893), .ZN(n7912) );
  AOI22_X1 U10261 ( .A1(SI_1_), .A2(keyinput_g31), .B1(P3_REG3_REG_15__SCAN_IN), .B2(keyinput_g63), .ZN(n7894) );
  OAI221_X1 U10262 ( .B1(SI_1_), .B2(keyinput_g31), .C1(
        P3_REG3_REG_15__SCAN_IN), .C2(keyinput_g63), .A(n7894), .ZN(n7901) );
  AOI22_X1 U10263 ( .A1(P3_DATAO_REG_2__SCAN_IN), .A2(keyinput_g94), .B1(
        P3_DATAO_REG_30__SCAN_IN), .B2(keyinput_g66), .ZN(n7895) );
  OAI221_X1 U10264 ( .B1(P3_DATAO_REG_2__SCAN_IN), .B2(keyinput_g94), .C1(
        P3_DATAO_REG_30__SCAN_IN), .C2(keyinput_g66), .A(n7895), .ZN(n7900) );
  AOI22_X1 U10265 ( .A1(P3_DATAO_REG_19__SCAN_IN), .A2(keyinput_g77), .B1(
        P3_DATAO_REG_8__SCAN_IN), .B2(keyinput_g88), .ZN(n7896) );
  OAI221_X1 U10266 ( .B1(P3_DATAO_REG_19__SCAN_IN), .B2(keyinput_g77), .C1(
        P3_DATAO_REG_8__SCAN_IN), .C2(keyinput_g88), .A(n7896), .ZN(n7899) );
  AOI22_X1 U10267 ( .A1(P1_IR_REG_16__SCAN_IN), .A2(keyinput_g123), .B1(
        P3_REG3_REG_27__SCAN_IN), .B2(keyinput_g36), .ZN(n7897) );
  OAI221_X1 U10268 ( .B1(P1_IR_REG_16__SCAN_IN), .B2(keyinput_g123), .C1(
        P3_REG3_REG_27__SCAN_IN), .C2(keyinput_g36), .A(n7897), .ZN(n7898) );
  NOR4_X1 U10269 ( .A1(n7901), .A2(n7900), .A3(n7899), .A4(n7898), .ZN(n7911)
         );
  AOI22_X1 U10270 ( .A1(P3_DATAO_REG_17__SCAN_IN), .A2(keyinput_g79), .B1(
        P1_IR_REG_5__SCAN_IN), .B2(keyinput_g112), .ZN(n7902) );
  OAI221_X1 U10271 ( .B1(P3_DATAO_REG_17__SCAN_IN), .B2(keyinput_g79), .C1(
        P1_IR_REG_5__SCAN_IN), .C2(keyinput_g112), .A(n7902), .ZN(n7909) );
  AOI22_X1 U10272 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(keyinput_g127), .B1(
        P1_IR_REG_11__SCAN_IN), .B2(keyinput_g118), .ZN(n7903) );
  OAI221_X1 U10273 ( .B1(P1_IR_REG_20__SCAN_IN), .B2(keyinput_g127), .C1(
        P1_IR_REG_11__SCAN_IN), .C2(keyinput_g118), .A(n7903), .ZN(n7908) );
  AOI22_X1 U10274 ( .A1(P3_REG3_REG_17__SCAN_IN), .A2(keyinput_g50), .B1(
        P3_REG3_REG_20__SCAN_IN), .B2(keyinput_g55), .ZN(n7904) );
  OAI221_X1 U10275 ( .B1(P3_REG3_REG_17__SCAN_IN), .B2(keyinput_g50), .C1(
        P3_REG3_REG_20__SCAN_IN), .C2(keyinput_g55), .A(n7904), .ZN(n7907) );
  AOI22_X1 U10276 ( .A1(P1_IR_REG_15__SCAN_IN), .A2(keyinput_g122), .B1(
        P3_REG3_REG_10__SCAN_IN), .B2(keyinput_g39), .ZN(n7905) );
  OAI221_X1 U10277 ( .B1(P1_IR_REG_15__SCAN_IN), .B2(keyinput_g122), .C1(
        P3_REG3_REG_10__SCAN_IN), .C2(keyinput_g39), .A(n7905), .ZN(n7906) );
  NOR4_X1 U10278 ( .A1(n7909), .A2(n7908), .A3(n7907), .A4(n7906), .ZN(n7910)
         );
  NAND4_X1 U10279 ( .A1(n7913), .A2(n7912), .A3(n7911), .A4(n7910), .ZN(n7999)
         );
  INV_X1 U10280 ( .A(P3_DATAO_REG_0__SCAN_IN), .ZN(n10633) );
  INV_X1 U10281 ( .A(P3_DATAO_REG_5__SCAN_IN), .ZN(n10624) );
  AOI22_X1 U10282 ( .A1(n10633), .A2(keyinput_g96), .B1(n10624), .B2(
        keyinput_g91), .ZN(n7914) );
  OAI221_X1 U10283 ( .B1(n10633), .B2(keyinput_g96), .C1(n10624), .C2(
        keyinput_g91), .A(n7914), .ZN(n7916) );
  INV_X1 U10284 ( .A(P3_DATAO_REG_9__SCAN_IN), .ZN(n10643) );
  XNOR2_X1 U10285 ( .A(n10643), .B(keyinput_g87), .ZN(n7915) );
  NOR2_X1 U10286 ( .A1(n7916), .A2(n7915), .ZN(n7925) );
  INV_X1 U10287 ( .A(P3_DATAO_REG_3__SCAN_IN), .ZN(n10627) );
  INV_X1 U10288 ( .A(P3_REG3_REG_24__SCAN_IN), .ZN(n7918) );
  AOI22_X1 U10289 ( .A1(n10627), .A2(keyinput_g93), .B1(n7918), .B2(
        keyinput_g51), .ZN(n7917) );
  OAI221_X1 U10290 ( .B1(n10627), .B2(keyinput_g93), .C1(n7918), .C2(
        keyinput_g51), .A(n7917), .ZN(n7919) );
  INV_X1 U10291 ( .A(n7919), .ZN(n7924) );
  AOI22_X1 U10292 ( .A1(P3_RD_REG_SCAN_IN), .A2(keyinput_g33), .B1(
        P3_REG3_REG_3__SCAN_IN), .B2(keyinput_g40), .ZN(n7920) );
  OAI221_X1 U10293 ( .B1(P3_RD_REG_SCAN_IN), .B2(keyinput_g33), .C1(
        P3_REG3_REG_3__SCAN_IN), .C2(keyinput_g40), .A(n7920), .ZN(n7921) );
  INV_X1 U10294 ( .A(n7921), .ZN(n7923) );
  XNOR2_X1 U10295 ( .A(P1_IR_REG_4__SCAN_IN), .B(keyinput_g111), .ZN(n7922) );
  AND4_X1 U10296 ( .A1(n7925), .A2(n7924), .A3(n7923), .A4(n7922), .ZN(n7955)
         );
  INV_X1 U10297 ( .A(P3_REG3_REG_25__SCAN_IN), .ZN(n9409) );
  AOI22_X1 U10298 ( .A1(n9409), .A2(keyinput_g47), .B1(keyinput_g97), .B2(
        n8141), .ZN(n7926) );
  OAI221_X1 U10299 ( .B1(n9409), .B2(keyinput_g47), .C1(n8141), .C2(
        keyinput_g97), .A(n7926), .ZN(n7934) );
  INV_X1 U10300 ( .A(P3_DATAO_REG_26__SCAN_IN), .ZN(n11063) );
  INV_X1 U10301 ( .A(P3_REG3_REG_28__SCAN_IN), .ZN(n8142) );
  AOI22_X1 U10302 ( .A1(n11063), .A2(keyinput_g70), .B1(n8142), .B2(
        keyinput_g42), .ZN(n7927) );
  OAI221_X1 U10303 ( .B1(n11063), .B2(keyinput_g70), .C1(n8142), .C2(
        keyinput_g42), .A(n7927), .ZN(n7933) );
  INV_X1 U10304 ( .A(P3_REG3_REG_6__SCAN_IN), .ZN(n10798) );
  AOI22_X1 U10305 ( .A1(n10798), .A2(keyinput_g61), .B1(keyinput_g120), .B2(
        n10456), .ZN(n7928) );
  OAI221_X1 U10306 ( .B1(n10798), .B2(keyinput_g61), .C1(n10456), .C2(
        keyinput_g120), .A(n7928), .ZN(n7932) );
  XNOR2_X1 U10307 ( .A(SI_7_), .B(keyinput_g25), .ZN(n7930) );
  XNOR2_X1 U10308 ( .A(SI_9_), .B(keyinput_g23), .ZN(n7929) );
  NAND2_X1 U10309 ( .A1(n7930), .A2(n7929), .ZN(n7931) );
  NOR4_X1 U10310 ( .A1(n7934), .A2(n7933), .A3(n7932), .A4(n7931), .ZN(n7954)
         );
  INV_X1 U10311 ( .A(P3_REG3_REG_23__SCAN_IN), .ZN(n13236) );
  INV_X1 U10312 ( .A(P3_REG3_REG_7__SCAN_IN), .ZN(n10866) );
  AOI22_X1 U10313 ( .A1(n13236), .A2(keyinput_g38), .B1(keyinput_g35), .B2(
        n10866), .ZN(n7935) );
  OAI221_X1 U10314 ( .B1(n13236), .B2(keyinput_g38), .C1(n10866), .C2(
        keyinput_g35), .A(n7935), .ZN(n7943) );
  INV_X1 U10315 ( .A(P3_DATAO_REG_7__SCAN_IN), .ZN(n10641) );
  AOI22_X1 U10316 ( .A1(n7138), .A2(keyinput_g101), .B1(keyinput_g89), .B2(
        n10641), .ZN(n7936) );
  OAI221_X1 U10317 ( .B1(n7138), .B2(keyinput_g101), .C1(n10641), .C2(
        keyinput_g89), .A(n7936), .ZN(n7942) );
  XNOR2_X1 U10318 ( .A(SI_14_), .B(keyinput_g18), .ZN(n7940) );
  XNOR2_X1 U10319 ( .A(P1_IR_REG_0__SCAN_IN), .B(keyinput_g107), .ZN(n7939) );
  XNOR2_X1 U10320 ( .A(P1_IR_REG_10__SCAN_IN), .B(keyinput_g117), .ZN(n7938)
         );
  XNOR2_X1 U10321 ( .A(P1_IR_REG_3__SCAN_IN), .B(keyinput_g110), .ZN(n7937) );
  NAND4_X1 U10322 ( .A1(n7940), .A2(n7939), .A3(n7938), .A4(n7937), .ZN(n7941)
         );
  NOR3_X1 U10323 ( .A1(n7943), .A2(n7942), .A3(n7941), .ZN(n7953) );
  INV_X1 U10324 ( .A(P3_B_REG_SCAN_IN), .ZN(n9734) );
  AOI22_X1 U10325 ( .A1(n10889), .A2(keyinput_g49), .B1(keyinput_g64), .B2(
        n9734), .ZN(n7944) );
  OAI221_X1 U10326 ( .B1(n10889), .B2(keyinput_g49), .C1(n9734), .C2(
        keyinput_g64), .A(n7944), .ZN(n7951) );
  INV_X1 U10327 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n10030) );
  AOI22_X1 U10328 ( .A1(n10030), .A2(keyinput_g115), .B1(keyinput_g99), .B2(
        n8106), .ZN(n7945) );
  OAI221_X1 U10329 ( .B1(n10030), .B2(keyinput_g115), .C1(n8106), .C2(
        keyinput_g99), .A(n7945), .ZN(n7950) );
  INV_X1 U10330 ( .A(P3_DATAO_REG_28__SCAN_IN), .ZN(n11342) );
  AOI22_X1 U10331 ( .A1(n8083), .A2(keyinput_g106), .B1(keyinput_g68), .B2(
        n11342), .ZN(n7946) );
  OAI221_X1 U10332 ( .B1(n8083), .B2(keyinput_g106), .C1(n11342), .C2(
        keyinput_g68), .A(n7946), .ZN(n7949) );
  INV_X1 U10333 ( .A(P3_REG3_REG_9__SCAN_IN), .ZN(n11335) );
  INV_X1 U10334 ( .A(P3_DATAO_REG_27__SCAN_IN), .ZN(n11198) );
  AOI22_X1 U10335 ( .A1(n11335), .A2(keyinput_g53), .B1(keyinput_g69), .B2(
        n11198), .ZN(n7947) );
  OAI221_X1 U10336 ( .B1(n11335), .B2(keyinput_g53), .C1(n11198), .C2(
        keyinput_g69), .A(n7947), .ZN(n7948) );
  NOR4_X1 U10337 ( .A1(n7951), .A2(n7950), .A3(n7949), .A4(n7948), .ZN(n7952)
         );
  NAND4_X1 U10338 ( .A1(n7955), .A2(n7954), .A3(n7953), .A4(n7952), .ZN(n7998)
         );
  INV_X1 U10339 ( .A(P3_DATAO_REG_22__SCAN_IN), .ZN(n10646) );
  INV_X1 U10340 ( .A(P3_REG3_REG_11__SCAN_IN), .ZN(n11902) );
  AOI22_X1 U10341 ( .A1(n10646), .A2(keyinput_g74), .B1(n11902), .B2(
        keyinput_g58), .ZN(n7956) );
  OAI221_X1 U10342 ( .B1(n10646), .B2(keyinput_g74), .C1(n11902), .C2(
        keyinput_g58), .A(n7956), .ZN(n7964) );
  INV_X1 U10343 ( .A(P3_REG3_REG_22__SCAN_IN), .ZN(n13314) );
  AOI22_X1 U10344 ( .A1(n8121), .A2(keyinput_g100), .B1(n13314), .B2(
        keyinput_g57), .ZN(n7957) );
  OAI221_X1 U10345 ( .B1(n8121), .B2(keyinput_g100), .C1(n13314), .C2(
        keyinput_g57), .A(n7957), .ZN(n7963) );
  XNOR2_X1 U10346 ( .A(SI_11_), .B(keyinput_g21), .ZN(n7961) );
  XNOR2_X1 U10347 ( .A(P1_IR_REG_17__SCAN_IN), .B(keyinput_g124), .ZN(n7960)
         );
  XNOR2_X1 U10348 ( .A(SI_4_), .B(keyinput_g28), .ZN(n7959) );
  XNOR2_X1 U10349 ( .A(SI_6_), .B(keyinput_g26), .ZN(n7958) );
  NAND4_X1 U10350 ( .A1(n7961), .A2(n7960), .A3(n7959), .A4(n7958), .ZN(n7962)
         );
  NOR3_X1 U10351 ( .A1(n7964), .A2(n7963), .A3(n7962), .ZN(n7996) );
  INV_X1 U10352 ( .A(P3_REG3_REG_19__SCAN_IN), .ZN(n7966) );
  INV_X1 U10353 ( .A(P3_DATAO_REG_4__SCAN_IN), .ZN(n10629) );
  AOI22_X1 U10354 ( .A1(n7966), .A2(keyinput_g41), .B1(keyinput_g92), .B2(
        n10629), .ZN(n7965) );
  OAI221_X1 U10355 ( .B1(n7966), .B2(keyinput_g41), .C1(n10629), .C2(
        keyinput_g92), .A(n7965), .ZN(n7974) );
  INV_X1 U10356 ( .A(P3_DATAO_REG_24__SCAN_IN), .ZN(n10666) );
  INV_X1 U10357 ( .A(SI_22_), .ZN(n9373) );
  AOI22_X1 U10358 ( .A1(n10666), .A2(keyinput_g72), .B1(n9373), .B2(
        keyinput_g10), .ZN(n7967) );
  OAI221_X1 U10359 ( .B1(n10666), .B2(keyinput_g72), .C1(n9373), .C2(
        keyinput_g10), .A(n7967), .ZN(n7973) );
  INV_X1 U10360 ( .A(SI_18_), .ZN(n10522) );
  AOI22_X1 U10361 ( .A1(n10250), .A2(keyinput_g16), .B1(n10522), .B2(
        keyinput_g14), .ZN(n7968) );
  OAI221_X1 U10362 ( .B1(n10250), .B2(keyinput_g16), .C1(n10522), .C2(
        keyinput_g14), .A(n7968), .ZN(n7972) );
  XNOR2_X1 U10363 ( .A(SI_5_), .B(keyinput_g27), .ZN(n7970) );
  XNOR2_X1 U10364 ( .A(SI_13_), .B(keyinput_g19), .ZN(n7969) );
  NAND2_X1 U10365 ( .A1(n7970), .A2(n7969), .ZN(n7971) );
  NOR4_X1 U10366 ( .A1(n7974), .A2(n7973), .A3(n7972), .A4(n7971), .ZN(n7995)
         );
  INV_X1 U10367 ( .A(P3_DATAO_REG_14__SCAN_IN), .ZN(n10327) );
  INV_X1 U10368 ( .A(P3_DATAO_REG_18__SCAN_IN), .ZN(n10561) );
  AOI22_X1 U10369 ( .A1(n10327), .A2(keyinput_g82), .B1(n10561), .B2(
        keyinput_g78), .ZN(n7975) );
  OAI221_X1 U10370 ( .B1(n10327), .B2(keyinput_g82), .C1(n10561), .C2(
        keyinput_g78), .A(n7975), .ZN(n7983) );
  INV_X1 U10371 ( .A(P3_DATAO_REG_23__SCAN_IN), .ZN(n10648) );
  AOI22_X1 U10372 ( .A1(n10648), .A2(keyinput_g73), .B1(n10682), .B2(
        keyinput_g59), .ZN(n7976) );
  OAI221_X1 U10373 ( .B1(n10648), .B2(keyinput_g73), .C1(n10682), .C2(
        keyinput_g59), .A(n7976), .ZN(n7982) );
  INV_X1 U10374 ( .A(SI_31_), .ZN(n7978) );
  INV_X1 U10375 ( .A(SI_23_), .ZN(n11600) );
  AOI22_X1 U10376 ( .A1(n7978), .A2(keyinput_g1), .B1(keyinput_g9), .B2(n11600), .ZN(n7977) );
  OAI221_X1 U10377 ( .B1(n7978), .B2(keyinput_g1), .C1(n11600), .C2(
        keyinput_g9), .A(n7977), .ZN(n7981) );
  INV_X1 U10378 ( .A(P3_DATAO_REG_20__SCAN_IN), .ZN(n10637) );
  AOI22_X1 U10379 ( .A1(n10637), .A2(keyinput_g76), .B1(n8104), .B2(
        keyinput_g105), .ZN(n7979) );
  OAI221_X1 U10380 ( .B1(n10637), .B2(keyinput_g76), .C1(n8104), .C2(
        keyinput_g105), .A(n7979), .ZN(n7980) );
  NOR4_X1 U10381 ( .A1(n7983), .A2(n7982), .A3(n7981), .A4(n7980), .ZN(n7994)
         );
  INV_X1 U10382 ( .A(P3_DATAO_REG_25__SCAN_IN), .ZN(n10859) );
  INV_X1 U10383 ( .A(P3_REG3_REG_4__SCAN_IN), .ZN(n10777) );
  AOI22_X1 U10384 ( .A1(n10859), .A2(keyinput_g71), .B1(n10777), .B2(
        keyinput_g52), .ZN(n7984) );
  OAI221_X1 U10385 ( .B1(n10859), .B2(keyinput_g71), .C1(n10777), .C2(
        keyinput_g52), .A(n7984), .ZN(n7988) );
  INV_X1 U10386 ( .A(P3_REG3_REG_12__SCAN_IN), .ZN(n11988) );
  AOI22_X1 U10387 ( .A1(n10983), .A2(keyinput_g43), .B1(n11988), .B2(
        keyinput_g46), .ZN(n7985) );
  OAI221_X1 U10388 ( .B1(n10983), .B2(keyinput_g43), .C1(n11988), .C2(
        keyinput_g46), .A(n7985), .ZN(n7987) );
  XOR2_X1 U10389 ( .A(SI_8_), .B(keyinput_g24), .Z(n7986) );
  OR3_X1 U10390 ( .A1(n7988), .A2(n7987), .A3(n7986), .ZN(n7992) );
  AOI22_X1 U10391 ( .A1(n9999), .A2(keyinput_g20), .B1(keyinput_g98), .B2(
        n8102), .ZN(n7989) );
  OAI221_X1 U10392 ( .B1(n9999), .B2(keyinput_g20), .C1(n8102), .C2(
        keyinput_g98), .A(n7989), .ZN(n7991) );
  INV_X1 U10393 ( .A(P3_DATAO_REG_31__SCAN_IN), .ZN(n11173) );
  XNOR2_X1 U10394 ( .A(n11173), .B(keyinput_g65), .ZN(n7990) );
  NOR3_X1 U10395 ( .A1(n7992), .A2(n7991), .A3(n7990), .ZN(n7993) );
  NAND4_X1 U10396 ( .A1(n7996), .A2(n7995), .A3(n7994), .A4(n7993), .ZN(n7997)
         );
  NOR4_X1 U10397 ( .A1(n8000), .A2(n7999), .A3(n7998), .A4(n7997), .ZN(n8173)
         );
  OAI22_X1 U10398 ( .A1(keyinput_f78), .A2(P3_DATAO_REG_18__SCAN_IN), .B1(
        keyinput_f87), .B2(P3_DATAO_REG_9__SCAN_IN), .ZN(n8001) );
  AOI221_X1 U10399 ( .B1(keyinput_f78), .B2(P3_DATAO_REG_18__SCAN_IN), .C1(
        P3_DATAO_REG_9__SCAN_IN), .C2(keyinput_f87), .A(n8001), .ZN(n8008) );
  OAI22_X1 U10400 ( .A1(P3_REG3_REG_26__SCAN_IN), .A2(keyinput_f62), .B1(SI_5_), .B2(keyinput_f27), .ZN(n8002) );
  AOI221_X1 U10401 ( .B1(P3_REG3_REG_26__SCAN_IN), .B2(keyinput_f62), .C1(
        keyinput_f27), .C2(SI_5_), .A(n8002), .ZN(n8007) );
  OAI22_X1 U10402 ( .A1(P3_REG3_REG_18__SCAN_IN), .A2(keyinput_f60), .B1(
        keyinput_f118), .B2(P1_IR_REG_11__SCAN_IN), .ZN(n8003) );
  AOI221_X1 U10403 ( .B1(P3_REG3_REG_18__SCAN_IN), .B2(keyinput_f60), .C1(
        P1_IR_REG_11__SCAN_IN), .C2(keyinput_f118), .A(n8003), .ZN(n8006) );
  OAI22_X1 U10404 ( .A1(P3_REG3_REG_19__SCAN_IN), .A2(keyinput_f41), .B1(
        P1_IR_REG_2__SCAN_IN), .B2(keyinput_f109), .ZN(n8004) );
  AOI221_X1 U10405 ( .B1(P3_REG3_REG_19__SCAN_IN), .B2(keyinput_f41), .C1(
        keyinput_f109), .C2(P1_IR_REG_2__SCAN_IN), .A(n8004), .ZN(n8005) );
  NAND4_X1 U10406 ( .A1(n8008), .A2(n8007), .A3(n8006), .A4(n8005), .ZN(n8037)
         );
  OAI22_X1 U10407 ( .A1(SI_25_), .A2(keyinput_f7), .B1(keyinput_f127), .B2(
        P1_IR_REG_20__SCAN_IN), .ZN(n8009) );
  AOI221_X1 U10408 ( .B1(SI_25_), .B2(keyinput_f7), .C1(P1_IR_REG_20__SCAN_IN), 
        .C2(keyinput_f127), .A(n8009), .ZN(n8016) );
  OAI22_X1 U10409 ( .A1(keyinput_f80), .A2(P3_DATAO_REG_16__SCAN_IN), .B1(
        keyinput_f94), .B2(P3_DATAO_REG_2__SCAN_IN), .ZN(n8010) );
  AOI221_X1 U10410 ( .B1(keyinput_f80), .B2(P3_DATAO_REG_16__SCAN_IN), .C1(
        P3_DATAO_REG_2__SCAN_IN), .C2(keyinput_f94), .A(n8010), .ZN(n8015) );
  OAI22_X1 U10411 ( .A1(P3_REG3_REG_24__SCAN_IN), .A2(keyinput_f51), .B1(
        keyinput_f102), .B2(P3_ADDR_REG_5__SCAN_IN), .ZN(n8011) );
  AOI221_X1 U10412 ( .B1(P3_REG3_REG_24__SCAN_IN), .B2(keyinput_f51), .C1(
        P3_ADDR_REG_5__SCAN_IN), .C2(keyinput_f102), .A(n8011), .ZN(n8014) );
  OAI22_X1 U10413 ( .A1(P1_IR_REG_12__SCAN_IN), .A2(keyinput_f119), .B1(
        keyinput_f116), .B2(P1_IR_REG_9__SCAN_IN), .ZN(n8012) );
  AOI221_X1 U10414 ( .B1(P1_IR_REG_12__SCAN_IN), .B2(keyinput_f119), .C1(
        P1_IR_REG_9__SCAN_IN), .C2(keyinput_f116), .A(n8012), .ZN(n8013) );
  NAND4_X1 U10415 ( .A1(n8016), .A2(n8015), .A3(n8014), .A4(n8013), .ZN(n8036)
         );
  OAI22_X1 U10416 ( .A1(P3_REG3_REG_27__SCAN_IN), .A2(keyinput_f36), .B1(
        P3_DATAO_REG_27__SCAN_IN), .B2(keyinput_f69), .ZN(n8017) );
  AOI221_X1 U10417 ( .B1(P3_REG3_REG_27__SCAN_IN), .B2(keyinput_f36), .C1(
        keyinput_f69), .C2(P3_DATAO_REG_27__SCAN_IN), .A(n8017), .ZN(n8024) );
  OAI22_X1 U10418 ( .A1(SI_1_), .A2(keyinput_f31), .B1(keyinput_f117), .B2(
        P1_IR_REG_10__SCAN_IN), .ZN(n8018) );
  AOI221_X1 U10419 ( .B1(SI_1_), .B2(keyinput_f31), .C1(P1_IR_REG_10__SCAN_IN), 
        .C2(keyinput_f117), .A(n8018), .ZN(n8023) );
  OAI22_X1 U10420 ( .A1(P3_REG3_REG_21__SCAN_IN), .A2(keyinput_f45), .B1(
        P1_IR_REG_7__SCAN_IN), .B2(keyinput_f114), .ZN(n8019) );
  AOI221_X1 U10421 ( .B1(P3_REG3_REG_21__SCAN_IN), .B2(keyinput_f45), .C1(
        keyinput_f114), .C2(P1_IR_REG_7__SCAN_IN), .A(n8019), .ZN(n8022) );
  OAI22_X1 U10422 ( .A1(P3_REG3_REG_8__SCAN_IN), .A2(keyinput_f43), .B1(
        P3_DATAO_REG_3__SCAN_IN), .B2(keyinput_f93), .ZN(n8020) );
  AOI221_X1 U10423 ( .B1(P3_REG3_REG_8__SCAN_IN), .B2(keyinput_f43), .C1(
        keyinput_f93), .C2(P3_DATAO_REG_3__SCAN_IN), .A(n8020), .ZN(n8021) );
  NAND4_X1 U10424 ( .A1(n8024), .A2(n8023), .A3(n8022), .A4(n8021), .ZN(n8035)
         );
  OAI22_X1 U10425 ( .A1(P3_REG3_REG_25__SCAN_IN), .A2(keyinput_f47), .B1(SI_8_), .B2(keyinput_f24), .ZN(n8025) );
  AOI221_X1 U10426 ( .B1(P3_REG3_REG_25__SCAN_IN), .B2(keyinput_f47), .C1(
        keyinput_f24), .C2(SI_8_), .A(n8025), .ZN(n8033) );
  OAI22_X1 U10427 ( .A1(P3_ADDR_REG_7__SCAN_IN), .A2(keyinput_f104), .B1(
        keyinput_f95), .B2(P3_DATAO_REG_1__SCAN_IN), .ZN(n8026) );
  AOI221_X1 U10428 ( .B1(P3_ADDR_REG_7__SCAN_IN), .B2(keyinput_f104), .C1(
        P3_DATAO_REG_1__SCAN_IN), .C2(keyinput_f95), .A(n8026), .ZN(n8032) );
  OAI22_X1 U10429 ( .A1(keyinput_f67), .A2(P3_DATAO_REG_29__SCAN_IN), .B1(
        P3_DATAO_REG_14__SCAN_IN), .B2(keyinput_f82), .ZN(n8027) );
  AOI221_X1 U10430 ( .B1(keyinput_f67), .B2(P3_DATAO_REG_29__SCAN_IN), .C1(
        keyinput_f82), .C2(P3_DATAO_REG_14__SCAN_IN), .A(n8027), .ZN(n8031) );
  XOR2_X1 U10431 ( .A(SI_0_), .B(keyinput_f32), .Z(n8029) );
  XNOR2_X1 U10432 ( .A(P1_IR_REG_8__SCAN_IN), .B(keyinput_f115), .ZN(n8028) );
  NOR2_X1 U10433 ( .A1(n8029), .A2(n8028), .ZN(n8030) );
  NAND4_X1 U10434 ( .A1(n8033), .A2(n8032), .A3(n8031), .A4(n8030), .ZN(n8034)
         );
  NOR4_X1 U10435 ( .A1(n8037), .A2(n8036), .A3(n8035), .A4(n8034), .ZN(n8167)
         );
  OAI22_X1 U10436 ( .A1(P3_REG3_REG_23__SCAN_IN), .A2(keyinput_f38), .B1(
        P3_REG3_REG_9__SCAN_IN), .B2(keyinput_f53), .ZN(n8038) );
  AOI221_X1 U10437 ( .B1(P3_REG3_REG_23__SCAN_IN), .B2(keyinput_f38), .C1(
        keyinput_f53), .C2(P3_REG3_REG_9__SCAN_IN), .A(n8038), .ZN(n8045) );
  OAI22_X1 U10438 ( .A1(P3_REG3_REG_3__SCAN_IN), .A2(keyinput_f40), .B1(
        keyinput_f88), .B2(P3_DATAO_REG_8__SCAN_IN), .ZN(n8039) );
  AOI221_X1 U10439 ( .B1(P3_REG3_REG_3__SCAN_IN), .B2(keyinput_f40), .C1(
        P3_DATAO_REG_8__SCAN_IN), .C2(keyinput_f88), .A(n8039), .ZN(n8044) );
  OAI22_X1 U10440 ( .A1(SI_26_), .A2(keyinput_f6), .B1(keyinput_f103), .B2(
        P3_ADDR_REG_6__SCAN_IN), .ZN(n8040) );
  AOI221_X1 U10441 ( .B1(SI_26_), .B2(keyinput_f6), .C1(P3_ADDR_REG_6__SCAN_IN), .C2(keyinput_f103), .A(n8040), .ZN(n8043) );
  OAI22_X1 U10442 ( .A1(P3_REG3_REG_10__SCAN_IN), .A2(keyinput_f39), .B1(
        P3_B_REG_SCAN_IN), .B2(keyinput_f64), .ZN(n8041) );
  AOI221_X1 U10443 ( .B1(P3_REG3_REG_10__SCAN_IN), .B2(keyinput_f39), .C1(
        keyinput_f64), .C2(P3_B_REG_SCAN_IN), .A(n8041), .ZN(n8042) );
  NAND4_X1 U10444 ( .A1(n8045), .A2(n8044), .A3(n8043), .A4(n8042), .ZN(n8165)
         );
  OAI22_X1 U10445 ( .A1(SI_19_), .A2(keyinput_f13), .B1(keyinput_f126), .B2(
        P1_IR_REG_19__SCAN_IN), .ZN(n8046) );
  AOI221_X1 U10446 ( .B1(SI_19_), .B2(keyinput_f13), .C1(P1_IR_REG_19__SCAN_IN), .C2(keyinput_f126), .A(n8046), .ZN(n8071) );
  OAI22_X1 U10447 ( .A1(SI_31_), .A2(keyinput_f1), .B1(keyinput_f52), .B2(
        P3_REG3_REG_4__SCAN_IN), .ZN(n8047) );
  AOI221_X1 U10448 ( .B1(SI_31_), .B2(keyinput_f1), .C1(P3_REG3_REG_4__SCAN_IN), .C2(keyinput_f52), .A(n8047), .ZN(n8050) );
  OAI22_X1 U10449 ( .A1(SI_11_), .A2(keyinput_f21), .B1(keyinput_f66), .B2(
        P3_DATAO_REG_30__SCAN_IN), .ZN(n8048) );
  AOI221_X1 U10450 ( .B1(SI_11_), .B2(keyinput_f21), .C1(
        P3_DATAO_REG_30__SCAN_IN), .C2(keyinput_f66), .A(n8048), .ZN(n8049) );
  OAI211_X1 U10451 ( .C1(n11902), .C2(keyinput_f58), .A(n8050), .B(n8049), 
        .ZN(n8051) );
  AOI21_X1 U10452 ( .B1(n11902), .B2(keyinput_f58), .A(n8051), .ZN(n8070) );
  AOI22_X1 U10453 ( .A1(P3_DATAO_REG_31__SCAN_IN), .A2(keyinput_f65), .B1(
        SI_14_), .B2(keyinput_f18), .ZN(n8052) );
  OAI221_X1 U10454 ( .B1(P3_DATAO_REG_31__SCAN_IN), .B2(keyinput_f65), .C1(
        SI_14_), .C2(keyinput_f18), .A(n8052), .ZN(n8059) );
  AOI22_X1 U10455 ( .A1(keyinput_f84), .A2(P3_DATAO_REG_12__SCAN_IN), .B1(
        P1_IR_REG_16__SCAN_IN), .B2(keyinput_f123), .ZN(n8053) );
  OAI221_X1 U10456 ( .B1(keyinput_f84), .B2(P3_DATAO_REG_12__SCAN_IN), .C1(
        P1_IR_REG_16__SCAN_IN), .C2(keyinput_f123), .A(n8053), .ZN(n8058) );
  AOI22_X1 U10457 ( .A1(keyinput_f75), .A2(P3_DATAO_REG_21__SCAN_IN), .B1(
        SI_15_), .B2(keyinput_f17), .ZN(n8054) );
  OAI221_X1 U10458 ( .B1(keyinput_f75), .B2(P3_DATAO_REG_21__SCAN_IN), .C1(
        SI_15_), .C2(keyinput_f17), .A(n8054), .ZN(n8057) );
  AOI22_X1 U10459 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(keyinput_f108), .B1(SI_7_), 
        .B2(keyinput_f25), .ZN(n8055) );
  OAI221_X1 U10460 ( .B1(P1_IR_REG_1__SCAN_IN), .B2(keyinput_f108), .C1(SI_7_), 
        .C2(keyinput_f25), .A(n8055), .ZN(n8056) );
  NOR4_X1 U10461 ( .A1(n8059), .A2(n8058), .A3(n8057), .A4(n8056), .ZN(n8069)
         );
  AOI22_X1 U10462 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(keyinput_f120), .B1(
        P3_REG3_REG_0__SCAN_IN), .B2(keyinput_f54), .ZN(n8060) );
  OAI221_X1 U10463 ( .B1(P1_IR_REG_13__SCAN_IN), .B2(keyinput_f120), .C1(
        P3_REG3_REG_0__SCAN_IN), .C2(keyinput_f54), .A(n8060), .ZN(n8067) );
  AOI22_X1 U10464 ( .A1(P3_ADDR_REG_4__SCAN_IN), .A2(keyinput_f101), .B1(SI_4_), .B2(keyinput_f28), .ZN(n8061) );
  OAI221_X1 U10465 ( .B1(P3_ADDR_REG_4__SCAN_IN), .B2(keyinput_f101), .C1(
        SI_4_), .C2(keyinput_f28), .A(n8061), .ZN(n8066) );
  AOI22_X1 U10466 ( .A1(keyinput_f83), .A2(P3_DATAO_REG_13__SCAN_IN), .B1(
        P1_IR_REG_15__SCAN_IN), .B2(keyinput_f122), .ZN(n8062) );
  OAI221_X1 U10467 ( .B1(keyinput_f83), .B2(P3_DATAO_REG_13__SCAN_IN), .C1(
        P1_IR_REG_15__SCAN_IN), .C2(keyinput_f122), .A(n8062), .ZN(n8065) );
  AOI22_X1 U10468 ( .A1(keyinput_f0), .A2(P3_WR_REG_SCAN_IN), .B1(SI_30_), 
        .B2(keyinput_f2), .ZN(n8063) );
  OAI221_X1 U10469 ( .B1(keyinput_f0), .B2(P3_WR_REG_SCAN_IN), .C1(SI_30_), 
        .C2(keyinput_f2), .A(n8063), .ZN(n8064) );
  NOR4_X1 U10470 ( .A1(n8067), .A2(n8066), .A3(n8065), .A4(n8064), .ZN(n8068)
         );
  NAND4_X1 U10471 ( .A1(n8071), .A2(n8070), .A3(n8069), .A4(n8068), .ZN(n8164)
         );
  AOI22_X1 U10472 ( .A1(n10648), .A2(keyinput_f73), .B1(n13314), .B2(
        keyinput_f57), .ZN(n8072) );
  OAI221_X1 U10473 ( .B1(n10648), .B2(keyinput_f73), .C1(n13314), .C2(
        keyinput_f57), .A(n8072), .ZN(n8081) );
  AOI22_X1 U10474 ( .A1(n13841), .A2(keyinput_f3), .B1(keyinput_f20), .B2(
        n9999), .ZN(n8073) );
  OAI221_X1 U10475 ( .B1(n13841), .B2(keyinput_f3), .C1(n9999), .C2(
        keyinput_f20), .A(n8073), .ZN(n8080) );
  INV_X1 U10476 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n8075) );
  AOI22_X1 U10477 ( .A1(n8075), .A2(keyinput_f121), .B1(n9373), .B2(
        keyinput_f10), .ZN(n8074) );
  OAI221_X1 U10478 ( .B1(n8075), .B2(keyinput_f121), .C1(n9373), .C2(
        keyinput_f10), .A(n8074), .ZN(n8079) );
  XNOR2_X1 U10479 ( .A(SI_3_), .B(keyinput_f29), .ZN(n8077) );
  XNOR2_X1 U10480 ( .A(SI_16_), .B(keyinput_f16), .ZN(n8076) );
  NAND2_X1 U10481 ( .A1(n8077), .A2(n8076), .ZN(n8078) );
  NOR4_X1 U10482 ( .A1(n8081), .A2(n8080), .A3(n8079), .A4(n8078), .ZN(n8116)
         );
  AOI22_X1 U10483 ( .A1(n8083), .A2(keyinput_f106), .B1(keyinput_f74), .B2(
        n10646), .ZN(n8082) );
  OAI221_X1 U10484 ( .B1(n8083), .B2(keyinput_f106), .C1(n10646), .C2(
        keyinput_f74), .A(n8082), .ZN(n8091) );
  AOI22_X1 U10485 ( .A1(n11600), .A2(keyinput_f9), .B1(keyinput_f76), .B2(
        n10637), .ZN(n8084) );
  OAI221_X1 U10486 ( .B1(n11600), .B2(keyinput_f9), .C1(n10637), .C2(
        keyinput_f76), .A(n8084), .ZN(n8090) );
  INV_X1 U10487 ( .A(P3_DATAO_REG_10__SCAN_IN), .ZN(n10635) );
  AOI22_X1 U10488 ( .A1(n10624), .A2(keyinput_f91), .B1(keyinput_f86), .B2(
        n10635), .ZN(n8085) );
  OAI221_X1 U10489 ( .B1(n10624), .B2(keyinput_f91), .C1(n10635), .C2(
        keyinput_f86), .A(n8085), .ZN(n8089) );
  XNOR2_X1 U10490 ( .A(P1_IR_REG_6__SCAN_IN), .B(keyinput_f113), .ZN(n8087) );
  XNOR2_X1 U10491 ( .A(SI_2_), .B(keyinput_f30), .ZN(n8086) );
  NAND2_X1 U10492 ( .A1(n8087), .A2(n8086), .ZN(n8088) );
  NOR4_X1 U10493 ( .A1(n8091), .A2(n8090), .A3(n8089), .A4(n8088), .ZN(n8115)
         );
  INV_X1 U10494 ( .A(P3_DATAO_REG_15__SCAN_IN), .ZN(n10559) );
  AOI22_X1 U10495 ( .A1(n10641), .A2(keyinput_f89), .B1(keyinput_f81), .B2(
        n10559), .ZN(n8092) );
  OAI221_X1 U10496 ( .B1(n10641), .B2(keyinput_f89), .C1(n10559), .C2(
        keyinput_f81), .A(n8092), .ZN(n8095) );
  XOR2_X1 U10497 ( .A(P1_IR_REG_4__SCAN_IN), .B(keyinput_f111), .Z(n8094) );
  XNOR2_X1 U10498 ( .A(n10666), .B(keyinput_f72), .ZN(n8093) );
  OR3_X1 U10499 ( .A1(n8095), .A2(n8094), .A3(n8093), .ZN(n8100) );
  AOI22_X1 U10500 ( .A1(n10798), .A2(keyinput_f61), .B1(keyinput_f44), .B2(
        n15728), .ZN(n8096) );
  OAI221_X1 U10501 ( .B1(n10798), .B2(keyinput_f61), .C1(n15728), .C2(
        keyinput_f44), .A(n8096), .ZN(n8099) );
  AOI22_X1 U10502 ( .A1(n9297), .A2(keyinput_f50), .B1(keyinput_f68), .B2(
        n11342), .ZN(n8097) );
  OAI221_X1 U10503 ( .B1(n9297), .B2(keyinput_f50), .C1(n11342), .C2(
        keyinput_f68), .A(n8097), .ZN(n8098) );
  NOR3_X1 U10504 ( .A1(n8100), .A2(n8099), .A3(n8098), .ZN(n8114) );
  AOI22_X1 U10505 ( .A1(n10629), .A2(keyinput_f92), .B1(n8102), .B2(
        keyinput_f98), .ZN(n8101) );
  OAI221_X1 U10506 ( .B1(n10629), .B2(keyinput_f92), .C1(n8102), .C2(
        keyinput_f98), .A(n8101), .ZN(n8112) );
  AOI22_X1 U10507 ( .A1(n8104), .A2(keyinput_f105), .B1(n10866), .B2(
        keyinput_f35), .ZN(n8103) );
  OAI221_X1 U10508 ( .B1(n8104), .B2(keyinput_f105), .C1(n10866), .C2(
        keyinput_f35), .A(n8103), .ZN(n8111) );
  INV_X1 U10509 ( .A(P3_REG3_REG_20__SCAN_IN), .ZN(n9343) );
  AOI22_X1 U10510 ( .A1(n8106), .A2(keyinput_f99), .B1(n9343), .B2(
        keyinput_f55), .ZN(n8105) );
  OAI221_X1 U10511 ( .B1(n8106), .B2(keyinput_f99), .C1(n9343), .C2(
        keyinput_f55), .A(n8105), .ZN(n8110) );
  XNOR2_X1 U10512 ( .A(P1_IR_REG_0__SCAN_IN), .B(keyinput_f107), .ZN(n8108) );
  XNOR2_X1 U10513 ( .A(P3_REG3_REG_16__SCAN_IN), .B(keyinput_f48), .ZN(n8107)
         );
  NAND2_X1 U10514 ( .A1(n8108), .A2(n8107), .ZN(n8109) );
  NOR4_X1 U10515 ( .A1(n8112), .A2(n8111), .A3(n8110), .A4(n8109), .ZN(n8113)
         );
  NAND4_X1 U10516 ( .A1(n8116), .A2(n8115), .A3(n8114), .A4(n8113), .ZN(n8163)
         );
  INV_X1 U10517 ( .A(SI_9_), .ZN(n9969) );
  AOI22_X1 U10518 ( .A1(n9969), .A2(keyinput_f23), .B1(n11988), .B2(
        keyinput_f46), .ZN(n8117) );
  OAI221_X1 U10519 ( .B1(n9969), .B2(keyinput_f23), .C1(n11988), .C2(
        keyinput_f46), .A(n8117), .ZN(n8125) );
  AOI22_X1 U10520 ( .A1(n10924), .A2(keyinput_f12), .B1(keyinput_f96), .B2(
        n10633), .ZN(n8118) );
  OAI221_X1 U10521 ( .B1(n10924), .B2(keyinput_f12), .C1(n10633), .C2(
        keyinput_f96), .A(n8118), .ZN(n8124) );
  AOI22_X1 U10522 ( .A1(n11063), .A2(keyinput_f70), .B1(n10016), .B2(
        keyinput_f19), .ZN(n8119) );
  OAI221_X1 U10523 ( .B1(n11063), .B2(keyinput_f70), .C1(n10016), .C2(
        keyinput_f19), .A(n8119), .ZN(n8123) );
  INV_X1 U10524 ( .A(P3_DATAO_REG_19__SCAN_IN), .ZN(n10565) );
  AOI22_X1 U10525 ( .A1(n10565), .A2(keyinput_f77), .B1(n8121), .B2(
        keyinput_f100), .ZN(n8120) );
  OAI221_X1 U10526 ( .B1(n10565), .B2(keyinput_f77), .C1(n8121), .C2(
        keyinput_f100), .A(n8120), .ZN(n8122) );
  NOR4_X1 U10527 ( .A1(n8125), .A2(n8124), .A3(n8123), .A4(n8122), .ZN(n8161)
         );
  INV_X1 U10528 ( .A(P3_REG3_REG_14__SCAN_IN), .ZN(n13226) );
  INV_X1 U10529 ( .A(SI_28_), .ZN(n8127) );
  AOI22_X1 U10530 ( .A1(n13226), .A2(keyinput_f37), .B1(keyinput_f4), .B2(
        n8127), .ZN(n8126) );
  OAI221_X1 U10531 ( .B1(n13226), .B2(keyinput_f37), .C1(n8127), .C2(
        keyinput_f4), .A(n8126), .ZN(n8135) );
  INV_X1 U10532 ( .A(P3_REG3_REG_15__SCAN_IN), .ZN(n13344) );
  AOI22_X1 U10533 ( .A1(n10522), .A2(keyinput_f14), .B1(n13344), .B2(
        keyinput_f63), .ZN(n8128) );
  OAI221_X1 U10534 ( .B1(n10522), .B2(keyinput_f14), .C1(n13344), .C2(
        keyinput_f63), .A(n8128), .ZN(n8134) );
  INV_X1 U10535 ( .A(SI_27_), .ZN(n13845) );
  INV_X2 U10536 ( .A(P3_STATE_REG_SCAN_IN), .ZN(P3_U3151) );
  AOI22_X1 U10537 ( .A1(n13845), .A2(keyinput_f5), .B1(P3_U3151), .B2(
        keyinput_f34), .ZN(n8129) );
  OAI221_X1 U10538 ( .B1(n13845), .B2(keyinput_f5), .C1(P3_U3151), .C2(
        keyinput_f34), .A(n8129), .ZN(n8133) );
  XNOR2_X1 U10539 ( .A(SI_6_), .B(keyinput_f26), .ZN(n8131) );
  XNOR2_X1 U10540 ( .A(SI_21_), .B(keyinput_f11), .ZN(n8130) );
  NAND2_X1 U10541 ( .A1(n8131), .A2(n8130), .ZN(n8132) );
  NOR4_X1 U10542 ( .A1(n8135), .A2(n8134), .A3(n8133), .A4(n8132), .ZN(n8160)
         );
  INV_X1 U10543 ( .A(P3_DATAO_REG_11__SCAN_IN), .ZN(n10639) );
  AOI22_X1 U10544 ( .A1(n10639), .A2(keyinput_f85), .B1(n10436), .B2(
        keyinput_f15), .ZN(n8136) );
  OAI221_X1 U10545 ( .B1(n10639), .B2(keyinput_f85), .C1(n10436), .C2(
        keyinput_f15), .A(n8136), .ZN(n8139) );
  XNOR2_X1 U10546 ( .A(n9846), .B(keyinput_f125), .ZN(n8138) );
  XNOR2_X1 U10547 ( .A(n10859), .B(keyinput_f71), .ZN(n8137) );
  OR3_X1 U10548 ( .A1(n8139), .A2(n8138), .A3(n8137), .ZN(n8146) );
  AOI22_X1 U10549 ( .A1(n8142), .A2(keyinput_f42), .B1(keyinput_f97), .B2(
        n8141), .ZN(n8140) );
  OAI221_X1 U10550 ( .B1(n8142), .B2(keyinput_f42), .C1(n8141), .C2(
        keyinput_f97), .A(n8140), .ZN(n8145) );
  INV_X1 U10551 ( .A(P3_DATAO_REG_6__SCAN_IN), .ZN(n10631) );
  AOI22_X1 U10552 ( .A1(n10631), .A2(keyinput_f90), .B1(n9235), .B2(
        keyinput_f56), .ZN(n8143) );
  OAI221_X1 U10553 ( .B1(n10631), .B2(keyinput_f90), .C1(n9235), .C2(
        keyinput_f56), .A(n8143), .ZN(n8144) );
  NOR3_X1 U10554 ( .A1(n8146), .A2(n8145), .A3(n8144), .ZN(n8159) );
  XNOR2_X1 U10555 ( .A(n9992), .B(keyinput_f112), .ZN(n8150) );
  XNOR2_X1 U10556 ( .A(n9794), .B(keyinput_f124), .ZN(n8149) );
  INV_X1 U10557 ( .A(SI_24_), .ZN(n8147) );
  XNOR2_X1 U10558 ( .A(keyinput_f8), .B(n8147), .ZN(n8148) );
  NOR3_X1 U10559 ( .A1(n8150), .A2(n8149), .A3(n8148), .ZN(n8153) );
  XOR2_X1 U10560 ( .A(n10682), .B(keyinput_f59), .Z(n8152) );
  XNOR2_X1 U10561 ( .A(P1_IR_REG_3__SCAN_IN), .B(keyinput_f110), .ZN(n8151) );
  NAND3_X1 U10562 ( .A1(n8153), .A2(n8152), .A3(n8151), .ZN(n8157) );
  INV_X1 U10563 ( .A(P3_RD_REG_SCAN_IN), .ZN(n15250) );
  AOI22_X1 U10564 ( .A1(n15250), .A2(keyinput_f33), .B1(n10889), .B2(
        keyinput_f49), .ZN(n8154) );
  OAI221_X1 U10565 ( .B1(n15250), .B2(keyinput_f33), .C1(n10889), .C2(
        keyinput_f49), .A(n8154), .ZN(n8156) );
  INV_X1 U10566 ( .A(P3_DATAO_REG_17__SCAN_IN), .ZN(n10325) );
  XNOR2_X1 U10567 ( .A(n10325), .B(keyinput_f79), .ZN(n8155) );
  NOR3_X1 U10568 ( .A1(n8157), .A2(n8156), .A3(n8155), .ZN(n8158) );
  NAND4_X1 U10569 ( .A1(n8161), .A2(n8160), .A3(n8159), .A4(n8158), .ZN(n8162)
         );
  NOR4_X1 U10570 ( .A1(n8165), .A2(n8164), .A3(n8163), .A4(n8162), .ZN(n8166)
         );
  NAND2_X1 U10571 ( .A1(n8167), .A2(n8166), .ZN(n8169) );
  AOI21_X1 U10572 ( .B1(keyinput_f22), .B2(n8169), .A(SI_10_), .ZN(n8171) );
  INV_X1 U10573 ( .A(keyinput_f22), .ZN(n8168) );
  AOI21_X1 U10574 ( .B1(n8169), .B2(n8168), .A(keyinput_g22), .ZN(n8170) );
  AOI22_X1 U10575 ( .A1(keyinput_g22), .A2(n8171), .B1(SI_10_), .B2(n8170), 
        .ZN(n8172) );
  AOI21_X1 U10576 ( .B1(n8174), .B2(n8173), .A(n8172), .ZN(n8175) );
  INV_X1 U10577 ( .A(n8175), .ZN(n8176) );
  AND3_X1 U10578 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .A3(P2_REG3_REG_5__SCAN_IN), .ZN(n8423) );
  NAND2_X1 U10579 ( .A1(n8423), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n8476) );
  NAND2_X1 U10580 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(P2_REG3_REG_7__SCAN_IN), 
        .ZN(n8179) );
  NOR2_X1 U10581 ( .A1(n8476), .A2(n8179), .ZN(n8474) );
  NAND2_X1 U10582 ( .A1(n8474), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n8513) );
  INV_X1 U10583 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n8512) );
  INV_X1 U10584 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n8528) );
  INV_X1 U10585 ( .A(n8548), .ZN(n8180) );
  NAND2_X1 U10586 ( .A1(n8180), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n8571) );
  INV_X1 U10587 ( .A(n8571), .ZN(n8181) );
  NAND2_X1 U10588 ( .A1(n8181), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n8587) );
  INV_X1 U10589 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n12258) );
  NAND2_X1 U10590 ( .A1(n8628), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n8665) );
  INV_X1 U10591 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n13942) );
  INV_X1 U10592 ( .A(n8684), .ZN(n8182) );
  NAND2_X1 U10593 ( .A1(n8182), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n8694) );
  INV_X1 U10594 ( .A(n8694), .ZN(n8183) );
  NAND2_X1 U10595 ( .A1(n8183), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n8718) );
  INV_X1 U10596 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n13874) );
  NAND2_X1 U10597 ( .A1(P2_REG3_REG_22__SCAN_IN), .A2(P2_REG3_REG_23__SCAN_IN), 
        .ZN(n8184) );
  INV_X1 U10598 ( .A(n8761), .ZN(n8185) );
  INV_X1 U10599 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n13882) );
  INV_X1 U10600 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n8186) );
  OAI21_X1 U10601 ( .B1(n8775), .B2(n13882), .A(n8186), .ZN(n8189) );
  INV_X1 U10602 ( .A(n8775), .ZN(n8188) );
  AND2_X1 U10603 ( .A1(P2_REG3_REG_26__SCAN_IN), .A2(P2_REG3_REG_25__SCAN_IN), 
        .ZN(n8187) );
  INV_X1 U10604 ( .A(n8793), .ZN(n8795) );
  NAND2_X1 U10605 ( .A1(n8189), .A2(n8795), .ZN(n14075) );
  NAND2_X1 U10606 ( .A1(n8342), .A2(n8193), .ZN(n8361) );
  NOR2_X1 U10607 ( .A1(P2_IR_REG_10__SCAN_IN), .A2(P2_IR_REG_14__SCAN_IN), 
        .ZN(n8199) );
  NAND4_X1 U10608 ( .A1(n8199), .A2(n8198), .A3(n8562), .A4(n8197), .ZN(n8323)
         );
  NAND4_X1 U10609 ( .A1(n8200), .A2(n8643), .A3(n8624), .A4(n7030), .ZN(n8201)
         );
  NOR2_X1 U10610 ( .A1(n8323), .A2(n8201), .ZN(n8202) );
  NOR2_X1 U10611 ( .A1(P2_IR_REG_23__SCAN_IN), .A2(P2_IR_REG_22__SCAN_IN), 
        .ZN(n8203) );
  NAND4_X1 U10612 ( .A1(n8203), .A2(n8837), .A3(n8833), .A4(n8830), .ZN(n8312)
         );
  NAND3_X1 U10613 ( .A1(n8204), .A2(n8230), .A3(n8313), .ZN(n8205) );
  NOR2_X1 U10614 ( .A1(n8312), .A2(n8205), .ZN(n8206) );
  NAND2_X1 U10615 ( .A1(n8210), .A2(n8207), .ZN(n14382) );
  OR2_X1 U10616 ( .A1(n14075), .A2(n8874), .ZN(n8223) );
  CLKBUF_X3 U10617 ( .A(n8384), .Z(n10131) );
  INV_X1 U10618 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n14257) );
  AND2_X2 U10619 ( .A1(n8217), .A2(n14388), .ZN(n8667) );
  CLKBUF_X3 U10620 ( .A(n8667), .Z(n8942) );
  NAND2_X1 U10621 ( .A1(n8942), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n8220) );
  NAND2_X1 U10622 ( .A1(n8941), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n8219) );
  OAI211_X1 U10623 ( .C1(n8945), .C2(n14257), .A(n8220), .B(n8219), .ZN(n8221)
         );
  INV_X1 U10624 ( .A(n8221), .ZN(n8222) );
  NAND2_X1 U10625 ( .A1(n8223), .A2(n8222), .ZN(n13963) );
  NAND2_X1 U10626 ( .A1(n8827), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8226) );
  NAND2_X1 U10627 ( .A1(n8229), .A2(n8230), .ZN(n8227) );
  NAND2_X1 U10628 ( .A1(n13099), .A2(n13158), .ZN(n8860) );
  INV_X1 U10629 ( .A(n11849), .ZN(n13122) );
  NAND2_X1 U10630 ( .A1(n13963), .A2(n6670), .ZN(n8785) );
  INV_X1 U10631 ( .A(n8785), .ZN(n8787) );
  INV_X1 U10632 ( .A(SI_1_), .ZN(n9955) );
  AND2_X1 U10633 ( .A1(P2_DATAO_REG_0__SCAN_IN), .A2(SI_0_), .ZN(n8235) );
  NAND2_X1 U10634 ( .A1(n7202), .A2(n8235), .ZN(n9872) );
  AND2_X1 U10635 ( .A1(SI_0_), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n8236) );
  NAND2_X1 U10636 ( .A1(n9975), .A2(n8236), .ZN(n8328) );
  NAND2_X1 U10637 ( .A1(n9872), .A2(n8328), .ZN(n8345) );
  MUX2_X1 U10638 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(P1_DATAO_REG_2__SCAN_IN), 
        .S(n9975), .Z(n8356) );
  INV_X1 U10639 ( .A(n8239), .ZN(n8240) );
  NAND2_X1 U10640 ( .A1(n8240), .A2(SI_2_), .ZN(n8241) );
  MUX2_X1 U10641 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(P1_DATAO_REG_3__SCAN_IN), 
        .S(n9975), .Z(n8242) );
  INV_X1 U10642 ( .A(SI_3_), .ZN(n9960) );
  NAND2_X1 U10643 ( .A1(n8242), .A2(SI_3_), .ZN(n8243) );
  MUX2_X1 U10644 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(P1_DATAO_REG_4__SCAN_IN), 
        .S(n9975), .Z(n8245) );
  XNOR2_X1 U10645 ( .A(n8245), .B(SI_4_), .ZN(n8394) );
  INV_X1 U10646 ( .A(n8394), .ZN(n8244) );
  NAND2_X1 U10647 ( .A1(n8245), .A2(SI_4_), .ZN(n8246) );
  MUX2_X1 U10648 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(P1_DATAO_REG_5__SCAN_IN), 
        .S(n9975), .Z(n8247) );
  XNOR2_X1 U10649 ( .A(n8247), .B(SI_5_), .ZN(n8410) );
  NAND2_X1 U10650 ( .A1(n8247), .A2(SI_5_), .ZN(n8248) );
  MUX2_X1 U10651 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(P1_DATAO_REG_6__SCAN_IN), 
        .S(n9950), .Z(n8250) );
  XNOR2_X1 U10652 ( .A(n8250), .B(SI_6_), .ZN(n8437) );
  INV_X1 U10653 ( .A(n8437), .ZN(n8249) );
  NAND2_X1 U10654 ( .A1(n8438), .A2(n8249), .ZN(n8252) );
  NAND2_X1 U10655 ( .A1(n8250), .A2(SI_6_), .ZN(n8251) );
  INV_X4 U10656 ( .A(n8253), .ZN(n9950) );
  MUX2_X1 U10657 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(P1_DATAO_REG_7__SCAN_IN), 
        .S(n9950), .Z(n8255) );
  INV_X1 U10658 ( .A(n8454), .ZN(n8254) );
  NAND2_X1 U10659 ( .A1(n8255), .A2(SI_7_), .ZN(n8256) );
  MUX2_X1 U10660 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(P1_DATAO_REG_8__SCAN_IN), 
        .S(n9950), .Z(n8257) );
  MUX2_X1 U10661 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(P1_DATAO_REG_9__SCAN_IN), 
        .S(n9950), .Z(n8259) );
  XNOR2_X1 U10662 ( .A(n8259), .B(SI_9_), .ZN(n8488) );
  INV_X1 U10663 ( .A(n8488), .ZN(n8258) );
  NAND2_X1 U10664 ( .A1(n8259), .A2(SI_9_), .ZN(n8260) );
  MUX2_X1 U10665 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(P1_DATAO_REG_10__SCAN_IN), 
        .S(n9950), .Z(n8262) );
  XNOR2_X1 U10666 ( .A(n8262), .B(SI_10_), .ZN(n8507) );
  INV_X1 U10667 ( .A(n8507), .ZN(n8261) );
  NAND2_X1 U10668 ( .A1(n8262), .A2(SI_10_), .ZN(n8263) );
  MUX2_X1 U10669 ( .A(n10246), .B(n10238), .S(n9950), .Z(n8264) );
  NAND2_X1 U10670 ( .A1(n8264), .A2(n9984), .ZN(n8267) );
  INV_X1 U10671 ( .A(n8264), .ZN(n8265) );
  NAND2_X1 U10672 ( .A1(n8265), .A2(SI_11_), .ZN(n8266) );
  NAND2_X1 U10673 ( .A1(n8267), .A2(n8266), .ZN(n8523) );
  MUX2_X1 U10674 ( .A(n10360), .B(n10352), .S(n9950), .Z(n8268) );
  INV_X1 U10675 ( .A(n8268), .ZN(n8269) );
  NAND2_X1 U10676 ( .A1(n8269), .A2(SI_12_), .ZN(n8270) );
  MUX2_X1 U10677 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(P1_DATAO_REG_13__SCAN_IN), 
        .S(n9950), .Z(n8559) );
  INV_X1 U10678 ( .A(n8559), .ZN(n8272) );
  MUX2_X1 U10679 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(P1_DATAO_REG_15__SCAN_IN), 
        .S(n9950), .Z(n8603) );
  NAND2_X1 U10680 ( .A1(n8603), .A2(SI_15_), .ZN(n8275) );
  MUX2_X1 U10681 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(P1_DATAO_REG_14__SCAN_IN), 
        .S(n9950), .Z(n8597) );
  NAND2_X1 U10682 ( .A1(n8597), .A2(SI_14_), .ZN(n8273) );
  NOR2_X1 U10683 ( .A1(n8597), .A2(SI_14_), .ZN(n8276) );
  INV_X1 U10684 ( .A(n8603), .ZN(n8274) );
  AOI22_X1 U10685 ( .A1(n8276), .A2(n8275), .B1(n8274), .B2(n10130), .ZN(n8277) );
  MUX2_X1 U10686 ( .A(n6925), .B(n10656), .S(n9950), .Z(n8278) );
  XNOR2_X1 U10687 ( .A(n8278), .B(SI_16_), .ZN(n8621) );
  NAND2_X1 U10688 ( .A1(n8622), .A2(n8621), .ZN(n8280) );
  NAND2_X1 U10689 ( .A1(n8278), .A2(n10250), .ZN(n8279) );
  MUX2_X1 U10690 ( .A(n10671), .B(n10652), .S(n9950), .Z(n8638) );
  NOR2_X1 U10691 ( .A1(n8281), .A2(SI_17_), .ZN(n8283) );
  NAND2_X1 U10692 ( .A1(n8281), .A2(SI_17_), .ZN(n8282) );
  MUX2_X1 U10693 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(P1_DATAO_REG_18__SCAN_IN), 
        .S(n9950), .Z(n8661) );
  NAND2_X1 U10694 ( .A1(n8284), .A2(SI_18_), .ZN(n8285) );
  MUX2_X1 U10695 ( .A(n11316), .B(n12566), .S(n9950), .Z(n8286) );
  INV_X1 U10696 ( .A(n8286), .ZN(n8287) );
  NAND2_X1 U10697 ( .A1(n8287), .A2(SI_19_), .ZN(n8288) );
  NAND2_X1 U10698 ( .A1(n8289), .A2(n8288), .ZN(n8677) );
  MUX2_X1 U10699 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(P1_DATAO_REG_21__SCAN_IN), 
        .S(n9950), .Z(n8713) );
  NOR2_X1 U10700 ( .A1(n8708), .A2(SI_20_), .ZN(n8290) );
  INV_X1 U10701 ( .A(n8708), .ZN(n8291) );
  NOR2_X1 U10702 ( .A1(n8291), .A2(n10924), .ZN(n8294) );
  INV_X1 U10703 ( .A(n8292), .ZN(n8293) );
  AOI22_X1 U10704 ( .A1(n8294), .A2(n8293), .B1(n8713), .B2(SI_21_), .ZN(n8295) );
  MUX2_X1 U10705 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(P1_DATAO_REG_22__SCAN_IN), 
        .S(n9950), .Z(n8733) );
  NAND2_X1 U10706 ( .A1(n8296), .A2(n8733), .ZN(n8299) );
  NAND2_X1 U10707 ( .A1(n8297), .A2(SI_22_), .ZN(n8298) );
  MUX2_X1 U10708 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(P1_DATAO_REG_23__SCAN_IN), 
        .S(n9950), .Z(n8301) );
  XNOR2_X1 U10709 ( .A(n8301), .B(SI_23_), .ZN(n8742) );
  INV_X1 U10710 ( .A(n8742), .ZN(n8300) );
  NAND2_X1 U10711 ( .A1(n8301), .A2(SI_23_), .ZN(n8302) );
  MUX2_X1 U10712 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(P1_DATAO_REG_24__SCAN_IN), 
        .S(n9950), .Z(n8757) );
  NAND2_X1 U10713 ( .A1(n8304), .A2(SI_24_), .ZN(n8305) );
  INV_X1 U10714 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n12481) );
  MUX2_X1 U10715 ( .A(n12481), .B(n12390), .S(n9950), .Z(n8307) );
  INV_X1 U10716 ( .A(SI_25_), .ZN(n12178) );
  NAND2_X1 U10717 ( .A1(n8307), .A2(n12178), .ZN(n8310) );
  INV_X1 U10718 ( .A(n8307), .ZN(n8308) );
  NAND2_X1 U10719 ( .A1(n8308), .A2(SI_25_), .ZN(n8309) );
  NAND2_X1 U10720 ( .A1(n8310), .A2(n8309), .ZN(n8771) );
  MUX2_X1 U10721 ( .A(n15240), .B(n14394), .S(n9950), .Z(n8788) );
  XNOR2_X1 U10722 ( .A(n7674), .B(n13849), .ZN(n8311) );
  XNOR2_X1 U10723 ( .A(n8789), .B(n8311), .ZN(n14393) );
  NAND2_X1 U10724 ( .A1(n8315), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8316) );
  NAND2_X1 U10725 ( .A1(n8381), .A2(n9975), .ZN(n8358) );
  INV_X2 U10726 ( .A(n8358), .ZN(n8412) );
  NAND2_X1 U10727 ( .A1(n14393), .A2(n8412), .ZN(n8320) );
  OR2_X1 U10728 ( .A1(n8379), .A2(n14394), .ZN(n8319) );
  AND2_X2 U10729 ( .A1(n8321), .A2(n11849), .ZN(n8325) );
  INV_X1 U10730 ( .A(n8323), .ZN(n8324) );
  NAND2_X1 U10731 ( .A1(n8508), .A2(n8324), .ZN(n8623) );
  INV_X1 U10732 ( .A(n8325), .ZN(n8326) );
  XNOR2_X1 U10733 ( .A(n14256), .B(n8369), .ZN(n8786) );
  INV_X1 U10734 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n10331) );
  NAND2_X1 U10735 ( .A1(n9975), .A2(SI_0_), .ZN(n8327) );
  NAND2_X1 U10736 ( .A1(n8327), .A2(n9039), .ZN(n8329) );
  AND2_X1 U10737 ( .A1(n8329), .A2(n8328), .ZN(n14397) );
  MUX2_X1 U10738 ( .A(P2_IR_REG_0__SCAN_IN), .B(n14397), .S(n8381), .Z(n12863)
         );
  OR2_X1 U10739 ( .A1(n15616), .A2(n8753), .ZN(n8334) );
  NAND2_X1 U10740 ( .A1(n8384), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n8333) );
  NAND2_X1 U10741 ( .A1(n8667), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n8331) );
  NAND2_X1 U10742 ( .A1(n8336), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n8330) );
  NAND2_X1 U10743 ( .A1(n8334), .A2(n13120), .ZN(n10354) );
  INV_X1 U10744 ( .A(n10354), .ZN(n8335) );
  NAND2_X1 U10745 ( .A1(n8384), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n8339) );
  NAND2_X1 U10746 ( .A1(n8336), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n8338) );
  NAND2_X1 U10747 ( .A1(n8667), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n8337) );
  NAND2_X1 U10748 ( .A1(n13988), .A2(n8753), .ZN(n8350) );
  NAND2_X1 U10749 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), 
        .ZN(n8341) );
  MUX2_X1 U10750 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8341), .S(
        P2_IR_REG_1__SCAN_IN), .Z(n8344) );
  INV_X1 U10751 ( .A(n8342), .ZN(n8343) );
  NAND2_X1 U10752 ( .A1(n8344), .A2(n8343), .ZN(n10261) );
  XNOR2_X1 U10753 ( .A(n8346), .B(n8345), .ZN(n9981) );
  OR2_X1 U10754 ( .A1(n8358), .A2(n9981), .ZN(n8348) );
  INV_X1 U10755 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n9982) );
  XNOR2_X1 U10756 ( .A(n8369), .B(n8886), .ZN(n8349) );
  NAND2_X1 U10757 ( .A1(n10404), .A2(n10405), .ZN(n10403) );
  INV_X1 U10758 ( .A(n8349), .ZN(n8351) );
  NAND2_X1 U10759 ( .A1(n8351), .A2(n8350), .ZN(n8352) );
  NAND2_X1 U10760 ( .A1(n10403), .A2(n8352), .ZN(n10413) );
  NAND2_X1 U10761 ( .A1(n8336), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n8355) );
  NAND2_X1 U10762 ( .A1(n8667), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n8354) );
  NAND2_X1 U10763 ( .A1(n8384), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n8353) );
  INV_X1 U10764 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n9977) );
  XNOR2_X1 U10765 ( .A(n8357), .B(n8356), .ZN(n9976) );
  INV_X1 U10766 ( .A(n10076), .ZN(n8365) );
  NOR2_X1 U10767 ( .A1(n8342), .A2(n14381), .ZN(n8359) );
  MUX2_X1 U10768 ( .A(n14381), .B(n8359), .S(P2_IR_REG_2__SCAN_IN), .Z(n8360)
         );
  INV_X1 U10769 ( .A(n8360), .ZN(n8363) );
  NAND2_X1 U10770 ( .A1(n8363), .A2(n8362), .ZN(n13990) );
  XNOR2_X1 U10771 ( .A(n12882), .B(n8382), .ZN(n8373) );
  INV_X1 U10772 ( .A(n8373), .ZN(n8370) );
  NAND2_X1 U10773 ( .A1(n8371), .A2(n8370), .ZN(n8374) );
  NAND2_X1 U10774 ( .A1(n8373), .A2(n8372), .ZN(n8375) );
  NAND2_X1 U10775 ( .A1(n10413), .A2(n10414), .ZN(n10412) );
  NAND2_X1 U10776 ( .A1(n8362), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8376) );
  MUX2_X1 U10777 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8376), .S(
        P2_IR_REG_3__SCAN_IN), .Z(n8377) );
  OR2_X1 U10778 ( .A1(n8362), .A2(P2_IR_REG_3__SCAN_IN), .ZN(n8413) );
  NAND2_X1 U10779 ( .A1(n8377), .A2(n8413), .ZN(n10166) );
  OR2_X1 U10780 ( .A1(n8379), .A2(n10531), .ZN(n8380) );
  XNOR2_X1 U10781 ( .A(n15652), .B(n8382), .ZN(n8389) );
  INV_X1 U10782 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n8383) );
  NAND2_X1 U10783 ( .A1(n8336), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n8387) );
  NAND2_X1 U10784 ( .A1(n8384), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n8386) );
  NAND2_X1 U10785 ( .A1(n8667), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n8385) );
  NAND2_X1 U10786 ( .A1(n13986), .A2(n6670), .ZN(n8390) );
  INV_X1 U10787 ( .A(n8389), .ZN(n8392) );
  INV_X1 U10788 ( .A(n8390), .ZN(n8391) );
  AOI21_X1 U10789 ( .B1(n8393), .B2(n6837), .A(n7731), .ZN(n10444) );
  XNOR2_X1 U10790 ( .A(n8395), .B(n8394), .ZN(n10945) );
  NAND2_X1 U10791 ( .A1(n10945), .A2(n8412), .ZN(n8398) );
  INV_X2 U10792 ( .A(n8379), .ZN(n8680) );
  INV_X2 U10793 ( .A(n10076), .ZN(n8679) );
  NAND2_X1 U10794 ( .A1(n8413), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8396) );
  XNOR2_X1 U10795 ( .A(n8396), .B(P2_IR_REG_4__SCAN_IN), .ZN(n10309) );
  XNOR2_X1 U10796 ( .A(n15659), .B(n8382), .ZN(n8404) );
  NAND2_X1 U10797 ( .A1(n8667), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n8403) );
  NAND2_X1 U10798 ( .A1(n8336), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n8402) );
  INV_X1 U10799 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n8399) );
  XNOR2_X1 U10800 ( .A(n8399), .B(P2_REG3_REG_3__SCAN_IN), .ZN(n11512) );
  NAND2_X1 U10801 ( .A1(n8817), .A2(n11512), .ZN(n8401) );
  NAND2_X1 U10802 ( .A1(n8384), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n8400) );
  NAND2_X1 U10803 ( .A1(n13985), .A2(n6670), .ZN(n8405) );
  NAND2_X1 U10804 ( .A1(n8404), .A2(n8405), .ZN(n8409) );
  INV_X1 U10805 ( .A(n8404), .ZN(n8407) );
  INV_X1 U10806 ( .A(n8405), .ZN(n8406) );
  NAND2_X1 U10807 ( .A1(n8407), .A2(n8406), .ZN(n8408) );
  AND2_X1 U10808 ( .A1(n8409), .A2(n8408), .ZN(n10443) );
  XNOR2_X1 U10809 ( .A(n8411), .B(n8410), .ZN(n11027) );
  NAND2_X1 U10810 ( .A1(n11027), .A2(n8412), .ZN(n8422) );
  INV_X1 U10811 ( .A(n8413), .ZN(n8415) );
  INV_X1 U10812 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n8414) );
  NAND2_X1 U10813 ( .A1(n8415), .A2(n8414), .ZN(n8417) );
  NAND2_X1 U10814 ( .A1(n8417), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8416) );
  MUX2_X1 U10815 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8416), .S(
        P2_IR_REG_5__SCAN_IN), .Z(n8420) );
  INV_X1 U10816 ( .A(n8417), .ZN(n8419) );
  NAND2_X1 U10817 ( .A1(n8419), .A2(n8418), .ZN(n8456) );
  AOI22_X1 U10818 ( .A1(n8680), .A2(P1_DATAO_REG_5__SCAN_IN), .B1(n8679), .B2(
        n10296), .ZN(n8421) );
  XNOR2_X1 U10819 ( .A(n12907), .B(n8382), .ZN(n8431) );
  NAND2_X1 U10820 ( .A1(n8942), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n8430) );
  NAND2_X1 U10821 ( .A1(n8336), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n8429) );
  INV_X1 U10822 ( .A(n8423), .ZN(n8443) );
  INV_X1 U10823 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n8425) );
  NAND2_X1 U10824 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n8424) );
  NAND2_X1 U10825 ( .A1(n8425), .A2(n8424), .ZN(n8426) );
  AND2_X1 U10826 ( .A1(n8443), .A2(n8426), .ZN(n11071) );
  NAND2_X1 U10827 ( .A1(n8817), .A2(n11071), .ZN(n8428) );
  NAND2_X1 U10828 ( .A1(n10131), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n8427) );
  NAND4_X1 U10829 ( .A1(n8430), .A2(n8429), .A3(n8428), .A4(n8427), .ZN(n13984) );
  NAND2_X1 U10830 ( .A1(n13984), .A2(n6670), .ZN(n8432) );
  NAND2_X1 U10831 ( .A1(n8431), .A2(n8432), .ZN(n8436) );
  INV_X1 U10832 ( .A(n8431), .ZN(n8434) );
  INV_X1 U10833 ( .A(n8432), .ZN(n8433) );
  NAND2_X1 U10834 ( .A1(n8434), .A2(n8433), .ZN(n8435) );
  AND2_X1 U10835 ( .A1(n8436), .A2(n8435), .ZN(n10535) );
  NAND2_X1 U10836 ( .A1(n10534), .A2(n10535), .ZN(n10533) );
  NAND2_X1 U10837 ( .A1(n11232), .A2(n8412), .ZN(n8441) );
  NAND2_X1 U10838 ( .A1(n8456), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8439) );
  XNOR2_X1 U10839 ( .A(n8439), .B(P2_IR_REG_6__SCAN_IN), .ZN(n15540) );
  AOI22_X1 U10840 ( .A1(n8680), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n8679), .B2(
        n15540), .ZN(n8440) );
  XNOR2_X1 U10841 ( .A(n15671), .B(n8382), .ZN(n8449) );
  NAND2_X1 U10842 ( .A1(n8941), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n8448) );
  NAND2_X1 U10843 ( .A1(n8942), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n8447) );
  INV_X1 U10844 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n8442) );
  NAND2_X1 U10845 ( .A1(n8443), .A2(n8442), .ZN(n8444) );
  AND2_X1 U10846 ( .A1(n8476), .A2(n8444), .ZN(n10568) );
  NAND2_X1 U10847 ( .A1(n8817), .A2(n10568), .ZN(n8446) );
  NAND2_X1 U10848 ( .A1(n10131), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n8445) );
  NAND2_X1 U10849 ( .A1(n13983), .A2(n6670), .ZN(n8450) );
  XNOR2_X1 U10850 ( .A(n8449), .B(n8450), .ZN(n10566) );
  INV_X1 U10851 ( .A(n8449), .ZN(n8452) );
  INV_X1 U10852 ( .A(n8450), .ZN(n8451) );
  NAND2_X1 U10853 ( .A1(n8452), .A2(n8451), .ZN(n8453) );
  NAND2_X1 U10854 ( .A1(n11343), .A2(n8412), .ZN(n8459) );
  OAI21_X1 U10855 ( .B1(n8456), .B2(P2_IR_REG_6__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n8457) );
  XNOR2_X1 U10856 ( .A(n8457), .B(P2_IR_REG_7__SCAN_IN), .ZN(n10143) );
  AOI22_X1 U10857 ( .A1(n8680), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n8679), .B2(
        n10143), .ZN(n8458) );
  NAND2_X2 U10858 ( .A1(n8459), .A2(n8458), .ZN(n12924) );
  XNOR2_X1 U10859 ( .A(n12924), .B(n8369), .ZN(n8466) );
  NAND2_X1 U10860 ( .A1(n8942), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n8463) );
  NAND2_X1 U10861 ( .A1(n10131), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n8462) );
  XNOR2_X1 U10862 ( .A(n8476), .B(P2_REG3_REG_7__SCAN_IN), .ZN(n11551) );
  NAND2_X1 U10863 ( .A1(n8817), .A2(n11551), .ZN(n8461) );
  NAND2_X1 U10864 ( .A1(n8941), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n8460) );
  NAND4_X1 U10865 ( .A1(n8463), .A2(n8462), .A3(n8461), .A4(n8460), .ZN(n13982) );
  NAND2_X1 U10866 ( .A1(n13982), .A2(n6670), .ZN(n8464) );
  XNOR2_X1 U10867 ( .A(n8466), .B(n8464), .ZN(n10721) );
  INV_X1 U10868 ( .A(n8464), .ZN(n8465) );
  NAND2_X1 U10869 ( .A1(n8466), .A2(n8465), .ZN(n8467) );
  XNOR2_X1 U10870 ( .A(n8469), .B(n8468), .ZN(n11395) );
  NAND2_X1 U10871 ( .A1(n11395), .A2(n8412), .ZN(n8473) );
  NAND2_X1 U10872 ( .A1(n8470), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8471) );
  XNOR2_X1 U10873 ( .A(n8471), .B(P2_IR_REG_8__SCAN_IN), .ZN(n10218) );
  AOI22_X1 U10874 ( .A1(n8680), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n8679), .B2(
        n10218), .ZN(n8472) );
  XNOR2_X1 U10875 ( .A(n12935), .B(n8382), .ZN(n8482) );
  NAND2_X1 U10876 ( .A1(n8941), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n8481) );
  NAND2_X1 U10877 ( .A1(n8942), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n8480) );
  INV_X1 U10878 ( .A(n8474), .ZN(n8494) );
  INV_X1 U10879 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n10080) );
  INV_X1 U10880 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n8475) );
  OAI21_X1 U10881 ( .B1(n8476), .B2(n10080), .A(n8475), .ZN(n8477) );
  AND2_X1 U10882 ( .A1(n8494), .A2(n8477), .ZN(n11135) );
  NAND2_X1 U10883 ( .A1(n8817), .A2(n11135), .ZN(n8479) );
  NAND2_X1 U10884 ( .A1(n10131), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n8478) );
  NAND4_X1 U10885 ( .A1(n8481), .A2(n8480), .A3(n8479), .A4(n8478), .ZN(n13981) );
  NAND2_X1 U10886 ( .A1(n13981), .A2(n6670), .ZN(n8483) );
  NAND2_X1 U10887 ( .A1(n8482), .A2(n8483), .ZN(n8487) );
  INV_X1 U10888 ( .A(n8482), .ZN(n8485) );
  INV_X1 U10889 ( .A(n8483), .ZN(n8484) );
  NAND2_X1 U10890 ( .A1(n8485), .A2(n8484), .ZN(n8486) );
  NAND2_X1 U10891 ( .A1(n11119), .A2(n8487), .ZN(n11265) );
  NAND2_X1 U10892 ( .A1(n11818), .A2(n8412), .ZN(n8493) );
  OR2_X1 U10893 ( .A1(n8490), .A2(n14381), .ZN(n8491) );
  XNOR2_X1 U10894 ( .A(n8491), .B(P2_IR_REG_9__SCAN_IN), .ZN(n10231) );
  AOI22_X1 U10895 ( .A1(n8680), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n8679), .B2(
        n10231), .ZN(n8492) );
  XNOR2_X1 U10896 ( .A(n12940), .B(n8382), .ZN(n8500) );
  NAND2_X1 U10897 ( .A1(n8941), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n8499) );
  NAND2_X1 U10898 ( .A1(n8942), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n8498) );
  INV_X1 U10899 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n11268) );
  NAND2_X1 U10900 ( .A1(n8494), .A2(n11268), .ZN(n8495) );
  AND2_X1 U10901 ( .A1(n8513), .A2(n8495), .ZN(n11271) );
  NAND2_X1 U10902 ( .A1(n8817), .A2(n11271), .ZN(n8497) );
  NAND2_X1 U10903 ( .A1(n10131), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n8496) );
  NAND4_X1 U10904 ( .A1(n8499), .A2(n8498), .A3(n8497), .A4(n8496), .ZN(n13980) );
  NAND2_X1 U10905 ( .A1(n13980), .A2(n6670), .ZN(n8501) );
  NAND2_X1 U10906 ( .A1(n8500), .A2(n8501), .ZN(n8505) );
  INV_X1 U10907 ( .A(n8500), .ZN(n8503) );
  INV_X1 U10908 ( .A(n8501), .ZN(n8502) );
  NAND2_X1 U10909 ( .A1(n8503), .A2(n8502), .ZN(n8504) );
  AND2_X1 U10910 ( .A1(n8505), .A2(n8504), .ZN(n11266) );
  NAND2_X1 U10911 ( .A1(n11265), .A2(n11266), .ZN(n11264) );
  XNOR2_X1 U10912 ( .A(n8506), .B(n8507), .ZN(n11934) );
  NAND2_X1 U10913 ( .A1(n11934), .A2(n8412), .ZN(n8511) );
  OR2_X1 U10914 ( .A1(n8508), .A2(n14381), .ZN(n8509) );
  XNOR2_X1 U10915 ( .A(n8509), .B(P2_IR_REG_10__SCAN_IN), .ZN(n10279) );
  AOI22_X1 U10916 ( .A1(n8680), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n8679), 
        .B2(n10279), .ZN(n8510) );
  XNOR2_X1 U10917 ( .A(n12947), .B(n8382), .ZN(n8520) );
  NAND2_X1 U10918 ( .A1(n8942), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n8518) );
  NAND2_X1 U10919 ( .A1(n8513), .A2(n8512), .ZN(n8514) );
  AND2_X1 U10920 ( .A1(n8529), .A2(n8514), .ZN(n11379) );
  NAND2_X1 U10921 ( .A1(n8817), .A2(n11379), .ZN(n8517) );
  NAND2_X1 U10922 ( .A1(n10131), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n8516) );
  NAND2_X1 U10923 ( .A1(n8941), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n8515) );
  NAND4_X1 U10924 ( .A1(n8518), .A2(n8517), .A3(n8516), .A4(n8515), .ZN(n13979) );
  NAND2_X1 U10925 ( .A1(n13979), .A2(n6670), .ZN(n8519) );
  XNOR2_X1 U10926 ( .A(n8520), .B(n8519), .ZN(n11307) );
  XNOR2_X1 U10927 ( .A(n8522), .B(n8523), .ZN(n12155) );
  NAND2_X1 U10928 ( .A1(n12155), .A2(n8412), .ZN(n8527) );
  INV_X1 U10929 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n8524) );
  NAND2_X1 U10930 ( .A1(n8508), .A2(n8524), .ZN(n8542) );
  NAND2_X1 U10931 ( .A1(n8542), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8525) );
  XNOR2_X1 U10932 ( .A(n8525), .B(P2_IR_REG_11__SCAN_IN), .ZN(n11679) );
  AOI22_X1 U10933 ( .A1(n8680), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n8679), 
        .B2(n11679), .ZN(n8526) );
  XNOR2_X1 U10934 ( .A(n15349), .B(n8382), .ZN(n8535) );
  NAND2_X1 U10935 ( .A1(n8942), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n8534) );
  NAND2_X1 U10936 ( .A1(n8529), .A2(n8528), .ZN(n8530) );
  NAND2_X1 U10937 ( .A1(n8548), .A2(n8530), .ZN(n15353) );
  INV_X1 U10938 ( .A(n15353), .ZN(n11630) );
  NAND2_X1 U10939 ( .A1(n8817), .A2(n11630), .ZN(n8533) );
  NAND2_X1 U10940 ( .A1(n10131), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n8532) );
  NAND2_X1 U10941 ( .A1(n8941), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n8531) );
  NAND4_X1 U10942 ( .A1(n8534), .A2(n8533), .A3(n8532), .A4(n8531), .ZN(n13978) );
  NAND2_X1 U10943 ( .A1(n13978), .A2(n6670), .ZN(n8536) );
  NAND2_X1 U10944 ( .A1(n8535), .A2(n8536), .ZN(n8540) );
  INV_X1 U10945 ( .A(n8535), .ZN(n8538) );
  INV_X1 U10946 ( .A(n8536), .ZN(n8537) );
  NAND2_X1 U10947 ( .A1(n8538), .A2(n8537), .ZN(n8539) );
  NAND2_X1 U10948 ( .A1(n8540), .A2(n8539), .ZN(n15342) );
  XNOR2_X1 U10949 ( .A(n8541), .B(n7735), .ZN(n12275) );
  NAND2_X1 U10950 ( .A1(n12275), .A2(n8412), .ZN(n8546) );
  NOR2_X1 U10951 ( .A1(n8542), .A2(P2_IR_REG_11__SCAN_IN), .ZN(n8563) );
  INV_X1 U10952 ( .A(n8563), .ZN(n8543) );
  NAND2_X1 U10953 ( .A1(n8543), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8544) );
  XNOR2_X1 U10954 ( .A(n8544), .B(P2_IR_REG_12__SCAN_IN), .ZN(n15555) );
  AOI22_X1 U10955 ( .A1(n8680), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n8679), 
        .B2(n15555), .ZN(n8545) );
  XNOR2_X1 U10956 ( .A(n12959), .B(n8382), .ZN(n8554) );
  NAND2_X1 U10957 ( .A1(n8941), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n8553) );
  NAND2_X1 U10958 ( .A1(n8942), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n8552) );
  INV_X1 U10959 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n8547) );
  NAND2_X1 U10960 ( .A1(n8548), .A2(n8547), .ZN(n8549) );
  AND2_X1 U10961 ( .A1(n8571), .A2(n8549), .ZN(n11714) );
  NAND2_X1 U10962 ( .A1(n8817), .A2(n11714), .ZN(n8551) );
  NAND2_X1 U10963 ( .A1(n10131), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n8550) );
  NAND4_X1 U10964 ( .A1(n8553), .A2(n8552), .A3(n8551), .A4(n8550), .ZN(n13977) );
  NAND2_X1 U10965 ( .A1(n13977), .A2(n6670), .ZN(n8555) );
  INV_X1 U10966 ( .A(n8554), .ZN(n8557) );
  INV_X1 U10967 ( .A(n8555), .ZN(n8556) );
  NAND2_X1 U10968 ( .A1(n8557), .A2(n8556), .ZN(n11699) );
  XNOR2_X1 U10969 ( .A(n8559), .B(n10016), .ZN(n8560) );
  XNOR2_X1 U10970 ( .A(n8561), .B(n8560), .ZN(n12326) );
  NAND2_X1 U10971 ( .A1(n12326), .A2(n8412), .ZN(n8570) );
  NAND2_X1 U10972 ( .A1(n8563), .A2(n8562), .ZN(n8565) );
  NAND2_X1 U10973 ( .A1(n8565), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8564) );
  MUX2_X1 U10974 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8564), .S(
        P2_IR_REG_13__SCAN_IN), .Z(n8568) );
  INV_X1 U10975 ( .A(n8565), .ZN(n8567) );
  INV_X1 U10976 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n8566) );
  NAND2_X1 U10977 ( .A1(n8567), .A2(n8566), .ZN(n8606) );
  AND2_X1 U10978 ( .A1(n8568), .A2(n8606), .ZN(n15568) );
  AOI22_X1 U10979 ( .A1(n8680), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n8679), 
        .B2(n15568), .ZN(n8569) );
  XNOR2_X1 U10980 ( .A(n12967), .B(n8369), .ZN(n8577) );
  NAND2_X1 U10981 ( .A1(n8942), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n8576) );
  NAND2_X1 U10982 ( .A1(n10131), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n8575) );
  INV_X1 U10983 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n11965) );
  NAND2_X1 U10984 ( .A1(n8571), .A2(n11965), .ZN(n8572) );
  AND2_X1 U10985 ( .A1(n8587), .A2(n8572), .ZN(n11968) );
  NAND2_X1 U10986 ( .A1(n8817), .A2(n11968), .ZN(n8574) );
  NAND2_X1 U10987 ( .A1(n8941), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n8573) );
  NAND4_X1 U10988 ( .A1(n8576), .A2(n8575), .A3(n8574), .A4(n8573), .ZN(n13976) );
  AND2_X1 U10989 ( .A1(n13976), .A2(n6670), .ZN(n8578) );
  NAND2_X1 U10990 ( .A1(n8577), .A2(n8578), .ZN(n8582) );
  INV_X1 U10991 ( .A(n8577), .ZN(n8580) );
  INV_X1 U10992 ( .A(n8578), .ZN(n8579) );
  NAND2_X1 U10993 ( .A1(n8580), .A2(n8579), .ZN(n8581) );
  AND2_X1 U10994 ( .A1(n8582), .A2(n8581), .ZN(n11963) );
  XNOR2_X1 U10995 ( .A(n8600), .B(SI_14_), .ZN(n8599) );
  INV_X1 U10996 ( .A(n8599), .ZN(n8583) );
  XNOR2_X1 U10997 ( .A(n8583), .B(n8597), .ZN(n12332) );
  NAND2_X1 U10998 ( .A1(n12332), .A2(n8412), .ZN(n8586) );
  NAND2_X1 U10999 ( .A1(n8606), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8584) );
  XNOR2_X1 U11000 ( .A(n8584), .B(P2_IR_REG_14__SCAN_IN), .ZN(n11669) );
  AOI22_X1 U11001 ( .A1(n8680), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n8679), 
        .B2(n11669), .ZN(n8585) );
  XNOR2_X1 U11002 ( .A(n12988), .B(n8369), .ZN(n8593) );
  NAND2_X1 U11003 ( .A1(n8942), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n8592) );
  NAND2_X1 U11004 ( .A1(n8941), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n8591) );
  NAND2_X1 U11005 ( .A1(n8587), .A2(n12132), .ZN(n8588) );
  AND2_X1 U11006 ( .A1(n8611), .A2(n8588), .ZN(n12135) );
  NAND2_X1 U11007 ( .A1(n8817), .A2(n12135), .ZN(n8590) );
  NAND2_X1 U11008 ( .A1(n10131), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n8589) );
  NAND4_X1 U11009 ( .A1(n8592), .A2(n8591), .A3(n8590), .A4(n8589), .ZN(n13975) );
  NAND2_X1 U11010 ( .A1(n13975), .A2(n6670), .ZN(n8594) );
  XNOR2_X1 U11011 ( .A(n8593), .B(n8594), .ZN(n12129) );
  INV_X1 U11012 ( .A(n8593), .ZN(n8595) );
  NAND2_X1 U11013 ( .A1(n8595), .A2(n8594), .ZN(n8596) );
  NAND2_X1 U11014 ( .A1(n12128), .A2(n8596), .ZN(n8617) );
  INV_X1 U11015 ( .A(n8597), .ZN(n8598) );
  NAND2_X1 U11016 ( .A1(n8599), .A2(n8598), .ZN(n8602) );
  INV_X1 U11017 ( .A(SI_14_), .ZN(n10029) );
  NAND2_X1 U11018 ( .A1(n8600), .A2(n10029), .ZN(n8601) );
  NAND2_X1 U11019 ( .A1(n8602), .A2(n8601), .ZN(n8605) );
  XNOR2_X1 U11020 ( .A(n8603), .B(n10130), .ZN(n8604) );
  XNOR2_X1 U11021 ( .A(n8605), .B(n8604), .ZN(n12345) );
  NAND2_X1 U11022 ( .A1(n12345), .A2(n8412), .ZN(n8609) );
  OAI21_X1 U11023 ( .B1(n8606), .B2(P2_IR_REG_14__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n8607) );
  XNOR2_X1 U11024 ( .A(n8607), .B(P2_IR_REG_15__SCAN_IN), .ZN(n15592) );
  AOI22_X1 U11025 ( .A1(n8680), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n15592), 
        .B2(n8679), .ZN(n8608) );
  NAND2_X2 U11026 ( .A1(n8609), .A2(n8608), .ZN(n12980) );
  XNOR2_X1 U11027 ( .A(n12980), .B(n8369), .ZN(n8618) );
  XNOR2_X1 U11028 ( .A(n8617), .B(n8618), .ZN(n12257) );
  NAND2_X1 U11029 ( .A1(n8941), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n8616) );
  NAND2_X1 U11030 ( .A1(n8942), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n8615) );
  INV_X1 U11031 ( .A(n8610), .ZN(n8630) );
  NAND2_X1 U11032 ( .A1(n8611), .A2(n12258), .ZN(n8612) );
  AND2_X1 U11033 ( .A1(n8630), .A2(n8612), .ZN(n12261) );
  NAND2_X1 U11034 ( .A1(n8817), .A2(n12261), .ZN(n8614) );
  NAND2_X1 U11035 ( .A1(n10131), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n8613) );
  NAND4_X1 U11036 ( .A1(n8616), .A2(n8615), .A3(n8614), .A4(n8613), .ZN(n13974) );
  AND2_X1 U11037 ( .A1(n13974), .A2(n6670), .ZN(n12256) );
  INV_X1 U11038 ( .A(n8617), .ZN(n8619) );
  NAND2_X1 U11039 ( .A1(n8619), .A2(n8618), .ZN(n8620) );
  XNOR2_X1 U11040 ( .A(n8622), .B(n8621), .ZN(n12394) );
  NAND2_X1 U11041 ( .A1(n12394), .A2(n8412), .ZN(n8627) );
  NAND2_X1 U11042 ( .A1(n8623), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8625) );
  XNOR2_X1 U11043 ( .A(n8625), .B(n8624), .ZN(n11690) );
  INV_X1 U11044 ( .A(n11690), .ZN(n15602) );
  AOI22_X1 U11045 ( .A1(n8680), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n8679), 
        .B2(n15602), .ZN(n8626) );
  XNOR2_X1 U11046 ( .A(n14376), .B(n8382), .ZN(n8637) );
  NAND2_X1 U11047 ( .A1(n8941), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n8635) );
  NAND2_X1 U11048 ( .A1(n8942), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n8634) );
  INV_X1 U11049 ( .A(n8628), .ZN(n8652) );
  INV_X1 U11050 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n8629) );
  NAND2_X1 U11051 ( .A1(n8630), .A2(n8629), .ZN(n8631) );
  AND2_X1 U11052 ( .A1(n8652), .A2(n8631), .ZN(n12207) );
  NAND2_X1 U11053 ( .A1(n8817), .A2(n12207), .ZN(n8633) );
  NAND2_X1 U11054 ( .A1(n10131), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n8632) );
  NAND4_X1 U11055 ( .A1(n8635), .A2(n8634), .A3(n8633), .A4(n8632), .ZN(n13973) );
  NAND2_X1 U11056 ( .A1(n13973), .A2(n6670), .ZN(n8636) );
  XNOR2_X1 U11057 ( .A(n8637), .B(n8636), .ZN(n13888) );
  NAND2_X1 U11058 ( .A1(n8637), .A2(n8636), .ZN(n13895) );
  XNOR2_X1 U11059 ( .A(n8638), .B(SI_17_), .ZN(n8639) );
  XNOR2_X1 U11060 ( .A(n8640), .B(n8639), .ZN(n12399) );
  NAND2_X1 U11061 ( .A1(n12399), .A2(n8412), .ZN(n8648) );
  INV_X1 U11062 ( .A(n8641), .ZN(n8642) );
  NAND2_X1 U11063 ( .A1(n8642), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8644) );
  MUX2_X1 U11064 ( .A(n8644), .B(P2_IR_REG_31__SCAN_IN), .S(n8643), .Z(n8646)
         );
  NAND2_X1 U11065 ( .A1(n8646), .A2(n8645), .ZN(n11884) );
  INV_X1 U11066 ( .A(n11884), .ZN(n11696) );
  AOI22_X1 U11067 ( .A1(n8680), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n8679), 
        .B2(n11696), .ZN(n8647) );
  NAND2_X2 U11068 ( .A1(n8648), .A2(n8647), .ZN(n14307) );
  XNOR2_X1 U11069 ( .A(n14307), .B(n8369), .ZN(n8656) );
  NAND2_X1 U11070 ( .A1(n8941), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n8650) );
  NAND2_X1 U11071 ( .A1(n8942), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n8649) );
  NAND2_X1 U11072 ( .A1(n8650), .A2(n8649), .ZN(n8655) );
  INV_X1 U11073 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n8651) );
  NAND2_X1 U11074 ( .A1(n8652), .A2(n8651), .ZN(n8653) );
  NAND2_X1 U11075 ( .A1(n8665), .A2(n8653), .ZN(n14225) );
  INV_X1 U11076 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n14308) );
  OAI22_X1 U11077 ( .A1(n14225), .A2(n8874), .B1(n8945), .B2(n14308), .ZN(
        n8654) );
  NAND2_X1 U11078 ( .A1(n13972), .A2(n6670), .ZN(n8657) );
  XNOR2_X1 U11079 ( .A(n8656), .B(n8657), .ZN(n13896) );
  INV_X1 U11080 ( .A(n8656), .ZN(n8658) );
  NAND2_X1 U11081 ( .A1(n8658), .A2(n8657), .ZN(n8659) );
  XNOR2_X1 U11082 ( .A(n8660), .B(n8661), .ZN(n12411) );
  NAND2_X1 U11083 ( .A1(n12411), .A2(n8412), .ZN(n8664) );
  NAND2_X1 U11084 ( .A1(n8645), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8662) );
  XNOR2_X1 U11085 ( .A(n8662), .B(P2_IR_REG_18__SCAN_IN), .ZN(n14004) );
  AOI22_X1 U11086 ( .A1(n8680), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n8679), 
        .B2(n14004), .ZN(n8663) );
  XNOR2_X1 U11087 ( .A(n14210), .B(n8369), .ZN(n8670) );
  NAND2_X1 U11088 ( .A1(n8665), .A2(n13942), .ZN(n8666) );
  NAND2_X1 U11089 ( .A1(n8684), .A2(n8666), .ZN(n13940) );
  AOI22_X1 U11090 ( .A1(n8941), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n8942), .B2(
        P2_REG0_REG_18__SCAN_IN), .ZN(n8669) );
  NAND2_X1 U11091 ( .A1(n10131), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n8668) );
  OAI211_X1 U11092 ( .C1(n13940), .C2(n8874), .A(n8669), .B(n8668), .ZN(n13971) );
  AND2_X1 U11093 ( .A1(n13971), .A2(n6670), .ZN(n8671) );
  NAND2_X1 U11094 ( .A1(n8670), .A2(n8671), .ZN(n8676) );
  INV_X1 U11095 ( .A(n8670), .ZN(n8673) );
  INV_X1 U11096 ( .A(n8671), .ZN(n8672) );
  NAND2_X1 U11097 ( .A1(n8673), .A2(n8672), .ZN(n8674) );
  NAND2_X1 U11098 ( .A1(n8676), .A2(n8674), .ZN(n13936) );
  XNOR2_X1 U11099 ( .A(n8678), .B(n8677), .ZN(n12414) );
  NAND2_X1 U11100 ( .A1(n12414), .A2(n8412), .ZN(n8682) );
  INV_X1 U11101 ( .A(n8859), .ZN(n13159) );
  AOI22_X1 U11102 ( .A1(n8680), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n13159), 
        .B2(n8679), .ZN(n8681) );
  XNOR2_X1 U11103 ( .A(n14295), .B(n8369), .ZN(n8688) );
  INV_X1 U11104 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n14296) );
  INV_X1 U11105 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n8683) );
  NAND2_X1 U11106 ( .A1(n8684), .A2(n8683), .ZN(n8685) );
  NAND2_X1 U11107 ( .A1(n8694), .A2(n8685), .ZN(n14188) );
  OR2_X1 U11108 ( .A1(n14188), .A2(n8874), .ZN(n8687) );
  AOI22_X1 U11109 ( .A1(n8941), .A2(P2_REG2_REG_19__SCAN_IN), .B1(n8942), .B2(
        P2_REG0_REG_19__SCAN_IN), .ZN(n8686) );
  OAI211_X1 U11110 ( .C1(n8945), .C2(n14296), .A(n8687), .B(n8686), .ZN(n13970) );
  NAND2_X1 U11111 ( .A1(n13970), .A2(n6670), .ZN(n8689) );
  XNOR2_X1 U11112 ( .A(n8688), .B(n8689), .ZN(n13860) );
  NAND2_X1 U11113 ( .A1(n13861), .A2(n13860), .ZN(n13859) );
  INV_X1 U11114 ( .A(n8688), .ZN(n8690) );
  NAND2_X1 U11115 ( .A1(n8690), .A2(n8689), .ZN(n13919) );
  NAND2_X1 U11116 ( .A1(n13859), .A2(n13919), .ZN(n8702) );
  XNOR2_X1 U11117 ( .A(n8710), .B(n10924), .ZN(n8707) );
  XNOR2_X1 U11118 ( .A(n8707), .B(n8708), .ZN(n12425) );
  NAND2_X1 U11119 ( .A1(n12425), .A2(n8412), .ZN(n8692) );
  OR2_X1 U11120 ( .A1(n8379), .A2(n11848), .ZN(n8691) );
  NAND2_X2 U11121 ( .A1(n8692), .A2(n8691), .ZN(n14289) );
  XNOR2_X1 U11122 ( .A(n14289), .B(n8369), .ZN(n8703) );
  INV_X1 U11123 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n8693) );
  NAND2_X1 U11124 ( .A1(n8694), .A2(n8693), .ZN(n8695) );
  NAND2_X1 U11125 ( .A1(n8718), .A2(n8695), .ZN(n14173) );
  OR2_X1 U11126 ( .A1(n14173), .A2(n8874), .ZN(n8701) );
  INV_X1 U11127 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n8698) );
  NAND2_X1 U11128 ( .A1(n8942), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n8697) );
  NAND2_X1 U11129 ( .A1(n8941), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n8696) );
  OAI211_X1 U11130 ( .C1(n8945), .C2(n8698), .A(n8697), .B(n8696), .ZN(n8699)
         );
  INV_X1 U11131 ( .A(n8699), .ZN(n8700) );
  NAND2_X1 U11132 ( .A1(n8701), .A2(n8700), .ZN(n13969) );
  NAND2_X1 U11133 ( .A1(n13969), .A2(n6670), .ZN(n8704) );
  XNOR2_X1 U11134 ( .A(n8703), .B(n8704), .ZN(n13918) );
  INV_X1 U11135 ( .A(n8703), .ZN(n8705) );
  NAND2_X1 U11136 ( .A1(n8705), .A2(n8704), .ZN(n8706) );
  INV_X1 U11137 ( .A(n8707), .ZN(n8709) );
  NAND2_X1 U11138 ( .A1(n8709), .A2(n8708), .ZN(n8712) );
  OR2_X1 U11139 ( .A1(n8710), .A2(n10924), .ZN(n8711) );
  NAND2_X1 U11140 ( .A1(n8712), .A2(n8711), .ZN(n8715) );
  XNOR2_X1 U11141 ( .A(n8713), .B(SI_21_), .ZN(n8714) );
  OR2_X1 U11142 ( .A1(n8379), .A2(n11960), .ZN(n8716) );
  XNOR2_X1 U11143 ( .A(n14285), .B(n8369), .ZN(n8725) );
  NAND2_X1 U11144 ( .A1(n8718), .A2(n13874), .ZN(n8719) );
  NAND2_X1 U11145 ( .A1(n8746), .A2(n8719), .ZN(n13873) );
  OR2_X1 U11146 ( .A1(n13873), .A2(n8874), .ZN(n8724) );
  INV_X1 U11147 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n14286) );
  NAND2_X1 U11148 ( .A1(n8941), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n8721) );
  NAND2_X1 U11149 ( .A1(n8942), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n8720) );
  OAI211_X1 U11150 ( .C1(n14286), .C2(n8945), .A(n8721), .B(n8720), .ZN(n8722)
         );
  INV_X1 U11151 ( .A(n8722), .ZN(n8723) );
  NAND2_X1 U11152 ( .A1(n8724), .A2(n8723), .ZN(n13968) );
  AND2_X1 U11153 ( .A1(n13968), .A2(n6670), .ZN(n8726) );
  NAND2_X1 U11154 ( .A1(n8725), .A2(n8726), .ZN(n8731) );
  INV_X1 U11155 ( .A(n8725), .ZN(n8728) );
  INV_X1 U11156 ( .A(n8726), .ZN(n8727) );
  NAND2_X1 U11157 ( .A1(n8728), .A2(n8727), .ZN(n8729) );
  NAND2_X1 U11158 ( .A1(n8731), .A2(n8729), .ZN(n13869) );
  INV_X1 U11159 ( .A(n13869), .ZN(n8730) );
  XNOR2_X1 U11160 ( .A(n8732), .B(n8733), .ZN(n12858) );
  NAND2_X1 U11161 ( .A1(n12858), .A2(n8412), .ZN(n8735) );
  INV_X1 U11162 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n12860) );
  OR2_X1 U11163 ( .A1(n8379), .A2(n12860), .ZN(n8734) );
  XNOR2_X1 U11164 ( .A(n8746), .B(P2_REG3_REG_22__SCAN_IN), .ZN(n14145) );
  NAND2_X1 U11165 ( .A1(n14145), .A2(n8817), .ZN(n8740) );
  INV_X1 U11166 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n14280) );
  NAND2_X1 U11167 ( .A1(n8941), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n8737) );
  NAND2_X1 U11168 ( .A1(n8942), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n8736) );
  OAI211_X1 U11169 ( .C1(n14280), .C2(n8945), .A(n8737), .B(n8736), .ZN(n8738)
         );
  INV_X1 U11170 ( .A(n8738), .ZN(n8739) );
  NAND2_X1 U11171 ( .A1(n8740), .A2(n8739), .ZN(n13967) );
  AND2_X1 U11172 ( .A1(n13967), .A2(n6670), .ZN(n13928) );
  NAND2_X1 U11173 ( .A1(n13926), .A2(n13928), .ZN(n8741) );
  XNOR2_X1 U11174 ( .A(n8743), .B(n8742), .ZN(n12457) );
  NAND2_X1 U11175 ( .A1(n12457), .A2(n8412), .ZN(n8745) );
  INV_X1 U11176 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n12060) );
  OR2_X1 U11177 ( .A1(n8379), .A2(n12060), .ZN(n8744) );
  XNOR2_X1 U11178 ( .A(n14274), .B(n8369), .ZN(n8755) );
  INV_X1 U11179 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n13930) );
  INV_X1 U11180 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n13854) );
  OAI21_X1 U11181 ( .B1(n8746), .B2(n13930), .A(n13854), .ZN(n8747) );
  AND2_X1 U11182 ( .A1(n8761), .A2(n8747), .ZN(n14129) );
  NAND2_X1 U11183 ( .A1(n14129), .A2(n8817), .ZN(n8752) );
  INV_X1 U11184 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n14275) );
  NAND2_X1 U11185 ( .A1(n8941), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n8749) );
  NAND2_X1 U11186 ( .A1(n8942), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n8748) );
  OAI211_X1 U11187 ( .C1(n14275), .C2(n8945), .A(n8749), .B(n8748), .ZN(n8750)
         );
  INV_X1 U11188 ( .A(n8750), .ZN(n8751) );
  NAND2_X1 U11189 ( .A1(n8752), .A2(n8751), .ZN(n13966) );
  INV_X1 U11190 ( .A(n13966), .ZN(n13048) );
  NOR2_X1 U11191 ( .A1(n13048), .A2(n14206), .ZN(n13853) );
  XNOR2_X1 U11192 ( .A(n8756), .B(n8757), .ZN(n12468) );
  NAND2_X1 U11193 ( .A1(n12468), .A2(n8412), .ZN(n8759) );
  INV_X1 U11194 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n12324) );
  OR2_X1 U11195 ( .A1(n8379), .A2(n12324), .ZN(n8758) );
  XNOR2_X1 U11196 ( .A(n14343), .B(n8369), .ZN(n8769) );
  INV_X1 U11197 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n8760) );
  NAND2_X1 U11198 ( .A1(n8761), .A2(n8760), .ZN(n8762) );
  NAND2_X1 U11199 ( .A1(n8775), .A2(n8762), .ZN(n14110) );
  OR2_X1 U11200 ( .A1(n14110), .A2(n8874), .ZN(n8767) );
  INV_X1 U11201 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n14267) );
  NAND2_X1 U11202 ( .A1(n8941), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n8764) );
  NAND2_X1 U11203 ( .A1(n8942), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n8763) );
  OAI211_X1 U11204 ( .C1(n14267), .C2(n8945), .A(n8764), .B(n8763), .ZN(n8765)
         );
  INV_X1 U11205 ( .A(n8765), .ZN(n8766) );
  NAND2_X1 U11206 ( .A1(n8767), .A2(n8766), .ZN(n13965) );
  AND2_X1 U11207 ( .A1(n13965), .A2(n6670), .ZN(n8768) );
  NAND2_X1 U11208 ( .A1(n8769), .A2(n8768), .ZN(n8770) );
  OAI21_X1 U11209 ( .B1(n8769), .B2(n8768), .A(n8770), .ZN(n13909) );
  XNOR2_X1 U11210 ( .A(n8772), .B(n8771), .ZN(n12480) );
  NAND2_X1 U11211 ( .A1(n12480), .A2(n8412), .ZN(n8774) );
  OR2_X1 U11212 ( .A1(n8379), .A2(n12390), .ZN(n8773) );
  XNOR2_X1 U11213 ( .A(n14262), .B(n8369), .ZN(n8782) );
  XNOR2_X1 U11214 ( .A(n8775), .B(P2_REG3_REG_25__SCAN_IN), .ZN(n14093) );
  NAND2_X1 U11215 ( .A1(n14093), .A2(n8817), .ZN(n8780) );
  INV_X1 U11216 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n14263) );
  NAND2_X1 U11217 ( .A1(n8942), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n8777) );
  NAND2_X1 U11218 ( .A1(n8941), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n8776) );
  OAI211_X1 U11219 ( .C1(n14263), .C2(n8945), .A(n8777), .B(n8776), .ZN(n8778)
         );
  INV_X1 U11220 ( .A(n8778), .ZN(n8779) );
  NAND2_X1 U11221 ( .A1(n8780), .A2(n8779), .ZN(n13964) );
  AND2_X1 U11222 ( .A1(n13964), .A2(n6670), .ZN(n8781) );
  NAND2_X1 U11223 ( .A1(n8782), .A2(n8781), .ZN(n8783) );
  OAI21_X1 U11224 ( .B1(n8782), .B2(n8781), .A(n8783), .ZN(n13879) );
  NOR2_X1 U11225 ( .A1(n13880), .A2(n13879), .ZN(n13878) );
  INV_X1 U11226 ( .A(n8783), .ZN(n8784) );
  XNOR2_X1 U11227 ( .A(n8786), .B(n8785), .ZN(n13948) );
  MUX2_X1 U11228 ( .A(n7339), .B(n12567), .S(n9950), .Z(n8806) );
  XNOR2_X1 U11229 ( .A(n8806), .B(SI_27_), .ZN(n8790) );
  XNOR2_X1 U11230 ( .A(n8809), .B(n8790), .ZN(n12555) );
  NAND2_X1 U11231 ( .A1(n12555), .A2(n8412), .ZN(n8792) );
  OR2_X1 U11232 ( .A1(n8379), .A2(n12567), .ZN(n8791) );
  XNOR2_X1 U11233 ( .A(n14329), .B(n8369), .ZN(n8803) );
  NAND2_X1 U11234 ( .A1(n8793), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n8815) );
  INV_X1 U11235 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n8794) );
  NAND2_X1 U11236 ( .A1(n8795), .A2(n8794), .ZN(n8796) );
  NAND2_X1 U11237 ( .A1(n8815), .A2(n8796), .ZN(n12849) );
  OR2_X1 U11238 ( .A1(n12849), .A2(n8874), .ZN(n8801) );
  INV_X1 U11239 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n14251) );
  NAND2_X1 U11240 ( .A1(n8942), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n8798) );
  NAND2_X1 U11241 ( .A1(n8941), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n8797) );
  OAI211_X1 U11242 ( .C1(n8945), .C2(n14251), .A(n8798), .B(n8797), .ZN(n8799)
         );
  INV_X1 U11243 ( .A(n8799), .ZN(n8800) );
  NAND2_X1 U11244 ( .A1(n8801), .A2(n8800), .ZN(n13962) );
  AND2_X1 U11245 ( .A1(n13962), .A2(n6670), .ZN(n8802) );
  NAND2_X1 U11246 ( .A1(n8803), .A2(n8802), .ZN(n8804) );
  OAI21_X1 U11247 ( .B1(n8803), .B2(n8802), .A(n8804), .ZN(n12846) );
  INV_X1 U11248 ( .A(n8804), .ZN(n8805) );
  NOR2_X1 U11249 ( .A1(n8807), .A2(SI_27_), .ZN(n8808) );
  INV_X1 U11250 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n14392) );
  MUX2_X1 U11251 ( .A(n15236), .B(n14392), .S(n9950), .Z(n8810) );
  NAND2_X1 U11252 ( .A1(n8810), .A2(n8127), .ZN(n8881) );
  INV_X1 U11253 ( .A(n8810), .ZN(n8811) );
  NAND2_X1 U11254 ( .A1(n8811), .A2(SI_28_), .ZN(n8812) );
  NAND2_X1 U11255 ( .A1(n8881), .A2(n8812), .ZN(n8882) );
  NAND2_X1 U11256 ( .A1(n15235), .A2(n8412), .ZN(n8814) );
  OR2_X1 U11257 ( .A1(n8379), .A2(n14392), .ZN(n8813) );
  INV_X1 U11258 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n8877) );
  NAND2_X1 U11259 ( .A1(n8815), .A2(n8877), .ZN(n8816) );
  NAND2_X1 U11260 ( .A1(n14049), .A2(n8817), .ZN(n8823) );
  INV_X1 U11261 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n8820) );
  NAND2_X1 U11262 ( .A1(n8941), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n8819) );
  NAND2_X1 U11263 ( .A1(n8942), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n8818) );
  OAI211_X1 U11264 ( .C1(n8820), .C2(n8945), .A(n8819), .B(n8818), .ZN(n8821)
         );
  INV_X1 U11265 ( .A(n8821), .ZN(n8822) );
  NAND2_X1 U11266 ( .A1(n8823), .A2(n8822), .ZN(n13961) );
  NAND2_X1 U11267 ( .A1(n13961), .A2(n6670), .ZN(n8824) );
  XOR2_X1 U11268 ( .A(n8369), .B(n8824), .Z(n8825) );
  XNOR2_X1 U11269 ( .A(n14247), .B(n8825), .ZN(n8826) );
  NOR2_X1 U11270 ( .A1(n8831), .A2(n14381), .ZN(n8828) );
  MUX2_X1 U11271 ( .A(n14381), .B(n8828), .S(P2_IR_REG_24__SCAN_IN), .Z(n8829)
         );
  XNOR2_X1 U11272 ( .A(n12322), .B(P2_B_REG_SCAN_IN), .ZN(n8835) );
  NAND2_X1 U11273 ( .A1(n8836), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8834) );
  NAND2_X1 U11274 ( .A1(n8835), .A2(n12388), .ZN(n8840) );
  INV_X1 U11275 ( .A(n14395), .ZN(n8839) );
  INV_X1 U11276 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n15631) );
  NAND2_X1 U11277 ( .A1(n15628), .A2(n15631), .ZN(n8842) );
  AND2_X1 U11278 ( .A1(n14395), .A2(n12322), .ZN(n15632) );
  INV_X1 U11279 ( .A(n15632), .ZN(n8841) );
  NAND2_X1 U11280 ( .A1(n8842), .A2(n8841), .ZN(n8995) );
  NOR2_X1 U11281 ( .A1(P2_D_REG_2__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .ZN(
        n8846) );
  NOR4_X1 U11282 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        P2_D_REG_4__SCAN_IN), .A4(P2_D_REG_5__SCAN_IN), .ZN(n8845) );
  NOR4_X1 U11283 ( .A1(P2_D_REG_10__SCAN_IN), .A2(P2_D_REG_11__SCAN_IN), .A3(
        P2_D_REG_12__SCAN_IN), .A4(P2_D_REG_13__SCAN_IN), .ZN(n8844) );
  NOR4_X1 U11284 ( .A1(P2_D_REG_6__SCAN_IN), .A2(P2_D_REG_7__SCAN_IN), .A3(
        P2_D_REG_8__SCAN_IN), .A4(P2_D_REG_9__SCAN_IN), .ZN(n8843) );
  AND4_X1 U11285 ( .A1(n8846), .A2(n8845), .A3(n8844), .A4(n8843), .ZN(n8852)
         );
  NOR4_X1 U11286 ( .A1(P2_D_REG_18__SCAN_IN), .A2(P2_D_REG_19__SCAN_IN), .A3(
        P2_D_REG_20__SCAN_IN), .A4(P2_D_REG_21__SCAN_IN), .ZN(n8850) );
  NOR4_X1 U11287 ( .A1(P2_D_REG_16__SCAN_IN), .A2(P2_D_REG_14__SCAN_IN), .A3(
        P2_D_REG_15__SCAN_IN), .A4(P2_D_REG_17__SCAN_IN), .ZN(n8849) );
  NOR4_X1 U11288 ( .A1(P2_D_REG_26__SCAN_IN), .A2(P2_D_REG_27__SCAN_IN), .A3(
        P2_D_REG_28__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n8848) );
  NOR4_X1 U11289 ( .A1(P2_D_REG_22__SCAN_IN), .A2(P2_D_REG_23__SCAN_IN), .A3(
        P2_D_REG_24__SCAN_IN), .A4(P2_D_REG_25__SCAN_IN), .ZN(n8847) );
  AND4_X1 U11290 ( .A1(n8850), .A2(n8849), .A3(n8848), .A4(n8847), .ZN(n8851)
         );
  NAND2_X1 U11291 ( .A1(n8852), .A2(n8851), .ZN(n8853) );
  AND2_X1 U11292 ( .A1(n15628), .A2(n8853), .ZN(n8994) );
  INV_X1 U11293 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n15634) );
  AND2_X1 U11294 ( .A1(n14395), .A2(n12388), .ZN(n8854) );
  AOI21_X1 U11295 ( .B1(n15628), .B2(n15634), .A(n8854), .ZN(n8867) );
  INV_X1 U11296 ( .A(n8855), .ZN(n8856) );
  NAND2_X1 U11297 ( .A1(n8856), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8858) );
  NAND2_X1 U11298 ( .A1(n8867), .A2(n15635), .ZN(n15633) );
  OR2_X1 U11299 ( .A1(n8952), .A2(n15633), .ZN(n8864) );
  INV_X1 U11300 ( .A(n8864), .ZN(n8876) );
  NAND2_X1 U11301 ( .A1(n8859), .A2(n11849), .ZN(n13157) );
  INV_X1 U11302 ( .A(n8860), .ZN(n8861) );
  NAND2_X1 U11303 ( .A1(n13157), .A2(n8861), .ZN(n15644) );
  INV_X1 U11304 ( .A(n10075), .ZN(n8862) );
  AND2_X1 U11305 ( .A1(n15644), .A2(n8862), .ZN(n8863) );
  OR2_X1 U11306 ( .A1(n8860), .A2(n11849), .ZN(n11069) );
  NAND2_X1 U11307 ( .A1(n13159), .A2(n11849), .ZN(n15620) );
  INV_X1 U11308 ( .A(n8865), .ZN(n8866) );
  OAI21_X2 U11309 ( .B1(n8864), .B2(n11069), .A(n15621), .ZN(n15350) );
  NAND2_X1 U11310 ( .A1(n14247), .A2(n15350), .ZN(n8880) );
  NAND2_X1 U11311 ( .A1(n8952), .A2(n8865), .ZN(n8869) );
  OR2_X1 U11312 ( .A1(n8867), .A2(n8866), .ZN(n8950) );
  NAND2_X1 U11313 ( .A1(n13157), .A2(n10075), .ZN(n8951) );
  NAND4_X1 U11314 ( .A1(n8869), .A2(n8868), .A3(n8950), .A4(n8951), .ZN(n10353) );
  NAND2_X1 U11315 ( .A1(n10353), .A2(P2_STATE_REG_SCAN_IN), .ZN(n15354) );
  INV_X1 U11316 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n8954) );
  NAND2_X1 U11317 ( .A1(n8941), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n8871) );
  NAND2_X1 U11318 ( .A1(n8942), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n8870) );
  OAI211_X1 U11319 ( .C1(n8954), .C2(n8945), .A(n8871), .B(n8870), .ZN(n8872)
         );
  INV_X1 U11320 ( .A(n8872), .ZN(n8873) );
  OAI21_X1 U11321 ( .B1(n14032), .B2(n8874), .A(n8873), .ZN(n13960) );
  INV_X1 U11322 ( .A(n13952), .ZN(n13915) );
  INV_X1 U11323 ( .A(n13915), .ZN(n12105) );
  INV_X1 U11324 ( .A(n8875), .ZN(n10081) );
  AOI22_X1 U11325 ( .A1(n13960), .A2(n12105), .B1(n13962), .B2(n13951), .ZN(
        n14045) );
  INV_X1 U11326 ( .A(n13157), .ZN(n13166) );
  OAI22_X1 U11327 ( .A1(n14045), .A2(n13953), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8877), .ZN(n8878) );
  AOI21_X1 U11328 ( .B1(n14049), .B2(n13944), .A(n8878), .ZN(n8879) );
  MUX2_X1 U11329 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(P1_DATAO_REG_29__SCAN_IN), 
        .S(n9950), .Z(n12558) );
  XNOR2_X1 U11330 ( .A(n12558), .B(n13841), .ZN(n12556) );
  NAND2_X1 U11331 ( .A1(n14386), .A2(n8412), .ZN(n8885) );
  INV_X1 U11332 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n14387) );
  OR2_X1 U11333 ( .A1(n8379), .A2(n14387), .ZN(n8884) );
  INV_X1 U11334 ( .A(n14329), .ZN(n14068) );
  NAND2_X1 U11335 ( .A1(n8887), .A2(n15616), .ZN(n11653) );
  OR2_X1 U11336 ( .A1(n11653), .A2(n12882), .ZN(n11157) );
  NOR2_X2 U11337 ( .A1(n11157), .A2(n15652), .ZN(n11511) );
  INV_X1 U11338 ( .A(n15659), .ZN(n11510) );
  NAND2_X1 U11339 ( .A1(n11511), .A2(n11510), .ZN(n11509) );
  OR2_X2 U11340 ( .A1(n11509), .A2(n12907), .ZN(n11113) );
  OR2_X1 U11341 ( .A1(n11113), .A2(n15671), .ZN(n11111) );
  NOR2_X2 U11342 ( .A1(n11111), .A2(n12924), .ZN(n11091) );
  INV_X1 U11343 ( .A(n12935), .ZN(n11137) );
  NAND2_X1 U11344 ( .A1(n11091), .A2(n11137), .ZN(n11150) );
  OR2_X2 U11345 ( .A1(n11150), .A2(n12940), .ZN(n11368) );
  INV_X1 U11346 ( .A(n15349), .ZN(n11783) );
  INV_X1 U11347 ( .A(n12959), .ZN(n15363) );
  INV_X1 U11348 ( .A(n14307), .ZN(n14229) );
  INV_X1 U11349 ( .A(n14274), .ZN(n14132) );
  INV_X1 U11350 ( .A(n13120), .ZN(n8890) );
  NAND2_X1 U11351 ( .A1(n8890), .A2(n11654), .ZN(n8893) );
  INV_X1 U11352 ( .A(n12874), .ZN(n8891) );
  NAND2_X1 U11353 ( .A1(n8891), .A2(n8886), .ZN(n8892) );
  INV_X1 U11354 ( .A(n13986), .ZN(n8957) );
  NAND2_X1 U11355 ( .A1(n8957), .A2(n15652), .ZN(n8896) );
  NAND2_X1 U11356 ( .A1(n11158), .A2(n13986), .ZN(n8895) );
  NAND2_X1 U11357 ( .A1(n8896), .A2(n8895), .ZN(n13124) );
  NAND2_X1 U11358 ( .A1(n11161), .A2(n11162), .ZN(n11160) );
  INV_X1 U11359 ( .A(n13985), .ZN(n10538) );
  NAND2_X1 U11360 ( .A1(n15659), .A2(n10538), .ZN(n8898) );
  OR2_X1 U11361 ( .A1(n10538), .A2(n15659), .ZN(n8897) );
  INV_X1 U11362 ( .A(n13126), .ZN(n11515) );
  NAND2_X1 U11363 ( .A1(n11518), .A2(n8898), .ZN(n10911) );
  INV_X1 U11364 ( .A(n13984), .ZN(n12909) );
  NAND2_X1 U11365 ( .A1(n12907), .A2(n12909), .ZN(n8900) );
  OR2_X1 U11366 ( .A1(n12907), .A2(n12909), .ZN(n8899) );
  NAND2_X1 U11367 ( .A1(n8900), .A2(n8899), .ZN(n13127) );
  INV_X1 U11368 ( .A(n13127), .ZN(n10912) );
  INV_X1 U11369 ( .A(n13983), .ZN(n10537) );
  NAND2_X1 U11370 ( .A1(n15671), .A2(n10537), .ZN(n8901) );
  INV_X1 U11371 ( .A(n13982), .ZN(n12926) );
  OR2_X1 U11372 ( .A1(n12924), .A2(n12926), .ZN(n8902) );
  NAND2_X1 U11373 ( .A1(n12924), .A2(n12926), .ZN(n8903) );
  INV_X1 U11374 ( .A(n13981), .ZN(n8904) );
  NAND2_X1 U11375 ( .A1(n12935), .A2(n8904), .ZN(n8905) );
  NAND2_X1 U11376 ( .A1(n8906), .A2(n8905), .ZN(n11145) );
  INV_X1 U11377 ( .A(n13980), .ZN(n8907) );
  XNOR2_X1 U11378 ( .A(n12940), .B(n8907), .ZN(n13133) );
  INV_X1 U11379 ( .A(n13133), .ZN(n11144) );
  INV_X1 U11380 ( .A(n13979), .ZN(n12949) );
  XNOR2_X1 U11381 ( .A(n12947), .B(n12949), .ZN(n13134) );
  OR2_X1 U11382 ( .A1(n12947), .A2(n12949), .ZN(n8909) );
  INV_X1 U11383 ( .A(n13978), .ZN(n8910) );
  XNOR2_X1 U11384 ( .A(n15349), .B(n8910), .ZN(n13135) );
  NAND2_X1 U11385 ( .A1(n15349), .A2(n8910), .ZN(n8911) );
  XNOR2_X1 U11386 ( .A(n12959), .B(n13977), .ZN(n13136) );
  INV_X1 U11387 ( .A(n13977), .ZN(n12961) );
  NAND2_X1 U11388 ( .A1(n12959), .A2(n12961), .ZN(n8912) );
  XNOR2_X1 U11389 ( .A(n12967), .B(n13976), .ZN(n13137) );
  INV_X1 U11390 ( .A(n13137), .ZN(n11804) );
  INV_X1 U11391 ( .A(n13976), .ZN(n8977) );
  OR2_X1 U11392 ( .A1(n12967), .A2(n8977), .ZN(n8914) );
  INV_X1 U11393 ( .A(n13975), .ZN(n8915) );
  XNOR2_X1 U11394 ( .A(n12988), .B(n8915), .ZN(n13141) );
  NAND2_X1 U11395 ( .A1(n12988), .A2(n8915), .ZN(n8916) );
  INV_X1 U11396 ( .A(n13974), .ZN(n8917) );
  NAND2_X1 U11397 ( .A1(n12980), .A2(n8917), .ZN(n8918) );
  XNOR2_X1 U11398 ( .A(n14376), .B(n13973), .ZN(n13139) );
  INV_X1 U11399 ( .A(n13973), .ZN(n8919) );
  OR2_X1 U11400 ( .A1(n14376), .A2(n8919), .ZN(n8920) );
  INV_X1 U11401 ( .A(n13972), .ZN(n8982) );
  NAND2_X1 U11402 ( .A1(n14307), .A2(n8982), .ZN(n8921) );
  OR2_X1 U11403 ( .A1(n14307), .A2(n8982), .ZN(n8922) );
  INV_X1 U11404 ( .A(n13971), .ZN(n13863) );
  NAND2_X1 U11405 ( .A1(n14210), .A2(n13863), .ZN(n8923) );
  INV_X1 U11406 ( .A(n13970), .ZN(n13914) );
  INV_X1 U11407 ( .A(n13969), .ZN(n13864) );
  NAND2_X1 U11408 ( .A1(n14289), .A2(n13864), .ZN(n8926) );
  OR2_X1 U11409 ( .A1(n14289), .A2(n13864), .ZN(n8925) );
  OR2_X1 U11410 ( .A1(n14285), .A2(n13916), .ZN(n8927) );
  INV_X1 U11411 ( .A(n13967), .ZN(n8928) );
  XNOR2_X1 U11412 ( .A(n14351), .B(n8928), .ZN(n13145) );
  OR2_X1 U11413 ( .A1(n14351), .A2(n8928), .ZN(n8929) );
  NAND2_X1 U11414 ( .A1(n14274), .A2(n13048), .ZN(n8987) );
  INV_X1 U11415 ( .A(n13965), .ZN(n8930) );
  XNOR2_X1 U11416 ( .A(n14262), .B(n13964), .ZN(n13146) );
  NAND2_X1 U11417 ( .A1(n14085), .A2(n13146), .ZN(n8932) );
  NAND2_X1 U11418 ( .A1(n14262), .A2(n7536), .ZN(n8931) );
  INV_X1 U11419 ( .A(n13963), .ZN(n8989) );
  OR2_X1 U11420 ( .A1(n14256), .A2(n8989), .ZN(n13118) );
  NAND2_X1 U11421 ( .A1(n14081), .A2(n13118), .ZN(n8933) );
  NAND2_X1 U11422 ( .A1(n14256), .A2(n8989), .ZN(n13117) );
  NAND2_X1 U11423 ( .A1(n8933), .A2(n13117), .ZN(n14058) );
  INV_X1 U11424 ( .A(n13962), .ZN(n8990) );
  XNOR2_X1 U11425 ( .A(n14329), .B(n8990), .ZN(n13149) );
  INV_X1 U11426 ( .A(n13961), .ZN(n8947) );
  OR2_X1 U11427 ( .A1(n14247), .A2(n8947), .ZN(n8935) );
  NAND2_X1 U11428 ( .A1(n14247), .A2(n8947), .ZN(n8934) );
  NAND2_X1 U11429 ( .A1(n8935), .A2(n8934), .ZN(n14041) );
  NAND2_X1 U11430 ( .A1(n14329), .A2(n8990), .ZN(n14044) );
  NAND3_X1 U11431 ( .A1(n14056), .A2(n7171), .A3(n14044), .ZN(n14043) );
  NAND2_X1 U11432 ( .A1(n14043), .A2(n8935), .ZN(n8936) );
  XNOR2_X1 U11433 ( .A(n14031), .B(n13960), .ZN(n13152) );
  NAND2_X1 U11434 ( .A1(n13159), .A2(n13169), .ZN(n8937) );
  NAND2_X1 U11435 ( .A1(n8321), .A2(n13122), .ZN(n13162) );
  INV_X1 U11436 ( .A(n13951), .ZN(n13913) );
  INV_X1 U11437 ( .A(P2_B_REG_SCAN_IN), .ZN(n8939) );
  OR2_X1 U11438 ( .A1(n8938), .A2(n8939), .ZN(n8940) );
  NAND2_X1 U11439 ( .A1(n13952), .A2(n8940), .ZN(n14022) );
  INV_X1 U11440 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n14243) );
  NAND2_X1 U11441 ( .A1(n8941), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n8944) );
  NAND2_X1 U11442 ( .A1(n8942), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n8943) );
  OAI211_X1 U11443 ( .C1(n8945), .C2(n14243), .A(n8944), .B(n8943), .ZN(n13959) );
  INV_X1 U11444 ( .A(n13959), .ZN(n8946) );
  INV_X1 U11445 ( .A(n15635), .ZN(n15629) );
  NOR2_X1 U11446 ( .A1(n8950), .A2(n15629), .ZN(n8997) );
  NOR2_X1 U11447 ( .A1(n8952), .A2(n8993), .ZN(n8953) );
  INV_X1 U11448 ( .A(n14256), .ZN(n14078) );
  NOR2_X1 U11449 ( .A1(n12866), .A2(n15616), .ZN(n11655) );
  OAI22_X1 U11450 ( .A1(n11655), .A2(n13121), .B1(n13988), .B2(n8886), .ZN(
        n10475) );
  NAND2_X1 U11451 ( .A1(n10475), .A2(n10476), .ZN(n8956) );
  NAND2_X1 U11452 ( .A1(n6962), .A2(n11501), .ZN(n8955) );
  NAND2_X1 U11453 ( .A1(n8956), .A2(n8955), .ZN(n11156) );
  NAND2_X1 U11454 ( .A1(n8957), .A2(n11158), .ZN(n8958) );
  NOR2_X1 U11455 ( .A1(n12907), .A2(n13984), .ZN(n8960) );
  NAND2_X1 U11456 ( .A1(n12907), .A2(n13984), .ZN(n8959) );
  INV_X1 U11457 ( .A(n13128), .ZN(n11103) );
  NAND2_X1 U11458 ( .A1(n11104), .A2(n11103), .ZN(n8962) );
  NAND2_X1 U11459 ( .A1(n15671), .A2(n13983), .ZN(n8961) );
  NAND2_X1 U11460 ( .A1(n8962), .A2(n8961), .ZN(n10896) );
  XNOR2_X1 U11461 ( .A(n12924), .B(n13982), .ZN(n13129) );
  INV_X1 U11462 ( .A(n13129), .ZN(n10899) );
  NAND2_X1 U11463 ( .A1(n10896), .A2(n10899), .ZN(n8964) );
  NAND2_X1 U11464 ( .A1(n12924), .A2(n13982), .ZN(n8963) );
  NAND2_X1 U11465 ( .A1(n8964), .A2(n8963), .ZN(n11090) );
  INV_X1 U11466 ( .A(n13130), .ZN(n11093) );
  NAND2_X1 U11467 ( .A1(n11090), .A2(n11093), .ZN(n8966) );
  NAND2_X1 U11468 ( .A1(n12935), .A2(n13981), .ZN(n8965) );
  NAND2_X1 U11469 ( .A1(n8966), .A2(n8965), .ZN(n11143) );
  NAND2_X1 U11470 ( .A1(n11143), .A2(n13133), .ZN(n8968) );
  NAND2_X1 U11471 ( .A1(n12940), .A2(n13980), .ZN(n8967) );
  NAND2_X1 U11472 ( .A1(n8968), .A2(n8967), .ZN(n11367) );
  NAND2_X1 U11473 ( .A1(n11367), .A2(n13134), .ZN(n8970) );
  NAND2_X1 U11474 ( .A1(n12947), .A2(n13979), .ZN(n8969) );
  AND2_X1 U11475 ( .A1(n15349), .A2(n13978), .ZN(n8971) );
  OR2_X1 U11476 ( .A1(n15349), .A2(n13978), .ZN(n8972) );
  NAND2_X1 U11477 ( .A1(n11712), .A2(n12961), .ZN(n8973) );
  NAND2_X1 U11478 ( .A1(n8973), .A2(n12959), .ZN(n8976) );
  NAND2_X1 U11479 ( .A1(n12988), .A2(n13975), .ZN(n8979) );
  OR2_X1 U11480 ( .A1(n12980), .A2(n13974), .ZN(n8980) );
  NAND2_X1 U11481 ( .A1(n14376), .A2(n13973), .ZN(n8981) );
  NAND2_X1 U11482 ( .A1(n12203), .A2(n8981), .ZN(n14224) );
  XNOR2_X1 U11483 ( .A(n14307), .B(n8982), .ZN(n14223) );
  NAND2_X1 U11484 ( .A1(n14307), .A2(n13972), .ZN(n8983) );
  XNOR2_X1 U11485 ( .A(n14210), .B(n13971), .ZN(n14198) );
  OR2_X1 U11486 ( .A1(n14210), .A2(n13971), .ZN(n8984) );
  INV_X1 U11487 ( .A(n14295), .ZN(n13868) );
  XNOR2_X1 U11488 ( .A(n14285), .B(n13916), .ZN(n14161) );
  OR2_X1 U11489 ( .A1(n14285), .A2(n13968), .ZN(n8985) );
  NAND2_X1 U11490 ( .A1(n14116), .A2(n8987), .ZN(n14125) );
  OR2_X1 U11491 ( .A1(n14274), .A2(n13966), .ZN(n8988) );
  XNOR2_X1 U11492 ( .A(n8991), .B(n13152), .ZN(n14040) );
  OR2_X1 U11493 ( .A1(n15620), .A2(n13169), .ZN(n15675) );
  NAND2_X1 U11494 ( .A1(n15688), .A2(n15366), .ZN(n14316) );
  NOR2_X1 U11495 ( .A1(n8994), .A2(n8993), .ZN(n8996) );
  NAND2_X1 U11496 ( .A1(n15680), .A2(n15366), .ZN(n14379) );
  NAND2_X1 U11497 ( .A1(n9001), .A2(n9000), .ZN(P2_U3496) );
  NOR2_X1 U11498 ( .A1(P3_IR_REG_18__SCAN_IN), .A2(P3_IR_REG_14__SCAN_IN), 
        .ZN(n9007) );
  NAND4_X1 U11499 ( .A1(n9499), .A2(n9010), .A3(n9009), .A4(n9008), .ZN(n9011)
         );
  NOR2_X2 U11500 ( .A1(n9015), .A2(P3_IR_REG_29__SCAN_IN), .ZN(n13830) );
  XNOR2_X2 U11501 ( .A(n9014), .B(P3_IR_REG_30__SCAN_IN), .ZN(n9018) );
  NAND2_X1 U11503 ( .A1(n9300), .A2(P3_REG3_REG_1__SCAN_IN), .ZN(n9024) );
  NAND2_X2 U11504 ( .A1(n13837), .A2(n9020), .ZN(n9346) );
  INV_X1 U11505 ( .A(P3_REG1_REG_1__SCAN_IN), .ZN(n9019) );
  OR2_X1 U11506 ( .A1(n9346), .A2(n9019), .ZN(n9023) );
  NAND2_X1 U11507 ( .A1(n9138), .A2(P3_REG0_REG_1__SCAN_IN), .ZN(n9022) );
  NAND2_X1 U11508 ( .A1(n9089), .A2(P3_REG2_REG_1__SCAN_IN), .ZN(n9021) );
  AND2_X1 U11509 ( .A1(n9039), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n9027) );
  OAI21_X1 U11510 ( .B1(n9028), .B2(n9027), .A(n9047), .ZN(n9954) );
  INV_X1 U11511 ( .A(n9954), .ZN(n9029) );
  NAND2_X1 U11512 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(P3_IR_REG_0__SCAN_IN), 
        .ZN(n9030) );
  INV_X1 U11513 ( .A(n9031), .ZN(n9032) );
  OR2_X1 U11514 ( .A1(n9733), .A2(n10826), .ZN(n9034) );
  NAND2_X1 U11515 ( .A1(n9300), .A2(P3_REG3_REG_0__SCAN_IN), .ZN(n9038) );
  INV_X1 U11516 ( .A(P3_REG1_REG_0__SCAN_IN), .ZN(n15689) );
  INV_X1 U11517 ( .A(SI_0_), .ZN(n9953) );
  OR2_X1 U11518 ( .A1(n9733), .A2(n10763), .ZN(n9040) );
  NAND2_X1 U11519 ( .A1(n6957), .A2(n9041), .ZN(n9544) );
  NAND2_X1 U11520 ( .A1(n10596), .A2(n9544), .ZN(n11050) );
  INV_X1 U11521 ( .A(P3_REG1_REG_2__SCAN_IN), .ZN(n10766) );
  OR2_X1 U11522 ( .A1(n9346), .A2(n10766), .ZN(n9045) );
  NAND2_X1 U11523 ( .A1(n9300), .A2(P3_REG3_REG_2__SCAN_IN), .ZN(n9044) );
  NAND2_X1 U11524 ( .A1(n9138), .A2(P3_REG0_REG_2__SCAN_IN), .ZN(n9043) );
  NAND2_X1 U11525 ( .A1(n6679), .A2(P3_REG2_REG_2__SCAN_IN), .ZN(n9042) );
  NAND4_X2 U11526 ( .A1(n9045), .A2(n9044), .A3(n9043), .A4(n9042), .ZN(n15718) );
  NAND2_X1 U11527 ( .A1(n9982), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n9046) );
  INV_X1 U11528 ( .A(n9057), .ZN(n9048) );
  XNOR2_X1 U11529 ( .A(n9058), .B(n9048), .ZN(n9957) );
  OR2_X1 U11530 ( .A1(n9733), .A2(n11194), .ZN(n9052) );
  INV_X1 U11531 ( .A(n10674), .ZN(n11051) );
  NAND2_X1 U11532 ( .A1(n10836), .A2(n11051), .ZN(n9548) );
  NAND2_X1 U11533 ( .A1(n11049), .A2(n9548), .ZN(n10998) );
  INV_X1 U11534 ( .A(P3_REG3_REG_3__SCAN_IN), .ZN(n10835) );
  NAND2_X1 U11535 ( .A1(n9300), .A2(n10835), .ZN(n9056) );
  NAND2_X1 U11536 ( .A1(n9138), .A2(P3_REG0_REG_3__SCAN_IN), .ZN(n9055) );
  NAND2_X1 U11537 ( .A1(n9089), .A2(P3_REG2_REG_3__SCAN_IN), .ZN(n9054) );
  INV_X1 U11538 ( .A(P3_REG1_REG_3__SCAN_IN), .ZN(n10735) );
  OR2_X1 U11539 ( .A1(n9346), .A2(n10735), .ZN(n9053) );
  NAND2_X1 U11540 ( .A1(n9977), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n9059) );
  INV_X1 U11541 ( .A(n9075), .ZN(n9060) );
  XNOR2_X1 U11542 ( .A(n9076), .B(n9060), .ZN(n9961) );
  NAND2_X1 U11543 ( .A1(n6668), .A2(n9961), .ZN(n9067) );
  OR2_X1 U11544 ( .A1(n9435), .A2(SI_3_), .ZN(n9066) );
  NAND2_X1 U11545 ( .A1(n9061), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9062) );
  MUX2_X1 U11546 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9062), .S(
        P3_IR_REG_3__SCAN_IN), .Z(n9064) );
  NAND2_X1 U11547 ( .A1(n11224), .A2(n10830), .ZN(n9556) );
  INV_X1 U11548 ( .A(n11224), .ZN(n10625) );
  AND2_X2 U11549 ( .A1(n9556), .A2(n9554), .ZN(n11000) );
  NAND2_X1 U11550 ( .A1(n10998), .A2(n11000), .ZN(n9068) );
  NAND2_X1 U11551 ( .A1(n9068), .A2(n9556), .ZN(n11219) );
  NAND2_X1 U11552 ( .A1(n9089), .A2(P3_REG2_REG_4__SCAN_IN), .ZN(n9073) );
  AND2_X1 U11553 ( .A1(P3_REG3_REG_4__SCAN_IN), .A2(P3_REG3_REG_3__SCAN_IN), 
        .ZN(n9069) );
  NOR2_X1 U11554 ( .A1(P3_REG3_REG_3__SCAN_IN), .A2(P3_REG3_REG_4__SCAN_IN), 
        .ZN(n9090) );
  OR2_X1 U11555 ( .A1(n9069), .A2(n9090), .ZN(n11229) );
  NAND2_X1 U11556 ( .A1(n9300), .A2(n11229), .ZN(n9072) );
  NAND2_X1 U11557 ( .A1(n9138), .A2(P3_REG0_REG_4__SCAN_IN), .ZN(n9071) );
  NAND4_X1 U11558 ( .A1(n9074), .A2(n9073), .A3(n9072), .A4(n9071), .ZN(n11425) );
  NAND2_X1 U11559 ( .A1(n9076), .A2(n9075), .ZN(n9078) );
  NAND2_X1 U11560 ( .A1(n10531), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n9077) );
  NAND2_X1 U11561 ( .A1(n9078), .A2(n9077), .ZN(n9098) );
  INV_X1 U11562 ( .A(n9097), .ZN(n9079) );
  XNOR2_X1 U11563 ( .A(n9098), .B(n9079), .ZN(n9971) );
  NAND2_X1 U11564 ( .A1(n9184), .A2(n9971), .ZN(n9086) );
  INV_X1 U11565 ( .A(n9080), .ZN(n9084) );
  NAND2_X1 U11566 ( .A1(n9081), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9082) );
  MUX2_X1 U11567 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9082), .S(
        P3_IR_REG_4__SCAN_IN), .Z(n9083) );
  INV_X1 U11568 ( .A(n10801), .ZN(n10741) );
  OR2_X1 U11569 ( .A1(n10748), .A2(n10741), .ZN(n9085) );
  OAI211_X1 U11570 ( .C1(n6678), .C2(SI_4_), .A(n9086), .B(n9085), .ZN(n11280)
         );
  INV_X1 U11571 ( .A(n11280), .ZN(n9087) );
  NAND2_X1 U11572 ( .A1(n11301), .A2(n9087), .ZN(n9088) );
  NAND2_X1 U11573 ( .A1(n9475), .A2(P3_REG2_REG_5__SCAN_IN), .ZN(n9096) );
  NAND2_X1 U11574 ( .A1(n9090), .A2(n10889), .ZN(n9107) );
  OR2_X1 U11575 ( .A1(n9090), .A2(n10889), .ZN(n9091) );
  NAND2_X1 U11576 ( .A1(n9107), .A2(n9091), .ZN(n11431) );
  NAND2_X1 U11577 ( .A1(n9300), .A2(n11431), .ZN(n9095) );
  NAND2_X1 U11578 ( .A1(n9138), .A2(P3_REG0_REG_5__SCAN_IN), .ZN(n9094) );
  INV_X1 U11579 ( .A(P3_REG1_REG_5__SCAN_IN), .ZN(n9092) );
  OR2_X1 U11580 ( .A1(n9346), .A2(n9092), .ZN(n9093) );
  NAND2_X1 U11582 ( .A1(n9098), .A2(n9097), .ZN(n9100) );
  NAND2_X1 U11583 ( .A1(n9985), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n9099) );
  XNOR2_X1 U11584 ( .A(n9115), .B(n7096), .ZN(n9959) );
  NAND2_X1 U11585 ( .A1(n9184), .A2(n9959), .ZN(n9106) );
  OR2_X1 U11586 ( .A1(n6678), .A2(SI_5_), .ZN(n9105) );
  NOR2_X1 U11587 ( .A1(n9080), .A2(n9682), .ZN(n9101) );
  MUX2_X1 U11588 ( .A(n9682), .B(n9101), .S(P3_IR_REG_5__SCAN_IN), .Z(n9103)
         );
  OR2_X1 U11589 ( .A1(n9103), .A2(n9102), .ZN(n10886) );
  INV_X1 U11590 ( .A(n10886), .ZN(n10802) );
  OR2_X1 U11591 ( .A1(n10748), .A2(n10802), .ZN(n9104) );
  AND3_X2 U11592 ( .A1(n9106), .A2(n9105), .A3(n9104), .ZN(n11432) );
  NAND2_X1 U11593 ( .A1(n11792), .A2(n11432), .ZN(n9562) );
  INV_X1 U11594 ( .A(n11792), .ZN(n11014) );
  NAND2_X1 U11595 ( .A1(n11014), .A2(n15753), .ZN(n9566) );
  NAND2_X1 U11596 ( .A1(n9475), .A2(P3_REG2_REG_6__SCAN_IN), .ZN(n9113) );
  NAND2_X1 U11597 ( .A1(n9107), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n9108) );
  NAND2_X1 U11598 ( .A1(n9121), .A2(n9108), .ZN(n15710) );
  NAND2_X1 U11599 ( .A1(n9300), .A2(n15710), .ZN(n9112) );
  NAND2_X1 U11600 ( .A1(n9138), .A2(P3_REG0_REG_6__SCAN_IN), .ZN(n9111) );
  INV_X1 U11601 ( .A(P3_REG1_REG_6__SCAN_IN), .ZN(n9109) );
  OR2_X1 U11602 ( .A1(n9479), .A2(n9109), .ZN(n9110) );
  INV_X1 U11603 ( .A(SI_6_), .ZN(n9973) );
  NAND2_X1 U11604 ( .A1(n9996), .A2(P2_DATAO_REG_5__SCAN_IN), .ZN(n9116) );
  XNOR2_X1 U11605 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .ZN(n9117) );
  XNOR2_X1 U11606 ( .A(n9129), .B(n9117), .ZN(n9972) );
  NAND2_X1 U11607 ( .A1(n9184), .A2(n9972), .ZN(n9120) );
  OR2_X1 U11608 ( .A1(n9102), .A2(n9682), .ZN(n9118) );
  XNOR2_X1 U11609 ( .A(n9118), .B(P3_IR_REG_6__SCAN_IN), .ZN(n10809) );
  OR2_X1 U11610 ( .A1(n10748), .A2(n10869), .ZN(n9119) );
  OAI211_X1 U11611 ( .C1(n6678), .C2(n9973), .A(n9120), .B(n9119), .ZN(n15708)
         );
  NAND2_X1 U11612 ( .A1(n11602), .A2(n15708), .ZN(n9570) );
  INV_X1 U11613 ( .A(n15708), .ZN(n11799) );
  NAND2_X1 U11614 ( .A1(n11751), .A2(n11799), .ZN(n9568) );
  NAND2_X1 U11615 ( .A1(n11789), .A2(n11790), .ZN(n11788) );
  NAND2_X1 U11616 ( .A1(n11788), .A2(n9570), .ZN(n11756) );
  NAND2_X1 U11617 ( .A1(n9476), .A2(P3_REG0_REG_7__SCAN_IN), .ZN(n9127) );
  AND2_X1 U11618 ( .A1(n9121), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n9122) );
  OR2_X1 U11619 ( .A1(n9122), .A2(n9136), .ZN(n11757) );
  NAND2_X1 U11620 ( .A1(n9300), .A2(n11757), .ZN(n9126) );
  NAND2_X1 U11621 ( .A1(n9475), .A2(P3_REG2_REG_7__SCAN_IN), .ZN(n9125) );
  INV_X1 U11622 ( .A(P3_REG1_REG_7__SCAN_IN), .ZN(n9123) );
  XNOR2_X1 U11623 ( .A(n9144), .B(n9143), .ZN(n9952) );
  NAND2_X1 U11624 ( .A1(n9184), .A2(n9952), .ZN(n9134) );
  OR2_X1 U11625 ( .A1(n6678), .A2(SI_7_), .ZN(n9133) );
  NAND2_X1 U11626 ( .A1(n9102), .A2(n9130), .ZN(n9148) );
  NAND2_X1 U11627 ( .A1(n9148), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9131) );
  OR2_X1 U11628 ( .A1(n10748), .A2(n10986), .ZN(n9132) );
  NAND2_X1 U11629 ( .A1(n11858), .A2(n11896), .ZN(n9574) );
  INV_X1 U11630 ( .A(n11896), .ZN(n11893) );
  INV_X1 U11631 ( .A(n11749), .ZN(n11755) );
  NAND2_X1 U11632 ( .A1(n11756), .A2(n11755), .ZN(n11754) );
  NAND2_X1 U11633 ( .A1(n9475), .A2(P3_REG2_REG_8__SCAN_IN), .ZN(n9142) );
  INV_X1 U11634 ( .A(P3_REG1_REG_8__SCAN_IN), .ZN(n9135) );
  OR2_X1 U11635 ( .A1(n9479), .A2(n9135), .ZN(n9141) );
  NOR2_X1 U11636 ( .A1(n9136), .A2(n10983), .ZN(n9137) );
  OR2_X1 U11637 ( .A1(n9155), .A2(n9137), .ZN(n12020) );
  NAND2_X1 U11638 ( .A1(n9300), .A2(n12020), .ZN(n9140) );
  NAND2_X1 U11639 ( .A1(n9476), .A2(P3_REG0_REG_8__SCAN_IN), .ZN(n9139) );
  NAND2_X1 U11640 ( .A1(n9144), .A2(n9143), .ZN(n9146) );
  NAND2_X1 U11641 ( .A1(n10013), .A2(P1_DATAO_REG_7__SCAN_IN), .ZN(n9145) );
  INV_X1 U11642 ( .A(n9159), .ZN(n9147) );
  XNOR2_X1 U11643 ( .A(n9160), .B(n9147), .ZN(n9965) );
  NAND2_X1 U11644 ( .A1(n9184), .A2(n9965), .ZN(n9153) );
  NAND2_X1 U11645 ( .A1(n9164), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9150) );
  OR2_X1 U11646 ( .A1(n10748), .A2(n11331), .ZN(n9152) );
  INV_X1 U11647 ( .A(SI_8_), .ZN(n9967) );
  OR2_X1 U11648 ( .A1(n6678), .A2(n9967), .ZN(n9151) );
  INV_X1 U11649 ( .A(n12173), .ZN(n11855) );
  NAND2_X1 U11650 ( .A1(n11640), .A2(n11855), .ZN(n9154) );
  NAND2_X1 U11651 ( .A1(n9475), .A2(P3_REG2_REG_9__SCAN_IN), .ZN(n9158) );
  INV_X1 U11652 ( .A(P3_REG1_REG_9__SCAN_IN), .ZN(n15780) );
  OR2_X1 U11653 ( .A1(n9155), .A2(n11335), .ZN(n9156) );
  NAND2_X1 U11654 ( .A1(n9173), .A2(n9156), .ZN(n12038) );
  NAND2_X1 U11655 ( .A1(n9476), .A2(P3_REG0_REG_9__SCAN_IN), .ZN(n9157) );
  NAND2_X1 U11656 ( .A1(n9160), .A2(n9159), .ZN(n9163) );
  NAND2_X1 U11657 ( .A1(n9161), .A2(P1_DATAO_REG_8__SCAN_IN), .ZN(n9162) );
  NAND2_X1 U11658 ( .A1(n9163), .A2(n9162), .ZN(n9180) );
  XNOR2_X1 U11659 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(P2_DATAO_REG_9__SCAN_IN), 
        .ZN(n9179) );
  XNOR2_X1 U11660 ( .A(n9180), .B(n9179), .ZN(n9968) );
  NAND2_X1 U11661 ( .A1(n9184), .A2(n9968), .ZN(n9170) );
  NOR2_X1 U11662 ( .A1(n9164), .A2(P3_IR_REG_8__SCAN_IN), .ZN(n9167) );
  OR2_X1 U11663 ( .A1(n9167), .A2(n9682), .ZN(n9165) );
  MUX2_X1 U11664 ( .A(n9165), .B(P3_IR_REG_31__SCAN_IN), .S(n9166), .Z(n9168)
         );
  NAND2_X1 U11665 ( .A1(n9167), .A2(n9166), .ZN(n9203) );
  NAND2_X1 U11666 ( .A1(n9168), .A2(n9203), .ZN(n11332) );
  OR2_X1 U11667 ( .A1(n10748), .A2(n11445), .ZN(n9169) );
  OAI211_X1 U11668 ( .C1(n6678), .C2(SI_9_), .A(n9170), .B(n9169), .ZN(n15759)
         );
  INV_X1 U11669 ( .A(n12018), .ZN(n9172) );
  INV_X1 U11670 ( .A(n15759), .ZN(n9582) );
  INV_X1 U11671 ( .A(n11995), .ZN(n9191) );
  NAND2_X1 U11672 ( .A1(n9476), .A2(P3_REG0_REG_10__SCAN_IN), .ZN(n9178) );
  NAND2_X1 U11673 ( .A1(n9173), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n9174) );
  NAND2_X1 U11674 ( .A1(n9192), .A2(n9174), .ZN(n12009) );
  NAND2_X1 U11675 ( .A1(n9300), .A2(n12009), .ZN(n9177) );
  NAND2_X1 U11676 ( .A1(n9475), .A2(P3_REG2_REG_10__SCAN_IN), .ZN(n9176) );
  INV_X1 U11677 ( .A(P3_REG1_REG_10__SCAN_IN), .ZN(n11451) );
  OR2_X1 U11678 ( .A1(n9479), .A2(n11451), .ZN(n9175) );
  NAND2_X1 U11679 ( .A1(n9180), .A2(n9179), .ZN(n9183) );
  NAND2_X1 U11680 ( .A1(n9181), .A2(P1_DATAO_REG_9__SCAN_IN), .ZN(n9182) );
  NAND2_X1 U11681 ( .A1(n9183), .A2(n9182), .ZN(n9200) );
  XNOR2_X1 U11682 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(P2_DATAO_REG_10__SCAN_IN), 
        .ZN(n9199) );
  XNOR2_X1 U11683 ( .A(n9200), .B(n9199), .ZN(n9978) );
  NAND2_X1 U11684 ( .A1(n9184), .A2(n9978), .ZN(n9189) );
  OR2_X1 U11685 ( .A1(n6678), .A2(SI_10_), .ZN(n9188) );
  NAND2_X1 U11686 ( .A1(n9203), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9186) );
  INV_X1 U11687 ( .A(P3_IR_REG_10__SCAN_IN), .ZN(n9185) );
  INV_X1 U11688 ( .A(n11914), .ZN(n11463) );
  OR2_X1 U11689 ( .A1(n10748), .A2(n11463), .ZN(n9187) );
  NAND2_X1 U11690 ( .A1(n12050), .A2(n15766), .ZN(n9586) );
  INV_X1 U11691 ( .A(n15766), .ZN(n12011) );
  NAND2_X1 U11692 ( .A1(n12145), .A2(n12011), .ZN(n9593) );
  NAND2_X1 U11693 ( .A1(n9586), .A2(n9593), .ZN(n12005) );
  INV_X1 U11694 ( .A(n12005), .ZN(n9190) );
  NAND2_X1 U11695 ( .A1(n9475), .A2(P3_REG2_REG_11__SCAN_IN), .ZN(n9198) );
  NAND2_X1 U11696 ( .A1(n9192), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n9193) );
  NAND2_X1 U11697 ( .A1(n9209), .A2(n9193), .ZN(n12144) );
  NAND2_X1 U11698 ( .A1(n9300), .A2(n12144), .ZN(n9197) );
  NAND2_X1 U11699 ( .A1(n9476), .A2(P3_REG0_REG_11__SCAN_IN), .ZN(n9196) );
  INV_X1 U11700 ( .A(P3_REG1_REG_11__SCAN_IN), .ZN(n9194) );
  OR2_X1 U11701 ( .A1(n9479), .A2(n9194), .ZN(n9195) );
  NAND2_X1 U11702 ( .A1(n9200), .A2(n9199), .ZN(n9202) );
  NAND2_X1 U11703 ( .A1(n10073), .A2(P1_DATAO_REG_10__SCAN_IN), .ZN(n9201) );
  XNOR2_X1 U11704 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(P2_DATAO_REG_11__SCAN_IN), 
        .ZN(n9216) );
  XNOR2_X1 U11705 ( .A(n9217), .B(n9216), .ZN(n9983) );
  NAND2_X1 U11706 ( .A1(n9184), .A2(n9983), .ZN(n9207) );
  OAI21_X1 U11707 ( .B1(n9203), .B2(P3_IR_REG_10__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n9205) );
  INV_X1 U11708 ( .A(P3_IR_REG_11__SCAN_IN), .ZN(n9204) );
  XNOR2_X1 U11709 ( .A(n9205), .B(n9204), .ZN(n11981) );
  INV_X1 U11710 ( .A(n11981), .ZN(n11977) );
  OR2_X1 U11711 ( .A1(n10748), .A2(n11977), .ZN(n9206) );
  OAI211_X1 U11712 ( .C1(n6678), .C2(SI_11_), .A(n9207), .B(n9206), .ZN(n15326) );
  NAND2_X1 U11713 ( .A1(n12377), .A2(n15326), .ZN(n12090) );
  INV_X1 U11714 ( .A(n15326), .ZN(n12143) );
  NAND2_X1 U11715 ( .A1(n12223), .A2(n12143), .ZN(n9208) );
  NAND2_X1 U11716 ( .A1(n12090), .A2(n9208), .ZN(n12048) );
  NAND2_X1 U11717 ( .A1(n12377), .A2(n12143), .ZN(n9588) );
  NAND2_X1 U11718 ( .A1(n9475), .A2(P3_REG2_REG_12__SCAN_IN), .ZN(n9215) );
  AND2_X1 U11719 ( .A1(n9209), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n9210) );
  OR2_X1 U11720 ( .A1(n9210), .A2(n9236), .ZN(n12374) );
  NAND2_X1 U11721 ( .A1(n9300), .A2(n12374), .ZN(n9214) );
  NAND2_X1 U11722 ( .A1(n9476), .A2(P3_REG0_REG_12__SCAN_IN), .ZN(n9213) );
  INV_X1 U11723 ( .A(P3_REG1_REG_12__SCAN_IN), .ZN(n9211) );
  OR2_X1 U11724 ( .A1(n9479), .A2(n9211), .ZN(n9212) );
  NAND2_X1 U11725 ( .A1(n9217), .A2(n9216), .ZN(n9219) );
  NAND2_X1 U11726 ( .A1(n10246), .A2(P1_DATAO_REG_11__SCAN_IN), .ZN(n9218) );
  NAND2_X1 U11727 ( .A1(n9219), .A2(n9218), .ZN(n9228) );
  XNOR2_X1 U11728 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(P2_DATAO_REG_12__SCAN_IN), 
        .ZN(n9229) );
  INV_X1 U11729 ( .A(n9229), .ZN(n9220) );
  XNOR2_X1 U11730 ( .A(n9228), .B(n9220), .ZN(n9997) );
  NAND2_X1 U11731 ( .A1(n9184), .A2(n9997), .ZN(n9226) );
  NAND2_X1 U11732 ( .A1(n9221), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9222) );
  MUX2_X1 U11733 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9222), .S(
        P3_IR_REG_12__SCAN_IN), .Z(n9224) );
  NAND2_X1 U11734 ( .A1(n9224), .A2(n9223), .ZN(n13377) );
  OR2_X1 U11735 ( .A1(n10748), .A2(n13377), .ZN(n9225) );
  OAI211_X1 U11736 ( .C1(n6678), .C2(n9999), .A(n9226), .B(n9225), .ZN(n15325)
         );
  NAND2_X1 U11737 ( .A1(n12230), .A2(n15325), .ZN(n9598) );
  INV_X1 U11738 ( .A(n15325), .ZN(n12096) );
  NAND2_X1 U11739 ( .A1(n13356), .A2(n12096), .ZN(n9596) );
  NAND2_X1 U11740 ( .A1(n9598), .A2(n9596), .ZN(n12089) );
  INV_X1 U11741 ( .A(n12089), .ZN(n9516) );
  NAND2_X1 U11742 ( .A1(n12087), .A2(n9516), .ZN(n9227) );
  NAND2_X1 U11743 ( .A1(n9229), .A2(n9228), .ZN(n9230) );
  XNOR2_X1 U11744 ( .A(n9242), .B(P1_DATAO_REG_13__SCAN_IN), .ZN(n10017) );
  NAND2_X1 U11745 ( .A1(n9223), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9231) );
  MUX2_X1 U11746 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9231), .S(
        P3_IR_REG_13__SCAN_IN), .Z(n9232) );
  NAND2_X1 U11747 ( .A1(n9232), .A2(n9259), .ZN(n13394) );
  INV_X1 U11748 ( .A(n13394), .ZN(n13388) );
  OAI22_X1 U11749 ( .A1(n6678), .A2(SI_13_), .B1(n13388), .B2(n10748), .ZN(
        n9233) );
  NAND2_X1 U11750 ( .A1(n9475), .A2(P3_REG2_REG_13__SCAN_IN), .ZN(n9241) );
  INV_X1 U11751 ( .A(P3_REG1_REG_13__SCAN_IN), .ZN(n9234) );
  OR2_X1 U11752 ( .A1(n9479), .A2(n9234), .ZN(n9240) );
  OR2_X1 U11753 ( .A1(n9236), .A2(n9235), .ZN(n9237) );
  NAND2_X1 U11754 ( .A1(n9249), .A2(n9237), .ZN(n12227) );
  NAND2_X1 U11755 ( .A1(n9300), .A2(n12227), .ZN(n9239) );
  NAND2_X1 U11756 ( .A1(n9476), .A2(P3_REG0_REG_13__SCAN_IN), .ZN(n9238) );
  NAND4_X1 U11757 ( .A1(n9241), .A2(n9240), .A3(n9239), .A4(n9238), .ZN(n13355) );
  AND2_X1 U11758 ( .A1(n15318), .A2(n13180), .ZN(n9601) );
  INV_X1 U11759 ( .A(n15318), .ZN(n12199) );
  NAND2_X1 U11760 ( .A1(n12199), .A2(n13355), .ZN(n9603) );
  NAND2_X1 U11761 ( .A1(n10458), .A2(n9243), .ZN(n9244) );
  XNOR2_X1 U11762 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(P2_DATAO_REG_14__SCAN_IN), 
        .ZN(n9255) );
  XNOR2_X1 U11763 ( .A(n9256), .B(n9255), .ZN(n10028) );
  NAND2_X1 U11764 ( .A1(n10028), .A2(n9184), .ZN(n9248) );
  NAND2_X1 U11765 ( .A1(n9259), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9245) );
  XNOR2_X1 U11766 ( .A(n9245), .B(n7307), .ZN(n13405) );
  INV_X1 U11767 ( .A(n13405), .ZN(n13390) );
  OAI22_X1 U11768 ( .A1(n6678), .A2(SI_14_), .B1(n13390), .B2(n10748), .ZN(
        n9246) );
  INV_X1 U11769 ( .A(n9246), .ZN(n9247) );
  NAND2_X1 U11770 ( .A1(n9475), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n9254) );
  INV_X1 U11771 ( .A(P3_REG1_REG_14__SCAN_IN), .ZN(n13775) );
  OR2_X1 U11772 ( .A1(n9479), .A2(n13775), .ZN(n9253) );
  NAND2_X1 U11773 ( .A1(n9249), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n9250) );
  NAND2_X1 U11774 ( .A1(n9264), .A2(n9250), .ZN(n13228) );
  NAND2_X1 U11775 ( .A1(n9300), .A2(n13228), .ZN(n9252) );
  NAND2_X1 U11776 ( .A1(n9476), .A2(P3_REG0_REG_14__SCAN_IN), .ZN(n9251) );
  NAND4_X1 U11777 ( .A1(n9254), .A2(n9253), .A3(n9252), .A4(n9251), .ZN(n13706) );
  NAND2_X1 U11778 ( .A1(n13824), .A2(n13706), .ZN(n9606) );
  OR2_X1 U11779 ( .A1(n13824), .A2(n13706), .ZN(n9607) );
  NAND2_X1 U11780 ( .A1(n10650), .A2(P1_DATAO_REG_14__SCAN_IN), .ZN(n9257) );
  XNOR2_X1 U11781 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(P2_DATAO_REG_15__SCAN_IN), 
        .ZN(n9272) );
  INV_X1 U11782 ( .A(n9272), .ZN(n9258) );
  XNOR2_X1 U11783 ( .A(n9273), .B(n9258), .ZN(n10128) );
  NAND2_X1 U11784 ( .A1(n10128), .A2(n9184), .ZN(n9263) );
  XNOR2_X1 U11785 ( .A(n9260), .B(P3_IR_REG_15__SCAN_IN), .ZN(n13449) );
  INV_X1 U11786 ( .A(n13449), .ZN(n13427) );
  OAI22_X1 U11787 ( .A1(n6678), .A2(n10130), .B1(n10748), .B2(n13427), .ZN(
        n9261) );
  INV_X1 U11788 ( .A(n9261), .ZN(n9262) );
  NAND2_X1 U11789 ( .A1(n9263), .A2(n9262), .ZN(n13187) );
  NAND2_X1 U11790 ( .A1(n9476), .A2(P3_REG0_REG_15__SCAN_IN), .ZN(n9270) );
  INV_X1 U11791 ( .A(n9280), .ZN(n9266) );
  NAND2_X1 U11792 ( .A1(n9264), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n9265) );
  NAND2_X1 U11793 ( .A1(n9266), .A2(n9265), .ZN(n13712) );
  NAND2_X1 U11794 ( .A1(n9300), .A2(n13712), .ZN(n9269) );
  NAND2_X1 U11795 ( .A1(n9475), .A2(P3_REG2_REG_15__SCAN_IN), .ZN(n9268) );
  INV_X1 U11796 ( .A(P3_REG1_REG_15__SCAN_IN), .ZN(n13429) );
  OR2_X1 U11797 ( .A1(n9479), .A2(n13429), .ZN(n9267) );
  OR2_X1 U11798 ( .A1(n13187), .A2(n13693), .ZN(n9610) );
  NAND2_X1 U11799 ( .A1(n13187), .A2(n13693), .ZN(n9615) );
  NAND2_X1 U11800 ( .A1(n13709), .A2(n13710), .ZN(n9271) );
  NAND2_X1 U11801 ( .A1(n9271), .A2(n9615), .ZN(n13697) );
  XNOR2_X1 U11802 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(P2_DATAO_REG_16__SCAN_IN), 
        .ZN(n9287) );
  INV_X1 U11803 ( .A(n9287), .ZN(n9274) );
  XNOR2_X1 U11804 ( .A(n9288), .B(n9274), .ZN(n10248) );
  NAND2_X1 U11805 ( .A1(n10248), .A2(n9184), .ZN(n9279) );
  OR2_X1 U11806 ( .A1(n9290), .A2(n9682), .ZN(n9276) );
  XNOR2_X1 U11807 ( .A(n9276), .B(n9289), .ZN(n13452) );
  OAI22_X1 U11808 ( .A1(n6678), .A2(n10250), .B1(n10748), .B2(n13452), .ZN(
        n9277) );
  INV_X1 U11809 ( .A(n9277), .ZN(n9278) );
  NAND2_X1 U11810 ( .A1(n9279), .A2(n9278), .ZN(n13699) );
  NAND2_X1 U11811 ( .A1(n9475), .A2(P3_REG2_REG_16__SCAN_IN), .ZN(n9285) );
  NOR2_X1 U11812 ( .A1(n9280), .A2(n13280), .ZN(n9281) );
  OR2_X1 U11813 ( .A1(n9298), .A2(n9281), .ZN(n13700) );
  NAND2_X1 U11814 ( .A1(n9300), .A2(n13700), .ZN(n9284) );
  NAND2_X1 U11815 ( .A1(n9476), .A2(P3_REG0_REG_16__SCAN_IN), .ZN(n9283) );
  INV_X1 U11816 ( .A(P3_REG1_REG_16__SCAN_IN), .ZN(n13767) );
  OR2_X1 U11817 ( .A1(n9479), .A2(n13767), .ZN(n9282) );
  OR2_X1 U11818 ( .A1(n13699), .A2(n13680), .ZN(n9617) );
  NAND2_X1 U11819 ( .A1(n13699), .A2(n13680), .ZN(n9616) );
  NAND2_X1 U11820 ( .A1(n9617), .A2(n9616), .ZN(n13689) );
  NAND2_X1 U11821 ( .A1(n13697), .A2(n7639), .ZN(n9286) );
  NAND2_X1 U11822 ( .A1(n9286), .A2(n9616), .ZN(n13675) );
  AOI22_X1 U11823 ( .A1(P2_DATAO_REG_17__SCAN_IN), .A2(n10652), .B1(
        P1_DATAO_REG_17__SCAN_IN), .B2(n10671), .ZN(n9306) );
  XOR2_X1 U11824 ( .A(n9307), .B(n9306), .Z(n10434) );
  INV_X1 U11825 ( .A(SI_17_), .ZN(n10436) );
  NOR2_X1 U11826 ( .A1(n9294), .A2(n9682), .ZN(n9291) );
  MUX2_X1 U11827 ( .A(n9682), .B(n9291), .S(P3_IR_REG_17__SCAN_IN), .Z(n9292)
         );
  INV_X1 U11828 ( .A(n9292), .ZN(n9295) );
  AND2_X1 U11829 ( .A1(n9295), .A2(n9326), .ZN(n13501) );
  OAI22_X1 U11830 ( .A1(n6678), .A2(n10436), .B1(n10748), .B2(n13494), .ZN(
        n9296) );
  NAND2_X1 U11831 ( .A1(n9475), .A2(P3_REG2_REG_17__SCAN_IN), .ZN(n9304) );
  INV_X1 U11832 ( .A(P3_REG1_REG_17__SCAN_IN), .ZN(n13468) );
  OR2_X1 U11833 ( .A1(n9479), .A2(n13468), .ZN(n9303) );
  OR2_X1 U11834 ( .A1(n9298), .A2(n9297), .ZN(n9299) );
  NAND2_X1 U11835 ( .A1(n9316), .A2(n9299), .ZN(n13682) );
  NAND2_X1 U11836 ( .A1(n9300), .A2(n13682), .ZN(n9302) );
  NAND2_X1 U11837 ( .A1(n9476), .A2(P3_REG0_REG_17__SCAN_IN), .ZN(n9301) );
  NAND4_X1 U11838 ( .A1(n9304), .A2(n9303), .A3(n9302), .A4(n9301), .ZN(n13326) );
  NAND2_X1 U11839 ( .A1(n13295), .A2(n13326), .ZN(n9621) );
  INV_X1 U11840 ( .A(n13295), .ZN(n13762) );
  NAND2_X1 U11841 ( .A1(n13762), .A2(n13695), .ZN(n9620) );
  NAND2_X1 U11842 ( .A1(n13675), .A2(n13677), .ZN(n9305) );
  NAND2_X1 U11843 ( .A1(n9305), .A2(n9620), .ZN(n13671) );
  AOI22_X1 U11844 ( .A1(P2_DATAO_REG_18__SCAN_IN), .A2(n11256), .B1(
        P1_DATAO_REG_18__SCAN_IN), .B2(n11262), .ZN(n9323) );
  INV_X1 U11845 ( .A(n9323), .ZN(n9310) );
  XNOR2_X1 U11846 ( .A(n9322), .B(n9310), .ZN(n10520) );
  NAND2_X1 U11847 ( .A1(n10520), .A2(n9184), .ZN(n9315) );
  NAND2_X1 U11848 ( .A1(n9326), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9312) );
  INV_X1 U11849 ( .A(P3_IR_REG_18__SCAN_IN), .ZN(n9311) );
  XNOR2_X1 U11850 ( .A(n9312), .B(n9311), .ZN(n13513) );
  OAI22_X1 U11851 ( .A1(n6678), .A2(n10522), .B1(n10748), .B2(n13513), .ZN(
        n9313) );
  INV_X1 U11852 ( .A(n9313), .ZN(n9314) );
  NAND2_X1 U11853 ( .A1(n9315), .A2(n9314), .ZN(n13670) );
  NAND2_X1 U11854 ( .A1(n9476), .A2(P3_REG0_REG_18__SCAN_IN), .ZN(n9321) );
  NAND2_X1 U11855 ( .A1(n9316), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n9317) );
  NAND2_X1 U11856 ( .A1(n9331), .A2(n9317), .ZN(n13666) );
  NAND2_X1 U11857 ( .A1(n9300), .A2(n13666), .ZN(n9320) );
  NAND2_X1 U11858 ( .A1(n9475), .A2(P3_REG2_REG_18__SCAN_IN), .ZN(n9319) );
  INV_X1 U11859 ( .A(P3_REG1_REG_18__SCAN_IN), .ZN(n13504) );
  OR2_X1 U11860 ( .A1(n9479), .A2(n13504), .ZN(n9318) );
  NAND2_X1 U11861 ( .A1(n13670), .A2(n13681), .ZN(n9628) );
  AOI22_X1 U11862 ( .A1(P2_DATAO_REG_19__SCAN_IN), .A2(n12566), .B1(
        P1_DATAO_REG_19__SCAN_IN), .B2(n11316), .ZN(n9338) );
  XNOR2_X1 U11863 ( .A(n9339), .B(n9338), .ZN(n10545) );
  NAND2_X1 U11864 ( .A1(n10545), .A2(n6668), .ZN(n9330) );
  OAI22_X1 U11865 ( .A1(n6678), .A2(SI_19_), .B1(n9769), .B2(n10748), .ZN(
        n9328) );
  INV_X1 U11866 ( .A(n9328), .ZN(n9329) );
  NAND2_X1 U11867 ( .A1(n9475), .A2(P3_REG2_REG_19__SCAN_IN), .ZN(n9336) );
  INV_X1 U11868 ( .A(P3_REG1_REG_19__SCAN_IN), .ZN(n13754) );
  OR2_X1 U11869 ( .A1(n9479), .A2(n13754), .ZN(n9335) );
  AND2_X1 U11870 ( .A1(n9331), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n9332) );
  OR2_X1 U11871 ( .A1(n9332), .A2(n9344), .ZN(n13655) );
  NAND2_X1 U11872 ( .A1(n9300), .A2(n13655), .ZN(n9334) );
  NAND2_X1 U11873 ( .A1(n9476), .A2(P3_REG0_REG_19__SCAN_IN), .ZN(n9333) );
  NAND4_X1 U11874 ( .A1(n9336), .A2(n9335), .A3(n9334), .A4(n9333), .ZN(n13308) );
  NAND2_X1 U11875 ( .A1(n13813), .A2(n13308), .ZN(n9633) );
  INV_X1 U11876 ( .A(n9633), .ZN(n9337) );
  OR2_X1 U11877 ( .A1(n13813), .A2(n13308), .ZN(n9634) );
  INV_X1 U11878 ( .A(n13642), .ZN(n9352) );
  XNOR2_X1 U11879 ( .A(n9354), .B(P2_DATAO_REG_20__SCAN_IN), .ZN(n10923) );
  NAND2_X1 U11880 ( .A1(n10923), .A2(n9184), .ZN(n9342) );
  OR2_X1 U11881 ( .A1(n6678), .A2(n10924), .ZN(n9341) );
  NOR2_X1 U11882 ( .A1(n9344), .A2(n9343), .ZN(n9345) );
  OR2_X1 U11883 ( .A1(n9362), .A2(n9345), .ZN(n13643) );
  NAND2_X1 U11884 ( .A1(n13643), .A2(n9300), .ZN(n9350) );
  INV_X1 U11885 ( .A(P3_REG1_REG_20__SCAN_IN), .ZN(n13750) );
  OR2_X1 U11886 ( .A1(n9479), .A2(n13750), .ZN(n9349) );
  NAND2_X1 U11887 ( .A1(n9476), .A2(P3_REG0_REG_20__SCAN_IN), .ZN(n9348) );
  NAND2_X1 U11888 ( .A1(n9475), .A2(P3_REG2_REG_20__SCAN_IN), .ZN(n9347) );
  NAND4_X1 U11889 ( .A1(n9350), .A2(n9349), .A3(n9348), .A4(n9347), .ZN(n13652) );
  NAND2_X1 U11890 ( .A1(n13809), .A2(n13652), .ZN(n9639) );
  INV_X1 U11891 ( .A(n13809), .ZN(n9351) );
  NAND2_X1 U11892 ( .A1(n9351), .A2(n13629), .ZN(n9638) );
  NAND2_X1 U11893 ( .A1(n13639), .A2(n9639), .ZN(n13622) );
  NAND2_X1 U11894 ( .A1(P1_DATAO_REG_20__SCAN_IN), .A2(n9353), .ZN(n9355) );
  INV_X1 U11895 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n12426) );
  AOI22_X1 U11896 ( .A1(P2_DATAO_REG_21__SCAN_IN), .A2(n11960), .B1(
        P1_DATAO_REG_21__SCAN_IN), .B2(n9370), .ZN(n9368) );
  INV_X1 U11897 ( .A(n9368), .ZN(n9356) );
  XNOR2_X1 U11898 ( .A(n9369), .B(n9356), .ZN(n11168) );
  NAND2_X1 U11899 ( .A1(n11168), .A2(n9184), .ZN(n9358) );
  INV_X1 U11900 ( .A(SI_21_), .ZN(n11170) );
  OR2_X1 U11901 ( .A1(n6678), .A2(n11170), .ZN(n9357) );
  NAND2_X1 U11902 ( .A1(n9475), .A2(P3_REG2_REG_21__SCAN_IN), .ZN(n9360) );
  INV_X1 U11903 ( .A(P3_REG1_REG_21__SCAN_IN), .ZN(n13746) );
  OR2_X1 U11904 ( .A1(n9479), .A2(n13746), .ZN(n9359) );
  AND2_X1 U11905 ( .A1(n9360), .A2(n9359), .ZN(n9366) );
  INV_X1 U11906 ( .A(P3_REG3_REG_21__SCAN_IN), .ZN(n9361) );
  OR2_X1 U11907 ( .A1(n9362), .A2(n9361), .ZN(n9363) );
  NAND2_X1 U11908 ( .A1(n9376), .A2(n9363), .ZN(n13631) );
  NAND2_X1 U11909 ( .A1(n13631), .A2(n9300), .ZN(n9365) );
  NAND2_X1 U11910 ( .A1(n9476), .A2(P3_REG0_REG_21__SCAN_IN), .ZN(n9364) );
  NAND2_X1 U11911 ( .A1(n13267), .A2(n13638), .ZN(n9537) );
  NAND2_X1 U11912 ( .A1(n13622), .A2(n9537), .ZN(n9367) );
  NAND2_X1 U11913 ( .A1(n9367), .A2(n9538), .ZN(n13614) );
  INV_X1 U11914 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n9372) );
  AOI22_X1 U11915 ( .A1(P2_DATAO_REG_22__SCAN_IN), .A2(
        P1_DATAO_REG_22__SCAN_IN), .B1(n12860), .B2(n9372), .ZN(n9382) );
  XNOR2_X1 U11916 ( .A(n9383), .B(n9382), .ZN(n11284) );
  NAND2_X1 U11917 ( .A1(n11284), .A2(n6668), .ZN(n9375) );
  NAND2_X1 U11918 ( .A1(n9376), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n9377) );
  NAND2_X1 U11919 ( .A1(n9386), .A2(n9377), .ZN(n13617) );
  NAND2_X1 U11920 ( .A1(n13617), .A2(n9300), .ZN(n9380) );
  AOI22_X1 U11921 ( .A1(n9388), .A2(P3_REG1_REG_22__SCAN_IN), .B1(n9475), .B2(
        P3_REG2_REG_22__SCAN_IN), .ZN(n9379) );
  NAND2_X1 U11922 ( .A1(n9476), .A2(P3_REG0_REG_22__SCAN_IN), .ZN(n9378) );
  NAND2_X1 U11923 ( .A1(n13318), .A2(n13630), .ZN(n9535) );
  NAND2_X1 U11924 ( .A1(n13614), .A2(n9535), .ZN(n9381) );
  NAND2_X1 U11925 ( .A1(n9381), .A2(n9536), .ZN(n13599) );
  INV_X1 U11926 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n12458) );
  AOI22_X1 U11927 ( .A1(P2_DATAO_REG_23__SCAN_IN), .A2(
        P1_DATAO_REG_23__SCAN_IN), .B1(n12060), .B2(n12458), .ZN(n9393) );
  XNOR2_X1 U11928 ( .A(n9394), .B(n9393), .ZN(n11597) );
  NAND2_X1 U11929 ( .A1(n11597), .A2(n6668), .ZN(n9385) );
  OR2_X1 U11930 ( .A1(n6678), .A2(n11600), .ZN(n9384) );
  INV_X1 U11931 ( .A(P3_REG0_REG_23__SCAN_IN), .ZN(n13795) );
  NAND2_X1 U11932 ( .A1(n9386), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n9387) );
  NAND2_X1 U11933 ( .A1(n9396), .A2(n9387), .ZN(n13606) );
  NAND2_X1 U11934 ( .A1(n13606), .A2(n9300), .ZN(n9390) );
  AOI22_X1 U11935 ( .A1(n9388), .A2(P3_REG1_REG_23__SCAN_IN), .B1(n9475), .B2(
        P3_REG2_REG_23__SCAN_IN), .ZN(n9389) );
  OAI211_X1 U11936 ( .C1(n9070), .C2(n13795), .A(n9390), .B(n9389), .ZN(n13298) );
  NAND2_X1 U11937 ( .A1(n13797), .A2(n13298), .ZN(n9531) );
  INV_X1 U11938 ( .A(n13797), .ZN(n13239) );
  NAND2_X1 U11939 ( .A1(n13239), .A2(n13613), .ZN(n9391) );
  NAND2_X1 U11940 ( .A1(n9531), .A2(n9391), .ZN(n13602) );
  INV_X1 U11941 ( .A(n13602), .ZN(n9721) );
  INV_X1 U11942 ( .A(n9531), .ZN(n9392) );
  AOI21_X2 U11943 ( .B1(n13599), .B2(n9721), .A(n9392), .ZN(n13593) );
  XOR2_X1 U11944 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(n9405), .Z(n12126) );
  NOR2_X1 U11945 ( .A1(n6678), .A2(n8147), .ZN(n9395) );
  INV_X1 U11946 ( .A(n9410), .ZN(n9398) );
  NAND2_X1 U11947 ( .A1(n9396), .A2(P3_REG3_REG_24__SCAN_IN), .ZN(n9397) );
  NAND2_X1 U11948 ( .A1(n9398), .A2(n9397), .ZN(n13594) );
  NAND2_X1 U11949 ( .A1(n13594), .A2(n9300), .ZN(n9403) );
  INV_X1 U11950 ( .A(P3_REG1_REG_24__SCAN_IN), .ZN(n13734) );
  NAND2_X1 U11951 ( .A1(n9475), .A2(P3_REG2_REG_24__SCAN_IN), .ZN(n9400) );
  NAND2_X1 U11952 ( .A1(n9476), .A2(P3_REG0_REG_24__SCAN_IN), .ZN(n9399) );
  OAI211_X1 U11953 ( .C1(n9479), .C2(n13734), .A(n9400), .B(n9399), .ZN(n9401)
         );
  INV_X1 U11954 ( .A(n9401), .ZN(n9402) );
  NAND2_X1 U11955 ( .A1(n13793), .A2(n13603), .ZN(n9532) );
  INV_X1 U11956 ( .A(n13793), .ZN(n13302) );
  NAND2_X1 U11957 ( .A1(n13302), .A2(n13580), .ZN(n9533) );
  NAND2_X1 U11958 ( .A1(n13593), .A2(n13592), .ZN(n13591) );
  NAND2_X1 U11959 ( .A1(P1_DATAO_REG_24__SCAN_IN), .A2(n9404), .ZN(n9406) );
  AOI22_X1 U11960 ( .A1(P2_DATAO_REG_25__SCAN_IN), .A2(
        P1_DATAO_REG_25__SCAN_IN), .B1(n12390), .B2(n12481), .ZN(n9419) );
  XNOR2_X1 U11961 ( .A(n9418), .B(n9419), .ZN(n12177) );
  NAND2_X1 U11962 ( .A1(n12177), .A2(n9184), .ZN(n9408) );
  NAND2_X1 U11963 ( .A1(n9410), .A2(n9409), .ZN(n9425) );
  OR2_X1 U11964 ( .A1(n9410), .A2(n9409), .ZN(n9411) );
  NAND2_X1 U11965 ( .A1(n9425), .A2(n9411), .ZN(n13582) );
  NAND2_X1 U11966 ( .A1(n13582), .A2(n9300), .ZN(n9416) );
  INV_X1 U11967 ( .A(P3_REG1_REG_25__SCAN_IN), .ZN(n13730) );
  NAND2_X1 U11968 ( .A1(n9475), .A2(P3_REG2_REG_25__SCAN_IN), .ZN(n9413) );
  NAND2_X1 U11969 ( .A1(n9476), .A2(P3_REG0_REG_25__SCAN_IN), .ZN(n9412) );
  OAI211_X1 U11970 ( .C1(n9479), .C2(n13730), .A(n9413), .B(n9412), .ZN(n9414)
         );
  INV_X1 U11971 ( .A(n9414), .ZN(n9415) );
  OR2_X1 U11972 ( .A1(n13581), .A2(n13590), .ZN(n9652) );
  NAND2_X1 U11973 ( .A1(n13581), .A2(n13590), .ZN(n9651) );
  NAND2_X1 U11974 ( .A1(n13573), .A2(n13574), .ZN(n9417) );
  NAND2_X2 U11975 ( .A1(n9417), .A2(n9651), .ZN(n13566) );
  NOR2_X1 U11976 ( .A1(n9419), .A2(n9418), .ZN(n9420) );
  AOI22_X1 U11977 ( .A1(P2_DATAO_REG_26__SCAN_IN), .A2(n14394), .B1(
        P1_DATAO_REG_26__SCAN_IN), .B2(n15240), .ZN(n9421) );
  INV_X1 U11978 ( .A(n9421), .ZN(n9422) );
  XNOR2_X1 U11979 ( .A(n9432), .B(n9422), .ZN(n13847) );
  NAND2_X1 U11980 ( .A1(n13847), .A2(n9184), .ZN(n9424) );
  NAND2_X1 U11981 ( .A1(n9425), .A2(P3_REG3_REG_26__SCAN_IN), .ZN(n9426) );
  NAND2_X1 U11982 ( .A1(n9438), .A2(n9426), .ZN(n13568) );
  NAND2_X1 U11983 ( .A1(n13568), .A2(n9300), .ZN(n9431) );
  INV_X1 U11984 ( .A(P3_REG1_REG_26__SCAN_IN), .ZN(n13726) );
  NAND2_X1 U11985 ( .A1(n9475), .A2(P3_REG2_REG_26__SCAN_IN), .ZN(n9428) );
  NAND2_X1 U11986 ( .A1(n9476), .A2(P3_REG0_REG_26__SCAN_IN), .ZN(n9427) );
  OAI211_X1 U11987 ( .C1(n9479), .C2(n13726), .A(n9428), .B(n9427), .ZN(n9429)
         );
  INV_X1 U11988 ( .A(n9429), .ZN(n9430) );
  NAND2_X1 U11989 ( .A1(n13338), .A2(n13548), .ZN(n9657) );
  AOI22_X1 U11990 ( .A1(P2_DATAO_REG_27__SCAN_IN), .A2(
        P1_DATAO_REG_27__SCAN_IN), .B1(n12567), .B2(n7339), .ZN(n9433) );
  INV_X1 U11991 ( .A(n9433), .ZN(n9434) );
  XNOR2_X1 U11992 ( .A(n9445), .B(n9434), .ZN(n13844) );
  NAND2_X1 U11993 ( .A1(n13844), .A2(n6668), .ZN(n9437) );
  INV_X1 U11994 ( .A(n9451), .ZN(n9440) );
  NAND2_X1 U11995 ( .A1(n9438), .A2(P3_REG3_REG_27__SCAN_IN), .ZN(n9439) );
  NAND2_X1 U11996 ( .A1(n9440), .A2(n9439), .ZN(n13557) );
  INV_X1 U11997 ( .A(P3_REG1_REG_27__SCAN_IN), .ZN(n9443) );
  NAND2_X1 U11998 ( .A1(n9475), .A2(P3_REG2_REG_27__SCAN_IN), .ZN(n9442) );
  NAND2_X1 U11999 ( .A1(n9476), .A2(P3_REG0_REG_27__SCAN_IN), .ZN(n9441) );
  OAI211_X1 U12000 ( .C1(n9479), .C2(n9443), .A(n9442), .B(n9441), .ZN(n9444)
         );
  OR2_X1 U12001 ( .A1(n13556), .A2(n13565), .ZN(n9660) );
  NAND2_X1 U12002 ( .A1(n13556), .A2(n13565), .ZN(n9662) );
  NOR2_X1 U12003 ( .A1(P1_DATAO_REG_27__SCAN_IN), .A2(n7339), .ZN(n9446) );
  AOI22_X1 U12004 ( .A1(P2_DATAO_REG_28__SCAN_IN), .A2(n14392), .B1(
        P1_DATAO_REG_28__SCAN_IN), .B2(n15236), .ZN(n9447) );
  INV_X1 U12005 ( .A(n9447), .ZN(n9448) );
  XNOR2_X1 U12006 ( .A(n9457), .B(n9448), .ZN(n13172) );
  NAND2_X1 U12007 ( .A1(n13172), .A2(n9184), .ZN(n9450) );
  NAND2_X2 U12008 ( .A1(n9450), .A2(n9449), .ZN(n13540) );
  NOR2_X1 U12009 ( .A1(n9451), .A2(n8142), .ZN(n9452) );
  INV_X1 U12010 ( .A(P3_REG1_REG_28__SCAN_IN), .ZN(n9455) );
  NAND2_X1 U12011 ( .A1(n9475), .A2(P3_REG2_REG_28__SCAN_IN), .ZN(n9454) );
  NAND2_X1 U12012 ( .A1(n9476), .A2(P3_REG0_REG_28__SCAN_IN), .ZN(n9453) );
  OAI211_X1 U12013 ( .C1(n9479), .C2(n9455), .A(n9454), .B(n9453), .ZN(n9456)
         );
  NAND2_X1 U12014 ( .A1(n13540), .A2(n6675), .ZN(n9663) );
  INV_X1 U12015 ( .A(n13537), .ZN(n9523) );
  INV_X1 U12016 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n15232) );
  AOI22_X1 U12017 ( .A1(P2_DATAO_REG_29__SCAN_IN), .A2(
        P1_DATAO_REG_29__SCAN_IN), .B1(n14387), .B2(n15232), .ZN(n9469) );
  INV_X1 U12018 ( .A(n9469), .ZN(n9458) );
  XNOR2_X1 U12019 ( .A(n9470), .B(n9458), .ZN(n13839) );
  NOR2_X1 U12020 ( .A1(n6678), .A2(n13841), .ZN(n9459) );
  AOI21_X2 U12021 ( .B1(n13839), .B2(n6668), .A(n9459), .ZN(n13176) );
  NAND2_X1 U12022 ( .A1(n15304), .A2(n9300), .ZN(n9482) );
  INV_X1 U12023 ( .A(P3_REG1_REG_29__SCAN_IN), .ZN(n9462) );
  NAND2_X1 U12024 ( .A1(n9475), .A2(P3_REG2_REG_29__SCAN_IN), .ZN(n9461) );
  NAND2_X1 U12025 ( .A1(n9476), .A2(P3_REG0_REG_29__SCAN_IN), .ZN(n9460) );
  OAI211_X1 U12026 ( .C1(n9479), .C2(n9462), .A(n9461), .B(n9460), .ZN(n9463)
         );
  INV_X1 U12027 ( .A(n9463), .ZN(n9464) );
  NAND2_X1 U12028 ( .A1(n9482), .A2(n9464), .ZN(n13354) );
  AND2_X1 U12029 ( .A1(n13176), .A2(n13354), .ZN(n9510) );
  INV_X1 U12030 ( .A(n9510), .ZN(n9665) );
  NAND2_X1 U12031 ( .A1(n9738), .A2(n9665), .ZN(n9498) );
  INV_X1 U12032 ( .A(P3_REG1_REG_31__SCAN_IN), .ZN(n15312) );
  NAND2_X1 U12033 ( .A1(n9475), .A2(P3_REG2_REG_31__SCAN_IN), .ZN(n9466) );
  NAND2_X1 U12034 ( .A1(n9476), .A2(P3_REG0_REG_31__SCAN_IN), .ZN(n9465) );
  OAI211_X1 U12035 ( .C1(n9479), .C2(n15312), .A(n9466), .B(n9465), .ZN(n9467)
         );
  INV_X1 U12036 ( .A(n9467), .ZN(n9468) );
  NAND2_X1 U12037 ( .A1(n9482), .A2(n9468), .ZN(n15303) );
  INV_X1 U12038 ( .A(n15303), .ZN(n9494) );
  INV_X1 U12039 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n12862) );
  OAI22_X1 U12040 ( .A1(n12862), .A2(n9487), .B1(P1_DATAO_REG_30__SCAN_IN), 
        .B2(P2_DATAO_REG_30__SCAN_IN), .ZN(n9485) );
  XOR2_X1 U12041 ( .A(n9486), .B(n9485), .Z(n13836) );
  INV_X1 U12042 ( .A(SI_30_), .ZN(n13835) );
  OR2_X1 U12043 ( .A1(n6678), .A2(n13835), .ZN(n9473) );
  OAI21_X1 U12044 ( .B1(n13836), .B2(n9474), .A(n9473), .ZN(n15314) );
  INV_X1 U12045 ( .A(P3_REG1_REG_30__SCAN_IN), .ZN(n15315) );
  NAND2_X1 U12046 ( .A1(n9475), .A2(P3_REG2_REG_30__SCAN_IN), .ZN(n9478) );
  NAND2_X1 U12047 ( .A1(n9476), .A2(P3_REG0_REG_30__SCAN_IN), .ZN(n9477) );
  OAI211_X1 U12048 ( .C1(n9479), .C2(n15315), .A(n9478), .B(n9477), .ZN(n9480)
         );
  INV_X1 U12049 ( .A(n9480), .ZN(n9481) );
  NAND2_X1 U12050 ( .A1(n15314), .A2(n11102), .ZN(n9526) );
  INV_X1 U12051 ( .A(n13176), .ZN(n9483) );
  INV_X1 U12052 ( .A(n13354), .ZN(n13533) );
  INV_X1 U12053 ( .A(n9509), .ZN(n9484) );
  NAND2_X1 U12054 ( .A1(n9526), .A2(n9484), .ZN(n9529) );
  NAND2_X1 U12055 ( .A1(n9486), .A2(n9485), .ZN(n9489) );
  NAND2_X1 U12056 ( .A1(n9489), .A2(n9488), .ZN(n9492) );
  INV_X1 U12057 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n13084) );
  INV_X1 U12058 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n10136) );
  AOI22_X1 U12059 ( .A1(P2_DATAO_REG_31__SCAN_IN), .A2(
        P1_DATAO_REG_31__SCAN_IN), .B1(n13084), .B2(n10136), .ZN(n9490) );
  INV_X1 U12060 ( .A(n9490), .ZN(n9491) );
  NOR2_X1 U12061 ( .A1(n6678), .A2(n7978), .ZN(n9493) );
  AOI211_X1 U12062 ( .C1(n9494), .C2(n15314), .A(n9529), .B(n9668), .ZN(n9497)
         );
  INV_X1 U12063 ( .A(n15309), .ZN(n15305) );
  NAND2_X1 U12064 ( .A1(n15305), .A2(n9494), .ZN(n9496) );
  OR2_X1 U12065 ( .A1(n15314), .A2(n11102), .ZN(n9495) );
  NAND2_X1 U12066 ( .A1(n9496), .A2(n9495), .ZN(n9508) );
  INV_X1 U12067 ( .A(n9499), .ZN(n9500) );
  NAND2_X1 U12068 ( .A1(n9504), .A2(n9506), .ZN(n9502) );
  NAND2_X1 U12069 ( .A1(n9502), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9501) );
  MUX2_X1 U12070 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9501), .S(
        P3_IR_REG_21__SCAN_IN), .Z(n9503) );
  INV_X1 U12071 ( .A(n9504), .ZN(n9505) );
  NAND2_X1 U12072 ( .A1(n9505), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9507) );
  INV_X1 U12073 ( .A(n10926), .ZN(n9767) );
  NAND2_X1 U12074 ( .A1(n10999), .A2(n9767), .ZN(n9732) );
  NAND2_X1 U12075 ( .A1(n11171), .A2(n9767), .ZN(n10591) );
  NAND2_X1 U12076 ( .A1(n9536), .A2(n9535), .ZN(n13615) );
  NAND2_X1 U12077 ( .A1(n9634), .A2(n9633), .ZN(n13650) );
  NAND2_X1 U12078 ( .A1(n9607), .A2(n9606), .ZN(n12266) );
  INV_X1 U12079 ( .A(n9603), .ZN(n9511) );
  AND2_X1 U12080 ( .A1(n9512), .A2(n10939), .ZN(n9540) );
  NOR2_X1 U12081 ( .A1(n6935), .A2(n9540), .ZN(n10584) );
  NAND4_X1 U12082 ( .A1(n10584), .A2(n11755), .A3(n11000), .A4(n11426), .ZN(
        n9514) );
  INV_X1 U12083 ( .A(n11790), .ZN(n9513) );
  NAND2_X1 U12084 ( .A1(n9545), .A2(n9544), .ZN(n15721) );
  NOR4_X1 U12085 ( .A1(n9514), .A2(n9513), .A3(n12034), .A4(n15721), .ZN(n9517) );
  NOR4_X1 U12086 ( .A1(n12016), .A2(n9695), .A3(n11222), .A4(n12005), .ZN(
        n9515) );
  AND4_X1 U12087 ( .A1(n9517), .A2(n9516), .A3(n9515), .A4(n12048), .ZN(n9518)
         );
  NAND4_X1 U12088 ( .A1(n13677), .A2(n7647), .A3(n7736), .A4(n9518), .ZN(n9519) );
  NOR4_X1 U12089 ( .A1(n13650), .A2(n7645), .A3(n13689), .A4(n9519), .ZN(n9520) );
  NAND4_X1 U12090 ( .A1(n9636), .A2(n13662), .A3(n13627), .A4(n9520), .ZN(
        n9521) );
  NAND4_X1 U12091 ( .A1(n13574), .A2(n13592), .A3(n9739), .A4(n9522), .ZN(
        n9524) );
  INV_X1 U12092 ( .A(n13552), .ZN(n13546) );
  NOR3_X1 U12093 ( .A1(n9524), .A2(n9523), .A3(n13546), .ZN(n9527) );
  INV_X1 U12094 ( .A(n9668), .ZN(n9525) );
  NAND4_X1 U12095 ( .A1(n9669), .A2(n9527), .A3(n9526), .A4(n9525), .ZN(n9528)
         );
  XNOR2_X1 U12096 ( .A(n9528), .B(n9671), .ZN(n9672) );
  INV_X1 U12097 ( .A(n9529), .ZN(n9667) );
  NAND2_X1 U12098 ( .A1(n9674), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9530) );
  AOI21_X1 U12099 ( .B1(n9532), .B2(n9531), .A(n10746), .ZN(n9534) );
  MUX2_X1 U12100 ( .A(n10746), .B(n9534), .S(n9533), .Z(n9650) );
  MUX2_X1 U12101 ( .A(n9536), .B(n9535), .S(n9771), .Z(n9645) );
  MUX2_X1 U12102 ( .A(n9538), .B(n9537), .S(n10746), .Z(n9643) );
  NAND2_X1 U12103 ( .A1(n9544), .A2(n9771), .ZN(n9539) );
  OAI21_X1 U12104 ( .B1(n15721), .B2(n9540), .A(n9539), .ZN(n9543) );
  INV_X1 U12105 ( .A(n9540), .ZN(n9541) );
  OAI211_X1 U12106 ( .C1(n6935), .C2(n10999), .A(n9541), .B(n9771), .ZN(n9542)
         );
  NAND2_X1 U12107 ( .A1(n9543), .A2(n9542), .ZN(n9547) );
  MUX2_X1 U12108 ( .A(n9545), .B(n9544), .S(n10746), .Z(n9546) );
  NAND3_X1 U12109 ( .A1(n9547), .A2(n11053), .A3(n9546), .ZN(n9551) );
  NAND2_X1 U12110 ( .A1(n9556), .A2(n9548), .ZN(n9549) );
  NAND2_X1 U12111 ( .A1(n9549), .A2(n9771), .ZN(n9550) );
  NAND2_X1 U12112 ( .A1(n9551), .A2(n9550), .ZN(n9555) );
  NAND2_X1 U12113 ( .A1(n15718), .A2(n10674), .ZN(n9552) );
  AOI21_X1 U12114 ( .B1(n9554), .B2(n9552), .A(n9771), .ZN(n9553) );
  AOI21_X1 U12115 ( .B1(n9555), .B2(n9554), .A(n9553), .ZN(n9561) );
  OAI21_X1 U12116 ( .B1(n9771), .B2(n9556), .A(n11218), .ZN(n9560) );
  NAND2_X1 U12117 ( .A1(n11425), .A2(n10746), .ZN(n9558) );
  NAND2_X1 U12118 ( .A1(n11301), .A2(n9771), .ZN(n9557) );
  MUX2_X1 U12119 ( .A(n9558), .B(n9557), .S(n9087), .Z(n9559) );
  OAI211_X1 U12120 ( .C1(n9561), .C2(n9560), .A(n11426), .B(n9559), .ZN(n9565)
         );
  NAND2_X1 U12121 ( .A1(n9570), .A2(n9562), .ZN(n9563) );
  NAND2_X1 U12122 ( .A1(n9563), .A2(n10746), .ZN(n9564) );
  NAND2_X1 U12123 ( .A1(n9565), .A2(n9564), .ZN(n9569) );
  AOI21_X1 U12124 ( .B1(n9568), .B2(n9566), .A(n10746), .ZN(n9567) );
  AOI21_X1 U12125 ( .B1(n9569), .B2(n9568), .A(n9567), .ZN(n9572) );
  NOR2_X1 U12126 ( .A1(n9570), .A2(n10746), .ZN(n9571) );
  OR3_X1 U12127 ( .A1(n9572), .A2(n9571), .A3(n11749), .ZN(n9576) );
  MUX2_X1 U12128 ( .A(n9574), .B(n9573), .S(n9771), .Z(n9575) );
  NAND3_X1 U12129 ( .A1(n9576), .A2(n12023), .A3(n9575), .ZN(n9581) );
  INV_X1 U12130 ( .A(n12034), .ZN(n9580) );
  NAND2_X1 U12131 ( .A1(n11855), .A2(n9771), .ZN(n9578) );
  NAND2_X1 U12132 ( .A1(n12173), .A2(n10746), .ZN(n9577) );
  MUX2_X1 U12133 ( .A(n9578), .B(n9577), .S(n13357), .Z(n9579) );
  NAND3_X1 U12134 ( .A1(n9581), .A2(n9580), .A3(n9579), .ZN(n9585) );
  NAND2_X1 U12135 ( .A1(n12018), .A2(n9582), .ZN(n9703) );
  MUX2_X1 U12136 ( .A(n12018), .B(n9582), .S(n10746), .Z(n9583) );
  AOI21_X1 U12137 ( .B1(n9703), .B2(n9583), .A(n12005), .ZN(n9584) );
  NAND3_X1 U12138 ( .A1(n9585), .A2(n9584), .A3(n12048), .ZN(n9592) );
  INV_X1 U12139 ( .A(n9586), .ZN(n9587) );
  NAND2_X1 U12140 ( .A1(n12048), .A2(n9587), .ZN(n9589) );
  NAND3_X1 U12141 ( .A1(n9589), .A2(n9598), .A3(n9588), .ZN(n9590) );
  NAND2_X1 U12142 ( .A1(n9590), .A2(n9771), .ZN(n9591) );
  NAND2_X1 U12143 ( .A1(n9592), .A2(n9591), .ZN(n9597) );
  NAND2_X1 U12144 ( .A1(n12048), .A2(n7473), .ZN(n9594) );
  OAI211_X1 U12145 ( .C1(n12377), .C2(n12143), .A(n9594), .B(n9596), .ZN(n9595) );
  AOI22_X1 U12146 ( .A1(n9597), .A2(n9596), .B1(n10746), .B2(n9595), .ZN(n9600) );
  NOR2_X1 U12147 ( .A1(n9598), .A2(n9771), .ZN(n9599) );
  OAI21_X1 U12148 ( .B1(n9600), .B2(n9599), .A(n7736), .ZN(n9605) );
  INV_X1 U12149 ( .A(n9601), .ZN(n9602) );
  MUX2_X1 U12150 ( .A(n9603), .B(n9602), .S(n10746), .Z(n9604) );
  NAND3_X1 U12151 ( .A1(n9605), .A2(n7647), .A3(n9604), .ZN(n9609) );
  MUX2_X1 U12152 ( .A(n9607), .B(n9606), .S(n10746), .Z(n9608) );
  NAND3_X1 U12153 ( .A1(n9609), .A2(n13710), .A3(n9608), .ZN(n9614) );
  NAND2_X1 U12154 ( .A1(n9617), .A2(n9610), .ZN(n9611) );
  NAND2_X1 U12155 ( .A1(n9611), .A2(n9771), .ZN(n9613) );
  INV_X1 U12156 ( .A(n9616), .ZN(n9612) );
  AOI21_X1 U12157 ( .B1(n9614), .B2(n9613), .A(n9612), .ZN(n9619) );
  AOI21_X1 U12158 ( .B1(n9616), .B2(n9615), .A(n9771), .ZN(n9618) );
  OAI22_X1 U12159 ( .A1(n9619), .A2(n9618), .B1(n9771), .B2(n9617), .ZN(n9627)
         );
  INV_X1 U12160 ( .A(n9620), .ZN(n9626) );
  INV_X1 U12161 ( .A(n9621), .ZN(n9622) );
  NAND2_X1 U12162 ( .A1(n9628), .A2(n9622), .ZN(n9624) );
  AND3_X1 U12163 ( .A1(n9624), .A2(n10746), .A3(n9623), .ZN(n9625) );
  NAND2_X1 U12164 ( .A1(n9625), .A2(n9633), .ZN(n9629) );
  AOI22_X1 U12165 ( .A1(n9627), .A2(n13677), .B1(n9626), .B2(n9629), .ZN(n9632) );
  NAND3_X1 U12166 ( .A1(n9634), .A2(n9771), .A3(n9628), .ZN(n9630) );
  NAND2_X1 U12167 ( .A1(n9630), .A2(n9629), .ZN(n9631) );
  OAI21_X1 U12168 ( .B1(n9632), .B2(n7651), .A(n9631), .ZN(n9637) );
  MUX2_X1 U12169 ( .A(n9634), .B(n9633), .S(n9771), .Z(n9635) );
  NAND3_X1 U12170 ( .A1(n9637), .A2(n9636), .A3(n9635), .ZN(n9641) );
  MUX2_X1 U12171 ( .A(n9639), .B(n9638), .S(n9771), .Z(n9640) );
  NAND3_X1 U12172 ( .A1(n9641), .A2(n13627), .A3(n9640), .ZN(n9642) );
  NAND3_X1 U12173 ( .A1(n7624), .A2(n9643), .A3(n9642), .ZN(n9644) );
  NAND3_X1 U12174 ( .A1(n9645), .A2(n9721), .A3(n9644), .ZN(n9647) );
  NAND3_X1 U12175 ( .A1(n13239), .A2(n13613), .A3(n10746), .ZN(n9646) );
  NAND2_X1 U12176 ( .A1(n9647), .A2(n9646), .ZN(n9648) );
  AND2_X1 U12177 ( .A1(n13592), .A2(n9648), .ZN(n9649) );
  NOR2_X1 U12178 ( .A1(n9650), .A2(n9649), .ZN(n9655) );
  MUX2_X1 U12179 ( .A(n9652), .B(n9651), .S(n9771), .Z(n9653) );
  INV_X1 U12180 ( .A(n9653), .ZN(n9654) );
  AOI21_X1 U12181 ( .B1(n9655), .B2(n13574), .A(n9654), .ZN(n9659) );
  MUX2_X1 U12182 ( .A(n9657), .B(n9656), .S(n10746), .Z(n9658) );
  OAI211_X1 U12183 ( .C1(n9659), .C2(n13567), .A(n13552), .B(n9658), .ZN(n9664) );
  NAND2_X1 U12184 ( .A1(n9664), .A2(n9660), .ZN(n9661) );
  AOI21_X1 U12185 ( .B1(n9670), .B2(n9669), .A(n9668), .ZN(n9673) );
  OR2_X1 U12186 ( .A1(n10745), .A2(P3_U3151), .ZN(n11598) );
  INV_X1 U12187 ( .A(n11598), .ZN(n9677) );
  NOR2_X1 U12188 ( .A1(n10594), .A2(n9771), .ZN(n10583) );
  INV_X1 U12189 ( .A(n9679), .ZN(n9680) );
  INV_X1 U12190 ( .A(n12180), .ZN(n9687) );
  OR2_X1 U12191 ( .A1(n9683), .A2(n9682), .ZN(n9685) );
  INV_X1 U12192 ( .A(n12124), .ZN(n9686) );
  NAND3_X1 U12193 ( .A1(n9687), .A2(n9748), .A3(n9686), .ZN(n10500) );
  NAND2_X1 U12194 ( .A1(n10583), .A2(n10934), .ZN(n10601) );
  NOR3_X1 U12195 ( .A1(n10601), .A2(n13517), .A3(n9689), .ZN(n9691) );
  OAI21_X1 U12196 ( .B1(n11598), .B2(n11285), .A(P3_B_REG_SCAN_IN), .ZN(n9690)
         );
  OR2_X1 U12197 ( .A1(n9691), .A2(n9690), .ZN(n9692) );
  INV_X1 U12198 ( .A(n13670), .ZN(n13760) );
  NAND2_X1 U12199 ( .A1(n9512), .A2(n9693), .ZN(n15720) );
  NAND2_X1 U12200 ( .A1(n6957), .A2(n15714), .ZN(n9694) );
  NAND2_X1 U12201 ( .A1(n7742), .A2(n9696), .ZN(n11001) );
  NAND2_X1 U12202 ( .A1(n10625), .A2(n10830), .ZN(n9697) );
  NAND2_X1 U12203 ( .A1(n11001), .A2(n9697), .ZN(n11223) );
  NAND2_X1 U12204 ( .A1(n11425), .A2(n9087), .ZN(n9698) );
  NAND2_X1 U12205 ( .A1(n11792), .A2(n15753), .ZN(n9699) );
  NAND2_X1 U12206 ( .A1(n11422), .A2(n9699), .ZN(n11791) );
  INV_X1 U12207 ( .A(n11791), .ZN(n9700) );
  NAND2_X1 U12208 ( .A1(n11751), .A2(n15708), .ZN(n11748) );
  NAND2_X1 U12209 ( .A1(n12145), .A2(n15766), .ZN(n9702) );
  AND2_X1 U12210 ( .A1(n12000), .A2(n9702), .ZN(n9701) );
  NAND2_X1 U12211 ( .A1(n12017), .A2(n11896), .ZN(n11998) );
  AND2_X1 U12212 ( .A1(n11748), .A2(n9706), .ZN(n9711) );
  INV_X1 U12213 ( .A(n9702), .ZN(n9705) );
  INV_X1 U12214 ( .A(n9703), .ZN(n9704) );
  NAND2_X1 U12215 ( .A1(n11640), .A2(n12173), .ZN(n12030) );
  INV_X1 U12216 ( .A(n9706), .ZN(n9707) );
  NAND2_X1 U12217 ( .A1(n13356), .A2(n15325), .ZN(n9712) );
  OAI21_X1 U12218 ( .B1(n15318), .B2(n13355), .A(n12193), .ZN(n9714) );
  NAND2_X1 U12219 ( .A1(n13355), .A2(n15318), .ZN(n9713) );
  INV_X1 U12220 ( .A(n13824), .ZN(n13232) );
  INV_X1 U12221 ( .A(n13187), .ZN(n13772) );
  OAI22_X1 U12222 ( .A1(n13678), .A2(n13677), .B1(n13695), .B2(n13295), .ZN(
        n13661) );
  NAND2_X1 U12223 ( .A1(n13636), .A2(n13641), .ZN(n9717) );
  NAND2_X1 U12224 ( .A1(n9717), .A2(n7728), .ZN(n13626) );
  NAND2_X1 U12225 ( .A1(n13805), .A2(n13638), .ZN(n9718) );
  NAND2_X1 U12226 ( .A1(n13801), .A2(n13630), .ZN(n9719) );
  NAND2_X1 U12227 ( .A1(n7747), .A2(n13602), .ZN(n13601) );
  OAI21_X1 U12228 ( .B1(n13613), .B2(n13797), .A(n13601), .ZN(n13588) );
  NAND2_X1 U12229 ( .A1(n13563), .A2(n9724), .ZN(n9727) );
  INV_X1 U12230 ( .A(n13567), .ZN(n9725) );
  NAND2_X1 U12231 ( .A1(n9725), .A2(n13338), .ZN(n9726) );
  NAND2_X1 U12232 ( .A1(n13782), .A2(n13565), .ZN(n9728) );
  NAND2_X1 U12233 ( .A1(n13535), .A2(n9730), .ZN(n9731) );
  XNOR2_X1 U12234 ( .A(n9731), .B(n9739), .ZN(n9737) );
  NAND2_X1 U12235 ( .A1(n9769), .A2(n11285), .ZN(n9777) );
  NAND2_X1 U12236 ( .A1(n10750), .A2(n13517), .ZN(n10760) );
  NAND2_X1 U12237 ( .A1(n10760), .A2(n10748), .ZN(n10600) );
  NOR2_X1 U12238 ( .A1(n9689), .A2(n9734), .ZN(n9735) );
  OR2_X1 U12239 ( .A1(n13696), .A2(n9735), .ZN(n15301) );
  OAI22_X1 U12240 ( .A1(n6675), .A2(n13694), .B1(n11102), .B2(n15301), .ZN(
        n9736) );
  NAND2_X1 U12241 ( .A1(n9671), .A2(n11171), .ZN(n9742) );
  NAND2_X1 U12242 ( .A1(n11171), .A2(n10926), .ZN(n9740) );
  XNOR2_X1 U12243 ( .A(n11285), .B(n9740), .ZN(n9741) );
  NAND2_X1 U12244 ( .A1(n9742), .A2(n9741), .ZN(n10508) );
  INV_X1 U12245 ( .A(n10594), .ZN(n9743) );
  NAND3_X1 U12246 ( .A1(n10508), .A2(n9743), .A3(n15758), .ZN(n9744) );
  OR3_X1 U12247 ( .A1(n9769), .A2(n9768), .A3(n10926), .ZN(n9772) );
  NAND2_X1 U12248 ( .A1(n13178), .A2(n15316), .ZN(n9745) );
  NAND2_X1 U12249 ( .A1(n13174), .A2(n9745), .ZN(n9784) );
  XNOR2_X1 U12250 ( .A(n12124), .B(P3_B_REG_SCAN_IN), .ZN(n9746) );
  INV_X1 U12251 ( .A(P3_D_REG_1__SCAN_IN), .ZN(n9747) );
  NAND2_X1 U12252 ( .A1(n9752), .A2(n9747), .ZN(n9750) );
  NAND2_X1 U12253 ( .A1(n13848), .A2(n12180), .ZN(n9749) );
  INV_X1 U12254 ( .A(P3_D_REG_0__SCAN_IN), .ZN(n9751) );
  XNOR2_X1 U12255 ( .A(n10592), .B(n13827), .ZN(n9766) );
  NOR2_X1 U12256 ( .A1(P3_D_REG_17__SCAN_IN), .A2(P3_D_REG_22__SCAN_IN), .ZN(
        n9758) );
  NOR4_X1 U12257 ( .A1(P3_D_REG_2__SCAN_IN), .A2(P3_D_REG_8__SCAN_IN), .A3(
        P3_D_REG_25__SCAN_IN), .A4(P3_D_REG_20__SCAN_IN), .ZN(n9757) );
  NOR4_X1 U12258 ( .A1(P3_D_REG_29__SCAN_IN), .A2(P3_D_REG_10__SCAN_IN), .A3(
        P3_D_REG_31__SCAN_IN), .A4(P3_D_REG_14__SCAN_IN), .ZN(n9756) );
  NOR4_X1 U12259 ( .A1(P3_D_REG_19__SCAN_IN), .A2(P3_D_REG_18__SCAN_IN), .A3(
        P3_D_REG_27__SCAN_IN), .A4(P3_D_REG_24__SCAN_IN), .ZN(n9755) );
  NAND4_X1 U12260 ( .A1(n9758), .A2(n9757), .A3(n9756), .A4(n9755), .ZN(n9764)
         );
  NOR4_X1 U12261 ( .A1(P3_D_REG_9__SCAN_IN), .A2(P3_D_REG_16__SCAN_IN), .A3(
        P3_D_REG_15__SCAN_IN), .A4(P3_D_REG_30__SCAN_IN), .ZN(n9762) );
  NOR4_X1 U12262 ( .A1(P3_D_REG_11__SCAN_IN), .A2(P3_D_REG_21__SCAN_IN), .A3(
        P3_D_REG_12__SCAN_IN), .A4(P3_D_REG_26__SCAN_IN), .ZN(n9761) );
  NOR4_X1 U12263 ( .A1(P3_D_REG_3__SCAN_IN), .A2(P3_D_REG_5__SCAN_IN), .A3(
        P3_D_REG_4__SCAN_IN), .A4(P3_D_REG_7__SCAN_IN), .ZN(n9760) );
  NOR4_X1 U12264 ( .A1(P3_D_REG_13__SCAN_IN), .A2(P3_D_REG_28__SCAN_IN), .A3(
        P3_D_REG_23__SCAN_IN), .A4(P3_D_REG_6__SCAN_IN), .ZN(n9759) );
  NAND4_X1 U12265 ( .A1(n9762), .A2(n9761), .A3(n9760), .A4(n9759), .ZN(n9763)
         );
  OAI21_X1 U12266 ( .B1(n9764), .B2(n9763), .A(n9752), .ZN(n9780) );
  AND2_X1 U12267 ( .A1(n10934), .A2(n9780), .ZN(n9765) );
  OAI22_X1 U12268 ( .A1(n9769), .A2(n9768), .B1(n9767), .B2(n15758), .ZN(n9770) );
  AOI21_X1 U12269 ( .B1(n9770), .B2(n10594), .A(n10746), .ZN(n9774) );
  NAND2_X1 U12270 ( .A1(n10594), .A2(n10746), .ZN(n10501) );
  NAND2_X1 U12271 ( .A1(n9772), .A2(n9771), .ZN(n10929) );
  NAND2_X1 U12272 ( .A1(n10501), .A2(n10929), .ZN(n10927) );
  NAND2_X1 U12273 ( .A1(n10927), .A2(n13827), .ZN(n9773) );
  OAI21_X1 U12274 ( .B1(n9774), .B2(n13827), .A(n9773), .ZN(n9775) );
  INV_X1 U12275 ( .A(n9775), .ZN(n9776) );
  AND3_X1 U12276 ( .A1(n6960), .A2(n13827), .A3(n9780), .ZN(n10513) );
  NOR2_X1 U12277 ( .A1(n9777), .A2(n10591), .ZN(n10509) );
  NAND2_X1 U12278 ( .A1(n10509), .A2(n10934), .ZN(n9778) );
  NAND2_X1 U12279 ( .A1(n10601), .A2(n9778), .ZN(n9779) );
  NAND2_X1 U12280 ( .A1(n10513), .A2(n9779), .ZN(n9783) );
  NAND2_X1 U12281 ( .A1(n10592), .A2(n9780), .ZN(n9781) );
  NAND3_X1 U12282 ( .A1(n10602), .A2(n10934), .A3(n10508), .ZN(n9782) );
  INV_X1 U12283 ( .A(n9785), .ZN(n9786) );
  OR2_X1 U12284 ( .A1(n15773), .A2(n15758), .ZN(n13825) );
  NAND2_X1 U12285 ( .A1(n9786), .A2(n7727), .ZN(P3_U3456) );
  INV_X1 U12286 ( .A(n9787), .ZN(n9788) );
  NAND2_X1 U12287 ( .A1(n9788), .A2(n12058), .ZN(n10079) );
  NOR2_X1 U12288 ( .A1(P1_IR_REG_5__SCAN_IN), .A2(P1_IR_REG_14__SCAN_IN), .ZN(
        n9790) );
  NAND4_X1 U12289 ( .A1(n10241), .A2(n9790), .A3(n10244), .A4(n10004), .ZN(
        n9792) );
  NOR2_X1 U12290 ( .A1(P1_IR_REG_25__SCAN_IN), .A2(P1_IR_REG_24__SCAN_IN), 
        .ZN(n9802) );
  NOR2_X1 U12291 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(P1_IR_REG_21__SCAN_IN), 
        .ZN(n9801) );
  NAND4_X1 U12292 ( .A1(n9802), .A2(n9801), .A3(n9810), .A4(n9829), .ZN(n9803)
         );
  INV_X1 U12293 ( .A(n9807), .ZN(n9804) );
  NAND2_X1 U12294 ( .A1(n9804), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9805) );
  MUX2_X1 U12295 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9805), .S(
        P1_IR_REG_26__SCAN_IN), .Z(n9808) );
  INV_X1 U12296 ( .A(n9814), .ZN(n9833) );
  NAND2_X1 U12297 ( .A1(n9900), .A2(n9905), .ZN(n9809) );
  NAND2_X1 U12298 ( .A1(n6823), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9811) );
  INV_X1 U12299 ( .A(n10500), .ZN(n9812) );
  XNOR2_X2 U12300 ( .A(n9818), .B(n9817), .ZN(n15234) );
  INV_X1 U12301 ( .A(n15234), .ZN(n9819) );
  INV_X1 U12302 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n14743) );
  NAND2_X1 U12303 ( .A1(n6677), .A2(n14743), .ZN(n9825) );
  NAND2_X1 U12304 ( .A1(n9865), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n9824) );
  NAND2_X1 U12305 ( .A1(n6878), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n9823) );
  NAND2_X1 U12306 ( .A1(n9864), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n9822) );
  AND4_X2 U12307 ( .A1(n9825), .A2(n9824), .A3(n9823), .A4(n9822), .ZN(n10954)
         );
  NAND2_X1 U12308 ( .A1(n9828), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9830) );
  NAND2_X4 U12309 ( .A1(n9844), .A2(n12592), .ZN(n14557) );
  XNOR2_X2 U12310 ( .A(n9832), .B(n9831), .ZN(n9941) );
  NAND2_X1 U12311 ( .A1(n9833), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9834) );
  INV_X1 U12312 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n9963) );
  OR2_X1 U12313 ( .A1(n9888), .A2(n9963), .ZN(n9843) );
  NAND2_X1 U12314 ( .A1(n9840), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9841) );
  XNOR2_X1 U12315 ( .A(n9841), .B(n9789), .ZN(n14750) );
  OAI22_X1 U12316 ( .A1(n10954), .A2(n14557), .B1(n11538), .B2(n6667), .ZN(
        n9852) );
  NAND2_X1 U12317 ( .A1(n11257), .A2(n9846), .ZN(n11260) );
  NAND2_X1 U12318 ( .A1(n12593), .A2(n15244), .ZN(n9849) );
  NAND2_X2 U12319 ( .A1(n9850), .A2(n9849), .ZN(n14445) );
  NOR2_X4 U12320 ( .A1(n9920), .A2(n12787), .ZN(n15291) );
  OAI22_X1 U12321 ( .A1(n10954), .A2(n6950), .B1(n11538), .B2(n14557), .ZN(
        n11023) );
  XNOR2_X1 U12322 ( .A(n11024), .B(n11023), .ZN(n9925) );
  NAND2_X1 U12323 ( .A1(n6680), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n9854) );
  NAND2_X1 U12324 ( .A1(n9880), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n9853) );
  NAND2_X1 U12325 ( .A1(n9865), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n9856) );
  AND2_X1 U12326 ( .A1(n9856), .A2(n9855), .ZN(n9857) );
  INV_X1 U12327 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n9859) );
  NAND2_X1 U12328 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), 
        .ZN(n9858) );
  XNOR2_X1 U12329 ( .A(n9859), .B(n9858), .ZN(n14710) );
  XNOR2_X1 U12330 ( .A(n9860), .B(n14445), .ZN(n9862) );
  OAI22_X1 U12331 ( .A1(n15092), .A2(n14555), .B1(n10686), .B2(n14557), .ZN(
        n9861) );
  NAND2_X1 U12332 ( .A1(n9864), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n9869) );
  NAND2_X1 U12333 ( .A1(n14707), .A2(n6676), .ZN(n9876) );
  INV_X1 U12334 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n14712) );
  INV_X1 U12335 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n9870) );
  OAI21_X1 U12336 ( .B1(n9950), .B2(n9953), .A(n9870), .ZN(n9871) );
  NAND2_X1 U12337 ( .A1(n9872), .A2(n9871), .ZN(n15245) );
  MUX2_X1 U12338 ( .A(n14712), .B(n15245), .S(n12448), .Z(n12591) );
  INV_X1 U12339 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n9873) );
  OAI22_X1 U12340 ( .A1(n6667), .A2(n12591), .B1(n9928), .B2(n9873), .ZN(n9874) );
  INV_X1 U12341 ( .A(n9874), .ZN(n9875) );
  NAND2_X1 U12342 ( .A1(n9876), .A2(n9875), .ZN(n10437) );
  INV_X4 U12343 ( .A(n14555), .ZN(n14517) );
  OAI22_X1 U12344 ( .A1(n14557), .A2(n12591), .B1(n9928), .B2(n14712), .ZN(
        n9877) );
  INV_X1 U12345 ( .A(n9878), .ZN(n9879) );
  NAND2_X1 U12346 ( .A1(n6681), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n9884) );
  NAND2_X1 U12347 ( .A1(n9865), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n9883) );
  NAND2_X1 U12348 ( .A1(n6878), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n9882) );
  NAND2_X1 U12349 ( .A1(n6677), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n9881) );
  INV_X2 U12350 ( .A(n10689), .ZN(n10688) );
  OR2_X1 U12351 ( .A1(n9885), .A2(n15227), .ZN(n9887) );
  XNOR2_X1 U12352 ( .A(n9887), .B(n9886), .ZN(n14734) );
  INV_X1 U12353 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n9962) );
  OR2_X1 U12354 ( .A1(n9889), .A2(n9976), .ZN(n9890) );
  OAI22_X1 U12355 ( .A1(n10688), .A2(n14557), .B1(n11544), .B2(n6667), .ZN(
        n9892) );
  NAND2_X1 U12356 ( .A1(n10689), .A2(n14517), .ZN(n9895) );
  NAND2_X1 U12357 ( .A1(n9893), .A2(n6669), .ZN(n9894) );
  NAND2_X1 U12358 ( .A1(n9895), .A2(n9894), .ZN(n9897) );
  OR2_X1 U12359 ( .A1(n9898), .A2(n9897), .ZN(n9899) );
  INV_X1 U12360 ( .A(n9906), .ZN(n12321) );
  NAND3_X1 U12361 ( .A1(n12321), .A2(n12387), .A3(P1_B_REG_SCAN_IN), .ZN(n9904) );
  INV_X1 U12362 ( .A(P1_B_REG_SCAN_IN), .ZN(n9902) );
  AOI21_X1 U12363 ( .B1(n9906), .B2(n9902), .A(n15242), .ZN(n9903) );
  OR2_X1 U12364 ( .A1(n10018), .A2(P1_D_REG_0__SCAN_IN), .ZN(n9907) );
  OR2_X1 U12365 ( .A1(n10018), .A2(P1_D_REG_1__SCAN_IN), .ZN(n9908) );
  NAND2_X1 U12366 ( .A1(n12387), .A2(n15242), .ZN(n10022) );
  NAND2_X1 U12367 ( .A1(n9908), .A2(n10022), .ZN(n11199) );
  NOR2_X1 U12368 ( .A1(n10711), .A2(n11199), .ZN(n9940) );
  NOR4_X1 U12369 ( .A1(P1_D_REG_18__SCAN_IN), .A2(P1_D_REG_19__SCAN_IN), .A3(
        P1_D_REG_20__SCAN_IN), .A4(P1_D_REG_21__SCAN_IN), .ZN(n9912) );
  NOR4_X1 U12370 ( .A1(P1_D_REG_16__SCAN_IN), .A2(P1_D_REG_14__SCAN_IN), .A3(
        P1_D_REG_15__SCAN_IN), .A4(P1_D_REG_17__SCAN_IN), .ZN(n9911) );
  NOR4_X1 U12371 ( .A1(P1_D_REG_26__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n9910) );
  NOR4_X1 U12372 ( .A1(P1_D_REG_22__SCAN_IN), .A2(P1_D_REG_23__SCAN_IN), .A3(
        P1_D_REG_24__SCAN_IN), .A4(P1_D_REG_25__SCAN_IN), .ZN(n9909) );
  NAND4_X1 U12373 ( .A1(n9912), .A2(n9911), .A3(n9910), .A4(n9909), .ZN(n9918)
         );
  NOR2_X1 U12374 ( .A1(P1_D_REG_2__SCAN_IN), .A2(P1_D_REG_3__SCAN_IN), .ZN(
        n9916) );
  NOR4_X1 U12375 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        P1_D_REG_4__SCAN_IN), .A4(P1_D_REG_5__SCAN_IN), .ZN(n9915) );
  NOR4_X1 U12376 ( .A1(P1_D_REG_10__SCAN_IN), .A2(P1_D_REG_11__SCAN_IN), .A3(
        P1_D_REG_12__SCAN_IN), .A4(P1_D_REG_13__SCAN_IN), .ZN(n9914) );
  NOR4_X1 U12377 ( .A1(P1_D_REG_6__SCAN_IN), .A2(P1_D_REG_7__SCAN_IN), .A3(
        P1_D_REG_8__SCAN_IN), .A4(P1_D_REG_9__SCAN_IN), .ZN(n9913) );
  NAND4_X1 U12378 ( .A1(n9916), .A2(n9915), .A3(n9914), .A4(n9913), .ZN(n9917)
         );
  NOR2_X1 U12379 ( .A1(n9918), .A2(n9917), .ZN(n9919) );
  OR2_X1 U12380 ( .A1(n10018), .A2(n9919), .ZN(n9937) );
  NAND2_X1 U12381 ( .A1(n9940), .A2(n9937), .ZN(n9926) );
  INV_X1 U12382 ( .A(n9926), .ZN(n9934) );
  INV_X1 U12383 ( .A(n10182), .ZN(n9935) );
  INV_X1 U12384 ( .A(n9920), .ZN(n15486) );
  NAND2_X1 U12385 ( .A1(n15486), .A2(n12787), .ZN(n9933) );
  NAND2_X1 U12386 ( .A1(n15486), .A2(n15048), .ZN(n9921) );
  NAND2_X1 U12387 ( .A1(n15244), .A2(n12594), .ZN(n12784) );
  INV_X1 U12388 ( .A(n12784), .ZN(n10184) );
  OR2_X1 U12389 ( .A1(n15495), .A2(n10184), .ZN(n9922) );
  NOR2_X1 U12390 ( .A1(n9935), .A2(n9922), .ZN(n9923) );
  AOI211_X1 U12391 ( .C1(n9925), .C2(n9924), .A(n15392), .B(n11079), .ZN(n9949) );
  NAND2_X1 U12392 ( .A1(n15291), .A2(n15048), .ZN(n10684) );
  NAND2_X1 U12393 ( .A1(n9926), .A2(n10684), .ZN(n9930) );
  OAI21_X1 U12394 ( .B1(n15048), .B2(n12787), .A(n10184), .ZN(n9927) );
  NAND2_X1 U12395 ( .A1(n9928), .A2(n9927), .ZN(n12841) );
  INV_X1 U12396 ( .A(n12841), .ZN(n9929) );
  NAND2_X1 U12397 ( .A1(n9930), .A2(n9929), .ZN(n10439) );
  NAND2_X1 U12398 ( .A1(n10439), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9932) );
  INV_X1 U12399 ( .A(n10183), .ZN(n9931) );
  NAND2_X1 U12400 ( .A1(n9931), .A2(P1_STATE_REG_SCAN_IN), .ZN(n12844) );
  MUX2_X1 U12401 ( .A(n14680), .B(P1_U3086), .S(P1_REG3_REG_3__SCAN_IN), .Z(
        n9948) );
  INV_X1 U12402 ( .A(n9933), .ZN(n11203) );
  NAND3_X1 U12403 ( .A1(n9934), .A2(n11203), .A3(n10182), .ZN(n9936) );
  NOR2_X1 U12404 ( .A1(n14683), .A2(n11538), .ZN(n9947) );
  NOR2_X1 U12405 ( .A1(n12841), .A2(n12840), .ZN(n9938) );
  NAND2_X1 U12406 ( .A1(n9938), .A2(n9937), .ZN(n11200) );
  INV_X1 U12407 ( .A(n11200), .ZN(n9939) );
  NAND2_X1 U12408 ( .A1(n9940), .A2(n9939), .ZN(n14668) );
  INV_X1 U12409 ( .A(n9941), .ZN(n14721) );
  NOR2_X2 U12410 ( .A1(n14668), .A2(n15069), .ZN(n14677) );
  INV_X1 U12411 ( .A(n14677), .ZN(n15387) );
  NAND2_X1 U12412 ( .A1(n9864), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n9945) );
  NAND2_X1 U12413 ( .A1(n6878), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n9944) );
  XNOR2_X1 U12414 ( .A(n14743), .B(P1_REG3_REG_4__SCAN_IN), .ZN(n11204) );
  NAND2_X1 U12415 ( .A1(n6677), .A2(n11204), .ZN(n9943) );
  NAND2_X1 U12416 ( .A1(n9865), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n9942) );
  INV_X1 U12417 ( .A(n14668), .ZN(n14574) );
  OAI22_X1 U12418 ( .A1(n15387), .A2(n10688), .B1(n11529), .B2(n15384), .ZN(
        n9946) );
  OR4_X1 U12419 ( .A1(n9949), .A2(n9948), .A3(n9947), .A4(n9946), .ZN(P1_U3218) );
  INV_X2 U12420 ( .A(n12056), .ZN(n15238) );
  OAI222_X1 U12421 ( .A1(n15239), .A2(n8234), .B1(n15238), .B2(n9981), .C1(
        n14710), .C2(P1_U3086), .ZN(P1_U3354) );
  NOR2_X1 U12422 ( .A1(n9975), .A2(P3_STATE_REG_SCAN_IN), .ZN(n13828) );
  INV_X2 U12423 ( .A(n13828), .ZN(n13851) );
  AND2_X1 U12424 ( .A1(n9975), .A2(P3_U3151), .ZN(n9964) );
  AOI22_X1 U12425 ( .A1(n10986), .A2(P3_STATE_REG_SCAN_IN), .B1(SI_7_), .B2(
        n9964), .ZN(n9951) );
  OAI21_X1 U12426 ( .B1(n9952), .B2(n13851), .A(n9951), .ZN(P3_U3288) );
  INV_X2 U12427 ( .A(n9964), .ZN(n13840) );
  OAI222_X1 U12428 ( .A1(n13851), .A2(n7734), .B1(n13840), .B2(n9953), .C1(
        P3_U3151), .C2(n10763), .ZN(P3_U3295) );
  OAI222_X1 U12429 ( .A1(n10826), .A2(P3_U3151), .B1(n13851), .B2(n9029), .C1(
        n9955), .C2(n13840), .ZN(P3_U3294) );
  INV_X1 U12430 ( .A(n11194), .ZN(n10731) );
  INV_X1 U12431 ( .A(SI_2_), .ZN(n9956) );
  OAI222_X1 U12432 ( .A1(n10731), .A2(P3_U3151), .B1(n13851), .B2(n9957), .C1(
        n9956), .C2(n13840), .ZN(P3_U3293) );
  INV_X1 U12433 ( .A(SI_5_), .ZN(n9958) );
  OAI222_X1 U12434 ( .A1(n10886), .A2(P3_U3151), .B1(n13851), .B2(n9959), .C1(
        n9958), .C2(n13840), .ZN(P3_U3290) );
  INV_X1 U12435 ( .A(n10768), .ZN(n10857) );
  OAI222_X1 U12436 ( .A1(n10857), .A2(P3_U3151), .B1(n13851), .B2(n9961), .C1(
        n9960), .C2(n13840), .ZN(P3_U3292) );
  OAI222_X1 U12437 ( .A1(n15239), .A2(n9962), .B1(n15238), .B2(n9976), .C1(
        n14734), .C2(P1_U3086), .ZN(P1_U3353) );
  INV_X1 U12438 ( .A(n9965), .ZN(n9966) );
  OAI222_X1 U12439 ( .A1(P3_U3151), .A2(n11331), .B1(n13840), .B2(n9967), .C1(
        n13851), .C2(n9966), .ZN(P3_U3287) );
  OAI222_X1 U12440 ( .A1(P3_U3151), .A2(n11332), .B1(n13840), .B2(n9969), .C1(
        n13851), .C2(n9968), .ZN(P3_U3286) );
  INV_X1 U12441 ( .A(SI_4_), .ZN(n9970) );
  OAI222_X1 U12442 ( .A1(n10801), .A2(P3_U3151), .B1(n13851), .B2(n9971), .C1(
        n9970), .C2(n13840), .ZN(P3_U3291) );
  INV_X1 U12443 ( .A(n9972), .ZN(n9974) );
  OAI222_X1 U12444 ( .A1(P3_U3151), .A2(n10869), .B1(n13851), .B2(n9974), .C1(
        n9973), .C2(n13840), .ZN(P3_U3289) );
  NOR2_X1 U12445 ( .A1(n9975), .A2(P2_STATE_REG_SCAN_IN), .ZN(n14384) );
  INV_X2 U12446 ( .A(n14384), .ZN(n12861) );
  AND2_X1 U12447 ( .A1(n9975), .A2(P2_U3088), .ZN(n14389) );
  INV_X2 U12448 ( .A(n14389), .ZN(n14396) );
  OAI222_X1 U12449 ( .A1(n12861), .A2(n9977), .B1(n14396), .B2(n9976), .C1(
        P2_U3088), .C2(n13990), .ZN(P2_U3325) );
  INV_X1 U12450 ( .A(SI_10_), .ZN(n9979) );
  OAI222_X1 U12451 ( .A1(P3_U3151), .A2(n11914), .B1(n13840), .B2(n9979), .C1(
        n13851), .C2(n9978), .ZN(P3_U3285) );
  OAI222_X1 U12452 ( .A1(n12861), .A2(n9982), .B1(n14396), .B2(n9981), .C1(
        P2_U3088), .C2(n10261), .ZN(P2_U3326) );
  OAI222_X1 U12453 ( .A1(P3_U3151), .A2(n11981), .B1(n13840), .B2(n9984), .C1(
        n13851), .C2(n9983), .ZN(P3_U3284) );
  INV_X1 U12454 ( .A(n10945), .ZN(n9988) );
  INV_X1 U12455 ( .A(n10309), .ZN(n10317) );
  OAI222_X1 U12456 ( .A1(n12861), .A2(n9985), .B1(n14396), .B2(n9988), .C1(
        P2_U3088), .C2(n10317), .ZN(P2_U3323) );
  NAND2_X1 U12457 ( .A1(n9986), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9987) );
  XNOR2_X1 U12458 ( .A(n9987), .B(P1_IR_REG_4__SCAN_IN), .ZN(n15456) );
  INV_X1 U12459 ( .A(n15456), .ZN(n9989) );
  INV_X1 U12460 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n10948) );
  OAI222_X1 U12461 ( .A1(n9989), .A2(P1_U3086), .B1(n15238), .B2(n9988), .C1(
        n10948), .C2(n15239), .ZN(P1_U3351) );
  INV_X1 U12462 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n9994) );
  INV_X1 U12463 ( .A(n11027), .ZN(n9995) );
  NOR2_X1 U12464 ( .A1(n9990), .A2(n15227), .ZN(n9991) );
  MUX2_X1 U12465 ( .A(n15227), .B(n9991), .S(P1_IR_REG_5__SCAN_IN), .Z(n9993)
         );
  AND2_X1 U12466 ( .A1(n9990), .A2(n9992), .ZN(n10005) );
  OR2_X1 U12467 ( .A1(n9993), .A2(n10005), .ZN(n14766) );
  OAI222_X1 U12468 ( .A1(n15239), .A2(n9994), .B1(n15238), .B2(n9995), .C1(
        n14766), .C2(P1_U3086), .ZN(P1_U3350) );
  INV_X1 U12469 ( .A(n10296), .ZN(n10303) );
  OAI222_X1 U12470 ( .A1(n12861), .A2(n9996), .B1(n14396), .B2(n9995), .C1(
        P2_U3088), .C2(n10303), .ZN(P2_U3322) );
  INV_X1 U12471 ( .A(n9997), .ZN(n9998) );
  OAI222_X1 U12472 ( .A1(P3_U3151), .A2(n13377), .B1(n13840), .B2(n9999), .C1(
        n13851), .C2(n9998), .ZN(P3_U3283) );
  NAND2_X1 U12473 ( .A1(n6960), .A2(n13826), .ZN(n10000) );
  OAI21_X1 U12474 ( .B1(n13826), .B2(n9751), .A(n10000), .ZN(P3_U3376) );
  INV_X1 U12475 ( .A(n11232), .ZN(n10009) );
  INV_X1 U12476 ( .A(n15540), .ZN(n10001) );
  OAI222_X1 U12477 ( .A1(n12861), .A2(n10002), .B1(n14396), .B2(n10009), .C1(
        P2_U3088), .C2(n10001), .ZN(P2_U3321) );
  NOR2_X1 U12478 ( .A1(n10005), .A2(n15227), .ZN(n10003) );
  MUX2_X1 U12479 ( .A(n15227), .B(n10003), .S(P1_IR_REG_6__SCAN_IN), .Z(n10007) );
  NAND2_X1 U12480 ( .A1(n10005), .A2(n10004), .ZN(n10243) );
  INV_X1 U12481 ( .A(n10243), .ZN(n10006) );
  OAI222_X1 U12482 ( .A1(n14782), .A2(P1_U3086), .B1(n15238), .B2(n10009), 
        .C1(n10008), .C2(n15239), .ZN(P1_U3349) );
  INV_X1 U12483 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n10010) );
  INV_X1 U12484 ( .A(n11343), .ZN(n10012) );
  INV_X1 U12485 ( .A(n10143), .ZN(n10127) );
  OAI222_X1 U12486 ( .A1(n12861), .A2(n10010), .B1(n14396), .B2(n10012), .C1(
        P2_U3088), .C2(n10127), .ZN(P2_U3320) );
  NAND2_X1 U12487 ( .A1(n10243), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10011) );
  XNOR2_X1 U12488 ( .A(n10011), .B(P1_IR_REG_7__SCAN_IN), .ZN(n11344) );
  INV_X1 U12489 ( .A(n11344), .ZN(n10557) );
  OAI222_X1 U12490 ( .A1(n15239), .A2(n10013), .B1(n15238), .B2(n10012), .C1(
        n10557), .C2(P1_U3086), .ZN(P1_U3348) );
  INV_X1 U12491 ( .A(n11395), .ZN(n10026) );
  OR2_X1 U12492 ( .A1(n10243), .A2(P1_IR_REG_7__SCAN_IN), .ZN(n10014) );
  NAND2_X1 U12493 ( .A1(n10014), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10031) );
  XNOR2_X1 U12494 ( .A(n10031), .B(P1_IR_REG_8__SCAN_IN), .ZN(n11396) );
  INV_X1 U12495 ( .A(n15239), .ZN(n15229) );
  AOI22_X1 U12496 ( .A1(n11396), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(n15229), .ZN(n10015) );
  OAI21_X1 U12497 ( .B1(n10026), .B2(n15238), .A(n10015), .ZN(P1_U3347) );
  OAI222_X1 U12498 ( .A1(n13394), .A2(P3_U3151), .B1(n13851), .B2(n10017), 
        .C1(n10016), .C2(n13840), .ZN(P3_U3282) );
  NAND2_X1 U12499 ( .A1(n10182), .A2(n10018), .ZN(n15478) );
  INV_X1 U12500 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n10021) );
  INV_X1 U12501 ( .A(n10019), .ZN(n10020) );
  AOI22_X1 U12502 ( .A1(n15478), .A2(n10021), .B1(n10024), .B2(n10020), .ZN(
        P1_U3445) );
  INV_X1 U12503 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n10025) );
  INV_X1 U12504 ( .A(n10022), .ZN(n10023) );
  AOI22_X1 U12505 ( .A1(n15478), .A2(n10025), .B1(n10024), .B2(n10023), .ZN(
        P1_U3446) );
  INV_X1 U12506 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n10027) );
  INV_X1 U12507 ( .A(n10218), .ZN(n10153) );
  OAI222_X1 U12508 ( .A1(n12861), .A2(n10027), .B1(n14396), .B2(n10026), .C1(
        P2_U3088), .C2(n10153), .ZN(P2_U3319) );
  OAI222_X1 U12509 ( .A1(P3_U3151), .A2(n13405), .B1(n13840), .B2(n10029), 
        .C1(n13851), .C2(n10028), .ZN(P3_U3281) );
  INV_X1 U12510 ( .A(n11818), .ZN(n10034) );
  NAND2_X1 U12511 ( .A1(n10031), .A2(n10030), .ZN(n10032) );
  NAND2_X1 U12512 ( .A1(n10032), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10070) );
  XNOR2_X1 U12513 ( .A(n10070), .B(P1_IR_REG_9__SCAN_IN), .ZN(n14800) );
  AOI22_X1 U12514 ( .A1(n14800), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_9__SCAN_IN), .B2(n15229), .ZN(n10033) );
  OAI21_X1 U12515 ( .B1(n10034), .B2(n15238), .A(n10033), .ZN(P1_U3346) );
  INV_X1 U12516 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n10035) );
  INV_X1 U12517 ( .A(n10231), .ZN(n10275) );
  OAI222_X1 U12518 ( .A1(n12861), .A2(n10035), .B1(n14396), .B2(n10034), .C1(
        P2_U3088), .C2(n10275), .ZN(P2_U3318) );
  INV_X1 U12519 ( .A(n13826), .ZN(n10036) );
  NOR2_X1 U12520 ( .A1(n10036), .A2(n9752), .ZN(n10038) );
  INV_X1 U12521 ( .A(P3_D_REG_23__SCAN_IN), .ZN(n10037) );
  NOR2_X1 U12522 ( .A1(n10068), .A2(n10037), .ZN(P3_U3242) );
  CLKBUF_X1 U12523 ( .A(n10038), .Z(n10068) );
  INV_X1 U12524 ( .A(P3_D_REG_2__SCAN_IN), .ZN(n10039) );
  NOR2_X1 U12525 ( .A1(n10068), .A2(n10039), .ZN(P3_U3263) );
  INV_X1 U12526 ( .A(P3_D_REG_22__SCAN_IN), .ZN(n10040) );
  NOR2_X1 U12527 ( .A1(n10038), .A2(n10040), .ZN(P3_U3243) );
  INV_X1 U12528 ( .A(P3_D_REG_31__SCAN_IN), .ZN(n10041) );
  NOR2_X1 U12529 ( .A1(n10038), .A2(n10041), .ZN(P3_U3234) );
  INV_X1 U12530 ( .A(P3_D_REG_29__SCAN_IN), .ZN(n10042) );
  NOR2_X1 U12531 ( .A1(n10038), .A2(n10042), .ZN(P3_U3236) );
  INV_X1 U12532 ( .A(P3_D_REG_15__SCAN_IN), .ZN(n10043) );
  NOR2_X1 U12533 ( .A1(n10068), .A2(n10043), .ZN(P3_U3250) );
  INV_X1 U12534 ( .A(P3_D_REG_5__SCAN_IN), .ZN(n10044) );
  NOR2_X1 U12535 ( .A1(n10038), .A2(n10044), .ZN(P3_U3260) );
  INV_X1 U12536 ( .A(P3_D_REG_16__SCAN_IN), .ZN(n10045) );
  NOR2_X1 U12537 ( .A1(n10068), .A2(n10045), .ZN(P3_U3249) );
  INV_X1 U12538 ( .A(P3_D_REG_17__SCAN_IN), .ZN(n10046) );
  NOR2_X1 U12539 ( .A1(n10068), .A2(n10046), .ZN(P3_U3248) );
  INV_X1 U12540 ( .A(P3_D_REG_18__SCAN_IN), .ZN(n10047) );
  NOR2_X1 U12541 ( .A1(n10068), .A2(n10047), .ZN(P3_U3247) );
  INV_X1 U12542 ( .A(P3_D_REG_19__SCAN_IN), .ZN(n10048) );
  NOR2_X1 U12543 ( .A1(n10068), .A2(n10048), .ZN(P3_U3246) );
  INV_X1 U12544 ( .A(P3_D_REG_20__SCAN_IN), .ZN(n10049) );
  NOR2_X1 U12545 ( .A1(n10038), .A2(n10049), .ZN(P3_U3245) );
  INV_X1 U12546 ( .A(P3_D_REG_24__SCAN_IN), .ZN(n10050) );
  NOR2_X1 U12547 ( .A1(n10038), .A2(n10050), .ZN(P3_U3241) );
  INV_X1 U12548 ( .A(P3_D_REG_25__SCAN_IN), .ZN(n10051) );
  NOR2_X1 U12549 ( .A1(n10038), .A2(n10051), .ZN(P3_U3240) );
  INV_X1 U12550 ( .A(P3_D_REG_26__SCAN_IN), .ZN(n10052) );
  NOR2_X1 U12551 ( .A1(n10038), .A2(n10052), .ZN(P3_U3239) );
  INV_X1 U12552 ( .A(P3_D_REG_27__SCAN_IN), .ZN(n10053) );
  NOR2_X1 U12553 ( .A1(n10038), .A2(n10053), .ZN(P3_U3238) );
  INV_X1 U12554 ( .A(P3_D_REG_28__SCAN_IN), .ZN(n10054) );
  NOR2_X1 U12555 ( .A1(n10038), .A2(n10054), .ZN(P3_U3237) );
  INV_X1 U12556 ( .A(P3_D_REG_13__SCAN_IN), .ZN(n10055) );
  NOR2_X1 U12557 ( .A1(n10068), .A2(n10055), .ZN(P3_U3252) );
  INV_X1 U12558 ( .A(P3_D_REG_30__SCAN_IN), .ZN(n10056) );
  NOR2_X1 U12559 ( .A1(n10038), .A2(n10056), .ZN(P3_U3235) );
  INV_X1 U12560 ( .A(P3_D_REG_12__SCAN_IN), .ZN(n10057) );
  NOR2_X1 U12561 ( .A1(n10068), .A2(n10057), .ZN(P3_U3253) );
  INV_X1 U12562 ( .A(P3_D_REG_4__SCAN_IN), .ZN(n10058) );
  NOR2_X1 U12563 ( .A1(n10068), .A2(n10058), .ZN(P3_U3261) );
  INV_X1 U12564 ( .A(P3_D_REG_3__SCAN_IN), .ZN(n10059) );
  NOR2_X1 U12565 ( .A1(n10068), .A2(n10059), .ZN(P3_U3262) );
  INV_X1 U12566 ( .A(P3_D_REG_10__SCAN_IN), .ZN(n10060) );
  NOR2_X1 U12567 ( .A1(n10068), .A2(n10060), .ZN(P3_U3255) );
  INV_X1 U12568 ( .A(P3_D_REG_9__SCAN_IN), .ZN(n10061) );
  NOR2_X1 U12569 ( .A1(n10068), .A2(n10061), .ZN(P3_U3256) );
  INV_X1 U12570 ( .A(P3_D_REG_8__SCAN_IN), .ZN(n10062) );
  NOR2_X1 U12571 ( .A1(n10068), .A2(n10062), .ZN(P3_U3257) );
  INV_X1 U12572 ( .A(P3_D_REG_21__SCAN_IN), .ZN(n10063) );
  NOR2_X1 U12573 ( .A1(n10068), .A2(n10063), .ZN(P3_U3244) );
  INV_X1 U12574 ( .A(P3_D_REG_11__SCAN_IN), .ZN(n10064) );
  NOR2_X1 U12575 ( .A1(n10068), .A2(n10064), .ZN(P3_U3254) );
  INV_X1 U12576 ( .A(P3_D_REG_14__SCAN_IN), .ZN(n10065) );
  NOR2_X1 U12577 ( .A1(n10068), .A2(n10065), .ZN(P3_U3251) );
  INV_X1 U12578 ( .A(P3_D_REG_7__SCAN_IN), .ZN(n10066) );
  NOR2_X1 U12579 ( .A1(n10068), .A2(n10066), .ZN(P3_U3258) );
  INV_X1 U12580 ( .A(P3_D_REG_6__SCAN_IN), .ZN(n10067) );
  NOR2_X1 U12581 ( .A1(n10068), .A2(n10067), .ZN(P3_U3259) );
  INV_X1 U12582 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n10069) );
  INV_X1 U12583 ( .A(n11934), .ZN(n10074) );
  INV_X1 U12584 ( .A(n10279), .ZN(n10349) );
  OAI222_X1 U12585 ( .A1(n12861), .A2(n10069), .B1(n14396), .B2(n10074), .C1(
        P2_U3088), .C2(n10349), .ZN(P2_U3317) );
  NAND2_X1 U12586 ( .A1(n10070), .A2(n10239), .ZN(n10071) );
  NAND2_X1 U12587 ( .A1(n10071), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10072) );
  XNOR2_X1 U12588 ( .A(n10072), .B(P1_IR_REG_10__SCAN_IN), .ZN(n11935) );
  INV_X1 U12589 ( .A(n11935), .ZN(n10474) );
  OAI222_X1 U12590 ( .A1(n10474), .A2(P1_U3086), .B1(n15238), .B2(n10074), 
        .C1(n10073), .C2(n15239), .ZN(P1_U3345) );
  NAND2_X1 U12591 ( .A1(n10075), .A2(n12058), .ZN(n10077) );
  NAND2_X1 U12592 ( .A1(n10077), .A2(n10076), .ZN(n10078) );
  NAND2_X1 U12593 ( .A1(n10079), .A2(n10078), .ZN(n10083) );
  AND2_X1 U12594 ( .A1(n10083), .A2(n8875), .ZN(n15579) );
  AND2_X1 U12595 ( .A1(n15579), .A2(P2_STATE_REG_SCAN_IN), .ZN(n15603) );
  OR2_X1 U12596 ( .A1(n10083), .A2(P2_U3088), .ZN(n15566) );
  INV_X1 U12597 ( .A(n15566), .ZN(n15601) );
  NOR2_X1 U12598 ( .A1(n10080), .A2(P2_STATE_REG_SCAN_IN), .ZN(n10101) );
  NAND2_X1 U12599 ( .A1(n10081), .A2(P2_STATE_REG_SCAN_IN), .ZN(n14390) );
  INV_X1 U12600 ( .A(n14390), .ZN(n10082) );
  NAND2_X1 U12601 ( .A1(n10083), .A2(n10082), .ZN(n10102) );
  INV_X1 U12602 ( .A(n10102), .ZN(n10084) );
  INV_X1 U12603 ( .A(n8938), .ZN(n13167) );
  AND2_X1 U12604 ( .A1(n10084), .A2(n13167), .ZN(n15604) );
  INV_X1 U12605 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n10086) );
  MUX2_X1 U12606 ( .A(n10086), .B(P2_REG2_REG_2__SCAN_IN), .S(n13990), .Z(
        n13996) );
  XNOR2_X1 U12607 ( .A(n10261), .B(P2_REG2_REG_1__SCAN_IN), .ZN(n10258) );
  AND2_X1 U12608 ( .A1(P2_REG2_REG_0__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), 
        .ZN(n10257) );
  NAND2_X1 U12609 ( .A1(n10258), .A2(n10257), .ZN(n10256) );
  INV_X1 U12610 ( .A(n10261), .ZN(n10103) );
  NAND2_X1 U12611 ( .A1(n10103), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n10085) );
  NAND2_X1 U12612 ( .A1(n10256), .A2(n10085), .ZN(n13995) );
  NAND2_X1 U12613 ( .A1(n13996), .A2(n13995), .ZN(n13994) );
  OR2_X1 U12614 ( .A1(n13990), .A2(n10086), .ZN(n10162) );
  NAND2_X1 U12615 ( .A1(n13994), .A2(n10162), .ZN(n10088) );
  INV_X1 U12616 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n11165) );
  MUX2_X1 U12617 ( .A(n11165), .B(P2_REG2_REG_3__SCAN_IN), .S(n10166), .Z(
        n10087) );
  NAND2_X1 U12618 ( .A1(n10088), .A2(n10087), .ZN(n10312) );
  OR2_X1 U12619 ( .A1(n10166), .A2(n11165), .ZN(n10311) );
  NAND2_X1 U12620 ( .A1(n10312), .A2(n10311), .ZN(n10090) );
  INV_X1 U12621 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n11521) );
  MUX2_X1 U12622 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n11521), .S(n10309), .Z(
        n10089) );
  NAND2_X1 U12623 ( .A1(n10090), .A2(n10089), .ZN(n10314) );
  NAND2_X1 U12624 ( .A1(n10309), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n10298) );
  NAND2_X1 U12625 ( .A1(n10314), .A2(n10298), .ZN(n10092) );
  INV_X1 U12626 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n11068) );
  MUX2_X1 U12627 ( .A(P2_REG2_REG_5__SCAN_IN), .B(n11068), .S(n10296), .Z(
        n10091) );
  NAND2_X1 U12628 ( .A1(n10092), .A2(n10091), .ZN(n10300) );
  NAND2_X1 U12629 ( .A1(n10296), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n10093) );
  NAND2_X1 U12630 ( .A1(n10300), .A2(n10093), .ZN(n15546) );
  INV_X1 U12631 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n11110) );
  MUX2_X1 U12632 ( .A(P2_REG2_REG_6__SCAN_IN), .B(n11110), .S(n15540), .Z(
        n15545) );
  NAND2_X1 U12633 ( .A1(n15546), .A2(n15545), .ZN(n15544) );
  NAND2_X1 U12634 ( .A1(n15540), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n10098) );
  NAND2_X1 U12635 ( .A1(n15544), .A2(n10098), .ZN(n10096) );
  INV_X1 U12636 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n10094) );
  MUX2_X1 U12637 ( .A(P2_REG2_REG_7__SCAN_IN), .B(n10094), .S(n10143), .Z(
        n10095) );
  NAND2_X1 U12638 ( .A1(n10096), .A2(n10095), .ZN(n10138) );
  MUX2_X1 U12639 ( .A(n10094), .B(P2_REG2_REG_7__SCAN_IN), .S(n10143), .Z(
        n10097) );
  NAND3_X1 U12640 ( .A1(n15544), .A2(n10098), .A3(n10097), .ZN(n10099) );
  AND3_X1 U12641 ( .A1(n15604), .A2(n10138), .A3(n10099), .ZN(n10100) );
  AOI211_X1 U12642 ( .C1(n15601), .C2(P2_ADDR_REG_7__SCAN_IN), .A(n10101), .B(
        n10100), .ZN(n10126) );
  XNOR2_X1 U12643 ( .A(n13990), .B(P2_REG1_REG_2__SCAN_IN), .ZN(n13991) );
  NAND2_X1 U12644 ( .A1(n10103), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n10106) );
  INV_X1 U12645 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n15683) );
  NAND2_X1 U12646 ( .A1(P2_REG1_REG_0__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), 
        .ZN(n10104) );
  AOI21_X1 U12647 ( .B1(n10261), .B2(n15683), .A(n10104), .ZN(n10105) );
  NAND2_X1 U12648 ( .A1(n10106), .A2(n10105), .ZN(n10253) );
  NAND2_X1 U12649 ( .A1(n10253), .A2(n10106), .ZN(n13992) );
  NAND2_X1 U12650 ( .A1(n13991), .A2(n13992), .ZN(n10109) );
  INV_X1 U12651 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n10107) );
  OR2_X1 U12652 ( .A1(n13990), .A2(n10107), .ZN(n10108) );
  NAND2_X1 U12653 ( .A1(n10109), .A2(n10108), .ZN(n10154) );
  INV_X1 U12654 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n10110) );
  MUX2_X1 U12655 ( .A(n10110), .B(P2_REG1_REG_3__SCAN_IN), .S(n10166), .Z(
        n10111) );
  NAND2_X1 U12656 ( .A1(n10154), .A2(n10111), .ZN(n10155) );
  INV_X1 U12657 ( .A(n10166), .ZN(n10112) );
  NAND2_X1 U12658 ( .A1(n10112), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n10113) );
  NAND2_X1 U12659 ( .A1(n10155), .A2(n10113), .ZN(n10306) );
  INV_X1 U12660 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n10114) );
  MUX2_X1 U12661 ( .A(P2_REG1_REG_4__SCAN_IN), .B(n10114), .S(n10309), .Z(
        n10305) );
  NAND2_X1 U12662 ( .A1(n10306), .A2(n10305), .ZN(n10304) );
  NAND2_X1 U12663 ( .A1(n10309), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n10291) );
  NAND2_X1 U12664 ( .A1(n10304), .A2(n10291), .ZN(n10116) );
  INV_X1 U12665 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n10289) );
  MUX2_X1 U12666 ( .A(P2_REG1_REG_5__SCAN_IN), .B(n10289), .S(n10296), .Z(
        n10115) );
  NAND2_X1 U12667 ( .A1(n10116), .A2(n10115), .ZN(n10293) );
  NAND2_X1 U12668 ( .A1(n10296), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n10117) );
  NAND2_X1 U12669 ( .A1(n10293), .A2(n10117), .ZN(n15543) );
  INV_X1 U12670 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n10118) );
  MUX2_X1 U12671 ( .A(P2_REG1_REG_6__SCAN_IN), .B(n10118), .S(n15540), .Z(
        n15542) );
  NAND2_X1 U12672 ( .A1(n15543), .A2(n15542), .ZN(n15541) );
  NAND2_X1 U12673 ( .A1(n15540), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n10123) );
  NAND2_X1 U12674 ( .A1(n15541), .A2(n10123), .ZN(n10121) );
  INV_X1 U12675 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n10119) );
  MUX2_X1 U12676 ( .A(P2_REG1_REG_7__SCAN_IN), .B(n10119), .S(n10143), .Z(
        n10120) );
  NAND2_X1 U12677 ( .A1(n10121), .A2(n10120), .ZN(n10149) );
  MUX2_X1 U12678 ( .A(n10119), .B(P2_REG1_REG_7__SCAN_IN), .S(n10143), .Z(
        n10122) );
  NAND3_X1 U12679 ( .A1(n15541), .A2(n10123), .A3(n10122), .ZN(n10124) );
  NAND3_X1 U12680 ( .A1(n15609), .A2(n10149), .A3(n10124), .ZN(n10125) );
  OAI211_X1 U12681 ( .C1(n10350), .C2(n10127), .A(n10126), .B(n10125), .ZN(
        P2_U3221) );
  INV_X1 U12682 ( .A(n10128), .ZN(n10129) );
  OAI222_X1 U12683 ( .A1(P3_U3151), .A2(n13427), .B1(n13840), .B2(n10130), 
        .C1(n13851), .C2(n10129), .ZN(P3_U3280) );
  NAND2_X1 U12684 ( .A1(n10131), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n10134) );
  NAND2_X1 U12685 ( .A1(n8941), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n10133) );
  NAND2_X1 U12686 ( .A1(n8942), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n10132) );
  INV_X1 U12687 ( .A(n14023), .ZN(n13098) );
  NAND2_X1 U12688 ( .A1(n6672), .A2(n13098), .ZN(n10135) );
  OAI21_X1 U12689 ( .B1(n6672), .B2(n10136), .A(n10135), .ZN(P2_U3562) );
  NAND2_X1 U12690 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(P2_U3088), .ZN(n11123) );
  NAND2_X1 U12691 ( .A1(n10143), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n10137) );
  NAND2_X1 U12692 ( .A1(n10138), .A2(n10137), .ZN(n10140) );
  INV_X1 U12693 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n11134) );
  MUX2_X1 U12694 ( .A(P2_REG2_REG_8__SCAN_IN), .B(n11134), .S(n10218), .Z(
        n10139) );
  NAND2_X1 U12695 ( .A1(n10140), .A2(n10139), .ZN(n10217) );
  OAI211_X1 U12696 ( .C1(n10140), .C2(n10139), .A(n15604), .B(n10217), .ZN(
        n10141) );
  NAND2_X1 U12697 ( .A1(n11123), .A2(n10141), .ZN(n10142) );
  AOI21_X1 U12698 ( .B1(n15601), .B2(P2_ADDR_REG_8__SCAN_IN), .A(n10142), .ZN(
        n10152) );
  NAND2_X1 U12699 ( .A1(n10143), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n10148) );
  NAND2_X1 U12700 ( .A1(n10149), .A2(n10148), .ZN(n10145) );
  MUX2_X1 U12701 ( .A(P2_REG1_REG_8__SCAN_IN), .B(n10146), .S(n10218), .Z(
        n10144) );
  NAND2_X1 U12702 ( .A1(n10145), .A2(n10144), .ZN(n10220) );
  INV_X1 U12703 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n10146) );
  MUX2_X1 U12704 ( .A(n10146), .B(P2_REG1_REG_8__SCAN_IN), .S(n10218), .Z(
        n10147) );
  NAND3_X1 U12705 ( .A1(n10149), .A2(n10148), .A3(n10147), .ZN(n10150) );
  NAND3_X1 U12706 ( .A1(n15609), .A2(n10220), .A3(n10150), .ZN(n10151) );
  OAI211_X1 U12707 ( .C1(n10350), .C2(n10153), .A(n10152), .B(n10151), .ZN(
        P2_U3222) );
  NAND2_X1 U12708 ( .A1(P2_U3088), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n10385) );
  INV_X1 U12709 ( .A(n10385), .ZN(n10160) );
  INV_X1 U12710 ( .A(n10154), .ZN(n10158) );
  MUX2_X1 U12711 ( .A(P2_REG1_REG_3__SCAN_IN), .B(n10110), .S(n10166), .Z(
        n10157) );
  INV_X1 U12712 ( .A(n10155), .ZN(n10156) );
  AOI211_X1 U12713 ( .C1(n10158), .C2(n10157), .A(n10156), .B(n14009), .ZN(
        n10159) );
  AOI211_X1 U12714 ( .C1(n15601), .C2(P2_ADDR_REG_3__SCAN_IN), .A(n10160), .B(
        n10159), .ZN(n10165) );
  MUX2_X1 U12715 ( .A(P2_REG2_REG_3__SCAN_IN), .B(n11165), .S(n10166), .Z(
        n10161) );
  NAND3_X1 U12716 ( .A1(n13994), .A2(n10162), .A3(n10161), .ZN(n10163) );
  NAND3_X1 U12717 ( .A1(n15604), .A2(n10312), .A3(n10163), .ZN(n10164) );
  OAI211_X1 U12718 ( .C1(n10350), .C2(n10166), .A(n10165), .B(n10164), .ZN(
        P2_U3217) );
  INV_X1 U12719 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n10167) );
  MUX2_X1 U12720 ( .A(n10167), .B(P1_REG1_REG_8__SCAN_IN), .S(n11396), .Z(
        n10180) );
  INV_X1 U12721 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n15532) );
  INV_X1 U12722 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n11652) );
  INV_X1 U12723 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n10168) );
  MUX2_X1 U12724 ( .A(n10168), .B(P1_REG1_REG_2__SCAN_IN), .S(n14734), .Z(
        n10173) );
  INV_X1 U12725 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n10169) );
  MUX2_X1 U12726 ( .A(n10169), .B(P1_REG1_REG_1__SCAN_IN), .S(n14710), .Z(
        n10171) );
  AND2_X1 U12727 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), 
        .ZN(n10170) );
  NAND2_X1 U12728 ( .A1(n10171), .A2(n10170), .ZN(n14731) );
  OR2_X1 U12729 ( .A1(n14710), .A2(n10169), .ZN(n14730) );
  NAND2_X1 U12730 ( .A1(n14731), .A2(n14730), .ZN(n10172) );
  NAND2_X1 U12731 ( .A1(n10173), .A2(n10172), .ZN(n14748) );
  INV_X1 U12732 ( .A(n14734), .ZN(n14729) );
  NAND2_X1 U12733 ( .A1(n14729), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n14746) );
  NAND2_X1 U12734 ( .A1(n14748), .A2(n14746), .ZN(n10175) );
  INV_X1 U12735 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n10176) );
  MUX2_X1 U12736 ( .A(n10176), .B(P1_REG1_REG_3__SCAN_IN), .S(n14750), .Z(
        n10174) );
  NAND2_X1 U12737 ( .A1(n10175), .A2(n10174), .ZN(n15446) );
  OR2_X1 U12738 ( .A1(n14750), .A2(n10176), .ZN(n15445) );
  INV_X1 U12739 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n10971) );
  MUX2_X1 U12740 ( .A(n10971), .B(P1_REG1_REG_4__SCAN_IN), .S(n15456), .Z(
        n15444) );
  AOI21_X1 U12741 ( .B1(n15446), .B2(n15445), .A(n15444), .ZN(n15448) );
  AND2_X1 U12742 ( .A1(n15456), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n10177) );
  NOR2_X1 U12743 ( .A1(n15448), .A2(n10177), .ZN(n14763) );
  INV_X1 U12744 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n15530) );
  MUX2_X1 U12745 ( .A(n15530), .B(P1_REG1_REG_5__SCAN_IN), .S(n14766), .Z(
        n14764) );
  NAND2_X1 U12746 ( .A1(n14763), .A2(n14764), .ZN(n14762) );
  NAND2_X1 U12747 ( .A1(n14766), .A2(n15530), .ZN(n10178) );
  NAND2_X1 U12748 ( .A1(n14762), .A2(n10178), .ZN(n14779) );
  MUX2_X1 U12749 ( .A(P1_REG1_REG_6__SCAN_IN), .B(n11652), .S(n14782), .Z(
        n14778) );
  OR2_X1 U12750 ( .A1(n14779), .A2(n14778), .ZN(n14781) );
  OAI21_X1 U12751 ( .B1(n11652), .B2(n14782), .A(n14781), .ZN(n10548) );
  MUX2_X1 U12752 ( .A(P1_REG1_REG_7__SCAN_IN), .B(n15532), .S(n11344), .Z(
        n10547) );
  NAND2_X1 U12753 ( .A1(n10548), .A2(n10547), .ZN(n10546) );
  OAI21_X1 U12754 ( .B1(n15532), .B2(n10557), .A(n10546), .ZN(n10179) );
  NOR2_X1 U12755 ( .A1(n10179), .A2(n10180), .ZN(n14797) );
  AOI21_X1 U12756 ( .B1(n10180), .B2(n10179), .A(n14797), .ZN(n10215) );
  INV_X1 U12757 ( .A(n12844), .ZN(n10181) );
  OR2_X1 U12758 ( .A1(n10182), .A2(n10181), .ZN(n10189) );
  NAND2_X1 U12759 ( .A1(n10184), .A2(n10183), .ZN(n10185) );
  NAND2_X1 U12760 ( .A1(n10185), .A2(n12448), .ZN(n10188) );
  INV_X1 U12761 ( .A(n10188), .ZN(n10186) );
  INV_X1 U12762 ( .A(n10193), .ZN(n10396) );
  NAND2_X1 U12763 ( .A1(n10396), .A2(n14718), .ZN(n15468) );
  NOR2_X2 U12764 ( .A1(n10193), .A2(n14721), .ZN(n15457) );
  NAND2_X1 U12765 ( .A1(n10189), .A2(n10188), .ZN(n15476) );
  NAND2_X1 U12766 ( .A1(P1_REG3_REG_8__SCAN_IN), .A2(P1_U3086), .ZN(n11772) );
  OAI21_X1 U12767 ( .B1(n15476), .B2(n10190), .A(n11772), .ZN(n10191) );
  AOI21_X1 U12768 ( .B1(n15457), .B2(n11396), .A(n10191), .ZN(n10214) );
  INV_X1 U12769 ( .A(n14718), .ZN(n12581) );
  NAND2_X1 U12770 ( .A1(n14721), .A2(n12581), .ZN(n10192) );
  NOR2_X2 U12771 ( .A1(n10193), .A2(n10192), .ZN(n14838) );
  INV_X1 U12772 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n10194) );
  MUX2_X1 U12773 ( .A(n10194), .B(P1_REG2_REG_5__SCAN_IN), .S(n14766), .Z(
        n10201) );
  INV_X1 U12774 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n14735) );
  MUX2_X1 U12775 ( .A(n14735), .B(P1_REG2_REG_2__SCAN_IN), .S(n14734), .Z(
        n10197) );
  INV_X1 U12776 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n10195) );
  MUX2_X1 U12777 ( .A(n10195), .B(P1_REG2_REG_1__SCAN_IN), .S(n14710), .Z(
        n14714) );
  AND2_X1 U12778 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n14720) );
  NAND2_X1 U12779 ( .A1(n14714), .A2(n14720), .ZN(n14737) );
  OR2_X1 U12780 ( .A1(n14710), .A2(n10195), .ZN(n14736) );
  NAND2_X1 U12781 ( .A1(n14737), .A2(n14736), .ZN(n10196) );
  NAND2_X1 U12782 ( .A1(n10197), .A2(n10196), .ZN(n14753) );
  NAND2_X1 U12783 ( .A1(n14729), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n14751) );
  NAND2_X1 U12784 ( .A1(n14753), .A2(n14751), .ZN(n10199) );
  INV_X1 U12785 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n11533) );
  MUX2_X1 U12786 ( .A(n11533), .B(P1_REG2_REG_3__SCAN_IN), .S(n14750), .Z(
        n10198) );
  NAND2_X1 U12787 ( .A1(n10199), .A2(n10198), .ZN(n15451) );
  OR2_X1 U12788 ( .A1(n14750), .A2(n11533), .ZN(n15450) );
  INV_X1 U12789 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n11206) );
  MUX2_X1 U12790 ( .A(n11206), .B(P1_REG2_REG_4__SCAN_IN), .S(n15456), .Z(
        n15449) );
  AOI21_X1 U12791 ( .B1(n15451), .B2(n15450), .A(n15449), .ZN(n15453) );
  AND2_X1 U12792 ( .A1(n15456), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n14767) );
  OR2_X1 U12793 ( .A1(n15453), .A2(n14767), .ZN(n10200) );
  NAND2_X1 U12794 ( .A1(n10201), .A2(n10200), .ZN(n14784) );
  INV_X1 U12795 ( .A(n14766), .ZN(n14761) );
  NAND2_X1 U12796 ( .A1(n14761), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n14783) );
  NAND2_X1 U12797 ( .A1(n14784), .A2(n14783), .ZN(n10203) );
  INV_X1 U12798 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n11588) );
  MUX2_X1 U12799 ( .A(n11588), .B(P1_REG2_REG_6__SCAN_IN), .S(n14782), .Z(
        n10202) );
  NAND2_X1 U12800 ( .A1(n10203), .A2(n10202), .ZN(n14787) );
  INV_X1 U12801 ( .A(n14782), .ZN(n14777) );
  NAND2_X1 U12802 ( .A1(n14777), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n10552) );
  NAND2_X1 U12803 ( .A1(n14787), .A2(n10552), .ZN(n10206) );
  INV_X1 U12804 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n10204) );
  MUX2_X1 U12805 ( .A(P1_REG2_REG_7__SCAN_IN), .B(n10204), .S(n11344), .Z(
        n10205) );
  NAND2_X1 U12806 ( .A1(n10206), .A2(n10205), .ZN(n10554) );
  NAND2_X1 U12807 ( .A1(n11344), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n10211) );
  NAND2_X1 U12808 ( .A1(n10554), .A2(n10211), .ZN(n10209) );
  INV_X1 U12809 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n10207) );
  MUX2_X1 U12810 ( .A(P1_REG2_REG_8__SCAN_IN), .B(n10207), .S(n11396), .Z(
        n10208) );
  NAND2_X1 U12811 ( .A1(n10209), .A2(n10208), .ZN(n14803) );
  MUX2_X1 U12812 ( .A(n10207), .B(P1_REG2_REG_8__SCAN_IN), .S(n11396), .Z(
        n10210) );
  NAND3_X1 U12813 ( .A1(n10554), .A2(n10211), .A3(n10210), .ZN(n10212) );
  NAND3_X1 U12814 ( .A1(n14838), .A2(n14803), .A3(n10212), .ZN(n10213) );
  OAI211_X1 U12815 ( .C1(n10215), .C2(n15468), .A(n10214), .B(n10213), .ZN(
        P1_U3251) );
  INV_X1 U12816 ( .A(n15604), .ZN(n11888) );
  INV_X1 U12817 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n10262) );
  NOR2_X1 U12818 ( .A1(n11888), .A2(n10262), .ZN(n10223) );
  NAND2_X1 U12819 ( .A1(n10218), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n10216) );
  NAND2_X1 U12820 ( .A1(n10217), .A2(n10216), .ZN(n10230) );
  INV_X1 U12821 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n10274) );
  NAND2_X1 U12822 ( .A1(n10218), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n10219) );
  NAND2_X1 U12823 ( .A1(n10220), .A2(n10219), .ZN(n10225) );
  INV_X1 U12824 ( .A(n10225), .ZN(n10221) );
  NOR3_X1 U12825 ( .A1(n14009), .A2(n10274), .A3(n10221), .ZN(n10222) );
  AOI211_X1 U12826 ( .C1(n10223), .C2(n10230), .A(n15603), .B(n10222), .ZN(
        n10237) );
  NOR2_X1 U12827 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n11268), .ZN(n10228) );
  MUX2_X1 U12828 ( .A(n10274), .B(P2_REG1_REG_9__SCAN_IN), .S(n10231), .Z(
        n10224) );
  OR2_X1 U12829 ( .A1(n10225), .A2(n10224), .ZN(n10277) );
  NAND3_X1 U12830 ( .A1(n10225), .A2(n10274), .A3(n10275), .ZN(n10226) );
  AOI21_X1 U12831 ( .B1(n10277), .B2(n10226), .A(n14009), .ZN(n10227) );
  AOI211_X1 U12832 ( .C1(n15601), .C2(P2_ADDR_REG_9__SCAN_IN), .A(n10228), .B(
        n10227), .ZN(n10236) );
  MUX2_X1 U12833 ( .A(n10262), .B(P2_REG2_REG_9__SCAN_IN), .S(n10231), .Z(
        n10229) );
  OR2_X1 U12834 ( .A1(n10230), .A2(n10229), .ZN(n10264) );
  INV_X1 U12835 ( .A(n10264), .ZN(n10234) );
  INV_X1 U12836 ( .A(n10230), .ZN(n10232) );
  NOR3_X1 U12837 ( .A1(n10232), .A2(P2_REG2_REG_9__SCAN_IN), .A3(n10231), .ZN(
        n10233) );
  OAI21_X1 U12838 ( .B1(n10234), .B2(n10233), .A(n15604), .ZN(n10235) );
  OAI211_X1 U12839 ( .C1(n10237), .C2(n10275), .A(n10236), .B(n10235), .ZN(
        P2_U3223) );
  INV_X1 U12840 ( .A(n12155), .ZN(n10247) );
  INV_X1 U12841 ( .A(n11679), .ZN(n10271) );
  OAI222_X1 U12842 ( .A1(n12861), .A2(n10238), .B1(n14396), .B2(n10247), .C1(
        P2_U3088), .C2(n10271), .ZN(P2_U3316) );
  NAND3_X1 U12843 ( .A1(n10241), .A2(n10240), .A3(n10239), .ZN(n10242) );
  NAND2_X1 U12844 ( .A1(n10358), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10245) );
  XNOR2_X1 U12845 ( .A(n10245), .B(n10244), .ZN(n10432) );
  OAI222_X1 U12846 ( .A1(n10432), .A2(P1_U3086), .B1(n15238), .B2(n10247), 
        .C1(n10246), .C2(n15239), .ZN(P1_U3344) );
  INV_X1 U12847 ( .A(n10248), .ZN(n10249) );
  OAI222_X1 U12848 ( .A1(n13840), .A2(n10250), .B1(n13851), .B2(n10249), .C1(
        n13452), .C2(P3_U3151), .ZN(P3_U3279) );
  INV_X1 U12849 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n11658) );
  NOR2_X1 U12850 ( .A1(n11658), .A2(P2_STATE_REG_SCAN_IN), .ZN(n10255) );
  INV_X1 U12851 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n15681) );
  MUX2_X1 U12852 ( .A(P2_REG1_REG_1__SCAN_IN), .B(n15683), .S(n10261), .Z(
        n10251) );
  OAI21_X1 U12853 ( .B1(n15681), .B2(n10331), .A(n10251), .ZN(n10252) );
  AND3_X1 U12854 ( .A1(n15609), .A2(n10253), .A3(n10252), .ZN(n10254) );
  AOI211_X1 U12855 ( .C1(n15601), .C2(P2_ADDR_REG_1__SCAN_IN), .A(n10255), .B(
        n10254), .ZN(n10260) );
  OAI211_X1 U12856 ( .C1(n10258), .C2(n10257), .A(n15604), .B(n10256), .ZN(
        n10259) );
  OAI211_X1 U12857 ( .C1(n10350), .C2(n10261), .A(n10260), .B(n10259), .ZN(
        P2_U3215) );
  NAND2_X1 U12858 ( .A1(n10275), .A2(n10262), .ZN(n10263) );
  NAND2_X1 U12859 ( .A1(n10264), .A2(n10263), .ZN(n10336) );
  INV_X1 U12860 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n10265) );
  MUX2_X1 U12861 ( .A(n10265), .B(P2_REG2_REG_10__SCAN_IN), .S(n10279), .Z(
        n10337) );
  OR2_X1 U12862 ( .A1(n10336), .A2(n10337), .ZN(n10338) );
  NAND2_X1 U12863 ( .A1(n10279), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n10266) );
  NAND2_X1 U12864 ( .A1(n10338), .A2(n10266), .ZN(n10270) );
  INV_X1 U12865 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n10267) );
  MUX2_X1 U12866 ( .A(n10267), .B(P2_REG2_REG_11__SCAN_IN), .S(n11679), .Z(
        n10269) );
  OR2_X1 U12867 ( .A1(n10270), .A2(n10269), .ZN(n15559) );
  INV_X1 U12868 ( .A(n15559), .ZN(n10268) );
  AOI21_X1 U12869 ( .B1(n10270), .B2(n10269), .A(n10268), .ZN(n10288) );
  NAND2_X1 U12870 ( .A1(P2_REG3_REG_11__SCAN_IN), .A2(P2_U3088), .ZN(n15351)
         );
  INV_X1 U12871 ( .A(n15351), .ZN(n10273) );
  NOR2_X1 U12872 ( .A1(n10350), .A2(n10271), .ZN(n10272) );
  AOI211_X1 U12873 ( .C1(n15601), .C2(P2_ADDR_REG_11__SCAN_IN), .A(n10273), 
        .B(n10272), .ZN(n10287) );
  NAND2_X1 U12874 ( .A1(n10275), .A2(n10274), .ZN(n10276) );
  NAND2_X1 U12875 ( .A1(n10277), .A2(n10276), .ZN(n10340) );
  INV_X1 U12876 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n10278) );
  MUX2_X1 U12877 ( .A(n10278), .B(P2_REG1_REG_10__SCAN_IN), .S(n10279), .Z(
        n10341) );
  OR2_X1 U12878 ( .A1(n10340), .A2(n10341), .ZN(n10342) );
  NAND2_X1 U12879 ( .A1(n10279), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n10284) );
  NAND2_X1 U12880 ( .A1(n10342), .A2(n10284), .ZN(n10282) );
  INV_X1 U12881 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n10280) );
  MUX2_X1 U12882 ( .A(P2_REG1_REG_11__SCAN_IN), .B(n10280), .S(n11679), .Z(
        n10281) );
  NAND2_X1 U12883 ( .A1(n10282), .A2(n10281), .ZN(n11681) );
  MUX2_X1 U12884 ( .A(n10280), .B(P2_REG1_REG_11__SCAN_IN), .S(n11679), .Z(
        n10283) );
  NAND3_X1 U12885 ( .A1(n10342), .A2(n10284), .A3(n10283), .ZN(n10285) );
  NAND3_X1 U12886 ( .A1(n15609), .A2(n11681), .A3(n10285), .ZN(n10286) );
  OAI211_X1 U12887 ( .C1(n10288), .C2(n11888), .A(n10287), .B(n10286), .ZN(
        P2_U3225) );
  MUX2_X1 U12888 ( .A(n10289), .B(P2_REG1_REG_5__SCAN_IN), .S(n10296), .Z(
        n10290) );
  NAND3_X1 U12889 ( .A1(n10304), .A2(n10291), .A3(n10290), .ZN(n10292) );
  NAND3_X1 U12890 ( .A1(n15609), .A2(n10293), .A3(n10292), .ZN(n10294) );
  NAND2_X1 U12891 ( .A1(P2_REG3_REG_5__SCAN_IN), .A2(P2_U3088), .ZN(n10539) );
  OAI211_X1 U12892 ( .C1(n15789), .C2(n15566), .A(n10294), .B(n10539), .ZN(
        n10295) );
  INV_X1 U12893 ( .A(n10295), .ZN(n10302) );
  MUX2_X1 U12894 ( .A(n11068), .B(P2_REG2_REG_5__SCAN_IN), .S(n10296), .Z(
        n10297) );
  NAND3_X1 U12895 ( .A1(n10314), .A2(n10298), .A3(n10297), .ZN(n10299) );
  NAND3_X1 U12896 ( .A1(n15604), .A2(n10300), .A3(n10299), .ZN(n10301) );
  OAI211_X1 U12897 ( .C1(n10350), .C2(n10303), .A(n10302), .B(n10301), .ZN(
        P2_U3219) );
  NAND2_X1 U12898 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_U3088), .ZN(n10448) );
  OAI211_X1 U12899 ( .C1(n10306), .C2(n10305), .A(n15609), .B(n10304), .ZN(
        n10307) );
  NAND2_X1 U12900 ( .A1(n10448), .A2(n10307), .ZN(n10308) );
  AOI21_X1 U12901 ( .B1(n15601), .B2(P2_ADDR_REG_4__SCAN_IN), .A(n10308), .ZN(
        n10316) );
  MUX2_X1 U12902 ( .A(n11521), .B(P2_REG2_REG_4__SCAN_IN), .S(n10309), .Z(
        n10310) );
  NAND3_X1 U12903 ( .A1(n10312), .A2(n10311), .A3(n10310), .ZN(n10313) );
  NAND3_X1 U12904 ( .A1(n15604), .A2(n10314), .A3(n10313), .ZN(n10315) );
  OAI211_X1 U12905 ( .C1(n10350), .C2(n10317), .A(n10316), .B(n10315), .ZN(
        P2_U3218) );
  NAND2_X1 U12906 ( .A1(n12519), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n10322) );
  NAND2_X1 U12907 ( .A1(n6680), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n10321) );
  NAND2_X1 U12908 ( .A1(n11039), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n11244) );
  NOR2_X1 U12909 ( .A1(n11244), .A2(n11243), .ZN(n11356) );
  NAND2_X1 U12910 ( .A1(n11356), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n11402) );
  INV_X1 U12911 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n11401) );
  INV_X1 U12912 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n11826) );
  INV_X1 U12913 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n11946) );
  OR2_X1 U12914 ( .A1(n11948), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n10318) );
  NAND2_X1 U12915 ( .A1(n11948), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n12289) );
  AND2_X1 U12916 ( .A1(n10318), .A2(n12289), .ZN(n12318) );
  NAND2_X1 U12917 ( .A1(n6677), .A2(n12318), .ZN(n10320) );
  NAND2_X1 U12918 ( .A1(n6683), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n10319) );
  MUX2_X1 U12919 ( .A(n10352), .B(n15385), .S(P1_U4016), .Z(n10323) );
  INV_X1 U12920 ( .A(n10323), .ZN(P1_U3572) );
  NAND2_X1 U12921 ( .A1(n13326), .A2(n10860), .ZN(n10324) );
  OAI21_X1 U12922 ( .B1(n10860), .B2(n10325), .A(n10324), .ZN(P3_U3508) );
  NAND2_X1 U12923 ( .A1(n13706), .A2(n10860), .ZN(n10326) );
  OAI21_X1 U12924 ( .B1(n10860), .B2(n10327), .A(n10326), .ZN(P3_U3505) );
  INV_X1 U12925 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n10328) );
  NAND2_X1 U12926 ( .A1(n15604), .A2(n10328), .ZN(n10329) );
  OAI211_X1 U12927 ( .C1(P2_REG1_REG_0__SCAN_IN), .C2(n14009), .A(n10350), .B(
        n10329), .ZN(n10330) );
  INV_X1 U12928 ( .A(n10330), .ZN(n10333) );
  AOI22_X1 U12929 ( .A1(P2_REG1_REG_0__SCAN_IN), .A2(n15609), .B1(n15604), 
        .B2(P2_REG2_REG_0__SCAN_IN), .ZN(n10332) );
  MUX2_X1 U12930 ( .A(n10333), .B(n10332), .S(n10331), .Z(n10335) );
  AOI22_X1 U12931 ( .A1(n15601), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3088), .ZN(n10334) );
  NAND2_X1 U12932 ( .A1(n10335), .A2(n10334), .ZN(P2_U3214) );
  AOI21_X1 U12933 ( .B1(n10337), .B2(n10336), .A(n11888), .ZN(n10339) );
  NAND2_X1 U12934 ( .A1(n10339), .A2(n10338), .ZN(n10345) );
  AOI21_X1 U12935 ( .B1(n10341), .B2(n10340), .A(n14009), .ZN(n10343) );
  NAND2_X1 U12936 ( .A1(n10343), .A2(n10342), .ZN(n10344) );
  NAND2_X1 U12937 ( .A1(n10345), .A2(n10344), .ZN(n10347) );
  NAND2_X1 U12938 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(P2_U3088), .ZN(n11311)
         );
  INV_X1 U12939 ( .A(n11311), .ZN(n10346) );
  AOI211_X1 U12940 ( .C1(n15601), .C2(P2_ADDR_REG_10__SCAN_IN), .A(n10347), 
        .B(n10346), .ZN(n10348) );
  OAI21_X1 U12941 ( .B1(n10350), .B2(n10349), .A(n10348), .ZN(P2_U3224) );
  NAND2_X1 U12942 ( .A1(n13358), .A2(P3_DATAO_REG_21__SCAN_IN), .ZN(n10351) );
  OAI21_X1 U12943 ( .B1(n13638), .B2(n13358), .A(n10351), .ZN(P3_U3512) );
  INV_X1 U12944 ( .A(n12275), .ZN(n10361) );
  INV_X1 U12945 ( .A(n15555), .ZN(n11684) );
  OAI222_X1 U12946 ( .A1(n14396), .A2(n10361), .B1(n11684), .B2(P2_U3088), 
        .C1(n10352), .C2(n12861), .ZN(P2_U3315) );
  NAND2_X1 U12947 ( .A1(n13988), .A2(n12105), .ZN(n15618) );
  OR2_X1 U12948 ( .A1(n10353), .A2(P2_U3088), .ZN(n10411) );
  AOI22_X1 U12949 ( .A1(n15350), .A2(n12863), .B1(n10411), .B2(
        P2_REG3_REG_0__SCAN_IN), .ZN(n10357) );
  NAND2_X1 U12950 ( .A1(n13989), .A2(n15616), .ZN(n13119) );
  NOR2_X1 U12951 ( .A1(n13119), .A2(n14206), .ZN(n10355) );
  OAI21_X1 U12952 ( .B1(n10355), .B2(n10354), .A(n15345), .ZN(n10356) );
  OAI211_X1 U12953 ( .C1(n15618), .C2(n13953), .A(n10357), .B(n10356), .ZN(
        P2_U3204) );
  NAND2_X1 U12954 ( .A1(n10359), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10454) );
  XNOR2_X1 U12955 ( .A(n10454), .B(P1_IR_REG_12__SCAN_IN), .ZN(n12276) );
  INV_X1 U12956 ( .A(n12276), .ZN(n10365) );
  OAI222_X1 U12957 ( .A1(P1_U3086), .A2(n10365), .B1(n15238), .B2(n10361), 
        .C1(n10360), .C2(n15239), .ZN(P1_U3343) );
  INV_X1 U12958 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n15415) );
  NOR2_X1 U12959 ( .A1(n11396), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n14795) );
  INV_X1 U12960 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n15535) );
  MUX2_X1 U12961 ( .A(P1_REG1_REG_9__SCAN_IN), .B(n15535), .S(n14800), .Z(
        n14796) );
  OAI21_X1 U12962 ( .B1(n14797), .B2(n14795), .A(n14796), .ZN(n14794) );
  OAI21_X1 U12963 ( .B1(n14800), .B2(P1_REG1_REG_9__SCAN_IN), .A(n14794), .ZN(
        n10461) );
  INV_X1 U12964 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n12086) );
  MUX2_X1 U12965 ( .A(n12086), .B(P1_REG1_REG_10__SCAN_IN), .S(n11935), .Z(
        n10462) );
  NOR2_X1 U12966 ( .A1(n10461), .A2(n10462), .ZN(n10460) );
  AOI21_X1 U12967 ( .B1(n11935), .B2(P1_REG1_REG_10__SCAN_IN), .A(n10460), 
        .ZN(n10427) );
  MUX2_X1 U12968 ( .A(n15415), .B(P1_REG1_REG_11__SCAN_IN), .S(n10432), .Z(
        n10362) );
  AND2_X1 U12969 ( .A1(n10427), .A2(n10362), .ZN(n10428) );
  AOI21_X1 U12970 ( .B1(n15415), .B2(n10432), .A(n10428), .ZN(n10364) );
  INV_X1 U12971 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n15275) );
  AOI22_X1 U12972 ( .A1(n12276), .A2(n15275), .B1(P1_REG1_REG_12__SCAN_IN), 
        .B2(n10365), .ZN(n10363) );
  NOR2_X1 U12973 ( .A1(n10364), .A2(n10363), .ZN(n10487) );
  AOI21_X1 U12974 ( .B1(n10364), .B2(n10363), .A(n10487), .ZN(n10383) );
  INV_X1 U12975 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n10366) );
  AOI22_X1 U12976 ( .A1(n12276), .A2(n10366), .B1(P1_REG2_REG_12__SCAN_IN), 
        .B2(n10365), .ZN(n10376) );
  INV_X1 U12977 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n10420) );
  NAND2_X1 U12978 ( .A1(n11396), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n14802) );
  NAND2_X1 U12979 ( .A1(n14803), .A2(n14802), .ZN(n10369) );
  INV_X1 U12980 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n10367) );
  MUX2_X1 U12981 ( .A(P1_REG2_REG_9__SCAN_IN), .B(n10367), .S(n14800), .Z(
        n10368) );
  NAND2_X1 U12982 ( .A1(n10369), .A2(n10368), .ZN(n14805) );
  NAND2_X1 U12983 ( .A1(n14800), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n10467) );
  NAND2_X1 U12984 ( .A1(n14805), .A2(n10467), .ZN(n10372) );
  INV_X1 U12985 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n10370) );
  MUX2_X1 U12986 ( .A(P1_REG2_REG_10__SCAN_IN), .B(n10370), .S(n11935), .Z(
        n10371) );
  NAND2_X1 U12987 ( .A1(n10372), .A2(n10371), .ZN(n10469) );
  NAND2_X1 U12988 ( .A1(n11935), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n10373) );
  NAND2_X1 U12989 ( .A1(n10469), .A2(n10373), .ZN(n10422) );
  MUX2_X1 U12990 ( .A(n10420), .B(P1_REG2_REG_11__SCAN_IN), .S(n10432), .Z(
        n10374) );
  NAND2_X1 U12991 ( .A1(n10422), .A2(n10374), .ZN(n10421) );
  OAI21_X1 U12992 ( .B1(n10432), .B2(n10420), .A(n10421), .ZN(n10375) );
  NOR2_X1 U12993 ( .A1(n10376), .A2(n10375), .ZN(n10491) );
  AOI21_X1 U12994 ( .B1(n10376), .B2(n10375), .A(n10491), .ZN(n10380) );
  INV_X1 U12995 ( .A(n14838), .ZN(n15470) );
  INV_X1 U12996 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n12315) );
  NOR2_X1 U12997 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n12315), .ZN(n10377) );
  AOI21_X1 U12998 ( .B1(n14819), .B2(P1_ADDR_REG_12__SCAN_IN), .A(n10377), 
        .ZN(n10379) );
  NAND2_X1 U12999 ( .A1(n15457), .A2(n12276), .ZN(n10378) );
  OAI211_X1 U13000 ( .C1(n10380), .C2(n15470), .A(n10379), .B(n10378), .ZN(
        n10381) );
  INV_X1 U13001 ( .A(n10381), .ZN(n10382) );
  OAI21_X1 U13002 ( .B1(n10383), .B2(n15468), .A(n10382), .ZN(P1_U3255) );
  OAI22_X1 U13003 ( .A1(n6962), .A2(n13913), .B1(n10538), .B2(n13915), .ZN(
        n11163) );
  INV_X1 U13004 ( .A(n11163), .ZN(n10387) );
  NAND2_X1 U13005 ( .A1(n13944), .A2(n8383), .ZN(n10386) );
  OAI211_X1 U13006 ( .C1(n10387), .C2(n13953), .A(n10386), .B(n10385), .ZN(
        n10388) );
  AOI21_X1 U13007 ( .B1(n15652), .B2(n15350), .A(n10388), .ZN(n10389) );
  OAI21_X1 U13008 ( .B1(n10390), .B2(n13935), .A(n10389), .ZN(P2_U3190) );
  INV_X1 U13009 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n10399) );
  NAND3_X1 U13010 ( .A1(n14833), .A2(P1_IR_REG_0__SCAN_IN), .A3(n9873), .ZN(
        n10398) );
  INV_X1 U13011 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n10391) );
  NAND2_X1 U13012 ( .A1(n12581), .A2(n10391), .ZN(n10392) );
  AND2_X1 U13013 ( .A1(n14721), .A2(n10392), .ZN(n14725) );
  INV_X1 U13014 ( .A(n14725), .ZN(n10394) );
  AOI21_X1 U13015 ( .B1(n9873), .B2(n14718), .A(n10394), .ZN(n10393) );
  MUX2_X1 U13016 ( .A(n10394), .B(n10393), .S(n14712), .Z(n10395) );
  AOI22_X1 U13017 ( .A1(n10396), .A2(n10395), .B1(P1_REG3_REG_0__SCAN_IN), 
        .B2(P1_U3086), .ZN(n10397) );
  OAI211_X1 U13018 ( .C1(n15476), .C2(n10399), .A(n10398), .B(n10397), .ZN(
        P1_U3243) );
  INV_X1 U13019 ( .A(n13953), .ZN(n15347) );
  OR2_X1 U13020 ( .A1(n12866), .A2(n13913), .ZN(n10401) );
  NAND2_X1 U13021 ( .A1(n13987), .A2(n12105), .ZN(n10400) );
  AND2_X1 U13022 ( .A1(n10401), .A2(n10400), .ZN(n11656) );
  INV_X1 U13023 ( .A(n11656), .ZN(n10402) );
  AOI22_X1 U13024 ( .A1(n15347), .A2(n10402), .B1(P2_REG3_REG_1__SCAN_IN), 
        .B2(n10411), .ZN(n10408) );
  OAI21_X1 U13025 ( .B1(n10405), .B2(n10404), .A(n10403), .ZN(n10406) );
  NAND2_X1 U13026 ( .A1(n15345), .A2(n10406), .ZN(n10407) );
  OAI211_X1 U13027 ( .C1(n8887), .C2(n13958), .A(n10408), .B(n10407), .ZN(
        P2_U3194) );
  NAND2_X1 U13028 ( .A1(n13988), .A2(n13951), .ZN(n10410) );
  NAND2_X1 U13029 ( .A1(n13986), .A2(n13952), .ZN(n10409) );
  NAND2_X1 U13030 ( .A1(n10410), .A2(n10409), .ZN(n10480) );
  AOI22_X1 U13031 ( .A1(n15347), .A2(n10480), .B1(P2_REG3_REG_2__SCAN_IN), 
        .B2(n10411), .ZN(n10417) );
  OAI21_X1 U13032 ( .B1(n10414), .B2(n10413), .A(n10412), .ZN(n10415) );
  NAND2_X1 U13033 ( .A1(n15345), .A2(n10415), .ZN(n10416) );
  OAI211_X1 U13034 ( .C1(n11501), .C2(n13958), .A(n10417), .B(n10416), .ZN(
        P2_U3209) );
  NOR3_X1 U13035 ( .A1(n10427), .A2(n15415), .A3(n15468), .ZN(n10419) );
  NOR3_X1 U13036 ( .A1(n15470), .A2(P1_REG2_REG_11__SCAN_IN), .A3(n10422), 
        .ZN(n10418) );
  NOR3_X1 U13037 ( .A1(n10419), .A2(n15457), .A3(n10418), .ZN(n10433) );
  INV_X1 U13038 ( .A(n10432), .ZN(n12156) );
  NOR2_X1 U13039 ( .A1(n12156), .A2(n10420), .ZN(n10423) );
  OAI211_X1 U13040 ( .C1(n10423), .C2(n10422), .A(n14838), .B(n10421), .ZN(
        n10424) );
  NAND2_X1 U13041 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_U3086), .ZN(n15399)
         );
  OAI211_X1 U13042 ( .C1(n10425), .C2(n15476), .A(n10424), .B(n15399), .ZN(
        n10426) );
  INV_X1 U13043 ( .A(n10426), .ZN(n10431) );
  NOR3_X1 U13044 ( .A1(n10427), .A2(P1_REG1_REG_11__SCAN_IN), .A3(n12156), 
        .ZN(n10429) );
  OAI21_X1 U13045 ( .B1(n10429), .B2(n10428), .A(n14833), .ZN(n10430) );
  OAI211_X1 U13046 ( .C1(n10433), .C2(n10432), .A(n10431), .B(n10430), .ZN(
        P1_U3254) );
  INV_X1 U13047 ( .A(n12326), .ZN(n10459) );
  INV_X1 U13048 ( .A(n15568), .ZN(n11685) );
  OAI222_X1 U13049 ( .A1(n14396), .A2(n10459), .B1(n11685), .B2(P2_U3088), 
        .C1(n7107), .C2(n12861), .ZN(P2_U3314) );
  INV_X1 U13050 ( .A(n10434), .ZN(n10435) );
  OAI222_X1 U13051 ( .A1(P3_U3151), .A2(n13494), .B1(n13840), .B2(n10436), 
        .C1(n13851), .C2(n10435), .ZN(P3_U3278) );
  XNOR2_X1 U13052 ( .A(n10438), .B(n6922), .ZN(n14719) );
  NOR2_X1 U13053 ( .A1(n10439), .A2(n12840), .ZN(n10664) );
  INV_X1 U13054 ( .A(n10664), .ZN(n10441) );
  OAI22_X1 U13055 ( .A1(n14683), .A2(n12591), .B1(n15092), .B2(n15384), .ZN(
        n10440) );
  AOI21_X1 U13056 ( .B1(n10441), .B2(P1_REG3_REG_0__SCAN_IN), .A(n10440), .ZN(
        n10442) );
  OAI21_X1 U13057 ( .B1(n15392), .B2(n14719), .A(n10442), .ZN(P1_U3232) );
  NAND2_X1 U13058 ( .A1(n10445), .A2(n15345), .ZN(n10452) );
  NAND2_X1 U13059 ( .A1(n13986), .A2(n13951), .ZN(n10447) );
  NAND2_X1 U13060 ( .A1(n13984), .A2(n12105), .ZN(n10446) );
  NAND2_X1 U13061 ( .A1(n10447), .A2(n10446), .ZN(n11519) );
  INV_X1 U13062 ( .A(n11519), .ZN(n10449) );
  OAI21_X1 U13063 ( .B1(n13953), .B2(n10449), .A(n10448), .ZN(n10450) );
  AOI21_X1 U13064 ( .B1(n11512), .B2(n13944), .A(n10450), .ZN(n10451) );
  OAI211_X1 U13065 ( .C1(n11510), .C2(n13958), .A(n10452), .B(n10451), .ZN(
        P2_U3202) );
  NAND2_X1 U13066 ( .A1(n10454), .A2(n10453), .ZN(n10455) );
  NAND2_X1 U13067 ( .A1(n10455), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10457) );
  NAND2_X1 U13068 ( .A1(n10457), .A2(n10456), .ZN(n10608) );
  OAI21_X1 U13069 ( .B1(n10457), .B2(n10456), .A(n10608), .ZN(n12327) );
  OAI222_X1 U13070 ( .A1(P1_U3086), .A2(n12327), .B1(n15238), .B2(n10459), 
        .C1(n10458), .C2(n15239), .ZN(P1_U3342) );
  AND2_X1 U13071 ( .A1(P1_U3086), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n12235) );
  AOI211_X1 U13072 ( .C1(n10462), .C2(n10461), .A(n15468), .B(n10460), .ZN(
        n10463) );
  INV_X1 U13073 ( .A(n10463), .ZN(n10464) );
  OAI21_X1 U13074 ( .B1(n10465), .B2(n15476), .A(n10464), .ZN(n10466) );
  NOR2_X1 U13075 ( .A1(n12235), .A2(n10466), .ZN(n10473) );
  INV_X1 U13076 ( .A(n14805), .ZN(n10471) );
  MUX2_X1 U13077 ( .A(n10370), .B(P1_REG2_REG_10__SCAN_IN), .S(n11935), .Z(
        n10468) );
  NAND2_X1 U13078 ( .A1(n10468), .A2(n10467), .ZN(n10470) );
  OAI211_X1 U13079 ( .C1(n10471), .C2(n10470), .A(n14838), .B(n10469), .ZN(
        n10472) );
  OAI211_X1 U13080 ( .C1(n15472), .C2(n10474), .A(n10473), .B(n10472), .ZN(
        P1_U3253) );
  INV_X1 U13081 ( .A(n8992), .ZN(n15663) );
  XNOR2_X1 U13082 ( .A(n10476), .B(n10475), .ZN(n11499) );
  INV_X1 U13083 ( .A(n11499), .ZN(n10483) );
  INV_X1 U13084 ( .A(n11157), .ZN(n10477) );
  AOI211_X1 U13085 ( .C1(n12882), .C2(n11653), .A(n6670), .B(n10477), .ZN(
        n11504) );
  AOI21_X1 U13086 ( .B1(n15672), .B2(n12882), .A(n11504), .ZN(n10482) );
  OAI21_X1 U13087 ( .B1(n6961), .B2(n10479), .A(n10478), .ZN(n10481) );
  AOI21_X1 U13088 ( .B1(n10481), .B2(n15617), .A(n10480), .ZN(n11507) );
  OAI211_X1 U13089 ( .C1(n10483), .C2(n15675), .A(n10482), .B(n11507), .ZN(
        n10484) );
  AOI21_X1 U13090 ( .B1(n15663), .B2(n11499), .A(n10484), .ZN(n15650) );
  NAND2_X1 U13091 ( .A1(n7435), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n10485) );
  OAI21_X1 U13092 ( .B1(n15650), .B2(n7435), .A(n10485), .ZN(P2_U3501) );
  NOR2_X1 U13093 ( .A1(n12276), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n10486) );
  NOR2_X1 U13094 ( .A1(n10487), .A2(n10486), .ZN(n10489) );
  MUX2_X1 U13095 ( .A(n15407), .B(P1_REG1_REG_13__SCAN_IN), .S(n12327), .Z(
        n10488) );
  NAND2_X1 U13096 ( .A1(n10489), .A2(n10488), .ZN(n10610) );
  OAI211_X1 U13097 ( .C1(n10489), .C2(n10488), .A(n14833), .B(n10610), .ZN(
        n10498) );
  NAND2_X1 U13098 ( .A1(P1_REG3_REG_13__SCAN_IN), .A2(P1_U3086), .ZN(n14640)
         );
  NOR2_X1 U13099 ( .A1(n12276), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n10490) );
  NOR2_X1 U13100 ( .A1(n10491), .A2(n10490), .ZN(n10494) );
  INV_X1 U13101 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n10492) );
  MUX2_X1 U13102 ( .A(n10492), .B(P1_REG2_REG_13__SCAN_IN), .S(n12327), .Z(
        n10493) );
  NAND2_X1 U13103 ( .A1(n10493), .A2(n10494), .ZN(n10615) );
  OAI211_X1 U13104 ( .C1(n10494), .C2(n10493), .A(n10615), .B(n14838), .ZN(
        n10495) );
  NAND2_X1 U13105 ( .A1(n14640), .A2(n10495), .ZN(n10496) );
  AOI21_X1 U13106 ( .B1(n14819), .B2(P1_ADDR_REG_13__SCAN_IN), .A(n10496), 
        .ZN(n10497) );
  OAI211_X1 U13107 ( .C1(n15472), .C2(n12327), .A(n10498), .B(n10497), .ZN(
        P1_U3256) );
  INV_X1 U13108 ( .A(n10508), .ZN(n10504) );
  INV_X1 U13109 ( .A(n10509), .ZN(n10499) );
  OR2_X1 U13110 ( .A1(n10602), .A2(n10499), .ZN(n10503) );
  AND3_X1 U13111 ( .A1(n10501), .A2(n10500), .A3(n10745), .ZN(n10502) );
  OAI211_X1 U13112 ( .C1(n10513), .C2(n10504), .A(n10503), .B(n10502), .ZN(
        n10505) );
  NAND2_X1 U13113 ( .A1(n10505), .A2(P3_STATE_REG_SCAN_IN), .ZN(n10507) );
  OR2_X1 U13114 ( .A1(n10602), .A2(n10601), .ZN(n10506) );
  NAND2_X2 U13115 ( .A1(n10507), .A2(n10506), .ZN(n13350) );
  NOR2_X1 U13116 ( .A1(n13350), .A2(P3_U3151), .ZN(n10683) );
  INV_X1 U13117 ( .A(P3_REG3_REG_0__SCAN_IN), .ZN(n15702) );
  INV_X1 U13118 ( .A(n10584), .ZN(n10518) );
  NAND3_X1 U13119 ( .A1(n10513), .A2(n10508), .A3(n15758), .ZN(n10511) );
  NAND2_X1 U13120 ( .A1(n10602), .A2(n10509), .ZN(n10510) );
  NAND2_X1 U13121 ( .A1(n10511), .A2(n10510), .ZN(n10512) );
  INV_X1 U13122 ( .A(n13352), .ZN(n13322) );
  OR2_X1 U13123 ( .A1(n10513), .A2(n15715), .ZN(n10515) );
  AND2_X1 U13124 ( .A1(n10934), .A2(n15765), .ZN(n10514) );
  INV_X1 U13125 ( .A(n10601), .ZN(n10516) );
  NAND3_X1 U13126 ( .A1(n10516), .A2(n10602), .A3(n10600), .ZN(n13346) );
  OAI22_X1 U13127 ( .A1(n13347), .A2(n10939), .B1(n6957), .B2(n13346), .ZN(
        n10517) );
  AOI21_X1 U13128 ( .B1(n10518), .B2(n13322), .A(n10517), .ZN(n10519) );
  OAI21_X1 U13129 ( .B1(n10683), .B2(n15702), .A(n10519), .ZN(P3_U3172) );
  INV_X1 U13130 ( .A(n10520), .ZN(n10521) );
  OAI222_X1 U13131 ( .A1(P3_U3151), .A2(n13513), .B1(n13840), .B2(n10522), 
        .C1(n13851), .C2(n10521), .ZN(P3_U3277) );
  INV_X1 U13132 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n12288) );
  INV_X1 U13133 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n12336) );
  NAND2_X1 U13134 ( .A1(n12362), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n12403) );
  INV_X1 U13135 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n12402) );
  INV_X1 U13136 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n10523) );
  AND2_X1 U13137 ( .A1(n12405), .A2(n10523), .ZN(n10524) );
  OR2_X1 U13138 ( .A1(n10524), .A2(n12418), .ZN(n15009) );
  NAND2_X1 U13139 ( .A1(n6683), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n10525) );
  OAI21_X1 U13140 ( .B1(n15009), .B2(n12451), .A(n10525), .ZN(n10529) );
  NAND2_X1 U13141 ( .A1(n6680), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n10527) );
  NAND2_X1 U13142 ( .A1(n12519), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n10526) );
  NAND2_X1 U13143 ( .A1(n10527), .A2(n10526), .ZN(n10528) );
  INV_X1 U13144 ( .A(P1_U4016), .ZN(n12391) );
  INV_X1 U13145 ( .A(n12391), .ZN(n14723) );
  MUX2_X1 U13146 ( .A(n11256), .B(n15022), .S(n14723), .Z(n10530) );
  INV_X1 U13147 ( .A(n10530), .ZN(P1_U3578) );
  MUX2_X1 U13148 ( .A(n10531), .B(n10954), .S(n14723), .Z(n10532) );
  INV_X1 U13149 ( .A(n10532), .ZN(P1_U3563) );
  INV_X1 U13150 ( .A(n12907), .ZN(n11073) );
  OAI21_X1 U13151 ( .B1(n10535), .B2(n10534), .A(n10533), .ZN(n10536) );
  NAND2_X1 U13152 ( .A1(n10536), .A2(n15345), .ZN(n10543) );
  OAI22_X1 U13153 ( .A1(n10538), .A2(n13913), .B1(n10537), .B2(n13915), .ZN(
        n10914) );
  INV_X1 U13154 ( .A(n10914), .ZN(n10540) );
  OAI21_X1 U13155 ( .B1(n13953), .B2(n10540), .A(n10539), .ZN(n10541) );
  AOI21_X1 U13156 ( .B1(n11071), .B2(n13944), .A(n10541), .ZN(n10542) );
  OAI211_X1 U13157 ( .C1(n11073), .C2(n13958), .A(n10543), .B(n10542), .ZN(
        P2_U3199) );
  OAI222_X1 U13158 ( .A1(n13851), .A2(n10545), .B1(n13840), .B2(n10544), .C1(
        P3_U3151), .C2(n9671), .ZN(P3_U3276) );
  NAND2_X1 U13159 ( .A1(P1_REG3_REG_7__SCAN_IN), .A2(P1_U3086), .ZN(n11362) );
  OAI211_X1 U13160 ( .C1(n10548), .C2(n10547), .A(n14833), .B(n10546), .ZN(
        n10549) );
  NAND2_X1 U13161 ( .A1(n11362), .A2(n10549), .ZN(n10550) );
  AOI21_X1 U13162 ( .B1(n14819), .B2(P1_ADDR_REG_7__SCAN_IN), .A(n10550), .ZN(
        n10556) );
  MUX2_X1 U13163 ( .A(n10204), .B(P1_REG2_REG_7__SCAN_IN), .S(n11344), .Z(
        n10551) );
  NAND3_X1 U13164 ( .A1(n14787), .A2(n10552), .A3(n10551), .ZN(n10553) );
  NAND3_X1 U13165 ( .A1(n14838), .A2(n10554), .A3(n10553), .ZN(n10555) );
  OAI211_X1 U13166 ( .C1(n15472), .C2(n10557), .A(n10556), .B(n10555), .ZN(
        P1_U3250) );
  INV_X1 U13167 ( .A(n13693), .ZN(n13227) );
  NAND2_X1 U13168 ( .A1(n13227), .A2(n10860), .ZN(n10558) );
  OAI21_X1 U13169 ( .B1(P3_U3897), .B2(n10559), .A(n10558), .ZN(P3_U3506) );
  NAND2_X1 U13170 ( .A1(n7656), .A2(n10860), .ZN(n10560) );
  OAI21_X1 U13171 ( .B1(P3_U3897), .B2(n10561), .A(n10560), .ZN(P3_U3509) );
  NAND2_X1 U13172 ( .A1(n13707), .A2(n10860), .ZN(n10562) );
  OAI21_X1 U13173 ( .B1(P3_U3897), .B2(n10563), .A(n10562), .ZN(P3_U3507) );
  NAND2_X1 U13174 ( .A1(n13308), .A2(n10860), .ZN(n10564) );
  OAI21_X1 U13175 ( .B1(P3_U3897), .B2(n10565), .A(n10564), .ZN(P3_U3510) );
  XNOR2_X1 U13176 ( .A(n10567), .B(n10566), .ZN(n10575) );
  INV_X1 U13177 ( .A(n10568), .ZN(n11114) );
  NOR2_X1 U13178 ( .A1(n15354), .A2(n11114), .ZN(n10573) );
  NAND2_X1 U13179 ( .A1(n13984), .A2(n13951), .ZN(n10570) );
  NAND2_X1 U13180 ( .A1(n13982), .A2(n12105), .ZN(n10569) );
  NAND2_X1 U13181 ( .A1(n10570), .A2(n10569), .ZN(n11108) );
  INV_X1 U13182 ( .A(n11108), .ZN(n10571) );
  NAND2_X1 U13183 ( .A1(P2_U3088), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n15538) );
  OAI21_X1 U13184 ( .B1(n13953), .B2(n10571), .A(n15538), .ZN(n10572) );
  AOI211_X1 U13185 ( .C1(n15671), .C2(n15350), .A(n10573), .B(n10572), .ZN(
        n10574) );
  OAI21_X1 U13186 ( .B1(n10575), .B2(n13935), .A(n10574), .ZN(P2_U3211) );
  INV_X1 U13187 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n14708) );
  OAI21_X1 U13188 ( .B1(n10578), .B2(n10577), .A(n10576), .ZN(n10579) );
  NAND2_X1 U13189 ( .A1(n10579), .A2(n14675), .ZN(n10582) );
  INV_X1 U13190 ( .A(n14707), .ZN(n15073) );
  OAI22_X1 U13191 ( .A1(n15387), .A2(n15073), .B1(n10688), .B2(n15384), .ZN(
        n10580) );
  AOI21_X1 U13192 ( .B1(n15085), .B2(n15397), .A(n10580), .ZN(n10581) );
  OAI211_X1 U13193 ( .C1(n10664), .C2(n14708), .A(n10582), .B(n10581), .ZN(
        P1_U3222) );
  OR3_X1 U13194 ( .A1(n10584), .A2(n15765), .A3(n10583), .ZN(n10587) );
  INV_X1 U13195 ( .A(n13696), .ZN(n15719) );
  NAND2_X1 U13196 ( .A1(n10585), .A2(n15719), .ZN(n10586) );
  NAND2_X1 U13197 ( .A1(n10587), .A2(n10586), .ZN(n10935) );
  INV_X1 U13198 ( .A(P3_REG0_REG_0__SCAN_IN), .ZN(n10588) );
  OAI22_X1 U13199 ( .A1(n10939), .A2(n13825), .B1(n15775), .B2(n10588), .ZN(
        n10589) );
  AOI21_X1 U13200 ( .B1(n10935), .B2(n15775), .A(n10589), .ZN(n10590) );
  INV_X1 U13201 ( .A(n10590), .ZN(P3_U3390) );
  INV_X1 U13202 ( .A(P3_REG3_REG_1__SCAN_IN), .ZN(n15728) );
  NAND2_X1 U13203 ( .A1(n10999), .A2(n10926), .ZN(n10593) );
  INV_X1 U13204 ( .A(n6935), .ZN(n10597) );
  NAND3_X1 U13205 ( .A1(n10597), .A2(n15721), .A3(n13254), .ZN(n10598) );
  OAI211_X1 U13206 ( .C1(n6842), .C2(n15720), .A(n10675), .B(n10598), .ZN(
        n10599) );
  NAND2_X1 U13207 ( .A1(n10599), .A2(n13322), .ZN(n10607) );
  NOR2_X1 U13208 ( .A1(n10601), .A2(n10600), .ZN(n10603) );
  NAND2_X1 U13209 ( .A1(n10603), .A2(n10602), .ZN(n13315) );
  OAI22_X1 U13210 ( .A1(n10836), .A2(n13346), .B1(n10604), .B2(n13315), .ZN(
        n10605) );
  AOI21_X1 U13211 ( .B1(n13337), .B2(n9041), .A(n10605), .ZN(n10606) );
  OAI211_X1 U13212 ( .C1(n10683), .C2(n15728), .A(n10607), .B(n10606), .ZN(
        P3_U3162) );
  NAND2_X1 U13213 ( .A1(n10608), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10609) );
  XNOR2_X1 U13214 ( .A(n10609), .B(P1_IR_REG_14__SCAN_IN), .ZN(n12333) );
  INV_X1 U13215 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n11728) );
  INV_X1 U13216 ( .A(n12333), .ZN(n11729) );
  AOI22_X1 U13217 ( .A1(n12333), .A2(n11728), .B1(P1_REG1_REG_14__SCAN_IN), 
        .B2(n11729), .ZN(n10612) );
  INV_X1 U13218 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n15407) );
  OAI21_X1 U13219 ( .B1(n15407), .B2(n12327), .A(n10610), .ZN(n10611) );
  NOR2_X1 U13220 ( .A1(n10612), .A2(n10611), .ZN(n11727) );
  AOI21_X1 U13221 ( .B1(n10612), .B2(n10611), .A(n11727), .ZN(n10621) );
  NAND2_X1 U13222 ( .A1(P1_REG3_REG_14__SCAN_IN), .A2(P1_U3086), .ZN(n15381)
         );
  OAI21_X1 U13223 ( .B1(n15476), .B2(n10613), .A(n15381), .ZN(n10614) );
  AOI21_X1 U13224 ( .B1(n15457), .B2(n12333), .A(n10614), .ZN(n10620) );
  OAI21_X1 U13225 ( .B1(n12327), .B2(n10492), .A(n10615), .ZN(n10618) );
  INV_X1 U13226 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n10616) );
  MUX2_X1 U13227 ( .A(P1_REG2_REG_14__SCAN_IN), .B(n10616), .S(n12333), .Z(
        n10617) );
  NAND2_X1 U13228 ( .A1(n10617), .A2(n10618), .ZN(n11720) );
  OAI211_X1 U13229 ( .C1(n10618), .C2(n10617), .A(n14838), .B(n11720), .ZN(
        n10619) );
  OAI211_X1 U13230 ( .C1(n10621), .C2(n15468), .A(n10620), .B(n10619), .ZN(
        P1_U3257) );
  INV_X1 U13231 ( .A(n12332), .ZN(n10651) );
  INV_X1 U13232 ( .A(n11669), .ZN(n15580) );
  INV_X1 U13233 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n10622) );
  OAI222_X1 U13234 ( .A1(n14396), .A2(n10651), .B1(n15580), .B2(P2_U3088), 
        .C1(n10622), .C2(n12861), .ZN(P2_U3313) );
  NAND2_X1 U13235 ( .A1(n11014), .A2(P3_U3897), .ZN(n10623) );
  OAI21_X1 U13236 ( .B1(n10860), .B2(n10624), .A(n10623), .ZN(P3_U3496) );
  NAND2_X1 U13237 ( .A1(n10625), .A2(P3_U3897), .ZN(n10626) );
  OAI21_X1 U13238 ( .B1(P3_U3897), .B2(n10627), .A(n10626), .ZN(P3_U3494) );
  NAND2_X1 U13239 ( .A1(n11425), .A2(P3_U3897), .ZN(n10628) );
  OAI21_X1 U13240 ( .B1(P3_U3897), .B2(n10629), .A(n10628), .ZN(P3_U3495) );
  NAND2_X1 U13241 ( .A1(n11751), .A2(P3_U3897), .ZN(n10630) );
  OAI21_X1 U13242 ( .B1(n10860), .B2(n10631), .A(n10630), .ZN(P3_U3497) );
  NAND2_X1 U13243 ( .A1(n9512), .A2(P3_U3897), .ZN(n10632) );
  OAI21_X1 U13244 ( .B1(n10860), .B2(n10633), .A(n10632), .ZN(P3_U3491) );
  NAND2_X1 U13245 ( .A1(n12145), .A2(P3_U3897), .ZN(n10634) );
  OAI21_X1 U13246 ( .B1(P3_U3897), .B2(n10635), .A(n10634), .ZN(P3_U3501) );
  NAND2_X1 U13247 ( .A1(n13652), .A2(P3_U3897), .ZN(n10636) );
  OAI21_X1 U13248 ( .B1(n10860), .B2(n10637), .A(n10636), .ZN(P3_U3511) );
  NAND2_X1 U13249 ( .A1(n12223), .A2(P3_U3897), .ZN(n10638) );
  OAI21_X1 U13250 ( .B1(P3_U3897), .B2(n10639), .A(n10638), .ZN(P3_U3502) );
  NAND2_X1 U13251 ( .A1(n12017), .A2(P3_U3897), .ZN(n10640) );
  OAI21_X1 U13252 ( .B1(n10860), .B2(n10641), .A(n10640), .ZN(P3_U3498) );
  NAND2_X1 U13253 ( .A1(n12018), .A2(P3_U3897), .ZN(n10642) );
  OAI21_X1 U13254 ( .B1(P3_U3897), .B2(n10643), .A(n10642), .ZN(P3_U3500) );
  INV_X1 U13255 ( .A(n13630), .ZN(n10644) );
  NAND2_X1 U13256 ( .A1(n10644), .A2(P3_U3897), .ZN(n10645) );
  OAI21_X1 U13257 ( .B1(P3_U3897), .B2(n10646), .A(n10645), .ZN(P3_U3513) );
  NAND2_X1 U13258 ( .A1(n13298), .A2(P3_U3897), .ZN(n10647) );
  OAI21_X1 U13259 ( .B1(P3_U3897), .B2(n10648), .A(n10647), .ZN(P3_U3514) );
  NAND2_X1 U13260 ( .A1(n10717), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10649) );
  XNOR2_X1 U13261 ( .A(n10649), .B(P1_IR_REG_16__SCAN_IN), .ZN(n12395) );
  INV_X1 U13262 ( .A(n12395), .ZN(n11738) );
  INV_X1 U13263 ( .A(n12394), .ZN(n10655) );
  OAI222_X1 U13264 ( .A1(P1_U3086), .A2(n11738), .B1(n15238), .B2(n10655), 
        .C1(n6925), .C2(n15239), .ZN(P1_U3339) );
  OAI222_X1 U13265 ( .A1(P1_U3086), .A2(n11729), .B1(n15238), .B2(n10651), 
        .C1(n10650), .C2(n15239), .ZN(P1_U3341) );
  INV_X1 U13266 ( .A(n12399), .ZN(n10672) );
  OAI222_X1 U13267 ( .A1(n14396), .A2(n10672), .B1(n11884), .B2(P2_U3088), 
        .C1(n10652), .C2(n12861), .ZN(P2_U3310) );
  OAI22_X1 U13268 ( .A1(n13777), .A2(n10939), .B1(n15784), .B2(n15689), .ZN(
        n10653) );
  AOI21_X1 U13269 ( .B1(n10935), .B2(n15784), .A(n10653), .ZN(n10654) );
  INV_X1 U13270 ( .A(n10654), .ZN(P3_U3459) );
  OAI222_X1 U13271 ( .A1(n12861), .A2(n10656), .B1(n11690), .B2(P2_U3088), 
        .C1(n14396), .C2(n10655), .ZN(P2_U3311) );
  INV_X1 U13272 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n14726) );
  OAI21_X1 U13273 ( .B1(n10659), .B2(n10658), .A(n10657), .ZN(n10660) );
  NAND2_X1 U13274 ( .A1(n10660), .A2(n14675), .ZN(n10663) );
  OAI22_X1 U13275 ( .A1(n15387), .A2(n15092), .B1(n10954), .B2(n15384), .ZN(
        n10661) );
  AOI21_X1 U13276 ( .B1(n6669), .B2(n15397), .A(n10661), .ZN(n10662) );
  OAI211_X1 U13277 ( .C1(n10664), .C2(n14726), .A(n10663), .B(n10662), .ZN(
        P1_U3237) );
  NAND2_X1 U13278 ( .A1(n13603), .A2(P3_U3897), .ZN(n10665) );
  OAI21_X1 U13279 ( .B1(P3_U3897), .B2(n10666), .A(n10665), .ZN(P3_U3515) );
  NAND2_X1 U13280 ( .A1(n10667), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10668) );
  MUX2_X1 U13281 ( .A(P1_IR_REG_31__SCAN_IN), .B(n10668), .S(
        P1_IR_REG_17__SCAN_IN), .Z(n10669) );
  INV_X1 U13282 ( .A(n10669), .ZN(n10670) );
  NOR2_X1 U13283 ( .A1(n10670), .A2(n11257), .ZN(n14811) );
  INV_X1 U13284 ( .A(n14811), .ZN(n11931) );
  OAI222_X1 U13285 ( .A1(P1_U3086), .A2(n11931), .B1(n15238), .B2(n10672), 
        .C1(n10671), .C2(n15239), .ZN(P1_U3338) );
  INV_X1 U13286 ( .A(n12345), .ZN(n10720) );
  INV_X1 U13287 ( .A(n15592), .ZN(n11688) );
  INV_X1 U13288 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n10673) );
  OAI222_X1 U13289 ( .A1(n14396), .A2(n10720), .B1(n11688), .B2(P2_U3088), 
        .C1(n10673), .C2(n12861), .ZN(P2_U3312) );
  INV_X1 U13290 ( .A(P3_REG3_REG_2__SCAN_IN), .ZN(n10682) );
  XNOR2_X1 U13291 ( .A(n10829), .B(n10674), .ZN(n10827) );
  XNOR2_X1 U13292 ( .A(n10836), .B(n10827), .ZN(n10677) );
  OAI21_X1 U13293 ( .B1(n10677), .B2(n10676), .A(n10832), .ZN(n10678) );
  NAND2_X1 U13294 ( .A1(n10678), .A2(n13322), .ZN(n10681) );
  OAI22_X1 U13295 ( .A1(n6957), .A2(n13315), .B1(n11224), .B2(n13346), .ZN(
        n10679) );
  AOI21_X1 U13296 ( .B1(n11051), .B2(n13337), .A(n10679), .ZN(n10680) );
  OAI211_X1 U13297 ( .C1(n10683), .C2(n10682), .A(n10681), .B(n10680), .ZN(
        P3_U3177) );
  NAND2_X1 U13298 ( .A1(n11199), .A2(n10684), .ZN(n10685) );
  OR2_X1 U13299 ( .A1(n11200), .A2(n10685), .ZN(n10712) );
  INV_X1 U13300 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n10710) );
  INV_X1 U13301 ( .A(n12591), .ZN(n15485) );
  NAND2_X1 U13302 ( .A1(n14707), .A2(n15485), .ZN(n15077) );
  NAND2_X1 U13303 ( .A1(n15092), .A2(n10686), .ZN(n10687) );
  NAND2_X1 U13304 ( .A1(n15079), .A2(n10687), .ZN(n10691) );
  NAND2_X1 U13305 ( .A1(n10688), .A2(n6669), .ZN(n10951) );
  NAND2_X1 U13306 ( .A1(n10689), .A2(n11544), .ZN(n10690) );
  NAND2_X1 U13307 ( .A1(n10951), .A2(n10690), .ZN(n12797) );
  NAND2_X1 U13308 ( .A1(n10691), .A2(n12797), .ZN(n10942) );
  OR2_X1 U13309 ( .A1(n10691), .A2(n12797), .ZN(n10692) );
  NAND2_X1 U13310 ( .A1(n10942), .A2(n10692), .ZN(n10702) );
  INV_X1 U13311 ( .A(n10702), .ZN(n11549) );
  INV_X1 U13312 ( .A(n15244), .ZN(n10693) );
  NAND2_X1 U13313 ( .A1(n10693), .A2(n12770), .ZN(n12783) );
  OR2_X1 U13314 ( .A1(n14707), .A2(n12591), .ZN(n12795) );
  NAND2_X1 U13315 ( .A1(n12597), .A2(n12795), .ZN(n10694) );
  AND2_X1 U13316 ( .A1(n10694), .A2(n12602), .ZN(n10695) );
  OAI21_X1 U13317 ( .B1(n10696), .B2(n10695), .A(n10952), .ZN(n10700) );
  NAND2_X1 U13318 ( .A1(n15048), .A2(n15244), .ZN(n10698) );
  NAND2_X1 U13319 ( .A1(n12594), .A2(n12787), .ZN(n10697) );
  OAI22_X1 U13320 ( .A1(n10954), .A2(n15091), .B1(n15092), .B2(n15069), .ZN(
        n10699) );
  AOI21_X1 U13321 ( .B1(n10700), .B2(n15280), .A(n10699), .ZN(n10704) );
  NAND2_X1 U13322 ( .A1(n12592), .A2(n15244), .ZN(n10701) );
  NAND2_X1 U13323 ( .A1(n14445), .A2(n10701), .ZN(n11210) );
  NAND2_X1 U13324 ( .A1(n10702), .A2(n15080), .ZN(n10703) );
  NAND2_X1 U13325 ( .A1(n10704), .A2(n10703), .ZN(n11542) );
  INV_X1 U13326 ( .A(n11542), .ZN(n10708) );
  NAND2_X1 U13327 ( .A1(n10686), .A2(n12591), .ZN(n15072) );
  NOR2_X1 U13328 ( .A1(n15072), .A2(n6669), .ZN(n11534) );
  NAND2_X1 U13329 ( .A1(n15072), .A2(n6669), .ZN(n10705) );
  NAND2_X1 U13330 ( .A1(n10705), .A2(n15291), .ZN(n10706) );
  NOR2_X1 U13331 ( .A1(n11534), .A2(n10706), .ZN(n11546) );
  AOI21_X1 U13332 ( .B1(n6669), .B2(n15495), .A(n11546), .ZN(n10707) );
  OAI211_X1 U13333 ( .C1(n11549), .C2(n15499), .A(n10708), .B(n10707), .ZN(
        n10713) );
  NAND2_X1 U13334 ( .A1(n10713), .A2(n15526), .ZN(n10709) );
  OAI21_X1 U13335 ( .B1(n15526), .B2(n10710), .A(n10709), .ZN(P1_U3465) );
  NAND2_X1 U13336 ( .A1(n10713), .A2(n15537), .ZN(n10714) );
  OAI21_X1 U13337 ( .B1(n15537), .B2(n10168), .A(n10714), .ZN(P1_U3530) );
  NAND2_X1 U13338 ( .A1(n10715), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10716) );
  MUX2_X1 U13339 ( .A(P1_IR_REG_31__SCAN_IN), .B(n10716), .S(
        P1_IR_REG_15__SCAN_IN), .Z(n10718) );
  AND2_X1 U13340 ( .A1(n10718), .A2(n10717), .ZN(n12346) );
  INV_X1 U13341 ( .A(n12346), .ZN(n15471) );
  OAI222_X1 U13342 ( .A1(P1_U3086), .A2(n15471), .B1(n15238), .B2(n10720), 
        .C1(n10719), .C2(n15239), .ZN(P1_U3340) );
  XNOR2_X1 U13343 ( .A(n10722), .B(n10721), .ZN(n10726) );
  AOI22_X1 U13344 ( .A1(n13951), .A2(n13983), .B1(n13981), .B2(n12105), .ZN(
        n10901) );
  OAI22_X1 U13345 ( .A1(n13953), .A2(n10901), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10080), .ZN(n10723) );
  AOI21_X1 U13346 ( .B1(n11551), .B2(n13944), .A(n10723), .ZN(n10725) );
  NAND2_X1 U13347 ( .A1(n15350), .A2(n12924), .ZN(n10724) );
  OAI211_X1 U13348 ( .C1(n10726), .C2(n13935), .A(n10725), .B(n10724), .ZN(
        P2_U3185) );
  MUX2_X1 U13349 ( .A(P3_REG2_REG_1__SCAN_IN), .B(P3_REG1_REG_1__SCAN_IN), .S(
        n6945), .Z(n10727) );
  NOR2_X1 U13350 ( .A1(n10727), .A2(n10826), .ZN(n10729) );
  AOI21_X1 U13351 ( .B1(n10727), .B2(n10826), .A(n10729), .ZN(n10822) );
  NOR2_X1 U13352 ( .A1(n10728), .A2(n10763), .ZN(n15697) );
  INV_X1 U13353 ( .A(n10729), .ZN(n11188) );
  INV_X1 U13354 ( .A(P3_REG2_REG_2__SCAN_IN), .ZN(n11059) );
  MUX2_X1 U13355 ( .A(n11059), .B(n10766), .S(n6945), .Z(n10730) );
  NAND2_X1 U13356 ( .A1(n10730), .A2(n11194), .ZN(n10734) );
  INV_X1 U13357 ( .A(n10730), .ZN(n10732) );
  NAND2_X1 U13358 ( .A1(n10732), .A2(n10731), .ZN(n10733) );
  NAND2_X1 U13359 ( .A1(n10734), .A2(n10733), .ZN(n11187) );
  INV_X1 U13360 ( .A(n10734), .ZN(n10842) );
  INV_X1 U13361 ( .A(P3_REG2_REG_3__SCAN_IN), .ZN(n10736) );
  MUX2_X1 U13362 ( .A(n10736), .B(n10735), .S(n6945), .Z(n10737) );
  NAND2_X1 U13363 ( .A1(n10737), .A2(n10768), .ZN(n10740) );
  INV_X1 U13364 ( .A(n10737), .ZN(n10738) );
  NAND2_X1 U13365 ( .A1(n10738), .A2(n10857), .ZN(n10739) );
  AND2_X1 U13366 ( .A1(n10740), .A2(n10739), .ZN(n10841) );
  OAI21_X1 U13367 ( .B1(n11186), .B2(n10842), .A(n10841), .ZN(n10840) );
  NAND2_X1 U13368 ( .A1(n10840), .A2(n10740), .ZN(n10743) );
  MUX2_X1 U13369 ( .A(P3_REG2_REG_4__SCAN_IN), .B(P3_REG1_REG_4__SCAN_IN), .S(
        n6945), .Z(n10792) );
  XNOR2_X1 U13370 ( .A(n10792), .B(n10741), .ZN(n10742) );
  NAND2_X1 U13371 ( .A1(n10743), .A2(n10742), .ZN(n10791) );
  OAI21_X1 U13372 ( .B1(n10743), .B2(n10742), .A(n10791), .ZN(n10783) );
  INV_X1 U13373 ( .A(n10934), .ZN(n10744) );
  NAND2_X1 U13374 ( .A1(n10744), .A2(n11598), .ZN(n10776) );
  NAND2_X1 U13375 ( .A1(n10746), .A2(n10745), .ZN(n10747) );
  NAND2_X1 U13376 ( .A1(n10748), .A2(n10747), .ZN(n10775) );
  INV_X1 U13377 ( .A(n10775), .ZN(n10749) );
  NAND2_X1 U13378 ( .A1(n10776), .A2(n10749), .ZN(n10773) );
  MUX2_X1 U13379 ( .A(n10773), .B(n13358), .S(n10750), .Z(n13521) );
  NOR2_X1 U13380 ( .A1(n13521), .A2(n10801), .ZN(n10782) );
  INV_X1 U13381 ( .A(P3_REG2_REG_0__SCAN_IN), .ZN(n15690) );
  NOR2_X1 U13382 ( .A1(n15690), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n10751) );
  NAND2_X1 U13383 ( .A1(n9031), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n10752) );
  OAI21_X1 U13384 ( .B1(n10826), .B2(n10751), .A(n10752), .ZN(n10813) );
  INV_X1 U13385 ( .A(P3_REG2_REG_1__SCAN_IN), .ZN(n15732) );
  NAND2_X1 U13386 ( .A1(n10815), .A2(n10752), .ZN(n11178) );
  NAND2_X1 U13387 ( .A1(n11178), .A2(n11179), .ZN(n11177) );
  OR2_X1 U13388 ( .A1(n11194), .A2(n11059), .ZN(n10754) );
  NAND2_X1 U13389 ( .A1(n10755), .A2(n10857), .ZN(n10756) );
  NAND2_X1 U13390 ( .A1(P3_REG2_REG_4__SCAN_IN), .A2(n10801), .ZN(n10757) );
  OAI21_X1 U13391 ( .B1(P3_REG2_REG_4__SCAN_IN), .B2(n10801), .A(n10757), .ZN(
        n10758) );
  AOI21_X1 U13392 ( .B1(n10759), .B2(n10758), .A(n10800), .ZN(n10780) );
  NAND2_X1 U13393 ( .A1(n10762), .A2(n10761), .ZN(n11175) );
  NAND2_X1 U13394 ( .A1(P3_REG1_REG_0__SCAN_IN), .A2(n10763), .ZN(n10764) );
  OR2_X1 U13395 ( .A1(P3_IR_REG_1__SCAN_IN), .A2(n10764), .ZN(n10765) );
  OR2_X1 U13396 ( .A1(n11194), .A2(n10766), .ZN(n10767) );
  NAND2_X1 U13397 ( .A1(n10769), .A2(n10857), .ZN(n10770) );
  NAND2_X1 U13398 ( .A1(P3_REG1_REG_4__SCAN_IN), .A2(n10801), .ZN(n10771) );
  AND2_X1 U13399 ( .A1(n6844), .A2(n10772), .ZN(n10774) );
  INV_X1 U13400 ( .A(n15693), .ZN(n13471) );
  OAI21_X1 U13401 ( .B1(n10786), .B2(n10774), .A(n13471), .ZN(n10779) );
  NOR2_X1 U13402 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n10777), .ZN(n11013) );
  AOI21_X1 U13403 ( .B1(n15698), .B2(P3_ADDR_REG_4__SCAN_IN), .A(n11013), .ZN(
        n10778) );
  OAI211_X1 U13404 ( .C1(n10780), .C2(n15694), .A(n10779), .B(n10778), .ZN(
        n10781) );
  AOI211_X1 U13405 ( .C1(n10783), .C2(n13529), .A(n10782), .B(n10781), .ZN(
        n10784) );
  INV_X1 U13406 ( .A(n10784), .ZN(P3_U3186) );
  NOR2_X1 U13407 ( .A1(n10802), .A2(n10787), .ZN(n10788) );
  XOR2_X1 U13408 ( .A(n10886), .B(n10787), .Z(n10884) );
  NOR2_X1 U13409 ( .A1(n9092), .A2(n10884), .ZN(n10883) );
  AOI22_X1 U13410 ( .A1(n10809), .A2(P3_REG1_REG_6__SCAN_IN), .B1(n9109), .B2(
        n10869), .ZN(n10789) );
  AOI21_X1 U13411 ( .B1(n10790), .B2(n10789), .A(n10861), .ZN(n10812) );
  OAI21_X1 U13412 ( .B1(n10792), .B2(n10801), .A(n10791), .ZN(n10878) );
  MUX2_X1 U13413 ( .A(P3_REG2_REG_5__SCAN_IN), .B(P3_REG1_REG_5__SCAN_IN), .S(
        n6945), .Z(n10793) );
  NAND2_X1 U13414 ( .A1(n10793), .A2(n10886), .ZN(n10879) );
  NAND2_X1 U13415 ( .A1(n10878), .A2(n10879), .ZN(n10877) );
  INV_X1 U13416 ( .A(n10793), .ZN(n10794) );
  NAND2_X1 U13417 ( .A1(n10794), .A2(n10802), .ZN(n10881) );
  NAND2_X1 U13418 ( .A1(n10877), .A2(n10881), .ZN(n10796) );
  MUX2_X1 U13419 ( .A(P3_REG2_REG_6__SCAN_IN), .B(P3_REG1_REG_6__SCAN_IN), .S(
        n6945), .Z(n10864) );
  XNOR2_X1 U13420 ( .A(n10864), .B(n10809), .ZN(n10795) );
  NAND2_X1 U13421 ( .A1(n10796), .A2(n10795), .ZN(n10863) );
  OAI21_X1 U13422 ( .B1(n10796), .B2(n10795), .A(n10863), .ZN(n10797) );
  NAND2_X1 U13423 ( .A1(n10797), .A2(n13529), .ZN(n10811) );
  INV_X1 U13424 ( .A(n15698), .ZN(n13492) );
  NOR2_X1 U13425 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n10798), .ZN(n11475) );
  INV_X1 U13426 ( .A(n11475), .ZN(n10799) );
  OAI21_X1 U13427 ( .B1(n13492), .B2(n7761), .A(n10799), .ZN(n10808) );
  INV_X1 U13428 ( .A(P3_REG2_REG_5__SCAN_IN), .ZN(n11434) );
  INV_X1 U13429 ( .A(P3_REG2_REG_6__SCAN_IN), .ZN(n15713) );
  AOI22_X1 U13430 ( .A1(n10809), .A2(P3_REG2_REG_6__SCAN_IN), .B1(n15713), 
        .B2(n10869), .ZN(n10804) );
  AOI21_X1 U13431 ( .B1(n10805), .B2(n10804), .A(n10868), .ZN(n10806) );
  NOR2_X1 U13432 ( .A1(n10806), .A2(n15694), .ZN(n10807) );
  AOI211_X1 U13433 ( .C1(n15699), .C2(n10809), .A(n10808), .B(n10807), .ZN(
        n10810) );
  OAI211_X1 U13434 ( .C1(n10812), .C2(n15693), .A(n10811), .B(n10810), .ZN(
        P3_U3188) );
  INV_X1 U13435 ( .A(n15694), .ZN(n11181) );
  NAND2_X1 U13436 ( .A1(n10813), .A2(n15732), .ZN(n10814) );
  NAND2_X1 U13437 ( .A1(n10815), .A2(n10814), .ZN(n10821) );
  NAND2_X1 U13438 ( .A1(n15698), .A2(P3_ADDR_REG_1__SCAN_IN), .ZN(n10816) );
  OAI21_X1 U13439 ( .B1(P3_STATE_REG_SCAN_IN), .B2(n15728), .A(n10816), .ZN(
        n10820) );
  AOI21_X1 U13440 ( .B1(n10818), .B2(n10817), .A(n15693), .ZN(n10819) );
  AOI211_X1 U13441 ( .C1(n11181), .C2(n10821), .A(n10820), .B(n10819), .ZN(
        n10825) );
  OAI21_X1 U13442 ( .B1(n10822), .B2(n15697), .A(n11189), .ZN(n10823) );
  NAND2_X1 U13443 ( .A1(n10823), .A2(n13529), .ZN(n10824) );
  OAI211_X1 U13444 ( .C1(n13521), .C2(n10826), .A(n10825), .B(n10824), .ZN(
        P3_U3183) );
  INV_X1 U13445 ( .A(n13350), .ZN(n11478) );
  INV_X1 U13446 ( .A(n10827), .ZN(n10828) );
  NAND2_X1 U13447 ( .A1(n10828), .A2(n10836), .ZN(n10831) );
  AND2_X1 U13448 ( .A1(n10832), .A2(n10831), .ZN(n10834) );
  OAI211_X1 U13449 ( .C1(n10834), .C2(n10833), .A(n13322), .B(n11008), .ZN(
        n10839) );
  NOR2_X1 U13450 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n10835), .ZN(n10850) );
  OAI22_X1 U13451 ( .A1(n13347), .A2(n15747), .B1(n10836), .B2(n13315), .ZN(
        n10837) );
  AOI211_X1 U13452 ( .C1(n13281), .C2(n11425), .A(n10850), .B(n10837), .ZN(
        n10838) );
  OAI211_X1 U13453 ( .C1(P3_REG3_REG_3__SCAN_IN), .C2(n11478), .A(n10839), .B(
        n10838), .ZN(P3_U3158) );
  INV_X1 U13454 ( .A(n10840), .ZN(n10844) );
  NOR3_X1 U13455 ( .A1(n11186), .A2(n10842), .A3(n10841), .ZN(n10843) );
  OAI21_X1 U13456 ( .B1(n10844), .B2(n10843), .A(n13529), .ZN(n10856) );
  OAI21_X1 U13457 ( .B1(n10846), .B2(P3_REG1_REG_3__SCAN_IN), .A(n10845), .ZN(
        n10854) );
  OAI21_X1 U13458 ( .B1(n10848), .B2(P3_REG2_REG_3__SCAN_IN), .A(n10847), .ZN(
        n10849) );
  NAND2_X1 U13459 ( .A1(n11181), .A2(n10849), .ZN(n10852) );
  INV_X1 U13460 ( .A(n10850), .ZN(n10851) );
  OAI211_X1 U13461 ( .C1(n13492), .C2(n8121), .A(n10852), .B(n10851), .ZN(
        n10853) );
  AOI21_X1 U13462 ( .B1(n13471), .B2(n10854), .A(n10853), .ZN(n10855) );
  OAI211_X1 U13463 ( .C1(n13521), .C2(n10857), .A(n10856), .B(n10855), .ZN(
        P3_U3185) );
  NAND2_X1 U13464 ( .A1(n13333), .A2(P3_U3897), .ZN(n10858) );
  OAI21_X1 U13465 ( .B1(n10860), .B2(n10859), .A(n10858), .ZN(P3_U3516) );
  AOI21_X1 U13466 ( .B1(n9123), .B2(n10862), .A(n10973), .ZN(n10876) );
  MUX2_X1 U13467 ( .A(P3_REG2_REG_7__SCAN_IN), .B(P3_REG1_REG_7__SCAN_IN), .S(
        n6945), .Z(n10978) );
  XNOR2_X1 U13468 ( .A(n10978), .B(n10986), .ZN(n10980) );
  XNOR2_X1 U13469 ( .A(n10981), .B(n10980), .ZN(n10865) );
  NAND2_X1 U13470 ( .A1(n10865), .A2(n13529), .ZN(n10875) );
  INV_X1 U13471 ( .A(P3_ADDR_REG_7__SCAN_IN), .ZN(n10867) );
  OR2_X1 U13472 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n10866), .ZN(n11638) );
  OAI21_X1 U13473 ( .B1(n13492), .B2(n10867), .A(n11638), .ZN(n10873) );
  INV_X1 U13474 ( .A(P3_REG2_REG_7__SCAN_IN), .ZN(n11759) );
  AOI21_X1 U13475 ( .B1(n11759), .B2(n10870), .A(n10987), .ZN(n10871) );
  NOR2_X1 U13476 ( .A1(n10871), .A2(n15694), .ZN(n10872) );
  AOI211_X1 U13477 ( .C1(n15699), .C2(n10986), .A(n10873), .B(n10872), .ZN(
        n10874) );
  OAI211_X1 U13478 ( .C1(n10876), .C2(n15693), .A(n10875), .B(n10874), .ZN(
        P3_U3189) );
  INV_X1 U13479 ( .A(n10877), .ZN(n10882) );
  AOI21_X1 U13480 ( .B1(n10881), .B2(n10879), .A(n10878), .ZN(n10880) );
  AOI21_X1 U13481 ( .B1(n10882), .B2(n10881), .A(n10880), .ZN(n10895) );
  AOI21_X1 U13482 ( .B1(n9092), .B2(n10884), .A(n10883), .ZN(n10885) );
  OAI22_X1 U13483 ( .A1(n13521), .A2(n10886), .B1(n10885), .B2(n15693), .ZN(
        n10893) );
  AOI21_X1 U13484 ( .B1(n11434), .B2(n10888), .A(n10887), .ZN(n10891) );
  NOR2_X1 U13485 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n10889), .ZN(n11303) );
  AOI21_X1 U13486 ( .B1(n15698), .B2(P3_ADDR_REG_5__SCAN_IN), .A(n11303), .ZN(
        n10890) );
  OAI21_X1 U13487 ( .B1(n10891), .B2(n15694), .A(n10890), .ZN(n10892) );
  NOR2_X1 U13488 ( .A1(n10893), .A2(n10892), .ZN(n10894) );
  OAI21_X1 U13489 ( .B1(n10895), .B2(n15692), .A(n10894), .ZN(P3_U3187) );
  XNOR2_X1 U13490 ( .A(n10896), .B(n13129), .ZN(n11557) );
  NAND2_X1 U13491 ( .A1(n11111), .A2(n12924), .ZN(n10897) );
  NAND2_X1 U13492 ( .A1(n10897), .A2(n14206), .ZN(n10898) );
  NOR2_X1 U13493 ( .A1(n11091), .A2(n10898), .ZN(n11550) );
  XNOR2_X1 U13494 ( .A(n10900), .B(n10899), .ZN(n10902) );
  OAI21_X1 U13495 ( .B1(n10902), .B2(n14220), .A(n10901), .ZN(n11554) );
  AOI211_X1 U13496 ( .C1(n15366), .C2(n11557), .A(n11550), .B(n11554), .ZN(
        n10907) );
  INV_X1 U13497 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n10903) );
  NOR2_X1 U13498 ( .A1(n15680), .A2(n10903), .ZN(n10904) );
  AOI21_X1 U13499 ( .B1(n14375), .B2(n12924), .A(n10904), .ZN(n10905) );
  OAI21_X1 U13500 ( .B1(n10907), .B2(n15678), .A(n10905), .ZN(P2_U3451) );
  AOI22_X1 U13501 ( .A1(n14313), .A2(n12924), .B1(n7435), .B2(
        P2_REG1_REG_7__SCAN_IN), .ZN(n10906) );
  OAI21_X1 U13502 ( .B1(n10907), .B2(n7435), .A(n10906), .ZN(P2_U3506) );
  INV_X1 U13503 ( .A(n15675), .ZN(n15662) );
  XNOR2_X1 U13504 ( .A(n10908), .B(n10912), .ZN(n11078) );
  INV_X1 U13505 ( .A(n11078), .ZN(n10917) );
  AOI21_X1 U13506 ( .B1(n11509), .B2(n12907), .A(n6670), .ZN(n10909) );
  AND2_X1 U13507 ( .A1(n10909), .A2(n11113), .ZN(n11075) );
  OAI21_X1 U13508 ( .B1(n10912), .B2(n10911), .A(n10910), .ZN(n10915) );
  NOR2_X1 U13509 ( .A1(n11078), .A2(n8992), .ZN(n10913) );
  AOI211_X1 U13510 ( .C1(n15617), .C2(n10915), .A(n10914), .B(n10913), .ZN(
        n11067) );
  INV_X1 U13511 ( .A(n11067), .ZN(n10916) );
  AOI211_X1 U13512 ( .C1(n15662), .C2(n10917), .A(n11075), .B(n10916), .ZN(
        n10922) );
  INV_X1 U13513 ( .A(n14375), .ZN(n14324) );
  INV_X1 U13514 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n10918) );
  OAI22_X1 U13515 ( .A1(n14324), .A2(n11073), .B1(n15680), .B2(n10918), .ZN(
        n10919) );
  INV_X1 U13516 ( .A(n10919), .ZN(n10920) );
  OAI21_X1 U13517 ( .B1(n10922), .B2(n15678), .A(n10920), .ZN(P2_U3445) );
  AOI22_X1 U13518 ( .A1(n14313), .A2(n12907), .B1(n7435), .B2(
        P2_REG1_REG_5__SCAN_IN), .ZN(n10921) );
  OAI21_X1 U13519 ( .B1(n10922), .B2(n7435), .A(n10921), .ZN(P2_U3504) );
  INV_X1 U13520 ( .A(n10923), .ZN(n10925) );
  OAI222_X1 U13521 ( .A1(P3_U3151), .A2(n10926), .B1(n13851), .B2(n10925), 
        .C1(n10924), .C2(n13840), .ZN(P3_U3275) );
  INV_X1 U13522 ( .A(n13827), .ZN(n10928) );
  NAND2_X1 U13523 ( .A1(n10928), .A2(n10927), .ZN(n10931) );
  NAND2_X1 U13524 ( .A1(n13827), .A2(n10929), .ZN(n10930) );
  MUX2_X1 U13525 ( .A(n10935), .B(P3_REG2_REG_0__SCAN_IN), .S(n15735), .Z(
        n10941) );
  INV_X1 U13526 ( .A(n10936), .ZN(n10938) );
  NOR2_X1 U13527 ( .A1(n15715), .A2(n15758), .ZN(n10937) );
  OAI22_X1 U13528 ( .A1(n13714), .A2(n10939), .B1(n15727), .B2(n15702), .ZN(
        n10940) );
  OR2_X1 U13529 ( .A1(n10941), .A2(n10940), .ZN(P3_U3233) );
  INV_X1 U13530 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n10968) );
  NAND2_X1 U13531 ( .A1(n10688), .A2(n11544), .ZN(n12613) );
  NAND2_X1 U13532 ( .A1(n10942), .A2(n12613), .ZN(n11525) );
  NAND2_X1 U13533 ( .A1(n10954), .A2(n15496), .ZN(n12617) );
  INV_X1 U13534 ( .A(n10954), .ZN(n10943) );
  NAND2_X1 U13535 ( .A1(n10943), .A2(n11538), .ZN(n12618) );
  NAND2_X1 U13536 ( .A1(n10954), .A2(n11538), .ZN(n10944) );
  NAND2_X1 U13537 ( .A1(n11524), .A2(n10944), .ZN(n10949) );
  INV_X2 U13538 ( .A(n9889), .ZN(n11026) );
  NAND2_X1 U13539 ( .A1(n10945), .A2(n11026), .ZN(n10947) );
  NAND2_X1 U13540 ( .A1(n12415), .A2(n15456), .ZN(n10946) );
  NAND2_X1 U13541 ( .A1(n11529), .A2(n12620), .ZN(n11387) );
  OAI21_X1 U13542 ( .B1(n10949), .B2(n10950), .A(n11412), .ZN(n11212) );
  INV_X1 U13543 ( .A(n11212), .ZN(n10966) );
  INV_X1 U13544 ( .A(n10950), .ZN(n12798) );
  NAND2_X1 U13545 ( .A1(n10952), .A2(n10951), .ZN(n11528) );
  NAND2_X1 U13546 ( .A1(n11528), .A2(n12616), .ZN(n11527) );
  NAND2_X1 U13547 ( .A1(n11527), .A2(n12617), .ZN(n10953) );
  NAND2_X1 U13548 ( .A1(n10953), .A2(n12798), .ZN(n11388) );
  OAI21_X1 U13549 ( .B1(n12798), .B2(n10953), .A(n11388), .ZN(n10963) );
  OR2_X1 U13550 ( .A1(n10954), .A2(n15069), .ZN(n10961) );
  NAND2_X1 U13551 ( .A1(n12519), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n10959) );
  NAND2_X1 U13552 ( .A1(n6680), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n10958) );
  AOI21_X1 U13553 ( .B1(P1_REG3_REG_4__SCAN_IN), .B2(P1_REG3_REG_3__SCAN_IN), 
        .A(P1_REG3_REG_5__SCAN_IN), .ZN(n10955) );
  NOR2_X1 U13554 ( .A1(n10955), .A2(n11039), .ZN(n11485) );
  NAND2_X1 U13555 ( .A1(n6677), .A2(n11485), .ZN(n10957) );
  NAND2_X1 U13556 ( .A1(n6878), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n10956) );
  NAND2_X1 U13557 ( .A1(n14704), .A2(n15002), .ZN(n10960) );
  AND2_X1 U13558 ( .A1(n10961), .A2(n10960), .ZN(n11086) );
  INV_X1 U13559 ( .A(n11086), .ZN(n10962) );
  AOI21_X1 U13560 ( .B1(n10963), .B2(n15280), .A(n10962), .ZN(n11215) );
  NAND2_X1 U13561 ( .A1(n11534), .A2(n11538), .ZN(n11535) );
  INV_X1 U13562 ( .A(n11483), .ZN(n10964) );
  AOI211_X1 U13563 ( .C1(n12620), .C2(n11535), .A(n15488), .B(n10964), .ZN(
        n11209) );
  AOI21_X1 U13564 ( .B1(n12620), .B2(n15495), .A(n11209), .ZN(n10965) );
  OAI211_X1 U13565 ( .C1(n10966), .C2(n15482), .A(n11215), .B(n10965), .ZN(
        n10969) );
  NAND2_X1 U13566 ( .A1(n10969), .A2(n15526), .ZN(n10967) );
  OAI21_X1 U13567 ( .B1(n15526), .B2(n10968), .A(n10967), .ZN(P1_U3471) );
  NAND2_X1 U13568 ( .A1(n10969), .A2(n15537), .ZN(n10970) );
  OAI21_X1 U13569 ( .B1(n15537), .B2(n10971), .A(n10970), .ZN(P1_U3532) );
  NOR2_X1 U13570 ( .A1(n10986), .A2(n10972), .ZN(n10974) );
  NAND2_X1 U13571 ( .A1(P3_REG1_REG_8__SCAN_IN), .A2(n11331), .ZN(n10975) );
  OAI21_X1 U13572 ( .B1(P3_REG1_REG_8__SCAN_IN), .B2(n11331), .A(n10975), .ZN(
        n10976) );
  AOI21_X1 U13573 ( .B1(n10977), .B2(n10976), .A(n11326), .ZN(n10997) );
  INV_X1 U13574 ( .A(n10978), .ZN(n10979) );
  MUX2_X1 U13575 ( .A(P3_REG2_REG_8__SCAN_IN), .B(P3_REG1_REG_8__SCAN_IN), .S(
        n6945), .Z(n11317) );
  XNOR2_X1 U13576 ( .A(n11317), .B(n11331), .ZN(n11318) );
  XNOR2_X1 U13577 ( .A(n11319), .B(n11318), .ZN(n10982) );
  NAND2_X1 U13578 ( .A1(n10982), .A2(n13529), .ZN(n10996) );
  INV_X1 U13579 ( .A(n11331), .ZN(n10994) );
  NOR2_X1 U13580 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n10983), .ZN(n11854) );
  INV_X1 U13581 ( .A(n11854), .ZN(n10984) );
  OAI21_X1 U13582 ( .B1(n13492), .B2(n8104), .A(n10984), .ZN(n10993) );
  NAND2_X1 U13583 ( .A1(P3_REG2_REG_8__SCAN_IN), .A2(n11331), .ZN(n10988) );
  OAI21_X1 U13584 ( .B1(P3_REG2_REG_8__SCAN_IN), .B2(n11331), .A(n10988), .ZN(
        n10989) );
  AOI21_X1 U13585 ( .B1(n10990), .B2(n10989), .A(n11330), .ZN(n10991) );
  NOR2_X1 U13586 ( .A1(n10991), .A2(n15694), .ZN(n10992) );
  AOI211_X1 U13587 ( .C1(n15699), .C2(n10994), .A(n10993), .B(n10992), .ZN(
        n10995) );
  OAI211_X1 U13588 ( .C1(n10997), .C2(n15693), .A(n10996), .B(n10995), .ZN(
        P3_U3190) );
  XOR2_X1 U13589 ( .A(n11000), .B(n10998), .Z(n15748) );
  AND2_X1 U13590 ( .A1(n15715), .A2(n10999), .ZN(n11216) );
  INV_X1 U13591 ( .A(n13561), .ZN(n15729) );
  INV_X1 U13592 ( .A(n13554), .ZN(n15764) );
  AOI22_X1 U13593 ( .A1(n15717), .A2(n15718), .B1(n11425), .B2(n15719), .ZN(
        n11003) );
  OAI211_X1 U13594 ( .C1(n7742), .C2(n9696), .A(n15722), .B(n11001), .ZN(
        n11002) );
  OAI211_X1 U13595 ( .C1(n15748), .C2(n15764), .A(n11003), .B(n11002), .ZN(
        n15750) );
  NAND2_X1 U13596 ( .A1(n15750), .A2(n15733), .ZN(n11006) );
  OAI22_X1 U13597 ( .A1(n13714), .A2(n15747), .B1(P3_REG3_REG_3__SCAN_IN), 
        .B2(n15727), .ZN(n11004) );
  AOI21_X1 U13598 ( .B1(n15735), .B2(P3_REG2_REG_3__SCAN_IN), .A(n11004), .ZN(
        n11005) );
  OAI211_X1 U13599 ( .C1(n15748), .C2(n15729), .A(n11006), .B(n11005), .ZN(
        P3_U3230) );
  XNOR2_X1 U13600 ( .A(n11280), .B(n13207), .ZN(n11009) );
  NAND2_X1 U13601 ( .A1(n11301), .A2(n11009), .ZN(n11297) );
  OAI21_X1 U13602 ( .B1(n11301), .B2(n11009), .A(n11297), .ZN(n11010) );
  AOI21_X1 U13603 ( .B1(n11011), .B2(n11010), .A(n11298), .ZN(n11017) );
  OAI22_X1 U13604 ( .A1(n13347), .A2(n11280), .B1(n11224), .B2(n13315), .ZN(
        n11012) );
  AOI211_X1 U13605 ( .C1(n13281), .C2(n11014), .A(n11013), .B(n11012), .ZN(
        n11016) );
  NAND2_X1 U13606 ( .A1(n13350), .A2(n11229), .ZN(n11015) );
  OAI211_X1 U13607 ( .C1(n11017), .C2(n13352), .A(n11016), .B(n11015), .ZN(
        P3_U3170) );
  NAND2_X1 U13608 ( .A1(n14705), .A2(n6676), .ZN(n11019) );
  INV_X2 U13609 ( .A(n6667), .ZN(n14511) );
  NAND2_X1 U13610 ( .A1(n14511), .A2(n12620), .ZN(n11018) );
  NAND2_X1 U13611 ( .A1(n11019), .A2(n11018), .ZN(n11020) );
  XNOR2_X1 U13612 ( .A(n11020), .B(n9851), .ZN(n11082) );
  NAND2_X1 U13613 ( .A1(n14705), .A2(n14517), .ZN(n11022) );
  NAND2_X1 U13614 ( .A1(n9893), .A2(n12620), .ZN(n11021) );
  NAND2_X1 U13615 ( .A1(n11024), .A2(n11023), .ZN(n11080) );
  OAI21_X1 U13616 ( .B1(n11082), .B2(n11081), .A(n11080), .ZN(n11025) );
  NAND2_X1 U13617 ( .A1(n14704), .A2(n9893), .ZN(n11031) );
  NAND2_X1 U13618 ( .A1(n11027), .A2(n11026), .ZN(n11029) );
  AOI22_X1 U13619 ( .A1(n7282), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n12415), 
        .B2(n14761), .ZN(n11028) );
  NAND2_X1 U13620 ( .A1(n11029), .A2(n11028), .ZN(n12629) );
  NAND2_X1 U13621 ( .A1(n12629), .A2(n14511), .ZN(n11030) );
  NAND2_X1 U13622 ( .A1(n11031), .A2(n11030), .ZN(n11032) );
  XNOR2_X1 U13623 ( .A(n11032), .B(n6921), .ZN(n11036) );
  NAND2_X1 U13624 ( .A1(n14704), .A2(n14517), .ZN(n11034) );
  NAND2_X1 U13625 ( .A1(n12629), .A2(n9893), .ZN(n11033) );
  NAND2_X1 U13626 ( .A1(n11034), .A2(n11033), .ZN(n11035) );
  NOR2_X1 U13627 ( .A1(n11036), .A2(n11035), .ZN(n11236) );
  INV_X1 U13628 ( .A(n11236), .ZN(n11037) );
  NAND2_X1 U13629 ( .A1(n11036), .A2(n11035), .ZN(n11235) );
  NAND2_X1 U13630 ( .A1(n11037), .A2(n11235), .ZN(n11038) );
  XNOR2_X1 U13631 ( .A(n11237), .B(n11038), .ZN(n11048) );
  INV_X1 U13632 ( .A(n12629), .ZN(n15505) );
  NOR2_X1 U13633 ( .A1(n14683), .A2(n15505), .ZN(n11046) );
  NAND2_X1 U13634 ( .A1(n12519), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n11043) );
  NAND2_X1 U13635 ( .A1(n9864), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n11042) );
  OAI21_X1 U13636 ( .B1(n11039), .B2(P1_REG3_REG_6__SCAN_IN), .A(n11244), .ZN(
        n11591) );
  INV_X1 U13637 ( .A(n11591), .ZN(n11252) );
  NAND2_X1 U13638 ( .A1(n6677), .A2(n11252), .ZN(n11041) );
  NAND2_X1 U13639 ( .A1(n6878), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n11040) );
  INV_X1 U13640 ( .A(n14703), .ZN(n11391) );
  NAND2_X1 U13641 ( .A1(n14677), .A2(n14705), .ZN(n11044) );
  NAND2_X1 U13642 ( .A1(P1_REG3_REG_5__SCAN_IN), .A2(P1_U3086), .ZN(n14758) );
  OAI211_X1 U13643 ( .C1(n11391), .C2(n15384), .A(n11044), .B(n14758), .ZN(
        n11045) );
  AOI211_X1 U13644 ( .C1(n11485), .C2(n14680), .A(n11046), .B(n11045), .ZN(
        n11047) );
  OAI21_X1 U13645 ( .B1(n11048), .B2(n15392), .A(n11047), .ZN(P1_U3227) );
  OAI21_X1 U13646 ( .B1(n11050), .B2(n11053), .A(n11049), .ZN(n15744) );
  INV_X1 U13647 ( .A(n15744), .ZN(n11061) );
  NAND2_X1 U13648 ( .A1(n11051), .A2(n15765), .ZN(n15741) );
  NOR2_X1 U13649 ( .A1(n15741), .A2(n15715), .ZN(n11057) );
  XNOR2_X1 U13650 ( .A(n11052), .B(n11053), .ZN(n11056) );
  OAI22_X1 U13651 ( .A1(n6957), .A2(n13694), .B1(n11224), .B2(n13696), .ZN(
        n11054) );
  AOI21_X1 U13652 ( .B1(n15744), .B2(n13554), .A(n11054), .ZN(n11055) );
  OAI21_X1 U13653 ( .B1(n13691), .B2(n11056), .A(n11055), .ZN(n15742) );
  AOI211_X1 U13654 ( .C1(n15709), .C2(P3_REG3_REG_2__SCAN_IN), .A(n11057), .B(
        n15742), .ZN(n11058) );
  MUX2_X1 U13655 ( .A(n11059), .B(n11058), .S(n15733), .Z(n11060) );
  OAI21_X1 U13656 ( .B1(n11061), .B2(n15729), .A(n11060), .ZN(P3_U3231) );
  NAND2_X1 U13657 ( .A1(n13577), .A2(P3_U3897), .ZN(n11062) );
  OAI21_X1 U13658 ( .B1(P3_U3897), .B2(n11063), .A(n11062), .ZN(P3_U3517) );
  INV_X1 U13659 ( .A(n15633), .ZN(n11065) );
  NAND2_X1 U13660 ( .A1(n11065), .A2(n11064), .ZN(n11129) );
  INV_X2 U13661 ( .A(n15627), .ZN(n14226) );
  AND2_X1 U13662 ( .A1(n13159), .A2(n8325), .ZN(n11066) );
  NAND2_X1 U13663 ( .A1(n14226), .A2(n11066), .ZN(n15623) );
  MUX2_X1 U13664 ( .A(n11068), .B(n11067), .S(n14226), .Z(n11077) );
  INV_X1 U13665 ( .A(n11069), .ZN(n11070) );
  INV_X1 U13666 ( .A(n11071), .ZN(n11072) );
  OAI22_X1 U13667 ( .A1(n14157), .A2(n11073), .B1(n11072), .B2(n15621), .ZN(
        n11074) );
  AOI21_X1 U13668 ( .B1(n14160), .B2(n11075), .A(n11074), .ZN(n11076) );
  OAI211_X1 U13669 ( .C1(n11078), .C2(n15623), .A(n11077), .B(n11076), .ZN(
        P2_U3260) );
  NAND2_X1 U13670 ( .A1(n7401), .A2(n11080), .ZN(n11084) );
  XNOR2_X1 U13671 ( .A(n11082), .B(n11081), .ZN(n11083) );
  XNOR2_X1 U13672 ( .A(n11084), .B(n11083), .ZN(n11085) );
  NAND2_X1 U13673 ( .A1(n11085), .A2(n14675), .ZN(n11089) );
  NAND2_X1 U13674 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_U3086), .ZN(n15460) );
  OAI21_X1 U13675 ( .B1(n11086), .B2(n14668), .A(n15460), .ZN(n11087) );
  AOI21_X1 U13676 ( .B1(n14680), .B2(n11204), .A(n11087), .ZN(n11088) );
  OAI211_X1 U13677 ( .C1(n11410), .C2(n14683), .A(n11089), .B(n11088), .ZN(
        P1_U3230) );
  XNOR2_X1 U13678 ( .A(n11090), .B(n13130), .ZN(n11131) );
  OR2_X1 U13679 ( .A1(n11091), .A2(n11137), .ZN(n11092) );
  AND3_X1 U13680 ( .A1(n11150), .A2(n11092), .A3(n14206), .ZN(n11139) );
  XNOR2_X1 U13681 ( .A(n11094), .B(n11093), .ZN(n11095) );
  AOI22_X1 U13682 ( .A1(n13951), .A2(n13982), .B1(n13980), .B2(n12105), .ZN(
        n11125) );
  OAI21_X1 U13683 ( .B1(n11095), .B2(n14220), .A(n11125), .ZN(n11132) );
  AOI211_X1 U13684 ( .C1(n15366), .C2(n11131), .A(n11139), .B(n11132), .ZN(
        n11100) );
  INV_X1 U13685 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n11096) );
  OAI22_X1 U13686 ( .A1(n14324), .A2(n11137), .B1(n15680), .B2(n11096), .ZN(
        n11097) );
  INV_X1 U13687 ( .A(n11097), .ZN(n11098) );
  OAI21_X1 U13688 ( .B1(n11100), .B2(n15678), .A(n11098), .ZN(P2_U3454) );
  AOI22_X1 U13689 ( .A1(n14313), .A2(n12935), .B1(n7435), .B2(
        P2_REG1_REG_8__SCAN_IN), .ZN(n11099) );
  OAI21_X1 U13690 ( .B1(n11100), .B2(n7435), .A(n11099), .ZN(P2_U3507) );
  NAND2_X1 U13691 ( .A1(n13358), .A2(P3_DATAO_REG_30__SCAN_IN), .ZN(n11101) );
  OAI21_X1 U13692 ( .B1(n11102), .B2(n13358), .A(n11101), .ZN(P3_U3521) );
  XNOR2_X1 U13693 ( .A(n11104), .B(n11103), .ZN(n15676) );
  OAI21_X1 U13694 ( .B1(n11106), .B2(n13128), .A(n11105), .ZN(n11109) );
  NOR2_X1 U13695 ( .A1(n15676), .A2(n8992), .ZN(n11107) );
  AOI211_X1 U13696 ( .C1(n15617), .C2(n11109), .A(n11108), .B(n11107), .ZN(
        n15674) );
  MUX2_X1 U13697 ( .A(n11110), .B(n15674), .S(n14226), .Z(n11118) );
  INV_X1 U13698 ( .A(n11111), .ZN(n11112) );
  AOI211_X1 U13699 ( .C1(n15671), .C2(n11113), .A(n6670), .B(n11112), .ZN(
        n15670) );
  INV_X1 U13700 ( .A(n15671), .ZN(n11115) );
  OAI22_X1 U13701 ( .A1(n14157), .A2(n11115), .B1(n15621), .B2(n11114), .ZN(
        n11116) );
  AOI21_X1 U13702 ( .B1(n15670), .B2(n14160), .A(n11116), .ZN(n11117) );
  OAI211_X1 U13703 ( .C1(n15676), .C2(n15623), .A(n11118), .B(n11117), .ZN(
        P2_U3259) );
  INV_X1 U13704 ( .A(n11119), .ZN(n11120) );
  AOI21_X1 U13705 ( .B1(n11122), .B2(n11121), .A(n11120), .ZN(n11128) );
  NAND2_X1 U13706 ( .A1(n13944), .A2(n11135), .ZN(n11124) );
  OAI211_X1 U13707 ( .C1(n11125), .C2(n13953), .A(n11124), .B(n11123), .ZN(
        n11126) );
  AOI21_X1 U13708 ( .B1(n12935), .B2(n15350), .A(n11126), .ZN(n11127) );
  OAI21_X1 U13709 ( .B1(n11128), .B2(n13935), .A(n11127), .ZN(P2_U3193) );
  OR2_X1 U13710 ( .A1(n11129), .A2(n8992), .ZN(n11130) );
  INV_X1 U13711 ( .A(n11131), .ZN(n11142) );
  INV_X1 U13712 ( .A(n11132), .ZN(n11133) );
  MUX2_X1 U13713 ( .A(n11134), .B(n11133), .S(n14226), .Z(n11141) );
  INV_X1 U13714 ( .A(n11135), .ZN(n11136) );
  OAI22_X1 U13715 ( .A1(n14157), .A2(n11137), .B1(n15621), .B2(n11136), .ZN(
        n11138) );
  AOI21_X1 U13716 ( .B1(n11139), .B2(n14160), .A(n11138), .ZN(n11140) );
  OAI211_X1 U13717 ( .C1(n14234), .C2(n11142), .A(n11141), .B(n11140), .ZN(
        P2_U3257) );
  XNOR2_X1 U13718 ( .A(n11143), .B(n11144), .ZN(n11290) );
  INV_X1 U13719 ( .A(n11290), .ZN(n11155) );
  XNOR2_X1 U13720 ( .A(n11145), .B(n13133), .ZN(n11148) );
  NAND2_X1 U13721 ( .A1(n13981), .A2(n13951), .ZN(n11147) );
  NAND2_X1 U13722 ( .A1(n13979), .A2(n13952), .ZN(n11146) );
  AND2_X1 U13723 ( .A1(n11147), .A2(n11146), .ZN(n11269) );
  OAI21_X1 U13724 ( .B1(n11148), .B2(n14220), .A(n11269), .ZN(n11288) );
  NAND2_X1 U13725 ( .A1(n11288), .A2(n14226), .ZN(n11154) );
  INV_X1 U13726 ( .A(n11368), .ZN(n11149) );
  AOI211_X1 U13727 ( .C1(n12940), .C2(n11150), .A(n6670), .B(n11149), .ZN(
        n11289) );
  INV_X1 U13728 ( .A(n12940), .ZN(n11292) );
  INV_X1 U13729 ( .A(n15621), .ZN(n14208) );
  AOI22_X1 U13730 ( .A1(n15627), .A2(P2_REG2_REG_9__SCAN_IN), .B1(n11271), 
        .B2(n14208), .ZN(n11151) );
  OAI21_X1 U13731 ( .B1(n11292), .B2(n14157), .A(n11151), .ZN(n11152) );
  AOI21_X1 U13732 ( .B1(n11289), .B2(n14160), .A(n11152), .ZN(n11153) );
  OAI211_X1 U13733 ( .C1(n14234), .C2(n11155), .A(n11154), .B(n11153), .ZN(
        P2_U3256) );
  XNOR2_X1 U13734 ( .A(n11156), .B(n11162), .ZN(n15655) );
  AOI211_X1 U13735 ( .C1(n15652), .C2(n11157), .A(n6670), .B(n11511), .ZN(
        n15651) );
  OAI22_X1 U13736 ( .A1(n14157), .A2(n11158), .B1(P2_REG3_REG_3__SCAN_IN), 
        .B2(n15621), .ZN(n11159) );
  AOI21_X1 U13737 ( .B1(n14160), .B2(n15651), .A(n11159), .ZN(n11167) );
  OAI21_X1 U13738 ( .B1(n11162), .B2(n11161), .A(n11160), .ZN(n11164) );
  AOI21_X1 U13739 ( .B1(n11164), .B2(n15617), .A(n11163), .ZN(n15653) );
  MUX2_X1 U13740 ( .A(n11165), .B(n15653), .S(n14226), .Z(n11166) );
  OAI211_X1 U13741 ( .C1(n14234), .C2(n15655), .A(n11167), .B(n11166), .ZN(
        P2_U3262) );
  INV_X1 U13742 ( .A(n11168), .ZN(n11169) );
  OAI222_X1 U13743 ( .A1(P3_U3151), .A2(n11171), .B1(n13840), .B2(n11170), 
        .C1(n13851), .C2(n11169), .ZN(P3_U3274) );
  NAND2_X1 U13744 ( .A1(n15303), .A2(P3_U3897), .ZN(n11172) );
  OAI21_X1 U13745 ( .B1(P3_U3897), .B2(n11173), .A(n11172), .ZN(P3_U3522) );
  NAND2_X1 U13746 ( .A1(n13471), .A2(n11176), .ZN(n11185) );
  OAI21_X1 U13747 ( .B1(n11179), .B2(n11178), .A(n11177), .ZN(n11180) );
  NAND2_X1 U13748 ( .A1(n11181), .A2(n11180), .ZN(n11184) );
  NOR2_X1 U13749 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n10682), .ZN(n11182) );
  AOI21_X1 U13750 ( .B1(n15698), .B2(P3_ADDR_REG_2__SCAN_IN), .A(n11182), .ZN(
        n11183) );
  NAND3_X1 U13751 ( .A1(n11185), .A2(n11184), .A3(n11183), .ZN(n11193) );
  INV_X1 U13752 ( .A(n11186), .ZN(n11191) );
  NAND3_X1 U13753 ( .A1(n11189), .A2(n11188), .A3(n11187), .ZN(n11190) );
  AOI21_X1 U13754 ( .B1(n11191), .B2(n11190), .A(n15692), .ZN(n11192) );
  AOI211_X1 U13755 ( .C1(n15699), .C2(n11194), .A(n11193), .B(n11192), .ZN(
        n11195) );
  INV_X1 U13756 ( .A(n11195), .ZN(P3_U3184) );
  INV_X1 U13757 ( .A(n13565), .ZN(n11196) );
  NAND2_X1 U13758 ( .A1(n11196), .A2(P3_U3897), .ZN(n11197) );
  OAI21_X1 U13759 ( .B1(P3_U3897), .B2(n11198), .A(n11197), .ZN(P3_U3518) );
  INV_X1 U13760 ( .A(n12584), .ZN(n11202) );
  NOR2_X1 U13761 ( .A1(n15013), .A2(n11410), .ZN(n11208) );
  INV_X1 U13762 ( .A(n11204), .ZN(n11205) );
  OAI22_X1 U13763 ( .A1(n15093), .A2(n11206), .B1(n11205), .B2(n15058), .ZN(
        n11207) );
  AOI211_X1 U13764 ( .C1(n11209), .C2(n15293), .A(n11208), .B(n11207), .ZN(
        n11214) );
  INV_X1 U13765 ( .A(n11210), .ZN(n11211) );
  NAND2_X1 U13766 ( .A1(n11212), .A2(n15294), .ZN(n11213) );
  OAI211_X1 U13767 ( .C1(n11215), .C2(n15067), .A(n11214), .B(n11213), .ZN(
        P1_U3289) );
  OR2_X1 U13768 ( .A1(n13554), .A2(n11216), .ZN(n15703) );
  OAI21_X1 U13769 ( .B1(n11219), .B2(n11218), .A(n11217), .ZN(n11220) );
  INV_X1 U13770 ( .A(n11220), .ZN(n11275) );
  INV_X1 U13771 ( .A(P3_REG2_REG_4__SCAN_IN), .ZN(n11228) );
  OAI211_X1 U13772 ( .C1(n11223), .C2(n11222), .A(n11221), .B(n15722), .ZN(
        n11227) );
  OAI22_X1 U13773 ( .A1(n11792), .A2(n13696), .B1(n11224), .B2(n13694), .ZN(
        n11225) );
  INV_X1 U13774 ( .A(n11225), .ZN(n11226) );
  AND2_X1 U13775 ( .A1(n11227), .A2(n11226), .ZN(n11274) );
  MUX2_X1 U13776 ( .A(n11228), .B(n11274), .S(n15733), .Z(n11231) );
  AOI22_X1 U13777 ( .A1(n15707), .A2(n9087), .B1(n15709), .B2(n11229), .ZN(
        n11230) );
  OAI211_X1 U13778 ( .C1(n13688), .C2(n11275), .A(n11231), .B(n11230), .ZN(
        P3_U3229) );
  NAND2_X1 U13779 ( .A1(n11232), .A2(n11026), .ZN(n11234) );
  AOI22_X1 U13780 ( .A1(n7282), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n12415), 
        .B2(n14777), .ZN(n11233) );
  NAND2_X1 U13781 ( .A1(n11234), .A2(n11233), .ZN(n12633) );
  INV_X1 U13782 ( .A(n12633), .ZN(n11592) );
  NAND2_X1 U13783 ( .A1(n12633), .A2(n14511), .ZN(n11239) );
  NAND2_X1 U13784 ( .A1(n14703), .A2(n9893), .ZN(n11238) );
  NAND2_X1 U13785 ( .A1(n11239), .A2(n11238), .ZN(n11240) );
  XNOR2_X1 U13786 ( .A(n11240), .B(n6921), .ZN(n11347) );
  AOI22_X1 U13787 ( .A1(n12633), .A2(n9893), .B1(n14517), .B2(n14703), .ZN(
        n11348) );
  XNOR2_X1 U13788 ( .A(n11347), .B(n11348), .ZN(n11241) );
  OAI211_X1 U13789 ( .C1(n11242), .C2(n11241), .A(n11351), .B(n14675), .ZN(
        n11254) );
  NAND2_X1 U13790 ( .A1(n12519), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n11249) );
  NAND2_X1 U13791 ( .A1(n9864), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n11248) );
  AND2_X1 U13792 ( .A1(n11244), .A2(n11243), .ZN(n11245) );
  NOR2_X1 U13793 ( .A1(n11356), .A2(n11245), .ZN(n11570) );
  NAND2_X1 U13794 ( .A1(n6677), .A2(n11570), .ZN(n11247) );
  NAND2_X1 U13795 ( .A1(n6878), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n11246) );
  NAND4_X1 U13796 ( .A1(n11249), .A2(n11248), .A3(n11247), .A4(n11246), .ZN(
        n14702) );
  NAND2_X1 U13797 ( .A1(n14677), .A2(n14704), .ZN(n11250) );
  NAND2_X1 U13798 ( .A1(P1_U3086), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n14774) );
  OAI211_X1 U13799 ( .C1(n11582), .C2(n15384), .A(n11250), .B(n14774), .ZN(
        n11251) );
  AOI21_X1 U13800 ( .B1(n14680), .B2(n11252), .A(n11251), .ZN(n11253) );
  OAI211_X1 U13801 ( .C1(n11592), .C2(n14683), .A(n11254), .B(n11253), .ZN(
        P1_U3239) );
  INV_X1 U13802 ( .A(n12411), .ZN(n11263) );
  INV_X1 U13803 ( .A(n14004), .ZN(n11255) );
  OAI222_X1 U13804 ( .A1(n12861), .A2(n11256), .B1(n14396), .B2(n11263), .C1(
        P2_U3088), .C2(n11255), .ZN(P2_U3309) );
  INV_X1 U13805 ( .A(n11257), .ZN(n11258) );
  NAND2_X1 U13806 ( .A1(n11258), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n11259) );
  MUX2_X1 U13807 ( .A(P1_IR_REG_31__SCAN_IN), .B(n11259), .S(
        P1_IR_REG_18__SCAN_IN), .Z(n11261) );
  AND2_X1 U13808 ( .A1(n11261), .A2(n11260), .ZN(n14828) );
  INV_X1 U13809 ( .A(n14828), .ZN(n14822) );
  OAI222_X1 U13810 ( .A1(n14822), .A2(P1_U3086), .B1(n15238), .B2(n11263), 
        .C1(n11262), .C2(n15239), .ZN(P1_U3337) );
  OAI21_X1 U13811 ( .B1(n11266), .B2(n11265), .A(n11264), .ZN(n11267) );
  NAND2_X1 U13812 ( .A1(n11267), .A2(n15345), .ZN(n11273) );
  OAI22_X1 U13813 ( .A1(n13953), .A2(n11269), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n11268), .ZN(n11270) );
  AOI21_X1 U13814 ( .B1(n11271), .B2(n13944), .A(n11270), .ZN(n11272) );
  OAI211_X1 U13815 ( .C1(n11292), .C2(n13958), .A(n11273), .B(n11272), .ZN(
        P2_U3203) );
  OAI21_X1 U13816 ( .B1(n11275), .B2(n15327), .A(n11274), .ZN(n11282) );
  INV_X1 U13817 ( .A(P3_REG0_REG_4__SCAN_IN), .ZN(n11276) );
  OAI22_X1 U13818 ( .A1(n11280), .A2(n13825), .B1(n15775), .B2(n11276), .ZN(
        n11277) );
  AOI21_X1 U13819 ( .B1(n11282), .B2(n15775), .A(n11277), .ZN(n11278) );
  INV_X1 U13820 ( .A(n11278), .ZN(P3_U3402) );
  INV_X1 U13821 ( .A(P3_REG1_REG_4__SCAN_IN), .ZN(n11279) );
  OAI22_X1 U13822 ( .A1(n13777), .A2(n11280), .B1(n15784), .B2(n11279), .ZN(
        n11281) );
  AOI21_X1 U13823 ( .B1(n11282), .B2(n15784), .A(n11281), .ZN(n11283) );
  INV_X1 U13824 ( .A(n11283), .ZN(P3_U3463) );
  INV_X1 U13825 ( .A(n11284), .ZN(n11287) );
  OAI22_X1 U13826 ( .A1(n11285), .A2(P3_U3151), .B1(SI_22_), .B2(n13840), .ZN(
        n11286) );
  AOI21_X1 U13827 ( .B1(n11287), .B2(n13828), .A(n11286), .ZN(P3_U3273) );
  AOI211_X1 U13828 ( .C1(n15366), .C2(n11290), .A(n11289), .B(n11288), .ZN(
        n11296) );
  INV_X1 U13829 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n11291) );
  OAI22_X1 U13830 ( .A1(n14324), .A2(n11292), .B1(n15680), .B2(n11291), .ZN(
        n11293) );
  INV_X1 U13831 ( .A(n11293), .ZN(n11294) );
  OAI21_X1 U13832 ( .B1(n11296), .B2(n15678), .A(n11294), .ZN(P2_U3457) );
  AOI22_X1 U13833 ( .A1(n14313), .A2(n12940), .B1(n7435), .B2(
        P2_REG1_REG_9__SCAN_IN), .ZN(n11295) );
  OAI21_X1 U13834 ( .B1(n11296), .B2(n7435), .A(n11295), .ZN(P2_U3508) );
  XNOR2_X1 U13835 ( .A(n11432), .B(n13254), .ZN(n11470) );
  XNOR2_X1 U13836 ( .A(n11470), .B(n11792), .ZN(n11299) );
  AOI21_X1 U13837 ( .B1(n11300), .B2(n11299), .A(n11612), .ZN(n11306) );
  OAI22_X1 U13838 ( .A1(n13347), .A2(n15753), .B1(n11301), .B2(n13315), .ZN(
        n11302) );
  AOI211_X1 U13839 ( .C1(n13281), .C2(n11751), .A(n11303), .B(n11302), .ZN(
        n11305) );
  NAND2_X1 U13840 ( .A1(n13350), .A2(n11431), .ZN(n11304) );
  OAI211_X1 U13841 ( .C1(n11306), .C2(n13352), .A(n11305), .B(n11304), .ZN(
        P3_U3167) );
  XNOR2_X1 U13842 ( .A(n11308), .B(n11307), .ZN(n11315) );
  NAND2_X1 U13843 ( .A1(n13980), .A2(n13951), .ZN(n11310) );
  NAND2_X1 U13844 ( .A1(n13978), .A2(n13952), .ZN(n11309) );
  AND2_X1 U13845 ( .A1(n11310), .A2(n11309), .ZN(n11370) );
  NAND2_X1 U13846 ( .A1(n13944), .A2(n11379), .ZN(n11312) );
  OAI211_X1 U13847 ( .C1(n11370), .C2(n13953), .A(n11312), .B(n11311), .ZN(
        n11313) );
  AOI21_X1 U13848 ( .B1(n12947), .B2(n15350), .A(n11313), .ZN(n11314) );
  OAI21_X1 U13849 ( .B1(n11315), .B2(n13935), .A(n11314), .ZN(P2_U3189) );
  INV_X1 U13850 ( .A(n12414), .ZN(n12565) );
  OAI222_X1 U13851 ( .A1(P1_U3086), .A2(n12593), .B1(n15238), .B2(n12565), 
        .C1(n11316), .C2(n15239), .ZN(P1_U3336) );
  MUX2_X1 U13852 ( .A(P3_REG2_REG_9__SCAN_IN), .B(P3_REG1_REG_9__SCAN_IN), .S(
        n6945), .Z(n11320) );
  NAND2_X1 U13853 ( .A1(n11320), .A2(n11332), .ZN(n11323) );
  INV_X1 U13854 ( .A(n11458), .ZN(n11325) );
  INV_X1 U13855 ( .A(n11320), .ZN(n11321) );
  NAND2_X1 U13856 ( .A1(n11321), .A2(n11445), .ZN(n11457) );
  AOI21_X1 U13857 ( .B1(n11457), .B2(n11323), .A(n11322), .ZN(n11324) );
  AOI21_X1 U13858 ( .B1(n11325), .B2(n11457), .A(n11324), .ZN(n11329) );
  AOI21_X1 U13859 ( .B1(n15780), .B2(n11327), .A(n11439), .ZN(n11328) );
  OAI22_X1 U13860 ( .A1(n11329), .A2(n15692), .B1(n11328), .B2(n15693), .ZN(
        n11340) );
  INV_X1 U13861 ( .A(P3_REG2_REG_9__SCAN_IN), .ZN(n11334) );
  AOI21_X1 U13862 ( .B1(n11334), .B2(n11333), .A(n11446), .ZN(n11338) );
  NOR2_X1 U13863 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11335), .ZN(n11616) );
  AOI21_X1 U13864 ( .B1(n15698), .B2(P3_ADDR_REG_9__SCAN_IN), .A(n11616), .ZN(
        n11337) );
  NAND2_X1 U13865 ( .A1(n15699), .A2(n11445), .ZN(n11336) );
  OAI211_X1 U13866 ( .C1(n11338), .C2(n15694), .A(n11337), .B(n11336), .ZN(
        n11339) );
  OR2_X1 U13867 ( .A1(n11340), .A2(n11339), .ZN(P3_U3191) );
  NAND2_X1 U13868 ( .A1(n9729), .A2(P3_U3897), .ZN(n11341) );
  OAI21_X1 U13869 ( .B1(P3_U3897), .B2(n11342), .A(n11341), .ZN(P3_U3519) );
  NAND2_X1 U13870 ( .A1(n11343), .A2(n11026), .ZN(n11346) );
  AOI22_X1 U13871 ( .A1(n7282), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n12415), 
        .B2(n11344), .ZN(n11345) );
  NAND2_X1 U13872 ( .A1(n11346), .A2(n11345), .ZN(n12637) );
  INV_X1 U13873 ( .A(n11348), .ZN(n11349) );
  NAND2_X1 U13874 ( .A1(n11351), .A2(n11350), .ZN(n11355) );
  OAI22_X1 U13875 ( .A1(n15511), .A2(n6667), .B1(n11582), .B2(n14557), .ZN(
        n11352) );
  XNOR2_X1 U13876 ( .A(n11352), .B(n6921), .ZN(n11764) );
  AND2_X1 U13877 ( .A1(n14517), .A2(n14702), .ZN(n11353) );
  AOI21_X1 U13878 ( .B1(n12637), .B2(n9893), .A(n11353), .ZN(n11766) );
  XNOR2_X1 U13879 ( .A(n11764), .B(n11766), .ZN(n11354) );
  OAI211_X1 U13880 ( .C1(n11355), .C2(n11354), .A(n11765), .B(n14675), .ZN(
        n11366) );
  NAND2_X1 U13881 ( .A1(n6681), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n11361) );
  NAND2_X1 U13882 ( .A1(n6683), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n11360) );
  OR2_X1 U13883 ( .A1(n11356), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n11357) );
  AND2_X1 U13884 ( .A1(n11402), .A2(n11357), .ZN(n11775) );
  NAND2_X1 U13885 ( .A1(n6677), .A2(n11775), .ZN(n11359) );
  NAND2_X1 U13886 ( .A1(n12519), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n11358) );
  NAND4_X1 U13887 ( .A1(n11361), .A2(n11360), .A3(n11359), .A4(n11358), .ZN(
        n14701) );
  INV_X1 U13888 ( .A(n14701), .ZN(n11821) );
  NAND2_X1 U13889 ( .A1(n14677), .A2(n14703), .ZN(n11363) );
  OAI211_X1 U13890 ( .C1(n11821), .C2(n15384), .A(n11363), .B(n11362), .ZN(
        n11364) );
  AOI21_X1 U13891 ( .B1(n14680), .B2(n11570), .A(n11364), .ZN(n11365) );
  OAI211_X1 U13892 ( .C1(n15511), .C2(n14683), .A(n11366), .B(n11365), .ZN(
        P1_U3213) );
  XOR2_X1 U13893 ( .A(n11367), .B(n13134), .Z(n11377) );
  AOI211_X1 U13894 ( .C1(n12947), .C2(n11368), .A(n6670), .B(n11628), .ZN(
        n11378) );
  OAI211_X1 U13895 ( .C1(n7725), .C2(n8908), .A(n15617), .B(n11369), .ZN(
        n11371) );
  NAND2_X1 U13896 ( .A1(n11371), .A2(n11370), .ZN(n11384) );
  AOI211_X1 U13897 ( .C1(n15366), .C2(n11377), .A(n11378), .B(n11384), .ZN(
        n11376) );
  AOI22_X1 U13898 ( .A1(n14313), .A2(n12947), .B1(n7435), .B2(
        P2_REG1_REG_10__SCAN_IN), .ZN(n11372) );
  OAI21_X1 U13899 ( .B1(n11376), .B2(n7435), .A(n11372), .ZN(P2_U3509) );
  INV_X1 U13900 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n11373) );
  NOR2_X1 U13901 ( .A1(n15680), .A2(n11373), .ZN(n11374) );
  AOI21_X1 U13902 ( .B1(n14375), .B2(n12947), .A(n11374), .ZN(n11375) );
  OAI21_X1 U13903 ( .B1(n11376), .B2(n15678), .A(n11375), .ZN(P2_U3460) );
  INV_X1 U13904 ( .A(n11377), .ZN(n11386) );
  INV_X1 U13905 ( .A(n12947), .ZN(n11382) );
  NAND2_X1 U13906 ( .A1(n11378), .A2(n14160), .ZN(n11381) );
  AOI22_X1 U13907 ( .A1(n15627), .A2(P2_REG2_REG_10__SCAN_IN), .B1(n11379), 
        .B2(n14208), .ZN(n11380) );
  OAI211_X1 U13908 ( .C1(n11382), .C2(n14157), .A(n11381), .B(n11380), .ZN(
        n11383) );
  AOI21_X1 U13909 ( .B1(n11384), .B2(n14226), .A(n11383), .ZN(n11385) );
  OAI21_X1 U13910 ( .B1(n11386), .B2(n14234), .A(n11385), .ZN(P2_U3255) );
  NAND2_X1 U13911 ( .A1(n11388), .A2(n11387), .ZN(n11488) );
  INV_X1 U13912 ( .A(n14704), .ZN(n11583) );
  NAND2_X1 U13913 ( .A1(n11583), .A2(n12629), .ZN(n11390) );
  NAND2_X1 U13914 ( .A1(n14704), .A2(n15505), .ZN(n11389) );
  NAND2_X1 U13915 ( .A1(n11390), .A2(n11389), .ZN(n12800) );
  INV_X1 U13916 ( .A(n12800), .ZN(n11489) );
  NAND2_X1 U13917 ( .A1(n11488), .A2(n11489), .ZN(n11487) );
  NAND2_X1 U13918 ( .A1(n11487), .A2(n11390), .ZN(n11580) );
  NAND2_X1 U13919 ( .A1(n12633), .A2(n11391), .ZN(n11393) );
  OR2_X1 U13920 ( .A1(n11391), .A2(n12633), .ZN(n11392) );
  NAND2_X1 U13921 ( .A1(n11393), .A2(n11392), .ZN(n12803) );
  INV_X1 U13922 ( .A(n12803), .ZN(n11581) );
  NAND2_X1 U13923 ( .A1(n11580), .A2(n11581), .ZN(n11579) );
  NAND2_X1 U13924 ( .A1(n11579), .A2(n11393), .ZN(n11562) );
  XNOR2_X1 U13925 ( .A(n12637), .B(n11582), .ZN(n12801) );
  INV_X1 U13926 ( .A(n12801), .ZN(n11561) );
  NAND2_X1 U13927 ( .A1(n11562), .A2(n11561), .ZN(n11560) );
  NAND2_X1 U13928 ( .A1(n12637), .A2(n11582), .ZN(n11394) );
  NAND2_X1 U13929 ( .A1(n11560), .A2(n11394), .ZN(n11399) );
  NAND2_X1 U13930 ( .A1(n11395), .A2(n11026), .ZN(n11398) );
  AOI22_X1 U13931 ( .A1(n7282), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n12415), 
        .B2(n11396), .ZN(n11397) );
  XNOR2_X1 U13932 ( .A(n12641), .B(n14701), .ZN(n12804) );
  AOI21_X1 U13933 ( .B1(n11399), .B2(n11416), .A(n15481), .ZN(n11409) );
  INV_X1 U13934 ( .A(n11399), .ZN(n11400) );
  NAND2_X1 U13935 ( .A1(n12519), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n11407) );
  NAND2_X1 U13936 ( .A1(n6681), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n11406) );
  NAND2_X1 U13937 ( .A1(n11402), .A2(n11401), .ZN(n11403) );
  AND2_X1 U13938 ( .A1(n11827), .A2(n11403), .ZN(n12074) );
  NAND2_X1 U13939 ( .A1(n6677), .A2(n12074), .ZN(n11405) );
  NAND2_X1 U13940 ( .A1(n6683), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n11404) );
  NAND4_X1 U13941 ( .A1(n11407), .A2(n11406), .A3(n11405), .A4(n11404), .ZN(
        n14700) );
  INV_X1 U13942 ( .A(n14700), .ZN(n12239) );
  OAI22_X1 U13943 ( .A1(n11582), .A2(n15069), .B1(n12239), .B2(n15091), .ZN(
        n11408) );
  AOI21_X1 U13944 ( .B1(n11409), .B2(n11823), .A(n11408), .ZN(n11742) );
  NAND2_X1 U13945 ( .A1(n11529), .A2(n11410), .ZN(n11411) );
  NAND2_X1 U13946 ( .A1(n11583), .A2(n15505), .ZN(n11413) );
  OR2_X1 U13947 ( .A1(n12633), .A2(n14703), .ZN(n11414) );
  OR2_X1 U13948 ( .A1(n12637), .A2(n14702), .ZN(n11415) );
  OAI21_X1 U13949 ( .B1(n11417), .B2(n11416), .A(n11834), .ZN(n11739) );
  INV_X1 U13950 ( .A(n11840), .ZN(n11842) );
  AOI211_X1 U13951 ( .C1(n12641), .C2(n11569), .A(n15488), .B(n11842), .ZN(
        n11740) );
  NAND2_X1 U13952 ( .A1(n11740), .A2(n15293), .ZN(n11419) );
  INV_X1 U13953 ( .A(n15058), .ZN(n15283) );
  AOI22_X1 U13954 ( .A1(n15067), .A2(P1_REG2_REG_8__SCAN_IN), .B1(n11775), 
        .B2(n15283), .ZN(n11418) );
  OAI211_X1 U13955 ( .C1(n7186), .C2(n15013), .A(n11419), .B(n11418), .ZN(
        n11420) );
  AOI21_X1 U13956 ( .B1(n11739), .B2(n15294), .A(n11420), .ZN(n11421) );
  OAI21_X1 U13957 ( .B1(n11742), .B2(n15067), .A(n11421), .ZN(P1_U3285) );
  INV_X1 U13958 ( .A(n11422), .ZN(n11423) );
  AOI21_X1 U13959 ( .B1(n11426), .B2(n11424), .A(n11423), .ZN(n11430) );
  AOI22_X1 U13960 ( .A1(n11751), .A2(n15719), .B1(n15717), .B2(n11425), .ZN(
        n11429) );
  XNOR2_X1 U13961 ( .A(n11427), .B(n11426), .ZN(n15752) );
  NAND2_X1 U13962 ( .A1(n15752), .A2(n13554), .ZN(n11428) );
  OAI211_X1 U13963 ( .C1(n11430), .C2(n13691), .A(n11429), .B(n11428), .ZN(
        n15756) );
  INV_X1 U13964 ( .A(n15756), .ZN(n11437) );
  AOI22_X1 U13965 ( .A1(n15707), .A2(n11432), .B1(n15709), .B2(n11431), .ZN(
        n11433) );
  OAI21_X1 U13966 ( .B1(n11434), .B2(n15733), .A(n11433), .ZN(n11435) );
  AOI21_X1 U13967 ( .B1(n15752), .B2(n13561), .A(n11435), .ZN(n11436) );
  OAI21_X1 U13968 ( .B1(n11437), .B2(n15735), .A(n11436), .ZN(P3_U3228) );
  NOR2_X1 U13969 ( .A1(n11445), .A2(n11438), .ZN(n11440) );
  NAND2_X1 U13970 ( .A1(P3_REG1_REG_10__SCAN_IN), .A2(n11914), .ZN(n11441) );
  OAI21_X1 U13971 ( .B1(P3_REG1_REG_10__SCAN_IN), .B2(n11914), .A(n11441), 
        .ZN(n11442) );
  AOI21_X1 U13972 ( .B1(n11443), .B2(n11442), .A(n11913), .ZN(n11469) );
  NOR2_X1 U13973 ( .A1(n11445), .A2(n11444), .ZN(n11447) );
  NAND2_X1 U13974 ( .A1(P3_REG2_REG_10__SCAN_IN), .A2(n11914), .ZN(n11448) );
  OAI21_X1 U13975 ( .B1(P3_REG2_REG_10__SCAN_IN), .B2(n11914), .A(n11448), 
        .ZN(n11449) );
  AOI21_X1 U13976 ( .B1(n11450), .B2(n11449), .A(n11900), .ZN(n11466) );
  INV_X1 U13977 ( .A(P3_REG2_REG_10__SCAN_IN), .ZN(n11452) );
  MUX2_X1 U13978 ( .A(n11452), .B(n11451), .S(n6945), .Z(n11453) );
  NAND2_X1 U13979 ( .A1(n11453), .A2(n11463), .ZN(n11905) );
  INV_X1 U13980 ( .A(n11453), .ZN(n11454) );
  NAND2_X1 U13981 ( .A1(n11454), .A2(n11914), .ZN(n11455) );
  NAND2_X1 U13982 ( .A1(n11905), .A2(n11455), .ZN(n11456) );
  AOI21_X1 U13983 ( .B1(n11458), .B2(n11457), .A(n11456), .ZN(n11907) );
  AND3_X1 U13984 ( .A1(n11458), .A2(n11457), .A3(n11456), .ZN(n11459) );
  OAI21_X1 U13985 ( .B1(n11907), .B2(n11459), .A(n13529), .ZN(n11465) );
  INV_X1 U13986 ( .A(P3_REG3_REG_10__SCAN_IN), .ZN(n11460) );
  NOR2_X1 U13987 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11460), .ZN(n11867) );
  NOR2_X1 U13988 ( .A1(n13492), .A2(n11461), .ZN(n11462) );
  AOI211_X1 U13989 ( .C1(n15699), .C2(n11463), .A(n11867), .B(n11462), .ZN(
        n11464) );
  OAI211_X1 U13990 ( .C1(n11466), .C2(n15694), .A(n11465), .B(n11464), .ZN(
        n11467) );
  INV_X1 U13991 ( .A(n11467), .ZN(n11468) );
  OAI21_X1 U13992 ( .B1(n11469), .B2(n15693), .A(n11468), .ZN(P3_U3192) );
  INV_X1 U13993 ( .A(n15710), .ZN(n11479) );
  NAND2_X1 U13994 ( .A1(n11470), .A2(n11792), .ZN(n11604) );
  INV_X1 U13995 ( .A(n11604), .ZN(n11471) );
  NOR2_X1 U13996 ( .A1(n11612), .A2(n11471), .ZN(n11473) );
  XNOR2_X1 U13997 ( .A(n15708), .B(n13207), .ZN(n11605) );
  XNOR2_X1 U13998 ( .A(n11602), .B(n11605), .ZN(n11472) );
  NAND2_X1 U13999 ( .A1(n11473), .A2(n11472), .ZN(n11637) );
  OAI211_X1 U14000 ( .C1(n11473), .C2(n11472), .A(n11637), .B(n13322), .ZN(
        n11477) );
  OAI22_X1 U14001 ( .A1(n13347), .A2(n11799), .B1(n11792), .B2(n13315), .ZN(
        n11474) );
  AOI211_X1 U14002 ( .C1(n13281), .C2(n12017), .A(n11475), .B(n11474), .ZN(
        n11476) );
  OAI211_X1 U14003 ( .C1(n11479), .C2(n11478), .A(n11477), .B(n11476), .ZN(
        P3_U3179) );
  NAND2_X1 U14004 ( .A1(n15048), .A2(n12592), .ZN(n12785) );
  OR2_X1 U14005 ( .A1(n11480), .A2(n12800), .ZN(n11481) );
  NAND2_X1 U14006 ( .A1(n11482), .A2(n11481), .ZN(n15503) );
  AOI21_X1 U14007 ( .B1(n11483), .B2(n12629), .A(n15488), .ZN(n11484) );
  NAND2_X1 U14008 ( .A1(n11484), .A2(n11590), .ZN(n15504) );
  AOI22_X1 U14009 ( .A1(n15285), .A2(n12629), .B1(n11485), .B2(n15283), .ZN(
        n11486) );
  OAI21_X1 U14010 ( .B1(n15504), .B2(n14994), .A(n11486), .ZN(n11497) );
  OAI21_X1 U14011 ( .B1(n11489), .B2(n11488), .A(n11487), .ZN(n11493) );
  NAND2_X1 U14012 ( .A1(n14705), .A2(n15001), .ZN(n11491) );
  NAND2_X1 U14013 ( .A1(n14703), .A2(n15002), .ZN(n11490) );
  NAND2_X1 U14014 ( .A1(n11491), .A2(n11490), .ZN(n11492) );
  AOI21_X1 U14015 ( .B1(n11493), .B2(n15280), .A(n11492), .ZN(n11495) );
  NAND2_X1 U14016 ( .A1(n15503), .A2(n15080), .ZN(n11494) );
  NAND2_X1 U14017 ( .A1(n11495), .A2(n11494), .ZN(n15508) );
  MUX2_X1 U14018 ( .A(P1_REG2_REG_5__SCAN_IN), .B(n15508), .S(n15093), .Z(
        n11496) );
  AOI211_X1 U14019 ( .C1(n15086), .C2(n15503), .A(n11497), .B(n11496), .ZN(
        n11498) );
  INV_X1 U14020 ( .A(n11498), .ZN(P1_U3288) );
  NAND2_X1 U14021 ( .A1(n14134), .A2(n11499), .ZN(n11506) );
  INV_X1 U14022 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n11500) );
  OAI22_X1 U14023 ( .A1(n14226), .A2(n10086), .B1(n11500), .B2(n15621), .ZN(
        n11503) );
  NOR2_X1 U14024 ( .A1(n14157), .A2(n11501), .ZN(n11502) );
  AOI211_X1 U14025 ( .C1(n11504), .C2(n14160), .A(n11503), .B(n11502), .ZN(
        n11505) );
  OAI211_X1 U14026 ( .C1(n15627), .C2(n11507), .A(n11506), .B(n11505), .ZN(
        P2_U3263) );
  XNOR2_X1 U14027 ( .A(n13126), .B(n11508), .ZN(n15664) );
  OAI211_X1 U14028 ( .C1(n11511), .C2(n11510), .A(n11509), .B(n14206), .ZN(
        n15661) );
  AOI22_X1 U14029 ( .A1(n14228), .A2(n15659), .B1(n14208), .B2(n11512), .ZN(
        n11513) );
  OAI21_X1 U14030 ( .B1(n14213), .B2(n15661), .A(n11513), .ZN(n11514) );
  AOI21_X1 U14031 ( .B1(n14134), .B2(n15664), .A(n11514), .ZN(n11523) );
  OR2_X1 U14032 ( .A1(n11516), .A2(n11515), .ZN(n11517) );
  NAND2_X1 U14033 ( .A1(n11518), .A2(n11517), .ZN(n11520) );
  AOI21_X1 U14034 ( .B1(n11520), .B2(n15617), .A(n11519), .ZN(n15668) );
  MUX2_X1 U14035 ( .A(n15668), .B(n11521), .S(n15627), .Z(n11522) );
  NAND2_X1 U14036 ( .A1(n11523), .A2(n11522), .ZN(P2_U3261) );
  OAI21_X1 U14037 ( .B1(n11525), .B2(n7055), .A(n11524), .ZN(n11526) );
  INV_X1 U14038 ( .A(n11526), .ZN(n15500) );
  INV_X1 U14039 ( .A(n15086), .ZN(n11596) );
  OAI21_X1 U14040 ( .B1(n12616), .B2(n11528), .A(n11527), .ZN(n11532) );
  OAI22_X1 U14041 ( .A1(n10688), .A2(n15069), .B1(n11529), .B2(n15091), .ZN(
        n11531) );
  NOR2_X1 U14042 ( .A1(n15500), .A2(n11584), .ZN(n11530) );
  AOI211_X1 U14043 ( .C1(n15280), .C2(n11532), .A(n11531), .B(n11530), .ZN(
        n15498) );
  MUX2_X1 U14044 ( .A(n11533), .B(n15498), .S(n15093), .Z(n11541) );
  INV_X1 U14045 ( .A(n11534), .ZN(n11537) );
  INV_X1 U14046 ( .A(n11535), .ZN(n11536) );
  AOI211_X1 U14047 ( .C1(n15496), .C2(n11537), .A(n15488), .B(n11536), .ZN(
        n15494) );
  OAI22_X1 U14048 ( .A1(n15013), .A2(n11538), .B1(P1_REG3_REG_3__SCAN_IN), 
        .B2(n15058), .ZN(n11539) );
  AOI21_X1 U14049 ( .B1(n15494), .B2(n15293), .A(n11539), .ZN(n11540) );
  OAI211_X1 U14050 ( .C1(n15500), .C2(n11596), .A(n11541), .B(n11540), .ZN(
        P1_U3290) );
  MUX2_X1 U14051 ( .A(n11542), .B(P1_REG2_REG_2__SCAN_IN), .S(n15067), .Z(
        n11543) );
  INV_X1 U14052 ( .A(n11543), .ZN(n11548) );
  OAI22_X1 U14053 ( .A1(n15013), .A2(n11544), .B1(n15058), .B2(n14726), .ZN(
        n11545) );
  AOI21_X1 U14054 ( .B1(n15293), .B2(n11546), .A(n11545), .ZN(n11547) );
  OAI211_X1 U14055 ( .C1(n11549), .C2(n11596), .A(n11548), .B(n11547), .ZN(
        P1_U3291) );
  INV_X1 U14056 ( .A(n11550), .ZN(n11553) );
  AOI22_X1 U14057 ( .A1(n14228), .A2(n12924), .B1(n11551), .B2(n14208), .ZN(
        n11552) );
  OAI21_X1 U14058 ( .B1(n11553), .B2(n14213), .A(n11552), .ZN(n11556) );
  MUX2_X1 U14059 ( .A(P2_REG2_REG_7__SCAN_IN), .B(n11554), .S(n14226), .Z(
        n11555) );
  AOI211_X1 U14060 ( .C1(n14134), .C2(n11557), .A(n11556), .B(n11555), .ZN(
        n11558) );
  INV_X1 U14061 ( .A(n11558), .ZN(P2_U3258) );
  XNOR2_X1 U14062 ( .A(n11559), .B(n12801), .ZN(n15513) );
  NAND2_X1 U14063 ( .A1(n15513), .A2(n15080), .ZN(n11568) );
  OAI21_X1 U14064 ( .B1(n11562), .B2(n11561), .A(n11560), .ZN(n11566) );
  NAND2_X1 U14065 ( .A1(n14703), .A2(n15001), .ZN(n11564) );
  NAND2_X1 U14066 ( .A1(n14701), .A2(n15002), .ZN(n11563) );
  NAND2_X1 U14067 ( .A1(n11564), .A2(n11563), .ZN(n11565) );
  AOI21_X1 U14068 ( .B1(n11566), .B2(n15280), .A(n11565), .ZN(n11567) );
  AND2_X1 U14069 ( .A1(n11568), .A2(n11567), .ZN(n15515) );
  OAI211_X1 U14070 ( .C1(n11589), .C2(n15511), .A(n15291), .B(n11569), .ZN(
        n15510) );
  INV_X1 U14071 ( .A(n11570), .ZN(n11571) );
  OAI22_X1 U14072 ( .A1(n15093), .A2(n10204), .B1(n11571), .B2(n15058), .ZN(
        n11572) );
  AOI21_X1 U14073 ( .B1(n15285), .B2(n12637), .A(n11572), .ZN(n11573) );
  OAI21_X1 U14074 ( .B1(n15510), .B2(n14994), .A(n11573), .ZN(n11574) );
  AOI21_X1 U14075 ( .B1(n15513), .B2(n15086), .A(n11574), .ZN(n11575) );
  OAI21_X1 U14076 ( .B1(n15515), .B2(n15067), .A(n11575), .ZN(P1_U3286) );
  OAI21_X1 U14077 ( .B1(n11577), .B2(n12803), .A(n11576), .ZN(n11578) );
  INV_X1 U14078 ( .A(n11578), .ZN(n11647) );
  OAI21_X1 U14079 ( .B1(n11581), .B2(n11580), .A(n11579), .ZN(n11587) );
  OAI22_X1 U14080 ( .A1(n11583), .A2(n15069), .B1(n11582), .B2(n15091), .ZN(
        n11586) );
  NOR2_X1 U14081 ( .A1(n11647), .A2(n11584), .ZN(n11585) );
  AOI211_X1 U14082 ( .C1(n15280), .C2(n11587), .A(n11586), .B(n11585), .ZN(
        n11646) );
  MUX2_X1 U14083 ( .A(n11588), .B(n11646), .S(n15093), .Z(n11595) );
  AOI211_X1 U14084 ( .C1(n12633), .C2(n11590), .A(n15488), .B(n11589), .ZN(
        n11644) );
  OAI22_X1 U14085 ( .A1(n15013), .A2(n11592), .B1(n15058), .B2(n11591), .ZN(
        n11593) );
  AOI21_X1 U14086 ( .B1(n11644), .B2(n15293), .A(n11593), .ZN(n11594) );
  OAI211_X1 U14087 ( .C1(n11647), .C2(n11596), .A(n11595), .B(n11594), .ZN(
        P1_U3287) );
  NAND2_X1 U14088 ( .A1(n11597), .A2(n13828), .ZN(n11599) );
  OAI211_X1 U14089 ( .C1(n11600), .C2(n13840), .A(n11599), .B(n11598), .ZN(
        P3_U3272) );
  XNOR2_X1 U14090 ( .A(n15759), .B(n13254), .ZN(n11862) );
  XNOR2_X1 U14091 ( .A(n11862), .B(n12018), .ZN(n11614) );
  XNOR2_X1 U14092 ( .A(n12173), .B(n13254), .ZN(n11608) );
  XNOR2_X1 U14093 ( .A(n11608), .B(n13357), .ZN(n11607) );
  INV_X1 U14094 ( .A(n11607), .ZN(n11852) );
  INV_X1 U14095 ( .A(n11605), .ZN(n11601) );
  NAND2_X1 U14096 ( .A1(n11602), .A2(n11601), .ZN(n11603) );
  NAND2_X1 U14097 ( .A1(n11751), .A2(n11605), .ZN(n11636) );
  OAI21_X1 U14098 ( .B1(n11607), .B2(n11636), .A(n11850), .ZN(n11610) );
  INV_X1 U14099 ( .A(n11850), .ZN(n11606) );
  OAI21_X1 U14100 ( .B1(n11607), .B2(n11858), .A(n11606), .ZN(n11609) );
  AOI22_X1 U14101 ( .A1(n11610), .A2(n11609), .B1(n11608), .B2(n13357), .ZN(
        n11611) );
  AOI21_X1 U14102 ( .B1(n11614), .B2(n11613), .A(n11864), .ZN(n11619) );
  OAI22_X1 U14103 ( .A1(n13347), .A2(n15759), .B1(n11640), .B2(n13315), .ZN(
        n11615) );
  AOI211_X1 U14104 ( .C1(n13281), .C2(n12145), .A(n11616), .B(n11615), .ZN(
        n11618) );
  NAND2_X1 U14105 ( .A1(n13350), .A2(n12038), .ZN(n11617) );
  OAI211_X1 U14106 ( .C1(n11619), .C2(n13352), .A(n11618), .B(n11617), .ZN(
        P3_U3171) );
  XOR2_X1 U14107 ( .A(n13135), .B(n11620), .Z(n11781) );
  INV_X1 U14108 ( .A(n11781), .ZN(n11635) );
  INV_X1 U14109 ( .A(n11621), .ZN(n11622) );
  AOI21_X1 U14110 ( .B1(n13135), .B2(n11623), .A(n11622), .ZN(n11627) );
  NAND2_X1 U14111 ( .A1(n13977), .A2(n12105), .ZN(n11625) );
  NAND2_X1 U14112 ( .A1(n13979), .A2(n13951), .ZN(n11624) );
  NAND2_X1 U14113 ( .A1(n11625), .A2(n11624), .ZN(n15348) );
  INV_X1 U14114 ( .A(n15348), .ZN(n11626) );
  OAI21_X1 U14115 ( .B1(n11627), .B2(n14220), .A(n11626), .ZN(n11779) );
  NAND2_X1 U14116 ( .A1(n11779), .A2(n14226), .ZN(n11634) );
  INV_X1 U14117 ( .A(n11628), .ZN(n11629) );
  AOI211_X1 U14118 ( .C1(n15349), .C2(n11629), .A(n6670), .B(n11713), .ZN(
        n11780) );
  AOI22_X1 U14119 ( .A1(n15627), .A2(P2_REG2_REG_11__SCAN_IN), .B1(n11630), 
        .B2(n14208), .ZN(n11631) );
  OAI21_X1 U14120 ( .B1(n11783), .B2(n14157), .A(n11631), .ZN(n11632) );
  AOI21_X1 U14121 ( .B1(n11780), .B2(n14160), .A(n11632), .ZN(n11633) );
  OAI211_X1 U14122 ( .C1(n14234), .C2(n11635), .A(n11634), .B(n11633), .ZN(
        P2_U3254) );
  NAND2_X1 U14123 ( .A1(n11637), .A2(n11636), .ZN(n11851) );
  XNOR2_X1 U14124 ( .A(n11851), .B(n11850), .ZN(n11643) );
  AOI22_X1 U14125 ( .A1(n11751), .A2(n13343), .B1(n11896), .B2(n13337), .ZN(
        n11639) );
  OAI211_X1 U14126 ( .C1(n11640), .C2(n13346), .A(n11639), .B(n11638), .ZN(
        n11641) );
  AOI21_X1 U14127 ( .B1(n11757), .B2(n13350), .A(n11641), .ZN(n11642) );
  OAI21_X1 U14128 ( .B1(n11643), .B2(n13352), .A(n11642), .ZN(P3_U3153) );
  INV_X1 U14129 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n11649) );
  AOI21_X1 U14130 ( .B1(n12633), .B2(n15495), .A(n11644), .ZN(n11645) );
  OAI211_X1 U14131 ( .C1(n11647), .C2(n15499), .A(n11646), .B(n11645), .ZN(
        n11650) );
  NAND2_X1 U14132 ( .A1(n11650), .A2(n15526), .ZN(n11648) );
  OAI21_X1 U14133 ( .B1(n15526), .B2(n11649), .A(n11648), .ZN(P1_U3477) );
  NAND2_X1 U14134 ( .A1(n11650), .A2(n15537), .ZN(n11651) );
  OAI21_X1 U14135 ( .B1(n15537), .B2(n11652), .A(n11651), .ZN(P1_U3534) );
  OAI211_X1 U14136 ( .C1(n8887), .C2(n15616), .A(n14206), .B(n11653), .ZN(
        n15643) );
  XNOR2_X1 U14137 ( .A(n11655), .B(n13121), .ZN(n15641) );
  XNOR2_X1 U14138 ( .A(n13121), .B(n13120), .ZN(n11657) );
  OAI21_X1 U14139 ( .B1(n11657), .B2(n14220), .A(n11656), .ZN(n15646) );
  AOI22_X1 U14140 ( .A1(n14134), .A2(n15641), .B1(n14226), .B2(n15646), .ZN(
        n11662) );
  INV_X1 U14141 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n11659) );
  OAI22_X1 U14142 ( .A1(n14226), .A2(n11659), .B1(n11658), .B2(n15621), .ZN(
        n11660) );
  AOI21_X1 U14143 ( .B1(n14228), .B2(n8886), .A(n11660), .ZN(n11661) );
  OAI211_X1 U14144 ( .C1(n14213), .C2(n15643), .A(n11662), .B(n11661), .ZN(
        P2_U3264) );
  NAND2_X1 U14145 ( .A1(n11696), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n11876) );
  INV_X1 U14146 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n11663) );
  NAND2_X1 U14147 ( .A1(n11884), .A2(n11663), .ZN(n11664) );
  AND2_X1 U14148 ( .A1(n11876), .A2(n11664), .ZN(n11676) );
  INV_X1 U14149 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n12208) );
  OR2_X1 U14150 ( .A1(n11690), .A2(n12208), .ZN(n11674) );
  XNOR2_X1 U14151 ( .A(n11690), .B(P2_REG2_REG_16__SCAN_IN), .ZN(n15606) );
  NAND2_X1 U14152 ( .A1(n15568), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n11668) );
  INV_X1 U14153 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n11665) );
  MUX2_X1 U14154 ( .A(n11665), .B(P2_REG2_REG_13__SCAN_IN), .S(n15568), .Z(
        n11666) );
  INV_X1 U14155 ( .A(n11666), .ZN(n15570) );
  INV_X1 U14156 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n11667) );
  OR2_X1 U14157 ( .A1(n11679), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n15557) );
  MUX2_X1 U14158 ( .A(n11667), .B(P2_REG2_REG_12__SCAN_IN), .S(n15555), .Z(
        n15558) );
  AOI21_X1 U14159 ( .B1(n15559), .B2(n15557), .A(n15558), .ZN(n15561) );
  AOI21_X1 U14160 ( .B1(n11667), .B2(n11684), .A(n15561), .ZN(n15571) );
  NAND2_X1 U14161 ( .A1(n15570), .A2(n15571), .ZN(n15569) );
  NAND2_X1 U14162 ( .A1(n11668), .A2(n15569), .ZN(n11670) );
  NAND2_X1 U14163 ( .A1(n11669), .A2(n11670), .ZN(n11671) );
  XNOR2_X1 U14164 ( .A(n11670), .B(n15580), .ZN(n15584) );
  NAND2_X1 U14165 ( .A1(P2_REG2_REG_14__SCAN_IN), .A2(n15584), .ZN(n15583) );
  NAND2_X1 U14166 ( .A1(n11671), .A2(n15583), .ZN(n11672) );
  NAND2_X1 U14167 ( .A1(n15592), .A2(n11672), .ZN(n11673) );
  XOR2_X1 U14168 ( .A(n15592), .B(n11672), .Z(n15594) );
  NAND2_X1 U14169 ( .A1(P2_REG2_REG_15__SCAN_IN), .A2(n15594), .ZN(n15593) );
  NAND2_X1 U14170 ( .A1(n11673), .A2(n15593), .ZN(n15607) );
  NAND2_X1 U14171 ( .A1(n15606), .A2(n15607), .ZN(n15605) );
  NAND2_X1 U14172 ( .A1(n11674), .A2(n15605), .ZN(n11675) );
  NAND2_X1 U14173 ( .A1(n11676), .A2(n11675), .ZN(n11875) );
  OAI211_X1 U14174 ( .C1(n11676), .C2(n11675), .A(n15604), .B(n11875), .ZN(
        n11678) );
  NAND2_X1 U14175 ( .A1(P2_U3088), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n13901)
         );
  NAND2_X1 U14176 ( .A1(n15601), .A2(P2_ADDR_REG_17__SCAN_IN), .ZN(n11677) );
  NAND3_X1 U14177 ( .A1(n11678), .A2(n13901), .A3(n11677), .ZN(n11695) );
  AOI22_X1 U14178 ( .A1(P2_REG1_REG_17__SCAN_IN), .A2(n11696), .B1(n11884), 
        .B2(n14308), .ZN(n11692) );
  INV_X1 U14179 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n14312) );
  XNOR2_X1 U14180 ( .A(n11690), .B(P2_REG1_REG_16__SCAN_IN), .ZN(n15610) );
  INV_X1 U14181 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n11686) );
  XNOR2_X1 U14182 ( .A(n15580), .B(P2_REG1_REG_14__SCAN_IN), .ZN(n15587) );
  INV_X1 U14183 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n15361) );
  INV_X1 U14184 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n15551) );
  NAND2_X1 U14185 ( .A1(n11679), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n11680) );
  NAND2_X1 U14186 ( .A1(n11681), .A2(n11680), .ZN(n15550) );
  MUX2_X1 U14187 ( .A(n15551), .B(P2_REG1_REG_12__SCAN_IN), .S(n15555), .Z(
        n11682) );
  OR2_X1 U14188 ( .A1(n15550), .A2(n11682), .ZN(n15552) );
  INV_X1 U14189 ( .A(n15552), .ZN(n11683) );
  AOI21_X1 U14190 ( .B1(n15551), .B2(n11684), .A(n11683), .ZN(n15574) );
  MUX2_X1 U14191 ( .A(P2_REG1_REG_13__SCAN_IN), .B(n15361), .S(n15568), .Z(
        n15573) );
  NAND2_X1 U14192 ( .A1(n15574), .A2(n15573), .ZN(n15572) );
  OAI21_X1 U14193 ( .B1(n11685), .B2(n15361), .A(n15572), .ZN(n15586) );
  NAND2_X1 U14194 ( .A1(n15587), .A2(n15586), .ZN(n15585) );
  OAI21_X1 U14195 ( .B1(n15580), .B2(n11686), .A(n15585), .ZN(n11687) );
  NAND2_X1 U14196 ( .A1(n15592), .A2(n11687), .ZN(n11689) );
  XNOR2_X1 U14197 ( .A(n11688), .B(n11687), .ZN(n15596) );
  NAND2_X1 U14198 ( .A1(P2_REG1_REG_15__SCAN_IN), .A2(n15596), .ZN(n15595) );
  NAND2_X1 U14199 ( .A1(n11689), .A2(n15595), .ZN(n15611) );
  NAND2_X1 U14200 ( .A1(n15610), .A2(n15611), .ZN(n15608) );
  OAI21_X1 U14201 ( .B1(n11690), .B2(n14312), .A(n15608), .ZN(n11691) );
  NAND2_X1 U14202 ( .A1(n11692), .A2(n11691), .ZN(n11883) );
  OAI21_X1 U14203 ( .B1(n11692), .B2(n11691), .A(n11883), .ZN(n11693) );
  NOR2_X1 U14204 ( .A1(n11693), .A2(n14009), .ZN(n11694) );
  AOI211_X1 U14205 ( .C1(n15603), .C2(n11696), .A(n11695), .B(n11694), .ZN(
        n11697) );
  INV_X1 U14206 ( .A(n11697), .ZN(P2_U3231) );
  NAND2_X1 U14207 ( .A1(n7733), .A2(n11699), .ZN(n11700) );
  XNOR2_X1 U14208 ( .A(n11698), .B(n11700), .ZN(n11707) );
  INV_X1 U14209 ( .A(n11714), .ZN(n11704) );
  NAND2_X1 U14210 ( .A1(n13976), .A2(n12105), .ZN(n11702) );
  NAND2_X1 U14211 ( .A1(n13978), .A2(n13951), .ZN(n11701) );
  NAND2_X1 U14212 ( .A1(n11702), .A2(n11701), .ZN(n11709) );
  AOI22_X1 U14213 ( .A1(n15347), .A2(n11709), .B1(P2_REG3_REG_12__SCAN_IN), 
        .B2(P2_U3088), .ZN(n11703) );
  OAI21_X1 U14214 ( .B1(n11704), .B2(n15354), .A(n11703), .ZN(n11705) );
  AOI21_X1 U14215 ( .B1(n12959), .B2(n15350), .A(n11705), .ZN(n11706) );
  OAI21_X1 U14216 ( .B1(n11707), .B2(n13935), .A(n11706), .ZN(P2_U3196) );
  XOR2_X1 U14217 ( .A(n11708), .B(n13136), .Z(n11711) );
  INV_X1 U14218 ( .A(n11709), .ZN(n11710) );
  OAI21_X1 U14219 ( .B1(n11711), .B2(n14220), .A(n11710), .ZN(n15364) );
  INV_X1 U14220 ( .A(n15364), .ZN(n11719) );
  XOR2_X1 U14221 ( .A(n13136), .B(n11712), .Z(n15367) );
  OAI211_X1 U14222 ( .C1(n11713), .C2(n15363), .A(n14206), .B(n11811), .ZN(
        n15362) );
  AOI22_X1 U14223 ( .A1(n15627), .A2(P2_REG2_REG_12__SCAN_IN), .B1(n11714), 
        .B2(n14208), .ZN(n11716) );
  NAND2_X1 U14224 ( .A1(n12959), .A2(n14228), .ZN(n11715) );
  OAI211_X1 U14225 ( .C1(n15362), .C2(n14213), .A(n11716), .B(n11715), .ZN(
        n11717) );
  AOI21_X1 U14226 ( .B1(n15367), .B2(n14134), .A(n11717), .ZN(n11718) );
  OAI21_X1 U14227 ( .B1(n11719), .B2(n15627), .A(n11718), .ZN(P2_U3253) );
  NAND2_X1 U14228 ( .A1(n12333), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n11721) );
  NAND2_X1 U14229 ( .A1(n11721), .A2(n11720), .ZN(n11722) );
  INV_X1 U14230 ( .A(n11722), .ZN(n11723) );
  XNOR2_X1 U14231 ( .A(n11722), .B(n12346), .ZN(n15464) );
  NOR2_X1 U14232 ( .A1(P1_REG2_REG_15__SCAN_IN), .A2(n15464), .ZN(n15463) );
  AOI21_X1 U14233 ( .B1(n11723), .B2(n15471), .A(n15463), .ZN(n11726) );
  INV_X1 U14234 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n11724) );
  MUX2_X1 U14235 ( .A(P1_REG2_REG_16__SCAN_IN), .B(n11724), .S(n12395), .Z(
        n11725) );
  NAND2_X1 U14236 ( .A1(n11725), .A2(n11726), .ZN(n11925) );
  OAI211_X1 U14237 ( .C1(n11726), .C2(n11725), .A(n14838), .B(n11925), .ZN(
        n11737) );
  NAND2_X1 U14238 ( .A1(P1_U3086), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n14597)
         );
  AOI21_X1 U14239 ( .B1(n11729), .B2(n11728), .A(n11727), .ZN(n11730) );
  INV_X1 U14240 ( .A(n11730), .ZN(n11731) );
  XNOR2_X1 U14241 ( .A(n11730), .B(n12346), .ZN(n15466) );
  NOR2_X1 U14242 ( .A1(P1_REG1_REG_15__SCAN_IN), .A2(n15466), .ZN(n15465) );
  AOI21_X1 U14243 ( .B1(n15471), .B2(n11731), .A(n15465), .ZN(n11733) );
  XOR2_X1 U14244 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n12395), .Z(n11732) );
  NAND2_X1 U14245 ( .A1(n11732), .A2(n11733), .ZN(n11920) );
  OAI211_X1 U14246 ( .C1(n11733), .C2(n11732), .A(n14833), .B(n11920), .ZN(
        n11734) );
  NAND2_X1 U14247 ( .A1(n14597), .A2(n11734), .ZN(n11735) );
  AOI21_X1 U14248 ( .B1(n14819), .B2(P1_ADDR_REG_16__SCAN_IN), .A(n11735), 
        .ZN(n11736) );
  OAI211_X1 U14249 ( .C1(n15472), .C2(n11738), .A(n11737), .B(n11736), .ZN(
        P1_U3259) );
  INV_X1 U14250 ( .A(n11739), .ZN(n11743) );
  AOI21_X1 U14251 ( .B1(n12641), .B2(n15495), .A(n11740), .ZN(n11741) );
  OAI211_X1 U14252 ( .C1(n11743), .C2(n15482), .A(n11742), .B(n11741), .ZN(
        n11745) );
  NAND2_X1 U14253 ( .A1(n11745), .A2(n15537), .ZN(n11744) );
  OAI21_X1 U14254 ( .B1(n15537), .B2(n10167), .A(n11744), .ZN(P1_U3536) );
  INV_X1 U14255 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n11747) );
  NAND2_X1 U14256 ( .A1(n11745), .A2(n15526), .ZN(n11746) );
  OAI21_X1 U14257 ( .B1(n15526), .B2(n11747), .A(n11746), .ZN(P1_U3483) );
  NAND2_X1 U14258 ( .A1(n11794), .A2(n11748), .ZN(n11750) );
  NAND2_X1 U14259 ( .A1(n11750), .A2(n11749), .ZN(n11999) );
  OAI211_X1 U14260 ( .C1(n11750), .C2(n11749), .A(n11999), .B(n15722), .ZN(
        n11753) );
  AOI22_X1 U14261 ( .A1(n11751), .A2(n15717), .B1(n15719), .B2(n13357), .ZN(
        n11752) );
  NAND2_X1 U14262 ( .A1(n11753), .A2(n11752), .ZN(n11890) );
  INV_X1 U14263 ( .A(n11890), .ZN(n11762) );
  OAI21_X1 U14264 ( .B1(n11756), .B2(n11755), .A(n11754), .ZN(n11891) );
  AOI22_X1 U14265 ( .A1(n15707), .A2(n11896), .B1(n15709), .B2(n11757), .ZN(
        n11758) );
  OAI21_X1 U14266 ( .B1(n11759), .B2(n15733), .A(n11758), .ZN(n11760) );
  AOI21_X1 U14267 ( .B1(n11891), .B2(n13716), .A(n11760), .ZN(n11761) );
  OAI21_X1 U14268 ( .B1(n11762), .B2(n15735), .A(n11761), .ZN(P3_U3226) );
  AOI22_X1 U14269 ( .A1(n12641), .A2(n14511), .B1(n9893), .B2(n14701), .ZN(
        n11763) );
  XNOR2_X1 U14270 ( .A(n11763), .B(n14445), .ZN(n12065) );
  AOI22_X1 U14271 ( .A1(n12641), .A2(n9893), .B1(n14517), .B2(n14701), .ZN(
        n12066) );
  XNOR2_X1 U14272 ( .A(n12065), .B(n12066), .ZN(n11771) );
  INV_X1 U14273 ( .A(n12068), .ZN(n11769) );
  AOI21_X1 U14274 ( .B1(n11771), .B2(n11770), .A(n11769), .ZN(n11778) );
  NAND2_X1 U14275 ( .A1(n14677), .A2(n14702), .ZN(n11773) );
  OAI211_X1 U14276 ( .C1(n12239), .C2(n15384), .A(n11773), .B(n11772), .ZN(
        n11774) );
  AOI21_X1 U14277 ( .B1(n14680), .B2(n11775), .A(n11774), .ZN(n11777) );
  NAND2_X1 U14278 ( .A1(n15397), .A2(n12641), .ZN(n11776) );
  OAI211_X1 U14279 ( .C1(n11778), .C2(n15392), .A(n11777), .B(n11776), .ZN(
        P1_U3221) );
  AOI211_X1 U14280 ( .C1(n15366), .C2(n11781), .A(n11780), .B(n11779), .ZN(
        n11787) );
  INV_X1 U14281 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n11782) );
  OAI22_X1 U14282 ( .A1(n11783), .A2(n14324), .B1(n15680), .B2(n11782), .ZN(
        n11784) );
  INV_X1 U14283 ( .A(n11784), .ZN(n11785) );
  OAI21_X1 U14284 ( .B1(n11787), .B2(n15678), .A(n11785), .ZN(P2_U3463) );
  AOI22_X1 U14285 ( .A1(n15349), .A2(n14313), .B1(n7435), .B2(
        P2_REG1_REG_11__SCAN_IN), .ZN(n11786) );
  OAI21_X1 U14286 ( .B1(n11787), .B2(n7435), .A(n11786), .ZN(P2_U3510) );
  OAI21_X1 U14287 ( .B1(n11789), .B2(n11790), .A(n11788), .ZN(n15704) );
  AOI21_X1 U14288 ( .B1(n11791), .B2(n11790), .A(n13691), .ZN(n11795) );
  OAI22_X1 U14289 ( .A1(n11858), .A2(n13696), .B1(n11792), .B2(n13694), .ZN(
        n11793) );
  AOI21_X1 U14290 ( .B1(n11795), .B2(n11794), .A(n11793), .ZN(n15706) );
  INV_X1 U14291 ( .A(n15706), .ZN(n11796) );
  AOI21_X1 U14292 ( .B1(n15316), .B2(n15704), .A(n11796), .ZN(n11802) );
  INV_X1 U14293 ( .A(n13777), .ZN(n11897) );
  AOI22_X1 U14294 ( .A1(n11897), .A2(n15708), .B1(n15782), .B2(
        P3_REG1_REG_6__SCAN_IN), .ZN(n11797) );
  OAI21_X1 U14295 ( .B1(n11802), .B2(n15782), .A(n11797), .ZN(P3_U3465) );
  INV_X1 U14296 ( .A(P3_REG0_REG_6__SCAN_IN), .ZN(n11798) );
  OAI22_X1 U14297 ( .A1(n11799), .A2(n13825), .B1(n15775), .B2(n11798), .ZN(
        n11800) );
  INV_X1 U14298 ( .A(n11800), .ZN(n11801) );
  OAI21_X1 U14299 ( .B1(n11802), .B2(n15773), .A(n11801), .ZN(P3_U3408) );
  XNOR2_X1 U14300 ( .A(n11803), .B(n13137), .ZN(n15355) );
  INV_X1 U14301 ( .A(n15355), .ZN(n11817) );
  NAND2_X1 U14302 ( .A1(n11805), .A2(n11804), .ZN(n11806) );
  NAND3_X1 U14303 ( .A1(n11807), .A2(n15617), .A3(n11806), .ZN(n11810) );
  NAND2_X1 U14304 ( .A1(n13975), .A2(n12105), .ZN(n11809) );
  NAND2_X1 U14305 ( .A1(n13977), .A2(n13951), .ZN(n11808) );
  AND2_X1 U14306 ( .A1(n11809), .A2(n11808), .ZN(n11966) );
  NAND2_X1 U14307 ( .A1(n11810), .A2(n11966), .ZN(n15359) );
  AOI21_X1 U14308 ( .B1(n11811), .B2(n12967), .A(n6670), .ZN(n11812) );
  NAND2_X1 U14309 ( .A1(n11812), .A2(n12110), .ZN(n15356) );
  AOI22_X1 U14310 ( .A1(n15627), .A2(P2_REG2_REG_13__SCAN_IN), .B1(n11968), 
        .B2(n14208), .ZN(n11814) );
  NAND2_X1 U14311 ( .A1(n12967), .A2(n14228), .ZN(n11813) );
  OAI211_X1 U14312 ( .C1(n15356), .C2(n14213), .A(n11814), .B(n11813), .ZN(
        n11815) );
  AOI21_X1 U14313 ( .B1(n15359), .B2(n14226), .A(n11815), .ZN(n11816) );
  OAI21_X1 U14314 ( .B1(n14234), .B2(n11817), .A(n11816), .ZN(P2_U3252) );
  NAND2_X1 U14315 ( .A1(n11818), .A2(n11026), .ZN(n11820) );
  AOI22_X1 U14316 ( .A1(n7282), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n12415), 
        .B2(n14800), .ZN(n11819) );
  XNOR2_X1 U14317 ( .A(n12650), .B(n14700), .ZN(n12805) );
  OR2_X1 U14318 ( .A1(n12641), .A2(n11821), .ZN(n11822) );
  INV_X1 U14319 ( .A(n11933), .ZN(n11824) );
  AOI21_X1 U14320 ( .B1(n11835), .B2(n11825), .A(n11824), .ZN(n11839) );
  NAND2_X1 U14321 ( .A1(n12519), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n11832) );
  NAND2_X1 U14322 ( .A1(n9864), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n11831) );
  NAND2_X1 U14323 ( .A1(n11827), .A2(n11826), .ZN(n11828) );
  AND2_X1 U14324 ( .A1(n11947), .A2(n11828), .ZN(n12234) );
  NAND2_X1 U14325 ( .A1(n6677), .A2(n12234), .ZN(n11830) );
  NAND2_X1 U14326 ( .A1(n6683), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n11829) );
  NAND4_X1 U14327 ( .A1(n11832), .A2(n11831), .A3(n11830), .A4(n11829), .ZN(
        n14699) );
  AOI22_X1 U14328 ( .A1(n15001), .A2(n14701), .B1(n14699), .B2(n15002), .ZN(
        n11838) );
  OR2_X1 U14329 ( .A1(n12641), .A2(n14701), .ZN(n11833) );
  OAI21_X1 U14330 ( .B1(n11836), .B2(n11835), .A(n11943), .ZN(n15522) );
  NAND2_X1 U14331 ( .A1(n15522), .A2(n15080), .ZN(n11837) );
  OAI211_X1 U14332 ( .C1(n11839), .C2(n15481), .A(n11838), .B(n11837), .ZN(
        n15520) );
  INV_X1 U14333 ( .A(n15520), .ZN(n11847) );
  INV_X1 U14334 ( .A(n12650), .ZN(n15519) );
  INV_X1 U14335 ( .A(n11945), .ZN(n11841) );
  OAI211_X1 U14336 ( .C1(n15519), .C2(n11842), .A(n11841), .B(n15291), .ZN(
        n15517) );
  AOI22_X1 U14337 ( .A1(n15067), .A2(P1_REG2_REG_9__SCAN_IN), .B1(n12074), 
        .B2(n15283), .ZN(n11844) );
  NAND2_X1 U14338 ( .A1(n12650), .A2(n15285), .ZN(n11843) );
  OAI211_X1 U14339 ( .C1(n15517), .C2(n14994), .A(n11844), .B(n11843), .ZN(
        n11845) );
  AOI21_X1 U14340 ( .B1(n15522), .B2(n15086), .A(n11845), .ZN(n11846) );
  OAI21_X1 U14341 ( .B1(n11847), .B2(n15067), .A(n11846), .ZN(P1_U3284) );
  INV_X1 U14342 ( .A(n12425), .ZN(n11874) );
  OAI222_X1 U14343 ( .A1(n14396), .A2(n11874), .B1(n11849), .B2(P2_U3088), 
        .C1(n11848), .C2(n12861), .ZN(P2_U3307) );
  MUX2_X1 U14344 ( .A(n12017), .B(n11851), .S(n11850), .Z(n11853) );
  XNOR2_X1 U14345 ( .A(n11853), .B(n11852), .ZN(n11861) );
  AOI21_X1 U14346 ( .B1(n13281), .B2(n12018), .A(n11854), .ZN(n11857) );
  NAND2_X1 U14347 ( .A1(n13337), .A2(n11855), .ZN(n11856) );
  OAI211_X1 U14348 ( .C1(n11858), .C2(n13315), .A(n11857), .B(n11856), .ZN(
        n11859) );
  AOI21_X1 U14349 ( .B1(n12020), .B2(n13350), .A(n11859), .ZN(n11860) );
  OAI21_X1 U14350 ( .B1(n11861), .B2(n13352), .A(n11860), .ZN(P3_U3161) );
  XNOR2_X1 U14351 ( .A(n15766), .B(n13254), .ZN(n12139) );
  XNOR2_X1 U14352 ( .A(n12139), .B(n12050), .ZN(n11866) );
  NOR2_X1 U14353 ( .A1(n11862), .A2(n12018), .ZN(n11863) );
  OR2_X1 U14354 ( .A1(n11864), .A2(n11863), .ZN(n11865) );
  AOI211_X1 U14355 ( .C1(n11866), .C2(n11865), .A(n13352), .B(n12140), .ZN(
        n11873) );
  AOI21_X1 U14356 ( .B1(n12223), .B2(n13281), .A(n11867), .ZN(n11871) );
  NAND2_X1 U14357 ( .A1(n13350), .A2(n12009), .ZN(n11870) );
  NAND2_X1 U14358 ( .A1(n13337), .A2(n15766), .ZN(n11869) );
  NAND2_X1 U14359 ( .A1(n13343), .A2(n12018), .ZN(n11868) );
  NAND4_X1 U14360 ( .A1(n11871), .A2(n11870), .A3(n11869), .A4(n11868), .ZN(
        n11872) );
  OR2_X1 U14361 ( .A1(n11873), .A2(n11872), .ZN(P3_U3157) );
  OAI222_X1 U14362 ( .A1(n12770), .A2(P1_U3086), .B1(n15238), .B2(n11874), 
        .C1(n12426), .C2(n15239), .ZN(P1_U3335) );
  NAND2_X1 U14363 ( .A1(n11876), .A2(n11875), .ZN(n11877) );
  NOR2_X1 U14364 ( .A1(n11877), .A2(n14004), .ZN(n14001) );
  AOI21_X1 U14365 ( .B1(n11877), .B2(n14004), .A(n14001), .ZN(n11878) );
  INV_X1 U14366 ( .A(n11878), .ZN(n11879) );
  NOR2_X1 U14367 ( .A1(P2_REG2_REG_18__SCAN_IN), .A2(n11879), .ZN(n14002) );
  AOI21_X1 U14368 ( .B1(n11879), .B2(P2_REG2_REG_18__SCAN_IN), .A(n14002), 
        .ZN(n11889) );
  INV_X1 U14369 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n11881) );
  NAND2_X1 U14370 ( .A1(P2_REG3_REG_18__SCAN_IN), .A2(P2_U3088), .ZN(n11880)
         );
  OAI21_X1 U14371 ( .B1(n15566), .B2(n11881), .A(n11880), .ZN(n11882) );
  AOI21_X1 U14372 ( .B1(n14004), .B2(n15603), .A(n11882), .ZN(n11887) );
  OAI21_X1 U14373 ( .B1(n14308), .B2(n11884), .A(n11883), .ZN(n14005) );
  XOR2_X1 U14374 ( .A(n14004), .B(n14005), .Z(n11885) );
  NAND2_X1 U14375 ( .A1(P2_REG1_REG_18__SCAN_IN), .A2(n11885), .ZN(n14007) );
  OAI211_X1 U14376 ( .C1(n11885), .C2(P2_REG1_REG_18__SCAN_IN), .A(n15609), 
        .B(n14007), .ZN(n11886) );
  OAI211_X1 U14377 ( .C1(n11889), .C2(n11888), .A(n11887), .B(n11886), .ZN(
        P2_U3232) );
  AOI21_X1 U14378 ( .B1(n15316), .B2(n11891), .A(n11890), .ZN(n11899) );
  INV_X1 U14379 ( .A(P3_REG0_REG_7__SCAN_IN), .ZN(n11892) );
  OAI22_X1 U14380 ( .A1(n11893), .A2(n13825), .B1(n15775), .B2(n11892), .ZN(
        n11894) );
  INV_X1 U14381 ( .A(n11894), .ZN(n11895) );
  OAI21_X1 U14382 ( .B1(n11899), .B2(n15773), .A(n11895), .ZN(P3_U3411) );
  AOI22_X1 U14383 ( .A1(n11897), .A2(n11896), .B1(n15782), .B2(
        P3_REG1_REG_7__SCAN_IN), .ZN(n11898) );
  OAI21_X1 U14384 ( .B1(n11899), .B2(n15782), .A(n11898), .ZN(P3_U3466) );
  INV_X1 U14385 ( .A(P3_REG2_REG_11__SCAN_IN), .ZN(n12052) );
  AOI21_X1 U14386 ( .B1(n12052), .B2(n11901), .A(n11972), .ZN(n11919) );
  NOR2_X1 U14387 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11902), .ZN(n12142) );
  INV_X1 U14388 ( .A(n12142), .ZN(n11903) );
  OAI21_X1 U14389 ( .B1(n13492), .B2(n11904), .A(n11903), .ZN(n11912) );
  INV_X1 U14390 ( .A(n11905), .ZN(n11906) );
  MUX2_X1 U14391 ( .A(P3_REG2_REG_11__SCAN_IN), .B(P3_REG1_REG_11__SCAN_IN), 
        .S(n6945), .Z(n11982) );
  XNOR2_X1 U14392 ( .A(n11982), .B(n11981), .ZN(n11908) );
  AOI21_X1 U14393 ( .B1(n11909), .B2(n11908), .A(n11985), .ZN(n11910) );
  NOR2_X1 U14394 ( .A1(n11910), .A2(n15692), .ZN(n11911) );
  AOI211_X1 U14395 ( .C1(n15699), .C2(n11977), .A(n11912), .B(n11911), .ZN(
        n11918) );
  AOI21_X1 U14396 ( .B1(n9194), .B2(n11915), .A(n11978), .ZN(n11916) );
  OR2_X1 U14397 ( .A1(n11916), .A2(n15693), .ZN(n11917) );
  OAI211_X1 U14398 ( .C1(n11919), .C2(n15694), .A(n11918), .B(n11917), .ZN(
        P3_U3193) );
  NAND2_X1 U14399 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n14606)
         );
  XNOR2_X1 U14400 ( .A(n11931), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n14813) );
  NAND2_X1 U14401 ( .A1(n12395), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n11921) );
  NAND2_X1 U14402 ( .A1(n11921), .A2(n11920), .ZN(n14812) );
  XOR2_X1 U14403 ( .A(n14813), .B(n14812), .Z(n11922) );
  NAND2_X1 U14404 ( .A1(n14833), .A2(n11922), .ZN(n11923) );
  NAND2_X1 U14405 ( .A1(n14606), .A2(n11923), .ZN(n11924) );
  AOI21_X1 U14406 ( .B1(n14819), .B2(P1_ADDR_REG_17__SCAN_IN), .A(n11924), 
        .ZN(n11930) );
  INV_X1 U14407 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n15030) );
  MUX2_X1 U14408 ( .A(P1_REG2_REG_17__SCAN_IN), .B(n15030), .S(n14811), .Z(
        n11928) );
  NAND2_X1 U14409 ( .A1(n12395), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n11926) );
  NAND2_X1 U14410 ( .A1(n11926), .A2(n11925), .ZN(n11927) );
  NAND2_X1 U14411 ( .A1(n11928), .A2(n11927), .ZN(n14810) );
  OAI211_X1 U14412 ( .C1(n11928), .C2(n11927), .A(n14838), .B(n14810), .ZN(
        n11929) );
  OAI211_X1 U14413 ( .C1(n15472), .C2(n11931), .A(n11930), .B(n11929), .ZN(
        P1_U3260) );
  NAND2_X1 U14414 ( .A1(n12650), .A2(n12239), .ZN(n11932) );
  NAND2_X1 U14415 ( .A1(n11933), .A2(n11932), .ZN(n11938) );
  NAND2_X1 U14416 ( .A1(n11934), .A2(n11026), .ZN(n11937) );
  AOI22_X1 U14417 ( .A1(n7282), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n12415), 
        .B2(n11935), .ZN(n11936) );
  XNOR2_X1 U14418 ( .A(n12654), .B(n15386), .ZN(n12809) );
  AOI21_X1 U14419 ( .B1(n11938), .B2(n12809), .A(n15481), .ZN(n11941) );
  INV_X1 U14420 ( .A(n11938), .ZN(n11940) );
  INV_X1 U14421 ( .A(n12809), .ZN(n11939) );
  NAND2_X1 U14422 ( .A1(n11940), .A2(n11939), .ZN(n12154) );
  AOI22_X1 U14423 ( .A1(n11941), .A2(n12154), .B1(n15001), .B2(n14700), .ZN(
        n12080) );
  OR2_X1 U14424 ( .A1(n12650), .A2(n14700), .ZN(n11942) );
  OAI21_X1 U14425 ( .B1(n11944), .B2(n12809), .A(n12161), .ZN(n12077) );
  INV_X1 U14426 ( .A(n12654), .ZN(n12243) );
  OAI21_X1 U14427 ( .B1(n11945), .B2(n12243), .A(n15291), .ZN(n11955) );
  NAND2_X1 U14428 ( .A1(n6681), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n11953) );
  AND2_X1 U14429 ( .A1(n11947), .A2(n11946), .ZN(n11949) );
  OR2_X1 U14430 ( .A1(n11949), .A2(n11948), .ZN(n15401) );
  INV_X1 U14431 ( .A(n15401), .ZN(n12163) );
  NAND2_X1 U14432 ( .A1(n6677), .A2(n12163), .ZN(n11952) );
  NAND2_X1 U14433 ( .A1(n6683), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n11951) );
  NAND2_X1 U14434 ( .A1(n12519), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n11950) );
  NAND4_X1 U14435 ( .A1(n11953), .A2(n11952), .A3(n11951), .A4(n11950), .ZN(
        n14698) );
  AND2_X1 U14436 ( .A1(n14698), .A2(n15002), .ZN(n12236) );
  INV_X1 U14437 ( .A(n12236), .ZN(n11954) );
  OAI21_X1 U14438 ( .B1(n11955), .B2(n12162), .A(n11954), .ZN(n12078) );
  NAND2_X1 U14439 ( .A1(n12078), .A2(n15293), .ZN(n11957) );
  AOI22_X1 U14440 ( .A1(n15067), .A2(P1_REG2_REG_10__SCAN_IN), .B1(n12234), 
        .B2(n15283), .ZN(n11956) );
  OAI211_X1 U14441 ( .C1(n12243), .C2(n15013), .A(n11957), .B(n11956), .ZN(
        n11958) );
  AOI21_X1 U14442 ( .B1(n12077), .B2(n15294), .A(n11958), .ZN(n11959) );
  OAI21_X1 U14443 ( .B1(n12080), .B2(n15067), .A(n11959), .ZN(P1_U3283) );
  INV_X1 U14444 ( .A(n12435), .ZN(n11961) );
  OAI222_X1 U14445 ( .A1(n12861), .A2(n11960), .B1(n14396), .B2(n11961), .C1(
        P2_U3088), .C2(n13158), .ZN(P2_U3306) );
  INV_X1 U14446 ( .A(n12594), .ZN(n12788) );
  OAI222_X1 U14447 ( .A1(P1_U3086), .A2(n12788), .B1(n15238), .B2(n11961), 
        .C1(n9370), .C2(n15239), .ZN(P1_U3334) );
  INV_X1 U14448 ( .A(n12967), .ZN(n15357) );
  OAI211_X1 U14449 ( .C1(n11964), .C2(n11963), .A(n11962), .B(n15345), .ZN(
        n11970) );
  OAI22_X1 U14450 ( .A1(n13953), .A2(n11966), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n11965), .ZN(n11967) );
  AOI21_X1 U14451 ( .B1(n11968), .B2(n13944), .A(n11967), .ZN(n11969) );
  OAI211_X1 U14452 ( .C1(n15357), .C2(n13958), .A(n11970), .B(n11969), .ZN(
        P2_U3206) );
  NOR2_X1 U14453 ( .A1(n11977), .A2(n11971), .ZN(n11973) );
  NAND2_X1 U14454 ( .A1(P3_REG2_REG_12__SCAN_IN), .A2(n13377), .ZN(n11974) );
  OAI21_X1 U14455 ( .B1(P3_REG2_REG_12__SCAN_IN), .B2(n13377), .A(n11974), 
        .ZN(n11975) );
  NOR2_X1 U14456 ( .A1(n11976), .A2(n11975), .ZN(n13359) );
  AOI21_X1 U14457 ( .B1(n11976), .B2(n11975), .A(n13359), .ZN(n11994) );
  NOR2_X1 U14458 ( .A1(n11977), .A2(n6765), .ZN(n11979) );
  NAND2_X1 U14459 ( .A1(P3_REG1_REG_12__SCAN_IN), .A2(n13377), .ZN(n11980) );
  OAI21_X1 U14460 ( .B1(P3_REG1_REG_12__SCAN_IN), .B2(n13377), .A(n11980), 
        .ZN(n13375) );
  XNOR2_X1 U14461 ( .A(n13376), .B(n13375), .ZN(n11992) );
  NOR2_X1 U14462 ( .A1(n11982), .A2(n11981), .ZN(n11984) );
  MUX2_X1 U14463 ( .A(P3_REG2_REG_12__SCAN_IN), .B(P3_REG1_REG_12__SCAN_IN), 
        .S(n6945), .Z(n13365) );
  XNOR2_X1 U14464 ( .A(n13365), .B(n13377), .ZN(n11983) );
  NOR3_X1 U14465 ( .A1(n11985), .A2(n11984), .A3(n11983), .ZN(n13370) );
  INV_X1 U14466 ( .A(n13370), .ZN(n11987) );
  OAI21_X1 U14467 ( .B1(n11985), .B2(n11984), .A(n11983), .ZN(n11986) );
  NAND3_X1 U14468 ( .A1(n11987), .A2(n13529), .A3(n11986), .ZN(n11990) );
  NOR2_X1 U14469 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11988), .ZN(n12373) );
  AOI21_X1 U14470 ( .B1(n15698), .B2(P3_ADDR_REG_12__SCAN_IN), .A(n12373), 
        .ZN(n11989) );
  OAI211_X1 U14471 ( .C1(n13521), .C2(n13377), .A(n11990), .B(n11989), .ZN(
        n11991) );
  AOI21_X1 U14472 ( .B1(n13471), .B2(n11992), .A(n11991), .ZN(n11993) );
  OAI21_X1 U14473 ( .B1(n11994), .B2(n15694), .A(n11993), .ZN(P3_U3194) );
  NAND2_X1 U14474 ( .A1(n11995), .A2(n12005), .ZN(n11996) );
  NAND2_X1 U14475 ( .A1(n11997), .A2(n11996), .ZN(n15770) );
  AND2_X1 U14476 ( .A1(n11999), .A2(n11998), .ZN(n12015) );
  NAND2_X1 U14477 ( .A1(n12015), .A2(n12000), .ZN(n12003) );
  AND2_X1 U14478 ( .A1(n12003), .A2(n12001), .ZN(n12006) );
  NAND2_X1 U14479 ( .A1(n12003), .A2(n12002), .ZN(n12004) );
  OAI211_X1 U14480 ( .C1(n12006), .C2(n12005), .A(n12004), .B(n15722), .ZN(
        n12008) );
  AOI22_X1 U14481 ( .A1(n12223), .A2(n15719), .B1(n15717), .B2(n12018), .ZN(
        n12007) );
  NAND2_X1 U14482 ( .A1(n12008), .A2(n12007), .ZN(n15772) );
  NAND2_X1 U14483 ( .A1(n15772), .A2(n15733), .ZN(n12014) );
  INV_X1 U14484 ( .A(n12009), .ZN(n12010) );
  OAI22_X1 U14485 ( .A1(n13714), .A2(n12011), .B1(n12010), .B2(n15727), .ZN(
        n12012) );
  AOI21_X1 U14486 ( .B1(P3_REG2_REG_10__SCAN_IN), .B2(n15735), .A(n12012), 
        .ZN(n12013) );
  OAI211_X1 U14487 ( .C1(n13688), .C2(n15770), .A(n12014), .B(n12013), .ZN(
        P3_U3223) );
  NAND2_X1 U14488 ( .A1(n12015), .A2(n12016), .ZN(n12032) );
  OAI21_X1 U14489 ( .B1(n12016), .B2(n12015), .A(n12032), .ZN(n12019) );
  AOI222_X1 U14490 ( .A1(n15722), .A2(n12019), .B1(n12018), .B2(n15719), .C1(
        n12017), .C2(n15717), .ZN(n12168) );
  INV_X1 U14491 ( .A(n12020), .ZN(n12021) );
  OAI22_X1 U14492 ( .A1(n13714), .A2(n12173), .B1(n12021), .B2(n15727), .ZN(
        n12027) );
  OAI21_X1 U14493 ( .B1(n12024), .B2(n12023), .A(n12022), .ZN(n12025) );
  INV_X1 U14494 ( .A(n12025), .ZN(n12169) );
  NOR2_X1 U14495 ( .A1(n12169), .A2(n13688), .ZN(n12026) );
  AOI211_X1 U14496 ( .C1(n15735), .C2(P3_REG2_REG_8__SCAN_IN), .A(n12027), .B(
        n12026), .ZN(n12028) );
  OAI21_X1 U14497 ( .B1(n12168), .B2(n15735), .A(n12028), .ZN(P3_U3225) );
  XNOR2_X1 U14498 ( .A(n12029), .B(n12034), .ZN(n15760) );
  AND2_X1 U14499 ( .A1(n12032), .A2(n12030), .ZN(n12035) );
  NAND2_X1 U14500 ( .A1(n12032), .A2(n12031), .ZN(n12033) );
  OAI211_X1 U14501 ( .C1(n12035), .C2(n12034), .A(n12033), .B(n15722), .ZN(
        n12037) );
  AOI22_X1 U14502 ( .A1(n12145), .A2(n15719), .B1(n15717), .B2(n13357), .ZN(
        n12036) );
  OAI211_X1 U14503 ( .C1(n15764), .C2(n15760), .A(n12037), .B(n12036), .ZN(
        n15762) );
  NAND2_X1 U14504 ( .A1(n15762), .A2(n15733), .ZN(n12042) );
  INV_X1 U14505 ( .A(n12038), .ZN(n12039) );
  OAI22_X1 U14506 ( .A1(n13714), .A2(n15759), .B1(n12039), .B2(n15727), .ZN(
        n12040) );
  AOI21_X1 U14507 ( .B1(P3_REG2_REG_9__SCAN_IN), .B2(n15735), .A(n12040), .ZN(
        n12041) );
  OAI211_X1 U14508 ( .C1(n15760), .C2(n15729), .A(n12042), .B(n12041), .ZN(
        P3_U3224) );
  INV_X1 U14509 ( .A(n12043), .ZN(n12044) );
  AOI21_X1 U14510 ( .B1(n7627), .B2(n12045), .A(n12044), .ZN(n15328) );
  INV_X1 U14511 ( .A(n12091), .ZN(n12046) );
  AOI21_X1 U14512 ( .B1(n12048), .B2(n12047), .A(n12046), .ZN(n12049) );
  OAI222_X1 U14513 ( .A1(n13696), .A2(n12230), .B1(n13694), .B2(n12050), .C1(
        n13691), .C2(n12049), .ZN(n15330) );
  NAND2_X1 U14514 ( .A1(n15330), .A2(n15733), .ZN(n12055) );
  INV_X1 U14515 ( .A(n12144), .ZN(n12051) );
  OAI22_X1 U14516 ( .A1(n15733), .A2(n12052), .B1(n12051), .B2(n15727), .ZN(
        n12053) );
  AOI21_X1 U14517 ( .B1(n12143), .B2(n15707), .A(n12053), .ZN(n12054) );
  OAI211_X1 U14518 ( .C1(n15328), .C2(n13688), .A(n12055), .B(n12054), .ZN(
        P3_U3222) );
  NAND2_X1 U14519 ( .A1(n12457), .A2(n12056), .ZN(n12057) );
  OAI211_X1 U14520 ( .C1(n12458), .C2(n15239), .A(n12057), .B(n12844), .ZN(
        P1_U3332) );
  NAND2_X1 U14521 ( .A1(n12457), .A2(n14389), .ZN(n12059) );
  OR2_X1 U14522 ( .A1(n12058), .A2(P2_U3088), .ZN(n13171) );
  OAI211_X1 U14523 ( .C1(n12060), .C2(n12861), .A(n12059), .B(n13171), .ZN(
        P2_U3304) );
  AND2_X1 U14524 ( .A1(n14517), .A2(n14700), .ZN(n12061) );
  AOI21_X1 U14525 ( .B1(n12650), .B2(n9893), .A(n12061), .ZN(n12240) );
  NAND2_X1 U14526 ( .A1(n12650), .A2(n14511), .ZN(n12063) );
  NAND2_X1 U14527 ( .A1(n14700), .A2(n9893), .ZN(n12062) );
  NAND2_X1 U14528 ( .A1(n12063), .A2(n12062), .ZN(n12064) );
  NAND2_X1 U14529 ( .A1(n12065), .A2(n12066), .ZN(n12067) );
  AOI211_X1 U14530 ( .C1(n12070), .C2(n12069), .A(n15392), .B(n6827), .ZN(
        n12071) );
  INV_X1 U14531 ( .A(n12071), .ZN(n12076) );
  NAND2_X1 U14532 ( .A1(n14677), .A2(n14701), .ZN(n12072) );
  NAND2_X1 U14533 ( .A1(P1_REG3_REG_9__SCAN_IN), .A2(P1_U3086), .ZN(n14791) );
  OAI211_X1 U14534 ( .C1(n15386), .C2(n15384), .A(n12072), .B(n14791), .ZN(
        n12073) );
  AOI21_X1 U14535 ( .B1(n14680), .B2(n12074), .A(n12073), .ZN(n12075) );
  OAI211_X1 U14536 ( .C1(n15519), .C2(n14683), .A(n12076), .B(n12075), .ZN(
        P1_U3231) );
  INV_X1 U14537 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n12083) );
  INV_X1 U14538 ( .A(n12077), .ZN(n12081) );
  AOI21_X1 U14539 ( .B1(n12654), .B2(n15495), .A(n12078), .ZN(n12079) );
  OAI211_X1 U14540 ( .C1(n12081), .C2(n15482), .A(n12080), .B(n12079), .ZN(
        n12084) );
  NAND2_X1 U14541 ( .A1(n12084), .A2(n15526), .ZN(n12082) );
  OAI21_X1 U14542 ( .B1(n15526), .B2(n12083), .A(n12082), .ZN(P1_U3489) );
  NAND2_X1 U14543 ( .A1(n12084), .A2(n15537), .ZN(n12085) );
  OAI21_X1 U14544 ( .B1(n15537), .B2(n12086), .A(n12085), .ZN(P1_U3538) );
  XNOR2_X1 U14545 ( .A(n12087), .B(n12089), .ZN(n15322) );
  NAND2_X1 U14546 ( .A1(n12088), .A2(n15722), .ZN(n12094) );
  AOI21_X1 U14547 ( .B1(n12091), .B2(n12090), .A(n12089), .ZN(n12093) );
  AOI22_X1 U14548 ( .A1(n12223), .A2(n15717), .B1(n15719), .B2(n13355), .ZN(
        n12092) );
  OAI21_X1 U14549 ( .B1(n12094), .B2(n12093), .A(n12092), .ZN(n15323) );
  AOI22_X1 U14550 ( .A1(n15735), .A2(P3_REG2_REG_12__SCAN_IN), .B1(n15709), 
        .B2(n12374), .ZN(n12095) );
  OAI21_X1 U14551 ( .B1(n12096), .B2(n13714), .A(n12095), .ZN(n12097) );
  AOI21_X1 U14552 ( .B1(n15323), .B2(n15733), .A(n12097), .ZN(n12098) );
  OAI21_X1 U14553 ( .B1(n13688), .B2(n15322), .A(n12098), .ZN(P3_U3221) );
  INV_X1 U14554 ( .A(n12099), .ZN(n12100) );
  AOI21_X1 U14555 ( .B1(n6966), .B2(n12101), .A(n12100), .ZN(n12120) );
  INV_X1 U14556 ( .A(n12120), .ZN(n12115) );
  INV_X1 U14557 ( .A(n12102), .ZN(n12103) );
  AOI21_X1 U14558 ( .B1(n13141), .B2(n12104), .A(n12103), .ZN(n12108) );
  NAND2_X1 U14559 ( .A1(n13974), .A2(n12105), .ZN(n12107) );
  NAND2_X1 U14560 ( .A1(n13976), .A2(n13951), .ZN(n12106) );
  AND2_X1 U14561 ( .A1(n12107), .A2(n12106), .ZN(n12133) );
  OAI21_X1 U14562 ( .B1(n12108), .B2(n14220), .A(n12133), .ZN(n12117) );
  NAND2_X1 U14563 ( .A1(n12117), .A2(n14226), .ZN(n12114) );
  AOI211_X1 U14564 ( .C1(n12988), .C2(n12110), .A(n6670), .B(n12109), .ZN(
        n12116) );
  INV_X1 U14565 ( .A(n12988), .ZN(n12138) );
  AOI22_X1 U14566 ( .A1(n15627), .A2(P2_REG2_REG_14__SCAN_IN), .B1(n12135), 
        .B2(n14208), .ZN(n12111) );
  OAI21_X1 U14567 ( .B1(n12138), .B2(n14157), .A(n12111), .ZN(n12112) );
  AOI21_X1 U14568 ( .B1(n12116), .B2(n14160), .A(n12112), .ZN(n12113) );
  OAI211_X1 U14569 ( .C1(n14234), .C2(n12115), .A(n12114), .B(n12113), .ZN(
        P2_U3251) );
  NOR2_X1 U14570 ( .A1(n12117), .A2(n12116), .ZN(n12123) );
  AOI22_X1 U14571 ( .A1(n12988), .A2(n14375), .B1(P2_REG0_REG_14__SCAN_IN), 
        .B2(n15678), .ZN(n12119) );
  NAND2_X1 U14572 ( .A1(n12120), .A2(n8998), .ZN(n12118) );
  OAI211_X1 U14573 ( .C1(n12123), .C2(n15678), .A(n12119), .B(n12118), .ZN(
        P2_U3472) );
  AOI22_X1 U14574 ( .A1(n12988), .A2(n14313), .B1(P2_REG1_REG_14__SCAN_IN), 
        .B2(n7435), .ZN(n12122) );
  INV_X1 U14575 ( .A(n14316), .ZN(n14277) );
  NAND2_X1 U14576 ( .A1(n12120), .A2(n14277), .ZN(n12121) );
  OAI211_X1 U14577 ( .C1(n12123), .C2(n7435), .A(n12122), .B(n12121), .ZN(
        P2_U3513) );
  OAI22_X1 U14578 ( .A1(n12124), .A2(P3_U3151), .B1(n8147), .B2(n13840), .ZN(
        n12125) );
  AOI21_X1 U14579 ( .B1(n12126), .B2(n13828), .A(n12125), .ZN(n12127) );
  INV_X1 U14580 ( .A(n12127), .ZN(P3_U3271) );
  OAI21_X1 U14581 ( .B1(n12130), .B2(n12129), .A(n12128), .ZN(n12131) );
  NAND2_X1 U14582 ( .A1(n12131), .A2(n15345), .ZN(n12137) );
  OAI22_X1 U14583 ( .A1(n13953), .A2(n12133), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n12132), .ZN(n12134) );
  AOI21_X1 U14584 ( .B1(n12135), .B2(n13944), .A(n12134), .ZN(n12136) );
  OAI211_X1 U14585 ( .C1(n12138), .C2(n13958), .A(n12137), .B(n12136), .ZN(
        P2_U3187) );
  INV_X1 U14586 ( .A(n12139), .ZN(n12141) );
  XNOR2_X1 U14587 ( .A(n15326), .B(n13254), .ZN(n12222) );
  XNOR2_X1 U14588 ( .A(n12224), .B(n12377), .ZN(n12151) );
  AOI21_X1 U14589 ( .B1(n13356), .B2(n13281), .A(n12142), .ZN(n12149) );
  NAND2_X1 U14590 ( .A1(n13337), .A2(n12143), .ZN(n12148) );
  NAND2_X1 U14591 ( .A1(n13350), .A2(n12144), .ZN(n12147) );
  NAND2_X1 U14592 ( .A1(n12145), .A2(n13343), .ZN(n12146) );
  NAND4_X1 U14593 ( .A1(n12149), .A2(n12148), .A3(n12147), .A4(n12146), .ZN(
        n12150) );
  AOI21_X1 U14594 ( .B1(n12151), .B2(n13322), .A(n12150), .ZN(n12152) );
  INV_X1 U14595 ( .A(n12152), .ZN(P3_U3176) );
  INV_X1 U14596 ( .A(n15385), .ZN(n12659) );
  OR2_X1 U14597 ( .A1(n12654), .A2(n15386), .ZN(n12153) );
  NAND2_X1 U14598 ( .A1(n12154), .A2(n12153), .ZN(n12286) );
  NAND2_X1 U14599 ( .A1(n12155), .A2(n11026), .ZN(n12158) );
  AOI22_X1 U14600 ( .A1(n7282), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n12415), 
        .B2(n12156), .ZN(n12157) );
  OR2_X1 U14601 ( .A1(n15398), .A2(n14698), .ZN(n12274) );
  NAND2_X1 U14602 ( .A1(n15398), .A2(n14698), .ZN(n12272) );
  NAND2_X1 U14603 ( .A1(n12274), .A2(n12272), .ZN(n12807) );
  XOR2_X1 U14604 ( .A(n12286), .B(n12807), .Z(n12159) );
  AOI222_X1 U14605 ( .A1(n14699), .A2(n15001), .B1(n12659), .B2(n15002), .C1(
        n15280), .C2(n12159), .ZN(n15410) );
  OR2_X1 U14606 ( .A1(n12654), .A2(n14699), .ZN(n12160) );
  XOR2_X1 U14607 ( .A(n12273), .B(n12807), .Z(n15414) );
  NAND2_X1 U14608 ( .A1(n12162), .A2(n15409), .ZN(n12280) );
  OAI211_X1 U14609 ( .C1(n12162), .C2(n15409), .A(n15291), .B(n12280), .ZN(
        n15408) );
  AOI22_X1 U14610 ( .A1(n15067), .A2(P1_REG2_REG_11__SCAN_IN), .B1(n12163), 
        .B2(n15283), .ZN(n12165) );
  NAND2_X1 U14611 ( .A1(n15398), .A2(n15285), .ZN(n12164) );
  OAI211_X1 U14612 ( .C1(n15408), .C2(n14994), .A(n12165), .B(n12164), .ZN(
        n12166) );
  AOI21_X1 U14613 ( .B1(n15414), .B2(n15294), .A(n12166), .ZN(n12167) );
  OAI21_X1 U14614 ( .B1(n15410), .B2(n15067), .A(n12167), .ZN(P1_U3282) );
  OAI21_X1 U14615 ( .B1(n15327), .B2(n12169), .A(n12168), .ZN(n12175) );
  INV_X1 U14616 ( .A(P3_REG0_REG_8__SCAN_IN), .ZN(n12170) );
  OAI22_X1 U14617 ( .A1(n12173), .A2(n13825), .B1(n15775), .B2(n12170), .ZN(
        n12171) );
  AOI21_X1 U14618 ( .B1(n12175), .B2(n15775), .A(n12171), .ZN(n12172) );
  INV_X1 U14619 ( .A(n12172), .ZN(P3_U3414) );
  OAI22_X1 U14620 ( .A1(n13777), .A2(n12173), .B1(n15784), .B2(n9135), .ZN(
        n12174) );
  AOI21_X1 U14621 ( .B1(n12175), .B2(n15784), .A(n12174), .ZN(n12176) );
  INV_X1 U14622 ( .A(n12176), .ZN(P3_U3467) );
  INV_X1 U14623 ( .A(n12177), .ZN(n12179) );
  OAI222_X1 U14624 ( .A1(P3_U3151), .A2(n12180), .B1(n13851), .B2(n12179), 
        .C1(n12178), .C2(n13840), .ZN(P3_U3270) );
  OAI211_X1 U14625 ( .C1(n6821), .C2(n12181), .A(n12213), .B(n15617), .ZN(
        n12184) );
  NAND2_X1 U14626 ( .A1(n13973), .A2(n13952), .ZN(n12183) );
  NAND2_X1 U14627 ( .A1(n13975), .A2(n13951), .ZN(n12182) );
  AND2_X1 U14628 ( .A1(n12183), .A2(n12182), .ZN(n12259) );
  NAND2_X1 U14629 ( .A1(n12184), .A2(n12259), .ZN(n12249) );
  AOI21_X1 U14630 ( .B1(n12261), .B2(n14208), .A(n12249), .ZN(n12192) );
  INV_X1 U14631 ( .A(n12205), .ZN(n12185) );
  AOI211_X1 U14632 ( .C1(n12980), .C2(n12186), .A(n6670), .B(n12185), .ZN(
        n12250) );
  INV_X1 U14633 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n12187) );
  OAI22_X1 U14634 ( .A1(n8888), .A2(n14157), .B1(n12187), .B2(n14226), .ZN(
        n12188) );
  AOI21_X1 U14635 ( .B1(n12250), .B2(n14160), .A(n12188), .ZN(n12191) );
  OAI21_X1 U14636 ( .B1(n7738), .B2(n13142), .A(n12189), .ZN(n12252) );
  NAND2_X1 U14637 ( .A1(n12252), .A2(n14134), .ZN(n12190) );
  OAI211_X1 U14638 ( .C1(n12192), .C2(n15627), .A(n12191), .B(n12190), .ZN(
        P2_U3250) );
  XNOR2_X1 U14639 ( .A(n12193), .B(n7736), .ZN(n12194) );
  NAND2_X1 U14640 ( .A1(n12194), .A2(n15722), .ZN(n12196) );
  AOI22_X1 U14641 ( .A1(n13356), .A2(n15717), .B1(n15719), .B2(n13706), .ZN(
        n12195) );
  NAND2_X1 U14642 ( .A1(n12196), .A2(n12195), .ZN(n15321) );
  INV_X1 U14643 ( .A(n15321), .ZN(n12202) );
  XNOR2_X1 U14644 ( .A(n12197), .B(n7736), .ZN(n15317) );
  AOI22_X1 U14645 ( .A1(n15735), .A2(P3_REG2_REG_13__SCAN_IN), .B1(n15709), 
        .B2(n12227), .ZN(n12198) );
  OAI21_X1 U14646 ( .B1(n12199), .B2(n13714), .A(n12198), .ZN(n12200) );
  AOI21_X1 U14647 ( .B1(n15317), .B2(n13716), .A(n12200), .ZN(n12201) );
  OAI21_X1 U14648 ( .B1(n12202), .B2(n15735), .A(n12201), .ZN(P3_U3220) );
  OAI21_X1 U14649 ( .B1(n12204), .B2(n12212), .A(n12203), .ZN(n14380) );
  AOI211_X1 U14650 ( .C1(n14376), .C2(n12205), .A(n6670), .B(n6816), .ZN(
        n14310) );
  INV_X1 U14651 ( .A(n14376), .ZN(n12206) );
  NOR2_X1 U14652 ( .A1(n12206), .A2(n14157), .ZN(n12210) );
  INV_X1 U14653 ( .A(n12207), .ZN(n13891) );
  OAI22_X1 U14654 ( .A1(n14226), .A2(n12208), .B1(n13891), .B2(n15621), .ZN(
        n12209) );
  AOI211_X1 U14655 ( .C1(n14310), .C2(n14160), .A(n12210), .B(n12209), .ZN(
        n12221) );
  NAND3_X1 U14656 ( .A1(n12213), .A2(n12212), .A3(n12211), .ZN(n12214) );
  NAND3_X1 U14657 ( .A1(n12215), .A2(n15617), .A3(n12214), .ZN(n12219) );
  NAND2_X1 U14658 ( .A1(n13972), .A2(n13952), .ZN(n12217) );
  NAND2_X1 U14659 ( .A1(n13974), .A2(n13951), .ZN(n12216) );
  NAND2_X1 U14660 ( .A1(n12217), .A2(n12216), .ZN(n13889) );
  INV_X1 U14661 ( .A(n13889), .ZN(n12218) );
  NAND2_X1 U14662 ( .A1(n12219), .A2(n12218), .ZN(n14311) );
  NAND2_X1 U14663 ( .A1(n14311), .A2(n14226), .ZN(n12220) );
  OAI211_X1 U14664 ( .C1(n14380), .C2(n14234), .A(n12221), .B(n12220), .ZN(
        P2_U3249) );
  XNOR2_X1 U14665 ( .A(n15325), .B(n13207), .ZN(n12225) );
  NOR2_X1 U14666 ( .A1(n13356), .A2(n12225), .ZN(n12378) );
  NAND2_X1 U14667 ( .A1(n13356), .A2(n12225), .ZN(n12379) );
  XNOR2_X1 U14668 ( .A(n15318), .B(n13207), .ZN(n13184) );
  XNOR2_X1 U14669 ( .A(n13184), .B(n13180), .ZN(n12226) );
  XNOR2_X1 U14670 ( .A(n13183), .B(n12226), .ZN(n12233) );
  NOR2_X1 U14671 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n9235), .ZN(n13362) );
  AOI21_X1 U14672 ( .B1(n13281), .B2(n13706), .A(n13362), .ZN(n12229) );
  NAND2_X1 U14673 ( .A1(n13350), .A2(n12227), .ZN(n12228) );
  OAI211_X1 U14674 ( .C1(n12230), .C2(n13315), .A(n12229), .B(n12228), .ZN(
        n12231) );
  AOI21_X1 U14675 ( .B1(n15318), .B2(n13337), .A(n12231), .ZN(n12232) );
  OAI21_X1 U14676 ( .B1(n12233), .B2(n13352), .A(n12232), .ZN(P3_U3174) );
  NAND2_X1 U14677 ( .A1(n14680), .A2(n12234), .ZN(n12238) );
  AOI21_X1 U14678 ( .B1(n14574), .B2(n12236), .A(n12235), .ZN(n12237) );
  OAI211_X1 U14679 ( .C1(n12239), .C2(n15387), .A(n12238), .B(n12237), .ZN(
        n12247) );
  AND2_X1 U14680 ( .A1(n14517), .A2(n14699), .ZN(n12242) );
  AOI21_X1 U14681 ( .B1(n12654), .B2(n9893), .A(n12242), .ZN(n12303) );
  OAI22_X1 U14682 ( .A1(n12243), .A2(n6667), .B1(n15386), .B2(n14557), .ZN(
        n12244) );
  XNOR2_X1 U14683 ( .A(n12244), .B(n6921), .ZN(n12302) );
  XOR2_X1 U14684 ( .A(n12303), .B(n12302), .Z(n12245) );
  AOI211_X1 U14685 ( .C1(n6717), .C2(n12245), .A(n15392), .B(n15391), .ZN(
        n12246) );
  AOI211_X1 U14686 ( .C1(n12654), .C2(n15397), .A(n12247), .B(n12246), .ZN(
        n12248) );
  INV_X1 U14687 ( .A(n12248), .ZN(P1_U3217) );
  AOI211_X1 U14688 ( .C1(n15672), .C2(n12980), .A(n12250), .B(n12249), .ZN(
        n12254) );
  AOI22_X1 U14689 ( .A1(n12252), .A2(n8998), .B1(P2_REG0_REG_15__SCAN_IN), 
        .B2(n15678), .ZN(n12251) );
  OAI21_X1 U14690 ( .B1(n12254), .B2(n15678), .A(n12251), .ZN(P2_U3475) );
  AOI22_X1 U14691 ( .A1(n12252), .A2(n14277), .B1(P2_REG1_REG_15__SCAN_IN), 
        .B2(n7435), .ZN(n12253) );
  OAI21_X1 U14692 ( .B1(n12254), .B2(n7435), .A(n12253), .ZN(P2_U3514) );
  OAI211_X1 U14693 ( .C1(n12257), .C2(n12256), .A(n12255), .B(n15345), .ZN(
        n12263) );
  OAI22_X1 U14694 ( .A1(n13953), .A2(n12259), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n12258), .ZN(n12260) );
  AOI21_X1 U14695 ( .B1(n12261), .B2(n13944), .A(n12260), .ZN(n12262) );
  OAI211_X1 U14696 ( .C1(n8888), .C2(n13958), .A(n12263), .B(n12262), .ZN(
        P2_U3213) );
  XNOR2_X1 U14697 ( .A(n12264), .B(n12266), .ZN(n12265) );
  OAI222_X1 U14698 ( .A1(n13694), .A2(n13180), .B1(n13696), .B2(n13693), .C1(
        n12265), .C2(n13691), .ZN(n13773) );
  INV_X1 U14699 ( .A(n13773), .ZN(n12271) );
  XNOR2_X1 U14700 ( .A(n12267), .B(n12266), .ZN(n13774) );
  AOI22_X1 U14701 ( .A1(n15735), .A2(P3_REG2_REG_14__SCAN_IN), .B1(n15709), 
        .B2(n13228), .ZN(n12268) );
  OAI21_X1 U14702 ( .B1(n13824), .B2(n13714), .A(n12268), .ZN(n12269) );
  AOI21_X1 U14703 ( .B1(n13774), .B2(n13716), .A(n12269), .ZN(n12270) );
  OAI21_X1 U14704 ( .B1(n12271), .B2(n15735), .A(n12270), .ZN(P3_U3219) );
  NAND2_X1 U14705 ( .A1(n12275), .A2(n11026), .ZN(n12278) );
  AOI22_X1 U14706 ( .A1(n7282), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n12415), 
        .B2(n12276), .ZN(n12277) );
  NAND2_X1 U14707 ( .A1(n12658), .A2(n15385), .ZN(n12279) );
  NAND2_X1 U14708 ( .A1(n15278), .A2(n12279), .ZN(n12810) );
  XNOR2_X1 U14709 ( .A(n12355), .B(n12810), .ZN(n15273) );
  AOI21_X1 U14710 ( .B1(n12280), .B2(n12658), .A(n15488), .ZN(n12281) );
  INV_X1 U14711 ( .A(n12360), .ZN(n15289) );
  NAND2_X1 U14712 ( .A1(n12281), .A2(n15289), .ZN(n15269) );
  INV_X1 U14713 ( .A(n12318), .ZN(n12282) );
  OAI22_X1 U14714 ( .A1(n15093), .A2(n10366), .B1(n12282), .B2(n15058), .ZN(
        n12283) );
  AOI21_X1 U14715 ( .B1(n12658), .B2(n15285), .A(n12283), .ZN(n12284) );
  OAI21_X1 U14716 ( .B1(n15269), .B2(n14994), .A(n12284), .ZN(n12300) );
  INV_X1 U14717 ( .A(n14698), .ZN(n12661) );
  NOR2_X1 U14718 ( .A1(n15398), .A2(n12661), .ZN(n12285) );
  AOI21_X1 U14719 ( .B1(n12287), .B2(n12810), .A(n15481), .ZN(n12298) );
  NAND2_X1 U14720 ( .A1(n14698), .A2(n15001), .ZN(n12296) );
  NAND2_X1 U14721 ( .A1(n12519), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n12294) );
  NAND2_X1 U14722 ( .A1(n9864), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n12293) );
  NAND2_X1 U14723 ( .A1(n12289), .A2(n12288), .ZN(n12290) );
  AND2_X1 U14724 ( .A1(n12337), .A2(n12290), .ZN(n15284) );
  NAND2_X1 U14725 ( .A1(n6677), .A2(n15284), .ZN(n12292) );
  NAND2_X1 U14726 ( .A1(n6683), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n12291) );
  NAND4_X1 U14727 ( .A1(n12294), .A2(n12293), .A3(n12292), .A4(n12291), .ZN(
        n14697) );
  NAND2_X1 U14728 ( .A1(n14697), .A2(n15002), .ZN(n12295) );
  AND2_X1 U14729 ( .A1(n12296), .A2(n12295), .ZN(n12316) );
  INV_X1 U14730 ( .A(n12316), .ZN(n12297) );
  AOI21_X1 U14731 ( .B1(n12298), .B2(n12325), .A(n12297), .ZN(n15270) );
  NOR2_X1 U14732 ( .A1(n15270), .A2(n15067), .ZN(n12299) );
  AOI211_X1 U14733 ( .C1(n15294), .C2(n15273), .A(n12300), .B(n12299), .ZN(
        n12301) );
  INV_X1 U14734 ( .A(n12301), .ZN(P1_U3281) );
  INV_X1 U14735 ( .A(n12302), .ZN(n12304) );
  NOR2_X1 U14736 ( .A1(n12304), .A2(n12303), .ZN(n15390) );
  NAND2_X1 U14737 ( .A1(n15398), .A2(n14511), .ZN(n12306) );
  NAND2_X1 U14738 ( .A1(n14698), .A2(n9893), .ZN(n12305) );
  NAND2_X1 U14739 ( .A1(n12306), .A2(n12305), .ZN(n12307) );
  XNOR2_X1 U14740 ( .A(n12307), .B(n9851), .ZN(n12310) );
  AND2_X1 U14741 ( .A1(n14517), .A2(n14698), .ZN(n12308) );
  AOI21_X1 U14742 ( .B1(n15398), .B2(n9893), .A(n12308), .ZN(n12309) );
  XNOR2_X1 U14743 ( .A(n12310), .B(n12309), .ZN(n15389) );
  OAI22_X1 U14744 ( .A1(n15271), .A2(n14557), .B1(n15385), .B2(n6950), .ZN(
        n14405) );
  OAI22_X1 U14745 ( .A1(n15271), .A2(n6667), .B1(n15385), .B2(n14557), .ZN(
        n12312) );
  XNOR2_X1 U14746 ( .A(n12312), .B(n6921), .ZN(n14406) );
  XOR2_X1 U14747 ( .A(n14405), .B(n14406), .Z(n12313) );
  NAND2_X1 U14748 ( .A1(n12314), .A2(n12313), .ZN(n14408) );
  OAI211_X1 U14749 ( .C1(n12314), .C2(n12313), .A(n14408), .B(n14675), .ZN(
        n12320) );
  OAI22_X1 U14750 ( .A1(n14668), .A2(n12316), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n12315), .ZN(n12317) );
  AOI21_X1 U14751 ( .B1(n14680), .B2(n12318), .A(n12317), .ZN(n12319) );
  OAI211_X1 U14752 ( .C1(n15271), .C2(n14683), .A(n12320), .B(n12319), .ZN(
        P1_U3224) );
  INV_X1 U14753 ( .A(n12468), .ZN(n12323) );
  INV_X1 U14754 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n12469) );
  OAI222_X1 U14755 ( .A1(P1_U3086), .A2(n12321), .B1(n15238), .B2(n12323), 
        .C1(n12469), .C2(n15239), .ZN(P1_U3331) );
  OAI222_X1 U14756 ( .A1(n12861), .A2(n12324), .B1(n14396), .B2(n12323), .C1(
        P2_U3088), .C2(n12322), .ZN(P2_U3303) );
  NAND2_X1 U14757 ( .A1(n12326), .A2(n11026), .ZN(n12330) );
  INV_X1 U14758 ( .A(n12327), .ZN(n12328) );
  AOI22_X1 U14759 ( .A1(n7282), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n12415), 
        .B2(n12328), .ZN(n12329) );
  XNOR2_X1 U14760 ( .A(n15286), .B(n15373), .ZN(n15288) );
  OR2_X1 U14761 ( .A1(n15286), .A2(n15373), .ZN(n12331) );
  NAND2_X1 U14762 ( .A1(n15277), .A2(n12331), .ZN(n15055) );
  NAND2_X1 U14763 ( .A1(n12332), .A2(n11026), .ZN(n12335) );
  AOI22_X1 U14764 ( .A1(n7282), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n12415), 
        .B2(n12333), .ZN(n12334) );
  AND2_X1 U14765 ( .A1(n12337), .A2(n12336), .ZN(n12338) );
  OR2_X1 U14766 ( .A1(n12338), .A2(n12349), .ZN(n15383) );
  INV_X1 U14767 ( .A(n15383), .ZN(n12339) );
  NAND2_X1 U14768 ( .A1(n6677), .A2(n12339), .ZN(n12343) );
  NAND2_X1 U14769 ( .A1(n9864), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n12342) );
  NAND2_X1 U14770 ( .A1(n6683), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n12341) );
  NAND2_X1 U14771 ( .A1(n12519), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n12340) );
  NAND2_X1 U14772 ( .A1(n15380), .A2(n14637), .ZN(n12677) );
  NAND2_X1 U14773 ( .A1(n15055), .A2(n12677), .ZN(n12344) );
  NAND2_X1 U14774 ( .A1(n12344), .A2(n12678), .ZN(n12393) );
  NAND2_X1 U14775 ( .A1(n12345), .A2(n11026), .ZN(n12348) );
  AOI22_X1 U14776 ( .A1(n7282), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n12415), 
        .B2(n12346), .ZN(n12347) );
  NAND2_X1 U14777 ( .A1(n12519), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n12354) );
  NAND2_X1 U14778 ( .A1(n6681), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n12353) );
  NOR2_X1 U14779 ( .A1(n12349), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n12350) );
  NAND2_X1 U14780 ( .A1(n6677), .A2(n6812), .ZN(n12352) );
  NAND2_X1 U14781 ( .A1(n6683), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n12351) );
  NAND2_X1 U14782 ( .A1(n15196), .A2(n15372), .ZN(n12682) );
  NAND2_X1 U14783 ( .A1(n12681), .A2(n12682), .ZN(n12813) );
  XNOR2_X1 U14784 ( .A(n12393), .B(n12392), .ZN(n15202) );
  NOR2_X1 U14785 ( .A1(n15067), .A2(n15481), .ZN(n15090) );
  INV_X1 U14786 ( .A(n15090), .ZN(n14887) );
  NAND2_X1 U14787 ( .A1(n15271), .A2(n15385), .ZN(n12356) );
  NAND2_X1 U14788 ( .A1(n15059), .A2(n15062), .ZN(n15061) );
  NAND2_X1 U14789 ( .A1(n15380), .A2(n14696), .ZN(n12357) );
  OAI21_X1 U14790 ( .B1(n12358), .B2(n12813), .A(n12534), .ZN(n15200) );
  INV_X1 U14791 ( .A(n15196), .ZN(n14684) );
  OR2_X1 U14792 ( .A1(n14684), .A2(n6815), .ZN(n12361) );
  NAND2_X1 U14793 ( .A1(n15045), .A2(n12361), .ZN(n15198) );
  NOR2_X1 U14794 ( .A1(n14994), .A2(n15488), .ZN(n15094) );
  INV_X1 U14795 ( .A(n15094), .ZN(n15034) );
  NOR2_X1 U14796 ( .A1(n15198), .A2(n15034), .ZN(n12371) );
  NAND2_X1 U14797 ( .A1(n12519), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n12367) );
  NAND2_X1 U14798 ( .A1(n9864), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n12366) );
  OR2_X1 U14799 ( .A1(n12362), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n12363) );
  AND2_X1 U14800 ( .A1(n12403), .A2(n12363), .ZN(n15046) );
  NAND2_X1 U14801 ( .A1(n6677), .A2(n15046), .ZN(n12365) );
  NAND2_X1 U14802 ( .A1(n6683), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n12364) );
  NAND4_X1 U14803 ( .A1(n12367), .A2(n12366), .A3(n12365), .A4(n12364), .ZN(
        n14694) );
  INV_X1 U14804 ( .A(n14694), .ZN(n15021) );
  OAI22_X1 U14805 ( .A1(n15021), .A2(n15091), .B1(n14637), .B2(n15069), .ZN(
        n15195) );
  AOI22_X1 U14806 ( .A1(n15195), .A2(n15093), .B1(n6812), .B2(n15283), .ZN(
        n12369) );
  NAND2_X1 U14807 ( .A1(n15067), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n12368) );
  OAI211_X1 U14808 ( .C1(n14684), .C2(n15013), .A(n12369), .B(n12368), .ZN(
        n12370) );
  AOI211_X1 U14809 ( .C1(n15200), .C2(n15294), .A(n12371), .B(n12370), .ZN(
        n12372) );
  OAI21_X1 U14810 ( .B1(n15202), .B2(n14887), .A(n12372), .ZN(P1_U3278) );
  AOI21_X1 U14811 ( .B1(n13281), .B2(n13355), .A(n12373), .ZN(n12376) );
  NAND2_X1 U14812 ( .A1(n13350), .A2(n12374), .ZN(n12375) );
  OAI211_X1 U14813 ( .C1(n12377), .C2(n13315), .A(n12376), .B(n12375), .ZN(
        n12385) );
  INV_X1 U14814 ( .A(n12378), .ZN(n12380) );
  NAND2_X1 U14815 ( .A1(n12380), .A2(n12379), .ZN(n12381) );
  XNOR2_X1 U14816 ( .A(n12382), .B(n12381), .ZN(n12383) );
  NOR2_X1 U14817 ( .A1(n12383), .A2(n13352), .ZN(n12384) );
  AOI211_X1 U14818 ( .C1(n13337), .C2(n15325), .A(n12385), .B(n12384), .ZN(
        n12386) );
  INV_X1 U14819 ( .A(n12386), .ZN(P3_U3164) );
  INV_X1 U14820 ( .A(n12480), .ZN(n12389) );
  OAI222_X1 U14821 ( .A1(P1_U3086), .A2(n12387), .B1(n15238), .B2(n12389), 
        .C1(n12481), .C2(n15239), .ZN(P1_U3330) );
  OAI222_X1 U14822 ( .A1(n12861), .A2(n12390), .B1(n14396), .B2(n12389), .C1(
        P2_U3088), .C2(n12388), .ZN(P2_U3302) );
  AND2_X1 U14823 ( .A1(n15476), .A2(n12391), .ZN(P1_U3085) );
  NAND2_X1 U14824 ( .A1(n12394), .A2(n11026), .ZN(n12397) );
  AOI22_X1 U14825 ( .A1(n7282), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n12415), 
        .B2(n12395), .ZN(n12396) );
  XNOR2_X1 U14826 ( .A(n15192), .B(n14694), .ZN(n15040) );
  INV_X1 U14827 ( .A(n15040), .ZN(n12535) );
  NAND2_X1 U14828 ( .A1(n15192), .A2(n15021), .ZN(n12398) );
  NAND2_X1 U14829 ( .A1(n12399), .A2(n11026), .ZN(n12401) );
  AOI22_X1 U14830 ( .A1(n7282), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n12415), 
        .B2(n14811), .ZN(n12400) );
  NAND2_X1 U14831 ( .A1(n12519), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n12409) );
  NAND2_X1 U14832 ( .A1(n6681), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n12408) );
  NAND2_X1 U14833 ( .A1(n12403), .A2(n12402), .ZN(n12404) );
  AND2_X1 U14834 ( .A1(n12405), .A2(n12404), .ZN(n15028) );
  NAND2_X1 U14835 ( .A1(n6677), .A2(n15028), .ZN(n12407) );
  NAND2_X1 U14836 ( .A1(n6683), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n12406) );
  NAND4_X1 U14837 ( .A1(n12409), .A2(n12408), .A3(n12407), .A4(n12406), .ZN(
        n15000) );
  OR2_X1 U14838 ( .A1(n15032), .A2(n15000), .ZN(n12538) );
  NAND2_X1 U14839 ( .A1(n15032), .A2(n15000), .ZN(n12540) );
  NAND2_X1 U14840 ( .A1(n12538), .A2(n12540), .ZN(n15018) );
  INV_X1 U14841 ( .A(n15018), .ZN(n15019) );
  NAND2_X1 U14842 ( .A1(n15184), .A2(n15000), .ZN(n12410) );
  NAND2_X1 U14843 ( .A1(n12411), .A2(n11026), .ZN(n12413) );
  AOI22_X1 U14844 ( .A1(n7282), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n12415), 
        .B2(n14828), .ZN(n12412) );
  XNOR2_X1 U14845 ( .A(n15180), .B(n15022), .ZN(n12814) );
  INV_X1 U14846 ( .A(n15022), .ZN(n14988) );
  NAND2_X1 U14847 ( .A1(n12414), .A2(n11026), .ZN(n12417) );
  AOI22_X1 U14848 ( .A1(n7282), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n15048), 
        .B2(n12415), .ZN(n12416) );
  NAND2_X1 U14849 ( .A1(n12418), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n12429) );
  OR2_X1 U14850 ( .A1(n12418), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n12419) );
  NAND2_X1 U14851 ( .A1(n12429), .A2(n12419), .ZN(n14990) );
  NAND2_X1 U14852 ( .A1(n9864), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n12421) );
  NAND2_X1 U14853 ( .A1(n12519), .A2(P1_REG1_REG_19__SCAN_IN), .ZN(n12420) );
  AND2_X1 U14854 ( .A1(n12421), .A2(n12420), .ZN(n12423) );
  NAND2_X1 U14855 ( .A1(n6683), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n12422) );
  OAI211_X1 U14856 ( .C1(n14990), .C2(n12451), .A(n12423), .B(n12422), .ZN(
        n15003) );
  XNOR2_X1 U14857 ( .A(n14448), .B(n15003), .ZN(n14985) );
  INV_X1 U14858 ( .A(n14985), .ZN(n12815) );
  INV_X1 U14859 ( .A(n15003), .ZN(n14657) );
  NAND2_X1 U14860 ( .A1(n14448), .A2(n14657), .ZN(n12424) );
  NAND2_X1 U14861 ( .A1(n12425), .A2(n11026), .ZN(n12428) );
  OR2_X1 U14862 ( .A1(n9888), .A2(n12426), .ZN(n12427) );
  INV_X1 U14863 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n14628) );
  NAND2_X1 U14864 ( .A1(n12429), .A2(n14628), .ZN(n12430) );
  NAND2_X1 U14865 ( .A1(n12439), .A2(n12430), .ZN(n14972) );
  OR2_X1 U14866 ( .A1(n14972), .A2(n12451), .ZN(n12433) );
  AOI22_X1 U14867 ( .A1(n12519), .A2(P1_REG1_REG_20__SCAN_IN), .B1(n6681), 
        .B2(P1_REG0_REG_20__SCAN_IN), .ZN(n12432) );
  NAND2_X1 U14868 ( .A1(n6683), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n12431) );
  INV_X1 U14869 ( .A(n14572), .ZN(n14989) );
  XNOR2_X1 U14870 ( .A(n14977), .B(n14989), .ZN(n14979) );
  NAND2_X1 U14871 ( .A1(n15166), .A2(n14989), .ZN(n12434) );
  NAND2_X2 U14872 ( .A1(n14967), .A2(n12434), .ZN(n14953) );
  NAND2_X1 U14873 ( .A1(n12435), .A2(n11026), .ZN(n12437) );
  OR2_X1 U14874 ( .A1(n9888), .A2(n9370), .ZN(n12436) );
  INV_X1 U14875 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n12438) );
  AND2_X1 U14876 ( .A1(n12439), .A2(n12438), .ZN(n12440) );
  OR2_X1 U14877 ( .A1(n12449), .A2(n12440), .ZN(n14956) );
  INV_X1 U14878 ( .A(P1_REG2_REG_21__SCAN_IN), .ZN(n12443) );
  NAND2_X1 U14879 ( .A1(n12519), .A2(P1_REG1_REG_21__SCAN_IN), .ZN(n12442) );
  NAND2_X1 U14880 ( .A1(n6681), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n12441) );
  OAI211_X1 U14881 ( .C1(n12443), .C2(n6684), .A(n12442), .B(n12441), .ZN(
        n12444) );
  INV_X1 U14882 ( .A(n12444), .ZN(n12445) );
  NAND2_X1 U14883 ( .A1(n15158), .A2(n14969), .ZN(n12446) );
  NAND2_X1 U14884 ( .A1(n12545), .A2(n12446), .ZN(n14963) );
  INV_X1 U14885 ( .A(n14969), .ZN(n14941) );
  OR2_X1 U14886 ( .A1(n8732), .A2(n9950), .ZN(n12447) );
  XNOR2_X1 U14887 ( .A(n12447), .B(P2_DATAO_REG_22__SCAN_IN), .ZN(n15243) );
  OR2_X1 U14888 ( .A1(n12449), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n12450) );
  NAND2_X1 U14889 ( .A1(n12449), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n12462) );
  NAND2_X1 U14890 ( .A1(n12450), .A2(n12462), .ZN(n14948) );
  OR2_X1 U14891 ( .A1(n14948), .A2(n12451), .ZN(n12456) );
  INV_X1 U14892 ( .A(P1_REG2_REG_22__SCAN_IN), .ZN(n14947) );
  NAND2_X1 U14893 ( .A1(n12519), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n12453) );
  NAND2_X1 U14894 ( .A1(n9864), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n12452) );
  OAI211_X1 U14895 ( .C1(n14947), .C2(n6684), .A(n12453), .B(n12452), .ZN(
        n12454) );
  INV_X1 U14896 ( .A(n12454), .ZN(n12455) );
  NAND2_X1 U14897 ( .A1(n12456), .A2(n12455), .ZN(n14693) );
  INV_X1 U14898 ( .A(n14693), .ZN(n14573) );
  XNOR2_X1 U14899 ( .A(n14946), .B(n14573), .ZN(n14936) );
  NAND2_X1 U14900 ( .A1(n12457), .A2(n11026), .ZN(n12460) );
  OR2_X1 U14901 ( .A1(n9888), .A2(n12458), .ZN(n12459) );
  NAND2_X1 U14902 ( .A1(n12519), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n12466) );
  NAND2_X1 U14903 ( .A1(n6681), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n12465) );
  INV_X1 U14904 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n14539) );
  INV_X1 U14905 ( .A(n12462), .ZN(n12461) );
  NAND2_X1 U14906 ( .A1(n12461), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n12473) );
  AOI21_X1 U14907 ( .B1(n14539), .B2(n12462), .A(n12472), .ZN(n14930) );
  NAND2_X1 U14908 ( .A1(n6677), .A2(n14930), .ZN(n12464) );
  NAND2_X1 U14909 ( .A1(n6683), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n12463) );
  NAND4_X1 U14910 ( .A1(n12466), .A2(n12465), .A3(n12464), .A4(n12463), .ZN(
        n14692) );
  XNOR2_X1 U14911 ( .A(n15148), .B(n14942), .ZN(n14921) );
  NAND2_X1 U14912 ( .A1(n15148), .A2(n14942), .ZN(n12467) );
  NAND2_X1 U14913 ( .A1(n14925), .A2(n12467), .ZN(n14909) );
  NAND2_X1 U14914 ( .A1(n12468), .A2(n11026), .ZN(n12471) );
  OR2_X1 U14915 ( .A1(n9888), .A2(n12469), .ZN(n12470) );
  NAND2_X1 U14916 ( .A1(n12519), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n12477) );
  NAND2_X1 U14917 ( .A1(n6681), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n12476) );
  INV_X1 U14918 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n14620) );
  NAND2_X1 U14919 ( .A1(n12472), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n12485) );
  INV_X1 U14920 ( .A(n12485), .ZN(n12484) );
  AOI21_X1 U14921 ( .B1(n14620), .B2(n12473), .A(n12484), .ZN(n14914) );
  NAND2_X1 U14922 ( .A1(n6677), .A2(n14914), .ZN(n12475) );
  NAND2_X1 U14923 ( .A1(n6683), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n12474) );
  NAND4_X1 U14924 ( .A1(n12477), .A2(n12476), .A3(n12475), .A4(n12474), .ZN(
        n14691) );
  INV_X1 U14925 ( .A(n14691), .ZN(n12478) );
  XNOR2_X1 U14926 ( .A(n15141), .B(n12478), .ZN(n14910) );
  OR2_X2 U14927 ( .A1(n14909), .A2(n14910), .ZN(n14907) );
  OR2_X1 U14928 ( .A1(n15141), .A2(n12478), .ZN(n12479) );
  NAND2_X1 U14929 ( .A1(n14907), .A2(n12479), .ZN(n14888) );
  NAND2_X1 U14930 ( .A1(n12480), .A2(n11026), .ZN(n12483) );
  OR2_X1 U14931 ( .A1(n9888), .A2(n12481), .ZN(n12482) );
  NAND2_X2 U14932 ( .A1(n12483), .A2(n12482), .ZN(n15133) );
  NAND2_X1 U14933 ( .A1(n12519), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n12489) );
  NAND2_X1 U14934 ( .A1(n6680), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n12488) );
  INV_X1 U14935 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n14588) );
  NAND2_X1 U14936 ( .A1(n12484), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n12495) );
  INV_X1 U14937 ( .A(n12495), .ZN(n12494) );
  AOI21_X1 U14938 ( .B1(n14588), .B2(n12485), .A(n12494), .ZN(n14890) );
  NAND2_X1 U14939 ( .A1(n6677), .A2(n14890), .ZN(n12487) );
  NAND2_X1 U14940 ( .A1(n6683), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n12486) );
  NAND4_X1 U14941 ( .A1(n12489), .A2(n12488), .A3(n12487), .A4(n12486), .ZN(
        n14690) );
  INV_X1 U14942 ( .A(n14690), .ZN(n12490) );
  XNOR2_X1 U14943 ( .A(n15133), .B(n12490), .ZN(n12818) );
  NAND2_X1 U14944 ( .A1(n15133), .A2(n12490), .ZN(n12491) );
  NAND2_X1 U14945 ( .A1(n14393), .A2(n11026), .ZN(n12493) );
  OR2_X1 U14946 ( .A1(n9888), .A2(n15240), .ZN(n12492) );
  NAND2_X1 U14947 ( .A1(n6681), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n12499) );
  NAND2_X1 U14948 ( .A1(n6683), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n12498) );
  INV_X1 U14949 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n14667) );
  NAND2_X1 U14950 ( .A1(n12494), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n12504) );
  INV_X1 U14951 ( .A(n12504), .ZN(n12506) );
  AOI21_X1 U14952 ( .B1(n14667), .B2(n12495), .A(n12506), .ZN(n14880) );
  NAND2_X1 U14953 ( .A1(n6677), .A2(n14880), .ZN(n12497) );
  NAND2_X1 U14954 ( .A1(n12519), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n12496) );
  NAND4_X1 U14955 ( .A1(n12499), .A2(n12498), .A3(n12497), .A4(n12496), .ZN(
        n14689) );
  INV_X1 U14956 ( .A(n14689), .ZN(n12500) );
  OR2_X1 U14957 ( .A1(n14516), .A2(n12500), .ZN(n12501) );
  NAND2_X1 U14958 ( .A1(n12555), .A2(n11026), .ZN(n12503) );
  OR2_X1 U14959 ( .A1(n9888), .A2(n7339), .ZN(n12502) );
  NAND2_X1 U14960 ( .A1(n12519), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n12511) );
  NAND2_X1 U14961 ( .A1(n9864), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n12510) );
  INV_X1 U14962 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n12505) );
  NAND2_X1 U14963 ( .A1(n12505), .A2(n12504), .ZN(n12507) );
  NAND2_X1 U14964 ( .A1(P1_REG3_REG_27__SCAN_IN), .A2(n12506), .ZN(n12521) );
  NAND2_X1 U14965 ( .A1(n6677), .A2(n14869), .ZN(n12509) );
  NAND2_X1 U14966 ( .A1(n6683), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n12508) );
  NAND2_X1 U14967 ( .A1(n15235), .A2(n11026), .ZN(n12513) );
  OR2_X1 U14968 ( .A1(n9888), .A2(n15236), .ZN(n12512) );
  NAND2_X1 U14969 ( .A1(n12519), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n12517) );
  NAND2_X1 U14970 ( .A1(n6681), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n12516) );
  XNOR2_X1 U14971 ( .A(n12521), .B(P1_REG3_REG_28__SCAN_IN), .ZN(n14566) );
  NAND2_X1 U14972 ( .A1(n6677), .A2(n14566), .ZN(n12515) );
  NAND2_X1 U14973 ( .A1(n6683), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n12514) );
  NAND4_X1 U14974 ( .A1(n12517), .A2(n12516), .A3(n12515), .A4(n12514), .ZN(
        n14687) );
  NAND2_X1 U14975 ( .A1(n15113), .A2(n14687), .ZN(n12569) );
  OR2_X1 U14976 ( .A1(n15113), .A2(n14687), .ZN(n12518) );
  NAND2_X1 U14977 ( .A1(n12569), .A2(n12518), .ZN(n12821) );
  NAND2_X1 U14978 ( .A1(n12519), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n12525) );
  NAND2_X1 U14979 ( .A1(n9864), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n12524) );
  INV_X1 U14980 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n12520) );
  NOR2_X1 U14981 ( .A1(n12521), .A2(n12520), .ZN(n12582) );
  NAND2_X1 U14982 ( .A1(n6677), .A2(n12582), .ZN(n12523) );
  NAND2_X1 U14983 ( .A1(n6683), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n12522) );
  INV_X1 U14984 ( .A(n14562), .ZN(n14686) );
  NAND2_X1 U14985 ( .A1(n14686), .A2(n15002), .ZN(n12527) );
  NAND2_X1 U14986 ( .A1(n14688), .A2(n15001), .ZN(n12526) );
  NOR2_X2 U14987 ( .A1(n14913), .A2(n15133), .ZN(n14899) );
  AOI211_X1 U14988 ( .C1(n15113), .C2(n14867), .A(n15488), .B(n12577), .ZN(
        n15112) );
  AOI22_X1 U14989 ( .A1(n15067), .A2(P1_REG2_REG_28__SCAN_IN), .B1(n14566), 
        .B2(n15283), .ZN(n12531) );
  OAI21_X1 U14990 ( .B1(n14563), .B2(n15013), .A(n12531), .ZN(n12532) );
  AOI21_X1 U14991 ( .B1(n15112), .B2(n15293), .A(n12532), .ZN(n12554) );
  INV_X1 U14992 ( .A(n15372), .ZN(n14695) );
  OR2_X1 U14993 ( .A1(n15196), .A2(n14695), .ZN(n12533) );
  OR2_X1 U14994 ( .A1(n15192), .A2(n14694), .ZN(n12536) );
  INV_X1 U14995 ( .A(n12538), .ZN(n12539) );
  AND2_X1 U14996 ( .A1(n15180), .A2(n14988), .ZN(n12710) );
  OR2_X1 U14997 ( .A1(n15180), .A2(n14988), .ZN(n12709) );
  NAND2_X1 U14998 ( .A1(n14983), .A2(n12815), .ZN(n12542) );
  OR2_X1 U14999 ( .A1(n14448), .A2(n15003), .ZN(n12541) );
  OR2_X1 U15000 ( .A1(n15166), .A2(n14572), .ZN(n12544) );
  INV_X1 U15001 ( .A(n14936), .ZN(n14938) );
  NAND2_X1 U15002 ( .A1(n14922), .A2(n14921), .ZN(n14920) );
  NAND2_X1 U15003 ( .A1(n15148), .A2(n14692), .ZN(n12546) );
  NAND2_X1 U15004 ( .A1(n14920), .A2(n12546), .ZN(n14904) );
  INV_X1 U15005 ( .A(n14910), .ZN(n12547) );
  OR2_X1 U15006 ( .A1(n15141), .A2(n14691), .ZN(n12548) );
  XNOR2_X1 U15007 ( .A(n14516), .B(n14689), .ZN(n12819) );
  NAND2_X1 U15008 ( .A1(n14877), .A2(n14876), .ZN(n14875) );
  NAND2_X1 U15009 ( .A1(n14516), .A2(n14689), .ZN(n12549) );
  OR2_X1 U15010 ( .A1(n14866), .A2(n14688), .ZN(n12550) );
  INV_X1 U15011 ( .A(n12821), .ZN(n12551) );
  NAND2_X1 U15012 ( .A1(n12552), .A2(n12821), .ZN(n15111) );
  NAND3_X1 U15013 ( .A1(n12570), .A2(n15294), .A3(n15111), .ZN(n12553) );
  OAI211_X1 U15014 ( .C1(n15115), .C2(n15067), .A(n12554), .B(n12553), .ZN(
        P1_U3265) );
  INV_X1 U15015 ( .A(n12555), .ZN(n12568) );
  OAI222_X1 U15016 ( .A1(n14718), .A2(P1_U3086), .B1(n15238), .B2(n12568), 
        .C1(n7339), .C2(n15239), .ZN(P1_U3328) );
  INV_X1 U15017 ( .A(n12558), .ZN(n12559) );
  NAND2_X1 U15018 ( .A1(n12559), .A2(n13841), .ZN(n12560) );
  MUX2_X1 U15019 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(P1_DATAO_REG_30__SCAN_IN), 
        .S(n9950), .Z(n12561) );
  NAND2_X1 U15020 ( .A1(n12561), .A2(SI_30_), .ZN(n12778) );
  OAI21_X1 U15021 ( .B1(n12561), .B2(SI_30_), .A(n12778), .ZN(n12562) );
  OAI222_X1 U15022 ( .A1(n14396), .A2(n13093), .B1(n12564), .B2(P2_U3088), 
        .C1(n9487), .C2(n12861), .ZN(P2_U3297) );
  OAI222_X1 U15023 ( .A1(n12861), .A2(n12566), .B1(n14396), .B2(n12565), .C1(
        P2_U3088), .C2(n8859), .ZN(P2_U3308) );
  OAI222_X1 U15024 ( .A1(n14396), .A2(n12568), .B1(n8938), .B2(P2_U3088), .C1(
        n12567), .C2(n12861), .ZN(P2_U3300) );
  NOR2_X1 U15025 ( .A1(n9888), .A2(n15232), .ZN(n12571) );
  INV_X1 U15026 ( .A(n12759), .ZN(n15104) );
  XNOR2_X1 U15027 ( .A(n15104), .B(n14562), .ZN(n12793) );
  NOR2_X1 U15028 ( .A1(n14563), .A2(n14687), .ZN(n12574) );
  INV_X1 U15029 ( .A(n14687), .ZN(n14556) );
  XNOR2_X1 U15030 ( .A(n12576), .B(n12793), .ZN(n15109) );
  OAI211_X1 U15031 ( .C1(n12759), .C2(n12577), .A(n15291), .B(n14851), .ZN(
        n15108) );
  NOR2_X1 U15032 ( .A1(n15108), .A2(n14994), .ZN(n12589) );
  NAND2_X1 U15033 ( .A1(n12519), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n12580) );
  NAND2_X1 U15034 ( .A1(n6683), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n12579) );
  NAND2_X1 U15035 ( .A1(n9864), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n12578) );
  AND3_X1 U15036 ( .A1(n12580), .A2(n12579), .A3(n12578), .ZN(n12769) );
  INV_X1 U15037 ( .A(n12769), .ZN(n14685) );
  AOI21_X1 U15038 ( .B1(n12581), .B2(P1_B_REG_SCAN_IN), .A(n15091), .ZN(n14847) );
  NAND2_X1 U15039 ( .A1(n14685), .A2(n14847), .ZN(n15105) );
  INV_X1 U15040 ( .A(n12582), .ZN(n12583) );
  OAI22_X1 U15041 ( .A1(n15105), .A2(n12584), .B1(n12583), .B2(n15058), .ZN(
        n12586) );
  NAND2_X1 U15042 ( .A1(n14687), .A2(n15001), .ZN(n15106) );
  NOR2_X1 U15043 ( .A1(n15067), .A2(n15106), .ZN(n12585) );
  AOI211_X1 U15044 ( .C1(n15067), .C2(P1_REG2_REG_29__SCAN_IN), .A(n12586), 
        .B(n12585), .ZN(n12587) );
  OAI21_X1 U15045 ( .B1(n12759), .B2(n15013), .A(n12587), .ZN(n12588) );
  AOI211_X1 U15046 ( .C1(n15109), .C2(n15090), .A(n12589), .B(n12588), .ZN(
        n12590) );
  OAI21_X1 U15047 ( .B1(n15110), .B2(n15063), .A(n12590), .ZN(P1_U3356) );
  NAND2_X1 U15048 ( .A1(n14707), .A2(n12591), .ZN(n12796) );
  NAND2_X1 U15049 ( .A1(n12796), .A2(n12592), .ZN(n12595) );
  MUX2_X1 U15050 ( .A(n12770), .B(n12594), .S(n12767), .Z(n12603) );
  NAND3_X1 U15051 ( .A1(n12595), .A2(n12795), .A3(n6674), .ZN(n12596) );
  NAND2_X1 U15052 ( .A1(n12596), .A2(n12597), .ZN(n12600) );
  INV_X1 U15053 ( .A(n12597), .ZN(n12598) );
  NAND2_X1 U15054 ( .A1(n12598), .A2(n6674), .ZN(n12599) );
  NAND2_X1 U15055 ( .A1(n12600), .A2(n12599), .ZN(n12607) );
  INV_X1 U15056 ( .A(n12795), .ZN(n12601) );
  NAND3_X1 U15057 ( .A1(n12601), .A2(n12789), .A3(n12602), .ZN(n12606) );
  INV_X1 U15058 ( .A(n12602), .ZN(n12604) );
  NAND2_X1 U15059 ( .A1(n12604), .A2(n6674), .ZN(n12605) );
  NAND2_X1 U15060 ( .A1(n12612), .A2(n12608), .ZN(n12611) );
  MUX2_X1 U15061 ( .A(n10689), .B(n6669), .S(n6674), .Z(n12610) );
  INV_X1 U15062 ( .A(n12612), .ZN(n12615) );
  MUX2_X1 U15063 ( .A(n12618), .B(n12617), .S(n6674), .Z(n12619) );
  MUX2_X1 U15064 ( .A(n14705), .B(n12620), .S(n6674), .Z(n12624) );
  NAND2_X1 U15065 ( .A1(n12623), .A2(n12624), .ZN(n12622) );
  NAND2_X1 U15066 ( .A1(n12622), .A2(n12621), .ZN(n12628) );
  INV_X1 U15067 ( .A(n12623), .ZN(n12626) );
  INV_X1 U15068 ( .A(n12624), .ZN(n12625) );
  NAND2_X1 U15069 ( .A1(n12626), .A2(n12625), .ZN(n12627) );
  MUX2_X1 U15070 ( .A(n14704), .B(n12629), .S(n6674), .Z(n12630) );
  INV_X1 U15071 ( .A(n12631), .ZN(n12632) );
  MUX2_X1 U15072 ( .A(n14703), .B(n12633), .S(n6674), .Z(n12636) );
  MUX2_X1 U15073 ( .A(n14702), .B(n12637), .S(n6674), .Z(n12638) );
  INV_X1 U15074 ( .A(n12639), .ZN(n12640) );
  MUX2_X1 U15075 ( .A(n14701), .B(n12641), .S(n6674), .Z(n12645) );
  NAND2_X1 U15076 ( .A1(n12644), .A2(n12645), .ZN(n12643) );
  NAND2_X1 U15077 ( .A1(n12643), .A2(n12642), .ZN(n12649) );
  INV_X1 U15078 ( .A(n12644), .ZN(n12647) );
  INV_X1 U15079 ( .A(n12645), .ZN(n12646) );
  NAND2_X1 U15080 ( .A1(n12647), .A2(n12646), .ZN(n12648) );
  NAND2_X1 U15081 ( .A1(n12649), .A2(n12648), .ZN(n12652) );
  MUX2_X1 U15082 ( .A(n14700), .B(n12650), .S(n6674), .Z(n12651) );
  MUX2_X1 U15083 ( .A(n14699), .B(n12654), .S(n6674), .Z(n12656) );
  MUX2_X1 U15084 ( .A(n14699), .B(n12654), .S(n12789), .Z(n12655) );
  INV_X1 U15085 ( .A(n12656), .ZN(n12657) );
  MUX2_X1 U15086 ( .A(n14698), .B(n15398), .S(n12789), .Z(n12663) );
  MUX2_X1 U15087 ( .A(n15385), .B(n15271), .S(n6674), .Z(n12669) );
  MUX2_X1 U15088 ( .A(n12659), .B(n12658), .S(n12789), .Z(n12668) );
  OAI22_X1 U15089 ( .A1(n12664), .A2(n12663), .B1(n12669), .B2(n12668), .ZN(
        n12660) );
  INV_X1 U15090 ( .A(n12660), .ZN(n12667) );
  MUX2_X1 U15091 ( .A(n12661), .B(n15409), .S(n6674), .Z(n12662) );
  AOI21_X1 U15092 ( .B1(n12664), .B2(n12663), .A(n12662), .ZN(n12665) );
  INV_X1 U15093 ( .A(n12665), .ZN(n12666) );
  NAND2_X1 U15094 ( .A1(n12669), .A2(n12668), .ZN(n12672) );
  MUX2_X1 U15095 ( .A(n14697), .B(n15286), .S(n12789), .Z(n12675) );
  NAND2_X1 U15096 ( .A1(n15373), .A2(n12789), .ZN(n12670) );
  OAI21_X1 U15097 ( .B1(n15286), .B2(n12789), .A(n12670), .ZN(n12676) );
  OAI211_X1 U15098 ( .C1(n12675), .C2(n12676), .A(n12678), .B(n12677), .ZN(
        n12671) );
  AND2_X1 U15099 ( .A1(n14696), .A2(n6674), .ZN(n12674) );
  OAI21_X1 U15100 ( .B1(n6674), .B2(n14696), .A(n15380), .ZN(n12673) );
  OAI21_X1 U15101 ( .B1(n12674), .B2(n15380), .A(n12673), .ZN(n12680) );
  NAND4_X1 U15102 ( .A1(n12678), .A2(n12677), .A3(n12676), .A4(n12675), .ZN(
        n12679) );
  NAND4_X1 U15103 ( .A1(n12681), .A2(n12682), .A3(n12680), .A4(n12679), .ZN(
        n12684) );
  MUX2_X1 U15104 ( .A(n12682), .B(n12681), .S(n12789), .Z(n12683) );
  MUX2_X1 U15105 ( .A(n14694), .B(n15192), .S(n6674), .Z(n12701) );
  NAND2_X1 U15106 ( .A1(n12701), .A2(n15000), .ZN(n12685) );
  NAND2_X1 U15107 ( .A1(n15021), .A2(n6674), .ZN(n12698) );
  AOI21_X1 U15108 ( .B1(n12685), .B2(n12698), .A(n15184), .ZN(n12690) );
  INV_X1 U15109 ( .A(n15000), .ZN(n14436) );
  NAND2_X1 U15110 ( .A1(n12701), .A2(n14436), .ZN(n12686) );
  OR2_X1 U15111 ( .A1(n15192), .A2(n6674), .ZN(n12692) );
  AOI21_X1 U15112 ( .B1(n12686), .B2(n12692), .A(n15032), .ZN(n12689) );
  NAND2_X1 U15113 ( .A1(n15000), .A2(n12789), .ZN(n12694) );
  OR2_X1 U15114 ( .A1(n15192), .A2(n12694), .ZN(n12688) );
  NOR2_X1 U15115 ( .A1(n15000), .A2(n12789), .ZN(n12699) );
  NAND2_X1 U15116 ( .A1(n12699), .A2(n15021), .ZN(n12687) );
  NAND2_X1 U15117 ( .A1(n12688), .A2(n12687), .ZN(n12696) );
  OR3_X1 U15118 ( .A1(n12690), .A2(n12689), .A3(n12696), .ZN(n12691) );
  INV_X1 U15119 ( .A(n12692), .ZN(n12693) );
  NAND2_X1 U15120 ( .A1(n12701), .A2(n12693), .ZN(n12695) );
  NAND2_X1 U15121 ( .A1(n12695), .A2(n12694), .ZN(n12697) );
  AOI22_X1 U15122 ( .A1(n12697), .A2(n15184), .B1(n12701), .B2(n12696), .ZN(
        n12705) );
  INV_X1 U15123 ( .A(n12698), .ZN(n12700) );
  AOI21_X1 U15124 ( .B1(n12701), .B2(n12700), .A(n12699), .ZN(n12702) );
  MUX2_X1 U15125 ( .A(n15022), .B(n15014), .S(n12789), .Z(n12708) );
  AOI21_X1 U15126 ( .B1(n12711), .B2(n12710), .A(n12815), .ZN(n12712) );
  NAND2_X1 U15127 ( .A1(n12713), .A2(n12712), .ZN(n12717) );
  NAND2_X1 U15128 ( .A1(n15003), .A2(n6674), .ZN(n12715) );
  NAND2_X1 U15129 ( .A1(n14657), .A2(n12789), .ZN(n12714) );
  MUX2_X1 U15130 ( .A(n12715), .B(n12714), .S(n14448), .Z(n12716) );
  NAND2_X1 U15131 ( .A1(n12717), .A2(n12716), .ZN(n12720) );
  MUX2_X1 U15132 ( .A(n14572), .B(n15166), .S(n6674), .Z(n12719) );
  MUX2_X1 U15133 ( .A(n14989), .B(n14977), .S(n12789), .Z(n12718) );
  NAND2_X1 U15134 ( .A1(n12720), .A2(n12719), .ZN(n12721) );
  MUX2_X1 U15135 ( .A(n14969), .B(n15158), .S(n6674), .Z(n12723) );
  INV_X1 U15136 ( .A(n12724), .ZN(n12725) );
  MUX2_X1 U15137 ( .A(n14693), .B(n15154), .S(n6674), .Z(n12728) );
  MUX2_X1 U15138 ( .A(n14693), .B(n15154), .S(n12789), .Z(n12726) );
  MUX2_X1 U15139 ( .A(n14692), .B(n15148), .S(n6674), .Z(n12729) );
  INV_X1 U15140 ( .A(n12730), .ZN(n12731) );
  MUX2_X1 U15141 ( .A(n14691), .B(n15141), .S(n6674), .Z(n12735) );
  NAND2_X1 U15142 ( .A1(n12734), .A2(n12735), .ZN(n12733) );
  MUX2_X1 U15143 ( .A(n14691), .B(n15141), .S(n12789), .Z(n12732) );
  INV_X1 U15144 ( .A(n12734), .ZN(n12737) );
  INV_X1 U15145 ( .A(n12735), .ZN(n12736) );
  NAND2_X1 U15146 ( .A1(n12744), .A2(n12743), .ZN(n12738) );
  NAND2_X1 U15147 ( .A1(n12738), .A2(n12741), .ZN(n12740) );
  MUX2_X1 U15148 ( .A(n14690), .B(n15133), .S(n6674), .Z(n12739) );
  NAND2_X1 U15149 ( .A1(n12740), .A2(n12739), .ZN(n12747) );
  INV_X1 U15150 ( .A(n12741), .ZN(n12742) );
  AND2_X1 U15151 ( .A1(n12743), .A2(n12742), .ZN(n12745) );
  NAND2_X1 U15152 ( .A1(n12745), .A2(n12744), .ZN(n12746) );
  MUX2_X1 U15153 ( .A(n14689), .B(n14516), .S(n6674), .Z(n12749) );
  INV_X1 U15154 ( .A(n12749), .ZN(n12750) );
  MUX2_X1 U15155 ( .A(n14688), .B(n14866), .S(n6674), .Z(n12751) );
  MUX2_X1 U15156 ( .A(n14687), .B(n15113), .S(n6674), .Z(n12754) );
  NAND2_X1 U15157 ( .A1(n12753), .A2(n12754), .ZN(n12758) );
  INV_X1 U15158 ( .A(n12753), .ZN(n12756) );
  INV_X1 U15159 ( .A(n12754), .ZN(n12755) );
  MUX2_X1 U15160 ( .A(n14562), .B(n12759), .S(n12789), .Z(n12760) );
  MUX2_X1 U15161 ( .A(n14562), .B(n12759), .S(n6674), .Z(n12761) );
  INV_X1 U15162 ( .A(n12774), .ZN(n12777) );
  OR2_X1 U15163 ( .A1(n9888), .A2(n12862), .ZN(n12762) );
  INV_X1 U15164 ( .A(P1_REG2_REG_31__SCAN_IN), .ZN(n12766) );
  NAND2_X1 U15165 ( .A1(n12519), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n12765) );
  NAND2_X1 U15166 ( .A1(n6680), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n12764) );
  OAI211_X1 U15167 ( .C1(n6684), .C2(n12766), .A(n12765), .B(n12764), .ZN(
        n14848) );
  AOI22_X1 U15168 ( .A1(n14848), .A2(n12789), .B1(n12767), .B2(n12788), .ZN(
        n12768) );
  OAI22_X1 U15169 ( .A1(n15103), .A2(n12789), .B1(n12769), .B2(n12768), .ZN(
        n12773) );
  INV_X1 U15170 ( .A(n12773), .ZN(n12776) );
  OAI21_X1 U15171 ( .B1(n14848), .B2(n12770), .A(n14685), .ZN(n12771) );
  MUX2_X1 U15172 ( .A(n15103), .B(n12771), .S(n6674), .Z(n12772) );
  INV_X1 U15173 ( .A(n12792), .ZN(n12839) );
  MUX2_X1 U15174 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n9950), .Z(n12779) );
  XNOR2_X1 U15175 ( .A(n12779), .B(SI_31_), .ZN(n12780) );
  OR2_X1 U15176 ( .A1(n9888), .A2(n10136), .ZN(n12782) );
  NAND2_X1 U15177 ( .A1(n12784), .A2(n12783), .ZN(n12786) );
  AND2_X1 U15178 ( .A1(n12786), .A2(n12785), .ZN(n12791) );
  INV_X1 U15179 ( .A(n12791), .ZN(n12826) );
  AND2_X1 U15180 ( .A1(n12788), .A2(n12787), .ZN(n12828) );
  INV_X1 U15181 ( .A(n12828), .ZN(n12835) );
  NAND2_X1 U15182 ( .A1(n12826), .A2(n12835), .ZN(n12825) );
  NAND2_X1 U15183 ( .A1(n14844), .A2(n12789), .ZN(n12833) );
  NOR2_X1 U15184 ( .A1(n12833), .A2(n14848), .ZN(n12790) );
  XNOR2_X1 U15185 ( .A(n14844), .B(n14848), .ZN(n12823) );
  NAND3_X1 U15186 ( .A1(n12792), .A2(n12823), .A3(n12791), .ZN(n12836) );
  INV_X1 U15187 ( .A(n15103), .ZN(n14843) );
  INV_X1 U15188 ( .A(n12793), .ZN(n12822) );
  NAND2_X1 U15189 ( .A1(n12796), .A2(n12795), .ZN(n15479) );
  NOR4_X1 U15190 ( .A1(n12794), .A2(n7055), .A3(n12797), .A4(n15479), .ZN(
        n12799) );
  NAND2_X1 U15191 ( .A1(n12799), .A2(n12798), .ZN(n12802) );
  NOR4_X1 U15192 ( .A1(n12803), .A2(n12802), .A3(n12801), .A4(n12800), .ZN(
        n12806) );
  NAND4_X1 U15193 ( .A1(n12807), .A2(n12806), .A3(n12805), .A4(n12804), .ZN(
        n12808) );
  NOR4_X1 U15194 ( .A1(n12810), .A2(n15288), .A3(n12809), .A4(n12808), .ZN(
        n12811) );
  NAND4_X1 U15195 ( .A1(n15060), .A2(n12811), .A3(n15018), .A4(n15040), .ZN(
        n12812) );
  NOR4_X1 U15196 ( .A1(n12815), .A2(n12814), .A3(n12813), .A4(n12812), .ZN(
        n12816) );
  NAND4_X1 U15197 ( .A1(n14936), .A2(n12816), .A3(n14963), .A4(n14979), .ZN(
        n12817) );
  NOR4_X1 U15198 ( .A1(n12818), .A2(n14910), .A3(n14921), .A4(n12817), .ZN(
        n12820) );
  NOR3_X1 U15199 ( .A1(n15100), .A2(n14848), .A3(n12825), .ZN(n12834) );
  NOR3_X1 U15200 ( .A1(n12833), .A2(n14848), .A3(n12826), .ZN(n12832) );
  INV_X1 U15201 ( .A(n14848), .ZN(n12829) );
  NOR4_X1 U15202 ( .A1(n12830), .A2(n12829), .A3(n12828), .A4(n14844), .ZN(
        n12831) );
  NOR4_X1 U15203 ( .A1(n12841), .A2(n15069), .A3(n14718), .A4(n12840), .ZN(
        n12843) );
  OAI21_X1 U15204 ( .B1(n12844), .B2(n15244), .A(P1_B_REG_SCAN_IN), .ZN(n12842) );
  OAI22_X1 U15205 ( .A1(n12845), .A2(n12844), .B1(n12843), .B2(n12842), .ZN(
        P1_U3242) );
  AND2_X1 U15206 ( .A1(n13963), .A2(n13951), .ZN(n12848) );
  AOI21_X1 U15207 ( .B1(n13961), .B2(n13952), .A(n12848), .ZN(n14060) );
  INV_X1 U15208 ( .A(n12849), .ZN(n14065) );
  AOI22_X1 U15209 ( .A1(n13944), .A2(n14065), .B1(P2_REG3_REG_27__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12850) );
  OAI21_X1 U15210 ( .B1(n14060), .B2(n13953), .A(n12850), .ZN(n12851) );
  INV_X1 U15211 ( .A(n12851), .ZN(n12852) );
  INV_X1 U15212 ( .A(n12857), .ZN(P2_U3186) );
  INV_X1 U15213 ( .A(n12858), .ZN(n12859) );
  OAI222_X1 U15214 ( .A1(n12861), .A2(n12860), .B1(n14396), .B2(n12859), .C1(
        P2_U3088), .C2(n13099), .ZN(P2_U3305) );
  OAI21_X1 U15215 ( .B1(n12863), .B2(n12871), .A(n8325), .ZN(n12864) );
  NAND2_X1 U15216 ( .A1(n13989), .A2(n12864), .ZN(n12870) );
  NAND2_X1 U15217 ( .A1(n13159), .A2(n13099), .ZN(n12865) );
  NAND2_X1 U15218 ( .A1(n12865), .A2(n8325), .ZN(n12867) );
  NAND3_X1 U15219 ( .A1(n12867), .A2(n12866), .A3(n15616), .ZN(n12869) );
  NAND3_X1 U15220 ( .A1(n12870), .A2(n12869), .A3(n12868), .ZN(n12877) );
  NAND2_X1 U15221 ( .A1(n8886), .A2(n12871), .ZN(n12873) );
  NAND2_X1 U15222 ( .A1(n13988), .A2(n12888), .ZN(n12872) );
  AOI22_X1 U15223 ( .A1(n13988), .A2(n12871), .B1(n8886), .B2(n12888), .ZN(
        n12875) );
  AOI21_X1 U15224 ( .B1(n12877), .B2(n12876), .A(n12875), .ZN(n12879) );
  NOR2_X1 U15225 ( .A1(n12877), .A2(n12876), .ZN(n12878) );
  NAND2_X1 U15226 ( .A1(n13987), .A2(n12871), .ZN(n12881) );
  NAND2_X1 U15227 ( .A1(n12882), .A2(n12888), .ZN(n12880) );
  NAND2_X1 U15228 ( .A1(n12881), .A2(n12880), .ZN(n12884) );
  AOI22_X1 U15229 ( .A1(n13987), .A2(n12888), .B1(n12882), .B2(n12891), .ZN(
        n12883) );
  AOI21_X1 U15230 ( .B1(n12885), .B2(n12884), .A(n12883), .ZN(n12887) );
  NOR2_X1 U15231 ( .A1(n12885), .A2(n12884), .ZN(n12886) );
  NAND2_X1 U15232 ( .A1(n13986), .A2(n12984), .ZN(n12890) );
  NAND2_X1 U15233 ( .A1(n15652), .A2(n13097), .ZN(n12889) );
  NAND2_X1 U15234 ( .A1(n12890), .A2(n12889), .ZN(n12897) );
  NAND2_X1 U15235 ( .A1(n12896), .A2(n12897), .ZN(n12895) );
  NAND2_X1 U15236 ( .A1(n13986), .A2(n12891), .ZN(n12893) );
  NAND2_X1 U15237 ( .A1(n15652), .A2(n13088), .ZN(n12892) );
  NAND2_X1 U15238 ( .A1(n12893), .A2(n12892), .ZN(n12894) );
  NAND2_X1 U15239 ( .A1(n12895), .A2(n12894), .ZN(n12901) );
  INV_X1 U15240 ( .A(n12896), .ZN(n12899) );
  NAND2_X1 U15241 ( .A1(n12899), .A2(n12898), .ZN(n12900) );
  NAND2_X1 U15242 ( .A1(n15659), .A2(n13096), .ZN(n12903) );
  NAND2_X1 U15243 ( .A1(n13985), .A2(n13097), .ZN(n12902) );
  AOI22_X1 U15244 ( .A1(n15659), .A2(n12891), .B1(n13088), .B2(n13985), .ZN(
        n12904) );
  NAND2_X1 U15245 ( .A1(n12907), .A2(n12891), .ZN(n12906) );
  NAND2_X1 U15246 ( .A1(n13984), .A2(n13088), .ZN(n12905) );
  NAND2_X1 U15247 ( .A1(n12906), .A2(n12905), .ZN(n12913) );
  NAND2_X1 U15248 ( .A1(n12907), .A2(n13088), .ZN(n12908) );
  OAI21_X1 U15249 ( .B1(n12909), .B2(n13088), .A(n12908), .ZN(n12910) );
  NAND2_X1 U15250 ( .A1(n12911), .A2(n12910), .ZN(n12917) );
  INV_X1 U15251 ( .A(n12912), .ZN(n12915) );
  NAND2_X1 U15252 ( .A1(n12915), .A2(n12914), .ZN(n12916) );
  NAND2_X1 U15253 ( .A1(n15671), .A2(n13088), .ZN(n12919) );
  NAND2_X1 U15254 ( .A1(n13983), .A2(n13097), .ZN(n12918) );
  NAND2_X1 U15255 ( .A1(n12919), .A2(n12918), .ZN(n12921) );
  AOI22_X1 U15256 ( .A1(n15671), .A2(n13097), .B1(n13088), .B2(n13983), .ZN(
        n12920) );
  NAND2_X1 U15257 ( .A1(n12924), .A2(n13097), .ZN(n12923) );
  NAND2_X1 U15258 ( .A1(n13982), .A2(n13088), .ZN(n12922) );
  NAND2_X1 U15259 ( .A1(n12923), .A2(n12922), .ZN(n12930) );
  NAND2_X1 U15260 ( .A1(n12929), .A2(n12930), .ZN(n12928) );
  NAND2_X1 U15261 ( .A1(n12924), .A2(n12984), .ZN(n12925) );
  OAI21_X1 U15262 ( .B1(n12926), .B2(n13096), .A(n12925), .ZN(n12927) );
  INV_X1 U15263 ( .A(n12929), .ZN(n12932) );
  NAND2_X1 U15264 ( .A1(n12935), .A2(n13088), .ZN(n12934) );
  NAND2_X1 U15265 ( .A1(n13981), .A2(n13097), .ZN(n12933) );
  NAND2_X1 U15266 ( .A1(n12934), .A2(n12933), .ZN(n12937) );
  AOI22_X1 U15267 ( .A1(n12935), .A2(n12891), .B1(n12984), .B2(n13981), .ZN(
        n12936) );
  NAND2_X1 U15268 ( .A1(n12940), .A2(n13097), .ZN(n12939) );
  NAND2_X1 U15269 ( .A1(n13980), .A2(n13088), .ZN(n12938) );
  NAND2_X1 U15270 ( .A1(n12939), .A2(n12938), .ZN(n12942) );
  AOI22_X1 U15271 ( .A1(n12940), .A2(n13096), .B1(n13097), .B2(n13980), .ZN(
        n12941) );
  AOI21_X1 U15272 ( .B1(n12943), .B2(n12942), .A(n12941), .ZN(n12944) );
  NAND2_X1 U15273 ( .A1(n12947), .A2(n13088), .ZN(n12946) );
  NAND2_X1 U15274 ( .A1(n13979), .A2(n12891), .ZN(n12945) );
  NAND2_X1 U15275 ( .A1(n12947), .A2(n13097), .ZN(n12948) );
  OAI21_X1 U15276 ( .B1(n12891), .B2(n12949), .A(n12948), .ZN(n12950) );
  NAND2_X1 U15277 ( .A1(n15349), .A2(n12891), .ZN(n12952) );
  NAND2_X1 U15278 ( .A1(n13978), .A2(n13088), .ZN(n12951) );
  NAND2_X1 U15279 ( .A1(n12952), .A2(n12951), .ZN(n12954) );
  AOI22_X1 U15280 ( .A1(n15349), .A2(n13096), .B1(n13097), .B2(n13978), .ZN(
        n12953) );
  AOI21_X1 U15281 ( .B1(n12955), .B2(n12954), .A(n12953), .ZN(n12956) );
  NAND2_X1 U15282 ( .A1(n12959), .A2(n13096), .ZN(n12958) );
  NAND2_X1 U15283 ( .A1(n13977), .A2(n12891), .ZN(n12957) );
  NAND2_X1 U15284 ( .A1(n12958), .A2(n12957), .ZN(n12963) );
  NAND2_X1 U15285 ( .A1(n12959), .A2(n13097), .ZN(n12960) );
  OAI21_X1 U15286 ( .B1(n13097), .B2(n12961), .A(n12960), .ZN(n12962) );
  INV_X1 U15287 ( .A(n12963), .ZN(n12964) );
  NAND2_X1 U15288 ( .A1(n12967), .A2(n13097), .ZN(n12966) );
  NAND2_X1 U15289 ( .A1(n13976), .A2(n12984), .ZN(n12965) );
  NAND2_X1 U15290 ( .A1(n12966), .A2(n12965), .ZN(n12969) );
  AOI22_X1 U15291 ( .A1(n12967), .A2(n13096), .B1(n13097), .B2(n13976), .ZN(
        n12968) );
  AOI21_X1 U15292 ( .B1(n12970), .B2(n12969), .A(n12968), .ZN(n12992) );
  NOR2_X1 U15293 ( .A1(n12970), .A2(n12969), .ZN(n12991) );
  AOI22_X1 U15294 ( .A1(n14307), .A2(n13088), .B1(n13097), .B2(n13972), .ZN(
        n12973) );
  NAND2_X1 U15295 ( .A1(n14307), .A2(n13097), .ZN(n12972) );
  NAND2_X1 U15296 ( .A1(n13972), .A2(n13096), .ZN(n12971) );
  NAND2_X1 U15297 ( .A1(n12972), .A2(n12971), .ZN(n13004) );
  NAND2_X1 U15298 ( .A1(n12973), .A2(n13004), .ZN(n12978) );
  AND2_X1 U15299 ( .A1(n13973), .A2(n13097), .ZN(n12974) );
  AOI21_X1 U15300 ( .B1(n14376), .B2(n12984), .A(n12974), .ZN(n12997) );
  NAND2_X1 U15301 ( .A1(n14376), .A2(n12891), .ZN(n12976) );
  NAND2_X1 U15302 ( .A1(n13973), .A2(n12984), .ZN(n12975) );
  NAND2_X1 U15303 ( .A1(n12976), .A2(n12975), .ZN(n12996) );
  NAND2_X1 U15304 ( .A1(n12997), .A2(n12996), .ZN(n12977) );
  AND2_X1 U15305 ( .A1(n12978), .A2(n12977), .ZN(n13001) );
  AND2_X1 U15306 ( .A1(n13974), .A2(n13097), .ZN(n12979) );
  AOI21_X1 U15307 ( .B1(n12980), .B2(n12984), .A(n12979), .ZN(n12999) );
  NAND2_X1 U15308 ( .A1(n12980), .A2(n13097), .ZN(n12982) );
  NAND2_X1 U15309 ( .A1(n13974), .A2(n12984), .ZN(n12981) );
  NAND2_X1 U15310 ( .A1(n12982), .A2(n12981), .ZN(n12998) );
  NAND2_X1 U15311 ( .A1(n12999), .A2(n12998), .ZN(n12983) );
  AND2_X1 U15312 ( .A1(n13001), .A2(n12983), .ZN(n12993) );
  NAND2_X1 U15313 ( .A1(n12988), .A2(n13088), .ZN(n12986) );
  NAND2_X1 U15314 ( .A1(n13975), .A2(n12891), .ZN(n12985) );
  AND2_X1 U15315 ( .A1(n13975), .A2(n13088), .ZN(n12987) );
  AOI21_X1 U15316 ( .B1(n12988), .B2(n13097), .A(n12987), .ZN(n12994) );
  NOR2_X1 U15317 ( .A1(n14307), .A2(n13972), .ZN(n13005) );
  INV_X1 U15318 ( .A(n12993), .ZN(n12995) );
  OR3_X1 U15319 ( .A1(n12995), .A2(n7737), .A3(n12989), .ZN(n13003) );
  OAI22_X1 U15320 ( .A1(n12999), .A2(n12998), .B1(n12997), .B2(n12996), .ZN(
        n13000) );
  NAND2_X1 U15321 ( .A1(n13001), .A2(n13000), .ZN(n13002) );
  OAI211_X1 U15322 ( .C1(n13005), .C2(n13004), .A(n13003), .B(n13002), .ZN(
        n13006) );
  INV_X1 U15323 ( .A(n13006), .ZN(n13007) );
  NAND2_X1 U15324 ( .A1(n13008), .A2(n13007), .ZN(n13012) );
  NAND2_X1 U15325 ( .A1(n14210), .A2(n13088), .ZN(n13010) );
  NAND2_X1 U15326 ( .A1(n13971), .A2(n13097), .ZN(n13009) );
  AOI22_X1 U15327 ( .A1(n14210), .A2(n12891), .B1(n12984), .B2(n13971), .ZN(
        n13011) );
  NAND2_X1 U15328 ( .A1(n14295), .A2(n12891), .ZN(n13014) );
  NAND2_X1 U15329 ( .A1(n13970), .A2(n13096), .ZN(n13013) );
  NAND2_X1 U15330 ( .A1(n14295), .A2(n13088), .ZN(n13016) );
  NAND2_X1 U15331 ( .A1(n13970), .A2(n13097), .ZN(n13015) );
  NAND2_X1 U15332 ( .A1(n13016), .A2(n13015), .ZN(n13017) );
  NAND2_X1 U15333 ( .A1(n13018), .A2(n13017), .ZN(n13022) );
  INV_X1 U15334 ( .A(n13019), .ZN(n13020) );
  NAND2_X1 U15335 ( .A1(n13020), .A2(n6771), .ZN(n13021) );
  NAND2_X1 U15336 ( .A1(n14289), .A2(n12984), .ZN(n13024) );
  NAND2_X1 U15337 ( .A1(n13969), .A2(n13097), .ZN(n13023) );
  NAND2_X1 U15338 ( .A1(n13024), .A2(n13023), .ZN(n13026) );
  AOI22_X1 U15339 ( .A1(n14289), .A2(n13097), .B1(n13096), .B2(n13969), .ZN(
        n13025) );
  NAND2_X1 U15340 ( .A1(n14285), .A2(n13097), .ZN(n13028) );
  NAND2_X1 U15341 ( .A1(n13968), .A2(n12984), .ZN(n13027) );
  NAND2_X1 U15342 ( .A1(n13028), .A2(n13027), .ZN(n13033) );
  NAND2_X1 U15343 ( .A1(n14285), .A2(n13096), .ZN(n13029) );
  OAI21_X1 U15344 ( .B1(n13916), .B2(n12984), .A(n13029), .ZN(n13030) );
  NAND2_X1 U15345 ( .A1(n13031), .A2(n13030), .ZN(n13037) );
  INV_X1 U15346 ( .A(n13032), .ZN(n13035) );
  NAND2_X1 U15347 ( .A1(n13035), .A2(n13034), .ZN(n13036) );
  NAND2_X1 U15348 ( .A1(n13037), .A2(n13036), .ZN(n13043) );
  NAND2_X1 U15349 ( .A1(n14351), .A2(n13088), .ZN(n13039) );
  NAND2_X1 U15350 ( .A1(n13967), .A2(n12891), .ZN(n13038) );
  NAND2_X1 U15351 ( .A1(n13039), .A2(n13038), .ZN(n13042) );
  AOI22_X1 U15352 ( .A1(n14351), .A2(n13097), .B1(n12984), .B2(n13967), .ZN(
        n13040) );
  AOI21_X1 U15353 ( .B1(n13043), .B2(n13042), .A(n13040), .ZN(n13041) );
  NOR2_X1 U15354 ( .A1(n13043), .A2(n13042), .ZN(n13044) );
  AND2_X1 U15355 ( .A1(n13966), .A2(n13088), .ZN(n13045) );
  AOI21_X1 U15356 ( .B1(n14274), .B2(n13097), .A(n13045), .ZN(n13050) );
  INV_X1 U15357 ( .A(n13050), .ZN(n13046) );
  NAND2_X1 U15358 ( .A1(n14274), .A2(n13088), .ZN(n13047) );
  OAI21_X1 U15359 ( .B1(n13048), .B2(n13096), .A(n13047), .ZN(n13049) );
  NAND2_X1 U15360 ( .A1(n14343), .A2(n12984), .ZN(n13052) );
  NAND2_X1 U15361 ( .A1(n13965), .A2(n13097), .ZN(n13051) );
  NAND2_X1 U15362 ( .A1(n13052), .A2(n13051), .ZN(n13054) );
  AOI22_X1 U15363 ( .A1(n14343), .A2(n12891), .B1(n13096), .B2(n13965), .ZN(
        n13053) );
  AOI21_X1 U15364 ( .B1(n13055), .B2(n13054), .A(n13053), .ZN(n13057) );
  NOR2_X1 U15365 ( .A1(n13055), .A2(n13054), .ZN(n13056) );
  NAND2_X1 U15366 ( .A1(n14262), .A2(n12891), .ZN(n13059) );
  NAND2_X1 U15367 ( .A1(n13964), .A2(n13096), .ZN(n13058) );
  NAND2_X1 U15368 ( .A1(n13059), .A2(n13058), .ZN(n13061) );
  AOI22_X1 U15369 ( .A1(n14262), .A2(n13088), .B1(n13097), .B2(n13964), .ZN(
        n13060) );
  AOI21_X1 U15370 ( .B1(n13062), .B2(n13061), .A(n13060), .ZN(n13064) );
  NOR2_X1 U15371 ( .A1(n13062), .A2(n13061), .ZN(n13063) );
  NAND2_X1 U15372 ( .A1(n14256), .A2(n13088), .ZN(n13066) );
  NAND2_X1 U15373 ( .A1(n13963), .A2(n13097), .ZN(n13065) );
  NAND2_X1 U15374 ( .A1(n13066), .A2(n13065), .ZN(n13071) );
  AND2_X1 U15375 ( .A1(n13962), .A2(n12984), .ZN(n13067) );
  AOI21_X1 U15376 ( .B1(n14329), .B2(n13097), .A(n13067), .ZN(n13076) );
  NAND2_X1 U15377 ( .A1(n14329), .A2(n13096), .ZN(n13069) );
  NAND2_X1 U15378 ( .A1(n13962), .A2(n13097), .ZN(n13068) );
  NAND2_X1 U15379 ( .A1(n13069), .A2(n13068), .ZN(n13075) );
  AOI22_X1 U15380 ( .A1(n14256), .A2(n13097), .B1(n13088), .B2(n13963), .ZN(
        n13070) );
  AND2_X1 U15381 ( .A1(n13961), .A2(n13096), .ZN(n13072) );
  AOI21_X1 U15382 ( .B1(n14247), .B2(n13097), .A(n13072), .ZN(n13080) );
  NAND2_X1 U15383 ( .A1(n14247), .A2(n13088), .ZN(n13074) );
  NAND2_X1 U15384 ( .A1(n13961), .A2(n12891), .ZN(n13073) );
  NAND2_X1 U15385 ( .A1(n13074), .A2(n13073), .ZN(n13079) );
  NAND2_X1 U15386 ( .A1(n13080), .A2(n13079), .ZN(n13078) );
  NAND2_X1 U15387 ( .A1(n13076), .A2(n13075), .ZN(n13077) );
  INV_X1 U15388 ( .A(n13079), .ZN(n13082) );
  INV_X1 U15389 ( .A(n13080), .ZN(n13081) );
  NAND2_X1 U15390 ( .A1(n13082), .A2(n13081), .ZN(n13092) );
  NAND2_X1 U15391 ( .A1(n13083), .A2(n8412), .ZN(n13086) );
  OR2_X1 U15392 ( .A1(n8379), .A2(n13084), .ZN(n13085) );
  XNOR2_X1 U15393 ( .A(n14020), .B(n14023), .ZN(n13151) );
  AND2_X1 U15394 ( .A1(n13960), .A2(n12984), .ZN(n13087) );
  AOI21_X1 U15395 ( .B1(n14031), .B2(n13097), .A(n13087), .ZN(n13104) );
  NAND2_X1 U15396 ( .A1(n14031), .A2(n12984), .ZN(n13090) );
  NAND2_X1 U15397 ( .A1(n13960), .A2(n13097), .ZN(n13089) );
  NAND2_X1 U15398 ( .A1(n13090), .A2(n13089), .ZN(n13103) );
  AND2_X1 U15399 ( .A1(n13104), .A2(n13103), .ZN(n13091) );
  MUX2_X1 U15400 ( .A(n13098), .B(n13097), .S(n14020), .Z(n13108) );
  NAND2_X1 U15401 ( .A1(n13098), .A2(n13097), .ZN(n13114) );
  OR2_X1 U15402 ( .A1(n8379), .A2(n9487), .ZN(n13094) );
  AND2_X1 U15403 ( .A1(n13959), .A2(n13097), .ZN(n13095) );
  AOI21_X1 U15404 ( .B1(n14019), .B2(n12984), .A(n13095), .ZN(n13110) );
  NAND2_X1 U15405 ( .A1(n14019), .A2(n13097), .ZN(n13102) );
  NAND2_X1 U15406 ( .A1(n13098), .A2(n13096), .ZN(n13112) );
  OR2_X1 U15407 ( .A1(n15620), .A2(n13099), .ZN(n13161) );
  NAND4_X1 U15408 ( .A1(n8321), .A2(n13112), .A3(n13161), .A4(n13157), .ZN(
        n13100) );
  NAND2_X1 U15409 ( .A1(n13100), .A2(n13959), .ZN(n13101) );
  INV_X1 U15410 ( .A(n13103), .ZN(n13106) );
  INV_X1 U15411 ( .A(n13104), .ZN(n13105) );
  AOI22_X1 U15412 ( .A1(n13110), .A2(n13109), .B1(n13106), .B2(n13105), .ZN(
        n13107) );
  AOI21_X1 U15413 ( .B1(n13108), .B2(n13114), .A(n13107), .ZN(n13111) );
  NAND2_X1 U15414 ( .A1(n13112), .A2(n13096), .ZN(n13113) );
  MUX2_X1 U15415 ( .A(n13114), .B(n13113), .S(n14020), .Z(n13115) );
  XOR2_X1 U15416 ( .A(n13959), .B(n14019), .Z(n13150) );
  AND2_X1 U15417 ( .A1(n13120), .A2(n13119), .ZN(n15636) );
  NAND4_X1 U15418 ( .A1(n15636), .A2(n6961), .A3(n13122), .A4(n13121), .ZN(
        n13125) );
  NOR4_X1 U15419 ( .A1(n13127), .A2(n13126), .A3(n13125), .A4(n13124), .ZN(
        n13131) );
  NAND4_X1 U15420 ( .A1(n13131), .A2(n13130), .A3(n13129), .A4(n13128), .ZN(
        n13132) );
  NOR4_X1 U15421 ( .A1(n13135), .A2(n13134), .A3(n13133), .A4(n13132), .ZN(
        n13138) );
  NAND4_X1 U15422 ( .A1(n13139), .A2(n13138), .A3(n13137), .A4(n13136), .ZN(
        n13140) );
  NOR4_X1 U15423 ( .A1(n13142), .A2(n14223), .A3(n13141), .A4(n13140), .ZN(
        n13143) );
  XNOR2_X1 U15424 ( .A(n14295), .B(n13970), .ZN(n14186) );
  NAND4_X1 U15425 ( .A1(n14170), .A2(n13143), .A3(n14198), .A4(n14186), .ZN(
        n13144) );
  NOR4_X1 U15426 ( .A1(n14125), .A2(n14161), .A3(n13145), .A4(n13144), .ZN(
        n13147) );
  NAND4_X1 U15427 ( .A1(n14080), .A2(n13147), .A3(n13146), .A4(n14104), .ZN(
        n13148) );
  NOR4_X1 U15428 ( .A1(n13150), .A2(n13149), .A3(n14041), .A4(n13148), .ZN(
        n13154) );
  INV_X1 U15429 ( .A(n13151), .ZN(n13153) );
  NAND3_X1 U15430 ( .A1(n13154), .A2(n13153), .A3(n13152), .ZN(n13155) );
  OAI211_X1 U15431 ( .C1(n13159), .C2(n13158), .A(n13157), .B(n13156), .ZN(
        n13160) );
  INV_X1 U15432 ( .A(n13160), .ZN(n13164) );
  OAI21_X1 U15433 ( .B1(n13162), .B2(n8859), .A(n13161), .ZN(n13163) );
  NAND4_X1 U15434 ( .A1(n15635), .A2(n13951), .A3(n13167), .A4(n13166), .ZN(
        n13168) );
  OAI211_X1 U15435 ( .C1(n13169), .C2(n13171), .A(n13168), .B(P2_B_REG_SCAN_IN), .ZN(n13170) );
  INV_X1 U15436 ( .A(n13172), .ZN(n13173) );
  OAI222_X1 U15437 ( .A1(n13851), .A2(n13173), .B1(n13840), .B2(n8127), .C1(
        P3_U3151), .C2(n9689), .ZN(P3_U3267) );
  AOI22_X1 U15438 ( .A1(n15304), .A2(n15709), .B1(P3_REG2_REG_29__SCAN_IN), 
        .B2(n15735), .ZN(n13175) );
  OAI21_X1 U15439 ( .B1(n13176), .B2(n13714), .A(n13175), .ZN(n13177) );
  AOI21_X1 U15440 ( .B1(n13178), .B2(n13716), .A(n13177), .ZN(n13179) );
  OAI21_X1 U15441 ( .B1(n13174), .B2(n15735), .A(n13179), .ZN(P3_U3204) );
  INV_X1 U15442 ( .A(n13184), .ZN(n13181) );
  NAND2_X1 U15443 ( .A1(n13181), .A2(n13180), .ZN(n13182) );
  XNOR2_X1 U15444 ( .A(n13824), .B(n13254), .ZN(n13186) );
  XOR2_X1 U15445 ( .A(n13706), .B(n13186), .Z(n13225) );
  XNOR2_X1 U15446 ( .A(n13187), .B(n13254), .ZN(n13188) );
  XOR2_X1 U15447 ( .A(n13693), .B(n13188), .Z(n13341) );
  INV_X1 U15448 ( .A(n13188), .ZN(n13189) );
  NAND2_X1 U15449 ( .A1(n13189), .A2(n13227), .ZN(n13190) );
  XNOR2_X1 U15450 ( .A(n13699), .B(n13254), .ZN(n13277) );
  NAND2_X1 U15451 ( .A1(n13277), .A2(n13680), .ZN(n13192) );
  XNOR2_X1 U15452 ( .A(n13295), .B(n13254), .ZN(n13193) );
  XNOR2_X1 U15453 ( .A(n13193), .B(n13326), .ZN(n13287) );
  NAND2_X1 U15454 ( .A1(n13193), .A2(n13326), .ZN(n13194) );
  XNOR2_X1 U15455 ( .A(n13670), .B(n13254), .ZN(n13195) );
  XOR2_X1 U15456 ( .A(n13681), .B(n13195), .Z(n13324) );
  INV_X1 U15457 ( .A(n13195), .ZN(n13196) );
  XNOR2_X1 U15458 ( .A(n13813), .B(n13254), .ZN(n13197) );
  XNOR2_X1 U15459 ( .A(n13197), .B(n13664), .ZN(n13244) );
  NAND2_X1 U15460 ( .A1(n13197), .A2(n13308), .ZN(n13198) );
  XNOR2_X1 U15461 ( .A(n13809), .B(n13254), .ZN(n13199) );
  XNOR2_X1 U15462 ( .A(n13199), .B(n13629), .ZN(n13306) );
  NAND2_X1 U15463 ( .A1(n13199), .A2(n13652), .ZN(n13200) );
  XNOR2_X1 U15464 ( .A(n13267), .B(n13254), .ZN(n13202) );
  XNOR2_X1 U15465 ( .A(n13202), .B(n13638), .ZN(n13263) );
  INV_X1 U15466 ( .A(n13263), .ZN(n13201) );
  XNOR2_X1 U15467 ( .A(n13318), .B(n13207), .ZN(n13203) );
  INV_X1 U15468 ( .A(n13203), .ZN(n13204) );
  XNOR2_X1 U15469 ( .A(n13797), .B(n13207), .ZN(n13208) );
  INV_X1 U15470 ( .A(n13208), .ZN(n13209) );
  OR2_X1 U15471 ( .A1(n13210), .A2(n13209), .ZN(n13211) );
  XNOR2_X1 U15472 ( .A(n13793), .B(n13254), .ZN(n13212) );
  INV_X1 U15473 ( .A(n13212), .ZN(n13213) );
  NAND2_X1 U15474 ( .A1(n13213), .A2(n13580), .ZN(n13214) );
  XNOR2_X1 U15475 ( .A(n13581), .B(n13254), .ZN(n13215) );
  XNOR2_X1 U15476 ( .A(n13215), .B(n13333), .ZN(n13271) );
  NAND2_X1 U15477 ( .A1(n13215), .A2(n13590), .ZN(n13216) );
  XNOR2_X1 U15478 ( .A(n13338), .B(n13254), .ZN(n13217) );
  XNOR2_X1 U15479 ( .A(n13217), .B(n13577), .ZN(n13332) );
  XNOR2_X1 U15480 ( .A(n13782), .B(n13254), .ZN(n13250) );
  INV_X1 U15481 ( .A(n13252), .ZN(n13218) );
  XNOR2_X1 U15482 ( .A(n13253), .B(n13218), .ZN(n13223) );
  AOI22_X1 U15483 ( .A1(n13577), .A2(n13343), .B1(P3_REG3_REG_27__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13220) );
  NAND2_X1 U15484 ( .A1(n13557), .A2(n13350), .ZN(n13219) );
  OAI211_X1 U15485 ( .C1(n6675), .C2(n13346), .A(n13220), .B(n13219), .ZN(
        n13221) );
  AOI21_X1 U15486 ( .B1(n13556), .B2(n13337), .A(n13221), .ZN(n13222) );
  OAI21_X1 U15487 ( .B1(n13223), .B2(n13352), .A(n13222), .ZN(P3_U3154) );
  XNOR2_X1 U15488 ( .A(n13224), .B(n13225), .ZN(n13234) );
  NOR2_X1 U15489 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n13226), .ZN(n13402) );
  AOI21_X1 U15490 ( .B1(n13227), .B2(n13281), .A(n13402), .ZN(n13230) );
  NAND2_X1 U15491 ( .A1(n13350), .A2(n13228), .ZN(n13229) );
  OAI211_X1 U15492 ( .C1(n13180), .C2(n13315), .A(n13230), .B(n13229), .ZN(
        n13231) );
  AOI21_X1 U15493 ( .B1(n13232), .B2(n13337), .A(n13231), .ZN(n13233) );
  OAI21_X1 U15494 ( .B1(n13234), .B2(n13352), .A(n13233), .ZN(P3_U3155) );
  XNOR2_X1 U15495 ( .A(n13235), .B(n13298), .ZN(n13242) );
  OAI22_X1 U15496 ( .A1(n13630), .A2(n13315), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n13236), .ZN(n13238) );
  NOR2_X1 U15497 ( .A1(n13580), .A2(n13346), .ZN(n13237) );
  AOI211_X1 U15498 ( .C1(n13606), .C2(n13350), .A(n13238), .B(n13237), .ZN(
        n13241) );
  NAND2_X1 U15499 ( .A1(n13239), .A2(n13337), .ZN(n13240) );
  OAI211_X1 U15500 ( .C1(n13242), .C2(n13352), .A(n13241), .B(n13240), .ZN(
        P3_U3156) );
  OAI211_X1 U15501 ( .C1(n13245), .C2(n13244), .A(n13243), .B(n13322), .ZN(
        n13249) );
  NAND2_X1 U15502 ( .A1(n7656), .A2(n13343), .ZN(n13246) );
  NAND2_X1 U15503 ( .A1(P3_U3151), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n13526)
         );
  OAI211_X1 U15504 ( .C1(n13629), .C2(n13346), .A(n13246), .B(n13526), .ZN(
        n13247) );
  AOI21_X1 U15505 ( .B1(n13655), .B2(n13350), .A(n13247), .ZN(n13248) );
  OAI211_X1 U15506 ( .C1(n13347), .C2(n13813), .A(n13249), .B(n13248), .ZN(
        P3_U3159) );
  INV_X1 U15507 ( .A(n13250), .ZN(n13251) );
  XNOR2_X1 U15508 ( .A(n13537), .B(n13254), .ZN(n13255) );
  XNOR2_X1 U15509 ( .A(n13256), .B(n13255), .ZN(n13261) );
  NOR2_X1 U15510 ( .A1(n13533), .A2(n13346), .ZN(n13259) );
  AOI22_X1 U15511 ( .A1(n13539), .A2(n13350), .B1(P3_REG3_REG_28__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13257) );
  OAI21_X1 U15512 ( .B1(n13565), .B2(n13315), .A(n13257), .ZN(n13258) );
  AOI211_X1 U15513 ( .C1(n13540), .C2(n13337), .A(n13259), .B(n13258), .ZN(
        n13260) );
  OAI21_X1 U15514 ( .B1(n13261), .B2(n13352), .A(n13260), .ZN(P3_U3160) );
  AOI21_X1 U15515 ( .B1(n13263), .B2(n13262), .A(n6822), .ZN(n13269) );
  AOI22_X1 U15516 ( .A1(n13343), .A2(n13652), .B1(P3_REG3_REG_21__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13265) );
  NAND2_X1 U15517 ( .A1(n13350), .A2(n13631), .ZN(n13264) );
  OAI211_X1 U15518 ( .C1(n13630), .C2(n13346), .A(n13265), .B(n13264), .ZN(
        n13266) );
  AOI21_X1 U15519 ( .B1(n13267), .B2(n13337), .A(n13266), .ZN(n13268) );
  OAI21_X1 U15520 ( .B1(n13269), .B2(n13352), .A(n13268), .ZN(P3_U3163) );
  XOR2_X1 U15521 ( .A(n13271), .B(n13270), .Z(n13276) );
  AOI22_X1 U15522 ( .A1(n13603), .A2(n13343), .B1(P3_REG3_REG_25__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13273) );
  NAND2_X1 U15523 ( .A1(n13582), .A2(n13350), .ZN(n13272) );
  OAI211_X1 U15524 ( .C1(n13548), .C2(n13346), .A(n13273), .B(n13272), .ZN(
        n13274) );
  AOI21_X1 U15525 ( .B1(n13581), .B2(n13337), .A(n13274), .ZN(n13275) );
  OAI21_X1 U15526 ( .B1(n13276), .B2(n13352), .A(n13275), .ZN(P3_U3165) );
  XNOR2_X1 U15527 ( .A(n13277), .B(n13707), .ZN(n13278) );
  XNOR2_X1 U15528 ( .A(n13279), .B(n13278), .ZN(n13286) );
  NOR2_X1 U15529 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n13280), .ZN(n13446) );
  AOI21_X1 U15530 ( .B1(n13281), .B2(n13326), .A(n13446), .ZN(n13283) );
  NAND2_X1 U15531 ( .A1(n13350), .A2(n13700), .ZN(n13282) );
  OAI211_X1 U15532 ( .C1(n13693), .C2(n13315), .A(n13283), .B(n13282), .ZN(
        n13284) );
  AOI21_X1 U15533 ( .B1(n13699), .B2(n13337), .A(n13284), .ZN(n13285) );
  OAI21_X1 U15534 ( .B1(n13286), .B2(n13352), .A(n13285), .ZN(P3_U3166) );
  AOI21_X1 U15535 ( .B1(n13288), .B2(n13287), .A(n13352), .ZN(n13290) );
  NAND2_X1 U15536 ( .A1(n13290), .A2(n13289), .ZN(n13294) );
  NAND2_X1 U15537 ( .A1(n13707), .A2(n13343), .ZN(n13291) );
  NAND2_X1 U15538 ( .A1(P3_U3151), .A2(P3_REG3_REG_17__SCAN_IN), .ZN(n13473)
         );
  OAI211_X1 U15539 ( .C1(n13681), .C2(n13346), .A(n13291), .B(n13473), .ZN(
        n13292) );
  AOI21_X1 U15540 ( .B1(n13682), .B2(n13350), .A(n13292), .ZN(n13293) );
  OAI211_X1 U15541 ( .C1(n13295), .C2(n13347), .A(n13294), .B(n13293), .ZN(
        P3_U3168) );
  XOR2_X1 U15542 ( .A(n13297), .B(n13296), .Z(n13304) );
  AOI22_X1 U15543 ( .A1(n13298), .A2(n13343), .B1(P3_REG3_REG_24__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13300) );
  NAND2_X1 U15544 ( .A1(n13594), .A2(n13350), .ZN(n13299) );
  OAI211_X1 U15545 ( .C1(n13590), .C2(n13346), .A(n13300), .B(n13299), .ZN(
        n13301) );
  AOI21_X1 U15546 ( .B1(n13302), .B2(n13337), .A(n13301), .ZN(n13303) );
  OAI21_X1 U15547 ( .B1(n13304), .B2(n13352), .A(n13303), .ZN(P3_U3169) );
  OAI211_X1 U15548 ( .C1(n13307), .C2(n13306), .A(n13305), .B(n13322), .ZN(
        n13312) );
  AOI22_X1 U15549 ( .A1(n13343), .A2(n13308), .B1(P3_REG3_REG_20__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13309) );
  OAI21_X1 U15550 ( .B1(n13638), .B2(n13346), .A(n13309), .ZN(n13310) );
  AOI21_X1 U15551 ( .B1(n13643), .B2(n13350), .A(n13310), .ZN(n13311) );
  OAI211_X1 U15552 ( .C1(n13809), .C2(n13347), .A(n13312), .B(n13311), .ZN(
        P3_U3173) );
  XOR2_X1 U15553 ( .A(n13313), .B(n13630), .Z(n13321) );
  OAI22_X1 U15554 ( .A1(n13638), .A2(n13315), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n13314), .ZN(n13317) );
  NOR2_X1 U15555 ( .A1(n13613), .A2(n13346), .ZN(n13316) );
  AOI211_X1 U15556 ( .C1(n13617), .C2(n13350), .A(n13317), .B(n13316), .ZN(
        n13320) );
  NAND2_X1 U15557 ( .A1(n13318), .A2(n13337), .ZN(n13319) );
  OAI211_X1 U15558 ( .C1(n13321), .C2(n13352), .A(n13320), .B(n13319), .ZN(
        P3_U3175) );
  OAI211_X1 U15559 ( .C1(n13325), .C2(n13324), .A(n13323), .B(n13322), .ZN(
        n13330) );
  NAND2_X1 U15560 ( .A1(n13343), .A2(n13326), .ZN(n13327) );
  NAND2_X1 U15561 ( .A1(P3_U3151), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n13490)
         );
  OAI211_X1 U15562 ( .C1(n13664), .C2(n13346), .A(n13327), .B(n13490), .ZN(
        n13328) );
  AOI21_X1 U15563 ( .B1(n13666), .B2(n13350), .A(n13328), .ZN(n13329) );
  OAI211_X1 U15564 ( .C1(n13760), .C2(n13347), .A(n13330), .B(n13329), .ZN(
        P3_U3178) );
  XOR2_X1 U15565 ( .A(n13332), .B(n13331), .Z(n13340) );
  AOI22_X1 U15566 ( .A1(n13333), .A2(n13343), .B1(P3_REG3_REG_26__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13335) );
  NAND2_X1 U15567 ( .A1(n13568), .A2(n13350), .ZN(n13334) );
  OAI211_X1 U15568 ( .C1(n13565), .C2(n13346), .A(n13335), .B(n13334), .ZN(
        n13336) );
  AOI21_X1 U15569 ( .B1(n13338), .B2(n13337), .A(n13336), .ZN(n13339) );
  OAI21_X1 U15570 ( .B1(n13340), .B2(n13352), .A(n13339), .ZN(P3_U3180) );
  XNOR2_X1 U15571 ( .A(n13342), .B(n13341), .ZN(n13353) );
  NAND2_X1 U15572 ( .A1(n13343), .A2(n13706), .ZN(n13345) );
  OR2_X1 U15573 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n13344), .ZN(n13414) );
  OAI211_X1 U15574 ( .C1(n13680), .C2(n13346), .A(n13345), .B(n13414), .ZN(
        n13349) );
  NOR2_X1 U15575 ( .A1(n13772), .A2(n13347), .ZN(n13348) );
  AOI211_X1 U15576 ( .C1(n13712), .C2(n13350), .A(n13349), .B(n13348), .ZN(
        n13351) );
  OAI21_X1 U15577 ( .B1(n13353), .B2(n13352), .A(n13351), .ZN(P3_U3181) );
  MUX2_X1 U15578 ( .A(n13354), .B(P3_DATAO_REG_29__SCAN_IN), .S(n13358), .Z(
        P3_U3520) );
  MUX2_X1 U15579 ( .A(n13355), .B(P3_DATAO_REG_13__SCAN_IN), .S(n13358), .Z(
        P3_U3504) );
  MUX2_X1 U15580 ( .A(P3_DATAO_REG_12__SCAN_IN), .B(n13356), .S(P3_U3897), .Z(
        P3_U3503) );
  MUX2_X1 U15581 ( .A(n13357), .B(P3_DATAO_REG_8__SCAN_IN), .S(n13358), .Z(
        P3_U3499) );
  MUX2_X1 U15582 ( .A(n15718), .B(P3_DATAO_REG_2__SCAN_IN), .S(n13358), .Z(
        P3_U3493) );
  MUX2_X1 U15583 ( .A(P3_DATAO_REG_1__SCAN_IN), .B(n10585), .S(P3_U3897), .Z(
        P3_U3492) );
  INV_X1 U15584 ( .A(P3_REG2_REG_13__SCAN_IN), .ZN(n13361) );
  AOI21_X1 U15585 ( .B1(n13361), .B2(n13360), .A(n13384), .ZN(n13382) );
  INV_X1 U15586 ( .A(n13362), .ZN(n13363) );
  OAI21_X1 U15587 ( .B1(n13492), .B2(n13364), .A(n13363), .ZN(n13374) );
  INV_X1 U15588 ( .A(n13365), .ZN(n13367) );
  INV_X1 U15589 ( .A(n13377), .ZN(n13366) );
  NOR2_X1 U15590 ( .A1(n13367), .A2(n13366), .ZN(n13369) );
  MUX2_X1 U15591 ( .A(P3_REG2_REG_13__SCAN_IN), .B(P3_REG1_REG_13__SCAN_IN), 
        .S(n6945), .Z(n13395) );
  XNOR2_X1 U15592 ( .A(n13395), .B(n13394), .ZN(n13368) );
  INV_X1 U15593 ( .A(n13400), .ZN(n13372) );
  OAI21_X1 U15594 ( .B1(n13370), .B2(n13369), .A(n13368), .ZN(n13371) );
  AOI21_X1 U15595 ( .B1(n13372), .B2(n13371), .A(n15692), .ZN(n13373) );
  AOI211_X1 U15596 ( .C1(n15699), .C2(n13388), .A(n13374), .B(n13373), .ZN(
        n13381) );
  AOI21_X1 U15597 ( .B1(n9234), .B2(n13378), .A(n13389), .ZN(n13379) );
  OR2_X1 U15598 ( .A1(n13379), .A2(n15693), .ZN(n13380) );
  OAI211_X1 U15599 ( .C1(n13382), .C2(n15694), .A(n13381), .B(n13380), .ZN(
        P3_U3195) );
  NOR2_X1 U15600 ( .A1(n13388), .A2(n13383), .ZN(n13385) );
  NAND2_X1 U15601 ( .A1(n13405), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n13417) );
  OAI21_X1 U15602 ( .B1(P3_REG2_REG_14__SCAN_IN), .B2(n13405), .A(n13417), 
        .ZN(n13397) );
  AOI21_X1 U15603 ( .B1(n13386), .B2(n13397), .A(n13410), .ZN(n13409) );
  AND2_X1 U15604 ( .A1(n13405), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n13425) );
  INV_X1 U15605 ( .A(n13425), .ZN(n13416) );
  NAND2_X1 U15606 ( .A1(n13390), .A2(n13775), .ZN(n13391) );
  NAND2_X1 U15607 ( .A1(n13416), .A2(n13391), .ZN(n13396) );
  AOI21_X1 U15608 ( .B1(n13392), .B2(n13396), .A(n13426), .ZN(n13393) );
  NOR2_X1 U15609 ( .A1(n13393), .A2(n15693), .ZN(n13407) );
  NOR2_X1 U15610 ( .A1(n13395), .A2(n13394), .ZN(n13399) );
  MUX2_X1 U15611 ( .A(n13397), .B(n13396), .S(n6945), .Z(n13398) );
  OAI21_X1 U15612 ( .B1(n13400), .B2(n13399), .A(n13398), .ZN(n13401) );
  NAND3_X1 U15613 ( .A1(n13401), .A2(n13529), .A3(n13419), .ZN(n13404) );
  AOI21_X1 U15614 ( .B1(n15698), .B2(P3_ADDR_REG_14__SCAN_IN), .A(n13402), 
        .ZN(n13403) );
  OAI211_X1 U15615 ( .C1(n13521), .C2(n13405), .A(n13404), .B(n13403), .ZN(
        n13406) );
  NOR2_X1 U15616 ( .A1(n13407), .A2(n13406), .ZN(n13408) );
  OAI21_X1 U15617 ( .B1(n13409), .B2(n15694), .A(n13408), .ZN(P3_U3196) );
  INV_X1 U15618 ( .A(P3_REG2_REG_15__SCAN_IN), .ZN(n13413) );
  INV_X1 U15619 ( .A(n13417), .ZN(n13411) );
  AOI21_X1 U15620 ( .B1(n13413), .B2(n13412), .A(n13450), .ZN(n13433) );
  OAI21_X1 U15621 ( .B1(n13492), .B2(n13415), .A(n13414), .ZN(n13424) );
  MUX2_X1 U15622 ( .A(n13417), .B(n13416), .S(n6945), .Z(n13418) );
  XNOR2_X1 U15623 ( .A(n13438), .B(n13427), .ZN(n13421) );
  MUX2_X1 U15624 ( .A(P3_REG2_REG_15__SCAN_IN), .B(P3_REG1_REG_15__SCAN_IN), 
        .S(n6945), .Z(n13420) );
  AOI21_X1 U15625 ( .B1(n13421), .B2(n13420), .A(n13439), .ZN(n13422) );
  NOR2_X1 U15626 ( .A1(n13422), .A2(n15692), .ZN(n13423) );
  AOI211_X1 U15627 ( .C1(n15699), .C2(n13449), .A(n13424), .B(n13423), .ZN(
        n13432) );
  AOI21_X1 U15628 ( .B1(n13429), .B2(n13428), .A(n13435), .ZN(n13430) );
  OR2_X1 U15629 ( .A1(n13430), .A2(n15693), .ZN(n13431) );
  OAI211_X1 U15630 ( .C1(n13433), .C2(n15694), .A(n13432), .B(n13431), .ZN(
        P3_U3197) );
  NAND2_X1 U15631 ( .A1(P3_REG1_REG_16__SCAN_IN), .A2(n13452), .ZN(n13465) );
  OAI21_X1 U15632 ( .B1(n13452), .B2(P3_REG1_REG_16__SCAN_IN), .A(n13465), 
        .ZN(n13437) );
  AOI21_X1 U15633 ( .B1(n6751), .B2(n13437), .A(n13467), .ZN(n13460) );
  INV_X1 U15634 ( .A(n13438), .ZN(n13440) );
  INV_X1 U15635 ( .A(P3_REG2_REG_16__SCAN_IN), .ZN(n13441) );
  MUX2_X1 U15636 ( .A(n13441), .B(n13767), .S(n6945), .Z(n13443) );
  INV_X1 U15637 ( .A(n13452), .ZN(n13442) );
  NOR2_X1 U15638 ( .A1(n13443), .A2(n13442), .ZN(n13477) );
  INV_X1 U15639 ( .A(n13477), .ZN(n13444) );
  NAND2_X1 U15640 ( .A1(n13443), .A2(n13442), .ZN(n13476) );
  NAND2_X1 U15641 ( .A1(n13444), .A2(n13476), .ZN(n13445) );
  XNOR2_X1 U15642 ( .A(n13478), .B(n13445), .ZN(n13458) );
  AOI21_X1 U15643 ( .B1(n15698), .B2(P3_ADDR_REG_16__SCAN_IN), .A(n13446), 
        .ZN(n13447) );
  OAI21_X1 U15644 ( .B1(n13521), .B2(n13452), .A(n13447), .ZN(n13457) );
  NOR2_X1 U15645 ( .A1(n13449), .A2(n13448), .ZN(n13451) );
  NAND2_X1 U15646 ( .A1(P3_REG2_REG_16__SCAN_IN), .A2(n13452), .ZN(n13461) );
  OAI21_X1 U15647 ( .B1(P3_REG2_REG_16__SCAN_IN), .B2(n13452), .A(n13461), 
        .ZN(n13453) );
  NOR2_X1 U15648 ( .A1(n13454), .A2(n13453), .ZN(n13463) );
  AOI21_X1 U15649 ( .B1(n13454), .B2(n13453), .A(n13463), .ZN(n13455) );
  NOR2_X1 U15650 ( .A1(n13455), .A2(n15694), .ZN(n13456) );
  AOI211_X1 U15651 ( .C1(n13529), .C2(n13458), .A(n13457), .B(n13456), .ZN(
        n13459) );
  OAI21_X1 U15652 ( .B1(n13460), .B2(n15693), .A(n13459), .ZN(P3_U3198) );
  INV_X1 U15653 ( .A(P3_REG2_REG_17__SCAN_IN), .ZN(n13684) );
  INV_X1 U15654 ( .A(n13461), .ZN(n13462) );
  AOI21_X1 U15655 ( .B1(n13684), .B2(n13464), .A(n13486), .ZN(n13484) );
  INV_X1 U15656 ( .A(n13465), .ZN(n13466) );
  XNOR2_X1 U15657 ( .A(n13500), .B(n13501), .ZN(n13469) );
  INV_X1 U15658 ( .A(n13469), .ZN(n13470) );
  NOR2_X1 U15659 ( .A1(n13470), .A2(P3_REG1_REG_17__SCAN_IN), .ZN(n13472) );
  OAI21_X1 U15660 ( .B1(n13502), .B2(n13472), .A(n13471), .ZN(n13474) );
  OAI211_X1 U15661 ( .C1(n13475), .C2(n13492), .A(n13474), .B(n13473), .ZN(
        n13482) );
  MUX2_X1 U15662 ( .A(P3_REG2_REG_17__SCAN_IN), .B(P3_REG1_REG_17__SCAN_IN), 
        .S(n6945), .Z(n13495) );
  XNOR2_X1 U15663 ( .A(n13495), .B(n13494), .ZN(n13480) );
  NOR2_X1 U15664 ( .A1(n13479), .A2(n13480), .ZN(n13493) );
  AOI211_X1 U15665 ( .C1(n13480), .C2(n13479), .A(n15692), .B(n13493), .ZN(
        n13481) );
  AOI211_X1 U15666 ( .C1(n15699), .C2(n13501), .A(n13482), .B(n13481), .ZN(
        n13483) );
  OAI21_X1 U15667 ( .B1(n13484), .B2(n15694), .A(n13483), .ZN(P3_U3199) );
  NOR2_X1 U15668 ( .A1(n13501), .A2(n13485), .ZN(n13487) );
  NAND2_X1 U15669 ( .A1(P3_REG2_REG_18__SCAN_IN), .A2(n13513), .ZN(n13488) );
  OAI21_X1 U15670 ( .B1(P3_REG2_REG_18__SCAN_IN), .B2(n13513), .A(n13488), 
        .ZN(n13489) );
  AOI21_X1 U15671 ( .B1(n6750), .B2(n13489), .A(n13512), .ZN(n13511) );
  INV_X1 U15672 ( .A(n13513), .ZN(n13515) );
  OAI21_X1 U15673 ( .B1(n13492), .B2(n13491), .A(n13490), .ZN(n13499) );
  MUX2_X1 U15674 ( .A(P3_REG2_REG_18__SCAN_IN), .B(P3_REG1_REG_18__SCAN_IN), 
        .S(n6945), .Z(n13497) );
  XOR2_X1 U15675 ( .A(n13513), .B(n13516), .Z(n13496) );
  NOR2_X1 U15676 ( .A1(n13496), .A2(n13497), .ZN(n13514) );
  AOI211_X1 U15677 ( .C1(n15699), .C2(n13515), .A(n13499), .B(n13498), .ZN(
        n13510) );
  NOR2_X1 U15678 ( .A1(n13501), .A2(n13500), .ZN(n13503) );
  NOR2_X1 U15679 ( .A1(n13515), .A2(n13504), .ZN(n13523) );
  INV_X1 U15680 ( .A(n13523), .ZN(n13505) );
  OAI21_X1 U15681 ( .B1(P3_REG1_REG_18__SCAN_IN), .B2(n13513), .A(n13505), 
        .ZN(n13506) );
  AOI21_X1 U15682 ( .B1(n13507), .B2(n13506), .A(n13522), .ZN(n13508) );
  OR2_X1 U15683 ( .A1(n13508), .A2(n15693), .ZN(n13509) );
  OAI211_X1 U15684 ( .C1(n13511), .C2(n15694), .A(n13510), .B(n13509), .ZN(
        P3_U3200) );
  XNOR2_X1 U15685 ( .A(n9671), .B(P3_REG2_REG_19__SCAN_IN), .ZN(n13518) );
  AOI21_X1 U15686 ( .B1(n13516), .B2(n13515), .A(n13514), .ZN(n13520) );
  XNOR2_X1 U15687 ( .A(n9671), .B(P3_REG1_REG_19__SCAN_IN), .ZN(n13524) );
  MUX2_X1 U15688 ( .A(n13524), .B(n13518), .S(n13517), .Z(n13519) );
  XNOR2_X1 U15689 ( .A(n13520), .B(n13519), .ZN(n13530) );
  NOR2_X1 U15690 ( .A1(n13521), .A2(n9671), .ZN(n13528) );
  INV_X1 U15691 ( .A(n13524), .ZN(n13525) );
  AOI21_X1 U15692 ( .B1(n13532), .B2(n13537), .A(n13691), .ZN(n13536) );
  OAI22_X1 U15693 ( .A1(n13533), .A2(n13696), .B1(n13565), .B2(n13694), .ZN(
        n13534) );
  AOI21_X1 U15694 ( .B1(n13536), .B2(n13535), .A(n13534), .ZN(n13718) );
  XNOR2_X1 U15695 ( .A(n13538), .B(n13537), .ZN(n13719) );
  AOI22_X1 U15696 ( .A1(n13539), .A2(n15709), .B1(n15735), .B2(
        P3_REG2_REG_28__SCAN_IN), .ZN(n13542) );
  NAND2_X1 U15697 ( .A1(n13540), .A2(n15707), .ZN(n13541) );
  OAI211_X1 U15698 ( .C1(n13719), .C2(n13688), .A(n13542), .B(n13541), .ZN(
        n13543) );
  INV_X1 U15699 ( .A(n13543), .ZN(n13544) );
  OAI21_X1 U15700 ( .B1(n13718), .B2(n15735), .A(n13544), .ZN(P3_U3205) );
  OAI21_X1 U15701 ( .B1(n13547), .B2(n13546), .A(n13545), .ZN(n13551) );
  OAI22_X1 U15702 ( .A1(n6675), .A2(n13696), .B1(n13548), .B2(n13694), .ZN(
        n13550) );
  AOI21_X1 U15703 ( .B1(n13551), .B2(n15722), .A(n13550), .ZN(n13555) );
  NAND2_X1 U15704 ( .A1(n13556), .A2(n15707), .ZN(n13559) );
  AOI22_X1 U15705 ( .A1(n13557), .A2(n15709), .B1(n15735), .B2(
        P3_REG2_REG_27__SCAN_IN), .ZN(n13558) );
  NAND2_X1 U15706 ( .A1(n13559), .A2(n13558), .ZN(n13560) );
  AOI21_X1 U15707 ( .B1(n13721), .B2(n13561), .A(n13560), .ZN(n13562) );
  OAI21_X1 U15708 ( .B1(n13722), .B2(n15735), .A(n13562), .ZN(P3_U3206) );
  XNOR2_X1 U15709 ( .A(n13563), .B(n13567), .ZN(n13564) );
  OAI222_X1 U15710 ( .A1(n13694), .A2(n13590), .B1(n13696), .B2(n13565), .C1(
        n13564), .C2(n13691), .ZN(n13724) );
  INV_X1 U15711 ( .A(n13724), .ZN(n13572) );
  XOR2_X1 U15712 ( .A(n13566), .B(n13567), .Z(n13725) );
  AOI22_X1 U15713 ( .A1(n13568), .A2(n15709), .B1(n15735), .B2(
        P3_REG2_REG_26__SCAN_IN), .ZN(n13569) );
  OAI21_X1 U15714 ( .B1(n9723), .B2(n13714), .A(n13569), .ZN(n13570) );
  AOI21_X1 U15715 ( .B1(n13725), .B2(n13716), .A(n13570), .ZN(n13571) );
  OAI21_X1 U15716 ( .B1(n13572), .B2(n15735), .A(n13571), .ZN(P3_U3207) );
  XNOR2_X1 U15717 ( .A(n13573), .B(n13574), .ZN(n13729) );
  INV_X1 U15718 ( .A(n13729), .ZN(n13586) );
  OAI211_X1 U15719 ( .C1(n13576), .C2(n9722), .A(n15722), .B(n13575), .ZN(
        n13579) );
  NAND2_X1 U15720 ( .A1(n13577), .A2(n15719), .ZN(n13578) );
  OAI211_X1 U15721 ( .C1(n13580), .C2(n13694), .A(n13579), .B(n13578), .ZN(
        n13728) );
  INV_X1 U15722 ( .A(n13581), .ZN(n13789) );
  AOI22_X1 U15723 ( .A1(n13582), .A2(n15709), .B1(n15735), .B2(
        P3_REG2_REG_25__SCAN_IN), .ZN(n13583) );
  OAI21_X1 U15724 ( .B1(n13789), .B2(n13714), .A(n13583), .ZN(n13584) );
  AOI21_X1 U15725 ( .B1(n13728), .B2(n15733), .A(n13584), .ZN(n13585) );
  OAI21_X1 U15726 ( .B1(n13688), .B2(n13586), .A(n13585), .ZN(P3_U3208) );
  AOI21_X1 U15727 ( .B1(n13592), .B2(n13588), .A(n13587), .ZN(n13589) );
  OAI222_X1 U15728 ( .A1(n13694), .A2(n13613), .B1(n13696), .B2(n13590), .C1(
        n13691), .C2(n13589), .ZN(n13732) );
  INV_X1 U15729 ( .A(n13732), .ZN(n13598) );
  OAI21_X1 U15730 ( .B1(n13593), .B2(n13592), .A(n13591), .ZN(n13733) );
  AOI22_X1 U15731 ( .A1(n13594), .A2(n15709), .B1(n15735), .B2(
        P3_REG2_REG_24__SCAN_IN), .ZN(n13595) );
  OAI21_X1 U15732 ( .B1(n13793), .B2(n13714), .A(n13595), .ZN(n13596) );
  AOI21_X1 U15733 ( .B1(n13733), .B2(n13716), .A(n13596), .ZN(n13597) );
  OAI21_X1 U15734 ( .B1(n13598), .B2(n15735), .A(n13597), .ZN(P3_U3209) );
  XNOR2_X1 U15735 ( .A(n13600), .B(n13602), .ZN(n13737) );
  INV_X1 U15736 ( .A(n13737), .ZN(n13610) );
  OAI211_X1 U15737 ( .C1(n7747), .C2(n13602), .A(n15722), .B(n13601), .ZN(
        n13605) );
  NAND2_X1 U15738 ( .A1(n13603), .A2(n15719), .ZN(n13604) );
  OAI211_X1 U15739 ( .C1(n13630), .C2(n13694), .A(n13605), .B(n13604), .ZN(
        n13736) );
  AOI22_X1 U15740 ( .A1(n15735), .A2(P3_REG2_REG_23__SCAN_IN), .B1(n15709), 
        .B2(n13606), .ZN(n13607) );
  OAI21_X1 U15741 ( .B1(n13797), .B2(n13714), .A(n13607), .ZN(n13608) );
  AOI21_X1 U15742 ( .B1(n13736), .B2(n15733), .A(n13608), .ZN(n13609) );
  OAI21_X1 U15743 ( .B1(n13610), .B2(n13688), .A(n13609), .ZN(P3_U3210) );
  XNOR2_X1 U15744 ( .A(n13611), .B(n7624), .ZN(n13612) );
  OAI222_X1 U15745 ( .A1(n13696), .A2(n13613), .B1(n13694), .B2(n13638), .C1(
        n13691), .C2(n13612), .ZN(n13740) );
  INV_X1 U15746 ( .A(n13740), .ZN(n13621) );
  XNOR2_X1 U15747 ( .A(n13616), .B(n13615), .ZN(n13741) );
  AOI22_X1 U15748 ( .A1(n15735), .A2(P3_REG2_REG_22__SCAN_IN), .B1(n15709), 
        .B2(n13617), .ZN(n13618) );
  OAI21_X1 U15749 ( .B1(n13801), .B2(n13714), .A(n13618), .ZN(n13619) );
  AOI21_X1 U15750 ( .B1(n13741), .B2(n13716), .A(n13619), .ZN(n13620) );
  OAI21_X1 U15751 ( .B1(n13621), .B2(n15735), .A(n13620), .ZN(P3_U3211) );
  XOR2_X1 U15752 ( .A(n13623), .B(n13627), .Z(n13745) );
  INV_X1 U15753 ( .A(n13745), .ZN(n13635) );
  INV_X1 U15754 ( .A(n13624), .ZN(n13625) );
  AOI21_X1 U15755 ( .B1(n13627), .B2(n13626), .A(n13625), .ZN(n13628) );
  OAI222_X1 U15756 ( .A1(n13696), .A2(n13630), .B1(n13694), .B2(n13629), .C1(
        n13691), .C2(n13628), .ZN(n13744) );
  AOI22_X1 U15757 ( .A1(n15735), .A2(P3_REG2_REG_21__SCAN_IN), .B1(n15709), 
        .B2(n13631), .ZN(n13632) );
  OAI21_X1 U15758 ( .B1(n13805), .B2(n13714), .A(n13632), .ZN(n13633) );
  AOI21_X1 U15759 ( .B1(n13744), .B2(n15733), .A(n13633), .ZN(n13634) );
  OAI21_X1 U15760 ( .B1(n13635), .B2(n13688), .A(n13634), .ZN(P3_U3212) );
  XNOR2_X1 U15761 ( .A(n13636), .B(n13641), .ZN(n13637) );
  OAI222_X1 U15762 ( .A1(n13696), .A2(n13638), .B1(n13694), .B2(n13664), .C1(
        n13637), .C2(n13691), .ZN(n13748) );
  INV_X1 U15763 ( .A(n13748), .ZN(n13647) );
  INV_X1 U15764 ( .A(n13639), .ZN(n13640) );
  AOI21_X1 U15765 ( .B1(n13642), .B2(n13641), .A(n13640), .ZN(n13749) );
  AOI22_X1 U15766 ( .A1(n15735), .A2(P3_REG2_REG_20__SCAN_IN), .B1(n15709), 
        .B2(n13643), .ZN(n13644) );
  OAI21_X1 U15767 ( .B1(n13809), .B2(n13714), .A(n13644), .ZN(n13645) );
  AOI21_X1 U15768 ( .B1(n13749), .B2(n13716), .A(n13645), .ZN(n13646) );
  OAI21_X1 U15769 ( .B1(n13647), .B2(n15735), .A(n13646), .ZN(P3_U3213) );
  XNOR2_X1 U15770 ( .A(n13648), .B(n13650), .ZN(n13753) );
  INV_X1 U15771 ( .A(n13753), .ZN(n13659) );
  OAI211_X1 U15772 ( .C1(n13651), .C2(n13650), .A(n13649), .B(n15722), .ZN(
        n13654) );
  NAND2_X1 U15773 ( .A1(n13652), .A2(n15719), .ZN(n13653) );
  OAI211_X1 U15774 ( .C1(n13681), .C2(n13694), .A(n13654), .B(n13653), .ZN(
        n13752) );
  AOI22_X1 U15775 ( .A1(n15735), .A2(P3_REG2_REG_19__SCAN_IN), .B1(n15709), 
        .B2(n13655), .ZN(n13656) );
  OAI21_X1 U15776 ( .B1(n13813), .B2(n13714), .A(n13656), .ZN(n13657) );
  AOI21_X1 U15777 ( .B1(n13752), .B2(n15733), .A(n13657), .ZN(n13658) );
  OAI21_X1 U15778 ( .B1(n13659), .B2(n13688), .A(n13658), .ZN(P3_U3214) );
  AOI21_X1 U15779 ( .B1(n13662), .B2(n13661), .A(n13660), .ZN(n13663) );
  OAI222_X1 U15780 ( .A1(n13696), .A2(n13664), .B1(n13694), .B2(n13695), .C1(
        n13691), .C2(n13663), .ZN(n13665) );
  INV_X1 U15781 ( .A(n13665), .ZN(n13759) );
  INV_X1 U15782 ( .A(P3_REG2_REG_18__SCAN_IN), .ZN(n13668) );
  INV_X1 U15783 ( .A(n13666), .ZN(n13667) );
  OAI22_X1 U15784 ( .A1(n15733), .A2(n13668), .B1(n13667), .B2(n15727), .ZN(
        n13669) );
  AOI21_X1 U15785 ( .B1(n13670), .B2(n15707), .A(n13669), .ZN(n13674) );
  NAND2_X1 U15786 ( .A1(n13672), .A2(n7651), .ZN(n13756) );
  NAND3_X1 U15787 ( .A1(n13757), .A2(n13756), .A3(n13716), .ZN(n13673) );
  OAI211_X1 U15788 ( .C1(n13759), .C2(n15735), .A(n13674), .B(n13673), .ZN(
        P3_U3215) );
  XOR2_X1 U15789 ( .A(n13676), .B(n13677), .Z(n13764) );
  XNOR2_X1 U15790 ( .A(n13678), .B(n13677), .ZN(n13679) );
  OAI222_X1 U15791 ( .A1(n13696), .A2(n13681), .B1(n13694), .B2(n13680), .C1(
        n13679), .C2(n13691), .ZN(n13761) );
  NAND2_X1 U15792 ( .A1(n13761), .A2(n15733), .ZN(n13687) );
  INV_X1 U15793 ( .A(n13682), .ZN(n13683) );
  OAI22_X1 U15794 ( .A1(n15733), .A2(n13684), .B1(n13683), .B2(n15727), .ZN(
        n13685) );
  AOI21_X1 U15795 ( .B1(n13762), .B2(n15707), .A(n13685), .ZN(n13686) );
  OAI211_X1 U15796 ( .C1(n13764), .C2(n13688), .A(n13687), .B(n13686), .ZN(
        P3_U3216) );
  XNOR2_X1 U15797 ( .A(n13690), .B(n13689), .ZN(n13692) );
  OAI222_X1 U15798 ( .A1(n13696), .A2(n13695), .B1(n13694), .B2(n13693), .C1(
        n13692), .C2(n13691), .ZN(n13765) );
  INV_X1 U15799 ( .A(n13765), .ZN(n13704) );
  XNOR2_X1 U15800 ( .A(n13698), .B(n7639), .ZN(n13766) );
  INV_X1 U15801 ( .A(n13699), .ZN(n13819) );
  AOI22_X1 U15802 ( .A1(n15735), .A2(P3_REG2_REG_16__SCAN_IN), .B1(n15709), 
        .B2(n13700), .ZN(n13701) );
  OAI21_X1 U15803 ( .B1(n13819), .B2(n13714), .A(n13701), .ZN(n13702) );
  AOI21_X1 U15804 ( .B1(n13766), .B2(n13716), .A(n13702), .ZN(n13703) );
  OAI21_X1 U15805 ( .B1(n13704), .B2(n15735), .A(n13703), .ZN(P3_U3217) );
  XOR2_X1 U15806 ( .A(n13705), .B(n13710), .Z(n13708) );
  AOI222_X1 U15807 ( .A1(n15722), .A2(n13708), .B1(n13707), .B2(n15719), .C1(
        n13706), .C2(n15717), .ZN(n13771) );
  XNOR2_X1 U15808 ( .A(n13711), .B(n13710), .ZN(n13769) );
  AOI22_X1 U15809 ( .A1(n15735), .A2(P3_REG2_REG_15__SCAN_IN), .B1(n15709), 
        .B2(n13712), .ZN(n13713) );
  OAI21_X1 U15810 ( .B1(n13772), .B2(n13714), .A(n13713), .ZN(n13715) );
  AOI21_X1 U15811 ( .B1(n13769), .B2(n13716), .A(n13715), .ZN(n13717) );
  OAI21_X1 U15812 ( .B1(n13771), .B2(n15735), .A(n13717), .ZN(P3_U3218) );
  OAI21_X1 U15813 ( .B1(n15327), .B2(n13719), .A(n13718), .ZN(n13778) );
  OAI21_X1 U15814 ( .B1(n13780), .B2(n13777), .A(n13720), .ZN(P3_U3487) );
  INV_X1 U15815 ( .A(n13721), .ZN(n13723) );
  AOI21_X1 U15816 ( .B1(n13725), .B2(n15316), .A(n13724), .ZN(n13783) );
  MUX2_X1 U15817 ( .A(n13726), .B(n13783), .S(n15784), .Z(n13727) );
  OAI21_X1 U15818 ( .B1(n9723), .B2(n13777), .A(n13727), .ZN(P3_U3485) );
  AOI21_X1 U15819 ( .B1(n13729), .B2(n15316), .A(n13728), .ZN(n13786) );
  MUX2_X1 U15820 ( .A(n13730), .B(n13786), .S(n15784), .Z(n13731) );
  OAI21_X1 U15821 ( .B1(n13789), .B2(n13777), .A(n13731), .ZN(P3_U3484) );
  AOI21_X1 U15822 ( .B1(n15316), .B2(n13733), .A(n13732), .ZN(n13790) );
  MUX2_X1 U15823 ( .A(n13734), .B(n13790), .S(n15784), .Z(n13735) );
  OAI21_X1 U15824 ( .B1(n13793), .B2(n13777), .A(n13735), .ZN(P3_U3483) );
  INV_X1 U15825 ( .A(P3_REG1_REG_23__SCAN_IN), .ZN(n13738) );
  AOI21_X1 U15826 ( .B1(n15316), .B2(n13737), .A(n13736), .ZN(n13794) );
  MUX2_X1 U15827 ( .A(n13738), .B(n13794), .S(n15784), .Z(n13739) );
  OAI21_X1 U15828 ( .B1(n13797), .B2(n13777), .A(n13739), .ZN(P3_U3482) );
  INV_X1 U15829 ( .A(P3_REG1_REG_22__SCAN_IN), .ZN(n13742) );
  AOI21_X1 U15830 ( .B1(n15316), .B2(n13741), .A(n13740), .ZN(n13798) );
  MUX2_X1 U15831 ( .A(n13742), .B(n13798), .S(n15784), .Z(n13743) );
  OAI21_X1 U15832 ( .B1(n13801), .B2(n13777), .A(n13743), .ZN(P3_U3481) );
  AOI21_X1 U15833 ( .B1(n15316), .B2(n13745), .A(n13744), .ZN(n13802) );
  MUX2_X1 U15834 ( .A(n13746), .B(n13802), .S(n15784), .Z(n13747) );
  OAI21_X1 U15835 ( .B1(n13805), .B2(n13777), .A(n13747), .ZN(P3_U3480) );
  AOI21_X1 U15836 ( .B1(n13749), .B2(n15316), .A(n13748), .ZN(n13806) );
  MUX2_X1 U15837 ( .A(n13750), .B(n13806), .S(n15784), .Z(n13751) );
  OAI21_X1 U15838 ( .B1(n13809), .B2(n13777), .A(n13751), .ZN(P3_U3479) );
  AOI21_X1 U15839 ( .B1(n15316), .B2(n13753), .A(n13752), .ZN(n13810) );
  MUX2_X1 U15840 ( .A(n13754), .B(n13810), .S(n15784), .Z(n13755) );
  OAI21_X1 U15841 ( .B1(n13777), .B2(n13813), .A(n13755), .ZN(P3_U3478) );
  NAND3_X1 U15842 ( .A1(n13757), .A2(n15316), .A3(n13756), .ZN(n13758) );
  OAI211_X1 U15843 ( .C1(n13760), .C2(n15758), .A(n13759), .B(n13758), .ZN(
        n13814) );
  MUX2_X1 U15844 ( .A(P3_REG1_REG_18__SCAN_IN), .B(n13814), .S(n15784), .Z(
        P3_U3477) );
  AOI21_X1 U15845 ( .B1(n15765), .B2(n13762), .A(n13761), .ZN(n13763) );
  OAI21_X1 U15846 ( .B1(n15327), .B2(n13764), .A(n13763), .ZN(n13815) );
  MUX2_X1 U15847 ( .A(P3_REG1_REG_17__SCAN_IN), .B(n13815), .S(n15784), .Z(
        P3_U3476) );
  AOI21_X1 U15848 ( .B1(n13766), .B2(n15316), .A(n13765), .ZN(n13816) );
  MUX2_X1 U15849 ( .A(n13767), .B(n13816), .S(n15784), .Z(n13768) );
  OAI21_X1 U15850 ( .B1(n13819), .B2(n13777), .A(n13768), .ZN(P3_U3475) );
  NAND2_X1 U15851 ( .A1(n13769), .A2(n15316), .ZN(n13770) );
  OAI211_X1 U15852 ( .C1(n13772), .C2(n15758), .A(n13771), .B(n13770), .ZN(
        n13820) );
  MUX2_X1 U15853 ( .A(P3_REG1_REG_15__SCAN_IN), .B(n13820), .S(n15784), .Z(
        P3_U3474) );
  AOI21_X1 U15854 ( .B1(n15316), .B2(n13774), .A(n13773), .ZN(n13821) );
  MUX2_X1 U15855 ( .A(n13775), .B(n13821), .S(n15784), .Z(n13776) );
  OAI21_X1 U15856 ( .B1(n13777), .B2(n13824), .A(n13776), .ZN(P3_U3473) );
  OAI21_X1 U15857 ( .B1(n13780), .B2(n13825), .A(n13779), .ZN(P3_U3455) );
  INV_X1 U15858 ( .A(P3_REG0_REG_26__SCAN_IN), .ZN(n13784) );
  MUX2_X1 U15859 ( .A(n13784), .B(n13783), .S(n15775), .Z(n13785) );
  OAI21_X1 U15860 ( .B1(n9723), .B2(n13825), .A(n13785), .ZN(P3_U3453) );
  INV_X1 U15861 ( .A(P3_REG0_REG_25__SCAN_IN), .ZN(n13787) );
  MUX2_X1 U15862 ( .A(n13787), .B(n13786), .S(n15775), .Z(n13788) );
  OAI21_X1 U15863 ( .B1(n13789), .B2(n13825), .A(n13788), .ZN(P3_U3452) );
  INV_X1 U15864 ( .A(P3_REG0_REG_24__SCAN_IN), .ZN(n13791) );
  MUX2_X1 U15865 ( .A(n13791), .B(n13790), .S(n15775), .Z(n13792) );
  OAI21_X1 U15866 ( .B1(n13793), .B2(n13825), .A(n13792), .ZN(P3_U3451) );
  MUX2_X1 U15867 ( .A(n13795), .B(n13794), .S(n15775), .Z(n13796) );
  OAI21_X1 U15868 ( .B1(n13797), .B2(n13825), .A(n13796), .ZN(P3_U3450) );
  INV_X1 U15869 ( .A(P3_REG0_REG_22__SCAN_IN), .ZN(n13799) );
  MUX2_X1 U15870 ( .A(n13799), .B(n13798), .S(n15775), .Z(n13800) );
  OAI21_X1 U15871 ( .B1(n13801), .B2(n13825), .A(n13800), .ZN(P3_U3449) );
  INV_X1 U15872 ( .A(P3_REG0_REG_21__SCAN_IN), .ZN(n13803) );
  MUX2_X1 U15873 ( .A(n13803), .B(n13802), .S(n15775), .Z(n13804) );
  OAI21_X1 U15874 ( .B1(n13805), .B2(n13825), .A(n13804), .ZN(P3_U3448) );
  INV_X1 U15875 ( .A(P3_REG0_REG_20__SCAN_IN), .ZN(n13807) );
  MUX2_X1 U15876 ( .A(n13807), .B(n13806), .S(n15775), .Z(n13808) );
  OAI21_X1 U15877 ( .B1(n13809), .B2(n13825), .A(n13808), .ZN(P3_U3447) );
  INV_X1 U15878 ( .A(P3_REG0_REG_19__SCAN_IN), .ZN(n13811) );
  MUX2_X1 U15879 ( .A(n13811), .B(n13810), .S(n15775), .Z(n13812) );
  OAI21_X1 U15880 ( .B1(n13825), .B2(n13813), .A(n13812), .ZN(P3_U3446) );
  MUX2_X1 U15881 ( .A(P3_REG0_REG_18__SCAN_IN), .B(n13814), .S(n15775), .Z(
        P3_U3444) );
  MUX2_X1 U15882 ( .A(P3_REG0_REG_17__SCAN_IN), .B(n13815), .S(n15775), .Z(
        P3_U3441) );
  INV_X1 U15883 ( .A(P3_REG0_REG_16__SCAN_IN), .ZN(n13817) );
  MUX2_X1 U15884 ( .A(n13817), .B(n13816), .S(n15775), .Z(n13818) );
  OAI21_X1 U15885 ( .B1(n13819), .B2(n13825), .A(n13818), .ZN(P3_U3438) );
  MUX2_X1 U15886 ( .A(P3_REG0_REG_15__SCAN_IN), .B(n13820), .S(n15775), .Z(
        P3_U3435) );
  INV_X1 U15887 ( .A(P3_REG0_REG_14__SCAN_IN), .ZN(n13822) );
  MUX2_X1 U15888 ( .A(n13822), .B(n13821), .S(n15775), .Z(n13823) );
  OAI21_X1 U15889 ( .B1(n13825), .B2(n13824), .A(n13823), .ZN(P3_U3432) );
  MUX2_X1 U15890 ( .A(P3_D_REG_1__SCAN_IN), .B(n13827), .S(n13826), .Z(
        P3_U3377) );
  NAND2_X1 U15891 ( .A1(n13829), .A2(n13828), .ZN(n13834) );
  INV_X1 U15892 ( .A(P3_IR_REG_30__SCAN_IN), .ZN(n13832) );
  NAND4_X1 U15893 ( .A1(n13831), .A2(P3_IR_REG_31__SCAN_IN), .A3(
        P3_STATE_REG_SCAN_IN), .A4(n13832), .ZN(n13833) );
  OAI211_X1 U15894 ( .C1(n7978), .C2(n13840), .A(n13834), .B(n13833), .ZN(
        P3_U3264) );
  OAI222_X1 U15895 ( .A1(P3_U3151), .A2(n13837), .B1(n13851), .B2(n13836), 
        .C1(n13835), .C2(n13840), .ZN(P3_U3265) );
  INV_X1 U15896 ( .A(n13839), .ZN(n13843) );
  OAI222_X1 U15897 ( .A1(n13851), .A2(n13843), .B1(P3_U3151), .B2(n13842), 
        .C1(n13841), .C2(n13840), .ZN(P3_U3266) );
  INV_X1 U15898 ( .A(n13844), .ZN(n13846) );
  OAI222_X1 U15899 ( .A1(n13851), .A2(n13846), .B1(n13840), .B2(n13845), .C1(
        P3_U3151), .C2(n6945), .ZN(P3_U3268) );
  INV_X1 U15900 ( .A(n13847), .ZN(n13850) );
  OAI222_X1 U15901 ( .A1(n13851), .A2(n13850), .B1(n13840), .B2(n13849), .C1(
        P3_U3151), .C2(n13848), .ZN(P3_U3269) );
  XOR2_X1 U15902 ( .A(n13853), .B(n13852), .Z(n13858) );
  AOI22_X1 U15903 ( .A1(n13965), .A2(n13952), .B1(n13951), .B2(n13967), .ZN(
        n14121) );
  OAI22_X1 U15904 ( .A1(n14121), .A2(n13953), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13854), .ZN(n13856) );
  NOR2_X1 U15905 ( .A1(n14132), .A2(n13958), .ZN(n13855) );
  AOI211_X1 U15906 ( .C1(n13944), .C2(n14129), .A(n13856), .B(n13855), .ZN(
        n13857) );
  OAI21_X1 U15907 ( .B1(n13858), .B2(n13935), .A(n13857), .ZN(P2_U3188) );
  OAI21_X1 U15908 ( .B1(n13861), .B2(n13860), .A(n13859), .ZN(n13862) );
  NAND2_X1 U15909 ( .A1(n13862), .A2(n15345), .ZN(n13867) );
  OAI22_X1 U15910 ( .A1(n13864), .A2(n13915), .B1(n13863), .B2(n13913), .ZN(
        n14183) );
  AND2_X1 U15911 ( .A1(P2_U3088), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n14016) );
  NOR2_X1 U15912 ( .A1(n15354), .A2(n14188), .ZN(n13865) );
  AOI211_X1 U15913 ( .C1(n15347), .C2(n14183), .A(n14016), .B(n13865), .ZN(
        n13866) );
  OAI211_X1 U15914 ( .C1(n13868), .C2(n13958), .A(n13867), .B(n13866), .ZN(
        P2_U3191) );
  INV_X1 U15915 ( .A(n14285), .ZN(n14158) );
  AOI21_X1 U15916 ( .B1(n13870), .B2(n13869), .A(n13935), .ZN(n13872) );
  NAND2_X1 U15917 ( .A1(n13872), .A2(n13871), .ZN(n13877) );
  INV_X1 U15918 ( .A(n13873), .ZN(n14155) );
  AOI22_X1 U15919 ( .A1(n13967), .A2(n13952), .B1(n13951), .B2(n13969), .ZN(
        n14163) );
  OAI22_X1 U15920 ( .A1(n13953), .A2(n14163), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13874), .ZN(n13875) );
  AOI21_X1 U15921 ( .B1(n14155), .B2(n13944), .A(n13875), .ZN(n13876) );
  OAI211_X1 U15922 ( .C1(n14158), .C2(n13958), .A(n13877), .B(n13876), .ZN(
        P2_U3195) );
  AOI211_X1 U15923 ( .C1(n13880), .C2(n13879), .A(n13935), .B(n13878), .ZN(
        n13881) );
  INV_X1 U15924 ( .A(n13881), .ZN(n13885) );
  AOI22_X1 U15925 ( .A1(n13963), .A2(n13952), .B1(n13951), .B2(n13965), .ZN(
        n14086) );
  OAI22_X1 U15926 ( .A1(n14086), .A2(n13953), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13882), .ZN(n13883) );
  AOI21_X1 U15927 ( .B1(n14093), .B2(n13944), .A(n13883), .ZN(n13884) );
  OAI211_X1 U15928 ( .C1(n8889), .C2(n13958), .A(n13885), .B(n13884), .ZN(
        P2_U3197) );
  INV_X1 U15929 ( .A(n13887), .ZN(n13897) );
  AOI21_X1 U15930 ( .B1(n13888), .B2(n13886), .A(n13897), .ZN(n13894) );
  AOI22_X1 U15931 ( .A1(n15347), .A2(n13889), .B1(P2_REG3_REG_16__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13890) );
  OAI21_X1 U15932 ( .B1(n13891), .B2(n15354), .A(n13890), .ZN(n13892) );
  AOI21_X1 U15933 ( .B1(n14376), .B2(n15350), .A(n13892), .ZN(n13893) );
  OAI21_X1 U15934 ( .B1(n13894), .B2(n13935), .A(n13893), .ZN(P2_U3198) );
  NOR3_X1 U15935 ( .A1(n13897), .A2(n7045), .A3(n13896), .ZN(n13900) );
  INV_X1 U15936 ( .A(n13898), .ZN(n13899) );
  OAI21_X1 U15937 ( .B1(n13900), .B2(n13899), .A(n15345), .ZN(n13905) );
  INV_X1 U15938 ( .A(n14225), .ZN(n13903) );
  AOI22_X1 U15939 ( .A1(n13971), .A2(n13952), .B1(n13951), .B2(n13973), .ZN(
        n14219) );
  OAI21_X1 U15940 ( .B1(n13953), .B2(n14219), .A(n13901), .ZN(n13902) );
  AOI21_X1 U15941 ( .B1(n13903), .B2(n13944), .A(n13902), .ZN(n13904) );
  OAI211_X1 U15942 ( .C1(n14229), .C2(n13958), .A(n13905), .B(n13904), .ZN(
        P2_U3200) );
  AOI22_X1 U15943 ( .A1(n13964), .A2(n13952), .B1(n13951), .B2(n13966), .ZN(
        n14101) );
  INV_X1 U15944 ( .A(n14110), .ZN(n13906) );
  AOI22_X1 U15945 ( .A1(n13944), .A2(n13906), .B1(P2_REG3_REG_24__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13907) );
  OAI21_X1 U15946 ( .B1(n14101), .B2(n13953), .A(n13907), .ZN(n13911) );
  AOI211_X1 U15947 ( .C1(n13909), .C2(n13908), .A(n13935), .B(n6757), .ZN(
        n13910) );
  AOI211_X1 U15948 ( .C1(n14343), .C2(n15350), .A(n13911), .B(n13910), .ZN(
        n13912) );
  INV_X1 U15949 ( .A(n13912), .ZN(P2_U3201) );
  OAI22_X1 U15950 ( .A1(n13916), .A2(n13915), .B1(n13914), .B2(n13913), .ZN(
        n14171) );
  AOI22_X1 U15951 ( .A1(n15347), .A2(n14171), .B1(P2_REG3_REG_20__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13917) );
  OAI21_X1 U15952 ( .B1(n14173), .B2(n15354), .A(n13917), .ZN(n13924) );
  INV_X1 U15953 ( .A(n13918), .ZN(n13920) );
  NAND3_X1 U15954 ( .A1(n13859), .A2(n13920), .A3(n13919), .ZN(n13921) );
  AOI21_X1 U15955 ( .B1(n13922), .B2(n13921), .A(n13935), .ZN(n13923) );
  AOI211_X1 U15956 ( .C1(n14289), .C2(n15350), .A(n13924), .B(n13923), .ZN(
        n13925) );
  INV_X1 U15957 ( .A(n13925), .ZN(P2_U3205) );
  XOR2_X1 U15958 ( .A(n13928), .B(n13927), .Z(n13934) );
  AND2_X1 U15959 ( .A1(n13968), .A2(n13951), .ZN(n13929) );
  AOI21_X1 U15960 ( .B1(n13966), .B2(n13952), .A(n13929), .ZN(n14141) );
  OAI22_X1 U15961 ( .A1(n13953), .A2(n14141), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13930), .ZN(n13931) );
  AOI21_X1 U15962 ( .B1(n14145), .B2(n13944), .A(n13931), .ZN(n13933) );
  NAND2_X1 U15963 ( .A1(n14351), .A2(n15350), .ZN(n13932) );
  OAI211_X1 U15964 ( .C1(n13934), .C2(n13935), .A(n13933), .B(n13932), .ZN(
        P2_U3207) );
  AOI21_X1 U15965 ( .B1(n13937), .B2(n13936), .A(n13935), .ZN(n13939) );
  NAND2_X1 U15966 ( .A1(n13939), .A2(n13938), .ZN(n13946) );
  INV_X1 U15967 ( .A(n13940), .ZN(n14209) );
  AND2_X1 U15968 ( .A1(n13972), .A2(n13951), .ZN(n13941) );
  AOI21_X1 U15969 ( .B1(n13970), .B2(n13952), .A(n13941), .ZN(n14202) );
  OAI22_X1 U15970 ( .A1(n13953), .A2(n14202), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13942), .ZN(n13943) );
  AOI21_X1 U15971 ( .B1(n14209), .B2(n13944), .A(n13943), .ZN(n13945) );
  OAI211_X1 U15972 ( .C1(n7151), .C2(n13958), .A(n13946), .B(n13945), .ZN(
        P2_U3210) );
  OAI21_X1 U15973 ( .B1(n13949), .B2(n13948), .A(n13947), .ZN(n13950) );
  NAND2_X1 U15974 ( .A1(n13950), .A2(n15345), .ZN(n13957) );
  NOR2_X1 U15975 ( .A1(n15354), .A2(n14075), .ZN(n13955) );
  AOI22_X1 U15976 ( .A1(n13962), .A2(n13952), .B1(n13951), .B2(n13964), .ZN(
        n14082) );
  NOR2_X1 U15977 ( .A1(n14082), .A2(n13953), .ZN(n13954) );
  AOI211_X1 U15978 ( .C1(P2_REG3_REG_26__SCAN_IN), .C2(P2_U3088), .A(n13955), 
        .B(n13954), .ZN(n13956) );
  OAI211_X1 U15979 ( .C1(n14078), .C2(n13958), .A(n13957), .B(n13956), .ZN(
        P2_U3212) );
  MUX2_X1 U15980 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(n13959), .S(n6672), .Z(
        P2_U3561) );
  MUX2_X1 U15981 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(n13960), .S(n6672), .Z(
        P2_U3560) );
  MUX2_X1 U15982 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(n13961), .S(n6672), .Z(
        P2_U3559) );
  MUX2_X1 U15983 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n13962), .S(n6672), .Z(
        P2_U3558) );
  MUX2_X1 U15984 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(n13963), .S(n6672), .Z(
        P2_U3557) );
  MUX2_X1 U15985 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n13964), .S(n6672), .Z(
        P2_U3556) );
  MUX2_X1 U15986 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(n13965), .S(n6672), .Z(
        P2_U3555) );
  MUX2_X1 U15987 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(n13966), .S(n6672), .Z(
        P2_U3554) );
  MUX2_X1 U15988 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n13967), .S(n6672), .Z(
        P2_U3553) );
  MUX2_X1 U15989 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n13968), .S(n6672), .Z(
        P2_U3552) );
  MUX2_X1 U15990 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n13969), .S(n6672), .Z(
        P2_U3551) );
  MUX2_X1 U15991 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n13970), .S(n6672), .Z(
        P2_U3550) );
  MUX2_X1 U15992 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(n13971), .S(n6672), .Z(
        P2_U3549) );
  MUX2_X1 U15993 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n13972), .S(n6672), .Z(
        P2_U3548) );
  MUX2_X1 U15994 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n13973), .S(n6672), .Z(
        P2_U3547) );
  MUX2_X1 U15995 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(n13974), .S(n6672), .Z(
        P2_U3546) );
  MUX2_X1 U15996 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(n13975), .S(n6672), .Z(
        P2_U3545) );
  MUX2_X1 U15997 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(n13976), .S(n6672), .Z(
        P2_U3544) );
  MUX2_X1 U15998 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(n13977), .S(n6672), .Z(
        P2_U3543) );
  MUX2_X1 U15999 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(n13978), .S(n6672), .Z(
        P2_U3542) );
  MUX2_X1 U16000 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(n13979), .S(n6672), .Z(
        P2_U3541) );
  MUX2_X1 U16001 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(n13980), .S(n6672), .Z(
        P2_U3540) );
  MUX2_X1 U16002 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(n13981), .S(n6672), .Z(
        P2_U3539) );
  MUX2_X1 U16003 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(n13982), .S(n6672), .Z(
        P2_U3538) );
  MUX2_X1 U16004 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(n13983), .S(n6672), .Z(
        P2_U3537) );
  MUX2_X1 U16005 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(n13984), .S(n6672), .Z(
        P2_U3536) );
  MUX2_X1 U16006 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(n13985), .S(n6672), .Z(
        P2_U3535) );
  MUX2_X1 U16007 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(n13986), .S(n6672), .Z(
        P2_U3534) );
  MUX2_X1 U16008 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(n13987), .S(n6672), .Z(
        P2_U3533) );
  MUX2_X1 U16009 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(n13988), .S(n6672), .Z(
        P2_U3532) );
  MUX2_X1 U16010 ( .A(P2_DATAO_REG_0__SCAN_IN), .B(n13989), .S(n6672), .Z(
        P2_U3531) );
  XOR2_X1 U16011 ( .A(n13992), .B(n13991), .Z(n13993) );
  AOI22_X1 U16012 ( .A1(n8364), .A2(n15603), .B1(n15609), .B2(n13993), .ZN(
        n14000) );
  OAI211_X1 U16013 ( .C1(n13996), .C2(n13995), .A(n15604), .B(n13994), .ZN(
        n13999) );
  NAND2_X1 U16014 ( .A1(n15601), .A2(P2_ADDR_REG_2__SCAN_IN), .ZN(n13998) );
  NAND2_X1 U16015 ( .A1(P2_U3088), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n13997) );
  NAND4_X1 U16016 ( .A1(n14000), .A2(n13999), .A3(n13998), .A4(n13997), .ZN(
        P2_U3216) );
  NOR2_X1 U16017 ( .A1(n14002), .A2(n14001), .ZN(n14003) );
  XOR2_X1 U16018 ( .A(n14003), .B(P2_REG2_REG_19__SCAN_IN), .Z(n14013) );
  INV_X1 U16019 ( .A(n14013), .ZN(n14011) );
  NAND2_X1 U16020 ( .A1(n14005), .A2(n14004), .ZN(n14006) );
  NAND2_X1 U16021 ( .A1(n14007), .A2(n14006), .ZN(n14008) );
  XOR2_X1 U16022 ( .A(n14008), .B(P2_REG1_REG_19__SCAN_IN), .Z(n14012) );
  NOR2_X1 U16023 ( .A1(n14012), .A2(n14009), .ZN(n14010) );
  AOI211_X1 U16024 ( .C1(n14011), .C2(n15604), .A(n15603), .B(n14010), .ZN(
        n14015) );
  AOI22_X1 U16025 ( .A1(n14013), .A2(n15604), .B1(n15609), .B2(n14012), .ZN(
        n14014) );
  MUX2_X1 U16026 ( .A(n14015), .B(n14014), .S(n8859), .Z(n14018) );
  AOI21_X1 U16027 ( .B1(n15601), .B2(P2_ADDR_REG_19__SCAN_IN), .A(n14016), 
        .ZN(n14017) );
  NAND2_X1 U16028 ( .A1(n14018), .A2(n14017), .ZN(P2_U3233) );
  NAND2_X1 U16029 ( .A1(n14325), .A2(n14027), .ZN(n14026) );
  XNOR2_X1 U16030 ( .A(n14026), .B(n14020), .ZN(n14021) );
  NAND2_X1 U16031 ( .A1(n14238), .A2(n14160), .ZN(n14025) );
  NOR2_X1 U16032 ( .A1(n14023), .A2(n14022), .ZN(n14237) );
  INV_X1 U16033 ( .A(n14237), .ZN(n14241) );
  NOR2_X1 U16034 ( .A1(n15627), .A2(n14241), .ZN(n14029) );
  AOI21_X1 U16035 ( .B1(n15627), .B2(P2_REG2_REG_31__SCAN_IN), .A(n14029), 
        .ZN(n14024) );
  OAI211_X1 U16036 ( .C1(n14320), .C2(n14157), .A(n14025), .B(n14024), .ZN(
        P2_U3234) );
  OAI211_X1 U16037 ( .C1(n14325), .C2(n14027), .A(n14206), .B(n14026), .ZN(
        n14242) );
  NOR2_X1 U16038 ( .A1(n14325), .A2(n14157), .ZN(n14028) );
  AOI211_X1 U16039 ( .C1(n15627), .C2(P2_REG2_REG_30__SCAN_IN), .A(n14029), 
        .B(n14028), .ZN(n14030) );
  OAI21_X1 U16040 ( .B1(n14213), .B2(n14242), .A(n14030), .ZN(P2_U3235) );
  INV_X1 U16041 ( .A(n14031), .ZN(n14035) );
  INV_X1 U16042 ( .A(n14032), .ZN(n14033) );
  AOI22_X1 U16043 ( .A1(n15627), .A2(P2_REG2_REG_29__SCAN_IN), .B1(n14033), 
        .B2(n14208), .ZN(n14034) );
  OAI21_X1 U16044 ( .B1(n14035), .B2(n14157), .A(n14034), .ZN(n14036) );
  AOI21_X1 U16045 ( .B1(n14037), .B2(n14160), .A(n14036), .ZN(n14039) );
  XNOR2_X1 U16046 ( .A(n14042), .B(n14041), .ZN(n14248) );
  NAND2_X1 U16047 ( .A1(n14043), .A2(n15617), .ZN(n14047) );
  AOI21_X1 U16048 ( .B1(n14056), .B2(n14044), .A(n7171), .ZN(n14046) );
  OAI21_X1 U16049 ( .B1(n14047), .B2(n14046), .A(n14045), .ZN(n14245) );
  INV_X1 U16050 ( .A(n14247), .ZN(n14052) );
  AOI211_X1 U16051 ( .C1(n14247), .C2(n14062), .A(n6670), .B(n14048), .ZN(
        n14246) );
  NAND2_X1 U16052 ( .A1(n14246), .A2(n14160), .ZN(n14051) );
  AOI22_X1 U16053 ( .A1(n14049), .A2(n14208), .B1(n15627), .B2(
        P2_REG2_REG_28__SCAN_IN), .ZN(n14050) );
  OAI211_X1 U16054 ( .C1(n14052), .C2(n14157), .A(n14051), .B(n14050), .ZN(
        n14053) );
  AOI21_X1 U16055 ( .B1(n14245), .B2(n14226), .A(n14053), .ZN(n14054) );
  OAI21_X1 U16056 ( .B1(n14248), .B2(n14234), .A(n14054), .ZN(P2_U3237) );
  XNOR2_X1 U16057 ( .A(n14055), .B(n14057), .ZN(n14332) );
  OAI21_X1 U16058 ( .B1(n14058), .B2(n14057), .A(n14056), .ZN(n14059) );
  NAND2_X1 U16059 ( .A1(n14059), .A2(n15617), .ZN(n14061) );
  NAND2_X1 U16060 ( .A1(n14061), .A2(n14060), .ZN(n14250) );
  INV_X1 U16061 ( .A(n14074), .ZN(n14064) );
  INV_X1 U16062 ( .A(n14062), .ZN(n14063) );
  AOI211_X1 U16063 ( .C1(n14329), .C2(n14064), .A(n6670), .B(n14063), .ZN(
        n14249) );
  NAND2_X1 U16064 ( .A1(n14249), .A2(n14160), .ZN(n14067) );
  AOI22_X1 U16065 ( .A1(n15627), .A2(P2_REG2_REG_27__SCAN_IN), .B1(n14065), 
        .B2(n14208), .ZN(n14066) );
  OAI211_X1 U16066 ( .C1(n14068), .C2(n14157), .A(n14067), .B(n14066), .ZN(
        n14069) );
  AOI21_X1 U16067 ( .B1(n14226), .B2(n14250), .A(n14069), .ZN(n14070) );
  OAI21_X1 U16068 ( .B1(n14332), .B2(n14234), .A(n14070), .ZN(P2_U3238) );
  XNOR2_X1 U16069 ( .A(n14071), .B(n14080), .ZN(n14336) );
  NAND2_X1 U16070 ( .A1(n14256), .A2(n14091), .ZN(n14072) );
  NAND2_X1 U16071 ( .A1(n14072), .A2(n14206), .ZN(n14073) );
  NOR2_X1 U16072 ( .A1(n14074), .A2(n14073), .ZN(n14255) );
  INV_X1 U16073 ( .A(n14075), .ZN(n14076) );
  AOI22_X1 U16074 ( .A1(n15627), .A2(P2_REG2_REG_26__SCAN_IN), .B1(n14076), 
        .B2(n14208), .ZN(n14077) );
  OAI21_X1 U16075 ( .B1(n14078), .B2(n14157), .A(n14077), .ZN(n14079) );
  AOI21_X1 U16076 ( .B1(n14255), .B2(n14160), .A(n14079), .ZN(n14084) );
  NAND2_X1 U16077 ( .A1(n14254), .A2(n14226), .ZN(n14083) );
  OAI211_X1 U16078 ( .C1(n14336), .C2(n14234), .A(n14084), .B(n14083), .ZN(
        P2_U3239) );
  XNOR2_X1 U16079 ( .A(n14085), .B(n14089), .ZN(n14087) );
  OAI21_X1 U16080 ( .B1(n14087), .B2(n14220), .A(n14086), .ZN(n14260) );
  INV_X1 U16081 ( .A(n14260), .ZN(n14098) );
  OAI21_X1 U16082 ( .B1(n6793), .B2(n14089), .A(n14088), .ZN(n14259) );
  INV_X1 U16083 ( .A(n14090), .ZN(n14108) );
  AOI21_X1 U16084 ( .B1(n14262), .B2(n14108), .A(n6670), .ZN(n14092) );
  AND2_X1 U16085 ( .A1(n14092), .A2(n14091), .ZN(n14261) );
  NAND2_X1 U16086 ( .A1(n14261), .A2(n14160), .ZN(n14095) );
  AOI22_X1 U16087 ( .A1(n15627), .A2(P2_REG2_REG_25__SCAN_IN), .B1(n14093), 
        .B2(n14208), .ZN(n14094) );
  OAI211_X1 U16088 ( .C1(n8889), .C2(n14157), .A(n14095), .B(n14094), .ZN(
        n14096) );
  AOI21_X1 U16089 ( .B1(n14259), .B2(n14134), .A(n14096), .ZN(n14097) );
  OAI21_X1 U16090 ( .B1(n15627), .B2(n14098), .A(n14097), .ZN(P2_U3240) );
  OAI21_X1 U16091 ( .B1(n14100), .B2(n14104), .A(n14099), .ZN(n14103) );
  INV_X1 U16092 ( .A(n14101), .ZN(n14102) );
  AOI21_X1 U16093 ( .B1(n14103), .B2(n15617), .A(n14102), .ZN(n14266) );
  AND2_X1 U16094 ( .A1(n14105), .A2(n14104), .ZN(n14106) );
  NOR2_X1 U16095 ( .A1(n14107), .A2(n14106), .ZN(n14344) );
  AOI21_X1 U16096 ( .B1(n14343), .B2(n14127), .A(n6670), .ZN(n14109) );
  NAND2_X1 U16097 ( .A1(n14109), .A2(n14108), .ZN(n14265) );
  INV_X1 U16098 ( .A(P2_REG2_REG_24__SCAN_IN), .ZN(n14111) );
  OAI22_X1 U16099 ( .A1(n14226), .A2(n14111), .B1(n14110), .B2(n15621), .ZN(
        n14112) );
  AOI21_X1 U16100 ( .B1(n14343), .B2(n14228), .A(n14112), .ZN(n14113) );
  OAI21_X1 U16101 ( .B1(n14265), .B2(n14213), .A(n14113), .ZN(n14114) );
  AOI21_X1 U16102 ( .B1(n14344), .B2(n14134), .A(n14114), .ZN(n14115) );
  OAI21_X1 U16103 ( .B1(n15627), .B2(n14266), .A(n14115), .ZN(P2_U3241) );
  INV_X1 U16104 ( .A(n14116), .ZN(n14117) );
  NOR2_X1 U16105 ( .A1(n14118), .A2(n14117), .ZN(n14123) );
  INV_X1 U16106 ( .A(n14125), .ZN(n14119) );
  OAI21_X1 U16107 ( .B1(n14120), .B2(n14119), .A(n15617), .ZN(n14122) );
  OAI21_X1 U16108 ( .B1(n14123), .B2(n14122), .A(n14121), .ZN(n14272) );
  INV_X1 U16109 ( .A(n14272), .ZN(n14136) );
  OAI21_X1 U16110 ( .B1(n14126), .B2(n14125), .A(n14124), .ZN(n14271) );
  OR2_X1 U16111 ( .A1(n6814), .A2(n14132), .ZN(n14128) );
  AND3_X1 U16112 ( .A1(n14128), .A2(n14127), .A3(n14206), .ZN(n14273) );
  NAND2_X1 U16113 ( .A1(n14273), .A2(n14160), .ZN(n14131) );
  AOI22_X1 U16114 ( .A1(n15627), .A2(P2_REG2_REG_23__SCAN_IN), .B1(n14129), 
        .B2(n14208), .ZN(n14130) );
  OAI211_X1 U16115 ( .C1(n14132), .C2(n14157), .A(n14131), .B(n14130), .ZN(
        n14133) );
  AOI21_X1 U16116 ( .B1(n14271), .B2(n14134), .A(n14133), .ZN(n14135) );
  OAI21_X1 U16117 ( .B1(n14136), .B2(n15627), .A(n14135), .ZN(P2_U3242) );
  AOI21_X1 U16118 ( .B1(n6986), .B2(n14138), .A(n14137), .ZN(n14352) );
  INV_X1 U16119 ( .A(n14352), .ZN(n14150) );
  OAI211_X1 U16120 ( .C1(n14140), .C2(n6986), .A(n14139), .B(n15617), .ZN(
        n14142) );
  NAND2_X1 U16121 ( .A1(n14142), .A2(n14141), .ZN(n14279) );
  NAND2_X1 U16122 ( .A1(n14153), .A2(n14351), .ZN(n14143) );
  NAND2_X1 U16123 ( .A1(n14143), .A2(n14206), .ZN(n14144) );
  NOR2_X1 U16124 ( .A1(n6814), .A2(n14144), .ZN(n14278) );
  NAND2_X1 U16125 ( .A1(n14278), .A2(n14160), .ZN(n14147) );
  AOI22_X1 U16126 ( .A1(n15627), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n14145), 
        .B2(n14208), .ZN(n14146) );
  OAI211_X1 U16127 ( .C1(n7144), .C2(n14157), .A(n14147), .B(n14146), .ZN(
        n14148) );
  AOI21_X1 U16128 ( .B1(n14279), .B2(n14226), .A(n14148), .ZN(n14149) );
  OAI21_X1 U16129 ( .B1(n14150), .B2(n14234), .A(n14149), .ZN(P2_U3243) );
  XOR2_X1 U16130 ( .A(n14161), .B(n14151), .Z(n14360) );
  INV_X1 U16131 ( .A(n14153), .ZN(n14154) );
  AOI211_X1 U16132 ( .C1(n14285), .C2(n14176), .A(n6670), .B(n14154), .ZN(
        n14284) );
  AOI22_X1 U16133 ( .A1(n15627), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n14155), 
        .B2(n14208), .ZN(n14156) );
  OAI21_X1 U16134 ( .B1(n14158), .B2(n14157), .A(n14156), .ZN(n14159) );
  AOI21_X1 U16135 ( .B1(n14284), .B2(n14160), .A(n14159), .ZN(n14166) );
  XNOR2_X1 U16136 ( .A(n14162), .B(n14161), .ZN(n14164) );
  OAI21_X1 U16137 ( .B1(n14164), .B2(n14220), .A(n14163), .ZN(n14283) );
  NAND2_X1 U16138 ( .A1(n14283), .A2(n14226), .ZN(n14165) );
  OAI211_X1 U16139 ( .C1(n14360), .C2(n14234), .A(n14166), .B(n14165), .ZN(
        P2_U3244) );
  XOR2_X1 U16140 ( .A(n14170), .B(n14167), .Z(n14292) );
  OAI21_X1 U16141 ( .B1(n14170), .B2(n14169), .A(n14168), .ZN(n14172) );
  AOI21_X1 U16142 ( .B1(n14172), .B2(n15617), .A(n14171), .ZN(n14291) );
  INV_X1 U16143 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n14174) );
  OAI22_X1 U16144 ( .A1(n14226), .A2(n14174), .B1(n14173), .B2(n15621), .ZN(
        n14175) );
  AOI21_X1 U16145 ( .B1(n14289), .B2(n14228), .A(n14175), .ZN(n14179) );
  AOI21_X1 U16146 ( .B1(n14289), .B2(n14192), .A(n6670), .ZN(n14177) );
  AND2_X1 U16147 ( .A1(n14177), .A2(n14176), .ZN(n14288) );
  NAND2_X1 U16148 ( .A1(n14288), .A2(n14160), .ZN(n14178) );
  OAI211_X1 U16149 ( .C1(n14291), .C2(n15627), .A(n14179), .B(n14178), .ZN(
        n14180) );
  INV_X1 U16150 ( .A(n14180), .ZN(n14181) );
  OAI21_X1 U16151 ( .B1(n14234), .B2(n14292), .A(n14181), .ZN(P2_U3245) );
  XOR2_X1 U16152 ( .A(n14182), .B(n14186), .Z(n14185) );
  INV_X1 U16153 ( .A(n14183), .ZN(n14184) );
  OAI21_X1 U16154 ( .B1(n14185), .B2(n14220), .A(n14184), .ZN(n14293) );
  XNOR2_X1 U16155 ( .A(n14187), .B(n14186), .ZN(n14365) );
  INV_X1 U16156 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n14189) );
  OAI22_X1 U16157 ( .A1(n14226), .A2(n14189), .B1(n14188), .B2(n15621), .ZN(
        n14190) );
  AOI21_X1 U16158 ( .B1(n14295), .B2(n14228), .A(n14190), .ZN(n14194) );
  AOI21_X1 U16159 ( .B1(n14295), .B2(n14207), .A(n6670), .ZN(n14191) );
  AND2_X1 U16160 ( .A1(n14192), .A2(n14191), .ZN(n14294) );
  NAND2_X1 U16161 ( .A1(n14294), .A2(n14160), .ZN(n14193) );
  OAI211_X1 U16162 ( .C1(n14365), .C2(n14234), .A(n14194), .B(n14193), .ZN(
        n14195) );
  AOI21_X1 U16163 ( .B1(n14226), .B2(n14293), .A(n14195), .ZN(n14196) );
  INV_X1 U16164 ( .A(n14196), .ZN(P2_U3246) );
  XNOR2_X1 U16165 ( .A(n14197), .B(n14198), .ZN(n14204) );
  NAND2_X1 U16166 ( .A1(n14199), .A2(n14198), .ZN(n14200) );
  NAND2_X1 U16167 ( .A1(n14201), .A2(n14200), .ZN(n14298) );
  NAND2_X1 U16168 ( .A1(n14298), .A2(n15663), .ZN(n14203) );
  OAI211_X1 U16169 ( .C1(n14220), .C2(n14204), .A(n14203), .B(n14202), .ZN(
        n14302) );
  INV_X1 U16170 ( .A(n14302), .ZN(n14217) );
  INV_X1 U16171 ( .A(n15623), .ZN(n14215) );
  NAND2_X1 U16172 ( .A1(n14231), .A2(n14210), .ZN(n14205) );
  NAND3_X1 U16173 ( .A1(n14207), .A2(n14206), .A3(n14205), .ZN(n14299) );
  AOI22_X1 U16174 ( .A1(n15627), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n14209), 
        .B2(n14208), .ZN(n14212) );
  NAND2_X1 U16175 ( .A1(n14210), .A2(n14228), .ZN(n14211) );
  OAI211_X1 U16176 ( .C1(n14299), .C2(n14213), .A(n14212), .B(n14211), .ZN(
        n14214) );
  AOI21_X1 U16177 ( .B1(n14298), .B2(n14215), .A(n14214), .ZN(n14216) );
  OAI21_X1 U16178 ( .B1(n14217), .B2(n15627), .A(n14216), .ZN(P2_U3247) );
  XOR2_X1 U16179 ( .A(n14218), .B(n14223), .Z(n14221) );
  OAI21_X1 U16180 ( .B1(n14221), .B2(n14220), .A(n14219), .ZN(n14305) );
  OAI21_X1 U16181 ( .B1(n14224), .B2(n14223), .A(n14222), .ZN(n14372) );
  OAI22_X1 U16182 ( .A1(n14226), .A2(n11663), .B1(n14225), .B2(n15621), .ZN(
        n14227) );
  AOI21_X1 U16183 ( .B1(n14307), .B2(n14228), .A(n14227), .ZN(n14233) );
  OR2_X1 U16184 ( .A1(n6816), .A2(n14229), .ZN(n14230) );
  AND3_X1 U16185 ( .A1(n14231), .A2(n14206), .A3(n14230), .ZN(n14306) );
  NAND2_X1 U16186 ( .A1(n14306), .A2(n14160), .ZN(n14232) );
  OAI211_X1 U16187 ( .C1(n14372), .C2(n14234), .A(n14233), .B(n14232), .ZN(
        n14235) );
  AOI21_X1 U16188 ( .B1(n14226), .B2(n14305), .A(n14235), .ZN(n14236) );
  INV_X1 U16189 ( .A(n14236), .ZN(P2_U3248) );
  INV_X1 U16190 ( .A(n14313), .ZN(n14270) );
  INV_X1 U16191 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n14239) );
  NOR2_X1 U16192 ( .A1(n14238), .A2(n14237), .ZN(n14317) );
  MUX2_X1 U16193 ( .A(n14239), .B(n14317), .S(n15688), .Z(n14240) );
  OAI21_X1 U16194 ( .B1(n14320), .B2(n14270), .A(n14240), .ZN(P2_U3530) );
  AND2_X1 U16195 ( .A1(n14242), .A2(n14241), .ZN(n14321) );
  MUX2_X1 U16196 ( .A(n14243), .B(n14321), .S(n15688), .Z(n14244) );
  OAI21_X1 U16197 ( .B1(n14325), .B2(n14270), .A(n14244), .ZN(P2_U3529) );
  INV_X1 U16198 ( .A(n15366), .ZN(n15656) );
  MUX2_X1 U16199 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n14326), .S(n15688), .Z(
        P2_U3527) );
  NOR2_X1 U16200 ( .A1(n14250), .A2(n14249), .ZN(n14327) );
  MUX2_X1 U16201 ( .A(n14251), .B(n14327), .S(n15688), .Z(n14253) );
  NAND2_X1 U16202 ( .A1(n14329), .A2(n14313), .ZN(n14252) );
  AOI211_X1 U16203 ( .C1(n15672), .C2(n14256), .A(n14255), .B(n14254), .ZN(
        n14333) );
  MUX2_X1 U16204 ( .A(n14257), .B(n14333), .S(n15688), .Z(n14258) );
  OAI21_X1 U16205 ( .B1(n14336), .B2(n14316), .A(n14258), .ZN(P2_U3525) );
  INV_X1 U16206 ( .A(n14259), .ZN(n14340) );
  AOI211_X1 U16207 ( .C1(n15672), .C2(n14262), .A(n14261), .B(n14260), .ZN(
        n14337) );
  MUX2_X1 U16208 ( .A(n14263), .B(n14337), .S(n15688), .Z(n14264) );
  OAI21_X1 U16209 ( .B1(n14340), .B2(n14316), .A(n14264), .ZN(P2_U3524) );
  AND2_X1 U16210 ( .A1(n14266), .A2(n14265), .ZN(n14342) );
  MUX2_X1 U16211 ( .A(n14342), .B(n14267), .S(n7435), .Z(n14269) );
  NAND2_X1 U16212 ( .A1(n14344), .A2(n14277), .ZN(n14268) );
  OAI211_X1 U16213 ( .C1(n7142), .C2(n14270), .A(n14269), .B(n14268), .ZN(
        P2_U3523) );
  INV_X1 U16214 ( .A(n14271), .ZN(n14350) );
  AOI211_X1 U16215 ( .C1(n15672), .C2(n14274), .A(n14273), .B(n14272), .ZN(
        n14347) );
  MUX2_X1 U16216 ( .A(n14275), .B(n14347), .S(n15688), .Z(n14276) );
  OAI21_X1 U16217 ( .B1(n14350), .B2(n14316), .A(n14276), .ZN(P2_U3522) );
  AOI22_X1 U16218 ( .A1(n14352), .A2(n14277), .B1(n14313), .B2(n14351), .ZN(
        n14282) );
  NOR2_X1 U16219 ( .A1(n14279), .A2(n14278), .ZN(n14354) );
  MUX2_X1 U16220 ( .A(n14354), .B(n14280), .S(n7435), .Z(n14281) );
  NAND2_X1 U16221 ( .A1(n14282), .A2(n14281), .ZN(P2_U3521) );
  AOI211_X1 U16222 ( .C1(n15672), .C2(n14285), .A(n14284), .B(n14283), .ZN(
        n14357) );
  MUX2_X1 U16223 ( .A(n14286), .B(n14357), .S(n15688), .Z(n14287) );
  OAI21_X1 U16224 ( .B1(n14316), .B2(n14360), .A(n14287), .ZN(P2_U3520) );
  AOI21_X1 U16225 ( .B1(n15672), .B2(n14289), .A(n14288), .ZN(n14290) );
  OAI211_X1 U16226 ( .C1(n14292), .C2(n15656), .A(n14291), .B(n14290), .ZN(
        n14361) );
  MUX2_X1 U16227 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n14361), .S(n15688), .Z(
        P2_U3519) );
  AOI211_X1 U16228 ( .C1(n15672), .C2(n14295), .A(n14294), .B(n14293), .ZN(
        n14362) );
  MUX2_X1 U16229 ( .A(n14296), .B(n14362), .S(n15688), .Z(n14297) );
  OAI21_X1 U16230 ( .B1(n14316), .B2(n14365), .A(n14297), .ZN(P2_U3518) );
  INV_X1 U16231 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n14303) );
  NAND2_X1 U16232 ( .A1(n14298), .A2(n15662), .ZN(n14300) );
  OAI211_X1 U16233 ( .C1(n7151), .C2(n15644), .A(n14300), .B(n14299), .ZN(
        n14301) );
  NOR2_X1 U16234 ( .A1(n14302), .A2(n14301), .ZN(n14366) );
  MUX2_X1 U16235 ( .A(n14303), .B(n14366), .S(n15688), .Z(n14304) );
  INV_X1 U16236 ( .A(n14304), .ZN(P2_U3517) );
  AOI211_X1 U16237 ( .C1(n15672), .C2(n14307), .A(n14306), .B(n14305), .ZN(
        n14369) );
  MUX2_X1 U16238 ( .A(n14308), .B(n14369), .S(n15688), .Z(n14309) );
  OAI21_X1 U16239 ( .B1(n14316), .B2(n14372), .A(n14309), .ZN(P2_U3516) );
  NOR2_X1 U16240 ( .A1(n14311), .A2(n14310), .ZN(n14373) );
  MUX2_X1 U16241 ( .A(n14312), .B(n14373), .S(n15688), .Z(n14315) );
  NAND2_X1 U16242 ( .A1(n14376), .A2(n14313), .ZN(n14314) );
  OAI211_X1 U16243 ( .C1(n14316), .C2(n14380), .A(n14315), .B(n14314), .ZN(
        P2_U3515) );
  INV_X1 U16244 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n14318) );
  MUX2_X1 U16245 ( .A(n14318), .B(n14317), .S(n15680), .Z(n14319) );
  OAI21_X1 U16246 ( .B1(n14320), .B2(n14324), .A(n14319), .ZN(P2_U3498) );
  INV_X1 U16247 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n14322) );
  MUX2_X1 U16248 ( .A(n14322), .B(n14321), .S(n15680), .Z(n14323) );
  OAI21_X1 U16249 ( .B1(n14325), .B2(n14324), .A(n14323), .ZN(P2_U3497) );
  MUX2_X1 U16250 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n14326), .S(n15680), .Z(
        P2_U3495) );
  INV_X1 U16251 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n14328) );
  MUX2_X1 U16252 ( .A(n14328), .B(n14327), .S(n15680), .Z(n14331) );
  NAND2_X1 U16253 ( .A1(n14329), .A2(n14375), .ZN(n14330) );
  INV_X1 U16254 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n14334) );
  MUX2_X1 U16255 ( .A(n14334), .B(n14333), .S(n15680), .Z(n14335) );
  OAI21_X1 U16256 ( .B1(n14336), .B2(n14379), .A(n14335), .ZN(P2_U3493) );
  INV_X1 U16257 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n14338) );
  MUX2_X1 U16258 ( .A(n14338), .B(n14337), .S(n15680), .Z(n14339) );
  OAI21_X1 U16259 ( .B1(n14340), .B2(n14379), .A(n14339), .ZN(P2_U3492) );
  INV_X1 U16260 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n14341) );
  MUX2_X1 U16261 ( .A(n14342), .B(n14341), .S(n15678), .Z(n14346) );
  AOI22_X1 U16262 ( .A1(n14344), .A2(n8998), .B1(n14375), .B2(n14343), .ZN(
        n14345) );
  NAND2_X1 U16263 ( .A1(n14346), .A2(n14345), .ZN(P2_U3491) );
  INV_X1 U16264 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n14348) );
  MUX2_X1 U16265 ( .A(n14348), .B(n14347), .S(n15680), .Z(n14349) );
  OAI21_X1 U16266 ( .B1(n14350), .B2(n14379), .A(n14349), .ZN(P2_U3490) );
  AOI22_X1 U16267 ( .A1(n14352), .A2(n8998), .B1(n14375), .B2(n14351), .ZN(
        n14356) );
  INV_X1 U16268 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n14353) );
  MUX2_X1 U16269 ( .A(n14354), .B(n14353), .S(n15678), .Z(n14355) );
  NAND2_X1 U16270 ( .A1(n14356), .A2(n14355), .ZN(P2_U3489) );
  INV_X1 U16271 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n14358) );
  MUX2_X1 U16272 ( .A(n14358), .B(n14357), .S(n15680), .Z(n14359) );
  OAI21_X1 U16273 ( .B1(n14360), .B2(n14379), .A(n14359), .ZN(P2_U3488) );
  MUX2_X1 U16274 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n14361), .S(n15680), .Z(
        P2_U3487) );
  INV_X1 U16275 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n14363) );
  MUX2_X1 U16276 ( .A(n14363), .B(n14362), .S(n15680), .Z(n14364) );
  OAI21_X1 U16277 ( .B1(n14365), .B2(n14379), .A(n14364), .ZN(P2_U3486) );
  INV_X1 U16278 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n14367) );
  MUX2_X1 U16279 ( .A(n14367), .B(n14366), .S(n15680), .Z(n14368) );
  INV_X1 U16280 ( .A(n14368), .ZN(P2_U3484) );
  INV_X1 U16281 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n14370) );
  MUX2_X1 U16282 ( .A(n14370), .B(n14369), .S(n15680), .Z(n14371) );
  OAI21_X1 U16283 ( .B1(n14372), .B2(n14379), .A(n14371), .ZN(P2_U3481) );
  INV_X1 U16284 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n14374) );
  MUX2_X1 U16285 ( .A(n14374), .B(n14373), .S(n15680), .Z(n14378) );
  NAND2_X1 U16286 ( .A1(n14376), .A2(n14375), .ZN(n14377) );
  OAI211_X1 U16287 ( .C1(n14380), .C2(n14379), .A(n14378), .B(n14377), .ZN(
        P2_U3478) );
  INV_X1 U16288 ( .A(n13083), .ZN(n15231) );
  NOR4_X1 U16289 ( .A1(n14382), .A2(P2_IR_REG_30__SCAN_IN), .A3(n14381), .A4(
        P2_U3088), .ZN(n14383) );
  AOI21_X1 U16290 ( .B1(P1_DATAO_REG_31__SCAN_IN), .B2(n14384), .A(n14383), 
        .ZN(n14385) );
  OAI21_X1 U16291 ( .B1(n15231), .B2(n14396), .A(n14385), .ZN(P2_U3296) );
  INV_X1 U16292 ( .A(n14386), .ZN(n15233) );
  OAI222_X1 U16293 ( .A1(n14396), .A2(n15233), .B1(n14388), .B2(P2_U3088), 
        .C1(n14387), .C2(n12861), .ZN(P2_U3298) );
  NAND2_X1 U16294 ( .A1(n15235), .A2(n14389), .ZN(n14391) );
  OAI211_X1 U16295 ( .C1(n12861), .C2(n14392), .A(n14391), .B(n14390), .ZN(
        P2_U3299) );
  INV_X1 U16296 ( .A(n14393), .ZN(n15241) );
  OAI222_X1 U16297 ( .A1(n14396), .A2(n15241), .B1(n14395), .B2(P2_U3088), 
        .C1(n14394), .C2(n12861), .ZN(P2_U3301) );
  MUX2_X1 U16298 ( .A(n14397), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3327) );
  NAND2_X1 U16299 ( .A1(n14866), .A2(n14511), .ZN(n14399) );
  NAND2_X1 U16300 ( .A1(n14688), .A2(n14515), .ZN(n14398) );
  NAND2_X1 U16301 ( .A1(n14399), .A2(n14398), .ZN(n14400) );
  XNOR2_X1 U16302 ( .A(n14400), .B(n14445), .ZN(n14404) );
  NAND2_X1 U16303 ( .A1(n14866), .A2(n14515), .ZN(n14402) );
  NAND2_X1 U16304 ( .A1(n14688), .A2(n14517), .ZN(n14401) );
  NAND2_X1 U16305 ( .A1(n14402), .A2(n14401), .ZN(n14403) );
  NOR2_X1 U16306 ( .A1(n14404), .A2(n14403), .ZN(n14552) );
  AOI21_X1 U16307 ( .B1(n14404), .B2(n14403), .A(n14552), .ZN(n14525) );
  NAND2_X1 U16308 ( .A1(n14406), .A2(n14405), .ZN(n14407) );
  NAND2_X1 U16309 ( .A1(n14408), .A2(n14407), .ZN(n14636) );
  AND2_X1 U16310 ( .A1(n14517), .A2(n14697), .ZN(n14409) );
  AOI21_X1 U16311 ( .B1(n15286), .B2(n9893), .A(n14409), .ZN(n14412) );
  AOI22_X1 U16312 ( .A1(n15286), .A2(n14511), .B1(n9893), .B2(n14697), .ZN(
        n14410) );
  XNOR2_X1 U16313 ( .A(n14410), .B(n14445), .ZN(n14411) );
  XOR2_X1 U16314 ( .A(n14412), .B(n14411), .Z(n14635) );
  INV_X1 U16315 ( .A(n14411), .ZN(n14414) );
  INV_X1 U16316 ( .A(n14412), .ZN(n14413) );
  NAND2_X1 U16317 ( .A1(n14414), .A2(n14413), .ZN(n14415) );
  AOI22_X1 U16318 ( .A1(n15380), .A2(n14511), .B1(n9893), .B2(n14696), .ZN(
        n14416) );
  XNOR2_X1 U16319 ( .A(n14416), .B(n14445), .ZN(n14419) );
  AOI22_X1 U16320 ( .A1(n15380), .A2(n9893), .B1(n14517), .B2(n14696), .ZN(
        n14418) );
  XNOR2_X1 U16321 ( .A(n14419), .B(n14418), .ZN(n15374) );
  INV_X1 U16322 ( .A(n15374), .ZN(n14417) );
  NAND2_X1 U16323 ( .A1(n14419), .A2(n14418), .ZN(n14420) );
  NAND2_X1 U16324 ( .A1(n15196), .A2(n14511), .ZN(n14422) );
  OR2_X1 U16325 ( .A1(n15372), .A2(n14557), .ZN(n14421) );
  NAND2_X1 U16326 ( .A1(n14422), .A2(n14421), .ZN(n14423) );
  XNOR2_X1 U16327 ( .A(n14423), .B(n14445), .ZN(n14424) );
  AOI22_X1 U16328 ( .A1(n15196), .A2(n14515), .B1(n14517), .B2(n14695), .ZN(
        n14674) );
  INV_X1 U16329 ( .A(n14424), .ZN(n14425) );
  NAND2_X1 U16330 ( .A1(n14426), .A2(n14425), .ZN(n14427) );
  NAND2_X1 U16331 ( .A1(n15192), .A2(n14511), .ZN(n14429) );
  NAND2_X1 U16332 ( .A1(n14694), .A2(n9893), .ZN(n14428) );
  NAND2_X1 U16333 ( .A1(n14429), .A2(n14428), .ZN(n14430) );
  XNOR2_X1 U16334 ( .A(n14430), .B(n14445), .ZN(n14431) );
  AOI22_X1 U16335 ( .A1(n15192), .A2(n14515), .B1(n14517), .B2(n14694), .ZN(
        n14432) );
  XNOR2_X1 U16336 ( .A(n14431), .B(n14432), .ZN(n14593) );
  NAND2_X1 U16337 ( .A1(n14594), .A2(n14593), .ZN(n14435) );
  INV_X1 U16338 ( .A(n14431), .ZN(n14433) );
  NAND2_X1 U16339 ( .A1(n14433), .A2(n14432), .ZN(n14434) );
  OAI22_X1 U16340 ( .A1(n15184), .A2(n6667), .B1(n14436), .B2(n14557), .ZN(
        n14437) );
  XNOR2_X1 U16341 ( .A(n14437), .B(n14445), .ZN(n14604) );
  OR2_X1 U16342 ( .A1(n15184), .A2(n14557), .ZN(n14439) );
  NAND2_X1 U16343 ( .A1(n15000), .A2(n14517), .ZN(n14438) );
  NAND2_X1 U16344 ( .A1(n14439), .A2(n14438), .ZN(n14603) );
  NOR2_X1 U16345 ( .A1(n14604), .A2(n14603), .ZN(n14441) );
  NAND2_X1 U16346 ( .A1(n14604), .A2(n14603), .ZN(n14440) );
  OAI22_X1 U16347 ( .A1(n15014), .A2(n6667), .B1(n15022), .B2(n14557), .ZN(
        n14442) );
  XNOR2_X1 U16348 ( .A(n14442), .B(n6921), .ZN(n14450) );
  OAI22_X1 U16349 ( .A1(n15014), .A2(n14557), .B1(n15022), .B2(n6950), .ZN(
        n14449) );
  XNOR2_X1 U16350 ( .A(n14450), .B(n14449), .ZN(n14656) );
  NAND2_X1 U16351 ( .A1(n14448), .A2(n14511), .ZN(n14444) );
  NAND2_X1 U16352 ( .A1(n15003), .A2(n14515), .ZN(n14443) );
  NAND2_X1 U16353 ( .A1(n14444), .A2(n14443), .ZN(n14446) );
  XNOR2_X1 U16354 ( .A(n14446), .B(n9851), .ZN(n14452) );
  AND2_X1 U16355 ( .A1(n15003), .A2(n14517), .ZN(n14447) );
  AOI21_X1 U16356 ( .B1(n14448), .B2(n14515), .A(n14447), .ZN(n14453) );
  XNOR2_X1 U16357 ( .A(n14452), .B(n14453), .ZN(n14544) );
  NOR2_X1 U16358 ( .A1(n14450), .A2(n14449), .ZN(n14545) );
  NOR2_X1 U16359 ( .A1(n14544), .A2(n14545), .ZN(n14451) );
  INV_X1 U16360 ( .A(n14452), .ZN(n14455) );
  INV_X1 U16361 ( .A(n14453), .ZN(n14454) );
  NAND2_X1 U16362 ( .A1(n14455), .A2(n14454), .ZN(n14625) );
  OAI22_X1 U16363 ( .A1(n15166), .A2(n6667), .B1(n14572), .B2(n14557), .ZN(
        n14456) );
  XNOR2_X1 U16364 ( .A(n14456), .B(n14445), .ZN(n14459) );
  OAI22_X1 U16365 ( .A1(n15166), .A2(n14557), .B1(n14572), .B2(n6950), .ZN(
        n14460) );
  NAND2_X1 U16366 ( .A1(n14459), .A2(n14460), .ZN(n14458) );
  AND2_X1 U16367 ( .A1(n14625), .A2(n14458), .ZN(n14457) );
  INV_X1 U16368 ( .A(n14458), .ZN(n14461) );
  XOR2_X1 U16369 ( .A(n14460), .B(n14459), .Z(n14626) );
  OR2_X1 U16370 ( .A1(n14461), .A2(n14626), .ZN(n14462) );
  NAND2_X1 U16371 ( .A1(n15158), .A2(n14511), .ZN(n14465) );
  NAND2_X1 U16372 ( .A1(n14969), .A2(n6676), .ZN(n14464) );
  NAND2_X1 U16373 ( .A1(n14465), .A2(n14464), .ZN(n14466) );
  XNOR2_X1 U16374 ( .A(n14466), .B(n9851), .ZN(n14469) );
  AND2_X1 U16375 ( .A1(n14969), .A2(n14517), .ZN(n14467) );
  AOI21_X1 U16376 ( .B1(n15158), .B2(n14515), .A(n14467), .ZN(n14468) );
  NAND2_X1 U16377 ( .A1(n14469), .A2(n14468), .ZN(n14644) );
  OAI21_X1 U16378 ( .B1(n14469), .B2(n14468), .A(n14644), .ZN(n14570) );
  INV_X1 U16379 ( .A(n14570), .ZN(n14470) );
  NAND2_X1 U16380 ( .A1(n15154), .A2(n14511), .ZN(n14472) );
  NAND2_X1 U16381 ( .A1(n14693), .A2(n14515), .ZN(n14471) );
  NAND2_X1 U16382 ( .A1(n14472), .A2(n14471), .ZN(n14473) );
  XNOR2_X1 U16383 ( .A(n14473), .B(n9851), .ZN(n14475) );
  AND2_X1 U16384 ( .A1(n14693), .A2(n14517), .ZN(n14474) );
  AOI21_X1 U16385 ( .B1(n15154), .B2(n14515), .A(n14474), .ZN(n14476) );
  NAND2_X1 U16386 ( .A1(n14475), .A2(n14476), .ZN(n14534) );
  INV_X1 U16387 ( .A(n14475), .ZN(n14478) );
  INV_X1 U16388 ( .A(n14476), .ZN(n14477) );
  NAND2_X1 U16389 ( .A1(n14478), .A2(n14477), .ZN(n14479) );
  AND2_X1 U16390 ( .A1(n14534), .A2(n14479), .ZN(n14645) );
  NAND2_X1 U16391 ( .A1(n14533), .A2(n14534), .ZN(n14489) );
  NAND2_X1 U16392 ( .A1(n15148), .A2(n14511), .ZN(n14481) );
  NAND2_X1 U16393 ( .A1(n14692), .A2(n14515), .ZN(n14480) );
  NAND2_X1 U16394 ( .A1(n14481), .A2(n14480), .ZN(n14482) );
  XNOR2_X1 U16395 ( .A(n14482), .B(n9851), .ZN(n14484) );
  AND2_X1 U16396 ( .A1(n14517), .A2(n14692), .ZN(n14483) );
  AOI21_X1 U16397 ( .B1(n15148), .B2(n14515), .A(n14483), .ZN(n14485) );
  NAND2_X1 U16398 ( .A1(n14484), .A2(n14485), .ZN(n14612) );
  INV_X1 U16399 ( .A(n14484), .ZN(n14487) );
  INV_X1 U16400 ( .A(n14485), .ZN(n14486) );
  NAND2_X1 U16401 ( .A1(n14487), .A2(n14486), .ZN(n14488) );
  AND2_X1 U16402 ( .A1(n14612), .A2(n14488), .ZN(n14535) );
  NAND2_X1 U16403 ( .A1(n14489), .A2(n14535), .ZN(n14537) );
  NAND2_X1 U16404 ( .A1(n14537), .A2(n14612), .ZN(n14499) );
  NAND2_X1 U16405 ( .A1(n15141), .A2(n14511), .ZN(n14491) );
  NAND2_X1 U16406 ( .A1(n14691), .A2(n14515), .ZN(n14490) );
  NAND2_X1 U16407 ( .A1(n14491), .A2(n14490), .ZN(n14492) );
  XNOR2_X1 U16408 ( .A(n14492), .B(n9851), .ZN(n14494) );
  AND2_X1 U16409 ( .A1(n14517), .A2(n14691), .ZN(n14493) );
  AOI21_X1 U16410 ( .B1(n15141), .B2(n14515), .A(n14493), .ZN(n14495) );
  NAND2_X1 U16411 ( .A1(n14494), .A2(n14495), .ZN(n14580) );
  INV_X1 U16412 ( .A(n14494), .ZN(n14497) );
  INV_X1 U16413 ( .A(n14495), .ZN(n14496) );
  NAND2_X1 U16414 ( .A1(n14497), .A2(n14496), .ZN(n14498) );
  AND2_X1 U16415 ( .A1(n14580), .A2(n14498), .ZN(n14613) );
  NAND2_X1 U16416 ( .A1(n14499), .A2(n14613), .ZN(n14579) );
  NAND2_X1 U16417 ( .A1(n14579), .A2(n14580), .ZN(n14509) );
  NAND2_X1 U16418 ( .A1(n15133), .A2(n14511), .ZN(n14501) );
  NAND2_X1 U16419 ( .A1(n14690), .A2(n14515), .ZN(n14500) );
  NAND2_X1 U16420 ( .A1(n14501), .A2(n14500), .ZN(n14502) );
  XNOR2_X1 U16421 ( .A(n14502), .B(n9851), .ZN(n14504) );
  AND2_X1 U16422 ( .A1(n14517), .A2(n14690), .ZN(n14503) );
  AOI21_X1 U16423 ( .B1(n15133), .B2(n14515), .A(n14503), .ZN(n14505) );
  NAND2_X1 U16424 ( .A1(n14504), .A2(n14505), .ZN(n14510) );
  INV_X1 U16425 ( .A(n14504), .ZN(n14507) );
  INV_X1 U16426 ( .A(n14505), .ZN(n14506) );
  NAND2_X1 U16427 ( .A1(n14507), .A2(n14506), .ZN(n14508) );
  NAND2_X1 U16428 ( .A1(n14509), .A2(n14581), .ZN(n14583) );
  NAND2_X1 U16429 ( .A1(n14516), .A2(n14511), .ZN(n14513) );
  NAND2_X1 U16430 ( .A1(n14689), .A2(n14515), .ZN(n14512) );
  NAND2_X1 U16431 ( .A1(n14513), .A2(n14512), .ZN(n14514) );
  XNOR2_X1 U16432 ( .A(n14514), .B(n14445), .ZN(n14521) );
  NAND2_X1 U16433 ( .A1(n14516), .A2(n14515), .ZN(n14519) );
  NAND2_X1 U16434 ( .A1(n14689), .A2(n14517), .ZN(n14518) );
  NAND2_X1 U16435 ( .A1(n14519), .A2(n14518), .ZN(n14520) );
  NOR2_X1 U16436 ( .A1(n14521), .A2(n14520), .ZN(n14522) );
  AOI21_X1 U16437 ( .B1(n14521), .B2(n14520), .A(n14522), .ZN(n14665) );
  INV_X1 U16438 ( .A(n14522), .ZN(n14523) );
  NAND2_X1 U16439 ( .A1(n14687), .A2(n15002), .ZN(n14527) );
  NAND2_X1 U16440 ( .A1(n14689), .A2(n15001), .ZN(n14526) );
  NAND2_X1 U16441 ( .A1(n14527), .A2(n14526), .ZN(n14863) );
  AOI22_X1 U16442 ( .A1(n14574), .A2(n14863), .B1(P1_REG3_REG_27__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14529) );
  NAND2_X1 U16443 ( .A1(n14680), .A2(n14869), .ZN(n14528) );
  OAI211_X1 U16444 ( .C1(n15121), .C2(n14683), .A(n14529), .B(n14528), .ZN(
        n14530) );
  AOI21_X1 U16445 ( .B1(n14531), .B2(n14675), .A(n14530), .ZN(n14532) );
  INV_X1 U16446 ( .A(n14532), .ZN(P1_U3214) );
  INV_X1 U16447 ( .A(n14533), .ZN(n14647) );
  INV_X1 U16448 ( .A(n14534), .ZN(n14536) );
  NOR3_X1 U16449 ( .A1(n14647), .A2(n14536), .A3(n14535), .ZN(n14538) );
  INV_X1 U16450 ( .A(n14537), .ZN(n14615) );
  OAI21_X1 U16451 ( .B1(n14538), .B2(n14615), .A(n14675), .ZN(n14542) );
  AOI22_X1 U16452 ( .A1(n14693), .A2(n15001), .B1(n15002), .B2(n14691), .ZN(
        n14929) );
  OAI22_X1 U16453 ( .A1(n14929), .A2(n14668), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14539), .ZN(n14540) );
  AOI21_X1 U16454 ( .B1(n14930), .B2(n14680), .A(n14540), .ZN(n14541) );
  OAI211_X1 U16455 ( .C1(n7193), .C2(n14683), .A(n14542), .B(n14541), .ZN(
        P1_U3216) );
  INV_X1 U16456 ( .A(n14543), .ZN(n14654) );
  OAI21_X1 U16457 ( .B1(n14654), .B2(n14545), .A(n14544), .ZN(n14547) );
  NAND3_X1 U16458 ( .A1(n14547), .A2(n14675), .A3(n14546), .ZN(n14551) );
  NAND2_X1 U16459 ( .A1(P1_U3086), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n14841)
         );
  OAI21_X1 U16460 ( .B1(n15384), .B2(n14572), .A(n14841), .ZN(n14549) );
  NOR2_X1 U16461 ( .A1(n15402), .A2(n14990), .ZN(n14548) );
  AOI211_X1 U16462 ( .C1(n14677), .C2(n14988), .A(n14549), .B(n14548), .ZN(
        n14550) );
  OAI211_X1 U16463 ( .C1(n15173), .C2(n14683), .A(n14551), .B(n14550), .ZN(
        P1_U3219) );
  OAI22_X1 U16464 ( .A1(n14563), .A2(n6667), .B1(n14556), .B2(n14557), .ZN(
        n14554) );
  XNOR2_X1 U16465 ( .A(n14554), .B(n14445), .ZN(n14559) );
  OAI22_X1 U16466 ( .A1(n14563), .A2(n14557), .B1(n14556), .B2(n6950), .ZN(
        n14558) );
  XNOR2_X1 U16467 ( .A(n14559), .B(n14558), .ZN(n14560) );
  AOI22_X1 U16468 ( .A1(n14677), .A2(n14688), .B1(P1_REG3_REG_28__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14561) );
  OAI21_X1 U16469 ( .B1(n14562), .B2(n15384), .A(n14561), .ZN(n14565) );
  NOR2_X1 U16470 ( .A1(n14563), .A2(n14683), .ZN(n14564) );
  AOI211_X1 U16471 ( .C1(n14566), .C2(n14680), .A(n14565), .B(n14564), .ZN(
        n14567) );
  OAI21_X1 U16472 ( .B1(n14568), .B2(n15392), .A(n14567), .ZN(P1_U3220) );
  AOI21_X1 U16473 ( .B1(n14571), .B2(n14570), .A(n6719), .ZN(n14578) );
  OAI22_X1 U16474 ( .A1(n14573), .A2(n15091), .B1(n14572), .B2(n15069), .ZN(
        n14954) );
  AOI22_X1 U16475 ( .A1(n14954), .A2(n14574), .B1(P1_REG3_REG_21__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14575) );
  OAI21_X1 U16476 ( .B1(n15402), .B2(n14956), .A(n14575), .ZN(n14576) );
  AOI21_X1 U16477 ( .B1(n15158), .B2(n15397), .A(n14576), .ZN(n14577) );
  OAI21_X1 U16478 ( .B1(n14578), .B2(n15392), .A(n14577), .ZN(P1_U3223) );
  INV_X1 U16479 ( .A(n15133), .ZN(n14592) );
  INV_X1 U16480 ( .A(n14579), .ZN(n14616) );
  INV_X1 U16481 ( .A(n14580), .ZN(n14582) );
  NOR3_X1 U16482 ( .A1(n14616), .A2(n14582), .A3(n14581), .ZN(n14585) );
  INV_X1 U16483 ( .A(n14583), .ZN(n14584) );
  OAI21_X1 U16484 ( .B1(n14585), .B2(n14584), .A(n14675), .ZN(n14591) );
  NAND2_X1 U16485 ( .A1(n14691), .A2(n15001), .ZN(n14587) );
  NAND2_X1 U16486 ( .A1(n14689), .A2(n15002), .ZN(n14586) );
  AND2_X1 U16487 ( .A1(n14587), .A2(n14586), .ZN(n15131) );
  OAI22_X1 U16488 ( .A1(n14668), .A2(n15131), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14588), .ZN(n14589) );
  AOI21_X1 U16489 ( .B1(n14680), .B2(n14890), .A(n14589), .ZN(n14590) );
  OAI211_X1 U16490 ( .C1(n14592), .C2(n14683), .A(n14591), .B(n14590), .ZN(
        P1_U3225) );
  XOR2_X1 U16491 ( .A(n14594), .B(n14593), .Z(n14601) );
  OR2_X1 U16492 ( .A1(n15372), .A2(n15069), .ZN(n14596) );
  NAND2_X1 U16493 ( .A1(n15000), .A2(n15002), .ZN(n14595) );
  AND2_X1 U16494 ( .A1(n14596), .A2(n14595), .ZN(n15041) );
  NAND2_X1 U16495 ( .A1(n14680), .A2(n15046), .ZN(n14598) );
  OAI211_X1 U16496 ( .C1(n15041), .C2(n14668), .A(n14598), .B(n14597), .ZN(
        n14599) );
  AOI21_X1 U16497 ( .B1(n15192), .B2(n15397), .A(n14599), .ZN(n14600) );
  OAI21_X1 U16498 ( .B1(n14601), .B2(n15392), .A(n14600), .ZN(P1_U3226) );
  XNOR2_X1 U16499 ( .A(n14604), .B(n14603), .ZN(n14605) );
  XNOR2_X1 U16500 ( .A(n14602), .B(n14605), .ZN(n14611) );
  NAND2_X1 U16501 ( .A1(n14677), .A2(n14694), .ZN(n14607) );
  OAI211_X1 U16502 ( .C1(n15022), .C2(n15384), .A(n14607), .B(n14606), .ZN(
        n14609) );
  NOR2_X1 U16503 ( .A1(n15184), .A2(n14683), .ZN(n14608) );
  AOI211_X1 U16504 ( .C1(n15028), .C2(n14680), .A(n14609), .B(n14608), .ZN(
        n14610) );
  OAI21_X1 U16505 ( .B1(n14611), .B2(n15392), .A(n14610), .ZN(P1_U3228) );
  INV_X1 U16506 ( .A(n15141), .ZN(n14917) );
  INV_X1 U16507 ( .A(n14612), .ZN(n14614) );
  NOR3_X1 U16508 ( .A1(n14615), .A2(n14614), .A3(n14613), .ZN(n14617) );
  OAI21_X1 U16509 ( .B1(n14617), .B2(n14616), .A(n14675), .ZN(n14624) );
  NAND2_X1 U16510 ( .A1(n14692), .A2(n15001), .ZN(n14619) );
  NAND2_X1 U16511 ( .A1(n14690), .A2(n15002), .ZN(n14618) );
  NAND2_X1 U16512 ( .A1(n14619), .A2(n14618), .ZN(n14912) );
  INV_X1 U16513 ( .A(n14912), .ZN(n14621) );
  OAI22_X1 U16514 ( .A1(n14621), .A2(n14668), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14620), .ZN(n14622) );
  AOI21_X1 U16515 ( .B1(n14680), .B2(n14914), .A(n14622), .ZN(n14623) );
  OAI211_X1 U16516 ( .C1(n14917), .C2(n14683), .A(n14624), .B(n14623), .ZN(
        P1_U3229) );
  NAND2_X1 U16517 ( .A1(n14546), .A2(n14625), .ZN(n14627) );
  XNOR2_X1 U16518 ( .A(n14627), .B(n14626), .ZN(n14633) );
  OAI22_X1 U16519 ( .A1(n14941), .A2(n15384), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14628), .ZN(n14629) );
  AOI21_X1 U16520 ( .B1(n14677), .B2(n15003), .A(n14629), .ZN(n14630) );
  OAI21_X1 U16521 ( .B1(n15402), .B2(n14972), .A(n14630), .ZN(n14631) );
  AOI21_X1 U16522 ( .B1(n14977), .B2(n15397), .A(n14631), .ZN(n14632) );
  OAI21_X1 U16523 ( .B1(n14633), .B2(n15392), .A(n14632), .ZN(P1_U3233) );
  OAI211_X1 U16524 ( .C1(n14636), .C2(n14635), .A(n14634), .B(n14675), .ZN(
        n14643) );
  OR2_X1 U16525 ( .A1(n14637), .A2(n15091), .ZN(n14639) );
  OR2_X1 U16526 ( .A1(n15385), .A2(n15069), .ZN(n14638) );
  AND2_X1 U16527 ( .A1(n14639), .A2(n14638), .ZN(n15281) );
  OAI21_X1 U16528 ( .B1(n15281), .B2(n14668), .A(n14640), .ZN(n14641) );
  AOI21_X1 U16529 ( .B1(n14680), .B2(n15284), .A(n14641), .ZN(n14642) );
  OAI211_X1 U16530 ( .C1(n12359), .C2(n14683), .A(n14643), .B(n14642), .ZN(
        P1_U3234) );
  INV_X1 U16531 ( .A(n14644), .ZN(n14646) );
  NOR3_X1 U16532 ( .A1(n6719), .A2(n14646), .A3(n14645), .ZN(n14648) );
  OAI21_X1 U16533 ( .B1(n14648), .B2(n14647), .A(n14675), .ZN(n14653) );
  INV_X1 U16534 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n14649) );
  OAI22_X1 U16535 ( .A1(n15384), .A2(n14942), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14649), .ZN(n14651) );
  NOR2_X1 U16536 ( .A1(n15402), .A2(n14948), .ZN(n14650) );
  AOI211_X1 U16537 ( .C1(n14677), .C2(n14969), .A(n14651), .B(n14650), .ZN(
        n14652) );
  OAI211_X1 U16538 ( .C1(n14683), .C2(n14946), .A(n14653), .B(n14652), .ZN(
        P1_U3235) );
  AOI21_X1 U16539 ( .B1(n14656), .B2(n14655), .A(n14654), .ZN(n14662) );
  NAND2_X1 U16540 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n14816)
         );
  OAI21_X1 U16541 ( .B1(n15384), .B2(n14657), .A(n14816), .ZN(n14658) );
  AOI21_X1 U16542 ( .B1(n14677), .B2(n15000), .A(n14658), .ZN(n14659) );
  OAI21_X1 U16543 ( .B1(n15402), .B2(n15009), .A(n14659), .ZN(n14660) );
  AOI21_X1 U16544 ( .B1(n15180), .B2(n15397), .A(n14660), .ZN(n14661) );
  OAI21_X1 U16545 ( .B1(n14662), .B2(n15392), .A(n14661), .ZN(P1_U3238) );
  OAI21_X1 U16546 ( .B1(n14665), .B2(n14664), .A(n14663), .ZN(n14666) );
  NAND2_X1 U16547 ( .A1(n14666), .A2(n14675), .ZN(n14671) );
  AOI22_X1 U16548 ( .A1(n15001), .A2(n14690), .B1(n14688), .B2(n15002), .ZN(
        n15123) );
  OAI22_X1 U16549 ( .A1(n15123), .A2(n14668), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14667), .ZN(n14669) );
  AOI21_X1 U16550 ( .B1(n14680), .B2(n14880), .A(n14669), .ZN(n14670) );
  OAI211_X1 U16551 ( .C1(n15125), .C2(n14683), .A(n14671), .B(n14670), .ZN(
        P1_U3240) );
  OAI21_X1 U16552 ( .B1(n14674), .B2(n14673), .A(n14672), .ZN(n14676) );
  NAND2_X1 U16553 ( .A1(n14676), .A2(n14675), .ZN(n14682) );
  NAND2_X1 U16554 ( .A1(n14677), .A2(n14696), .ZN(n14678) );
  NAND2_X1 U16555 ( .A1(P1_U3086), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n15474)
         );
  OAI211_X1 U16556 ( .C1(n15021), .C2(n15384), .A(n14678), .B(n15474), .ZN(
        n14679) );
  AOI21_X1 U16557 ( .B1(n14680), .B2(n6812), .A(n14679), .ZN(n14681) );
  OAI211_X1 U16558 ( .C1(n14684), .C2(n14683), .A(n14682), .B(n14681), .ZN(
        P1_U3241) );
  MUX2_X1 U16559 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(n14848), .S(n14723), .Z(
        P1_U3591) );
  MUX2_X1 U16560 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n14685), .S(n14723), .Z(
        P1_U3590) );
  MUX2_X1 U16561 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n14686), .S(n14723), .Z(
        P1_U3589) );
  MUX2_X1 U16562 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n14687), .S(n14723), .Z(
        P1_U3588) );
  MUX2_X1 U16563 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n14688), .S(n14723), .Z(
        P1_U3587) );
  MUX2_X1 U16564 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n14689), .S(n14723), .Z(
        P1_U3586) );
  MUX2_X1 U16565 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n14690), .S(n14723), .Z(
        P1_U3585) );
  MUX2_X1 U16566 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n14691), .S(n14723), .Z(
        P1_U3584) );
  MUX2_X1 U16567 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n14692), .S(n14723), .Z(
        P1_U3583) );
  MUX2_X1 U16568 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n14693), .S(n14723), .Z(
        P1_U3582) );
  MUX2_X1 U16569 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n14969), .S(n14723), .Z(
        P1_U3581) );
  MUX2_X1 U16570 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n14989), .S(n14723), .Z(
        P1_U3580) );
  MUX2_X1 U16571 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n15003), .S(n14723), .Z(
        P1_U3579) );
  MUX2_X1 U16572 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n15000), .S(n14723), .Z(
        P1_U3577) );
  MUX2_X1 U16573 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n14694), .S(P1_U4016), .Z(
        P1_U3576) );
  MUX2_X1 U16574 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n14695), .S(P1_U4016), .Z(
        P1_U3575) );
  MUX2_X1 U16575 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n14696), .S(P1_U4016), .Z(
        P1_U3574) );
  MUX2_X1 U16576 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n14697), .S(P1_U4016), .Z(
        P1_U3573) );
  MUX2_X1 U16577 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n14698), .S(P1_U4016), .Z(
        P1_U3571) );
  MUX2_X1 U16578 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n14699), .S(P1_U4016), .Z(
        P1_U3570) );
  MUX2_X1 U16579 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n14700), .S(P1_U4016), .Z(
        P1_U3569) );
  MUX2_X1 U16580 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n14701), .S(P1_U4016), .Z(
        P1_U3568) );
  MUX2_X1 U16581 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n14702), .S(P1_U4016), .Z(
        P1_U3567) );
  MUX2_X1 U16582 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n14703), .S(P1_U4016), .Z(
        P1_U3566) );
  MUX2_X1 U16583 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n14704), .S(P1_U4016), .Z(
        P1_U3565) );
  MUX2_X1 U16584 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n14705), .S(P1_U4016), .Z(
        P1_U3564) );
  MUX2_X1 U16585 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n10689), .S(P1_U4016), .Z(
        P1_U3562) );
  MUX2_X1 U16586 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n14706), .S(P1_U4016), .Z(
        P1_U3561) );
  MUX2_X1 U16587 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(n14707), .S(P1_U4016), .Z(
        P1_U3560) );
  OAI22_X1 U16588 ( .A1(n15476), .A2(n7748), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14708), .ZN(n14709) );
  AOI21_X1 U16589 ( .B1(n7341), .B2(n15457), .A(n14709), .ZN(n14717) );
  MUX2_X1 U16590 ( .A(P1_REG1_REG_1__SCAN_IN), .B(n10169), .S(n14710), .Z(
        n14711) );
  OAI21_X1 U16591 ( .B1(n9873), .B2(n14712), .A(n14711), .ZN(n14713) );
  NAND3_X1 U16592 ( .A1(n14833), .A2(n14731), .A3(n14713), .ZN(n14716) );
  OAI211_X1 U16593 ( .C1(n14720), .C2(n14714), .A(n14838), .B(n14737), .ZN(
        n14715) );
  NAND3_X1 U16594 ( .A1(n14717), .A2(n14716), .A3(n14715), .ZN(P1_U3244) );
  MUX2_X1 U16595 ( .A(n14720), .B(n14719), .S(n14718), .Z(n14722) );
  NAND2_X1 U16596 ( .A1(n14722), .A2(n14721), .ZN(n14724) );
  OAI211_X1 U16597 ( .C1(P1_IR_REG_0__SCAN_IN), .C2(n14725), .A(n14724), .B(
        n14723), .ZN(n15458) );
  INV_X1 U16598 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n14727) );
  OAI22_X1 U16599 ( .A1(n15476), .A2(n14727), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14726), .ZN(n14728) );
  AOI21_X1 U16600 ( .B1(n14729), .B2(n15457), .A(n14728), .ZN(n14742) );
  MUX2_X1 U16601 ( .A(P1_REG1_REG_2__SCAN_IN), .B(n10168), .S(n14734), .Z(
        n14732) );
  NAND3_X1 U16602 ( .A1(n14732), .A2(n14731), .A3(n14730), .ZN(n14733) );
  NAND3_X1 U16603 ( .A1(n14833), .A2(n14748), .A3(n14733), .ZN(n14741) );
  MUX2_X1 U16604 ( .A(P1_REG2_REG_2__SCAN_IN), .B(n14735), .S(n14734), .Z(
        n14738) );
  NAND3_X1 U16605 ( .A1(n14738), .A2(n14737), .A3(n14736), .ZN(n14739) );
  NAND3_X1 U16606 ( .A1(n14838), .A2(n14753), .A3(n14739), .ZN(n14740) );
  NAND4_X1 U16607 ( .A1(n15458), .A2(n14742), .A3(n14741), .A4(n14740), .ZN(
        P1_U3245) );
  INV_X1 U16608 ( .A(n14750), .ZN(n14745) );
  OAI22_X1 U16609 ( .A1(n15476), .A2(n7804), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14743), .ZN(n14744) );
  AOI21_X1 U16610 ( .B1(n14745), .B2(n15457), .A(n14744), .ZN(n14757) );
  MUX2_X1 U16611 ( .A(P1_REG1_REG_3__SCAN_IN), .B(n10176), .S(n14750), .Z(
        n14747) );
  NAND3_X1 U16612 ( .A1(n14748), .A2(n14747), .A3(n14746), .ZN(n14749) );
  NAND3_X1 U16613 ( .A1(n14833), .A2(n15446), .A3(n14749), .ZN(n14756) );
  MUX2_X1 U16614 ( .A(P1_REG2_REG_3__SCAN_IN), .B(n11533), .S(n14750), .Z(
        n14752) );
  NAND3_X1 U16615 ( .A1(n14753), .A2(n14752), .A3(n14751), .ZN(n14754) );
  NAND3_X1 U16616 ( .A1(n14838), .A2(n15451), .A3(n14754), .ZN(n14755) );
  NAND3_X1 U16617 ( .A1(n14757), .A2(n14756), .A3(n14755), .ZN(P1_U3246) );
  OAI21_X1 U16618 ( .B1(n15476), .B2(n14759), .A(n14758), .ZN(n14760) );
  AOI21_X1 U16619 ( .B1(n15457), .B2(n14761), .A(n14760), .ZN(n14773) );
  OAI21_X1 U16620 ( .B1(n14764), .B2(n14763), .A(n14762), .ZN(n14765) );
  NAND2_X1 U16621 ( .A1(n14833), .A2(n14765), .ZN(n14772) );
  MUX2_X1 U16622 ( .A(P1_REG2_REG_5__SCAN_IN), .B(n10194), .S(n14766), .Z(
        n14769) );
  INV_X1 U16623 ( .A(n14767), .ZN(n14768) );
  NAND2_X1 U16624 ( .A1(n14769), .A2(n14768), .ZN(n14770) );
  OAI211_X1 U16625 ( .C1(n15453), .C2(n14770), .A(n14838), .B(n14784), .ZN(
        n14771) );
  NAND3_X1 U16626 ( .A1(n14773), .A2(n14772), .A3(n14771), .ZN(P1_U3248) );
  INV_X1 U16627 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n14775) );
  OAI21_X1 U16628 ( .B1(n15476), .B2(n14775), .A(n14774), .ZN(n14776) );
  AOI21_X1 U16629 ( .B1(n15457), .B2(n14777), .A(n14776), .ZN(n14790) );
  NAND2_X1 U16630 ( .A1(n14779), .A2(n14778), .ZN(n14780) );
  NAND3_X1 U16631 ( .A1(n14833), .A2(n14781), .A3(n14780), .ZN(n14789) );
  MUX2_X1 U16632 ( .A(P1_REG2_REG_6__SCAN_IN), .B(n11588), .S(n14782), .Z(
        n14785) );
  NAND3_X1 U16633 ( .A1(n14785), .A2(n14784), .A3(n14783), .ZN(n14786) );
  NAND3_X1 U16634 ( .A1(n14838), .A2(n14787), .A3(n14786), .ZN(n14788) );
  NAND3_X1 U16635 ( .A1(n14790), .A2(n14789), .A3(n14788), .ZN(P1_U3249) );
  OAI21_X1 U16636 ( .B1(n15476), .B2(n14792), .A(n14791), .ZN(n14793) );
  AOI21_X1 U16637 ( .B1(n15457), .B2(n14800), .A(n14793), .ZN(n14808) );
  INV_X1 U16638 ( .A(n14794), .ZN(n14799) );
  NOR3_X1 U16639 ( .A1(n14797), .A2(n14796), .A3(n14795), .ZN(n14798) );
  OAI21_X1 U16640 ( .B1(n14799), .B2(n14798), .A(n14833), .ZN(n14807) );
  MUX2_X1 U16641 ( .A(n10367), .B(P1_REG2_REG_9__SCAN_IN), .S(n14800), .Z(
        n14801) );
  NAND3_X1 U16642 ( .A1(n14803), .A2(n14802), .A3(n14801), .ZN(n14804) );
  NAND3_X1 U16643 ( .A1(n14838), .A2(n14805), .A3(n14804), .ZN(n14806) );
  NAND3_X1 U16644 ( .A1(n14808), .A2(n14807), .A3(n14806), .ZN(P1_U3252) );
  NAND2_X1 U16645 ( .A1(n14811), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n14809) );
  NAND2_X1 U16646 ( .A1(n14810), .A2(n14809), .ZN(n14829) );
  XNOR2_X1 U16647 ( .A(n14829), .B(n14822), .ZN(n14827) );
  XNOR2_X1 U16648 ( .A(n14827), .B(P1_REG2_REG_18__SCAN_IN), .ZN(n14821) );
  AOI22_X1 U16649 ( .A1(n14813), .A2(n14812), .B1(n14811), .B2(
        P1_REG1_REG_17__SCAN_IN), .ZN(n14823) );
  XNOR2_X1 U16650 ( .A(n14823), .B(n14828), .ZN(n14814) );
  NAND2_X1 U16651 ( .A1(n14814), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n14825) );
  OAI211_X1 U16652 ( .C1(P1_REG1_REG_18__SCAN_IN), .C2(n14814), .A(n14833), 
        .B(n14825), .ZN(n14815) );
  NAND2_X1 U16653 ( .A1(n14816), .A2(n14815), .ZN(n14818) );
  NOR2_X1 U16654 ( .A1(n15472), .A2(n14822), .ZN(n14817) );
  AOI211_X1 U16655 ( .C1(n14819), .C2(P1_ADDR_REG_18__SCAN_IN), .A(n14818), 
        .B(n14817), .ZN(n14820) );
  OAI21_X1 U16656 ( .B1(n14821), .B2(n15470), .A(n14820), .ZN(P1_U3261) );
  OR2_X1 U16657 ( .A1(n14823), .A2(n14822), .ZN(n14824) );
  NAND2_X1 U16658 ( .A1(n14825), .A2(n14824), .ZN(n14826) );
  XOR2_X1 U16659 ( .A(n14826), .B(P1_REG1_REG_19__SCAN_IN), .Z(n14835) );
  NAND2_X1 U16660 ( .A1(n14827), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n14831) );
  NAND2_X1 U16661 ( .A1(n14829), .A2(n14828), .ZN(n14830) );
  NAND2_X1 U16662 ( .A1(n14831), .A2(n14830), .ZN(n14832) );
  XOR2_X1 U16663 ( .A(n14832), .B(P1_REG2_REG_19__SCAN_IN), .Z(n14834) );
  AOI22_X1 U16664 ( .A1(n14835), .A2(n14833), .B1(n14838), .B2(n14834), .ZN(
        n14840) );
  INV_X1 U16665 ( .A(n14834), .ZN(n14837) );
  NOR2_X1 U16666 ( .A1(n14835), .A2(n15468), .ZN(n14836) );
  AOI211_X1 U16667 ( .C1(n14838), .C2(n14837), .A(n15457), .B(n14836), .ZN(
        n14839) );
  MUX2_X1 U16668 ( .A(n14840), .B(n14839), .S(n15048), .Z(n14842) );
  OAI211_X1 U16669 ( .C1(n8233), .C2(n15476), .A(n14842), .B(n14841), .ZN(
        P1_U3262) );
  NOR2_X1 U16670 ( .A1(n14843), .A2(n14851), .ZN(n14845) );
  XNOR2_X1 U16671 ( .A(n14845), .B(n14844), .ZN(n14846) );
  NAND2_X1 U16672 ( .A1(n14846), .A2(n15291), .ZN(n15099) );
  NAND2_X1 U16673 ( .A1(n14848), .A2(n14847), .ZN(n15101) );
  NOR2_X1 U16674 ( .A1(n15067), .A2(n15101), .ZN(n14854) );
  NOR2_X1 U16675 ( .A1(n15100), .A2(n15013), .ZN(n14849) );
  AOI211_X1 U16676 ( .C1(n15067), .C2(P1_REG2_REG_31__SCAN_IN), .A(n14854), 
        .B(n14849), .ZN(n14850) );
  OAI21_X1 U16677 ( .B1(n15099), .B2(n14994), .A(n14850), .ZN(P1_U3263) );
  XNOR2_X1 U16678 ( .A(n15103), .B(n14851), .ZN(n14852) );
  NAND2_X1 U16679 ( .A1(n14852), .A2(n15291), .ZN(n15102) );
  NOR2_X1 U16680 ( .A1(n15103), .A2(n15013), .ZN(n14853) );
  AOI211_X1 U16681 ( .C1(n15067), .C2(P1_REG2_REG_30__SCAN_IN), .A(n14854), 
        .B(n14853), .ZN(n14855) );
  OAI21_X1 U16682 ( .B1(n14994), .B2(n15102), .A(n14855), .ZN(P1_U3264) );
  XNOR2_X1 U16683 ( .A(n14856), .B(n14857), .ZN(n14858) );
  NAND2_X1 U16684 ( .A1(n14858), .A2(n15280), .ZN(n14865) );
  NAND2_X1 U16685 ( .A1(n14860), .A2(n14859), .ZN(n14861) );
  NAND2_X1 U16686 ( .A1(n14862), .A2(n14861), .ZN(n15118) );
  AOI21_X1 U16687 ( .B1(n14866), .B2(n14879), .A(n15488), .ZN(n14868) );
  NAND2_X1 U16688 ( .A1(n14868), .A2(n14867), .ZN(n15119) );
  NOR2_X1 U16689 ( .A1(n15119), .A2(n14994), .ZN(n14872) );
  AOI22_X1 U16690 ( .A1(n15067), .A2(P1_REG2_REG_27__SCAN_IN), .B1(n14869), 
        .B2(n15283), .ZN(n14870) );
  OAI21_X1 U16691 ( .B1(n15121), .B2(n15013), .A(n14870), .ZN(n14871) );
  AOI211_X1 U16692 ( .C1(n15118), .C2(n15086), .A(n14872), .B(n14871), .ZN(
        n14873) );
  OAI21_X1 U16693 ( .B1(n6740), .B2(n15067), .A(n14873), .ZN(P1_U3266) );
  XNOR2_X1 U16694 ( .A(n14874), .B(n14876), .ZN(n15129) );
  OAI21_X1 U16695 ( .B1(n14877), .B2(n14876), .A(n14875), .ZN(n14878) );
  INV_X1 U16696 ( .A(n14878), .ZN(n15127) );
  OAI211_X1 U16697 ( .C1(n15125), .C2(n14899), .A(n15291), .B(n14879), .ZN(
        n15124) );
  INV_X1 U16698 ( .A(n14880), .ZN(n14881) );
  OAI22_X1 U16699 ( .A1(n15067), .A2(n15123), .B1(n14881), .B2(n15058), .ZN(
        n14883) );
  NOR2_X1 U16700 ( .A1(n15125), .A2(n15013), .ZN(n14882) );
  AOI211_X1 U16701 ( .C1(n15067), .C2(P1_REG2_REG_26__SCAN_IN), .A(n14883), 
        .B(n14882), .ZN(n14884) );
  OAI21_X1 U16702 ( .B1(n14994), .B2(n15124), .A(n14884), .ZN(n14885) );
  AOI21_X1 U16703 ( .B1(n15127), .B2(n15294), .A(n14885), .ZN(n14886) );
  OAI21_X1 U16704 ( .B1(n15129), .B2(n14887), .A(n14886), .ZN(P1_U3267) );
  OAI21_X1 U16705 ( .B1(n7267), .B2(n7266), .A(n14889), .ZN(n15130) );
  NAND2_X1 U16706 ( .A1(n15130), .A2(n15090), .ZN(n14903) );
  INV_X1 U16707 ( .A(P1_REG2_REG_25__SCAN_IN), .ZN(n14894) );
  NAND2_X1 U16708 ( .A1(n15283), .A2(n14890), .ZN(n14891) );
  NAND2_X1 U16709 ( .A1(n15131), .A2(n14891), .ZN(n14892) );
  NAND2_X1 U16710 ( .A1(n14892), .A2(n15093), .ZN(n14893) );
  OAI21_X1 U16711 ( .B1(n15093), .B2(n14894), .A(n14893), .ZN(n14895) );
  AOI21_X1 U16712 ( .B1(n15133), .B2(n15285), .A(n14895), .ZN(n14902) );
  NAND2_X1 U16713 ( .A1(n14897), .A2(n7266), .ZN(n15134) );
  NAND3_X1 U16714 ( .A1(n14896), .A2(n15134), .A3(n15294), .ZN(n14901) );
  AND2_X1 U16715 ( .A1(n15133), .A2(n14913), .ZN(n14898) );
  NOR2_X1 U16716 ( .A1(n14899), .A2(n14898), .ZN(n15135) );
  NAND2_X1 U16717 ( .A1(n15135), .A2(n15094), .ZN(n14900) );
  NAND4_X1 U16718 ( .A1(n14903), .A2(n14902), .A3(n14901), .A4(n14900), .ZN(
        P1_U3268) );
  INV_X1 U16719 ( .A(n14904), .ZN(n14906) );
  OAI21_X1 U16720 ( .B1(n14906), .B2(n14910), .A(n14905), .ZN(n15140) );
  INV_X1 U16721 ( .A(n14907), .ZN(n14908) );
  AOI211_X1 U16722 ( .C1(n14910), .C2(n14909), .A(n15481), .B(n14908), .ZN(
        n14911) );
  AOI211_X1 U16723 ( .C1(n15080), .C2(n15140), .A(n14912), .B(n14911), .ZN(
        n15144) );
  AOI21_X1 U16724 ( .B1(n15141), .B2(n14923), .A(n12530), .ZN(n15142) );
  NAND2_X1 U16725 ( .A1(n15142), .A2(n15094), .ZN(n14916) );
  AOI22_X1 U16726 ( .A1(n15067), .A2(P1_REG2_REG_24__SCAN_IN), .B1(n14914), 
        .B2(n15283), .ZN(n14915) );
  OAI211_X1 U16727 ( .C1(n14917), .C2(n15013), .A(n14916), .B(n14915), .ZN(
        n14918) );
  AOI21_X1 U16728 ( .B1(n15140), .B2(n15086), .A(n14918), .ZN(n14919) );
  OAI21_X1 U16729 ( .B1(n15144), .B2(n15067), .A(n14919), .ZN(P1_U3269) );
  OAI21_X1 U16730 ( .B1(n14922), .B2(n14921), .A(n14920), .ZN(n15151) );
  INV_X1 U16731 ( .A(n14923), .ZN(n14924) );
  AOI211_X1 U16732 ( .C1(n15148), .C2(n14944), .A(n15488), .B(n14924), .ZN(
        n15146) );
  INV_X1 U16733 ( .A(n15146), .ZN(n14932) );
  OAI21_X1 U16734 ( .B1(n14927), .B2(n14926), .A(n14925), .ZN(n14928) );
  NAND2_X1 U16735 ( .A1(n14928), .A2(n15280), .ZN(n15150) );
  INV_X1 U16736 ( .A(n14929), .ZN(n15147) );
  AOI21_X1 U16737 ( .B1(n14930), .B2(n15283), .A(n15147), .ZN(n14931) );
  OAI211_X1 U16738 ( .C1(n15048), .C2(n14932), .A(n15150), .B(n14931), .ZN(
        n14933) );
  NAND2_X1 U16739 ( .A1(n14933), .A2(n15093), .ZN(n14935) );
  AOI22_X1 U16740 ( .A1(n15148), .A2(n15285), .B1(P1_REG2_REG_23__SCAN_IN), 
        .B2(n15067), .ZN(n14934) );
  OAI211_X1 U16741 ( .C1(n15151), .C2(n15063), .A(n14935), .B(n14934), .ZN(
        P1_U3270) );
  XNOR2_X1 U16742 ( .A(n14937), .B(n14936), .ZN(n15156) );
  XNOR2_X1 U16743 ( .A(n14939), .B(n14938), .ZN(n14940) );
  OAI222_X1 U16744 ( .A1(n15091), .A2(n14942), .B1(n15069), .B2(n14941), .C1(
        n15481), .C2(n14940), .ZN(n15152) );
  NAND2_X1 U16745 ( .A1(n15152), .A2(n15093), .ZN(n14952) );
  INV_X1 U16746 ( .A(n14944), .ZN(n14945) );
  AOI211_X1 U16747 ( .C1(n15154), .C2(n7197), .A(n15488), .B(n14945), .ZN(
        n15153) );
  NOR2_X1 U16748 ( .A1(n14946), .A2(n15013), .ZN(n14950) );
  OAI22_X1 U16749 ( .A1(n14948), .A2(n15058), .B1(n15093), .B2(n14947), .ZN(
        n14949) );
  AOI211_X1 U16750 ( .C1(n15153), .C2(n15293), .A(n14950), .B(n14949), .ZN(
        n14951) );
  OAI211_X1 U16751 ( .C1(n15156), .C2(n15063), .A(n14952), .B(n14951), .ZN(
        P1_U3271) );
  XOR2_X1 U16752 ( .A(n14953), .B(n14963), .Z(n14955) );
  AOI21_X1 U16753 ( .B1(n14955), .B2(n15280), .A(n14954), .ZN(n15160) );
  AOI211_X1 U16754 ( .C1(n15158), .C2(n14974), .A(n15488), .B(n14943), .ZN(
        n15157) );
  INV_X1 U16755 ( .A(n15158), .ZN(n14959) );
  INV_X1 U16756 ( .A(n14956), .ZN(n14957) );
  AOI22_X1 U16757 ( .A1(n15067), .A2(P1_REG2_REG_21__SCAN_IN), .B1(n14957), 
        .B2(n15283), .ZN(n14958) );
  OAI21_X1 U16758 ( .B1(n14959), .B2(n15013), .A(n14958), .ZN(n14965) );
  INV_X1 U16759 ( .A(n14960), .ZN(n14961) );
  AOI21_X1 U16760 ( .B1(n14963), .B2(n14962), .A(n14961), .ZN(n15161) );
  NOR2_X1 U16761 ( .A1(n15161), .A2(n15063), .ZN(n14964) );
  AOI211_X1 U16762 ( .C1(n15157), .C2(n15293), .A(n14965), .B(n14964), .ZN(
        n14966) );
  OAI21_X1 U16763 ( .B1(n15067), .B2(n15160), .A(n14966), .ZN(P1_U3272) );
  OAI211_X1 U16764 ( .C1(n14968), .C2(n14979), .A(n14967), .B(n15280), .ZN(
        n14971) );
  AOI22_X1 U16765 ( .A1(n14969), .A2(n15002), .B1(n15001), .B2(n15003), .ZN(
        n14970) );
  NAND2_X1 U16766 ( .A1(n14971), .A2(n14970), .ZN(n15168) );
  INV_X1 U16767 ( .A(n15168), .ZN(n14982) );
  INV_X1 U16768 ( .A(P1_REG2_REG_20__SCAN_IN), .ZN(n14973) );
  OAI22_X1 U16769 ( .A1(n15093), .A2(n14973), .B1(n14972), .B2(n15058), .ZN(
        n14976) );
  OAI211_X1 U16770 ( .C1(n15166), .C2(n14986), .A(n15291), .B(n14974), .ZN(
        n15164) );
  NOR2_X1 U16771 ( .A1(n15164), .A2(n14994), .ZN(n14975) );
  AOI211_X1 U16772 ( .C1(n15285), .C2(n14977), .A(n14976), .B(n14975), .ZN(
        n14981) );
  NAND2_X1 U16773 ( .A1(n14978), .A2(n14979), .ZN(n15162) );
  NAND3_X1 U16774 ( .A1(n15163), .A2(n15162), .A3(n15294), .ZN(n14980) );
  OAI211_X1 U16775 ( .C1(n14982), .C2(n15067), .A(n14981), .B(n14980), .ZN(
        P1_U3273) );
  XNOR2_X1 U16776 ( .A(n14983), .B(n14985), .ZN(n15177) );
  OAI21_X1 U16777 ( .B1(n7740), .B2(n14985), .A(n14984), .ZN(n15175) );
  NOR2_X1 U16778 ( .A1(n15007), .A2(n15173), .ZN(n14987) );
  AOI22_X1 U16779 ( .A1(n14989), .A2(n15002), .B1(n15001), .B2(n14988), .ZN(
        n15171) );
  OAI22_X1 U16780 ( .A1(n15171), .A2(n15067), .B1(n14990), .B2(n15058), .ZN(
        n14992) );
  NOR2_X1 U16781 ( .A1(n15173), .A2(n15013), .ZN(n14991) );
  AOI211_X1 U16782 ( .C1(n15067), .C2(P1_REG2_REG_19__SCAN_IN), .A(n14992), 
        .B(n14991), .ZN(n14993) );
  OAI21_X1 U16783 ( .B1(n14994), .B2(n15172), .A(n14993), .ZN(n14995) );
  AOI21_X1 U16784 ( .B1(n15175), .B2(n15090), .A(n14995), .ZN(n14996) );
  OAI21_X1 U16785 ( .B1(n15063), .B2(n15177), .A(n14996), .ZN(P1_U3274) );
  XNOR2_X1 U16786 ( .A(n14997), .B(n14999), .ZN(n15178) );
  XNOR2_X1 U16787 ( .A(n14998), .B(n14999), .ZN(n15005) );
  AOI22_X1 U16788 ( .A1(n15003), .A2(n15002), .B1(n15001), .B2(n15000), .ZN(
        n15004) );
  OAI21_X1 U16789 ( .B1(n15005), .B2(n15481), .A(n15004), .ZN(n15006) );
  AOI21_X1 U16790 ( .B1(n15080), .B2(n15178), .A(n15006), .ZN(n15182) );
  INV_X1 U16791 ( .A(n15027), .ZN(n15008) );
  AOI211_X1 U16792 ( .C1(n15180), .C2(n15008), .A(n15488), .B(n15007), .ZN(
        n15179) );
  NAND2_X1 U16793 ( .A1(n15179), .A2(n15293), .ZN(n15012) );
  INV_X1 U16794 ( .A(n15009), .ZN(n15010) );
  AOI22_X1 U16795 ( .A1(n15067), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n15010), 
        .B2(n15283), .ZN(n15011) );
  OAI211_X1 U16796 ( .C1(n15014), .C2(n15013), .A(n15012), .B(n15011), .ZN(
        n15015) );
  AOI21_X1 U16797 ( .B1(n15178), .B2(n15086), .A(n15015), .ZN(n15016) );
  OAI21_X1 U16798 ( .B1(n15182), .B2(n15067), .A(n15016), .ZN(P1_U3275) );
  XNOR2_X1 U16799 ( .A(n15017), .B(n15018), .ZN(n15189) );
  AOI21_X1 U16800 ( .B1(n15020), .B2(n15019), .A(n15481), .ZN(n15025) );
  OAI22_X1 U16801 ( .A1(n15022), .A2(n15091), .B1(n15021), .B2(n15069), .ZN(
        n15023) );
  AOI21_X1 U16802 ( .B1(n15025), .B2(n15024), .A(n15023), .ZN(n15188) );
  INV_X1 U16803 ( .A(n15188), .ZN(n15036) );
  AND2_X1 U16804 ( .A1(n15043), .A2(n15032), .ZN(n15026) );
  OR2_X1 U16805 ( .A1(n15027), .A2(n15026), .ZN(n15185) );
  INV_X1 U16806 ( .A(n15028), .ZN(n15029) );
  OAI22_X1 U16807 ( .A1(n15093), .A2(n15030), .B1(n15029), .B2(n15058), .ZN(
        n15031) );
  AOI21_X1 U16808 ( .B1(n15032), .B2(n15285), .A(n15031), .ZN(n15033) );
  OAI21_X1 U16809 ( .B1(n15185), .B2(n15034), .A(n15033), .ZN(n15035) );
  AOI21_X1 U16810 ( .B1(n15036), .B2(n15093), .A(n15035), .ZN(n15037) );
  OAI21_X1 U16811 ( .B1(n15063), .B2(n15189), .A(n15037), .ZN(P1_U3276) );
  XNOR2_X1 U16812 ( .A(n15038), .B(n15040), .ZN(n15194) );
  XNOR2_X1 U16813 ( .A(n15039), .B(n15040), .ZN(n15042) );
  OAI21_X1 U16814 ( .B1(n15042), .B2(n15481), .A(n15041), .ZN(n15190) );
  INV_X1 U16815 ( .A(n15043), .ZN(n15044) );
  AOI211_X1 U16816 ( .C1(n15192), .C2(n15045), .A(n15488), .B(n15044), .ZN(
        n15191) );
  INV_X1 U16817 ( .A(n15191), .ZN(n15049) );
  INV_X1 U16818 ( .A(n15046), .ZN(n15047) );
  OAI22_X1 U16819 ( .A1(n15049), .A2(n15048), .B1(n15058), .B2(n15047), .ZN(
        n15050) );
  OAI21_X1 U16820 ( .B1(n15190), .B2(n15050), .A(n15093), .ZN(n15052) );
  AOI22_X1 U16821 ( .A1(n15192), .A2(n15285), .B1(P1_REG2_REG_16__SCAN_IN), 
        .B2(n15067), .ZN(n15051) );
  OAI211_X1 U16822 ( .C1(n15194), .C2(n15063), .A(n15052), .B(n15051), .ZN(
        P1_U3277) );
  NAND2_X1 U16823 ( .A1(n15380), .A2(n15290), .ZN(n15053) );
  NAND2_X1 U16824 ( .A1(n15053), .A2(n15291), .ZN(n15054) );
  NOR2_X1 U16825 ( .A1(n6815), .A2(n15054), .ZN(n15203) );
  OAI22_X1 U16826 ( .A1(n15373), .A2(n15069), .B1(n15372), .B2(n15091), .ZN(
        n15204) );
  XOR2_X1 U16827 ( .A(n15060), .B(n15055), .Z(n15056) );
  NAND2_X1 U16828 ( .A1(n15056), .A2(n15280), .ZN(n15206) );
  INV_X1 U16829 ( .A(n15206), .ZN(n15057) );
  AOI211_X1 U16830 ( .C1(n15203), .C2(n12593), .A(n15204), .B(n15057), .ZN(
        n15068) );
  OAI22_X1 U16831 ( .A1(n15093), .A2(n10616), .B1(n15383), .B2(n15058), .ZN(
        n15065) );
  INV_X1 U16832 ( .A(n15060), .ZN(n15062) );
  OAI21_X1 U16833 ( .B1(n15059), .B2(n15062), .A(n15061), .ZN(n15207) );
  NOR2_X1 U16834 ( .A1(n15207), .A2(n15063), .ZN(n15064) );
  AOI211_X1 U16835 ( .C1(n15285), .C2(n15380), .A(n15065), .B(n15064), .ZN(
        n15066) );
  OAI21_X1 U16836 ( .B1(n15068), .B2(n15067), .A(n15066), .ZN(P1_U3279) );
  OAI21_X1 U16837 ( .B1(n12794), .B2(n15073), .A(n15280), .ZN(n15070) );
  NAND2_X1 U16838 ( .A1(n15070), .A2(n15069), .ZN(n15076) );
  NAND2_X1 U16839 ( .A1(n15485), .A2(n15085), .ZN(n15071) );
  NAND2_X1 U16840 ( .A1(n15072), .A2(n15071), .ZN(n15489) );
  XNOR2_X1 U16841 ( .A(n15092), .B(n15489), .ZN(n15074) );
  OAI21_X1 U16842 ( .B1(n15074), .B2(n15481), .A(n15073), .ZN(n15075) );
  NAND2_X1 U16843 ( .A1(n15076), .A2(n15075), .ZN(n15082) );
  OR2_X1 U16844 ( .A1(n12794), .A2(n15077), .ZN(n15078) );
  NAND2_X1 U16845 ( .A1(n15079), .A2(n15078), .ZN(n15492) );
  NAND2_X1 U16846 ( .A1(n15492), .A2(n15080), .ZN(n15081) );
  OAI211_X1 U16847 ( .C1(n10688), .C2(n15091), .A(n15082), .B(n15081), .ZN(
        n15490) );
  MUX2_X1 U16848 ( .A(n15490), .B(P1_REG2_REG_1__SCAN_IN), .S(n15067), .Z(
        n15083) );
  INV_X1 U16849 ( .A(n15083), .ZN(n15089) );
  INV_X1 U16850 ( .A(n15489), .ZN(n15084) );
  AOI22_X1 U16851 ( .A1(n15094), .A2(n15084), .B1(P1_REG3_REG_1__SCAN_IN), 
        .B2(n15283), .ZN(n15088) );
  AOI22_X1 U16852 ( .A1(n15086), .A2(n15492), .B1(n15285), .B2(n15085), .ZN(
        n15087) );
  NAND3_X1 U16853 ( .A1(n15089), .A2(n15088), .A3(n15087), .ZN(P1_U3292) );
  OAI21_X1 U16854 ( .B1(n15090), .B2(n15294), .A(n15479), .ZN(n15098) );
  NOR2_X1 U16855 ( .A1(n15092), .A2(n15091), .ZN(n15484) );
  AOI22_X1 U16856 ( .A1(n15484), .A2(n15093), .B1(P1_REG3_REG_0__SCAN_IN), 
        .B2(n15283), .ZN(n15097) );
  OAI21_X1 U16857 ( .B1(n15094), .B2(n15285), .A(n15485), .ZN(n15096) );
  NAND2_X1 U16858 ( .A1(n15067), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n15095) );
  NAND4_X1 U16859 ( .A1(n15098), .A2(n15097), .A3(n15096), .A4(n15095), .ZN(
        P1_U3293) );
  OAI211_X1 U16860 ( .C1(n15100), .C2(n15518), .A(n15099), .B(n15101), .ZN(
        n15208) );
  MUX2_X1 U16861 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n15208), .S(n15537), .Z(
        P1_U3559) );
  OAI211_X1 U16862 ( .C1(n15103), .C2(n15518), .A(n15102), .B(n15101), .ZN(
        n15209) );
  MUX2_X1 U16863 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n15209), .S(n15537), .Z(
        P1_U3558) );
  NAND2_X1 U16864 ( .A1(n15104), .A2(n15495), .ZN(n15107) );
  NAND2_X1 U16865 ( .A1(n15111), .A2(n15413), .ZN(n15116) );
  AOI21_X1 U16866 ( .B1(n15113), .B2(n15495), .A(n15112), .ZN(n15114) );
  OAI211_X1 U16867 ( .C1(n15117), .C2(n15116), .A(n15115), .B(n15114), .ZN(
        n15210) );
  MUX2_X1 U16868 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n15210), .S(n15537), .Z(
        P1_U3556) );
  INV_X1 U16869 ( .A(n15499), .ZN(n15523) );
  NAND2_X1 U16870 ( .A1(n15118), .A2(n15523), .ZN(n15120) );
  OAI211_X1 U16871 ( .C1(n15121), .C2(n15518), .A(n15120), .B(n15119), .ZN(
        n15122) );
  OAI211_X1 U16872 ( .C1(n15125), .C2(n15518), .A(n15124), .B(n15123), .ZN(
        n15126) );
  AOI21_X1 U16873 ( .B1(n15127), .B2(n15413), .A(n15126), .ZN(n15128) );
  OAI21_X1 U16874 ( .B1(n15129), .B2(n15481), .A(n15128), .ZN(n15212) );
  MUX2_X1 U16875 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n15212), .S(n15537), .Z(
        P1_U3554) );
  NAND2_X1 U16876 ( .A1(n15130), .A2(n15280), .ZN(n15139) );
  INV_X1 U16877 ( .A(n15131), .ZN(n15132) );
  AOI21_X1 U16878 ( .B1(n15133), .B2(n15495), .A(n15132), .ZN(n15138) );
  NAND3_X1 U16879 ( .A1(n14896), .A2(n15413), .A3(n15134), .ZN(n15137) );
  NAND2_X1 U16880 ( .A1(n15135), .A2(n15291), .ZN(n15136) );
  NAND4_X1 U16881 ( .A1(n15139), .A2(n15138), .A3(n15137), .A4(n15136), .ZN(
        n15213) );
  MUX2_X1 U16882 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n15213), .S(n15537), .Z(
        P1_U3553) );
  INV_X1 U16883 ( .A(n15140), .ZN(n15145) );
  AOI22_X1 U16884 ( .A1(n15142), .A2(n15291), .B1(n15141), .B2(n15495), .ZN(
        n15143) );
  OAI211_X1 U16885 ( .C1(n15145), .C2(n15499), .A(n15144), .B(n15143), .ZN(
        n15214) );
  MUX2_X1 U16886 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n15214), .S(n15537), .Z(
        P1_U3552) );
  AOI211_X1 U16887 ( .C1(n15148), .C2(n15495), .A(n15147), .B(n15146), .ZN(
        n15149) );
  OAI211_X1 U16888 ( .C1(n15151), .C2(n15482), .A(n15150), .B(n15149), .ZN(
        n15215) );
  MUX2_X1 U16889 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n15215), .S(n15537), .Z(
        P1_U3551) );
  AOI211_X1 U16890 ( .C1(n15154), .C2(n15495), .A(n15153), .B(n15152), .ZN(
        n15155) );
  OAI21_X1 U16891 ( .B1(n15482), .B2(n15156), .A(n15155), .ZN(n15216) );
  MUX2_X1 U16892 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n15216), .S(n15537), .Z(
        P1_U3550) );
  AOI21_X1 U16893 ( .B1(n15158), .B2(n15495), .A(n15157), .ZN(n15159) );
  OAI211_X1 U16894 ( .C1(n15161), .C2(n15482), .A(n15160), .B(n15159), .ZN(
        n15217) );
  MUX2_X1 U16895 ( .A(n15217), .B(P1_REG1_REG_21__SCAN_IN), .S(n15534), .Z(
        P1_U3549) );
  INV_X1 U16896 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n15169) );
  NAND3_X1 U16897 ( .A1(n15163), .A2(n15162), .A3(n15413), .ZN(n15165) );
  OAI211_X1 U16898 ( .C1(n15166), .C2(n15518), .A(n15165), .B(n15164), .ZN(
        n15167) );
  NOR2_X1 U16899 ( .A1(n15168), .A2(n15167), .ZN(n15218) );
  MUX2_X1 U16900 ( .A(n15169), .B(n15218), .S(n15537), .Z(n15170) );
  INV_X1 U16901 ( .A(n15170), .ZN(P1_U3548) );
  OAI211_X1 U16902 ( .C1(n15173), .C2(n15518), .A(n15172), .B(n15171), .ZN(
        n15174) );
  AOI21_X1 U16903 ( .B1(n15175), .B2(n15280), .A(n15174), .ZN(n15176) );
  OAI21_X1 U16904 ( .B1(n15482), .B2(n15177), .A(n15176), .ZN(n15221) );
  MUX2_X1 U16905 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n15221), .S(n15537), .Z(
        P1_U3547) );
  INV_X1 U16906 ( .A(n15178), .ZN(n15183) );
  AOI21_X1 U16907 ( .B1(n15180), .B2(n15495), .A(n15179), .ZN(n15181) );
  OAI211_X1 U16908 ( .C1(n15183), .C2(n15499), .A(n15182), .B(n15181), .ZN(
        n15222) );
  MUX2_X1 U16909 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n15222), .S(n15537), .Z(
        P1_U3546) );
  OAI22_X1 U16910 ( .A1(n15185), .A2(n15488), .B1(n15184), .B2(n15518), .ZN(
        n15186) );
  INV_X1 U16911 ( .A(n15186), .ZN(n15187) );
  OAI211_X1 U16912 ( .C1(n15482), .C2(n15189), .A(n15188), .B(n15187), .ZN(
        n15223) );
  MUX2_X1 U16913 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n15223), .S(n15537), .Z(
        P1_U3545) );
  AOI211_X1 U16914 ( .C1(n15192), .C2(n15495), .A(n15191), .B(n15190), .ZN(
        n15193) );
  OAI21_X1 U16915 ( .B1(n15482), .B2(n15194), .A(n15193), .ZN(n15224) );
  MUX2_X1 U16916 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n15224), .S(n15537), .Z(
        P1_U3544) );
  AOI21_X1 U16917 ( .B1(n15196), .B2(n15495), .A(n15195), .ZN(n15197) );
  OAI21_X1 U16918 ( .B1(n15198), .B2(n15488), .A(n15197), .ZN(n15199) );
  AOI21_X1 U16919 ( .B1(n15200), .B2(n15413), .A(n15199), .ZN(n15201) );
  OAI21_X1 U16920 ( .B1(n15481), .B2(n15202), .A(n15201), .ZN(n15225) );
  MUX2_X1 U16921 ( .A(P1_REG1_REG_15__SCAN_IN), .B(n15225), .S(n15537), .Z(
        P1_U3543) );
  AOI211_X1 U16922 ( .C1(n15380), .C2(n15495), .A(n15204), .B(n15203), .ZN(
        n15205) );
  OAI211_X1 U16923 ( .C1(n15482), .C2(n15207), .A(n15206), .B(n15205), .ZN(
        n15226) );
  MUX2_X1 U16924 ( .A(n15226), .B(P1_REG1_REG_14__SCAN_IN), .S(n15534), .Z(
        P1_U3542) );
  MUX2_X1 U16925 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n15208), .S(n15526), .Z(
        P1_U3527) );
  MUX2_X1 U16926 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n15209), .S(n15526), .Z(
        P1_U3526) );
  MUX2_X1 U16927 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n15210), .S(n15526), .Z(
        P1_U3524) );
  MUX2_X1 U16928 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n15212), .S(n15526), .Z(
        P1_U3522) );
  MUX2_X1 U16929 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n15213), .S(n15526), .Z(
        P1_U3521) );
  MUX2_X1 U16930 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n15214), .S(n15526), .Z(
        P1_U3520) );
  MUX2_X1 U16931 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n15215), .S(n15526), .Z(
        P1_U3519) );
  MUX2_X1 U16932 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n15216), .S(n15526), .Z(
        P1_U3518) );
  MUX2_X1 U16933 ( .A(n15217), .B(P1_REG0_REG_21__SCAN_IN), .S(n15524), .Z(
        P1_U3517) );
  INV_X1 U16934 ( .A(P1_REG0_REG_20__SCAN_IN), .ZN(n15219) );
  MUX2_X1 U16935 ( .A(n15219), .B(n15218), .S(n15526), .Z(n15220) );
  INV_X1 U16936 ( .A(n15220), .ZN(P1_U3516) );
  MUX2_X1 U16937 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n15221), .S(n15526), .Z(
        P1_U3515) );
  MUX2_X1 U16938 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n15222), .S(n15526), .Z(
        P1_U3513) );
  MUX2_X1 U16939 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n15223), .S(n15526), .Z(
        P1_U3510) );
  MUX2_X1 U16940 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n15224), .S(n15526), .Z(
        P1_U3507) );
  MUX2_X1 U16941 ( .A(P1_REG0_REG_15__SCAN_IN), .B(n15225), .S(n15526), .Z(
        P1_U3504) );
  MUX2_X1 U16942 ( .A(n15226), .B(P1_REG0_REG_14__SCAN_IN), .S(n15524), .Z(
        P1_U3501) );
  NOR4_X1 U16943 ( .A1(n7722), .A2(P1_IR_REG_30__SCAN_IN), .A3(P1_U3086), .A4(
        n15227), .ZN(n15228) );
  AOI21_X1 U16944 ( .B1(P2_DATAO_REG_31__SCAN_IN), .B2(n15229), .A(n15228), 
        .ZN(n15230) );
  OAI21_X1 U16945 ( .B1(n15231), .B2(n15238), .A(n15230), .ZN(P1_U3324) );
  INV_X1 U16946 ( .A(n15235), .ZN(n15237) );
  OAI222_X1 U16947 ( .A1(n15242), .A2(P1_U3086), .B1(n15238), .B2(n15241), 
        .C1(n15240), .C2(n15239), .ZN(P1_U3329) );
  MUX2_X1 U16948 ( .A(n15244), .B(n15243), .S(P1_U3086), .Z(P1_U3333) );
  INV_X1 U16949 ( .A(n15245), .ZN(n15246) );
  MUX2_X1 U16950 ( .A(n15246), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  AOI21_X1 U16951 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(
        P3_WR_REG_SCAN_IN), .ZN(n15249) );
  OAI21_X1 U16952 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(n15249), 
        .ZN(U28) );
  INV_X1 U16953 ( .A(P2_RD_REG_SCAN_IN), .ZN(n15251) );
  OAI221_X1 U16954 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .C1(
        n15251), .C2(n7140), .A(n15250), .ZN(U29) );
  OAI21_X1 U16955 ( .B1(n15253), .B2(n6693), .A(n15252), .ZN(n15254) );
  XNOR2_X1 U16956 ( .A(n15254), .B(P2_ADDR_REG_2__SCAN_IN), .ZN(SUB_1596_U61)
         );
  AOI21_X1 U16957 ( .B1(n15257), .B2(n15256), .A(n15255), .ZN(SUB_1596_U57) );
  AOI21_X1 U16958 ( .B1(n15260), .B2(n15259), .A(n15258), .ZN(SUB_1596_U55) );
  AOI21_X1 U16959 ( .B1(n15263), .B2(n15262), .A(n15261), .ZN(n15264) );
  XOR2_X1 U16960 ( .A(P2_ADDR_REG_9__SCAN_IN), .B(n15264), .Z(SUB_1596_U54) );
  OAI21_X1 U16961 ( .B1(n15267), .B2(n15266), .A(n15265), .ZN(n15268) );
  XNOR2_X1 U16962 ( .A(n15268), .B(P2_ADDR_REG_10__SCAN_IN), .ZN(SUB_1596_U70)
         );
  OAI211_X1 U16963 ( .C1(n15271), .C2(n15518), .A(n15270), .B(n15269), .ZN(
        n15272) );
  AOI21_X1 U16964 ( .B1(n15413), .B2(n15273), .A(n15272), .ZN(n15276) );
  INV_X1 U16965 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n15274) );
  AOI22_X1 U16966 ( .A1(n15526), .A2(n15276), .B1(n15274), .B2(n15524), .ZN(
        P1_U3495) );
  AOI22_X1 U16967 ( .A1(n15537), .A2(n15276), .B1(n15275), .B2(n15534), .ZN(
        P1_U3540) );
  NAND3_X1 U16968 ( .A1(n12325), .A2(n15288), .A3(n15278), .ZN(n15279) );
  NAND3_X1 U16969 ( .A1(n15277), .A2(n15280), .A3(n15279), .ZN(n15282) );
  AND2_X1 U16970 ( .A1(n15282), .A2(n15281), .ZN(n15404) );
  AOI222_X1 U16971 ( .A1(n15286), .A2(n15285), .B1(P1_REG2_REG_13__SCAN_IN), 
        .B2(n15067), .C1(n15284), .C2(n15283), .ZN(n15296) );
  XNOR2_X1 U16972 ( .A(n15287), .B(n15288), .ZN(n15406) );
  OAI211_X1 U16973 ( .C1(n12360), .C2(n12359), .A(n15291), .B(n15290), .ZN(
        n15403) );
  INV_X1 U16974 ( .A(n15403), .ZN(n15292) );
  AOI22_X1 U16975 ( .A1(n15406), .A2(n15294), .B1(n15293), .B2(n15292), .ZN(
        n15295) );
  OAI211_X1 U16976 ( .C1(n15067), .C2(n15404), .A(n15296), .B(n15295), .ZN(
        P1_U3280) );
  AOI21_X1 U16977 ( .B1(n15299), .B2(n15298), .A(n15297), .ZN(n15300) );
  XOR2_X1 U16978 ( .A(P2_ADDR_REG_17__SCAN_IN), .B(n15300), .Z(SUB_1596_U63)
         );
  INV_X1 U16979 ( .A(n15301), .ZN(n15302) );
  AOI22_X1 U16980 ( .A1(n15304), .A2(n15709), .B1(n15313), .B2(n15733), .ZN(
        n15308) );
  AOI22_X1 U16981 ( .A1(n15305), .A2(n15707), .B1(P3_REG2_REG_31__SCAN_IN), 
        .B2(n15735), .ZN(n15306) );
  NAND2_X1 U16982 ( .A1(n15308), .A2(n15306), .ZN(P3_U3202) );
  AOI22_X1 U16983 ( .A1(n15314), .A2(n15707), .B1(P3_REG2_REG_30__SCAN_IN), 
        .B2(n15735), .ZN(n15307) );
  NAND2_X1 U16984 ( .A1(n15308), .A2(n15307), .ZN(P3_U3203) );
  OR2_X1 U16985 ( .A1(n15309), .A2(n15758), .ZN(n15311) );
  INV_X1 U16986 ( .A(n15313), .ZN(n15310) );
  AOI22_X1 U16987 ( .A1(n15784), .A2(n15332), .B1(n15312), .B2(n15782), .ZN(
        P3_U3490) );
  AOI21_X1 U16988 ( .B1(n15314), .B2(n15765), .A(n15313), .ZN(n15334) );
  AOI22_X1 U16989 ( .A1(n15784), .A2(n15334), .B1(n15315), .B2(n15782), .ZN(
        P3_U3489) );
  AND2_X1 U16990 ( .A1(n15317), .A2(n15316), .ZN(n15320) );
  AND2_X1 U16991 ( .A1(n15318), .A2(n15765), .ZN(n15319) );
  NOR3_X1 U16992 ( .A1(n15321), .A2(n15320), .A3(n15319), .ZN(n15336) );
  AOI22_X1 U16993 ( .A1(n15784), .A2(n15336), .B1(n9234), .B2(n15782), .ZN(
        P3_U3472) );
  NOR2_X1 U16994 ( .A1(n15322), .A2(n15327), .ZN(n15324) );
  AOI211_X1 U16995 ( .C1(n15765), .C2(n15325), .A(n15324), .B(n15323), .ZN(
        n15338) );
  AOI22_X1 U16996 ( .A1(n15784), .A2(n15338), .B1(n9211), .B2(n15782), .ZN(
        P3_U3471) );
  OAI22_X1 U16997 ( .A1(n15328), .A2(n15327), .B1(n15326), .B2(n15758), .ZN(
        n15329) );
  NOR2_X1 U16998 ( .A1(n15330), .A2(n15329), .ZN(n15340) );
  AOI22_X1 U16999 ( .A1(n15784), .A2(n15340), .B1(n9194), .B2(n15782), .ZN(
        P3_U3470) );
  INV_X1 U17000 ( .A(P3_REG0_REG_31__SCAN_IN), .ZN(n15331) );
  AOI22_X1 U17001 ( .A1(n15775), .A2(n15332), .B1(n15331), .B2(n15773), .ZN(
        P3_U3458) );
  INV_X1 U17002 ( .A(P3_REG0_REG_30__SCAN_IN), .ZN(n15333) );
  AOI22_X1 U17003 ( .A1(n15775), .A2(n15334), .B1(n15333), .B2(n15773), .ZN(
        P3_U3457) );
  INV_X1 U17004 ( .A(P3_REG0_REG_13__SCAN_IN), .ZN(n15335) );
  AOI22_X1 U17005 ( .A1(n15775), .A2(n15336), .B1(n15335), .B2(n15773), .ZN(
        P3_U3429) );
  INV_X1 U17006 ( .A(P3_REG0_REG_12__SCAN_IN), .ZN(n15337) );
  AOI22_X1 U17007 ( .A1(n15775), .A2(n15338), .B1(n15337), .B2(n15773), .ZN(
        P3_U3426) );
  INV_X1 U17008 ( .A(P3_REG0_REG_11__SCAN_IN), .ZN(n15339) );
  AOI22_X1 U17009 ( .A1(n15775), .A2(n15340), .B1(n15339), .B2(n15773), .ZN(
        P3_U3423) );
  NAND2_X1 U17010 ( .A1(n15343), .A2(n15342), .ZN(n15344) );
  NAND2_X1 U17011 ( .A1(n15341), .A2(n15344), .ZN(n15346) );
  AOI222_X1 U17012 ( .A1(n15350), .A2(n15349), .B1(n15348), .B2(n15347), .C1(
        n15346), .C2(n15345), .ZN(n15352) );
  OAI211_X1 U17013 ( .C1(n15354), .C2(n15353), .A(n15352), .B(n15351), .ZN(
        P2_U3208) );
  AND2_X1 U17014 ( .A1(n15355), .A2(n15366), .ZN(n15360) );
  OAI21_X1 U17015 ( .B1(n15357), .B2(n15644), .A(n15356), .ZN(n15358) );
  NOR3_X1 U17016 ( .A1(n15360), .A2(n15359), .A3(n15358), .ZN(n15369) );
  AOI22_X1 U17017 ( .A1(n15688), .A2(n15369), .B1(n15361), .B2(n7435), .ZN(
        P2_U3512) );
  OAI21_X1 U17018 ( .B1(n15363), .B2(n15644), .A(n15362), .ZN(n15365) );
  AOI211_X1 U17019 ( .C1(n15367), .C2(n15366), .A(n15365), .B(n15364), .ZN(
        n15371) );
  AOI22_X1 U17020 ( .A1(n15688), .A2(n15371), .B1(n15551), .B2(n7435), .ZN(
        P2_U3511) );
  INV_X1 U17021 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n15368) );
  AOI22_X1 U17022 ( .A1(n15680), .A2(n15369), .B1(n15368), .B2(n15678), .ZN(
        P2_U3469) );
  INV_X1 U17023 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n15370) );
  AOI22_X1 U17024 ( .A1(n15680), .A2(n15371), .B1(n15370), .B2(n15678), .ZN(
        P2_U3466) );
  OAI22_X1 U17025 ( .A1(n15387), .A2(n15373), .B1(n15372), .B2(n15384), .ZN(
        n15379) );
  NAND2_X1 U17026 ( .A1(n15375), .A2(n15374), .ZN(n15376) );
  AOI21_X1 U17027 ( .B1(n15377), .B2(n15376), .A(n15392), .ZN(n15378) );
  AOI211_X1 U17028 ( .C1(n15380), .C2(n15397), .A(n15379), .B(n15378), .ZN(
        n15382) );
  OAI211_X1 U17029 ( .C1(n15402), .C2(n15383), .A(n15382), .B(n15381), .ZN(
        P1_U3215) );
  OAI22_X1 U17030 ( .A1(n15387), .A2(n15386), .B1(n15385), .B2(n15384), .ZN(
        n15396) );
  INV_X1 U17031 ( .A(n15388), .ZN(n15394) );
  OAI21_X1 U17032 ( .B1(n15391), .B2(n15390), .A(n15389), .ZN(n15393) );
  AOI21_X1 U17033 ( .B1(n15394), .B2(n15393), .A(n15392), .ZN(n15395) );
  AOI211_X1 U17034 ( .C1(n15398), .C2(n15397), .A(n15396), .B(n15395), .ZN(
        n15400) );
  OAI211_X1 U17035 ( .C1(n15402), .C2(n15401), .A(n15400), .B(n15399), .ZN(
        P1_U3236) );
  OAI211_X1 U17036 ( .C1(n12359), .C2(n15518), .A(n15404), .B(n15403), .ZN(
        n15405) );
  AOI21_X1 U17037 ( .B1(n15406), .B2(n15413), .A(n15405), .ZN(n15417) );
  AOI22_X1 U17038 ( .A1(n15537), .A2(n15417), .B1(n15407), .B2(n15534), .ZN(
        P1_U3541) );
  OAI21_X1 U17039 ( .B1(n15409), .B2(n15518), .A(n15408), .ZN(n15412) );
  INV_X1 U17040 ( .A(n15410), .ZN(n15411) );
  AOI211_X1 U17041 ( .C1(n15414), .C2(n15413), .A(n15412), .B(n15411), .ZN(
        n15419) );
  AOI22_X1 U17042 ( .A1(n15537), .A2(n15419), .B1(n15415), .B2(n15534), .ZN(
        P1_U3539) );
  INV_X1 U17043 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n15416) );
  AOI22_X1 U17044 ( .A1(n15526), .A2(n15417), .B1(n15416), .B2(n15524), .ZN(
        P1_U3498) );
  INV_X1 U17045 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n15418) );
  AOI22_X1 U17046 ( .A1(n15526), .A2(n15419), .B1(n15418), .B2(n15524), .ZN(
        P1_U3492) );
  OAI21_X1 U17047 ( .B1(n15422), .B2(n15421), .A(n15420), .ZN(n15423) );
  XNOR2_X1 U17048 ( .A(n15423), .B(P2_ADDR_REG_11__SCAN_IN), .ZN(SUB_1596_U69)
         );
  OAI222_X1 U17049 ( .A1(n15567), .A2(n15427), .B1(n15567), .B2(n15426), .C1(
        n15425), .C2(n15424), .ZN(SUB_1596_U68) );
  OAI21_X1 U17050 ( .B1(n15430), .B2(n15429), .A(n15428), .ZN(n15431) );
  XNOR2_X1 U17051 ( .A(n15431), .B(P2_ADDR_REG_13__SCAN_IN), .ZN(SUB_1596_U67)
         );
  OAI21_X1 U17052 ( .B1(n15434), .B2(n15433), .A(n15432), .ZN(n15435) );
  XNOR2_X1 U17053 ( .A(n15435), .B(P2_ADDR_REG_14__SCAN_IN), .ZN(SUB_1596_U66)
         );
  OAI21_X1 U17054 ( .B1(n15438), .B2(n15437), .A(n15436), .ZN(n15439) );
  XNOR2_X1 U17055 ( .A(n15439), .B(P2_ADDR_REG_15__SCAN_IN), .ZN(SUB_1596_U65)
         );
  OAI21_X1 U17056 ( .B1(n15442), .B2(n15441), .A(n15440), .ZN(n15443) );
  XNOR2_X1 U17057 ( .A(n15443), .B(P2_ADDR_REG_16__SCAN_IN), .ZN(SUB_1596_U64)
         );
  AND3_X1 U17058 ( .A1(n15446), .A2(n15445), .A3(n15444), .ZN(n15447) );
  NOR3_X1 U17059 ( .A1(n15468), .A2(n15448), .A3(n15447), .ZN(n15455) );
  AND3_X1 U17060 ( .A1(n15451), .A2(n15450), .A3(n15449), .ZN(n15452) );
  NOR3_X1 U17061 ( .A1(n15470), .A2(n15453), .A3(n15452), .ZN(n15454) );
  AOI211_X1 U17062 ( .C1(n15457), .C2(n15456), .A(n15455), .B(n15454), .ZN(
        n15459) );
  AND2_X1 U17063 ( .A1(n15459), .A2(n15458), .ZN(n15461) );
  OAI211_X1 U17064 ( .C1(n15476), .C2(n15462), .A(n15461), .B(n15460), .ZN(
        P1_U3247) );
  AOI21_X1 U17065 ( .B1(n15464), .B2(P1_REG2_REG_15__SCAN_IN), .A(n15463), 
        .ZN(n15469) );
  AOI21_X1 U17066 ( .B1(n15466), .B2(P1_REG1_REG_15__SCAN_IN), .A(n15465), 
        .ZN(n15467) );
  OAI222_X1 U17067 ( .A1(n15472), .A2(n15471), .B1(n15470), .B2(n15469), .C1(
        n15468), .C2(n15467), .ZN(n15473) );
  INV_X1 U17068 ( .A(n15473), .ZN(n15475) );
  OAI211_X1 U17069 ( .C1(n15477), .C2(n15476), .A(n15475), .B(n15474), .ZN(
        P1_U3258) );
  AND2_X1 U17070 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n15478), .ZN(P1_U3294) );
  AND2_X1 U17071 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n15478), .ZN(P1_U3295) );
  AND2_X1 U17072 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n15478), .ZN(P1_U3296) );
  AND2_X1 U17073 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n15478), .ZN(P1_U3297) );
  AND2_X1 U17074 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n15478), .ZN(P1_U3298) );
  AND2_X1 U17075 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n15478), .ZN(P1_U3299) );
  AND2_X1 U17076 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n15478), .ZN(P1_U3300) );
  AND2_X1 U17077 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n15478), .ZN(P1_U3301) );
  AND2_X1 U17078 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n15478), .ZN(P1_U3302) );
  AND2_X1 U17079 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n15478), .ZN(P1_U3303) );
  AND2_X1 U17080 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n15478), .ZN(P1_U3304) );
  AND2_X1 U17081 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n15478), .ZN(P1_U3305) );
  AND2_X1 U17082 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n15478), .ZN(P1_U3306) );
  AND2_X1 U17083 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n15478), .ZN(P1_U3307) );
  AND2_X1 U17084 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n15478), .ZN(P1_U3308) );
  AND2_X1 U17085 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n15478), .ZN(P1_U3309) );
  AND2_X1 U17086 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n15478), .ZN(P1_U3310) );
  AND2_X1 U17087 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n15478), .ZN(P1_U3311) );
  AND2_X1 U17088 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n15478), .ZN(P1_U3312) );
  AND2_X1 U17089 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n15478), .ZN(P1_U3313) );
  AND2_X1 U17090 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n15478), .ZN(P1_U3314) );
  AND2_X1 U17091 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n15478), .ZN(P1_U3315) );
  AND2_X1 U17092 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n15478), .ZN(P1_U3316) );
  AND2_X1 U17093 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n15478), .ZN(P1_U3317) );
  AND2_X1 U17094 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n15478), .ZN(P1_U3318) );
  AND2_X1 U17095 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n15478), .ZN(P1_U3319) );
  AND2_X1 U17096 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n15478), .ZN(P1_U3320) );
  AND2_X1 U17097 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n15478), .ZN(P1_U3321) );
  AND2_X1 U17098 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n15478), .ZN(P1_U3322) );
  AND2_X1 U17099 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n15478), .ZN(P1_U3323) );
  INV_X1 U17100 ( .A(n15479), .ZN(n15480) );
  AOI21_X1 U17101 ( .B1(n15482), .B2(n15481), .A(n15480), .ZN(n15483) );
  AOI211_X1 U17102 ( .C1(n15486), .C2(n15485), .A(n15484), .B(n15483), .ZN(
        n15527) );
  INV_X1 U17103 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n15487) );
  AOI22_X1 U17104 ( .A1(n15526), .A2(n15527), .B1(n15487), .B2(n15524), .ZN(
        P1_U3459) );
  OAI22_X1 U17105 ( .A1(n15489), .A2(n15488), .B1(n10686), .B2(n15518), .ZN(
        n15491) );
  AOI211_X1 U17106 ( .C1(n15523), .C2(n15492), .A(n15491), .B(n15490), .ZN(
        n15528) );
  INV_X1 U17107 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n15493) );
  AOI22_X1 U17108 ( .A1(n15526), .A2(n15528), .B1(n15493), .B2(n15524), .ZN(
        P1_U3462) );
  AOI21_X1 U17109 ( .B1(n15496), .B2(n15495), .A(n15494), .ZN(n15497) );
  OAI211_X1 U17110 ( .C1(n15500), .C2(n15499), .A(n15498), .B(n15497), .ZN(
        n15501) );
  INV_X1 U17111 ( .A(n15501), .ZN(n15529) );
  INV_X1 U17112 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n15502) );
  AOI22_X1 U17113 ( .A1(n15526), .A2(n15529), .B1(n15502), .B2(n15524), .ZN(
        P1_U3468) );
  AND2_X1 U17114 ( .A1(n15503), .A2(n15523), .ZN(n15507) );
  OAI21_X1 U17115 ( .B1(n15505), .B2(n15518), .A(n15504), .ZN(n15506) );
  NOR3_X1 U17116 ( .A1(n15508), .A2(n15507), .A3(n15506), .ZN(n15531) );
  INV_X1 U17117 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n15509) );
  AOI22_X1 U17118 ( .A1(n15526), .A2(n15531), .B1(n15509), .B2(n15524), .ZN(
        P1_U3474) );
  OAI21_X1 U17119 ( .B1(n15511), .B2(n15518), .A(n15510), .ZN(n15512) );
  AOI21_X1 U17120 ( .B1(n15513), .B2(n15523), .A(n15512), .ZN(n15514) );
  INV_X1 U17121 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n15516) );
  AOI22_X1 U17122 ( .A1(n15526), .A2(n15533), .B1(n15516), .B2(n15524), .ZN(
        P1_U3480) );
  OAI21_X1 U17123 ( .B1(n15519), .B2(n15518), .A(n15517), .ZN(n15521) );
  AOI211_X1 U17124 ( .C1(n15523), .C2(n15522), .A(n15521), .B(n15520), .ZN(
        n15536) );
  INV_X1 U17125 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n15525) );
  AOI22_X1 U17126 ( .A1(n15526), .A2(n15536), .B1(n15525), .B2(n15524), .ZN(
        P1_U3486) );
  AOI22_X1 U17127 ( .A1(n15537), .A2(n15527), .B1(n9873), .B2(n15534), .ZN(
        P1_U3528) );
  AOI22_X1 U17128 ( .A1(n15537), .A2(n15528), .B1(n10169), .B2(n15534), .ZN(
        P1_U3529) );
  AOI22_X1 U17129 ( .A1(n15537), .A2(n15529), .B1(n10176), .B2(n15534), .ZN(
        P1_U3531) );
  AOI22_X1 U17130 ( .A1(n15537), .A2(n15531), .B1(n15530), .B2(n15534), .ZN(
        P1_U3533) );
  AOI22_X1 U17131 ( .A1(n15537), .A2(n15533), .B1(n15532), .B2(n15534), .ZN(
        P1_U3535) );
  AOI22_X1 U17132 ( .A1(n15537), .A2(n15536), .B1(n15535), .B2(n15534), .ZN(
        P1_U3537) );
  NOR2_X1 U17133 ( .A1(n15601), .A2(n6672), .ZN(P2_U3087) );
  OAI21_X1 U17134 ( .B1(n15566), .B2(n7822), .A(n15538), .ZN(n15539) );
  AOI21_X1 U17135 ( .B1(n15540), .B2(n15603), .A(n15539), .ZN(n15549) );
  OAI211_X1 U17136 ( .C1(n15543), .C2(n15542), .A(n15609), .B(n15541), .ZN(
        n15548) );
  OAI211_X1 U17137 ( .C1(n15546), .C2(n15545), .A(n15604), .B(n15544), .ZN(
        n15547) );
  NAND3_X1 U17138 ( .A1(n15549), .A2(n15548), .A3(n15547), .ZN(P2_U3220) );
  INV_X1 U17139 ( .A(n15550), .ZN(n15554) );
  MUX2_X1 U17140 ( .A(P2_REG1_REG_12__SCAN_IN), .B(n15551), .S(n15555), .Z(
        n15553) );
  OAI21_X1 U17141 ( .B1(n15554), .B2(n15553), .A(n15552), .ZN(n15556) );
  AOI22_X1 U17142 ( .A1(n15556), .A2(n15609), .B1(n15555), .B2(n15603), .ZN(
        n15563) );
  AND3_X1 U17143 ( .A1(n15559), .A2(n15558), .A3(n15557), .ZN(n15560) );
  OAI21_X1 U17144 ( .B1(n15561), .B2(n15560), .A(n15604), .ZN(n15562) );
  AND2_X1 U17145 ( .A1(n15563), .A2(n15562), .ZN(n15565) );
  NAND2_X1 U17146 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(P2_U3088), .ZN(n15564)
         );
  OAI211_X1 U17147 ( .C1(n15567), .C2(n15566), .A(n15565), .B(n15564), .ZN(
        P2_U3226) );
  AOI22_X1 U17148 ( .A1(n15601), .A2(P2_ADDR_REG_13__SCAN_IN), .B1(
        P2_REG3_REG_13__SCAN_IN), .B2(P2_U3088), .ZN(n15578) );
  NAND2_X1 U17149 ( .A1(n15568), .A2(n15603), .ZN(n15577) );
  OAI211_X1 U17150 ( .C1(n15571), .C2(n15570), .A(n15604), .B(n15569), .ZN(
        n15576) );
  OAI211_X1 U17151 ( .C1(n15574), .C2(n15573), .A(n15609), .B(n15572), .ZN(
        n15575) );
  NAND4_X1 U17152 ( .A1(n15578), .A2(n15577), .A3(n15576), .A4(n15575), .ZN(
        P2_U3227) );
  INV_X1 U17153 ( .A(n15579), .ZN(n15581) );
  OAI21_X1 U17154 ( .B1(n15581), .B2(n15580), .A(P2_STATE_REG_SCAN_IN), .ZN(
        n15582) );
  OAI21_X1 U17155 ( .B1(P2_STATE_REG_SCAN_IN), .B2(P2_REG3_REG_14__SCAN_IN), 
        .A(n15582), .ZN(n15591) );
  OAI211_X1 U17156 ( .C1(n15584), .C2(P2_REG2_REG_14__SCAN_IN), .A(n15604), 
        .B(n15583), .ZN(n15590) );
  OAI211_X1 U17157 ( .C1(n15587), .C2(n15586), .A(n15609), .B(n15585), .ZN(
        n15589) );
  NAND2_X1 U17158 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(n15601), .ZN(n15588) );
  NAND4_X1 U17159 ( .A1(n15591), .A2(n15590), .A3(n15589), .A4(n15588), .ZN(
        P2_U3228) );
  AOI22_X1 U17160 ( .A1(n15601), .A2(P2_ADDR_REG_15__SCAN_IN), .B1(
        P2_REG3_REG_15__SCAN_IN), .B2(P2_U3088), .ZN(n15600) );
  NAND2_X1 U17161 ( .A1(n15603), .A2(n15592), .ZN(n15599) );
  OAI211_X1 U17162 ( .C1(n15594), .C2(P2_REG2_REG_15__SCAN_IN), .A(n15604), 
        .B(n15593), .ZN(n15598) );
  OAI211_X1 U17163 ( .C1(P2_REG1_REG_15__SCAN_IN), .C2(n15596), .A(n15609), 
        .B(n15595), .ZN(n15597) );
  NAND4_X1 U17164 ( .A1(n15600), .A2(n15599), .A3(n15598), .A4(n15597), .ZN(
        P2_U3229) );
  AOI22_X1 U17165 ( .A1(n15601), .A2(P2_ADDR_REG_16__SCAN_IN), .B1(
        P2_REG3_REG_16__SCAN_IN), .B2(P2_U3088), .ZN(n15615) );
  NAND2_X1 U17166 ( .A1(n15603), .A2(n15602), .ZN(n15614) );
  OAI211_X1 U17167 ( .C1(n15607), .C2(n15606), .A(n15605), .B(n15604), .ZN(
        n15613) );
  OAI211_X1 U17168 ( .C1(n15611), .C2(n15610), .A(n15609), .B(n15608), .ZN(
        n15612) );
  NAND4_X1 U17169 ( .A1(n15615), .A2(n15614), .A3(n15613), .A4(n15612), .ZN(
        P2_U3230) );
  NOR2_X1 U17170 ( .A1(n15616), .A2(n8860), .ZN(n15638) );
  NOR2_X1 U17171 ( .A1(n15663), .A2(n15617), .ZN(n15619) );
  OAI21_X1 U17172 ( .B1(n15636), .B2(n15619), .A(n15618), .ZN(n15637) );
  AOI21_X1 U17173 ( .B1(n15638), .B2(n15620), .A(n15637), .ZN(n15626) );
  INV_X1 U17174 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n15622) );
  OAI22_X1 U17175 ( .A1(n15623), .A2(n15636), .B1(n15622), .B2(n15621), .ZN(
        n15624) );
  INV_X1 U17176 ( .A(n15624), .ZN(n15625) );
  OAI221_X1 U17177 ( .B1(n15627), .B2(n15626), .C1(n14226), .C2(n10328), .A(
        n15625), .ZN(P2_U3265) );
  AND2_X1 U17178 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n15630), .ZN(P2_U3266) );
  AND2_X1 U17179 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n15630), .ZN(P2_U3267) );
  AND2_X1 U17180 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n15630), .ZN(P2_U3268) );
  AND2_X1 U17181 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n15630), .ZN(P2_U3269) );
  AND2_X1 U17182 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n15630), .ZN(P2_U3270) );
  AND2_X1 U17183 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n15630), .ZN(P2_U3271) );
  AND2_X1 U17184 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n15630), .ZN(P2_U3272) );
  AND2_X1 U17185 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n15630), .ZN(P2_U3273) );
  AND2_X1 U17186 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n15630), .ZN(P2_U3274) );
  AND2_X1 U17187 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n15630), .ZN(P2_U3275) );
  AND2_X1 U17188 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n15630), .ZN(P2_U3276) );
  AND2_X1 U17189 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n15630), .ZN(P2_U3277) );
  AND2_X1 U17190 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n15630), .ZN(P2_U3278) );
  AND2_X1 U17191 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n15630), .ZN(P2_U3279) );
  AND2_X1 U17192 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n15630), .ZN(P2_U3280) );
  AND2_X1 U17193 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n15630), .ZN(P2_U3281) );
  AND2_X1 U17194 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n15630), .ZN(P2_U3282) );
  AND2_X1 U17195 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n15630), .ZN(P2_U3283) );
  AND2_X1 U17196 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n15630), .ZN(P2_U3284) );
  AND2_X1 U17197 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n15630), .ZN(P2_U3285) );
  AND2_X1 U17198 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n15630), .ZN(P2_U3286) );
  AND2_X1 U17199 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n15630), .ZN(P2_U3287) );
  AND2_X1 U17200 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n15630), .ZN(P2_U3288) );
  AND2_X1 U17201 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n15630), .ZN(P2_U3289) );
  AND2_X1 U17202 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n15630), .ZN(P2_U3290) );
  AND2_X1 U17203 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n15630), .ZN(P2_U3291) );
  AND2_X1 U17204 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n15630), .ZN(P2_U3292) );
  AND2_X1 U17205 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n15630), .ZN(P2_U3293) );
  AND2_X1 U17206 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n15630), .ZN(P2_U3294) );
  AND2_X1 U17207 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n15630), .ZN(P2_U3295) );
  AOI22_X1 U17208 ( .A1(n15635), .A2(n15632), .B1(n15631), .B2(n15630), .ZN(
        P2_U3416) );
  OAI21_X1 U17209 ( .B1(n15635), .B2(n15634), .A(n15633), .ZN(P2_U3417) );
  INV_X1 U17210 ( .A(n15636), .ZN(n15639) );
  AOI211_X1 U17211 ( .C1(n15662), .C2(n15639), .A(n15638), .B(n15637), .ZN(
        n15682) );
  INV_X1 U17212 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n15640) );
  AOI22_X1 U17213 ( .A1(n15680), .A2(n15682), .B1(n15640), .B2(n15678), .ZN(
        P2_U3430) );
  INV_X1 U17214 ( .A(n15641), .ZN(n15642) );
  AOI21_X1 U17215 ( .B1(n15675), .B2(n8992), .A(n15642), .ZN(n15647) );
  OAI21_X1 U17216 ( .B1(n8887), .B2(n15644), .A(n15643), .ZN(n15645) );
  NOR3_X1 U17217 ( .A1(n15647), .A2(n15646), .A3(n15645), .ZN(n15684) );
  INV_X1 U17218 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n15648) );
  AOI22_X1 U17219 ( .A1(n15680), .A2(n15684), .B1(n15648), .B2(n15678), .ZN(
        P2_U3433) );
  INV_X1 U17220 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n15649) );
  AOI22_X1 U17221 ( .A1(n15680), .A2(n15650), .B1(n15649), .B2(n15678), .ZN(
        P2_U3436) );
  AOI21_X1 U17222 ( .B1(n15672), .B2(n15652), .A(n15651), .ZN(n15654) );
  OAI211_X1 U17223 ( .C1(n15656), .C2(n15655), .A(n15654), .B(n15653), .ZN(
        n15657) );
  INV_X1 U17224 ( .A(n15657), .ZN(n15685) );
  INV_X1 U17225 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n15658) );
  AOI22_X1 U17226 ( .A1(n15680), .A2(n15685), .B1(n15658), .B2(n15678), .ZN(
        P2_U3439) );
  NAND2_X1 U17227 ( .A1(n15659), .A2(n15672), .ZN(n15660) );
  AND2_X1 U17228 ( .A1(n15661), .A2(n15660), .ZN(n15667) );
  NAND2_X1 U17229 ( .A1(n15664), .A2(n15662), .ZN(n15666) );
  NAND2_X1 U17230 ( .A1(n15664), .A2(n15663), .ZN(n15665) );
  INV_X1 U17231 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n15669) );
  AOI22_X1 U17232 ( .A1(n15680), .A2(n15686), .B1(n15669), .B2(n15678), .ZN(
        P2_U3442) );
  AOI21_X1 U17233 ( .B1(n15672), .B2(n15671), .A(n15670), .ZN(n15673) );
  OAI211_X1 U17234 ( .C1(n15676), .C2(n15675), .A(n15674), .B(n15673), .ZN(
        n15677) );
  INV_X1 U17235 ( .A(n15677), .ZN(n15687) );
  INV_X1 U17236 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n15679) );
  AOI22_X1 U17237 ( .A1(n15680), .A2(n15687), .B1(n15679), .B2(n15678), .ZN(
        P2_U3448) );
  AOI22_X1 U17238 ( .A1(n15688), .A2(n15682), .B1(n15681), .B2(n7435), .ZN(
        P2_U3499) );
  AOI22_X1 U17239 ( .A1(n15688), .A2(n15684), .B1(n15683), .B2(n7435), .ZN(
        P2_U3500) );
  AOI22_X1 U17240 ( .A1(n15688), .A2(n15685), .B1(n10110), .B2(n7435), .ZN(
        P2_U3502) );
  AOI22_X1 U17241 ( .A1(n15688), .A2(n15686), .B1(n10114), .B2(n7435), .ZN(
        P2_U3503) );
  AOI22_X1 U17242 ( .A1(n15688), .A2(n15687), .B1(n10118), .B2(n7435), .ZN(
        P2_U3505) );
  NOR2_X1 U17243 ( .A1(P3_U3897), .A2(n15698), .ZN(P3_U3150) );
  MUX2_X1 U17244 ( .A(n15690), .B(n15689), .S(n6945), .Z(n15691) );
  NOR2_X1 U17245 ( .A1(n15691), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n15696) );
  NAND3_X1 U17246 ( .A1(n15694), .A2(n15693), .A3(n15692), .ZN(n15695) );
  OAI21_X1 U17247 ( .B1(n15697), .B2(n15696), .A(n15695), .ZN(n15701) );
  AOI22_X1 U17248 ( .A1(n15699), .A2(P3_IR_REG_0__SCAN_IN), .B1(n15698), .B2(
        P3_ADDR_REG_0__SCAN_IN), .ZN(n15700) );
  OAI211_X1 U17249 ( .C1(P3_STATE_REG_SCAN_IN), .C2(n15702), .A(n15701), .B(
        n15700), .ZN(P3_U3182) );
  NAND2_X1 U17250 ( .A1(n15704), .A2(n15703), .ZN(n15705) );
  NAND2_X1 U17251 ( .A1(n15706), .A2(n15705), .ZN(n15711) );
  AOI222_X1 U17252 ( .A1(n15733), .A2(n15711), .B1(n15710), .B2(n15709), .C1(
        n15708), .C2(n15707), .ZN(n15712) );
  OAI21_X1 U17253 ( .B1(n15733), .B2(n15713), .A(n15712), .ZN(P3_U3227) );
  NOR2_X1 U17254 ( .A1(n15714), .A2(n15758), .ZN(n15738) );
  INV_X1 U17255 ( .A(n15715), .ZN(n15726) );
  XNOR2_X1 U17256 ( .A(n6935), .B(n15721), .ZN(n15736) );
  AOI22_X1 U17257 ( .A1(n15719), .A2(n15718), .B1(n9512), .B2(n15717), .ZN(
        n15725) );
  XNOR2_X1 U17258 ( .A(n15721), .B(n15720), .ZN(n15723) );
  NAND2_X1 U17259 ( .A1(n15723), .A2(n15722), .ZN(n15724) );
  OAI211_X1 U17260 ( .C1(n15736), .C2(n15764), .A(n15725), .B(n15724), .ZN(
        n15737) );
  AOI21_X1 U17261 ( .B1(n15738), .B2(n15726), .A(n15737), .ZN(n15734) );
  OAI22_X1 U17262 ( .A1(n15736), .A2(n15729), .B1(n15728), .B2(n15727), .ZN(
        n15730) );
  INV_X1 U17263 ( .A(n15730), .ZN(n15731) );
  OAI221_X1 U17264 ( .B1(n15735), .B2(n15734), .C1(n15733), .C2(n15732), .A(
        n15731), .ZN(P3_U3232) );
  INV_X1 U17265 ( .A(n15736), .ZN(n15739) );
  AOI211_X1 U17266 ( .C1(n15745), .C2(n15739), .A(n15738), .B(n15737), .ZN(
        n15776) );
  INV_X1 U17267 ( .A(P3_REG0_REG_1__SCAN_IN), .ZN(n15740) );
  AOI22_X1 U17268 ( .A1(n15775), .A2(n15776), .B1(n15740), .B2(n15773), .ZN(
        P3_U3393) );
  INV_X1 U17269 ( .A(n15741), .ZN(n15743) );
  AOI211_X1 U17270 ( .C1(n15745), .C2(n15744), .A(n15743), .B(n15742), .ZN(
        n15777) );
  INV_X1 U17271 ( .A(P3_REG0_REG_2__SCAN_IN), .ZN(n15746) );
  AOI22_X1 U17272 ( .A1(n15775), .A2(n15777), .B1(n15746), .B2(n15773), .ZN(
        P3_U3396) );
  OAI22_X1 U17273 ( .A1(n15748), .A2(n15769), .B1(n15747), .B2(n15758), .ZN(
        n15749) );
  NOR2_X1 U17274 ( .A1(n15750), .A2(n15749), .ZN(n15778) );
  INV_X1 U17275 ( .A(P3_REG0_REG_3__SCAN_IN), .ZN(n15751) );
  AOI22_X1 U17276 ( .A1(n15775), .A2(n15778), .B1(n15751), .B2(n15773), .ZN(
        P3_U3399) );
  INV_X1 U17277 ( .A(n15752), .ZN(n15754) );
  OAI22_X1 U17278 ( .A1(n15754), .A2(n15769), .B1(n15753), .B2(n15758), .ZN(
        n15755) );
  NOR2_X1 U17279 ( .A1(n15756), .A2(n15755), .ZN(n15779) );
  INV_X1 U17280 ( .A(P3_REG0_REG_5__SCAN_IN), .ZN(n15757) );
  AOI22_X1 U17281 ( .A1(n15775), .A2(n15779), .B1(n15757), .B2(n15773), .ZN(
        P3_U3405) );
  OAI22_X1 U17282 ( .A1(n15760), .A2(n15769), .B1(n15759), .B2(n15758), .ZN(
        n15761) );
  NOR2_X1 U17283 ( .A1(n15762), .A2(n15761), .ZN(n15781) );
  INV_X1 U17284 ( .A(P3_REG0_REG_9__SCAN_IN), .ZN(n15763) );
  AOI22_X1 U17285 ( .A1(n15775), .A2(n15781), .B1(n15763), .B2(n15773), .ZN(
        P3_U3417) );
  OR2_X1 U17286 ( .A1(n15770), .A2(n15764), .ZN(n15768) );
  NAND2_X1 U17287 ( .A1(n15766), .A2(n15765), .ZN(n15767) );
  OAI211_X1 U17288 ( .C1(n15770), .C2(n15769), .A(n15768), .B(n15767), .ZN(
        n15771) );
  NOR2_X1 U17289 ( .A1(n15772), .A2(n15771), .ZN(n15783) );
  INV_X1 U17290 ( .A(P3_REG0_REG_10__SCAN_IN), .ZN(n15774) );
  AOI22_X1 U17291 ( .A1(n15775), .A2(n15783), .B1(n15774), .B2(n15773), .ZN(
        P3_U3420) );
  AOI22_X1 U17292 ( .A1(n15784), .A2(n15776), .B1(n9019), .B2(n15782), .ZN(
        P3_U3460) );
  AOI22_X1 U17293 ( .A1(n15784), .A2(n15777), .B1(n10766), .B2(n15782), .ZN(
        P3_U3461) );
  AOI22_X1 U17294 ( .A1(n15784), .A2(n15778), .B1(n10735), .B2(n15782), .ZN(
        P3_U3462) );
  AOI22_X1 U17295 ( .A1(n15784), .A2(n15779), .B1(n9092), .B2(n15782), .ZN(
        P3_U3464) );
  AOI22_X1 U17296 ( .A1(n15784), .A2(n15781), .B1(n15780), .B2(n15782), .ZN(
        P3_U3468) );
  AOI22_X1 U17297 ( .A1(n15784), .A2(n15783), .B1(n11451), .B2(n15782), .ZN(
        P3_U3469) );
  AOI21_X1 U17298 ( .B1(n15787), .B2(n15786), .A(n15785), .ZN(SUB_1596_U59) );
  OAI21_X1 U17299 ( .B1(n15790), .B2(n15789), .A(n15788), .ZN(SUB_1596_U58) );
  XOR2_X1 U17300 ( .A(P2_ADDR_REG_0__SCAN_IN), .B(n15791), .Z(SUB_1596_U53) );
  OAI21_X1 U17301 ( .B1(n15794), .B2(n15793), .A(n15792), .ZN(SUB_1596_U56) );
  AOI21_X1 U17302 ( .B1(n15797), .B2(n15796), .A(n15795), .ZN(n15798) );
  XOR2_X1 U17303 ( .A(P2_ADDR_REG_3__SCAN_IN), .B(n15798), .Z(SUB_1596_U60) );
  AOI21_X1 U17304 ( .B1(n15801), .B2(n15800), .A(n15799), .ZN(SUB_1596_U5) );
  XNOR2_X1 U11502 ( .A(n9017), .B(P3_IR_REG_29__SCAN_IN), .ZN(n9020) );
  BUF_X2 U7417 ( .A(n9865), .Z(n12519) );
  CLKBUF_X1 U7427 ( .A(n14555), .Z(n6950) );
  CLKBUF_X1 U7431 ( .A(n9893), .Z(n14515) );
  CLKBUF_X2 U7432 ( .A(n9733), .Z(n10748) );
  AND4_X1 U7493 ( .A1(n9096), .A2(n9095), .A3(n9094), .A4(n9093), .ZN(n11792)
         );
  OR2_X1 U7524 ( .A1(n8379), .A2(n9982), .ZN(n8347) );
  CLKBUF_X2 U7723 ( .A(n12609), .Z(n6669) );
endmodule

