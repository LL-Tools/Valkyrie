

module b21_C_SARLock_k_64_7 ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, 
        P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, 
        P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, 
        P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, 
        P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, 
        P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, 
        P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, 
        P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, 
        P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, 
        P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, 
        P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, 
        P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, 
        P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, 
        P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, 
        P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, 
        P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, 
        P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, 
        P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, 
        P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, 
        P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, 
        P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, 
        P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, 
        P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, 
        P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, 
        P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3, 
        keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9, 
        keyinput10, keyinput11, keyinput12, keyinput13, keyinput14, keyinput15, 
        keyinput16, keyinput17, keyinput18, keyinput19, keyinput20, keyinput21, 
        keyinput22, keyinput23, keyinput24, keyinput25, keyinput26, keyinput27, 
        keyinput28, keyinput29, keyinput30, keyinput31, keyinput32, keyinput33, 
        keyinput34, keyinput35, keyinput36, keyinput37, keyinput38, keyinput39, 
        keyinput40, keyinput41, keyinput42, keyinput43, keyinput44, keyinput45, 
        keyinput46, keyinput47, keyinput48, keyinput49, keyinput50, keyinput51, 
        keyinput52, keyinput53, keyinput54, keyinput55, keyinput56, keyinput57, 
        keyinput58, keyinput59, keyinput60, keyinput61, keyinput62, keyinput63, 
        ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, ADD_1071_U57, ADD_1071_U58, 
        ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, ADD_1071_U62, ADD_1071_U63, 
        ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, ADD_1071_U50, ADD_1071_U51, 
        ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, ADD_1071_U5, ADD_1071_U46, 
        U126, U123, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349, P1_U3348, 
        P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342, P1_U3341, 
        P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335, P1_U3334, 
        P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328, P1_U3327, 
        P1_U3326, P1_U3325, P1_U3324, P1_U3323, P1_U3322, P1_U3440, P1_U3441, 
        P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316, P1_U3315, 
        P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309, P1_U3308, 
        P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302, P1_U3301, 
        P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295, P1_U3294, 
        P1_U3293, P1_U3292, P1_U3454, P1_U3457, P1_U3460, P1_U3463, P1_U3466, 
        P1_U3469, P1_U3472, P1_U3475, P1_U3478, P1_U3481, P1_U3484, P1_U3487, 
        P1_U3490, P1_U3493, P1_U3496, P1_U3499, P1_U3502, P1_U3505, P1_U3508, 
        P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515, P1_U3516, 
        P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, P1_U3523, 
        P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, P1_U3530, 
        P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, P1_U3537, 
        P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, P1_U3544, 
        P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, P1_U3551, 
        P1_U3552, P1_U3553, P1_U3554, P1_U3291, P1_U3290, P1_U3289, P1_U3288, 
        P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282, P1_U3281, 
        P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275, P1_U3274, 
        P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268, P1_U3267, 
        P1_U3266, P1_U3265, P1_U3264, P1_U3263, P1_U3355, P1_U3262, P1_U3261, 
        P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255, P1_U3254, 
        P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248, P1_U3247, 
        P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3242, P1_U3241, P1_U3555, 
        P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561, P1_U3562, 
        P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, P1_U3569, 
        P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, P1_U3576, 
        P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, P1_U3583, 
        P1_U3584, P1_U3585, P1_U3586, P1_U3240, P1_U3239, P1_U3238, P1_U3237, 
        P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231, P1_U3230, 
        P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224, P1_U3223, 
        P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, P1_U3216, 
        P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, P1_U3084, P1_U3083, 
        P1_U4006, P2_U3358, P2_U3357, P2_U3356, P2_U3355, P2_U3354, P2_U3353, 
        P2_U3352, P2_U3351, P2_U3350, P2_U3349, P2_U3348, P2_U3347, P2_U3346, 
        P2_U3345, P2_U3344, P2_U3343, P2_U3342, P2_U3341, P2_U3340, P2_U3339, 
        P2_U3338, P2_U3337, P2_U3336, P2_U3335, P2_U3334, P2_U3333, P2_U3332, 
        P2_U3331, P2_U3330, P2_U3329, P2_U3328, P2_U3327, P2_U3437, P2_U3438, 
        P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321, P2_U3320, 
        P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314, P2_U3313, 
        P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307, P2_U3306, 
        P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300, P2_U3299, 
        P2_U3298, P2_U3297, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463, 
        P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484, 
        P2_U3487, P2_U3490, P2_U3493, P2_U3496, P2_U3499, P2_U3502, P2_U3505, 
        P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, 
        P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, 
        P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527, 
        P2_U3528, P2_U3529, P2_U3530, P2_U3531, P2_U3532, P2_U3533, P2_U3534, 
        P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540, P2_U3541, 
        P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547, P2_U3548, 
        P2_U3549, P2_U3550, P2_U3551, P2_U3296, P2_U3295, P2_U3294, P2_U3293, 
        P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, 
        P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, 
        P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, 
        P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, 
        P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258, 
        P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251, 
        P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3552, 
        P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559, 
        P2_U3560, P2_U3561, P2_U3562, P2_U3563, P2_U3564, P2_U3565, P2_U3566, 
        P2_U3567, P2_U3568, P2_U3569, P2_U3570, P2_U3571, P2_U3572, P2_U3573, 
        P2_U3574, P2_U3575, P2_U3576, P2_U3577, P2_U3578, P2_U3579, P2_U3580, 
        P2_U3581, P2_U3582, P2_U3583, P2_U3244, P2_U3243, P2_U3242, P2_U3241, 
        P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, 
        P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, 
        P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, 
        P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3152, P2_U3151, 
        P2_U3966 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN,
         P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN,
         P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN,
         P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN,
         P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN,
         P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN,
         P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN,
         P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN,
         P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN,
         P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN,
         P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN,
         P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN,
         P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN,
         P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN,
         P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN,
         P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN,
         P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN,
         P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN,
         P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN,
         P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN,
         P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN,
         P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63;
  output ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, ADD_1071_U57, ADD_1071_U58,
         ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, ADD_1071_U62, ADD_1071_U63,
         ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, ADD_1071_U50, ADD_1071_U51,
         ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, ADD_1071_U5, ADD_1071_U46,
         U126, U123, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349,
         P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342,
         P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335,
         P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328,
         P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, P1_U3322, P1_U3440,
         P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316,
         P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309,
         P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302,
         P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295,
         P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, P1_U3460, P1_U3463,
         P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, P1_U3481, P1_U3484,
         P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, P1_U3502, P1_U3505,
         P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515,
         P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522,
         P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529,
         P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536,
         P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543,
         P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550,
         P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, P1_U3290, P1_U3289,
         P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282,
         P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275,
         P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268,
         P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, P1_U3355, P1_U3262,
         P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255,
         P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248,
         P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3242, P1_U3241,
         P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561,
         P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568,
         P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575,
         P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582,
         P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, P1_U3239, P1_U3238,
         P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231,
         P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224,
         P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217,
         P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, P1_U3084,
         P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, P2_U3355, P2_U3354,
         P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, P2_U3348, P2_U3347,
         P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, P2_U3341, P2_U3340,
         P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, P2_U3334, P2_U3333,
         P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, P2_U3327, P2_U3437,
         P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321,
         P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314,
         P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307,
         P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300,
         P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, P2_U3457, P2_U3460,
         P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481,
         P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, P2_U3499, P2_U3502,
         P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512,
         P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519,
         P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526,
         P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, P2_U3532, P2_U3533,
         P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540,
         P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547,
         P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, P2_U3295, P2_U3294,
         P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287,
         P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280,
         P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273,
         P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266,
         P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259,
         P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252,
         P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245,
         P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558,
         P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, P2_U3564, P2_U3565,
         P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, P2_U3571, P2_U3572,
         P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, P2_U3578, P2_U3579,
         P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, P2_U3243, P2_U3242,
         P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235,
         P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228,
         P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221,
         P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3152,
         P2_U3151, P2_U3966;
  wire   n10047, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283,
         n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293,
         n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303,
         n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313,
         n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323,
         n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333,
         n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343,
         n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353,
         n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363,
         n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373,
         n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383,
         n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393,
         n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403,
         n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413,
         n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423,
         n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433,
         n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443,
         n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453,
         n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463,
         n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473,
         n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483,
         n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493,
         n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503,
         n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513,
         n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523,
         n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533,
         n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543,
         n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553,
         n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563,
         n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573,
         n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583,
         n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593,
         n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603,
         n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613,
         n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623,
         n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633,
         n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643,
         n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653,
         n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663,
         n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673,
         n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683,
         n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693,
         n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703,
         n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713,
         n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723,
         n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733,
         n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743,
         n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753,
         n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763,
         n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773,
         n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783,
         n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793,
         n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803,
         n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813,
         n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823,
         n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833,
         n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843,
         n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853,
         n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863,
         n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873,
         n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883,
         n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893,
         n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903,
         n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913,
         n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923,
         n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933,
         n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943,
         n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953,
         n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963,
         n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973,
         n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983,
         n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993,
         n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003,
         n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013,
         n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023,
         n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033,
         n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043,
         n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053,
         n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063,
         n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073,
         n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083,
         n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093,
         n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103,
         n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113,
         n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123,
         n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133,
         n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143,
         n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153,
         n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163,
         n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173,
         n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183,
         n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193,
         n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203,
         n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213,
         n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223,
         n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233,
         n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243,
         n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253,
         n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263,
         n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273,
         n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283,
         n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293,
         n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303,
         n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313,
         n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323,
         n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333,
         n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343,
         n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353,
         n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363,
         n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373,
         n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383,
         n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393,
         n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403,
         n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413,
         n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423,
         n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433,
         n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443,
         n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453,
         n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463,
         n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473,
         n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483,
         n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493,
         n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503,
         n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513,
         n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523,
         n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533,
         n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543,
         n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553,
         n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563,
         n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573,
         n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583,
         n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593,
         n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603,
         n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613,
         n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623,
         n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633,
         n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643,
         n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653,
         n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663,
         n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673,
         n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683,
         n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693,
         n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703,
         n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713,
         n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723,
         n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733,
         n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743,
         n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753,
         n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763,
         n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773,
         n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783,
         n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793,
         n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803,
         n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813,
         n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823,
         n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833,
         n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843,
         n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853,
         n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863,
         n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873,
         n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883,
         n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893,
         n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903,
         n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913,
         n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923,
         n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933,
         n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943,
         n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953,
         n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963,
         n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973,
         n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983,
         n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993,
         n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003,
         n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013,
         n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023,
         n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033,
         n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043,
         n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053,
         n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063,
         n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073,
         n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083,
         n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093,
         n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103,
         n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113,
         n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123,
         n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133,
         n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143,
         n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153,
         n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163,
         n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173,
         n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183,
         n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193,
         n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203,
         n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213,
         n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223,
         n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233,
         n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243,
         n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253,
         n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263,
         n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273,
         n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283,
         n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293,
         n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303,
         n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313,
         n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323,
         n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333,
         n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343,
         n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353,
         n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363,
         n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373,
         n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383,
         n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393,
         n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403,
         n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413,
         n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423,
         n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433,
         n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443,
         n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453,
         n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463,
         n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473,
         n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483,
         n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493,
         n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503,
         n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513,
         n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523,
         n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533,
         n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543,
         n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553,
         n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563,
         n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573,
         n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583,
         n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593,
         n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603,
         n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613,
         n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623,
         n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633,
         n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643,
         n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653,
         n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663,
         n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673,
         n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683,
         n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693,
         n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703,
         n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713,
         n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723,
         n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733,
         n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743,
         n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753,
         n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763,
         n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773,
         n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783,
         n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793,
         n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803,
         n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813,
         n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823,
         n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833,
         n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843,
         n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853,
         n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863,
         n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873,
         n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883,
         n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893,
         n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903,
         n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913,
         n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923,
         n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933,
         n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943,
         n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953,
         n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963,
         n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973,
         n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983,
         n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993,
         n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003,
         n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013,
         n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023,
         n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033,
         n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043,
         n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053,
         n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063,
         n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073,
         n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083,
         n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093,
         n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103,
         n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113,
         n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123,
         n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133,
         n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143,
         n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153,
         n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163,
         n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173,
         n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183,
         n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193,
         n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203,
         n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213,
         n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223,
         n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233,
         n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243,
         n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253,
         n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263,
         n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273,
         n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283,
         n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293,
         n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303,
         n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313,
         n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323,
         n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333,
         n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343,
         n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353,
         n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363,
         n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373,
         n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383,
         n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393,
         n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403,
         n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413,
         n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423,
         n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433,
         n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443,
         n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453,
         n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463,
         n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473,
         n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483,
         n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493,
         n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503,
         n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513,
         n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523,
         n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533,
         n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543,
         n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553,
         n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563,
         n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573,
         n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583,
         n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593,
         n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603,
         n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613,
         n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623,
         n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633,
         n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643,
         n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653,
         n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663,
         n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673,
         n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683,
         n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693,
         n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703,
         n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713,
         n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723,
         n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733,
         n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743,
         n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753,
         n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763,
         n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773,
         n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783,
         n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793,
         n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803,
         n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813,
         n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823,
         n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833,
         n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843,
         n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853,
         n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863,
         n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873,
         n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883,
         n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893,
         n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903,
         n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913,
         n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923,
         n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933,
         n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943,
         n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7953, n7954,
         n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964,
         n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974,
         n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984,
         n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994,
         n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004,
         n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014,
         n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024,
         n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034,
         n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044,
         n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054,
         n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064,
         n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074,
         n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084,
         n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094,
         n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104,
         n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114,
         n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124,
         n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134,
         n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144,
         n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154,
         n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164,
         n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174,
         n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184,
         n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194,
         n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204,
         n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214,
         n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224,
         n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234,
         n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244,
         n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254,
         n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264,
         n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274,
         n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284,
         n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294,
         n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304,
         n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314,
         n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324,
         n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334,
         n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344,
         n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354,
         n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364,
         n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374,
         n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384,
         n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394,
         n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404,
         n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414,
         n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424,
         n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434,
         n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444,
         n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454,
         n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464,
         n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474,
         n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484,
         n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494,
         n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504,
         n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514,
         n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524,
         n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534,
         n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544,
         n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554,
         n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564,
         n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574,
         n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584,
         n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594,
         n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604,
         n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614,
         n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624,
         n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634,
         n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644,
         n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654,
         n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664,
         n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674,
         n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684,
         n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694,
         n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704,
         n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714,
         n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724,
         n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734,
         n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744,
         n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754,
         n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764,
         n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774,
         n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784,
         n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794,
         n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804,
         n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814,
         n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824,
         n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834,
         n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844,
         n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854,
         n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864,
         n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874,
         n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884,
         n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894,
         n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904,
         n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914,
         n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924,
         n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934,
         n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944,
         n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954,
         n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964,
         n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974,
         n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984,
         n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994,
         n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004,
         n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014,
         n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024,
         n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034,
         n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044,
         n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054,
         n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064,
         n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074,
         n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084,
         n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094,
         n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104,
         n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114,
         n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124,
         n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134,
         n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144,
         n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154,
         n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164,
         n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174,
         n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184,
         n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194,
         n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204,
         n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214,
         n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224,
         n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234,
         n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244,
         n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254,
         n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264,
         n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274,
         n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284,
         n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294,
         n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304,
         n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314,
         n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324,
         n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334,
         n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344,
         n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354,
         n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364,
         n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374,
         n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384,
         n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394,
         n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404,
         n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414,
         n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424,
         n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434,
         n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444,
         n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454,
         n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464,
         n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474,
         n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484,
         n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494,
         n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504,
         n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514,
         n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524,
         n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534,
         n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544,
         n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554,
         n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564,
         n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574,
         n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584,
         n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594,
         n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604,
         n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614,
         n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624,
         n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634,
         n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644,
         n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654,
         n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664,
         n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674,
         n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684,
         n9685, n9686, n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695,
         n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705,
         n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715,
         n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725,
         n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735,
         n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745,
         n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755,
         n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765,
         n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775,
         n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785,
         n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795,
         n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805,
         n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815,
         n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825,
         n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835,
         n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845,
         n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855,
         n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865,
         n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875,
         n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885,
         n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895,
         n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905,
         n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915,
         n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925,
         n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935,
         n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945,
         n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955,
         n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965,
         n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975,
         n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985,
         n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995,
         n9996, n9997, n9998, n9999, n10000, n10001, n10002, n10003, n10004,
         n10005, n10006, n10007, n10008, n10009, n10010, n10011, n10012,
         n10013, n10014, n10015, n10016, n10017, n10018, n10019, n10020,
         n10021, n10022, n10023, n10024, n10025, n10026, n10027, n10028,
         n10029, n10030, n10031, n10032, n10033, n10034, n10035, n10036,
         n10037, n10038, n10039, n10040, n10041, n10042, n10043, n10044;

  INV_X4 U4779 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3152) );
  NAND2_X1 U4780 ( .A1(n8293), .A2(n8295), .ZN(n8684) );
  NAND2_X1 U4781 ( .A1(n5866), .A2(n5865), .ZN(n7062) );
  AND2_X1 U4782 ( .A1(n8194), .A2(n8210), .ZN(n8346) );
  OR2_X1 U4783 ( .A1(n8530), .A2(n9792), .ZN(n8189) );
  CLKBUF_X2 U4784 ( .A(n5035), .Z(n5466) );
  NAND2_X2 U4785 ( .A1(n5731), .A2(n5730), .ZN(n8165) );
  INV_X2 U4786 ( .A(n9821), .ZN(n5731) );
  BUF_X2 U4788 ( .A(n5788), .Z(n5843) );
  AND3_X2 U4789 ( .A1(n5740), .A2(n5739), .A3(n5738), .ZN(n9785) );
  NAND2_X1 U4790 ( .A1(n5721), .A2(n5720), .ZN(n8407) );
  XNOR2_X1 U4791 ( .A(n5703), .B(P2_IR_REG_29__SCAN_IN), .ZN(n5706) );
  CLKBUF_X1 U4792 ( .A(n10047), .Z(P2_U3966) );
  NOR2_X1 U4793 ( .A1(n6473), .A2(n6204), .ZN(n10047) );
  MUX2_X1 U4794 ( .A(n5521), .B(n5520), .S(n9278), .Z(n5522) );
  INV_X1 U4795 ( .A(n8035), .ZN(n6132) );
  NAND2_X1 U4796 ( .A1(n7951), .A2(n6626), .ZN(n7117) );
  INV_X1 U4797 ( .A(n8743), .ZN(n7762) );
  NAND2_X1 U4798 ( .A1(n5842), .A2(n5841), .ZN(n8219) );
  INV_X2 U4799 ( .A(n7936), .ZN(n6860) );
  AND2_X1 U4800 ( .A1(n4843), .A2(n8071), .ZN(n5020) );
  OAI22_X1 U4801 ( .A1(n7006), .A2(n7007), .B1(n5913), .B2(n5912), .ZN(n7271)
         );
  CLKBUF_X2 U4802 ( .A(n5823), .Z(n8013) );
  AND2_X2 U4803 ( .A1(n5706), .A2(n8878), .ZN(n5828) );
  INV_X1 U4804 ( .A(n5767), .ZN(n6097) );
  INV_X1 U4805 ( .A(n7238), .ZN(n6748) );
  XNOR2_X1 U4806 ( .A(n5701), .B(P2_IR_REG_30__SCAN_IN), .ZN(n5741) );
  INV_X4 U4807 ( .A(n6359), .ZN(n7939) );
  INV_X1 U4808 ( .A(n5030), .ZN(n5480) );
  NAND2_X1 U4809 ( .A1(n4415), .A2(n4947), .ZN(n5345) );
  NAND2_X1 U4810 ( .A1(n4939), .A2(n4938), .ZN(n5272) );
  NAND2_X1 U4811 ( .A1(n6993), .A2(n5898), .ZN(n7006) );
  NAND2_X1 U4812 ( .A1(n7774), .A2(n7771), .ZN(n7784) );
  CLKBUF_X2 U4813 ( .A(n5828), .Z(n8034) );
  BUF_X1 U4814 ( .A(n5741), .Z(n8878) );
  BUF_X1 U4815 ( .A(n5715), .Z(n5720) );
  NAND2_X1 U4816 ( .A1(n5334), .A2(n5333), .ZN(n9319) );
  NAND4_X2 U4817 ( .A1(n5774), .A2(n5773), .A3(n5772), .A4(n5771), .ZN(n8530)
         );
  INV_X1 U4819 ( .A(n5706), .ZN(n7781) );
  INV_X1 U4820 ( .A(n4968), .ZN(n6213) );
  OR2_X1 U4822 ( .A1(n7117), .A2(n8373), .ZN(n9821) );
  NAND4_X4 U4823 ( .A1(n5003), .A2(n5002), .A3(n5001), .A4(n5000), .ZN(n6897)
         );
  NAND3_X1 U4824 ( .A1(n5710), .A2(n5709), .A3(n5708), .ZN(n6644) );
  AOI211_X1 U4825 ( .C1(n9087), .C2(n9278), .A(n5499), .B(n5619), .ZN(n5523)
         );
  CLKBUF_X1 U4826 ( .A(n5020), .Z(n4277) );
  BUF_X4 U4827 ( .A(n5020), .Z(n4278) );
  INV_X2 U4828 ( .A(n6213), .ZN(n4279) );
  INV_X2 U4829 ( .A(n6213), .ZN(n4280) );
  CLKBUF_X1 U4830 ( .A(n7764), .Z(n4281) );
  OAI21_X2 U4831 ( .B1(n5272), .B2(n4944), .A(n4943), .ZN(n5288) );
  AOI21_X1 U4832 ( .B1(n4432), .B2(n4805), .A(n5474), .ZN(n5514) );
  NAND2_X1 U4833 ( .A1(n4320), .A2(n4380), .ZN(n8741) );
  NAND2_X1 U4834 ( .A1(n5995), .A2(n5994), .ZN(n7771) );
  NAND2_X1 U4835 ( .A1(n7650), .A2(n7649), .ZN(n7748) );
  AOI21_X1 U4836 ( .B1(n4719), .B2(n7785), .A(n4717), .ZN(n4716) );
  INV_X1 U4837 ( .A(n4719), .ZN(n4718) );
  NAND2_X1 U4838 ( .A1(n5352), .A2(n5351), .ZN(n9324) );
  AND2_X1 U4839 ( .A1(n6081), .A2(n6080), .ZN(n8692) );
  XNOR2_X1 U4840 ( .A(n5317), .B(n5316), .ZN(n7003) );
  NAND2_X1 U4841 ( .A1(n6825), .A2(n6824), .ZN(n4712) );
  OAI21_X1 U4842 ( .B1(n7294), .B2(n4609), .A(n4606), .ZN(n7355) );
  NAND2_X1 U4843 ( .A1(n7956), .A2(n7957), .ZN(n7955) );
  OAI21_X1 U4844 ( .B1(n5237), .B2(n5236), .A(n4932), .ZN(n5254) );
  NAND2_X1 U4845 ( .A1(n5919), .A2(n5918), .ZN(n9818) );
  NAND2_X1 U4846 ( .A1(n5161), .A2(n5160), .ZN(n9433) );
  NAND2_X1 U4847 ( .A1(n8225), .A2(n8224), .ZN(n8345) );
  INV_X2 U4848 ( .A(n8734), .ZN(n9772) );
  NAND2_X1 U4849 ( .A1(n6166), .A2(n6165), .ZN(n8511) );
  AND2_X1 U4850 ( .A1(n5779), .A2(n5766), .ZN(n4715) );
  AND2_X1 U4851 ( .A1(n5822), .A2(n5821), .ZN(n7965) );
  NAND2_X1 U4852 ( .A1(n9007), .A2(n9633), .ZN(n5599) );
  NAND2_X2 U4853 ( .A1(n6660), .A2(P1_STATE_REG_SCAN_IN), .ZN(n8989) );
  NAND2_X1 U4854 ( .A1(n8197), .A2(n8185), .ZN(n8342) );
  INV_X2 U4855 ( .A(n9600), .ZN(n4283) );
  NAND4_X1 U4856 ( .A1(n5793), .A2(n5792), .A3(n5791), .A4(n5790), .ZN(n8529)
         );
  INV_X2 U4857 ( .A(n6630), .ZN(n6629) );
  NAND4_X1 U4858 ( .A1(n5806), .A2(n5805), .A3(n5804), .A4(n5803), .ZN(n8528)
         );
  INV_X1 U4859 ( .A(n6937), .ZN(n9612) );
  NOR2_X2 U4860 ( .A1(n6384), .A2(n6355), .ZN(n7904) );
  INV_X1 U4861 ( .A(n9761), .ZN(n6733) );
  INV_X1 U4862 ( .A(n8166), .ZN(n8167) );
  INV_X2 U4863 ( .A(n5753), .ZN(n6253) );
  INV_X2 U4864 ( .A(n6384), .ZN(n7933) );
  AND2_X2 U4865 ( .A1(n6280), .A2(P1_STATE_REG_SCAN_IN), .ZN(P1_U4006) );
  BUF_X2 U4866 ( .A(n5119), .Z(n5492) );
  INV_X2 U4867 ( .A(n5027), .ZN(n5509) );
  INV_X2 U4868 ( .A(n6283), .ZN(n5303) );
  MUX2_X1 U4869 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5719), .S(
        P2_IR_REG_27__SCAN_IN), .Z(n5721) );
  NAND2_X1 U4870 ( .A1(n8874), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5701) );
  XNOR2_X1 U4871 ( .A(n5729), .B(P2_IR_REG_19__SCAN_IN), .ZN(n7764) );
  XNOR2_X1 U4872 ( .A(n4841), .B(P1_IR_REG_29__SCAN_IN), .ZN(n4852) );
  INV_X2 U4873 ( .A(n7059), .ZN(n4284) );
  AND2_X2 U4874 ( .A1(n4687), .A2(n4686), .ZN(n4968) );
  NAND2_X1 U4875 ( .A1(n4869), .A2(n4868), .ZN(n4687) );
  NAND2_X1 U4876 ( .A1(n4865), .A2(P1_ADDR_REG_19__SCAN_IN), .ZN(n4686) );
  AND2_X1 U4877 ( .A1(n5028), .A2(n4823), .ZN(n5059) );
  AND2_X1 U4878 ( .A1(n4463), .A2(n4462), .ZN(n5754) );
  INV_X1 U4879 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n5980) );
  INV_X1 U4880 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n6134) );
  INV_X1 U4881 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n5723) );
  INV_X1 U4882 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n5914) );
  NOR2_X1 U4883 ( .A1(P2_IR_REG_11__SCAN_IN), .A2(P2_IR_REG_15__SCAN_IN), .ZN(
        n5688) );
  INV_X4 U4884 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3084) );
  NOR2_X1 U4885 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5028) );
  INV_X1 U4886 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n5861) );
  NOR2_X1 U4887 ( .A1(P2_IR_REG_2__SCAN_IN), .A2(P2_IR_REG_3__SCAN_IN), .ZN(
        n4790) );
  INV_X1 U4888 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n5839) );
  NOR2_X2 U4889 ( .A1(n7802), .A2(n8074), .ZN(n8129) );
  XNOR2_X2 U4890 ( .A(n5726), .B(P2_IR_REG_21__SCAN_IN), .ZN(n5733) );
  XNOR2_X2 U4891 ( .A(n5717), .B(n5716), .ZN(n6183) );
  AOI21_X1 U4892 ( .B1(n8769), .B2(n8676), .A(n4628), .ZN(n4627) );
  NAND2_X1 U4893 ( .A1(n4383), .A2(n4385), .ZN(n4910) );
  INV_X1 U4894 ( .A(n4386), .ZN(n4385) );
  OAI21_X1 U4895 ( .B1(n4388), .B2(n4387), .A(n4817), .ZN(n4386) );
  AND2_X1 U4896 ( .A1(n5617), .A2(n9281), .ZN(n4349) );
  AOI21_X1 U4897 ( .B1(n4662), .B2(n4664), .A(n4316), .ZN(n4660) );
  AOI21_X1 U4898 ( .B1(n4709), .B2(n4707), .A(n4340), .ZN(n4706) );
  INV_X1 U4899 ( .A(n8009), .ZN(n4707) );
  NAND2_X1 U4900 ( .A1(n4483), .A2(n8686), .ZN(n4397) );
  NAND2_X1 U4901 ( .A1(n8669), .A2(n8672), .ZN(n4398) );
  NAND2_X1 U4902 ( .A1(n4843), .A2(n4852), .ZN(n5035) );
  NAND2_X1 U4903 ( .A1(n7855), .A2(n4852), .ZN(n5119) );
  NAND2_X1 U4904 ( .A1(n5516), .A2(n5515), .ZN(n5531) );
  NOR2_X1 U4905 ( .A1(n9289), .A2(n9114), .ZN(n8097) );
  OR2_X1 U4906 ( .A1(n8762), .A2(n8162), .ZN(n8331) );
  INV_X1 U4907 ( .A(n4642), .ZN(n4641) );
  OAI21_X1 U4908 ( .B1(n8392), .B2(n4643), .A(n8365), .ZN(n4642) );
  OR2_X1 U4909 ( .A1(n8785), .A2(n8459), .ZN(n8307) );
  NOR2_X1 U4910 ( .A1(n8392), .A2(n4785), .ZN(n4783) );
  OR2_X1 U4911 ( .A1(n8806), .A2(n8686), .ZN(n8298) );
  NAND2_X1 U4912 ( .A1(n8246), .A2(n4395), .ZN(n4795) );
  OR2_X1 U4913 ( .A1(n8848), .A2(n4396), .ZN(n4395) );
  AND2_X1 U4914 ( .A1(n8521), .A2(n7453), .ZN(n4396) );
  OR2_X1 U4915 ( .A1(n8848), .A2(n9818), .ZN(n4490) );
  OR2_X1 U4916 ( .A1(n8848), .A2(n7453), .ZN(n8245) );
  NAND2_X1 U4917 ( .A1(n8528), .A2(n6748), .ZN(n8210) );
  NAND2_X1 U4918 ( .A1(n4321), .A2(n5723), .ZN(n4723) );
  OAI21_X1 U4919 ( .B1(n5512), .B2(n5515), .A(n5516), .ZN(n5617) );
  AND2_X1 U4920 ( .A1(n9070), .A2(n4657), .ZN(n5619) );
  NAND2_X1 U4921 ( .A1(n9066), .A2(n8998), .ZN(n4657) );
  BUF_X1 U4922 ( .A(n4842), .Z(n4843) );
  NAND2_X1 U4923 ( .A1(n9284), .A2(n8999), .ZN(n8122) );
  NAND2_X1 U4924 ( .A1(n4290), .A2(n4295), .ZN(n4753) );
  NAND2_X1 U4925 ( .A1(n9167), .A2(n8089), .ZN(n4746) );
  NOR2_X1 U4926 ( .A1(n9408), .A2(n4766), .ZN(n4765) );
  NOR2_X1 U4927 ( .A1(n7695), .A2(n7697), .ZN(n4766) );
  OR2_X1 U4928 ( .A1(n9008), .A2(n9618), .ZN(n5638) );
  NAND2_X1 U4929 ( .A1(n5458), .A2(n5457), .ZN(n5460) );
  NAND2_X1 U4930 ( .A1(n5365), .A2(n5364), .ZN(n4975) );
  INV_X1 U4931 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n4832) );
  INV_X1 U4932 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n4768) );
  NAND2_X1 U4933 ( .A1(n4402), .A2(n4924), .ZN(n5237) );
  OR2_X1 U4934 ( .A1(n5194), .A2(n4925), .ZN(n4402) );
  XNOR2_X1 U4935 ( .A(n4892), .B(SI_7_), .ZN(n5104) );
  XNOR2_X1 U4936 ( .A(n4889), .B(SI_6_), .ZN(n5087) );
  NAND2_X1 U4937 ( .A1(n4887), .A2(n4886), .ZN(n5088) );
  INV_X1 U4938 ( .A(n5004), .ZN(n4655) );
  NAND2_X1 U4939 ( .A1(n4706), .A2(n4703), .ZN(n4702) );
  NAND2_X1 U4940 ( .A1(n4708), .A2(n4704), .ZN(n4703) );
  AND2_X1 U4941 ( .A1(n5897), .A2(n5880), .ZN(n4711) );
  XNOR2_X1 U4942 ( .A(n8035), .B(n9785), .ZN(n5748) );
  OR2_X1 U4943 ( .A1(n7111), .A2(n6158), .ZN(n6182) );
  NAND2_X1 U4944 ( .A1(n8383), .A2(n4281), .ZN(n8372) );
  INV_X1 U4945 ( .A(n8034), .ZN(n8001) );
  AND2_X1 U4946 ( .A1(n5706), .A2(n5707), .ZN(n5923) );
  NOR2_X1 U4947 ( .A1(n8587), .A2(n8586), .ZN(n8585) );
  AND2_X1 U4948 ( .A1(n8030), .A2(n8029), .ZN(n8583) );
  OR2_X1 U4949 ( .A1(n4652), .A2(n8613), .ZN(n4647) );
  OR2_X1 U4950 ( .A1(n8785), .A2(n8604), .ZN(n8395) );
  OR2_X1 U4951 ( .A1(n8705), .A2(n8722), .ZN(n8292) );
  AND2_X1 U4952 ( .A1(n8705), .A2(n8516), .ZN(n4803) );
  NAND2_X1 U4953 ( .A1(n7748), .A2(n4788), .ZN(n4380) );
  OR2_X1 U4954 ( .A1(n8848), .A2(n8521), .ZN(n7326) );
  AND2_X1 U4955 ( .A1(n6646), .A2(n6163), .ZN(n8849) );
  NAND2_X1 U4956 ( .A1(n5727), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5728) );
  XNOR2_X1 U4957 ( .A(n6653), .B(n6860), .ZN(n6716) );
  NAND2_X1 U4958 ( .A1(n6652), .A2(n6651), .ZN(n6653) );
  OAI21_X1 U4959 ( .B1(n4286), .B2(n4565), .A(n4564), .ZN(n4563) );
  NOR2_X1 U4960 ( .A1(n4567), .A2(n4566), .ZN(n4565) );
  NAND2_X1 U4961 ( .A1(n4286), .A2(n8882), .ZN(n4564) );
  NAND2_X1 U4962 ( .A1(n6283), .A2(n4499), .ZN(n5030) );
  NAND2_X1 U4963 ( .A1(n6283), .A2(n4280), .ZN(n5027) );
  NAND2_X1 U4964 ( .A1(n8926), .A2(n8924), .ZN(n4550) );
  OR2_X1 U4965 ( .A1(n9111), .A2(n6359), .ZN(n7928) );
  OR2_X1 U4966 ( .A1(n6976), .A2(n9277), .ZN(n6388) );
  INV_X2 U4967 ( .A(n5019), .ZN(n5484) );
  INV_X2 U4968 ( .A(n4278), .ZN(n5419) );
  NOR2_X1 U4969 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(P1_IR_REG_2__SCAN_IN), .ZN(
        n4823) );
  NAND2_X1 U4970 ( .A1(n9084), .A2(n8122), .ZN(n4496) );
  NAND2_X1 U4971 ( .A1(n4742), .A2(n4746), .ZN(n4741) );
  OR2_X1 U4972 ( .A1(n9437), .A2(n8077), .ZN(n4815) );
  OR2_X1 U4973 ( .A1(n8074), .A2(n9260), .ZN(n8075) );
  OR2_X1 U4974 ( .A1(n9575), .A2(n9639), .ZN(n5574) );
  OR2_X1 U4975 ( .A1(n4839), .A2(n4838), .ZN(n4841) );
  INV_X1 U4976 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n5524) );
  AND2_X1 U4977 ( .A1(n6255), .A2(n6193), .ZN(n8753) );
  INV_X1 U4978 ( .A(n8411), .ZN(n4629) );
  AOI21_X1 U4979 ( .B1(n5175), .B2(n5174), .A(n5173), .ZN(n4351) );
  OAI21_X1 U4980 ( .B1(n5607), .B2(n8117), .A(n8118), .ZN(n5405) );
  OR2_X1 U4981 ( .A1(n9134), .A2(n8114), .ZN(n5400) );
  AOI21_X1 U4982 ( .B1(n4682), .B2(n4684), .A(SI_29_), .ZN(n4681) );
  NOR2_X1 U4983 ( .A1(n4580), .A2(n4576), .ZN(n4575) );
  INV_X1 U4984 ( .A(n7885), .ZN(n4576) );
  INV_X1 U4985 ( .A(n4581), .ZN(n4580) );
  INV_X1 U4986 ( .A(n5475), .ZN(n4684) );
  AND2_X1 U4987 ( .A1(n5208), .A2(n5211), .ZN(n4921) );
  INV_X1 U4988 ( .A(n4921), .ZN(n4675) );
  INV_X1 U4989 ( .A(n4637), .ZN(n4636) );
  OAI21_X1 U4990 ( .B1(n4641), .B2(n4638), .A(n4314), .ZN(n4637) );
  INV_X1 U4991 ( .A(n8613), .ZN(n4651) );
  INV_X1 U4992 ( .A(n4649), .ZN(n4633) );
  AOI21_X1 U4993 ( .B1(n8310), .B2(n4650), .A(n8313), .ZN(n4649) );
  INV_X1 U4994 ( .A(n8307), .ZN(n4650) );
  NOR2_X1 U4995 ( .A1(n4638), .A2(n4643), .ZN(n4635) );
  AOI21_X1 U4996 ( .B1(n4622), .B2(n4623), .A(n4621), .ZN(n4620) );
  NAND2_X1 U4997 ( .A1(n8295), .A2(n4626), .ZN(n4621) );
  INV_X1 U4998 ( .A(n4820), .ZN(n4622) );
  INV_X1 U4999 ( .A(n8672), .ZN(n4626) );
  NOR2_X1 U5000 ( .A1(n8684), .A2(n4624), .ZN(n4623) );
  INV_X1 U5001 ( .A(n8292), .ZN(n4624) );
  OR2_X1 U5002 ( .A1(n8810), .A2(n8700), .ZN(n8293) );
  AOI21_X1 U5003 ( .B1(n4615), .B2(n4617), .A(n4614), .ZN(n4613) );
  INV_X1 U5004 ( .A(n8262), .ZN(n4614) );
  OR2_X1 U5005 ( .A1(n7647), .A2(n8050), .ZN(n8262) );
  INV_X1 U5006 ( .A(n4490), .ZN(n4489) );
  NAND2_X1 U5007 ( .A1(n7445), .A2(n8245), .ZN(n7330) );
  INV_X1 U5008 ( .A(n8241), .ZN(n4599) );
  INV_X1 U5009 ( .A(n4598), .ZN(n4597) );
  OAI21_X1 U5010 ( .B1(n8234), .B2(n4599), .A(n8242), .ZN(n4598) );
  OR2_X1 U5011 ( .A1(n9818), .A2(n7442), .ZN(n8242) );
  NAND2_X1 U5012 ( .A1(n7355), .A2(n8233), .ZN(n7077) );
  NOR2_X1 U5013 ( .A1(n8345), .A2(n4611), .ZN(n4610) );
  INV_X1 U5014 ( .A(n7049), .ZN(n4611) );
  INV_X1 U5015 ( .A(n7048), .ZN(n4608) );
  NAND2_X1 U5016 ( .A1(n6852), .A2(n7238), .ZN(n8194) );
  NAND2_X1 U5017 ( .A1(n6578), .A2(n6629), .ZN(n8197) );
  NAND2_X1 U5018 ( .A1(n9785), .A2(n6630), .ZN(n8185) );
  INV_X1 U5019 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n4588) );
  INV_X1 U5020 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n4799) );
  AND2_X1 U5021 ( .A1(n7893), .A2(n4583), .ZN(n4582) );
  INV_X1 U5022 ( .A(n8909), .ZN(n4583) );
  AOI21_X1 U5023 ( .B1(n4582), .B2(n7894), .A(n4333), .ZN(n4581) );
  INV_X1 U5024 ( .A(n6719), .ZN(n4356) );
  INV_X1 U5025 ( .A(n6437), .ZN(n4408) );
  NOR2_X1 U5026 ( .A1(n4527), .A2(n8117), .ZN(n4526) );
  INV_X1 U5027 ( .A(n4529), .ZN(n4527) );
  NAND2_X1 U5028 ( .A1(n9125), .A2(n9151), .ZN(n4473) );
  AND2_X1 U5029 ( .A1(n8113), .A2(n5403), .ZN(n4531) );
  NOR2_X1 U5030 ( .A1(n4739), .A2(n4735), .ZN(n4734) );
  INV_X1 U5031 ( .A(n4744), .ZN(n4735) );
  NAND2_X1 U5032 ( .A1(n4746), .A2(n4304), .ZN(n4740) );
  NOR2_X1 U5033 ( .A1(n8088), .A2(n4745), .ZN(n4744) );
  INV_X1 U5034 ( .A(n4811), .ZN(n4745) );
  AND2_X1 U5035 ( .A1(n5538), .A2(n9224), .ZN(n8107) );
  OR2_X1 U5036 ( .A1(n9334), .A2(n8928), .ZN(n5538) );
  OAI21_X1 U5037 ( .B1(n4504), .B2(n9249), .A(n8103), .ZN(n4502) );
  INV_X1 U5038 ( .A(n7799), .ZN(n4508) );
  NAND2_X1 U5039 ( .A1(n7795), .A2(n4761), .ZN(n4760) );
  INV_X1 U5040 ( .A(n4762), .ZN(n4761) );
  AND2_X1 U5041 ( .A1(n5539), .A2(n7797), .ZN(n9400) );
  AND2_X1 U5042 ( .A1(n7580), .A2(n7578), .ZN(n7419) );
  AND2_X1 U5043 ( .A1(n5139), .A2(n5563), .ZN(n4540) );
  AOI21_X1 U5044 ( .B1(n4514), .B2(n4517), .A(n4511), .ZN(n4510) );
  INV_X1 U5045 ( .A(n4514), .ZN(n4512) );
  INV_X1 U5046 ( .A(n5574), .ZN(n4517) );
  NAND2_X1 U5047 ( .A1(n5573), .A2(n5599), .ZN(n5078) );
  OR2_X1 U5048 ( .A1(n6448), .A2(n9612), .ZN(n5541) );
  XNOR2_X1 U5049 ( .A(n6897), .B(n6795), .ZN(n6895) );
  AND2_X1 U5050 ( .A1(n5534), .A2(n9168), .ZN(n8113) );
  AND2_X1 U5051 ( .A1(n9314), .A2(n8089), .ZN(n8112) );
  XNOR2_X1 U5052 ( .A(n5503), .B(n5502), .ZN(n5500) );
  NAND2_X1 U5053 ( .A1(n5438), .A2(n5437), .ZN(n5458) );
  NAND2_X1 U5054 ( .A1(n4667), .A2(n4665), .ZN(n5438) );
  AOI21_X1 U5055 ( .B1(n4668), .B2(n4327), .A(n4666), .ZN(n4665) );
  INV_X1 U5056 ( .A(n4669), .ZN(n4668) );
  OAI21_X1 U5057 ( .B1(n4672), .B2(n4327), .A(n5409), .ZN(n4669) );
  AND2_X1 U5058 ( .A1(n4962), .A2(n4961), .ZN(n5329) );
  AND2_X1 U5059 ( .A1(n4938), .A2(n4937), .ZN(n5253) );
  NOR2_X1 U5060 ( .A1(n5177), .A2(n4678), .ZN(n4677) );
  INV_X1 U5061 ( .A(n4913), .ZN(n4678) );
  NAND2_X1 U5062 ( .A1(n4382), .A2(n5156), .ZN(n4679) );
  AND2_X1 U5063 ( .A1(n4816), .A2(n4393), .ZN(n4388) );
  INV_X1 U5064 ( .A(n5108), .ZN(n4393) );
  INV_X1 U5065 ( .A(n4903), .ZN(n4390) );
  INV_X1 U5066 ( .A(n4897), .ZN(n4391) );
  INV_X1 U5067 ( .A(n5087), .ZN(n4888) );
  OAI211_X1 U5068 ( .C1(n4686), .C2(n4436), .A(n4434), .B(n4433), .ZN(n4878)
         );
  NAND2_X1 U5069 ( .A1(n4435), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n4434) );
  OAI211_X1 U5070 ( .C1(n4687), .C2(n4495), .A(n4494), .B(n4493), .ZN(n5004)
         );
  OR2_X1 U5071 ( .A1(n8008), .A2(n8007), .ZN(n8009) );
  NAND2_X1 U5072 ( .A1(n5920), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n5938) );
  NAND2_X1 U5073 ( .A1(n6009), .A2(n6008), .ZN(n7782) );
  NAND2_X1 U5074 ( .A1(n5884), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n5904) );
  INV_X1 U5075 ( .A(n5886), .ZN(n5884) );
  AND2_X1 U5076 ( .A1(n8432), .A2(n6057), .ZN(n6058) );
  INV_X1 U5077 ( .A(n5826), .ZN(n5824) );
  OR2_X1 U5078 ( .A1(n8338), .A2(n8373), .ZN(n8376) );
  OAI21_X1 U5079 ( .B1(n8156), .B2(n8765), .A(n8150), .ZN(n8158) );
  AND2_X1 U5080 ( .A1(n8006), .A2(n8005), .ZN(n8459) );
  NAND2_X1 U5081 ( .A1(n9719), .A2(n6527), .ZN(n4455) );
  NAND2_X1 U5082 ( .A1(n4455), .A2(n4454), .ZN(n4453) );
  INV_X1 U5083 ( .A(n6529), .ZN(n4454) );
  XNOR2_X1 U5084 ( .A(n7152), .B(n8564), .ZN(n8562) );
  NAND2_X1 U5085 ( .A1(n7611), .A2(n7610), .ZN(n9742) );
  NOR3_X1 U5086 ( .A1(n8617), .A2(n8770), .A3(n4479), .ZN(n8574) );
  NAND2_X1 U5087 ( .A1(n4481), .A2(n4480), .ZN(n4479) );
  NOR2_X1 U5088 ( .A1(n8598), .A2(n8775), .ZN(n8582) );
  OAI21_X1 U5089 ( .B1(n8173), .B2(n8613), .A(n8307), .ZN(n4646) );
  OR2_X1 U5090 ( .A1(n8785), .A2(n8633), .ZN(n8617) );
  XNOR2_X1 U5091 ( .A(n8779), .B(n8503), .ZN(n8601) );
  INV_X1 U5092 ( .A(n8173), .ZN(n4638) );
  NAND2_X1 U5093 ( .A1(n4644), .A2(n4641), .ZN(n4652) );
  NAND2_X1 U5094 ( .A1(n8393), .A2(n8644), .ZN(n8394) );
  NAND2_X1 U5095 ( .A1(n8307), .A2(n8308), .ZN(n8613) );
  OR2_X1 U5096 ( .A1(n6186), .A2(n6185), .ZN(n7999) );
  AOI21_X1 U5097 ( .B1(n4783), .B2(n8662), .A(n4317), .ZN(n4781) );
  INV_X1 U5098 ( .A(n4783), .ZN(n4782) );
  NOR2_X1 U5099 ( .A1(n4818), .A2(n8799), .ZN(n8655) );
  NAND2_X1 U5100 ( .A1(n8654), .A2(n8653), .ZN(n8652) );
  INV_X1 U5101 ( .A(n6084), .ZN(n6082) );
  NAND2_X1 U5102 ( .A1(n8692), .A2(n8700), .ZN(n4801) );
  AND2_X1 U5103 ( .A1(n8810), .A2(n8515), .ZN(n4800) );
  AND2_X1 U5104 ( .A1(n6109), .A2(n6108), .ZN(n8686) );
  NAND2_X1 U5105 ( .A1(n8716), .A2(n4820), .ZN(n4625) );
  NAND2_X1 U5106 ( .A1(n8717), .A2(n8718), .ZN(n8716) );
  NAND2_X1 U5107 ( .A1(n6050), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n6066) );
  INV_X1 U5108 ( .A(n6052), .ZN(n6050) );
  NOR2_X1 U5109 ( .A1(n7673), .A2(n7647), .ZN(n7660) );
  AND4_X1 U5110 ( .A1(n6007), .A2(n6006), .A3(n6005), .A4(n6004), .ZN(n7745)
         );
  NAND2_X1 U5111 ( .A1(n7677), .A2(n7597), .ZN(n7681) );
  NOR2_X1 U5112 ( .A1(n8356), .A2(n4798), .ZN(n4796) );
  INV_X1 U5113 ( .A(n7326), .ZN(n4798) );
  NAND2_X1 U5114 ( .A1(n8246), .A2(n8245), .ZN(n7430) );
  NAND2_X1 U5115 ( .A1(n7431), .A2(n7430), .ZN(n7429) );
  AND4_X1 U5116 ( .A1(n5909), .A2(n5908), .A3(n5907), .A4(n5906), .ZN(n7376)
         );
  AND2_X1 U5117 ( .A1(n8234), .A2(n8235), .ZN(n7075) );
  NAND2_X1 U5118 ( .A1(n7357), .A2(n8349), .ZN(n7356) );
  AND4_X1 U5119 ( .A1(n5875), .A2(n5874), .A3(n5873), .A4(n5872), .ZN(n7296)
         );
  NAND2_X1 U5120 ( .A1(n4296), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5729) );
  INV_X1 U5121 ( .A(n4723), .ZN(n4721) );
  INV_X1 U5122 ( .A(n7208), .ZN(n8341) );
  NAND2_X1 U5123 ( .A1(n6038), .A2(n6037), .ZN(n8827) );
  NAND2_X1 U5124 ( .A1(n5936), .A2(n5935), .ZN(n8848) );
  NAND2_X1 U5125 ( .A1(n6327), .A2(n6129), .ZN(n5936) );
  AND2_X1 U5126 ( .A1(n5722), .A2(n5723), .ZN(n6015) );
  INV_X1 U5127 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n5687) );
  NAND2_X1 U5128 ( .A1(n4584), .A2(n4299), .ZN(n7825) );
  NAND2_X1 U5129 ( .A1(n7638), .A2(n4585), .ZN(n4584) );
  AND2_X1 U5130 ( .A1(n4586), .A2(n7635), .ZN(n4585) );
  NAND2_X1 U5131 ( .A1(n4547), .A2(n7877), .ZN(n4546) );
  INV_X1 U5132 ( .A(n8923), .ZN(n4547) );
  INV_X1 U5133 ( .A(n8960), .ZN(n4548) );
  NOR2_X1 U5134 ( .A1(n4549), .A2(n4542), .ZN(n4541) );
  INV_X1 U5135 ( .A(n8924), .ZN(n4542) );
  NOR2_X1 U5136 ( .A1(n7877), .A2(n8960), .ZN(n4549) );
  OAI21_X1 U5137 ( .B1(n7172), .B2(n7171), .A(n7170), .ZN(n7179) );
  OR2_X1 U5138 ( .A1(n6795), .A2(n6384), .ZN(n6385) );
  NAND2_X1 U5139 ( .A1(n7550), .A2(n7549), .ZN(n7633) );
  AOI21_X1 U5140 ( .B1(n6778), .B2(n7933), .A(n6361), .ZN(n6362) );
  NAND2_X1 U5141 ( .A1(n8900), .A2(n8901), .ZN(n7886) );
  NAND2_X1 U5142 ( .A1(n7342), .A2(n7343), .ZN(n7341) );
  AND2_X1 U5143 ( .A1(n7189), .A2(n7393), .ZN(n4551) );
  NAND2_X1 U5144 ( .A1(n7393), .A2(n4557), .ZN(n4556) );
  INV_X1 U5145 ( .A(n7390), .ZN(n4557) );
  NOR4_X1 U5146 ( .A1(n5661), .A2(n5660), .A3(n5627), .A4(n5554), .ZN(n5555)
         );
  AND2_X1 U5147 ( .A1(n5663), .A2(n5662), .ZN(n5666) );
  AND4_X1 U5148 ( .A1(n4857), .A2(n4856), .A3(n4855), .A4(n4854), .ZN(n7947)
         );
  AND4_X1 U5149 ( .A1(n5427), .A2(n5426), .A3(n5425), .A4(n5424), .ZN(n8094)
         );
  AND4_X1 U5150 ( .A1(n5151), .A2(n5150), .A3(n5149), .A4(n5148), .ZN(n9424)
         );
  NAND2_X1 U5151 ( .A1(n4417), .A2(n4416), .ZN(n4418) );
  AOI21_X1 U5152 ( .B1(n4419), .B2(n9487), .A(n9502), .ZN(n4416) );
  NAND2_X1 U5153 ( .A1(n9488), .A2(n4419), .ZN(n4417) );
  NAND2_X1 U5154 ( .A1(n6695), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n4409) );
  NAND2_X1 U5155 ( .A1(n4405), .A2(n4403), .ZN(n6805) );
  NAND2_X1 U5156 ( .A1(n4407), .A2(n4404), .ZN(n4403) );
  NAND2_X1 U5157 ( .A1(n6435), .A2(n4406), .ZN(n4405) );
  INV_X1 U5158 ( .A(n4409), .ZN(n4404) );
  NAND2_X1 U5159 ( .A1(n6435), .A2(n4330), .ZN(n4410) );
  OR2_X1 U5160 ( .A1(n7730), .A2(n7729), .ZN(n4428) );
  NAND2_X1 U5161 ( .A1(n4428), .A2(n4427), .ZN(n4426) );
  NAND2_X1 U5162 ( .A1(n9039), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n4427) );
  NAND2_X1 U5163 ( .A1(n4426), .A2(n4425), .ZN(n9052) );
  INV_X1 U5164 ( .A(n9042), .ZN(n4425) );
  AND4_X1 U5165 ( .A1(n5471), .A2(n5470), .A3(n5469), .A4(n5468), .ZN(n8999)
         );
  NAND2_X1 U5166 ( .A1(n9083), .A2(n4310), .ZN(n9084) );
  NAND2_X1 U5167 ( .A1(n5612), .A2(n8122), .ZN(n9075) );
  NAND2_X1 U5168 ( .A1(n4748), .A2(n4311), .ZN(n9076) );
  NAND2_X1 U5169 ( .A1(n9133), .A2(n4308), .ZN(n4748) );
  INV_X1 U5170 ( .A(n4754), .ZN(n4752) );
  NAND2_X1 U5171 ( .A1(n9082), .A2(n5610), .ZN(n9100) );
  AOI21_X1 U5172 ( .B1(n9112), .B2(n8121), .A(n8120), .ZN(n9101) );
  NAND2_X1 U5173 ( .A1(n4749), .A2(n4753), .ZN(n9107) );
  AOI21_X1 U5174 ( .B1(n4526), .B2(n4524), .A(n4523), .ZN(n4522) );
  INV_X1 U5175 ( .A(n8116), .ZN(n4523) );
  INV_X1 U5176 ( .A(n4531), .ZN(n4524) );
  INV_X1 U5177 ( .A(n4526), .ZN(n4525) );
  NAND2_X1 U5178 ( .A1(n8118), .A2(n8119), .ZN(n9126) );
  AOI21_X1 U5179 ( .B1(n8112), .B2(n5403), .A(n4530), .ZN(n4529) );
  NAND2_X1 U5180 ( .A1(n9169), .A2(n4531), .ZN(n4528) );
  INV_X1 U5181 ( .A(n4740), .ZN(n4739) );
  OR2_X1 U5182 ( .A1(n9319), .A2(n8087), .ZN(n9168) );
  OR2_X1 U5183 ( .A1(n9178), .A2(n9314), .ZN(n9162) );
  NAND2_X1 U5184 ( .A1(n5551), .A2(n4747), .ZN(n4742) );
  OAI21_X1 U5185 ( .B1(n9198), .B2(n8110), .A(n8109), .ZN(n9186) );
  OR2_X1 U5186 ( .A1(n9197), .A2(n8902), .ZN(n4811) );
  OAI21_X1 U5187 ( .B1(n9212), .B2(n9211), .A(n8108), .ZN(n9198) );
  NOR2_X1 U5188 ( .A1(n9329), .A2(n9228), .ZN(n8084) );
  AOI21_X1 U5189 ( .B1(n9218), .B2(n9226), .A(n8083), .ZN(n9205) );
  AND2_X1 U5190 ( .A1(n9334), .A2(n9244), .ZN(n8083) );
  INV_X1 U5191 ( .A(n4505), .ZN(n4504) );
  OAI21_X1 U5192 ( .B1(n4294), .B2(n4506), .A(n8100), .ZN(n4505) );
  NAND2_X1 U5193 ( .A1(n5244), .A2(n5243), .ZN(n8074) );
  AND4_X1 U5194 ( .A1(n5266), .A2(n5265), .A3(n5264), .A4(n5263), .ZN(n8079)
         );
  OR2_X1 U5195 ( .A1(n7719), .A2(n9401), .ZN(n7799) );
  NAND2_X1 U5196 ( .A1(n4765), .A2(n7697), .ZN(n4762) );
  NOR2_X1 U5197 ( .A1(n4764), .A2(n9000), .ZN(n4763) );
  INV_X1 U5198 ( .A(n7695), .ZN(n4764) );
  NAND2_X1 U5199 ( .A1(n4772), .A2(n4770), .ZN(n4769) );
  AND2_X1 U5200 ( .A1(n4297), .A2(n7575), .ZN(n4773) );
  INV_X1 U5201 ( .A(n7574), .ZN(n4772) );
  NAND2_X1 U5202 ( .A1(n5144), .A2(n5143), .ZN(n7571) );
  NAND2_X1 U5203 ( .A1(n7418), .A2(n4297), .ZN(n7573) );
  NAND2_X1 U5204 ( .A1(n4540), .A2(n5124), .ZN(n7487) );
  NAND2_X1 U5205 ( .A1(n4319), .A2(n7413), .ZN(n4729) );
  AND2_X1 U5206 ( .A1(n5116), .A2(n5115), .ZN(n7176) );
  NAND2_X1 U5207 ( .A1(n9593), .A2(n4731), .ZN(n7412) );
  NOR2_X1 U5208 ( .A1(n6952), .A2(n4732), .ZN(n4731) );
  INV_X1 U5209 ( .A(n6948), .ZN(n4732) );
  AND2_X1 U5210 ( .A1(n5574), .A2(n6977), .ZN(n6952) );
  NAND2_X1 U5211 ( .A1(n9578), .A2(n5599), .ZN(n6951) );
  INV_X1 U5212 ( .A(n5078), .ZN(n9596) );
  NAND2_X1 U5213 ( .A1(n4728), .A2(n4727), .ZN(n6947) );
  AND2_X1 U5214 ( .A1(n6946), .A2(n6913), .ZN(n4726) );
  INV_X1 U5215 ( .A(n9618), .ZN(n6921) );
  NAND2_X1 U5216 ( .A1(n5638), .A2(n5559), .ZN(n6911) );
  NAND2_X1 U5217 ( .A1(n6780), .A2(n5017), .ZN(n6929) );
  INV_X1 U5218 ( .A(n9576), .ZN(n9261) );
  AND2_X1 U5219 ( .A1(n6795), .A2(n6794), .ZN(n6936) );
  XNOR2_X1 U5220 ( .A(n6388), .B(n6387), .ZN(n4374) );
  NOR2_X1 U5221 ( .A1(n6360), .A2(n6794), .ZN(n6781) );
  NAND2_X1 U5222 ( .A1(n5482), .A2(n5481), .ZN(n9281) );
  INV_X1 U5223 ( .A(n9111), .ZN(n9294) );
  AND2_X1 U5224 ( .A1(n5107), .A2(n5106), .ZN(n9646) );
  AND3_X1 U5225 ( .A1(n5093), .A2(n5092), .A3(n5091), .ZN(n9639) );
  AND3_X1 U5226 ( .A1(n5064), .A2(n5063), .A3(n5062), .ZN(n9627) );
  NAND2_X2 U5227 ( .A1(n6239), .A2(n5680), .ZN(n6357) );
  NOR2_X1 U5228 ( .A1(n7459), .A2(n7165), .ZN(n5680) );
  XNOR2_X1 U5229 ( .A(n5508), .B(n5507), .ZN(n8872) );
  NAND2_X1 U5230 ( .A1(n5678), .A2(n4777), .ZN(n4776) );
  INV_X1 U5231 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n5674) );
  XNOR2_X1 U5232 ( .A(n5436), .B(n5435), .ZN(n7995) );
  OAI21_X1 U5233 ( .B1(n4975), .B2(n4327), .A(n4668), .ZN(n5436) );
  INV_X1 U5234 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n5676) );
  XNOR2_X1 U5235 ( .A(n5411), .B(n5410), .ZN(n7991) );
  NAND2_X1 U5236 ( .A1(n4671), .A2(n4978), .ZN(n5411) );
  OAI21_X1 U5237 ( .B1(n5288), .B2(n4412), .A(n4411), .ZN(n5365) );
  AOI21_X1 U5238 ( .B1(n4413), .B2(n5287), .A(n4289), .ZN(n4411) );
  INV_X1 U5239 ( .A(n4413), .ZN(n4412) );
  AND2_X1 U5240 ( .A1(n5315), .A2(n5314), .ZN(n5317) );
  AOI21_X1 U5241 ( .B1(n4858), .B2(P1_IR_REG_31__SCAN_IN), .A(n4370), .ZN(
        n4369) );
  NAND2_X1 U5242 ( .A1(n4371), .A2(n5524), .ZN(n4370) );
  NAND2_X1 U5243 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), 
        .ZN(n4371) );
  NAND2_X1 U5244 ( .A1(n4858), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5626) );
  INV_X1 U5245 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n4862) );
  NAND2_X1 U5246 ( .A1(n4372), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4863) );
  XNOR2_X1 U5247 ( .A(n4381), .B(n5177), .ZN(n6327) );
  NAND2_X1 U5248 ( .A1(n4679), .A2(n4913), .ZN(n4381) );
  NAND2_X1 U5249 ( .A1(n4883), .A2(n4882), .ZN(n5073) );
  XNOR2_X1 U5250 ( .A(n4878), .B(SI_3_), .ZN(n5041) );
  NAND2_X1 U5251 ( .A1(n4378), .A2(n4876), .ZN(n5042) );
  XNOR2_X1 U5252 ( .A(n5006), .B(P1_IR_REG_1__SCAN_IN), .ZN(n6289) );
  NOR2_X1 U5253 ( .A1(n4699), .A2(n8511), .ZN(n4697) );
  NAND2_X1 U5254 ( .A1(n4701), .A2(n4705), .ZN(n4700) );
  NAND2_X1 U5255 ( .A1(n4709), .A2(n8038), .ZN(n4705) );
  NAND2_X1 U5256 ( .A1(n5858), .A2(n5857), .ZN(n6825) );
  INV_X1 U5257 ( .A(n9785), .ZN(n6578) );
  AND2_X1 U5258 ( .A1(n6073), .A2(n6072), .ZN(n8722) );
  INV_X1 U5259 ( .A(n9764), .ZN(n5732) );
  AND2_X1 U5260 ( .A1(n7451), .A2(n4693), .ZN(n4692) );
  NAND2_X1 U5261 ( .A1(n7305), .A2(n4694), .ZN(n4693) );
  AND2_X1 U5262 ( .A1(n6125), .A2(n6124), .ZN(n8674) );
  NAND2_X1 U5263 ( .A1(n5762), .A2(n7970), .ZN(n7980) );
  AND3_X1 U5264 ( .A1(n6029), .A2(n6028), .A3(n6027), .ZN(n8494) );
  AND2_X1 U5265 ( .A1(n6180), .A2(n6178), .ZN(n8509) );
  AND2_X1 U5266 ( .A1(n6735), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8496) );
  AND2_X1 U5267 ( .A1(n6473), .A2(n9783), .ZN(n9774) );
  INV_X1 U5268 ( .A(n8459), .ZN(n8604) );
  NAND2_X1 U5269 ( .A1(n8013), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n5805) );
  NAND2_X1 U5270 ( .A1(n9732), .A2(n6556), .ZN(n6705) );
  NOR2_X1 U5271 ( .A1(n6705), .A2(n6704), .ZN(n6703) );
  INV_X1 U5272 ( .A(n7614), .ZN(n8057) );
  AND2_X1 U5273 ( .A1(n6479), .A2(n6478), .ZN(n9748) );
  OAI21_X1 U5274 ( .B1(n8065), .B2(n9692), .A(n4459), .ZN(n4458) );
  AOI21_X1 U5275 ( .B1(n8066), .B2(n9748), .A(n9747), .ZN(n4459) );
  OAI21_X1 U5276 ( .B1(n8068), .B2(n4866), .A(n8429), .ZN(n4457) );
  XNOR2_X1 U5277 ( .A(n4379), .B(n8368), .ZN(n8773) );
  NAND2_X1 U5278 ( .A1(n8579), .A2(n8397), .ZN(n4379) );
  AOI211_X1 U5279 ( .C1(n4482), .C2(n8770), .A(n8574), .B(n4275), .ZN(n8769)
         );
  INV_X1 U5280 ( .A(n8582), .ZN(n4482) );
  NAND2_X1 U5281 ( .A1(n8410), .A2(n8409), .ZN(n4631) );
  AOI22_X1 U5282 ( .A1(n8603), .A2(n8753), .B1(n8570), .B2(n8513), .ZN(n8409)
         );
  NOR3_X1 U5283 ( .A1(n8591), .A2(n8590), .A3(n8589), .ZN(n8777) );
  AND2_X1 U5284 ( .A1(n8615), .A2(n8753), .ZN(n8589) );
  NAND2_X1 U5285 ( .A1(n6020), .A2(n6019), .ZN(n8834) );
  NAND2_X1 U5286 ( .A1(n8734), .A2(n7118), .ZN(n9768) );
  NAND2_X1 U5287 ( .A1(n8734), .A2(n7115), .ZN(n8761) );
  NOR2_X1 U5288 ( .A1(n4561), .A2(n8984), .ZN(n4559) );
  AND2_X1 U5289 ( .A1(n4325), .A2(n4563), .ZN(n4561) );
  NAND2_X1 U5290 ( .A1(n4563), .A2(n4334), .ZN(n4562) );
  NAND2_X1 U5291 ( .A1(n5462), .A2(n5461), .ZN(n9284) );
  OR2_X1 U5292 ( .A1(n7179), .A2(n7178), .ZN(n7345) );
  NAND2_X1 U5293 ( .A1(n7861), .A2(n7860), .ZN(n8926) );
  AND2_X1 U5294 ( .A1(n7347), .A2(n9345), .ZN(n8968) );
  AND4_X1 U5295 ( .A1(n4998), .A2(n4997), .A3(n4996), .A4(n4995), .ZN(n8977)
         );
  NAND2_X1 U5296 ( .A1(n4360), .A2(n4358), .ZN(n8971) );
  NAND2_X1 U5297 ( .A1(n4359), .A2(n4328), .ZN(n4358) );
  INV_X1 U5298 ( .A(n8917), .ZN(n4359) );
  NAND2_X2 U5299 ( .A1(n5040), .A2(n5039), .ZN(n9008) );
  OR2_X1 U5300 ( .A1(n5419), .A2(n6268), .ZN(n5040) );
  AND3_X1 U5301 ( .A1(n5038), .A2(n5037), .A3(n5036), .ZN(n5039) );
  NOR2_X1 U5302 ( .A1(n6315), .A2(n6276), .ZN(n6279) );
  NOR2_X1 U5303 ( .A1(n6279), .A2(n6278), .ZN(n6430) );
  INV_X1 U5304 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n4868) );
  OAI21_X1 U5305 ( .B1(n9060), .B2(n9551), .A(n4424), .ZN(n4423) );
  AND2_X1 U5306 ( .A1(n9059), .A2(n9538), .ZN(n4424) );
  XNOR2_X1 U5307 ( .A(n9064), .B(n9270), .ZN(n9269) );
  AOI21_X1 U5308 ( .B1(n9269), .B2(n9572), .A(n4469), .ZN(n4468) );
  OAI21_X1 U5309 ( .B1(n9270), .B2(n9658), .A(n9274), .ZN(n4469) );
  MUX2_X1 U5310 ( .A(n5235), .B(n5234), .S(n5483), .Z(n5252) );
  AOI21_X1 U5311 ( .B1(n5232), .B2(n5546), .A(n5231), .ZN(n5233) );
  AND2_X1 U5312 ( .A1(n9242), .A2(n5286), .ZN(n4347) );
  AND2_X1 U5313 ( .A1(n5537), .A2(n5538), .ZN(n4352) );
  AOI21_X1 U5314 ( .B1(n5406), .B2(n5483), .A(n4821), .ZN(n5407) );
  AND2_X1 U5315 ( .A1(n8116), .A2(n5403), .ZN(n5607) );
  NAND2_X1 U5316 ( .A1(n5402), .A2(n7917), .ZN(n5404) );
  INV_X1 U5317 ( .A(n5155), .ZN(n4539) );
  OR2_X1 U5318 ( .A1(n8770), .A2(n8588), .ZN(n8326) );
  INV_X1 U5319 ( .A(n4616), .ZN(n4615) );
  OAI21_X1 U5320 ( .B1(n7597), .B2(n4617), .A(n8259), .ZN(n4616) );
  INV_X1 U5321 ( .A(n8257), .ZN(n4617) );
  OR2_X1 U5322 ( .A1(n9281), .A2(n9087), .ZN(n4431) );
  NAND2_X1 U5323 ( .A1(n9281), .A2(n5483), .ZN(n4430) );
  NAND2_X1 U5324 ( .A1(n5514), .A2(n4349), .ZN(n5519) );
  NOR2_X1 U5325 ( .A1(n8097), .A2(n4756), .ZN(n4755) );
  INV_X1 U5326 ( .A(n8096), .ZN(n4756) );
  INV_X1 U5327 ( .A(n5404), .ZN(n8117) );
  OR2_X1 U5328 ( .A1(n7571), .A2(n9424), .ZN(n7580) );
  AND2_X1 U5329 ( .A1(n5601), .A2(n4515), .ZN(n4514) );
  NAND2_X1 U5330 ( .A1(n5574), .A2(n4516), .ZN(n4515) );
  INV_X1 U5331 ( .A(n5562), .ZN(n4511) );
  NAND2_X1 U5332 ( .A1(n7581), .A2(n7580), .ZN(n9422) );
  OAI21_X1 U5333 ( .B1(n5124), .B2(n4539), .A(n4537), .ZN(n7581) );
  INV_X1 U5334 ( .A(n4538), .ZN(n4537) );
  OAI21_X1 U5335 ( .B1(n4540), .B2(n4539), .A(n7578), .ZN(n4538) );
  AOI21_X1 U5336 ( .B1(n4683), .B2(n5475), .A(n4342), .ZN(n4682) );
  INV_X1 U5337 ( .A(n5459), .ZN(n4683) );
  INV_X1 U5338 ( .A(n5435), .ZN(n4666) );
  NAND2_X1 U5339 ( .A1(n4900), .A2(n4899), .ZN(n4903) );
  INV_X1 U5340 ( .A(n4663), .ZN(n4662) );
  OAI21_X1 U5341 ( .B1(n4888), .B2(n4664), .A(n4891), .ZN(n4663) );
  INV_X1 U5342 ( .A(n4890), .ZN(n4664) );
  NAND2_X1 U5343 ( .A1(n4864), .A2(P2_ADDR_REG_19__SCAN_IN), .ZN(n4865) );
  INV_X1 U5344 ( .A(P2_RD_REG_SCAN_IN), .ZN(n4864) );
  AND2_X1 U5345 ( .A1(n4448), .A2(n6501), .ZN(n4440) );
  OR3_X1 U5346 ( .A1(n8028), .A2(n8027), .A3(n8026), .ZN(n8029) );
  OR2_X1 U5347 ( .A1(n8775), .A2(n8416), .ZN(n8401) );
  NOR2_X1 U5348 ( .A1(n8705), .A2(n8823), .ZN(n4484) );
  AND2_X1 U5349 ( .A1(n7747), .A2(n7756), .ZN(n4788) );
  NOR2_X1 U5350 ( .A1(n7215), .A2(n6747), .ZN(n6770) );
  NAND2_X1 U5351 ( .A1(n8645), .A2(n8393), .ZN(n8633) );
  AND2_X1 U5352 ( .A1(n4654), .A2(n8655), .ZN(n8645) );
  NAND2_X1 U5353 ( .A1(n8725), .A2(n4285), .ZN(n8687) );
  AND2_X1 U5354 ( .A1(n4602), .A2(n4799), .ZN(n4600) );
  NOR2_X1 U5355 ( .A1(P2_IR_REG_26__SCAN_IN), .A2(P2_IR_REG_27__SCAN_IN), .ZN(
        n4602) );
  NOR2_X1 U5356 ( .A1(n4723), .A2(n4725), .ZN(n4722) );
  INV_X1 U5357 ( .A(n5724), .ZN(n4725) );
  OR3_X1 U5358 ( .A1(n5933), .A2(P2_IR_REG_11__SCAN_IN), .A3(
        P2_IR_REG_10__SCAN_IN), .ZN(n5948) );
  NAND2_X1 U5359 ( .A1(n7706), .A2(n7705), .ZN(n4586) );
  AOI21_X1 U5360 ( .B1(n4581), .B2(n4579), .A(n4578), .ZN(n4577) );
  NAND2_X1 U5361 ( .A1(n7886), .A2(n4575), .ZN(n4574) );
  INV_X1 U5362 ( .A(n4582), .ZN(n4579) );
  AND2_X1 U5363 ( .A1(n9281), .A2(n7947), .ZN(n5654) );
  AND2_X1 U5364 ( .A1(n9270), .A2(n9066), .ZN(n5661) );
  AND2_X1 U5365 ( .A1(n4330), .A2(n4407), .ZN(n4406) );
  INV_X1 U5366 ( .A(n6697), .ZN(n4407) );
  OR2_X1 U5367 ( .A1(n9284), .A2(n8999), .ZN(n5612) );
  AOI21_X1 U5368 ( .B1(n9100), .B2(n4757), .A(n8097), .ZN(n4754) );
  NAND2_X1 U5369 ( .A1(n4755), .A2(n4751), .ZN(n4750) );
  INV_X1 U5370 ( .A(n4753), .ZN(n4751) );
  AND2_X1 U5371 ( .A1(n9294), .A2(n8094), .ZN(n8120) );
  OR2_X1 U5372 ( .A1(n9294), .A2(n8094), .ZN(n8121) );
  AND2_X1 U5373 ( .A1(n9324), .A2(n8902), .ZN(n8110) );
  OR2_X1 U5374 ( .A1(n9324), .A2(n8902), .ZN(n8109) );
  NOR2_X1 U5375 ( .A1(n9339), .A2(n9344), .ZN(n4476) );
  AND2_X1 U5376 ( .A1(n5245), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n5260) );
  NAND2_X1 U5377 ( .A1(n7575), .A2(n4771), .ZN(n4770) );
  INV_X1 U5378 ( .A(n7572), .ZN(n4771) );
  OR2_X1 U5379 ( .A1(n7408), .A2(n7409), .ZN(n7413) );
  OR2_X1 U5380 ( .A1(n7484), .A2(n5138), .ZN(n5155) );
  NAND2_X1 U5381 ( .A1(n5563), .A2(n5581), .ZN(n7406) );
  NOR2_X1 U5382 ( .A1(n9573), .A2(n7026), .ZN(n6982) );
  INV_X1 U5383 ( .A(n4978), .ZN(n4670) );
  NOR2_X1 U5384 ( .A1(n4979), .A2(n4673), .ZN(n4672) );
  INV_X1 U5385 ( .A(n4974), .ZN(n4673) );
  INV_X1 U5386 ( .A(n4966), .ZN(n4967) );
  NOR2_X1 U5387 ( .A1(n4960), .A2(n4414), .ZN(n4413) );
  INV_X1 U5388 ( .A(n4947), .ZN(n4414) );
  OR2_X1 U5389 ( .A1(n5313), .A2(n5316), .ZN(n4960) );
  OR2_X1 U5390 ( .A1(n5328), .A2(n4965), .ZN(n5313) );
  OR2_X1 U5391 ( .A1(n4965), .A2(n4964), .ZN(n5314) );
  AND2_X1 U5392 ( .A1(n5329), .A2(n5331), .ZN(n4964) );
  AND4_X1 U5393 ( .A1(n4830), .A2(n5239), .A3(n4829), .A4(n4828), .ZN(n4807)
         );
  INV_X1 U5394 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n4830) );
  INV_X1 U5395 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n4829) );
  INV_X1 U5396 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n4828) );
  INV_X1 U5397 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n5239) );
  AOI21_X1 U5398 ( .B1(n4910), .B2(n4401), .A(n4674), .ZN(n5194) );
  AND2_X1 U5399 ( .A1(n4676), .A2(n4909), .ZN(n4401) );
  AND2_X1 U5400 ( .A1(n5156), .A2(n4921), .ZN(n4676) );
  NOR2_X1 U5401 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(P1_IR_REG_7__SCAN_IN), .ZN(
        n4826) );
  NOR2_X1 U5402 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_11__SCAN_IN), .ZN(
        n4824) );
  NOR2_X1 U5403 ( .A1(P1_IR_REG_6__SCAN_IN), .A2(P1_IR_REG_10__SCAN_IN), .ZN(
        n4825) );
  NAND2_X1 U5404 ( .A1(n4897), .A2(n4896), .ZN(n5108) );
  XNOR2_X1 U5405 ( .A(n4881), .B(SI_4_), .ZN(n5055) );
  INV_X1 U5406 ( .A(n5041), .ZN(n4877) );
  NAND2_X1 U5407 ( .A1(n4867), .A2(n4866), .ZN(n4869) );
  INV_X1 U5408 ( .A(P1_RD_REG_SCAN_IN), .ZN(n4867) );
  INV_X1 U5409 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n4866) );
  OR2_X1 U5410 ( .A1(n5904), .A2(n5903), .ZN(n5921) );
  NAND2_X1 U5411 ( .A1(n8500), .A2(n8009), .ZN(n4710) );
  AND2_X1 U5412 ( .A1(n5852), .A2(n5838), .ZN(n4713) );
  NAND2_X1 U5413 ( .A1(n5867), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n5886) );
  INV_X1 U5414 ( .A(n5869), .ZN(n5867) );
  OR2_X1 U5415 ( .A1(n6066), .A2(n6065), .ZN(n6084) );
  INV_X1 U5416 ( .A(n7304), .ZN(n4694) );
  NOR2_X1 U5417 ( .A1(n4695), .A2(n4690), .ZN(n4689) );
  INV_X1 U5418 ( .A(n5931), .ZN(n4690) );
  INV_X1 U5419 ( .A(n7305), .ZN(n4695) );
  NAND2_X1 U5420 ( .A1(n8441), .A2(n6096), .ZN(n6112) );
  NOR2_X1 U5421 ( .A1(n7811), .A2(n4720), .ZN(n4719) );
  INV_X1 U5422 ( .A(n6014), .ZN(n4720) );
  INV_X1 U5423 ( .A(n6034), .ZN(n4717) );
  AND2_X1 U5424 ( .A1(n6057), .A2(n6046), .ZN(n8482) );
  INV_X1 U5425 ( .A(n5801), .ZN(n5799) );
  INV_X1 U5426 ( .A(n8502), .ZN(n8491) );
  OR2_X1 U5427 ( .A1(n5968), .A2(n5967), .ZN(n5986) );
  OR2_X1 U5428 ( .A1(n4446), .A2(n6502), .ZN(n4444) );
  INV_X1 U5429 ( .A(n6503), .ZN(n4447) );
  CLKBUF_X1 U5430 ( .A(n5808), .Z(n5809) );
  OAI21_X1 U5431 ( .B1(n9693), .B2(n4442), .A(n4437), .ZN(n9708) );
  AOI21_X1 U5432 ( .B1(n4439), .B2(n4438), .A(n9707), .ZN(n4437) );
  INV_X1 U5433 ( .A(n4440), .ZN(n4438) );
  NAND2_X1 U5434 ( .A1(n9693), .A2(n4440), .ZN(n4443) );
  OR2_X1 U5435 ( .A1(n5859), .A2(P2_IR_REG_7__SCAN_IN), .ZN(n5860) );
  NOR2_X1 U5436 ( .A1(n5860), .A2(P2_IR_REG_8__SCAN_IN), .ZN(n5900) );
  NOR2_X1 U5437 ( .A1(n7150), .A2(n7151), .ZN(n7152) );
  AOI21_X1 U5438 ( .B1(n9742), .B2(n9743), .A(n7613), .ZN(n7616) );
  NAND2_X1 U5439 ( .A1(n7616), .A2(n7615), .ZN(n7614) );
  OR2_X1 U5440 ( .A1(n8585), .A2(n8145), .ZN(n8404) );
  NAND2_X1 U5441 ( .A1(n8368), .A2(n8401), .ZN(n8145) );
  INV_X1 U5442 ( .A(n4648), .ZN(n8587) );
  AND2_X1 U5443 ( .A1(n4649), .A2(n4635), .ZN(n4634) );
  NOR2_X1 U5444 ( .A1(n4636), .A2(n4633), .ZN(n4632) );
  NAND2_X1 U5445 ( .A1(n8595), .A2(n8396), .ZN(n8580) );
  NAND2_X1 U5446 ( .A1(n4480), .A2(n8503), .ZN(n8396) );
  NAND2_X1 U5447 ( .A1(n8580), .A2(n8586), .ZN(n8579) );
  NAND2_X1 U5448 ( .A1(n8401), .A2(n8320), .ZN(n8586) );
  NAND2_X1 U5449 ( .A1(n6614), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n8028) );
  INV_X1 U5450 ( .A(n7999), .ZN(n6614) );
  AOI21_X1 U5451 ( .B1(n4781), .B2(n4782), .A(n8365), .ZN(n4779) );
  NAND2_X1 U5452 ( .A1(n8654), .A2(n4781), .ZN(n4780) );
  INV_X1 U5453 ( .A(n6118), .ZN(n6116) );
  AOI21_X1 U5454 ( .B1(n4619), .B2(n4623), .A(n4618), .ZN(n8141) );
  INV_X1 U5455 ( .A(n4620), .ZN(n4618) );
  NAND2_X1 U5456 ( .A1(n8298), .A2(n8296), .ZN(n8672) );
  NAND2_X1 U5457 ( .A1(n8725), .A2(n8390), .ZN(n8726) );
  AND2_X1 U5458 ( .A1(n8292), .A2(n8290), .ZN(n8709) );
  AND2_X1 U5459 ( .A1(n6091), .A2(n6090), .ZN(n8700) );
  AND2_X1 U5460 ( .A1(n8288), .A2(n8695), .ZN(n8718) );
  AOI21_X1 U5461 ( .B1(n8741), .B2(n8389), .A(n8388), .ZN(n8715) );
  NAND2_X1 U5462 ( .A1(n6000), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n6025) );
  INV_X1 U5463 ( .A(n6002), .ZN(n6000) );
  AND2_X1 U5464 ( .A1(n7660), .A2(n7734), .ZN(n7761) );
  NAND2_X1 U5465 ( .A1(n5985), .A2(n5984), .ZN(n7647) );
  OAI21_X1 U5466 ( .B1(n8356), .B2(n4795), .A(n7600), .ZN(n4794) );
  NOR2_X1 U5467 ( .A1(n7377), .A2(n4487), .ZN(n4486) );
  NAND2_X1 U5468 ( .A1(n4488), .A2(n4489), .ZN(n7675) );
  NOR2_X1 U5469 ( .A1(n7377), .A2(n7599), .ZN(n4488) );
  NAND2_X1 U5470 ( .A1(n5951), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n5968) );
  INV_X1 U5471 ( .A(n5952), .ZN(n5951) );
  AND2_X1 U5472 ( .A1(n8355), .A2(n4596), .ZN(n4594) );
  NAND2_X1 U5473 ( .A1(n7327), .A2(n4597), .ZN(n4595) );
  NAND2_X1 U5474 ( .A1(n4597), .A2(n4599), .ZN(n4596) );
  NAND2_X1 U5475 ( .A1(n7374), .A2(n8241), .ZN(n7441) );
  NOR2_X1 U5476 ( .A1(n4490), .A2(n7377), .ZN(n7434) );
  NOR2_X1 U5477 ( .A1(n7377), .A2(n9818), .ZN(n7433) );
  NAND2_X1 U5478 ( .A1(n7327), .A2(n8234), .ZN(n7374) );
  AND4_X1 U5479 ( .A1(n5927), .A2(n5926), .A3(n5925), .A4(n5924), .ZN(n7442)
         );
  AOI21_X1 U5480 ( .B1(n4608), .B2(n4610), .A(n4607), .ZN(n4606) );
  INV_X1 U5481 ( .A(n4610), .ZN(n4609) );
  INV_X1 U5482 ( .A(n8224), .ZN(n4607) );
  NOR2_X1 U5483 ( .A1(n7282), .A2(n7040), .ZN(n7033) );
  NAND2_X1 U5484 ( .A1(n7299), .A2(n7049), .ZN(n7073) );
  AND4_X1 U5485 ( .A1(n5891), .A2(n5890), .A3(n5889), .A4(n5888), .ZN(n7078)
         );
  NAND2_X1 U5486 ( .A1(n7294), .A2(n7048), .ZN(n7299) );
  OR2_X1 U5487 ( .A1(n7231), .A2(n7314), .ZN(n7286) );
  NAND2_X1 U5488 ( .A1(n8346), .A2(n7238), .ZN(n7037) );
  NAND2_X1 U5489 ( .A1(n8346), .A2(n4592), .ZN(n4591) );
  INV_X1 U5490 ( .A(n8346), .ZN(n7227) );
  AND2_X1 U5491 ( .A1(n8183), .A2(n8185), .ZN(n6637) );
  NAND2_X1 U5492 ( .A1(n8149), .A2(n8148), .ZN(n8765) );
  OR2_X1 U5493 ( .A1(n9777), .A2(n6145), .ZN(n7111) );
  NOR2_X1 U5494 ( .A1(n5715), .A2(P2_IR_REG_28__SCAN_IN), .ZN(n5702) );
  INV_X1 U5495 ( .A(n4605), .ZN(n4603) );
  INV_X1 U5496 ( .A(n5733), .ZN(n6626) );
  INV_X1 U5497 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n4463) );
  NOR2_X1 U5498 ( .A1(n8883), .A2(n4568), .ZN(n4567) );
  INV_X1 U5499 ( .A(n7932), .ZN(n4568) );
  NAND3_X1 U5500 ( .A1(n4572), .A2(n4571), .A3(n7913), .ZN(n8892) );
  NAND2_X1 U5501 ( .A1(n8950), .A2(n8951), .ZN(n4572) );
  OR2_X1 U5502 ( .A1(n5130), .A2(n5129), .ZN(n5146) );
  NOR2_X1 U5503 ( .A1(n4553), .A2(n4554), .ZN(n4552) );
  INV_X1 U5504 ( .A(n7345), .ZN(n4553) );
  INV_X1 U5505 ( .A(n5306), .ZN(n5355) );
  NAND2_X1 U5506 ( .A1(P1_REG3_REG_20__SCAN_IN), .A2(n5355), .ZN(n5354) );
  NAND2_X1 U5507 ( .A1(n4376), .A2(n4375), .ZN(n8950) );
  AND2_X1 U5508 ( .A1(n4581), .A2(n4578), .ZN(n4375) );
  NAND2_X1 U5509 ( .A1(n8944), .A2(n4582), .ZN(n4376) );
  NOR2_X1 U5510 ( .A1(n10003), .A2(n5293), .ZN(n5307) );
  INV_X1 U5511 ( .A(n7904), .ZN(n7942) );
  AND2_X1 U5512 ( .A1(n6864), .A2(n6657), .ZN(n4357) );
  NAND2_X1 U5513 ( .A1(n4355), .A2(n4345), .ZN(n4354) );
  NAND2_X1 U5514 ( .A1(n4356), .A2(n6864), .ZN(n4355) );
  NAND2_X1 U5515 ( .A1(n8892), .A2(n4365), .ZN(n4362) );
  NOR2_X1 U5516 ( .A1(n8935), .A2(n4366), .ZN(n4365) );
  INV_X1 U5517 ( .A(n8893), .ZN(n4366) );
  NAND2_X1 U5518 ( .A1(n8891), .A2(n4367), .ZN(n4361) );
  INV_X1 U5519 ( .A(n8935), .ZN(n4367) );
  NAND2_X1 U5520 ( .A1(n7841), .A2(n7840), .ZN(n8983) );
  AND2_X1 U5521 ( .A1(n7839), .A2(n7838), .ZN(n7840) );
  AND4_X1 U5522 ( .A1(n5191), .A2(n5190), .A3(n5189), .A4(n5188), .ZN(n9425)
         );
  NAND2_X1 U5523 ( .A1(n6265), .A2(n9015), .ZN(n6406) );
  OR2_X1 U5524 ( .A1(n9488), .A2(n9487), .ZN(n4420) );
  OR2_X1 U5525 ( .A1(n5089), .A2(P1_IR_REG_5__SCAN_IN), .ZN(n5180) );
  AND2_X1 U5526 ( .A1(n4418), .A2(n4329), .ZN(n9514) );
  AND2_X1 U5527 ( .A1(n6432), .A2(n9528), .ZN(n9544) );
  NOR2_X1 U5528 ( .A1(n9544), .A2(n9545), .ZN(n9542) );
  NAND2_X1 U5529 ( .A1(n4685), .A2(n5511), .ZN(n5516) );
  NAND2_X1 U5530 ( .A1(n8872), .A2(n5509), .ZN(n4685) );
  NAND2_X1 U5531 ( .A1(n4658), .A2(n5498), .ZN(n9070) );
  NAND2_X1 U5532 ( .A1(n8146), .A2(n5509), .ZN(n4658) );
  AND2_X1 U5533 ( .A1(n8135), .A2(n9077), .ZN(n9069) );
  OR2_X1 U5534 ( .A1(n9289), .A2(n10020), .ZN(n9082) );
  INV_X1 U5535 ( .A(n9075), .ZN(n9085) );
  NOR2_X1 U5536 ( .A1(n9284), .A2(n9094), .ZN(n9077) );
  OR2_X1 U5537 ( .A1(n9108), .A2(n9289), .ZN(n9094) );
  AOI21_X1 U5538 ( .B1(n4521), .B2(n4519), .A(n4518), .ZN(n9112) );
  NOR2_X1 U5539 ( .A1(n4525), .A2(n4520), .ZN(n4519) );
  OAI21_X1 U5540 ( .B1(n4522), .B2(n4520), .A(n8118), .ZN(n4518) );
  OR2_X1 U5541 ( .A1(n4473), .A2(n9294), .ZN(n4472) );
  NOR3_X1 U5542 ( .A1(n9162), .A2(n5402), .A3(n9308), .ZN(n9139) );
  NAND2_X1 U5543 ( .A1(n4847), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n5393) );
  INV_X1 U5544 ( .A(n5391), .ZN(n4847) );
  AOI21_X1 U5545 ( .B1(n4741), .B2(n4740), .A(n4339), .ZN(n4738) );
  NOR2_X1 U5546 ( .A1(n9162), .A2(n9308), .ZN(n9149) );
  NOR2_X1 U5547 ( .A1(n9206), .A2(n9324), .ZN(n9193) );
  AOI21_X1 U5548 ( .B1(n9225), .B2(n8107), .A(n8106), .ZN(n9212) );
  NAND2_X1 U5549 ( .A1(n4288), .A2(n8129), .ZN(n9219) );
  INV_X1 U5550 ( .A(n4500), .ZN(n9241) );
  NAND2_X1 U5551 ( .A1(n9258), .A2(n4507), .ZN(n4503) );
  INV_X1 U5552 ( .A(n4502), .ZN(n4501) );
  NAND2_X1 U5553 ( .A1(n8129), .A2(n4476), .ZN(n9234) );
  AND2_X1 U5554 ( .A1(n9344), .A2(n9243), .ZN(n8080) );
  AND2_X1 U5555 ( .A1(n8129), .A2(n9257), .ZN(n9251) );
  NOR2_X1 U5556 ( .A1(n7719), .A2(n9433), .ZN(n4465) );
  INV_X1 U5557 ( .A(n9413), .ZN(n4464) );
  AOI21_X1 U5558 ( .B1(n7696), .B2(n4303), .A(n4759), .ZN(n8076) );
  NAND2_X1 U5559 ( .A1(n4760), .A2(n4309), .ZN(n4759) );
  OR2_X1 U5560 ( .A1(n5218), .A2(n5217), .ZN(n5220) );
  NOR2_X1 U5561 ( .A1(n5220), .A2(n5202), .ZN(n5245) );
  NAND2_X1 U5562 ( .A1(n4343), .A2(n9414), .ZN(n9394) );
  AND2_X1 U5563 ( .A1(n9414), .A2(n7590), .ZN(n9392) );
  NOR2_X1 U5564 ( .A1(n9413), .A2(n9433), .ZN(n9414) );
  OR2_X1 U5565 ( .A1(n5146), .A2(n7394), .ZN(n5163) );
  OR2_X1 U5566 ( .A1(n7480), .A2(n7571), .ZN(n9413) );
  NAND2_X1 U5567 ( .A1(n7487), .A2(n5155), .ZN(n7579) );
  NOR2_X1 U5568 ( .A1(n5096), .A2(n5095), .ZN(n5117) );
  BUF_X1 U5569 ( .A(n5152), .Z(n7097) );
  INV_X1 U5570 ( .A(n7406), .ZN(n7096) );
  NAND2_X1 U5571 ( .A1(n6982), .A2(n9646), .ZN(n7102) );
  NAND2_X1 U5572 ( .A1(n5081), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n5096) );
  AND3_X1 U5573 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .A3(P1_REG3_REG_5__SCAN_IN), .ZN(n5081) );
  NAND2_X1 U5574 ( .A1(n5541), .A2(n5634), .ZN(n6930) );
  AND2_X1 U5575 ( .A1(n6283), .A2(n4498), .ZN(n4497) );
  OAI22_X1 U5576 ( .A1(n6220), .A2(n4499), .B1(n6221), .B2(n4279), .ZN(n4498)
         );
  INV_X1 U5577 ( .A(n6895), .ZN(n6782) );
  NAND2_X1 U5578 ( .A1(n6782), .A2(n6781), .ZN(n6780) );
  AOI21_X1 U5579 ( .B1(n9169), .B2(n8113), .A(n8112), .ZN(n9154) );
  INV_X1 U5580 ( .A(n9373), .ZN(n4477) );
  NOR3_X2 U5581 ( .A1(n5667), .A2(n4774), .A3(n4835), .ZN(n4839) );
  NAND2_X1 U5582 ( .A1(n4775), .A2(n4836), .ZN(n4774) );
  INV_X1 U5583 ( .A(n4776), .ZN(n4775) );
  XNOR2_X1 U5584 ( .A(n4837), .B(P1_IR_REG_30__SCAN_IN), .ZN(n4842) );
  NAND2_X1 U5585 ( .A1(n9367), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4837) );
  XNOR2_X1 U5586 ( .A(n5500), .B(SI_30_), .ZN(n8146) );
  XNOR2_X1 U5587 ( .A(n5496), .B(n5479), .ZN(n8142) );
  XNOR2_X1 U5588 ( .A(n5476), .B(n5475), .ZN(n8023) );
  XNOR2_X1 U5589 ( .A(n5458), .B(n5457), .ZN(n8010) );
  XNOR2_X1 U5590 ( .A(n5385), .B(n5386), .ZN(n7163) );
  XNOR2_X1 U5591 ( .A(n5332), .B(n5331), .ZN(n6974) );
  NAND2_X1 U5592 ( .A1(n5330), .A2(n5329), .ZN(n5332) );
  XNOR2_X1 U5593 ( .A(n5350), .B(n5349), .ZN(n6972) );
  NAND2_X1 U5594 ( .A1(n5347), .A2(n5346), .ZN(n5350) );
  NAND2_X1 U5595 ( .A1(n4679), .A2(n4677), .ZN(n5209) );
  OR2_X1 U5596 ( .A1(n5141), .A2(P1_IR_REG_9__SCAN_IN), .ZN(n5158) );
  NAND2_X1 U5597 ( .A1(n4384), .A2(n4389), .ZN(n5140) );
  NAND2_X1 U5598 ( .A1(n4394), .A2(n4388), .ZN(n4384) );
  OR2_X1 U5599 ( .A1(n5113), .A2(P1_IR_REG_8__SCAN_IN), .ZN(n5141) );
  XNOR2_X1 U5600 ( .A(n5125), .B(n4816), .ZN(n6245) );
  NAND2_X1 U5601 ( .A1(n4392), .A2(n4897), .ZN(n5125) );
  OR2_X1 U5602 ( .A1(n5109), .A2(n5108), .ZN(n4392) );
  NAND2_X1 U5603 ( .A1(n5088), .A2(n4888), .ZN(n4661) );
  NAND2_X1 U5604 ( .A1(n6115), .A2(n6114), .ZN(n8799) );
  NAND2_X1 U5605 ( .A1(n7980), .A2(n5766), .ZN(n6208) );
  NAND2_X1 U5606 ( .A1(n5932), .A2(n5931), .ZN(n7306) );
  NAND2_X1 U5607 ( .A1(n5999), .A2(n5998), .ZN(n7791) );
  NAND2_X1 U5608 ( .A1(n7782), .A2(n6014), .ZN(n7812) );
  NAND2_X1 U5609 ( .A1(n6205), .A2(n5795), .ZN(n6846) );
  AND3_X1 U5610 ( .A1(n6056), .A2(n6055), .A3(n6054), .ZN(n8701) );
  AND2_X1 U5611 ( .A1(n6078), .A2(n6062), .ZN(n4714) );
  NAND2_X1 U5612 ( .A1(n8426), .A2(n6062), .ZN(n8466) );
  AND4_X1 U5613 ( .A1(n5943), .A2(n5942), .A3(n5941), .A4(n5940), .ZN(n7453)
         );
  NAND2_X1 U5614 ( .A1(n4691), .A2(n7305), .ZN(n7450) );
  NAND2_X1 U5615 ( .A1(n7306), .A2(n7304), .ZN(n4691) );
  OR2_X1 U5616 ( .A1(n7960), .A2(n8721), .ZN(n8502) );
  INV_X1 U5617 ( .A(n8504), .ZN(n8493) );
  INV_X1 U5618 ( .A(n8509), .ZN(n8499) );
  NAND2_X1 U5619 ( .A1(n4822), .A2(n8377), .ZN(n8378) );
  NAND2_X1 U5620 ( .A1(n5923), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n5708) );
  AND2_X1 U5621 ( .A1(n5705), .A2(n5704), .ZN(n5710) );
  NAND2_X1 U5622 ( .A1(n4445), .A2(n6501), .ZN(n6545) );
  NAND2_X1 U5623 ( .A1(n4443), .A2(n4444), .ZN(n6523) );
  INV_X1 U5624 ( .A(n4453), .ZN(n6553) );
  INV_X1 U5625 ( .A(n4455), .ZN(n6530) );
  NAND2_X1 U5626 ( .A1(n4453), .A2(n4336), .ZN(n6610) );
  NOR2_X1 U5627 ( .A1(n6703), .A2(n6558), .ZN(n6590) );
  NAND2_X1 U5628 ( .A1(n6590), .A2(n4449), .ZN(n6588) );
  NOR2_X1 U5629 ( .A1(n4451), .A2(n4450), .ZN(n4449) );
  NOR2_X1 U5630 ( .A1(n6586), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n4450) );
  INV_X1 U5631 ( .A(n6559), .ZN(n4451) );
  NOR2_X1 U5632 ( .A1(n6667), .A2(n4452), .ZN(n6671) );
  NOR2_X1 U5633 ( .A1(n6575), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n4452) );
  NOR2_X1 U5634 ( .A1(n6671), .A2(n6670), .ZN(n7150) );
  AND2_X1 U5635 ( .A1(n6257), .A2(n6256), .ZN(n8068) );
  NAND2_X1 U5636 ( .A1(n6015), .A2(n6017), .ZN(n6035) );
  AND2_X1 U5637 ( .A1(n6496), .A2(n6183), .ZN(n9747) );
  NAND2_X1 U5638 ( .A1(n8160), .A2(n8159), .ZN(n8762) );
  NAND2_X1 U5639 ( .A1(n4647), .A2(n4645), .ZN(n8602) );
  INV_X1 U5640 ( .A(n4646), .ZN(n4645) );
  NOR2_X1 U5641 ( .A1(n4639), .A2(n4638), .ZN(n8612) );
  INV_X1 U5642 ( .A(n4652), .ZN(n4639) );
  NAND2_X1 U5643 ( .A1(n7997), .A2(n7996), .ZN(n8785) );
  NAND2_X1 U5644 ( .A1(n7993), .A2(n7992), .ZN(n8790) );
  NAND2_X1 U5645 ( .A1(n4640), .A2(n4653), .ZN(n8630) );
  OR2_X1 U5646 ( .A1(n8642), .A2(n8641), .ZN(n4640) );
  NAND2_X1 U5647 ( .A1(n8652), .A2(n4784), .ZN(n8640) );
  NAND2_X1 U5648 ( .A1(n4625), .A2(n8292), .ZN(n8683) );
  INV_X1 U5649 ( .A(n4802), .ZN(n8682) );
  NOR2_X1 U5650 ( .A1(n8710), .A2(n8709), .ZN(n8816) );
  NAND2_X1 U5651 ( .A1(n4789), .A2(n7751), .ZN(n7752) );
  NAND2_X1 U5652 ( .A1(n7681), .A2(n8257), .ZN(n7655) );
  NAND2_X1 U5653 ( .A1(n4797), .A2(n7600), .ZN(n7672) );
  NAND2_X1 U5654 ( .A1(n7429), .A2(n7326), .ZN(n7601) );
  NAND2_X1 U5655 ( .A1(n7356), .A2(n7070), .ZN(n7071) );
  NAND2_X1 U5656 ( .A1(n7216), .A2(n8189), .ZN(n6768) );
  OR2_X1 U5657 ( .A1(n5753), .A2(n5737), .ZN(n5738) );
  INV_X1 U5658 ( .A(n9837), .ZN(n9836) );
  INV_X1 U5659 ( .A(n4631), .ZN(n8772) );
  XNOR2_X1 U5660 ( .A(n6138), .B(n6137), .ZN(n7199) );
  INV_X1 U5661 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n6217) );
  XNOR2_X1 U5662 ( .A(n4461), .B(n4460), .ZN(n8548) );
  INV_X1 U5663 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n4460) );
  NOR2_X1 U5664 ( .A1(n5754), .A2(n8873), .ZN(n4461) );
  NAND2_X1 U5665 ( .A1(n6655), .A2(n6654), .ZN(n6656) );
  AND3_X1 U5666 ( .A1(n5049), .A2(n5048), .A3(n5047), .ZN(n9618) );
  NAND2_X1 U5667 ( .A1(n6656), .A2(n6657), .ZN(n6720) );
  INV_X1 U5668 ( .A(n4545), .ZN(n4544) );
  NAND2_X1 U5669 ( .A1(n8926), .A2(n4541), .ZN(n4353) );
  OAI21_X1 U5670 ( .B1(n7875), .B2(n4548), .A(n4546), .ZN(n4545) );
  OAI21_X1 U5671 ( .B1(n8944), .B2(n7894), .A(n7893), .ZN(n8908) );
  NAND2_X1 U5672 ( .A1(n7633), .A2(n7634), .ZN(n7638) );
  NAND2_X1 U5673 ( .A1(n4990), .A2(n4989), .ZN(n9299) );
  AND3_X1 U5674 ( .A1(n5077), .A2(n5076), .A3(n5075), .ZN(n9633) );
  OR2_X1 U5675 ( .A1(n5027), .A2(n6225), .ZN(n5077) );
  AND2_X1 U5676 ( .A1(n4364), .A2(n4363), .ZN(n8934) );
  NAND2_X1 U5677 ( .A1(n8892), .A2(n8893), .ZN(n4363) );
  NAND2_X1 U5678 ( .A1(n6720), .A2(n6719), .ZN(n6865) );
  NAND2_X1 U5679 ( .A1(n5319), .A2(n5318), .ZN(n9314) );
  NAND2_X1 U5680 ( .A1(n4373), .A2(n4555), .ZN(n7550) );
  AND2_X1 U5681 ( .A1(n7470), .A2(n4556), .ZN(n4555) );
  NAND3_X1 U5682 ( .A1(n5033), .A2(n5032), .A3(n5031), .ZN(n6937) );
  NAND2_X1 U5683 ( .A1(n4550), .A2(n8923), .ZN(n4543) );
  NAND2_X1 U5684 ( .A1(n5291), .A2(n5290), .ZN(n9334) );
  INV_X1 U5685 ( .A(n8963), .ZN(n8994) );
  NOR2_X1 U5686 ( .A1(n5624), .A2(n5664), .ZN(n4656) );
  NOR2_X1 U5687 ( .A1(n5671), .A2(n5670), .ZN(n5672) );
  AND2_X1 U5688 ( .A1(n5665), .A2(n5664), .ZN(n5671) );
  XNOR2_X1 U5689 ( .A(n4861), .B(P1_IR_REG_22__SCAN_IN), .ZN(n6387) );
  OR2_X1 U5690 ( .A1(n5466), .A2(n6920), .ZN(n5051) );
  OR2_X1 U5691 ( .A1(n5035), .A2(n6468), .ZN(n5024) );
  OR2_X1 U5692 ( .A1(n5119), .A2(n6287), .ZN(n5023) );
  OR2_X1 U5693 ( .A1(n5035), .A2(n6796), .ZN(n5003) );
  OR2_X1 U5694 ( .A1(n5119), .A2(n6288), .ZN(n5000) );
  OR2_X1 U5695 ( .A1(n5119), .A2(n9473), .ZN(n5011) );
  XNOR2_X1 U5696 ( .A(n6289), .B(n6264), .ZN(n9017) );
  NAND2_X1 U5697 ( .A1(n9017), .A2(n9016), .ZN(n9015) );
  NOR2_X1 U5698 ( .A1(n5061), .A2(n5060), .ZN(n9484) );
  AND2_X1 U5699 ( .A1(n4420), .A2(n4419), .ZN(n9503) );
  NOR2_X1 U5700 ( .A1(n6430), .A2(n4335), .ZN(n9530) );
  NAND2_X1 U5701 ( .A1(n9530), .A2(n9529), .ZN(n9528) );
  NAND2_X1 U5702 ( .A1(n6435), .A2(n9558), .ZN(n9557) );
  AND2_X1 U5703 ( .A1(n4410), .A2(n4409), .ZN(n6698) );
  NOR2_X1 U5704 ( .A1(n7727), .A2(n4429), .ZN(n7730) );
  AND2_X1 U5705 ( .A1(n7728), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n4429) );
  INV_X1 U5706 ( .A(n4428), .ZN(n9038) );
  INV_X1 U5707 ( .A(n4426), .ZN(n9043) );
  INV_X1 U5708 ( .A(n5516), .ZN(n9270) );
  INV_X1 U5709 ( .A(n9070), .ZN(n9276) );
  XNOR2_X1 U5710 ( .A(n8099), .B(n8098), .ZN(n9283) );
  INV_X1 U5711 ( .A(n8128), .ZN(n9282) );
  XNOR2_X1 U5712 ( .A(n4496), .B(n8098), .ZN(n8127) );
  AOI21_X1 U5713 ( .B1(n9107), .B2(n8096), .A(n8095), .ZN(n9093) );
  AND2_X1 U5714 ( .A1(n5417), .A2(n5416), .ZN(n9111) );
  OAI21_X1 U5715 ( .B1(n9169), .B2(n4525), .A(n4522), .ZN(n9127) );
  INV_X1 U5716 ( .A(n9299), .ZN(n9125) );
  NAND2_X1 U5717 ( .A1(n4528), .A2(n4529), .ZN(n9136) );
  INV_X1 U5718 ( .A(n4736), .ZN(n9147) );
  AOI21_X1 U5719 ( .B1(n4743), .B2(n4737), .A(n4739), .ZN(n4736) );
  INV_X1 U5720 ( .A(n4741), .ZN(n4737) );
  NAND2_X1 U5721 ( .A1(n4743), .A2(n4742), .ZN(n9161) );
  NAND2_X1 U5722 ( .A1(n8086), .A2(n4811), .ZN(n9177) );
  OAI21_X1 U5723 ( .B1(n9398), .B2(n4506), .A(n4504), .ZN(n9259) );
  NAND2_X1 U5724 ( .A1(n4509), .A2(n7799), .ZN(n8102) );
  NAND2_X1 U5725 ( .A1(n9398), .A2(n4294), .ZN(n4509) );
  NAND2_X1 U5726 ( .A1(n4758), .A2(n4762), .ZN(n7796) );
  NAND2_X1 U5727 ( .A1(n7696), .A2(n4292), .ZN(n4758) );
  AND2_X1 U5728 ( .A1(n7696), .A2(n7695), .ZN(n9391) );
  NAND2_X1 U5729 ( .A1(n5183), .A2(n5182), .ZN(n7694) );
  NAND2_X1 U5730 ( .A1(n7573), .A2(n7572), .ZN(n9412) );
  AND2_X1 U5731 ( .A1(n7418), .A2(n7417), .ZN(n7421) );
  AND2_X1 U5732 ( .A1(n5124), .A2(n5563), .ZN(n4804) );
  INV_X1 U5733 ( .A(n7176), .ZN(n7405) );
  NAND2_X1 U5734 ( .A1(n6951), .A2(n5574), .ZN(n6978) );
  NAND2_X1 U5735 ( .A1(n9593), .A2(n6948), .ZN(n6950) );
  INV_X1 U5736 ( .A(n9639), .ZN(n7026) );
  INV_X1 U5737 ( .A(n6947), .ZN(n9595) );
  NAND2_X1 U5738 ( .A1(n6914), .A2(n6913), .ZN(n6944) );
  INV_X1 U5739 ( .A(n9627), .ZN(n6945) );
  INV_X1 U5740 ( .A(n6794), .ZN(n6778) );
  INV_X1 U5741 ( .A(n9256), .ZN(n9434) );
  AND2_X1 U5742 ( .A1(n9600), .A2(n6762), .ZN(n9417) );
  NAND2_X1 U5743 ( .A1(n9282), .A2(n4534), .ZN(n9352) );
  NOR2_X1 U5744 ( .A1(n9280), .A2(n4535), .ZN(n4534) );
  OAI21_X1 U5745 ( .B1(n9283), .B2(n9374), .A(n4536), .ZN(n4535) );
  NAND2_X1 U5746 ( .A1(n9281), .A2(n9345), .ZN(n4536) );
  AND2_X1 U5747 ( .A1(n6357), .A2(n5681), .ZN(n9602) );
  INV_X1 U5748 ( .A(n4852), .ZN(n8071) );
  XNOR2_X1 U5749 ( .A(n4985), .B(n4836), .ZN(n5682) );
  OR2_X1 U5750 ( .A1(n4984), .A2(n4838), .ZN(n4985) );
  NAND2_X1 U5751 ( .A1(n5673), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5675) );
  XNOR2_X1 U5752 ( .A(n5365), .B(n5364), .ZN(n7060) );
  INV_X1 U5753 ( .A(n6387), .ZN(n7004) );
  NAND2_X1 U5754 ( .A1(n5527), .A2(n5526), .ZN(n6976) );
  OAI21_X1 U5755 ( .B1(n4858), .B2(P1_IR_REG_20__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5525) );
  INV_X1 U5756 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n9901) );
  NAND2_X1 U5757 ( .A1(n7955), .A2(n5838), .ZN(n6683) );
  NAND2_X1 U5758 ( .A1(n4700), .A2(n8473), .ZN(n4698) );
  NAND2_X1 U5759 ( .A1(n4712), .A2(n5880), .ZN(n6996) );
  OAI21_X1 U5760 ( .B1(n8067), .B2(n4282), .A(n4456), .ZN(P2_U3264) );
  AOI21_X1 U5761 ( .B1(n4458), .B2(n4282), .A(n4457), .ZN(n4456) );
  NAND2_X1 U5762 ( .A1(n4630), .A2(n4627), .ZN(P2_U3267) );
  NAND2_X1 U5763 ( .A1(n4631), .A2(n8734), .ZN(n4630) );
  OAI21_X1 U5764 ( .B1(n8773), .B2(n8761), .A(n4629), .ZN(n4628) );
  NOR2_X1 U5765 ( .A1(n8777), .A2(n9772), .ZN(n8592) );
  NAND2_X1 U5766 ( .A1(n4562), .A2(n8973), .ZN(n4560) );
  OAI21_X1 U5767 ( .B1(n9062), .B2(n9592), .A(n4421), .ZN(P1_U3260) );
  AOI21_X1 U5768 ( .B1(n4423), .B2(n9592), .A(n4422), .ZN(n4421) );
  OAI21_X1 U5769 ( .B1(n9571), .B2(n4868), .A(n9063), .ZN(n4422) );
  INV_X1 U5770 ( .A(n4468), .ZN(n9350) );
  NAND2_X1 U5771 ( .A1(n4533), .A2(n4532), .ZN(P1_U3552) );
  OR2_X1 U5772 ( .A1(n9678), .A2(n4853), .ZN(n4532) );
  NAND2_X1 U5773 ( .A1(n9352), .A2(n9678), .ZN(n4533) );
  NAND2_X1 U5774 ( .A1(n9666), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n4467) );
  AND2_X1 U5775 ( .A1(n4484), .A2(n8692), .ZN(n4285) );
  XOR2_X1 U5776 ( .A(n7945), .B(n7944), .Z(n4286) );
  NAND2_X1 U5777 ( .A1(n6357), .A2(n6388), .ZN(n6384) );
  AND2_X1 U5778 ( .A1(n9151), .A2(n9172), .ZN(n8115) );
  AND2_X1 U5779 ( .A1(n4807), .A2(n4312), .ZN(n4287) );
  AND2_X1 U5780 ( .A1(n4476), .A2(n4475), .ZN(n4288) );
  INV_X1 U5781 ( .A(n8119), .ZN(n4520) );
  NAND2_X1 U5782 ( .A1(n4543), .A2(n7877), .ZN(n8959) );
  NAND2_X1 U5783 ( .A1(n8282), .A2(n8176), .ZN(n8653) );
  NAND2_X1 U5784 ( .A1(n4654), .A2(n8663), .ZN(n4653) );
  INV_X1 U5785 ( .A(n4653), .ZN(n4643) );
  NAND2_X1 U5786 ( .A1(n5276), .A2(n5275), .ZN(n9339) );
  INV_X1 U5787 ( .A(n8692), .ZN(n8810) );
  OR2_X1 U5788 ( .A1(n4819), .A2(n4967), .ZN(n4289) );
  NAND2_X1 U5789 ( .A1(n9126), .A2(n5399), .ZN(n4290) );
  AND2_X1 U5790 ( .A1(n4591), .A2(n8210), .ZN(n4291) );
  NAND2_X1 U5791 ( .A1(n7392), .A2(n7393), .ZN(n7471) );
  NAND2_X1 U5792 ( .A1(n8025), .A2(n8024), .ZN(n8775) );
  INV_X1 U5793 ( .A(n8775), .ZN(n4481) );
  NAND2_X1 U5794 ( .A1(n8086), .A2(n4744), .ZN(n4743) );
  AND2_X2 U5795 ( .A1(n5753), .A2(n4279), .ZN(n5819) );
  CLKBUF_X3 U5796 ( .A(n5819), .Z(n8147) );
  NAND4_X1 U5797 ( .A1(n5012), .A2(n5011), .A3(n5010), .A4(n5009), .ZN(n6360)
         );
  NAND4_X1 U5798 ( .A1(n5024), .A2(n5023), .A3(n5022), .A4(n5021), .ZN(n6448)
         );
  NAND2_X1 U5799 ( .A1(n5388), .A2(n5387), .ZN(n5402) );
  OR2_X1 U5800 ( .A1(n4765), .A2(n4763), .ZN(n4292) );
  AND2_X1 U5801 ( .A1(n5029), .A2(n6289), .ZN(n4293) );
  AND2_X1 U5802 ( .A1(n7798), .A2(n7797), .ZN(n4294) );
  NAND2_X1 U5803 ( .A1(n9125), .A2(n8977), .ZN(n4295) );
  OR2_X1 U5804 ( .A1(n8790), .A2(n8644), .ZN(n8173) );
  NAND2_X1 U5805 ( .A1(n5722), .A2(n4721), .ZN(n4296) );
  INV_X1 U5806 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n4838) );
  AND2_X1 U5807 ( .A1(n7420), .A2(n7417), .ZN(n4297) );
  AND2_X1 U5808 ( .A1(n4295), .A2(n8093), .ZN(n4298) );
  NAND2_X1 U5809 ( .A1(n5707), .A2(n5706), .ZN(n6169) );
  NAND2_X1 U5810 ( .A1(n5216), .A2(n5215), .ZN(n9408) );
  INV_X1 U5811 ( .A(n9408), .ZN(n4767) );
  OR2_X1 U5812 ( .A1(n7706), .A2(n7705), .ZN(n4299) );
  INV_X1 U5813 ( .A(n8114), .ZN(n4530) );
  INV_X1 U5814 ( .A(n4279), .ZN(n4499) );
  OR3_X1 U5815 ( .A1(P2_IR_REG_2__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .A3(
        P2_IR_REG_0__SCAN_IN), .ZN(n4300) );
  AND2_X1 U5816 ( .A1(n4625), .A2(n4623), .ZN(n4301) );
  AND2_X1 U5817 ( .A1(n4574), .A2(n4577), .ZN(n4302) );
  AND2_X1 U5818 ( .A1(n7795), .A2(n4292), .ZN(n4303) );
  NAND2_X1 U5819 ( .A1(n5367), .A2(n5366), .ZN(n9308) );
  INV_X1 U5820 ( .A(n9308), .ZN(n9151) );
  NAND2_X1 U5821 ( .A1(n6099), .A2(n6098), .ZN(n8806) );
  INV_X1 U5822 ( .A(n8806), .ZN(n4483) );
  AND2_X1 U5823 ( .A1(n9314), .A2(n9187), .ZN(n4304) );
  OR2_X1 U5824 ( .A1(n5496), .A2(n5495), .ZN(n4305) );
  NAND2_X1 U5825 ( .A1(n8971), .A2(n8974), .ZN(n8972) );
  OR2_X1 U5826 ( .A1(n5529), .A2(n7004), .ZN(n4306) );
  OR2_X1 U5827 ( .A1(n6453), .A2(n6452), .ZN(n4307) );
  NAND2_X1 U5828 ( .A1(n4790), .A2(n5754), .ZN(n5782) );
  AND2_X1 U5829 ( .A1(n4755), .A2(n4298), .ZN(n4308) );
  NAND2_X1 U5830 ( .A1(n5445), .A2(n5444), .ZN(n9289) );
  OR2_X1 U5831 ( .A1(n7719), .A2(n7794), .ZN(n4309) );
  NAND2_X1 U5832 ( .A1(n5258), .A2(n5257), .ZN(n9344) );
  INV_X1 U5833 ( .A(n8356), .ZN(n7329) );
  AND2_X1 U5834 ( .A1(n8251), .A2(n8250), .ZN(n8356) );
  INV_X1 U5835 ( .A(n4507), .ZN(n4506) );
  NOR2_X1 U5836 ( .A1(n8101), .A2(n4508), .ZN(n4507) );
  AND2_X1 U5837 ( .A1(n6049), .A2(n6048), .ZN(n8390) );
  INV_X1 U5838 ( .A(n8390), .ZN(n8823) );
  AND2_X1 U5839 ( .A1(n9085), .A2(n9082), .ZN(n4310) );
  INV_X1 U5840 ( .A(n4785), .ZN(n4784) );
  INV_X1 U5841 ( .A(n4478), .ZN(n8598) );
  NOR2_X1 U5842 ( .A1(n8617), .A2(n8779), .ZN(n4478) );
  AND2_X1 U5843 ( .A1(n4752), .A2(n4750), .ZN(n4311) );
  AND2_X1 U5844 ( .A1(n4832), .A2(n4768), .ZN(n4312) );
  NAND2_X1 U5845 ( .A1(n8173), .A2(n8171), .ZN(n8629) );
  INV_X1 U5846 ( .A(n8629), .ZN(n8365) );
  AND2_X1 U5847 ( .A1(n8346), .A2(n8189), .ZN(n4313) );
  NAND2_X1 U5848 ( .A1(n5305), .A2(n5304), .ZN(n9329) );
  INV_X1 U5849 ( .A(n9329), .ZN(n4474) );
  AND2_X1 U5850 ( .A1(n8310), .A2(n4651), .ZN(n4314) );
  INV_X1 U5851 ( .A(n8088), .ZN(n4747) );
  INV_X1 U5852 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n4724) );
  OR2_X1 U5853 ( .A1(n8834), .A2(n8754), .ZN(n4315) );
  AND2_X1 U5854 ( .A1(n4892), .A2(SI_7_), .ZN(n4316) );
  NOR2_X1 U5855 ( .A1(n8796), .A2(n8663), .ZN(n4317) );
  OR2_X1 U5856 ( .A1(n5667), .A2(P1_IR_REG_23__SCAN_IN), .ZN(n4318) );
  OR2_X1 U5857 ( .A1(n9299), .A2(n8977), .ZN(n8118) );
  INV_X1 U5858 ( .A(n4442), .ZN(n4439) );
  NAND2_X1 U5859 ( .A1(n4444), .A2(n4338), .ZN(n4442) );
  OAI21_X1 U5860 ( .B1(n4677), .B2(n4675), .A(n5210), .ZN(n4674) );
  NAND2_X1 U5861 ( .A1(n7415), .A2(n7414), .ZN(n4319) );
  AND2_X2 U5862 ( .A1(n9279), .A2(n6388), .ZN(n7936) );
  AND2_X1 U5863 ( .A1(n4786), .A2(n4315), .ZN(n4320) );
  AND2_X1 U5864 ( .A1(n6017), .A2(n4724), .ZN(n4321) );
  INV_X1 U5865 ( .A(n8891), .ZN(n4364) );
  INV_X1 U5866 ( .A(n4389), .ZN(n4387) );
  AOI21_X1 U5867 ( .B1(n4816), .B2(n4391), .A(n4390), .ZN(n4389) );
  AND2_X1 U5868 ( .A1(n5819), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n4322) );
  AND2_X1 U5869 ( .A1(n9092), .A2(n5455), .ZN(n4323) );
  INV_X1 U5870 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n8873) );
  INV_X1 U5871 ( .A(n7189), .ZN(n4554) );
  INV_X1 U5872 ( .A(n6502), .ZN(n4448) );
  AND2_X1 U5873 ( .A1(n4285), .A2(n4483), .ZN(n4324) );
  NAND2_X1 U5874 ( .A1(n4286), .A2(n4567), .ZN(n4325) );
  INV_X1 U5875 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n4495) );
  NAND2_X1 U5876 ( .A1(n4706), .A2(n4704), .ZN(n4326) );
  NAND2_X1 U5877 ( .A1(n6131), .A2(n6130), .ZN(n8796) );
  INV_X1 U5878 ( .A(n8796), .ZN(n4654) );
  OR2_X1 U5879 ( .A1(n5410), .A2(n4670), .ZN(n4327) );
  NAND2_X1 U5880 ( .A1(n8486), .A2(n6058), .ZN(n8426) );
  NAND2_X1 U5881 ( .A1(n8326), .A2(n8327), .ZN(n8402) );
  NAND2_X1 U5882 ( .A1(n7782), .A2(n4719), .ZN(n7813) );
  AND2_X1 U5883 ( .A1(n8019), .A2(n8018), .ZN(n8503) );
  AND2_X1 U5884 ( .A1(n5811), .A2(n5810), .ZN(n6524) );
  INV_X1 U5885 ( .A(n5599), .ZN(n4516) );
  NAND2_X1 U5886 ( .A1(n7926), .A2(n7925), .ZN(n4328) );
  INV_X1 U5887 ( .A(n7909), .ZN(n4578) );
  OR2_X1 U5888 ( .A1(n9500), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n4329) );
  AND2_X1 U5889 ( .A1(n9558), .A2(n4408), .ZN(n4330) );
  NAND2_X1 U5890 ( .A1(n7638), .A2(n7635), .ZN(n7707) );
  NAND2_X1 U5891 ( .A1(n4353), .A2(n4544), .ZN(n8900) );
  NOR2_X1 U5892 ( .A1(n5614), .A2(n5654), .ZN(n8123) );
  INV_X1 U5893 ( .A(n8882), .ZN(n4566) );
  INV_X1 U5894 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n4860) );
  OR2_X1 U5895 ( .A1(n4604), .A2(n4605), .ZN(n4331) );
  OR2_X1 U5896 ( .A1(n5273), .A2(P1_IR_REG_17__SCAN_IN), .ZN(n4332) );
  AND2_X1 U5897 ( .A1(n7903), .A2(n7902), .ZN(n4333) );
  INV_X1 U5898 ( .A(n5287), .ZN(n4945) );
  NAND2_X1 U5899 ( .A1(n8012), .A2(n8011), .ZN(n8779) );
  INV_X1 U5900 ( .A(n8779), .ZN(n4480) );
  NOR2_X1 U5901 ( .A1(n8743), .A2(n8827), .ZN(n8725) );
  NAND2_X1 U5902 ( .A1(n4831), .A2(n4807), .ZN(n5273) );
  NAND2_X1 U5903 ( .A1(n4550), .A2(n7875), .ZN(n8958) );
  OR2_X1 U5904 ( .A1(n4286), .A2(n4566), .ZN(n4334) );
  NOR3_X1 U5905 ( .A1(n9162), .A2(n4472), .A3(n5402), .ZN(n4470) );
  NAND2_X1 U5906 ( .A1(n8144), .A2(n8143), .ZN(n8770) );
  INV_X1 U5907 ( .A(n4471), .ZN(n9120) );
  NOR3_X1 U5908 ( .A1(n9162), .A2(n5402), .A3(n4473), .ZN(n4471) );
  NAND2_X1 U5909 ( .A1(n8725), .A2(n4484), .ZN(n4485) );
  AND2_X1 U5910 ( .A1(n6431), .A2(n7101), .ZN(n4335) );
  OR2_X1 U5911 ( .A1(n6554), .A2(n6528), .ZN(n4336) );
  AND2_X1 U5912 ( .A1(n8951), .A2(n4573), .ZN(n4337) );
  OR2_X1 U5913 ( .A1(n6510), .A2(n7236), .ZN(n4338) );
  NOR2_X1 U5914 ( .A1(n9308), .A2(n9172), .ZN(n4339) );
  AND3_X1 U5915 ( .A1(n4826), .A2(n4825), .A3(n4824), .ZN(n5178) );
  AND2_X1 U5916 ( .A1(n8022), .A2(n8021), .ZN(n4340) );
  INV_X1 U5917 ( .A(n8095), .ZN(n4757) );
  AND2_X1 U5918 ( .A1(n9294), .A2(n9128), .ZN(n8095) );
  INV_X1 U5919 ( .A(n4709), .ZN(n4708) );
  AND2_X1 U5920 ( .A1(n4710), .A2(n8413), .ZN(n4709) );
  AND2_X1 U5921 ( .A1(n4328), .A2(n4368), .ZN(n4341) );
  INV_X1 U5922 ( .A(n8511), .ZN(n8473) );
  AOI21_X1 U5923 ( .B1(n6656), .B2(n4357), .A(n4354), .ZN(n6961) );
  NAND2_X1 U5924 ( .A1(n5966), .A2(n5965), .ZN(n8843) );
  INV_X1 U5925 ( .A(n8843), .ZN(n4491) );
  NAND2_X1 U5926 ( .A1(n5201), .A2(n5200), .ZN(n7719) );
  INV_X1 U5927 ( .A(n7719), .ZN(n4466) );
  NAND2_X1 U5928 ( .A1(n4730), .A2(n4729), .ZN(n7479) );
  INV_X1 U5929 ( .A(n9334), .ZN(n4475) );
  INV_X1 U5930 ( .A(n9578), .ZN(n4513) );
  NAND2_X1 U5931 ( .A1(n4552), .A2(n7341), .ZN(n7391) );
  NAND2_X1 U5932 ( .A1(n5950), .A2(n5949), .ZN(n7599) );
  AND2_X1 U5933 ( .A1(n5478), .A2(n9900), .ZN(n4342) );
  AND2_X1 U5934 ( .A1(n4767), .A2(n7590), .ZN(n4343) );
  NOR3_X1 U5935 ( .A1(n6388), .A2(n9592), .A3(n7004), .ZN(n4344) );
  INV_X1 U5936 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n4777) );
  NAND2_X1 U5937 ( .A1(n6363), .A2(n6362), .ZN(n6390) );
  NAND2_X1 U5938 ( .A1(n6725), .A2(n6724), .ZN(n4345) );
  NAND2_X1 U5939 ( .A1(n4443), .A2(n4439), .ZN(n4346) );
  INV_X1 U5940 ( .A(n9707), .ZN(n4441) );
  INV_X1 U5941 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n4462) );
  INV_X1 U5942 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n4436) );
  NAND2_X1 U5943 ( .A1(n4374), .A2(n9141), .ZN(n9279) );
  INV_X1 U5944 ( .A(P2_U3966), .ZN(n8531) );
  NAND2_X2 U5945 ( .A1(n6784), .A2(n6783), .ZN(n9427) );
  NAND3_X1 U5946 ( .A1(n5430), .A2(n5428), .A3(n5429), .ZN(n5433) );
  NAND2_X1 U5947 ( .A1(n4348), .A2(n4347), .ZN(n5302) );
  NAND2_X1 U5948 ( .A1(n5270), .A2(n5269), .ZN(n4348) );
  MUX2_X1 U5949 ( .A(n5384), .B(n5383), .S(n5483), .Z(n5408) );
  OAI21_X1 U5950 ( .B1(n5514), .B2(n4431), .A(n4430), .ZN(n5499) );
  NAND2_X1 U5951 ( .A1(n5456), .A2(n4323), .ZN(n4432) );
  AOI21_X1 U5952 ( .B1(n5381), .B2(n8111), .A(n5380), .ZN(n5382) );
  XNOR2_X1 U5953 ( .A(n4872), .B(SI_1_), .ZN(n5005) );
  NAND2_X1 U5954 ( .A1(n5079), .A2(n9580), .ZN(n9578) );
  NAND2_X1 U5955 ( .A1(n4350), .A2(n5686), .ZN(P1_U3240) );
  NAND2_X1 U5956 ( .A1(n4399), .A2(n5672), .ZN(n4350) );
  NAND2_X1 U5957 ( .A1(n5176), .A2(n4351), .ZN(n5230) );
  NAND2_X1 U5958 ( .A1(n5377), .A2(n4352), .ZN(n5378) );
  INV_X1 U5959 ( .A(n5055), .ZN(n4880) );
  NAND2_X1 U5960 ( .A1(n7770), .A2(n7769), .ZN(n7774) );
  NAND2_X1 U5961 ( .A1(n4661), .A2(n4890), .ZN(n5105) );
  NAND2_X1 U5962 ( .A1(n4377), .A2(n4879), .ZN(n5056) );
  NAND2_X1 U5963 ( .A1(n4688), .A2(n4692), .ZN(n7449) );
  NAND3_X1 U5964 ( .A1(n4362), .A2(n4361), .A3(n4368), .ZN(n8916) );
  NAND3_X1 U5965 ( .A1(n4361), .A2(n4362), .A3(n4341), .ZN(n4360) );
  OR2_X1 U5966 ( .A1(n7919), .A2(n7918), .ZN(n4368) );
  INV_X1 U5967 ( .A(n4369), .ZN(n5527) );
  INV_X1 U5968 ( .A(n4831), .ZN(n5195) );
  NAND2_X1 U5969 ( .A1(n4287), .A2(n4831), .ZN(n4372) );
  AND3_X2 U5970 ( .A1(n5178), .A2(n4827), .A3(n5059), .ZN(n4831) );
  NAND3_X1 U5971 ( .A1(n7341), .A2(n7345), .A3(n4551), .ZN(n4373) );
  NAND2_X1 U5972 ( .A1(n5042), .A2(n4877), .ZN(n4377) );
  NAND2_X1 U5973 ( .A1(n4874), .A2(n5025), .ZN(n4378) );
  INV_X1 U5974 ( .A(n5157), .ZN(n4382) );
  INV_X1 U5975 ( .A(n5109), .ZN(n4394) );
  NAND2_X1 U5976 ( .A1(n5109), .A2(n4389), .ZN(n4383) );
  NAND2_X1 U5977 ( .A1(n8848), .A2(n7453), .ZN(n8246) );
  AND2_X2 U5978 ( .A1(n4398), .A2(n4397), .ZN(n8654) );
  AOI21_X2 U5979 ( .B1(n4802), .B2(n4801), .A(n4800), .ZN(n8669) );
  OR2_X2 U5980 ( .A1(n8816), .A2(n4803), .ZN(n4802) );
  MUX2_X1 U5981 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(P2_DATAO_REG_2__SCAN_IN), 
        .S(n4968), .Z(n4875) );
  NAND2_X1 U5982 ( .A1(n4400), .A2(n4656), .ZN(n4399) );
  NAND2_X1 U5983 ( .A1(n5625), .A2(n4306), .ZN(n4400) );
  NAND2_X1 U5984 ( .A1(n4910), .A2(n4909), .ZN(n5157) );
  INV_X1 U5985 ( .A(n4410), .ZN(n6694) );
  NAND2_X1 U5986 ( .A1(n5288), .A2(n4945), .ZN(n4415) );
  INV_X1 U5987 ( .A(n4420), .ZN(n9486) );
  INV_X1 U5988 ( .A(n4418), .ZN(n9501) );
  NAND2_X1 U5989 ( .A1(n6270), .A2(n6269), .ZN(n4419) );
  NAND3_X1 U5990 ( .A1(n4686), .A2(n4687), .A3(P2_DATAO_REG_3__SCAN_IN), .ZN(
        n4433) );
  INV_X1 U5991 ( .A(n4687), .ZN(n4435) );
  OR2_X1 U5992 ( .A1(n9693), .A2(n6542), .ZN(n4445) );
  AOI21_X1 U5993 ( .B1(n6542), .B2(n6501), .A(n4447), .ZN(n4446) );
  NAND4_X1 U5994 ( .A1(n4767), .A2(n4465), .A3(n4464), .A4(n7590), .ZN(n7802)
         );
  OAI21_X1 U5995 ( .B1(n4468), .B2(n9666), .A(n4467), .ZN(P1_U3522) );
  INV_X1 U5996 ( .A(n4470), .ZN(n9108) );
  NAND3_X1 U5997 ( .A1(n4474), .A2(n4288), .A3(n8129), .ZN(n9206) );
  MUX2_X1 U5998 ( .A(n9474), .B(n4477), .S(n6283), .Z(n6794) );
  NAND2_X1 U6000 ( .A1(n4324), .A2(n8725), .ZN(n4818) );
  INV_X1 U6001 ( .A(n4485), .ZN(n8702) );
  NAND2_X1 U6002 ( .A1(n9382), .A2(n4491), .ZN(n4487) );
  NAND2_X1 U6003 ( .A1(n4489), .A2(n4486), .ZN(n7673) );
  OAI21_X1 U6004 ( .B1(n4809), .B2(n6097), .A(n5769), .ZN(n4492) );
  OR2_X2 U6005 ( .A1(n4322), .A2(n4492), .ZN(n7215) );
  INV_X2 U6006 ( .A(n7215), .ZN(n9792) );
  NAND3_X1 U6007 ( .A1(n4865), .A2(P1_ADDR_REG_19__SCAN_IN), .A3(
        P1_DATAO_REG_1__SCAN_IN), .ZN(n4493) );
  NAND3_X1 U6008 ( .A1(n4687), .A2(P2_DATAO_REG_1__SCAN_IN), .A3(n4686), .ZN(
        n4494) );
  NOR2_X4 U6009 ( .A1(n4293), .A2(n4497), .ZN(n6795) );
  OAI21_X1 U6010 ( .B1(n9398), .B2(n4503), .A(n4501), .ZN(n4500) );
  OAI21_X2 U6011 ( .B1(n4513), .B2(n4512), .A(n4510), .ZN(n5152) );
  INV_X1 U6012 ( .A(n9169), .ZN(n4521) );
  NAND3_X2 U6013 ( .A1(n4831), .A2(n4808), .A3(n4287), .ZN(n5667) );
  OAI21_X2 U6014 ( .B1(n6929), .B2(n5034), .A(n5634), .ZN(n6904) );
  NAND2_X1 U6015 ( .A1(n7391), .A2(n7390), .ZN(n7392) );
  NAND2_X1 U6016 ( .A1(n8972), .A2(n4559), .ZN(n4558) );
  OAI211_X1 U6017 ( .C1(n8972), .C2(n4560), .A(n4558), .B(n7950), .ZN(P1_U3218) );
  NAND2_X1 U6018 ( .A1(n8972), .A2(n7932), .ZN(n8885) );
  NAND2_X1 U6019 ( .A1(n4302), .A2(n4573), .ZN(n4570) );
  NAND2_X1 U6020 ( .A1(n8950), .A2(n4337), .ZN(n4569) );
  NAND2_X1 U6021 ( .A1(n4570), .A2(n4569), .ZN(n8891) );
  INV_X1 U6022 ( .A(n4302), .ZN(n4571) );
  INV_X1 U6023 ( .A(n7913), .ZN(n4573) );
  NAND2_X1 U6024 ( .A1(n7886), .A2(n7885), .ZN(n8944) );
  INV_X1 U6025 ( .A(n7825), .ZN(n7822) );
  OAI21_X2 U6026 ( .B1(n5667), .B2(n4776), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n5677) );
  XNOR2_X1 U6027 ( .A(n5675), .B(n5674), .ZN(n6235) );
  INV_X1 U6028 ( .A(n6235), .ZN(n6239) );
  NAND4_X1 U6029 ( .A1(n5724), .A2(n6137), .A3(n5723), .A4(n6159), .ZN(n5697)
         );
  AND2_X2 U6030 ( .A1(n4588), .A2(n4587), .ZN(n5724) );
  INV_X2 U6031 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n4587) );
  NAND2_X1 U6032 ( .A1(n4589), .A2(n4291), .ZN(n7044) );
  NAND3_X1 U6033 ( .A1(n4313), .A2(n7216), .A3(n4593), .ZN(n4589) );
  INV_X1 U6034 ( .A(n8343), .ZN(n4593) );
  NAND2_X1 U6035 ( .A1(n4590), .A2(n8209), .ZN(n7226) );
  NAND3_X1 U6036 ( .A1(n7216), .A2(n4593), .A3(n8189), .ZN(n4590) );
  INV_X1 U6037 ( .A(n8209), .ZN(n4592) );
  NAND2_X1 U6038 ( .A1(n4595), .A2(n4594), .ZN(n7445) );
  NAND3_X1 U6039 ( .A1(n5808), .A2(n5694), .A3(n4799), .ZN(n4605) );
  NAND4_X1 U6040 ( .A1(n5698), .A2(n5808), .A3(n5694), .A4(n4600), .ZN(n5715)
         );
  NAND2_X1 U6041 ( .A1(n4603), .A2(n4601), .ZN(n5718) );
  AND2_X1 U6042 ( .A1(n5698), .A2(n5699), .ZN(n4601) );
  INV_X1 U6043 ( .A(n5698), .ZN(n4604) );
  NAND2_X1 U6044 ( .A1(n4612), .A2(n4613), .ZN(n7754) );
  NAND2_X1 U6045 ( .A1(n7677), .A2(n4615), .ZN(n4612) );
  INV_X1 U6046 ( .A(n8716), .ZN(n4619) );
  NAND2_X1 U6047 ( .A1(n8642), .A2(n4653), .ZN(n4644) );
  AOI21_X1 U6048 ( .B1(n8642), .B2(n4634), .A(n4632), .ZN(n4648) );
  OAI21_X2 U6049 ( .B1(n5005), .B2(n4655), .A(n4873), .ZN(n5025) );
  NAND2_X1 U6050 ( .A1(n5088), .A2(n4662), .ZN(n4659) );
  NAND2_X1 U6051 ( .A1(n4659), .A2(n4660), .ZN(n5109) );
  NAND2_X1 U6052 ( .A1(n4975), .A2(n4668), .ZN(n4667) );
  NAND2_X1 U6053 ( .A1(n4975), .A2(n4672), .ZN(n4671) );
  NAND2_X1 U6054 ( .A1(n4975), .A2(n4974), .ZN(n5385) );
  NAND2_X1 U6055 ( .A1(n5460), .A2(n4682), .ZN(n4680) );
  OAI21_X1 U6056 ( .B1(n5460), .B2(n4684), .A(n4682), .ZN(n5496) );
  NAND2_X1 U6057 ( .A1(n4680), .A2(n4681), .ZN(n5494) );
  NAND2_X1 U6058 ( .A1(n5460), .A2(n5459), .ZN(n5476) );
  NAND3_X1 U6059 ( .A1(n4686), .A2(n4687), .A3(n4870), .ZN(n5015) );
  NAND2_X1 U6060 ( .A1(n5932), .A2(n4689), .ZN(n4688) );
  OAI211_X1 U6061 ( .C1(n8501), .C2(n4698), .A(n8042), .B(n4696), .ZN(P2_U3222) );
  NAND2_X1 U6062 ( .A1(n8501), .A2(n4697), .ZN(n4696) );
  AND2_X1 U6063 ( .A1(n4701), .A2(n4326), .ZN(n4699) );
  OAI21_X1 U6064 ( .B1(n4706), .B2(n8038), .A(n4702), .ZN(n4701) );
  INV_X1 U6065 ( .A(n8038), .ZN(n4704) );
  OAI21_X1 U6066 ( .B1(n8501), .B2(n8500), .A(n8009), .ZN(n8412) );
  NAND2_X1 U6068 ( .A1(n7955), .A2(n4713), .ZN(n5858) );
  NAND2_X1 U6069 ( .A1(n8426), .A2(n4714), .ZN(n8437) );
  NAND2_X1 U6070 ( .A1(n7980), .A2(n4715), .ZN(n6205) );
  OAI21_X1 U6071 ( .B1(n6009), .B2(n4718), .A(n4716), .ZN(n6047) );
  NAND2_X1 U6072 ( .A1(n5722), .A2(n4722), .ZN(n5725) );
  XNOR2_X2 U6073 ( .A(n4988), .B(P1_IR_REG_27__SCAN_IN), .ZN(n5683) );
  NAND2_X1 U6074 ( .A1(n6914), .A2(n4726), .ZN(n4728) );
  NAND3_X1 U6075 ( .A1(n9579), .A2(n6946), .A3(n5600), .ZN(n4727) );
  NAND2_X1 U6076 ( .A1(n9579), .A2(n5600), .ZN(n6943) );
  NAND2_X1 U6077 ( .A1(n7411), .A2(n7412), .ZN(n4730) );
  NAND2_X1 U6078 ( .A1(n8086), .A2(n4734), .ZN(n4733) );
  NAND2_X1 U6079 ( .A1(n4733), .A2(n4738), .ZN(n8091) );
  NAND2_X1 U6080 ( .A1(n9133), .A2(n4298), .ZN(n4749) );
  AOI21_X1 U6081 ( .B1(n9133), .B2(n8093), .A(n8092), .ZN(n9119) );
  AOI21_X1 U6082 ( .B1(n7418), .B2(n4773), .A(n4769), .ZN(n7576) );
  NOR3_X1 U6083 ( .A1(n5667), .A2(n4776), .A3(n4835), .ZN(n4984) );
  NAND2_X1 U6084 ( .A1(n4778), .A2(n8350), .ZN(n7041) );
  NAND2_X1 U6085 ( .A1(n7283), .A2(n4778), .ZN(n7285) );
  NAND2_X1 U6086 ( .A1(n7038), .A2(n7039), .ZN(n4778) );
  OAI21_X1 U6087 ( .B1(n8654), .B2(n4782), .A(n4781), .ZN(n8625) );
  NAND2_X1 U6088 ( .A1(n4780), .A2(n4779), .ZN(n8624) );
  NOR2_X1 U6089 ( .A1(n8659), .A2(n8674), .ZN(n4785) );
  NAND2_X1 U6090 ( .A1(n7748), .A2(n7747), .ZN(n4789) );
  NAND2_X1 U6091 ( .A1(n4787), .A2(n7756), .ZN(n4786) );
  INV_X1 U6092 ( .A(n7751), .ZN(n4787) );
  NAND2_X1 U6093 ( .A1(n7752), .A2(n7756), .ZN(n8387) );
  NAND3_X1 U6094 ( .A1(n5754), .A2(n4790), .A3(n5687), .ZN(n5781) );
  NAND2_X1 U6095 ( .A1(n4793), .A2(n4791), .ZN(n7650) );
  NAND2_X1 U6096 ( .A1(n4796), .A2(n4792), .ZN(n4791) );
  INV_X1 U6097 ( .A(n7431), .ZN(n4792) );
  NOR2_X1 U6098 ( .A1(n4794), .A2(n8253), .ZN(n4793) );
  NAND2_X1 U6099 ( .A1(n7429), .A2(n4796), .ZN(n4797) );
  NAND3_X1 U6100 ( .A1(n7356), .A2(n7070), .A3(n8352), .ZN(n7324) );
  AND2_X1 U6101 ( .A1(n5808), .A2(n5694), .ZN(n5722) );
  NAND3_X1 U6102 ( .A1(n5808), .A2(n5698), .A3(n5694), .ZN(n6140) );
  OAI21_X1 U6103 ( .B1(n8585), .B2(n8403), .A(n8402), .ZN(n8405) );
  NAND2_X1 U6104 ( .A1(n6580), .A2(n6581), .ZN(n6579) );
  NAND2_X1 U6105 ( .A1(n6644), .A2(n9761), .ZN(n9764) );
  OAI21_X1 U6106 ( .B1(n8163), .B2(n8168), .A(n8169), .ZN(n8164) );
  INV_X1 U6107 ( .A(n6015), .ZN(n6016) );
  NAND2_X1 U6108 ( .A1(n8165), .A2(n6630), .ZN(n5749) );
  XNOR2_X1 U6109 ( .A(n5088), .B(n5087), .ZN(n6227) );
  NAND2_X1 U6110 ( .A1(n5725), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5726) );
  INV_X1 U6111 ( .A(n5992), .ZN(n5995) );
  NAND2_X1 U6112 ( .A1(n5992), .A2(n5993), .ZN(n7770) );
  AND2_X1 U6113 ( .A1(n6128), .A2(n6127), .ZN(n7984) );
  OR2_X1 U6114 ( .A1(n5702), .A2(n8873), .ZN(n5703) );
  OAI21_X2 U6115 ( .B1(n8454), .B2(n8450), .A(n8453), .ZN(n8501) );
  INV_X1 U6116 ( .A(n4842), .ZN(n7855) );
  NAND2_X1 U6117 ( .A1(n7208), .A2(n7209), .ZN(n7207) );
  OAI222_X1 U6118 ( .A1(n9581), .A2(n8127), .B1(n5532), .B2(n8126), .C1(n8999), 
        .C2(n9423), .ZN(n8128) );
  AND2_X1 U6119 ( .A1(n7983), .A2(n7981), .ZN(n8424) );
  NAND2_X1 U6120 ( .A1(n8010), .A2(n6129), .ZN(n8012) );
  AND2_X1 U6121 ( .A1(n9085), .A2(n5472), .ZN(n4805) );
  OR2_X1 U6122 ( .A1(n5876), .A2(n8167), .ZN(n4806) );
  AND4_X1 U6123 ( .A1(n4862), .A2(n4859), .A3(n5524), .A4(n4860), .ZN(n4808)
         );
  XOR2_X1 U6124 ( .A(n5042), .B(n5041), .Z(n4809) );
  OR2_X1 U6125 ( .A1(n7988), .A2(n7987), .ZN(n4810) );
  OR2_X1 U6126 ( .A1(n9081), .A2(n8999), .ZN(n4812) );
  AND2_X1 U6127 ( .A1(n6787), .A2(n6786), .ZN(n9586) );
  AND2_X1 U6128 ( .A1(n7982), .A2(n7981), .ZN(n4813) );
  OR2_X1 U6129 ( .A1(n9151), .A2(n8090), .ZN(n4814) );
  AND4_X1 U6130 ( .A1(n5454), .A2(n5453), .A3(n5452), .A4(n5451), .ZN(n10020)
         );
  AND2_X1 U6131 ( .A1(n4903), .A2(n4902), .ZN(n4816) );
  AND2_X1 U6132 ( .A1(n4909), .A2(n4908), .ZN(n4817) );
  INV_X1 U6133 ( .A(n7486), .ZN(n5139) );
  NOR2_X1 U6134 ( .A1(n5316), .A2(n5314), .ZN(n4819) );
  INV_X1 U6135 ( .A(n8644), .ZN(n8614) );
  AND2_X1 U6136 ( .A1(n6192), .A2(n6191), .ZN(n8644) );
  AND2_X1 U6137 ( .A1(n8709), .A2(n8695), .ZN(n4820) );
  INV_X1 U6138 ( .A(n8790), .ZN(n8393) );
  AND2_X1 U6139 ( .A1(n5405), .A2(n9278), .ZN(n4821) );
  OR2_X1 U6140 ( .A1(n8376), .A2(n8339), .ZN(n4822) );
  INV_X1 U6141 ( .A(n9646), .ZN(n7091) );
  NAND2_X1 U6142 ( .A1(n5431), .A2(n9278), .ZN(n5432) );
  NAND2_X1 U6143 ( .A1(n5433), .A2(n5432), .ZN(n5434) );
  INV_X1 U6144 ( .A(n5473), .ZN(n5474) );
  OR2_X1 U6145 ( .A1(n7986), .A2(n8663), .ZN(n7982) );
  NOR3_X1 U6146 ( .A1(P1_IR_REG_4__SCAN_IN), .A2(P1_IR_REG_12__SCAN_IN), .A3(
        P1_IR_REG_5__SCAN_IN), .ZN(n4827) );
  INV_X1 U6147 ( .A(n8170), .ZN(n8155) );
  NAND2_X1 U6148 ( .A1(n9008), .A2(n7939), .ZN(n6651) );
  NAND2_X1 U6149 ( .A1(n4834), .A2(n4833), .ZN(n4835) );
  NOR2_X1 U6150 ( .A1(n6112), .A2(n6111), .ZN(n6113) );
  INV_X1 U6151 ( .A(n5921), .ZN(n5920) );
  INV_X1 U6152 ( .A(n6025), .ZN(n6023) );
  NAND2_X1 U6153 ( .A1(n7047), .A2(n7046), .ZN(n7294) );
  INV_X1 U6154 ( .A(n5354), .ZN(n4844) );
  INV_X1 U6155 ( .A(n5338), .ZN(n4845) );
  INV_X1 U6156 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n5095) );
  INV_X1 U6157 ( .A(n5369), .ZN(n4846) );
  OR2_X1 U6158 ( .A1(n7176), .A2(n9005), .ZN(n5563) );
  INV_X1 U6159 ( .A(n9401), .ZN(n7794) );
  OR2_X1 U6160 ( .A1(n5344), .A2(n5348), .ZN(n5328) );
  INV_X1 U6161 ( .A(n5104), .ZN(n4891) );
  INV_X1 U6162 ( .A(n5846), .ZN(n5844) );
  INV_X1 U6163 ( .A(n7785), .ZN(n6008) );
  NAND2_X1 U6164 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n5801) );
  INV_X1 U6165 ( .A(n4282), .ZN(n5730) );
  NAND2_X1 U6166 ( .A1(n6082), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n6101) );
  NAND2_X1 U6167 ( .A1(n6116), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n6186) );
  AND2_X1 U6168 ( .A1(n6594), .A2(n6593), .ZN(n6591) );
  NAND2_X1 U6169 ( .A1(n6023), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n6039) );
  NAND2_X1 U6170 ( .A1(n7217), .A2(n8341), .ZN(n7216) );
  INV_X1 U6171 ( .A(n8653), .ZN(n8662) );
  NAND2_X1 U6172 ( .A1(n7328), .A2(n8356), .ZN(n7677) );
  INV_X1 U6173 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n5700) );
  NAND2_X1 U6174 ( .A1(n4844), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n5338) );
  NAND2_X1 U6175 ( .A1(n5260), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n5279) );
  AND2_X1 U6176 ( .A1(n7846), .A2(n7847), .ZN(n7844) );
  NAND2_X1 U6177 ( .A1(n4845), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n5369) );
  OR2_X1 U6178 ( .A1(n5279), .A2(n5278), .ZN(n5293) );
  NAND2_X1 U6179 ( .A1(n4846), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n5391) );
  NAND2_X1 U6180 ( .A1(n9399), .A2(n9400), .ZN(n9398) );
  NOR2_X1 U6181 ( .A1(n5163), .A2(n5162), .ZN(n5185) );
  INV_X1 U6182 ( .A(n7419), .ZN(n7420) );
  INV_X1 U6183 ( .A(n6982), .ZN(n6981) );
  INV_X1 U6184 ( .A(n5193), .ZN(n4925) );
  NAND2_X1 U6185 ( .A1(n4894), .A2(n4893), .ZN(n4897) );
  NAND2_X1 U6186 ( .A1(n5844), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n5869) );
  OR2_X1 U6187 ( .A1(n5938), .A2(n5937), .ZN(n5952) );
  NAND2_X1 U6188 ( .A1(n5799), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n5826) );
  OR2_X1 U6189 ( .A1(n6101), .A2(n6100), .ZN(n6118) );
  NAND2_X1 U6190 ( .A1(n5824), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5846) );
  OR2_X1 U6191 ( .A1(n5986), .A2(n9998), .ZN(n6002) );
  NAND2_X1 U6192 ( .A1(n8376), .A2(n8375), .ZN(n8377) );
  OR2_X1 U6193 ( .A1(n8620), .A2(n8001), .ZN(n8006) );
  OR2_X1 U6194 ( .A1(n6039), .A2(n7626), .ZN(n6052) );
  NAND2_X1 U6195 ( .A1(n5828), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n5747) );
  OR2_X1 U6196 ( .A1(n6628), .A2(n6193), .ZN(n8721) );
  NAND2_X1 U6197 ( .A1(n7930), .A2(n7931), .ZN(n7932) );
  AND2_X1 U6198 ( .A1(n7900), .A2(n7901), .ZN(n8909) );
  AND2_X1 U6199 ( .A1(n9319), .A2(n9200), .ZN(n8088) );
  INV_X1 U6200 ( .A(n8123), .ZN(n8098) );
  INV_X1 U6201 ( .A(n9660), .ZN(n9572) );
  XNOR2_X1 U6202 ( .A(n4911), .B(SI_11_), .ZN(n5156) );
  AND2_X1 U6203 ( .A1(n8462), .A2(n8753), .ZN(n8504) );
  INV_X1 U6204 ( .A(n8013), .ZN(n8154) );
  AND4_X1 U6205 ( .A1(n5957), .A2(n5956), .A3(n5955), .A4(n5954), .ZN(n7679)
         );
  INV_X1 U6206 ( .A(n9692), .ZN(n9744) );
  INV_X1 U6207 ( .A(n9768), .ZN(n8736) );
  AND2_X1 U6208 ( .A1(n8729), .A2(n9381), .ZN(n9798) );
  NAND2_X1 U6209 ( .A1(n9778), .A2(n6144), .ZN(n9773) );
  INV_X1 U6210 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n6137) );
  AND2_X1 U6211 ( .A1(n5864), .A2(n5863), .ZN(n6563) );
  AND2_X1 U6212 ( .A1(n6380), .A2(n6760), .ZN(n9345) );
  AND4_X1 U6213 ( .A1(n5343), .A2(n5342), .A3(n5341), .A4(n5340), .ZN(n8087)
         );
  AND4_X1 U6214 ( .A1(n5299), .A2(n5298), .A3(n5297), .A4(n5296), .ZN(n8928)
         );
  AND4_X1 U6215 ( .A1(n5225), .A2(n5224), .A3(n5223), .A4(n5222), .ZN(n7697)
         );
  INV_X1 U6216 ( .A(n9100), .ZN(n9092) );
  NAND2_X1 U6217 ( .A1(n9168), .A2(n8111), .ZN(n9185) );
  AOI21_X1 U6218 ( .B1(n9250), .B2(n9249), .A(n8080), .ZN(n9233) );
  INV_X1 U6219 ( .A(n9345), .ZN(n9658) );
  AND2_X1 U6220 ( .A1(n9405), .A2(n9404), .ZN(n9450) );
  OR3_X1 U6221 ( .A1(n6235), .A2(n6238), .A3(n6237), .ZN(n9601) );
  AND2_X1 U6222 ( .A1(n5114), .A2(n5141), .ZN(n6301) );
  XNOR2_X1 U6223 ( .A(n4884), .B(SI_5_), .ZN(n5072) );
  OR3_X1 U6224 ( .A1(n7199), .A2(n7524), .A3(n7458), .ZN(n6473) );
  INV_X1 U6225 ( .A(n6197), .ZN(n6198) );
  INV_X1 U6226 ( .A(n8503), .ZN(n8615) );
  INV_X1 U6227 ( .A(n8700), .ZN(n8515) );
  AND4_X1 U6228 ( .A1(n5991), .A2(n5990), .A3(n5989), .A4(n5988), .ZN(n8050)
         );
  INV_X1 U6229 ( .A(n9840), .ZN(n9837) );
  OR3_X1 U6230 ( .A1(n8821), .A2(n8820), .A3(n8819), .ZN(n8865) );
  OR2_X1 U6231 ( .A1(n6814), .A2(n6625), .ZN(n9827) );
  AND2_X1 U6232 ( .A1(n6252), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9783) );
  INV_X1 U6233 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n9941) );
  INV_X1 U6234 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n9914) );
  INV_X1 U6235 ( .A(n8094), .ZN(n9128) );
  AND4_X1 U6236 ( .A1(n5207), .A2(n5206), .A3(n5205), .A4(n5204), .ZN(n9401)
         );
  OR2_X1 U6237 ( .A1(n9272), .A2(n9271), .ZN(n9676) );
  AND2_X1 U6238 ( .A1(n9450), .A2(n9449), .ZN(n9468) );
  AND2_X1 U6239 ( .A1(n9462), .A2(n9461), .ZN(n9471) );
  OR2_X1 U6240 ( .A1(n9272), .A2(n6379), .ZN(n9666) );
  INV_X1 U6241 ( .A(n9604), .ZN(n9603) );
  INV_X1 U6242 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n9989) );
  INV_X1 U6243 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n4859) );
  INV_X1 U6244 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n5678) );
  NAND2_X1 U6245 ( .A1(n5676), .A2(n5674), .ZN(n4986) );
  INV_X1 U6246 ( .A(n4986), .ZN(n4834) );
  INV_X1 U6247 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n4833) );
  INV_X1 U6248 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n4836) );
  INV_X1 U6249 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n4840) );
  NAND2_X1 U6250 ( .A1(n4839), .A2(n4840), .ZN(n9367) );
  NAND2_X2 U6251 ( .A1(n7855), .A2(n8071), .ZN(n5019) );
  NAND2_X1 U6252 ( .A1(n5484), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n4857) );
  INV_X1 U6253 ( .A(P1_REG2_REG_29__SCAN_IN), .ZN(n8134) );
  OR2_X1 U6254 ( .A1(n5419), .A2(n8134), .ZN(n4856) );
  INV_X1 U6255 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n10003) );
  NAND2_X1 U6256 ( .A1(n5117), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n5130) );
  INV_X1 U6257 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n5129) );
  INV_X1 U6258 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n7394) );
  INV_X1 U6259 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n5162) );
  NAND2_X1 U6260 ( .A1(n5185), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n5218) );
  INV_X1 U6261 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n5217) );
  INV_X1 U6262 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n5202) );
  INV_X1 U6263 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n5278) );
  NAND2_X1 U6264 ( .A1(P1_REG3_REG_19__SCAN_IN), .A2(n5307), .ZN(n5306) );
  INV_X1 U6265 ( .A(n5393), .ZN(n4848) );
  NAND2_X1 U6266 ( .A1(n4848), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n5421) );
  INV_X1 U6267 ( .A(n5421), .ZN(n4849) );
  NAND2_X1 U6268 ( .A1(n4849), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n5448) );
  INV_X1 U6269 ( .A(n5448), .ZN(n4850) );
  NAND2_X1 U6270 ( .A1(n4850), .A2(P1_REG3_REG_27__SCAN_IN), .ZN(n5464) );
  INV_X1 U6271 ( .A(n5464), .ZN(n4851) );
  NAND2_X1 U6272 ( .A1(n4851), .A2(P1_REG3_REG_28__SCAN_IN), .ZN(n8133) );
  OR2_X1 U6273 ( .A1(n5466), .A2(n8133), .ZN(n4855) );
  INV_X1 U6274 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n4853) );
  OR2_X1 U6275 ( .A1(n5492), .A2(n4853), .ZN(n4854) );
  INV_X1 U6276 ( .A(n7947), .ZN(n9087) );
  NAND2_X1 U6277 ( .A1(n4863), .A2(n4862), .ZN(n4858) );
  NAND2_X1 U6278 ( .A1(n5527), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4861) );
  XNOR2_X1 U6279 ( .A(n4863), .B(n4862), .ZN(n9141) );
  INV_X1 U6280 ( .A(n9141), .ZN(n9592) );
  NAND2_X1 U6281 ( .A1(n7004), .A2(n9592), .ZN(n9278) );
  AND2_X1 U6282 ( .A1(SI_0_), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n4870) );
  AND2_X1 U6283 ( .A1(SI_0_), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n4871) );
  NAND2_X1 U6284 ( .A1(n6213), .A2(n4871), .ZN(n5713) );
  NAND2_X1 U6285 ( .A1(n5015), .A2(n5713), .ZN(n4872) );
  NAND2_X1 U6286 ( .A1(n4872), .A2(SI_1_), .ZN(n4873) );
  XNOR2_X1 U6287 ( .A(n4875), .B(SI_2_), .ZN(n5026) );
  INV_X1 U6288 ( .A(n5026), .ZN(n4874) );
  NAND2_X1 U6289 ( .A1(n4875), .A2(SI_2_), .ZN(n4876) );
  NAND2_X1 U6290 ( .A1(n4878), .A2(SI_3_), .ZN(n4879) );
  MUX2_X1 U6291 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(P2_DATAO_REG_4__SCAN_IN), 
        .S(n4279), .Z(n4881) );
  NAND2_X1 U6292 ( .A1(n5056), .A2(n4880), .ZN(n4883) );
  NAND2_X1 U6293 ( .A1(n4881), .A2(SI_4_), .ZN(n4882) );
  MUX2_X1 U6294 ( .A(n6217), .B(n9901), .S(n4279), .Z(n4884) );
  NAND2_X1 U6295 ( .A1(n5073), .A2(n5072), .ZN(n4887) );
  INV_X1 U6296 ( .A(n4884), .ZN(n4885) );
  NAND2_X1 U6297 ( .A1(n4885), .A2(SI_5_), .ZN(n4886) );
  MUX2_X1 U6298 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .S(n4280), .Z(n4889) );
  NAND2_X1 U6299 ( .A1(n4889), .A2(SI_6_), .ZN(n4890) );
  MUX2_X1 U6300 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .S(n4279), .Z(n4892) );
  MUX2_X1 U6301 ( .A(n9914), .B(n9989), .S(n4279), .Z(n4894) );
  INV_X1 U6302 ( .A(SI_8_), .ZN(n4893) );
  INV_X1 U6303 ( .A(n4894), .ZN(n4895) );
  NAND2_X1 U6304 ( .A1(n4895), .A2(SI_8_), .ZN(n4896) );
  INV_X1 U6305 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n4898) );
  MUX2_X1 U6306 ( .A(n9941), .B(n4898), .S(n4280), .Z(n4900) );
  INV_X1 U6307 ( .A(SI_9_), .ZN(n4899) );
  INV_X1 U6308 ( .A(n4900), .ZN(n4901) );
  NAND2_X1 U6309 ( .A1(n4901), .A2(SI_9_), .ZN(n4902) );
  INV_X1 U6310 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n6251) );
  INV_X1 U6311 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n4904) );
  MUX2_X1 U6312 ( .A(n6251), .B(n4904), .S(n4279), .Z(n4906) );
  INV_X1 U6313 ( .A(SI_10_), .ZN(n4905) );
  NAND2_X1 U6314 ( .A1(n4906), .A2(n4905), .ZN(n4909) );
  INV_X1 U6315 ( .A(n4906), .ZN(n4907) );
  NAND2_X1 U6316 ( .A1(n4907), .A2(SI_10_), .ZN(n4908) );
  INV_X1 U6317 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n6312) );
  INV_X1 U6318 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n6263) );
  MUX2_X1 U6319 ( .A(n6312), .B(n6263), .S(n4280), .Z(n4911) );
  INV_X1 U6320 ( .A(n4911), .ZN(n4912) );
  NAND2_X1 U6321 ( .A1(n4912), .A2(SI_11_), .ZN(n4913) );
  INV_X1 U6322 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n6330) );
  INV_X1 U6323 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n6328) );
  MUX2_X1 U6324 ( .A(n6330), .B(n6328), .S(n4280), .Z(n4915) );
  INV_X1 U6325 ( .A(SI_12_), .ZN(n4914) );
  NAND2_X1 U6326 ( .A1(n4915), .A2(n4914), .ZN(n5208) );
  INV_X1 U6327 ( .A(n4915), .ZN(n4916) );
  NAND2_X1 U6328 ( .A1(n4916), .A2(SI_12_), .ZN(n4917) );
  NAND2_X1 U6329 ( .A1(n5208), .A2(n4917), .ZN(n5177) );
  INV_X1 U6330 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n6336) );
  INV_X1 U6331 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n6334) );
  MUX2_X1 U6332 ( .A(n6336), .B(n6334), .S(n4280), .Z(n4919) );
  INV_X1 U6333 ( .A(SI_13_), .ZN(n4918) );
  NAND2_X1 U6334 ( .A1(n4919), .A2(n4918), .ZN(n5211) );
  INV_X1 U6335 ( .A(n4919), .ZN(n4920) );
  NAND2_X1 U6336 ( .A1(n4920), .A2(SI_13_), .ZN(n5210) );
  INV_X1 U6337 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n6375) );
  INV_X1 U6338 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n6338) );
  MUX2_X1 U6339 ( .A(n6375), .B(n6338), .S(n4279), .Z(n4922) );
  XNOR2_X1 U6340 ( .A(n4922), .B(SI_14_), .ZN(n5193) );
  INV_X1 U6341 ( .A(n4922), .ZN(n4923) );
  NAND2_X1 U6342 ( .A1(n4923), .A2(SI_14_), .ZN(n4924) );
  INV_X1 U6343 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n4927) );
  INV_X1 U6344 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n4926) );
  MUX2_X1 U6345 ( .A(n4927), .B(n4926), .S(n4280), .Z(n4929) );
  INV_X1 U6346 ( .A(SI_15_), .ZN(n4928) );
  NAND2_X1 U6347 ( .A1(n4929), .A2(n4928), .ZN(n4932) );
  INV_X1 U6348 ( .A(n4929), .ZN(n4930) );
  NAND2_X1 U6349 ( .A1(n4930), .A2(SI_15_), .ZN(n4931) );
  NAND2_X1 U6350 ( .A1(n4932), .A2(n4931), .ZN(n5236) );
  INV_X1 U6351 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n6549) );
  INV_X1 U6352 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n4933) );
  MUX2_X1 U6353 ( .A(n6549), .B(n4933), .S(n4280), .Z(n4935) );
  INV_X1 U6354 ( .A(SI_16_), .ZN(n4934) );
  NAND2_X1 U6355 ( .A1(n4935), .A2(n4934), .ZN(n4938) );
  INV_X1 U6356 ( .A(n4935), .ZN(n4936) );
  NAND2_X1 U6357 ( .A1(n4936), .A2(SI_16_), .ZN(n4937) );
  NAND2_X1 U6358 ( .A1(n5254), .A2(n5253), .ZN(n4939) );
  INV_X1 U6359 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n6649) );
  INV_X1 U6360 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n4940) );
  MUX2_X1 U6361 ( .A(n6649), .B(n4940), .S(n4280), .Z(n4941) );
  XNOR2_X1 U6362 ( .A(n4941), .B(SI_17_), .ZN(n5271) );
  INV_X1 U6363 ( .A(n5271), .ZN(n4944) );
  INV_X1 U6364 ( .A(n4941), .ZN(n4942) );
  NAND2_X1 U6365 ( .A1(n4942), .A2(SI_17_), .ZN(n4943) );
  MUX2_X1 U6366 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .S(n4279), .Z(n4946) );
  XNOR2_X1 U6367 ( .A(n4946), .B(SI_18_), .ZN(n5287) );
  NAND2_X1 U6368 ( .A1(n4946), .A2(SI_18_), .ZN(n4947) );
  INV_X1 U6369 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n6891) );
  INV_X1 U6370 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n6893) );
  MUX2_X1 U6371 ( .A(n6891), .B(n6893), .S(n4280), .Z(n4948) );
  INV_X1 U6372 ( .A(SI_19_), .ZN(n9988) );
  NAND2_X1 U6373 ( .A1(n4948), .A2(n9988), .ZN(n5346) );
  INV_X1 U6374 ( .A(n4948), .ZN(n4949) );
  NAND2_X1 U6375 ( .A1(n4949), .A2(SI_19_), .ZN(n4950) );
  NAND2_X1 U6376 ( .A1(n5346), .A2(n4950), .ZN(n5344) );
  INV_X1 U6377 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n9997) );
  INV_X1 U6378 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n6973) );
  MUX2_X1 U6379 ( .A(n9997), .B(n6973), .S(n4280), .Z(n4952) );
  INV_X1 U6380 ( .A(SI_20_), .ZN(n4951) );
  NAND2_X1 U6381 ( .A1(n4952), .A2(n4951), .ZN(n4961) );
  INV_X1 U6382 ( .A(n4952), .ZN(n4953) );
  NAND2_X1 U6383 ( .A1(n4953), .A2(SI_20_), .ZN(n4954) );
  NAND2_X1 U6384 ( .A1(n4961), .A2(n4954), .ZN(n5348) );
  INV_X1 U6385 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n6992) );
  INV_X1 U6386 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n6975) );
  MUX2_X1 U6387 ( .A(n6992), .B(n6975), .S(n4279), .Z(n4963) );
  INV_X1 U6388 ( .A(n4963), .ZN(n4955) );
  AND2_X1 U6389 ( .A1(n4955), .A2(SI_21_), .ZN(n4965) );
  INV_X1 U6390 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n7954) );
  INV_X1 U6391 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n7005) );
  MUX2_X1 U6392 ( .A(n7954), .B(n7005), .S(n4280), .Z(n4957) );
  INV_X1 U6393 ( .A(SI_22_), .ZN(n4956) );
  NAND2_X1 U6394 ( .A1(n4957), .A2(n4956), .ZN(n4966) );
  INV_X1 U6395 ( .A(n4957), .ZN(n4958) );
  NAND2_X1 U6396 ( .A1(n4958), .A2(SI_22_), .ZN(n4959) );
  NAND2_X1 U6397 ( .A1(n4966), .A2(n4959), .ZN(n5316) );
  OR2_X1 U6398 ( .A1(n5348), .A2(n5346), .ZN(n4962) );
  XNOR2_X1 U6399 ( .A(n4963), .B(SI_21_), .ZN(n5331) );
  INV_X1 U6400 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n9961) );
  INV_X1 U6401 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n4969) );
  MUX2_X1 U6402 ( .A(n9961), .B(n4969), .S(n4279), .Z(n4971) );
  INV_X1 U6403 ( .A(SI_23_), .ZN(n4970) );
  NAND2_X1 U6404 ( .A1(n4971), .A2(n4970), .ZN(n4974) );
  INV_X1 U6405 ( .A(n4971), .ZN(n4972) );
  NAND2_X1 U6406 ( .A1(n4972), .A2(SI_23_), .ZN(n4973) );
  AND2_X1 U6407 ( .A1(n4974), .A2(n4973), .ZN(n5364) );
  INV_X1 U6408 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n7197) );
  INV_X1 U6409 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n7164) );
  MUX2_X1 U6410 ( .A(n7197), .B(n7164), .S(n4279), .Z(n4976) );
  XNOR2_X1 U6411 ( .A(n4976), .B(SI_24_), .ZN(n5386) );
  INV_X1 U6412 ( .A(n5386), .ZN(n4979) );
  INV_X1 U6413 ( .A(n4976), .ZN(n4977) );
  NAND2_X1 U6414 ( .A1(n4977), .A2(SI_24_), .ZN(n4978) );
  INV_X1 U6415 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n10000) );
  INV_X1 U6416 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n7461) );
  MUX2_X1 U6417 ( .A(n10000), .B(n7461), .S(n4280), .Z(n4981) );
  INV_X1 U6418 ( .A(SI_25_), .ZN(n4980) );
  NAND2_X1 U6419 ( .A1(n4981), .A2(n4980), .ZN(n5409) );
  INV_X1 U6420 ( .A(n4981), .ZN(n4982) );
  NAND2_X1 U6421 ( .A1(n4982), .A2(SI_25_), .ZN(n4983) );
  NAND2_X1 U6422 ( .A1(n5409), .A2(n4983), .ZN(n5410) );
  NAND2_X1 U6423 ( .A1(n4986), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4987) );
  NAND2_X1 U6424 ( .A1(n5677), .A2(n4987), .ZN(n4988) );
  NAND2_X1 U6425 ( .A1(n7991), .A2(n5509), .ZN(n4990) );
  NAND2_X1 U6426 ( .A1(n5480), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n4989) );
  NAND2_X1 U6427 ( .A1(n4278), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n4998) );
  INV_X1 U6428 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n4991) );
  OR2_X1 U6429 ( .A1(n5492), .A2(n4991), .ZN(n4997) );
  INV_X1 U6430 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n4992) );
  NAND2_X1 U6431 ( .A1(n5393), .A2(n4992), .ZN(n4993) );
  NAND2_X1 U6432 ( .A1(n5421), .A2(n4993), .ZN(n9122) );
  OR2_X1 U6433 ( .A1(n5466), .A2(n9122), .ZN(n4996) );
  INV_X1 U6434 ( .A(P1_REG0_REG_25__SCAN_IN), .ZN(n4994) );
  OR2_X1 U6435 ( .A1(n5019), .A2(n4994), .ZN(n4995) );
  INV_X1 U6436 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n6796) );
  NAND2_X1 U6437 ( .A1(n4277), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n5002) );
  INV_X1 U6438 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n4999) );
  OR2_X1 U6439 ( .A1(n5019), .A2(n4999), .ZN(n5001) );
  INV_X1 U6440 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n6288) );
  XNOR2_X1 U6441 ( .A(n5005), .B(n5004), .ZN(n5735) );
  INV_X1 U6442 ( .A(n5735), .ZN(n6220) );
  INV_X1 U6443 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n6221) );
  INV_X1 U6444 ( .A(n6283), .ZN(n5029) );
  NAND2_X1 U6445 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5006) );
  INV_X1 U6446 ( .A(n5035), .ZN(n5007) );
  NAND2_X1 U6447 ( .A1(n5007), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n5012) );
  INV_X1 U6448 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n9473) );
  NAND2_X1 U6449 ( .A1(n4278), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n5010) );
  INV_X1 U6450 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n5008) );
  OR2_X1 U6451 ( .A1(n5019), .A2(n5008), .ZN(n5009) );
  INV_X1 U6452 ( .A(SI_0_), .ZN(n5014) );
  INV_X1 U6453 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n5013) );
  OAI21_X1 U6454 ( .B1(n4499), .B2(n5014), .A(n5013), .ZN(n5016) );
  AND2_X1 U6455 ( .A1(n5016), .A2(n5015), .ZN(n9373) );
  OR2_X1 U6456 ( .A1(n6897), .A2(n6795), .ZN(n5017) );
  INV_X1 U6457 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n6468) );
  INV_X1 U6458 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n6287) );
  INV_X1 U6459 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n5018) );
  OR2_X1 U6460 ( .A1(n5019), .A2(n5018), .ZN(n5022) );
  NAND2_X1 U6461 ( .A1(n4278), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n5021) );
  XNOR2_X1 U6462 ( .A(n5026), .B(n5025), .ZN(n5752) );
  INV_X1 U6463 ( .A(n5752), .ZN(n6218) );
  OR2_X1 U6464 ( .A1(n5027), .A2(n6218), .ZN(n5033) );
  OR2_X1 U6465 ( .A1(n5028), .A2(n4838), .ZN(n5044) );
  XNOR2_X1 U6466 ( .A(n5044), .B(P1_IR_REG_2__SCAN_IN), .ZN(n6291) );
  NAND2_X1 U6467 ( .A1(n5029), .A2(n6291), .ZN(n5032) );
  INV_X1 U6468 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n6219) );
  OR2_X1 U6469 ( .A1(n5030), .A2(n6219), .ZN(n5031) );
  INV_X1 U6470 ( .A(n5541), .ZN(n5034) );
  NAND2_X1 U6471 ( .A1(n6448), .A2(n9612), .ZN(n5634) );
  INV_X1 U6472 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n6268) );
  OR2_X1 U6473 ( .A1(n5035), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n5038) );
  INV_X1 U6474 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n6293) );
  OR2_X1 U6475 ( .A1(n5119), .A2(n6293), .ZN(n5037) );
  NAND2_X1 U6476 ( .A1(n5484), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n5036) );
  OR2_X1 U6477 ( .A1(n5027), .A2(n4809), .ZN(n5049) );
  INV_X1 U6478 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n6226) );
  OR2_X1 U6479 ( .A1(n5030), .A2(n6226), .ZN(n5048) );
  INV_X1 U6480 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n5043) );
  NAND2_X1 U6481 ( .A1(n5044), .A2(n5043), .ZN(n5045) );
  NAND2_X1 U6482 ( .A1(n5045), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5046) );
  XNOR2_X1 U6483 ( .A(n5046), .B(P1_IR_REG_3__SCAN_IN), .ZN(n6294) );
  NAND2_X1 U6484 ( .A1(n5303), .A2(n6294), .ZN(n5047) );
  NAND2_X1 U6485 ( .A1(n9008), .A2(n9618), .ZN(n5559) );
  OAI21_X1 U6486 ( .B1(n6904), .B2(n6911), .A(n5638), .ZN(n6916) );
  NAND2_X1 U6487 ( .A1(n5484), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n5054) );
  INV_X1 U6488 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n6269) );
  OR2_X1 U6489 ( .A1(n5419), .A2(n6269), .ZN(n5053) );
  INV_X1 U6490 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n5050) );
  OR2_X1 U6491 ( .A1(n5119), .A2(n5050), .ZN(n5052) );
  XNOR2_X1 U6492 ( .A(P1_REG3_REG_3__SCAN_IN), .B(P1_REG3_REG_4__SCAN_IN), 
        .ZN(n6920) );
  NAND4_X1 U6493 ( .A1(n5054), .A2(n5053), .A3(n5052), .A4(n5051), .ZN(n9585)
         );
  XNOR2_X1 U6494 ( .A(n5056), .B(n5055), .ZN(n5780) );
  INV_X1 U6495 ( .A(n5780), .ZN(n6222) );
  OR2_X1 U6496 ( .A1(n5027), .A2(n6222), .ZN(n5064) );
  INV_X1 U6497 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n6223) );
  OR2_X1 U6498 ( .A1(n5030), .A2(n6223), .ZN(n5063) );
  NOR2_X1 U6499 ( .A1(n5059), .A2(n4838), .ZN(n5057) );
  MUX2_X1 U6500 ( .A(n4838), .B(n5057), .S(P1_IR_REG_4__SCAN_IN), .Z(n5061) );
  INV_X1 U6501 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n5058) );
  NAND2_X1 U6502 ( .A1(n5059), .A2(n5058), .ZN(n5089) );
  INV_X1 U6503 ( .A(n5089), .ZN(n5060) );
  NAND2_X1 U6504 ( .A1(n5303), .A2(n9484), .ZN(n5062) );
  NAND2_X1 U6505 ( .A1(n9585), .A2(n9627), .ZN(n5600) );
  NAND2_X1 U6506 ( .A1(n6916), .A2(n5600), .ZN(n9580) );
  AOI21_X1 U6507 ( .B1(P1_REG3_REG_4__SCAN_IN), .B2(P1_REG3_REG_3__SCAN_IN), 
        .A(P1_REG3_REG_5__SCAN_IN), .ZN(n5065) );
  NOR2_X1 U6508 ( .A1(n5065), .A2(n5081), .ZN(n9587) );
  NAND2_X1 U6509 ( .A1(n5007), .A2(n9587), .ZN(n5071) );
  INV_X1 U6510 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n6271) );
  OR2_X1 U6511 ( .A1(n5419), .A2(n6271), .ZN(n5070) );
  INV_X1 U6512 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n5066) );
  OR2_X1 U6513 ( .A1(n5119), .A2(n5066), .ZN(n5069) );
  INV_X1 U6514 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n5067) );
  OR2_X1 U6515 ( .A1(n5019), .A2(n5067), .ZN(n5068) );
  NAND4_X1 U6516 ( .A1(n5071), .A2(n5070), .A3(n5069), .A4(n5068), .ZN(n9007)
         );
  XNOR2_X1 U6517 ( .A(n5073), .B(n5072), .ZN(n6225) );
  OR2_X1 U6518 ( .A1(n5030), .A2(n9901), .ZN(n5076) );
  NAND2_X1 U6519 ( .A1(n5089), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5074) );
  XNOR2_X1 U6520 ( .A(n5074), .B(P1_IR_REG_5__SCAN_IN), .ZN(n9500) );
  NAND2_X1 U6521 ( .A1(n5303), .A2(n9500), .ZN(n5075) );
  OR2_X1 U6522 ( .A1(n9007), .A2(n9633), .ZN(n5573) );
  OR2_X1 U6523 ( .A1(n9585), .A2(n9627), .ZN(n9579) );
  INV_X1 U6524 ( .A(n9579), .ZN(n5575) );
  NOR2_X1 U6525 ( .A1(n5078), .A2(n5575), .ZN(n5079) );
  NAND2_X1 U6526 ( .A1(n4278), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n5086) );
  INV_X1 U6527 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n5080) );
  OR2_X1 U6528 ( .A1(n5019), .A2(n5080), .ZN(n5085) );
  OAI21_X1 U6529 ( .B1(n5081), .B2(P1_REG3_REG_6__SCAN_IN), .A(n5096), .ZN(
        n7024) );
  OR2_X1 U6530 ( .A1(n5466), .A2(n7024), .ZN(n5084) );
  INV_X1 U6531 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n5082) );
  OR2_X1 U6532 ( .A1(n5119), .A2(n5082), .ZN(n5083) );
  NAND4_X1 U6533 ( .A1(n5086), .A2(n5085), .A3(n5084), .A4(n5083), .ZN(n9575)
         );
  NAND2_X1 U6534 ( .A1(n5509), .A2(n6227), .ZN(n5093) );
  INV_X1 U6535 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n6228) );
  OR2_X1 U6536 ( .A1(n5030), .A2(n6228), .ZN(n5092) );
  NAND2_X1 U6537 ( .A1(n5180), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5090) );
  XNOR2_X1 U6538 ( .A(n5090), .B(P1_IR_REG_6__SCAN_IN), .ZN(n9507) );
  NAND2_X1 U6539 ( .A1(n5303), .A2(n9507), .ZN(n5091) );
  NAND2_X1 U6540 ( .A1(n9575), .A2(n9639), .ZN(n6977) );
  NAND2_X1 U6541 ( .A1(n5484), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n5102) );
  INV_X1 U6542 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n5094) );
  OR2_X1 U6543 ( .A1(n5419), .A2(n5094), .ZN(n5101) );
  AND2_X1 U6544 ( .A1(n5096), .A2(n5095), .ZN(n5097) );
  OR2_X1 U6545 ( .A1(n5097), .A2(n5117), .ZN(n6985) );
  OR2_X1 U6546 ( .A1(n5466), .A2(n6985), .ZN(n5100) );
  INV_X1 U6547 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n5098) );
  OR2_X1 U6548 ( .A1(n5492), .A2(n5098), .ZN(n5099) );
  NAND4_X1 U6549 ( .A1(n5102), .A2(n5101), .A3(n5100), .A4(n5099), .ZN(n9006)
         );
  NOR2_X1 U6550 ( .A1(n5180), .A2(P1_IR_REG_6__SCAN_IN), .ZN(n5111) );
  OR2_X1 U6551 ( .A1(n5111), .A2(n4838), .ZN(n5103) );
  XNOR2_X1 U6552 ( .A(n5103), .B(P1_IR_REG_7__SCAN_IN), .ZN(n6300) );
  AOI22_X1 U6553 ( .A1(n5480), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n5303), .B2(
        n6300), .ZN(n5107) );
  XNOR2_X1 U6554 ( .A(n5105), .B(n5104), .ZN(n6231) );
  NAND2_X1 U6555 ( .A1(n6231), .A2(n5509), .ZN(n5106) );
  NAND2_X1 U6556 ( .A1(n9006), .A2(n9646), .ZN(n5543) );
  AND2_X1 U6557 ( .A1(n6977), .A2(n5543), .ZN(n5601) );
  OR2_X1 U6558 ( .A1(n9006), .A2(n9646), .ZN(n5562) );
  XNOR2_X1 U6559 ( .A(n5109), .B(n5108), .ZN(n6243) );
  NAND2_X1 U6560 ( .A1(n6243), .A2(n5509), .ZN(n5116) );
  INV_X1 U6561 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n5110) );
  NAND2_X1 U6562 ( .A1(n5111), .A2(n5110), .ZN(n5113) );
  NAND2_X1 U6563 ( .A1(n5113), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5112) );
  MUX2_X1 U6564 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5112), .S(
        P1_IR_REG_8__SCAN_IN), .Z(n5114) );
  AOI22_X1 U6565 ( .A1(n5480), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n5303), .B2(
        n6301), .ZN(n5115) );
  NAND2_X1 U6566 ( .A1(n5484), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n5123) );
  INV_X1 U6567 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n7101) );
  OR2_X1 U6568 ( .A1(n5419), .A2(n7101), .ZN(n5122) );
  OR2_X1 U6569 ( .A1(n5117), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n5118) );
  NAND2_X1 U6570 ( .A1(n5130), .A2(n5118), .ZN(n7351) );
  OR2_X1 U6571 ( .A1(n5466), .A2(n7351), .ZN(n5121) );
  INV_X1 U6572 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n6418) );
  OR2_X1 U6573 ( .A1(n5119), .A2(n6418), .ZN(n5120) );
  NAND4_X1 U6574 ( .A1(n5123), .A2(n5122), .A3(n5121), .A4(n5120), .ZN(n9005)
         );
  NAND2_X1 U6575 ( .A1(n7176), .A2(n9005), .ZN(n5581) );
  NAND2_X1 U6576 ( .A1(n5152), .A2(n5581), .ZN(n5124) );
  NAND2_X1 U6577 ( .A1(n6245), .A2(n5509), .ZN(n5128) );
  NAND2_X1 U6578 ( .A1(n5141), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5126) );
  XNOR2_X1 U6579 ( .A(n5126), .B(P1_IR_REG_9__SCAN_IN), .ZN(n9527) );
  AOI22_X1 U6580 ( .A1(n5480), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n5303), .B2(
        n9527), .ZN(n5127) );
  NAND2_X2 U6581 ( .A1(n5128), .A2(n5127), .ZN(n7484) );
  NAND2_X1 U6582 ( .A1(n5484), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n5137) );
  NAND2_X1 U6583 ( .A1(n5130), .A2(n5129), .ZN(n5131) );
  NAND2_X1 U6584 ( .A1(n5146), .A2(n5131), .ZN(n7482) );
  OR2_X1 U6585 ( .A1(n5466), .A2(n7482), .ZN(n5136) );
  INV_X1 U6586 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n5132) );
  OR2_X1 U6587 ( .A1(n5419), .A2(n5132), .ZN(n5135) );
  INV_X1 U6588 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n5133) );
  OR2_X1 U6589 ( .A1(n5492), .A2(n5133), .ZN(n5134) );
  NAND4_X1 U6590 ( .A1(n5137), .A2(n5136), .A3(n5135), .A4(n5134), .ZN(n9004)
         );
  INV_X1 U6591 ( .A(n9004), .ZN(n5138) );
  NAND2_X1 U6592 ( .A1(n7484), .A2(n5138), .ZN(n5565) );
  NAND2_X1 U6593 ( .A1(n5155), .A2(n5565), .ZN(n7486) );
  INV_X1 U6594 ( .A(n9278), .ZN(n5483) );
  XNOR2_X1 U6595 ( .A(n5140), .B(n4817), .ZN(n6248) );
  NAND2_X1 U6596 ( .A1(n6248), .A2(n5509), .ZN(n5144) );
  NAND2_X1 U6597 ( .A1(n5158), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5142) );
  XNOR2_X1 U6598 ( .A(n5142), .B(P1_IR_REG_10__SCAN_IN), .ZN(n9536) );
  AOI22_X1 U6599 ( .A1(n5480), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n5303), .B2(
        n9536), .ZN(n5143) );
  NAND2_X1 U6600 ( .A1(n4278), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n5151) );
  INV_X1 U6601 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n5145) );
  OR2_X1 U6602 ( .A1(n5019), .A2(n5145), .ZN(n5150) );
  NAND2_X1 U6603 ( .A1(n5146), .A2(n7394), .ZN(n5147) );
  NAND2_X1 U6604 ( .A1(n5163), .A2(n5147), .ZN(n7423) );
  OR2_X1 U6605 ( .A1(n5466), .A2(n7423), .ZN(n5149) );
  INV_X1 U6606 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n6421) );
  OR2_X1 U6607 ( .A1(n5492), .A2(n6421), .ZN(n5148) );
  NAND2_X1 U6608 ( .A1(n7571), .A2(n9424), .ZN(n7578) );
  NAND3_X1 U6609 ( .A1(n7579), .A2(n5483), .A3(n7578), .ZN(n5176) );
  INV_X1 U6610 ( .A(n5563), .ZN(n5153) );
  OAI21_X1 U6611 ( .B1(n7097), .B2(n5153), .A(n5581), .ZN(n5154) );
  NAND2_X1 U6612 ( .A1(n5154), .A2(n5565), .ZN(n5175) );
  NAND2_X1 U6613 ( .A1(n7580), .A2(n5155), .ZN(n5583) );
  NOR2_X1 U6614 ( .A1(n5583), .A2(n5483), .ZN(n5174) );
  XNOR2_X1 U6615 ( .A(n5157), .B(n5156), .ZN(n6262) );
  NAND2_X1 U6616 ( .A1(n6262), .A2(n5509), .ZN(n5161) );
  OAI21_X1 U6617 ( .B1(n5158), .B2(P1_IR_REG_10__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5159) );
  XNOR2_X1 U6618 ( .A(n5159), .B(P1_IR_REG_11__SCAN_IN), .ZN(n9552) );
  AOI22_X1 U6619 ( .A1(n5480), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n5303), .B2(
        n9552), .ZN(n5160) );
  NAND2_X1 U6620 ( .A1(n5484), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n5168) );
  INV_X1 U6621 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n9550) );
  OR2_X1 U6622 ( .A1(n5419), .A2(n9550), .ZN(n5167) );
  AND2_X1 U6623 ( .A1(n5163), .A2(n5162), .ZN(n5164) );
  OR2_X1 U6624 ( .A1(n5164), .A2(n5185), .ZN(n9419) );
  OR2_X1 U6625 ( .A1(n5466), .A2(n9419), .ZN(n5166) );
  INV_X1 U6626 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n6422) );
  OR2_X1 U6627 ( .A1(n5492), .A2(n6422), .ZN(n5165) );
  NAND4_X1 U6628 ( .A1(n5168), .A2(n5167), .A3(n5166), .A4(n5165), .ZN(n9002)
         );
  NOR2_X1 U6629 ( .A1(n9433), .A2(n9002), .ZN(n7574) );
  NAND2_X1 U6630 ( .A1(n9433), .A2(n9002), .ZN(n7575) );
  INV_X1 U6631 ( .A(n7575), .ZN(n5169) );
  OR2_X1 U6632 ( .A1(n7574), .A2(n5169), .ZN(n9411) );
  NOR2_X1 U6633 ( .A1(n9424), .A2(n9278), .ZN(n5171) );
  INV_X1 U6634 ( .A(n9424), .ZN(n9003) );
  OAI21_X1 U6635 ( .B1(n5483), .B2(n9003), .A(n7571), .ZN(n5170) );
  OAI21_X1 U6636 ( .B1(n5171), .B2(n7571), .A(n5170), .ZN(n5172) );
  NAND2_X1 U6637 ( .A1(n9411), .A2(n5172), .ZN(n5173) );
  NAND2_X1 U6638 ( .A1(n6327), .A2(n5509), .ZN(n5183) );
  INV_X1 U6639 ( .A(n5178), .ZN(n5179) );
  OAI21_X1 U6640 ( .B1(n5180), .B2(n5179), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n5181) );
  XNOR2_X1 U6641 ( .A(n5181), .B(P1_IR_REG_12__SCAN_IN), .ZN(n6695) );
  AOI22_X1 U6642 ( .A1(n5480), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n5303), .B2(
        n6695), .ZN(n5182) );
  NAND2_X1 U6643 ( .A1(n4278), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n5191) );
  INV_X1 U6644 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n5184) );
  OR2_X1 U6645 ( .A1(n5492), .A2(n5184), .ZN(n5190) );
  OR2_X1 U6646 ( .A1(n5185), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n5186) );
  NAND2_X1 U6647 ( .A1(n5218), .A2(n5186), .ZN(n7641) );
  OR2_X1 U6648 ( .A1(n5466), .A2(n7641), .ZN(n5189) );
  INV_X1 U6649 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n5187) );
  OR2_X1 U6650 ( .A1(n5019), .A2(n5187), .ZN(n5188) );
  OR2_X1 U6651 ( .A1(n7694), .A2(n9425), .ZN(n5546) );
  INV_X1 U6652 ( .A(n9002), .ZN(n7395) );
  OR2_X1 U6653 ( .A1(n9433), .A2(n7395), .ZN(n7583) );
  AND2_X1 U6654 ( .A1(n5546), .A2(n7583), .ZN(n7686) );
  NAND2_X1 U6655 ( .A1(n5230), .A2(n7686), .ZN(n5192) );
  NAND2_X1 U6656 ( .A1(n7694), .A2(n9425), .ZN(n7688) );
  NAND2_X1 U6657 ( .A1(n5192), .A2(n7688), .ZN(n5228) );
  XNOR2_X1 U6658 ( .A(n5194), .B(n5193), .ZN(n6337) );
  NAND2_X1 U6659 ( .A1(n6337), .A2(n5509), .ZN(n5201) );
  OR2_X1 U6660 ( .A1(n5195), .A2(P1_IR_REG_13__SCAN_IN), .ZN(n5197) );
  NAND2_X1 U6661 ( .A1(n5197), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5196) );
  MUX2_X1 U6662 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5196), .S(
        P1_IR_REG_14__SCAN_IN), .Z(n5199) );
  NOR2_X1 U6663 ( .A1(n5197), .A2(P1_IR_REG_14__SCAN_IN), .ZN(n5240) );
  INV_X1 U6664 ( .A(n5240), .ZN(n5198) );
  NAND2_X1 U6665 ( .A1(n5199), .A2(n5198), .ZN(n7258) );
  INV_X1 U6666 ( .A(n7258), .ZN(n6807) );
  AOI22_X1 U6667 ( .A1(n5480), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n5303), .B2(
        n6807), .ZN(n5200) );
  NAND2_X1 U6668 ( .A1(n5484), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n5207) );
  INV_X1 U6669 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n7698) );
  OR2_X1 U6670 ( .A1(n5419), .A2(n7698), .ZN(n5206) );
  AND2_X1 U6671 ( .A1(n5220), .A2(n5202), .ZN(n5203) );
  OR2_X1 U6672 ( .A1(n5203), .A2(n5245), .ZN(n7717) );
  OR2_X1 U6673 ( .A1(n5466), .A2(n7717), .ZN(n5205) );
  INV_X1 U6674 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n7257) );
  OR2_X1 U6675 ( .A1(n5492), .A2(n7257), .ZN(n5204) );
  NAND2_X1 U6676 ( .A1(n5209), .A2(n5208), .ZN(n5213) );
  AND2_X1 U6677 ( .A1(n5211), .A2(n5210), .ZN(n5212) );
  XNOR2_X1 U6678 ( .A(n5213), .B(n5212), .ZN(n6333) );
  NAND2_X1 U6679 ( .A1(n6333), .A2(n5509), .ZN(n5216) );
  NAND2_X1 U6680 ( .A1(n5195), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5214) );
  XNOR2_X1 U6681 ( .A(n5214), .B(P1_IR_REG_13__SCAN_IN), .ZN(n6806) );
  AOI22_X1 U6682 ( .A1(n5480), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n5303), .B2(
        n6806), .ZN(n5215) );
  NAND2_X1 U6683 ( .A1(n5484), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n5225) );
  INV_X1 U6684 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n9397) );
  OR2_X1 U6685 ( .A1(n5419), .A2(n9397), .ZN(n5224) );
  NAND2_X1 U6686 ( .A1(n5218), .A2(n5217), .ZN(n5219) );
  NAND2_X1 U6687 ( .A1(n5220), .A2(n5219), .ZN(n9396) );
  OR2_X1 U6688 ( .A1(n5466), .A2(n9396), .ZN(n5223) );
  INV_X1 U6689 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n5221) );
  OR2_X1 U6690 ( .A1(n5492), .A2(n5221), .ZN(n5222) );
  OR2_X1 U6691 ( .A1(n9408), .A2(n7697), .ZN(n5539) );
  NAND2_X1 U6692 ( .A1(n7799), .A2(n5539), .ZN(n5589) );
  INV_X1 U6693 ( .A(n5589), .ZN(n5227) );
  NAND2_X1 U6694 ( .A1(n7719), .A2(n9401), .ZN(n5588) );
  NAND2_X1 U6695 ( .A1(n9408), .A2(n7697), .ZN(n7797) );
  NAND2_X1 U6696 ( .A1(n5588), .A2(n7797), .ZN(n5226) );
  AOI22_X1 U6697 ( .A1(n5228), .A2(n5227), .B1(n7799), .B2(n5226), .ZN(n5235)
         );
  NAND2_X1 U6698 ( .A1(n9433), .A2(n7395), .ZN(n7582) );
  NAND2_X1 U6699 ( .A1(n7688), .A2(n7582), .ZN(n5568) );
  INV_X1 U6700 ( .A(n5568), .ZN(n5229) );
  NAND2_X1 U6701 ( .A1(n5230), .A2(n5229), .ZN(n5232) );
  INV_X1 U6702 ( .A(n7797), .ZN(n5231) );
  OAI21_X1 U6703 ( .B1(n5233), .B2(n5589), .A(n5588), .ZN(n5234) );
  XNOR2_X1 U6704 ( .A(n5237), .B(n5236), .ZN(n6442) );
  NAND2_X1 U6705 ( .A1(n6442), .A2(n5509), .ZN(n5244) );
  NOR2_X1 U6706 ( .A1(n5240), .A2(n4838), .ZN(n5238) );
  MUX2_X1 U6707 ( .A(n4838), .B(n5238), .S(P1_IR_REG_15__SCAN_IN), .Z(n5242)
         );
  NAND2_X1 U6708 ( .A1(n5240), .A2(n5239), .ZN(n5255) );
  INV_X1 U6709 ( .A(n5255), .ZN(n5241) );
  NOR2_X1 U6710 ( .A1(n5242), .A2(n5241), .ZN(n7533) );
  AOI22_X1 U6711 ( .A1(n5480), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n5303), .B2(
        n7533), .ZN(n5243) );
  NAND2_X1 U6712 ( .A1(n5484), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n5251) );
  INV_X1 U6713 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n7804) );
  OR2_X1 U6714 ( .A1(n5419), .A2(n7804), .ZN(n5250) );
  NOR2_X1 U6715 ( .A1(n5245), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n5246) );
  OR2_X1 U6716 ( .A1(n5260), .A2(n5246), .ZN(n8988) );
  OR2_X1 U6717 ( .A1(n5466), .A2(n8988), .ZN(n5249) );
  INV_X1 U6718 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n5247) );
  OR2_X1 U6719 ( .A1(n5492), .A2(n5247), .ZN(n5248) );
  NAND4_X1 U6720 ( .A1(n5251), .A2(n5250), .A3(n5249), .A4(n5248), .ZN(n9260)
         );
  XNOR2_X1 U6721 ( .A(n8074), .B(n9260), .ZN(n7800) );
  NAND2_X1 U6722 ( .A1(n5252), .A2(n7800), .ZN(n5270) );
  XNOR2_X1 U6723 ( .A(n5254), .B(n5253), .ZN(n6446) );
  NAND2_X1 U6724 ( .A1(n6446), .A2(n5509), .ZN(n5258) );
  NAND2_X1 U6725 ( .A1(n5255), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5256) );
  XNOR2_X1 U6726 ( .A(n5256), .B(P1_IR_REG_16__SCAN_IN), .ZN(n7728) );
  AOI22_X1 U6727 ( .A1(n5480), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n5303), .B2(
        n7728), .ZN(n5257) );
  NAND2_X1 U6728 ( .A1(n5484), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n5266) );
  INV_X1 U6729 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n5259) );
  OR2_X1 U6730 ( .A1(n5419), .A2(n5259), .ZN(n5265) );
  OR2_X1 U6731 ( .A1(n5260), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n5261) );
  NAND2_X1 U6732 ( .A1(n5279), .A2(n5261), .ZN(n9253) );
  OR2_X1 U6733 ( .A1(n5466), .A2(n9253), .ZN(n5264) );
  INV_X1 U6734 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n5262) );
  OR2_X1 U6735 ( .A1(n5492), .A2(n5262), .ZN(n5263) );
  OR2_X1 U6736 ( .A1(n9344), .A2(n8079), .ZN(n5593) );
  NAND2_X1 U6737 ( .A1(n9344), .A2(n8079), .ZN(n8103) );
  NAND2_X1 U6738 ( .A1(n5593), .A2(n8103), .ZN(n9249) );
  INV_X1 U6739 ( .A(n9260), .ZN(n8077) );
  NOR2_X1 U6740 ( .A1(n8074), .A2(n8077), .ZN(n8101) );
  NAND2_X1 U6741 ( .A1(n8074), .A2(n8077), .ZN(n8100) );
  INV_X1 U6742 ( .A(n8100), .ZN(n5267) );
  MUX2_X1 U6743 ( .A(n8101), .B(n5267), .S(n5483), .Z(n5268) );
  NOR2_X1 U6744 ( .A1(n9249), .A2(n5268), .ZN(n5269) );
  XNOR2_X1 U6745 ( .A(n5272), .B(n5271), .ZN(n6620) );
  NAND2_X1 U6746 ( .A1(n6620), .A2(n5509), .ZN(n5276) );
  NAND2_X1 U6747 ( .A1(n5273), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5274) );
  XNOR2_X1 U6748 ( .A(n5274), .B(P1_IR_REG_17__SCAN_IN), .ZN(n9039) );
  AOI22_X1 U6749 ( .A1(n5480), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n5303), .B2(
        n9039), .ZN(n5275) );
  NAND2_X1 U6750 ( .A1(n5484), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n5285) );
  INV_X1 U6751 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n5277) );
  OR2_X1 U6752 ( .A1(n5419), .A2(n5277), .ZN(n5284) );
  NAND2_X1 U6753 ( .A1(n5279), .A2(n5278), .ZN(n5280) );
  NAND2_X1 U6754 ( .A1(n5293), .A2(n5280), .ZN(n9237) );
  OR2_X1 U6755 ( .A1(n5466), .A2(n9237), .ZN(n5283) );
  INV_X1 U6756 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n5281) );
  OR2_X1 U6757 ( .A1(n5492), .A2(n5281), .ZN(n5282) );
  NAND4_X1 U6758 ( .A1(n5285), .A2(n5284), .A3(n5283), .A4(n5282), .ZN(n9262)
         );
  INV_X1 U6759 ( .A(n9262), .ZN(n8081) );
  OR2_X1 U6760 ( .A1(n9339), .A2(n8081), .ZN(n9224) );
  NAND2_X1 U6761 ( .A1(n9339), .A2(n8081), .ZN(n8104) );
  AND2_X1 U6762 ( .A1(n9224), .A2(n8104), .ZN(n9242) );
  MUX2_X1 U6763 ( .A(n5593), .B(n8103), .S(n9278), .Z(n5286) );
  XNOR2_X1 U6764 ( .A(n5288), .B(n5287), .ZN(n6776) );
  NAND2_X1 U6765 ( .A1(n6776), .A2(n5509), .ZN(n5291) );
  NAND2_X1 U6766 ( .A1(n4332), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5289) );
  XNOR2_X1 U6767 ( .A(n5289), .B(P1_IR_REG_18__SCAN_IN), .ZN(n9055) );
  AOI22_X1 U6768 ( .A1(n5480), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n5303), .B2(
        n9055), .ZN(n5290) );
  NAND2_X1 U6769 ( .A1(n4278), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n5299) );
  INV_X1 U6770 ( .A(P1_REG0_REG_18__SCAN_IN), .ZN(n5292) );
  OR2_X1 U6771 ( .A1(n5019), .A2(n5292), .ZN(n5298) );
  NAND2_X1 U6772 ( .A1(n5293), .A2(n10003), .ZN(n5295) );
  INV_X1 U6773 ( .A(n5307), .ZN(n5294) );
  NAND2_X1 U6774 ( .A1(n5295), .A2(n5294), .ZN(n9221) );
  OR2_X1 U6775 ( .A1(n5466), .A2(n9221), .ZN(n5297) );
  INV_X1 U6776 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n9034) );
  OR2_X1 U6777 ( .A1(n5492), .A2(n9034), .ZN(n5296) );
  NAND2_X1 U6778 ( .A1(n9334), .A2(n8928), .ZN(n8105) );
  AND2_X1 U6779 ( .A1(n8105), .A2(n8104), .ZN(n5300) );
  MUX2_X1 U6780 ( .A(n8107), .B(n5300), .S(n5483), .Z(n5301) );
  NAND2_X1 U6781 ( .A1(n5302), .A2(n5301), .ZN(n5377) );
  XNOR2_X1 U6782 ( .A(n5345), .B(n5344), .ZN(n6890) );
  NAND2_X1 U6783 ( .A1(n6890), .A2(n5509), .ZN(n5305) );
  AOI22_X1 U6784 ( .A1(n5480), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n9592), .B2(
        n5303), .ZN(n5304) );
  NAND2_X1 U6785 ( .A1(n5484), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n5311) );
  INV_X1 U6786 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n9053) );
  OR2_X1 U6787 ( .A1(n5419), .A2(n9053), .ZN(n5310) );
  INV_X1 U6788 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n9986) );
  OR2_X1 U6789 ( .A1(n5492), .A2(n9986), .ZN(n5309) );
  OAI21_X1 U6790 ( .B1(P1_REG3_REG_19__SCAN_IN), .B2(n5307), .A(n5306), .ZN(
        n9208) );
  OR2_X1 U6791 ( .A1(n5466), .A2(n9208), .ZN(n5308) );
  NAND4_X1 U6792 ( .A1(n5311), .A2(n5310), .A3(n5309), .A4(n5308), .ZN(n9228)
         );
  INV_X1 U6793 ( .A(n9228), .ZN(n8962) );
  NAND2_X1 U6794 ( .A1(n9329), .A2(n8962), .ZN(n8108) );
  NAND2_X1 U6795 ( .A1(n8108), .A2(n8105), .ZN(n5577) );
  INV_X1 U6796 ( .A(n5577), .ZN(n5312) );
  AND2_X1 U6797 ( .A1(n5377), .A2(n5312), .ZN(n5376) );
  OR2_X1 U6798 ( .A1(n5345), .A2(n5313), .ZN(n5315) );
  NAND2_X1 U6799 ( .A1(n7003), .A2(n5509), .ZN(n5319) );
  NAND2_X1 U6800 ( .A1(n5480), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n5318) );
  NAND2_X1 U6801 ( .A1(n5484), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n5327) );
  INV_X1 U6802 ( .A(P1_REG2_REG_22__SCAN_IN), .ZN(n5320) );
  OR2_X1 U6803 ( .A1(n5419), .A2(n5320), .ZN(n5326) );
  INV_X1 U6804 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n5321) );
  NAND2_X1 U6805 ( .A1(n5338), .A2(n5321), .ZN(n5322) );
  NAND2_X1 U6806 ( .A1(n5369), .A2(n5322), .ZN(n9164) );
  OR2_X1 U6807 ( .A1(n5466), .A2(n9164), .ZN(n5325) );
  INV_X1 U6808 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n5323) );
  OR2_X1 U6809 ( .A1(n5492), .A2(n5323), .ZN(n5324) );
  NAND4_X1 U6810 ( .A1(n5327), .A2(n5326), .A3(n5325), .A4(n5324), .ZN(n9187)
         );
  INV_X1 U6811 ( .A(n9187), .ZN(n8089) );
  OR2_X1 U6812 ( .A1(n9314), .A2(n8089), .ZN(n5534) );
  OR2_X1 U6813 ( .A1(n5345), .A2(n5328), .ZN(n5330) );
  NAND2_X1 U6814 ( .A1(n6974), .A2(n5509), .ZN(n5334) );
  NAND2_X1 U6815 ( .A1(n5480), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n5333) );
  NAND2_X1 U6816 ( .A1(n5484), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n5343) );
  INV_X1 U6817 ( .A(P1_REG2_REG_21__SCAN_IN), .ZN(n5335) );
  OR2_X1 U6818 ( .A1(n5419), .A2(n5335), .ZN(n5342) );
  INV_X1 U6819 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n5336) );
  NAND2_X1 U6820 ( .A1(n5354), .A2(n5336), .ZN(n5337) );
  NAND2_X1 U6821 ( .A1(n5338), .A2(n5337), .ZN(n9181) );
  OR2_X1 U6822 ( .A1(n5466), .A2(n9181), .ZN(n5341) );
  INV_X1 U6823 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n5339) );
  OR2_X1 U6824 ( .A1(n5492), .A2(n5339), .ZN(n5340) );
  OR2_X1 U6825 ( .A1(n5345), .A2(n5344), .ZN(n5347) );
  INV_X1 U6826 ( .A(n5348), .ZN(n5349) );
  NAND2_X1 U6827 ( .A1(n6972), .A2(n5509), .ZN(n5352) );
  NAND2_X1 U6828 ( .A1(n5480), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n5351) );
  NAND2_X1 U6829 ( .A1(n5484), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n5360) );
  INV_X1 U6830 ( .A(P1_REG2_REG_20__SCAN_IN), .ZN(n5353) );
  OR2_X1 U6831 ( .A1(n5419), .A2(n5353), .ZN(n5359) );
  OAI21_X1 U6832 ( .B1(P1_REG3_REG_20__SCAN_IN), .B2(n5355), .A(n5354), .ZN(
        n9194) );
  OR2_X1 U6833 ( .A1(n5466), .A2(n9194), .ZN(n5358) );
  INV_X1 U6834 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n5356) );
  OR2_X1 U6835 ( .A1(n5492), .A2(n5356), .ZN(n5357) );
  NAND4_X1 U6836 ( .A1(n5360), .A2(n5359), .A3(n5358), .A4(n5357), .ZN(n9213)
         );
  INV_X1 U6837 ( .A(n9213), .ZN(n8902) );
  OR2_X1 U6838 ( .A1(n9329), .A2(n8962), .ZN(n5537) );
  AND2_X1 U6839 ( .A1(n8109), .A2(n5537), .ZN(n5361) );
  NAND2_X1 U6840 ( .A1(n8113), .A2(n5361), .ZN(n5580) );
  NAND2_X1 U6841 ( .A1(n9168), .A2(n8110), .ZN(n5557) );
  NAND2_X1 U6842 ( .A1(n9319), .A2(n8087), .ZN(n8111) );
  NAND2_X1 U6843 ( .A1(n5557), .A2(n8111), .ZN(n5362) );
  OR2_X1 U6844 ( .A1(n8112), .A2(n5362), .ZN(n5363) );
  NAND2_X1 U6845 ( .A1(n5363), .A2(n5534), .ZN(n5578) );
  NAND2_X1 U6846 ( .A1(n7060), .A2(n5509), .ZN(n5367) );
  NAND2_X1 U6847 ( .A1(n5480), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n5366) );
  NAND2_X1 U6848 ( .A1(n5484), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n5375) );
  INV_X1 U6849 ( .A(P1_REG2_REG_23__SCAN_IN), .ZN(n9150) );
  OR2_X1 U6850 ( .A1(n5419), .A2(n9150), .ZN(n5374) );
  INV_X1 U6851 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n5368) );
  NAND2_X1 U6852 ( .A1(n5369), .A2(n5368), .ZN(n5370) );
  NAND2_X1 U6853 ( .A1(n5391), .A2(n5370), .ZN(n9157) );
  OR2_X1 U6854 ( .A1(n5466), .A2(n9157), .ZN(n5373) );
  INV_X1 U6855 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n5371) );
  OR2_X1 U6856 ( .A1(n5492), .A2(n5371), .ZN(n5372) );
  NAND4_X1 U6857 ( .A1(n5375), .A2(n5374), .A3(n5373), .A4(n5372), .ZN(n9172)
         );
  INV_X1 U6858 ( .A(n9172), .ZN(n8090) );
  NAND2_X1 U6859 ( .A1(n9308), .A2(n8090), .ZN(n8114) );
  OAI211_X1 U6860 ( .C1(n5376), .C2(n5580), .A(n5578), .B(n8114), .ZN(n5384)
         );
  INV_X1 U6861 ( .A(n8110), .ZN(n5536) );
  NAND3_X1 U6862 ( .A1(n5378), .A2(n5536), .A3(n8108), .ZN(n5379) );
  NAND2_X1 U6863 ( .A1(n5379), .A2(n8109), .ZN(n5381) );
  INV_X1 U6864 ( .A(n8113), .ZN(n5380) );
  INV_X1 U6865 ( .A(n8115), .ZN(n5403) );
  OAI21_X1 U6866 ( .B1(n5382), .B2(n8112), .A(n5403), .ZN(n5383) );
  NAND2_X1 U6867 ( .A1(n7163), .A2(n5509), .ZN(n5388) );
  NAND2_X1 U6868 ( .A1(n5480), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n5387) );
  NAND2_X1 U6869 ( .A1(n4278), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n5398) );
  INV_X1 U6870 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n5389) );
  OR2_X1 U6871 ( .A1(n5492), .A2(n5389), .ZN(n5397) );
  INV_X1 U6872 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n5390) );
  NAND2_X1 U6873 ( .A1(n5391), .A2(n5390), .ZN(n5392) );
  NAND2_X1 U6874 ( .A1(n5393), .A2(n5392), .ZN(n9143) );
  OR2_X1 U6875 ( .A1(n5466), .A2(n9143), .ZN(n5396) );
  INV_X1 U6876 ( .A(P1_REG0_REG_24__SCAN_IN), .ZN(n5394) );
  OR2_X1 U6877 ( .A1(n5019), .A2(n5394), .ZN(n5395) );
  NAND4_X1 U6878 ( .A1(n5398), .A2(n5397), .A3(n5396), .A4(n5395), .ZN(n9155)
         );
  AND2_X1 U6879 ( .A1(n5402), .A2(n9155), .ZN(n8092) );
  INV_X1 U6880 ( .A(n8092), .ZN(n5399) );
  OR2_X1 U6881 ( .A1(n5402), .A2(n9155), .ZN(n8093) );
  AND2_X1 U6882 ( .A1(n5399), .A2(n8093), .ZN(n9134) );
  NAND2_X1 U6883 ( .A1(n9299), .A2(n8977), .ZN(n8119) );
  INV_X1 U6884 ( .A(n9155), .ZN(n7917) );
  NAND2_X1 U6885 ( .A1(n8119), .A2(n5404), .ZN(n5606) );
  INV_X1 U6886 ( .A(n5606), .ZN(n5401) );
  NAND2_X1 U6887 ( .A1(n5401), .A2(n5400), .ZN(n5406) );
  OR2_X1 U6888 ( .A1(n5402), .A2(n7917), .ZN(n8116) );
  OAI21_X1 U6889 ( .B1(n5408), .B2(n9134), .A(n5407), .ZN(n5430) );
  INV_X1 U6890 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n9932) );
  INV_X1 U6891 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n7542) );
  MUX2_X1 U6892 ( .A(n9932), .B(n7542), .S(n4280), .Z(n5413) );
  INV_X1 U6893 ( .A(SI_26_), .ZN(n5412) );
  NAND2_X1 U6894 ( .A1(n5413), .A2(n5412), .ZN(n5437) );
  INV_X1 U6895 ( .A(n5413), .ZN(n5414) );
  NAND2_X1 U6896 ( .A1(n5414), .A2(SI_26_), .ZN(n5415) );
  AND2_X1 U6897 ( .A1(n5437), .A2(n5415), .ZN(n5435) );
  NAND2_X1 U6898 ( .A1(n7995), .A2(n5509), .ZN(n5417) );
  NAND2_X1 U6899 ( .A1(n5480), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n5416) );
  NAND2_X1 U6900 ( .A1(n5484), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n5427) );
  INV_X1 U6901 ( .A(P1_REG2_REG_26__SCAN_IN), .ZN(n5418) );
  OR2_X1 U6902 ( .A1(n5419), .A2(n5418), .ZN(n5426) );
  INV_X1 U6903 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n5420) );
  NAND2_X1 U6904 ( .A1(n5421), .A2(n5420), .ZN(n5422) );
  NAND2_X1 U6905 ( .A1(n5448), .A2(n5422), .ZN(n8975) );
  OR2_X1 U6906 ( .A1(n5466), .A2(n8975), .ZN(n5425) );
  INV_X1 U6907 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n5423) );
  OR2_X1 U6908 ( .A1(n5492), .A2(n5423), .ZN(n5424) );
  XNOR2_X1 U6909 ( .A(n9111), .B(n8094), .ZN(n5429) );
  NAND2_X1 U6910 ( .A1(n4520), .A2(n9278), .ZN(n5428) );
  INV_X1 U6911 ( .A(n8121), .ZN(n5431) );
  OAI21_X1 U6912 ( .B1(n9278), .B2(n8118), .A(n5434), .ZN(n5456) );
  INV_X1 U6913 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n10021) );
  INV_X1 U6914 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n5439) );
  MUX2_X1 U6915 ( .A(n10021), .B(n5439), .S(n4279), .Z(n5441) );
  INV_X1 U6916 ( .A(SI_27_), .ZN(n5440) );
  NAND2_X1 U6917 ( .A1(n5441), .A2(n5440), .ZN(n5459) );
  INV_X1 U6918 ( .A(n5441), .ZN(n5442) );
  NAND2_X1 U6919 ( .A1(n5442), .A2(SI_27_), .ZN(n5443) );
  AND2_X1 U6920 ( .A1(n5459), .A2(n5443), .ZN(n5457) );
  NAND2_X1 U6921 ( .A1(n8010), .A2(n5509), .ZN(n5445) );
  NAND2_X1 U6922 ( .A1(n5480), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n5444) );
  NAND2_X1 U6923 ( .A1(n4278), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n5454) );
  INV_X1 U6924 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n5446) );
  OR2_X1 U6925 ( .A1(n5019), .A2(n5446), .ZN(n5453) );
  INV_X1 U6926 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n5447) );
  NAND2_X1 U6927 ( .A1(n5448), .A2(n5447), .ZN(n5449) );
  NAND2_X1 U6928 ( .A1(n5464), .A2(n5449), .ZN(n9096) );
  OR2_X1 U6929 ( .A1(n5466), .A2(n9096), .ZN(n5452) );
  INV_X1 U6930 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n5450) );
  OR2_X1 U6931 ( .A1(n5492), .A2(n5450), .ZN(n5451) );
  NAND2_X1 U6932 ( .A1(n9289), .A2(n10020), .ZN(n5610) );
  NAND2_X1 U6933 ( .A1(n8120), .A2(n5483), .ZN(n5455) );
  MUX2_X1 U6934 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(P2_DATAO_REG_28__SCAN_IN), 
        .S(n4280), .Z(n5477) );
  INV_X1 U6935 ( .A(SI_28_), .ZN(n9900) );
  XNOR2_X1 U6936 ( .A(n5477), .B(n9900), .ZN(n5475) );
  NAND2_X1 U6937 ( .A1(n8023), .A2(n5509), .ZN(n5462) );
  NAND2_X1 U6938 ( .A1(n5480), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n5461) );
  NAND2_X1 U6939 ( .A1(n4278), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n5471) );
  INV_X1 U6940 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n9946) );
  OR2_X1 U6941 ( .A1(n5019), .A2(n9946), .ZN(n5470) );
  INV_X1 U6942 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n5463) );
  NAND2_X1 U6943 ( .A1(n5464), .A2(n5463), .ZN(n5465) );
  NAND2_X1 U6944 ( .A1(n8133), .A2(n5465), .ZN(n9078) );
  OR2_X1 U6945 ( .A1(n5466), .A2(n9078), .ZN(n5469) );
  INV_X1 U6946 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n5467) );
  OR2_X1 U6947 ( .A1(n5492), .A2(n5467), .ZN(n5468) );
  MUX2_X1 U6948 ( .A(n5610), .B(n9082), .S(n5483), .Z(n5472) );
  MUX2_X1 U6949 ( .A(n8122), .B(n5612), .S(n9278), .Z(n5473) );
  INV_X1 U6950 ( .A(n5477), .ZN(n5478) );
  MUX2_X1 U6951 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(P2_DATAO_REG_29__SCAN_IN), 
        .S(n4280), .Z(n5493) );
  INV_X1 U6952 ( .A(SI_29_), .ZN(n5495) );
  XNOR2_X1 U6953 ( .A(n5493), .B(n5495), .ZN(n5479) );
  NAND2_X1 U6954 ( .A1(n8142), .A2(n5509), .ZN(n5482) );
  NAND2_X1 U6955 ( .A1(n5480), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n5481) );
  INV_X1 U6956 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n5487) );
  NAND2_X1 U6957 ( .A1(n4278), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n5486) );
  NAND2_X1 U6958 ( .A1(n5484), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n5485) );
  OAI211_X1 U6959 ( .C1(n5492), .C2(n5487), .A(n5486), .B(n5485), .ZN(n8998)
         );
  INV_X1 U6960 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n5491) );
  NAND2_X1 U6961 ( .A1(n4278), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n5490) );
  INV_X1 U6962 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n5488) );
  OR2_X1 U6963 ( .A1(n5019), .A2(n5488), .ZN(n5489) );
  OAI211_X1 U6964 ( .C1(n5492), .C2(n5491), .A(n5490), .B(n5489), .ZN(n9066)
         );
  NAND2_X1 U6965 ( .A1(n5494), .A2(n5493), .ZN(n5497) );
  NAND2_X1 U6966 ( .A1(n5497), .A2(n4305), .ZN(n5503) );
  MUX2_X1 U6967 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(P1_DATAO_REG_30__SCAN_IN), 
        .S(n4499), .Z(n5502) );
  INV_X1 U6968 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n7856) );
  OR2_X1 U6969 ( .A1(n5030), .A2(n7856), .ZN(n5498) );
  INV_X1 U6970 ( .A(n8998), .ZN(n5532) );
  OR2_X1 U6971 ( .A1(n9070), .A2(n5532), .ZN(n5530) );
  INV_X1 U6972 ( .A(n5530), .ZN(n5512) );
  INV_X1 U6973 ( .A(n9066), .ZN(n5515) );
  INV_X1 U6974 ( .A(n5500), .ZN(n5501) );
  NAND2_X1 U6975 ( .A1(n5501), .A2(SI_30_), .ZN(n5505) );
  NAND2_X1 U6976 ( .A1(n5503), .A2(n5502), .ZN(n5504) );
  NAND2_X1 U6977 ( .A1(n5505), .A2(n5504), .ZN(n5508) );
  MUX2_X1 U6978 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n4499), .Z(n5506) );
  XNOR2_X1 U6979 ( .A(n5506), .B(SI_31_), .ZN(n5507) );
  INV_X1 U6980 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n5510) );
  OR2_X1 U6981 ( .A1(n5030), .A2(n5510), .ZN(n5511) );
  NAND2_X1 U6982 ( .A1(n5514), .A2(n9087), .ZN(n5513) );
  OAI21_X1 U6983 ( .B1(n5619), .B2(n5513), .A(n5617), .ZN(n5521) );
  INV_X1 U6984 ( .A(n5619), .ZN(n5518) );
  INV_X1 U6985 ( .A(n5531), .ZN(n5517) );
  AOI21_X1 U6986 ( .B1(n5519), .B2(n5518), .A(n5517), .ZN(n5520) );
  AOI21_X1 U6987 ( .B1(n5523), .B2(n5617), .A(n5522), .ZN(n5529) );
  NAND2_X1 U6988 ( .A1(n6387), .A2(n9592), .ZN(n6784) );
  OR2_X1 U6989 ( .A1(n5525), .A2(n5524), .ZN(n5526) );
  NOR2_X1 U6990 ( .A1(n5661), .A2(n6976), .ZN(n5621) );
  INV_X1 U6991 ( .A(n5621), .ZN(n5528) );
  AOI21_X1 U6992 ( .B1(n5529), .B2(n6784), .A(n5528), .ZN(n5625) );
  NAND2_X1 U6993 ( .A1(n5531), .A2(n5530), .ZN(n5660) );
  AND2_X1 U6994 ( .A1(n9070), .A2(n5532), .ZN(n5627) );
  NOR2_X1 U6995 ( .A1(n9281), .A2(n7947), .ZN(n5614) );
  INV_X1 U6996 ( .A(n8120), .ZN(n5533) );
  NAND2_X1 U6997 ( .A1(n8121), .A2(n5533), .ZN(n9113) );
  NOR2_X1 U6998 ( .A1(n8115), .A2(n4530), .ZN(n9153) );
  INV_X1 U6999 ( .A(n8112), .ZN(n5535) );
  AND2_X1 U7000 ( .A1(n5535), .A2(n5534), .ZN(n9171) );
  INV_X1 U7001 ( .A(n9185), .ZN(n5551) );
  NAND2_X1 U7002 ( .A1(n5536), .A2(n8109), .ZN(n9199) );
  NAND2_X1 U7003 ( .A1(n5537), .A2(n8108), .ZN(n9211) );
  NAND2_X1 U7004 ( .A1(n5538), .A2(n8105), .ZN(n9226) );
  INV_X1 U7005 ( .A(n9249), .ZN(n9258) );
  NAND2_X1 U7006 ( .A1(n7799), .A2(n5588), .ZN(n7795) );
  INV_X1 U7007 ( .A(n9400), .ZN(n9390) );
  INV_X1 U7008 ( .A(n6781), .ZN(n5540) );
  NAND2_X1 U7009 ( .A1(n6360), .A2(n6794), .ZN(n5633) );
  NAND2_X1 U7010 ( .A1(n5540), .A2(n5633), .ZN(n6382) );
  NOR4_X1 U7011 ( .A1(n6382), .A2(n6930), .A3(n6943), .A4(n6911), .ZN(n5542)
         );
  NAND4_X1 U7012 ( .A1(n5542), .A2(n9596), .A3(n6952), .A4(n6782), .ZN(n5544)
         );
  NAND2_X1 U7013 ( .A1(n5562), .A2(n5543), .ZN(n7415) );
  NOR4_X1 U7014 ( .A1(n5544), .A2(n7486), .A3(n7406), .A4(n7415), .ZN(n5545)
         );
  NAND3_X1 U7015 ( .A1(n5545), .A2(n7419), .A3(n9411), .ZN(n5547) );
  NAND2_X1 U7016 ( .A1(n5546), .A2(n7688), .ZN(n7584) );
  NOR4_X1 U7017 ( .A1(n7795), .A2(n9390), .A3(n5547), .A4(n7584), .ZN(n5548)
         );
  NAND4_X1 U7018 ( .A1(n9242), .A2(n9258), .A3(n5548), .A4(n7800), .ZN(n5549)
         );
  NOR4_X1 U7019 ( .A1(n9199), .A2(n9211), .A3(n9226), .A4(n5549), .ZN(n5550)
         );
  NAND4_X1 U7020 ( .A1(n9153), .A2(n9171), .A3(n5551), .A4(n5550), .ZN(n5552)
         );
  NOR4_X1 U7021 ( .A1(n9113), .A2(n9134), .A3(n9126), .A4(n5552), .ZN(n5553)
         );
  NAND4_X1 U7022 ( .A1(n8123), .A2(n9092), .A3(n9085), .A4(n5553), .ZN(n5554)
         );
  INV_X1 U7023 ( .A(n6976), .ZN(n6201) );
  NOR2_X1 U7024 ( .A1(n5555), .A2(n6201), .ZN(n5623) );
  NOR2_X1 U7025 ( .A1(n5606), .A2(n4530), .ZN(n5631) );
  INV_X1 U7026 ( .A(n5638), .ZN(n5605) );
  AND4_X1 U7027 ( .A1(n8108), .A2(n8105), .A3(n8103), .A4(n8104), .ZN(n5556)
         );
  NAND3_X1 U7028 ( .A1(n5557), .A2(n5556), .A3(n8111), .ZN(n5558) );
  NOR2_X1 U7029 ( .A1(n8112), .A2(n5558), .ZN(n5595) );
  INV_X1 U7030 ( .A(n5595), .ZN(n5572) );
  INV_X1 U7031 ( .A(n6904), .ZN(n5561) );
  AND2_X1 U7032 ( .A1(n5600), .A2(n5559), .ZN(n5635) );
  NAND2_X1 U7033 ( .A1(n4516), .A2(n5574), .ZN(n5560) );
  AND2_X1 U7034 ( .A1(n5560), .A2(n5601), .ZN(n5639) );
  NAND3_X1 U7035 ( .A1(n5561), .A2(n5635), .A3(n5639), .ZN(n5564) );
  NAND4_X1 U7036 ( .A1(n7797), .A2(n5564), .A3(n5563), .A4(n5562), .ZN(n5569)
         );
  NAND2_X1 U7037 ( .A1(n7578), .A2(n5565), .ZN(n5566) );
  AND2_X1 U7038 ( .A1(n5566), .A2(n7580), .ZN(n5567) );
  OR2_X1 U7039 ( .A1(n5568), .A2(n5567), .ZN(n5586) );
  NOR2_X1 U7040 ( .A1(n5569), .A2(n5586), .ZN(n5570) );
  NAND3_X1 U7041 ( .A1(n8100), .A2(n5570), .A3(n5588), .ZN(n5571) );
  NOR2_X1 U7042 ( .A1(n5572), .A2(n5571), .ZN(n5641) );
  INV_X1 U7043 ( .A(n5641), .ZN(n5576) );
  NAND2_X1 U7044 ( .A1(n5574), .A2(n5573), .ZN(n5598) );
  OR3_X1 U7045 ( .A1(n5576), .A2(n5575), .A3(n5598), .ZN(n5644) );
  NOR2_X1 U7046 ( .A1(n5577), .A2(n8107), .ZN(n5579) );
  OAI21_X1 U7047 ( .B1(n5580), .B2(n5579), .A(n5578), .ZN(n5597) );
  INV_X1 U7048 ( .A(n8101), .ZN(n5592) );
  INV_X1 U7049 ( .A(n5581), .ZN(n5582) );
  NOR2_X1 U7050 ( .A1(n5583), .A2(n5582), .ZN(n5585) );
  INV_X1 U7051 ( .A(n7688), .ZN(n5584) );
  OAI22_X1 U7052 ( .A1(n5586), .A2(n5585), .B1(n7686), .B2(n5584), .ZN(n5587)
         );
  AND2_X1 U7053 ( .A1(n5587), .A2(n7797), .ZN(n5590) );
  OAI211_X1 U7054 ( .C1(n5590), .C2(n5589), .A(n8100), .B(n5588), .ZN(n5591)
         );
  NAND3_X1 U7055 ( .A1(n5593), .A2(n5592), .A3(n5591), .ZN(n5594) );
  NAND2_X1 U7056 ( .A1(n5595), .A2(n5594), .ZN(n5596) );
  AND2_X1 U7057 ( .A1(n5597), .A2(n5596), .ZN(n5643) );
  AOI21_X1 U7058 ( .B1(n5600), .B2(n5599), .A(n5598), .ZN(n5603) );
  INV_X1 U7059 ( .A(n5601), .ZN(n5602) );
  OAI21_X1 U7060 ( .B1(n5603), .B2(n5602), .A(n5641), .ZN(n5604) );
  OAI211_X1 U7061 ( .C1(n5605), .C2(n5644), .A(n5643), .B(n5604), .ZN(n5609)
         );
  OAI211_X1 U7062 ( .C1(n5607), .C2(n5606), .A(n8121), .B(n8118), .ZN(n5650)
         );
  INV_X1 U7063 ( .A(n9082), .ZN(n5608) );
  AOI211_X1 U7064 ( .C1(n5631), .C2(n5609), .A(n5650), .B(n5608), .ZN(n5611)
         );
  AND2_X1 U7065 ( .A1(n9082), .A2(n8120), .ZN(n5630) );
  NAND2_X1 U7066 ( .A1(n8122), .A2(n5610), .ZN(n5629) );
  NOR3_X1 U7067 ( .A1(n5611), .A2(n5630), .A3(n5629), .ZN(n5616) );
  INV_X1 U7068 ( .A(n5612), .ZN(n5613) );
  OR2_X1 U7069 ( .A1(n5614), .A2(n5613), .ZN(n5628) );
  INV_X1 U7070 ( .A(n5654), .ZN(n5615) );
  OAI21_X1 U7071 ( .B1(n5616), .B2(n5628), .A(n5615), .ZN(n5618) );
  OAI21_X1 U7072 ( .B1(n5619), .B2(n5618), .A(n5617), .ZN(n5620) );
  AOI21_X1 U7073 ( .B1(n5621), .B2(n5620), .A(n5623), .ZN(n5622) );
  MUX2_X1 U7074 ( .A(n5623), .B(n5622), .S(n9141), .Z(n5624) );
  XNOR2_X1 U7075 ( .A(n5626), .B(P1_IR_REG_20__SCAN_IN), .ZN(n9277) );
  INV_X1 U7076 ( .A(n5627), .ZN(n5658) );
  INV_X1 U7077 ( .A(n5628), .ZN(n5656) );
  INV_X1 U7078 ( .A(n5629), .ZN(n5653) );
  INV_X1 U7079 ( .A(n5630), .ZN(n5652) );
  INV_X1 U7080 ( .A(n5631), .ZN(n5648) );
  NAND2_X1 U7081 ( .A1(n6897), .A2(n6795), .ZN(n5632) );
  NAND4_X1 U7082 ( .A1(n5634), .A2(n5633), .A3(n6201), .A4(n5632), .ZN(n5637)
         );
  INV_X1 U7083 ( .A(n5635), .ZN(n5636) );
  AOI21_X1 U7084 ( .B1(n5638), .B2(n5637), .A(n5636), .ZN(n5645) );
  INV_X1 U7085 ( .A(n5639), .ZN(n5640) );
  NAND2_X1 U7086 ( .A1(n5641), .A2(n5640), .ZN(n5642) );
  OAI211_X1 U7087 ( .C1(n5645), .C2(n5644), .A(n5643), .B(n5642), .ZN(n5646)
         );
  INV_X1 U7088 ( .A(n5646), .ZN(n5647) );
  NOR2_X1 U7089 ( .A1(n5648), .A2(n5647), .ZN(n5649) );
  OR3_X1 U7090 ( .A1(n9100), .A2(n5650), .A3(n5649), .ZN(n5651) );
  NAND3_X1 U7091 ( .A1(n5653), .A2(n5652), .A3(n5651), .ZN(n5655) );
  AOI21_X1 U7092 ( .B1(n5656), .B2(n5655), .A(n5654), .ZN(n5657) );
  AND2_X1 U7093 ( .A1(n5658), .A2(n5657), .ZN(n5659) );
  OR2_X1 U7094 ( .A1(n5660), .A2(n5659), .ZN(n5663) );
  INV_X1 U7095 ( .A(n5661), .ZN(n5662) );
  NOR2_X1 U7096 ( .A1(n5666), .A2(n9141), .ZN(n5665) );
  INV_X1 U7097 ( .A(n9277), .ZN(n5664) );
  INV_X1 U7098 ( .A(n5666), .ZN(n5669) );
  AND2_X1 U7099 ( .A1(n5664), .A2(n9141), .ZN(n6354) );
  INV_X1 U7100 ( .A(n6354), .ZN(n6760) );
  NAND2_X1 U7101 ( .A1(n5667), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5668) );
  XNOR2_X1 U7102 ( .A(n5668), .B(n4777), .ZN(n6352) );
  OR2_X1 U7103 ( .A1(n6352), .A2(P1_U3084), .ZN(n5685) );
  INV_X1 U7104 ( .A(n5685), .ZN(n7013) );
  OAI21_X1 U7105 ( .B1(n5669), .B2(n6760), .A(n7013), .ZN(n5670) );
  NAND2_X1 U7106 ( .A1(n5677), .A2(n5676), .ZN(n5673) );
  XNOR2_X1 U7107 ( .A(n5677), .B(n5676), .ZN(n7459) );
  NAND2_X1 U7108 ( .A1(n4318), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5679) );
  XNOR2_X1 U7109 ( .A(n5679), .B(n5678), .ZN(n7165) );
  AND2_X1 U7110 ( .A1(n6352), .A2(P1_STATE_REG_SCAN_IN), .ZN(n5681) );
  INV_X1 U7111 ( .A(n5682), .ZN(n6786) );
  INV_X1 U7112 ( .A(n5683), .ZN(n8124) );
  NAND4_X1 U7113 ( .A1(n9602), .A2(n4344), .A3(n6786), .A4(n8124), .ZN(n5684)
         );
  OAI211_X1 U7114 ( .C1(n6387), .C2(n5685), .A(n5684), .B(P1_B_REG_SCAN_IN), 
        .ZN(n5686) );
  NOR2_X2 U7115 ( .A1(n5781), .A2(P2_IR_REG_5__SCAN_IN), .ZN(n5808) );
  NOR2_X1 U7116 ( .A1(P2_IR_REG_9__SCAN_IN), .A2(P2_IR_REG_13__SCAN_IN), .ZN(
        n5689) );
  NAND4_X1 U7117 ( .A1(n5689), .A2(n5688), .A3(n5839), .A4(n5914), .ZN(n5693)
         );
  INV_X1 U7118 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n5691) );
  INV_X1 U7119 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n5690) );
  NAND4_X1 U7120 ( .A1(n5691), .A2(n5980), .A3(n5861), .A4(n5690), .ZN(n5692)
         );
  NOR2_X1 U7121 ( .A1(n5693), .A2(n5692), .ZN(n5694) );
  INV_X1 U7122 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n6159) );
  INV_X1 U7123 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n5695) );
  INV_X1 U7124 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n6017) );
  NAND4_X1 U7125 ( .A1(n6134), .A2(n5695), .A3(n4724), .A4(n6017), .ZN(n5696)
         );
  NOR2_X1 U7126 ( .A1(n5697), .A2(n5696), .ZN(n5698) );
  INV_X1 U7127 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n5699) );
  NAND2_X1 U7128 ( .A1(n5702), .A2(n5700), .ZN(n8874) );
  AND2_X2 U7129 ( .A1(n5741), .A2(n7781), .ZN(n5788) );
  NAND2_X1 U7130 ( .A1(n5788), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n5705) );
  INV_X1 U7131 ( .A(n5741), .ZN(n5707) );
  AND2_X2 U7132 ( .A1(n5707), .A2(n7781), .ZN(n5823) );
  NAND2_X1 U7133 ( .A1(n5823), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n5704) );
  NAND2_X1 U7134 ( .A1(n5828), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n5709) );
  NAND2_X1 U7135 ( .A1(n4499), .A2(SI_0_), .ZN(n5712) );
  INV_X1 U7136 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n5711) );
  NAND2_X1 U7137 ( .A1(n5712), .A2(n5711), .ZN(n5714) );
  AND2_X1 U7138 ( .A1(n5714), .A2(n5713), .ZN(n8881) );
  NAND2_X2 U7139 ( .A1(n5720), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5717) );
  INV_X1 U7140 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n5716) );
  NAND2_X1 U7141 ( .A1(n5718), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5719) );
  NAND2_X2 U7142 ( .A1(n6183), .A2(n8407), .ZN(n5753) );
  MUX2_X1 U7143 ( .A(P2_IR_REG_0__SCAN_IN), .B(n8881), .S(n5753), .Z(n9761) );
  OAI21_X2 U7144 ( .B1(n5725), .B2(P2_IR_REG_21__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n6135) );
  XNOR2_X2 U7145 ( .A(n6135), .B(n6134), .ZN(n7951) );
  NAND2_X1 U7146 ( .A1(n5729), .A2(n4587), .ZN(n5727) );
  XNOR2_X2 U7147 ( .A(n5728), .B(P2_IR_REG_20__SCAN_IN), .ZN(n8373) );
  NAND2_X1 U7148 ( .A1(n5732), .A2(n8165), .ZN(n6732) );
  INV_X1 U7149 ( .A(n7951), .ZN(n8383) );
  NAND2_X1 U7150 ( .A1(n7117), .A2(n8372), .ZN(n8339) );
  NAND2_X1 U7151 ( .A1(n5733), .A2(n8373), .ZN(n8166) );
  OR2_X4 U7152 ( .A1(n8339), .A2(n8167), .ZN(n8035) );
  NAND2_X1 U7153 ( .A1(n6733), .A2(n8035), .ZN(n5734) );
  AND2_X1 U7154 ( .A1(n6732), .A2(n5734), .ZN(n6580) );
  NAND2_X1 U7155 ( .A1(n5819), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n5740) );
  AND2_X1 U7156 ( .A1(n5753), .A2(n4499), .ZN(n5767) );
  NAND2_X1 U7157 ( .A1(n5767), .A2(n5735), .ZN(n5739) );
  NAND2_X1 U7158 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n5736) );
  XNOR2_X1 U7159 ( .A(n5736), .B(P2_IR_REG_1__SCAN_IN), .ZN(n8535) );
  INV_X1 U7160 ( .A(n8535), .ZN(n5737) );
  NAND2_X1 U7161 ( .A1(n5823), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n5746) );
  NAND2_X1 U7162 ( .A1(n5788), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n5745) );
  INV_X1 U7163 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n5742) );
  NOR2_X1 U7164 ( .A1(n7781), .A2(n5742), .ZN(n5743) );
  NAND2_X1 U7165 ( .A1(n5707), .A2(n5743), .ZN(n5744) );
  NAND4_X2 U7166 ( .A1(n5747), .A2(n5746), .A3(n5745), .A4(n5744), .ZN(n6630)
         );
  XNOR2_X1 U7167 ( .A(n5748), .B(n5749), .ZN(n6581) );
  INV_X1 U7168 ( .A(n5748), .ZN(n5750) );
  NAND2_X1 U7169 ( .A1(n5750), .A2(n5749), .ZN(n5751) );
  NAND2_X1 U7170 ( .A1(n6579), .A2(n5751), .ZN(n5762) );
  NAND2_X1 U7171 ( .A1(n5767), .A2(n5752), .ZN(n5757) );
  NAND2_X1 U7172 ( .A1(n5819), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n5756) );
  NAND2_X1 U7173 ( .A1(n6253), .A2(n8548), .ZN(n5755) );
  AND3_X2 U7174 ( .A1(n5757), .A2(n5756), .A3(n5755), .ZN(n6739) );
  XNOR2_X1 U7175 ( .A(n6739), .B(n8035), .ZN(n5763) );
  NAND2_X1 U7176 ( .A1(n5828), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n5761) );
  NAND2_X1 U7177 ( .A1(n4276), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n5760) );
  NAND2_X1 U7178 ( .A1(n5923), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n5759) );
  NAND2_X1 U7179 ( .A1(n5823), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n5758) );
  NAND4_X1 U7180 ( .A1(n5761), .A2(n5760), .A3(n5759), .A4(n5758), .ZN(n6632)
         );
  NAND2_X1 U7181 ( .A1(n6632), .A2(n8165), .ZN(n5764) );
  XNOR2_X1 U7182 ( .A(n5763), .B(n5764), .ZN(n7970) );
  INV_X1 U7183 ( .A(n5763), .ZN(n5765) );
  NAND2_X1 U7184 ( .A1(n5765), .A2(n5764), .ZN(n5766) );
  NAND2_X1 U7185 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(n4300), .ZN(n5768) );
  XNOR2_X1 U7186 ( .A(n5768), .B(P2_IR_REG_3__SCAN_IN), .ZN(n9688) );
  NAND2_X1 U7187 ( .A1(n6253), .A2(n9688), .ZN(n5769) );
  XNOR2_X1 U7188 ( .A(n9792), .B(n8035), .ZN(n5775) );
  INV_X1 U7189 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n5770) );
  NAND2_X1 U7190 ( .A1(n5828), .A2(n5770), .ZN(n5774) );
  NAND2_X1 U7191 ( .A1(n5843), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n5773) );
  INV_X2 U7192 ( .A(n6169), .ZN(n5871) );
  NAND2_X1 U7193 ( .A1(n5871), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n5772) );
  NAND2_X1 U7194 ( .A1(n5823), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n5771) );
  AND2_X1 U7195 ( .A1(n8530), .A2(n8165), .ZN(n5776) );
  NAND2_X1 U7196 ( .A1(n5775), .A2(n5776), .ZN(n5794) );
  INV_X1 U7197 ( .A(n5775), .ZN(n6836) );
  INV_X1 U7198 ( .A(n5776), .ZN(n5777) );
  NAND2_X1 U7199 ( .A1(n6836), .A2(n5777), .ZN(n5778) );
  NAND2_X1 U7200 ( .A1(n5794), .A2(n5778), .ZN(n6207) );
  INV_X1 U7201 ( .A(n6207), .ZN(n5779) );
  NAND2_X1 U7202 ( .A1(n5767), .A2(n5780), .ZN(n5787) );
  NAND2_X1 U7203 ( .A1(n8147), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n5786) );
  NAND2_X1 U7204 ( .A1(n5782), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5783) );
  MUX2_X1 U7205 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5783), .S(
        P2_IR_REG_4__SCAN_IN), .Z(n5784) );
  AND2_X1 U7206 ( .A1(n5781), .A2(n5784), .ZN(n6541) );
  NAND2_X1 U7207 ( .A1(n6253), .A2(n6541), .ZN(n5785) );
  AND3_X2 U7208 ( .A1(n5787), .A2(n5786), .A3(n5785), .ZN(n7124) );
  XNOR2_X1 U7209 ( .A(n7124), .B(n8035), .ZN(n5796) );
  NAND2_X1 U7210 ( .A1(n5843), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n5793) );
  NAND2_X1 U7211 ( .A1(n8013), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n5792) );
  OAI21_X1 U7212 ( .B1(P2_REG3_REG_3__SCAN_IN), .B2(P2_REG3_REG_4__SCAN_IN), 
        .A(n5801), .ZN(n7120) );
  INV_X1 U7213 ( .A(n7120), .ZN(n5789) );
  NAND2_X1 U7214 ( .A1(n8034), .A2(n5789), .ZN(n5791) );
  NAND2_X1 U7215 ( .A1(n5871), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n5790) );
  NAND2_X1 U7216 ( .A1(n8529), .A2(n8165), .ZN(n5797) );
  XNOR2_X1 U7217 ( .A(n5796), .B(n5797), .ZN(n6837) );
  AND2_X1 U7218 ( .A1(n6837), .A2(n5794), .ZN(n5795) );
  INV_X1 U7219 ( .A(n5796), .ZN(n5798) );
  NAND2_X1 U7220 ( .A1(n5798), .A2(n5797), .ZN(n6845) );
  NAND2_X1 U7221 ( .A1(n5843), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n5806) );
  INV_X1 U7222 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n5800) );
  NAND2_X1 U7223 ( .A1(n5801), .A2(n5800), .ZN(n5802) );
  AND2_X1 U7224 ( .A1(n5826), .A2(n5802), .ZN(n7234) );
  NAND2_X1 U7225 ( .A1(n5828), .A2(n7234), .ZN(n5804) );
  NAND2_X1 U7226 ( .A1(n5923), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n5803) );
  AND2_X1 U7227 ( .A1(n8528), .A2(n8165), .ZN(n5815) );
  INV_X1 U7228 ( .A(n5815), .ZN(n5814) );
  NAND2_X1 U7229 ( .A1(n5819), .A2(P1_DATAO_REG_5__SCAN_IN), .ZN(n5813) );
  NAND2_X1 U7230 ( .A1(n5781), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5807) );
  MUX2_X1 U7231 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5807), .S(
        P2_IR_REG_5__SCAN_IN), .Z(n5811) );
  INV_X1 U7232 ( .A(n5809), .ZN(n5810) );
  NAND2_X1 U7233 ( .A1(n6253), .A2(n6524), .ZN(n5812) );
  OAI211_X2 U7234 ( .C1(n6225), .C2(n6097), .A(n5813), .B(n5812), .ZN(n7238)
         );
  XNOR2_X1 U7235 ( .A(n6132), .B(n7238), .ZN(n5816) );
  INV_X1 U7236 ( .A(n5816), .ZN(n6851) );
  NAND2_X1 U7237 ( .A1(n5814), .A2(n6851), .ZN(n6848) );
  AND2_X1 U7238 ( .A1(n6845), .A2(n6848), .ZN(n5818) );
  NAND2_X1 U7239 ( .A1(n5816), .A2(n5815), .ZN(n6844) );
  INV_X1 U7240 ( .A(n6844), .ZN(n5817) );
  AOI21_X1 U7241 ( .B1(n6846), .B2(n5818), .A(n5817), .ZN(n7956) );
  OR2_X1 U7242 ( .A1(n5809), .A2(n8873), .ZN(n5820) );
  XNOR2_X1 U7243 ( .A(n5820), .B(P2_IR_REG_6__SCAN_IN), .ZN(n9703) );
  AOI22_X1 U7244 ( .A1(n8147), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n6253), .B2(
        n9703), .ZN(n5822) );
  NAND2_X1 U7245 ( .A1(n6227), .A2(n5767), .ZN(n5821) );
  XNOR2_X1 U7246 ( .A(n7965), .B(n6132), .ZN(n5833) );
  NAND2_X1 U7247 ( .A1(n5823), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n5832) );
  NAND2_X1 U7248 ( .A1(n5843), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n5831) );
  INV_X1 U7249 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n5825) );
  NAND2_X1 U7250 ( .A1(n5826), .A2(n5825), .ZN(n5827) );
  AND2_X1 U7251 ( .A1(n5846), .A2(n5827), .ZN(n7962) );
  NAND2_X1 U7252 ( .A1(n5828), .A2(n7962), .ZN(n5830) );
  NAND2_X1 U7253 ( .A1(n5871), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n5829) );
  NAND4_X1 U7254 ( .A1(n5832), .A2(n5831), .A3(n5830), .A4(n5829), .ZN(n8527)
         );
  NAND2_X1 U7255 ( .A1(n8527), .A2(n8165), .ZN(n5834) );
  NAND2_X1 U7256 ( .A1(n5833), .A2(n5834), .ZN(n5838) );
  INV_X1 U7257 ( .A(n5833), .ZN(n5836) );
  INV_X1 U7258 ( .A(n5834), .ZN(n5835) );
  NAND2_X1 U7259 ( .A1(n5836), .A2(n5835), .ZN(n5837) );
  AND2_X1 U7260 ( .A1(n5838), .A2(n5837), .ZN(n7957) );
  NAND2_X1 U7261 ( .A1(n6231), .A2(n6129), .ZN(n5842) );
  NAND2_X1 U7262 ( .A1(n5809), .A2(n5839), .ZN(n5859) );
  NAND2_X1 U7263 ( .A1(n5859), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5840) );
  XNOR2_X1 U7264 ( .A(n5840), .B(P2_IR_REG_7__SCAN_IN), .ZN(n9715) );
  AOI22_X1 U7265 ( .A1(n8147), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n6253), .B2(
        n9715), .ZN(n5841) );
  XNOR2_X1 U7266 ( .A(n8219), .B(n8035), .ZN(n5853) );
  NAND2_X1 U7267 ( .A1(n8013), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n5851) );
  NAND2_X1 U7268 ( .A1(n5843), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n5850) );
  INV_X1 U7269 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n5845) );
  NAND2_X1 U7270 ( .A1(n5846), .A2(n5845), .ZN(n5847) );
  AND2_X1 U7271 ( .A1(n5869), .A2(n5847), .ZN(n7289) );
  NAND2_X1 U7272 ( .A1(n8034), .A2(n7289), .ZN(n5849) );
  NAND2_X1 U7273 ( .A1(n5923), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n5848) );
  NAND4_X1 U7274 ( .A1(n5851), .A2(n5850), .A3(n5849), .A4(n5848), .ZN(n8526)
         );
  NAND2_X1 U7275 ( .A1(n8526), .A2(n8165), .ZN(n5854) );
  XNOR2_X1 U7276 ( .A(n5853), .B(n5854), .ZN(n6682) );
  INV_X1 U7277 ( .A(n6682), .ZN(n5852) );
  INV_X1 U7278 ( .A(n5853), .ZN(n5856) );
  INV_X1 U7279 ( .A(n5854), .ZN(n5855) );
  NAND2_X1 U7280 ( .A1(n5856), .A2(n5855), .ZN(n5857) );
  NAND2_X1 U7281 ( .A1(n6243), .A2(n6129), .ZN(n5866) );
  INV_X1 U7282 ( .A(n5900), .ZN(n5864) );
  NAND2_X1 U7283 ( .A1(n5860), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5862) );
  MUX2_X1 U7284 ( .A(n5862), .B(P2_IR_REG_31__SCAN_IN), .S(n5861), .Z(n5863)
         );
  AOI22_X1 U7285 ( .A1(n8147), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n6253), .B2(
        n6563), .ZN(n5865) );
  XNOR2_X1 U7286 ( .A(n7062), .B(n8035), .ZN(n5877) );
  NAND2_X1 U7287 ( .A1(n8013), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n5875) );
  NAND2_X1 U7288 ( .A1(n5843), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n5874) );
  INV_X1 U7289 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n5868) );
  NAND2_X1 U7290 ( .A1(n5869), .A2(n5868), .ZN(n5870) );
  AND2_X1 U7291 ( .A1(n5886), .A2(n5870), .ZN(n7241) );
  NAND2_X1 U7292 ( .A1(n8034), .A2(n7241), .ZN(n5873) );
  NAND2_X1 U7293 ( .A1(n5871), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n5872) );
  INV_X1 U7294 ( .A(n8165), .ZN(n5876) );
  NOR2_X1 U7295 ( .A1(n7296), .A2(n5876), .ZN(n5878) );
  XNOR2_X1 U7296 ( .A(n5877), .B(n5878), .ZN(n6824) );
  INV_X1 U7297 ( .A(n5877), .ZN(n5879) );
  NAND2_X1 U7298 ( .A1(n5879), .A2(n5878), .ZN(n5880) );
  NAND2_X1 U7299 ( .A1(n6245), .A2(n6129), .ZN(n5883) );
  OR2_X1 U7300 ( .A1(n5900), .A2(n8873), .ZN(n5881) );
  XNOR2_X1 U7301 ( .A(n5881), .B(P2_IR_REG_9__SCAN_IN), .ZN(n6564) );
  AOI22_X1 U7302 ( .A1(n8147), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n6253), .B2(
        n6564), .ZN(n5882) );
  NAND2_X1 U7303 ( .A1(n5883), .A2(n5882), .ZN(n7366) );
  XNOR2_X1 U7304 ( .A(n7366), .B(n8035), .ZN(n5892) );
  NAND2_X1 U7305 ( .A1(n5843), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n5891) );
  NAND2_X1 U7306 ( .A1(n8013), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n5890) );
  INV_X1 U7307 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n5885) );
  NAND2_X1 U7308 ( .A1(n5886), .A2(n5885), .ZN(n5887) );
  AND2_X1 U7309 ( .A1(n5904), .A2(n5887), .ZN(n7365) );
  NAND2_X1 U7310 ( .A1(n8034), .A2(n7365), .ZN(n5889) );
  NAND2_X1 U7311 ( .A1(n5871), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n5888) );
  OR2_X1 U7312 ( .A1(n7078), .A2(n5876), .ZN(n5893) );
  NAND2_X1 U7313 ( .A1(n5892), .A2(n5893), .ZN(n5898) );
  INV_X1 U7314 ( .A(n5892), .ZN(n5895) );
  INV_X1 U7315 ( .A(n5893), .ZN(n5894) );
  NAND2_X1 U7316 ( .A1(n5895), .A2(n5894), .ZN(n5896) );
  NAND2_X1 U7317 ( .A1(n5898), .A2(n5896), .ZN(n6995) );
  INV_X1 U7318 ( .A(n6995), .ZN(n5897) );
  NAND2_X1 U7319 ( .A1(n6248), .A2(n6129), .ZN(n5902) );
  INV_X1 U7320 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n5899) );
  NAND2_X1 U7321 ( .A1(n5900), .A2(n5899), .ZN(n5933) );
  NAND2_X1 U7322 ( .A1(n5933), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5915) );
  XNOR2_X1 U7323 ( .A(n5915), .B(P2_IR_REG_10__SCAN_IN), .ZN(n9728) );
  AOI22_X1 U7324 ( .A1(n8147), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n6253), .B2(
        n9728), .ZN(n5901) );
  NAND2_X1 U7325 ( .A1(n5902), .A2(n5901), .ZN(n7322) );
  XNOR2_X1 U7326 ( .A(n7322), .B(n6132), .ZN(n5910) );
  NAND2_X1 U7327 ( .A1(n8013), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n5909) );
  NAND2_X1 U7328 ( .A1(n5843), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n5908) );
  INV_X1 U7329 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n5903) );
  NAND2_X1 U7330 ( .A1(n5904), .A2(n5903), .ZN(n5905) );
  AND2_X1 U7331 ( .A1(n5921), .A2(n5905), .ZN(n7132) );
  NAND2_X1 U7332 ( .A1(n8034), .A2(n7132), .ZN(n5907) );
  NAND2_X1 U7333 ( .A1(n5871), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n5906) );
  NOR2_X1 U7334 ( .A1(n7376), .A2(n5876), .ZN(n5911) );
  XNOR2_X1 U7335 ( .A(n5910), .B(n5911), .ZN(n7007) );
  INV_X1 U7336 ( .A(n5910), .ZN(n5913) );
  INV_X1 U7337 ( .A(n5911), .ZN(n5912) );
  NAND2_X1 U7338 ( .A1(n6262), .A2(n6129), .ZN(n5919) );
  NAND2_X1 U7339 ( .A1(n5915), .A2(n5914), .ZN(n5916) );
  NAND2_X1 U7340 ( .A1(n5916), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5917) );
  XNOR2_X1 U7341 ( .A(n5917), .B(P2_IR_REG_11__SCAN_IN), .ZN(n6562) );
  AOI22_X1 U7342 ( .A1(n8147), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n6253), .B2(
        n6562), .ZN(n5918) );
  XNOR2_X1 U7343 ( .A(n9818), .B(n8035), .ZN(n5928) );
  NAND2_X1 U7344 ( .A1(n8013), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n5927) );
  NAND2_X1 U7345 ( .A1(n5843), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n5926) );
  INV_X1 U7346 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n7273) );
  NAND2_X1 U7347 ( .A1(n5921), .A2(n7273), .ZN(n5922) );
  AND2_X1 U7348 ( .A1(n5938), .A2(n5922), .ZN(n7379) );
  NAND2_X1 U7349 ( .A1(n8034), .A2(n7379), .ZN(n5925) );
  NAND2_X1 U7350 ( .A1(n5923), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n5924) );
  NOR2_X1 U7351 ( .A1(n7442), .A2(n5876), .ZN(n5929) );
  XNOR2_X1 U7352 ( .A(n5928), .B(n5929), .ZN(n7272) );
  NAND2_X1 U7353 ( .A1(n7271), .A2(n7272), .ZN(n5932) );
  INV_X1 U7354 ( .A(n5928), .ZN(n5930) );
  NAND2_X1 U7355 ( .A1(n5930), .A2(n5929), .ZN(n5931) );
  NAND2_X1 U7356 ( .A1(n5948), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5934) );
  XNOR2_X1 U7357 ( .A(n5934), .B(P2_IR_REG_12__SCAN_IN), .ZN(n6586) );
  AOI22_X1 U7358 ( .A1(n8147), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n6253), .B2(
        n6586), .ZN(n5935) );
  XNOR2_X1 U7359 ( .A(n8848), .B(n8035), .ZN(n5944) );
  NAND2_X1 U7360 ( .A1(n8013), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n5943) );
  NAND2_X1 U7361 ( .A1(n4276), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n5942) );
  INV_X1 U7362 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n5937) );
  NAND2_X1 U7363 ( .A1(n5938), .A2(n5937), .ZN(n5939) );
  AND2_X1 U7364 ( .A1(n5952), .A2(n5939), .ZN(n7436) );
  NAND2_X1 U7365 ( .A1(n8034), .A2(n7436), .ZN(n5941) );
  NAND2_X1 U7366 ( .A1(n5871), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n5940) );
  OR2_X1 U7367 ( .A1(n7453), .A2(n5876), .ZN(n5945) );
  NAND2_X1 U7368 ( .A1(n5944), .A2(n5945), .ZN(n7304) );
  INV_X1 U7369 ( .A(n5944), .ZN(n5947) );
  INV_X1 U7370 ( .A(n5945), .ZN(n5946) );
  NAND2_X1 U7371 ( .A1(n5947), .A2(n5946), .ZN(n7305) );
  NAND2_X1 U7372 ( .A1(n6333), .A2(n6129), .ZN(n5950) );
  OAI21_X1 U7373 ( .B1(n5948), .B2(P2_IR_REG_12__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5963) );
  XNOR2_X1 U7374 ( .A(n5963), .B(P2_IR_REG_13__SCAN_IN), .ZN(n6575) );
  AOI22_X1 U7375 ( .A1(n8147), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n6253), .B2(
        n6575), .ZN(n5949) );
  XNOR2_X1 U7376 ( .A(n7599), .B(n6132), .ZN(n8043) );
  INV_X1 U7377 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n6570) );
  NAND2_X1 U7378 ( .A1(n5952), .A2(n6570), .ZN(n5953) );
  AND2_X1 U7379 ( .A1(n5968), .A2(n5953), .ZN(n7455) );
  NAND2_X1 U7380 ( .A1(n8034), .A2(n7455), .ZN(n5957) );
  NAND2_X1 U7381 ( .A1(n5843), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n5956) );
  NAND2_X1 U7382 ( .A1(n5871), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n5955) );
  NAND2_X1 U7383 ( .A1(n8013), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n5954) );
  NOR2_X1 U7384 ( .A1(n7679), .A2(n5876), .ZN(n5958) );
  NAND2_X1 U7385 ( .A1(n8043), .A2(n5958), .ZN(n5974) );
  INV_X1 U7386 ( .A(n8043), .ZN(n5960) );
  INV_X1 U7387 ( .A(n5958), .ZN(n5959) );
  NAND2_X1 U7388 ( .A1(n5960), .A2(n5959), .ZN(n5961) );
  AND2_X1 U7389 ( .A1(n5974), .A2(n5961), .ZN(n7451) );
  INV_X2 U7390 ( .A(n6097), .ZN(n6129) );
  NAND2_X1 U7391 ( .A1(n6337), .A2(n6129), .ZN(n5966) );
  INV_X1 U7392 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n5962) );
  NAND2_X1 U7393 ( .A1(n5963), .A2(n5962), .ZN(n5964) );
  NAND2_X1 U7394 ( .A1(n5964), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5981) );
  XNOR2_X1 U7395 ( .A(n5981), .B(P2_IR_REG_14__SCAN_IN), .ZN(n7149) );
  AOI22_X1 U7396 ( .A1(n7149), .A2(n6253), .B1(n5819), .B2(
        P1_DATAO_REG_14__SCAN_IN), .ZN(n5965) );
  XNOR2_X1 U7397 ( .A(n8843), .B(n6132), .ZN(n5976) );
  NAND2_X1 U7398 ( .A1(n8013), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n5973) );
  NAND2_X1 U7399 ( .A1(n4276), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n5972) );
  INV_X1 U7400 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n5967) );
  NAND2_X1 U7401 ( .A1(n5968), .A2(n5967), .ZN(n5969) );
  AND2_X1 U7402 ( .A1(n5986), .A2(n5969), .ZN(n8053) );
  NAND2_X1 U7403 ( .A1(n8034), .A2(n8053), .ZN(n5971) );
  NAND2_X1 U7404 ( .A1(n5871), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n5970) );
  NAND4_X1 U7405 ( .A1(n5973), .A2(n5972), .A3(n5971), .A4(n5970), .ZN(n8519)
         );
  NAND2_X1 U7406 ( .A1(n8519), .A2(n8165), .ZN(n5977) );
  XNOR2_X1 U7407 ( .A(n5976), .B(n5977), .ZN(n8045) );
  AND2_X1 U7408 ( .A1(n8045), .A2(n5974), .ZN(n5975) );
  NAND2_X1 U7409 ( .A1(n7449), .A2(n5975), .ZN(n8056) );
  INV_X1 U7410 ( .A(n5976), .ZN(n5978) );
  NAND2_X1 U7411 ( .A1(n5978), .A2(n5977), .ZN(n5979) );
  NAND2_X1 U7412 ( .A1(n8056), .A2(n5979), .ZN(n5992) );
  NAND2_X1 U7413 ( .A1(n6442), .A2(n6129), .ZN(n5985) );
  NAND2_X1 U7414 ( .A1(n5981), .A2(n5980), .ZN(n5982) );
  NAND2_X1 U7415 ( .A1(n5982), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5983) );
  XNOR2_X1 U7416 ( .A(n5983), .B(P2_IR_REG_15__SCAN_IN), .ZN(n8564) );
  AOI22_X1 U7417 ( .A1(n8564), .A2(n6253), .B1(n5819), .B2(
        P1_DATAO_REG_15__SCAN_IN), .ZN(n5984) );
  XNOR2_X1 U7418 ( .A(n7647), .B(n8035), .ZN(n5993) );
  NAND2_X1 U7419 ( .A1(n5843), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n5991) );
  NAND2_X1 U7420 ( .A1(n5871), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n5990) );
  INV_X1 U7421 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n9998) );
  NAND2_X1 U7422 ( .A1(n5986), .A2(n9998), .ZN(n5987) );
  AND2_X1 U7423 ( .A1(n6002), .A2(n5987), .ZN(n7778) );
  NAND2_X1 U7424 ( .A1(n8034), .A2(n7778), .ZN(n5989) );
  NAND2_X1 U7425 ( .A1(n8013), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n5988) );
  NOR2_X1 U7426 ( .A1(n8050), .A2(n5876), .ZN(n7769) );
  INV_X1 U7427 ( .A(n5993), .ZN(n5994) );
  INV_X1 U7428 ( .A(n7784), .ZN(n6009) );
  NAND2_X1 U7429 ( .A1(n6446), .A2(n6129), .ZN(n5999) );
  NOR2_X1 U7430 ( .A1(n5722), .A2(n8873), .ZN(n5996) );
  MUX2_X1 U7431 ( .A(n8873), .B(n5996), .S(P2_IR_REG_16__SCAN_IN), .Z(n5997)
         );
  OR2_X1 U7432 ( .A1(n5997), .A2(n6015), .ZN(n7620) );
  INV_X1 U7433 ( .A(n7620), .ZN(n7156) );
  AOI22_X1 U7434 ( .A1(n8147), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n6253), .B2(
        n7156), .ZN(n5998) );
  XNOR2_X1 U7435 ( .A(n7791), .B(n6132), .ZN(n6010) );
  INV_X1 U7436 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n6001) );
  NAND2_X1 U7437 ( .A1(n6002), .A2(n6001), .ZN(n6003) );
  AND2_X1 U7438 ( .A1(n6025), .A2(n6003), .ZN(n7662) );
  NAND2_X1 U7439 ( .A1(n7662), .A2(n8034), .ZN(n6007) );
  NAND2_X1 U7440 ( .A1(n5843), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n6006) );
  NAND2_X1 U7441 ( .A1(n8013), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n6005) );
  NAND2_X1 U7442 ( .A1(n5871), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n6004) );
  NOR2_X1 U7443 ( .A1(n7745), .A2(n5876), .ZN(n6011) );
  XNOR2_X1 U7444 ( .A(n6010), .B(n6011), .ZN(n7785) );
  INV_X1 U7445 ( .A(n6010), .ZN(n6013) );
  INV_X1 U7446 ( .A(n6011), .ZN(n6012) );
  NAND2_X1 U7447 ( .A1(n6013), .A2(n6012), .ZN(n6014) );
  NAND2_X1 U7448 ( .A1(n6620), .A2(n6129), .ZN(n6020) );
  NAND2_X1 U7449 ( .A1(n6016), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6018) );
  XNOR2_X1 U7450 ( .A(n6018), .B(n6017), .ZN(n7622) );
  INV_X1 U7451 ( .A(n7622), .ZN(n9746) );
  AOI22_X1 U7452 ( .A1(n8147), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n6253), .B2(
        n9746), .ZN(n6019) );
  XNOR2_X1 U7453 ( .A(n8834), .B(n6132), .ZN(n6030) );
  NAND2_X1 U7454 ( .A1(n8013), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n6022) );
  NAND2_X1 U7455 ( .A1(n4276), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n6021) );
  AND2_X1 U7456 ( .A1(n6022), .A2(n6021), .ZN(n6029) );
  INV_X1 U7457 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n6024) );
  NAND2_X1 U7458 ( .A1(n6025), .A2(n6024), .ZN(n6026) );
  NAND2_X1 U7459 ( .A1(n6039), .A2(n6026), .ZN(n7815) );
  OR2_X1 U7460 ( .A1(n7815), .A2(n8001), .ZN(n6028) );
  NAND2_X1 U7461 ( .A1(n5871), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n6027) );
  NOR2_X1 U7462 ( .A1(n8494), .A2(n5876), .ZN(n6031) );
  NAND2_X1 U7463 ( .A1(n6030), .A2(n6031), .ZN(n6034) );
  INV_X1 U7464 ( .A(n6030), .ZN(n8485) );
  INV_X1 U7465 ( .A(n6031), .ZN(n6032) );
  NAND2_X1 U7466 ( .A1(n8485), .A2(n6032), .ZN(n6033) );
  NAND2_X1 U7467 ( .A1(n6034), .A2(n6033), .ZN(n7811) );
  NAND2_X1 U7468 ( .A1(n6776), .A2(n6129), .ZN(n6038) );
  NAND2_X1 U7469 ( .A1(n6035), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6036) );
  XNOR2_X1 U7470 ( .A(n6036), .B(P2_IR_REG_18__SCAN_IN), .ZN(n7629) );
  AOI22_X1 U7471 ( .A1(n5819), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n6253), .B2(
        n7629), .ZN(n6037) );
  XNOR2_X1 U7472 ( .A(n8827), .B(n6132), .ZN(n6043) );
  INV_X1 U7473 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n7626) );
  NAND2_X1 U7474 ( .A1(n6039), .A2(n7626), .ZN(n6040) );
  NAND2_X1 U7475 ( .A1(n6052), .A2(n6040), .ZN(n8489) );
  AOI22_X1 U7476 ( .A1(n8013), .A2(P2_REG0_REG_18__SCAN_IN), .B1(n5843), .B2(
        P2_REG2_REG_18__SCAN_IN), .ZN(n6042) );
  NAND2_X1 U7477 ( .A1(n5871), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n6041) );
  OAI211_X1 U7478 ( .C1(n8489), .C2(n8001), .A(n6042), .B(n6041), .ZN(n8517)
         );
  AND2_X1 U7479 ( .A1(n8517), .A2(n8165), .ZN(n6044) );
  NAND2_X1 U7480 ( .A1(n6043), .A2(n6044), .ZN(n6057) );
  INV_X1 U7481 ( .A(n6043), .ZN(n8431) );
  INV_X1 U7482 ( .A(n6044), .ZN(n6045) );
  NAND2_X1 U7483 ( .A1(n8431), .A2(n6045), .ZN(n6046) );
  NAND2_X1 U7484 ( .A1(n6047), .A2(n8482), .ZN(n8486) );
  NAND2_X1 U7485 ( .A1(n6890), .A2(n6129), .ZN(n6049) );
  AOI22_X1 U7486 ( .A1(n5819), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n6253), .B2(
        n4282), .ZN(n6048) );
  XNOR2_X1 U7487 ( .A(n8390), .B(n8035), .ZN(n6059) );
  INV_X1 U7488 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n6051) );
  NAND2_X1 U7489 ( .A1(n6052), .A2(n6051), .ZN(n6053) );
  NAND2_X1 U7490 ( .A1(n6066), .A2(n6053), .ZN(n8732) );
  OR2_X1 U7491 ( .A1(n8732), .A2(n8001), .ZN(n6056) );
  AOI22_X1 U7492 ( .A1(n8013), .A2(P2_REG0_REG_19__SCAN_IN), .B1(n4276), .B2(
        P2_REG2_REG_19__SCAN_IN), .ZN(n6055) );
  NAND2_X1 U7493 ( .A1(n5871), .A2(P2_REG1_REG_19__SCAN_IN), .ZN(n6054) );
  INV_X1 U7494 ( .A(n8701), .ZN(n8756) );
  NAND2_X1 U7495 ( .A1(n8756), .A2(n8165), .ZN(n6060) );
  XNOR2_X1 U7496 ( .A(n6059), .B(n6060), .ZN(n8432) );
  INV_X1 U7497 ( .A(n6059), .ZN(n6061) );
  NAND2_X1 U7498 ( .A1(n6061), .A2(n6060), .ZN(n6062) );
  NAND2_X1 U7499 ( .A1(n6972), .A2(n6129), .ZN(n6064) );
  NAND2_X1 U7500 ( .A1(n8147), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n6063) );
  NAND2_X2 U7501 ( .A1(n6064), .A2(n6063), .ZN(n8705) );
  XNOR2_X1 U7502 ( .A(n8705), .B(n6132), .ZN(n6074) );
  INV_X1 U7503 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n6065) );
  NAND2_X1 U7504 ( .A1(n6066), .A2(n6065), .ZN(n6067) );
  AND2_X1 U7505 ( .A1(n6084), .A2(n6067), .ZN(n8704) );
  NAND2_X1 U7506 ( .A1(n8704), .A2(n8034), .ZN(n6073) );
  INV_X1 U7507 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n6070) );
  NAND2_X1 U7508 ( .A1(n4276), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n6069) );
  NAND2_X1 U7509 ( .A1(n5871), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n6068) );
  OAI211_X1 U7510 ( .C1(n6070), .C2(n8154), .A(n6069), .B(n6068), .ZN(n6071)
         );
  INV_X1 U7511 ( .A(n6071), .ZN(n6072) );
  NOR2_X1 U7512 ( .A1(n8722), .A2(n5876), .ZN(n6075) );
  NAND2_X1 U7513 ( .A1(n6074), .A2(n6075), .ZN(n6079) );
  INV_X1 U7514 ( .A(n6074), .ZN(n8440) );
  INV_X1 U7515 ( .A(n6075), .ZN(n6076) );
  NAND2_X1 U7516 ( .A1(n8440), .A2(n6076), .ZN(n6077) );
  NAND2_X1 U7517 ( .A1(n6079), .A2(n6077), .ZN(n8465) );
  INV_X1 U7518 ( .A(n8465), .ZN(n6078) );
  NAND2_X1 U7519 ( .A1(n8437), .A2(n6079), .ZN(n6092) );
  NAND2_X1 U7520 ( .A1(n6974), .A2(n6129), .ZN(n6081) );
  NAND2_X1 U7521 ( .A1(n8147), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n6080) );
  XNOR2_X1 U7522 ( .A(n8692), .B(n8035), .ZN(n6095) );
  INV_X1 U7523 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n6083) );
  NAND2_X1 U7524 ( .A1(n6084), .A2(n6083), .ZN(n6085) );
  NAND2_X1 U7525 ( .A1(n6101), .A2(n6085), .ZN(n8444) );
  OR2_X1 U7526 ( .A1(n8444), .A2(n8001), .ZN(n6091) );
  INV_X1 U7527 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n6088) );
  NAND2_X1 U7528 ( .A1(n5871), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n6087) );
  NAND2_X1 U7529 ( .A1(n5843), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n6086) );
  OAI211_X1 U7530 ( .C1(n8154), .C2(n6088), .A(n6087), .B(n6086), .ZN(n6089)
         );
  INV_X1 U7531 ( .A(n6089), .ZN(n6090) );
  NAND2_X1 U7532 ( .A1(n8515), .A2(n8165), .ZN(n6093) );
  XNOR2_X1 U7533 ( .A(n6095), .B(n6093), .ZN(n8438) );
  NAND2_X1 U7534 ( .A1(n6092), .A2(n8438), .ZN(n8441) );
  INV_X1 U7535 ( .A(n6093), .ZN(n6094) );
  NAND2_X1 U7536 ( .A1(n6095), .A2(n6094), .ZN(n6096) );
  NAND2_X1 U7537 ( .A1(n7003), .A2(n6129), .ZN(n6099) );
  NAND2_X1 U7538 ( .A1(n8147), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n6098) );
  XNOR2_X1 U7539 ( .A(n8806), .B(n8035), .ZN(n6110) );
  INV_X1 U7541 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n6100) );
  NAND2_X1 U7542 ( .A1(n6101), .A2(n6100), .ZN(n6102) );
  AND2_X1 U7543 ( .A1(n6118), .A2(n6102), .ZN(n8677) );
  NAND2_X1 U7544 ( .A1(n8677), .A2(n8034), .ZN(n6109) );
  INV_X1 U7545 ( .A(n5788), .ZN(n6106) );
  INV_X1 U7546 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n6105) );
  NAND2_X1 U7547 ( .A1(n8013), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n6104) );
  NAND2_X1 U7548 ( .A1(n5871), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n6103) );
  OAI211_X1 U7549 ( .C1(n6106), .C2(n6105), .A(n6104), .B(n6103), .ZN(n6107)
         );
  INV_X1 U7550 ( .A(n6107), .ZN(n6108) );
  OR2_X1 U7551 ( .A1(n8686), .A2(n5876), .ZN(n8474) );
  INV_X1 U7552 ( .A(n6110), .ZN(n6111) );
  NAND2_X1 U7554 ( .A1(n7060), .A2(n6129), .ZN(n6115) );
  NAND2_X1 U7555 ( .A1(n8147), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n6114) );
  XNOR2_X1 U7556 ( .A(n8799), .B(n8035), .ZN(n6126) );
  XNOR2_X1 U7557 ( .A(n6128), .B(n6126), .ZN(n7983) );
  INV_X1 U7558 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n6117) );
  NAND2_X1 U7559 ( .A1(n6118), .A2(n6117), .ZN(n6119) );
  NAND2_X1 U7560 ( .A1(n6186), .A2(n6119), .ZN(n8656) );
  OR2_X1 U7561 ( .A1(n8656), .A2(n8001), .ZN(n6125) );
  INV_X1 U7562 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n6122) );
  NAND2_X1 U7563 ( .A1(n4276), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n6121) );
  NAND2_X1 U7564 ( .A1(n5871), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n6120) );
  OAI211_X1 U7565 ( .C1(n6122), .C2(n8154), .A(n6121), .B(n6120), .ZN(n6123)
         );
  INV_X1 U7566 ( .A(n6123), .ZN(n6124) );
  NOR2_X1 U7567 ( .A1(n8674), .A2(n5876), .ZN(n7981) );
  INV_X1 U7568 ( .A(n6126), .ZN(n6127) );
  NOR2_X1 U7569 ( .A1(n8424), .A2(n7984), .ZN(n6133) );
  NAND2_X1 U7570 ( .A1(n7163), .A2(n6129), .ZN(n6131) );
  NAND2_X1 U7571 ( .A1(n5819), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n6130) );
  XNOR2_X1 U7572 ( .A(n8796), .B(n6132), .ZN(n7986) );
  INV_X1 U7573 ( .A(n7986), .ZN(n7988) );
  XNOR2_X1 U7574 ( .A(n6133), .B(n7988), .ZN(n6174) );
  NAND2_X1 U7575 ( .A1(n6135), .A2(n6134), .ZN(n6136) );
  NAND2_X1 U7576 ( .A1(n6136), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6160) );
  NAND2_X1 U7577 ( .A1(n6160), .A2(n6159), .ZN(n6162) );
  NAND2_X1 U7578 ( .A1(n6162), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6138) );
  NAND2_X1 U7579 ( .A1(n4331), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6139) );
  XNOR2_X1 U7580 ( .A(n6139), .B(P2_IR_REG_26__SCAN_IN), .ZN(n9778) );
  INV_X1 U7581 ( .A(n9778), .ZN(n7524) );
  AND2_X1 U7582 ( .A1(n7199), .A2(n7524), .ZN(n9777) );
  INV_X1 U7583 ( .A(n7199), .ZN(n6142) );
  INV_X1 U7584 ( .A(P2_B_REG_SCAN_IN), .ZN(n9966) );
  NAND2_X1 U7585 ( .A1(n6140), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6141) );
  XNOR2_X1 U7586 ( .A(n6141), .B(P2_IR_REG_25__SCAN_IN), .ZN(n9779) );
  AOI221_X1 U7587 ( .B1(n6142), .B2(P2_B_REG_SCAN_IN), .C1(n7199), .C2(n9966), 
        .A(n9779), .ZN(n6143) );
  INV_X1 U7588 ( .A(n6143), .ZN(n6144) );
  NOR2_X1 U7589 ( .A1(n9773), .A2(P2_D_REG_0__SCAN_IN), .ZN(n6145) );
  NOR4_X1 U7590 ( .A1(P2_D_REG_2__SCAN_IN), .A2(P2_D_REG_4__SCAN_IN), .A3(
        P2_D_REG_5__SCAN_IN), .A4(P2_D_REG_6__SCAN_IN), .ZN(n6154) );
  NOR4_X1 U7591 ( .A1(P2_D_REG_9__SCAN_IN), .A2(P2_D_REG_11__SCAN_IN), .A3(
        P2_D_REG_12__SCAN_IN), .A4(P2_D_REG_13__SCAN_IN), .ZN(n6153) );
  INV_X1 U7592 ( .A(P2_D_REG_8__SCAN_IN), .ZN(n9905) );
  INV_X1 U7593 ( .A(P2_D_REG_3__SCAN_IN), .ZN(n9920) );
  INV_X1 U7594 ( .A(P2_D_REG_7__SCAN_IN), .ZN(n9958) );
  INV_X1 U7595 ( .A(P2_D_REG_10__SCAN_IN), .ZN(n10006) );
  NAND4_X1 U7596 ( .A1(n9905), .A2(n9920), .A3(n9958), .A4(n10006), .ZN(n6151)
         );
  NOR4_X1 U7597 ( .A1(P2_D_REG_18__SCAN_IN), .A2(P2_D_REG_19__SCAN_IN), .A3(
        P2_D_REG_20__SCAN_IN), .A4(P2_D_REG_21__SCAN_IN), .ZN(n6149) );
  NOR4_X1 U7598 ( .A1(P2_D_REG_16__SCAN_IN), .A2(P2_D_REG_14__SCAN_IN), .A3(
        P2_D_REG_15__SCAN_IN), .A4(P2_D_REG_17__SCAN_IN), .ZN(n6148) );
  NOR4_X1 U7599 ( .A1(P2_D_REG_26__SCAN_IN), .A2(P2_D_REG_27__SCAN_IN), .A3(
        P2_D_REG_28__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n6147) );
  NOR4_X1 U7600 ( .A1(P2_D_REG_22__SCAN_IN), .A2(P2_D_REG_23__SCAN_IN), .A3(
        P2_D_REG_24__SCAN_IN), .A4(P2_D_REG_25__SCAN_IN), .ZN(n6146) );
  NAND4_X1 U7601 ( .A1(n6149), .A2(n6148), .A3(n6147), .A4(n6146), .ZN(n6150)
         );
  NOR4_X1 U7602 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        n6151), .A4(n6150), .ZN(n6152) );
  AND3_X1 U7603 ( .A1(n6154), .A2(n6153), .A3(n6152), .ZN(n6155) );
  NOR2_X1 U7604 ( .A1(n6155), .A2(n9773), .ZN(n6624) );
  OR2_X1 U7605 ( .A1(n9773), .A2(P2_D_REG_1__SCAN_IN), .ZN(n6157) );
  OR2_X1 U7606 ( .A1(n9778), .A2(n9779), .ZN(n6156) );
  NAND2_X1 U7607 ( .A1(n6157), .A2(n6156), .ZN(n6622) );
  NOR2_X1 U7608 ( .A1(n6624), .A2(n6622), .ZN(n7108) );
  INV_X1 U7609 ( .A(n7108), .ZN(n6158) );
  INV_X1 U7610 ( .A(n6182), .ZN(n6166) );
  INV_X1 U7611 ( .A(n9779), .ZN(n7458) );
  OR2_X1 U7612 ( .A1(n6160), .A2(n6159), .ZN(n6161) );
  NAND2_X1 U7613 ( .A1(n6162), .A2(n6161), .ZN(n6252) );
  INV_X1 U7614 ( .A(n7117), .ZN(n6646) );
  INV_X1 U7615 ( .A(n8373), .ZN(n7116) );
  AND2_X1 U7616 ( .A1(n7116), .A2(n5730), .ZN(n8380) );
  INV_X1 U7617 ( .A(n8380), .ZN(n6163) );
  NAND2_X1 U7618 ( .A1(n8383), .A2(n5733), .ZN(n6628) );
  INV_X1 U7619 ( .A(n6628), .ZN(n6255) );
  NOR2_X1 U7620 ( .A1(n8849), .A2(n6255), .ZN(n6164) );
  AND2_X1 U7621 ( .A1(n9774), .A2(n6164), .ZN(n6165) );
  XNOR2_X1 U7622 ( .A(n6186), .B(P2_REG3_REG_24__SCAN_IN), .ZN(n8647) );
  NAND2_X1 U7623 ( .A1(n8647), .A2(n8034), .ZN(n6173) );
  INV_X1 U7624 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n6170) );
  NAND2_X1 U7625 ( .A1(n4276), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n6168) );
  NAND2_X1 U7626 ( .A1(n8013), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n6167) );
  OAI211_X1 U7627 ( .C1(n6170), .C2(n6169), .A(n6168), .B(n6167), .ZN(n6171)
         );
  INV_X1 U7628 ( .A(n6171), .ZN(n6172) );
  NAND2_X1 U7629 ( .A1(n6173), .A2(n6172), .ZN(n8663) );
  INV_X1 U7630 ( .A(n8663), .ZN(n8458) );
  OR2_X1 U7631 ( .A1(n8511), .A2(n5876), .ZN(n8484) );
  OAI22_X1 U7632 ( .A1(n6174), .A2(n8511), .B1(n8458), .B2(n8484), .ZN(n6177)
         );
  INV_X1 U7633 ( .A(n6174), .ZN(n6175) );
  AND2_X1 U7634 ( .A1(n8663), .A2(n8165), .ZN(n7985) );
  INV_X1 U7635 ( .A(n7985), .ZN(n7987) );
  NAND2_X1 U7636 ( .A1(n6175), .A2(n7985), .ZN(n6176) );
  NAND2_X1 U7637 ( .A1(n6177), .A2(n6176), .ZN(n6199) );
  NAND2_X1 U7638 ( .A1(n7951), .A2(n4282), .ZN(n8179) );
  OR2_X1 U7639 ( .A1(n8179), .A2(n8373), .ZN(n9381) );
  OR2_X1 U7640 ( .A1(n9381), .A2(n5733), .ZN(n7112) );
  NAND2_X1 U7641 ( .A1(n6182), .A2(n7112), .ZN(n6180) );
  AND2_X1 U7642 ( .A1(n9774), .A2(n8849), .ZN(n6178) );
  OR2_X1 U7643 ( .A1(n8380), .A2(n6628), .ZN(n7109) );
  AND3_X1 U7644 ( .A1(n6473), .A2(n6252), .A3(n7109), .ZN(n6179) );
  NAND2_X1 U7645 ( .A1(n6180), .A2(n6179), .ZN(n6735) );
  NAND2_X1 U7646 ( .A1(n9774), .A2(n8380), .ZN(n6181) );
  NOR2_X1 U7647 ( .A1(n6182), .A2(n6181), .ZN(n8462) );
  INV_X1 U7648 ( .A(n6183), .ZN(n6193) );
  INV_X1 U7649 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n6184) );
  OAI22_X1 U7650 ( .A1(n8674), .A2(n8493), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n6184), .ZN(n6195) );
  INV_X1 U7651 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n8460) );
  OAI21_X1 U7652 ( .B1(n6186), .B2(n6184), .A(n8460), .ZN(n6187) );
  NAND2_X1 U7653 ( .A1(P2_REG3_REG_25__SCAN_IN), .A2(P2_REG3_REG_24__SCAN_IN), 
        .ZN(n6185) );
  NAND2_X1 U7654 ( .A1(n6187), .A2(n7999), .ZN(n8628) );
  OR2_X1 U7655 ( .A1(n8628), .A2(n8001), .ZN(n6192) );
  INV_X1 U7656 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n9926) );
  NAND2_X1 U7657 ( .A1(n5871), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n6189) );
  NAND2_X1 U7658 ( .A1(n5843), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n6188) );
  OAI211_X1 U7659 ( .C1(n8154), .C2(n9926), .A(n6189), .B(n6188), .ZN(n6190)
         );
  INV_X1 U7660 ( .A(n6190), .ZN(n6191) );
  INV_X1 U7661 ( .A(n8462), .ZN(n7960) );
  NOR2_X1 U7662 ( .A1(n8644), .A2(n8502), .ZN(n6194) );
  AOI211_X1 U7663 ( .C1(n8496), .C2(n8647), .A(n6195), .B(n6194), .ZN(n6196)
         );
  OAI21_X1 U7664 ( .B1(n4654), .B2(n8499), .A(n6196), .ZN(n6197) );
  NAND2_X1 U7665 ( .A1(n6199), .A2(n6198), .ZN(P2_U3231) );
  INV_X1 U7666 ( .A(n6352), .ZN(n6200) );
  NOR2_X1 U7667 ( .A1(n6357), .A2(n6200), .ZN(n6280) );
  NAND2_X1 U7668 ( .A1(n6387), .A2(n6201), .ZN(n6785) );
  NAND2_X1 U7669 ( .A1(n6357), .A2(n6785), .ZN(n6202) );
  NAND2_X1 U7670 ( .A1(n6202), .A2(n6352), .ZN(n6285) );
  NAND2_X1 U7671 ( .A1(n6285), .A2(n6283), .ZN(n6203) );
  NAND2_X1 U7672 ( .A1(n6203), .A2(P1_STATE_REG_SCAN_IN), .ZN(P1_U3083) );
  INV_X1 U7673 ( .A(n9783), .ZN(n6204) );
  INV_X1 U7674 ( .A(n6205), .ZN(n6206) );
  AOI211_X1 U7675 ( .C1(n6208), .C2(n6207), .A(n8511), .B(n6206), .ZN(n6212)
         );
  INV_X1 U7676 ( .A(n8496), .ZN(n8506) );
  NOR2_X1 U7677 ( .A1(n8506), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n6211) );
  OAI22_X1 U7678 ( .A1(n8499), .A2(n9792), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n5770), .ZN(n6210) );
  INV_X1 U7679 ( .A(n6632), .ZN(n7219) );
  INV_X1 U7680 ( .A(n8529), .ZN(n7218) );
  OAI22_X1 U7681 ( .A1(n8493), .A2(n7219), .B1(n7218), .B2(n8502), .ZN(n6209)
         );
  OR4_X1 U7682 ( .A1(n6212), .A2(n6211), .A3(n6210), .A4(n6209), .ZN(P2_U3220)
         );
  AND2_X1 U7683 ( .A1(n4499), .A2(P2_U3152), .ZN(n7059) );
  NOR2_X1 U7684 ( .A1(n4499), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8877) );
  AOI22_X1 U7685 ( .A1(n8877), .A2(P1_DATAO_REG_1__SCAN_IN), .B1(n8535), .B2(
        P2_STATE_REG_SCAN_IN), .ZN(n6214) );
  OAI21_X1 U7686 ( .B1(n6220), .B2(n4284), .A(n6214), .ZN(P2_U3357) );
  AOI22_X1 U7687 ( .A1(n8877), .A2(P1_DATAO_REG_2__SCAN_IN), .B1(n8548), .B2(
        P2_STATE_REG_SCAN_IN), .ZN(n6215) );
  OAI21_X1 U7688 ( .B1(n6218), .B2(n4284), .A(n6215), .ZN(P2_U3356) );
  INV_X1 U7689 ( .A(n8877), .ZN(n7969) );
  INV_X1 U7690 ( .A(n9688), .ZN(n6499) );
  OAI222_X1 U7691 ( .A1(n7969), .A2(n4436), .B1(n4284), .B2(n4809), .C1(
        P2_U3152), .C2(n6499), .ZN(P2_U3355) );
  AOI22_X1 U7692 ( .A1(n6541), .A2(P2_STATE_REG_SCAN_IN), .B1(n8877), .B2(
        P1_DATAO_REG_4__SCAN_IN), .ZN(n6216) );
  OAI21_X1 U7693 ( .B1(n6222), .B2(n4284), .A(n6216), .ZN(P2_U3354) );
  INV_X1 U7694 ( .A(n6524), .ZN(n6510) );
  OAI222_X1 U7695 ( .A1(n7969), .A2(n6217), .B1(n4284), .B2(n6225), .C1(
        P2_U3152), .C2(n6510), .ZN(P2_U3353) );
  NOR2_X1 U7696 ( .A1(n4279), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9369) );
  INV_X1 U7697 ( .A(n9369), .ZN(n8069) );
  NAND2_X1 U7698 ( .A1(n4280), .A2(P1_U3084), .ZN(n8073) );
  CLKBUF_X1 U7699 ( .A(n8073), .Z(n9371) );
  INV_X1 U7700 ( .A(n6291), .ZN(n6412) );
  OAI222_X1 U7701 ( .A1(n8069), .A2(n6219), .B1(n9371), .B2(n6218), .C1(
        P1_U3084), .C2(n6412), .ZN(P1_U3351) );
  INV_X1 U7702 ( .A(n6289), .ZN(n9010) );
  OAI222_X1 U7703 ( .A1(n8069), .A2(n6221), .B1(n9371), .B2(n6220), .C1(
        P1_U3084), .C2(n9010), .ZN(P1_U3352) );
  INV_X1 U7704 ( .A(n9484), .ZN(n6270) );
  OAI222_X1 U7705 ( .A1(n8069), .A2(n6223), .B1(n9371), .B2(n6222), .C1(
        P1_U3084), .C2(n6270), .ZN(P1_U3349) );
  INV_X1 U7706 ( .A(n9500), .ZN(n6224) );
  OAI222_X1 U7707 ( .A1(n8069), .A2(n9901), .B1(n9371), .B2(n6225), .C1(
        P1_U3084), .C2(n6224), .ZN(P1_U3348) );
  INV_X1 U7708 ( .A(n6294), .ZN(n9023) );
  OAI222_X1 U7709 ( .A1(n8069), .A2(n6226), .B1(n9371), .B2(n4809), .C1(
        P1_U3084), .C2(n9023), .ZN(P1_U3350) );
  INV_X1 U7710 ( .A(n6227), .ZN(n6229) );
  INV_X1 U7711 ( .A(n9507), .ZN(n6273) );
  OAI222_X1 U7712 ( .A1(n8069), .A2(n6228), .B1(n9371), .B2(n6229), .C1(
        P1_U3084), .C2(n6273), .ZN(P1_U3347) );
  INV_X1 U7713 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n6230) );
  INV_X1 U7714 ( .A(n9703), .ZN(n6526) );
  OAI222_X1 U7715 ( .A1(n7969), .A2(n6230), .B1(n4284), .B2(n6229), .C1(
        P2_U3152), .C2(n6526), .ZN(P2_U3352) );
  INV_X1 U7716 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n6232) );
  INV_X1 U7717 ( .A(n6231), .ZN(n6234) );
  INV_X1 U7718 ( .A(n6300), .ZN(n6321) );
  OAI222_X1 U7719 ( .A1(n8069), .A2(n6232), .B1(n9371), .B2(n6234), .C1(
        P1_U3084), .C2(n6321), .ZN(P1_U3346) );
  INV_X1 U7720 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n9897) );
  INV_X1 U7721 ( .A(n9715), .ZN(n6233) );
  OAI222_X1 U7722 ( .A1(n7969), .A2(n9897), .B1(n4284), .B2(n6234), .C1(
        P2_U3152), .C2(n6233), .ZN(P2_U3351) );
  INV_X1 U7723 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n6242) );
  AND3_X1 U7724 ( .A1(n7459), .A2(P1_B_REG_SCAN_IN), .A3(n7165), .ZN(n6238) );
  INV_X1 U7725 ( .A(n7165), .ZN(n6240) );
  INV_X1 U7726 ( .A(P1_B_REG_SCAN_IN), .ZN(n6236) );
  AND2_X1 U7727 ( .A1(n6240), .A2(n6236), .ZN(n6237) );
  OAI22_X1 U7728 ( .A1(n9601), .A2(P1_D_REG_0__SCAN_IN), .B1(n6239), .B2(n6240), .ZN(n9271) );
  INV_X1 U7729 ( .A(n9271), .ZN(n6379) );
  NAND2_X1 U7730 ( .A1(n6379), .A2(n9602), .ZN(n6241) );
  OAI21_X1 U7731 ( .B1(n9602), .B2(n6242), .A(n6241), .ZN(P1_U3440) );
  INV_X1 U7732 ( .A(n6243), .ZN(n6244) );
  INV_X1 U7733 ( .A(n6563), .ZN(n6554) );
  OAI222_X1 U7734 ( .A1(n7969), .A2(n9914), .B1(n4284), .B2(n6244), .C1(
        P2_U3152), .C2(n6554), .ZN(P2_U3350) );
  INV_X1 U7735 ( .A(n6301), .ZN(n6431) );
  OAI222_X1 U7736 ( .A1(n8069), .A2(n9989), .B1(n9371), .B2(n6244), .C1(
        P1_U3084), .C2(n6431), .ZN(P1_U3345) );
  INV_X1 U7737 ( .A(n6245), .ZN(n6247) );
  AOI22_X1 U7738 ( .A1(n9527), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_9__SCAN_IN), .B2(n9369), .ZN(n6246) );
  OAI21_X1 U7739 ( .B1(n6247), .B2(n9371), .A(n6246), .ZN(P1_U3344) );
  INV_X1 U7740 ( .A(n6564), .ZN(n6613) );
  OAI222_X1 U7741 ( .A1(n7969), .A2(n9941), .B1(n4284), .B2(n6247), .C1(n6613), 
        .C2(P2_U3152), .ZN(P2_U3349) );
  INV_X1 U7742 ( .A(n6248), .ZN(n6250) );
  AOI22_X1 U7743 ( .A1(n9536), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n9369), .ZN(n6249) );
  OAI21_X1 U7744 ( .B1(n6250), .B2(n9371), .A(n6249), .ZN(P1_U3343) );
  INV_X1 U7745 ( .A(n9728), .ZN(n6566) );
  OAI222_X1 U7746 ( .A1(n7969), .A2(n6251), .B1(n4284), .B2(n6250), .C1(n6566), 
        .C2(P2_U3152), .ZN(P2_U3348) );
  OR2_X1 U7747 ( .A1(n6252), .A2(P2_U3152), .ZN(n8385) );
  INV_X1 U7748 ( .A(n8385), .ZN(n6254) );
  OAI21_X1 U7749 ( .B1(n9774), .B2(n6254), .A(n6253), .ZN(n6257) );
  NAND2_X1 U7750 ( .A1(n9774), .A2(n6255), .ZN(n6256) );
  INV_X1 U7751 ( .A(n8068), .ZN(n9741) );
  NOR2_X1 U7752 ( .A1(n9741), .A2(P2_U3966), .ZN(P2_U3151) );
  NAND2_X1 U7753 ( .A1(n5871), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n6260) );
  NAND2_X1 U7754 ( .A1(n4276), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n6259) );
  NAND2_X1 U7755 ( .A1(n8013), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n6258) );
  AND3_X1 U7756 ( .A1(n6260), .A2(n6259), .A3(n6258), .ZN(n8162) );
  INV_X1 U7757 ( .A(n8162), .ZN(n8571) );
  NAND2_X1 U7758 ( .A1(n8571), .A2(P2_U3966), .ZN(n6261) );
  OAI21_X1 U7759 ( .B1(P2_U3966), .B2(n5510), .A(n6261), .ZN(P2_U3583) );
  INV_X1 U7760 ( .A(n6262), .ZN(n6311) );
  INV_X1 U7761 ( .A(n9552), .ZN(n6434) );
  OAI222_X1 U7762 ( .A1(n8073), .A2(n6311), .B1(n6434), .B2(P1_U3084), .C1(
        n6263), .C2(n8069), .ZN(P1_U3342) );
  NOR2_X1 U7763 ( .A1(n6300), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n6276) );
  AOI22_X1 U7764 ( .A1(n6300), .A2(n5094), .B1(P1_REG2_REG_7__SCAN_IN), .B2(
        n6321), .ZN(n6317) );
  NAND2_X1 U7765 ( .A1(n9507), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n6275) );
  INV_X1 U7766 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n6264) );
  AND2_X1 U7767 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(
        n9016) );
  NAND2_X1 U7768 ( .A1(n6289), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n6265) );
  INV_X1 U7769 ( .A(n6406), .ZN(n6267) );
  XNOR2_X1 U7770 ( .A(n6291), .B(P1_REG2_REG_2__SCAN_IN), .ZN(n6405) );
  INV_X1 U7771 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n6266) );
  OAI22_X1 U7772 ( .A1(n6267), .A2(n6405), .B1(n6412), .B2(n6266), .ZN(n9026)
         );
  MUX2_X1 U7773 ( .A(P1_REG2_REG_3__SCAN_IN), .B(n6268), .S(n6294), .Z(n9027)
         );
  NAND2_X1 U7774 ( .A1(n9026), .A2(n9027), .ZN(n9025) );
  OAI21_X1 U7775 ( .B1(n9023), .B2(n6268), .A(n9025), .ZN(n9488) );
  MUX2_X1 U7776 ( .A(n6269), .B(P1_REG2_REG_4__SCAN_IN), .S(n9484), .Z(n9487)
         );
  MUX2_X1 U7777 ( .A(n6271), .B(P1_REG2_REG_5__SCAN_IN), .S(n9500), .Z(n9502)
         );
  INV_X1 U7778 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n6274) );
  INV_X1 U7779 ( .A(n6275), .ZN(n6272) );
  AOI21_X1 U7780 ( .B1(n6274), .B2(n6273), .A(n6272), .ZN(n9515) );
  NAND2_X1 U7781 ( .A1(n9514), .A2(n9515), .ZN(n9513) );
  NAND2_X1 U7782 ( .A1(n6275), .A2(n9513), .ZN(n6316) );
  NOR2_X1 U7783 ( .A1(n6317), .A2(n6316), .ZN(n6315) );
  MUX2_X1 U7784 ( .A(P1_REG2_REG_8__SCAN_IN), .B(n7101), .S(n6301), .Z(n6277)
         );
  INV_X1 U7785 ( .A(n6277), .ZN(n6278) );
  AOI21_X1 U7786 ( .B1(n6279), .B2(n6278), .A(n6430), .ZN(n6310) );
  NOR2_X1 U7787 ( .A1(n5683), .A2(P1_U3084), .ZN(n7544) );
  NAND2_X1 U7788 ( .A1(n6285), .A2(n7544), .ZN(n9551) );
  OR2_X1 U7789 ( .A1(n9551), .A2(n5682), .ZN(n9543) );
  INV_X1 U7790 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n6307) );
  OR2_X1 U7791 ( .A1(P1_U3083), .A2(n6280), .ZN(n9571) );
  INV_X1 U7792 ( .A(n9551), .ZN(n6281) );
  AND2_X1 U7793 ( .A1(n6281), .A2(n5682), .ZN(n9553) );
  INV_X1 U7794 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n6282) );
  NOR2_X1 U7795 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6282), .ZN(n7348) );
  AOI21_X1 U7796 ( .B1(n9553), .B2(n6301), .A(n7348), .ZN(n6306) );
  AND2_X1 U7797 ( .A1(n6283), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6284) );
  AND2_X1 U7798 ( .A1(n6285), .A2(n6284), .ZN(n9477) );
  NAND2_X1 U7799 ( .A1(n9477), .A2(n5683), .ZN(n9522) );
  INV_X1 U7800 ( .A(n9522), .ZN(n9566) );
  NOR2_X1 U7801 ( .A1(n6300), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n6286) );
  AOI21_X1 U7802 ( .B1(P1_REG1_REG_7__SCAN_IN), .B2(n6300), .A(n6286), .ZN(
        n6320) );
  XNOR2_X1 U7803 ( .A(n9507), .B(P1_REG1_REG_6__SCAN_IN), .ZN(n9511) );
  XNOR2_X1 U7804 ( .A(n6291), .B(n6287), .ZN(n6409) );
  XNOR2_X1 U7805 ( .A(n6289), .B(n6288), .ZN(n9014) );
  AND2_X1 U7806 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(
        n9013) );
  NAND2_X1 U7807 ( .A1(n9014), .A2(n9013), .ZN(n9012) );
  NAND2_X1 U7808 ( .A1(n6289), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n6290) );
  NAND2_X1 U7809 ( .A1(n9012), .A2(n6290), .ZN(n6408) );
  NAND2_X1 U7810 ( .A1(n6409), .A2(n6408), .ZN(n6407) );
  NAND2_X1 U7811 ( .A1(n6291), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n6292) );
  NAND2_X1 U7812 ( .A1(n6407), .A2(n6292), .ZN(n9029) );
  XNOR2_X1 U7813 ( .A(n6294), .B(n6293), .ZN(n9030) );
  NAND2_X1 U7814 ( .A1(n9029), .A2(n9030), .ZN(n9028) );
  NAND2_X1 U7815 ( .A1(n6294), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n6295) );
  NAND2_X1 U7816 ( .A1(n9028), .A2(n6295), .ZN(n9479) );
  XNOR2_X1 U7817 ( .A(n9484), .B(P1_REG1_REG_4__SCAN_IN), .ZN(n9480) );
  OR2_X1 U7818 ( .A1(n9479), .A2(n9480), .ZN(n9481) );
  OR2_X1 U7819 ( .A1(n9484), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n6296) );
  NAND2_X1 U7820 ( .A1(n9481), .A2(n6296), .ZN(n9497) );
  OR2_X1 U7821 ( .A1(n9500), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n6298) );
  NAND2_X1 U7822 ( .A1(n9500), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n6297) );
  NAND2_X1 U7823 ( .A1(n6298), .A2(n6297), .ZN(n9496) );
  NOR2_X1 U7824 ( .A1(n9497), .A2(n9496), .ZN(n9495) );
  AOI21_X1 U7825 ( .B1(P1_REG1_REG_5__SCAN_IN), .B2(n9500), .A(n9495), .ZN(
        n6299) );
  INV_X1 U7826 ( .A(n6299), .ZN(n9510) );
  OAI22_X1 U7827 ( .A1(n9511), .A2(n9510), .B1(n9507), .B2(
        P1_REG1_REG_6__SCAN_IN), .ZN(n6319) );
  NAND2_X1 U7828 ( .A1(n6320), .A2(n6319), .ZN(n6318) );
  OAI21_X1 U7829 ( .B1(n6300), .B2(P1_REG1_REG_7__SCAN_IN), .A(n6318), .ZN(
        n6303) );
  MUX2_X1 U7830 ( .A(P1_REG1_REG_8__SCAN_IN), .B(n6418), .S(n6301), .Z(n6302)
         );
  NAND2_X1 U7831 ( .A1(n6302), .A2(n6303), .ZN(n6416) );
  OAI21_X1 U7832 ( .B1(n6303), .B2(n6302), .A(n6416), .ZN(n6304) );
  NAND2_X1 U7833 ( .A1(n9566), .A2(n6304), .ZN(n6305) );
  OAI211_X1 U7834 ( .C1(n6307), .C2(n9571), .A(n6306), .B(n6305), .ZN(n6308)
         );
  INV_X1 U7835 ( .A(n6308), .ZN(n6309) );
  OAI21_X1 U7836 ( .B1(n6310), .B2(n9543), .A(n6309), .ZN(P1_U3249) );
  INV_X1 U7837 ( .A(n6562), .ZN(n6712) );
  OAI222_X1 U7838 ( .A1(n7969), .A2(n6312), .B1(n4284), .B2(n6311), .C1(n6712), 
        .C2(P2_U3152), .ZN(P2_U3347) );
  NAND2_X1 U7839 ( .A1(P2_DATAO_REG_15__SCAN_IN), .A2(n8531), .ZN(n6313) );
  OAI21_X1 U7840 ( .B1(n8050), .B2(n8531), .A(n6313), .ZN(P2_U3567) );
  INV_X1 U7841 ( .A(P1_U4006), .ZN(n9009) );
  NAND2_X1 U7842 ( .A1(n9009), .A2(P1_DATAO_REG_14__SCAN_IN), .ZN(n6314) );
  OAI21_X1 U7843 ( .B1(n9401), .B2(n9009), .A(n6314), .ZN(P1_U3569) );
  AOI21_X1 U7844 ( .B1(n6317), .B2(n6316), .A(n6315), .ZN(n6326) );
  OAI21_X1 U7845 ( .B1(n6320), .B2(n6319), .A(n6318), .ZN(n6323) );
  AND2_X1 U7846 ( .A1(P1_U3084), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n6884) );
  INV_X1 U7847 ( .A(n9553), .ZN(n9538) );
  NOR2_X1 U7848 ( .A1(n9538), .A2(n6321), .ZN(n6322) );
  AOI211_X1 U7849 ( .C1(n9566), .C2(n6323), .A(n6884), .B(n6322), .ZN(n6325)
         );
  INV_X1 U7850 ( .A(n9571), .ZN(n9508) );
  NAND2_X1 U7851 ( .A1(n9508), .A2(P1_ADDR_REG_7__SCAN_IN), .ZN(n6324) );
  OAI211_X1 U7852 ( .C1(n6326), .C2(n9543), .A(n6325), .B(n6324), .ZN(P1_U3248) );
  INV_X1 U7853 ( .A(n6327), .ZN(n6329) );
  INV_X1 U7854 ( .A(n6695), .ZN(n6423) );
  OAI222_X1 U7855 ( .A1(n8069), .A2(n6328), .B1(n9371), .B2(n6329), .C1(
        P1_U3084), .C2(n6423), .ZN(P1_U3341) );
  INV_X1 U7856 ( .A(n6586), .ZN(n6600) );
  OAI222_X1 U7857 ( .A1(n7969), .A2(n6330), .B1(n4284), .B2(n6329), .C1(
        P2_U3152), .C2(n6600), .ZN(P2_U3346) );
  INV_X1 U7858 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n6332) );
  NAND2_X1 U7859 ( .A1(n9066), .A2(P1_U4006), .ZN(n6331) );
  OAI21_X1 U7860 ( .B1(P1_U4006), .B2(n6332), .A(n6331), .ZN(P1_U3586) );
  INV_X1 U7861 ( .A(n6333), .ZN(n6335) );
  INV_X1 U7862 ( .A(n6806), .ZN(n6690) );
  OAI222_X1 U7863 ( .A1(n9371), .A2(n6335), .B1(n6690), .B2(P1_U3084), .C1(
        n6334), .C2(n8069), .ZN(P1_U3340) );
  INV_X1 U7864 ( .A(n6575), .ZN(n6674) );
  OAI222_X1 U7865 ( .A1(n7969), .A2(n6336), .B1(n4284), .B2(n6335), .C1(n6674), 
        .C2(P2_U3152), .ZN(P2_U3345) );
  INV_X1 U7866 ( .A(n6337), .ZN(n6374) );
  OAI222_X1 U7867 ( .A1(n9371), .A2(n6374), .B1(n7258), .B2(P1_U3084), .C1(
        n6338), .C2(n8069), .ZN(P1_U3339) );
  INV_X1 U7868 ( .A(n7459), .ZN(n6339) );
  OAI22_X1 U7869 ( .A1(n9601), .A2(P1_D_REG_1__SCAN_IN), .B1(n6239), .B2(n6339), .ZN(n6754) );
  INV_X1 U7870 ( .A(n9601), .ZN(n6350) );
  NOR4_X1 U7871 ( .A1(P1_D_REG_3__SCAN_IN), .A2(P1_D_REG_4__SCAN_IN), .A3(
        P1_D_REG_5__SCAN_IN), .A4(P1_D_REG_6__SCAN_IN), .ZN(n6348) );
  NOR4_X1 U7872 ( .A1(P1_D_REG_9__SCAN_IN), .A2(P1_D_REG_10__SCAN_IN), .A3(
        P1_D_REG_11__SCAN_IN), .A4(P1_D_REG_12__SCAN_IN), .ZN(n6347) );
  INV_X1 U7873 ( .A(P1_D_REG_2__SCAN_IN), .ZN(n9898) );
  INV_X1 U7874 ( .A(P1_D_REG_7__SCAN_IN), .ZN(n9913) );
  INV_X1 U7875 ( .A(P1_D_REG_13__SCAN_IN), .ZN(n9944) );
  INV_X1 U7876 ( .A(P1_D_REG_8__SCAN_IN), .ZN(n9979) );
  NAND4_X1 U7877 ( .A1(n9898), .A2(n9913), .A3(n9944), .A4(n9979), .ZN(n6345)
         );
  NOR4_X1 U7878 ( .A1(P1_D_REG_18__SCAN_IN), .A2(P1_D_REG_19__SCAN_IN), .A3(
        P1_D_REG_20__SCAN_IN), .A4(P1_D_REG_21__SCAN_IN), .ZN(n6343) );
  NOR4_X1 U7879 ( .A1(P1_D_REG_16__SCAN_IN), .A2(P1_D_REG_14__SCAN_IN), .A3(
        P1_D_REG_15__SCAN_IN), .A4(P1_D_REG_17__SCAN_IN), .ZN(n6342) );
  NOR4_X1 U7880 ( .A1(P1_D_REG_26__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n6341) );
  NOR4_X1 U7881 ( .A1(P1_D_REG_22__SCAN_IN), .A2(P1_D_REG_23__SCAN_IN), .A3(
        P1_D_REG_24__SCAN_IN), .A4(P1_D_REG_25__SCAN_IN), .ZN(n6340) );
  NAND4_X1 U7882 ( .A1(n6343), .A2(n6342), .A3(n6341), .A4(n6340), .ZN(n6344)
         );
  NOR4_X1 U7883 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        n6345), .A4(n6344), .ZN(n6346) );
  NAND3_X1 U7884 ( .A1(n6348), .A2(n6347), .A3(n6346), .ZN(n6349) );
  NAND2_X1 U7885 ( .A1(n6350), .A2(n6349), .ZN(n6377) );
  INV_X1 U7886 ( .A(n6377), .ZN(n6351) );
  OR3_X1 U7887 ( .A1(n9271), .A2(n6754), .A3(n6351), .ZN(n6371) );
  NAND2_X1 U7888 ( .A1(n7004), .A2(n6976), .ZN(n6761) );
  NOR2_X1 U7889 ( .A1(n6761), .A2(n5664), .ZN(n9590) );
  OR2_X1 U7890 ( .A1(n6785), .A2(n6354), .ZN(n6376) );
  NAND3_X1 U7891 ( .A1(n6376), .A2(n6357), .A3(n6352), .ZN(n6353) );
  AOI21_X1 U7892 ( .B1(n6371), .B2(n9590), .A(n6353), .ZN(n6659) );
  AND2_X1 U7893 ( .A1(n6659), .A2(P1_STATE_REG_SCAN_IN), .ZN(n7347) );
  INV_X1 U7894 ( .A(n6761), .ZN(n6380) );
  NAND2_X1 U7895 ( .A1(n6371), .A2(n9658), .ZN(n6658) );
  AND2_X1 U7896 ( .A1(n7347), .A2(n6658), .ZN(n6469) );
  INV_X1 U7897 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n6758) );
  AND2_X1 U7898 ( .A1(n7004), .A2(n6354), .ZN(n6355) );
  NAND2_X1 U7899 ( .A1(n6360), .A2(n7904), .ZN(n6365) );
  INV_X1 U7900 ( .A(n6388), .ZN(n6356) );
  NAND2_X2 U7901 ( .A1(n6357), .A2(n6356), .ZN(n6359) );
  INV_X1 U7902 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n9474) );
  NOR2_X1 U7903 ( .A1(n6357), .A2(n9474), .ZN(n6358) );
  AOI21_X1 U7904 ( .B1(n6778), .B2(n7939), .A(n6358), .ZN(n6364) );
  AND2_X1 U7905 ( .A1(n6365), .A2(n6364), .ZN(n6366) );
  NAND2_X1 U7906 ( .A1(n6360), .A2(n7939), .ZN(n6363) );
  NOR2_X1 U7907 ( .A1(n6357), .A2(n9473), .ZN(n6361) );
  NAND3_X1 U7908 ( .A1(n6365), .A2(n6390), .A3(n6364), .ZN(n6392) );
  OAI21_X1 U7909 ( .B1(n6366), .B2(n6390), .A(n6392), .ZN(n6402) );
  INV_X1 U7910 ( .A(n6371), .ZN(n6369) );
  NAND2_X1 U7911 ( .A1(n9602), .A2(n6785), .ZN(n6367) );
  NOR2_X1 U7912 ( .A1(n6367), .A2(n9345), .ZN(n6368) );
  NAND2_X1 U7913 ( .A1(n6369), .A2(n6368), .ZN(n8984) );
  INV_X1 U7914 ( .A(n8984), .ZN(n8973) );
  AOI22_X1 U7915 ( .A1(n6402), .A2(n8973), .B1(n8968), .B2(n6778), .ZN(n6373)
         );
  NAND2_X1 U7916 ( .A1(n9602), .A2(n4344), .ZN(n6370) );
  NOR2_X1 U7917 ( .A1(n6371), .A2(n6370), .ZN(n6397) );
  NAND2_X1 U7918 ( .A1(n6397), .A2(n5682), .ZN(n8963) );
  NAND2_X1 U7919 ( .A1(n8994), .A2(n6897), .ZN(n6372) );
  OAI211_X1 U7920 ( .C1(n6469), .C2(n6758), .A(n6373), .B(n6372), .ZN(P1_U3230) );
  INV_X1 U7921 ( .A(n7149), .ZN(n7141) );
  OAI222_X1 U7922 ( .A1(n7969), .A2(n6375), .B1(n4284), .B2(n6374), .C1(n7141), 
        .C2(P2_U3152), .ZN(P2_U3344) );
  NAND3_X1 U7923 ( .A1(n6377), .A2(n9602), .A3(n6376), .ZN(n6755) );
  OR2_X1 U7924 ( .A1(n6761), .A2(n9277), .ZN(n9660) );
  OAI21_X1 U7925 ( .B1(n9660), .B2(n9141), .A(n6754), .ZN(n6378) );
  OR2_X1 U7926 ( .A1(n6755), .A2(n6378), .ZN(n9272) );
  INV_X2 U7927 ( .A(n9666), .ZN(n9470) );
  NOR2_X1 U7928 ( .A1(n4344), .A2(n6380), .ZN(n6381) );
  OR2_X1 U7929 ( .A1(n6785), .A2(n6786), .ZN(n9576) );
  AOI22_X1 U7930 ( .A1(n6382), .A2(n6381), .B1(n9261), .B2(n6897), .ZN(n6757)
         );
  OAI21_X1 U7931 ( .B1(n6794), .B2(n6761), .A(n6757), .ZN(n9349) );
  NAND2_X1 U7932 ( .A1(n9349), .A2(n9470), .ZN(n6383) );
  OAI21_X1 U7933 ( .B1(n9470), .B2(n5008), .A(n6383), .ZN(P1_U3454) );
  NAND2_X1 U7934 ( .A1(n6897), .A2(n7939), .ZN(n6386) );
  NAND2_X1 U7935 ( .A1(n6386), .A2(n6385), .ZN(n6389) );
  XNOR2_X1 U7936 ( .A(n6389), .B(n7936), .ZN(n6454) );
  INV_X1 U7937 ( .A(n6454), .ZN(n6458) );
  INV_X1 U7938 ( .A(n6390), .ZN(n6391) );
  NAND2_X1 U7939 ( .A1(n6391), .A2(n6860), .ZN(n6393) );
  NAND2_X1 U7940 ( .A1(n6393), .A2(n6392), .ZN(n6457) );
  NAND2_X1 U7941 ( .A1(n6897), .A2(n7904), .ZN(n6395) );
  INV_X1 U7942 ( .A(n6795), .ZN(n6896) );
  NAND2_X1 U7943 ( .A1(n6896), .A2(n7939), .ZN(n6394) );
  NAND2_X1 U7944 ( .A1(n6395), .A2(n6394), .ZN(n6455) );
  XNOR2_X1 U7945 ( .A(n6457), .B(n6455), .ZN(n6396) );
  XNOR2_X1 U7946 ( .A(n6458), .B(n6396), .ZN(n6401) );
  NOR2_X1 U7947 ( .A1(n6795), .A2(n9658), .ZN(n9605) );
  AND2_X2 U7948 ( .A1(n6397), .A2(n6786), .ZN(n8965) );
  INV_X1 U7949 ( .A(n8965), .ZN(n8991) );
  INV_X1 U7950 ( .A(n6360), .ZN(n6789) );
  INV_X1 U7951 ( .A(n6448), .ZN(n6788) );
  OAI22_X1 U7952 ( .A1(n8991), .A2(n6789), .B1(n6788), .B2(n8963), .ZN(n6399)
         );
  NOR2_X1 U7953 ( .A1(n6469), .A2(n6796), .ZN(n6398) );
  AOI211_X1 U7954 ( .C1(n7347), .C2(n9605), .A(n6399), .B(n6398), .ZN(n6400)
         );
  OAI21_X1 U7955 ( .B1(n8984), .B2(n6401), .A(n6400), .ZN(P1_U3220) );
  MUX2_X1 U7956 ( .A(n9474), .B(n6402), .S(n5683), .Z(n6404) );
  OAI21_X1 U7957 ( .B1(n5683), .B2(P1_REG2_REG_0__SCAN_IN), .A(n6786), .ZN(
        n9472) );
  NAND2_X1 U7958 ( .A1(n9472), .A2(n9474), .ZN(n6403) );
  OAI211_X1 U7959 ( .C1(n6404), .C2(n9472), .A(P1_U4006), .B(n6403), .ZN(n9492) );
  XOR2_X1 U7960 ( .A(n6406), .B(n6405), .Z(n6411) );
  OAI211_X1 U7961 ( .C1(n6409), .C2(n6408), .A(n9566), .B(n6407), .ZN(n6410)
         );
  OAI21_X1 U7962 ( .B1(n6411), .B2(n9543), .A(n6410), .ZN(n6414) );
  OAI22_X1 U7963 ( .A1(n9538), .A2(n6412), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n6468), .ZN(n6413) );
  AOI211_X1 U7964 ( .C1(n9508), .C2(P1_ADDR_REG_2__SCAN_IN), .A(n6414), .B(
        n6413), .ZN(n6415) );
  NAND2_X1 U7965 ( .A1(n9492), .A2(n6415), .ZN(P1_U3243) );
  INV_X1 U7966 ( .A(n6416), .ZN(n6417) );
  AOI21_X1 U7967 ( .B1(n6418), .B2(n6431), .A(n6417), .ZN(n9521) );
  INV_X1 U7968 ( .A(n9521), .ZN(n6420) );
  MUX2_X1 U7969 ( .A(n5133), .B(P1_REG1_REG_9__SCAN_IN), .S(n9527), .Z(n9520)
         );
  INV_X1 U7970 ( .A(n9520), .ZN(n6419) );
  NAND2_X1 U7971 ( .A1(n6420), .A2(n6419), .ZN(n9524) );
  OAI21_X1 U7972 ( .B1(n9527), .B2(P1_REG1_REG_9__SCAN_IN), .A(n9524), .ZN(
        n9534) );
  MUX2_X1 U7973 ( .A(P1_REG1_REG_10__SCAN_IN), .B(n6421), .S(n9536), .Z(n9535)
         );
  NAND2_X1 U7974 ( .A1(n9534), .A2(n9535), .ZN(n9533) );
  OAI21_X1 U7975 ( .B1(n9536), .B2(P1_REG1_REG_10__SCAN_IN), .A(n9533), .ZN(
        n9563) );
  MUX2_X1 U7976 ( .A(P1_REG1_REG_11__SCAN_IN), .B(n6422), .S(n9552), .Z(n9564)
         );
  NAND2_X1 U7977 ( .A1(n9563), .A2(n9564), .ZN(n9562) );
  OAI21_X1 U7978 ( .B1(P1_REG1_REG_11__SCAN_IN), .B2(n9552), .A(n9562), .ZN(
        n6425) );
  AOI22_X1 U7979 ( .A1(n6695), .A2(P1_REG1_REG_12__SCAN_IN), .B1(n5184), .B2(
        n6423), .ZN(n6424) );
  NAND2_X1 U7980 ( .A1(n6424), .A2(n6425), .ZN(n6689) );
  OAI21_X1 U7981 ( .B1(n6425), .B2(n6424), .A(n6689), .ZN(n6440) );
  INV_X1 U7982 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n6428) );
  NAND2_X1 U7983 ( .A1(P1_REG3_REG_12__SCAN_IN), .A2(P1_U3084), .ZN(n7640) );
  INV_X1 U7984 ( .A(n7640), .ZN(n6426) );
  AOI21_X1 U7985 ( .B1(n9553), .B2(n6695), .A(n6426), .ZN(n6427) );
  OAI21_X1 U7986 ( .B1(n9571), .B2(n6428), .A(n6427), .ZN(n6439) );
  NAND2_X1 U7987 ( .A1(n9527), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n6432) );
  MUX2_X1 U7988 ( .A(n5132), .B(P1_REG2_REG_9__SCAN_IN), .S(n9527), .Z(n6429)
         );
  INV_X1 U7989 ( .A(n6429), .ZN(n9529) );
  INV_X1 U7990 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n6433) );
  MUX2_X1 U7991 ( .A(n6433), .B(P1_REG2_REG_10__SCAN_IN), .S(n9536), .Z(n9545)
         );
  AOI21_X1 U7992 ( .B1(P1_REG2_REG_10__SCAN_IN), .B2(n9536), .A(n9542), .ZN(
        n9555) );
  OAI21_X1 U7993 ( .B1(n9550), .B2(n6434), .A(n9555), .ZN(n6435) );
  OR2_X1 U7994 ( .A1(n9552), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n9558) );
  NAND2_X1 U7995 ( .A1(n6695), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n6436) );
  OAI21_X1 U7996 ( .B1(n6695), .B2(P1_REG2_REG_12__SCAN_IN), .A(n6436), .ZN(
        n6437) );
  AOI211_X1 U7997 ( .C1(n9557), .C2(n6437), .A(n6694), .B(n9543), .ZN(n6438)
         );
  AOI211_X1 U7998 ( .C1(n6440), .C2(n9566), .A(n6439), .B(n6438), .ZN(n6441)
         );
  INV_X1 U7999 ( .A(n6441), .ZN(P1_U3253) );
  INV_X1 U8000 ( .A(n6442), .ZN(n6445) );
  AOI22_X1 U8001 ( .A1(n7533), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_15__SCAN_IN), .B2(n9369), .ZN(n6443) );
  OAI21_X1 U8002 ( .B1(n6445), .B2(n9371), .A(n6443), .ZN(P1_U3338) );
  AOI22_X1 U8003 ( .A1(n8564), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_15__SCAN_IN), .B2(n8877), .ZN(n6444) );
  OAI21_X1 U8004 ( .B1(n6445), .B2(n4284), .A(n6444), .ZN(P2_U3343) );
  INV_X1 U8005 ( .A(n6446), .ZN(n6550) );
  AOI22_X1 U8006 ( .A1(n7728), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(n9369), .ZN(n6447) );
  OAI21_X1 U8007 ( .B1(n6550), .B2(n9371), .A(n6447), .ZN(P1_U3337) );
  NAND2_X1 U8008 ( .A1(n6448), .A2(n7939), .ZN(n6450) );
  NAND2_X1 U8009 ( .A1(n6937), .A2(n7933), .ZN(n6449) );
  NAND2_X1 U8010 ( .A1(n6450), .A2(n6449), .ZN(n6451) );
  XNOR2_X1 U8011 ( .A(n6451), .B(n7936), .ZN(n6453) );
  AOI22_X1 U8012 ( .A1(n6448), .A2(n7904), .B1(n6937), .B2(n7939), .ZN(n6452)
         );
  NAND2_X1 U8013 ( .A1(n6453), .A2(n6452), .ZN(n6654) );
  NAND2_X1 U8014 ( .A1(n6654), .A2(n4307), .ZN(n6463) );
  NAND2_X1 U8015 ( .A1(n6454), .A2(n6457), .ZN(n6456) );
  NAND2_X1 U8016 ( .A1(n6456), .A2(n6455), .ZN(n6461) );
  INV_X1 U8017 ( .A(n6457), .ZN(n6459) );
  NAND2_X1 U8018 ( .A1(n6459), .A2(n6458), .ZN(n6460) );
  NAND2_X1 U8019 ( .A1(n6461), .A2(n6460), .ZN(n6462) );
  INV_X1 U8020 ( .A(n6462), .ZN(n6465) );
  INV_X1 U8021 ( .A(n6463), .ZN(n6464) );
  NAND2_X1 U8022 ( .A1(n6465), .A2(n6464), .ZN(n6655) );
  INV_X1 U8023 ( .A(n6655), .ZN(n6466) );
  AOI21_X1 U8024 ( .B1(n6463), .B2(n6462), .A(n6466), .ZN(n6472) );
  AOI22_X1 U8025 ( .A1(n8994), .A2(n9008), .B1(n8965), .B2(n6897), .ZN(n6467)
         );
  OAI21_X1 U8026 ( .B1(n6469), .B2(n6468), .A(n6467), .ZN(n6470) );
  AOI21_X1 U8027 ( .B1(n8968), .B2(n6937), .A(n6470), .ZN(n6471) );
  OAI21_X1 U8028 ( .B1(n6472), .B2(n8984), .A(n6471), .ZN(P1_U3235) );
  NAND2_X1 U8029 ( .A1(n9774), .A2(n6628), .ZN(n6476) );
  OR2_X1 U8030 ( .A1(n6183), .A2(P2_U3152), .ZN(n7671) );
  OAI21_X1 U8031 ( .B1(n6473), .B2(n7671), .A(n8385), .ZN(n6474) );
  INV_X1 U8032 ( .A(n6474), .ZN(n6475) );
  NAND2_X1 U8033 ( .A1(n6476), .A2(n6475), .ZN(n6479) );
  NAND2_X1 U8034 ( .A1(n6479), .A2(n5753), .ZN(n6477) );
  NAND2_X1 U8035 ( .A1(n6477), .A2(n8531), .ZN(n6496) );
  INV_X1 U8036 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n6494) );
  AND2_X1 U8037 ( .A1(n5753), .A2(n8407), .ZN(n6478) );
  INV_X1 U8038 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n9831) );
  MUX2_X1 U8039 ( .A(n9831), .B(P2_REG1_REG_5__SCAN_IN), .S(n6524), .Z(n6488)
         );
  INV_X1 U8040 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n6480) );
  MUX2_X1 U8041 ( .A(P2_REG1_REG_2__SCAN_IN), .B(n6480), .S(n8548), .Z(n6482)
         );
  MUX2_X1 U8042 ( .A(P2_REG1_REG_1__SCAN_IN), .B(n5742), .S(n8535), .Z(n8536)
         );
  AND2_X1 U8043 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(
        n8537) );
  NAND2_X1 U8044 ( .A1(n8536), .A2(n8537), .ZN(n8549) );
  NAND2_X1 U8045 ( .A1(n8535), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n8550) );
  NAND2_X1 U8046 ( .A1(n8549), .A2(n8550), .ZN(n6481) );
  NAND2_X1 U8047 ( .A1(n6482), .A2(n6481), .ZN(n8553) );
  NAND2_X1 U8048 ( .A1(n8548), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n6483) );
  NAND2_X1 U8049 ( .A1(n8553), .A2(n6483), .ZN(n9691) );
  INV_X1 U8050 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n6484) );
  MUX2_X1 U8051 ( .A(P2_REG1_REG_3__SCAN_IN), .B(n6484), .S(n9688), .Z(n9690)
         );
  NAND2_X1 U8052 ( .A1(n9691), .A2(n9690), .ZN(n9689) );
  NAND2_X1 U8053 ( .A1(n9688), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n6535) );
  NAND2_X1 U8054 ( .A1(n9689), .A2(n6535), .ZN(n6487) );
  INV_X1 U8055 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n6485) );
  MUX2_X1 U8056 ( .A(P2_REG1_REG_4__SCAN_IN), .B(n6485), .S(n6541), .Z(n6486)
         );
  NAND2_X1 U8057 ( .A1(n6487), .A2(n6486), .ZN(n6537) );
  NAND2_X1 U8058 ( .A1(n6541), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n6489) );
  NAND3_X1 U8059 ( .A1(n6488), .A2(n6537), .A3(n6489), .ZN(n6492) );
  NAND2_X1 U8060 ( .A1(n6537), .A2(n6489), .ZN(n6491) );
  MUX2_X1 U8061 ( .A(P2_REG1_REG_5__SCAN_IN), .B(n9831), .S(n6524), .Z(n6490)
         );
  NAND2_X1 U8062 ( .A1(n6491), .A2(n6490), .ZN(n6509) );
  NAND3_X1 U8063 ( .A1(n9748), .A2(n6492), .A3(n6509), .ZN(n6493) );
  NAND2_X1 U8064 ( .A1(P2_REG3_REG_5__SCAN_IN), .A2(P2_U3152), .ZN(n6849) );
  OAI211_X1 U8065 ( .C1(n8068), .C2(n6494), .A(n6493), .B(n6849), .ZN(n6506)
         );
  NOR2_X1 U8066 ( .A1(n6183), .A2(n8407), .ZN(n6495) );
  NAND2_X1 U8067 ( .A1(n6496), .A2(n6495), .ZN(n9692) );
  NAND2_X1 U8068 ( .A1(n8535), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n8544) );
  INV_X1 U8069 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n6497) );
  MUX2_X1 U8070 ( .A(P2_REG2_REG_1__SCAN_IN), .B(n6497), .S(n8535), .Z(n8533)
         );
  NAND3_X1 U8071 ( .A1(n8533), .A2(P2_REG2_REG_0__SCAN_IN), .A3(
        P2_IR_REG_0__SCAN_IN), .ZN(n8543) );
  INV_X1 U8072 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n6498) );
  MUX2_X1 U8073 ( .A(n6498), .B(P2_REG2_REG_2__SCAN_IN), .S(n8548), .Z(n8545)
         );
  AOI21_X1 U8074 ( .B1(n8544), .B2(n8543), .A(n8545), .ZN(n8542) );
  AOI21_X1 U8075 ( .B1(n8548), .B2(P2_REG2_REG_2__SCAN_IN), .A(n8542), .ZN(
        n9695) );
  INV_X1 U8076 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n7210) );
  MUX2_X1 U8077 ( .A(n7210), .B(P2_REG2_REG_3__SCAN_IN), .S(n9688), .Z(n9694)
         );
  NOR2_X1 U8078 ( .A1(n9695), .A2(n9694), .ZN(n9693) );
  NOR2_X1 U8079 ( .A1(n6499), .A2(n7210), .ZN(n6542) );
  INV_X1 U8080 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n6500) );
  MUX2_X1 U8081 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n6500), .S(n6541), .Z(n6501)
         );
  NAND2_X1 U8082 ( .A1(n6541), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n6503) );
  INV_X1 U8083 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n7236) );
  MUX2_X1 U8084 ( .A(n7236), .B(P2_REG2_REG_5__SCAN_IN), .S(n6524), .Z(n6502)
         );
  AND3_X1 U8085 ( .A1(n6545), .A2(n6503), .A3(n6502), .ZN(n6504) );
  NOR3_X1 U8086 ( .A1(n9692), .A2(n6504), .A3(n6523), .ZN(n6505) );
  AOI211_X1 U8087 ( .C1(n9747), .C2(n6524), .A(n6506), .B(n6505), .ZN(n6507)
         );
  INV_X1 U8088 ( .A(n6507), .ZN(P2_U3250) );
  INV_X1 U8089 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n6520) );
  NAND2_X1 U8090 ( .A1(n9715), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n6512) );
  INV_X1 U8091 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n6508) );
  MUX2_X1 U8092 ( .A(P2_REG1_REG_7__SCAN_IN), .B(n6508), .S(n9715), .Z(n9717)
         );
  INV_X1 U8093 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n6511) );
  OAI21_X1 U8094 ( .B1(n9831), .B2(n6510), .A(n6509), .ZN(n9706) );
  MUX2_X1 U8095 ( .A(P2_REG1_REG_6__SCAN_IN), .B(n6511), .S(n9703), .Z(n9705)
         );
  NAND2_X1 U8096 ( .A1(n9706), .A2(n9705), .ZN(n9704) );
  OAI21_X1 U8097 ( .B1(n6526), .B2(n6511), .A(n9704), .ZN(n9718) );
  NAND2_X1 U8098 ( .A1(n9717), .A2(n9718), .ZN(n9716) );
  NAND2_X1 U8099 ( .A1(n6512), .A2(n9716), .ZN(n6515) );
  INV_X1 U8100 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n6513) );
  MUX2_X1 U8101 ( .A(P2_REG1_REG_8__SCAN_IN), .B(n6513), .S(n6563), .Z(n6514)
         );
  NAND2_X1 U8102 ( .A1(n6515), .A2(n6514), .ZN(n6603) );
  INV_X1 U8103 ( .A(n6515), .ZN(n6517) );
  MUX2_X1 U8104 ( .A(n6513), .B(P2_REG1_REG_8__SCAN_IN), .S(n6563), .Z(n6516)
         );
  NAND2_X1 U8105 ( .A1(n6517), .A2(n6516), .ZN(n6518) );
  NAND3_X1 U8106 ( .A1(n9748), .A2(n6603), .A3(n6518), .ZN(n6519) );
  NAND2_X1 U8107 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(P2_U3152), .ZN(n6826) );
  OAI211_X1 U8108 ( .C1(n8068), .C2(n6520), .A(n6519), .B(n6826), .ZN(n6532)
         );
  NAND2_X1 U8109 ( .A1(n9715), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n6527) );
  INV_X1 U8110 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n6521) );
  MUX2_X1 U8111 ( .A(n6521), .B(P2_REG2_REG_7__SCAN_IN), .S(n9715), .Z(n6522)
         );
  INV_X1 U8112 ( .A(n6522), .ZN(n9720) );
  INV_X1 U8113 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n6525) );
  MUX2_X1 U8114 ( .A(n6525), .B(P2_REG2_REG_6__SCAN_IN), .S(n9703), .Z(n9707)
         );
  OAI21_X1 U8115 ( .B1(n6526), .B2(n6525), .A(n9708), .ZN(n9721) );
  NAND2_X1 U8116 ( .A1(n9720), .A2(n9721), .ZN(n9719) );
  INV_X1 U8117 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n6528) );
  MUX2_X1 U8118 ( .A(n6528), .B(P2_REG2_REG_8__SCAN_IN), .S(n6563), .Z(n6529)
         );
  AOI211_X1 U8119 ( .C1(n6530), .C2(n6529), .A(n6553), .B(n9692), .ZN(n6531)
         );
  AOI211_X1 U8120 ( .C1(n9747), .C2(n6563), .A(n6532), .B(n6531), .ZN(n6533)
         );
  INV_X1 U8121 ( .A(n6533), .ZN(P2_U3253) );
  INV_X1 U8122 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n6539) );
  MUX2_X1 U8123 ( .A(n6485), .B(P2_REG1_REG_4__SCAN_IN), .S(n6541), .Z(n6534)
         );
  NAND3_X1 U8124 ( .A1(n9689), .A2(n6535), .A3(n6534), .ZN(n6536) );
  NAND3_X1 U8125 ( .A1(n9748), .A2(n6537), .A3(n6536), .ZN(n6538) );
  NAND2_X1 U8126 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_U3152), .ZN(n6834) );
  OAI211_X1 U8127 ( .C1(n8068), .C2(n6539), .A(n6538), .B(n6834), .ZN(n6540)
         );
  AOI21_X1 U8128 ( .B1(n6541), .B2(n9747), .A(n6540), .ZN(n6548) );
  MUX2_X1 U8129 ( .A(n6500), .B(P2_REG2_REG_4__SCAN_IN), .S(n6541), .Z(n6544)
         );
  INV_X1 U8130 ( .A(n6542), .ZN(n6543) );
  NAND2_X1 U8131 ( .A1(n6544), .A2(n6543), .ZN(n6546) );
  OAI211_X1 U8132 ( .C1(n9693), .C2(n6546), .A(n9744), .B(n6545), .ZN(n6547)
         );
  NAND2_X1 U8133 ( .A1(n6548), .A2(n6547), .ZN(P2_U3249) );
  OAI222_X1 U8134 ( .A1(P2_U3152), .A2(n7620), .B1(n4284), .B2(n6550), .C1(
        n6549), .C2(n7969), .ZN(P2_U3342) );
  NAND2_X1 U8135 ( .A1(n6586), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n6559) );
  INV_X1 U8136 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n6587) );
  NOR2_X1 U8137 ( .A1(P2_REG2_REG_11__SCAN_IN), .A2(n6562), .ZN(n6558) );
  NAND2_X1 U8138 ( .A1(n9728), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n6556) );
  INV_X1 U8139 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n6551) );
  MUX2_X1 U8140 ( .A(n6551), .B(P2_REG2_REG_10__SCAN_IN), .S(n9728), .Z(n6552)
         );
  INV_X1 U8141 ( .A(n6552), .ZN(n9734) );
  INV_X1 U8142 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n6555) );
  MUX2_X1 U8143 ( .A(P2_REG2_REG_9__SCAN_IN), .B(n6555), .S(n6564), .Z(n6609)
         );
  NAND2_X1 U8144 ( .A1(n6609), .A2(n6610), .ZN(n6608) );
  OAI21_X1 U8145 ( .B1(n6613), .B2(n6555), .A(n6608), .ZN(n9733) );
  NAND2_X1 U8146 ( .A1(n9734), .A2(n9733), .ZN(n9732) );
  INV_X1 U8147 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n6557) );
  AOI22_X1 U8148 ( .A1(P2_REG2_REG_11__SCAN_IN), .A2(n6712), .B1(n6562), .B2(
        n6557), .ZN(n6704) );
  NAND2_X1 U8149 ( .A1(n6559), .A2(n6588), .ZN(n6561) );
  INV_X1 U8150 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n6668) );
  AOI22_X1 U8151 ( .A1(P2_REG2_REG_13__SCAN_IN), .A2(n6674), .B1(n6575), .B2(
        n6668), .ZN(n6560) );
  NOR2_X1 U8152 ( .A1(n6561), .A2(n6560), .ZN(n6667) );
  AOI21_X1 U8153 ( .B1(n6561), .B2(n6560), .A(n6667), .ZN(n6577) );
  INV_X1 U8154 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n9972) );
  MUX2_X1 U8155 ( .A(P2_REG1_REG_12__SCAN_IN), .B(n9972), .S(n6586), .Z(n6594)
         );
  INV_X1 U8156 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n9838) );
  MUX2_X1 U8157 ( .A(P2_REG1_REG_11__SCAN_IN), .B(n9838), .S(n6562), .Z(n6709)
         );
  INV_X1 U8158 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n7088) );
  MUX2_X1 U8159 ( .A(P2_REG1_REG_10__SCAN_IN), .B(n7088), .S(n9728), .Z(n9730)
         );
  INV_X1 U8160 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n9834) );
  NAND2_X1 U8161 ( .A1(n6563), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n6602) );
  MUX2_X1 U8162 ( .A(n9834), .B(P2_REG1_REG_9__SCAN_IN), .S(n6564), .Z(n6601)
         );
  AOI21_X1 U8163 ( .B1(n6603), .B2(n6602), .A(n6601), .ZN(n6605) );
  INV_X1 U8164 ( .A(n6605), .ZN(n6565) );
  OAI21_X1 U8165 ( .B1(n9834), .B2(n6613), .A(n6565), .ZN(n9731) );
  NAND2_X1 U8166 ( .A1(n9730), .A2(n9731), .ZN(n9729) );
  OAI21_X1 U8167 ( .B1(n6566), .B2(n7088), .A(n9729), .ZN(n6708) );
  NAND2_X1 U8168 ( .A1(n6709), .A2(n6708), .ZN(n6707) );
  OAI21_X1 U8169 ( .B1(n6712), .B2(n9838), .A(n6707), .ZN(n6567) );
  INV_X1 U8170 ( .A(n6567), .ZN(n6593) );
  AOI21_X1 U8171 ( .B1(n9972), .B2(n6600), .A(n6591), .ZN(n6569) );
  INV_X1 U8172 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n9388) );
  AOI22_X1 U8173 ( .A1(P2_REG1_REG_13__SCAN_IN), .A2(n6674), .B1(n6575), .B2(
        n9388), .ZN(n6568) );
  NOR2_X1 U8174 ( .A1(n6569), .A2(n6568), .ZN(n6673) );
  AOI21_X1 U8175 ( .B1(n6569), .B2(n6568), .A(n6673), .ZN(n6573) );
  INV_X1 U8176 ( .A(n9748), .ZN(n9681) );
  NOR2_X1 U8177 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6570), .ZN(n6571) );
  AOI21_X1 U8178 ( .B1(n9741), .B2(P2_ADDR_REG_13__SCAN_IN), .A(n6571), .ZN(
        n6572) );
  OAI21_X1 U8179 ( .B1(n6573), .B2(n9681), .A(n6572), .ZN(n6574) );
  AOI21_X1 U8180 ( .B1(n6575), .B2(n9747), .A(n6574), .ZN(n6576) );
  OAI21_X1 U8181 ( .B1(n6577), .B2(n9692), .A(n6576), .ZN(P2_U3258) );
  NOR2_X1 U8182 ( .A1(n6735), .A2(P2_U3152), .ZN(n7976) );
  INV_X1 U8183 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n6585) );
  INV_X1 U8184 ( .A(n6644), .ZN(n6636) );
  INV_X1 U8185 ( .A(n8753), .ZN(n8719) );
  OAI22_X1 U8186 ( .A1(n6636), .A2(n8719), .B1(n7219), .B2(n8721), .ZN(n9757)
         );
  AOI22_X1 U8187 ( .A1(n8509), .A2(n6578), .B1(n8462), .B2(n9757), .ZN(n6584)
         );
  OAI21_X1 U8188 ( .B1(n6581), .B2(n6580), .A(n6579), .ZN(n6582) );
  NAND2_X1 U8189 ( .A1(n6582), .A2(n8473), .ZN(n6583) );
  OAI211_X1 U8190 ( .C1(n7976), .C2(n6585), .A(n6584), .B(n6583), .ZN(P2_U3224) );
  INV_X1 U8191 ( .A(n9747), .ZN(n9680) );
  MUX2_X1 U8192 ( .A(P2_REG2_REG_12__SCAN_IN), .B(n6587), .S(n6586), .Z(n6589)
         );
  OAI211_X1 U8193 ( .C1(n6590), .C2(n6589), .A(n6588), .B(n9744), .ZN(n6599)
         );
  INV_X1 U8194 ( .A(n6591), .ZN(n6592) );
  OAI21_X1 U8195 ( .B1(n6594), .B2(n6593), .A(n6592), .ZN(n6597) );
  INV_X1 U8196 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n6595) );
  NAND2_X1 U8197 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(P2_U3152), .ZN(n7308) );
  OAI21_X1 U8198 ( .B1(n8068), .B2(n6595), .A(n7308), .ZN(n6596) );
  AOI21_X1 U8199 ( .B1(n9748), .B2(n6597), .A(n6596), .ZN(n6598) );
  OAI211_X1 U8200 ( .C1(n9680), .C2(n6600), .A(n6599), .B(n6598), .ZN(P2_U3257) );
  NAND2_X1 U8201 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(P2_U3152), .ZN(n6997) );
  INV_X1 U8202 ( .A(n6997), .ZN(n6607) );
  AND3_X1 U8203 ( .A1(n6603), .A2(n6602), .A3(n6601), .ZN(n6604) );
  NOR3_X1 U8204 ( .A1(n9681), .A2(n6605), .A3(n6604), .ZN(n6606) );
  AOI211_X1 U8205 ( .C1(P2_ADDR_REG_9__SCAN_IN), .C2(n9741), .A(n6607), .B(
        n6606), .ZN(n6612) );
  OAI211_X1 U8206 ( .C1(n6610), .C2(n6609), .A(n9744), .B(n6608), .ZN(n6611)
         );
  OAI211_X1 U8207 ( .C1(n9680), .C2(n6613), .A(n6612), .B(n6611), .ZN(P2_U3254) );
  INV_X1 U8208 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n8027) );
  INV_X1 U8209 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n8026) );
  INV_X1 U8210 ( .A(n8029), .ZN(n8398) );
  INV_X1 U8211 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n6617) );
  NAND2_X1 U8212 ( .A1(n5871), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n6616) );
  NAND2_X1 U8213 ( .A1(n4276), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n6615) );
  OAI211_X1 U8214 ( .C1(n8154), .C2(n6617), .A(n6616), .B(n6615), .ZN(n6618)
         );
  AOI21_X1 U8215 ( .B1(n8398), .B2(n8034), .A(n6618), .ZN(n8588) );
  NAND2_X1 U8216 ( .A1(P2_DATAO_REG_29__SCAN_IN), .A2(n8531), .ZN(n6619) );
  OAI21_X1 U8217 ( .B1(n8588), .B2(n8531), .A(n6619), .ZN(P2_U3581) );
  INV_X1 U8218 ( .A(n6620), .ZN(n6650) );
  AOI22_X1 U8219 ( .A1(n9039), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n9369), .ZN(n6621) );
  OAI21_X1 U8220 ( .B1(n6650), .B2(n9371), .A(n6621), .ZN(P1_U3336) );
  NAND4_X1 U8221 ( .A1(n9774), .A2(n7109), .A3(n7112), .A4(n6622), .ZN(n6623)
         );
  OR2_X1 U8222 ( .A1(n6624), .A2(n6623), .ZN(n6814) );
  INV_X1 U8223 ( .A(n7111), .ZN(n6625) );
  INV_X2 U8224 ( .A(n9827), .ZN(n9828) );
  INV_X1 U8225 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n6643) );
  OAI21_X1 U8226 ( .B1(n8373), .B2(n6626), .A(n7951), .ZN(n6627) );
  NAND3_X1 U8227 ( .A1(n6628), .A2(n6627), .A3(n5730), .ZN(n8729) );
  NAND2_X1 U8228 ( .A1(n8342), .A2(n9764), .ZN(n9763) );
  NAND2_X1 U8229 ( .A1(n6629), .A2(n9785), .ZN(n6631) );
  NAND2_X1 U8230 ( .A1(n9763), .A2(n6631), .ZN(n6633) );
  OR2_X1 U8231 ( .A1(n6632), .A2(n6739), .ZN(n8198) );
  NAND2_X1 U8232 ( .A1(n6632), .A2(n6739), .ZN(n8199) );
  NAND2_X1 U8233 ( .A1(n8198), .A2(n8199), .ZN(n6635) );
  NAND2_X1 U8234 ( .A1(n6633), .A2(n6635), .ZN(n6741) );
  OAI21_X1 U8235 ( .B1(n6633), .B2(n6635), .A(n6741), .ZN(n6634) );
  INV_X1 U8236 ( .A(n6634), .ZN(n7206) );
  NAND2_X1 U8237 ( .A1(n8372), .A2(n8166), .ZN(n9759) );
  INV_X1 U8238 ( .A(n6635), .ZN(n6638) );
  NAND2_X1 U8239 ( .A1(n6636), .A2(n9761), .ZN(n9756) );
  NAND2_X1 U8240 ( .A1(n8197), .A2(n9756), .ZN(n8183) );
  NAND2_X1 U8241 ( .A1(n6638), .A2(n6637), .ZN(n6750) );
  OAI21_X1 U8242 ( .B1(n6638), .B2(n6637), .A(n6750), .ZN(n6639) );
  INV_X1 U8243 ( .A(n8721), .ZN(n8755) );
  AOI222_X1 U8244 ( .A1(n9759), .A2(n6639), .B1(n6630), .B2(n8753), .C1(n8530), 
        .C2(n8755), .ZN(n7200) );
  NAND3_X1 U8245 ( .A1(n9785), .A2(n6739), .A3(n6733), .ZN(n6747) );
  INV_X1 U8246 ( .A(n6747), .ZN(n7212) );
  AOI21_X1 U8247 ( .B1(n9785), .B2(n6733), .A(n6739), .ZN(n6640) );
  NOR2_X1 U8248 ( .A1(n7212), .A2(n6640), .ZN(n7201) );
  INV_X1 U8249 ( .A(n6739), .ZN(n7972) );
  AOI22_X1 U8250 ( .A1(n7201), .A2(n5731), .B1(n8849), .B2(n7972), .ZN(n6641)
         );
  OAI211_X1 U8251 ( .C1(n9798), .C2(n7206), .A(n7200), .B(n6641), .ZN(n6815)
         );
  NAND2_X1 U8252 ( .A1(n9828), .A2(n6815), .ZN(n6642) );
  OAI21_X1 U8253 ( .B1(n9828), .B2(n6643), .A(n6642), .ZN(P2_U3457) );
  INV_X1 U8254 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n9943) );
  NAND2_X1 U8255 ( .A1(n6644), .A2(n6733), .ZN(n8177) );
  AND2_X1 U8256 ( .A1(n9756), .A2(n8177), .ZN(n8340) );
  INV_X1 U8257 ( .A(n8340), .ZN(n6645) );
  AOI22_X1 U8258 ( .A1(n6645), .A2(n9759), .B1(n8755), .B2(n6630), .ZN(n7265)
         );
  NAND2_X1 U8259 ( .A1(n9761), .A2(n6646), .ZN(n6647) );
  OAI211_X1 U8260 ( .C1(n8340), .C2(n9798), .A(n7265), .B(n6647), .ZN(n6817)
         );
  NAND2_X1 U8261 ( .A1(n9828), .A2(n6817), .ZN(n6648) );
  OAI21_X1 U8262 ( .B1(n9828), .B2(n9943), .A(n6648), .ZN(P2_U3451) );
  OAI222_X1 U8263 ( .A1(P2_U3152), .A2(n7622), .B1(n4284), .B2(n6650), .C1(
        n6649), .C2(n7969), .ZN(P2_U3341) );
  NAND2_X1 U8264 ( .A1(n6921), .A2(n7933), .ZN(n6652) );
  AOI22_X1 U8265 ( .A1(n9008), .A2(n7904), .B1(n6921), .B2(n7939), .ZN(n6717)
         );
  XNOR2_X1 U8266 ( .A(n6716), .B(n6717), .ZN(n6657) );
  OAI21_X1 U8267 ( .B1(n6657), .B2(n6656), .A(n6720), .ZN(n6665) );
  INV_X1 U8268 ( .A(n8968), .ZN(n8997) );
  NOR2_X1 U8269 ( .A1(n8997), .A2(n9618), .ZN(n6664) );
  NAND2_X1 U8270 ( .A1(n6659), .A2(n6658), .ZN(n6660) );
  INV_X1 U8271 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n6902) );
  NOR2_X1 U8272 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6902), .ZN(n9021) );
  AOI21_X1 U8273 ( .B1(n8965), .B2(n6448), .A(n9021), .ZN(n6662) );
  NAND2_X1 U8274 ( .A1(n8994), .A2(n9585), .ZN(n6661) );
  OAI211_X1 U8275 ( .C1(P1_REG3_REG_3__SCAN_IN), .C2(n8989), .A(n6662), .B(
        n6661), .ZN(n6663) );
  AOI211_X1 U8276 ( .C1(n6665), .C2(n8973), .A(n6664), .B(n6663), .ZN(n6666)
         );
  INV_X1 U8277 ( .A(n6666), .ZN(P1_U3216) );
  INV_X1 U8278 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n6669) );
  AOI22_X1 U8279 ( .A1(P2_REG2_REG_14__SCAN_IN), .A2(n7141), .B1(n7149), .B2(
        n6669), .ZN(n6670) );
  AOI21_X1 U8280 ( .B1(n6671), .B2(n6670), .A(n7150), .ZN(n6681) );
  INV_X1 U8281 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n6672) );
  NAND2_X1 U8282 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(P2_U3152), .ZN(n8048) );
  OAI21_X1 U8283 ( .B1(n8068), .B2(n6672), .A(n8048), .ZN(n6679) );
  AOI21_X1 U8284 ( .B1(n9388), .B2(n6674), .A(n6673), .ZN(n6676) );
  INV_X1 U8285 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n7142) );
  AOI22_X1 U8286 ( .A1(P2_REG1_REG_14__SCAN_IN), .A2(n7141), .B1(n7149), .B2(
        n7142), .ZN(n6675) );
  NOR2_X1 U8287 ( .A1(n6676), .A2(n6675), .ZN(n7140) );
  AOI21_X1 U8288 ( .B1(n6676), .B2(n6675), .A(n7140), .ZN(n6677) );
  NOR2_X1 U8289 ( .A1(n6677), .A2(n9681), .ZN(n6678) );
  AOI211_X1 U8290 ( .C1(n9747), .C2(n7149), .A(n6679), .B(n6678), .ZN(n6680)
         );
  OAI21_X1 U8291 ( .B1(n6681), .B2(n9692), .A(n6680), .ZN(P2_U3259) );
  XNOR2_X1 U8292 ( .A(n6683), .B(n6682), .ZN(n6688) );
  INV_X1 U8293 ( .A(n8219), .ZN(n9807) );
  NOR2_X1 U8294 ( .A1(n8499), .A2(n9807), .ZN(n6686) );
  NAND2_X1 U8295 ( .A1(n8504), .A2(n8527), .ZN(n6684) );
  NAND2_X1 U8296 ( .A1(P2_U3152), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n9713) );
  OAI211_X1 U8297 ( .C1(n7296), .C2(n8502), .A(n6684), .B(n9713), .ZN(n6685)
         );
  AOI211_X1 U8298 ( .C1(n8496), .C2(n7289), .A(n6686), .B(n6685), .ZN(n6687)
         );
  OAI21_X1 U8299 ( .B1(n6688), .B2(n8511), .A(n6687), .ZN(P2_U3215) );
  INV_X1 U8300 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n6702) );
  OAI21_X1 U8301 ( .B1(n6695), .B2(P1_REG1_REG_12__SCAN_IN), .A(n6689), .ZN(
        n6692) );
  AOI22_X1 U8302 ( .A1(n6806), .A2(P1_REG1_REG_13__SCAN_IN), .B1(n5221), .B2(
        n6690), .ZN(n6691) );
  NAND2_X1 U8303 ( .A1(n6691), .A2(n6692), .ZN(n6800) );
  OAI21_X1 U8304 ( .B1(n6692), .B2(n6691), .A(n6800), .ZN(n6693) );
  NAND2_X1 U8305 ( .A1(n6693), .A2(n9566), .ZN(n6701) );
  AND2_X1 U8306 ( .A1(P1_U3084), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n7566) );
  NAND2_X1 U8307 ( .A1(n6806), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n6696) );
  OAI21_X1 U8308 ( .B1(n6806), .B2(P1_REG2_REG_13__SCAN_IN), .A(n6696), .ZN(
        n6697) );
  AOI211_X1 U8309 ( .C1(n6698), .C2(n6697), .A(n6805), .B(n9543), .ZN(n6699)
         );
  AOI211_X1 U8310 ( .C1(n6806), .C2(n9553), .A(n7566), .B(n6699), .ZN(n6700)
         );
  OAI211_X1 U8311 ( .C1(n9571), .C2(n6702), .A(n6701), .B(n6700), .ZN(P1_U3254) );
  AOI21_X1 U8312 ( .B1(n6705), .B2(n6704), .A(n6703), .ZN(n6715) );
  NOR2_X1 U8313 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7273), .ZN(n6706) );
  AOI21_X1 U8314 ( .B1(n9741), .B2(P2_ADDR_REG_11__SCAN_IN), .A(n6706), .ZN(
        n6711) );
  OAI211_X1 U8315 ( .C1(n6709), .C2(n6708), .A(n9748), .B(n6707), .ZN(n6710)
         );
  OAI211_X1 U8316 ( .C1(n9680), .C2(n6712), .A(n6711), .B(n6710), .ZN(n6713)
         );
  INV_X1 U8317 ( .A(n6713), .ZN(n6714) );
  OAI21_X1 U8318 ( .B1(n6715), .B2(n9692), .A(n6714), .ZN(P2_U3256) );
  INV_X1 U8319 ( .A(n6716), .ZN(n6718) );
  NAND2_X1 U8320 ( .A1(n6718), .A2(n6717), .ZN(n6719) );
  NAND2_X1 U8321 ( .A1(n9585), .A2(n7939), .ZN(n6722) );
  NAND2_X1 U8322 ( .A1(n6945), .A2(n7933), .ZN(n6721) );
  NAND2_X1 U8323 ( .A1(n6722), .A2(n6721), .ZN(n6723) );
  XNOR2_X1 U8324 ( .A(n6723), .B(n7936), .ZN(n6725) );
  AOI22_X1 U8325 ( .A1(n9585), .A2(n7904), .B1(n6945), .B2(n7939), .ZN(n6724)
         );
  OR2_X1 U8326 ( .A1(n6725), .A2(n6724), .ZN(n6864) );
  NAND2_X1 U8327 ( .A1(n4345), .A2(n6864), .ZN(n6726) );
  XNOR2_X1 U8328 ( .A(n6865), .B(n6726), .ZN(n6731) );
  AND2_X1 U8329 ( .A1(P1_U3084), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n9491) );
  AOI21_X1 U8330 ( .B1(n8965), .B2(n9008), .A(n9491), .ZN(n6728) );
  NAND2_X1 U8331 ( .A1(n8994), .A2(n9007), .ZN(n6727) );
  OAI211_X1 U8332 ( .C1(n8989), .C2(n6920), .A(n6728), .B(n6727), .ZN(n6729)
         );
  AOI21_X1 U8333 ( .B1(n8968), .B2(n6945), .A(n6729), .ZN(n6730) );
  OAI21_X1 U8334 ( .B1(n6731), .B2(n8984), .A(n6730), .ZN(P1_U3228) );
  INV_X1 U8335 ( .A(n6732), .ZN(n6738) );
  INV_X1 U8336 ( .A(n8484), .ZN(n8472) );
  AOI22_X1 U8337 ( .A1(n8472), .A2(n6644), .B1(n9761), .B2(n8473), .ZN(n6737)
         );
  INV_X1 U8338 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n7266) );
  NOR2_X1 U8339 ( .A1(n7266), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9679) );
  OAI22_X1 U8340 ( .A1(n8499), .A2(n6733), .B1(n8502), .B2(n6629), .ZN(n6734)
         );
  AOI211_X1 U8341 ( .C1(P2_REG3_REG_0__SCAN_IN), .C2(n6735), .A(n9679), .B(
        n6734), .ZN(n6736) );
  OAI21_X1 U8342 ( .B1(n6738), .B2(n6737), .A(n6736), .ZN(P2_U3234) );
  NAND2_X1 U8343 ( .A1(n8530), .A2(n9792), .ZN(n8208) );
  NAND2_X1 U8344 ( .A1(n8189), .A2(n8208), .ZN(n7208) );
  NAND2_X1 U8345 ( .A1(n7219), .A2(n6739), .ZN(n6740) );
  NAND2_X1 U8346 ( .A1(n6741), .A2(n6740), .ZN(n7209) );
  INV_X1 U8347 ( .A(n8530), .ZN(n6742) );
  NAND2_X1 U8348 ( .A1(n6742), .A2(n9792), .ZN(n6743) );
  NAND2_X1 U8349 ( .A1(n7207), .A2(n6743), .ZN(n6767) );
  OR2_X1 U8350 ( .A1(n8529), .A2(n7124), .ZN(n8191) );
  NAND2_X1 U8351 ( .A1(n8529), .A2(n7124), .ZN(n8209) );
  NAND2_X1 U8352 ( .A1(n8191), .A2(n8209), .ZN(n8343) );
  NAND2_X1 U8353 ( .A1(n6767), .A2(n8343), .ZN(n6766) );
  NAND2_X1 U8354 ( .A1(n7218), .A2(n7124), .ZN(n6744) );
  NAND2_X1 U8355 ( .A1(n6766), .A2(n6744), .ZN(n7029) );
  NOR2_X1 U8356 ( .A1(n8528), .A2(n7238), .ZN(n7031) );
  OR2_X1 U8357 ( .A1(n7029), .A2(n7031), .ZN(n6745) );
  INV_X1 U8358 ( .A(n8528), .ZN(n6852) );
  NAND2_X1 U8359 ( .A1(n6745), .A2(n7037), .ZN(n6746) );
  OR2_X1 U8360 ( .A1(n8527), .A2(n7965), .ZN(n8215) );
  NAND2_X1 U8361 ( .A1(n8527), .A2(n7965), .ZN(n8211) );
  NAND2_X1 U8362 ( .A1(n8215), .A2(n8211), .ZN(n7045) );
  XNOR2_X1 U8363 ( .A(n6746), .B(n7046), .ZN(n7320) );
  INV_X1 U8364 ( .A(n9798), .ZN(n9825) );
  AND2_X1 U8365 ( .A1(n6770), .A2(n7124), .ZN(n7232) );
  NAND2_X1 U8366 ( .A1(n7232), .A2(n6748), .ZN(n7231) );
  INV_X1 U8367 ( .A(n7965), .ZN(n7314) );
  NAND2_X1 U8368 ( .A1(n7231), .A2(n7314), .ZN(n6749) );
  NAND2_X1 U8369 ( .A1(n7286), .A2(n6749), .ZN(n7316) );
  INV_X1 U8370 ( .A(n8849), .ZN(n9819) );
  OAI22_X1 U8371 ( .A1(n7316), .A2(n4275), .B1(n7965), .B2(n9819), .ZN(n6752)
         );
  NAND2_X1 U8372 ( .A1(n6750), .A2(n8198), .ZN(n7217) );
  XNOR2_X1 U8373 ( .A(n7044), .B(n7046), .ZN(n6751) );
  INV_X1 U8374 ( .A(n9759), .ZN(n8698) );
  AOI22_X1 U8375 ( .A1(n8753), .A2(n8528), .B1(n8526), .B2(n8755), .ZN(n7959)
         );
  OAI21_X1 U8376 ( .B1(n6751), .B2(n8698), .A(n7959), .ZN(n7317) );
  AOI211_X1 U8377 ( .C1(n7320), .C2(n9825), .A(n6752), .B(n7317), .ZN(n6820)
         );
  NAND2_X1 U8378 ( .A1(n9827), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n6753) );
  OAI21_X1 U8379 ( .B1(n6820), .B2(n9827), .A(n6753), .ZN(P2_U3469) );
  INV_X1 U8380 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n6765) );
  INV_X1 U8381 ( .A(n6754), .ZN(n9366) );
  NAND2_X1 U8382 ( .A1(n9366), .A2(n9271), .ZN(n6756) );
  OR2_X1 U8383 ( .A1(n6756), .A2(n6755), .ZN(n6984) );
  NAND3_X1 U8384 ( .A1(n9602), .A2(n9572), .A3(n9592), .ZN(n9418) );
  NAND2_X2 U8385 ( .A1(n6984), .A2(n9418), .ZN(n9600) );
  OAI21_X1 U8386 ( .B1(n6758), .B2(n9418), .A(n6757), .ZN(n6759) );
  NAND2_X1 U8387 ( .A1(n6759), .A2(n9600), .ZN(n6764) );
  NAND2_X1 U8388 ( .A1(n9600), .A2(n9590), .ZN(n9256) );
  NOR2_X1 U8389 ( .A1(n6761), .A2(n6760), .ZN(n6762) );
  OAI21_X1 U8390 ( .B1(n9434), .B2(n9417), .A(n6778), .ZN(n6763) );
  OAI211_X1 U8391 ( .C1(n6765), .C2(n9600), .A(n6764), .B(n6763), .ZN(P1_U3291) );
  INV_X1 U8392 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n6775) );
  OAI21_X1 U8393 ( .B1(n6767), .B2(n8343), .A(n6766), .ZN(n7126) );
  INV_X1 U8394 ( .A(n7126), .ZN(n6773) );
  XOR2_X1 U8395 ( .A(n6768), .B(n8343), .Z(n6769) );
  AOI222_X1 U8396 ( .A1(n9759), .A2(n6769), .B1(n8528), .B2(n8755), .C1(n8530), 
        .C2(n8753), .ZN(n7128) );
  INV_X1 U8397 ( .A(n7124), .ZN(n6771) );
  INV_X1 U8398 ( .A(n6770), .ZN(n7211) );
  AOI211_X1 U8399 ( .C1(n6771), .C2(n7211), .A(n4275), .B(n7232), .ZN(n7122)
         );
  AOI21_X1 U8400 ( .B1(n8849), .B2(n6771), .A(n7122), .ZN(n6772) );
  OAI211_X1 U8401 ( .C1(n9798), .C2(n6773), .A(n7128), .B(n6772), .ZN(n6822)
         );
  NAND2_X1 U8402 ( .A1(n6822), .A2(n9828), .ZN(n6774) );
  OAI21_X1 U8403 ( .B1(n9828), .B2(n6775), .A(n6774), .ZN(P2_U3463) );
  INV_X1 U8404 ( .A(n6776), .ZN(n6832) );
  AOI22_X1 U8405 ( .A1(n9055), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n9369), .ZN(n6777) );
  OAI21_X1 U8406 ( .B1(n6832), .B2(n9371), .A(n6777), .ZN(P1_U3335) );
  NAND2_X1 U8407 ( .A1(n6360), .A2(n6778), .ZN(n6894) );
  XNOR2_X1 U8408 ( .A(n6782), .B(n6894), .ZN(n9609) );
  NOR2_X1 U8409 ( .A1(n7936), .A2(n4344), .ZN(n6779) );
  NAND2_X1 U8410 ( .A1(n9600), .A2(n6779), .ZN(n9268) );
  OAI21_X1 U8411 ( .B1(n6782), .B2(n6781), .A(n6780), .ZN(n6791) );
  OR2_X1 U8412 ( .A1(n6976), .A2(n5664), .ZN(n6783) );
  INV_X1 U8413 ( .A(n6785), .ZN(n6787) );
  INV_X1 U8414 ( .A(n9586), .ZN(n9423) );
  OAI22_X1 U8415 ( .A1(n6789), .A2(n9423), .B1(n6788), .B2(n9576), .ZN(n6790)
         );
  AOI21_X1 U8416 ( .B1(n6791), .B2(n9427), .A(n6790), .ZN(n6792) );
  OAI21_X1 U8417 ( .B1(n9609), .B2(n9279), .A(n6792), .ZN(n9611) );
  INV_X1 U8418 ( .A(n6936), .ZN(n6793) );
  OAI211_X1 U8419 ( .C1(n6795), .C2(n6794), .A(n6793), .B(n9572), .ZN(n9607)
         );
  OAI22_X1 U8420 ( .A1(n9607), .A2(n9592), .B1(n9418), .B2(n6796), .ZN(n6797)
         );
  OAI21_X1 U8421 ( .B1(n9611), .B2(n6797), .A(n9600), .ZN(n6799) );
  AOI22_X1 U8422 ( .A1(n9434), .A2(n6896), .B1(n4283), .B2(
        P1_REG2_REG_1__SCAN_IN), .ZN(n6798) );
  OAI211_X1 U8423 ( .C1(n9609), .C2(n9268), .A(n6799), .B(n6798), .ZN(P1_U3290) );
  INV_X1 U8424 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n6813) );
  OAI21_X1 U8425 ( .B1(P1_REG1_REG_13__SCAN_IN), .B2(n6806), .A(n6800), .ZN(
        n6803) );
  NOR2_X1 U8426 ( .A1(n7258), .A2(n7257), .ZN(n6801) );
  AOI21_X1 U8427 ( .B1(n7257), .B2(n7258), .A(n6801), .ZN(n6802) );
  NAND2_X1 U8428 ( .A1(n6802), .A2(n6803), .ZN(n7255) );
  OAI21_X1 U8429 ( .B1(n6803), .B2(n6802), .A(n7255), .ZN(n6804) );
  NAND2_X1 U8430 ( .A1(n6804), .A2(n9566), .ZN(n6812) );
  INV_X1 U8431 ( .A(n9543), .ZN(n9556) );
  AOI21_X1 U8432 ( .B1(P1_REG2_REG_13__SCAN_IN), .B2(n6806), .A(n6805), .ZN(
        n7250) );
  XNOR2_X1 U8433 ( .A(n6807), .B(n7250), .ZN(n6808) );
  NAND2_X1 U8434 ( .A1(n6808), .A2(n7698), .ZN(n7251) );
  OAI21_X1 U8435 ( .B1(n6808), .B2(n7698), .A(n7251), .ZN(n6810) );
  NAND2_X1 U8436 ( .A1(P1_REG3_REG_14__SCAN_IN), .A2(P1_U3084), .ZN(n7714) );
  OAI21_X1 U8437 ( .B1(n9538), .B2(n7258), .A(n7714), .ZN(n6809) );
  AOI21_X1 U8438 ( .B1(n9556), .B2(n6810), .A(n6809), .ZN(n6811) );
  OAI211_X1 U8439 ( .C1(n9571), .C2(n6813), .A(n6812), .B(n6811), .ZN(P1_U3255) );
  NOR2_X2 U8440 ( .A1(n6814), .A2(n7111), .ZN(n9840) );
  NAND2_X1 U8441 ( .A1(n9836), .A2(n6815), .ZN(n6816) );
  OAI21_X1 U8442 ( .B1(n9836), .B2(n6480), .A(n6816), .ZN(P2_U3522) );
  INV_X1 U8443 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n6819) );
  NAND2_X1 U8444 ( .A1(n9836), .A2(n6817), .ZN(n6818) );
  OAI21_X1 U8445 ( .B1(n9836), .B2(n6819), .A(n6818), .ZN(P2_U3520) );
  OR2_X1 U8446 ( .A1(n6820), .A2(n9837), .ZN(n6821) );
  OAI21_X1 U8447 ( .B1(n9836), .B2(n6511), .A(n6821), .ZN(P2_U3526) );
  NAND2_X1 U8448 ( .A1(n6822), .A2(n9836), .ZN(n6823) );
  OAI21_X1 U8449 ( .B1(n9836), .B2(n6485), .A(n6823), .ZN(P2_U3524) );
  XNOR2_X1 U8450 ( .A(n6825), .B(n6824), .ZN(n6831) );
  INV_X1 U8451 ( .A(n7062), .ZN(n7243) );
  NOR2_X1 U8452 ( .A1(n8499), .A2(n7243), .ZN(n6829) );
  NAND2_X1 U8453 ( .A1(n8504), .A2(n8526), .ZN(n6827) );
  OAI211_X1 U8454 ( .C1(n7078), .C2(n8502), .A(n6827), .B(n6826), .ZN(n6828)
         );
  AOI211_X1 U8455 ( .C1(n8496), .C2(n7241), .A(n6829), .B(n6828), .ZN(n6830)
         );
  OAI21_X1 U8456 ( .B1(n6831), .B2(n8511), .A(n6830), .ZN(P2_U3223) );
  INV_X1 U8457 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n6833) );
  INV_X1 U8458 ( .A(n7629), .ZN(n7615) );
  OAI222_X1 U8459 ( .A1(n7969), .A2(n6833), .B1(n4284), .B2(n6832), .C1(
        P2_U3152), .C2(n7615), .ZN(P2_U3340) );
  OAI21_X1 U8460 ( .B1(n6837), .B2(n6205), .A(n6846), .ZN(n6842) );
  OAI21_X1 U8461 ( .B1(n8499), .B2(n7124), .A(n6834), .ZN(n6835) );
  AOI21_X1 U8462 ( .B1(n8491), .B2(n8528), .A(n6835), .ZN(n6840) );
  NOR3_X1 U8463 ( .A1(n8484), .A2(n6837), .A3(n6836), .ZN(n6838) );
  OAI21_X1 U8464 ( .B1(n6838), .B2(n8504), .A(n8530), .ZN(n6839) );
  OAI211_X1 U8465 ( .C1(n8506), .C2(n7120), .A(n6840), .B(n6839), .ZN(n6841)
         );
  AOI21_X1 U8466 ( .B1(n8473), .B2(n6842), .A(n6841), .ZN(n6843) );
  INV_X1 U8467 ( .A(n6843), .ZN(P2_U3232) );
  NAND2_X1 U8468 ( .A1(n6844), .A2(n6848), .ZN(n6847) );
  NAND2_X1 U8469 ( .A1(n6846), .A2(n6845), .ZN(n6853) );
  MUX2_X1 U8470 ( .A(n6848), .B(n6847), .S(n6853), .Z(n6857) );
  AOI22_X1 U8471 ( .A1(n8491), .A2(n8527), .B1(n8504), .B2(n8529), .ZN(n6850)
         );
  OAI211_X1 U8472 ( .C1(n6748), .C2(n8499), .A(n6850), .B(n6849), .ZN(n6855)
         );
  NOR4_X1 U8473 ( .A1(n6853), .A2(n6852), .A3(n6851), .A4(n8484), .ZN(n6854)
         );
  AOI211_X1 U8474 ( .C1(n8496), .C2(n7234), .A(n6855), .B(n6854), .ZN(n6856)
         );
  OAI21_X1 U8475 ( .B1(n6857), .B2(n8511), .A(n6856), .ZN(P2_U3229) );
  NAND2_X1 U8476 ( .A1(n9006), .A2(n7939), .ZN(n6859) );
  OR2_X1 U8477 ( .A1(n9646), .A2(n6384), .ZN(n6858) );
  NAND2_X1 U8478 ( .A1(n6859), .A2(n6858), .ZN(n6861) );
  XNOR2_X1 U8479 ( .A(n6861), .B(n6860), .ZN(n7166) );
  NAND2_X1 U8480 ( .A1(n9006), .A2(n7904), .ZN(n6863) );
  OR2_X1 U8481 ( .A1(n9646), .A2(n6359), .ZN(n6862) );
  NAND2_X1 U8482 ( .A1(n6863), .A2(n6862), .ZN(n7167) );
  XNOR2_X1 U8483 ( .A(n7166), .B(n7167), .ZN(n7171) );
  NAND2_X1 U8484 ( .A1(n9007), .A2(n7939), .ZN(n6867) );
  INV_X1 U8485 ( .A(n9633), .ZN(n9589) );
  NAND2_X1 U8486 ( .A1(n9589), .A2(n7933), .ZN(n6866) );
  NAND2_X1 U8487 ( .A1(n6867), .A2(n6866), .ZN(n6868) );
  XNOR2_X1 U8488 ( .A(n6868), .B(n7936), .ZN(n6962) );
  NAND2_X1 U8489 ( .A1(n9007), .A2(n7904), .ZN(n6870) );
  NAND2_X1 U8490 ( .A1(n9589), .A2(n7939), .ZN(n6869) );
  AND2_X1 U8491 ( .A1(n6870), .A2(n6869), .ZN(n6964) );
  NAND2_X1 U8492 ( .A1(n9575), .A2(n7939), .ZN(n6872) );
  NAND2_X1 U8493 ( .A1(n7026), .A2(n7933), .ZN(n6871) );
  NAND2_X1 U8494 ( .A1(n6872), .A2(n6871), .ZN(n6873) );
  XNOR2_X1 U8495 ( .A(n6873), .B(n7936), .ZN(n7019) );
  NAND2_X1 U8496 ( .A1(n9575), .A2(n7904), .ZN(n6875) );
  NAND2_X1 U8497 ( .A1(n7026), .A2(n7939), .ZN(n6874) );
  AND2_X1 U8498 ( .A1(n6875), .A2(n6874), .ZN(n7018) );
  AOI22_X1 U8499 ( .A1(n6962), .A2(n6964), .B1(n7019), .B2(n7018), .ZN(n6876)
         );
  NAND2_X1 U8500 ( .A1(n6961), .A2(n6876), .ZN(n6883) );
  OAI21_X1 U8501 ( .B1(n6962), .B2(n6964), .A(n7018), .ZN(n6881) );
  INV_X1 U8502 ( .A(n7019), .ZN(n6880) );
  INV_X1 U8503 ( .A(n6964), .ZN(n6878) );
  INV_X1 U8504 ( .A(n7018), .ZN(n6877) );
  AND2_X1 U8505 ( .A1(n6878), .A2(n6877), .ZN(n6879) );
  INV_X1 U8506 ( .A(n6962), .ZN(n7017) );
  AOI22_X1 U8507 ( .A1(n6881), .A2(n6880), .B1(n6879), .B2(n7017), .ZN(n6882)
         );
  NAND2_X1 U8508 ( .A1(n6883), .A2(n6882), .ZN(n7172) );
  XOR2_X1 U8509 ( .A(n7171), .B(n7172), .Z(n6889) );
  AOI21_X1 U8510 ( .B1(n8994), .B2(n9005), .A(n6884), .ZN(n6886) );
  NAND2_X1 U8511 ( .A1(n8965), .A2(n9575), .ZN(n6885) );
  OAI211_X1 U8512 ( .C1(n8989), .C2(n6985), .A(n6886), .B(n6885), .ZN(n6887)
         );
  AOI21_X1 U8513 ( .B1(n8968), .B2(n7091), .A(n6887), .ZN(n6888) );
  OAI21_X1 U8514 ( .B1(n6889), .B2(n8984), .A(n6888), .ZN(P1_U3211) );
  INV_X1 U8515 ( .A(n6890), .ZN(n6892) );
  OAI222_X1 U8516 ( .A1(n7969), .A2(n6891), .B1(n4284), .B2(n6892), .C1(
        P2_U3152), .C2(n5730), .ZN(P2_U3339) );
  OAI222_X1 U8517 ( .A1(n8069), .A2(n6893), .B1(n9371), .B2(n6892), .C1(
        P1_U3084), .C2(n9141), .ZN(P1_U3334) );
  INV_X1 U8518 ( .A(n9268), .ZN(n9597) );
  NAND2_X1 U8519 ( .A1(n6895), .A2(n6894), .ZN(n6899) );
  OR2_X1 U8520 ( .A1(n6897), .A2(n6896), .ZN(n6898) );
  NAND2_X1 U8521 ( .A1(n6899), .A2(n6898), .ZN(n6931) );
  NAND2_X1 U8522 ( .A1(n6931), .A2(n6930), .ZN(n6901) );
  OR2_X1 U8523 ( .A1(n6448), .A2(n6937), .ZN(n6900) );
  NAND2_X1 U8524 ( .A1(n6901), .A2(n6900), .ZN(n6912) );
  XNOR2_X1 U8525 ( .A(n6912), .B(n6911), .ZN(n9621) );
  INV_X1 U8526 ( .A(n9417), .ZN(n7807) );
  NAND2_X1 U8527 ( .A1(n6936), .A2(n9612), .ZN(n6935) );
  XNOR2_X1 U8528 ( .A(n6935), .B(n6921), .ZN(n9619) );
  INV_X1 U8529 ( .A(n9418), .ZN(n9588) );
  AOI22_X1 U8530 ( .A1(n9434), .A2(n6921), .B1(n6902), .B2(n9588), .ZN(n6903)
         );
  OAI21_X1 U8531 ( .B1(n7807), .B2(n9619), .A(n6903), .ZN(n6909) );
  XNOR2_X1 U8532 ( .A(n6904), .B(n6911), .ZN(n6905) );
  NAND2_X1 U8533 ( .A1(n6905), .A2(n9427), .ZN(n6907) );
  AOI22_X1 U8534 ( .A1(n9261), .A2(n9585), .B1(n6448), .B2(n9586), .ZN(n6906)
         );
  NAND2_X1 U8535 ( .A1(n6907), .A2(n6906), .ZN(n9617) );
  MUX2_X1 U8536 ( .A(n9617), .B(P1_REG2_REG_3__SCAN_IN), .S(n4283), .Z(n6908)
         );
  AOI211_X1 U8537 ( .C1(n9597), .C2(n9621), .A(n6909), .B(n6908), .ZN(n6910)
         );
  INV_X1 U8538 ( .A(n6910), .ZN(P1_U3288) );
  NAND2_X1 U8539 ( .A1(n6912), .A2(n6911), .ZN(n6914) );
  OR2_X1 U8540 ( .A1(n9008), .A2(n6921), .ZN(n6913) );
  INV_X1 U8541 ( .A(n6943), .ZN(n6915) );
  XNOR2_X1 U8542 ( .A(n6944), .B(n6915), .ZN(n9625) );
  XNOR2_X1 U8543 ( .A(n6916), .B(n6915), .ZN(n6917) );
  NAND2_X1 U8544 ( .A1(n6917), .A2(n9427), .ZN(n6919) );
  AOI22_X1 U8545 ( .A1(n9261), .A2(n9007), .B1(n9008), .B2(n9586), .ZN(n6918)
         );
  OAI211_X1 U8546 ( .C1(n9625), .C2(n9279), .A(n6919), .B(n6918), .ZN(n9631)
         );
  NAND2_X1 U8547 ( .A1(n9631), .A2(n9600), .ZN(n6928) );
  OAI22_X1 U8548 ( .A1(n9600), .A2(n6269), .B1(n6920), .B2(n9418), .ZN(n6926)
         );
  OAI21_X1 U8549 ( .B1(n6935), .B2(n6921), .A(n6945), .ZN(n6922) );
  INV_X1 U8550 ( .A(n6922), .ZN(n6924) );
  NAND2_X1 U8551 ( .A1(n9618), .A2(n9627), .ZN(n6923) );
  NOR2_X1 U8552 ( .A1(n6935), .A2(n6923), .ZN(n9574) );
  OR2_X1 U8553 ( .A1(n6924), .A2(n9574), .ZN(n9628) );
  NOR2_X1 U8554 ( .A1(n9628), .A2(n7807), .ZN(n6925) );
  AOI211_X1 U8555 ( .C1(n9434), .C2(n6945), .A(n6926), .B(n6925), .ZN(n6927)
         );
  OAI211_X1 U8556 ( .C1(n9625), .C2(n9268), .A(n6928), .B(n6927), .ZN(P1_U3287) );
  XNOR2_X1 U8557 ( .A(n6929), .B(n6930), .ZN(n6934) );
  INV_X1 U8558 ( .A(n9427), .ZN(n9581) );
  XNOR2_X1 U8559 ( .A(n6931), .B(n6930), .ZN(n9616) );
  INV_X1 U8560 ( .A(n9279), .ZN(n9420) );
  NAND2_X1 U8561 ( .A1(n9616), .A2(n9420), .ZN(n6933) );
  AOI22_X1 U8562 ( .A1(n9586), .A2(n6897), .B1(n9008), .B2(n9261), .ZN(n6932)
         );
  OAI211_X1 U8563 ( .C1(n6934), .C2(n9581), .A(n6933), .B(n6932), .ZN(n9614)
         );
  INV_X1 U8564 ( .A(n9614), .ZN(n6942) );
  OAI21_X1 U8565 ( .B1(n6936), .B2(n9612), .A(n6935), .ZN(n9613) );
  AOI22_X1 U8566 ( .A1(n4283), .A2(P1_REG2_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(n9588), .ZN(n6939) );
  NAND2_X1 U8567 ( .A1(n9434), .A2(n6937), .ZN(n6938) );
  OAI211_X1 U8568 ( .C1(n7807), .C2(n9613), .A(n6939), .B(n6938), .ZN(n6940)
         );
  AOI21_X1 U8569 ( .B1(n9616), .B2(n9597), .A(n6940), .ZN(n6941) );
  OAI21_X1 U8570 ( .B1(n6942), .B2(n4283), .A(n6941), .ZN(P1_U3289) );
  OR2_X1 U8571 ( .A1(n9585), .A2(n6945), .ZN(n6946) );
  NAND2_X1 U8572 ( .A1(n6947), .A2(n5078), .ZN(n9593) );
  NAND2_X1 U8573 ( .A1(n9007), .A2(n9589), .ZN(n6948) );
  INV_X1 U8574 ( .A(n7412), .ZN(n6949) );
  AOI21_X1 U8575 ( .B1(n6952), .B2(n6950), .A(n6949), .ZN(n9638) );
  AOI22_X1 U8576 ( .A1(n9586), .A2(n9007), .B1(n9006), .B2(n9261), .ZN(n6955)
         );
  XOR2_X1 U8577 ( .A(n6952), .B(n6951), .Z(n6953) );
  NAND2_X1 U8578 ( .A1(n6953), .A2(n9427), .ZN(n6954) );
  OAI211_X1 U8579 ( .C1(n9638), .C2(n9279), .A(n6955), .B(n6954), .ZN(n9641)
         );
  NAND2_X1 U8580 ( .A1(n9641), .A2(n9600), .ZN(n6960) );
  OAI22_X1 U8581 ( .A1(n9600), .A2(n6274), .B1(n7024), .B2(n9418), .ZN(n6958)
         );
  NAND2_X1 U8582 ( .A1(n9574), .A2(n9633), .ZN(n9573) );
  NAND2_X1 U8583 ( .A1(n9573), .A2(n7026), .ZN(n6956) );
  NAND2_X1 U8584 ( .A1(n6981), .A2(n6956), .ZN(n9640) );
  NOR2_X1 U8585 ( .A1(n9640), .A2(n7807), .ZN(n6957) );
  AOI211_X1 U8586 ( .C1(n9434), .C2(n7026), .A(n6958), .B(n6957), .ZN(n6959)
         );
  OAI211_X1 U8587 ( .C1(n9638), .C2(n9268), .A(n6960), .B(n6959), .ZN(P1_U3285) );
  XNOR2_X1 U8588 ( .A(n6961), .B(n6962), .ZN(n6963) );
  NAND2_X1 U8589 ( .A1(n6963), .A2(n6964), .ZN(n7016) );
  OAI21_X1 U8590 ( .B1(n6964), .B2(n6963), .A(n7016), .ZN(n6970) );
  NOR2_X1 U8591 ( .A1(n8997), .A2(n9633), .ZN(n6969) );
  INV_X1 U8592 ( .A(n9587), .ZN(n6967) );
  AND2_X1 U8593 ( .A1(P1_U3084), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n9499) );
  AOI21_X1 U8594 ( .B1(n8965), .B2(n9585), .A(n9499), .ZN(n6966) );
  NAND2_X1 U8595 ( .A1(n8994), .A2(n9575), .ZN(n6965) );
  OAI211_X1 U8596 ( .C1(n8989), .C2(n6967), .A(n6966), .B(n6965), .ZN(n6968)
         );
  AOI211_X1 U8597 ( .C1(n6970), .C2(n8973), .A(n6969), .B(n6968), .ZN(n6971)
         );
  INV_X1 U8598 ( .A(n6971), .ZN(P1_U3225) );
  INV_X1 U8599 ( .A(n6972), .ZN(n6990) );
  OAI222_X1 U8600 ( .A1(n9371), .A2(n6990), .B1(n5664), .B2(P1_U3084), .C1(
        n6973), .C2(n8069), .ZN(P1_U3333) );
  INV_X1 U8601 ( .A(n6974), .ZN(n6991) );
  OAI222_X1 U8602 ( .A1(n8073), .A2(n6991), .B1(n6976), .B2(P1_U3084), .C1(
        n6975), .C2(n8069), .ZN(P1_U3332) );
  NAND2_X1 U8603 ( .A1(n6978), .A2(n6977), .ZN(n6979) );
  XNOR2_X1 U8604 ( .A(n6979), .B(n7415), .ZN(n6980) );
  AOI222_X1 U8605 ( .A1(n9427), .A2(n6980), .B1(n9005), .B2(n9261), .C1(n9575), 
        .C2(n9586), .ZN(n9645) );
  OR2_X1 U8606 ( .A1(n9575), .A2(n7026), .ZN(n7410) );
  NAND2_X1 U8607 ( .A1(n7412), .A2(n7410), .ZN(n7090) );
  XNOR2_X1 U8608 ( .A(n7090), .B(n7415), .ZN(n9648) );
  AOI21_X1 U8609 ( .B1(n6981), .B2(n7091), .A(n9660), .ZN(n6983) );
  NAND2_X1 U8610 ( .A1(n6983), .A2(n7102), .ZN(n9644) );
  NOR2_X1 U8611 ( .A1(n6984), .A2(n9592), .ZN(n9266) );
  INV_X1 U8612 ( .A(n9266), .ZN(n7700) );
  OAI22_X1 U8613 ( .A1(n9600), .A2(n5094), .B1(n6985), .B2(n9418), .ZN(n6986)
         );
  AOI21_X1 U8614 ( .B1(n9434), .B2(n7091), .A(n6986), .ZN(n6987) );
  OAI21_X1 U8615 ( .B1(n9644), .B2(n7700), .A(n6987), .ZN(n6988) );
  AOI21_X1 U8616 ( .B1(n9648), .B2(n9597), .A(n6988), .ZN(n6989) );
  OAI21_X1 U8617 ( .B1(n9645), .B2(n4283), .A(n6989), .ZN(P1_U3284) );
  OAI222_X1 U8618 ( .A1(n7969), .A2(n9997), .B1(n4284), .B2(n6990), .C1(n7116), 
        .C2(P2_U3152), .ZN(P2_U3338) );
  OAI222_X1 U8619 ( .A1(n7969), .A2(n6992), .B1(n4284), .B2(n6991), .C1(n6626), 
        .C2(P2_U3152), .ZN(P2_U3337) );
  INV_X1 U8620 ( .A(n6993), .ZN(n6994) );
  AOI21_X1 U8621 ( .B1(n6996), .B2(n6995), .A(n6994), .ZN(n7002) );
  INV_X1 U8622 ( .A(n7366), .ZN(n9811) );
  NOR2_X1 U8623 ( .A1(n8499), .A2(n9811), .ZN(n7000) );
  INV_X1 U8624 ( .A(n7296), .ZN(n8525) );
  NAND2_X1 U8625 ( .A1(n8504), .A2(n8525), .ZN(n6998) );
  OAI211_X1 U8626 ( .C1(n7376), .C2(n8502), .A(n6998), .B(n6997), .ZN(n6999)
         );
  AOI211_X1 U8627 ( .C1(n8496), .C2(n7365), .A(n7000), .B(n6999), .ZN(n7001)
         );
  OAI21_X1 U8628 ( .B1(n7002), .B2(n8511), .A(n7001), .ZN(P2_U3233) );
  INV_X1 U8629 ( .A(n7003), .ZN(n7953) );
  OAI222_X1 U8630 ( .A1(n8069), .A2(n7005), .B1(n9371), .B2(n7953), .C1(
        P1_U3084), .C2(n7004), .ZN(P1_U3331) );
  XNOR2_X1 U8631 ( .A(n7006), .B(n7007), .ZN(n7012) );
  INV_X1 U8632 ( .A(n7078), .ZN(n8524) );
  NAND2_X1 U8633 ( .A1(n8504), .A2(n8524), .ZN(n7008) );
  NAND2_X1 U8634 ( .A1(P2_U3152), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n9726) );
  OAI211_X1 U8635 ( .C1(n7442), .C2(n8502), .A(n7008), .B(n9726), .ZN(n7010)
         );
  INV_X1 U8636 ( .A(n7322), .ZN(n7134) );
  NOR2_X1 U8637 ( .A1(n7134), .A2(n8499), .ZN(n7009) );
  AOI211_X1 U8638 ( .C1(n8496), .C2(n7132), .A(n7010), .B(n7009), .ZN(n7011)
         );
  OAI21_X1 U8639 ( .B1(n7012), .B2(n8511), .A(n7011), .ZN(P2_U3219) );
  INV_X1 U8640 ( .A(n7060), .ZN(n7015) );
  AOI21_X1 U8641 ( .B1(P2_DATAO_REG_23__SCAN_IN), .B2(n9369), .A(n7013), .ZN(
        n7014) );
  OAI21_X1 U8642 ( .B1(n7015), .B2(n8073), .A(n7014), .ZN(P1_U3330) );
  OAI21_X1 U8643 ( .B1(n6961), .B2(n7017), .A(n7016), .ZN(n7021) );
  XNOR2_X1 U8644 ( .A(n7019), .B(n7018), .ZN(n7020) );
  XNOR2_X1 U8645 ( .A(n7021), .B(n7020), .ZN(n7028) );
  INV_X1 U8646 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n9933) );
  NOR2_X1 U8647 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n9933), .ZN(n9509) );
  AOI21_X1 U8648 ( .B1(n8965), .B2(n9007), .A(n9509), .ZN(n7023) );
  NAND2_X1 U8649 ( .A1(n8994), .A2(n9006), .ZN(n7022) );
  OAI211_X1 U8650 ( .C1(n8989), .C2(n7024), .A(n7023), .B(n7022), .ZN(n7025)
         );
  AOI21_X1 U8651 ( .B1(n8968), .B2(n7026), .A(n7025), .ZN(n7027) );
  OAI21_X1 U8652 ( .B1(n7028), .B2(n8984), .A(n7027), .ZN(P1_U3237) );
  INV_X1 U8653 ( .A(n7029), .ZN(n7034) );
  NAND2_X1 U8654 ( .A1(n8527), .A2(n7314), .ZN(n7036) );
  INV_X1 U8655 ( .A(n7036), .ZN(n7030) );
  NOR2_X1 U8656 ( .A1(n7045), .A2(n7030), .ZN(n7035) );
  OR2_X1 U8657 ( .A1(n7031), .A2(n7035), .ZN(n7282) );
  INV_X1 U8658 ( .A(n8526), .ZN(n7050) );
  NAND2_X1 U8659 ( .A1(n7050), .A2(n9807), .ZN(n7032) );
  INV_X1 U8660 ( .A(n7032), .ZN(n7040) );
  NAND2_X1 U8661 ( .A1(n7034), .A2(n7033), .ZN(n7065) );
  INV_X1 U8662 ( .A(n7035), .ZN(n7039) );
  NAND2_X1 U8663 ( .A1(n7037), .A2(n7036), .ZN(n7038) );
  XNOR2_X1 U8664 ( .A(n8219), .B(n8526), .ZN(n7284) );
  INV_X1 U8665 ( .A(n7284), .ZN(n8350) );
  NAND2_X1 U8666 ( .A1(n7041), .A2(n7032), .ZN(n7063) );
  NAND2_X1 U8667 ( .A1(n7065), .A2(n7063), .ZN(n7043) );
  OR2_X1 U8668 ( .A1(n7062), .A2(n7296), .ZN(n8225) );
  NAND2_X1 U8669 ( .A1(n7062), .A2(n7296), .ZN(n8224) );
  NAND2_X1 U8670 ( .A1(n7043), .A2(n8345), .ZN(n7042) );
  OAI21_X1 U8671 ( .B1(n7043), .B2(n8345), .A(n7042), .ZN(n7244) );
  INV_X1 U8672 ( .A(n7044), .ZN(n7047) );
  INV_X1 U8673 ( .A(n7045), .ZN(n7046) );
  AND2_X1 U8674 ( .A1(n8215), .A2(n7284), .ZN(n7048) );
  NAND2_X1 U8675 ( .A1(n9807), .A2(n8526), .ZN(n7049) );
  XNOR2_X1 U8676 ( .A(n7073), .B(n8345), .ZN(n7053) );
  OAI22_X1 U8677 ( .A1(n7050), .A2(n8719), .B1(n7078), .B2(n8721), .ZN(n7052)
         );
  NOR2_X1 U8678 ( .A1(n7244), .A2(n8729), .ZN(n7051) );
  AOI211_X1 U8679 ( .C1(n9759), .C2(n7053), .A(n7052), .B(n7051), .ZN(n7249)
         );
  OR2_X1 U8680 ( .A1(n7286), .A2(n8219), .ZN(n7287) );
  NOR2_X2 U8681 ( .A1(n7287), .A2(n7062), .ZN(n7362) );
  AOI21_X1 U8682 ( .B1(n7062), .B2(n7287), .A(n7362), .ZN(n7247) );
  AOI22_X1 U8683 ( .A1(n7247), .A2(n5731), .B1(n8849), .B2(n7062), .ZN(n7054)
         );
  OAI211_X1 U8684 ( .C1(n9381), .C2(n7244), .A(n7249), .B(n7054), .ZN(n7056)
         );
  NAND2_X1 U8685 ( .A1(n7056), .A2(n9836), .ZN(n7055) );
  OAI21_X1 U8686 ( .B1(n9836), .B2(n6513), .A(n7055), .ZN(P2_U3528) );
  INV_X1 U8687 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n7058) );
  NAND2_X1 U8688 ( .A1(n7056), .A2(n9828), .ZN(n7057) );
  OAI21_X1 U8689 ( .B1(n9828), .B2(n7058), .A(n7057), .ZN(P2_U3475) );
  NAND2_X1 U8690 ( .A1(n7060), .A2(n7059), .ZN(n7061) );
  OAI211_X1 U8691 ( .C1(n9961), .C2(n7969), .A(n7061), .B(n8385), .ZN(P2_U3335) );
  INV_X1 U8692 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n7085) );
  NAND2_X1 U8693 ( .A1(n7062), .A2(n8525), .ZN(n7066) );
  AND2_X1 U8694 ( .A1(n7063), .A2(n7066), .ZN(n7064) );
  NAND2_X1 U8695 ( .A1(n7065), .A2(n7064), .ZN(n7069) );
  INV_X1 U8696 ( .A(n7066), .ZN(n7067) );
  OR2_X1 U8697 ( .A1(n7067), .A2(n8345), .ZN(n7068) );
  NAND2_X1 U8698 ( .A1(n7069), .A2(n7068), .ZN(n7357) );
  OR2_X1 U8699 ( .A1(n7366), .A2(n7078), .ZN(n8233) );
  NAND2_X1 U8700 ( .A1(n7366), .A2(n7078), .ZN(n8229) );
  NAND2_X1 U8701 ( .A1(n8233), .A2(n8229), .ZN(n8349) );
  OR2_X1 U8702 ( .A1(n7366), .A2(n8524), .ZN(n7070) );
  OR2_X1 U8703 ( .A1(n7322), .A2(n7376), .ZN(n8234) );
  NAND2_X1 U8704 ( .A1(n7322), .A2(n7376), .ZN(n8235) );
  NAND2_X1 U8705 ( .A1(n7071), .A2(n7075), .ZN(n7072) );
  NAND2_X1 U8706 ( .A1(n7324), .A2(n7072), .ZN(n7139) );
  NAND2_X1 U8707 ( .A1(n7077), .A2(n8229), .ZN(n7074) );
  INV_X1 U8708 ( .A(n7075), .ZN(n8352) );
  AOI21_X1 U8709 ( .B1(n7074), .B2(n8352), .A(n8698), .ZN(n7080) );
  AND2_X1 U8710 ( .A1(n8229), .A2(n7075), .ZN(n7076) );
  NAND2_X1 U8711 ( .A1(n7077), .A2(n7076), .ZN(n7327) );
  OAI22_X1 U8712 ( .A1(n7078), .A2(n8719), .B1(n7442), .B2(n8721), .ZN(n7079)
         );
  AOI21_X1 U8713 ( .B1(n7080), .B2(n7327), .A(n7079), .ZN(n7081) );
  OAI21_X1 U8714 ( .B1(n7139), .B2(n8729), .A(n7081), .ZN(n7131) );
  NAND2_X1 U8715 ( .A1(n7362), .A2(n9811), .ZN(n7364) );
  OR2_X1 U8716 ( .A1(n7364), .A2(n7322), .ZN(n7377) );
  NAND2_X1 U8717 ( .A1(n7364), .A2(n7322), .ZN(n7082) );
  AND2_X1 U8718 ( .A1(n7377), .A2(n7082), .ZN(n7136) );
  AOI22_X1 U8719 ( .A1(n7136), .A2(n5731), .B1(n8849), .B2(n7322), .ZN(n7083)
         );
  OAI21_X1 U8720 ( .B1(n7139), .B2(n9381), .A(n7083), .ZN(n7084) );
  NOR2_X1 U8721 ( .A1(n7131), .A2(n7084), .ZN(n7087) );
  MUX2_X1 U8722 ( .A(n7085), .B(n7087), .S(n9828), .Z(n7086) );
  INV_X1 U8723 ( .A(n7086), .ZN(P2_U3481) );
  MUX2_X1 U8724 ( .A(n7088), .B(n7087), .S(n9836), .Z(n7089) );
  INV_X1 U8725 ( .A(n7089), .ZN(P2_U3530) );
  NAND2_X1 U8726 ( .A1(n7090), .A2(n7415), .ZN(n7092) );
  OR2_X1 U8727 ( .A1(n9006), .A2(n7091), .ZN(n7407) );
  NAND2_X1 U8728 ( .A1(n7092), .A2(n7407), .ZN(n7093) );
  OR2_X1 U8729 ( .A1(n7093), .A2(n7096), .ZN(n7095) );
  NAND2_X1 U8730 ( .A1(n7093), .A2(n7096), .ZN(n7094) );
  NAND2_X1 U8731 ( .A1(n7095), .A2(n7094), .ZN(n9650) );
  AOI22_X1 U8732 ( .A1(n9586), .A2(n9006), .B1(n9004), .B2(n9261), .ZN(n7100)
         );
  XNOR2_X1 U8733 ( .A(n7097), .B(n7096), .ZN(n7098) );
  NAND2_X1 U8734 ( .A1(n7098), .A2(n9427), .ZN(n7099) );
  OAI211_X1 U8735 ( .C1(n9650), .C2(n9279), .A(n7100), .B(n7099), .ZN(n9653)
         );
  NAND2_X1 U8736 ( .A1(n9653), .A2(n9600), .ZN(n7107) );
  OAI22_X1 U8737 ( .A1(n9600), .A2(n7101), .B1(n7351), .B2(n9418), .ZN(n7105)
         );
  AND2_X1 U8738 ( .A1(n7102), .A2(n7405), .ZN(n7103) );
  NOR2_X1 U8739 ( .A1(n7102), .A2(n7405), .ZN(n7481) );
  OR2_X1 U8740 ( .A1(n7103), .A2(n7481), .ZN(n9652) );
  NOR2_X1 U8741 ( .A1(n9652), .A2(n7807), .ZN(n7104) );
  AOI211_X1 U8742 ( .C1(n9434), .C2(n7405), .A(n7105), .B(n7104), .ZN(n7106)
         );
  OAI211_X1 U8743 ( .C1(n9650), .C2(n9268), .A(n7107), .B(n7106), .ZN(P1_U3283) );
  AND2_X1 U8744 ( .A1(n7109), .A2(n7108), .ZN(n7110) );
  NAND3_X1 U8745 ( .A1(n9774), .A2(n7111), .A3(n7110), .ZN(n7119) );
  INV_X1 U8746 ( .A(n7112), .ZN(n7113) );
  NAND2_X1 U8747 ( .A1(n9774), .A2(n7113), .ZN(n8731) );
  NAND2_X2 U8748 ( .A1(n7119), .A2(n8731), .ZN(n8734) );
  NAND2_X1 U8749 ( .A1(n5733), .A2(n4282), .ZN(n7114) );
  OR2_X1 U8750 ( .A1(n7114), .A2(n8373), .ZN(n7129) );
  NAND2_X1 U8751 ( .A1(n8729), .A2(n7129), .ZN(n7115) );
  INV_X1 U8752 ( .A(n8761), .ZN(n9765) );
  NOR2_X1 U8753 ( .A1(n7117), .A2(n7116), .ZN(n7118) );
  OR2_X1 U8754 ( .A1(n7119), .A2(n4282), .ZN(n7293) );
  INV_X1 U8755 ( .A(n7293), .ZN(n8676) );
  OAI22_X1 U8756 ( .A1(n8734), .A2(n6500), .B1(n7120), .B2(n8731), .ZN(n7121)
         );
  AOI21_X1 U8757 ( .B1(n7122), .B2(n8676), .A(n7121), .ZN(n7123) );
  OAI21_X1 U8758 ( .B1(n7124), .B2(n9768), .A(n7123), .ZN(n7125) );
  AOI21_X1 U8759 ( .B1(n9765), .B2(n7126), .A(n7125), .ZN(n7127) );
  OAI21_X1 U8760 ( .B1(n7128), .B2(n9772), .A(n7127), .ZN(P2_U3292) );
  INV_X1 U8761 ( .A(n7129), .ZN(n7130) );
  NAND2_X1 U8762 ( .A1(n8734), .A2(n7130), .ZN(n8739) );
  NAND2_X1 U8763 ( .A1(n7131), .A2(n8734), .ZN(n7138) );
  NOR2_X1 U8764 ( .A1(n7293), .A2(n4275), .ZN(n9762) );
  INV_X1 U8765 ( .A(n8731), .ZN(n9760) );
  AOI22_X1 U8766 ( .A1(n9772), .A2(P2_REG2_REG_10__SCAN_IN), .B1(n7132), .B2(
        n9760), .ZN(n7133) );
  OAI21_X1 U8767 ( .B1(n7134), .B2(n9768), .A(n7133), .ZN(n7135) );
  AOI21_X1 U8768 ( .B1(n7136), .B2(n9762), .A(n7135), .ZN(n7137) );
  OAI211_X1 U8769 ( .C1(n7139), .C2(n8739), .A(n7138), .B(n7137), .ZN(P2_U3286) );
  AOI21_X1 U8770 ( .B1(n7142), .B2(n7141), .A(n7140), .ZN(n7143) );
  NAND2_X1 U8771 ( .A1(n8564), .A2(n7143), .ZN(n7144) );
  XOR2_X1 U8772 ( .A(n8564), .B(n7143), .Z(n8559) );
  NAND2_X1 U8773 ( .A1(P2_REG1_REG_15__SCAN_IN), .A2(n8559), .ZN(n8558) );
  NAND2_X1 U8774 ( .A1(n7144), .A2(n8558), .ZN(n7146) );
  INV_X1 U8775 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n9977) );
  XNOR2_X1 U8776 ( .A(n7620), .B(n9977), .ZN(n7145) );
  NOR2_X1 U8777 ( .A1(n7146), .A2(n7145), .ZN(n7619) );
  AOI21_X1 U8778 ( .B1(n7146), .B2(n7145), .A(n7619), .ZN(n7162) );
  INV_X1 U8779 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n7147) );
  NAND2_X1 U8780 ( .A1(P2_REG3_REG_16__SCAN_IN), .A2(P2_U3152), .ZN(n7788) );
  OAI21_X1 U8781 ( .B1(n8068), .B2(n7147), .A(n7788), .ZN(n7148) );
  AOI21_X1 U8782 ( .B1(n7156), .B2(n9747), .A(n7148), .ZN(n7161) );
  NOR2_X1 U8783 ( .A1(P2_REG2_REG_14__SCAN_IN), .A2(n7149), .ZN(n7151) );
  NOR2_X1 U8784 ( .A1(n8564), .A2(n7152), .ZN(n7153) );
  NOR2_X1 U8785 ( .A1(P2_REG2_REG_15__SCAN_IN), .A2(n8562), .ZN(n8561) );
  NOR2_X1 U8786 ( .A1(n7153), .A2(n8561), .ZN(n7159) );
  NAND2_X1 U8787 ( .A1(n7620), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n7154) );
  OAI21_X1 U8788 ( .B1(n7620), .B2(P2_REG2_REG_16__SCAN_IN), .A(n7154), .ZN(
        n7158) );
  INV_X1 U8789 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n7155) );
  NAND2_X1 U8790 ( .A1(n7620), .A2(n7155), .ZN(n7157) );
  NAND2_X1 U8791 ( .A1(n7156), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n7610) );
  NAND3_X1 U8792 ( .A1(n7159), .A2(n7157), .A3(n7610), .ZN(n7611) );
  OAI211_X1 U8793 ( .C1(n7159), .C2(n7158), .A(n7611), .B(n9744), .ZN(n7160)
         );
  OAI211_X1 U8794 ( .C1(n7162), .C2(n9681), .A(n7161), .B(n7160), .ZN(P2_U3261) );
  INV_X1 U8795 ( .A(n7163), .ZN(n7198) );
  OAI222_X1 U8796 ( .A1(n8073), .A2(n7198), .B1(P1_U3084), .B2(n7165), .C1(
        n7164), .C2(n8069), .ZN(P1_U3329) );
  INV_X1 U8797 ( .A(n7166), .ZN(n7169) );
  INV_X1 U8798 ( .A(n7167), .ZN(n7168) );
  NAND2_X1 U8799 ( .A1(n7169), .A2(n7168), .ZN(n7170) );
  OR2_X1 U8800 ( .A1(n7176), .A2(n6359), .ZN(n7174) );
  NAND2_X1 U8801 ( .A1(n9005), .A2(n7904), .ZN(n7173) );
  AND2_X1 U8802 ( .A1(n7174), .A2(n7173), .ZN(n7178) );
  NAND2_X1 U8803 ( .A1(n7179), .A2(n7178), .ZN(n7342) );
  NAND2_X1 U8804 ( .A1(n9005), .A2(n7939), .ZN(n7175) );
  OAI21_X1 U8805 ( .B1(n7176), .B2(n6384), .A(n7175), .ZN(n7177) );
  XNOR2_X1 U8806 ( .A(n7177), .B(n6860), .ZN(n7343) );
  NAND2_X1 U8807 ( .A1(n7484), .A2(n7933), .ZN(n7181) );
  NAND2_X1 U8808 ( .A1(n9004), .A2(n7939), .ZN(n7180) );
  NAND2_X1 U8809 ( .A1(n7181), .A2(n7180), .ZN(n7182) );
  XNOR2_X1 U8810 ( .A(n7182), .B(n7936), .ZN(n7184) );
  AND2_X1 U8811 ( .A1(n9004), .A2(n7904), .ZN(n7183) );
  AOI21_X1 U8812 ( .B1(n7484), .B2(n7939), .A(n7183), .ZN(n7185) );
  NAND2_X1 U8813 ( .A1(n7184), .A2(n7185), .ZN(n7390) );
  INV_X1 U8814 ( .A(n7184), .ZN(n7187) );
  INV_X1 U8815 ( .A(n7185), .ZN(n7186) );
  NAND2_X1 U8816 ( .A1(n7187), .A2(n7186), .ZN(n7188) );
  AND2_X1 U8817 ( .A1(n7390), .A2(n7188), .ZN(n7189) );
  INV_X1 U8818 ( .A(n7391), .ZN(n7191) );
  AOI21_X1 U8819 ( .B1(n7341), .B2(n7345), .A(n7189), .ZN(n7190) );
  OAI21_X1 U8820 ( .B1(n7191), .B2(n7190), .A(n8973), .ZN(n7196) );
  AND2_X1 U8821 ( .A1(P1_U3084), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n9526) );
  AOI21_X1 U8822 ( .B1(n8965), .B2(n9005), .A(n9526), .ZN(n7193) );
  OR2_X1 U8823 ( .A1(n8963), .A2(n9424), .ZN(n7192) );
  OAI211_X1 U8824 ( .C1(n8989), .C2(n7482), .A(n7193), .B(n7192), .ZN(n7194)
         );
  AOI21_X1 U8825 ( .B1(n8968), .B2(n7484), .A(n7194), .ZN(n7195) );
  NAND2_X1 U8826 ( .A1(n7196), .A2(n7195), .ZN(P1_U3229) );
  OAI222_X1 U8827 ( .A1(P2_U3152), .A2(n7199), .B1(n4284), .B2(n7198), .C1(
        n7197), .C2(n7969), .ZN(P2_U3334) );
  MUX2_X1 U8828 ( .A(n6498), .B(n7200), .S(n8734), .Z(n7205) );
  INV_X1 U8829 ( .A(n9762), .ZN(n8708) );
  INV_X1 U8830 ( .A(n7201), .ZN(n7202) );
  INV_X1 U8831 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n7975) );
  OAI22_X1 U8832 ( .A1(n8708), .A2(n7202), .B1(n7975), .B2(n8731), .ZN(n7203)
         );
  AOI21_X1 U8833 ( .B1(n8736), .B2(n7972), .A(n7203), .ZN(n7204) );
  OAI211_X1 U8834 ( .C1(n7206), .C2(n8761), .A(n7205), .B(n7204), .ZN(P2_U3294) );
  OAI21_X1 U8835 ( .B1(n7209), .B2(n7208), .A(n7207), .ZN(n9796) );
  INV_X1 U8836 ( .A(n9796), .ZN(n7225) );
  OAI22_X1 U8837 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(n8731), .B1(n8734), .B2(
        n7210), .ZN(n7214) );
  OAI21_X1 U8838 ( .B1(n9792), .B2(n7212), .A(n7211), .ZN(n9793) );
  NOR2_X1 U8839 ( .A1(n8708), .A2(n9793), .ZN(n7213) );
  AOI211_X1 U8840 ( .C1(n8736), .C2(n7215), .A(n7214), .B(n7213), .ZN(n7224)
         );
  OAI21_X1 U8841 ( .B1(n8341), .B2(n7217), .A(n7216), .ZN(n7221) );
  OAI22_X1 U8842 ( .A1(n7219), .A2(n8719), .B1(n7218), .B2(n8721), .ZN(n7220)
         );
  AOI21_X1 U8843 ( .B1(n7221), .B2(n9759), .A(n7220), .ZN(n7222) );
  OAI21_X1 U8844 ( .B1(n7225), .B2(n8729), .A(n7222), .ZN(n9794) );
  NAND2_X1 U8845 ( .A1(n9794), .A2(n8734), .ZN(n7223) );
  OAI211_X1 U8846 ( .C1(n7225), .C2(n8739), .A(n7224), .B(n7223), .ZN(P2_U3293) );
  XNOR2_X1 U8847 ( .A(n8346), .B(n7029), .ZN(n9799) );
  XNOR2_X1 U8848 ( .A(n7227), .B(n7226), .ZN(n7228) );
  NAND2_X1 U8849 ( .A1(n7228), .A2(n9759), .ZN(n7230) );
  AOI22_X1 U8850 ( .A1(n8753), .A2(n8529), .B1(n8527), .B2(n8755), .ZN(n7229)
         );
  NAND2_X1 U8851 ( .A1(n7230), .A2(n7229), .ZN(n9802) );
  OAI211_X1 U8852 ( .C1(n7232), .C2(n6748), .A(n5731), .B(n7231), .ZN(n9800)
         );
  NOR2_X1 U8853 ( .A1(n9800), .A2(n4282), .ZN(n7233) );
  OAI21_X1 U8854 ( .B1(n9802), .B2(n7233), .A(n8734), .ZN(n7240) );
  INV_X1 U8855 ( .A(n7234), .ZN(n7235) );
  OAI22_X1 U8856 ( .A1(n8734), .A2(n7236), .B1(n7235), .B2(n8731), .ZN(n7237)
         );
  AOI21_X1 U8857 ( .B1(n8736), .B2(n7238), .A(n7237), .ZN(n7239) );
  OAI211_X1 U8858 ( .C1(n9799), .C2(n8761), .A(n7240), .B(n7239), .ZN(P2_U3291) );
  AOI22_X1 U8859 ( .A1(n9772), .A2(P2_REG2_REG_8__SCAN_IN), .B1(n7241), .B2(
        n9760), .ZN(n7242) );
  OAI21_X1 U8860 ( .B1(n7243), .B2(n9768), .A(n7242), .ZN(n7246) );
  NOR2_X1 U8861 ( .A1(n7244), .A2(n8739), .ZN(n7245) );
  AOI211_X1 U8862 ( .C1(n7247), .C2(n9762), .A(n7246), .B(n7245), .ZN(n7248)
         );
  OAI21_X1 U8863 ( .B1(n7249), .B2(n9772), .A(n7248), .ZN(P2_U3288) );
  INV_X1 U8864 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n7264) );
  NAND2_X1 U8865 ( .A1(n7250), .A2(n7258), .ZN(n7252) );
  NAND2_X1 U8866 ( .A1(n7252), .A2(n7251), .ZN(n7525) );
  XOR2_X1 U8867 ( .A(n7533), .B(n7525), .Z(n7253) );
  NOR2_X1 U8868 ( .A1(n7253), .A2(n7804), .ZN(n7526) );
  AOI211_X1 U8869 ( .C1(n7253), .C2(n7804), .A(n9543), .B(n7526), .ZN(n7254)
         );
  INV_X1 U8870 ( .A(n7254), .ZN(n7263) );
  NAND2_X1 U8871 ( .A1(P1_U3084), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n8990) );
  INV_X1 U8872 ( .A(n8990), .ZN(n7261) );
  INV_X1 U8873 ( .A(n7255), .ZN(n7256) );
  AOI21_X1 U8874 ( .B1(n7258), .B2(n7257), .A(n7256), .ZN(n7534) );
  XNOR2_X1 U8875 ( .A(n7533), .B(n7534), .ZN(n7259) );
  NOR2_X1 U8876 ( .A1(n7259), .A2(n5247), .ZN(n7532) );
  AOI211_X1 U8877 ( .C1(n5247), .C2(n7259), .A(n7532), .B(n9522), .ZN(n7260)
         );
  AOI211_X1 U8878 ( .C1(n7533), .C2(n9553), .A(n7261), .B(n7260), .ZN(n7262)
         );
  OAI211_X1 U8879 ( .C1(n9571), .C2(n7264), .A(n7263), .B(n7262), .ZN(P1_U3256) );
  OAI21_X1 U8880 ( .B1(n7266), .B2(n8731), .A(n7265), .ZN(n7268) );
  INV_X1 U8881 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n8532) );
  NOR2_X1 U8882 ( .A1(n8734), .A2(n8532), .ZN(n7267) );
  AOI21_X1 U8883 ( .B1(n7268), .B2(n8734), .A(n7267), .ZN(n7270) );
  OAI21_X1 U8884 ( .B1(n9762), .B2(n8736), .A(n9761), .ZN(n7269) );
  OAI211_X1 U8885 ( .C1(n8340), .C2(n8761), .A(n7270), .B(n7269), .ZN(P2_U3296) );
  XOR2_X1 U8886 ( .A(n7271), .B(n7272), .Z(n7280) );
  NAND2_X1 U8887 ( .A1(n9818), .A2(n8509), .ZN(n7278) );
  OAI22_X1 U8888 ( .A1(n8502), .A2(n7453), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7273), .ZN(n7274) );
  INV_X1 U8889 ( .A(n7274), .ZN(n7277) );
  NAND2_X1 U8890 ( .A1(n8496), .A2(n7379), .ZN(n7276) );
  INV_X1 U8891 ( .A(n7376), .ZN(n8523) );
  NAND2_X1 U8892 ( .A1(n8504), .A2(n8523), .ZN(n7275) );
  NAND4_X1 U8893 ( .A1(n7278), .A2(n7277), .A3(n7276), .A4(n7275), .ZN(n7279)
         );
  AOI21_X1 U8894 ( .B1(n7280), .B2(n8473), .A(n7279), .ZN(n7281) );
  INV_X1 U8895 ( .A(n7281), .ZN(P2_U3238) );
  OR2_X1 U8896 ( .A1(n7029), .A2(n7282), .ZN(n7283) );
  XNOR2_X1 U8897 ( .A(n7285), .B(n7284), .ZN(n9809) );
  AOI21_X1 U8898 ( .B1(n7286), .B2(n8219), .A(n4275), .ZN(n7288) );
  NAND2_X1 U8899 ( .A1(n7288), .A2(n7287), .ZN(n9805) );
  INV_X1 U8900 ( .A(n7289), .ZN(n7290) );
  OAI22_X1 U8901 ( .A1(n8734), .A2(n6521), .B1(n7290), .B2(n8731), .ZN(n7291)
         );
  AOI21_X1 U8902 ( .B1(n8736), .B2(n8219), .A(n7291), .ZN(n7292) );
  OAI21_X1 U8903 ( .B1(n9805), .B2(n7293), .A(n7292), .ZN(n7302) );
  NAND2_X1 U8904 ( .A1(n7294), .A2(n8215), .ZN(n7295) );
  AOI21_X1 U8905 ( .B1(n7295), .B2(n8350), .A(n8698), .ZN(n7300) );
  INV_X1 U8906 ( .A(n8527), .ZN(n7297) );
  OAI22_X1 U8907 ( .A1(n7297), .A2(n8719), .B1(n7296), .B2(n8721), .ZN(n7298)
         );
  AOI21_X1 U8908 ( .B1(n7300), .B2(n7299), .A(n7298), .ZN(n9806) );
  NOR2_X1 U8909 ( .A1(n9806), .A2(n9772), .ZN(n7301) );
  AOI211_X1 U8910 ( .C1(n9765), .C2(n9809), .A(n7302), .B(n7301), .ZN(n7303)
         );
  INV_X1 U8911 ( .A(n7303), .ZN(P2_U3289) );
  NAND2_X1 U8912 ( .A1(n7305), .A2(n7304), .ZN(n7307) );
  XOR2_X1 U8913 ( .A(n7307), .B(n7306), .Z(n7313) );
  INV_X1 U8914 ( .A(n7442), .ZN(n8522) );
  NAND2_X1 U8915 ( .A1(n8504), .A2(n8522), .ZN(n7309) );
  OAI211_X1 U8916 ( .C1(n7679), .C2(n8502), .A(n7309), .B(n7308), .ZN(n7311)
         );
  INV_X1 U8917 ( .A(n8848), .ZN(n7438) );
  NOR2_X1 U8918 ( .A1(n7438), .A2(n8499), .ZN(n7310) );
  AOI211_X1 U8919 ( .C1(n8496), .C2(n7436), .A(n7311), .B(n7310), .ZN(n7312)
         );
  OAI21_X1 U8920 ( .B1(n7313), .B2(n8511), .A(n7312), .ZN(P2_U3226) );
  AOI22_X1 U8921 ( .A1(n8736), .A2(n7314), .B1(n7962), .B2(n9760), .ZN(n7315)
         );
  OAI21_X1 U8922 ( .B1(n7316), .B2(n8708), .A(n7315), .ZN(n7319) );
  MUX2_X1 U8923 ( .A(P2_REG2_REG_6__SCAN_IN), .B(n7317), .S(n8734), .Z(n7318)
         );
  AOI211_X1 U8924 ( .C1(n9765), .C2(n7320), .A(n7319), .B(n7318), .ZN(n7321)
         );
  INV_X1 U8925 ( .A(n7321), .ZN(P2_U3290) );
  NAND2_X1 U8926 ( .A1(n7322), .A2(n8523), .ZN(n7323) );
  NAND2_X1 U8927 ( .A1(n7324), .A2(n7323), .ZN(n7373) );
  NAND2_X1 U8928 ( .A1(n9818), .A2(n7442), .ZN(n8241) );
  NAND2_X1 U8929 ( .A1(n8242), .A2(n8241), .ZN(n7372) );
  AND2_X1 U8930 ( .A1(n9818), .A2(n8522), .ZN(n7325) );
  AOI21_X2 U8931 ( .B1(n7373), .B2(n7372), .A(n7325), .ZN(n7431) );
  INV_X1 U8932 ( .A(n7453), .ZN(n8521) );
  OR2_X1 U8933 ( .A1(n7599), .A2(n7679), .ZN(n8251) );
  NAND2_X1 U8934 ( .A1(n7599), .A2(n7679), .ZN(n8250) );
  XNOR2_X1 U8935 ( .A(n7601), .B(n7329), .ZN(n9385) );
  INV_X1 U8936 ( .A(n8729), .ZN(n7358) );
  INV_X1 U8937 ( .A(n7430), .ZN(n8355) );
  INV_X1 U8938 ( .A(n7330), .ZN(n7328) );
  NAND2_X1 U8939 ( .A1(n7330), .A2(n7329), .ZN(n7331) );
  NAND2_X1 U8940 ( .A1(n7677), .A2(n7331), .ZN(n7332) );
  NAND2_X1 U8941 ( .A1(n7332), .A2(n9759), .ZN(n7334) );
  AOI22_X1 U8942 ( .A1(n8521), .A2(n8753), .B1(n8755), .B2(n8519), .ZN(n7333)
         );
  NAND2_X1 U8943 ( .A1(n7334), .A2(n7333), .ZN(n7335) );
  AOI21_X1 U8944 ( .B1(n9385), .B2(n7358), .A(n7335), .ZN(n9387) );
  INV_X1 U8945 ( .A(n8739), .ZN(n7666) );
  INV_X1 U8946 ( .A(n7599), .ZN(n9382) );
  OR2_X1 U8947 ( .A1(n7434), .A2(n9382), .ZN(n7336) );
  NAND2_X1 U8948 ( .A1(n7675), .A2(n7336), .ZN(n9383) );
  AOI22_X1 U8949 ( .A1(n9772), .A2(P2_REG2_REG_13__SCAN_IN), .B1(n7455), .B2(
        n9760), .ZN(n7338) );
  NAND2_X1 U8950 ( .A1(n7599), .A2(n8736), .ZN(n7337) );
  OAI211_X1 U8951 ( .C1(n9383), .C2(n8708), .A(n7338), .B(n7337), .ZN(n7339)
         );
  AOI21_X1 U8952 ( .B1(n9385), .B2(n7666), .A(n7339), .ZN(n7340) );
  OAI21_X1 U8953 ( .B1(n9387), .B2(n9772), .A(n7340), .ZN(P2_U3283) );
  INV_X1 U8954 ( .A(n7341), .ZN(n7346) );
  AOI21_X1 U8955 ( .B1(n7345), .B2(n7342), .A(n7343), .ZN(n7344) );
  AOI211_X1 U8956 ( .C1(n7346), .C2(n7345), .A(n8984), .B(n7344), .ZN(n7354)
         );
  INV_X1 U8957 ( .A(n7347), .ZN(n7646) );
  NAND2_X1 U8958 ( .A1(n7405), .A2(n9345), .ZN(n9651) );
  NOR2_X1 U8959 ( .A1(n7646), .A2(n9651), .ZN(n7353) );
  AOI21_X1 U8960 ( .B1(n8994), .B2(n9004), .A(n7348), .ZN(n7350) );
  NAND2_X1 U8961 ( .A1(n8965), .A2(n9006), .ZN(n7349) );
  OAI211_X1 U8962 ( .C1(n8989), .C2(n7351), .A(n7350), .B(n7349), .ZN(n7352)
         );
  OR3_X1 U8963 ( .A1(n7354), .A2(n7353), .A3(n7352), .ZN(P1_U3219) );
  XNOR2_X1 U8964 ( .A(n7355), .B(n8349), .ZN(n7361) );
  OAI21_X1 U8965 ( .B1(n7357), .B2(n8349), .A(n7356), .ZN(n9815) );
  NAND2_X1 U8966 ( .A1(n9815), .A2(n7358), .ZN(n7360) );
  AOI22_X1 U8967 ( .A1(n8753), .A2(n8525), .B1(n8523), .B2(n8755), .ZN(n7359)
         );
  OAI211_X1 U8968 ( .C1(n8698), .C2(n7361), .A(n7360), .B(n7359), .ZN(n9813)
         );
  INV_X1 U8969 ( .A(n9813), .ZN(n7371) );
  OR2_X1 U8970 ( .A1(n7362), .A2(n9811), .ZN(n7363) );
  NAND2_X1 U8971 ( .A1(n7364), .A2(n7363), .ZN(n9812) );
  AOI22_X1 U8972 ( .A1(n9772), .A2(P2_REG2_REG_9__SCAN_IN), .B1(n7365), .B2(
        n9760), .ZN(n7368) );
  NAND2_X1 U8973 ( .A1(n8736), .A2(n7366), .ZN(n7367) );
  OAI211_X1 U8974 ( .C1(n9812), .C2(n8708), .A(n7368), .B(n7367), .ZN(n7369)
         );
  AOI21_X1 U8975 ( .B1(n9815), .B2(n7666), .A(n7369), .ZN(n7370) );
  OAI21_X1 U8976 ( .B1(n7371), .B2(n9772), .A(n7370), .ZN(P2_U3287) );
  INV_X1 U8977 ( .A(n7372), .ZN(n8354) );
  XNOR2_X1 U8978 ( .A(n7373), .B(n8354), .ZN(n9826) );
  INV_X1 U8979 ( .A(n9826), .ZN(n7385) );
  XNOR2_X1 U8980 ( .A(n7374), .B(n8354), .ZN(n7375) );
  OAI222_X1 U8981 ( .A1(n8721), .A2(n7453), .B1(n8719), .B2(n7376), .C1(n8698), 
        .C2(n7375), .ZN(n9823) );
  AND2_X1 U8982 ( .A1(n7377), .A2(n9818), .ZN(n7378) );
  OR2_X1 U8983 ( .A1(n7378), .A2(n7433), .ZN(n9822) );
  INV_X1 U8984 ( .A(n7379), .ZN(n7380) );
  OAI22_X1 U8985 ( .A1(n8734), .A2(n6557), .B1(n7380), .B2(n8731), .ZN(n7381)
         );
  AOI21_X1 U8986 ( .B1(n9818), .B2(n8736), .A(n7381), .ZN(n7382) );
  OAI21_X1 U8987 ( .B1(n9822), .B2(n8708), .A(n7382), .ZN(n7383) );
  AOI21_X1 U8988 ( .B1(n9823), .B2(n8734), .A(n7383), .ZN(n7384) );
  OAI21_X1 U8989 ( .B1(n8761), .B2(n7385), .A(n7384), .ZN(P2_U3285) );
  NAND2_X1 U8990 ( .A1(n7571), .A2(n7933), .ZN(n7387) );
  OR2_X1 U8991 ( .A1(n9424), .A2(n6359), .ZN(n7386) );
  NAND2_X1 U8992 ( .A1(n7387), .A2(n7386), .ZN(n7388) );
  XNOR2_X1 U8993 ( .A(n7388), .B(n6860), .ZN(n7462) );
  NOR2_X1 U8994 ( .A1(n9424), .A2(n7942), .ZN(n7389) );
  AOI21_X1 U8995 ( .B1(n7571), .B2(n7939), .A(n7389), .ZN(n7463) );
  XNOR2_X1 U8996 ( .A(n7462), .B(n7463), .ZN(n7393) );
  OAI21_X1 U8997 ( .B1(n7393), .B2(n7392), .A(n7471), .ZN(n7400) );
  INV_X1 U8998 ( .A(n7571), .ZN(n9376) );
  NOR2_X1 U8999 ( .A1(n8997), .A2(n9376), .ZN(n7399) );
  NOR2_X1 U9000 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7394), .ZN(n9540) );
  AOI21_X1 U9001 ( .B1(n8965), .B2(n9004), .A(n9540), .ZN(n7397) );
  OR2_X1 U9002 ( .A1(n8963), .A2(n7395), .ZN(n7396) );
  OAI211_X1 U9003 ( .C1(n8989), .C2(n7423), .A(n7397), .B(n7396), .ZN(n7398)
         );
  AOI211_X1 U9004 ( .C1(n7400), .C2(n8973), .A(n7399), .B(n7398), .ZN(n7401)
         );
  INV_X1 U9005 ( .A(n7401), .ZN(P1_U3215) );
  XNOR2_X1 U9006 ( .A(n7579), .B(n7420), .ZN(n7402) );
  NAND2_X1 U9007 ( .A1(n7402), .A2(n9427), .ZN(n7404) );
  AOI22_X1 U9008 ( .A1(n9261), .A2(n9002), .B1(n9004), .B2(n9586), .ZN(n7403)
         );
  NAND2_X1 U9009 ( .A1(n7404), .A2(n7403), .ZN(n9377) );
  INV_X1 U9010 ( .A(n9377), .ZN(n7428) );
  NAND2_X1 U9011 ( .A1(n7405), .A2(n9005), .ZN(n7414) );
  INV_X1 U9012 ( .A(n7414), .ZN(n7409) );
  AND2_X1 U9013 ( .A1(n7407), .A2(n7406), .ZN(n7408) );
  AND2_X1 U9014 ( .A1(n7410), .A2(n7413), .ZN(n7411) );
  OR2_X1 U9015 ( .A1(n7484), .A2(n9004), .ZN(n7416) );
  NAND2_X1 U9016 ( .A1(n7479), .A2(n7416), .ZN(n7418) );
  NAND2_X1 U9017 ( .A1(n7484), .A2(n9004), .ZN(n7417) );
  OAI21_X1 U9018 ( .B1(n7421), .B2(n7420), .A(n7573), .ZN(n9379) );
  INV_X1 U9019 ( .A(n7484), .ZN(n9659) );
  NAND2_X1 U9020 ( .A1(n7481), .A2(n9659), .ZN(n7480) );
  INV_X1 U9021 ( .A(n7480), .ZN(n7422) );
  OAI211_X1 U9022 ( .C1(n7422), .C2(n9376), .A(n9572), .B(n9413), .ZN(n9375)
         );
  OAI22_X1 U9023 ( .A1(n9600), .A2(n6433), .B1(n7423), .B2(n9418), .ZN(n7424)
         );
  AOI21_X1 U9024 ( .B1(n7571), .B2(n9434), .A(n7424), .ZN(n7425) );
  OAI21_X1 U9025 ( .B1(n9375), .B2(n7700), .A(n7425), .ZN(n7426) );
  AOI21_X1 U9026 ( .B1(n9379), .B2(n9597), .A(n7426), .ZN(n7427) );
  OAI21_X1 U9027 ( .B1(n4283), .B2(n7428), .A(n7427), .ZN(P1_U3281) );
  OAI21_X1 U9028 ( .B1(n7431), .B2(n7430), .A(n7429), .ZN(n7432) );
  INV_X1 U9029 ( .A(n7432), .ZN(n8853) );
  INV_X1 U9030 ( .A(n7433), .ZN(n7435) );
  AOI21_X1 U9031 ( .B1(n8848), .B2(n7435), .A(n7434), .ZN(n8850) );
  AOI22_X1 U9032 ( .A1(n9772), .A2(P2_REG2_REG_12__SCAN_IN), .B1(n7436), .B2(
        n9760), .ZN(n7437) );
  OAI21_X1 U9033 ( .B1(n7438), .B2(n9768), .A(n7437), .ZN(n7447) );
  INV_X1 U9034 ( .A(n8242), .ZN(n7439) );
  NOR2_X1 U9035 ( .A1(n8355), .A2(n7439), .ZN(n7440) );
  AOI21_X1 U9036 ( .B1(n7441), .B2(n7440), .A(n8698), .ZN(n7444) );
  OAI22_X1 U9037 ( .A1(n7679), .A2(n8721), .B1(n7442), .B2(n8719), .ZN(n7443)
         );
  AOI21_X1 U9038 ( .B1(n7445), .B2(n7444), .A(n7443), .ZN(n8852) );
  NOR2_X1 U9039 ( .A1(n8852), .A2(n9772), .ZN(n7446) );
  AOI211_X1 U9040 ( .C1(n8850), .C2(n9762), .A(n7447), .B(n7446), .ZN(n7448)
         );
  OAI21_X1 U9041 ( .B1(n8853), .B2(n8761), .A(n7448), .ZN(P2_U3284) );
  OAI211_X1 U9042 ( .C1(n7451), .C2(n7450), .A(n7449), .B(n8473), .ZN(n7457)
         );
  AOI22_X1 U9043 ( .A1(n8491), .A2(n8519), .B1(P2_REG3_REG_13__SCAN_IN), .B2(
        P2_U3152), .ZN(n7452) );
  OAI21_X1 U9044 ( .B1(n7453), .B2(n8493), .A(n7452), .ZN(n7454) );
  AOI21_X1 U9045 ( .B1(n7455), .B2(n8496), .A(n7454), .ZN(n7456) );
  OAI211_X1 U9046 ( .C1(n9382), .C2(n8499), .A(n7457), .B(n7456), .ZN(P2_U3236) );
  INV_X1 U9047 ( .A(n7991), .ZN(n7460) );
  OAI222_X1 U9048 ( .A1(n7969), .A2(n10000), .B1(n4284), .B2(n7460), .C1(n7458), .C2(P2_U3152), .ZN(P2_U3333) );
  OAI222_X1 U9049 ( .A1(n8069), .A2(n7461), .B1(n9371), .B2(n7460), .C1(n7459), 
        .C2(P1_U3084), .ZN(P1_U3328) );
  INV_X1 U9050 ( .A(n9433), .ZN(n9457) );
  INV_X1 U9051 ( .A(n7462), .ZN(n7464) );
  NAND2_X1 U9052 ( .A1(n7464), .A2(n7463), .ZN(n7469) );
  AND2_X1 U9053 ( .A1(n7471), .A2(n7469), .ZN(n7473) );
  NAND2_X1 U9054 ( .A1(n9433), .A2(n7933), .ZN(n7466) );
  NAND2_X1 U9055 ( .A1(n9002), .A2(n7939), .ZN(n7465) );
  NAND2_X1 U9056 ( .A1(n7466), .A2(n7465), .ZN(n7467) );
  XNOR2_X1 U9057 ( .A(n7467), .B(n6860), .ZN(n7548) );
  AND2_X1 U9058 ( .A1(n9002), .A2(n7904), .ZN(n7468) );
  AOI21_X1 U9059 ( .B1(n9433), .B2(n7939), .A(n7468), .ZN(n7546) );
  XNOR2_X1 U9060 ( .A(n7548), .B(n7546), .ZN(n7472) );
  AND2_X1 U9061 ( .A1(n7472), .A2(n7469), .ZN(n7470) );
  OAI211_X1 U9062 ( .C1(n7473), .C2(n7472), .A(n8973), .B(n7550), .ZN(n7478)
         );
  INV_X1 U9063 ( .A(n9419), .ZN(n7476) );
  INV_X1 U9064 ( .A(n8989), .ZN(n8979) );
  AND2_X1 U9065 ( .A1(P1_U3084), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n9569) );
  AOI21_X1 U9066 ( .B1(n8965), .B2(n9003), .A(n9569), .ZN(n7474) );
  OAI21_X1 U9067 ( .B1(n9425), .B2(n8963), .A(n7474), .ZN(n7475) );
  AOI21_X1 U9068 ( .B1(n7476), .B2(n8979), .A(n7475), .ZN(n7477) );
  OAI211_X1 U9069 ( .C1(n9457), .C2(n8997), .A(n7478), .B(n7477), .ZN(P1_U3234) );
  XOR2_X1 U9070 ( .A(n7486), .B(n7479), .Z(n9665) );
  OAI21_X1 U9071 ( .B1(n7481), .B2(n9659), .A(n7480), .ZN(n9661) );
  INV_X1 U9072 ( .A(n7482), .ZN(n7483) );
  AOI22_X1 U9073 ( .A1(n9434), .A2(n7484), .B1(n9588), .B2(n7483), .ZN(n7485)
         );
  OAI21_X1 U9074 ( .B1(n9661), .B2(n7807), .A(n7485), .ZN(n7491) );
  OAI211_X1 U9075 ( .C1(n4804), .C2(n5139), .A(n9427), .B(n7487), .ZN(n7489)
         );
  AOI22_X1 U9076 ( .A1(n9003), .A2(n9261), .B1(n9586), .B2(n9005), .ZN(n7488)
         );
  NAND2_X1 U9077 ( .A1(n7489), .A2(n7488), .ZN(n9662) );
  MUX2_X1 U9078 ( .A(P1_REG2_REG_9__SCAN_IN), .B(n9662), .S(n9600), .Z(n7490)
         );
  AOI211_X1 U9079 ( .C1(n9597), .C2(n9665), .A(n7491), .B(n7490), .ZN(n7492)
         );
  INV_X1 U9080 ( .A(n7492), .ZN(P1_U3282) );
  INV_X1 U9081 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n10031) );
  NOR2_X1 U9082 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n7493) );
  AOI21_X1 U9083 ( .B1(P1_ADDR_REG_17__SCAN_IN), .B2(P2_ADDR_REG_17__SCAN_IN), 
        .A(n7493), .ZN(n9847) );
  NOR2_X1 U9084 ( .A1(P1_ADDR_REG_16__SCAN_IN), .A2(P2_ADDR_REG_16__SCAN_IN), 
        .ZN(n7494) );
  AOI21_X1 U9085 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(P1_ADDR_REG_16__SCAN_IN), 
        .A(n7494), .ZN(n9850) );
  NOR2_X1 U9086 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n7495) );
  AOI21_X1 U9087 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(P2_ADDR_REG_15__SCAN_IN), 
        .A(n7495), .ZN(n9853) );
  NOR2_X1 U9088 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n7496) );
  AOI21_X1 U9089 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(P2_ADDR_REG_14__SCAN_IN), 
        .A(n7496), .ZN(n9856) );
  NOR2_X1 U9090 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n7497) );
  AOI21_X1 U9091 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(P2_ADDR_REG_13__SCAN_IN), 
        .A(n7497), .ZN(n9859) );
  NOR2_X1 U9092 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n7504) );
  XNOR2_X1 U9093 ( .A(P1_ADDR_REG_4__SCAN_IN), .B(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n10044) );
  NAND2_X1 U9094 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n7502) );
  XOR2_X1 U9095 ( .A(P1_ADDR_REG_3__SCAN_IN), .B(P2_ADDR_REG_3__SCAN_IN), .Z(
        n10042) );
  NAND2_X1 U9096 ( .A1(P2_ADDR_REG_2__SCAN_IN), .A2(P1_ADDR_REG_2__SCAN_IN), 
        .ZN(n7500) );
  XOR2_X1 U9097 ( .A(P2_ADDR_REG_2__SCAN_IN), .B(P1_ADDR_REG_2__SCAN_IN), .Z(
        n10040) );
  AOI21_X1 U9098 ( .B1(P2_ADDR_REG_0__SCAN_IN), .B2(P1_ADDR_REG_0__SCAN_IN), 
        .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n9841) );
  INV_X1 U9099 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n7498) );
  NAND3_X1 U9100 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .A3(P1_ADDR_REG_1__SCAN_IN), .ZN(n9843) );
  OAI21_X1 U9101 ( .B1(n9841), .B2(n7498), .A(n9843), .ZN(n10039) );
  NAND2_X1 U9102 ( .A1(n10040), .A2(n10039), .ZN(n7499) );
  NAND2_X1 U9103 ( .A1(n7500), .A2(n7499), .ZN(n10041) );
  NAND2_X1 U9104 ( .A1(n10042), .A2(n10041), .ZN(n7501) );
  NAND2_X1 U9105 ( .A1(n7502), .A2(n7501), .ZN(n10043) );
  NOR2_X1 U9106 ( .A1(n10044), .A2(n10043), .ZN(n7503) );
  NOR2_X1 U9107 ( .A1(n7504), .A2(n7503), .ZN(n7505) );
  NOR2_X1 U9108 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n7505), .ZN(n10025) );
  AND2_X1 U9109 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n7505), .ZN(n10026) );
  NOR2_X1 U9110 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n10026), .ZN(n7506) );
  NOR2_X1 U9111 ( .A1(n10025), .A2(n7506), .ZN(n7507) );
  NAND2_X1 U9112 ( .A1(n7507), .A2(P1_ADDR_REG_6__SCAN_IN), .ZN(n7509) );
  XOR2_X1 U9113 ( .A(n7507), .B(P1_ADDR_REG_6__SCAN_IN), .Z(n10024) );
  NAND2_X1 U9114 ( .A1(n10024), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n7508) );
  NAND2_X1 U9115 ( .A1(n7509), .A2(n7508), .ZN(n7510) );
  NAND2_X1 U9116 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(n7510), .ZN(n7512) );
  XOR2_X1 U9117 ( .A(P2_ADDR_REG_7__SCAN_IN), .B(n7510), .Z(n10038) );
  NAND2_X1 U9118 ( .A1(P1_ADDR_REG_7__SCAN_IN), .A2(n10038), .ZN(n7511) );
  NAND2_X1 U9119 ( .A1(n7512), .A2(n7511), .ZN(n7513) );
  NAND2_X1 U9120 ( .A1(P1_ADDR_REG_8__SCAN_IN), .A2(n7513), .ZN(n7515) );
  XOR2_X1 U9121 ( .A(P1_ADDR_REG_8__SCAN_IN), .B(n7513), .Z(n10036) );
  NAND2_X1 U9122 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(n10036), .ZN(n7514) );
  NAND2_X1 U9123 ( .A1(n7515), .A2(n7514), .ZN(n7516) );
  AND2_X1 U9124 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(n7516), .ZN(n7517) );
  INV_X1 U9125 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n10035) );
  XNOR2_X1 U9126 ( .A(P2_ADDR_REG_9__SCAN_IN), .B(n7516), .ZN(n10034) );
  NOR2_X1 U9127 ( .A1(n10035), .A2(n10034), .ZN(n10033) );
  NOR2_X1 U9128 ( .A1(n7517), .A2(n10033), .ZN(n9868) );
  NAND2_X1 U9129 ( .A1(P1_ADDR_REG_10__SCAN_IN), .A2(P2_ADDR_REG_10__SCAN_IN), 
        .ZN(n7518) );
  OAI21_X1 U9130 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(P2_ADDR_REG_10__SCAN_IN), 
        .A(n7518), .ZN(n9867) );
  NOR2_X1 U9131 ( .A1(n9868), .A2(n9867), .ZN(n9866) );
  AOI21_X1 U9132 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(P1_ADDR_REG_10__SCAN_IN), 
        .A(n9866), .ZN(n9865) );
  NAND2_X1 U9133 ( .A1(P1_ADDR_REG_11__SCAN_IN), .A2(P2_ADDR_REG_11__SCAN_IN), 
        .ZN(n7519) );
  OAI21_X1 U9134 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(P2_ADDR_REG_11__SCAN_IN), 
        .A(n7519), .ZN(n9864) );
  NOR2_X1 U9135 ( .A1(n9865), .A2(n9864), .ZN(n9863) );
  AOI21_X1 U9136 ( .B1(P2_ADDR_REG_11__SCAN_IN), .B2(P1_ADDR_REG_11__SCAN_IN), 
        .A(n9863), .ZN(n9862) );
  NOR2_X1 U9137 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n7520) );
  AOI21_X1 U9138 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(P2_ADDR_REG_12__SCAN_IN), 
        .A(n7520), .ZN(n9861) );
  NAND2_X1 U9139 ( .A1(n9862), .A2(n9861), .ZN(n9860) );
  OAI21_X1 U9140 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(P1_ADDR_REG_12__SCAN_IN), 
        .A(n9860), .ZN(n9858) );
  NAND2_X1 U9141 ( .A1(n9859), .A2(n9858), .ZN(n9857) );
  OAI21_X1 U9142 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(P1_ADDR_REG_13__SCAN_IN), 
        .A(n9857), .ZN(n9855) );
  NAND2_X1 U9143 ( .A1(n9856), .A2(n9855), .ZN(n9854) );
  OAI21_X1 U9144 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(P1_ADDR_REG_14__SCAN_IN), 
        .A(n9854), .ZN(n9852) );
  NAND2_X1 U9145 ( .A1(n9853), .A2(n9852), .ZN(n9851) );
  OAI21_X1 U9146 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(P1_ADDR_REG_15__SCAN_IN), 
        .A(n9851), .ZN(n9849) );
  NAND2_X1 U9147 ( .A1(n9850), .A2(n9849), .ZN(n9848) );
  OAI21_X1 U9148 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(P2_ADDR_REG_16__SCAN_IN), 
        .A(n9848), .ZN(n9846) );
  NAND2_X1 U9149 ( .A1(n9847), .A2(n9846), .ZN(n9845) );
  OAI21_X1 U9150 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(P1_ADDR_REG_17__SCAN_IN), 
        .A(n9845), .ZN(n10030) );
  NOR2_X1 U9151 ( .A1(n10031), .A2(n10030), .ZN(n7521) );
  NAND2_X1 U9152 ( .A1(n10031), .A2(n10030), .ZN(n10029) );
  OAI21_X1 U9153 ( .B1(P1_ADDR_REG_18__SCAN_IN), .B2(n7521), .A(n10029), .ZN(
        n7523) );
  XNOR2_X1 U9154 ( .A(n4866), .B(P1_ADDR_REG_19__SCAN_IN), .ZN(n7522) );
  XNOR2_X1 U9155 ( .A(n7523), .B(n7522), .ZN(ADD_1071_U4) );
  INV_X1 U9156 ( .A(n7995), .ZN(n7543) );
  OAI222_X1 U9157 ( .A1(P2_U3152), .A2(n7524), .B1(n4284), .B2(n7543), .C1(
        n9932), .C2(n7969), .ZN(P2_U3332) );
  INV_X1 U9158 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n7541) );
  INV_X1 U9159 ( .A(n7525), .ZN(n7527) );
  AOI21_X1 U9160 ( .B1(n7533), .B2(n7527), .A(n7526), .ZN(n7530) );
  NAND2_X1 U9161 ( .A1(n7728), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n7528) );
  OAI21_X1 U9162 ( .B1(n7728), .B2(P1_REG2_REG_16__SCAN_IN), .A(n7528), .ZN(
        n7529) );
  NOR2_X1 U9163 ( .A1(n7530), .A2(n7529), .ZN(n7727) );
  AOI211_X1 U9164 ( .C1(n7530), .C2(n7529), .A(n7727), .B(n9543), .ZN(n7531)
         );
  INV_X1 U9165 ( .A(n7531), .ZN(n7540) );
  NAND2_X1 U9166 ( .A1(P1_U3084), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n7850) );
  INV_X1 U9167 ( .A(n7850), .ZN(n7538) );
  AOI21_X1 U9168 ( .B1(n7534), .B2(n7533), .A(n7532), .ZN(n7536) );
  XNOR2_X1 U9169 ( .A(n7728), .B(P1_REG1_REG_16__SCAN_IN), .ZN(n7535) );
  NOR2_X1 U9170 ( .A1(n7536), .A2(n7535), .ZN(n7724) );
  AOI211_X1 U9171 ( .C1(n7536), .C2(n7535), .A(n7724), .B(n9522), .ZN(n7537)
         );
  AOI211_X1 U9172 ( .C1(n7728), .C2(n9553), .A(n7538), .B(n7537), .ZN(n7539)
         );
  OAI211_X1 U9173 ( .C1(n9571), .C2(n7541), .A(n7540), .B(n7539), .ZN(P1_U3257) );
  OAI222_X1 U9174 ( .A1(n8073), .A2(n7543), .B1(P1_U3084), .B2(n6235), .C1(
        n7542), .C2(n8069), .ZN(P1_U3327) );
  INV_X1 U9175 ( .A(n8010), .ZN(n7968) );
  AOI21_X1 U9176 ( .B1(n9369), .B2(P2_DATAO_REG_27__SCAN_IN), .A(n7544), .ZN(
        n7545) );
  OAI21_X1 U9177 ( .B1(n7968), .B2(n8073), .A(n7545), .ZN(P1_U3326) );
  INV_X1 U9178 ( .A(n7546), .ZN(n7547) );
  NAND2_X1 U9179 ( .A1(n7548), .A2(n7547), .ZN(n7549) );
  NAND2_X1 U9180 ( .A1(n7694), .A2(n7933), .ZN(n7552) );
  OR2_X1 U9181 ( .A1(n9425), .A2(n6359), .ZN(n7551) );
  NAND2_X1 U9182 ( .A1(n7552), .A2(n7551), .ZN(n7553) );
  XNOR2_X1 U9183 ( .A(n7553), .B(n7936), .ZN(n7555) );
  NOR2_X1 U9184 ( .A1(n9425), .A2(n7942), .ZN(n7554) );
  AOI21_X1 U9185 ( .B1(n7694), .B2(n7939), .A(n7554), .ZN(n7556) );
  NAND2_X1 U9186 ( .A1(n7555), .A2(n7556), .ZN(n7634) );
  INV_X1 U9187 ( .A(n7555), .ZN(n7558) );
  INV_X1 U9188 ( .A(n7556), .ZN(n7557) );
  NAND2_X1 U9189 ( .A1(n7558), .A2(n7557), .ZN(n7635) );
  NAND2_X1 U9190 ( .A1(n9408), .A2(n7939), .ZN(n7560) );
  OR2_X1 U9191 ( .A1(n7697), .A2(n7942), .ZN(n7559) );
  NAND2_X1 U9192 ( .A1(n7560), .A2(n7559), .ZN(n7705) );
  NAND2_X1 U9193 ( .A1(n9408), .A2(n7933), .ZN(n7562) );
  OR2_X1 U9194 ( .A1(n7697), .A2(n6359), .ZN(n7561) );
  NAND2_X1 U9195 ( .A1(n7562), .A2(n7561), .ZN(n7563) );
  XNOR2_X1 U9196 ( .A(n7563), .B(n6860), .ZN(n7706) );
  XOR2_X1 U9197 ( .A(n7705), .B(n7706), .Z(n7564) );
  XNOR2_X1 U9198 ( .A(n7707), .B(n7564), .ZN(n7570) );
  INV_X1 U9199 ( .A(n9425), .ZN(n9001) );
  NOR2_X1 U9200 ( .A1(n8963), .A2(n9401), .ZN(n7565) );
  AOI211_X1 U9201 ( .C1(n8965), .C2(n9001), .A(n7566), .B(n7565), .ZN(n7567)
         );
  OAI21_X1 U9202 ( .B1(n9396), .B2(n8989), .A(n7567), .ZN(n7568) );
  AOI21_X1 U9203 ( .B1(n9408), .B2(n8968), .A(n7568), .ZN(n7569) );
  OAI21_X1 U9204 ( .B1(n7570), .B2(n8984), .A(n7569), .ZN(P1_U3232) );
  OR2_X1 U9205 ( .A1(n7571), .A2(n9003), .ZN(n7572) );
  NAND2_X1 U9206 ( .A1(n7576), .A2(n7584), .ZN(n7696) );
  OR2_X1 U9207 ( .A1(n7576), .A2(n7584), .ZN(n7577) );
  AND2_X1 U9208 ( .A1(n7696), .A2(n7577), .ZN(n9454) );
  NAND2_X1 U9209 ( .A1(n9422), .A2(n7582), .ZN(n7687) );
  NAND2_X1 U9210 ( .A1(n7687), .A2(n7583), .ZN(n7585) );
  XNOR2_X1 U9211 ( .A(n7585), .B(n7584), .ZN(n7586) );
  NAND2_X1 U9212 ( .A1(n7586), .A2(n9427), .ZN(n7588) );
  INV_X1 U9213 ( .A(n7697), .ZN(n9000) );
  AOI22_X1 U9214 ( .A1(n9000), .A2(n9261), .B1(n9586), .B2(n9002), .ZN(n7587)
         );
  NAND2_X1 U9215 ( .A1(n7588), .A2(n7587), .ZN(n7589) );
  AOI21_X1 U9216 ( .B1(n9454), .B2(n9420), .A(n7589), .ZN(n9456) );
  INV_X1 U9217 ( .A(n7694), .ZN(n7590) );
  OAI21_X1 U9218 ( .B1(n9414), .B2(n7590), .A(n9572), .ZN(n7591) );
  OR2_X1 U9219 ( .A1(n7591), .A2(n9392), .ZN(n9452) );
  INV_X1 U9220 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n7592) );
  OAI22_X1 U9221 ( .A1(n9600), .A2(n7592), .B1(n7641), .B2(n9418), .ZN(n7593)
         );
  AOI21_X1 U9222 ( .B1(n7694), .B2(n9434), .A(n7593), .ZN(n7594) );
  OAI21_X1 U9223 ( .B1(n9452), .B2(n7700), .A(n7594), .ZN(n7595) );
  AOI21_X1 U9224 ( .B1(n9454), .B2(n9597), .A(n7595), .ZN(n7596) );
  OAI21_X1 U9225 ( .B1(n9456), .B2(n4283), .A(n7596), .ZN(P1_U3279) );
  INV_X1 U9226 ( .A(n8519), .ZN(n8255) );
  XNOR2_X1 U9227 ( .A(n8843), .B(n8519), .ZN(n8253) );
  AND2_X1 U9228 ( .A1(n8253), .A2(n8250), .ZN(n7597) );
  OR2_X1 U9229 ( .A1(n8843), .A2(n8255), .ZN(n8257) );
  NAND2_X1 U9230 ( .A1(n7647), .A2(n8050), .ZN(n8261) );
  NAND2_X1 U9231 ( .A1(n8262), .A2(n8261), .ZN(n8358) );
  INV_X1 U9232 ( .A(n8358), .ZN(n8259) );
  XNOR2_X1 U9233 ( .A(n7655), .B(n8259), .ZN(n7598) );
  OAI222_X1 U9234 ( .A1(n8721), .A2(n7745), .B1(n8719), .B2(n8255), .C1(n8698), 
        .C2(n7598), .ZN(n8839) );
  INV_X1 U9235 ( .A(n8839), .ZN(n7609) );
  INV_X1 U9236 ( .A(n7679), .ZN(n8520) );
  NAND2_X1 U9237 ( .A1(n7599), .A2(n8520), .ZN(n7600) );
  OR2_X1 U9238 ( .A1(n8843), .A2(n8519), .ZN(n7648) );
  NAND2_X1 U9239 ( .A1(n7650), .A2(n7648), .ZN(n7603) );
  NAND2_X1 U9240 ( .A1(n7603), .A2(n8358), .ZN(n7602) );
  OAI21_X1 U9241 ( .B1(n7603), .B2(n8358), .A(n7602), .ZN(n8841) );
  AND2_X1 U9242 ( .A1(n7673), .A2(n7647), .ZN(n7604) );
  OR2_X1 U9243 ( .A1(n7604), .A2(n7660), .ZN(n8838) );
  AOI22_X1 U9244 ( .A1(n9772), .A2(P2_REG2_REG_15__SCAN_IN), .B1(n7778), .B2(
        n9760), .ZN(n7606) );
  NAND2_X1 U9245 ( .A1(n7647), .A2(n8736), .ZN(n7605) );
  OAI211_X1 U9246 ( .C1(n8838), .C2(n8708), .A(n7606), .B(n7605), .ZN(n7607)
         );
  AOI21_X1 U9247 ( .B1(n8841), .B2(n9765), .A(n7607), .ZN(n7608) );
  OAI21_X1 U9248 ( .B1(n7609), .B2(n9772), .A(n7608), .ZN(P2_U3281) );
  XNOR2_X1 U9249 ( .A(n7622), .B(P2_REG2_REG_17__SCAN_IN), .ZN(n9743) );
  INV_X1 U9250 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n7612) );
  NOR2_X1 U9251 ( .A1(n7622), .A2(n7612), .ZN(n7613) );
  OAI21_X1 U9252 ( .B1(n7616), .B2(n7615), .A(n7614), .ZN(n7617) );
  NOR2_X1 U9253 ( .A1(P2_REG2_REG_18__SCAN_IN), .A2(n7617), .ZN(n8058) );
  AOI21_X1 U9254 ( .B1(n7617), .B2(P2_REG2_REG_18__SCAN_IN), .A(n8058), .ZN(
        n7632) );
  OR2_X1 U9255 ( .A1(n7629), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n8060) );
  NAND2_X1 U9256 ( .A1(n7629), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n7618) );
  AND2_X1 U9257 ( .A1(n8060), .A2(n7618), .ZN(n7625) );
  INV_X1 U9258 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n7621) );
  AOI21_X1 U9259 ( .B1(n9977), .B2(n7620), .A(n7619), .ZN(n9751) );
  XNOR2_X1 U9260 ( .A(n7622), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n9750) );
  NAND2_X1 U9261 ( .A1(n9751), .A2(n9750), .ZN(n9749) );
  OAI21_X1 U9262 ( .B1(n7622), .B2(n7621), .A(n9749), .ZN(n7623) );
  INV_X1 U9263 ( .A(n7623), .ZN(n7624) );
  NAND2_X1 U9264 ( .A1(n7625), .A2(n7624), .ZN(n8061) );
  OAI21_X1 U9265 ( .B1(n7625), .B2(n7624), .A(n8061), .ZN(n7628) );
  NOR2_X1 U9266 ( .A1(n7626), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8490) );
  NOR2_X1 U9267 ( .A1(n8068), .A2(n10031), .ZN(n7627) );
  AOI211_X1 U9268 ( .C1(n9748), .C2(n7628), .A(n8490), .B(n7627), .ZN(n7631)
         );
  NAND2_X1 U9269 ( .A1(n9747), .A2(n7629), .ZN(n7630) );
  OAI211_X1 U9270 ( .C1(n7632), .C2(n9692), .A(n7631), .B(n7630), .ZN(P2_U3263) );
  NAND2_X1 U9271 ( .A1(n7694), .A2(n9345), .ZN(n9451) );
  INV_X1 U9272 ( .A(n7635), .ZN(n7639) );
  AOI21_X1 U9273 ( .B1(n7635), .B2(n7634), .A(n7633), .ZN(n7636) );
  NOR2_X1 U9274 ( .A1(n7636), .A2(n8984), .ZN(n7637) );
  OAI21_X1 U9275 ( .B1(n7639), .B2(n7638), .A(n7637), .ZN(n7645) );
  OAI21_X1 U9276 ( .B1(n8963), .B2(n7697), .A(n7640), .ZN(n7643) );
  NOR2_X1 U9277 ( .A1(n8989), .A2(n7641), .ZN(n7642) );
  AOI211_X1 U9278 ( .C1(n8965), .C2(n9002), .A(n7643), .B(n7642), .ZN(n7644)
         );
  OAI211_X1 U9279 ( .C1(n9451), .C2(n7646), .A(n7645), .B(n7644), .ZN(P1_U3222) );
  INV_X1 U9280 ( .A(n7647), .ZN(n8837) );
  NAND2_X1 U9281 ( .A1(n8837), .A2(n8050), .ZN(n7651) );
  AND2_X1 U9282 ( .A1(n7648), .A2(n7651), .ZN(n7649) );
  INV_X1 U9283 ( .A(n7651), .ZN(n7652) );
  OR2_X1 U9284 ( .A1(n7652), .A2(n8358), .ZN(n7746) );
  NAND2_X1 U9285 ( .A1(n7748), .A2(n7746), .ZN(n7654) );
  OR2_X1 U9286 ( .A1(n7791), .A2(n7745), .ZN(n8268) );
  NAND2_X1 U9287 ( .A1(n7791), .A2(n7745), .ZN(n8267) );
  NAND2_X1 U9288 ( .A1(n8268), .A2(n8267), .ZN(n8360) );
  NAND2_X1 U9289 ( .A1(n7654), .A2(n8360), .ZN(n7653) );
  OAI21_X1 U9290 ( .B1(n7654), .B2(n8360), .A(n7653), .ZN(n7738) );
  OR2_X1 U9291 ( .A1(n7738), .A2(n8729), .ZN(n7659) );
  XNOR2_X1 U9292 ( .A(n7754), .B(n8360), .ZN(n7657) );
  OAI22_X1 U9293 ( .A1(n8494), .A2(n8721), .B1(n8050), .B2(n8719), .ZN(n7656)
         );
  AOI21_X1 U9294 ( .B1(n7657), .B2(n9759), .A(n7656), .ZN(n7658) );
  NAND2_X1 U9295 ( .A1(n7659), .A2(n7658), .ZN(n7740) );
  INV_X1 U9296 ( .A(n7740), .ZN(n7669) );
  INV_X1 U9297 ( .A(n7738), .ZN(n7667) );
  INV_X1 U9298 ( .A(n7791), .ZN(n7734) );
  NOR2_X1 U9299 ( .A1(n7660), .A2(n7734), .ZN(n7661) );
  OR2_X1 U9300 ( .A1(n7761), .A2(n7661), .ZN(n7735) );
  INV_X1 U9301 ( .A(n7662), .ZN(n7786) );
  OAI22_X1 U9302 ( .A1(n8734), .A2(n7155), .B1(n7786), .B2(n8731), .ZN(n7663)
         );
  AOI21_X1 U9303 ( .B1(n7791), .B2(n8736), .A(n7663), .ZN(n7664) );
  OAI21_X1 U9304 ( .B1(n7735), .B2(n8708), .A(n7664), .ZN(n7665) );
  AOI21_X1 U9305 ( .B1(n7667), .B2(n7666), .A(n7665), .ZN(n7668) );
  OAI21_X1 U9306 ( .B1(n7669), .B2(n9772), .A(n7668), .ZN(P2_U3280) );
  INV_X1 U9307 ( .A(n8023), .ZN(n7967) );
  NAND2_X1 U9308 ( .A1(n8877), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n7670) );
  OAI211_X1 U9309 ( .C1(n7967), .C2(n4284), .A(n7671), .B(n7670), .ZN(P2_U3330) );
  INV_X1 U9310 ( .A(n8253), .ZN(n8359) );
  XNOR2_X1 U9311 ( .A(n7672), .B(n8359), .ZN(n8847) );
  INV_X1 U9312 ( .A(n7673), .ZN(n7674) );
  AOI21_X1 U9313 ( .B1(n8843), .B2(n7675), .A(n7674), .ZN(n8844) );
  AOI22_X1 U9314 ( .A1(n9772), .A2(P2_REG2_REG_14__SCAN_IN), .B1(n8053), .B2(
        n9760), .ZN(n7676) );
  OAI21_X1 U9315 ( .B1(n4491), .B2(n9768), .A(n7676), .ZN(n7684) );
  NAND2_X1 U9316 ( .A1(n7677), .A2(n8250), .ZN(n7678) );
  AOI21_X1 U9317 ( .B1(n7678), .B2(n8359), .A(n8698), .ZN(n7682) );
  OAI22_X1 U9318 ( .A1(n8050), .A2(n8721), .B1(n7679), .B2(n8719), .ZN(n7680)
         );
  AOI21_X1 U9319 ( .B1(n7682), .B2(n7681), .A(n7680), .ZN(n8846) );
  NOR2_X1 U9320 ( .A1(n8846), .A2(n9772), .ZN(n7683) );
  AOI211_X1 U9321 ( .C1(n8844), .C2(n9762), .A(n7684), .B(n7683), .ZN(n7685)
         );
  OAI21_X1 U9322 ( .B1(n8847), .B2(n8761), .A(n7685), .ZN(P2_U3282) );
  NAND2_X1 U9323 ( .A1(n7687), .A2(n7686), .ZN(n7689) );
  NAND2_X1 U9324 ( .A1(n7689), .A2(n7688), .ZN(n9399) );
  NAND2_X1 U9325 ( .A1(n9398), .A2(n7797), .ZN(n7690) );
  INV_X1 U9326 ( .A(n7795), .ZN(n7798) );
  XNOR2_X1 U9327 ( .A(n7690), .B(n7798), .ZN(n7693) );
  NAND2_X1 U9328 ( .A1(n9260), .A2(n9261), .ZN(n7691) );
  OAI21_X1 U9329 ( .B1(n7697), .B2(n9423), .A(n7691), .ZN(n7692) );
  AOI21_X1 U9330 ( .B1(n7693), .B2(n9427), .A(n7692), .ZN(n9443) );
  NAND2_X1 U9331 ( .A1(n7694), .A2(n9001), .ZN(n7695) );
  XNOR2_X1 U9332 ( .A(n7796), .B(n7795), .ZN(n9445) );
  NAND2_X1 U9333 ( .A1(n9445), .A2(n9597), .ZN(n7704) );
  OAI22_X1 U9334 ( .A1(n9600), .A2(n7698), .B1(n7717), .B2(n9418), .ZN(n7702)
         );
  INV_X1 U9335 ( .A(n9394), .ZN(n7699) );
  OAI211_X1 U9336 ( .C1(n7699), .C2(n4466), .A(n9572), .B(n7802), .ZN(n9442)
         );
  NOR2_X1 U9337 ( .A1(n9442), .A2(n7700), .ZN(n7701) );
  AOI211_X1 U9338 ( .C1(n9434), .C2(n7719), .A(n7702), .B(n7701), .ZN(n7703)
         );
  OAI211_X1 U9339 ( .C1(n4283), .C2(n9443), .A(n7704), .B(n7703), .ZN(P1_U3277) );
  NAND2_X1 U9340 ( .A1(n7719), .A2(n7933), .ZN(n7709) );
  OR2_X1 U9341 ( .A1(n9401), .A2(n6359), .ZN(n7708) );
  NAND2_X1 U9342 ( .A1(n7709), .A2(n7708), .ZN(n7710) );
  XNOR2_X1 U9343 ( .A(n7710), .B(n7936), .ZN(n7834) );
  NAND2_X1 U9344 ( .A1(n7719), .A2(n7939), .ZN(n7712) );
  OR2_X1 U9345 ( .A1(n9401), .A2(n7942), .ZN(n7711) );
  NAND2_X1 U9346 ( .A1(n7712), .A2(n7711), .ZN(n7823) );
  XNOR2_X1 U9347 ( .A(n7834), .B(n7823), .ZN(n7713) );
  XNOR2_X1 U9348 ( .A(n7822), .B(n7713), .ZN(n7721) );
  OAI21_X1 U9349 ( .B1(n8963), .B2(n8077), .A(n7714), .ZN(n7715) );
  AOI21_X1 U9350 ( .B1(n8965), .B2(n9000), .A(n7715), .ZN(n7716) );
  OAI21_X1 U9351 ( .B1(n7717), .B2(n8989), .A(n7716), .ZN(n7718) );
  AOI21_X1 U9352 ( .B1(n7719), .B2(n8968), .A(n7718), .ZN(n7720) );
  OAI21_X1 U9353 ( .B1(n7721), .B2(n8984), .A(n7720), .ZN(P1_U3213) );
  INV_X1 U9354 ( .A(n9039), .ZN(n7723) );
  NAND2_X1 U9355 ( .A1(P1_U3084), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n8927) );
  NAND2_X1 U9356 ( .A1(n9508), .A2(P1_ADDR_REG_17__SCAN_IN), .ZN(n7722) );
  OAI211_X1 U9357 ( .C1(n9538), .C2(n7723), .A(n8927), .B(n7722), .ZN(n7733)
         );
  AOI21_X1 U9358 ( .B1(n7728), .B2(P1_REG1_REG_16__SCAN_IN), .A(n7724), .ZN(
        n7726) );
  XNOR2_X1 U9359 ( .A(n9039), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n7725) );
  NOR2_X1 U9360 ( .A1(n7726), .A2(n7725), .ZN(n9035) );
  AOI211_X1 U9361 ( .C1(n7726), .C2(n7725), .A(n9035), .B(n9522), .ZN(n7732)
         );
  XNOR2_X1 U9362 ( .A(n9039), .B(P1_REG2_REG_17__SCAN_IN), .ZN(n7729) );
  AOI211_X1 U9363 ( .C1(n7730), .C2(n7729), .A(n9038), .B(n9543), .ZN(n7731)
         );
  OR3_X1 U9364 ( .A1(n7733), .A2(n7732), .A3(n7731), .ZN(P1_U3258) );
  OAI22_X1 U9365 ( .A1(n7735), .A2(n4275), .B1(n7734), .B2(n9819), .ZN(n7736)
         );
  INV_X1 U9366 ( .A(n7736), .ZN(n7737) );
  OAI21_X1 U9367 ( .B1(n7738), .B2(n9381), .A(n7737), .ZN(n7739) );
  NOR2_X1 U9368 ( .A1(n7740), .A2(n7739), .ZN(n7742) );
  MUX2_X1 U9369 ( .A(n9977), .B(n7742), .S(n9836), .Z(n7741) );
  INV_X1 U9370 ( .A(n7741), .ZN(P2_U3536) );
  INV_X1 U9371 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n7743) );
  MUX2_X1 U9372 ( .A(n7743), .B(n7742), .S(n9828), .Z(n7744) );
  INV_X1 U9373 ( .A(n7744), .ZN(P2_U3499) );
  INV_X1 U9374 ( .A(n7745), .ZN(n8518) );
  NAND2_X1 U9375 ( .A1(n7791), .A2(n8518), .ZN(n7749) );
  AND2_X1 U9376 ( .A1(n7746), .A2(n7749), .ZN(n7747) );
  INV_X1 U9377 ( .A(n7749), .ZN(n7750) );
  OR2_X1 U9378 ( .A1(n7750), .A2(n8360), .ZN(n7751) );
  XNOR2_X1 U9379 ( .A(n8834), .B(n8494), .ZN(n7756) );
  OAI21_X1 U9380 ( .B1(n7752), .B2(n7756), .A(n8387), .ZN(n7753) );
  INV_X1 U9381 ( .A(n7753), .ZN(n8836) );
  AOI22_X1 U9382 ( .A1(n8834), .A2(n8736), .B1(n9772), .B2(
        P2_REG2_REG_17__SCAN_IN), .ZN(n7768) );
  INV_X1 U9383 ( .A(n7754), .ZN(n7755) );
  NAND2_X1 U9384 ( .A1(n7755), .A2(n8265), .ZN(n7758) );
  AND2_X1 U9385 ( .A1(n7758), .A2(n8267), .ZN(n7759) );
  INV_X1 U9386 ( .A(n7756), .ZN(n8361) );
  AND2_X1 U9387 ( .A1(n8361), .A2(n8267), .ZN(n7757) );
  NAND2_X1 U9388 ( .A1(n7758), .A2(n7757), .ZN(n8747) );
  OAI211_X1 U9389 ( .C1(n7759), .C2(n8361), .A(n8747), .B(n9759), .ZN(n7760)
         );
  AOI22_X1 U9390 ( .A1(n8755), .A2(n8517), .B1(n8518), .B2(n8753), .ZN(n7816)
         );
  NAND2_X1 U9391 ( .A1(n7760), .A2(n7816), .ZN(n8832) );
  INV_X1 U9392 ( .A(n7761), .ZN(n7763) );
  INV_X1 U9393 ( .A(n8834), .ZN(n7821) );
  NAND2_X1 U9394 ( .A1(n7761), .A2(n7821), .ZN(n8743) );
  AOI211_X1 U9395 ( .C1(n8834), .C2(n7763), .A(n4275), .B(n7762), .ZN(n8833)
         );
  INV_X1 U9396 ( .A(n8833), .ZN(n7765) );
  OAI22_X1 U9397 ( .A1(n7765), .A2(n4282), .B1(n8731), .B2(n7815), .ZN(n7766)
         );
  OAI21_X1 U9398 ( .B1(n8832), .B2(n7766), .A(n8734), .ZN(n7767) );
  OAI211_X1 U9399 ( .C1(n8836), .C2(n8761), .A(n7768), .B(n7767), .ZN(P2_U3279) );
  INV_X1 U9400 ( .A(n7771), .ZN(n7775) );
  AOI21_X1 U9401 ( .B1(n7771), .B2(n7770), .A(n7769), .ZN(n7772) );
  NOR2_X1 U9402 ( .A1(n7772), .A2(n8511), .ZN(n7773) );
  OAI21_X1 U9403 ( .B1(n7775), .B2(n7774), .A(n7773), .ZN(n7780) );
  AOI22_X1 U9404 ( .A1(n8491), .A2(n8518), .B1(P2_REG3_REG_15__SCAN_IN), .B2(
        P2_U3152), .ZN(n7776) );
  OAI21_X1 U9405 ( .B1(n8255), .B2(n8493), .A(n7776), .ZN(n7777) );
  AOI21_X1 U9406 ( .B1(n7778), .B2(n8496), .A(n7777), .ZN(n7779) );
  OAI211_X1 U9407 ( .C1(n8837), .C2(n8499), .A(n7780), .B(n7779), .ZN(P2_U3243) );
  INV_X1 U9408 ( .A(n8142), .ZN(n8072) );
  INV_X1 U9409 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n9975) );
  OAI222_X1 U9410 ( .A1(n7781), .A2(P2_U3152), .B1(n4284), .B2(n8072), .C1(
        n9975), .C2(n7969), .ZN(P2_U3329) );
  INV_X1 U9411 ( .A(n7782), .ZN(n7783) );
  AOI21_X1 U9412 ( .B1(n7785), .B2(n7784), .A(n7783), .ZN(n7793) );
  NOR2_X1 U9413 ( .A1(n8506), .A2(n7786), .ZN(n7790) );
  INV_X1 U9414 ( .A(n8494), .ZN(n8754) );
  NAND2_X1 U9415 ( .A1(n8491), .A2(n8754), .ZN(n7787) );
  OAI211_X1 U9416 ( .C1(n8493), .C2(n8050), .A(n7788), .B(n7787), .ZN(n7789)
         );
  AOI211_X1 U9417 ( .C1(n7791), .C2(n8509), .A(n7790), .B(n7789), .ZN(n7792)
         );
  OAI21_X1 U9418 ( .B1(n7793), .B2(n8511), .A(n7792), .ZN(P2_U3228) );
  XNOR2_X1 U9419 ( .A(n8076), .B(n7800), .ZN(n9441) );
  INV_X1 U9420 ( .A(n9441), .ZN(n7810) );
  XNOR2_X1 U9421 ( .A(n8102), .B(n7800), .ZN(n7801) );
  OAI222_X1 U9422 ( .A1(n9576), .A2(n8079), .B1(n9423), .B2(n9401), .C1(n7801), 
        .C2(n9581), .ZN(n9440) );
  INV_X1 U9423 ( .A(n8074), .ZN(n9437) );
  INV_X1 U9424 ( .A(n7802), .ZN(n7803) );
  INV_X1 U9425 ( .A(n8129), .ZN(n9252) );
  OAI21_X1 U9426 ( .B1(n9437), .B2(n7803), .A(n9252), .ZN(n9438) );
  OAI22_X1 U9427 ( .A1(n9600), .A2(n7804), .B1(n8988), .B2(n9418), .ZN(n7805)
         );
  AOI21_X1 U9428 ( .B1(n8074), .B2(n9434), .A(n7805), .ZN(n7806) );
  OAI21_X1 U9429 ( .B1(n9438), .B2(n7807), .A(n7806), .ZN(n7808) );
  AOI21_X1 U9430 ( .B1(n9440), .B2(n9600), .A(n7808), .ZN(n7809) );
  OAI21_X1 U9431 ( .B1(n7810), .B2(n9268), .A(n7809), .ZN(P1_U3276) );
  AOI21_X1 U9432 ( .B1(n7812), .B2(n7811), .A(n8511), .ZN(n7814) );
  NAND2_X1 U9433 ( .A1(n7814), .A2(n7813), .ZN(n7820) );
  INV_X1 U9434 ( .A(n7815), .ZN(n7818) );
  NAND2_X1 U9435 ( .A1(P2_U3152), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n9739) );
  OAI21_X1 U9436 ( .B1(n7960), .B2(n7816), .A(n9739), .ZN(n7817) );
  AOI21_X1 U9437 ( .B1(n7818), .B2(n8496), .A(n7817), .ZN(n7819) );
  OAI211_X1 U9438 ( .C1(n7821), .C2(n8499), .A(n7820), .B(n7819), .ZN(P2_U3230) );
  INV_X1 U9439 ( .A(n9344), .ZN(n9257) );
  NAND2_X1 U9440 ( .A1(n7822), .A2(n7823), .ZN(n7839) );
  NAND2_X1 U9441 ( .A1(n7839), .A2(n7834), .ZN(n7829) );
  INV_X1 U9442 ( .A(n7823), .ZN(n7824) );
  NAND2_X1 U9443 ( .A1(n7825), .A2(n7824), .ZN(n7836) );
  NAND2_X1 U9444 ( .A1(n8074), .A2(n7933), .ZN(n7827) );
  NAND2_X1 U9445 ( .A1(n9260), .A2(n7939), .ZN(n7826) );
  NAND2_X1 U9446 ( .A1(n7827), .A2(n7826), .ZN(n7828) );
  XNOR2_X1 U9447 ( .A(n7828), .B(n6860), .ZN(n7837) );
  NAND3_X1 U9448 ( .A1(n7829), .A2(n7836), .A3(n7837), .ZN(n7846) );
  NAND2_X1 U9449 ( .A1(n9344), .A2(n7933), .ZN(n7831) );
  OR2_X1 U9450 ( .A1(n8079), .A2(n6359), .ZN(n7830) );
  NAND2_X1 U9451 ( .A1(n7831), .A2(n7830), .ZN(n7832) );
  XNOR2_X1 U9452 ( .A(n7832), .B(n6860), .ZN(n7857) );
  NOR2_X1 U9453 ( .A1(n8079), .A2(n7942), .ZN(n7833) );
  AOI21_X1 U9454 ( .B1(n9344), .B2(n7939), .A(n7833), .ZN(n7858) );
  XNOR2_X1 U9455 ( .A(n7857), .B(n7858), .ZN(n7847) );
  INV_X1 U9456 ( .A(n7834), .ZN(n7835) );
  NAND2_X1 U9457 ( .A1(n7836), .A2(n7835), .ZN(n7841) );
  INV_X1 U9458 ( .A(n7837), .ZN(n7838) );
  NAND2_X1 U9459 ( .A1(n8074), .A2(n7939), .ZN(n7843) );
  NAND2_X1 U9460 ( .A1(n9260), .A2(n7904), .ZN(n7842) );
  NAND2_X1 U9461 ( .A1(n7843), .A2(n7842), .ZN(n8982) );
  NAND2_X1 U9462 ( .A1(n8983), .A2(n8982), .ZN(n7845) );
  NAND2_X1 U9463 ( .A1(n7844), .A2(n7845), .ZN(n7861) );
  INV_X1 U9464 ( .A(n7861), .ZN(n7849) );
  AOI21_X1 U9465 ( .B1(n7845), .B2(n7846), .A(n7847), .ZN(n7848) );
  OAI21_X1 U9466 ( .B1(n7849), .B2(n7848), .A(n8973), .ZN(n7854) );
  NOR2_X1 U9467 ( .A1(n8989), .A2(n9253), .ZN(n7852) );
  OAI21_X1 U9468 ( .B1(n8991), .B2(n8077), .A(n7850), .ZN(n7851) );
  AOI211_X1 U9469 ( .C1(n8994), .C2(n9262), .A(n7852), .B(n7851), .ZN(n7853)
         );
  OAI211_X1 U9470 ( .C1(n9257), .C2(n8997), .A(n7854), .B(n7853), .ZN(P1_U3224) );
  INV_X1 U9471 ( .A(n8146), .ZN(n8880) );
  OAI222_X1 U9472 ( .A1(n8069), .A2(n7856), .B1(n9371), .B2(n8880), .C1(
        P1_U3084), .C2(n7855), .ZN(P1_U3323) );
  AOI22_X1 U9473 ( .A1(n9308), .A2(n7939), .B1(n7904), .B2(n9172), .ZN(n8893)
         );
  INV_X1 U9474 ( .A(n7857), .ZN(n7859) );
  NAND2_X1 U9475 ( .A1(n7859), .A2(n7858), .ZN(n7860) );
  NAND2_X1 U9476 ( .A1(n9339), .A2(n7933), .ZN(n7863) );
  NAND2_X1 U9477 ( .A1(n9262), .A2(n7939), .ZN(n7862) );
  NAND2_X1 U9478 ( .A1(n7863), .A2(n7862), .ZN(n7864) );
  XNOR2_X1 U9479 ( .A(n7864), .B(n6860), .ZN(n7870) );
  NAND2_X1 U9480 ( .A1(n9339), .A2(n7939), .ZN(n7866) );
  NAND2_X1 U9481 ( .A1(n9262), .A2(n7904), .ZN(n7865) );
  NAND2_X1 U9482 ( .A1(n7866), .A2(n7865), .ZN(n7871) );
  NAND2_X1 U9483 ( .A1(n7870), .A2(n7871), .ZN(n8924) );
  NAND2_X1 U9484 ( .A1(n9334), .A2(n7933), .ZN(n7868) );
  OR2_X1 U9485 ( .A1(n8928), .A2(n6359), .ZN(n7867) );
  NAND2_X1 U9486 ( .A1(n7868), .A2(n7867), .ZN(n7869) );
  XNOR2_X1 U9487 ( .A(n7869), .B(n7936), .ZN(n7877) );
  INV_X1 U9488 ( .A(n7877), .ZN(n7874) );
  INV_X1 U9489 ( .A(n7870), .ZN(n7873) );
  INV_X1 U9490 ( .A(n7871), .ZN(n7872) );
  NAND2_X1 U9491 ( .A1(n7873), .A2(n7872), .ZN(n8923) );
  AND2_X1 U9492 ( .A1(n7874), .A2(n8923), .ZN(n7875) );
  NOR2_X1 U9493 ( .A1(n8928), .A2(n7942), .ZN(n7876) );
  AOI21_X1 U9494 ( .B1(n9334), .B2(n7939), .A(n7876), .ZN(n8960) );
  NAND2_X1 U9495 ( .A1(n9329), .A2(n7933), .ZN(n7879) );
  NAND2_X1 U9496 ( .A1(n9228), .A2(n7939), .ZN(n7878) );
  NAND2_X1 U9497 ( .A1(n7879), .A2(n7878), .ZN(n7880) );
  XNOR2_X1 U9498 ( .A(n7880), .B(n6860), .ZN(n7882) );
  AND2_X1 U9499 ( .A1(n9228), .A2(n7904), .ZN(n7881) );
  AOI21_X1 U9500 ( .B1(n9329), .B2(n7939), .A(n7881), .ZN(n7883) );
  XNOR2_X1 U9501 ( .A(n7882), .B(n7883), .ZN(n8901) );
  INV_X1 U9502 ( .A(n7882), .ZN(n7884) );
  NAND2_X1 U9503 ( .A1(n7884), .A2(n7883), .ZN(n7885) );
  NAND2_X1 U9504 ( .A1(n9324), .A2(n7933), .ZN(n7888) );
  NAND2_X1 U9505 ( .A1(n9213), .A2(n7939), .ZN(n7887) );
  NAND2_X1 U9506 ( .A1(n7888), .A2(n7887), .ZN(n7889) );
  XNOR2_X1 U9507 ( .A(n7889), .B(n7936), .ZN(n8942) );
  AND2_X1 U9508 ( .A1(n9213), .A2(n7904), .ZN(n7890) );
  AOI21_X1 U9509 ( .B1(n9324), .B2(n7939), .A(n7890), .ZN(n8941) );
  AND2_X1 U9510 ( .A1(n8942), .A2(n8941), .ZN(n7894) );
  INV_X1 U9511 ( .A(n8942), .ZN(n7892) );
  INV_X1 U9512 ( .A(n8941), .ZN(n7891) );
  NAND2_X1 U9513 ( .A1(n7892), .A2(n7891), .ZN(n7893) );
  NAND2_X1 U9514 ( .A1(n9319), .A2(n7933), .ZN(n7896) );
  OR2_X1 U9515 ( .A1(n8087), .A2(n6359), .ZN(n7895) );
  NAND2_X1 U9516 ( .A1(n7896), .A2(n7895), .ZN(n7897) );
  XNOR2_X1 U9517 ( .A(n7897), .B(n6860), .ZN(n7900) );
  NAND2_X1 U9518 ( .A1(n9319), .A2(n7939), .ZN(n7899) );
  OR2_X1 U9519 ( .A1(n8087), .A2(n7942), .ZN(n7898) );
  NAND2_X1 U9520 ( .A1(n7899), .A2(n7898), .ZN(n7901) );
  INV_X1 U9521 ( .A(n7900), .ZN(n7903) );
  INV_X1 U9522 ( .A(n7901), .ZN(n7902) );
  AND2_X1 U9523 ( .A1(n9187), .A2(n7904), .ZN(n7905) );
  AOI21_X1 U9524 ( .B1(n9314), .B2(n7939), .A(n7905), .ZN(n7909) );
  NAND2_X1 U9525 ( .A1(n9314), .A2(n7933), .ZN(n7907) );
  NAND2_X1 U9526 ( .A1(n9187), .A2(n7939), .ZN(n7906) );
  NAND2_X1 U9527 ( .A1(n7907), .A2(n7906), .ZN(n7908) );
  XNOR2_X1 U9528 ( .A(n7908), .B(n7936), .ZN(n8951) );
  NAND2_X1 U9529 ( .A1(n9308), .A2(n7933), .ZN(n7911) );
  NAND2_X1 U9530 ( .A1(n9172), .A2(n7939), .ZN(n7910) );
  NAND2_X1 U9531 ( .A1(n7911), .A2(n7910), .ZN(n7912) );
  XNOR2_X1 U9532 ( .A(n7912), .B(n6860), .ZN(n7913) );
  NAND2_X1 U9533 ( .A1(n5402), .A2(n7933), .ZN(n7915) );
  NAND2_X1 U9534 ( .A1(n9155), .A2(n7939), .ZN(n7914) );
  NAND2_X1 U9535 ( .A1(n7915), .A2(n7914), .ZN(n7916) );
  XNOR2_X1 U9536 ( .A(n7916), .B(n6860), .ZN(n7919) );
  INV_X1 U9537 ( .A(n5402), .ZN(n8130) );
  OAI22_X1 U9538 ( .A1(n8130), .A2(n6359), .B1(n7917), .B2(n7942), .ZN(n7918)
         );
  XNOR2_X1 U9539 ( .A(n7919), .B(n7918), .ZN(n8935) );
  OAI22_X1 U9540 ( .A1(n9125), .A2(n6359), .B1(n8977), .B2(n7942), .ZN(n7924)
         );
  NAND2_X1 U9541 ( .A1(n9299), .A2(n7933), .ZN(n7921) );
  OR2_X1 U9542 ( .A1(n8977), .A2(n6359), .ZN(n7920) );
  NAND2_X1 U9543 ( .A1(n7921), .A2(n7920), .ZN(n7922) );
  XNOR2_X1 U9544 ( .A(n7922), .B(n6860), .ZN(n7923) );
  XOR2_X1 U9545 ( .A(n7924), .B(n7923), .Z(n8917) );
  INV_X1 U9546 ( .A(n7923), .ZN(n7926) );
  INV_X1 U9547 ( .A(n7924), .ZN(n7925) );
  OR2_X1 U9548 ( .A1(n8094), .A2(n7942), .ZN(n7927) );
  NAND2_X1 U9549 ( .A1(n7928), .A2(n7927), .ZN(n7931) );
  OAI22_X1 U9550 ( .A1(n9111), .A2(n6384), .B1(n8094), .B2(n6359), .ZN(n7929)
         );
  XNOR2_X1 U9551 ( .A(n7929), .B(n6860), .ZN(n7930) );
  XOR2_X1 U9552 ( .A(n7931), .B(n7930), .Z(n8974) );
  NAND2_X1 U9553 ( .A1(n9289), .A2(n7933), .ZN(n7935) );
  OR2_X1 U9554 ( .A1(n10020), .A2(n6359), .ZN(n7934) );
  NAND2_X1 U9555 ( .A1(n7935), .A2(n7934), .ZN(n7937) );
  XNOR2_X1 U9556 ( .A(n7937), .B(n7936), .ZN(n7941) );
  NOR2_X1 U9557 ( .A1(n10020), .A2(n7942), .ZN(n7938) );
  AOI21_X1 U9558 ( .B1(n9289), .B2(n7939), .A(n7938), .ZN(n7940) );
  NOR2_X1 U9559 ( .A1(n7941), .A2(n7940), .ZN(n8883) );
  NAND2_X1 U9560 ( .A1(n7941), .A2(n7940), .ZN(n8882) );
  INV_X1 U9561 ( .A(n9284), .ZN(n9081) );
  OAI22_X1 U9562 ( .A1(n9081), .A2(n6359), .B1(n8999), .B2(n7942), .ZN(n7943)
         );
  XNOR2_X1 U9563 ( .A(n7943), .B(n6860), .ZN(n7945) );
  OAI22_X1 U9564 ( .A1(n9081), .A2(n6384), .B1(n8999), .B2(n6359), .ZN(n7944)
         );
  NOR2_X1 U9565 ( .A1(n8989), .A2(n9078), .ZN(n7949) );
  INV_X1 U9566 ( .A(n10020), .ZN(n9114) );
  AOI22_X1 U9567 ( .A1(n8965), .A2(n9114), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3084), .ZN(n7946) );
  OAI21_X1 U9568 ( .B1(n7947), .B2(n8963), .A(n7946), .ZN(n7948) );
  AOI211_X1 U9569 ( .C1(n9284), .C2(n8968), .A(n7949), .B(n7948), .ZN(n7950)
         );
  OAI222_X1 U9570 ( .A1(n7969), .A2(n7954), .B1(n4284), .B2(n7953), .C1(
        P2_U3152), .C2(n7951), .ZN(P2_U3336) );
  OAI21_X1 U9571 ( .B1(n7957), .B2(n7956), .A(n7955), .ZN(n7958) );
  NAND2_X1 U9572 ( .A1(n7958), .A2(n8473), .ZN(n7964) );
  NAND2_X1 U9573 ( .A1(P2_U3152), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n9701) );
  OAI21_X1 U9574 ( .B1(n7960), .B2(n7959), .A(n9701), .ZN(n7961) );
  AOI21_X1 U9575 ( .B1(n7962), .B2(n8496), .A(n7961), .ZN(n7963) );
  OAI211_X1 U9576 ( .C1(n7965), .C2(n8499), .A(n7964), .B(n7963), .ZN(P2_U3241) );
  INV_X1 U9577 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n7966) );
  OAI222_X1 U9578 ( .A1(n8073), .A2(n7967), .B1(n5682), .B2(P1_U3084), .C1(
        n7966), .C2(n8069), .ZN(P1_U3325) );
  OAI222_X1 U9579 ( .A1(n7969), .A2(n10021), .B1(n4284), .B2(n7968), .C1(n8407), .C2(P2_U3152), .ZN(P2_U3331) );
  AOI22_X1 U9580 ( .A1(n8472), .A2(n6630), .B1(n8473), .B2(n5748), .ZN(n7971)
         );
  NOR2_X1 U9581 ( .A1(n7971), .A2(n7970), .ZN(n7978) );
  AOI22_X1 U9582 ( .A1(n8491), .A2(n8530), .B1(n8509), .B2(n7972), .ZN(n7974)
         );
  NAND2_X1 U9583 ( .A1(n8504), .A2(n6630), .ZN(n7973) );
  OAI211_X1 U9584 ( .C1(n7976), .C2(n7975), .A(n7974), .B(n7973), .ZN(n7977)
         );
  AOI21_X1 U9585 ( .B1(n7978), .B2(n6579), .A(n7977), .ZN(n7979) );
  OAI21_X1 U9586 ( .B1(n7980), .B2(n8511), .A(n7979), .ZN(P2_U3239) );
  NAND2_X1 U9587 ( .A1(n7983), .A2(n4813), .ZN(n7990) );
  OAI21_X1 U9588 ( .B1(n7986), .B2(n7985), .A(n7984), .ZN(n7989) );
  NAND3_X1 U9589 ( .A1(n7990), .A2(n7989), .A3(n4810), .ZN(n8454) );
  NAND2_X1 U9590 ( .A1(n7991), .A2(n6129), .ZN(n7993) );
  NAND2_X1 U9591 ( .A1(n8147), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n7992) );
  XNOR2_X1 U9592 ( .A(n8790), .B(n8035), .ZN(n8452) );
  NAND2_X1 U9593 ( .A1(n8614), .A2(n8165), .ZN(n7994) );
  NOR2_X1 U9594 ( .A1(n8452), .A2(n7994), .ZN(n8450) );
  NAND2_X1 U9595 ( .A1(n8452), .A2(n7994), .ZN(n8453) );
  NAND2_X1 U9596 ( .A1(n7995), .A2(n6129), .ZN(n7997) );
  NAND2_X1 U9597 ( .A1(n8147), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n7996) );
  XNOR2_X1 U9598 ( .A(n8785), .B(n8035), .ZN(n8008) );
  INV_X1 U9599 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n7998) );
  NAND2_X1 U9600 ( .A1(n7999), .A2(n7998), .ZN(n8000) );
  NAND2_X1 U9601 ( .A1(n8028), .A2(n8000), .ZN(n8620) );
  INV_X1 U9602 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n9974) );
  NAND2_X1 U9603 ( .A1(n5871), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n8003) );
  NAND2_X1 U9604 ( .A1(n5843), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n8002) );
  OAI211_X1 U9605 ( .C1(n8154), .C2(n9974), .A(n8003), .B(n8002), .ZN(n8004)
         );
  INV_X1 U9606 ( .A(n8004), .ZN(n8005) );
  NAND2_X1 U9607 ( .A1(n8604), .A2(n8165), .ZN(n8007) );
  XNOR2_X1 U9608 ( .A(n8008), .B(n8007), .ZN(n8500) );
  NAND2_X1 U9609 ( .A1(n8147), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n8011) );
  XNOR2_X1 U9610 ( .A(n8779), .B(n8035), .ZN(n8020) );
  XNOR2_X1 U9611 ( .A(n8028), .B(P2_REG3_REG_27__SCAN_IN), .ZN(n8599) );
  NAND2_X1 U9612 ( .A1(n8599), .A2(n8034), .ZN(n8019) );
  INV_X1 U9613 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n8016) );
  NAND2_X1 U9614 ( .A1(n8013), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n8015) );
  NAND2_X1 U9615 ( .A1(n5871), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n8014) );
  OAI211_X1 U9616 ( .C1(n6106), .C2(n8016), .A(n8015), .B(n8014), .ZN(n8017)
         );
  INV_X1 U9617 ( .A(n8017), .ZN(n8018) );
  NOR2_X1 U9618 ( .A1(n8503), .A2(n5876), .ZN(n8021) );
  XNOR2_X1 U9619 ( .A(n8020), .B(n8021), .ZN(n8413) );
  INV_X1 U9620 ( .A(n8020), .ZN(n8022) );
  NAND2_X1 U9621 ( .A1(n8023), .A2(n6129), .ZN(n8025) );
  NAND2_X1 U9622 ( .A1(n8147), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n8024) );
  OAI21_X1 U9623 ( .B1(n8028), .B2(n8027), .A(n8026), .ZN(n8030) );
  INV_X1 U9624 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n9929) );
  NAND2_X1 U9625 ( .A1(n5843), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n8032) );
  NAND2_X1 U9626 ( .A1(n5871), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n8031) );
  OAI211_X1 U9627 ( .C1(n9929), .C2(n8154), .A(n8032), .B(n8031), .ZN(n8033)
         );
  AOI21_X1 U9628 ( .B1(n8583), .B2(n8034), .A(n8033), .ZN(n8416) );
  INV_X1 U9629 ( .A(n8416), .ZN(n8603) );
  NAND2_X1 U9630 ( .A1(n8603), .A2(n8165), .ZN(n8036) );
  XNOR2_X1 U9631 ( .A(n8036), .B(n8035), .ZN(n8037) );
  XNOR2_X1 U9632 ( .A(n8775), .B(n8037), .ZN(n8038) );
  NAND2_X1 U9633 ( .A1(n8615), .A2(n8504), .ZN(n8040) );
  AOI22_X1 U9634 ( .A1(n8583), .A2(n8496), .B1(P2_REG3_REG_28__SCAN_IN), .B2(
        P2_U3152), .ZN(n8039) );
  OAI211_X1 U9635 ( .C1(n8588), .C2(n8502), .A(n8040), .B(n8039), .ZN(n8041)
         );
  AOI21_X1 U9636 ( .B1(n8775), .B2(n8509), .A(n8041), .ZN(n8042) );
  NAND3_X1 U9637 ( .A1(n8043), .A2(n8472), .A3(n8520), .ZN(n8044) );
  OAI21_X1 U9638 ( .B1(n7449), .B2(n8511), .A(n8044), .ZN(n8047) );
  INV_X1 U9639 ( .A(n8045), .ZN(n8046) );
  NAND2_X1 U9640 ( .A1(n8047), .A2(n8046), .ZN(n8055) );
  NAND2_X1 U9641 ( .A1(n8504), .A2(n8520), .ZN(n8049) );
  OAI211_X1 U9642 ( .C1(n8050), .C2(n8502), .A(n8049), .B(n8048), .ZN(n8052)
         );
  NOR2_X1 U9643 ( .A1(n4491), .A2(n8499), .ZN(n8051) );
  AOI211_X1 U9644 ( .C1(n8496), .C2(n8053), .A(n8052), .B(n8051), .ZN(n8054)
         );
  OAI211_X1 U9645 ( .C1(n8511), .C2(n8056), .A(n8055), .B(n8054), .ZN(P2_U3217) );
  NOR2_X1 U9646 ( .A1(n8058), .A2(n8057), .ZN(n8059) );
  XOR2_X1 U9647 ( .A(n8059), .B(P2_REG2_REG_19__SCAN_IN), .Z(n8065) );
  NAND2_X1 U9648 ( .A1(n8061), .A2(n8060), .ZN(n8063) );
  INV_X1 U9649 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n8062) );
  XNOR2_X1 U9650 ( .A(n8063), .B(n8062), .ZN(n8066) );
  INV_X1 U9651 ( .A(n8066), .ZN(n8064) );
  AOI22_X1 U9652 ( .A1(n8065), .A2(n9744), .B1(n8064), .B2(n9748), .ZN(n8067)
         );
  NAND2_X1 U9653 ( .A1(P2_U3152), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n8429) );
  INV_X1 U9654 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n8070) );
  OAI222_X1 U9655 ( .A1(n8073), .A2(n8072), .B1(n8071), .B2(P1_U3084), .C1(
        n8070), .C2(n8069), .ZN(P1_U3324) );
  NAND2_X1 U9656 ( .A1(n8076), .A2(n8075), .ZN(n8078) );
  NAND2_X1 U9657 ( .A1(n8078), .A2(n4815), .ZN(n9250) );
  INV_X1 U9658 ( .A(n8079), .ZN(n9243) );
  NOR2_X1 U9659 ( .A1(n9339), .A2(n9262), .ZN(n8082) );
  INV_X1 U9660 ( .A(n9339), .ZN(n9240) );
  OAI22_X1 U9661 ( .A1(n9233), .A2(n8082), .B1(n9240), .B2(n8081), .ZN(n9218)
         );
  INV_X1 U9662 ( .A(n8928), .ZN(n9244) );
  NAND2_X1 U9663 ( .A1(n9329), .A2(n9228), .ZN(n8085) );
  AOI21_X1 U9664 ( .B1(n9205), .B2(n8085), .A(n8084), .ZN(n9192) );
  OAI21_X1 U9665 ( .B1(n9213), .B2(n9324), .A(n9192), .ZN(n8086) );
  INV_X1 U9666 ( .A(n9324), .ZN(n9197) );
  INV_X1 U9667 ( .A(n8087), .ZN(n9200) );
  INV_X1 U9668 ( .A(n9314), .ZN(n9167) );
  NAND2_X1 U9669 ( .A1(n8091), .A2(n4814), .ZN(n9133) );
  NAND2_X1 U9670 ( .A1(n9111), .A2(n8094), .ZN(n8096) );
  INV_X1 U9671 ( .A(n9289), .ZN(n9099) );
  NAND2_X1 U9672 ( .A1(n9076), .A2(n9075), .ZN(n9074) );
  NAND2_X1 U9673 ( .A1(n9074), .A2(n4812), .ZN(n8099) );
  NAND2_X1 U9674 ( .A1(n9241), .A2(n8104), .ZN(n9225) );
  INV_X1 U9675 ( .A(n8105), .ZN(n8106) );
  NAND2_X1 U9676 ( .A1(n9186), .A2(n8111), .ZN(n9169) );
  NAND2_X1 U9677 ( .A1(n9101), .A2(n9092), .ZN(n9083) );
  AND2_X1 U9678 ( .A1(n8124), .A2(P1_B_REG_SCAN_IN), .ZN(n8125) );
  NOR2_X1 U9679 ( .A1(n9576), .A2(n8125), .ZN(n9065) );
  INV_X1 U9680 ( .A(n9065), .ZN(n8126) );
  INV_X1 U9681 ( .A(n9319), .ZN(n9184) );
  NAND2_X1 U9682 ( .A1(n9193), .A2(n9184), .ZN(n9178) );
  INV_X1 U9683 ( .A(n9077), .ZN(n8131) );
  INV_X1 U9684 ( .A(n9281), .ZN(n8135) );
  AOI211_X1 U9685 ( .C1(n9281), .C2(n8131), .A(n9660), .B(n9069), .ZN(n9280)
         );
  NAND2_X1 U9686 ( .A1(n9280), .A2(n9141), .ZN(n8132) );
  OAI211_X1 U9687 ( .C1(n8133), .C2(n9418), .A(n9282), .B(n8132), .ZN(n8137)
         );
  OAI22_X1 U9688 ( .A1(n8135), .A2(n9256), .B1(n8134), .B2(n9600), .ZN(n8136)
         );
  AOI21_X1 U9689 ( .B1(n8137), .B2(n9600), .A(n8136), .ZN(n8138) );
  OAI21_X1 U9690 ( .B1(n9283), .B2(n9268), .A(n8138), .ZN(P1_U3355) );
  INV_X1 U9691 ( .A(n8517), .ZN(n8720) );
  OR2_X1 U9692 ( .A1(n8827), .A2(n8720), .ZN(n8276) );
  NAND2_X1 U9693 ( .A1(n8827), .A2(n8720), .ZN(n8286) );
  NAND2_X1 U9694 ( .A1(n8276), .A2(n8286), .ZN(n8748) );
  NOR2_X1 U9695 ( .A1(n8834), .A2(n8494), .ZN(n8749) );
  NOR2_X1 U9696 ( .A1(n8748), .A2(n8749), .ZN(n8139) );
  NAND2_X1 U9697 ( .A1(n8747), .A2(n8139), .ZN(n8751) );
  NAND2_X1 U9698 ( .A1(n8751), .A2(n8286), .ZN(n8717) );
  OR2_X1 U9699 ( .A1(n8823), .A2(n8701), .ZN(n8288) );
  NAND2_X1 U9700 ( .A1(n8823), .A2(n8701), .ZN(n8695) );
  NAND2_X1 U9701 ( .A1(n8705), .A2(n8722), .ZN(n8290) );
  NAND2_X1 U9702 ( .A1(n8810), .A2(n8700), .ZN(n8295) );
  INV_X1 U9703 ( .A(n8295), .ZN(n8670) );
  NAND2_X1 U9704 ( .A1(n8806), .A2(n8686), .ZN(n8296) );
  INV_X1 U9705 ( .A(n8298), .ZN(n8140) );
  NOR2_X1 U9706 ( .A1(n8141), .A2(n8140), .ZN(n8661) );
  OR2_X1 U9707 ( .A1(n8799), .A2(n8674), .ZN(n8282) );
  NAND2_X1 U9708 ( .A1(n8799), .A2(n8674), .ZN(n8176) );
  NAND2_X1 U9709 ( .A1(n8661), .A2(n8662), .ZN(n8660) );
  NAND2_X1 U9710 ( .A1(n8660), .A2(n8176), .ZN(n8642) );
  XNOR2_X1 U9711 ( .A(n8796), .B(n8663), .ZN(n8392) );
  INV_X1 U9712 ( .A(n8392), .ZN(n8641) );
  NAND2_X1 U9713 ( .A1(n8790), .A2(n8644), .ZN(n8171) );
  NAND2_X1 U9714 ( .A1(n8785), .A2(n8459), .ZN(n8308) );
  INV_X1 U9715 ( .A(n8601), .ZN(n8310) );
  NOR2_X1 U9716 ( .A1(n8779), .A2(n8503), .ZN(n8313) );
  NAND2_X1 U9717 ( .A1(n8775), .A2(n8416), .ZN(n8320) );
  NAND2_X1 U9718 ( .A1(n8142), .A2(n6129), .ZN(n8144) );
  NAND2_X1 U9719 ( .A1(n8147), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n8143) );
  NAND2_X1 U9720 ( .A1(n8770), .A2(n8588), .ZN(n8327) );
  INV_X1 U9721 ( .A(n8402), .ZN(n8368) );
  NAND2_X1 U9722 ( .A1(n8404), .A2(n8327), .ZN(n8156) );
  NAND2_X1 U9723 ( .A1(n8146), .A2(n6129), .ZN(n8149) );
  NAND2_X1 U9724 ( .A1(n8147), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n8148) );
  NOR2_X1 U9725 ( .A1(n8571), .A2(n6626), .ZN(n8150) );
  INV_X1 U9726 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n8153) );
  NAND2_X1 U9727 ( .A1(n5843), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n8152) );
  NAND2_X1 U9728 ( .A1(n5871), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n8151) );
  OAI211_X1 U9729 ( .C1(n8154), .C2(n8153), .A(n8152), .B(n8151), .ZN(n8513)
         );
  INV_X1 U9730 ( .A(n8513), .ZN(n8161) );
  NOR2_X1 U9731 ( .A1(n8765), .A2(n8161), .ZN(n8170) );
  NAND2_X1 U9732 ( .A1(n8156), .A2(n8155), .ZN(n8157) );
  NAND2_X1 U9733 ( .A1(n8158), .A2(n8157), .ZN(n8163) );
  NAND2_X1 U9734 ( .A1(n8872), .A2(n6129), .ZN(n8160) );
  NAND2_X1 U9735 ( .A1(n5819), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(n8159) );
  NAND2_X1 U9736 ( .A1(n8765), .A2(n8161), .ZN(n8330) );
  NAND2_X1 U9737 ( .A1(n8331), .A2(n8330), .ZN(n8168) );
  NAND2_X1 U9738 ( .A1(n8762), .A2(n8162), .ZN(n8169) );
  XNOR2_X1 U9739 ( .A(n8164), .B(n4282), .ZN(n8379) );
  INV_X1 U9740 ( .A(n8168), .ZN(n8369) );
  INV_X1 U9741 ( .A(n8169), .ZN(n8334) );
  NOR2_X1 U9742 ( .A1(n8334), .A2(n8170), .ZN(n8370) );
  OR2_X1 U9743 ( .A1(n8179), .A2(n6626), .ZN(n8332) );
  MUX2_X1 U9744 ( .A(n8369), .B(n8370), .S(n8332), .Z(n8337) );
  INV_X1 U9745 ( .A(n8171), .ZN(n8172) );
  OR2_X1 U9746 ( .A1(n8613), .A2(n8172), .ZN(n8175) );
  NAND2_X1 U9747 ( .A1(n8307), .A2(n8173), .ZN(n8174) );
  INV_X1 U9748 ( .A(n8332), .ZN(n8325) );
  MUX2_X1 U9749 ( .A(n8175), .B(n8174), .S(n8325), .Z(n8312) );
  INV_X1 U9750 ( .A(n8176), .ZN(n8285) );
  AND2_X1 U9751 ( .A1(n8177), .A2(n5733), .ZN(n8181) );
  INV_X1 U9752 ( .A(n8181), .ZN(n8178) );
  NAND2_X1 U9753 ( .A1(n8178), .A2(n8332), .ZN(n8184) );
  INV_X1 U9754 ( .A(n8179), .ZN(n8180) );
  NAND3_X1 U9755 ( .A1(n8181), .A2(n8180), .A3(n8185), .ZN(n8182) );
  OAI21_X1 U9756 ( .B1(n8184), .B2(n8183), .A(n8182), .ZN(n8201) );
  NAND2_X1 U9757 ( .A1(n8185), .A2(n8199), .ZN(n8186) );
  OR2_X1 U9758 ( .A1(n8201), .A2(n8186), .ZN(n8188) );
  AND2_X1 U9759 ( .A1(n8198), .A2(n8332), .ZN(n8187) );
  NAND2_X1 U9760 ( .A1(n8188), .A2(n8187), .ZN(n8203) );
  NAND2_X1 U9761 ( .A1(n8191), .A2(n8189), .ZN(n8190) );
  AOI21_X1 U9762 ( .B1(n8203), .B2(n8341), .A(n8190), .ZN(n8195) );
  NAND2_X1 U9763 ( .A1(n8194), .A2(n8191), .ZN(n8193) );
  NAND2_X1 U9764 ( .A1(n8210), .A2(n8209), .ZN(n8192) );
  MUX2_X1 U9765 ( .A(n8193), .B(n8192), .S(n8332), .Z(n8213) );
  OAI211_X1 U9766 ( .C1(n8195), .C2(n8213), .A(n8215), .B(n8194), .ZN(n8196)
         );
  NAND2_X1 U9767 ( .A1(n8196), .A2(n8332), .ZN(n8206) );
  INV_X1 U9768 ( .A(n8213), .ZN(n8204) );
  NAND2_X1 U9769 ( .A1(n8198), .A2(n8197), .ZN(n8200) );
  OAI21_X1 U9770 ( .B1(n8201), .B2(n8200), .A(n8199), .ZN(n8202) );
  NAND4_X1 U9771 ( .A1(n8204), .A2(n8341), .A3(n8203), .A4(n8202), .ZN(n8205)
         );
  NAND2_X1 U9772 ( .A1(n8206), .A2(n8205), .ZN(n8207) );
  NAND2_X1 U9773 ( .A1(n8207), .A2(n8211), .ZN(n8218) );
  AND2_X1 U9774 ( .A1(n8209), .A2(n8208), .ZN(n8212) );
  OAI211_X1 U9775 ( .C1(n8213), .C2(n8212), .A(n8211), .B(n8210), .ZN(n8214)
         );
  NAND2_X1 U9776 ( .A1(n8214), .A2(n8325), .ZN(n8217) );
  OAI21_X1 U9777 ( .B1(n8215), .B2(n8332), .A(n7284), .ZN(n8216) );
  AOI21_X1 U9778 ( .B1(n8218), .B2(n8217), .A(n8216), .ZN(n8223) );
  AND2_X1 U9779 ( .A1(n8219), .A2(n8332), .ZN(n8221) );
  NOR2_X1 U9780 ( .A1(n8219), .A2(n8332), .ZN(n8220) );
  MUX2_X1 U9781 ( .A(n8221), .B(n8220), .S(n8526), .Z(n8222) );
  OR3_X1 U9782 ( .A1(n8223), .A2(n8222), .A3(n8345), .ZN(n8228) );
  MUX2_X1 U9783 ( .A(n8225), .B(n8224), .S(n8325), .Z(n8226) );
  AND2_X1 U9784 ( .A1(n8226), .A2(n8229), .ZN(n8227) );
  NAND2_X1 U9785 ( .A1(n8228), .A2(n8227), .ZN(n8238) );
  AND2_X1 U9786 ( .A1(n8235), .A2(n8229), .ZN(n8232) );
  INV_X1 U9787 ( .A(n8235), .ZN(n8230) );
  OAI211_X1 U9788 ( .C1(n8230), .C2(n8233), .A(n8242), .B(n8234), .ZN(n8231)
         );
  AOI21_X1 U9789 ( .B1(n8238), .B2(n8232), .A(n8231), .ZN(n8240) );
  AND2_X1 U9790 ( .A1(n8234), .A2(n8233), .ZN(n8237) );
  NAND2_X1 U9791 ( .A1(n8241), .A2(n8235), .ZN(n8236) );
  AOI21_X1 U9792 ( .B1(n8238), .B2(n8237), .A(n8236), .ZN(n8239) );
  MUX2_X1 U9793 ( .A(n8240), .B(n8239), .S(n8325), .Z(n8249) );
  NAND2_X1 U9794 ( .A1(n8246), .A2(n8241), .ZN(n8244) );
  NAND2_X1 U9795 ( .A1(n8245), .A2(n8242), .ZN(n8243) );
  MUX2_X1 U9796 ( .A(n8244), .B(n8243), .S(n8325), .Z(n8248) );
  MUX2_X1 U9797 ( .A(n8246), .B(n8245), .S(n8332), .Z(n8247) );
  OAI211_X1 U9798 ( .C1(n8249), .C2(n8248), .A(n8356), .B(n8247), .ZN(n8254)
         );
  MUX2_X1 U9799 ( .A(n8251), .B(n8250), .S(n8332), .Z(n8252) );
  NAND3_X1 U9800 ( .A1(n8254), .A2(n8253), .A3(n8252), .ZN(n8260) );
  NAND2_X1 U9801 ( .A1(n8843), .A2(n8255), .ZN(n8256) );
  MUX2_X1 U9802 ( .A(n8257), .B(n8256), .S(n8325), .Z(n8258) );
  NAND3_X1 U9803 ( .A1(n8260), .A2(n8259), .A3(n8258), .ZN(n8264) );
  MUX2_X1 U9804 ( .A(n8262), .B(n8261), .S(n8332), .Z(n8263) );
  NAND2_X1 U9805 ( .A1(n8264), .A2(n8263), .ZN(n8266) );
  INV_X1 U9806 ( .A(n8360), .ZN(n8265) );
  NAND2_X1 U9807 ( .A1(n8266), .A2(n8265), .ZN(n8270) );
  MUX2_X1 U9808 ( .A(n8268), .B(n8267), .S(n8332), .Z(n8269) );
  NAND3_X1 U9809 ( .A1(n8270), .A2(n8361), .A3(n8269), .ZN(n8275) );
  INV_X1 U9810 ( .A(n8749), .ZN(n8273) );
  NAND2_X1 U9811 ( .A1(n8834), .A2(n8494), .ZN(n8271) );
  AND2_X1 U9812 ( .A1(n8286), .A2(n8271), .ZN(n8272) );
  MUX2_X1 U9813 ( .A(n8273), .B(n8272), .S(n8325), .Z(n8274) );
  NAND3_X1 U9814 ( .A1(n8275), .A2(n8274), .A3(n8276), .ZN(n8287) );
  NAND2_X1 U9815 ( .A1(n8287), .A2(n8276), .ZN(n8277) );
  NAND2_X1 U9816 ( .A1(n8277), .A2(n8695), .ZN(n8278) );
  NAND3_X1 U9817 ( .A1(n8278), .A2(n8292), .A3(n8288), .ZN(n8279) );
  NAND3_X1 U9818 ( .A1(n8279), .A2(n8295), .A3(n8290), .ZN(n8280) );
  NAND3_X1 U9819 ( .A1(n8298), .A2(n8280), .A3(n8293), .ZN(n8281) );
  NAND2_X1 U9820 ( .A1(n8281), .A2(n8296), .ZN(n8283) );
  OAI21_X1 U9821 ( .B1(n8653), .B2(n8283), .A(n8282), .ZN(n8284) );
  MUX2_X1 U9822 ( .A(n8285), .B(n8284), .S(n8325), .Z(n8305) );
  NAND2_X1 U9823 ( .A1(n8287), .A2(n8286), .ZN(n8289) );
  NAND2_X1 U9824 ( .A1(n8289), .A2(n8288), .ZN(n8291) );
  NAND3_X1 U9825 ( .A1(n8291), .A2(n8290), .A3(n8695), .ZN(n8294) );
  NAND3_X1 U9826 ( .A1(n8294), .A2(n8293), .A3(n8292), .ZN(n8297) );
  NAND3_X1 U9827 ( .A1(n8297), .A2(n8296), .A3(n8295), .ZN(n8299) );
  NAND3_X1 U9828 ( .A1(n8299), .A2(n8298), .A3(n8332), .ZN(n8300) );
  OAI21_X1 U9829 ( .B1(n8653), .B2(n8300), .A(n8392), .ZN(n8304) );
  NAND2_X1 U9830 ( .A1(n8663), .A2(n8332), .ZN(n8302) );
  OR2_X1 U9831 ( .A1(n8663), .A2(n8332), .ZN(n8301) );
  MUX2_X1 U9832 ( .A(n8302), .B(n8301), .S(n8796), .Z(n8303) );
  OAI211_X1 U9833 ( .C1(n8305), .C2(n8304), .A(n8365), .B(n8303), .ZN(n8306)
         );
  INV_X1 U9834 ( .A(n8306), .ZN(n8311) );
  MUX2_X1 U9835 ( .A(n8308), .B(n8307), .S(n8332), .Z(n8309) );
  OAI211_X1 U9836 ( .C1(n8312), .C2(n8311), .A(n8310), .B(n8309), .ZN(n8318)
         );
  INV_X1 U9837 ( .A(n8313), .ZN(n8314) );
  NAND2_X1 U9838 ( .A1(n8314), .A2(n8401), .ZN(n8315) );
  NAND2_X1 U9839 ( .A1(n8315), .A2(n8325), .ZN(n8317) );
  INV_X1 U9840 ( .A(n8320), .ZN(n8316) );
  AOI21_X1 U9841 ( .B1(n8318), .B2(n8317), .A(n8316), .ZN(n8324) );
  NAND2_X1 U9842 ( .A1(n8779), .A2(n8503), .ZN(n8319) );
  AOI21_X1 U9843 ( .B1(n8320), .B2(n8319), .A(n8325), .ZN(n8323) );
  NOR2_X1 U9844 ( .A1(n8401), .A2(n8325), .ZN(n8321) );
  NOR2_X1 U9845 ( .A1(n8402), .A2(n8321), .ZN(n8322) );
  OAI21_X1 U9846 ( .B1(n8324), .B2(n8323), .A(n8322), .ZN(n8329) );
  MUX2_X1 U9847 ( .A(n8327), .B(n8326), .S(n8325), .Z(n8328) );
  NAND4_X1 U9848 ( .A1(n8155), .A2(n8330), .A3(n8329), .A4(n8328), .ZN(n8336)
         );
  INV_X1 U9849 ( .A(n8331), .ZN(n8333) );
  MUX2_X1 U9850 ( .A(n8334), .B(n8333), .S(n8332), .Z(n8335) );
  AOI21_X1 U9851 ( .B1(n8337), .B2(n8336), .A(n8335), .ZN(n8338) );
  INV_X1 U9852 ( .A(n8709), .ZN(n8696) );
  INV_X1 U9853 ( .A(n8748), .ZN(n8740) );
  NAND3_X1 U9854 ( .A1(n8341), .A2(n8373), .A3(n8340), .ZN(n8344) );
  NOR4_X1 U9855 ( .A1(n8344), .A2(n8343), .A3(n8342), .A4(n6635), .ZN(n8348)
         );
  INV_X1 U9856 ( .A(n8345), .ZN(n8347) );
  NAND4_X1 U9857 ( .A1(n8348), .A2(n8347), .A3(n7046), .A4(n8346), .ZN(n8351)
         );
  NOR4_X1 U9858 ( .A1(n8352), .A2(n8351), .A3(n8350), .A4(n8349), .ZN(n8353)
         );
  NAND4_X1 U9859 ( .A1(n8356), .A2(n8355), .A3(n8354), .A4(n8353), .ZN(n8357)
         );
  NOR4_X1 U9860 ( .A1(n8360), .A2(n8359), .A3(n8358), .A4(n8357), .ZN(n8362)
         );
  NAND4_X1 U9861 ( .A1(n8718), .A2(n8740), .A3(n8362), .A4(n8361), .ZN(n8363)
         );
  NOR4_X1 U9862 ( .A1(n8672), .A2(n8684), .A3(n8696), .A4(n8363), .ZN(n8364)
         );
  NAND4_X1 U9863 ( .A1(n8365), .A2(n8662), .A3(n8364), .A4(n8392), .ZN(n8366)
         );
  NOR4_X1 U9864 ( .A1(n8586), .A2(n8601), .A3(n8613), .A4(n8366), .ZN(n8367)
         );
  NAND4_X1 U9865 ( .A1(n8370), .A2(n8369), .A3(n8368), .A4(n8367), .ZN(n8371)
         );
  XNOR2_X1 U9866 ( .A(n8371), .B(n5730), .ZN(n8374) );
  OAI22_X1 U9867 ( .A1(n8374), .A2(n5733), .B1(n8373), .B2(n8372), .ZN(n8375)
         );
  AOI21_X1 U9868 ( .B1(n8379), .B2(n4806), .A(n8378), .ZN(n8386) );
  INV_X1 U9869 ( .A(n8407), .ZN(n8381) );
  NAND4_X1 U9870 ( .A1(n9774), .A2(n8381), .A3(n8380), .A4(n8753), .ZN(n8382)
         );
  OAI211_X1 U9871 ( .C1(n8383), .C2(n8385), .A(n8382), .B(P2_B_REG_SCAN_IN), 
        .ZN(n8384) );
  OAI21_X1 U9872 ( .B1(n8386), .B2(n8385), .A(n8384), .ZN(P2_U3244) );
  INV_X1 U9873 ( .A(n8799), .ZN(n8659) );
  INV_X1 U9874 ( .A(n8722), .ZN(n8516) );
  NAND2_X1 U9875 ( .A1(n8827), .A2(n8517), .ZN(n8389) );
  NOR2_X1 U9876 ( .A1(n8827), .A2(n8517), .ZN(n8388) );
  NOR2_X1 U9877 ( .A1(n8390), .A2(n8701), .ZN(n8391) );
  OAI22_X1 U9878 ( .A1(n8715), .A2(n8391), .B1(n8756), .B2(n8823), .ZN(n8710)
         );
  NAND2_X1 U9879 ( .A1(n8624), .A2(n8394), .ZN(n8610) );
  NAND2_X1 U9880 ( .A1(n8610), .A2(n8613), .ZN(n8609) );
  NAND2_X1 U9881 ( .A1(n8609), .A2(n8395), .ZN(n8596) );
  NAND2_X1 U9882 ( .A1(n8596), .A2(n8601), .ZN(n8595) );
  NAND2_X1 U9883 ( .A1(n4481), .A2(n8416), .ZN(n8397) );
  INV_X1 U9884 ( .A(n8770), .ZN(n8400) );
  AOI22_X1 U9885 ( .A1(n8398), .A2(n9760), .B1(P2_REG2_REG_29__SCAN_IN), .B2(
        n9772), .ZN(n8399) );
  OAI21_X1 U9886 ( .B1(n8400), .B2(n9768), .A(n8399), .ZN(n8411) );
  INV_X1 U9887 ( .A(n8401), .ZN(n8403) );
  NAND2_X1 U9888 ( .A1(n8405), .A2(n8404), .ZN(n8406) );
  NAND2_X1 U9889 ( .A1(n8406), .A2(n9759), .ZN(n8410) );
  NOR2_X1 U9890 ( .A1(n8407), .A2(n9966), .ZN(n8408) );
  NOR2_X1 U9891 ( .A1(n8721), .A2(n8408), .ZN(n8570) );
  XNOR2_X1 U9892 ( .A(n8412), .B(n8413), .ZN(n8419) );
  AOI22_X1 U9893 ( .A1(n8604), .A2(n8504), .B1(P2_REG3_REG_27__SCAN_IN), .B2(
        P2_U3152), .ZN(n8415) );
  NAND2_X1 U9894 ( .A1(n8599), .A2(n8496), .ZN(n8414) );
  OAI211_X1 U9895 ( .C1(n8416), .C2(n8502), .A(n8415), .B(n8414), .ZN(n8417)
         );
  AOI21_X1 U9896 ( .B1(n8779), .B2(n8509), .A(n8417), .ZN(n8418) );
  OAI21_X1 U9897 ( .B1(n8419), .B2(n8511), .A(n8418), .ZN(P2_U3216) );
  INV_X1 U9898 ( .A(n8674), .ZN(n8514) );
  AOI22_X1 U9899 ( .A1(n7983), .A2(n8473), .B1(n8472), .B2(n8514), .ZN(n8425)
         );
  NOR2_X1 U9900 ( .A1(n8458), .A2(n8502), .ZN(n8422) );
  INV_X1 U9901 ( .A(n8686), .ZN(n8664) );
  AOI22_X1 U9902 ( .A1(n8664), .A2(n8504), .B1(P2_REG3_REG_23__SCAN_IN), .B2(
        P2_U3152), .ZN(n8420) );
  OAI21_X1 U9903 ( .B1(n8656), .B2(n8506), .A(n8420), .ZN(n8421) );
  AOI211_X1 U9904 ( .C1(n8799), .C2(n8509), .A(n8422), .B(n8421), .ZN(n8423)
         );
  OAI21_X1 U9905 ( .B1(n8425), .B2(n8424), .A(n8423), .ZN(P2_U3218) );
  OAI21_X1 U9906 ( .B1(n8432), .B2(n8486), .A(n8426), .ZN(n8427) );
  NAND2_X1 U9907 ( .A1(n8427), .A2(n8473), .ZN(n8436) );
  NAND2_X1 U9908 ( .A1(n8491), .A2(n8516), .ZN(n8428) );
  OAI211_X1 U9909 ( .C1(n8506), .C2(n8732), .A(n8429), .B(n8428), .ZN(n8430)
         );
  AOI21_X1 U9910 ( .B1(n8823), .B2(n8509), .A(n8430), .ZN(n8435) );
  NOR3_X1 U9911 ( .A1(n8432), .A2(n8431), .A3(n8484), .ZN(n8433) );
  OAI21_X1 U9912 ( .B1(n8433), .B2(n8504), .A(n8517), .ZN(n8434) );
  NAND3_X1 U9913 ( .A1(n8436), .A2(n8435), .A3(n8434), .ZN(P2_U3221) );
  INV_X1 U9914 ( .A(n8438), .ZN(n8439) );
  AOI21_X1 U9915 ( .B1(n8437), .B2(n8439), .A(n8511), .ZN(n8443) );
  NOR3_X1 U9916 ( .A1(n8440), .A2(n8722), .A3(n8484), .ZN(n8442) );
  OAI21_X1 U9917 ( .B1(n8443), .B2(n8442), .A(n8441), .ZN(n8448) );
  INV_X1 U9918 ( .A(n8444), .ZN(n8689) );
  AOI22_X1 U9919 ( .A1(n8664), .A2(n8491), .B1(P2_REG3_REG_21__SCAN_IN), .B2(
        P2_U3152), .ZN(n8445) );
  OAI21_X1 U9920 ( .B1(n8722), .B2(n8493), .A(n8445), .ZN(n8446) );
  AOI21_X1 U9921 ( .B1(n8689), .B2(n8496), .A(n8446), .ZN(n8447) );
  OAI211_X1 U9922 ( .C1(n8692), .C2(n8499), .A(n8448), .B(n8447), .ZN(P2_U3225) );
  INV_X1 U9923 ( .A(n8453), .ZN(n8449) );
  NOR3_X1 U9924 ( .A1(n8450), .A2(n8449), .A3(n8511), .ZN(n8456) );
  NAND2_X1 U9925 ( .A1(n8614), .A2(n8472), .ZN(n8451) );
  OAI22_X1 U9926 ( .A1(n8453), .A2(n8511), .B1(n8452), .B2(n8451), .ZN(n8455)
         );
  MUX2_X1 U9927 ( .A(n8456), .B(n8455), .S(n8454), .Z(n8457) );
  INV_X1 U9928 ( .A(n8457), .ZN(n8464) );
  OAI22_X1 U9929 ( .A1(n8459), .A2(n8721), .B1(n8458), .B2(n8719), .ZN(n8631)
         );
  OAI22_X1 U9930 ( .A1(n8628), .A2(n8506), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8460), .ZN(n8461) );
  AOI21_X1 U9931 ( .B1(n8631), .B2(n8462), .A(n8461), .ZN(n8463) );
  OAI211_X1 U9932 ( .C1(n8393), .C2(n8499), .A(n8464), .B(n8463), .ZN(P2_U3227) );
  INV_X1 U9933 ( .A(n8705), .ZN(n8817) );
  AOI21_X1 U9934 ( .B1(n8466), .B2(n8465), .A(n8511), .ZN(n8467) );
  NAND2_X1 U9935 ( .A1(n8467), .A2(n8437), .ZN(n8471) );
  AOI22_X1 U9936 ( .A1(n8515), .A2(n8491), .B1(P2_REG3_REG_20__SCAN_IN), .B2(
        P2_U3152), .ZN(n8468) );
  OAI21_X1 U9937 ( .B1(n8701), .B2(n8493), .A(n8468), .ZN(n8469) );
  AOI21_X1 U9938 ( .B1(n8704), .B2(n8496), .A(n8469), .ZN(n8470) );
  OAI211_X1 U9939 ( .C1(n8817), .C2(n8499), .A(n8471), .B(n8470), .ZN(P2_U3235) );
  NAND2_X1 U9940 ( .A1(n8664), .A2(n8472), .ZN(n8477) );
  NAND2_X1 U9941 ( .A1(n8474), .A2(n8473), .ZN(n8476) );
  MUX2_X1 U9942 ( .A(n8477), .B(n8476), .S(n8475), .Z(n8481) );
  AOI22_X1 U9943 ( .A1(n8515), .A2(n8504), .B1(P2_REG3_REG_22__SCAN_IN), .B2(
        P2_U3152), .ZN(n8478) );
  OAI21_X1 U9944 ( .B1(n8674), .B2(n8502), .A(n8478), .ZN(n8479) );
  AOI21_X1 U9945 ( .B1(n8677), .B2(n8496), .A(n8479), .ZN(n8480) );
  OAI211_X1 U9946 ( .C1(n4483), .C2(n8499), .A(n8481), .B(n8480), .ZN(P2_U3237) );
  INV_X1 U9947 ( .A(n8827), .ZN(n8746) );
  INV_X1 U9948 ( .A(n8482), .ZN(n8483) );
  AOI21_X1 U9949 ( .B1(n7813), .B2(n8483), .A(n8511), .ZN(n8488) );
  NOR3_X1 U9950 ( .A1(n8485), .A2(n8494), .A3(n8484), .ZN(n8487) );
  OAI21_X1 U9951 ( .B1(n8488), .B2(n8487), .A(n8486), .ZN(n8498) );
  INV_X1 U9952 ( .A(n8489), .ZN(n8744) );
  AOI21_X1 U9953 ( .B1(n8491), .B2(n8756), .A(n8490), .ZN(n8492) );
  OAI21_X1 U9954 ( .B1(n8494), .B2(n8493), .A(n8492), .ZN(n8495) );
  AOI21_X1 U9955 ( .B1(n8744), .B2(n8496), .A(n8495), .ZN(n8497) );
  OAI211_X1 U9956 ( .C1(n8746), .C2(n8499), .A(n8498), .B(n8497), .ZN(P2_U3240) );
  XNOR2_X1 U9957 ( .A(n8501), .B(n8500), .ZN(n8512) );
  NOR2_X1 U9958 ( .A1(n8503), .A2(n8502), .ZN(n8508) );
  AOI22_X1 U9959 ( .A1(n8614), .A2(n8504), .B1(P2_REG3_REG_26__SCAN_IN), .B2(
        P2_U3152), .ZN(n8505) );
  OAI21_X1 U9960 ( .B1(n8620), .B2(n8506), .A(n8505), .ZN(n8507) );
  AOI211_X1 U9961 ( .C1(n8785), .C2(n8509), .A(n8508), .B(n8507), .ZN(n8510)
         );
  OAI21_X1 U9962 ( .B1(n8512), .B2(n8511), .A(n8510), .ZN(P2_U3242) );
  MUX2_X1 U9963 ( .A(n8513), .B(P2_DATAO_REG_30__SCAN_IN), .S(n8531), .Z(
        P2_U3582) );
  MUX2_X1 U9964 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(n8603), .S(P2_U3966), .Z(
        P2_U3580) );
  MUX2_X1 U9965 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n8615), .S(P2_U3966), .Z(
        P2_U3579) );
  MUX2_X1 U9966 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(n8604), .S(P2_U3966), .Z(
        P2_U3578) );
  MUX2_X1 U9967 ( .A(n8614), .B(P2_DATAO_REG_25__SCAN_IN), .S(n8531), .Z(
        P2_U3577) );
  MUX2_X1 U9968 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(n8663), .S(P2_U3966), .Z(
        P2_U3576) );
  MUX2_X1 U9969 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(n8514), .S(P2_U3966), .Z(
        P2_U3575) );
  MUX2_X1 U9970 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n8664), .S(P2_U3966), .Z(
        P2_U3574) );
  MUX2_X1 U9971 ( .A(n8515), .B(P2_DATAO_REG_21__SCAN_IN), .S(n8531), .Z(
        P2_U3573) );
  MUX2_X1 U9972 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n8516), .S(P2_U3966), .Z(
        P2_U3572) );
  MUX2_X1 U9973 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n8756), .S(P2_U3966), .Z(
        P2_U3571) );
  MUX2_X1 U9974 ( .A(n8517), .B(P2_DATAO_REG_18__SCAN_IN), .S(n8531), .Z(
        P2_U3570) );
  MUX2_X1 U9975 ( .A(n8754), .B(P2_DATAO_REG_17__SCAN_IN), .S(n8531), .Z(
        P2_U3569) );
  MUX2_X1 U9976 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n8518), .S(P2_U3966), .Z(
        P2_U3568) );
  MUX2_X1 U9977 ( .A(n8519), .B(P2_DATAO_REG_14__SCAN_IN), .S(n8531), .Z(
        P2_U3566) );
  MUX2_X1 U9978 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(n8520), .S(P2_U3966), .Z(
        P2_U3565) );
  MUX2_X1 U9979 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(n8521), .S(P2_U3966), .Z(
        P2_U3564) );
  MUX2_X1 U9980 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(n8522), .S(P2_U3966), .Z(
        P2_U3563) );
  MUX2_X1 U9981 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(n8523), .S(P2_U3966), .Z(
        P2_U3562) );
  MUX2_X1 U9982 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(n8524), .S(P2_U3966), .Z(
        P2_U3561) );
  MUX2_X1 U9983 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(n8525), .S(P2_U3966), .Z(
        P2_U3560) );
  MUX2_X1 U9984 ( .A(n8526), .B(P2_DATAO_REG_7__SCAN_IN), .S(n8531), .Z(
        P2_U3559) );
  MUX2_X1 U9985 ( .A(n8527), .B(P2_DATAO_REG_6__SCAN_IN), .S(n8531), .Z(
        P2_U3558) );
  MUX2_X1 U9986 ( .A(n8528), .B(P2_DATAO_REG_5__SCAN_IN), .S(n8531), .Z(
        P2_U3557) );
  MUX2_X1 U9987 ( .A(n8529), .B(P2_DATAO_REG_4__SCAN_IN), .S(n8531), .Z(
        P2_U3556) );
  MUX2_X1 U9988 ( .A(n8530), .B(P2_DATAO_REG_3__SCAN_IN), .S(n8531), .Z(
        P2_U3555) );
  MUX2_X1 U9989 ( .A(n6632), .B(P2_DATAO_REG_2__SCAN_IN), .S(n8531), .Z(
        P2_U3554) );
  MUX2_X1 U9990 ( .A(n6630), .B(P2_DATAO_REG_1__SCAN_IN), .S(n8531), .Z(
        P2_U3553) );
  MUX2_X1 U9991 ( .A(n6644), .B(P2_DATAO_REG_0__SCAN_IN), .S(n8531), .Z(
        P2_U3552) );
  NOR2_X1 U9992 ( .A1(n4462), .A2(n8532), .ZN(n8534) );
  OAI211_X1 U9993 ( .C1(n8534), .C2(n8533), .A(n9744), .B(n8543), .ZN(n8541)
         );
  AOI22_X1 U9994 ( .A1(n9741), .A2(P2_ADDR_REG_1__SCAN_IN), .B1(
        P2_REG3_REG_1__SCAN_IN), .B2(P2_U3152), .ZN(n8540) );
  NAND2_X1 U9995 ( .A1(n9747), .A2(n8535), .ZN(n8539) );
  OAI211_X1 U9996 ( .C1(n8537), .C2(n8536), .A(n9748), .B(n8549), .ZN(n8538)
         );
  NAND4_X1 U9997 ( .A1(n8541), .A2(n8540), .A3(n8539), .A4(n8538), .ZN(
        P2_U3246) );
  INV_X1 U9998 ( .A(n8542), .ZN(n8547) );
  NAND3_X1 U9999 ( .A1(n8545), .A2(n8544), .A3(n8543), .ZN(n8546) );
  NAND3_X1 U10000 ( .A1(n9744), .A2(n8547), .A3(n8546), .ZN(n8557) );
  AOI22_X1 U10001 ( .A1(n9741), .A2(P2_ADDR_REG_2__SCAN_IN), .B1(
        P2_REG3_REG_2__SCAN_IN), .B2(P2_U3152), .ZN(n8556) );
  NAND2_X1 U10002 ( .A1(n9747), .A2(n8548), .ZN(n8555) );
  MUX2_X1 U10003 ( .A(n6480), .B(P2_REG1_REG_2__SCAN_IN), .S(n8548), .Z(n8551)
         );
  NAND3_X1 U10004 ( .A1(n8551), .A2(n8550), .A3(n8549), .ZN(n8552) );
  NAND3_X1 U10005 ( .A1(n9748), .A2(n8553), .A3(n8552), .ZN(n8554) );
  NAND4_X1 U10006 ( .A1(n8557), .A2(n8556), .A3(n8555), .A4(n8554), .ZN(
        P2_U3247) );
  OAI211_X1 U10007 ( .C1(n8559), .C2(P2_REG1_REG_15__SCAN_IN), .A(n9748), .B(
        n8558), .ZN(n8568) );
  NOR2_X1 U10008 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9998), .ZN(n8560) );
  AOI21_X1 U10009 ( .B1(n9741), .B2(P2_ADDR_REG_15__SCAN_IN), .A(n8560), .ZN(
        n8567) );
  AOI21_X1 U10010 ( .B1(P2_REG2_REG_15__SCAN_IN), .B2(n8562), .A(n8561), .ZN(
        n8563) );
  OR2_X1 U10011 ( .A1(n8563), .A2(n9692), .ZN(n8566) );
  NAND2_X1 U10012 ( .A1(n9747), .A2(n8564), .ZN(n8565) );
  NAND4_X1 U10013 ( .A1(n8568), .A2(n8567), .A3(n8566), .A4(n8565), .ZN(
        P2_U3260) );
  INV_X1 U10014 ( .A(n8765), .ZN(n8575) );
  NAND2_X1 U10015 ( .A1(n8575), .A2(n8574), .ZN(n8569) );
  XNOR2_X1 U10016 ( .A(n8569), .B(n8762), .ZN(n8764) );
  NAND2_X1 U10017 ( .A1(n8571), .A2(n8570), .ZN(n8767) );
  NOR2_X1 U10018 ( .A1(n9772), .A2(n8767), .ZN(n8577) );
  AOI21_X1 U10019 ( .B1(n9772), .B2(P2_REG2_REG_31__SCAN_IN), .A(n8577), .ZN(
        n8573) );
  NAND2_X1 U10020 ( .A1(n8762), .A2(n8736), .ZN(n8572) );
  OAI211_X1 U10021 ( .C1(n8764), .C2(n8708), .A(n8573), .B(n8572), .ZN(
        P2_U3265) );
  XNOR2_X1 U10022 ( .A(n8575), .B(n8574), .ZN(n8768) );
  NOR2_X1 U10023 ( .A1(n8575), .A2(n9768), .ZN(n8576) );
  AOI211_X1 U10024 ( .C1(n9772), .C2(P2_REG2_REG_30__SCAN_IN), .A(n8577), .B(
        n8576), .ZN(n8578) );
  OAI21_X1 U10025 ( .B1(n8768), .B2(n8708), .A(n8578), .ZN(P2_U3266) );
  OAI21_X1 U10026 ( .B1(n8580), .B2(n8586), .A(n8579), .ZN(n8581) );
  INV_X1 U10027 ( .A(n8581), .ZN(n8778) );
  AOI211_X1 U10028 ( .C1(n8775), .C2(n8598), .A(n4275), .B(n8582), .ZN(n8774)
         );
  AOI22_X1 U10029 ( .A1(n8583), .A2(n9760), .B1(P2_REG2_REG_28__SCAN_IN), .B2(
        n9772), .ZN(n8584) );
  OAI21_X1 U10030 ( .B1(n4481), .B2(n9768), .A(n8584), .ZN(n8593) );
  AOI211_X1 U10031 ( .C1(n8587), .C2(n8586), .A(n8698), .B(n8585), .ZN(n8591)
         );
  NOR2_X1 U10032 ( .A1(n8588), .A2(n8721), .ZN(n8590) );
  AOI211_X1 U10033 ( .C1(n8774), .C2(n8676), .A(n8593), .B(n8592), .ZN(n8594)
         );
  OAI21_X1 U10034 ( .B1(n8778), .B2(n8761), .A(n8594), .ZN(P2_U3268) );
  OAI21_X1 U10035 ( .B1(n8596), .B2(n8601), .A(n8595), .ZN(n8597) );
  INV_X1 U10036 ( .A(n8597), .ZN(n8783) );
  AOI21_X1 U10037 ( .B1(n8779), .B2(n8617), .A(n4478), .ZN(n8780) );
  AOI22_X1 U10038 ( .A1(n8599), .A2(n9760), .B1(P2_REG2_REG_27__SCAN_IN), .B2(
        n9772), .ZN(n8600) );
  OAI21_X1 U10039 ( .B1(n4480), .B2(n9768), .A(n8600), .ZN(n8607) );
  XNOR2_X1 U10040 ( .A(n8602), .B(n8601), .ZN(n8605) );
  AOI222_X1 U10041 ( .A1(n9759), .A2(n8605), .B1(n8604), .B2(n8753), .C1(n8603), .C2(n8755), .ZN(n8782) );
  NOR2_X1 U10042 ( .A1(n8782), .A2(n9772), .ZN(n8606) );
  AOI211_X1 U10043 ( .C1(n8780), .C2(n9762), .A(n8607), .B(n8606), .ZN(n8608)
         );
  OAI21_X1 U10044 ( .B1(n8783), .B2(n8761), .A(n8608), .ZN(P2_U3269) );
  OAI21_X1 U10045 ( .B1(n8610), .B2(n8613), .A(n8609), .ZN(n8611) );
  INV_X1 U10046 ( .A(n8611), .ZN(n8788) );
  AOI22_X1 U10047 ( .A1(n8785), .A2(n8736), .B1(n9772), .B2(
        P2_REG2_REG_26__SCAN_IN), .ZN(n8623) );
  XOR2_X1 U10048 ( .A(n8613), .B(n8612), .Z(n8616) );
  AOI222_X1 U10049 ( .A1(n9759), .A2(n8616), .B1(n8615), .B2(n8755), .C1(n8614), .C2(n8753), .ZN(n8787) );
  INV_X1 U10050 ( .A(n8617), .ZN(n8618) );
  AOI211_X1 U10051 ( .C1(n8785), .C2(n8633), .A(n4275), .B(n8618), .ZN(n8784)
         );
  NAND2_X1 U10052 ( .A1(n8784), .A2(n5730), .ZN(n8619) );
  OAI211_X1 U10053 ( .C1(n8731), .C2(n8620), .A(n8787), .B(n8619), .ZN(n8621)
         );
  NAND2_X1 U10054 ( .A1(n8621), .A2(n8734), .ZN(n8622) );
  OAI211_X1 U10055 ( .C1(n8788), .C2(n8761), .A(n8623), .B(n8622), .ZN(
        P2_U3270) );
  OAI21_X1 U10056 ( .B1(n8625), .B2(n8629), .A(n8624), .ZN(n8626) );
  INV_X1 U10057 ( .A(n8626), .ZN(n8793) );
  INV_X1 U10058 ( .A(P2_REG2_REG_25__SCAN_IN), .ZN(n8627) );
  OAI22_X1 U10059 ( .A1(n8628), .A2(n8731), .B1(n8627), .B2(n8734), .ZN(n8638)
         );
  XNOR2_X1 U10060 ( .A(n8630), .B(n8629), .ZN(n8632) );
  AOI21_X1 U10061 ( .B1(n8632), .B2(n9759), .A(n8631), .ZN(n8792) );
  INV_X1 U10062 ( .A(n8645), .ZN(n8635) );
  INV_X1 U10063 ( .A(n8633), .ZN(n8634) );
  AOI211_X1 U10064 ( .C1(n8790), .C2(n8635), .A(n4275), .B(n8634), .ZN(n8789)
         );
  NAND2_X1 U10065 ( .A1(n8789), .A2(n5730), .ZN(n8636) );
  AOI21_X1 U10066 ( .B1(n8792), .B2(n8636), .A(n9772), .ZN(n8637) );
  AOI211_X1 U10067 ( .C1(n8736), .C2(n8790), .A(n8638), .B(n8637), .ZN(n8639)
         );
  OAI21_X1 U10068 ( .B1(n8793), .B2(n8761), .A(n8639), .ZN(P2_U3271) );
  XNOR2_X1 U10069 ( .A(n8640), .B(n8641), .ZN(n8798) );
  XNOR2_X1 U10070 ( .A(n8642), .B(n8641), .ZN(n8643) );
  OAI222_X1 U10071 ( .A1(n8721), .A2(n8644), .B1(n8719), .B2(n8674), .C1(n8698), .C2(n8643), .ZN(n8794) );
  INV_X1 U10072 ( .A(n8655), .ZN(n8646) );
  AOI211_X1 U10073 ( .C1(n8796), .C2(n8646), .A(n4275), .B(n8645), .ZN(n8795)
         );
  NAND2_X1 U10074 ( .A1(n8795), .A2(n8676), .ZN(n8649) );
  AOI22_X1 U10075 ( .A1(n8647), .A2(n9760), .B1(P2_REG2_REG_24__SCAN_IN), .B2(
        n9772), .ZN(n8648) );
  OAI211_X1 U10076 ( .C1(n4654), .C2(n9768), .A(n8649), .B(n8648), .ZN(n8650)
         );
  AOI21_X1 U10077 ( .B1(n8794), .B2(n8734), .A(n8650), .ZN(n8651) );
  OAI21_X1 U10078 ( .B1(n8798), .B2(n8761), .A(n8651), .ZN(P2_U3272) );
  OAI21_X1 U10079 ( .B1(n8654), .B2(n8653), .A(n8652), .ZN(n8803) );
  AOI21_X1 U10080 ( .B1(n8799), .B2(n4818), .A(n8655), .ZN(n8800) );
  INV_X1 U10081 ( .A(n8656), .ZN(n8657) );
  AOI22_X1 U10082 ( .A1(n8657), .A2(n9760), .B1(P2_REG2_REG_23__SCAN_IN), .B2(
        n9772), .ZN(n8658) );
  OAI21_X1 U10083 ( .B1(n8659), .B2(n9768), .A(n8658), .ZN(n8667) );
  OAI21_X1 U10084 ( .B1(n8662), .B2(n8661), .A(n8660), .ZN(n8665) );
  AOI222_X1 U10085 ( .A1(n9759), .A2(n8665), .B1(n8664), .B2(n8753), .C1(n8663), .C2(n8755), .ZN(n8802) );
  NOR2_X1 U10086 ( .A1(n8802), .A2(n9772), .ZN(n8666) );
  AOI211_X1 U10087 ( .C1(n8800), .C2(n9762), .A(n8667), .B(n8666), .ZN(n8668)
         );
  OAI21_X1 U10088 ( .B1(n8761), .B2(n8803), .A(n8668), .ZN(P2_U3273) );
  XOR2_X1 U10089 ( .A(n8672), .B(n8669), .Z(n8808) );
  NOR2_X1 U10090 ( .A1(n4301), .A2(n8670), .ZN(n8671) );
  XOR2_X1 U10091 ( .A(n8672), .B(n8671), .Z(n8673) );
  OAI222_X1 U10092 ( .A1(n8719), .A2(n8700), .B1(n8721), .B2(n8674), .C1(n8673), .C2(n8698), .ZN(n8804) );
  INV_X1 U10093 ( .A(n4818), .ZN(n8675) );
  AOI211_X1 U10094 ( .C1(n8806), .C2(n8687), .A(n4275), .B(n8675), .ZN(n8805)
         );
  NAND2_X1 U10095 ( .A1(n8805), .A2(n8676), .ZN(n8679) );
  AOI22_X1 U10096 ( .A1(n8677), .A2(n9760), .B1(n9772), .B2(
        P2_REG2_REG_22__SCAN_IN), .ZN(n8678) );
  OAI211_X1 U10097 ( .C1(n4483), .C2(n9768), .A(n8679), .B(n8678), .ZN(n8680)
         );
  AOI21_X1 U10098 ( .B1(n8804), .B2(n8734), .A(n8680), .ZN(n8681) );
  OAI21_X1 U10099 ( .B1(n8808), .B2(n8761), .A(n8681), .ZN(P2_U3274) );
  XOR2_X1 U10100 ( .A(n8684), .B(n8682), .Z(n8814) );
  AOI21_X1 U10101 ( .B1(n8684), .B2(n8683), .A(n4301), .ZN(n8685) );
  OAI222_X1 U10102 ( .A1(n8719), .A2(n8722), .B1(n8721), .B2(n8686), .C1(n8698), .C2(n8685), .ZN(n8809) );
  INV_X1 U10103 ( .A(n8687), .ZN(n8688) );
  AOI21_X1 U10104 ( .B1(n8810), .B2(n4485), .A(n8688), .ZN(n8811) );
  NAND2_X1 U10105 ( .A1(n8811), .A2(n9762), .ZN(n8691) );
  AOI22_X1 U10106 ( .A1(n8689), .A2(n9760), .B1(n9772), .B2(
        P2_REG2_REG_21__SCAN_IN), .ZN(n8690) );
  OAI211_X1 U10107 ( .C1(n8692), .C2(n9768), .A(n8691), .B(n8690), .ZN(n8693)
         );
  AOI21_X1 U10108 ( .B1(n8809), .B2(n8734), .A(n8693), .ZN(n8694) );
  OAI21_X1 U10109 ( .B1(n8814), .B2(n8761), .A(n8694), .ZN(P2_U3275) );
  NAND2_X1 U10110 ( .A1(n8716), .A2(n8695), .ZN(n8697) );
  XNOR2_X1 U10111 ( .A(n8697), .B(n8696), .ZN(n8699) );
  OAI222_X1 U10112 ( .A1(n8719), .A2(n8701), .B1(n8721), .B2(n8700), .C1(n8699), .C2(n8698), .ZN(n8820) );
  AND2_X1 U10113 ( .A1(n8726), .A2(n8705), .ZN(n8703) );
  OR2_X1 U10114 ( .A1(n8703), .A2(n8702), .ZN(n8818) );
  AOI22_X1 U10115 ( .A1(n9772), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n8704), .B2(
        n9760), .ZN(n8707) );
  NAND2_X1 U10116 ( .A1(n8705), .A2(n8736), .ZN(n8706) );
  OAI211_X1 U10117 ( .C1(n8818), .C2(n8708), .A(n8707), .B(n8706), .ZN(n8712)
         );
  AND2_X1 U10118 ( .A1(n8710), .A2(n8709), .ZN(n8815) );
  NOR3_X1 U10119 ( .A1(n8816), .A2(n8815), .A3(n8761), .ZN(n8711) );
  AOI211_X1 U10120 ( .C1(n8734), .C2(n8820), .A(n8712), .B(n8711), .ZN(n8713)
         );
  INV_X1 U10121 ( .A(n8713), .ZN(P2_U3276) );
  INV_X1 U10122 ( .A(n8718), .ZN(n8714) );
  XNOR2_X1 U10123 ( .A(n8715), .B(n8714), .ZN(n8826) );
  OAI21_X1 U10124 ( .B1(n8718), .B2(n8717), .A(n8716), .ZN(n8724) );
  OAI22_X1 U10125 ( .A1(n8722), .A2(n8721), .B1(n8720), .B2(n8719), .ZN(n8723)
         );
  AOI21_X1 U10126 ( .B1(n8724), .B2(n9759), .A(n8723), .ZN(n8825) );
  INV_X1 U10127 ( .A(n8725), .ZN(n8742) );
  INV_X1 U10128 ( .A(n8726), .ZN(n8727) );
  AOI211_X1 U10129 ( .C1(n8823), .C2(n8742), .A(n4275), .B(n8727), .ZN(n8822)
         );
  NAND2_X1 U10130 ( .A1(n8822), .A2(n5730), .ZN(n8728) );
  OAI211_X1 U10131 ( .C1(n8826), .C2(n8729), .A(n8825), .B(n8728), .ZN(n8730)
         );
  NAND2_X1 U10132 ( .A1(n8730), .A2(n8734), .ZN(n8738) );
  INV_X1 U10133 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n8733) );
  OAI22_X1 U10134 ( .A1(n8734), .A2(n8733), .B1(n8732), .B2(n8731), .ZN(n8735)
         );
  AOI21_X1 U10135 ( .B1(n8823), .B2(n8736), .A(n8735), .ZN(n8737) );
  OAI211_X1 U10136 ( .C1(n8826), .C2(n8739), .A(n8738), .B(n8737), .ZN(
        P2_U3277) );
  XNOR2_X1 U10137 ( .A(n8741), .B(n8740), .ZN(n8831) );
  AOI21_X1 U10138 ( .B1(n8827), .B2(n8743), .A(n8725), .ZN(n8828) );
  AOI22_X1 U10139 ( .A1(n9772), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n8744), .B2(
        n9760), .ZN(n8745) );
  OAI21_X1 U10140 ( .B1(n8746), .B2(n9768), .A(n8745), .ZN(n8759) );
  INV_X1 U10141 ( .A(n8747), .ZN(n8750) );
  OAI21_X1 U10142 ( .B1(n8750), .B2(n8749), .A(n8748), .ZN(n8752) );
  NAND2_X1 U10143 ( .A1(n8752), .A2(n8751), .ZN(n8757) );
  AOI222_X1 U10144 ( .A1(n9759), .A2(n8757), .B1(n8756), .B2(n8755), .C1(n8754), .C2(n8753), .ZN(n8830) );
  NOR2_X1 U10145 ( .A1(n8830), .A2(n9772), .ZN(n8758) );
  AOI211_X1 U10146 ( .C1(n8828), .C2(n9762), .A(n8759), .B(n8758), .ZN(n8760)
         );
  OAI21_X1 U10147 ( .B1(n8831), .B2(n8761), .A(n8760), .ZN(P2_U3278) );
  NAND2_X1 U10148 ( .A1(n8762), .A2(n8849), .ZN(n8763) );
  OAI211_X1 U10149 ( .C1(n8764), .C2(n4275), .A(n8763), .B(n8767), .ZN(n8854)
         );
  MUX2_X1 U10150 ( .A(P2_REG1_REG_31__SCAN_IN), .B(n8854), .S(n9840), .Z(
        P2_U3551) );
  NAND2_X1 U10151 ( .A1(n8765), .A2(n8849), .ZN(n8766) );
  OAI211_X1 U10152 ( .C1(n8768), .C2(n4275), .A(n8767), .B(n8766), .ZN(n8855)
         );
  MUX2_X1 U10153 ( .A(P2_REG1_REG_30__SCAN_IN), .B(n8855), .S(n9836), .Z(
        P2_U3550) );
  AOI21_X1 U10154 ( .B1(n8849), .B2(n8770), .A(n8769), .ZN(n8771) );
  OAI211_X1 U10155 ( .C1(n8773), .C2(n9798), .A(n8772), .B(n8771), .ZN(n8856)
         );
  MUX2_X1 U10156 ( .A(P2_REG1_REG_29__SCAN_IN), .B(n8856), .S(n9836), .Z(
        P2_U3549) );
  AOI21_X1 U10157 ( .B1(n8849), .B2(n8775), .A(n8774), .ZN(n8776) );
  OAI211_X1 U10158 ( .C1(n8778), .C2(n9798), .A(n8777), .B(n8776), .ZN(n8857)
         );
  MUX2_X1 U10159 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n8857), .S(n9836), .Z(
        P2_U3548) );
  AOI22_X1 U10160 ( .A1(n8780), .A2(n5731), .B1(n8849), .B2(n8779), .ZN(n8781)
         );
  OAI211_X1 U10161 ( .C1(n8783), .C2(n9798), .A(n8782), .B(n8781), .ZN(n8858)
         );
  MUX2_X1 U10162 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n8858), .S(n9836), .Z(
        P2_U3547) );
  AOI21_X1 U10163 ( .B1(n8849), .B2(n8785), .A(n8784), .ZN(n8786) );
  OAI211_X1 U10164 ( .C1(n8788), .C2(n9798), .A(n8787), .B(n8786), .ZN(n8859)
         );
  MUX2_X1 U10165 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n8859), .S(n9836), .Z(
        P2_U3546) );
  AOI21_X1 U10166 ( .B1(n8849), .B2(n8790), .A(n8789), .ZN(n8791) );
  OAI211_X1 U10167 ( .C1(n8793), .C2(n9798), .A(n8792), .B(n8791), .ZN(n8860)
         );
  MUX2_X1 U10168 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n8860), .S(n9836), .Z(
        P2_U3545) );
  AOI211_X1 U10169 ( .C1(n8849), .C2(n8796), .A(n8795), .B(n8794), .ZN(n8797)
         );
  OAI21_X1 U10170 ( .B1(n8798), .B2(n9798), .A(n8797), .ZN(n8861) );
  MUX2_X1 U10171 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n8861), .S(n9840), .Z(
        P2_U3544) );
  AOI22_X1 U10172 ( .A1(n8800), .A2(n5731), .B1(n8849), .B2(n8799), .ZN(n8801)
         );
  OAI211_X1 U10173 ( .C1(n8803), .C2(n9798), .A(n8802), .B(n8801), .ZN(n8862)
         );
  MUX2_X1 U10174 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n8862), .S(n9840), .Z(
        P2_U3543) );
  AOI211_X1 U10175 ( .C1(n8849), .C2(n8806), .A(n8805), .B(n8804), .ZN(n8807)
         );
  OAI21_X1 U10176 ( .B1(n8808), .B2(n9798), .A(n8807), .ZN(n8863) );
  MUX2_X1 U10177 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n8863), .S(n9840), .Z(
        P2_U3542) );
  INV_X1 U10178 ( .A(n8809), .ZN(n8813) );
  AOI22_X1 U10179 ( .A1(n8811), .A2(n5731), .B1(n8849), .B2(n8810), .ZN(n8812)
         );
  OAI211_X1 U10180 ( .C1(n8814), .C2(n9798), .A(n8813), .B(n8812), .ZN(n8864)
         );
  MUX2_X1 U10181 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n8864), .S(n9840), .Z(
        P2_U3541) );
  NOR3_X1 U10182 ( .A1(n8816), .A2(n8815), .A3(n9798), .ZN(n8821) );
  OAI22_X1 U10183 ( .A1(n8818), .A2(n4275), .B1(n8817), .B2(n9819), .ZN(n8819)
         );
  MUX2_X1 U10184 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n8865), .S(n9840), .Z(
        P2_U3540) );
  AOI21_X1 U10185 ( .B1(n8849), .B2(n8823), .A(n8822), .ZN(n8824) );
  OAI211_X1 U10186 ( .C1(n8826), .C2(n9798), .A(n8825), .B(n8824), .ZN(n8866)
         );
  MUX2_X1 U10187 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n8866), .S(n9840), .Z(
        P2_U3539) );
  AOI22_X1 U10188 ( .A1(n8828), .A2(n5731), .B1(n8849), .B2(n8827), .ZN(n8829)
         );
  OAI211_X1 U10189 ( .C1(n9798), .C2(n8831), .A(n8830), .B(n8829), .ZN(n8867)
         );
  MUX2_X1 U10190 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n8867), .S(n9840), .Z(
        P2_U3538) );
  AOI211_X1 U10191 ( .C1(n8849), .C2(n8834), .A(n8833), .B(n8832), .ZN(n8835)
         );
  OAI21_X1 U10192 ( .B1(n9798), .B2(n8836), .A(n8835), .ZN(n8868) );
  MUX2_X1 U10193 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n8868), .S(n9840), .Z(
        P2_U3537) );
  OAI22_X1 U10194 ( .A1(n8838), .A2(n4275), .B1(n8837), .B2(n9819), .ZN(n8840)
         );
  AOI211_X1 U10195 ( .C1(n9825), .C2(n8841), .A(n8840), .B(n8839), .ZN(n8842)
         );
  INV_X1 U10196 ( .A(n8842), .ZN(n8869) );
  MUX2_X1 U10197 ( .A(P2_REG1_REG_15__SCAN_IN), .B(n8869), .S(n9840), .Z(
        P2_U3535) );
  AOI22_X1 U10198 ( .A1(n8844), .A2(n5731), .B1(n8849), .B2(n8843), .ZN(n8845)
         );
  OAI211_X1 U10199 ( .C1(n8847), .C2(n9798), .A(n8846), .B(n8845), .ZN(n8870)
         );
  MUX2_X1 U10200 ( .A(P2_REG1_REG_14__SCAN_IN), .B(n8870), .S(n9840), .Z(
        P2_U3534) );
  AOI22_X1 U10201 ( .A1(n8850), .A2(n5731), .B1(n8849), .B2(n8848), .ZN(n8851)
         );
  OAI211_X1 U10202 ( .C1(n8853), .C2(n9798), .A(n8852), .B(n8851), .ZN(n8871)
         );
  MUX2_X1 U10203 ( .A(P2_REG1_REG_12__SCAN_IN), .B(n8871), .S(n9840), .Z(
        P2_U3532) );
  MUX2_X1 U10204 ( .A(P2_REG0_REG_31__SCAN_IN), .B(n8854), .S(n9828), .Z(
        P2_U3519) );
  MUX2_X1 U10205 ( .A(P2_REG0_REG_30__SCAN_IN), .B(n8855), .S(n9828), .Z(
        P2_U3518) );
  MUX2_X1 U10206 ( .A(P2_REG0_REG_29__SCAN_IN), .B(n8856), .S(n9828), .Z(
        P2_U3517) );
  MUX2_X1 U10207 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n8857), .S(n9828), .Z(
        P2_U3516) );
  MUX2_X1 U10208 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n8858), .S(n9828), .Z(
        P2_U3515) );
  MUX2_X1 U10209 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n8859), .S(n9828), .Z(
        P2_U3514) );
  MUX2_X1 U10210 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n8860), .S(n9828), .Z(
        P2_U3513) );
  MUX2_X1 U10211 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n8861), .S(n9828), .Z(
        P2_U3512) );
  MUX2_X1 U10212 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n8862), .S(n9828), .Z(
        P2_U3511) );
  MUX2_X1 U10213 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n8863), .S(n9828), .Z(
        P2_U3510) );
  MUX2_X1 U10214 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n8864), .S(n9828), .Z(
        P2_U3509) );
  MUX2_X1 U10215 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n8865), .S(n9828), .Z(
        P2_U3508) );
  MUX2_X1 U10216 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n8866), .S(n9828), .Z(
        P2_U3507) );
  MUX2_X1 U10217 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n8867), .S(n9828), .Z(
        P2_U3505) );
  MUX2_X1 U10218 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n8868), .S(n9828), .Z(
        P2_U3502) );
  MUX2_X1 U10219 ( .A(P2_REG0_REG_15__SCAN_IN), .B(n8869), .S(n9828), .Z(
        P2_U3496) );
  MUX2_X1 U10220 ( .A(P2_REG0_REG_14__SCAN_IN), .B(n8870), .S(n9828), .Z(
        P2_U3493) );
  MUX2_X1 U10221 ( .A(P2_REG0_REG_12__SCAN_IN), .B(n8871), .S(n9828), .Z(
        P2_U3487) );
  INV_X1 U10222 ( .A(n8872), .ZN(n9372) );
  NOR4_X1 U10223 ( .A1(n8874), .A2(P2_IR_REG_30__SCAN_IN), .A3(n8873), .A4(
        P2_U3152), .ZN(n8875) );
  AOI21_X1 U10224 ( .B1(n8877), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n8875), .ZN(
        n8876) );
  OAI21_X1 U10225 ( .B1(n9372), .B2(n4284), .A(n8876), .ZN(P2_U3327) );
  AOI22_X1 U10226 ( .A1(n8878), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_30__SCAN_IN), .B2(n8877), .ZN(n8879) );
  OAI21_X1 U10227 ( .B1(n8880), .B2(n4284), .A(n8879), .ZN(P2_U3328) );
  MUX2_X1 U10228 ( .A(n8881), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3358) );
  NOR2_X1 U10229 ( .A1(n8883), .A2(n4566), .ZN(n8884) );
  XNOR2_X1 U10230 ( .A(n8885), .B(n8884), .ZN(n8890) );
  NOR2_X1 U10231 ( .A1(n8989), .A2(n9096), .ZN(n8888) );
  AOI22_X1 U10232 ( .A1(n8965), .A2(n9128), .B1(P1_REG3_REG_27__SCAN_IN), .B2(
        P1_U3084), .ZN(n8886) );
  OAI21_X1 U10233 ( .B1(n8999), .B2(n8963), .A(n8886), .ZN(n8887) );
  AOI211_X1 U10234 ( .C1(n9289), .C2(n8968), .A(n8888), .B(n8887), .ZN(n8889)
         );
  OAI21_X1 U10235 ( .B1(n8890), .B2(n8984), .A(n8889), .ZN(P1_U3212) );
  NAND2_X1 U10236 ( .A1(n4364), .A2(n8892), .ZN(n8894) );
  XNOR2_X1 U10237 ( .A(n8894), .B(n8893), .ZN(n8899) );
  AOI22_X1 U10238 ( .A1(n8994), .A2(n9155), .B1(P1_REG3_REG_23__SCAN_IN), .B2(
        P1_U3084), .ZN(n8896) );
  NAND2_X1 U10239 ( .A1(n8965), .A2(n9187), .ZN(n8895) );
  OAI211_X1 U10240 ( .C1(n8989), .C2(n9157), .A(n8896), .B(n8895), .ZN(n8897)
         );
  AOI21_X1 U10241 ( .B1(n9308), .B2(n8968), .A(n8897), .ZN(n8898) );
  OAI21_X1 U10242 ( .B1(n8899), .B2(n8984), .A(n8898), .ZN(P1_U3214) );
  XOR2_X1 U10243 ( .A(n8900), .B(n8901), .Z(n8907) );
  NAND2_X1 U10244 ( .A1(P1_U3084), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n9063) );
  OAI21_X1 U10245 ( .B1(n8963), .B2(n8902), .A(n9063), .ZN(n8903) );
  AOI21_X1 U10246 ( .B1(n8965), .B2(n9244), .A(n8903), .ZN(n8904) );
  OAI21_X1 U10247 ( .B1(n9208), .B2(n8989), .A(n8904), .ZN(n8905) );
  AOI21_X1 U10248 ( .B1(n9329), .B2(n8968), .A(n8905), .ZN(n8906) );
  OAI21_X1 U10249 ( .B1(n8907), .B2(n8984), .A(n8906), .ZN(P1_U3217) );
  NOR2_X1 U10250 ( .A1(n4333), .A2(n8909), .ZN(n8910) );
  XNOR2_X1 U10251 ( .A(n8908), .B(n8910), .ZN(n8915) );
  AOI22_X1 U10252 ( .A1(n8994), .A2(n9187), .B1(P1_REG3_REG_21__SCAN_IN), .B2(
        P1_U3084), .ZN(n8912) );
  NAND2_X1 U10253 ( .A1(n8965), .A2(n9213), .ZN(n8911) );
  OAI211_X1 U10254 ( .C1(n8989), .C2(n9181), .A(n8912), .B(n8911), .ZN(n8913)
         );
  AOI21_X1 U10255 ( .B1(n9319), .B2(n8968), .A(n8913), .ZN(n8914) );
  OAI21_X1 U10256 ( .B1(n8915), .B2(n8984), .A(n8914), .ZN(P1_U3221) );
  XOR2_X1 U10257 ( .A(n8917), .B(n8916), .Z(n8922) );
  AOI22_X1 U10258 ( .A1(n8994), .A2(n9128), .B1(P1_REG3_REG_25__SCAN_IN), .B2(
        P1_U3084), .ZN(n8919) );
  NAND2_X1 U10259 ( .A1(n8965), .A2(n9155), .ZN(n8918) );
  OAI211_X1 U10260 ( .C1(n8989), .C2(n9122), .A(n8919), .B(n8918), .ZN(n8920)
         );
  AOI21_X1 U10261 ( .B1(n9299), .B2(n8968), .A(n8920), .ZN(n8921) );
  OAI21_X1 U10262 ( .B1(n8922), .B2(n8984), .A(n8921), .ZN(P1_U3223) );
  NAND2_X1 U10263 ( .A1(n8924), .A2(n8923), .ZN(n8925) );
  XNOR2_X1 U10264 ( .A(n8926), .B(n8925), .ZN(n8933) );
  OAI21_X1 U10265 ( .B1(n8963), .B2(n8928), .A(n8927), .ZN(n8929) );
  AOI21_X1 U10266 ( .B1(n8965), .B2(n9243), .A(n8929), .ZN(n8930) );
  OAI21_X1 U10267 ( .B1(n9237), .B2(n8989), .A(n8930), .ZN(n8931) );
  AOI21_X1 U10268 ( .B1(n9339), .B2(n8968), .A(n8931), .ZN(n8932) );
  OAI21_X1 U10269 ( .B1(n8933), .B2(n8984), .A(n8932), .ZN(P1_U3226) );
  XOR2_X1 U10270 ( .A(n8935), .B(n8934), .Z(n8940) );
  INV_X1 U10271 ( .A(n8977), .ZN(n9137) );
  AOI22_X1 U10272 ( .A1(n8994), .A2(n9137), .B1(P1_REG3_REG_24__SCAN_IN), .B2(
        P1_U3084), .ZN(n8937) );
  NAND2_X1 U10273 ( .A1(n8965), .A2(n9172), .ZN(n8936) );
  OAI211_X1 U10274 ( .C1(n8989), .C2(n9143), .A(n8937), .B(n8936), .ZN(n8938)
         );
  AOI21_X1 U10275 ( .B1(n5402), .B2(n8968), .A(n8938), .ZN(n8939) );
  OAI21_X1 U10276 ( .B1(n8940), .B2(n8984), .A(n8939), .ZN(P1_U3227) );
  XNOR2_X1 U10277 ( .A(n8942), .B(n8941), .ZN(n8943) );
  XNOR2_X1 U10278 ( .A(n8944), .B(n8943), .ZN(n8949) );
  AOI22_X1 U10279 ( .A1(n8994), .A2(n9200), .B1(P1_REG3_REG_20__SCAN_IN), .B2(
        P1_U3084), .ZN(n8946) );
  NAND2_X1 U10280 ( .A1(n8965), .A2(n9228), .ZN(n8945) );
  OAI211_X1 U10281 ( .C1(n8989), .C2(n9194), .A(n8946), .B(n8945), .ZN(n8947)
         );
  AOI21_X1 U10282 ( .B1(n9324), .B2(n8968), .A(n8947), .ZN(n8948) );
  OAI21_X1 U10283 ( .B1(n8949), .B2(n8984), .A(n8948), .ZN(P1_U3231) );
  NAND2_X1 U10284 ( .A1(n8950), .A2(n4571), .ZN(n8952) );
  XNOR2_X1 U10285 ( .A(n8952), .B(n8951), .ZN(n8957) );
  AOI22_X1 U10286 ( .A1(n8994), .A2(n9172), .B1(P1_REG3_REG_22__SCAN_IN), .B2(
        P1_U3084), .ZN(n8954) );
  NAND2_X1 U10287 ( .A1(n8965), .A2(n9200), .ZN(n8953) );
  OAI211_X1 U10288 ( .C1(n8989), .C2(n9164), .A(n8954), .B(n8953), .ZN(n8955)
         );
  AOI21_X1 U10289 ( .B1(n9314), .B2(n8968), .A(n8955), .ZN(n8956) );
  OAI21_X1 U10290 ( .B1(n8957), .B2(n8984), .A(n8956), .ZN(P1_U3233) );
  NAND2_X1 U10291 ( .A1(n8958), .A2(n8959), .ZN(n8961) );
  XNOR2_X1 U10292 ( .A(n8961), .B(n8960), .ZN(n8970) );
  NAND2_X1 U10293 ( .A1(P1_U3084), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n9046) );
  OAI21_X1 U10294 ( .B1(n8963), .B2(n8962), .A(n9046), .ZN(n8964) );
  AOI21_X1 U10295 ( .B1(n8965), .B2(n9262), .A(n8964), .ZN(n8966) );
  OAI21_X1 U10296 ( .B1(n9221), .B2(n8989), .A(n8966), .ZN(n8967) );
  AOI21_X1 U10297 ( .B1(n9334), .B2(n8968), .A(n8967), .ZN(n8969) );
  OAI21_X1 U10298 ( .B1(n8970), .B2(n8984), .A(n8969), .ZN(P1_U3236) );
  OAI211_X1 U10299 ( .C1(n8971), .C2(n8974), .A(n8972), .B(n8973), .ZN(n8981)
         );
  INV_X1 U10300 ( .A(n8975), .ZN(n9109) );
  AOI22_X1 U10301 ( .A1(n8994), .A2(n9114), .B1(P1_REG3_REG_26__SCAN_IN), .B2(
        P1_U3084), .ZN(n8976) );
  OAI21_X1 U10302 ( .B1(n8977), .B2(n8991), .A(n8976), .ZN(n8978) );
  AOI21_X1 U10303 ( .B1(n9109), .B2(n8979), .A(n8978), .ZN(n8980) );
  OAI211_X1 U10304 ( .C1(n9111), .C2(n8997), .A(n8981), .B(n8980), .ZN(
        P1_U3238) );
  INV_X1 U10305 ( .A(n7846), .ZN(n8987) );
  AOI21_X1 U10306 ( .B1(n7846), .B2(n8983), .A(n8982), .ZN(n8985) );
  NOR2_X1 U10307 ( .A1(n8985), .A2(n8984), .ZN(n8986) );
  OAI21_X1 U10308 ( .B1(n8987), .B2(n7845), .A(n8986), .ZN(n8996) );
  NOR2_X1 U10309 ( .A1(n8989), .A2(n8988), .ZN(n8993) );
  OAI21_X1 U10310 ( .B1(n8991), .B2(n9401), .A(n8990), .ZN(n8992) );
  AOI211_X1 U10311 ( .C1(n8994), .C2(n9243), .A(n8993), .B(n8992), .ZN(n8995)
         );
  OAI211_X1 U10312 ( .C1(n9437), .C2(n8997), .A(n8996), .B(n8995), .ZN(
        P1_U3239) );
  MUX2_X1 U10313 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n8998), .S(P1_U4006), .Z(
        P1_U3585) );
  MUX2_X1 U10314 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n9087), .S(P1_U4006), .Z(
        P1_U3584) );
  INV_X1 U10315 ( .A(n8999), .ZN(n9102) );
  MUX2_X1 U10316 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n9102), .S(P1_U4006), .Z(
        P1_U3583) );
  MUX2_X1 U10317 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n9128), .S(P1_U4006), .Z(
        P1_U3581) );
  MUX2_X1 U10318 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n9137), .S(P1_U4006), .Z(
        P1_U3580) );
  MUX2_X1 U10319 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n9155), .S(P1_U4006), .Z(
        P1_U3579) );
  MUX2_X1 U10320 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n9172), .S(P1_U4006), .Z(
        P1_U3578) );
  MUX2_X1 U10321 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n9187), .S(P1_U4006), .Z(
        P1_U3577) );
  MUX2_X1 U10322 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n9200), .S(P1_U4006), .Z(
        P1_U3576) );
  MUX2_X1 U10323 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n9213), .S(P1_U4006), .Z(
        P1_U3575) );
  MUX2_X1 U10324 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n9228), .S(P1_U4006), .Z(
        P1_U3574) );
  MUX2_X1 U10325 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n9244), .S(P1_U4006), .Z(
        P1_U3573) );
  MUX2_X1 U10326 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n9262), .S(P1_U4006), .Z(
        P1_U3572) );
  MUX2_X1 U10327 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n9243), .S(P1_U4006), .Z(
        P1_U3571) );
  MUX2_X1 U10328 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n9260), .S(P1_U4006), .Z(
        P1_U3570) );
  MUX2_X1 U10329 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n9000), .S(P1_U4006), .Z(
        P1_U3568) );
  MUX2_X1 U10330 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n9001), .S(P1_U4006), .Z(
        P1_U3567) );
  MUX2_X1 U10331 ( .A(n9002), .B(P1_DATAO_REG_11__SCAN_IN), .S(n9009), .Z(
        P1_U3566) );
  MUX2_X1 U10332 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n9003), .S(P1_U4006), .Z(
        P1_U3565) );
  MUX2_X1 U10333 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n9004), .S(P1_U4006), .Z(
        P1_U3564) );
  MUX2_X1 U10334 ( .A(n9005), .B(P1_DATAO_REG_8__SCAN_IN), .S(n9009), .Z(
        P1_U3563) );
  MUX2_X1 U10335 ( .A(n9006), .B(P1_DATAO_REG_7__SCAN_IN), .S(n9009), .Z(
        P1_U3562) );
  MUX2_X1 U10336 ( .A(n9575), .B(P1_DATAO_REG_6__SCAN_IN), .S(n9009), .Z(
        P1_U3561) );
  MUX2_X1 U10337 ( .A(n9007), .B(P1_DATAO_REG_5__SCAN_IN), .S(n9009), .Z(
        P1_U3560) );
  MUX2_X1 U10338 ( .A(n9585), .B(P1_DATAO_REG_4__SCAN_IN), .S(n9009), .Z(
        P1_U3559) );
  MUX2_X1 U10339 ( .A(n9008), .B(P1_DATAO_REG_3__SCAN_IN), .S(n9009), .Z(
        P1_U3558) );
  MUX2_X1 U10340 ( .A(n6448), .B(P1_DATAO_REG_2__SCAN_IN), .S(n9009), .Z(
        P1_U3557) );
  MUX2_X1 U10341 ( .A(n6897), .B(P1_DATAO_REG_1__SCAN_IN), .S(n9009), .Z(
        P1_U3556) );
  MUX2_X1 U10342 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(n6360), .S(P1_U4006), .Z(
        P1_U3555) );
  OAI22_X1 U10343 ( .A1(n9538), .A2(n9010), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n6796), .ZN(n9011) );
  AOI21_X1 U10344 ( .B1(n9508), .B2(P1_ADDR_REG_1__SCAN_IN), .A(n9011), .ZN(
        n9020) );
  OAI211_X1 U10345 ( .C1(n9014), .C2(n9013), .A(n9566), .B(n9012), .ZN(n9019)
         );
  OAI211_X1 U10346 ( .C1(n9017), .C2(n9016), .A(n9556), .B(n9015), .ZN(n9018)
         );
  NAND3_X1 U10347 ( .A1(n9020), .A2(n9019), .A3(n9018), .ZN(P1_U3242) );
  INV_X1 U10348 ( .A(n9021), .ZN(n9022) );
  OAI21_X1 U10349 ( .B1(n9538), .B2(n9023), .A(n9022), .ZN(n9024) );
  AOI21_X1 U10350 ( .B1(n9508), .B2(P1_ADDR_REG_3__SCAN_IN), .A(n9024), .ZN(
        n9033) );
  OAI211_X1 U10351 ( .C1(n9027), .C2(n9026), .A(n9556), .B(n9025), .ZN(n9032)
         );
  OAI211_X1 U10352 ( .C1(n9030), .C2(n9029), .A(n9566), .B(n9028), .ZN(n9031)
         );
  NAND3_X1 U10353 ( .A1(n9033), .A2(n9032), .A3(n9031), .ZN(P1_U3244) );
  INV_X1 U10354 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n9050) );
  XNOR2_X1 U10355 ( .A(n9055), .B(n9034), .ZN(n9037) );
  AOI21_X1 U10356 ( .B1(n9039), .B2(P1_REG1_REG_17__SCAN_IN), .A(n9035), .ZN(
        n9036) );
  NAND2_X1 U10357 ( .A1(n9037), .A2(n9036), .ZN(n9057) );
  OAI21_X1 U10358 ( .B1(n9037), .B2(n9036), .A(n9057), .ZN(n9045) );
  NAND2_X1 U10359 ( .A1(n9055), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n9051) );
  OR2_X1 U10360 ( .A1(n9055), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n9040) );
  NAND2_X1 U10361 ( .A1(n9051), .A2(n9040), .ZN(n9042) );
  INV_X1 U10362 ( .A(n9052), .ZN(n9041) );
  AOI211_X1 U10363 ( .C1(n9043), .C2(n9042), .A(n9041), .B(n9543), .ZN(n9044)
         );
  AOI21_X1 U10364 ( .B1(n9566), .B2(n9045), .A(n9044), .ZN(n9049) );
  INV_X1 U10365 ( .A(n9046), .ZN(n9047) );
  AOI21_X1 U10366 ( .B1(n9553), .B2(n9055), .A(n9047), .ZN(n9048) );
  OAI211_X1 U10367 ( .C1(n9571), .C2(n9050), .A(n9049), .B(n9048), .ZN(
        P1_U3259) );
  NAND2_X1 U10368 ( .A1(n9052), .A2(n9051), .ZN(n9054) );
  XNOR2_X1 U10369 ( .A(n9054), .B(n9053), .ZN(n9060) );
  OR2_X1 U10370 ( .A1(n9055), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n9056) );
  NAND2_X1 U10371 ( .A1(n9057), .A2(n9056), .ZN(n9058) );
  XNOR2_X1 U10372 ( .A(n9058), .B(P1_REG1_REG_19__SCAN_IN), .ZN(n9061) );
  OR2_X1 U10373 ( .A1(n9522), .A2(n9061), .ZN(n9059) );
  AOI22_X1 U10374 ( .A1(n9566), .A2(n9061), .B1(n9556), .B2(n9060), .ZN(n9062)
         );
  NAND2_X1 U10375 ( .A1(n9276), .A2(n9069), .ZN(n9064) );
  NAND2_X1 U10376 ( .A1(n9269), .A2(n9417), .ZN(n9068) );
  NAND2_X1 U10377 ( .A1(n9066), .A2(n9065), .ZN(n9274) );
  NOR2_X1 U10378 ( .A1(n4283), .A2(n9274), .ZN(n9071) );
  AOI21_X1 U10379 ( .B1(n4283), .B2(P1_REG2_REG_31__SCAN_IN), .A(n9071), .ZN(
        n9067) );
  OAI211_X1 U10380 ( .C1(n9270), .C2(n9256), .A(n9068), .B(n9067), .ZN(
        P1_U3261) );
  XNOR2_X1 U10381 ( .A(n9070), .B(n9069), .ZN(n9273) );
  NAND2_X1 U10382 ( .A1(n9273), .A2(n9417), .ZN(n9073) );
  AOI21_X1 U10383 ( .B1(n4283), .B2(P1_REG2_REG_30__SCAN_IN), .A(n9071), .ZN(
        n9072) );
  OAI211_X1 U10384 ( .C1(n9276), .C2(n9256), .A(n9073), .B(n9072), .ZN(
        P1_U3262) );
  OAI21_X1 U10385 ( .B1(n9076), .B2(n9075), .A(n9074), .ZN(n9288) );
  AOI21_X1 U10386 ( .B1(n9284), .B2(n9094), .A(n9077), .ZN(n9285) );
  INV_X1 U10387 ( .A(n9078), .ZN(n9079) );
  AOI22_X1 U10388 ( .A1(n4283), .A2(P1_REG2_REG_28__SCAN_IN), .B1(n9079), .B2(
        n9588), .ZN(n9080) );
  OAI21_X1 U10389 ( .B1(n9081), .B2(n9256), .A(n9080), .ZN(n9090) );
  AND2_X1 U10390 ( .A1(n9083), .A2(n9082), .ZN(n9086) );
  OAI21_X1 U10391 ( .B1(n9086), .B2(n9085), .A(n9084), .ZN(n9088) );
  AOI222_X1 U10392 ( .A1(n9427), .A2(n9088), .B1(n9087), .B2(n9261), .C1(n9114), .C2(n9586), .ZN(n9287) );
  NOR2_X1 U10393 ( .A1(n9287), .A2(n4283), .ZN(n9089) );
  AOI211_X1 U10394 ( .C1(n9417), .C2(n9285), .A(n9090), .B(n9089), .ZN(n9091)
         );
  OAI21_X1 U10395 ( .B1(n9288), .B2(n9268), .A(n9091), .ZN(P1_U3263) );
  XNOR2_X1 U10396 ( .A(n9093), .B(n9092), .ZN(n9293) );
  INV_X1 U10397 ( .A(n9094), .ZN(n9095) );
  AOI21_X1 U10398 ( .B1(n9289), .B2(n9108), .A(n9095), .ZN(n9290) );
  INV_X1 U10399 ( .A(n9096), .ZN(n9097) );
  AOI22_X1 U10400 ( .A1(n4283), .A2(P1_REG2_REG_27__SCAN_IN), .B1(n9097), .B2(
        n9588), .ZN(n9098) );
  OAI21_X1 U10401 ( .B1(n9099), .B2(n9256), .A(n9098), .ZN(n9105) );
  XNOR2_X1 U10402 ( .A(n9101), .B(n9100), .ZN(n9103) );
  AOI222_X1 U10403 ( .A1(n9427), .A2(n9103), .B1(n9102), .B2(n9261), .C1(n9128), .C2(n9586), .ZN(n9292) );
  NOR2_X1 U10404 ( .A1(n9292), .A2(n4283), .ZN(n9104) );
  AOI211_X1 U10405 ( .C1(n9417), .C2(n9290), .A(n9105), .B(n9104), .ZN(n9106)
         );
  OAI21_X1 U10406 ( .B1(n9293), .B2(n9268), .A(n9106), .ZN(P1_U3264) );
  XNOR2_X1 U10407 ( .A(n9107), .B(n9113), .ZN(n9298) );
  AOI21_X1 U10408 ( .B1(n9294), .B2(n9120), .A(n4470), .ZN(n9295) );
  AOI22_X1 U10409 ( .A1(n4283), .A2(P1_REG2_REG_26__SCAN_IN), .B1(n9109), .B2(
        n9588), .ZN(n9110) );
  OAI21_X1 U10410 ( .B1(n9111), .B2(n9256), .A(n9110), .ZN(n9117) );
  XOR2_X1 U10411 ( .A(n9113), .B(n9112), .Z(n9115) );
  AOI222_X1 U10412 ( .A1(n9427), .A2(n9115), .B1(n9114), .B2(n9261), .C1(n9137), .C2(n9586), .ZN(n9297) );
  NOR2_X1 U10413 ( .A1(n9297), .A2(n4283), .ZN(n9116) );
  AOI211_X1 U10414 ( .C1(n9417), .C2(n9295), .A(n9117), .B(n9116), .ZN(n9118)
         );
  OAI21_X1 U10415 ( .B1(n9298), .B2(n9268), .A(n9118), .ZN(P1_U3265) );
  XOR2_X1 U10416 ( .A(n9126), .B(n9119), .Z(n9303) );
  INV_X1 U10417 ( .A(n9139), .ZN(n9121) );
  AOI21_X1 U10418 ( .B1(n9299), .B2(n9121), .A(n4471), .ZN(n9300) );
  INV_X1 U10419 ( .A(n9122), .ZN(n9123) );
  AOI22_X1 U10420 ( .A1(n4283), .A2(P1_REG2_REG_25__SCAN_IN), .B1(n9123), .B2(
        n9588), .ZN(n9124) );
  OAI21_X1 U10421 ( .B1(n9125), .B2(n9256), .A(n9124), .ZN(n9131) );
  XNOR2_X1 U10422 ( .A(n9127), .B(n9126), .ZN(n9129) );
  AOI222_X1 U10423 ( .A1(n9427), .A2(n9129), .B1(n9128), .B2(n9261), .C1(n9155), .C2(n9586), .ZN(n9302) );
  NOR2_X1 U10424 ( .A1(n9302), .A2(n4283), .ZN(n9130) );
  AOI211_X1 U10425 ( .C1(n9300), .C2(n9417), .A(n9131), .B(n9130), .ZN(n9132)
         );
  OAI21_X1 U10426 ( .B1(n9303), .B2(n9268), .A(n9132), .ZN(P1_U3266) );
  XNOR2_X1 U10427 ( .A(n9133), .B(n9134), .ZN(n9307) );
  AOI22_X1 U10428 ( .A1(n5402), .A2(n9434), .B1(P1_REG2_REG_24__SCAN_IN), .B2(
        n4283), .ZN(n9146) );
  INV_X1 U10429 ( .A(n9134), .ZN(n9135) );
  XNOR2_X1 U10430 ( .A(n9136), .B(n9135), .ZN(n9138) );
  AOI222_X1 U10431 ( .A1(n9427), .A2(n9138), .B1(n9172), .B2(n9586), .C1(n9137), .C2(n9261), .ZN(n9306) );
  INV_X1 U10432 ( .A(n9149), .ZN(n9140) );
  AOI211_X1 U10433 ( .C1(n5402), .C2(n9140), .A(n9660), .B(n9139), .ZN(n9304)
         );
  NAND2_X1 U10434 ( .A1(n9304), .A2(n9141), .ZN(n9142) );
  OAI211_X1 U10435 ( .C1(n9418), .C2(n9143), .A(n9306), .B(n9142), .ZN(n9144)
         );
  NAND2_X1 U10436 ( .A1(n9144), .A2(n9600), .ZN(n9145) );
  OAI211_X1 U10437 ( .C1(n9307), .C2(n9268), .A(n9146), .B(n9145), .ZN(
        P1_U3267) );
  XOR2_X1 U10438 ( .A(n9153), .B(n9147), .Z(n9312) );
  AND2_X1 U10439 ( .A1(n9162), .A2(n9308), .ZN(n9148) );
  NOR2_X1 U10440 ( .A1(n9149), .A2(n9148), .ZN(n9309) );
  OAI22_X1 U10441 ( .A1(n9151), .A2(n9256), .B1(n9150), .B2(n9600), .ZN(n9152)
         );
  AOI21_X1 U10442 ( .B1(n9309), .B2(n9417), .A(n9152), .ZN(n9160) );
  XOR2_X1 U10443 ( .A(n9154), .B(n9153), .Z(n9156) );
  AOI222_X1 U10444 ( .A1(n9427), .A2(n9156), .B1(n9187), .B2(n9586), .C1(n9155), .C2(n9261), .ZN(n9311) );
  OAI21_X1 U10445 ( .B1(n9157), .B2(n9418), .A(n9311), .ZN(n9158) );
  NAND2_X1 U10446 ( .A1(n9158), .A2(n9600), .ZN(n9159) );
  OAI211_X1 U10447 ( .C1(n9312), .C2(n9268), .A(n9160), .B(n9159), .ZN(
        P1_U3268) );
  XNOR2_X1 U10448 ( .A(n9161), .B(n9171), .ZN(n9317) );
  INV_X1 U10449 ( .A(n9162), .ZN(n9163) );
  AOI211_X1 U10450 ( .C1(n9314), .C2(n9178), .A(n9660), .B(n9163), .ZN(n9313)
         );
  INV_X1 U10451 ( .A(n9164), .ZN(n9165) );
  AOI22_X1 U10452 ( .A1(n4283), .A2(P1_REG2_REG_22__SCAN_IN), .B1(n9165), .B2(
        n9588), .ZN(n9166) );
  OAI21_X1 U10453 ( .B1(n9167), .B2(n9256), .A(n9166), .ZN(n9175) );
  NAND2_X1 U10454 ( .A1(n9169), .A2(n9168), .ZN(n9170) );
  XOR2_X1 U10455 ( .A(n9171), .B(n9170), .Z(n9173) );
  AOI222_X1 U10456 ( .A1(n9427), .A2(n9173), .B1(n9200), .B2(n9586), .C1(n9172), .C2(n9261), .ZN(n9316) );
  NOR2_X1 U10457 ( .A1(n9316), .A2(n4283), .ZN(n9174) );
  AOI211_X1 U10458 ( .C1(n9313), .C2(n9266), .A(n9175), .B(n9174), .ZN(n9176)
         );
  OAI21_X1 U10459 ( .B1(n9268), .B2(n9317), .A(n9176), .ZN(P1_U3269) );
  XNOR2_X1 U10460 ( .A(n9177), .B(n9185), .ZN(n9322) );
  INV_X1 U10461 ( .A(n9193), .ZN(n9180) );
  INV_X1 U10462 ( .A(n9178), .ZN(n9179) );
  AOI211_X1 U10463 ( .C1(n9319), .C2(n9180), .A(n9660), .B(n9179), .ZN(n9318)
         );
  INV_X1 U10464 ( .A(n9181), .ZN(n9182) );
  AOI22_X1 U10465 ( .A1(n4283), .A2(P1_REG2_REG_21__SCAN_IN), .B1(n9182), .B2(
        n9588), .ZN(n9183) );
  OAI21_X1 U10466 ( .B1(n9184), .B2(n9256), .A(n9183), .ZN(n9190) );
  XNOR2_X1 U10467 ( .A(n9186), .B(n9185), .ZN(n9188) );
  AOI222_X1 U10468 ( .A1(n9427), .A2(n9188), .B1(n9187), .B2(n9261), .C1(n9213), .C2(n9586), .ZN(n9321) );
  NOR2_X1 U10469 ( .A1(n9321), .A2(n4283), .ZN(n9189) );
  AOI211_X1 U10470 ( .C1(n9266), .C2(n9318), .A(n9190), .B(n9189), .ZN(n9191)
         );
  OAI21_X1 U10471 ( .B1(n9268), .B2(n9322), .A(n9191), .ZN(P1_U3270) );
  XNOR2_X1 U10472 ( .A(n9192), .B(n9199), .ZN(n9327) );
  AOI211_X1 U10473 ( .C1(n9324), .C2(n9206), .A(n9660), .B(n9193), .ZN(n9323)
         );
  INV_X1 U10474 ( .A(n9194), .ZN(n9195) );
  AOI22_X1 U10475 ( .A1(n4283), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n9195), .B2(
        n9588), .ZN(n9196) );
  OAI21_X1 U10476 ( .B1(n9197), .B2(n9256), .A(n9196), .ZN(n9203) );
  XOR2_X1 U10477 ( .A(n9199), .B(n9198), .Z(n9201) );
  AOI222_X1 U10478 ( .A1(n9427), .A2(n9201), .B1(n9200), .B2(n9261), .C1(n9228), .C2(n9586), .ZN(n9326) );
  NOR2_X1 U10479 ( .A1(n9326), .A2(n4283), .ZN(n9202) );
  AOI211_X1 U10480 ( .C1(n9266), .C2(n9323), .A(n9203), .B(n9202), .ZN(n9204)
         );
  OAI21_X1 U10481 ( .B1(n9327), .B2(n9268), .A(n9204), .ZN(P1_U3271) );
  XOR2_X1 U10482 ( .A(n9211), .B(n9205), .Z(n9332) );
  INV_X1 U10483 ( .A(n9206), .ZN(n9207) );
  AOI211_X1 U10484 ( .C1(n9329), .C2(n9219), .A(n9660), .B(n9207), .ZN(n9328)
         );
  INV_X1 U10485 ( .A(n9208), .ZN(n9209) );
  AOI22_X1 U10486 ( .A1(n4283), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n9209), .B2(
        n9588), .ZN(n9210) );
  OAI21_X1 U10487 ( .B1(n4474), .B2(n9256), .A(n9210), .ZN(n9216) );
  XNOR2_X1 U10488 ( .A(n9212), .B(n9211), .ZN(n9214) );
  AOI222_X1 U10489 ( .A1(n9427), .A2(n9214), .B1(n9213), .B2(n9261), .C1(n9244), .C2(n9586), .ZN(n9331) );
  NOR2_X1 U10490 ( .A1(n9331), .A2(n4283), .ZN(n9215) );
  AOI211_X1 U10491 ( .C1(n9328), .C2(n9266), .A(n9216), .B(n9215), .ZN(n9217)
         );
  OAI21_X1 U10492 ( .B1(n9332), .B2(n9268), .A(n9217), .ZN(P1_U3272) );
  XNOR2_X1 U10493 ( .A(n9218), .B(n9226), .ZN(n9337) );
  INV_X1 U10494 ( .A(n9219), .ZN(n9220) );
  AOI211_X1 U10495 ( .C1(n9334), .C2(n9234), .A(n9660), .B(n9220), .ZN(n9333)
         );
  INV_X1 U10496 ( .A(n9221), .ZN(n9222) );
  AOI22_X1 U10497 ( .A1(n4283), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n9222), .B2(
        n9588), .ZN(n9223) );
  OAI21_X1 U10498 ( .B1(n4475), .B2(n9256), .A(n9223), .ZN(n9231) );
  NAND2_X1 U10499 ( .A1(n9225), .A2(n9224), .ZN(n9227) );
  XNOR2_X1 U10500 ( .A(n9227), .B(n9226), .ZN(n9229) );
  AOI222_X1 U10501 ( .A1(n9427), .A2(n9229), .B1(n9228), .B2(n9261), .C1(n9262), .C2(n9586), .ZN(n9336) );
  NOR2_X1 U10502 ( .A1(n9336), .A2(n4283), .ZN(n9230) );
  AOI211_X1 U10503 ( .C1(n9333), .C2(n9266), .A(n9231), .B(n9230), .ZN(n9232)
         );
  OAI21_X1 U10504 ( .B1(n9268), .B2(n9337), .A(n9232), .ZN(P1_U3273) );
  XNOR2_X1 U10505 ( .A(n9233), .B(n9242), .ZN(n9342) );
  INV_X1 U10506 ( .A(n9251), .ZN(n9236) );
  INV_X1 U10507 ( .A(n9234), .ZN(n9235) );
  AOI211_X1 U10508 ( .C1(n9339), .C2(n9236), .A(n9660), .B(n9235), .ZN(n9338)
         );
  INV_X1 U10509 ( .A(n9237), .ZN(n9238) );
  AOI22_X1 U10510 ( .A1(n4283), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n9238), .B2(
        n9588), .ZN(n9239) );
  OAI21_X1 U10511 ( .B1(n9240), .B2(n9256), .A(n9239), .ZN(n9247) );
  XOR2_X1 U10512 ( .A(n9242), .B(n9241), .Z(n9245) );
  AOI222_X1 U10513 ( .A1(n9427), .A2(n9245), .B1(n9244), .B2(n9261), .C1(n9243), .C2(n9586), .ZN(n9341) );
  NOR2_X1 U10514 ( .A1(n9341), .A2(n4283), .ZN(n9246) );
  AOI211_X1 U10515 ( .C1(n9338), .C2(n9266), .A(n9247), .B(n9246), .ZN(n9248)
         );
  OAI21_X1 U10516 ( .B1(n9268), .B2(n9342), .A(n9248), .ZN(P1_U3274) );
  XNOR2_X1 U10517 ( .A(n9250), .B(n9249), .ZN(n9348) );
  AOI211_X1 U10518 ( .C1(n9344), .C2(n9252), .A(n9660), .B(n9251), .ZN(n9343)
         );
  INV_X1 U10519 ( .A(n9253), .ZN(n9254) );
  AOI22_X1 U10520 ( .A1(n4283), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n9254), .B2(
        n9588), .ZN(n9255) );
  OAI21_X1 U10521 ( .B1(n9257), .B2(n9256), .A(n9255), .ZN(n9265) );
  XNOR2_X1 U10522 ( .A(n9259), .B(n9258), .ZN(n9263) );
  AOI222_X1 U10523 ( .A1(n9427), .A2(n9263), .B1(n9262), .B2(n9261), .C1(n9260), .C2(n9586), .ZN(n9347) );
  NOR2_X1 U10524 ( .A1(n9347), .A2(n4283), .ZN(n9264) );
  AOI211_X1 U10525 ( .C1(n9343), .C2(n9266), .A(n9265), .B(n9264), .ZN(n9267)
         );
  OAI21_X1 U10526 ( .B1(n9268), .B2(n9348), .A(n9267), .ZN(P1_U3275) );
  MUX2_X1 U10527 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n9350), .S(n9678), .Z(
        P1_U3554) );
  NAND2_X1 U10528 ( .A1(n9273), .A2(n9572), .ZN(n9275) );
  OAI211_X1 U10529 ( .C1(n9276), .C2(n9658), .A(n9275), .B(n9274), .ZN(n9351)
         );
  MUX2_X1 U10530 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n9351), .S(n9678), .Z(
        P1_U3553) );
  OR2_X1 U10531 ( .A1(n9278), .A2(n9277), .ZN(n9608) );
  AND2_X1 U10532 ( .A1(n9279), .A2(n9608), .ZN(n9374) );
  AOI22_X1 U10533 ( .A1(n9285), .A2(n9572), .B1(n9345), .B2(n9284), .ZN(n9286)
         );
  OAI211_X1 U10534 ( .C1(n9288), .C2(n9374), .A(n9287), .B(n9286), .ZN(n9353)
         );
  MUX2_X1 U10535 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n9353), .S(n9678), .Z(
        P1_U3551) );
  AOI22_X1 U10536 ( .A1(n9290), .A2(n9572), .B1(n9345), .B2(n9289), .ZN(n9291)
         );
  OAI211_X1 U10537 ( .C1(n9293), .C2(n9374), .A(n9292), .B(n9291), .ZN(n9354)
         );
  MUX2_X1 U10538 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n9354), .S(n9678), .Z(
        P1_U3550) );
  AOI22_X1 U10539 ( .A1(n9295), .A2(n9572), .B1(n9345), .B2(n9294), .ZN(n9296)
         );
  OAI211_X1 U10540 ( .C1(n9298), .C2(n9374), .A(n9297), .B(n9296), .ZN(n9355)
         );
  MUX2_X1 U10541 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n9355), .S(n9678), .Z(
        P1_U3549) );
  AOI22_X1 U10542 ( .A1(n9300), .A2(n9572), .B1(n9345), .B2(n9299), .ZN(n9301)
         );
  OAI211_X1 U10543 ( .C1(n9303), .C2(n9374), .A(n9302), .B(n9301), .ZN(n9356)
         );
  MUX2_X1 U10544 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n9356), .S(n9678), .Z(
        P1_U3548) );
  AOI21_X1 U10545 ( .B1(n9345), .B2(n5402), .A(n9304), .ZN(n9305) );
  OAI211_X1 U10546 ( .C1(n9307), .C2(n9374), .A(n9306), .B(n9305), .ZN(n9357)
         );
  MUX2_X1 U10547 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n9357), .S(n9678), .Z(
        P1_U3547) );
  AOI22_X1 U10548 ( .A1(n9309), .A2(n9572), .B1(n9345), .B2(n9308), .ZN(n9310)
         );
  OAI211_X1 U10549 ( .C1(n9312), .C2(n9374), .A(n9311), .B(n9310), .ZN(n9358)
         );
  MUX2_X1 U10550 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n9358), .S(n9678), .Z(
        P1_U3546) );
  AOI21_X1 U10551 ( .B1(n9345), .B2(n9314), .A(n9313), .ZN(n9315) );
  OAI211_X1 U10552 ( .C1(n9317), .C2(n9374), .A(n9316), .B(n9315), .ZN(n9359)
         );
  MUX2_X1 U10553 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n9359), .S(n9678), .Z(
        P1_U3545) );
  AOI21_X1 U10554 ( .B1(n9345), .B2(n9319), .A(n9318), .ZN(n9320) );
  OAI211_X1 U10555 ( .C1(n9322), .C2(n9374), .A(n9321), .B(n9320), .ZN(n9360)
         );
  MUX2_X1 U10556 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n9360), .S(n9678), .Z(
        P1_U3544) );
  AOI21_X1 U10557 ( .B1(n9345), .B2(n9324), .A(n9323), .ZN(n9325) );
  OAI211_X1 U10558 ( .C1(n9327), .C2(n9374), .A(n9326), .B(n9325), .ZN(n9361)
         );
  MUX2_X1 U10559 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n9361), .S(n9678), .Z(
        P1_U3543) );
  AOI21_X1 U10560 ( .B1(n9345), .B2(n9329), .A(n9328), .ZN(n9330) );
  OAI211_X1 U10561 ( .C1(n9332), .C2(n9374), .A(n9331), .B(n9330), .ZN(n9362)
         );
  INV_X2 U10562 ( .A(n9676), .ZN(n9678) );
  MUX2_X1 U10563 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n9362), .S(n9678), .Z(
        P1_U3542) );
  AOI21_X1 U10564 ( .B1(n9345), .B2(n9334), .A(n9333), .ZN(n9335) );
  OAI211_X1 U10565 ( .C1(n9337), .C2(n9374), .A(n9336), .B(n9335), .ZN(n9363)
         );
  MUX2_X1 U10566 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n9363), .S(n9678), .Z(
        P1_U3541) );
  AOI21_X1 U10567 ( .B1(n9345), .B2(n9339), .A(n9338), .ZN(n9340) );
  OAI211_X1 U10568 ( .C1(n9342), .C2(n9374), .A(n9341), .B(n9340), .ZN(n9364)
         );
  MUX2_X1 U10569 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n9364), .S(n9678), .Z(
        P1_U3540) );
  AOI21_X1 U10570 ( .B1(n9345), .B2(n9344), .A(n9343), .ZN(n9346) );
  OAI211_X1 U10571 ( .C1(n9348), .C2(n9374), .A(n9347), .B(n9346), .ZN(n9365)
         );
  MUX2_X1 U10572 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n9365), .S(n9678), .Z(
        P1_U3539) );
  MUX2_X1 U10573 ( .A(P1_REG1_REG_0__SCAN_IN), .B(n9349), .S(n9678), .Z(
        P1_U3523) );
  MUX2_X1 U10574 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n9351), .S(n9470), .Z(
        P1_U3521) );
  MUX2_X1 U10575 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n9352), .S(n9470), .Z(
        P1_U3520) );
  MUX2_X1 U10576 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n9353), .S(n9470), .Z(
        P1_U3519) );
  MUX2_X1 U10577 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n9354), .S(n9470), .Z(
        P1_U3518) );
  MUX2_X1 U10578 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n9355), .S(n9470), .Z(
        P1_U3517) );
  MUX2_X1 U10579 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n9356), .S(n9470), .Z(
        P1_U3516) );
  MUX2_X1 U10580 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n9357), .S(n9470), .Z(
        P1_U3515) );
  MUX2_X1 U10581 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n9358), .S(n9470), .Z(
        P1_U3514) );
  MUX2_X1 U10582 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n9359), .S(n9470), .Z(
        P1_U3513) );
  MUX2_X1 U10583 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n9360), .S(n9470), .Z(
        P1_U3512) );
  MUX2_X1 U10584 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n9361), .S(n9470), .Z(
        P1_U3511) );
  MUX2_X1 U10585 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n9362), .S(n9470), .Z(
        P1_U3510) );
  MUX2_X1 U10586 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n9363), .S(n9470), .Z(
        P1_U3508) );
  MUX2_X1 U10587 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n9364), .S(n9470), .Z(
        P1_U3505) );
  MUX2_X1 U10588 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n9365), .S(n9470), .Z(
        P1_U3502) );
  MUX2_X1 U10589 ( .A(P1_D_REG_1__SCAN_IN), .B(n9366), .S(n9602), .Z(P1_U3441)
         );
  NOR4_X1 U10590 ( .A1(n9367), .A2(P1_IR_REG_30__SCAN_IN), .A3(P1_U3084), .A4(
        n4838), .ZN(n9368) );
  AOI21_X1 U10591 ( .B1(n9369), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n9368), .ZN(
        n9370) );
  OAI21_X1 U10592 ( .B1(n9372), .B2(n9371), .A(n9370), .ZN(P1_U3322) );
  MUX2_X1 U10593 ( .A(n9373), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3353) );
  INV_X1 U10594 ( .A(n9374), .ZN(n9664) );
  OAI21_X1 U10595 ( .B1(n9376), .B2(n9658), .A(n9375), .ZN(n9378) );
  AOI211_X1 U10596 ( .C1(n9664), .C2(n9379), .A(n9378), .B(n9377), .ZN(n9380)
         );
  AOI22_X1 U10597 ( .A1(n9470), .A2(n9380), .B1(n5145), .B2(n9666), .ZN(
        P1_U3484) );
  AOI22_X1 U10598 ( .A1(n9678), .A2(n9380), .B1(n6421), .B2(n9676), .ZN(
        P1_U3533) );
  INV_X1 U10599 ( .A(n9381), .ZN(n9816) );
  OAI22_X1 U10600 ( .A1(n9383), .A2(n4275), .B1(n9382), .B2(n9819), .ZN(n9384)
         );
  AOI21_X1 U10601 ( .B1(n9385), .B2(n9816), .A(n9384), .ZN(n9386) );
  AND2_X1 U10602 ( .A1(n9387), .A2(n9386), .ZN(n9389) );
  AOI22_X1 U10603 ( .A1(n9836), .A2(n9389), .B1(n9388), .B2(n9837), .ZN(
        P2_U3533) );
  INV_X1 U10604 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n9930) );
  AOI22_X1 U10605 ( .A1(n9828), .A2(n9389), .B1(n9930), .B2(n9827), .ZN(
        P2_U3490) );
  XNOR2_X1 U10606 ( .A(n9391), .B(n9390), .ZN(n9448) );
  OR2_X1 U10607 ( .A1(n9392), .A2(n4767), .ZN(n9393) );
  NAND2_X1 U10608 ( .A1(n9394), .A2(n9393), .ZN(n9446) );
  INV_X1 U10609 ( .A(n9446), .ZN(n9395) );
  AOI22_X1 U10610 ( .A1(n9448), .A2(n9597), .B1(n9417), .B2(n9395), .ZN(n9410)
         );
  OAI22_X1 U10611 ( .A1(n9600), .A2(n9397), .B1(n9396), .B2(n9418), .ZN(n9407)
         );
  NAND2_X1 U10612 ( .A1(n9448), .A2(n9420), .ZN(n9405) );
  OAI21_X1 U10613 ( .B1(n9400), .B2(n9399), .A(n9398), .ZN(n9403) );
  OAI22_X1 U10614 ( .A1(n9401), .A2(n9576), .B1(n9425), .B2(n9423), .ZN(n9402)
         );
  AOI21_X1 U10615 ( .B1(n9403), .B2(n9427), .A(n9402), .ZN(n9404) );
  NOR2_X1 U10616 ( .A1(n9450), .A2(n4283), .ZN(n9406) );
  AOI211_X1 U10617 ( .C1(n9434), .C2(n9408), .A(n9407), .B(n9406), .ZN(n9409)
         );
  NAND2_X1 U10618 ( .A1(n9410), .A2(n9409), .ZN(P1_U3278) );
  INV_X1 U10619 ( .A(n9411), .ZN(n9421) );
  XNOR2_X1 U10620 ( .A(n9412), .B(n9421), .ZN(n9460) );
  AND2_X1 U10621 ( .A1(n9413), .A2(n9433), .ZN(n9415) );
  OR2_X1 U10622 ( .A1(n9415), .A2(n9414), .ZN(n9458) );
  INV_X1 U10623 ( .A(n9458), .ZN(n9416) );
  AOI22_X1 U10624 ( .A1(n9460), .A2(n9597), .B1(n9417), .B2(n9416), .ZN(n9436)
         );
  OAI22_X1 U10625 ( .A1(n9600), .A2(n9550), .B1(n9419), .B2(n9418), .ZN(n9432)
         );
  NAND2_X1 U10626 ( .A1(n9460), .A2(n9420), .ZN(n9430) );
  XNOR2_X1 U10627 ( .A(n9422), .B(n9421), .ZN(n9428) );
  OAI22_X1 U10628 ( .A1(n9425), .A2(n9576), .B1(n9424), .B2(n9423), .ZN(n9426)
         );
  AOI21_X1 U10629 ( .B1(n9428), .B2(n9427), .A(n9426), .ZN(n9429) );
  AND2_X1 U10630 ( .A1(n9430), .A2(n9429), .ZN(n9462) );
  NOR2_X1 U10631 ( .A1(n9462), .A2(n4283), .ZN(n9431) );
  AOI211_X1 U10632 ( .C1(n9434), .C2(n9433), .A(n9432), .B(n9431), .ZN(n9435)
         );
  NAND2_X1 U10633 ( .A1(n9436), .A2(n9435), .ZN(P1_U3280) );
  OAI22_X1 U10634 ( .A1(n9438), .A2(n9660), .B1(n9437), .B2(n9658), .ZN(n9439)
         );
  AOI211_X1 U10635 ( .C1(n9441), .C2(n9664), .A(n9440), .B(n9439), .ZN(n9464)
         );
  AOI22_X1 U10636 ( .A1(n9678), .A2(n9464), .B1(n5247), .B2(n9676), .ZN(
        P1_U3538) );
  OAI211_X1 U10637 ( .C1(n4466), .C2(n9658), .A(n9443), .B(n9442), .ZN(n9444)
         );
  AOI21_X1 U10638 ( .B1(n9445), .B2(n9664), .A(n9444), .ZN(n9466) );
  AOI22_X1 U10639 ( .A1(n9678), .A2(n9466), .B1(n7257), .B2(n9676), .ZN(
        P1_U3537) );
  INV_X1 U10640 ( .A(n9608), .ZN(n9656) );
  OAI22_X1 U10641 ( .A1(n9446), .A2(n9660), .B1(n4767), .B2(n9658), .ZN(n9447)
         );
  AOI21_X1 U10642 ( .B1(n9448), .B2(n9656), .A(n9447), .ZN(n9449) );
  AOI22_X1 U10643 ( .A1(n9678), .A2(n9468), .B1(n5221), .B2(n9676), .ZN(
        P1_U3536) );
  NAND2_X1 U10644 ( .A1(n9452), .A2(n9451), .ZN(n9453) );
  AOI21_X1 U10645 ( .B1(n9454), .B2(n9656), .A(n9453), .ZN(n9455) );
  AND2_X1 U10646 ( .A1(n9456), .A2(n9455), .ZN(n9469) );
  AOI22_X1 U10647 ( .A1(n9678), .A2(n9469), .B1(n5184), .B2(n9676), .ZN(
        P1_U3535) );
  OAI22_X1 U10648 ( .A1(n9458), .A2(n9660), .B1(n9457), .B2(n9658), .ZN(n9459)
         );
  AOI21_X1 U10649 ( .B1(n9460), .B2(n9656), .A(n9459), .ZN(n9461) );
  AOI22_X1 U10650 ( .A1(n9678), .A2(n9471), .B1(n6422), .B2(n9676), .ZN(
        P1_U3534) );
  INV_X1 U10651 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n9463) );
  AOI22_X1 U10652 ( .A1(n9470), .A2(n9464), .B1(n9463), .B2(n9666), .ZN(
        P1_U3499) );
  INV_X1 U10653 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n9465) );
  AOI22_X1 U10654 ( .A1(n9470), .A2(n9466), .B1(n9465), .B2(n9666), .ZN(
        P1_U3496) );
  INV_X1 U10655 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n9467) );
  AOI22_X1 U10656 ( .A1(n9470), .A2(n9468), .B1(n9467), .B2(n9666), .ZN(
        P1_U3493) );
  AOI22_X1 U10657 ( .A1(n9470), .A2(n9469), .B1(n5187), .B2(n9666), .ZN(
        P1_U3490) );
  INV_X1 U10658 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n9911) );
  AOI22_X1 U10659 ( .A1(n9470), .A2(n9471), .B1(n9911), .B2(n9666), .ZN(
        P1_U3487) );
  XNOR2_X1 U10660 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  XNOR2_X1 U10661 ( .A(P1_RD_REG_SCAN_IN), .B(P2_RD_REG_SCAN_IN), .ZN(U126) );
  AOI21_X1 U10662 ( .B1(n5683), .B2(n9473), .A(n9472), .ZN(n9475) );
  XNOR2_X1 U10663 ( .A(n9475), .B(n9474), .ZN(n9476) );
  AOI22_X1 U10664 ( .A1(n9477), .A2(n9476), .B1(n9508), .B2(
        P1_ADDR_REG_0__SCAN_IN), .ZN(n9478) );
  OAI21_X1 U10665 ( .B1(P1_STATE_REG_SCAN_IN), .B2(n6758), .A(n9478), .ZN(
        P1_U3241) );
  INV_X1 U10666 ( .A(n9479), .ZN(n9483) );
  INV_X1 U10667 ( .A(n9480), .ZN(n9482) );
  OAI21_X1 U10668 ( .B1(n9483), .B2(n9482), .A(n9481), .ZN(n9485) );
  AOI22_X1 U10669 ( .A1(n9566), .A2(n9485), .B1(n9553), .B2(n9484), .ZN(n9494)
         );
  AOI21_X1 U10670 ( .B1(n9488), .B2(n9487), .A(n9486), .ZN(n9489) );
  NOR2_X1 U10671 ( .A1(n9543), .A2(n9489), .ZN(n9490) );
  AOI211_X1 U10672 ( .C1(P1_ADDR_REG_4__SCAN_IN), .C2(n9508), .A(n9491), .B(
        n9490), .ZN(n9493) );
  NAND3_X1 U10673 ( .A1(n9494), .A2(n9493), .A3(n9492), .ZN(P1_U3245) );
  INV_X1 U10674 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n10027) );
  AOI211_X1 U10675 ( .C1(n9497), .C2(n9496), .A(n9495), .B(n9522), .ZN(n9498)
         );
  AOI211_X1 U10676 ( .C1(n9553), .C2(n9500), .A(n9499), .B(n9498), .ZN(n9506)
         );
  AOI21_X1 U10677 ( .B1(n9503), .B2(n9502), .A(n9501), .ZN(n9504) );
  OR2_X1 U10678 ( .A1(n9543), .A2(n9504), .ZN(n9505) );
  OAI211_X1 U10679 ( .C1(n10027), .C2(n9571), .A(n9506), .B(n9505), .ZN(
        P1_U3246) );
  AOI22_X1 U10680 ( .A1(n9508), .A2(P1_ADDR_REG_6__SCAN_IN), .B1(n9553), .B2(
        n9507), .ZN(n9519) );
  INV_X1 U10681 ( .A(n9509), .ZN(n9518) );
  XNOR2_X1 U10682 ( .A(n9511), .B(n9510), .ZN(n9512) );
  NAND2_X1 U10683 ( .A1(n9566), .A2(n9512), .ZN(n9517) );
  OAI211_X1 U10684 ( .C1(n9515), .C2(n9514), .A(n9556), .B(n9513), .ZN(n9516)
         );
  NAND4_X1 U10685 ( .A1(n9519), .A2(n9518), .A3(n9517), .A4(n9516), .ZN(
        P1_U3247) );
  NAND2_X1 U10686 ( .A1(n9521), .A2(n9520), .ZN(n9523) );
  AOI21_X1 U10687 ( .B1(n9524), .B2(n9523), .A(n9522), .ZN(n9525) );
  AOI211_X1 U10688 ( .C1(n9553), .C2(n9527), .A(n9526), .B(n9525), .ZN(n9532)
         );
  OAI211_X1 U10689 ( .C1(n9530), .C2(n9529), .A(n9556), .B(n9528), .ZN(n9531)
         );
  OAI211_X1 U10690 ( .C1(n10035), .C2(n9571), .A(n9532), .B(n9531), .ZN(
        P1_U3250) );
  INV_X1 U10691 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n9549) );
  OAI21_X1 U10692 ( .B1(n9535), .B2(n9534), .A(n9533), .ZN(n9541) );
  INV_X1 U10693 ( .A(n9536), .ZN(n9537) );
  NOR2_X1 U10694 ( .A1(n9538), .A2(n9537), .ZN(n9539) );
  AOI211_X1 U10695 ( .C1(n9566), .C2(n9541), .A(n9540), .B(n9539), .ZN(n9548)
         );
  AOI211_X1 U10696 ( .C1(n9545), .C2(n9544), .A(n9543), .B(n9542), .ZN(n9546)
         );
  INV_X1 U10697 ( .A(n9546), .ZN(n9547) );
  OAI211_X1 U10698 ( .C1(n9549), .C2(n9571), .A(n9548), .B(n9547), .ZN(
        P1_U3251) );
  INV_X1 U10699 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n9964) );
  NOR3_X1 U10700 ( .A1(n9555), .A2(n9551), .A3(n9550), .ZN(n9554) );
  OAI21_X1 U10701 ( .B1(n9554), .B2(n9553), .A(n9552), .ZN(n9561) );
  INV_X1 U10702 ( .A(n9555), .ZN(n9559) );
  OAI211_X1 U10703 ( .C1(n9559), .C2(n9558), .A(n9557), .B(n9556), .ZN(n9560)
         );
  NAND2_X1 U10704 ( .A1(n9561), .A2(n9560), .ZN(n9568) );
  OAI21_X1 U10705 ( .B1(n9564), .B2(n9563), .A(n9562), .ZN(n9565) );
  AND2_X1 U10706 ( .A1(n9566), .A2(n9565), .ZN(n9567) );
  NOR3_X1 U10707 ( .A1(n9569), .A2(n9568), .A3(n9567), .ZN(n9570) );
  OAI21_X1 U10708 ( .B1(n9571), .B2(n9964), .A(n9570), .ZN(P1_U3252) );
  OAI211_X1 U10709 ( .C1(n9574), .C2(n9633), .A(n9573), .B(n9572), .ZN(n9632)
         );
  INV_X1 U10710 ( .A(n9575), .ZN(n9577) );
  NOR2_X1 U10711 ( .A1(n9577), .A2(n9576), .ZN(n9584) );
  AOI21_X1 U10712 ( .B1(n9580), .B2(n9579), .A(n9596), .ZN(n9582) );
  NOR3_X1 U10713 ( .A1(n4513), .A2(n9582), .A3(n9581), .ZN(n9583) );
  AOI211_X1 U10714 ( .C1(n9586), .C2(n9585), .A(n9584), .B(n9583), .ZN(n9634)
         );
  AOI22_X1 U10715 ( .A1(n9590), .A2(n9589), .B1(n9588), .B2(n9587), .ZN(n9591)
         );
  OAI211_X1 U10716 ( .C1(n9592), .C2(n9632), .A(n9634), .B(n9591), .ZN(n9598)
         );
  INV_X1 U10717 ( .A(n9593), .ZN(n9594) );
  AOI21_X1 U10718 ( .B1(n9596), .B2(n9595), .A(n9594), .ZN(n9637) );
  AOI22_X1 U10719 ( .A1(n9598), .A2(n9600), .B1(n9637), .B2(n9597), .ZN(n9599)
         );
  OAI21_X1 U10720 ( .B1(n6271), .B2(n9600), .A(n9599), .ZN(P1_U3286) );
  AND2_X1 U10721 ( .A1(n9602), .A2(n9601), .ZN(n9604) );
  AND2_X1 U10722 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n9603), .ZN(P1_U3292) );
  AND2_X1 U10723 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n9603), .ZN(P1_U3293) );
  AND2_X1 U10724 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n9603), .ZN(P1_U3294) );
  AND2_X1 U10725 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n9603), .ZN(P1_U3295) );
  AND2_X1 U10726 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n9603), .ZN(P1_U3296) );
  AND2_X1 U10727 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n9603), .ZN(P1_U3297) );
  AND2_X1 U10728 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n9603), .ZN(P1_U3298) );
  AND2_X1 U10729 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n9603), .ZN(P1_U3299) );
  AND2_X1 U10730 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n9603), .ZN(P1_U3300) );
  AND2_X1 U10731 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n9603), .ZN(P1_U3301) );
  AND2_X1 U10732 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n9603), .ZN(P1_U3302) );
  AND2_X1 U10733 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n9603), .ZN(P1_U3303) );
  AND2_X1 U10734 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n9603), .ZN(P1_U3304) );
  AND2_X1 U10735 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n9603), .ZN(P1_U3305) );
  AND2_X1 U10736 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n9603), .ZN(P1_U3306) );
  AND2_X1 U10737 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n9603), .ZN(P1_U3307) );
  AND2_X1 U10738 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n9603), .ZN(P1_U3308) );
  AND2_X1 U10739 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n9603), .ZN(P1_U3309) );
  NOR2_X1 U10740 ( .A1(n9604), .A2(n9944), .ZN(P1_U3310) );
  AND2_X1 U10741 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n9603), .ZN(P1_U3311) );
  AND2_X1 U10742 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n9603), .ZN(P1_U3312) );
  AND2_X1 U10743 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n9603), .ZN(P1_U3313) );
  AND2_X1 U10744 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n9603), .ZN(P1_U3314) );
  NOR2_X1 U10745 ( .A1(n9604), .A2(n9979), .ZN(P1_U3315) );
  NOR2_X1 U10746 ( .A1(n9604), .A2(n9913), .ZN(P1_U3316) );
  AND2_X1 U10747 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n9603), .ZN(P1_U3317) );
  AND2_X1 U10748 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n9603), .ZN(P1_U3318) );
  AND2_X1 U10749 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n9603), .ZN(P1_U3319) );
  AND2_X1 U10750 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n9603), .ZN(P1_U3320) );
  NOR2_X1 U10751 ( .A1(n9604), .A2(n9898), .ZN(P1_U3321) );
  INV_X1 U10752 ( .A(n9605), .ZN(n9606) );
  OAI211_X1 U10753 ( .C1(n9609), .C2(n9608), .A(n9607), .B(n9606), .ZN(n9610)
         );
  NOR2_X1 U10754 ( .A1(n9611), .A2(n9610), .ZN(n9668) );
  AOI22_X1 U10755 ( .A1(n9470), .A2(n9668), .B1(n4999), .B2(n9666), .ZN(
        P1_U3457) );
  OAI22_X1 U10756 ( .A1(n9613), .A2(n9660), .B1(n9612), .B2(n9658), .ZN(n9615)
         );
  AOI211_X1 U10757 ( .C1(n9656), .C2(n9616), .A(n9615), .B(n9614), .ZN(n9669)
         );
  AOI22_X1 U10758 ( .A1(n9470), .A2(n9669), .B1(n5018), .B2(n9666), .ZN(
        P1_U3460) );
  INV_X1 U10759 ( .A(n9617), .ZN(n9623) );
  OAI22_X1 U10760 ( .A1(n9619), .A2(n9660), .B1(n9618), .B2(n9658), .ZN(n9620)
         );
  AOI21_X1 U10761 ( .B1(n9621), .B2(n9664), .A(n9620), .ZN(n9622) );
  AND2_X1 U10762 ( .A1(n9623), .A2(n9622), .ZN(n9670) );
  INV_X1 U10763 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n9624) );
  AOI22_X1 U10764 ( .A1(n9470), .A2(n9670), .B1(n9624), .B2(n9666), .ZN(
        P1_U3463) );
  INV_X1 U10765 ( .A(n9625), .ZN(n9626) );
  AND2_X1 U10766 ( .A1(n9626), .A2(n9656), .ZN(n9630) );
  OAI22_X1 U10767 ( .A1(n9628), .A2(n9660), .B1(n9627), .B2(n9658), .ZN(n9629)
         );
  NOR3_X1 U10768 ( .A1(n9631), .A2(n9630), .A3(n9629), .ZN(n9671) );
  INV_X1 U10769 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n9903) );
  AOI22_X1 U10770 ( .A1(n9470), .A2(n9671), .B1(n9903), .B2(n9666), .ZN(
        P1_U3466) );
  OAI21_X1 U10771 ( .B1(n9633), .B2(n9658), .A(n9632), .ZN(n9636) );
  INV_X1 U10772 ( .A(n9634), .ZN(n9635) );
  AOI211_X1 U10773 ( .C1(n9637), .C2(n9664), .A(n9636), .B(n9635), .ZN(n9672)
         );
  AOI22_X1 U10774 ( .A1(n9470), .A2(n9672), .B1(n5067), .B2(n9666), .ZN(
        P1_U3469) );
  INV_X1 U10775 ( .A(n9638), .ZN(n9643) );
  OAI22_X1 U10776 ( .A1(n9640), .A2(n9660), .B1(n9639), .B2(n9658), .ZN(n9642)
         );
  AOI211_X1 U10777 ( .C1(n9656), .C2(n9643), .A(n9642), .B(n9641), .ZN(n9673)
         );
  AOI22_X1 U10778 ( .A1(n9470), .A2(n9673), .B1(n5080), .B2(n9666), .ZN(
        P1_U3472) );
  OAI211_X1 U10779 ( .C1(n9646), .C2(n9658), .A(n9645), .B(n9644), .ZN(n9647)
         );
  AOI21_X1 U10780 ( .B1(n9664), .B2(n9648), .A(n9647), .ZN(n9674) );
  INV_X1 U10781 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n9649) );
  AOI22_X1 U10782 ( .A1(n9470), .A2(n9674), .B1(n9649), .B2(n9666), .ZN(
        P1_U3475) );
  INV_X1 U10783 ( .A(n9650), .ZN(n9655) );
  OAI21_X1 U10784 ( .B1(n9652), .B2(n9660), .A(n9651), .ZN(n9654) );
  AOI211_X1 U10785 ( .C1(n9656), .C2(n9655), .A(n9654), .B(n9653), .ZN(n9675)
         );
  INV_X1 U10786 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n9657) );
  AOI22_X1 U10787 ( .A1(n9470), .A2(n9675), .B1(n9657), .B2(n9666), .ZN(
        P1_U3478) );
  OAI22_X1 U10788 ( .A1(n9661), .A2(n9660), .B1(n9659), .B2(n9658), .ZN(n9663)
         );
  AOI211_X1 U10789 ( .C1(n9665), .C2(n9664), .A(n9663), .B(n9662), .ZN(n9677)
         );
  INV_X1 U10790 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n9667) );
  AOI22_X1 U10791 ( .A1(n9470), .A2(n9677), .B1(n9667), .B2(n9666), .ZN(
        P1_U3481) );
  AOI22_X1 U10792 ( .A1(n9678), .A2(n9668), .B1(n6288), .B2(n9676), .ZN(
        P1_U3524) );
  AOI22_X1 U10793 ( .A1(n9678), .A2(n9669), .B1(n6287), .B2(n9676), .ZN(
        P1_U3525) );
  AOI22_X1 U10794 ( .A1(n9678), .A2(n9670), .B1(n6293), .B2(n9676), .ZN(
        P1_U3526) );
  AOI22_X1 U10795 ( .A1(n9678), .A2(n9671), .B1(n5050), .B2(n9676), .ZN(
        P1_U3527) );
  AOI22_X1 U10796 ( .A1(n9678), .A2(n9672), .B1(n5066), .B2(n9676), .ZN(
        P1_U3528) );
  AOI22_X1 U10797 ( .A1(n9678), .A2(n9673), .B1(n5082), .B2(n9676), .ZN(
        P1_U3529) );
  AOI22_X1 U10798 ( .A1(n9678), .A2(n9674), .B1(n5098), .B2(n9676), .ZN(
        P1_U3530) );
  AOI22_X1 U10799 ( .A1(n9678), .A2(n9675), .B1(n6418), .B2(n9676), .ZN(
        P1_U3531) );
  AOI22_X1 U10800 ( .A1(n9678), .A2(n9677), .B1(n5133), .B2(n9676), .ZN(
        P1_U3532) );
  AOI22_X1 U10801 ( .A1(n9744), .A2(P2_REG2_REG_0__SCAN_IN), .B1(
        P2_REG1_REG_0__SCAN_IN), .B2(n9748), .ZN(n9686) );
  AOI21_X1 U10802 ( .B1(n9741), .B2(P2_ADDR_REG_0__SCAN_IN), .A(n9679), .ZN(
        n9685) );
  OAI21_X1 U10803 ( .B1(P2_REG1_REG_0__SCAN_IN), .B2(n9681), .A(n9680), .ZN(
        n9683) );
  NOR2_X1 U10804 ( .A1(n9692), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n9682) );
  OAI21_X1 U10805 ( .B1(n9683), .B2(n9682), .A(P2_IR_REG_0__SCAN_IN), .ZN(
        n9684) );
  OAI211_X1 U10806 ( .C1(P2_IR_REG_0__SCAN_IN), .C2(n9686), .A(n9685), .B(
        n9684), .ZN(P2_U3245) );
  AOI22_X1 U10807 ( .A1(n9741), .A2(P2_ADDR_REG_3__SCAN_IN), .B1(
        P2_REG3_REG_3__SCAN_IN), .B2(P2_U3152), .ZN(n9700) );
  NAND2_X1 U10808 ( .A1(n9747), .A2(n9688), .ZN(n9699) );
  OAI211_X1 U10809 ( .C1(n9691), .C2(n9690), .A(n9748), .B(n9689), .ZN(n9698)
         );
  AOI211_X1 U10810 ( .C1(n9695), .C2(n9694), .A(n9693), .B(n9692), .ZN(n9696)
         );
  INV_X1 U10811 ( .A(n9696), .ZN(n9697) );
  NAND4_X1 U10812 ( .A1(n9700), .A2(n9699), .A3(n9698), .A4(n9697), .ZN(
        P2_U3248) );
  INV_X1 U10813 ( .A(n9701), .ZN(n9702) );
  AOI21_X1 U10814 ( .B1(n9741), .B2(P2_ADDR_REG_6__SCAN_IN), .A(n9702), .ZN(
        n9712) );
  NAND2_X1 U10815 ( .A1(n9747), .A2(n9703), .ZN(n9711) );
  OAI211_X1 U10816 ( .C1(n9706), .C2(n9705), .A(n9748), .B(n9704), .ZN(n9710)
         );
  OAI211_X1 U10817 ( .C1(n4346), .C2(n4441), .A(n9744), .B(n9708), .ZN(n9709)
         );
  NAND4_X1 U10818 ( .A1(n9712), .A2(n9711), .A3(n9710), .A4(n9709), .ZN(
        P2_U3251) );
  INV_X1 U10819 ( .A(n9713), .ZN(n9714) );
  AOI21_X1 U10820 ( .B1(n9741), .B2(P2_ADDR_REG_7__SCAN_IN), .A(n9714), .ZN(
        n9725) );
  NAND2_X1 U10821 ( .A1(n9747), .A2(n9715), .ZN(n9724) );
  OAI211_X1 U10822 ( .C1(n9718), .C2(n9717), .A(n9748), .B(n9716), .ZN(n9723)
         );
  OAI211_X1 U10823 ( .C1(n9721), .C2(n9720), .A(n9744), .B(n9719), .ZN(n9722)
         );
  NAND4_X1 U10824 ( .A1(n9725), .A2(n9724), .A3(n9723), .A4(n9722), .ZN(
        P2_U3252) );
  INV_X1 U10825 ( .A(n9726), .ZN(n9727) );
  AOI21_X1 U10826 ( .B1(n9741), .B2(P2_ADDR_REG_10__SCAN_IN), .A(n9727), .ZN(
        n9738) );
  NAND2_X1 U10827 ( .A1(n9747), .A2(n9728), .ZN(n9737) );
  OAI211_X1 U10828 ( .C1(n9731), .C2(n9730), .A(n9729), .B(n9748), .ZN(n9736)
         );
  OAI211_X1 U10829 ( .C1(n9734), .C2(n9733), .A(n9744), .B(n9732), .ZN(n9735)
         );
  NAND4_X1 U10830 ( .A1(n9738), .A2(n9737), .A3(n9736), .A4(n9735), .ZN(
        P2_U3255) );
  INV_X1 U10831 ( .A(n9739), .ZN(n9740) );
  AOI21_X1 U10832 ( .B1(n9741), .B2(P2_ADDR_REG_17__SCAN_IN), .A(n9740), .ZN(
        n9755) );
  XOR2_X1 U10833 ( .A(n9743), .B(n9742), .Z(n9745) );
  NAND2_X1 U10834 ( .A1(n9745), .A2(n9744), .ZN(n9754) );
  NAND2_X1 U10835 ( .A1(n9747), .A2(n9746), .ZN(n9753) );
  OAI211_X1 U10836 ( .C1(n9751), .C2(n9750), .A(n9749), .B(n9748), .ZN(n9752)
         );
  NAND4_X1 U10837 ( .A1(n9755), .A2(n9754), .A3(n9753), .A4(n9752), .ZN(
        P2_U3262) );
  XNOR2_X1 U10838 ( .A(n9756), .B(n8342), .ZN(n9758) );
  AOI21_X1 U10839 ( .B1(n9759), .B2(n9758), .A(n9757), .ZN(n9787) );
  AOI22_X1 U10840 ( .A1(P2_REG2_REG_1__SCAN_IN), .A2(n9772), .B1(
        P2_REG3_REG_1__SCAN_IN), .B2(n9760), .ZN(n9771) );
  XNOR2_X1 U10841 ( .A(n9785), .B(n9761), .ZN(n9784) );
  NAND2_X1 U10842 ( .A1(n9762), .A2(n9784), .ZN(n9767) );
  OAI21_X1 U10843 ( .B1(n8342), .B2(n9764), .A(n9763), .ZN(n9790) );
  NAND2_X1 U10844 ( .A1(n9765), .A2(n9790), .ZN(n9766) );
  OAI211_X1 U10845 ( .C1(n9785), .C2(n9768), .A(n9767), .B(n9766), .ZN(n9769)
         );
  INV_X1 U10846 ( .A(n9769), .ZN(n9770) );
  OAI211_X1 U10847 ( .C1(n9772), .C2(n9787), .A(n9771), .B(n9770), .ZN(
        P2_U3295) );
  NAND2_X1 U10848 ( .A1(n9774), .A2(n9773), .ZN(n9780) );
  AND2_X1 U10849 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n9780), .ZN(P2_U3297) );
  AND2_X1 U10850 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n9780), .ZN(P2_U3298) );
  AND2_X1 U10851 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n9780), .ZN(P2_U3299) );
  AND2_X1 U10852 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n9780), .ZN(P2_U3300) );
  AND2_X1 U10853 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n9780), .ZN(P2_U3301) );
  AND2_X1 U10854 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n9780), .ZN(P2_U3302) );
  AND2_X1 U10855 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n9780), .ZN(P2_U3303) );
  AND2_X1 U10856 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n9780), .ZN(P2_U3304) );
  AND2_X1 U10857 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n9780), .ZN(P2_U3305) );
  AND2_X1 U10858 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n9780), .ZN(P2_U3306) );
  AND2_X1 U10859 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n9780), .ZN(P2_U3307) );
  AND2_X1 U10860 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n9780), .ZN(P2_U3308) );
  AND2_X1 U10861 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n9780), .ZN(P2_U3309) );
  AND2_X1 U10862 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n9780), .ZN(P2_U3310) );
  AND2_X1 U10863 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n9780), .ZN(P2_U3311) );
  AND2_X1 U10864 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n9780), .ZN(P2_U3312) );
  AND2_X1 U10865 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n9780), .ZN(P2_U3313) );
  AND2_X1 U10866 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n9780), .ZN(P2_U3314) );
  AND2_X1 U10867 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n9780), .ZN(P2_U3315) );
  AND2_X1 U10868 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n9780), .ZN(P2_U3316) );
  AND2_X1 U10869 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n9780), .ZN(P2_U3317) );
  INV_X1 U10870 ( .A(n9780), .ZN(n9775) );
  NOR2_X1 U10871 ( .A1(n9775), .A2(n10006), .ZN(P2_U3318) );
  AND2_X1 U10872 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n9780), .ZN(P2_U3319) );
  NOR2_X1 U10873 ( .A1(n9775), .A2(n9905), .ZN(P2_U3320) );
  NOR2_X1 U10874 ( .A1(n9775), .A2(n9958), .ZN(P2_U3321) );
  AND2_X1 U10875 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n9780), .ZN(P2_U3322) );
  AND2_X1 U10876 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n9780), .ZN(P2_U3323) );
  AND2_X1 U10877 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n9780), .ZN(P2_U3324) );
  NOR2_X1 U10878 ( .A1(n9775), .A2(n9920), .ZN(P2_U3325) );
  AND2_X1 U10879 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n9780), .ZN(P2_U3326) );
  INV_X1 U10880 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n9776) );
  AOI22_X1 U10881 ( .A1(n9783), .A2(n9777), .B1(n9776), .B2(n9780), .ZN(
        P2_U3437) );
  NOR2_X1 U10882 ( .A1(n9779), .A2(n9778), .ZN(n9782) );
  INV_X1 U10883 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n9781) );
  AOI22_X1 U10884 ( .A1(n9783), .A2(n9782), .B1(n9781), .B2(n9780), .ZN(
        P2_U3438) );
  INV_X1 U10885 ( .A(n9784), .ZN(n9786) );
  OAI22_X1 U10886 ( .A1(n9786), .A2(n4275), .B1(n9785), .B2(n9819), .ZN(n9789)
         );
  INV_X1 U10887 ( .A(n9787), .ZN(n9788) );
  AOI211_X1 U10888 ( .C1(n9825), .C2(n9790), .A(n9789), .B(n9788), .ZN(n9829)
         );
  INV_X1 U10889 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n9791) );
  AOI22_X1 U10890 ( .A1(n9828), .A2(n9829), .B1(n9791), .B2(n9827), .ZN(
        P2_U3454) );
  OAI22_X1 U10891 ( .A1(n9793), .A2(n4275), .B1(n9792), .B2(n9819), .ZN(n9795)
         );
  AOI211_X1 U10892 ( .C1(n9816), .C2(n9796), .A(n9795), .B(n9794), .ZN(n9830)
         );
  INV_X1 U10893 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n9797) );
  AOI22_X1 U10894 ( .A1(n9828), .A2(n9830), .B1(n9797), .B2(n9827), .ZN(
        P2_U3460) );
  NOR2_X1 U10895 ( .A1(n9799), .A2(n9798), .ZN(n9803) );
  OAI21_X1 U10896 ( .B1(n6748), .B2(n9819), .A(n9800), .ZN(n9801) );
  NOR3_X1 U10897 ( .A1(n9803), .A2(n9802), .A3(n9801), .ZN(n9832) );
  INV_X1 U10898 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n9804) );
  AOI22_X1 U10899 ( .A1(n9828), .A2(n9832), .B1(n9804), .B2(n9827), .ZN(
        P2_U3466) );
  OAI211_X1 U10900 ( .C1(n9807), .C2(n9819), .A(n9806), .B(n9805), .ZN(n9808)
         );
  AOI21_X1 U10901 ( .B1(n9825), .B2(n9809), .A(n9808), .ZN(n9833) );
  INV_X1 U10902 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n9810) );
  AOI22_X1 U10903 ( .A1(n9828), .A2(n9833), .B1(n9810), .B2(n9827), .ZN(
        P2_U3472) );
  OAI22_X1 U10904 ( .A1(n9812), .A2(n4275), .B1(n9811), .B2(n9819), .ZN(n9814)
         );
  AOI211_X1 U10905 ( .C1(n9816), .C2(n9815), .A(n9814), .B(n9813), .ZN(n9835)
         );
  INV_X1 U10906 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n9817) );
  AOI22_X1 U10907 ( .A1(n9828), .A2(n9835), .B1(n9817), .B2(n9827), .ZN(
        P2_U3478) );
  INV_X1 U10908 ( .A(n9818), .ZN(n9820) );
  OAI22_X1 U10909 ( .A1(n9822), .A2(n4275), .B1(n9820), .B2(n9819), .ZN(n9824)
         );
  AOI211_X1 U10910 ( .C1(n9826), .C2(n9825), .A(n9824), .B(n9823), .ZN(n9839)
         );
  INV_X1 U10911 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n9917) );
  AOI22_X1 U10912 ( .A1(n9828), .A2(n9839), .B1(n9917), .B2(n9827), .ZN(
        P2_U3484) );
  AOI22_X1 U10913 ( .A1(n9836), .A2(n9829), .B1(n5742), .B2(n9837), .ZN(
        P2_U3521) );
  AOI22_X1 U10914 ( .A1(n9836), .A2(n9830), .B1(n6484), .B2(n9837), .ZN(
        P2_U3523) );
  AOI22_X1 U10915 ( .A1(n9836), .A2(n9832), .B1(n9831), .B2(n9837), .ZN(
        P2_U3525) );
  AOI22_X1 U10916 ( .A1(n9836), .A2(n9833), .B1(n6508), .B2(n9837), .ZN(
        P2_U3527) );
  AOI22_X1 U10917 ( .A1(n9836), .A2(n9835), .B1(n9834), .B2(n9837), .ZN(
        P2_U3529) );
  AOI22_X1 U10918 ( .A1(n9840), .A2(n9839), .B1(n9838), .B2(n9837), .ZN(
        P2_U3531) );
  INV_X1 U10919 ( .A(n9841), .ZN(n9842) );
  NAND2_X1 U10920 ( .A1(n9843), .A2(n9842), .ZN(n9844) );
  XNOR2_X1 U10921 ( .A(P2_ADDR_REG_1__SCAN_IN), .B(n9844), .ZN(ADD_1071_U5) );
  XOR2_X1 U10922 ( .A(P1_ADDR_REG_0__SCAN_IN), .B(P2_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1071_U46) );
  OAI21_X1 U10923 ( .B1(n9847), .B2(n9846), .A(n9845), .ZN(ADD_1071_U56) );
  OAI21_X1 U10924 ( .B1(n9850), .B2(n9849), .A(n9848), .ZN(ADD_1071_U57) );
  OAI21_X1 U10925 ( .B1(n9853), .B2(n9852), .A(n9851), .ZN(ADD_1071_U58) );
  OAI21_X1 U10926 ( .B1(n9856), .B2(n9855), .A(n9854), .ZN(ADD_1071_U59) );
  OAI21_X1 U10927 ( .B1(n9859), .B2(n9858), .A(n9857), .ZN(ADD_1071_U60) );
  OAI21_X1 U10928 ( .B1(n9862), .B2(n9861), .A(n9860), .ZN(ADD_1071_U61) );
  AOI21_X1 U10929 ( .B1(n9865), .B2(n9864), .A(n9863), .ZN(ADD_1071_U62) );
  AOI21_X1 U10930 ( .B1(n9868), .B2(n9867), .A(n9866), .ZN(ADD_1071_U63) );
  NAND2_X1 U10931 ( .A1(keyinput18), .A2(keyinput30), .ZN(n9874) );
  NOR2_X1 U10932 ( .A1(keyinput52), .A2(keyinput47), .ZN(n9872) );
  NAND3_X1 U10933 ( .A1(keyinput32), .A2(keyinput36), .A3(keyinput25), .ZN(
        n9870) );
  NAND3_X1 U10934 ( .A1(keyinput39), .A2(keyinput46), .A3(keyinput54), .ZN(
        n9869) );
  NOR4_X1 U10935 ( .A1(keyinput21), .A2(keyinput5), .A3(n9870), .A4(n9869), 
        .ZN(n9871) );
  NAND4_X1 U10936 ( .A1(keyinput0), .A2(keyinput7), .A3(n9872), .A4(n9871), 
        .ZN(n9873) );
  NOR4_X1 U10937 ( .A1(keyinput40), .A2(keyinput6), .A3(n9874), .A4(n9873), 
        .ZN(n10019) );
  NAND3_X1 U10938 ( .A1(keyinput8), .A2(keyinput41), .A3(keyinput3), .ZN(n9895) );
  NOR3_X1 U10939 ( .A1(keyinput62), .A2(keyinput15), .A3(keyinput63), .ZN(
        n9878) );
  NOR4_X1 U10940 ( .A1(keyinput42), .A2(keyinput49), .A3(keyinput48), .A4(
        keyinput61), .ZN(n9877) );
  NAND2_X1 U10941 ( .A1(keyinput56), .A2(keyinput43), .ZN(n9875) );
  NOR3_X1 U10942 ( .A1(keyinput45), .A2(keyinput4), .A3(n9875), .ZN(n9876) );
  NAND4_X1 U10943 ( .A1(keyinput1), .A2(n9878), .A3(n9877), .A4(n9876), .ZN(
        n9894) );
  NOR3_X1 U10944 ( .A1(keyinput13), .A2(keyinput20), .A3(keyinput59), .ZN(
        n9892) );
  NAND3_X1 U10945 ( .A1(keyinput44), .A2(keyinput50), .A3(keyinput27), .ZN(
        n9883) );
  NOR2_X1 U10946 ( .A1(keyinput17), .A2(keyinput26), .ZN(n9879) );
  NAND3_X1 U10947 ( .A1(keyinput28), .A2(keyinput58), .A3(n9879), .ZN(n9882)
         );
  NOR2_X1 U10948 ( .A1(keyinput14), .A2(keyinput37), .ZN(n9880) );
  NAND3_X1 U10949 ( .A1(keyinput9), .A2(keyinput57), .A3(n9880), .ZN(n9881) );
  NOR4_X1 U10950 ( .A1(keyinput60), .A2(n9883), .A3(n9882), .A4(n9881), .ZN(
        n9891) );
  INV_X1 U10951 ( .A(keyinput16), .ZN(n9884) );
  NAND3_X1 U10952 ( .A1(keyinput24), .A2(keyinput53), .A3(n9884), .ZN(n9889)
         );
  NAND4_X1 U10953 ( .A1(keyinput11), .A2(keyinput23), .A3(keyinput19), .A4(
        keyinput33), .ZN(n9888) );
  NOR3_X1 U10954 ( .A1(keyinput55), .A2(keyinput51), .A3(keyinput12), .ZN(
        n9886) );
  NOR3_X1 U10955 ( .A1(keyinput34), .A2(keyinput2), .A3(keyinput38), .ZN(n9885) );
  NAND4_X1 U10956 ( .A1(keyinput22), .A2(n9886), .A3(keyinput35), .A4(n9885), 
        .ZN(n9887) );
  NOR4_X1 U10957 ( .A1(keyinput10), .A2(n9889), .A3(n9888), .A4(n9887), .ZN(
        n9890) );
  NAND4_X1 U10958 ( .A1(keyinput31), .A2(n9892), .A3(n9891), .A4(n9890), .ZN(
        n9893) );
  NOR4_X1 U10959 ( .A1(keyinput29), .A2(n9895), .A3(n9894), .A4(n9893), .ZN(
        n10018) );
  AOI22_X1 U10960 ( .A1(n9898), .A2(keyinput32), .B1(keyinput36), .B2(n9897), 
        .ZN(n9896) );
  OAI221_X1 U10961 ( .B1(n9898), .B2(keyinput32), .C1(n9897), .C2(keyinput36), 
        .A(n9896), .ZN(n9909) );
  AOI22_X1 U10962 ( .A1(n9901), .A2(keyinput25), .B1(keyinput21), .B2(n9900), 
        .ZN(n9899) );
  OAI221_X1 U10963 ( .B1(n9901), .B2(keyinput25), .C1(n9900), .C2(keyinput21), 
        .A(n9899), .ZN(n9908) );
  AOI22_X1 U10964 ( .A1(n9903), .A2(keyinput18), .B1(n5098), .B2(keyinput40), 
        .ZN(n9902) );
  OAI221_X1 U10965 ( .B1(n9903), .B2(keyinput18), .C1(n5098), .C2(keyinput40), 
        .A(n9902), .ZN(n9907) );
  AOI22_X1 U10966 ( .A1(n9905), .A2(keyinput30), .B1(n5080), .B2(keyinput6), 
        .ZN(n9904) );
  OAI221_X1 U10967 ( .B1(n9905), .B2(keyinput30), .C1(n5080), .C2(keyinput6), 
        .A(n9904), .ZN(n9906) );
  NOR4_X1 U10968 ( .A1(n9909), .A2(n9908), .A3(n9907), .A4(n9906), .ZN(n9956)
         );
  AOI22_X1 U10969 ( .A1(n6585), .A2(keyinput52), .B1(n9911), .B2(keyinput0), 
        .ZN(n9910) );
  OAI221_X1 U10970 ( .B1(n6585), .B2(keyinput52), .C1(n9911), .C2(keyinput0), 
        .A(n9910), .ZN(n9924) );
  AOI22_X1 U10971 ( .A1(n9914), .A2(keyinput7), .B1(n9913), .B2(keyinput47), 
        .ZN(n9912) );
  OAI221_X1 U10972 ( .B1(n9914), .B2(keyinput7), .C1(n9913), .C2(keyinput47), 
        .A(n9912), .ZN(n9923) );
  INV_X1 U10973 ( .A(SI_7_), .ZN(n9916) );
  AOI22_X1 U10974 ( .A1(n9917), .A2(keyinput5), .B1(n9916), .B2(keyinput39), 
        .ZN(n9915) );
  OAI221_X1 U10975 ( .B1(n9917), .B2(keyinput5), .C1(n9916), .C2(keyinput39), 
        .A(n9915), .ZN(n9922) );
  INV_X1 U10976 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n9919) );
  AOI22_X1 U10977 ( .A1(n9920), .A2(keyinput46), .B1(n9919), .B2(keyinput54), 
        .ZN(n9918) );
  OAI221_X1 U10978 ( .B1(n9920), .B2(keyinput46), .C1(n9919), .C2(keyinput54), 
        .A(n9918), .ZN(n9921) );
  NOR4_X1 U10979 ( .A1(n9924), .A2(n9923), .A3(n9922), .A4(n9921), .ZN(n9955)
         );
  INV_X1 U10980 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n9927) );
  AOI22_X1 U10981 ( .A1(n9927), .A2(keyinput42), .B1(keyinput49), .B2(n9926), 
        .ZN(n9925) );
  OAI221_X1 U10982 ( .B1(n9927), .B2(keyinput42), .C1(n9926), .C2(keyinput49), 
        .A(n9925), .ZN(n9939) );
  AOI22_X1 U10983 ( .A1(n9930), .A2(keyinput63), .B1(n9929), .B2(keyinput1), 
        .ZN(n9928) );
  OAI221_X1 U10984 ( .B1(n9930), .B2(keyinput63), .C1(n9929), .C2(keyinput1), 
        .A(n9928), .ZN(n9938) );
  AOI22_X1 U10985 ( .A1(n9933), .A2(keyinput62), .B1(n9932), .B2(keyinput15), 
        .ZN(n9931) );
  OAI221_X1 U10986 ( .B1(n9933), .B2(keyinput62), .C1(n9932), .C2(keyinput15), 
        .A(n9931), .ZN(n9937) );
  XOR2_X1 U10987 ( .A(n6105), .B(keyinput61), .Z(n9935) );
  XNOR2_X1 U10988 ( .A(P1_IR_REG_13__SCAN_IN), .B(keyinput48), .ZN(n9934) );
  NAND2_X1 U10989 ( .A1(n9935), .A2(n9934), .ZN(n9936) );
  NOR4_X1 U10990 ( .A1(n9939), .A2(n9938), .A3(n9937), .A4(n9936), .ZN(n9954)
         );
  AOI22_X1 U10991 ( .A1(n9941), .A2(keyinput45), .B1(keyinput43), .B2(n6421), 
        .ZN(n9940) );
  OAI221_X1 U10992 ( .B1(n9941), .B2(keyinput45), .C1(n6421), .C2(keyinput43), 
        .A(n9940), .ZN(n9952) );
  AOI22_X1 U10993 ( .A1(n9944), .A2(keyinput4), .B1(keyinput56), .B2(n9943), 
        .ZN(n9942) );
  OAI221_X1 U10994 ( .B1(n9944), .B2(keyinput4), .C1(n9943), .C2(keyinput56), 
        .A(n9942), .ZN(n9951) );
  AOI22_X1 U10995 ( .A1(n8627), .A2(keyinput41), .B1(n9946), .B2(keyinput3), 
        .ZN(n9945) );
  OAI221_X1 U10996 ( .B1(n8627), .B2(keyinput41), .C1(n9946), .C2(keyinput3), 
        .A(n9945), .ZN(n9950) );
  XOR2_X1 U10997 ( .A(n8016), .B(keyinput29), .Z(n9948) );
  XNOR2_X1 U10998 ( .A(P1_IR_REG_28__SCAN_IN), .B(keyinput8), .ZN(n9947) );
  NAND2_X1 U10999 ( .A1(n9948), .A2(n9947), .ZN(n9949) );
  NOR4_X1 U11000 ( .A1(n9952), .A2(n9951), .A3(n9950), .A4(n9949), .ZN(n9953)
         );
  NAND4_X1 U11001 ( .A1(n9956), .A2(n9955), .A3(n9954), .A4(n9953), .ZN(n10017) );
  INV_X1 U11002 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n9959) );
  AOI22_X1 U11003 ( .A1(n9959), .A2(keyinput31), .B1(keyinput59), .B2(n9958), 
        .ZN(n9957) );
  OAI221_X1 U11004 ( .B1(n9959), .B2(keyinput31), .C1(n9958), .C2(keyinput59), 
        .A(n9957), .ZN(n9970) );
  AOI22_X1 U11005 ( .A1(n9961), .A2(keyinput13), .B1(keyinput20), .B2(n5937), 
        .ZN(n9960) );
  OAI221_X1 U11006 ( .B1(n9961), .B2(keyinput13), .C1(n5937), .C2(keyinput20), 
        .A(n9960), .ZN(n9969) );
  INV_X1 U11007 ( .A(SI_14_), .ZN(n9963) );
  AOI22_X1 U11008 ( .A1(n9964), .A2(keyinput37), .B1(n9963), .B2(keyinput57), 
        .ZN(n9962) );
  OAI221_X1 U11009 ( .B1(n9964), .B2(keyinput37), .C1(n9963), .C2(keyinput57), 
        .A(n9962), .ZN(n9968) );
  AOI22_X1 U11010 ( .A1(n6497), .A2(keyinput14), .B1(keyinput9), .B2(n9966), 
        .ZN(n9965) );
  OAI221_X1 U11011 ( .B1(n6497), .B2(keyinput14), .C1(n9966), .C2(keyinput9), 
        .A(n9965), .ZN(n9967) );
  NOR4_X1 U11012 ( .A1(n9970), .A2(n9969), .A3(n9968), .A4(n9967), .ZN(n10015)
         );
  AOI22_X1 U11013 ( .A1(n9972), .A2(keyinput60), .B1(keyinput27), .B2(n6539), 
        .ZN(n9971) );
  OAI221_X1 U11014 ( .B1(n9972), .B2(keyinput60), .C1(n6539), .C2(keyinput27), 
        .A(n9971), .ZN(n9983) );
  AOI22_X1 U11015 ( .A1(n9975), .A2(keyinput44), .B1(keyinput50), .B2(n9974), 
        .ZN(n9973) );
  OAI221_X1 U11016 ( .B1(n9975), .B2(keyinput44), .C1(n9974), .C2(keyinput50), 
        .A(n9973), .ZN(n9982) );
  AOI22_X1 U11017 ( .A1(n4587), .A2(keyinput58), .B1(keyinput26), .B2(n9977), 
        .ZN(n9976) );
  OAI221_X1 U11018 ( .B1(n4587), .B2(keyinput58), .C1(n9977), .C2(keyinput26), 
        .A(n9976), .ZN(n9981) );
  INV_X1 U11019 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n10037) );
  AOI22_X1 U11020 ( .A1(n10037), .A2(keyinput17), .B1(n9979), .B2(keyinput28), 
        .ZN(n9978) );
  OAI221_X1 U11021 ( .B1(n10037), .B2(keyinput17), .C1(n9979), .C2(keyinput28), 
        .A(n9978), .ZN(n9980) );
  NOR4_X1 U11022 ( .A1(n9983), .A2(n9982), .A3(n9981), .A4(n9980), .ZN(n10014)
         );
  AOI22_X1 U11023 ( .A1(n5043), .A2(keyinput35), .B1(keyinput34), .B2(n7541), 
        .ZN(n9984) );
  OAI221_X1 U11024 ( .B1(n5043), .B2(keyinput35), .C1(n7541), .C2(keyinput34), 
        .A(n9984), .ZN(n9995) );
  AOI22_X1 U11025 ( .A1(n9986), .A2(keyinput11), .B1(n5463), .B2(keyinput23), 
        .ZN(n9985) );
  OAI221_X1 U11026 ( .B1(n9986), .B2(keyinput11), .C1(n5463), .C2(keyinput23), 
        .A(n9985), .ZN(n9994) );
  AOI22_X1 U11027 ( .A1(n9989), .A2(keyinput19), .B1(n9988), .B2(keyinput33), 
        .ZN(n9987) );
  OAI221_X1 U11028 ( .B1(n9989), .B2(keyinput19), .C1(n9988), .C2(keyinput33), 
        .A(n9987), .ZN(n9993) );
  XNOR2_X1 U11029 ( .A(P2_REG1_REG_24__SCAN_IN), .B(keyinput2), .ZN(n9991) );
  XNOR2_X1 U11030 ( .A(SI_0_), .B(keyinput38), .ZN(n9990) );
  NAND2_X1 U11031 ( .A1(n9991), .A2(n9990), .ZN(n9992) );
  NOR4_X1 U11032 ( .A1(n9995), .A2(n9994), .A3(n9993), .A4(n9992), .ZN(n10013)
         );
  AOI22_X1 U11033 ( .A1(n9998), .A2(keyinput22), .B1(n9997), .B2(keyinput12), 
        .ZN(n9996) );
  OAI221_X1 U11034 ( .B1(n9998), .B2(keyinput22), .C1(n9997), .C2(keyinput12), 
        .A(n9996), .ZN(n10011) );
  INV_X1 U11035 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n10001) );
  AOI22_X1 U11036 ( .A1(n10001), .A2(keyinput55), .B1(n10000), .B2(keyinput51), 
        .ZN(n9999) );
  OAI221_X1 U11037 ( .B1(n10001), .B2(keyinput55), .C1(n10000), .C2(keyinput51), .A(n9999), .ZN(n10010) );
  INV_X1 U11038 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n10004) );
  AOI22_X1 U11039 ( .A1(n10004), .A2(keyinput16), .B1(n10003), .B2(keyinput53), 
        .ZN(n10002) );
  OAI221_X1 U11040 ( .B1(n10004), .B2(keyinput16), .C1(n10003), .C2(keyinput53), .A(n10002), .ZN(n10009) );
  INV_X1 U11041 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n10007) );
  AOI22_X1 U11042 ( .A1(n10007), .A2(keyinput24), .B1(keyinput10), .B2(n10006), 
        .ZN(n10005) );
  OAI221_X1 U11043 ( .B1(n10007), .B2(keyinput24), .C1(n10006), .C2(keyinput10), .A(n10005), .ZN(n10008) );
  NOR4_X1 U11044 ( .A1(n10011), .A2(n10010), .A3(n10009), .A4(n10008), .ZN(
        n10012) );
  NAND4_X1 U11045 ( .A1(n10015), .A2(n10014), .A3(n10013), .A4(n10012), .ZN(
        n10016) );
  AOI211_X1 U11046 ( .C1(n10019), .C2(n10018), .A(n10017), .B(n10016), .ZN(
        n10023) );
  MUX2_X1 U11047 ( .A(n10021), .B(n10020), .S(P1_U4006), .Z(n10022) );
  XNOR2_X1 U11048 ( .A(n10023), .B(n10022), .ZN(P1_U3582) );
  XOR2_X1 U11049 ( .A(n10024), .B(P2_ADDR_REG_6__SCAN_IN), .Z(ADD_1071_U50) );
  NOR2_X1 U11050 ( .A1(n10026), .A2(n10025), .ZN(n10028) );
  XNOR2_X1 U11051 ( .A(n10028), .B(n10027), .ZN(ADD_1071_U51) );
  OAI21_X1 U11052 ( .B1(n10031), .B2(n10030), .A(n10029), .ZN(n10032) );
  XNOR2_X1 U11053 ( .A(n10032), .B(P1_ADDR_REG_18__SCAN_IN), .ZN(ADD_1071_U55)
         );
  AOI21_X1 U11054 ( .B1(n10035), .B2(n10034), .A(n10033), .ZN(ADD_1071_U47) );
  XOR2_X1 U11055 ( .A(P2_ADDR_REG_8__SCAN_IN), .B(n10036), .Z(ADD_1071_U48) );
  XNOR2_X1 U11056 ( .A(n10038), .B(n10037), .ZN(ADD_1071_U49) );
  XOR2_X1 U11057 ( .A(n10040), .B(n10039), .Z(ADD_1071_U54) );
  XOR2_X1 U11058 ( .A(n10042), .B(n10041), .Z(ADD_1071_U53) );
  XNOR2_X1 U11059 ( .A(n10044), .B(n10043), .ZN(ADD_1071_U52) );
  BUF_X1 U4787 ( .A(n5788), .Z(n4276) );
  CLKBUF_X2 U4821 ( .A(n9821), .Z(n4275) );
  NAND2_X1 U6067 ( .A1(n4712), .A2(n4711), .ZN(n6993) );
  XNOR2_X1 U7540 ( .A(n6112), .B(n6110), .ZN(n8475) );
  AOI21_X1 U7553 ( .B1(n8475), .B2(n8474), .A(n6113), .ZN(n6128) );
  NAND2_X1 U4818 ( .A1(n5682), .A2(n5683), .ZN(n6283) );
  CLKBUF_X1 U5999 ( .A(n7764), .Z(n4282) );
endmodule

