

module b22_C_2inp_gates_syn ( P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN, 
        P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN, 
        P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN, 
        P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN, 
        P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN, 
        P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN, 
        P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN, 
        P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN, 
        P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN, 
        P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN, P3_REG3_REG_0__SCAN_IN, 
        P3_REG3_REG_20__SCAN_IN, P3_REG3_REG_13__SCAN_IN, 
        P3_REG3_REG_22__SCAN_IN, P3_REG3_REG_11__SCAN_IN, 
        P3_REG3_REG_2__SCAN_IN, P3_REG3_REG_18__SCAN_IN, 
        P3_REG3_REG_6__SCAN_IN, P3_REG3_REG_26__SCAN_IN, 
        P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_ADDR_REG_0__SCAN_IN, 
        P3_ADDR_REG_1__SCAN_IN, P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN, 
        P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN, P3_ADDR_REG_6__SCAN_IN, 
        P3_ADDR_REG_7__SCAN_IN, P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, 
        P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, 
        P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, 
        P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, 
        P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, 
        P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, 
        P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, 
        P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, 
        P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, 
        P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, 
        P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, 
        P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, 
        P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, 
        P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, 
        P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, 
        P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, 
        P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, 
        P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, 
        P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, 
        P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, 
        P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, 
        P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, 
        P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, 
        P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, 
        P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, 
        P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, 
        P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN, 
        P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN, 
        P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN, 
        P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN, 
        P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN, 
        P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN, 
        P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN, 
        P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN, 
        P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN, 
        P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN, 
        P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN, 
        P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN, 
        P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN, 
        P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN, 
        P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN, 
        P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN, 
        P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN, 
        P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_4__SCAN_IN, 
        P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_17__SCAN_IN, 
        P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_16__SCAN_IN, 
        P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_12__SCAN_IN, 
        P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_1__SCAN_IN, 
        P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_28__SCAN_IN, 
        P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_3__SCAN_IN, 
        P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_23__SCAN_IN, 
        P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_27__SCAN_IN, 
        P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN, P2_RD_REG_SCAN_IN, 
        P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN, P3_IR_REG_1__SCAN_IN, 
        P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN, P3_IR_REG_4__SCAN_IN, 
        P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN, P3_IR_REG_7__SCAN_IN, 
        P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN, P3_IR_REG_10__SCAN_IN, 
        P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN, P3_IR_REG_13__SCAN_IN, 
        P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN, P3_IR_REG_16__SCAN_IN, 
        P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN, P3_IR_REG_19__SCAN_IN, 
        P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN, P3_IR_REG_22__SCAN_IN, 
        P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN, P3_IR_REG_25__SCAN_IN, 
        P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN, P3_IR_REG_28__SCAN_IN, 
        P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN, P3_IR_REG_31__SCAN_IN, 
        P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN, P3_D_REG_2__SCAN_IN, 
        P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN, P3_D_REG_5__SCAN_IN, 
        P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN, P3_D_REG_8__SCAN_IN, 
        P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN, P3_D_REG_11__SCAN_IN, 
        P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN, P3_D_REG_14__SCAN_IN, 
        P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN, P3_D_REG_17__SCAN_IN, 
        P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN, P3_D_REG_20__SCAN_IN, 
        P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN, P3_D_REG_23__SCAN_IN, 
        P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN, P3_D_REG_26__SCAN_IN, 
        P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN, P3_D_REG_29__SCAN_IN, 
        P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN, P3_REG0_REG_0__SCAN_IN, 
        P3_REG0_REG_1__SCAN_IN, P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN, 
        P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN, P3_REG0_REG_6__SCAN_IN, 
        P3_REG0_REG_7__SCAN_IN, P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN, 
        P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN, 
        P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN, 
        P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN, 
        P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN, 
        P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN, 
        P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN, 
        P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN, 
        P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN, 
        P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN, 
        P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN, 
        P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN, 
        P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN, P3_REG1_REG_2__SCAN_IN, 
        P3_REG1_REG_3__SCAN_IN, P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN, 
        P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN, P3_REG1_REG_8__SCAN_IN, 
        P3_REG1_REG_9__SCAN_IN, P3_REG1_REG_10__SCAN_IN, 
        P3_REG1_REG_11__SCAN_IN, P3_REG1_REG_12__SCAN_IN, 
        P3_REG1_REG_13__SCAN_IN, P3_REG1_REG_14__SCAN_IN, 
        P3_REG1_REG_15__SCAN_IN, P3_REG1_REG_16__SCAN_IN, 
        P3_REG1_REG_17__SCAN_IN, P3_REG1_REG_18__SCAN_IN, 
        P3_REG1_REG_19__SCAN_IN, P3_REG1_REG_20__SCAN_IN, 
        P3_REG1_REG_21__SCAN_IN, P3_REG1_REG_22__SCAN_IN, 
        P3_REG1_REG_23__SCAN_IN, P3_REG1_REG_24__SCAN_IN, 
        P3_REG1_REG_25__SCAN_IN, P3_REG1_REG_26__SCAN_IN, 
        P3_REG1_REG_27__SCAN_IN, P3_REG1_REG_28__SCAN_IN, 
        P3_REG1_REG_29__SCAN_IN, P3_REG1_REG_30__SCAN_IN, 
        P3_REG1_REG_31__SCAN_IN, P3_REG2_REG_0__SCAN_IN, 
        P3_REG2_REG_1__SCAN_IN, P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN, 
        P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN, P3_REG2_REG_6__SCAN_IN, 
        P3_REG2_REG_7__SCAN_IN, P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN, 
        P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN, 
        P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN, 
        P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN, 
        P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN, 
        P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN, 
        P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN, 
        P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN, 
        P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN, 
        P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN, 
        P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN, 
        P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN, 
        P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN, 
        P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN, 
        P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN, 
        P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN, 
        P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, SUB_1596_U4, 
        SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65, SUB_1596_U66, 
        SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70, SUB_1596_U54, 
        SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58, SUB_1596_U59, 
        SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53, U29, U28, 
        P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349, 
        P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342, 
        P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335, 
        P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328, 
        P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446, P1_U3323, 
        P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316, 
        P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309, 
        P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302, 
        P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295, 
        P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471, P1_U3474, 
        P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492, P1_U3495, 
        P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513, P1_U3515, 
        P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, 
        P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, 
        P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, 
        P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, 
        P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, 
        P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556, P1_U3557, 
        P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290, P1_U3289, 
        P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282, 
        P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275, 
        P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268, 
        P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, P1_U3262, 
        P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255, 
        P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248, 
        P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560, P1_U3561, 
        P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, 
        P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, 
        P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, 
        P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588, P1_U3589, 
        P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239, P1_U3238, 
        P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231, 
        P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224, 
        P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, 
        P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, P1_U4016, 
        P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321, 
        P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314, 
        P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307, 
        P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300, 
        P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417, P2_U3295, 
        P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, 
        P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, 
        P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, 
        P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, 
        P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442, P2_U3445, 
        P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463, P2_U3466, 
        P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484, P2_U3486, 
        P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492, P2_U3493, 
        P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499, P2_U3500, 
        P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506, P2_U3507, 
        P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, P2_U3514, 
        P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, P2_U3521, 
        P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527, P2_U3528, 
        P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, 
        P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, 
        P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, 
        P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241, P2_U3240, 
        P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, 
        P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, 
        P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, 
        P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531, P2_U3532, 
        P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, 
        P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, 
        P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552, P2_U3553, 
        P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559, P2_U3560, 
        P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211, P2_U3210, 
        P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, 
        P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, 
        P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, 
        P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087, P2_U3947, 
        P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290, P3_U3289, 
        P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283, P3_U3282, 
        P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276, P3_U3275, 
        P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269, P3_U3268, 
        P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377, P3_U3263, 
        P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257, P3_U3256, 
        P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250, P3_U3249, 
        P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243, P3_U3242, 
        P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236, P3_U3235, 
        P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402, P3_U3405, 
        P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423, P3_U3426, 
        P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444, P3_U3446, 
        P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452, P3_U3453, 
        P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459, P3_U3460, 
        P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466, P3_U3467, 
        P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473, P3_U3474, 
        P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480, P3_U3481, 
        P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487, P3_U3488, 
        P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230, P3_U3229, 
        P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223, P3_U3222, 
        P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216, P3_U3215, 
        P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209, P3_U3208, 
        P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202, P3_U3201, 
        P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195, P3_U3194, 
        P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188, P3_U3187, 
        P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491, P3_U3492, 
        P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498, P3_U3499, 
        P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505, P3_U3506, 
        P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512, P3_U3513, 
        P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519, P3_U3520, 
        P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179, P3_U3178, 
        P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172, P3_U3171, 
        P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165, P3_U3164, 
        P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158, P3_U3157, 
        P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150, P3_U3897, 
        keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, 
        keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, 
        keyinput12, keyinput13, keyinput14, keyinput15, keyinput16, keyinput17, 
        keyinput18, keyinput19, keyinput20, keyinput21, keyinput22, keyinput23, 
        keyinput24, keyinput25, keyinput26, keyinput27, keyinput28, keyinput29, 
        keyinput30, keyinput31, keyinput32, keyinput33, keyinput34, keyinput35, 
        keyinput36, keyinput37, keyinput38, keyinput39, keyinput40, keyinput41, 
        keyinput42, keyinput43, keyinput44, keyinput45, keyinput46, keyinput47, 
        keyinput48, keyinput49, keyinput50, keyinput51, keyinput52, keyinput53, 
        keyinput54, keyinput55, keyinput56, keyinput57, keyinput58, keyinput59, 
        keyinput60, keyinput61, keyinput62, keyinput63, keyinput64, keyinput65, 
        keyinput66, keyinput67, keyinput68, keyinput69, keyinput70, keyinput71, 
        keyinput72, keyinput73, keyinput74, keyinput75, keyinput76, keyinput77, 
        keyinput78, keyinput79, keyinput80, keyinput81, keyinput82, keyinput83, 
        keyinput84, keyinput85, keyinput86, keyinput87, keyinput88, keyinput89, 
        keyinput90, keyinput91, keyinput92, keyinput93, keyinput94, keyinput95, 
        keyinput96, keyinput97, keyinput98, keyinput99, keyinput100, 
        keyinput101, keyinput102, keyinput103, keyinput104, keyinput105, 
        keyinput106, keyinput107, keyinput108, keyinput109, keyinput110, 
        keyinput111, keyinput112, keyinput113, keyinput114, keyinput115, 
        keyinput116, keyinput117, keyinput118, keyinput119, keyinput120, 
        keyinput121, keyinput122, keyinput123, keyinput124, keyinput125, 
        keyinput126, keyinput127 );
  input P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN,
         P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN,
         P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN,
         P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN,
         P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN,
         P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN,
         P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN,
         P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN,
         P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN,
         P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN,
         P3_REG3_REG_0__SCAN_IN, P3_REG3_REG_20__SCAN_IN,
         P3_REG3_REG_13__SCAN_IN, P3_REG3_REG_22__SCAN_IN,
         P3_REG3_REG_11__SCAN_IN, P3_REG3_REG_2__SCAN_IN,
         P3_REG3_REG_18__SCAN_IN, P3_REG3_REG_6__SCAN_IN,
         P3_REG3_REG_26__SCAN_IN, P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN,
         P3_DATAO_REG_31__SCAN_IN, P3_DATAO_REG_30__SCAN_IN,
         P3_DATAO_REG_29__SCAN_IN, P3_DATAO_REG_28__SCAN_IN,
         P3_DATAO_REG_27__SCAN_IN, P3_DATAO_REG_26__SCAN_IN,
         P3_DATAO_REG_25__SCAN_IN, P3_DATAO_REG_24__SCAN_IN,
         P3_DATAO_REG_23__SCAN_IN, P3_DATAO_REG_22__SCAN_IN,
         P3_DATAO_REG_21__SCAN_IN, P3_DATAO_REG_20__SCAN_IN,
         P3_DATAO_REG_19__SCAN_IN, P3_DATAO_REG_18__SCAN_IN,
         P3_DATAO_REG_17__SCAN_IN, P3_DATAO_REG_16__SCAN_IN,
         P3_DATAO_REG_15__SCAN_IN, P3_DATAO_REG_14__SCAN_IN,
         P3_DATAO_REG_13__SCAN_IN, P3_DATAO_REG_12__SCAN_IN,
         P3_DATAO_REG_11__SCAN_IN, P3_DATAO_REG_10__SCAN_IN,
         P3_DATAO_REG_9__SCAN_IN, P3_DATAO_REG_8__SCAN_IN,
         P3_DATAO_REG_7__SCAN_IN, P3_DATAO_REG_6__SCAN_IN,
         P3_DATAO_REG_5__SCAN_IN, P3_DATAO_REG_4__SCAN_IN,
         P3_DATAO_REG_3__SCAN_IN, P3_DATAO_REG_2__SCAN_IN,
         P3_DATAO_REG_1__SCAN_IN, P3_DATAO_REG_0__SCAN_IN,
         P3_ADDR_REG_0__SCAN_IN, P3_ADDR_REG_1__SCAN_IN,
         P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN,
         P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN,
         P3_ADDR_REG_6__SCAN_IN, P3_ADDR_REG_7__SCAN_IN,
         P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, P1_IR_REG_0__SCAN_IN,
         P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN,
         P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN,
         P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN,
         P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN,
         P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN,
         P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN,
         P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN,
         P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN,
         P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN,
         P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN,
         P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN,
         P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN,
         P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN,
         P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN,
         P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN,
         P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN,
         P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN,
         P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN,
         P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN,
         P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN,
         P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN,
         P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN,
         P2_RD_REG_SCAN_IN, P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN,
         P3_IR_REG_1__SCAN_IN, P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN,
         P3_IR_REG_4__SCAN_IN, P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN,
         P3_IR_REG_7__SCAN_IN, P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN,
         P3_IR_REG_10__SCAN_IN, P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN,
         P3_IR_REG_13__SCAN_IN, P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN,
         P3_IR_REG_16__SCAN_IN, P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN,
         P3_IR_REG_19__SCAN_IN, P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN,
         P3_IR_REG_22__SCAN_IN, P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN,
         P3_IR_REG_25__SCAN_IN, P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN,
         P3_IR_REG_28__SCAN_IN, P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN,
         P3_IR_REG_31__SCAN_IN, P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN,
         P3_D_REG_2__SCAN_IN, P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN,
         P3_D_REG_5__SCAN_IN, P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN,
         P3_D_REG_8__SCAN_IN, P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN,
         P3_D_REG_11__SCAN_IN, P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN,
         P3_D_REG_14__SCAN_IN, P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN,
         P3_D_REG_17__SCAN_IN, P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN,
         P3_D_REG_20__SCAN_IN, P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN,
         P3_D_REG_23__SCAN_IN, P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN,
         P3_D_REG_26__SCAN_IN, P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN,
         P3_D_REG_29__SCAN_IN, P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN,
         P3_REG0_REG_0__SCAN_IN, P3_REG0_REG_1__SCAN_IN,
         P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN,
         P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN,
         P3_REG0_REG_6__SCAN_IN, P3_REG0_REG_7__SCAN_IN,
         P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN,
         P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN,
         P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN,
         P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN,
         P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN,
         P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN,
         P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN,
         P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN,
         P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN,
         P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN,
         P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN,
         P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN,
         P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN,
         P3_REG1_REG_2__SCAN_IN, P3_REG1_REG_3__SCAN_IN,
         P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN,
         P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN,
         P3_REG1_REG_8__SCAN_IN, P3_REG1_REG_9__SCAN_IN,
         P3_REG1_REG_10__SCAN_IN, P3_REG1_REG_11__SCAN_IN,
         P3_REG1_REG_12__SCAN_IN, P3_REG1_REG_13__SCAN_IN,
         P3_REG1_REG_14__SCAN_IN, P3_REG1_REG_15__SCAN_IN,
         P3_REG1_REG_16__SCAN_IN, P3_REG1_REG_17__SCAN_IN,
         P3_REG1_REG_18__SCAN_IN, P3_REG1_REG_19__SCAN_IN,
         P3_REG1_REG_20__SCAN_IN, P3_REG1_REG_21__SCAN_IN,
         P3_REG1_REG_22__SCAN_IN, P3_REG1_REG_23__SCAN_IN,
         P3_REG1_REG_24__SCAN_IN, P3_REG1_REG_25__SCAN_IN,
         P3_REG1_REG_26__SCAN_IN, P3_REG1_REG_27__SCAN_IN,
         P3_REG1_REG_28__SCAN_IN, P3_REG1_REG_29__SCAN_IN,
         P3_REG1_REG_30__SCAN_IN, P3_REG1_REG_31__SCAN_IN,
         P3_REG2_REG_0__SCAN_IN, P3_REG2_REG_1__SCAN_IN,
         P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN,
         P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN,
         P3_REG2_REG_6__SCAN_IN, P3_REG2_REG_7__SCAN_IN,
         P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN,
         P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN,
         P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN,
         P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN,
         P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN,
         P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN,
         P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN,
         P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN,
         P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN,
         P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN,
         P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN,
         P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN,
         P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN,
         P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN,
         P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN,
         P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN,
         P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, keyinput0,
         keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, keyinput6,
         keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, keyinput12,
         keyinput13, keyinput14, keyinput15, keyinput16, keyinput17,
         keyinput18, keyinput19, keyinput20, keyinput21, keyinput22,
         keyinput23, keyinput24, keyinput25, keyinput26, keyinput27,
         keyinput28, keyinput29, keyinput30, keyinput31, keyinput32,
         keyinput33, keyinput34, keyinput35, keyinput36, keyinput37,
         keyinput38, keyinput39, keyinput40, keyinput41, keyinput42,
         keyinput43, keyinput44, keyinput45, keyinput46, keyinput47,
         keyinput48, keyinput49, keyinput50, keyinput51, keyinput52,
         keyinput53, keyinput54, keyinput55, keyinput56, keyinput57,
         keyinput58, keyinput59, keyinput60, keyinput61, keyinput62,
         keyinput63, keyinput64, keyinput65, keyinput66, keyinput67,
         keyinput68, keyinput69, keyinput70, keyinput71, keyinput72,
         keyinput73, keyinput74, keyinput75, keyinput76, keyinput77,
         keyinput78, keyinput79, keyinput80, keyinput81, keyinput82,
         keyinput83, keyinput84, keyinput85, keyinput86, keyinput87,
         keyinput88, keyinput89, keyinput90, keyinput91, keyinput92,
         keyinput93, keyinput94, keyinput95, keyinput96, keyinput97,
         keyinput98, keyinput99, keyinput100, keyinput101, keyinput102,
         keyinput103, keyinput104, keyinput105, keyinput106, keyinput107,
         keyinput108, keyinput109, keyinput110, keyinput111, keyinput112,
         keyinput113, keyinput114, keyinput115, keyinput116, keyinput117,
         keyinput118, keyinput119, keyinput120, keyinput121, keyinput122,
         keyinput123, keyinput124, keyinput125, keyinput126, keyinput127;
  output SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65,
         SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70,
         SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58,
         SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53,
         U29, U28, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350,
         P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343,
         P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336,
         P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329,
         P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446,
         P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317,
         P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310,
         P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303,
         P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296,
         P1_U3295, P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471,
         P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492,
         P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556,
         P1_U3557, P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290,
         P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283,
         P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276,
         P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269,
         P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263,
         P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256,
         P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249,
         P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588,
         P1_U3589, P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239,
         P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232,
         P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085,
         P1_U4016, P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322,
         P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315,
         P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308,
         P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301,
         P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417,
         P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289,
         P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282,
         P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275,
         P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268,
         P2_U3267, P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442,
         P2_U3445, P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463,
         P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484,
         P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492,
         P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499,
         P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506,
         P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513,
         P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520,
         P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527,
         P2_U3528, P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262,
         P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255,
         P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248,
         P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241,
         P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234,
         P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227,
         P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220,
         P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531,
         P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538,
         P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545,
         P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552,
         P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559,
         P2_U3560, P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204,
         P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197,
         P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190,
         P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087,
         P2_U3947, P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290,
         P3_U3289, P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283,
         P3_U3282, P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276,
         P3_U3275, P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269,
         P3_U3268, P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377,
         P3_U3263, P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257,
         P3_U3256, P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250,
         P3_U3249, P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243,
         P3_U3242, P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236,
         P3_U3235, P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402,
         P3_U3405, P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423,
         P3_U3426, P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444,
         P3_U3446, P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452,
         P3_U3453, P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459,
         P3_U3460, P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466,
         P3_U3467, P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473,
         P3_U3474, P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480,
         P3_U3481, P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487,
         P3_U3488, P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230,
         P3_U3229, P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223,
         P3_U3222, P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216,
         P3_U3215, P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209,
         P3_U3208, P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202,
         P3_U3201, P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195,
         P3_U3194, P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188,
         P3_U3187, P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491,
         P3_U3492, P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498,
         P3_U3499, P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505,
         P3_U3506, P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512,
         P3_U3513, P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519,
         P3_U3520, P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179,
         P3_U3178, P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172,
         P3_U3171, P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165,
         P3_U3164, P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158,
         P3_U3157, P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150,
         P3_U3897;
  wire   n6522, n6523, n6525, n6527, n6528, n6529, n6530, n6531, n6532, n6533,
         n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543,
         n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553,
         n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563,
         n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573,
         n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583,
         n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593,
         n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603,
         n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613,
         n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623,
         n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633,
         n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643,
         n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653,
         n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663,
         n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673,
         n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683,
         n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693,
         n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703,
         n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713,
         n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723,
         n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733,
         n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743,
         n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753,
         n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763,
         n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773,
         n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783,
         n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793,
         n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803,
         n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813,
         n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823,
         n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833,
         n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843,
         n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853,
         n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863,
         n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873,
         n6874, n6875, n6876, n6877, n6878, n6879, n6881, n6882, n6883, n6884,
         n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894,
         n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904,
         n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914,
         n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924,
         n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934,
         n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944,
         n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954,
         n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964,
         n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974,
         n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984,
         n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994,
         n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004,
         n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014,
         n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024,
         n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034,
         n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044,
         n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054,
         n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064,
         n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074,
         n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084,
         n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094,
         n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104,
         n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114,
         n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124,
         n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134,
         n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144,
         n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154,
         n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164,
         n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174,
         n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184,
         n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194,
         n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204,
         n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214,
         n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224,
         n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234,
         n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244,
         n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254,
         n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264,
         n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274,
         n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284,
         n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294,
         n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304,
         n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314,
         n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324,
         n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334,
         n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344,
         n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354,
         n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364,
         n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374,
         n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384,
         n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394,
         n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404,
         n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414,
         n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424,
         n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434,
         n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444,
         n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454,
         n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464,
         n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474,
         n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484,
         n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494,
         n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504,
         n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514,
         n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524,
         n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534,
         n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544,
         n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554,
         n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564,
         n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574,
         n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584,
         n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594,
         n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604,
         n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614,
         n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624,
         n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634,
         n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644,
         n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654,
         n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664,
         n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674,
         n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684,
         n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694,
         n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704,
         n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714,
         n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724,
         n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734,
         n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744,
         n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754,
         n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764,
         n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774,
         n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784,
         n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794,
         n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804,
         n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814,
         n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824,
         n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834,
         n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844,
         n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854,
         n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864,
         n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874,
         n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884,
         n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894,
         n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904,
         n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914,
         n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924,
         n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934,
         n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944,
         n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954,
         n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964,
         n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974,
         n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984,
         n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994,
         n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004,
         n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014,
         n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024,
         n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034,
         n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044,
         n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054,
         n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064,
         n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074,
         n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084,
         n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094,
         n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104,
         n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114,
         n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124,
         n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134,
         n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144,
         n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154,
         n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164,
         n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174,
         n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184,
         n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194,
         n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204,
         n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214,
         n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224,
         n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234,
         n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244,
         n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254,
         n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264,
         n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274,
         n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284,
         n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294,
         n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304,
         n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314,
         n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324,
         n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334,
         n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344,
         n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354,
         n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364,
         n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374,
         n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384,
         n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394,
         n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404,
         n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414,
         n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424,
         n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434,
         n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444,
         n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454,
         n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464,
         n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474,
         n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484,
         n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494,
         n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504,
         n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514,
         n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524,
         n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534,
         n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544,
         n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554,
         n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564,
         n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574,
         n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584,
         n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594,
         n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604,
         n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614,
         n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624,
         n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634,
         n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644,
         n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654,
         n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664,
         n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674,
         n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684,
         n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694,
         n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704,
         n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714,
         n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724,
         n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734,
         n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744,
         n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754,
         n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764,
         n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774,
         n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784,
         n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794,
         n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804,
         n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814,
         n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824,
         n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834,
         n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844,
         n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854,
         n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864,
         n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874,
         n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884,
         n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894,
         n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904,
         n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914,
         n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924,
         n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934,
         n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944,
         n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954,
         n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964,
         n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974,
         n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984,
         n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994,
         n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004,
         n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014,
         n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024,
         n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034,
         n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044,
         n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054,
         n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064,
         n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074,
         n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084,
         n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094,
         n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104,
         n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114,
         n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124,
         n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134,
         n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144,
         n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154,
         n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164,
         n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174,
         n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184,
         n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194,
         n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204,
         n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214,
         n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224,
         n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234,
         n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244,
         n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254,
         n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264,
         n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274,
         n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284,
         n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294,
         n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304,
         n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314,
         n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324,
         n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334,
         n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344,
         n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354,
         n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364,
         n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374,
         n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384,
         n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394,
         n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404,
         n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414,
         n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424,
         n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434,
         n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444,
         n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454,
         n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464,
         n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474,
         n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484,
         n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494,
         n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504,
         n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514,
         n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524,
         n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534,
         n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544,
         n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554,
         n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564,
         n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574,
         n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584,
         n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594,
         n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604,
         n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614,
         n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624,
         n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634,
         n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644,
         n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654,
         n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664,
         n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674,
         n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684,
         n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694,
         n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704,
         n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714,
         n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724,
         n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734,
         n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744,
         n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754,
         n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764,
         n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774,
         n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784,
         n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794,
         n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804,
         n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814,
         n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824,
         n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834,
         n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844,
         n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854,
         n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864,
         n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874,
         n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884,
         n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894,
         n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904,
         n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914,
         n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924,
         n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934,
         n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944,
         n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954,
         n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964,
         n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974,
         n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984,
         n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994,
         n9995, n9996, n9997, n9998, n9999, n10000, n10001, n10002, n10003,
         n10004, n10005, n10006, n10007, n10008, n10009, n10010, n10011,
         n10012, n10013, n10014, n10015, n10016, n10017, n10018, n10019,
         n10020, n10021, n10022, n10023, n10024, n10025, n10026, n10027,
         n10028, n10029, n10030, n10031, n10032, n10033, n10034, n10035,
         n10036, n10037, n10038, n10039, n10040, n10041, n10042, n10043,
         n10044, n10045, n10046, n10047, n10048, n10049, n10050, n10051,
         n10052, n10053, n10054, n10055, n10056, n10057, n10058, n10059,
         n10060, n10061, n10062, n10063, n10064, n10065, n10066, n10067,
         n10068, n10069, n10070, n10071, n10072, n10073, n10074, n10075,
         n10076, n10077, n10078, n10079, n10080, n10081, n10082, n10083,
         n10084, n10085, n10086, n10087, n10088, n10089, n10090, n10091,
         n10092, n10093, n10094, n10095, n10096, n10097, n10098, n10099,
         n10100, n10101, n10102, n10103, n10104, n10105, n10106, n10107,
         n10108, n10109, n10110, n10111, n10112, n10113, n10114, n10115,
         n10116, n10117, n10118, n10119, n10120, n10121, n10122, n10123,
         n10124, n10125, n10126, n10127, n10128, n10129, n10130, n10131,
         n10132, n10133, n10134, n10135, n10136, n10137, n10138, n10139,
         n10140, n10141, n10142, n10143, n10144, n10145, n10146, n10147,
         n10148, n10149, n10150, n10151, n10152, n10153, n10154, n10155,
         n10156, n10157, n10158, n10159, n10160, n10161, n10162, n10163,
         n10164, n10165, n10166, n10167, n10168, n10169, n10170, n10171,
         n10172, n10173, n10174, n10175, n10176, n10177, n10178, n10179,
         n10180, n10181, n10182, n10183, n10184, n10185, n10186, n10187,
         n10188, n10189, n10190, n10191, n10192, n10193, n10194, n10195,
         n10196, n10197, n10198, n10199, n10200, n10201, n10202, n10203,
         n10204, n10205, n10206, n10207, n10208, n10209, n10210, n10211,
         n10212, n10213, n10214, n10215, n10216, n10217, n10218, n10219,
         n10220, n10221, n10222, n10223, n10224, n10225, n10226, n10227,
         n10228, n10229, n10230, n10231, n10232, n10233, n10234, n10235,
         n10236, n10237, n10238, n10239, n10240, n10241, n10242, n10243,
         n10244, n10245, n10246, n10247, n10248, n10249, n10250, n10251,
         n10252, n10253, n10254, n10255, n10256, n10257, n10258, n10259,
         n10260, n10261, n10262, n10263, n10264, n10265, n10266, n10267,
         n10268, n10269, n10270, n10271, n10272, n10273, n10274, n10275,
         n10276, n10277, n10278, n10279, n10280, n10281, n10282, n10283,
         n10284, n10285, n10286, n10287, n10288, n10289, n10290, n10291,
         n10292, n10293, n10294, n10295, n10296, n10297, n10298, n10299,
         n10300, n10301, n10302, n10303, n10304, n10305, n10306, n10307,
         n10308, n10309, n10310, n10311, n10312, n10313, n10314, n10315,
         n10316, n10317, n10318, n10319, n10320, n10321, n10322, n10323,
         n10324, n10325, n10326, n10327, n10328, n10329, n10330, n10331,
         n10332, n10333, n10334, n10335, n10336, n10337, n10338, n10339,
         n10340, n10341, n10342, n10343, n10344, n10345, n10346, n10347,
         n10348, n10349, n10350, n10351, n10352, n10353, n10354, n10355,
         n10356, n10357, n10358, n10359, n10360, n10361, n10362, n10363,
         n10364, n10365, n10366, n10367, n10368, n10369, n10370, n10371,
         n10372, n10373, n10374, n10375, n10376, n10377, n10378, n10379,
         n10380, n10381, n10382, n10383, n10384, n10385, n10386, n10387,
         n10388, n10389, n10390, n10391, n10392, n10393, n10394, n10395,
         n10396, n10397, n10398, n10399, n10400, n10401, n10402, n10403,
         n10404, n10405, n10406, n10407, n10408, n10409, n10410, n10411,
         n10412, n10413, n10414, n10415, n10416, n10417, n10418, n10419,
         n10420, n10421, n10422, n10423, n10424, n10425, n10426, n10427,
         n10428, n10429, n10430, n10431, n10432, n10433, n10434, n10435,
         n10436, n10437, n10438, n10439, n10440, n10441, n10442, n10443,
         n10444, n10445, n10446, n10447, n10448, n10449, n10450, n10451,
         n10452, n10453, n10454, n10455, n10456, n10457, n10458, n10459,
         n10460, n10461, n10462, n10463, n10464, n10465, n10466, n10467,
         n10468, n10469, n10470, n10471, n10472, n10473, n10474, n10475,
         n10476, n10477, n10478, n10479, n10480, n10481, n10482, n10483,
         n10484, n10485, n10486, n10487, n10488, n10489, n10490, n10491,
         n10492, n10493, n10494, n10495, n10496, n10497, n10498, n10499,
         n10500, n10501, n10502, n10503, n10504, n10505, n10506, n10507,
         n10508, n10509, n10510, n10511, n10512, n10513, n10514, n10515,
         n10516, n10517, n10518, n10519, n10520, n10521, n10522, n10523,
         n10524, n10525, n10526, n10527, n10528, n10529, n10530, n10531,
         n10532, n10533, n10534, n10535, n10536, n10537, n10538, n10539,
         n10540, n10541, n10542, n10543, n10544, n10545, n10546, n10547,
         n10548, n10549, n10550, n10551, n10552, n10553, n10554, n10555,
         n10556, n10557, n10558, n10559, n10560, n10561, n10562, n10563,
         n10564, n10565, n10566, n10567, n10568, n10569, n10570, n10571,
         n10572, n10573, n10574, n10575, n10576, n10577, n10578, n10579,
         n10580, n10581, n10582, n10583, n10584, n10585, n10586, n10587,
         n10588, n10589, n10590, n10591, n10592, n10593, n10594, n10595,
         n10596, n10597, n10598, n10599, n10600, n10601, n10602, n10603,
         n10604, n10605, n10606, n10607, n10608, n10609, n10610, n10611,
         n10612, n10613, n10614, n10615, n10616, n10617, n10618, n10619,
         n10620, n10621, n10622, n10623, n10624, n10625, n10626, n10627,
         n10628, n10629, n10630, n10631, n10632, n10633, n10634, n10635,
         n10636, n10637, n10638, n10639, n10640, n10641, n10642, n10643,
         n10644, n10645, n10646, n10647, n10648, n10649, n10650, n10651,
         n10652, n10653, n10654, n10655, n10656, n10657, n10658, n10659,
         n10660, n10661, n10662, n10663, n10664, n10665, n10666, n10667,
         n10668, n10669, n10670, n10671, n10672, n10673, n10674, n10675,
         n10676, n10677, n10678, n10679, n10680, n10681, n10682, n10683,
         n10684, n10685, n10686, n10687, n10688, n10689, n10690, n10691,
         n10692, n10693, n10694, n10695, n10696, n10697, n10698, n10699,
         n10700, n10701, n10702, n10703, n10704, n10705, n10706, n10707,
         n10708, n10709, n10710, n10711, n10712, n10713, n10714, n10715,
         n10716, n10717, n10718, n10719, n10720, n10721, n10722, n10723,
         n10724, n10725, n10726, n10727, n10728, n10729, n10730, n10731,
         n10732, n10733, n10734, n10735, n10736, n10737, n10738, n10739,
         n10740, n10741, n10742, n10743, n10744, n10745, n10746, n10747,
         n10748, n10749, n10750, n10751, n10752, n10753, n10754, n10755,
         n10756, n10757, n10758, n10759, n10760, n10761, n10762, n10763,
         n10764, n10765, n10766, n10767, n10768, n10769, n10770, n10771,
         n10772, n10773, n10774, n10775, n10776, n10777, n10778, n10779,
         n10780, n10781, n10782, n10783, n10784, n10785, n10786, n10787,
         n10788, n10789, n10790, n10791, n10792, n10793, n10794, n10795,
         n10796, n10797, n10798, n10799, n10800, n10801, n10802, n10803,
         n10804, n10805, n10806, n10807, n10808, n10809, n10810, n10811,
         n10812, n10813, n10814, n10815, n10816, n10817, n10818, n10819,
         n10820, n10821, n10822, n10823, n10824, n10825, n10826, n10827,
         n10828, n10829, n10830, n10831, n10832, n10833, n10834, n10835,
         n10836, n10837, n10838, n10839, n10840, n10841, n10842, n10843,
         n10844, n10845, n10846, n10847, n10848, n10849, n10850, n10851,
         n10852, n10853, n10854, n10855, n10856, n10857, n10858, n10859,
         n10860, n10861, n10862, n10863, n10864, n10865, n10866, n10867,
         n10868, n10869, n10870, n10871, n10872, n10873, n10874, n10875,
         n10876, n10877, n10878, n10879, n10880, n10881, n10882, n10883,
         n10884, n10885, n10886, n10887, n10888, n10889, n10890, n10891,
         n10892, n10893, n10894, n10895, n10896, n10897, n10898, n10899,
         n10900, n10901, n10902, n10903, n10904, n10905, n10906, n10907,
         n10908, n10909, n10910, n10911, n10912, n10913, n10914, n10915,
         n10916, n10917, n10918, n10919, n10920, n10921, n10922, n10923,
         n10924, n10925, n10926, n10927, n10928, n10929, n10930, n10931,
         n10932, n10933, n10934, n10935, n10936, n10937, n10938, n10939,
         n10940, n10941, n10942, n10943, n10944, n10945, n10946, n10947,
         n10948, n10949, n10950, n10951, n10952, n10953, n10954, n10955,
         n10956, n10957, n10958, n10959, n10960, n10961, n10962, n10963,
         n10964, n10965, n10966, n10967, n10968, n10969, n10970, n10971,
         n10972, n10973, n10974, n10975, n10976, n10977, n10978, n10979,
         n10980, n10981, n10982, n10983, n10984, n10985, n10986, n10987,
         n10988, n10989, n10990, n10991, n10992, n10993, n10994, n10995,
         n10996, n10997, n10998, n10999, n11000, n11001, n11002, n11003,
         n11004, n11005, n11006, n11007, n11008, n11009, n11010, n11011,
         n11012, n11013, n11014, n11015, n11016, n11017, n11018, n11019,
         n11020, n11021, n11022, n11023, n11024, n11025, n11026, n11027,
         n11028, n11029, n11030, n11031, n11032, n11033, n11034, n11035,
         n11036, n11037, n11038, n11039, n11040, n11041, n11042, n11043,
         n11044, n11045, n11046, n11047, n11048, n11049, n11050, n11051,
         n11052, n11053, n11054, n11055, n11056, n11057, n11058, n11059,
         n11060, n11061, n11062, n11063, n11064, n11065, n11066, n11067,
         n11068, n11069, n11070, n11071, n11072, n11073, n11074, n11075,
         n11076, n11077, n11078, n11079, n11080, n11081, n11082, n11083,
         n11084, n11085, n11086, n11087, n11088, n11089, n11090, n11091,
         n11092, n11093, n11094, n11095, n11096, n11097, n11098, n11099,
         n11100, n11101, n11102, n11103, n11104, n11105, n11106, n11107,
         n11108, n11109, n11110, n11111, n11112, n11113, n11114, n11115,
         n11116, n11117, n11118, n11119, n11120, n11121, n11122, n11123,
         n11124, n11125, n11126, n11127, n11128, n11129, n11130, n11131,
         n11132, n11133, n11134, n11135, n11136, n11137, n11138, n11139,
         n11140, n11141, n11142, n11143, n11144, n11145, n11146, n11147,
         n11148, n11149, n11150, n11151, n11152, n11153, n11154, n11155,
         n11156, n11157, n11158, n11159, n11160, n11161, n11162, n11163,
         n11164, n11165, n11166, n11167, n11168, n11169, n11170, n11171,
         n11172, n11173, n11174, n11175, n11176, n11177, n11178, n11179,
         n11180, n11181, n11182, n11183, n11184, n11185, n11186, n11187,
         n11188, n11189, n11190, n11191, n11192, n11193, n11194, n11195,
         n11196, n11197, n11198, n11199, n11200, n11201, n11202, n11203,
         n11204, n11205, n11206, n11207, n11208, n11209, n11210, n11211,
         n11212, n11213, n11214, n11215, n11216, n11217, n11218, n11219,
         n11220, n11221, n11222, n11223, n11224, n11225, n11226, n11227,
         n11228, n11229, n11230, n11231, n11232, n11233, n11234, n11235,
         n11236, n11237, n11238, n11239, n11240, n11241, n11242, n11243,
         n11244, n11245, n11246, n11247, n11248, n11249, n11250, n11251,
         n11252, n11253, n11254, n11255, n11256, n11257, n11258, n11259,
         n11260, n11261, n11262, n11263, n11264, n11265, n11266, n11267,
         n11268, n11269, n11270, n11271, n11272, n11273, n11274, n11275,
         n11276, n11277, n11278, n11279, n11280, n11281, n11282, n11283,
         n11284, n11285, n11286, n11287, n11288, n11289, n11290, n11291,
         n11292, n11293, n11294, n11295, n11296, n11297, n11298, n11299,
         n11300, n11301, n11302, n11303, n11304, n11305, n11306, n11307,
         n11308, n11309, n11310, n11311, n11312, n11313, n11314, n11315,
         n11316, n11317, n11318, n11319, n11320, n11321, n11322, n11323,
         n11324, n11325, n11326, n11327, n11328, n11329, n11330, n11331,
         n11332, n11333, n11334, n11335, n11336, n11337, n11338, n11339,
         n11340, n11341, n11342, n11343, n11344, n11345, n11346, n11347,
         n11348, n11349, n11350, n11351, n11352, n11353, n11354, n11355,
         n11356, n11357, n11358, n11359, n11360, n11361, n11362, n11363,
         n11364, n11365, n11366, n11367, n11368, n11369, n11370, n11371,
         n11372, n11373, n11374, n11375, n11376, n11377, n11378, n11379,
         n11380, n11381, n11382, n11383, n11384, n11385, n11386, n11387,
         n11388, n11389, n11390, n11391, n11392, n11393, n11394, n11395,
         n11396, n11397, n11398, n11399, n11400, n11401, n11402, n11403,
         n11404, n11405, n11406, n11407, n11408, n11409, n11410, n11411,
         n11412, n11413, n11414, n11415, n11416, n11417, n11418, n11419,
         n11420, n11421, n11422, n11423, n11424, n11425, n11426, n11427,
         n11428, n11429, n11430, n11431, n11432, n11433, n11434, n11435,
         n11436, n11437, n11438, n11439, n11440, n11441, n11442, n11443,
         n11444, n11445, n11446, n11447, n11448, n11449, n11450, n11451,
         n11452, n11453, n11454, n11455, n11456, n11457, n11458, n11459,
         n11460, n11461, n11462, n11463, n11464, n11465, n11466, n11467,
         n11468, n11469, n11470, n11471, n11472, n11473, n11474, n11475,
         n11476, n11477, n11478, n11479, n11480, n11481, n11482, n11483,
         n11484, n11485, n11486, n11487, n11488, n11489, n11490, n11491,
         n11492, n11493, n11494, n11495, n11496, n11497, n11498, n11499,
         n11500, n11501, n11502, n11503, n11504, n11505, n11506, n11507,
         n11508, n11509, n11510, n11511, n11512, n11513, n11514, n11515,
         n11516, n11517, n11518, n11519, n11520, n11521, n11522, n11523,
         n11524, n11525, n11526, n11527, n11528, n11529, n11530, n11531,
         n11532, n11533, n11534, n11535, n11536, n11537, n11538, n11539,
         n11540, n11541, n11542, n11543, n11544, n11545, n11546, n11547,
         n11548, n11549, n11550, n11551, n11552, n11553, n11554, n11555,
         n11556, n11557, n11558, n11559, n11560, n11561, n11562, n11563,
         n11564, n11565, n11566, n11567, n11568, n11569, n11570, n11571,
         n11572, n11573, n11574, n11575, n11576, n11577, n11578, n11579,
         n11580, n11581, n11582, n11583, n11584, n11585, n11586, n11587,
         n11588, n11589, n11590, n11591, n11592, n11593, n11594, n11595,
         n11596, n11597, n11598, n11599, n11600, n11601, n11602, n11603,
         n11604, n11605, n11606, n11607, n11608, n11609, n11610, n11611,
         n11612, n11613, n11614, n11615, n11616, n11617, n11618, n11619,
         n11620, n11621, n11622, n11623, n11624, n11625, n11626, n11627,
         n11628, n11629, n11630, n11631, n11632, n11633, n11634, n11635,
         n11636, n11637, n11638, n11639, n11640, n11641, n11642, n11643,
         n11644, n11645, n11646, n11647, n11648, n11649, n11650, n11651,
         n11652, n11653, n11654, n11655, n11656, n11657, n11658, n11659,
         n11660, n11661, n11662, n11663, n11664, n11665, n11666, n11667,
         n11668, n11669, n11670, n11671, n11672, n11673, n11674, n11675,
         n11676, n11677, n11678, n11679, n11680, n11681, n11682, n11683,
         n11684, n11685, n11686, n11687, n11688, n11689, n11690, n11691,
         n11692, n11693, n11694, n11695, n11696, n11697, n11698, n11699,
         n11700, n11701, n11702, n11703, n11704, n11705, n11706, n11707,
         n11708, n11709, n11710, n11711, n11712, n11713, n11714, n11715,
         n11716, n11717, n11718, n11719, n11720, n11721, n11722, n11723,
         n11724, n11725, n11726, n11727, n11728, n11729, n11730, n11731,
         n11732, n11733, n11734, n11735, n11736, n11737, n11738, n11739,
         n11740, n11741, n11742, n11743, n11744, n11745, n11746, n11747,
         n11748, n11749, n11750, n11751, n11752, n11753, n11754, n11755,
         n11756, n11757, n11758, n11759, n11760, n11761, n11762, n11763,
         n11764, n11765, n11766, n11767, n11768, n11769, n11770, n11771,
         n11772, n11773, n11774, n11775, n11776, n11777, n11778, n11779,
         n11780, n11781, n11782, n11783, n11784, n11785, n11786, n11787,
         n11788, n11789, n11790, n11791, n11792, n11793, n11794, n11795,
         n11796, n11797, n11798, n11799, n11800, n11801, n11802, n11803,
         n11804, n11805, n11806, n11807, n11808, n11809, n11810, n11811,
         n11812, n11813, n11814, n11815, n11816, n11817, n11818, n11819,
         n11820, n11821, n11822, n11823, n11824, n11825, n11826, n11827,
         n11828, n11829, n11830, n11831, n11832, n11833, n11834, n11835,
         n11836, n11837, n11838, n11839, n11840, n11841, n11842, n11843,
         n11844, n11845, n11846, n11847, n11848, n11849, n11850, n11851,
         n11852, n11853, n11854, n11855, n11856, n11857, n11858, n11859,
         n11860, n11861, n11862, n11863, n11864, n11865, n11866, n11867,
         n11868, n11869, n11870, n11871, n11872, n11873, n11874, n11875,
         n11876, n11877, n11878, n11879, n11880, n11881, n11882, n11883,
         n11884, n11885, n11886, n11887, n11888, n11889, n11890, n11891,
         n11892, n11893, n11894, n11895, n11896, n11897, n11898, n11899,
         n11900, n11901, n11902, n11903, n11904, n11905, n11906, n11907,
         n11908, n11909, n11910, n11911, n11912, n11913, n11914, n11915,
         n11916, n11917, n11918, n11919, n11920, n11921, n11922, n11923,
         n11924, n11925, n11926, n11927, n11928, n11929, n11930, n11931,
         n11932, n11933, n11934, n11935, n11936, n11937, n11938, n11939,
         n11940, n11941, n11942, n11943, n11944, n11945, n11946, n11947,
         n11948, n11949, n11950, n11951, n11952, n11953, n11954, n11955,
         n11956, n11957, n11958, n11959, n11960, n11961, n11962, n11963,
         n11964, n11965, n11966, n11967, n11968, n11969, n11970, n11971,
         n11972, n11973, n11974, n11975, n11976, n11977, n11978, n11979,
         n11980, n11981, n11982, n11983, n11984, n11985, n11986, n11987,
         n11988, n11989, n11990, n11991, n11992, n11993, n11994, n11995,
         n11996, n11997, n11998, n11999, n12000, n12001, n12002, n12003,
         n12004, n12005, n12006, n12007, n12008, n12009, n12010, n12011,
         n12012, n12013, n12014, n12015, n12016, n12017, n12018, n12019,
         n12020, n12021, n12022, n12023, n12024, n12025, n12026, n12027,
         n12028, n12029, n12030, n12031, n12032, n12033, n12034, n12035,
         n12036, n12037, n12038, n12039, n12040, n12041, n12042, n12043,
         n12044, n12045, n12046, n12047, n12048, n12049, n12050, n12051,
         n12052, n12053, n12054, n12055, n12056, n12057, n12058, n12059,
         n12060, n12061, n12062, n12063, n12064, n12065, n12066, n12067,
         n12068, n12069, n12070, n12071, n12072, n12073, n12074, n12075,
         n12076, n12077, n12078, n12079, n12080, n12081, n12082, n12083,
         n12084, n12085, n12086, n12087, n12088, n12089, n12090, n12091,
         n12092, n12093, n12094, n12095, n12096, n12097, n12098, n12099,
         n12100, n12101, n12102, n12103, n12104, n12105, n12106, n12107,
         n12108, n12109, n12110, n12111, n12112, n12113, n12114, n12115,
         n12116, n12117, n12118, n12119, n12120, n12121, n12122, n12123,
         n12124, n12125, n12126, n12127, n12128, n12129, n12130, n12131,
         n12132, n12133, n12134, n12135, n12136, n12137, n12138, n12139,
         n12140, n12141, n12142, n12143, n12144, n12145, n12146, n12147,
         n12148, n12149, n12150, n12151, n12152, n12153, n12154, n12155,
         n12156, n12157, n12158, n12159, n12160, n12161, n12162, n12163,
         n12164, n12165, n12166, n12167, n12168, n12169, n12170, n12171,
         n12172, n12173, n12174, n12175, n12176, n12177, n12178, n12179,
         n12180, n12181, n12182, n12183, n12184, n12185, n12186, n12187,
         n12188, n12189, n12190, n12191, n12192, n12193, n12194, n12195,
         n12196, n12197, n12198, n12199, n12200, n12201, n12202, n12203,
         n12204, n12205, n12206, n12207, n12208, n12209, n12210, n12211,
         n12212, n12213, n12214, n12215, n12216, n12217, n12218, n12219,
         n12220, n12221, n12222, n12223, n12224, n12225, n12226, n12227,
         n12228, n12229, n12230, n12231, n12232, n12233, n12234, n12235,
         n12236, n12237, n12238, n12239, n12240, n12241, n12242, n12243,
         n12244, n12245, n12246, n12247, n12248, n12249, n12250, n12251,
         n12252, n12253, n12254, n12255, n12256, n12257, n12258, n12259,
         n12260, n12261, n12262, n12263, n12264, n12265, n12266, n12267,
         n12268, n12269, n12270, n12271, n12272, n12273, n12274, n12275,
         n12276, n12277, n12278, n12279, n12280, n12281, n12282, n12283,
         n12284, n12285, n12286, n12287, n12288, n12289, n12290, n12291,
         n12292, n12293, n12294, n12295, n12296, n12297, n12298, n12299,
         n12300, n12301, n12302, n12303, n12304, n12305, n12306, n12307,
         n12308, n12309, n12310, n12311, n12312, n12313, n12314, n12315,
         n12316, n12317, n12318, n12319, n12320, n12321, n12322, n12323,
         n12324, n12325, n12326, n12327, n12328, n12329, n12330, n12331,
         n12332, n12333, n12334, n12335, n12336, n12337, n12338, n12339,
         n12340, n12341, n12342, n12343, n12344, n12345, n12346, n12347,
         n12348, n12349, n12350, n12351, n12352, n12353, n12354, n12355,
         n12356, n12357, n12358, n12359, n12360, n12361, n12362, n12363,
         n12364, n12365, n12366, n12367, n12368, n12369, n12370, n12371,
         n12372, n12373, n12374, n12375, n12376, n12377, n12378, n12379,
         n12380, n12381, n12382, n12383, n12384, n12385, n12386, n12387,
         n12388, n12389, n12390, n12391, n12392, n12393, n12394, n12395,
         n12396, n12397, n12398, n12399, n12400, n12401, n12402, n12403,
         n12404, n12405, n12406, n12407, n12408, n12409, n12410, n12411,
         n12412, n12413, n12414, n12415, n12416, n12417, n12418, n12419,
         n12420, n12421, n12422, n12423, n12424, n12425, n12426, n12427,
         n12428, n12429, n12430, n12431, n12432, n12433, n12434, n12435,
         n12436, n12437, n12438, n12439, n12440, n12441, n12442, n12443,
         n12444, n12445, n12446, n12447, n12448, n12449, n12450, n12451,
         n12452, n12453, n12454, n12455, n12456, n12457, n12458, n12459,
         n12460, n12461, n12462, n12463, n12464, n12465, n12466, n12467,
         n12468, n12469, n12470, n12471, n12472, n12473, n12474, n12475,
         n12476, n12477, n12478, n12479, n12480, n12481, n12482, n12483,
         n12484, n12485, n12486, n12487, n12488, n12489, n12490, n12491,
         n12492, n12493, n12494, n12495, n12496, n12497, n12498, n12499,
         n12500, n12501, n12502, n12503, n12504, n12505, n12506, n12507,
         n12508, n12509, n12510, n12511, n12512, n12513, n12514, n12515,
         n12516, n12517, n12518, n12519, n12520, n12521, n12522, n12523,
         n12524, n12525, n12526, n12527, n12528, n12529, n12530, n12531,
         n12532, n12533, n12534, n12535, n12536, n12537, n12538, n12539,
         n12540, n12541, n12542, n12543, n12544, n12545, n12546, n12547,
         n12548, n12549, n12550, n12551, n12552, n12553, n12554, n12555,
         n12556, n12557, n12558, n12559, n12560, n12561, n12562, n12563,
         n12564, n12565, n12566, n12567, n12568, n12569, n12570, n12571,
         n12572, n12573, n12574, n12575, n12576, n12577, n12578, n12579,
         n12580, n12581, n12582, n12583, n12584, n12585, n12586, n12587,
         n12588, n12589, n12590, n12591, n12592, n12593, n12594, n12595,
         n12596, n12597, n12598, n12599, n12600, n12601, n12602, n12603,
         n12604, n12605, n12606, n12607, n12608, n12609, n12610, n12611,
         n12612, n12613, n12614, n12615, n12616, n12617, n12618, n12619,
         n12620, n12621, n12622, n12623, n12624, n12625, n12626, n12627,
         n12628, n12629, n12630, n12631, n12632, n12633, n12634, n12635,
         n12636, n12637, n12638, n12639, n12640, n12641, n12642, n12643,
         n12644, n12645, n12646, n12647, n12648, n12649, n12650, n12651,
         n12652, n12653, n12654, n12655, n12656, n12657, n12658, n12659,
         n12660, n12661, n12662, n12663, n12664, n12665, n12666, n12667,
         n12668, n12669, n12670, n12671, n12672, n12673, n12674, n12675,
         n12676, n12677, n12678, n12679, n12680, n12681, n12682, n12683,
         n12684, n12685, n12686, n12687, n12688, n12689, n12690, n12691,
         n12692, n12693, n12694, n12695, n12696, n12697, n12698, n12699,
         n12700, n12701, n12702, n12703, n12704, n12705, n12706, n12707,
         n12708, n12709, n12710, n12711, n12712, n12713, n12714, n12715,
         n12716, n12717, n12718, n12719, n12720, n12721, n12722, n12723,
         n12724, n12725, n12726, n12727, n12728, n12729, n12730, n12731,
         n12732, n12733, n12734, n12735, n12736, n12737, n12738, n12739,
         n12740, n12741, n12742, n12743, n12744, n12745, n12746, n12747,
         n12748, n12749, n12750, n12751, n12752, n12753, n12754, n12755,
         n12756, n12757, n12758, n12759, n12760, n12761, n12762, n12763,
         n12764, n12765, n12766, n12767, n12768, n12769, n12770, n12771,
         n12772, n12773, n12774, n12775, n12776, n12777, n12778, n12779,
         n12780, n12781, n12782, n12783, n12784, n12785, n12786, n12787,
         n12788, n12789, n12790, n12791, n12792, n12793, n12794, n12795,
         n12796, n12797, n12798, n12799, n12800, n12801, n12802, n12803,
         n12804, n12805, n12806, n12807, n12808, n12809, n12810, n12811,
         n12812, n12813, n12814, n12815, n12816, n12817, n12818, n12819,
         n12820, n12821, n12822, n12823, n12824, n12825, n12826, n12827,
         n12828, n12829, n12830, n12831, n12832, n12833, n12834, n12835,
         n12836, n12837, n12838, n12839, n12840, n12841, n12842, n12843,
         n12844, n12845, n12846, n12847, n12848, n12849, n12850, n12851,
         n12852, n12853, n12854, n12855, n12856, n12857, n12858, n12859,
         n12860, n12861, n12862, n12863, n12864, n12865, n12866, n12867,
         n12868, n12869, n12870, n12871, n12872, n12873, n12874, n12875,
         n12876, n12877, n12878, n12879, n12880, n12881, n12882, n12883,
         n12884, n12885, n12886, n12887, n12888, n12889, n12890, n12891,
         n12892, n12893, n12894, n12895, n12896, n12897, n12898, n12899,
         n12900, n12901, n12902, n12903, n12904, n12905, n12906, n12907,
         n12908, n12909, n12910, n12911, n12912, n12913, n12914, n12915,
         n12916, n12917, n12918, n12919, n12920, n12921, n12922, n12923,
         n12924, n12925, n12926, n12927, n12929, n12930, n12931, n12932,
         n12933, n12934, n12935, n12936, n12937, n12938, n12939, n12940,
         n12941, n12942, n12943, n12944, n12945, n12946, n12947, n12948,
         n12949, n12950, n12951, n12952, n12953, n12954, n12955, n12956,
         n12957, n12958, n12959, n12960, n12961, n12962, n12963, n12964,
         n12965, n12966, n12967, n12968, n12969, n12970, n12971, n12972,
         n12973, n12974, n12975, n12976, n12977, n12978, n12979, n12980,
         n12981, n12982, n12983, n12984, n12985, n12986, n12987, n12988,
         n12989, n12990, n12991, n12992, n12993, n12994, n12995, n12996,
         n12997, n12998, n12999, n13000, n13001, n13002, n13003, n13004,
         n13005, n13006, n13007, n13008, n13009, n13010, n13011, n13012,
         n13013, n13014, n13015, n13016, n13017, n13018, n13019, n13020,
         n13021, n13022, n13023, n13024, n13025, n13026, n13027, n13028,
         n13029, n13030, n13031, n13032, n13033, n13034, n13035, n13036,
         n13037, n13038, n13039, n13040, n13041, n13042, n13043, n13044,
         n13045, n13046, n13047, n13048, n13049, n13050, n13051, n13052,
         n13053, n13054, n13055, n13056, n13057, n13058, n13059, n13060,
         n13061, n13062, n13063, n13064, n13065, n13066, n13067, n13068,
         n13069, n13070, n13071, n13072, n13073, n13074, n13075, n13076,
         n13077, n13078, n13079, n13080, n13081, n13082, n13083, n13084,
         n13085, n13086, n13087, n13088, n13089, n13090, n13091, n13092,
         n13093, n13094, n13095, n13096, n13097, n13098, n13099, n13100,
         n13101, n13102, n13103, n13104, n13105, n13106, n13107, n13108,
         n13109, n13110, n13111, n13112, n13113, n13114, n13115, n13116,
         n13117, n13118, n13119, n13120, n13121, n13122, n13123, n13124,
         n13125, n13126, n13127, n13128, n13129, n13130, n13131, n13132,
         n13133, n13134, n13135, n13136, n13137, n13138, n13139, n13140,
         n13141, n13142, n13143, n13144, n13145, n13146, n13147, n13148,
         n13149, n13150, n13151, n13152, n13153, n13154, n13155, n13156,
         n13157, n13158, n13159, n13160, n13161, n13162, n13163, n13164,
         n13165, n13166, n13167, n13168, n13169, n13170, n13171, n13172,
         n13173, n13174, n13175, n13176, n13177, n13178, n13179, n13180,
         n13181, n13182, n13183, n13184, n13185, n13186, n13187, n13188,
         n13189, n13190, n13191, n13192, n13193, n13194, n13195, n13196,
         n13197, n13198, n13199, n13200, n13201, n13202, n13203, n13204,
         n13205, n13206, n13207, n13208, n13209, n13210, n13211, n13212,
         n13213, n13214, n13215, n13216, n13217, n13218, n13219, n13220,
         n13221, n13222, n13223, n13224, n13225, n13226, n13227, n13228,
         n13229, n13230, n13231, n13232, n13233, n13234, n13235, n13236,
         n13237, n13238, n13239, n13240, n13241, n13242, n13243, n13244,
         n13245, n13246, n13247, n13248, n13249, n13250, n13251, n13252,
         n13253, n13254, n13255, n13256, n13257, n13258, n13259, n13260,
         n13261, n13262, n13263, n13264, n13265, n13266, n13267, n13268,
         n13269, n13270, n13271, n13272, n13273, n13274, n13275, n13276,
         n13277, n13278, n13279, n13280, n13281, n13282, n13283, n13284,
         n13285, n13286, n13287, n13288, n13289, n13290, n13291, n13292,
         n13293, n13294, n13295, n13296, n13297, n13298, n13299, n13300,
         n13301, n13302, n13303, n13304, n13305, n13306, n13307, n13308,
         n13309, n13310, n13311, n13312, n13313, n13314, n13315, n13316,
         n13317, n13318, n13319, n13320, n13321, n13322, n13323, n13324,
         n13325, n13326, n13327, n13328, n13329, n13330, n13331, n13332,
         n13333, n13334, n13335, n13336, n13337, n13338, n13339, n13340,
         n13341, n13342, n13343, n13344, n13345, n13346, n13347, n13348,
         n13349, n13350, n13351, n13352, n13353, n13354, n13355, n13356,
         n13357, n13358, n13359, n13360, n13361, n13362, n13363, n13364,
         n13365, n13366, n13367, n13368, n13369, n13370, n13371, n13372,
         n13373, n13374, n13375, n13376, n13377, n13378, n13379, n13380,
         n13381, n13382, n13383, n13384, n13385, n13386, n13387, n13388,
         n13389, n13390, n13391, n13392, n13393, n13394, n13395, n13396,
         n13397, n13398, n13399, n13400, n13401, n13402, n13403, n13404,
         n13405, n13406, n13407, n13408, n13409, n13410, n13411, n13412,
         n13413, n13414, n13415, n13416, n13417, n13418, n13419, n13420,
         n13421, n13422, n13423, n13424, n13425, n13426, n13427, n13428,
         n13429, n13430, n13431, n13432, n13433, n13434, n13435, n13436,
         n13437, n13438, n13439, n13440, n13441, n13442, n13443, n13444,
         n13445, n13446, n13447, n13448, n13449, n13450, n13451, n13452,
         n13453, n13454, n13455, n13456, n13457, n13458, n13459, n13460,
         n13461, n13462, n13463, n13464, n13465, n13466, n13467, n13468,
         n13469, n13470, n13471, n13472, n13473, n13474, n13475, n13476,
         n13477, n13478, n13479, n13480, n13481, n13482, n13483, n13484,
         n13485, n13486, n13487, n13488, n13489, n13490, n13491, n13492,
         n13493, n13494, n13495, n13496, n13497, n13498, n13499, n13500,
         n13501, n13502, n13503, n13504, n13505, n13506, n13507, n13508,
         n13509, n13510, n13511, n13512, n13513, n13514, n13515, n13516,
         n13517, n13518, n13519, n13520, n13521, n13522, n13523, n13524,
         n13525, n13526, n13527, n13528, n13529, n13530, n13531, n13532,
         n13533, n13534, n13535, n13536, n13537, n13538, n13539, n13540,
         n13541, n13542, n13543, n13544, n13545, n13546, n13547, n13548,
         n13549, n13550, n13551, n13552, n13553, n13554, n13555, n13556,
         n13557, n13558, n13559, n13560, n13561, n13562, n13563, n13564,
         n13565, n13566, n13567, n13568, n13569, n13570, n13571, n13572,
         n13573, n13574, n13575, n13576, n13577, n13578, n13579, n13580,
         n13581, n13582, n13583, n13584, n13585, n13586, n13587, n13588,
         n13589, n13590, n13591, n13592, n13593, n13594, n13595, n13596,
         n13597, n13598, n13599, n13600, n13601, n13602, n13603, n13604,
         n13605, n13606, n13607, n13608, n13609, n13610, n13611, n13612,
         n13613, n13614, n13615, n13616, n13617, n13618, n13619, n13620,
         n13621, n13622, n13623, n13624, n13625, n13626, n13627, n13628,
         n13629, n13630, n13631, n13632, n13633, n13634, n13635, n13636,
         n13637, n13638, n13639, n13640, n13641, n13642, n13643, n13644,
         n13645, n13646, n13647, n13648, n13649, n13650, n13651, n13652,
         n13653, n13654, n13655, n13656, n13657, n13658, n13659, n13660,
         n13661, n13662, n13663, n13664, n13665, n13666, n13667, n13668,
         n13669, n13670, n13671, n13672, n13673, n13674, n13675, n13676,
         n13677, n13678, n13679, n13680, n13681, n13682, n13683, n13684,
         n13685, n13686, n13687, n13688, n13689, n13690, n13691, n13692,
         n13693, n13694, n13695, n13696, n13697, n13698, n13699, n13700,
         n13701, n13702, n13703, n13704, n13705, n13706, n13707, n13708,
         n13709, n13710, n13711, n13712, n13713, n13714, n13715, n13716,
         n13717, n13718, n13719, n13720, n13721, n13722, n13723, n13724,
         n13725, n13726, n13727, n13728, n13729, n13730, n13731, n13732,
         n13733, n13734, n13735, n13736, n13737, n13738, n13739, n13740,
         n13741, n13742, n13743, n13744, n13745, n13746, n13747, n13748,
         n13749, n13750, n13751, n13752, n13753, n13754, n13755, n13756,
         n13757, n13758, n13759, n13760, n13761, n13762, n13763, n13764,
         n13765, n13766, n13767, n13768, n13769, n13770, n13771, n13772,
         n13773, n13774, n13775, n13776, n13777, n13778, n13779, n13780,
         n13781, n13782, n13783, n13784, n13785, n13786, n13787, n13788,
         n13789, n13790, n13791, n13792, n13793, n13794, n13795, n13796,
         n13797, n13798, n13799, n13800, n13801, n13802, n13803, n13804,
         n13805, n13806, n13807, n13808, n13809, n13810, n13811, n13812,
         n13813, n13814, n13815, n13816, n13817, n13818, n13819, n13820,
         n13821, n13822, n13823, n13824, n13825, n13826, n13827, n13828,
         n13829, n13830, n13831, n13832, n13833, n13834, n13835, n13836,
         n13837, n13838, n13839, n13840, n13841, n13842, n13843, n13844,
         n13845, n13846, n13847, n13848, n13849, n13850, n13851, n13852,
         n13853, n13854, n13855, n13856, n13857, n13858, n13859, n13860,
         n13861, n13862, n13863, n13864, n13865, n13866, n13867, n13868,
         n13869, n13870, n13871, n13872, n13873, n13874, n13875, n13876,
         n13877, n13878, n13879, n13880, n13881, n13882, n13883, n13884,
         n13885, n13886, n13887, n13888, n13889, n13890, n13891, n13892,
         n13893, n13894, n13895, n13896, n13897, n13898, n13899, n13900,
         n13901, n13902, n13903, n13904, n13905, n13906, n13907, n13908,
         n13909, n13910, n13911, n13912, n13913, n13914, n13915, n13916,
         n13917, n13918, n13919, n13920, n13921, n13922, n13923, n13924,
         n13925, n13926, n13927, n13928, n13929, n13930, n13931, n13932,
         n13933, n13934, n13935, n13936, n13937, n13938, n13939, n13940,
         n13941, n13942, n13943, n13944, n13945, n13946, n13947, n13948,
         n13949, n13950, n13951, n13952, n13953, n13954, n13955, n13956,
         n13957, n13958, n13959, n13960, n13961, n13962, n13963, n13964,
         n13965, n13966, n13967, n13968, n13969, n13970, n13971, n13972,
         n13973, n13974, n13975, n13976, n13977, n13978, n13979, n13980,
         n13981, n13982, n13983, n13984, n13985, n13986, n13987, n13988,
         n13989, n13990, n13991, n13992, n13993, n13994, n13995, n13996,
         n13997, n13998, n13999, n14000, n14001, n14002, n14003, n14004,
         n14005, n14006, n14007, n14008, n14009, n14010, n14011, n14012,
         n14013, n14014, n14015, n14016, n14017, n14018, n14019, n14020,
         n14021, n14022, n14023, n14024, n14025, n14026, n14027, n14028,
         n14029, n14030, n14031, n14032, n14033, n14034, n14035, n14036,
         n14037, n14038, n14039, n14040, n14041, n14042, n14043, n14044,
         n14045, n14046, n14047, n14048, n14049, n14050, n14051, n14052,
         n14053, n14054, n14055, n14056, n14057, n14058, n14059, n14060,
         n14061, n14062, n14063, n14064, n14065, n14066, n14067, n14068,
         n14069, n14070, n14071, n14072, n14073, n14074, n14075, n14076,
         n14077, n14078, n14079, n14080, n14081, n14082, n14083, n14084,
         n14085, n14086, n14087, n14088, n14089, n14090, n14091, n14092,
         n14093, n14094, n14095, n14096, n14097, n14098, n14099, n14100,
         n14101, n14102, n14103, n14104, n14105, n14106, n14107, n14108,
         n14109, n14110, n14111, n14112, n14113, n14114, n14115, n14116,
         n14117, n14118, n14119, n14120, n14121, n14122, n14123, n14124,
         n14125, n14126, n14127, n14128, n14129, n14130, n14131, n14132,
         n14133, n14134, n14135, n14136, n14137, n14138, n14139, n14140,
         n14141, n14142, n14143, n14144, n14145, n14146, n14147, n14148,
         n14149, n14150, n14151, n14152, n14153, n14154, n14155, n14156,
         n14157, n14158, n14159, n14160, n14161, n14162, n14163, n14164,
         n14165, n14166, n14167, n14168, n14169, n14170, n14171, n14172,
         n14173, n14174, n14175, n14176, n14177, n14178, n14179, n14180,
         n14181, n14182, n14183, n14184, n14185, n14186, n14187, n14188,
         n14189, n14190, n14191, n14192, n14193, n14194, n14195, n14196,
         n14197, n14198, n14199, n14200, n14201, n14202, n14203, n14204,
         n14205, n14206, n14207, n14208, n14209, n14210, n14211, n14212,
         n14213, n14214, n14215, n14216, n14217, n14218, n14219, n14220,
         n14221, n14222, n14223, n14224, n14225, n14226, n14227, n14228,
         n14229, n14230, n14231, n14232, n14233, n14234, n14235, n14236,
         n14237, n14238, n14239, n14240, n14241, n14242, n14243, n14244,
         n14245, n14246, n14247, n14248, n14249, n14250, n14251, n14252,
         n14253, n14254, n14255, n14256, n14257, n14258, n14259, n14260,
         n14261, n14262, n14263, n14264, n14265, n14266, n14267, n14268,
         n14269, n14270, n14271, n14272, n14273, n14274, n14275, n14276,
         n14277, n14278, n14279, n14280, n14281, n14282, n14283, n14284,
         n14285, n14286, n14287, n14288, n14289, n14290, n14291, n14292,
         n14293, n14294, n14295, n14296, n14297, n14298, n14299, n14300,
         n14301, n14302, n14303, n14304, n14305, n14306, n14307, n14308,
         n14309, n14310, n14311, n14312, n14313, n14314, n14315, n14316,
         n14317, n14318, n14319, n14320, n14321, n14322, n14323, n14324,
         n14325, n14326, n14327, n14328, n14329, n14330, n14331, n14332,
         n14333, n14334, n14335, n14336, n14337, n14338, n14339, n14340,
         n14341, n14342, n14343, n14344, n14345, n14346, n14347, n14348,
         n14349, n14350, n14351, n14352, n14353, n14354, n14355, n14356,
         n14357, n14358, n14359, n14360, n14361, n14362, n14363, n14364,
         n14365, n14366, n14367, n14368, n14369, n14370, n14371, n14372,
         n14373, n14374, n14375, n14376, n14377, n14378, n14379, n14380,
         n14381, n14382, n14383, n14384, n14385, n14386, n14387, n14388,
         n14389, n14390, n14391, n14392, n14393, n14394, n14395, n14396,
         n14397, n14398, n14399, n14400, n14401, n14402, n14403, n14404,
         n14405, n14406, n14407, n14408, n14409, n14410, n14411, n14412,
         n14413, n14414, n14415, n14416, n14417, n14418, n14419, n14420,
         n14421, n14422, n14423, n14424, n14425, n14426, n14427, n14428,
         n14429, n14430, n14431, n14432, n14433, n14434, n14435, n14436,
         n14437, n14438, n14439, n14440, n14441, n14442, n14443, n14444,
         n14445, n14446, n14447, n14448, n14449, n14450, n14451, n14452,
         n14453, n14454, n14455, n14456, n14457, n14458, n14459, n14460,
         n14461, n14462, n14463, n14464, n14465, n14466, n14467, n14468,
         n14470, n14471, n14472, n14473, n14474, n14475, n14476, n14477,
         n14478, n14479, n14480, n14481, n14482, n14483, n14484, n14485,
         n14486, n14487, n14488, n14489, n14490, n14491, n14492, n14493,
         n14494, n14495, n14496, n14497, n14498, n14499, n14500, n14501,
         n14502, n14503, n14504, n14505, n14506, n14507, n14508, n14509,
         n14510, n14511, n14512, n14513, n14514, n14515, n14516, n14517,
         n14518, n14519, n14520, n14521, n14522, n14523, n14524, n14525,
         n14526, n14527, n14528, n14529, n14530, n14531, n14532, n14533,
         n14534, n14535, n14536, n14537, n14538, n14539, n14540, n14541,
         n14542, n14543, n14544, n14545, n14546, n14547, n14548, n14549,
         n14550, n14551, n14552, n14553, n14554, n14555, n14556, n14557,
         n14558, n14559, n14560, n14561, n14562, n14563, n14564, n14565,
         n14566, n14567, n14568, n14569, n14570, n14571, n14572, n14573,
         n14574, n14575, n14576, n14577, n14578, n14579, n14580, n14581,
         n14582, n14583, n14584, n14585, n14586, n14587, n14588, n14589,
         n14590, n14591, n14592, n14593, n14594, n14595, n14596, n14597,
         n14598, n14599, n14600, n14601, n14602, n14603, n14604, n14605,
         n14606, n14607, n14608, n14609, n14610, n14611, n14612, n14613,
         n14614, n14615, n14616, n14617, n14618, n14619, n14620, n14621,
         n14622, n14623, n14624, n14625, n14626, n14627, n14628, n14629,
         n14630, n14631, n14632, n14633, n14634, n14635, n14636, n14637,
         n14638, n14639, n14640, n14641, n14642, n14643, n14644, n14645,
         n14646, n14647, n14648, n14649, n14650, n14651, n14652, n14653,
         n14654, n14655, n14656, n14657, n14658, n14659, n14660, n14661,
         n14662, n14663, n14664, n14665, n14666, n14667, n14668, n14669,
         n14670, n14671, n14672, n14673, n14674, n14675, n14676, n14677,
         n14678, n14679, n14680, n14681, n14682, n14683, n14684, n14685,
         n14686, n14687, n14688, n14689, n14690, n14691, n14692, n14693,
         n14694, n14695, n14696, n14697, n14698, n14699, n14700, n14701,
         n14702, n14703, n14704, n14705, n14706, n14707, n14708, n14709,
         n14710, n14711, n14712, n14713, n14714, n14715, n14716, n14717,
         n14718, n14719, n14720, n14721, n14722, n14723, n14724, n14725,
         n14726, n14727, n14728, n14729, n14730, n14731, n14732, n14733,
         n14734, n14735, n14736, n14737, n14738, n14739, n14740, n14741,
         n14742, n14743, n14744, n14745, n14746, n14747, n14748, n14749,
         n14750, n14751, n14752, n14753, n14754, n14755, n14756, n14757,
         n14758, n14759, n14760, n14761, n14762, n14763, n14764, n14765,
         n14766, n14767, n14768, n14769, n14770, n14771, n14772, n14773,
         n14774, n14775, n14776, n14777, n14778, n14779, n14780, n14781,
         n14782, n14783, n14784, n14785, n14786, n14787, n14788, n14789,
         n14790, n14791, n14792, n14793, n14794, n14795, n14796, n14797,
         n14798, n14799, n14800, n14801, n14802, n14803, n14804, n14805,
         n14806, n14807, n14808, n14809, n14810, n14811, n14812, n14813,
         n14814, n14815, n14816, n14817, n14818, n14819, n14820, n14821,
         n14822, n14823, n14824, n14825, n14826, n14827, n14828, n14829,
         n14830, n14831, n14832, n14833, n14834, n14835, n14836, n14837,
         n14838, n14839, n14840, n14841, n14842, n14843, n14844, n14845,
         n14846, n14847, n14848, n14849, n14850, n14851, n14852, n14853,
         n14854, n14855, n14856, n14857, n14858, n14859, n14860, n14861,
         n14862, n14863, n14864, n14865, n14866, n14867, n14868, n14869,
         n14870, n14871, n14872, n14873, n14874, n14875, n14876, n14877,
         n14878, n14879, n14880, n14881, n14882, n14883, n14884, n14885,
         n14886, n14887, n14888, n14889, n14890, n14891, n14892, n14893,
         n14894, n14895, n14896, n14897, n14898, n14899, n14900, n14901,
         n14902, n14903, n14904, n14905, n14906, n14907, n14908, n14909,
         n14910, n14911, n14912, n14913, n14914, n14915, n14916, n14917,
         n14918, n14919, n14920, n14921, n14922, n14923, n14924, n14925,
         n14926, n14927, n14928, n14929, n14930, n14931, n14932, n14933,
         n14934, n14935, n14936, n14937, n14938, n14939, n14940, n14941,
         n14942, n14943, n14944, n14945, n14946, n14947, n14948, n14949,
         n14950, n14951, n14952, n14953, n14954, n14955, n14956, n14957,
         n14958, n14959, n14960, n14961, n14962, n14963, n14964, n14965,
         n14966, n14967, n14968, n14969, n14970, n14971, n14972, n14973,
         n14974, n14975, n14976, n14977, n14978, n14979, n14980, n14981,
         n14982, n14983, n14984, n14985, n14986, n14987, n14988, n14989,
         n14990, n14991, n14992, n14993, n14994, n14995, n14996, n14997,
         n14998, n14999, n15000, n15001, n15002, n15003, n15004, n15005,
         n15006, n15007, n15008, n15009, n15010, n15011, n15012, n15013,
         n15014, n15015, n15016, n15017, n15018, n15019, n15020, n15021,
         n15022, n15023, n15024, n15025, n15026, n15027, n15028, n15029,
         n15030, n15031, n15032, n15033, n15034, n15035, n15036, n15037,
         n15038, n15039, n15040, n15041, n15042, n15043, n15044, n15045,
         n15046, n15047, n15048, n15049, n15050, n15051, n15052, n15053,
         n15054, n15055, n15056, n15057, n15058, n15059, n15060, n15061,
         n15062, n15063, n15064, n15065, n15066, n15067, n15068, n15069,
         n15070, n15071, n15072, n15073, n15074, n15075, n15076, n15077,
         n15078, n15079, n15080, n15081, n15082, n15083, n15084, n15085,
         n15086, n15087, n15088, n15089, n15090, n15091, n15092, n15093,
         n15094, n15095, n15096, n15097, n15098, n15099, n15100, n15101,
         n15102, n15103, n15104, n15105, n15106, n15107, n15108, n15109,
         n15110, n15111, n15112, n15113, n15114, n15115, n15116, n15117,
         n15118, n15119, n15120, n15121, n15122, n15123, n15124, n15125,
         n15126, n15127, n15128, n15129, n15130, n15131, n15132, n15133,
         n15134, n15135, n15136, n15137, n15138, n15139, n15140, n15141,
         n15142, n15143, n15144, n15145, n15146, n15147, n15148, n15149,
         n15150, n15151, n15152, n15153, n15154, n15155, n15156, n15157,
         n15158, n15159, n15160, n15161, n15162, n15163, n15164, n15165,
         n15166, n15167, n15168, n15169, n15170, n15171, n15172, n15173,
         n15174, n15175, n15176, n15177, n15178, n15179, n15180, n15181,
         n15182, n15183, n15184, n15185, n15186, n15187, n15188, n15189,
         n15190, n15191, n15192, n15193, n15194, n15195, n15196, n15197,
         n15198, n15199, n15200, n15201, n15202, n15203, n15204, n15205,
         n15206, n15207, n15208, n15209, n15210, n15211, n15212, n15213,
         n15214, n15215, n15216, n15217, n15218, n15219, n15220, n15221,
         n15222, n15223, n15224, n15225, n15226, n15227, n15228, n15229,
         n15230, n15231, n15232, n15233, n15234, n15235, n15236, n15237,
         n15238, n15239, n15240, n15241, n15242, n15243, n15244, n15245,
         n15246, n15247, n15248, n15249, n15250, n15251, n15252, n15253,
         n15254, n15255, n15256, n15257, n15258, n15259, n15260, n15261,
         n15262, n15263, n15264, n15265, n15266, n15267, n15268, n15269,
         n15270, n15271, n15272, n15273, n15274, n15275, n15276, n15277,
         n15278, n15279, n15280, n15281, n15282, n15283, n15284, n15285,
         n15286, n15287, n15288, n15289, n15290, n15291, n15292, n15293,
         n15294, n15295, n15296, n15297, n15298, n15299, n15300, n15301,
         n15302, n15303, n15304, n15305, n15306, n15307, n15308, n15309,
         n15310, n15311, n15312, n15313, n15314, n15315, n15316, n15317,
         n15318, n15319, n15320, n15321, n15322, n15323, n15324, n15325,
         n15326, n15327, n15328, n15329, n15330, n15331, n15332, n15333,
         n15334, n15335, n15336, n15337, n15338, n15339, n15340, n15341,
         n15342, n15343, n15344, n15345, n15346, n15347, n15348, n15349,
         n15350, n15351, n15352, n15353, n15354, n15355, n15356, n15357,
         n15358, n15359, n15360, n15361, n15362, n15363, n15364, n15365,
         n15366, n15367, n15368, n15369, n15370, n15371, n15372, n15373,
         n15374, n15375, n15376, n15377, n15378, n15379, n15380, n15381,
         n15382, n15383, n15384, n15385, n15386, n15387, n15388, n15389,
         n15390, n15391, n15392, n15393, n15394, n15395, n15396, n15397,
         n15398, n15399, n15400, n15401, n15402, n15403, n15404, n15405,
         n15406, n15407, n15408, n15409, n15410, n15411, n15412, n15413,
         n15414, n15415, n15416, n15417, n15418, n15419, n15420, n15421,
         n15422, n15423, n15424, n15425, n15426, n15427, n15428, n15429,
         n15430, n15431, n15432, n15433, n15434, n15435, n15436, n15437,
         n15438, n15439, n15440, n15441, n15442, n15443, n15444, n15445,
         n15446, n15447, n15448, n15449, n15450, n15451, n15452, n15453,
         n15454, n15455, n15456, n15457, n15458, n15459, n15460, n15461,
         n15462, n15463, n15464, n15465, n15466, n15467, n15468, n15469,
         n15470, n15471, n15472, n15473, n15474, n15475, n15476, n15477,
         n15478, n15479, n15480, n15481, n15482, n15483, n15484, n15485,
         n15486, n15487, n15488, n15489, n15490, n15491, n15492, n15493,
         n15494, n15495, n15496, n15497, n15498, n15499, n15500, n15501,
         n15502, n15503, n15504, n15505, n15506, n15507, n15508, n15509,
         n15510, n15511, n15512, n15513, n15514, n15515, n15516, n15517,
         n15518, n15519, n15520, n15521, n15522, n15523, n15525, n15526,
         n15527, n15528, n15529, n15530, n15531, n15532, n15533, n15534,
         n15535, n15536, n15537, n15538, n15539, n15540, n15541, n15542,
         n15543, n15544, n15545, n15546, n15547, n15548, n15549, n15550,
         n15551, n15552, n15553, n15554, n15555, n15556, n15557, n15558,
         n15559, n15560, n15561, n15562, n15563, n15564, n15565, n15566,
         n15567, n15568, n15569, n15570, n15571, n15572, n15573, n15574,
         n15575, n15576, n15577, n15578, n15579, n15580, n15581, n15582,
         n15583, n15584, n15585, n15586, n15587, n15588, n15589, n15590,
         n15591, n15592, n15593, n15594, n15595, n15596, n15597, n15598,
         n15599, n15600, n15601, n15602, n15603, n15604, n15605, n15606,
         n15607, n15608, n15609, n15610, n15611, n15612, n15613, n15614,
         n15615, n15616, n15617, n15618, n15619, n15620, n15621, n15622,
         n15623, n15624, n15625, n15626, n15627, n15628, n15629, n15630,
         n15631, n15632, n15633, n15634, n15635, n15636, n15637, n15638,
         n15639, n15640, n15641, n15642, n15643, n15644, n15645, n15646,
         n15647, n15648, n15649, n15650, n15651, n15652, n15653, n15654,
         n15655, n15656, n15657, n15658, n15659, n15660, n15661, n15662,
         n15663, n15664, n15665, n15666, n15667, n15668, n15669, n15670,
         n15671, n15672, n15673, n15674, n15675, n15676, n15677, n15678,
         n15679, n15680, n15681, n15682, n15683, n15684, n15685, n15686,
         n15687, n15688, n15689, n15690, n15691, n15692, n15693, n15694,
         n15695, n15696, n15697, n15698, n15699, n15700, n15701, n15702,
         n15703, n15704, n15705, n15706, n15707, n15708, n15709, n15710,
         n15711, n15712, n15713, n15714, n15715, n15716, n15717, n15718,
         n15719, n15720, n15721, n15722, n15723, n15724, n15725, n15726,
         n15727, n15728, n15729, n15730, n15731, n15732, n15733, n15734,
         n15735, n15736, n15737, n15738, n15739, n15740, n15741, n15742,
         n15743, n15744, n15745, n15746, n15747, n15748, n15749, n15750,
         n15751, n15752, n15753, n15754, n15755, n15756, n15757, n15758,
         n15759, n15760, n15761, n15762, n15763, n15764, n15765, n15766,
         n15767, n15768, n15769, n15770, n15771, n15772, n15773, n15774,
         n15775, n15776, n15777, n15778, n15779, n15780, n15781, n15782,
         n15783, n15784, n15785, n15786, n15787, n15788, n15789, n15790,
         n15791, n15792, n15793, n15794, n15795, n15796, n15797, n15798,
         n15799, n15800, n15801, n15802, n15803, n15804, n15805, n15806,
         n15807, n15808, n15809, n15810, n15811, n15812, n15813, n15814,
         n15815, n15816, n15817, n15818, n15819, n15820, n15821, n15822,
         n15823, n15824, n15825, n15826, n15827, n15828, n15829, n15830,
         n15831, n15832, n15833, n15834, n15835, n15836, n15837, n15838,
         n15839, n15840, n15841, n15842, n15843, n15844, n15845, n15846,
         n15847, n15848, n15849, n15850, n15851, n15852, n15853, n15854,
         n15855, n15856, n15857, n15858, n15859, n15860, n15861, n15862,
         n15863, n15864, n15865, n15866, n15867, n15868, n15869, n15870,
         n15871, n15872, n15873, n15874, n15875, n15876, n15877, n15878,
         n15879, n15880, n15881, n15882, n15883, n15884, n15885, n15886,
         n15887, n15888, n15889, n15890, n15891, n15892, n15893, n15894,
         n15895, n15896, n15897, n15898, n15899, n15900, n15901, n15902,
         n15903, n15904, n15905, n15906, n15907, n15908, n15909, n15910,
         n15911, n15912, n15913, n15914, n15915, n15916, n15917, n15918,
         n15919, n15920, n15921, n15922, n15923, n15924, n15925, n15926,
         n15927, n15928, n15929, n15930, n15931, n15932, n15933, n15934,
         n15935, n15936, n15937, n15938, n15939, n15940, n15941, n15942,
         n15943, n15944, n15945, n15946, n15947, n15948, n15949, n15950,
         n15951, n15952, n15953, n15954, n15955, n15956, n15957, n15958,
         n15959, n15960, n15961, n15962, n15963, n15964, n15965, n15966,
         n15967, n15968, n15969, n15970, n15971, n15972, n15973, n15974,
         n15975, n15976, n15977, n15978, n15979, n15980, n15981, n15982,
         n15983, n15984, n15985, n15986;

  NAND2_X1 U7270 ( .A1(n8612), .A2(n12616), .ZN(n12397) );
  AND2_X1 U7271 ( .A1(n10495), .A2(n10494), .ZN(n14823) );
  OR2_X1 U7272 ( .A1(n10531), .A2(n10530), .ZN(n15132) );
  INV_X1 U7273 ( .A(n15200), .ZN(n15191) );
  OR2_X1 U7274 ( .A1(n15194), .A2(n15212), .ZN(n12729) );
  NAND2_X1 U7275 ( .A1(n10338), .A2(n10337), .ZN(n14478) );
  OR2_X1 U7276 ( .A1(n9014), .A2(n9013), .ZN(n9035) );
  AND3_X1 U7277 ( .A1(n9565), .A2(n9564), .A3(n9563), .ZN(n11506) );
  NAND2_X2 U7278 ( .A1(n14706), .A2(n9178), .ZN(n14529) );
  INV_X1 U7279 ( .A(n8214), .ZN(n12423) );
  INV_X2 U7280 ( .A(n9856), .ZN(n6529) );
  NOR2_X1 U7281 ( .A1(n15550), .A2(n15542), .ZN(n9217) );
  INV_X1 U7282 ( .A(n12461), .ZN(n13128) );
  NAND2_X1 U7283 ( .A1(n8746), .A2(n8747), .ZN(n14725) );
  INV_X2 U7284 ( .A(P3_ADDR_REG_2__SCAN_IN), .ZN(n15556) );
  INV_X1 U7285 ( .A(n14834), .ZN(n10533) );
  CLKBUF_X1 U7286 ( .A(n10692), .Z(n6523) );
  AND2_X1 U7287 ( .A1(n8216), .A2(n7782), .ZN(n6984) );
  INV_X1 U7288 ( .A(n14719), .ZN(n14824) );
  INV_X1 U7290 ( .A(n12626), .ZN(n12598) );
  XNOR2_X1 U7291 ( .A(n14299), .B(n13787), .ZN(n14018) );
  NAND2_X1 U7292 ( .A1(n6749), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n9183) );
  NAND2_X1 U7293 ( .A1(n6545), .A2(n15191), .ZN(n6842) );
  NAND3_X1 U7294 ( .A1(n7940), .A2(n7939), .A3(n8722), .ZN(n8997) );
  NOR2_X1 U7295 ( .A1(P1_ADDR_REG_2__SCAN_IN), .A2(n15556), .ZN(n15558) );
  INV_X1 U7296 ( .A(n12832), .ZN(n12792) );
  INV_X1 U7297 ( .A(n8287), .ZN(n8492) );
  NAND2_X1 U7298 ( .A1(n6847), .A2(n6846), .ZN(n13197) );
  NAND3_X1 U7299 ( .A1(n8242), .A2(n7313), .A3(n7312), .ZN(n11761) );
  XNOR2_X1 U7300 ( .A(n13423), .B(n12939), .ZN(n12615) );
  INV_X1 U7301 ( .A(n8214), .ZN(n12410) );
  NAND2_X1 U7302 ( .A1(n8602), .A2(n12580), .ZN(n13297) );
  NAND2_X1 U7303 ( .A1(n7828), .A2(n7826), .ZN(n8213) );
  NAND2_X1 U7305 ( .A1(n9904), .A2(n9903), .ZN(n14299) );
  INV_X1 U7306 ( .A(n11930), .ZN(n10197) );
  CLKBUF_X2 U7307 ( .A(n14307), .Z(n15891) );
  INV_X1 U7308 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n14451) );
  NAND2_X1 U7310 ( .A1(n8958), .A2(n8871), .ZN(n8907) );
  NAND2_X1 U7311 ( .A1(n7444), .A2(n7443), .ZN(n8788) );
  INV_X1 U7312 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n8645) );
  AOI21_X1 U7313 ( .B1(P1_ADDR_REG_2__SCAN_IN), .B2(n15556), .A(n15558), .ZN(
        n15584) );
  OAI21_X1 U7314 ( .B1(n15650), .B2(P2_ADDR_REG_8__SCAN_IN), .A(n6600), .ZN(
        n7394) );
  NAND2_X1 U7315 ( .A1(n8532), .A2(n8531), .ZN(n13423) );
  OAI21_X1 U7316 ( .B1(n8213), .B2(n8084), .A(n8083), .ZN(n8264) );
  NAND2_X1 U7317 ( .A1(n7440), .A2(n7357), .ZN(n9493) );
  XNOR2_X1 U7318 ( .A(n15252), .B(n15409), .ZN(n15262) );
  NAND2_X1 U7319 ( .A1(n15135), .A2(n15294), .ZN(n15312) );
  AND2_X1 U7320 ( .A1(n7397), .A2(n7396), .ZN(n15682) );
  INV_X1 U7321 ( .A(n12493), .ZN(n12490) );
  NAND2_X1 U7322 ( .A1(n10540), .A2(n10539), .ZN(n15139) );
  INV_X1 U7323 ( .A(n11849), .ZN(n14969) );
  INV_X2 U7324 ( .A(n15312), .ZN(n15286) );
  OR2_X1 U7325 ( .A1(n12637), .A2(n12636), .ZN(n6522) );
  OR2_X2 U7326 ( .A1(n12217), .A2(n8600), .ZN(n7781) );
  XNOR2_X2 U7327 ( .A(n13015), .B(n13027), .ZN(n13017) );
  AOI22_X2 U7328 ( .A1(n13010), .A2(n13009), .B1(P3_REG1_REG_12__SCAN_IN), 
        .B2(n13008), .ZN(n13015) );
  NAND2_X2 U7329 ( .A1(n12736), .A2(n12735), .ZN(n15153) );
  NOR2_X2 U7330 ( .A1(n15694), .A2(n7389), .ZN(n15661) );
  NAND2_X2 U7331 ( .A1(n12973), .A2(n12972), .ZN(n13010) );
  XNOR2_X2 U7332 ( .A(n12792), .B(n11760), .ZN(n11802) );
  NAND4_X4 U7333 ( .A1(n8716), .A2(n8715), .A3(n8714), .A4(n8713), .ZN(n14970)
         );
  NAND3_X2 U7334 ( .A1(n8643), .A2(n7879), .A3(n8938), .ZN(n7308) );
  AOI21_X2 U7335 ( .B1(n15366), .B2(n15812), .A(n6655), .ZN(n8042) );
  AOI211_X1 U7336 ( .C1(n14725), .C2(n15701), .A(n11889), .B(n11886), .ZN(
        n11749) );
  AOI21_X2 U7337 ( .B1(n12511), .B2(n11267), .A(n8165), .ZN(n11301) );
  AOI21_X2 U7338 ( .B1(n15171), .B2(n15170), .A(n15169), .ZN(n15380) );
  NOR2_X2 U7339 ( .A1(n15045), .A2(n15743), .ZN(n15046) );
  XNOR2_X1 U7340 ( .A(n9520), .B(n9521), .ZN(n10692) );
  NAND2_X2 U7341 ( .A1(n9561), .A2(n9567), .ZN(n13830) );
  XNOR2_X2 U7342 ( .A(n13807), .B(n11506), .ZN(n11463) );
  XNOR2_X1 U7344 ( .A(n8414), .B(P3_IR_REG_19__SCAN_IN), .ZN(n12461) );
  BUF_X4 U7345 ( .A(n10580), .Z(n6532) );
  XNOR2_X2 U7347 ( .A(n8543), .B(P3_IR_REG_22__SCAN_IN), .ZN(n12644) );
  XNOR2_X2 U7352 ( .A(n9028), .B(n9027), .ZN(n11877) );
  XNOR2_X1 U7354 ( .A(n15611), .B(n15610), .ZN(n15650) );
  NAND2_X2 U7355 ( .A1(n8913), .A2(n8912), .ZN(n14772) );
  OAI21_X2 U7356 ( .B1(n7155), .B2(n8738), .A(n7153), .ZN(n8751) );
  NAND2_X1 U7357 ( .A1(n8760), .A2(n8759), .ZN(n14729) );
  INV_X4 U7358 ( .A(n8139), .ZN(n8517) );
  AOI211_X2 U7359 ( .C1(n15798), .C2(n15274), .A(n15273), .B(n15272), .ZN(
        n15432) );
  NAND2_X2 U7360 ( .A1(n9217), .A2(n9220), .ZN(n10549) );
  OAI22_X2 U7361 ( .A1(n8413), .A2(n8412), .B1(P1_DATAO_REG_19__SCAN_IN), .B2(
        n11878), .ZN(n8428) );
  NAND2_X1 U7362 ( .A1(n15222), .A2(n15220), .ZN(n15221) );
  NAND3_X1 U7363 ( .A1(n7141), .A2(n10462), .A3(n6751), .ZN(n14562) );
  AND2_X1 U7364 ( .A1(n7204), .A2(n7203), .ZN(n12821) );
  NAND2_X1 U7365 ( .A1(n9990), .A2(n9989), .ZN(n14405) );
  NAND2_X1 U7366 ( .A1(n9068), .A2(n9067), .ZN(n15405) );
  XNOR2_X1 U7367 ( .A(n13881), .B(n12302), .ZN(n13880) );
  NAND2_X1 U7368 ( .A1(n9000), .A2(n8999), .ZN(n15438) );
  NAND2_X1 U7369 ( .A1(n14257), .A2(n10161), .ZN(n14241) );
  NAND2_X1 U7370 ( .A1(n8875), .A2(n8874), .ZN(n15480) );
  NAND2_X1 U7371 ( .A1(n7483), .A2(n9635), .ZN(n14264) );
  AND3_X1 U7372 ( .A1(n8727), .A2(n8726), .A3(n8725), .ZN(n11283) );
  INV_X1 U7374 ( .A(n14968), .ZN(n14481) );
  INV_X4 U7375 ( .A(n9947), .ZN(n10091) );
  NAND2_X1 U7378 ( .A1(n14709), .A2(n14699), .ZN(n9144) );
  INV_X4 U7379 ( .A(n14529), .ZN(n10287) );
  NAND4_X1 U7381 ( .A1(n8180), .A2(n8179), .A3(n8178), .A4(n8177), .ZN(n12954)
         );
  AND3_X1 U7382 ( .A1(n8186), .A2(n8185), .A3(n8184), .ZN(n11310) );
  XNOR2_X1 U7383 ( .A(n8538), .B(P3_IR_REG_21__SCAN_IN), .ZN(n12493) );
  AOI21_X1 U7384 ( .B1(n7154), .B2(n8739), .A(n6626), .ZN(n7153) );
  OAI22_X1 U7385 ( .A1(n15580), .A2(n15562), .B1(P1_ADDR_REG_4__SCAN_IN), .B2(
        n15563), .ZN(n7500) );
  INV_X1 U7386 ( .A(n11371), .ZN(n11497) );
  AND3_X1 U7387 ( .A1(n7357), .A2(n6701), .A3(n7795), .ZN(n7792) );
  CLKBUF_X2 U7388 ( .A(n8149), .Z(n8216) );
  NAND2_X1 U7389 ( .A1(n9192), .A2(n7342), .ZN(n15183) );
  NOR2_X1 U7391 ( .A1(n6738), .A2(n12638), .ZN(n12647) );
  NAND2_X1 U7392 ( .A1(n6765), .A2(n6522), .ZN(n6738) );
  NAND2_X1 U7393 ( .A1(n7160), .A2(n7159), .ZN(n12388) );
  OR2_X1 U7394 ( .A1(n12639), .A2(n12640), .ZN(n6765) );
  AOI21_X1 U7395 ( .B1(n13939), .B2(n15866), .A(n15850), .ZN(n7575) );
  NAND2_X1 U7396 ( .A1(n6591), .A2(n12383), .ZN(n13965) );
  OAI21_X1 U7397 ( .B1(n12374), .B2(n7484), .A(n12387), .ZN(n7161) );
  XNOR2_X1 U7398 ( .A(n6757), .B(n14099), .ZN(n13939) );
  NAND2_X1 U7399 ( .A1(n14602), .A2(n7919), .ZN(n14579) );
  NAND2_X1 U7400 ( .A1(n12377), .A2(n6595), .ZN(n12383) );
  CLKBUF_X1 U7401 ( .A(n15247), .Z(n7336) );
  OAI21_X1 U7402 ( .B1(n6907), .B2(n6906), .A(n7980), .ZN(n9919) );
  AOI21_X1 U7403 ( .B1(n15102), .B2(n15745), .A(n7581), .ZN(n7580) );
  AOI21_X1 U7404 ( .B1(n13108), .B2(n6558), .A(n6780), .ZN(n6779) );
  CLKBUF_X1 U7405 ( .A(n9166), .Z(n7284) );
  AOI21_X1 U7406 ( .B1(n6831), .B2(n6833), .A(n6830), .ZN(n6829) );
  OR2_X1 U7407 ( .A1(n15101), .A2(n15742), .ZN(n7581) );
  NOR2_X1 U7408 ( .A1(n14887), .A2(n14890), .ZN(n14913) );
  NAND2_X1 U7409 ( .A1(n6876), .A2(n6874), .ZN(n13976) );
  AND2_X1 U7410 ( .A1(n15159), .A2(n6688), .ZN(n15130) );
  AND2_X1 U7411 ( .A1(n7355), .A2(n6603), .ZN(n12385) );
  OAI21_X1 U7412 ( .B1(n7642), .B2(n7420), .A(n10248), .ZN(n6875) );
  AND2_X1 U7413 ( .A1(n12616), .A2(n12620), .ZN(n13153) );
  NAND2_X1 U7414 ( .A1(n15268), .A2(n7997), .ZN(n15259) );
  NAND2_X1 U7415 ( .A1(n12692), .A2(n12691), .ZN(n13739) );
  AND2_X1 U7416 ( .A1(n7007), .A2(n6676), .ZN(n14803) );
  NOR2_X1 U7417 ( .A1(n14521), .A2(n7890), .ZN(n7889) );
  NAND2_X1 U7418 ( .A1(n14845), .A2(n14844), .ZN(n15114) );
  CLKBUF_X1 U7419 ( .A(n13254), .Z(n13296) );
  NAND2_X2 U7420 ( .A1(n10479), .A2(n10478), .ZN(n15379) );
  NAND2_X1 U7421 ( .A1(n10055), .A2(n10054), .ZN(n14401) );
  NAND2_X1 U7422 ( .A1(n9940), .A2(n9939), .ZN(n13972) );
  AOI21_X1 U7423 ( .B1(n7798), .B2(n7800), .A(n7797), .ZN(n7796) );
  NAND2_X1 U7424 ( .A1(n9965), .A2(n7237), .ZN(n14854) );
  NAND2_X1 U7425 ( .A1(n8516), .A2(n8515), .ZN(n13358) );
  NAND2_X1 U7426 ( .A1(n14091), .A2(n7665), .ZN(n7664) );
  AND2_X1 U7427 ( .A1(n7065), .A2(n7696), .ZN(n7064) );
  CLKBUF_X1 U7428 ( .A(n14142), .Z(n6741) );
  NAND2_X1 U7429 ( .A1(n10006), .A2(n10005), .ZN(n13995) );
  CLKBUF_X1 U7430 ( .A(n14299), .Z(n7324) );
  XNOR2_X1 U7431 ( .A(n9988), .B(n9987), .ZN(n14460) );
  OAI21_X1 U7432 ( .B1(n14106), .B2(n10235), .A(n10234), .ZN(n14091) );
  XNOR2_X1 U7433 ( .A(n9951), .B(n9950), .ZN(n14456) );
  INV_X1 U7434 ( .A(n15262), .ZN(n6530) );
  AND2_X1 U7435 ( .A1(n8490), .A2(n8489), .ZN(n13440) );
  NOR2_X1 U7436 ( .A1(n15077), .A2(n6764), .ZN(n15087) );
  NAND2_X1 U7437 ( .A1(n9860), .A2(n9859), .ZN(n14320) );
  XNOR2_X1 U7438 ( .A(n10021), .B(n9923), .ZN(n14471) );
  NAND2_X2 U7439 ( .A1(n9033), .A2(n9032), .ZN(n15252) );
  INV_X1 U7440 ( .A(n15313), .ZN(n6531) );
  NAND2_X1 U7441 ( .A1(n9103), .A2(n9102), .ZN(n15194) );
  NAND2_X1 U7442 ( .A1(n9836), .A2(n9835), .ZN(n14097) );
  AND2_X1 U7443 ( .A1(n6805), .A2(n6804), .ZN(n14170) );
  NAND2_X1 U7444 ( .A1(n9847), .A2(n9846), .ZN(n14325) );
  NAND2_X1 U7445 ( .A1(n9052), .A2(n9051), .ZN(n15413) );
  NAND2_X1 U7446 ( .A1(n9876), .A2(n9875), .ZN(n14417) );
  XNOR2_X1 U7447 ( .A(n9066), .B(n9065), .ZN(n12050) );
  NAND2_X1 U7448 ( .A1(n15682), .A2(n7723), .ZN(n7722) );
  NAND2_X1 U7449 ( .A1(n9120), .A2(n9119), .ZN(n10022) );
  OAI21_X1 U7450 ( .B1(n15615), .B2(n7398), .A(n15679), .ZN(n7396) );
  XNOR2_X1 U7451 ( .A(n15325), .B(n15458), .ZN(n15324) );
  NAND2_X1 U7452 ( .A1(n9026), .A2(n9025), .ZN(n9028) );
  OAI21_X1 U7453 ( .B1(n13094), .B2(n13093), .A(n13092), .ZN(n13095) );
  OAI22_X1 U7454 ( .A1(n15741), .A2(P1_REG1_REG_15__SCAN_IN), .B1(n15743), 
        .B2(n15038), .ZN(n15039) );
  AND2_X1 U7455 ( .A1(n9189), .A2(n9188), .ZN(n14816) );
  NAND2_X2 U7456 ( .A1(n7603), .A2(n9765), .ZN(n14351) );
  XNOR2_X1 U7457 ( .A(n15037), .B(n7595), .ZN(n15741) );
  NAND2_X1 U7458 ( .A1(n8942), .A2(n8941), .ZN(n15325) );
  OAI21_X1 U7459 ( .B1(n7715), .B2(n7714), .A(n7713), .ZN(n7712) );
  NAND2_X1 U7460 ( .A1(n9734), .A2(n9733), .ZN(n14341) );
  NAND2_X1 U7461 ( .A1(n15035), .A2(n7596), .ZN(n15037) );
  XNOR2_X1 U7462 ( .A(n9050), .B(SI_18_), .ZN(n9024) );
  NAND2_X1 U7463 ( .A1(n7021), .A2(n7558), .ZN(n14748) );
  NAND2_X1 U7464 ( .A1(n9009), .A2(n9008), .ZN(n9050) );
  NAND2_X1 U7465 ( .A1(n14241), .A2(n14240), .ZN(n14239) );
  NAND2_X1 U7466 ( .A1(n9097), .A2(n9096), .ZN(n15383) );
  INV_X1 U7467 ( .A(n14368), .ZN(n14197) );
  NAND2_X1 U7468 ( .A1(n9718), .A2(n9717), .ZN(n14362) );
  OAI21_X1 U7469 ( .B1(n7729), .B2(n7728), .A(n6656), .ZN(n7727) );
  XNOR2_X1 U7470 ( .A(n8924), .B(n8959), .ZN(n11446) );
  OAI211_X1 U7471 ( .C1(n8907), .C2(n8906), .A(n8905), .B(n8904), .ZN(n8924)
         );
  NAND2_X1 U7472 ( .A1(n12003), .A2(n10214), .ZN(n12021) );
  NAND2_X1 U7473 ( .A1(n9687), .A2(n9686), .ZN(n14443) );
  NAND2_X1 U7474 ( .A1(n9672), .A2(n9671), .ZN(n14379) );
  NAND2_X1 U7475 ( .A1(n7442), .A2(n8834), .ZN(n15495) );
  NOR3_X1 U7476 ( .A1(n12978), .A2(n12977), .A3(n12976), .ZN(n13002) );
  NAND2_X1 U7477 ( .A1(n11576), .A2(n11575), .ZN(n11595) );
  NAND2_X1 U7478 ( .A1(n11241), .A2(n11240), .ZN(n11477) );
  OR2_X1 U7479 ( .A1(n10883), .A2(n10882), .ZN(n11179) );
  NAND2_X1 U7480 ( .A1(n9651), .A2(n9650), .ZN(n14386) );
  AOI22_X1 U7481 ( .A1(n11238), .A2(n11237), .B1(n11236), .B2(n12258), .ZN(
        n11241) );
  NAND2_X1 U7482 ( .A1(n13608), .A2(n13607), .ZN(n13606) );
  AND2_X1 U7483 ( .A1(n6689), .A2(n6892), .ZN(n7655) );
  AND3_X1 U7484 ( .A1(n11417), .A2(n7323), .A3(n6678), .ZN(n13608) );
  AND2_X1 U7485 ( .A1(n7582), .A2(n6684), .ZN(n15022) );
  NAND2_X1 U7486 ( .A1(n15603), .A2(n15602), .ZN(n15605) );
  INV_X1 U7487 ( .A(n11283), .ZN(n7945) );
  NAND2_X1 U7488 ( .A1(n10801), .A2(n10735), .ZN(n12931) );
  NAND2_X1 U7489 ( .A1(n9572), .A2(n9571), .ZN(n11930) );
  NAND2_X1 U7490 ( .A1(n6835), .A2(n14705), .ZN(n11637) );
  BUF_X1 U7491 ( .A(n15700), .Z(n6534) );
  OAI21_X1 U7492 ( .B1(n14699), .B2(n14709), .A(n9144), .ZN(n14923) );
  INV_X1 U7493 ( .A(n14695), .ZN(n10309) );
  NAND2_X1 U7494 ( .A1(n8544), .A2(n10706), .ZN(n13336) );
  NAND2_X1 U7495 ( .A1(n12518), .A2(n8590), .ZN(n12511) );
  AND2_X1 U7496 ( .A1(n10279), .A2(n7130), .ZN(n10296) );
  AND4_X2 U7497 ( .A1(n8690), .A2(n8689), .A3(n8688), .A4(n8687), .ZN(n14709)
         );
  NAND4_X1 U7498 ( .A1(n9580), .A2(n9579), .A3(n9578), .A4(n9577), .ZN(n13806)
         );
  INV_X2 U7499 ( .A(n10290), .ZN(n14531) );
  AND3_X2 U7500 ( .A1(n6605), .A2(n7082), .A3(n7081), .ZN(n14699) );
  AND4_X2 U7501 ( .A1(n8695), .A2(n8696), .A3(n7538), .A4(n7537), .ZN(n14695)
         );
  CLKBUF_X1 U7502 ( .A(n10782), .Z(n10707) );
  NAND4_X2 U7503 ( .A1(n9527), .A2(n9526), .A3(n9525), .A4(n9524), .ZN(n13809)
         );
  NAND2_X1 U7504 ( .A1(n8224), .A2(n8223), .ZN(n11974) );
  NAND4_X1 U7505 ( .A1(n8190), .A2(n8189), .A3(n8188), .A4(n8187), .ZN(n10796)
         );
  NAND4_X1 U7506 ( .A1(n8157), .A2(n8156), .A3(n8155), .A4(n8154), .ZN(n12952)
         );
  AOI21_X1 U7507 ( .B1(n12493), .B2(n11753), .A(n12632), .ZN(n10781) );
  NAND2_X1 U7508 ( .A1(n10252), .A2(n10251), .ZN(n14270) );
  NAND4_X2 U7509 ( .A1(n8144), .A2(n8143), .A3(n8142), .A4(n8141), .ZN(n12344)
         );
  NAND4_X1 U7510 ( .A1(n8236), .A2(n8235), .A3(n8234), .A4(n8233), .ZN(n12949)
         );
  INV_X1 U7511 ( .A(n7500), .ZN(n15565) );
  BUF_X2 U7512 ( .A(n8198), .Z(n8521) );
  BUF_X2 U7513 ( .A(n8197), .Z(n12398) );
  XNOR2_X1 U7515 ( .A(n8541), .B(n7332), .ZN(n11753) );
  NAND2_X1 U7516 ( .A1(n9210), .A2(n9214), .ZN(n15550) );
  NAND2_X1 U7517 ( .A1(n9131), .A2(n9204), .ZN(n11962) );
  NAND2_X4 U7518 ( .A1(n10102), .A2(n14462), .ZN(n10552) );
  NAND2_X1 U7519 ( .A1(n9497), .A2(n9498), .ZN(n11964) );
  NAND2_X1 U7520 ( .A1(n7791), .A2(n7790), .ZN(n14462) );
  XNOR2_X1 U7521 ( .A(n8059), .B(n7782), .ZN(n13510) );
  NAND2_X1 U7522 ( .A1(n8151), .A2(n8150), .ZN(n10976) );
  XNOR2_X1 U7523 ( .A(n8774), .B(SI_6_), .ZN(n8772) );
  OR2_X1 U7524 ( .A1(n9130), .A2(n8645), .ZN(n9128) );
  XNOR2_X1 U7525 ( .A(n7090), .B(n8661), .ZN(n9190) );
  XNOR2_X1 U7526 ( .A(n8130), .B(n8129), .ZN(n13515) );
  NAND2_X1 U7527 ( .A1(n8553), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8414) );
  INV_X4 U7528 ( .A(n6533), .ZN(n10579) );
  NAND2_X1 U7529 ( .A1(n7091), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7090) );
  OR2_X1 U7530 ( .A1(n7792), .A2(n7958), .ZN(n7957) );
  NAND2_X1 U7532 ( .A1(n7373), .A2(n7371), .ZN(n15583) );
  INV_X1 U7533 ( .A(n9207), .ZN(n8642) );
  AND3_X1 U7534 ( .A1(n8371), .A2(n8149), .A3(n8051), .ZN(n7089) );
  AND2_X1 U7536 ( .A1(n10097), .A2(n9478), .ZN(n7794) );
  AND3_X1 U7537 ( .A1(n8047), .A2(n8046), .A3(n8206), .ZN(n8149) );
  AND2_X1 U7538 ( .A1(n15717), .A2(n7599), .ZN(n8673) );
  AND3_X1 U7539 ( .A1(n9474), .A2(n9473), .A3(n9475), .ZN(n6785) );
  NAND2_X1 U7541 ( .A1(n15919), .A2(n6783), .ZN(n10902) );
  AND2_X1 U7542 ( .A1(n9477), .A2(n9476), .ZN(n9500) );
  AND3_X1 U7543 ( .A1(n8049), .A2(n8050), .A3(n8048), .ZN(n8371) );
  AND2_X1 U7544 ( .A1(n8795), .A2(n8638), .ZN(n7557) );
  INV_X4 U7545 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  INV_X1 U7546 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n9201) );
  INV_X1 U7548 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n8830) );
  INV_X1 U7549 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n10097) );
  INV_X1 U7550 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n7057) );
  INV_X4 U7551 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3088) );
  INV_X1 U7552 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n8795) );
  NOR2_X2 U7553 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_2__SCAN_IN), .ZN(
        n7940) );
  INV_X1 U7554 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n8661) );
  NOR2_X1 U7555 ( .A1(P2_IR_REG_18__SCAN_IN), .A2(P2_IR_REG_17__SCAN_IN), .ZN(
        n7977) );
  INV_X1 U7556 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n9559) );
  NOR2_X1 U7557 ( .A1(P2_IR_REG_22__SCAN_IN), .A2(P2_IR_REG_21__SCAN_IN), .ZN(
        n7976) );
  NOR2_X1 U7558 ( .A1(P2_IR_REG_20__SCAN_IN), .A2(P2_IR_REG_19__SCAN_IN), .ZN(
        n7975) );
  INV_X4 U7559 ( .A(P3_STATE_REG_SCAN_IN), .ZN(P3_U3151) );
  NAND2_X1 U7560 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_28__SCAN_IN), 
        .ZN(n7958) );
  INV_X1 U7561 ( .A(P3_IR_REG_1__SCAN_IN), .ZN(n6783) );
  OAI21_X2 U7562 ( .B1(n11538), .B2(n7776), .A(n7775), .ZN(n11949) );
  NAND3_X1 U7563 ( .A1(n7527), .A2(n6949), .A3(n7795), .ZN(n9498) );
  INV_X2 U7564 ( .A(n15783), .ZN(n11166) );
  NOR2_X2 U7565 ( .A1(n11646), .A2(n6534), .ZN(n11512) );
  NOR2_X2 U7566 ( .A1(n11565), .A2(n15890), .ZN(n11564) );
  INV_X2 U7567 ( .A(n10053), .ZN(n9834) );
  NAND2_X1 U7568 ( .A1(n12728), .A2(n8038), .ZN(n12736) );
  NOR2_X2 U7569 ( .A1(n9053), .A2(n14626), .ZN(n7319) );
  NAND2_X4 U7570 ( .A1(n14851), .A2(n10549), .ZN(n10295) );
  BUF_X4 U7571 ( .A(n10580), .Z(n6533) );
  NAND2_X2 U7572 ( .A1(n7460), .A2(n7459), .ZN(n10580) );
  OAI211_X1 U7573 ( .C1(n8697), .C2(n10590), .A(n8711), .B(n8710), .ZN(n15700)
         );
  NOR2_X2 U7574 ( .A1(n12133), .A2(n12132), .ZN(n15044) );
  NOR2_X2 U7575 ( .A1(n9090), .A2(n9428), .ZN(n6749) );
  NAND2_X1 U7576 ( .A1(n9089), .A2(n6532), .ZN(n6535) );
  NAND2_X1 U7577 ( .A1(n9089), .A2(n6532), .ZN(n6536) );
  NAND2_X1 U7578 ( .A1(n9089), .A2(n6533), .ZN(n8724) );
  AND2_X4 U7579 ( .A1(n12771), .A2(n14455), .ZN(n9552) );
  INV_X1 U7580 ( .A(n7339), .ZN(n7338) );
  OAI21_X1 U7581 ( .B1(n12616), .B2(n12626), .A(n12615), .ZN(n7339) );
  AOI21_X1 U7582 ( .B1(n7690), .B2(n7692), .A(n6634), .ZN(n7689) );
  OR2_X1 U7583 ( .A1(n7493), .A2(P3_REG1_REG_1__SCAN_IN), .ZN(n7086) );
  OR2_X1 U7584 ( .A1(n7490), .A2(P3_REG1_REG_1__SCAN_IN), .ZN(n7085) );
  NAND2_X1 U7585 ( .A1(n13275), .A2(n8424), .ZN(n8426) );
  NOR2_X1 U7586 ( .A1(P3_IR_REG_21__SCAN_IN), .A2(P3_IR_REG_20__SCAN_IN), .ZN(
        n8550) );
  NOR2_X1 U7587 ( .A1(P3_IR_REG_22__SCAN_IN), .A2(P3_IR_REG_23__SCAN_IN), .ZN(
        n8551) );
  NAND2_X1 U7588 ( .A1(n6647), .A2(n10075), .ZN(n7293) );
  AOI21_X1 U7589 ( .B1(n13976), .B2(n7933), .A(n10250), .ZN(n10253) );
  AOI21_X1 U7590 ( .B1(n7163), .B2(n7162), .A(n6710), .ZN(n7169) );
  NAND2_X1 U7591 ( .A1(n7168), .A2(n7167), .ZN(n7166) );
  AND2_X1 U7592 ( .A1(n9494), .A2(n9501), .ZN(n7262) );
  NOR2_X1 U7593 ( .A1(P2_IR_REG_18__SCAN_IN), .A2(P2_IR_REG_19__SCAN_IN), .ZN(
        n9494) );
  NAND2_X1 U7594 ( .A1(n10501), .A2(n10500), .ZN(n7917) );
  NAND2_X1 U7595 ( .A1(n9173), .A2(n9172), .ZN(n12728) );
  INV_X1 U7596 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n8637) );
  INV_X1 U7597 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n8638) );
  NAND2_X1 U7598 ( .A1(n7923), .A2(n9928), .ZN(n10004) );
  NAND2_X1 U7599 ( .A1(n10022), .A2(n9922), .ZN(n7923) );
  XNOR2_X1 U7600 ( .A(n8845), .B(SI_10_), .ZN(n8843) );
  NAND2_X1 U7601 ( .A1(n6740), .A2(n7351), .ZN(n7204) );
  AND2_X1 U7602 ( .A1(n8068), .A2(n8060), .ZN(n8198) );
  AOI21_X1 U7603 ( .B1(n6848), .B2(n6851), .A(n13193), .ZN(n6846) );
  XNOR2_X1 U7604 ( .A(n14295), .B(n13786), .ZN(n14013) );
  BUF_X1 U7605 ( .A(n10056), .Z(n10140) );
  OR2_X1 U7606 ( .A1(n15495), .A2(n12249), .ZN(n8842) );
  AOI21_X1 U7607 ( .B1(n9625), .B2(n9624), .A(n9623), .ZN(n9627) );
  INV_X1 U7608 ( .A(n13419), .ZN(n12460) );
  NAND2_X1 U7609 ( .A1(n11674), .A2(n12950), .ZN(n12528) );
  NAND2_X1 U7610 ( .A1(n12954), .A2(n11310), .ZN(n12495) );
  AND2_X1 U7611 ( .A1(n14815), .A2(n7542), .ZN(n7354) );
  AND2_X1 U7612 ( .A1(n15262), .A2(n7697), .ZN(n7696) );
  OR2_X1 U7613 ( .A1(n15271), .A2(n7698), .ZN(n7697) );
  INV_X1 U7614 ( .A(n9934), .ZN(n7922) );
  NAND2_X1 U7615 ( .A1(n7274), .A2(n12626), .ZN(n7273) );
  OR2_X1 U7616 ( .A1(n12460), .A2(n13144), .ZN(n12630) );
  INV_X1 U7617 ( .A(n13510), .ZN(n8060) );
  INV_X1 U7618 ( .A(n10923), .ZN(n10922) );
  INV_X1 U7619 ( .A(n10931), .ZN(n7489) );
  NAND2_X1 U7620 ( .A1(n10946), .A2(n10945), .ZN(n10962) );
  OAI21_X1 U7621 ( .B1(n6894), .B2(n10970), .A(n6775), .ZN(n7401) );
  INV_X1 U7622 ( .A(n6776), .ZN(n6775) );
  OAI21_X1 U7623 ( .B1(n10971), .B2(n10970), .A(n6657), .ZN(n6776) );
  NAND2_X1 U7624 ( .A1(n12089), .A2(P3_REG2_REG_10__SCAN_IN), .ZN(n7650) );
  NAND2_X1 U7625 ( .A1(n11598), .A2(n7652), .ZN(n6770) );
  NAND2_X1 U7626 ( .A1(n11580), .A2(n6772), .ZN(n6771) );
  NAND2_X1 U7627 ( .A1(n12994), .A2(n13018), .ZN(n7399) );
  AOI21_X1 U7628 ( .B1(n13018), .B2(n12995), .A(n13026), .ZN(n7400) );
  OR2_X1 U7629 ( .A1(n12953), .A2(n11339), .ZN(n12504) );
  OR2_X1 U7630 ( .A1(n13451), .A2(n13246), .ZN(n12467) );
  AND2_X1 U7631 ( .A1(n7769), .A2(n6596), .ZN(n7766) );
  OR2_X1 U7632 ( .A1(n13381), .A2(n13247), .ZN(n12472) );
  OR2_X1 U7633 ( .A1(n13384), .A2(n13266), .ZN(n12587) );
  OR2_X1 U7634 ( .A1(n13469), .A2(n12869), .ZN(n13255) );
  NOR2_X1 U7635 ( .A1(n8102), .A2(n7855), .ZN(n7854) );
  INV_X1 U7636 ( .A(n8100), .ZN(n7855) );
  NOR2_X1 U7637 ( .A1(P3_IR_REG_14__SCAN_IN), .A2(P3_IR_REG_16__SCAN_IN), .ZN(
        n8049) );
  NOR2_X1 U7638 ( .A1(P3_IR_REG_15__SCAN_IN), .A2(P3_IR_REG_13__SCAN_IN), .ZN(
        n8050) );
  INV_X1 U7639 ( .A(P3_IR_REG_12__SCAN_IN), .ZN(n8048) );
  NAND2_X1 U7640 ( .A1(n6856), .A2(n6602), .ZN(n8088) );
  NOR2_X1 U7641 ( .A1(P3_IR_REG_9__SCAN_IN), .A2(P3_IR_REG_11__SCAN_IN), .ZN(
        n8044) );
  AND2_X1 U7642 ( .A1(n6692), .A2(n8085), .ZN(n7848) );
  NOR2_X1 U7643 ( .A1(n8243), .A2(n7835), .ZN(n7834) );
  NOR2_X1 U7644 ( .A1(P3_IR_REG_4__SCAN_IN), .A2(P3_IR_REG_1__SCAN_IN), .ZN(
        n8047) );
  NOR2_X1 U7645 ( .A1(P3_IR_REG_0__SCAN_IN), .A2(P3_IR_REG_3__SCAN_IN), .ZN(
        n8046) );
  NOR2_X1 U7646 ( .A1(n10079), .A2(n10019), .ZN(n10046) );
  NAND2_X1 U7647 ( .A1(n6761), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n10009) );
  NOR2_X1 U7648 ( .A1(n10029), .A2(n13659), .ZN(n6761) );
  INV_X1 U7649 ( .A(n10183), .ZN(n7809) );
  NAND2_X1 U7650 ( .A1(n9877), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n9908) );
  INV_X1 U7651 ( .A(n9878), .ZN(n9877) );
  INV_X1 U7652 ( .A(n10172), .ZN(n7481) );
  NAND2_X1 U7653 ( .A1(n10170), .A2(n7810), .ZN(n14142) );
  AND2_X1 U7654 ( .A1(n10169), .A2(n10171), .ZN(n7810) );
  INV_X1 U7655 ( .A(n14175), .ZN(n6884) );
  XNOR2_X1 U7656 ( .A(n14351), .B(n13670), .ZN(n10230) );
  INV_X1 U7657 ( .A(n7473), .ZN(n7471) );
  NAND2_X1 U7658 ( .A1(n11462), .A2(n11463), .ZN(n7802) );
  AND2_X1 U7659 ( .A1(n13808), .A2(n15890), .ZN(n10147) );
  NAND2_X1 U7660 ( .A1(n7434), .A2(n7433), .ZN(n12003) );
  NOR2_X1 U7661 ( .A1(n12000), .A2(n7432), .ZN(n7433) );
  INV_X1 U7662 ( .A(n10212), .ZN(n7432) );
  NAND2_X1 U7663 ( .A1(n6919), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6918) );
  NAND2_X1 U7664 ( .A1(n6921), .A2(n6920), .ZN(n6919) );
  NOR2_X1 U7665 ( .A1(P2_IR_REG_14__SCAN_IN), .A2(P2_IR_REG_13__SCAN_IN), .ZN(
        n9476) );
  NOR2_X1 U7666 ( .A1(P2_IR_REG_16__SCAN_IN), .A2(P2_IR_REG_15__SCAN_IN), .ZN(
        n9477) );
  NOR2_X1 U7667 ( .A1(P2_IR_REG_6__SCAN_IN), .A2(P2_IR_REG_10__SCAN_IN), .ZN(
        n9474) );
  NOR2_X1 U7668 ( .A1(P2_IR_REG_9__SCAN_IN), .A2(P2_IR_REG_11__SCAN_IN), .ZN(
        n9473) );
  NOR2_X1 U7669 ( .A1(P2_IR_REG_8__SCAN_IN), .A2(P2_IR_REG_7__SCAN_IN), .ZN(
        n9475) );
  NOR2_X1 U7670 ( .A1(P2_IR_REG_2__SCAN_IN), .A2(P2_IR_REG_3__SCAN_IN), .ZN(
        n6909) );
  NOR2_X1 U7671 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n6908) );
  AOI21_X1 U7672 ( .B1(n10309), .B2(n14526), .A(n10313), .ZN(n10315) );
  AND2_X1 U7673 ( .A1(n7905), .A2(n10466), .ZN(n7904) );
  NAND2_X1 U7674 ( .A1(n7320), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n10531) );
  AOI21_X1 U7675 ( .B1(n7689), .B2(n7067), .A(n6628), .ZN(n7066) );
  INV_X1 U7676 ( .A(n7690), .ZN(n7067) );
  NOR2_X1 U7677 ( .A1(n8010), .A2(n8009), .ZN(n8008) );
  INV_X1 U7678 ( .A(n14766), .ZN(n8009) );
  OR2_X1 U7679 ( .A1(n15480), .A2(n15466), .ZN(n14766) );
  NAND2_X1 U7680 ( .A1(n14481), .A2(n14729), .ZN(n8771) );
  NOR2_X1 U7681 ( .A1(n8015), .A2(n11850), .ZN(n8012) );
  INV_X1 U7682 ( .A(n8785), .ZN(n8015) );
  NAND2_X1 U7683 ( .A1(n10048), .A2(n9957), .ZN(n9964) );
  AND2_X1 U7684 ( .A1(n10024), .A2(n7173), .ZN(n7164) );
  XNOR2_X1 U7685 ( .A(n10022), .B(SI_24_), .ZN(n10021) );
  OR2_X1 U7686 ( .A1(n7924), .A2(n7186), .ZN(n7185) );
  NOR2_X1 U7687 ( .A1(n7928), .A2(n7186), .ZN(n7181) );
  AOI21_X1 U7688 ( .B1(n7606), .B2(n7607), .A(n6638), .ZN(n7604) );
  INV_X1 U7689 ( .A(n8829), .ZN(n7607) );
  AOI21_X1 U7690 ( .B1(n7446), .B2(n7448), .A(n6636), .ZN(n7443) );
  NAND2_X1 U7691 ( .A1(n6863), .A2(n8717), .ZN(n7155) );
  INV_X1 U7692 ( .A(n7030), .ZN(n15569) );
  OAI21_X1 U7693 ( .B1(n15609), .B2(P1_ADDR_REG_8__SCAN_IN), .A(n6585), .ZN(
        n7030) );
  AOI21_X1 U7694 ( .B1(n15629), .B2(n15630), .A(n7507), .ZN(n7506) );
  NOR2_X1 U7695 ( .A1(n15631), .A2(P1_ADDR_REG_16__SCAN_IN), .ZN(n7507) );
  XNOR2_X1 U7696 ( .A(n12829), .B(n13181), .ZN(n12831) );
  INV_X1 U7697 ( .A(n12823), .ZN(n7203) );
  NAND2_X1 U7698 ( .A1(n8066), .A2(n8065), .ZN(n8633) );
  NOR2_X1 U7699 ( .A1(n12904), .A2(n12905), .ZN(n12903) );
  NOR2_X1 U7700 ( .A1(n7641), .A2(n10961), .ZN(n7640) );
  INV_X1 U7701 ( .A(n10939), .ZN(n7641) );
  NOR2_X1 U7702 ( .A1(n7648), .A2(n7405), .ZN(n7404) );
  INV_X1 U7703 ( .A(P3_REG2_REG_11__SCAN_IN), .ZN(n7405) );
  OR2_X1 U7704 ( .A1(n13000), .A2(n13001), .ZN(n7496) );
  OAI22_X1 U7705 ( .A1(n13192), .A2(n7866), .B1(n7867), .B2(n8510), .ZN(n13168) );
  NAND2_X1 U7706 ( .A1(n8509), .A2(n8497), .ZN(n7866) );
  INV_X1 U7707 ( .A(n7868), .ZN(n7867) );
  OR2_X1 U7708 ( .A1(n12920), .A2(n13196), .ZN(n8609) );
  NAND2_X1 U7709 ( .A1(n6986), .A2(n6985), .ZN(n13275) );
  AOI21_X1 U7710 ( .B1(n6988), .B2(n6990), .A(n6709), .ZN(n6985) );
  AND4_X1 U7711 ( .A1(n8324), .A2(n8323), .A3(n8322), .A4(n8321), .ZN(n12216)
         );
  AOI21_X1 U7712 ( .B1(n7777), .B2(n7779), .A(n12565), .ZN(n7775) );
  INV_X1 U7713 ( .A(n7777), .ZN(n7776) );
  INV_X1 U7714 ( .A(n12636), .ZN(n10731) );
  INV_X1 U7715 ( .A(n7772), .ZN(n7771) );
  INV_X1 U7716 ( .A(n13153), .ZN(n13150) );
  NAND2_X1 U7717 ( .A1(n8384), .A2(n6992), .ZN(n6987) );
  OR2_X1 U7718 ( .A1(n13477), .A2(n13313), .ZN(n13286) );
  INV_X1 U7719 ( .A(n6981), .ZN(n6980) );
  AOI21_X1 U7720 ( .B1(n6981), .B2(n6979), .A(n6561), .ZN(n6978) );
  NOR2_X1 U7721 ( .A1(n6982), .A2(n8365), .ZN(n6981) );
  INV_X2 U7722 ( .A(n8488), .ZN(n12422) );
  INV_X1 U7723 ( .A(n8312), .ZN(n8052) );
  AND4_X1 U7724 ( .A1(n8054), .A2(n7857), .A3(n7329), .A4(n8053), .ZN(n8055)
         );
  INV_X1 U7725 ( .A(P3_IR_REG_26__SCAN_IN), .ZN(n8053) );
  AND2_X1 U7726 ( .A1(n7270), .A2(n8371), .ZN(n7231) );
  AND2_X1 U7727 ( .A1(n7785), .A2(n8051), .ZN(n7270) );
  AND2_X1 U7728 ( .A1(n8129), .A2(n7494), .ZN(n7785) );
  NAND2_X1 U7729 ( .A1(n8485), .A2(n8118), .ZN(n8499) );
  NAND2_X1 U7730 ( .A1(n8095), .A2(n8094), .ZN(n8353) );
  AND2_X1 U7731 ( .A1(n10659), .A2(P1_DATAO_REG_8__SCAN_IN), .ZN(n8084) );
  INV_X1 U7732 ( .A(n8192), .ZN(n8181) );
  NOR2_X1 U7733 ( .A1(n7610), .A2(n6941), .ZN(n6940) );
  INV_X1 U7734 ( .A(n13705), .ZN(n6941) );
  NAND2_X1 U7735 ( .A1(n6943), .A2(n6942), .ZN(n13586) );
  AOI21_X1 U7736 ( .B1(n6944), .B2(n6946), .A(n6565), .ZN(n6942) );
  INV_X1 U7737 ( .A(n9552), .ZN(n10035) );
  AND2_X1 U7738 ( .A1(n9482), .A2(n9483), .ZN(n9599) );
  NOR2_X1 U7739 ( .A1(n15859), .A2(n6951), .ZN(n13938) );
  OR2_X1 U7740 ( .A1(n14405), .A2(n13784), .ZN(n10129) );
  NOR2_X1 U7741 ( .A1(n14018), .A2(n7807), .ZN(n7806) );
  INV_X1 U7742 ( .A(n10185), .ZN(n7807) );
  INV_X1 U7743 ( .A(n14005), .ZN(n7355) );
  NAND2_X1 U7744 ( .A1(n14047), .A2(n10182), .ZN(n10184) );
  NAND2_X1 U7745 ( .A1(n6659), .A2(n10218), .ZN(n7439) );
  NOR2_X1 U7746 ( .A1(n10160), .A2(n6879), .ZN(n6878) );
  INV_X1 U7747 ( .A(n10217), .ZN(n6879) );
  AND2_X1 U7748 ( .A1(n10160), .A2(n10158), .ZN(n7461) );
  NAND2_X1 U7749 ( .A1(n10552), .A2(n6533), .ZN(n9557) );
  NOR2_X1 U7750 ( .A1(n13971), .A2(n6869), .ZN(n6868) );
  INV_X1 U7751 ( .A(n13622), .ZN(n6869) );
  NAND2_X1 U7752 ( .A1(n7240), .A2(n6865), .ZN(n6870) );
  INV_X1 U7753 ( .A(n10254), .ZN(n6865) );
  INV_X1 U7754 ( .A(n10552), .ZN(n9833) );
  NAND2_X1 U7755 ( .A1(n10552), .A2(n10579), .ZN(n9562) );
  AND2_X1 U7756 ( .A1(n11126), .A2(n11014), .ZN(n14387) );
  AND2_X1 U7757 ( .A1(n12056), .A2(n12052), .ZN(n11126) );
  XNOR2_X1 U7758 ( .A(n9480), .B(n9479), .ZN(n9482) );
  INV_X1 U7759 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n9479) );
  OR2_X1 U7760 ( .A1(n14449), .A2(n14451), .ZN(n9480) );
  XNOR2_X1 U7761 ( .A(n9481), .B(P2_IR_REG_29__SCAN_IN), .ZN(n9483) );
  OAI21_X1 U7762 ( .B1(n9493), .B2(n7989), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n9481) );
  OR2_X1 U7763 ( .A1(n6671), .A2(n7916), .ZN(n7912) );
  INV_X1 U7764 ( .A(n7917), .ZN(n7916) );
  NAND2_X1 U7765 ( .A1(n8654), .A2(n8650), .ZN(n8692) );
  OR2_X1 U7766 ( .A1(n11379), .A2(n11210), .ZN(n10525) );
  OR2_X1 U7767 ( .A1(n10522), .A2(P1_U3086), .ZN(n10526) );
  AND2_X1 U7768 ( .A1(n9193), .A2(n15552), .ZN(n10631) );
  NOR2_X1 U7769 ( .A1(n12135), .A2(n7597), .ZN(n12137) );
  AND2_X1 U7770 ( .A1(n12136), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n7597) );
  NAND2_X1 U7771 ( .A1(n12137), .A2(n12138), .ZN(n15035) );
  AND2_X1 U7772 ( .A1(n8996), .A2(n8995), .ZN(n7879) );
  NAND2_X1 U7773 ( .A1(n15153), .A2(n7709), .ZN(n15128) );
  NOR2_X1 U7774 ( .A1(n12715), .A2(n12714), .ZN(n12716) );
  NOR2_X1 U7775 ( .A1(n7127), .A2(n14963), .ZN(n12715) );
  XNOR2_X1 U7776 ( .A(n15350), .B(n14961), .ZN(n15144) );
  NAND2_X1 U7777 ( .A1(n15199), .A2(n9176), .ZN(n15167) );
  NAND2_X1 U7778 ( .A1(n7236), .A2(n7702), .ZN(n15216) );
  AOI21_X1 U7779 ( .B1(n7704), .B2(n7703), .A(n6630), .ZN(n7702) );
  NAND2_X1 U7780 ( .A1(n15235), .A2(n9061), .ZN(n15220) );
  NAND2_X1 U7781 ( .A1(n15259), .A2(n7449), .ZN(n15235) );
  NOR2_X1 U7782 ( .A1(n14945), .A2(n7450), .ZN(n7449) );
  INV_X1 U7783 ( .A(n9042), .ZN(n7450) );
  NAND2_X1 U7784 ( .A1(n11877), .A2(n8743), .ZN(n9033) );
  OAI21_X1 U7785 ( .B1(n15307), .B2(n8003), .A(n8000), .ZN(n15270) );
  AOI21_X1 U7786 ( .B1(n8002), .B2(n8004), .A(n8001), .ZN(n8000) );
  INV_X1 U7787 ( .A(n14780), .ZN(n8001) );
  INV_X1 U7788 ( .A(n14835), .ZN(n10536) );
  NAND2_X1 U7789 ( .A1(n8984), .A2(n8986), .ZN(n15308) );
  OR2_X1 U7790 ( .A1(n15471), .A2(n14572), .ZN(n14768) );
  NAND2_X1 U7791 ( .A1(n14932), .A2(n8842), .ZN(n7998) );
  NAND2_X1 U7792 ( .A1(n12112), .A2(n8842), .ZN(n6844) );
  INV_X1 U7793 ( .A(n9089), .ZN(n10629) );
  NAND2_X1 U7794 ( .A1(n15447), .A2(n15103), .ZN(n11381) );
  NAND2_X1 U7795 ( .A1(n10487), .A2(n10486), .ZN(n15373) );
  INV_X1 U7796 ( .A(n15801), .ZN(n15467) );
  AND2_X1 U7797 ( .A1(n10631), .A2(n15533), .ZN(n15801) );
  OR2_X1 U7798 ( .A1(n8697), .A2(n10592), .ZN(n7082) );
  OR2_X1 U7799 ( .A1(n6536), .A2(n10575), .ZN(n7081) );
  XNOR2_X1 U7800 ( .A(n8937), .B(n8936), .ZN(n11495) );
  OR2_X1 U7801 ( .A1(n8931), .A2(SI_14_), .ZN(n8932) );
  NAND2_X1 U7802 ( .A1(n7453), .A2(n7191), .ZN(n7451) );
  XNOR2_X1 U7803 ( .A(n15569), .B(n15570), .ZN(n15612) );
  AOI21_X1 U7804 ( .B1(n7258), .B2(n7257), .A(n6734), .ZN(n15626) );
  INV_X1 U7805 ( .A(n15621), .ZN(n7257) );
  INV_X1 U7806 ( .A(n15620), .ZN(n7258) );
  AOI21_X1 U7807 ( .B1(n12912), .B2(n12913), .A(n7748), .ZN(n7200) );
  NAND2_X1 U7808 ( .A1(n6973), .A2(n6971), .ZN(n13361) );
  INV_X1 U7809 ( .A(n6972), .ZN(n6971) );
  OR2_X1 U7810 ( .A1(n13179), .A2(n13245), .ZN(n6973) );
  OAI22_X1 U7811 ( .A1(n13181), .A2(n13267), .B1(n13265), .B2(n13180), .ZN(
        n6972) );
  NAND2_X1 U7812 ( .A1(n7317), .A2(n7316), .ZN(n7315) );
  NOR2_X1 U7813 ( .A1(n8549), .A2(n15970), .ZN(n7316) );
  NAND2_X1 U7814 ( .A1(n7862), .A2(n13336), .ZN(n7317) );
  NOR2_X1 U7815 ( .A1(n7932), .A2(n10135), .ZN(n10137) );
  AND2_X1 U7816 ( .A1(n10556), .A2(n12378), .ZN(n15866) );
  NAND2_X1 U7817 ( .A1(n7230), .A2(n13990), .ZN(n14288) );
  NAND2_X1 U7818 ( .A1(n6555), .A2(n14270), .ZN(n7230) );
  NAND2_X1 U7819 ( .A1(n7642), .A2(n7421), .ZN(n13989) );
  INV_X1 U7820 ( .A(n15183), .ZN(n9200) );
  NAND2_X1 U7821 ( .A1(n15615), .A2(n7398), .ZN(n7397) );
  INV_X1 U7822 ( .A(n7510), .ZN(n15619) );
  OR2_X1 U7823 ( .A1(n15687), .A2(P2_ADDR_REG_14__SCAN_IN), .ZN(n7718) );
  NAND2_X1 U7824 ( .A1(n7722), .A2(n7719), .ZN(n7717) );
  AOI21_X1 U7825 ( .B1(n15687), .B2(P2_ADDR_REG_14__SCAN_IN), .A(n7720), .ZN(
        n7719) );
  NAND2_X1 U7826 ( .A1(n10196), .A2(n11002), .ZN(n9507) );
  NOR2_X1 U7827 ( .A1(n8030), .A2(n6563), .ZN(n6912) );
  NAND2_X1 U7828 ( .A1(n9595), .A2(n9596), .ZN(n6913) );
  OR2_X1 U7829 ( .A1(n14726), .A2(n14728), .ZN(n7562) );
  INV_X1 U7830 ( .A(n14726), .ZN(n7564) );
  INV_X1 U7831 ( .A(n14728), .ZN(n14727) );
  NAND2_X1 U7832 ( .A1(n7363), .A2(n12626), .ZN(n7362) );
  INV_X1 U7833 ( .A(n12583), .ZN(n7363) );
  INV_X1 U7834 ( .A(n9626), .ZN(n7532) );
  INV_X1 U7835 ( .A(n9627), .ZN(n7533) );
  NAND2_X1 U7836 ( .A1(n14734), .A2(n14736), .ZN(n7560) );
  NAND2_X1 U7837 ( .A1(n6543), .A2(n7016), .ZN(n14734) );
  AND2_X1 U7838 ( .A1(n6685), .A2(n7019), .ZN(n7018) );
  NAND2_X1 U7839 ( .A1(n14738), .A2(n14741), .ZN(n7019) );
  OAI22_X1 U7840 ( .A1(n9713), .A2(n9714), .B1(n9695), .B2(n9696), .ZN(n7983)
         );
  NAND2_X1 U7841 ( .A1(n9831), .A2(n7621), .ZN(n7620) );
  INV_X1 U7842 ( .A(n14775), .ZN(n7549) );
  MUX2_X1 U7843 ( .A(n15310), .B(n15453), .S(n14824), .Z(n14782) );
  NOR2_X1 U7844 ( .A1(n15289), .A2(n14774), .ZN(n14783) );
  AND2_X1 U7845 ( .A1(n13198), .A2(n12603), .ZN(n7367) );
  NAND2_X1 U7846 ( .A1(n7979), .A2(n9858), .ZN(n7602) );
  INV_X1 U7847 ( .A(n9857), .ZN(n7978) );
  NAND2_X1 U7848 ( .A1(n6925), .A2(n6923), .ZN(n7979) );
  OAI21_X1 U7849 ( .B1(n6926), .B2(n7616), .A(n7614), .ZN(n6925) );
  OAI21_X1 U7850 ( .B1(n6926), .B2(n7622), .A(n6924), .ZN(n6923) );
  NAND2_X1 U7851 ( .A1(n7617), .A2(n9845), .ZN(n7616) );
  MUX2_X1 U7852 ( .A(n15435), .B(n15280), .S(n14824), .Z(n14790) );
  NOR2_X1 U7853 ( .A1(n14796), .A2(n14795), .ZN(n14799) );
  NOR2_X1 U7854 ( .A1(n14792), .A2(n14791), .ZN(n14796) );
  NAND2_X1 U7855 ( .A1(n8898), .A2(SI_13_), .ZN(n8926) );
  INV_X1 U7856 ( .A(n10243), .ZN(n7428) );
  INV_X1 U7857 ( .A(n14477), .ZN(n7894) );
  NAND2_X1 U7858 ( .A1(n10397), .A2(n7885), .ZN(n7884) );
  INV_X1 U7859 ( .A(n14631), .ZN(n7885) );
  INV_X1 U7860 ( .A(n15106), .ZN(n7307) );
  INV_X1 U7861 ( .A(n9048), .ZN(n7929) );
  NOR2_X1 U7862 ( .A1(n9049), .A2(n7931), .ZN(n7930) );
  INV_X1 U7863 ( .A(n9008), .ZN(n7931) );
  INV_X1 U7864 ( .A(n9043), .ZN(n9045) );
  INV_X1 U7865 ( .A(n8903), .ZN(n8927) );
  NAND2_X1 U7866 ( .A1(n8846), .A2(n10633), .ZN(n8867) );
  OAI21_X1 U7867 ( .B1(n6532), .B2(n10589), .A(n8721), .ZN(n8741) );
  NAND2_X1 U7868 ( .A1(n10580), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n8721) );
  INV_X1 U7869 ( .A(n15599), .ZN(n7038) );
  INV_X1 U7870 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n7037) );
  NAND2_X1 U7871 ( .A1(n7504), .A2(P3_ADDR_REG_7__SCAN_IN), .ZN(n7503) );
  INV_X1 U7872 ( .A(n12926), .ZN(n7216) );
  NOR2_X1 U7873 ( .A1(n7751), .A2(n12854), .ZN(n7217) );
  AND2_X1 U7874 ( .A1(n12854), .A2(n7215), .ZN(n7214) );
  NAND2_X1 U7875 ( .A1(n7216), .A2(n7750), .ZN(n7215) );
  INV_X1 U7876 ( .A(n11069), .ZN(n6797) );
  NOR2_X1 U7877 ( .A1(n11040), .A2(n11192), .ZN(n11201) );
  AOI21_X1 U7878 ( .B1(n11194), .B2(n6789), .A(n6788), .ZN(n6787) );
  INV_X1 U7879 ( .A(n11571), .ZN(n6788) );
  NOR2_X1 U7880 ( .A1(n13039), .A2(n6813), .ZN(n6812) );
  INV_X1 U7881 ( .A(P3_REG1_REG_13__SCAN_IN), .ZN(n6813) );
  OR2_X1 U7882 ( .A1(n13358), .A2(n13181), .ZN(n12611) );
  NOR2_X1 U7883 ( .A1(n13185), .A2(n7101), .ZN(n7100) );
  INV_X1 U7884 ( .A(n12463), .ZN(n7101) );
  NAND2_X1 U7885 ( .A1(n6977), .A2(n6974), .ZN(n12532) );
  NAND2_X1 U7886 ( .A1(n12532), .A2(n12528), .ZN(n8594) );
  INV_X1 U7887 ( .A(P3_REG3_REG_6__SCAN_IN), .ZN(n7105) );
  INV_X1 U7888 ( .A(P3_REG3_REG_5__SCAN_IN), .ZN(n7107) );
  NAND2_X1 U7889 ( .A1(n12496), .A2(n12495), .ZN(n10784) );
  INV_X1 U7890 ( .A(n11753), .ZN(n10705) );
  INV_X1 U7891 ( .A(n12644), .ZN(n8618) );
  NOR2_X1 U7892 ( .A1(P3_IR_REG_27__SCAN_IN), .A2(P3_IR_REG_31__SCAN_IN), .ZN(
        n7491) );
  NAND2_X1 U7893 ( .A1(n8441), .A2(n8109), .ZN(n8111) );
  INV_X1 U7894 ( .A(n8540), .ZN(n8539) );
  INV_X1 U7895 ( .A(n7854), .ZN(n7851) );
  INV_X1 U7896 ( .A(n8104), .ZN(n7850) );
  OR2_X1 U7897 ( .A1(n8353), .A2(n8352), .ZN(n8098) );
  INV_X1 U7898 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n8868) );
  NAND2_X1 U7899 ( .A1(n10625), .A2(P2_DATAO_REG_6__SCAN_IN), .ZN(n8082) );
  INV_X1 U7900 ( .A(P3_IR_REG_2__SCAN_IN), .ZN(n8206) );
  INV_X1 U7901 ( .A(n13653), .ZN(n13550) );
  NOR2_X1 U7902 ( .A1(n13632), .A2(n6948), .ZN(n6947) );
  INV_X1 U7903 ( .A(n13538), .ZN(n6948) );
  INV_X1 U7904 ( .A(n10069), .ZN(n7292) );
  INV_X1 U7905 ( .A(n10070), .ZN(n7291) );
  OR2_X1 U7906 ( .A1(n10071), .A2(n10001), .ZN(n10079) );
  OR2_X1 U7907 ( .A1(n9901), .A2(n9902), .ZN(n7980) );
  NAND2_X1 U7908 ( .A1(n7525), .A2(n7981), .ZN(n6906) );
  AND2_X1 U7909 ( .A1(n7152), .A2(n13993), .ZN(n6877) );
  AND2_X1 U7910 ( .A1(n7645), .A2(n14013), .ZN(n7152) );
  AND4_X1 U7911 ( .A1(n7973), .A2(n14114), .A3(n6608), .A4(n10202), .ZN(n14025) );
  INV_X1 U7912 ( .A(n14417), .ZN(n7971) );
  NAND2_X1 U7913 ( .A1(n7480), .A2(n10173), .ZN(n7478) );
  INV_X1 U7914 ( .A(n7799), .ZN(n7798) );
  OAI21_X1 U7915 ( .B1(n14110), .B2(n7800), .A(n10176), .ZN(n7799) );
  NOR2_X1 U7916 ( .A1(n9821), .A2(n9820), .ZN(n6762) );
  NOR2_X1 U7917 ( .A1(n14379), .A2(n14386), .ZN(n7969) );
  INV_X1 U7918 ( .A(n14260), .ZN(n10199) );
  XNOR2_X1 U7919 ( .A(n14264), .B(n7482), .ZN(n10160) );
  NAND2_X1 U7921 ( .A1(n9498), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9495) );
  INV_X1 U7922 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n9501) );
  NOR2_X1 U7923 ( .A1(n7888), .A2(n7140), .ZN(n7139) );
  INV_X1 U7924 ( .A(n10433), .ZN(n7140) );
  INV_X1 U7925 ( .A(n7888), .ZN(n6753) );
  INV_X1 U7926 ( .A(n14663), .ZN(n6752) );
  INV_X1 U7927 ( .A(n14851), .ZN(n14706) );
  AND2_X1 U7928 ( .A1(n7883), .A2(n7143), .ZN(n7142) );
  NAND2_X1 U7929 ( .A1(n7144), .A2(n7146), .ZN(n7143) );
  AND2_X1 U7930 ( .A1(n7884), .A2(n14487), .ZN(n7883) );
  OR2_X1 U7931 ( .A1(n14819), .A2(n14821), .ZN(n7024) );
  NOR2_X1 U7932 ( .A1(n7354), .A2(n6637), .ZN(n7029) );
  OR2_X1 U7933 ( .A1(n14892), .A2(n14885), .ZN(n14887) );
  NAND2_X1 U7934 ( .A1(n7304), .A2(n6611), .ZN(n14886) );
  NOR2_X1 U7935 ( .A1(n7594), .A2(n11480), .ZN(n7590) );
  NAND2_X1 U7936 ( .A1(n6545), .A2(n6841), .ZN(n6840) );
  AND2_X1 U7937 ( .A1(n14951), .A2(n12732), .ZN(n15148) );
  NAND2_X1 U7938 ( .A1(n15280), .A2(n7123), .ZN(n7122) );
  INV_X1 U7939 ( .A(n15438), .ZN(n7123) );
  AND2_X1 U7940 ( .A1(n7951), .A2(n7950), .ZN(n7949) );
  NAND2_X1 U7941 ( .A1(n7693), .A2(n7694), .ZN(n15247) );
  AOI21_X1 U7942 ( .B1(n7696), .B2(n7698), .A(n6629), .ZN(n7694) );
  AND2_X1 U7943 ( .A1(n15236), .A2(n15421), .ZN(n7951) );
  INV_X1 U7944 ( .A(n7689), .ZN(n7068) );
  OR2_X1 U7945 ( .A1(n15438), .A2(n15311), .ZN(n14779) );
  OAI21_X1 U7946 ( .B1(n14939), .B2(n8010), .A(n8921), .ZN(n8006) );
  INV_X1 U7947 ( .A(n14698), .ZN(n6838) );
  AOI21_X1 U7948 ( .B1(n14926), .B2(n8728), .A(n6620), .ZN(n7999) );
  NAND2_X1 U7949 ( .A1(n14695), .A2(n6534), .ZN(n14698) );
  NAND2_X1 U7950 ( .A1(n11212), .A2(n9141), .ZN(n6835) );
  NAND2_X1 U7951 ( .A1(n14835), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n8688) );
  XNOR2_X1 U7952 ( .A(n14742), .B(n14513), .ZN(n14933) );
  AND2_X2 U7953 ( .A1(n9193), .A2(n11962), .ZN(n14851) );
  AND2_X1 U7954 ( .A1(n9224), .A2(n9223), .ZN(n9239) );
  AOI21_X1 U7955 ( .B1(n7180), .B2(n7177), .A(n6704), .ZN(n10048) );
  NOR3_X1 U7956 ( .A1(n7179), .A2(n9950), .A3(n7178), .ZN(n7177) );
  INV_X1 U7957 ( .A(n9952), .ZN(n7176) );
  AOI21_X1 U7958 ( .B1(n6571), .B2(n9921), .A(n7921), .ZN(n7920) );
  INV_X1 U7959 ( .A(n9933), .ZN(n7921) );
  NAND2_X1 U7960 ( .A1(n10023), .A2(n6571), .ZN(n7180) );
  INV_X1 U7961 ( .A(n10025), .ZN(n7168) );
  INV_X1 U7962 ( .A(n10024), .ZN(n7163) );
  NOR2_X1 U7963 ( .A1(n7308), .A2(n9207), .ZN(n9209) );
  NAND2_X1 U7964 ( .A1(n8989), .A2(n8988), .ZN(n9007) );
  NAND2_X1 U7965 ( .A1(n7193), .A2(n8790), .ZN(n8807) );
  INV_X1 U7966 ( .A(n15572), .ZN(n7041) );
  INV_X1 U7967 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n7045) );
  XNOR2_X1 U7968 ( .A(n7506), .B(n15637), .ZN(n15638) );
  AOI21_X1 U7969 ( .B1(n7217), .B2(n7216), .A(n12932), .ZN(n7212) );
  INV_X1 U7970 ( .A(n7217), .ZN(n7213) );
  NAND2_X1 U7971 ( .A1(n7211), .A2(n7210), .ZN(n7209) );
  INV_X1 U7972 ( .A(n7212), .ZN(n7211) );
  INV_X1 U7973 ( .A(n7214), .ZN(n7210) );
  NAND2_X1 U7974 ( .A1(n7214), .A2(n7751), .ZN(n7206) );
  OAI21_X1 U7975 ( .B1(n12435), .B2(n12434), .A(n12433), .ZN(n12640) );
  AND2_X1 U7976 ( .A1(n12432), .A2(n12431), .ZN(n12433) );
  AOI21_X1 U7977 ( .B1(n12631), .B2(n12630), .A(n12629), .ZN(n12637) );
  NAND2_X1 U7978 ( .A1(n7273), .A2(n7272), .ZN(n12631) );
  NAND2_X1 U7979 ( .A1(n12627), .A2(n12598), .ZN(n7272) );
  NOR2_X1 U7980 ( .A1(n12462), .A2(n7838), .ZN(n7837) );
  AND4_X1 U7981 ( .A1(n12403), .A2(n8537), .A3(n8536), .A4(n8535), .ZN(n13157)
         );
  AOI21_X1 U7982 ( .B1(n13293), .B2(n8466), .A(n8411), .ZN(n12869) );
  NAND2_X1 U7983 ( .A1(n8466), .A2(n11668), .ZN(n6976) );
  INV_X1 U7984 ( .A(n10921), .ZN(n12955) );
  NAND2_X1 U7985 ( .A1(n7060), .A2(n7058), .ZN(n11076) );
  INV_X1 U7986 ( .A(n7059), .ZN(n7058) );
  NAND2_X1 U7987 ( .A1(n7062), .A2(n12962), .ZN(n7060) );
  XNOR2_X1 U7988 ( .A(n10962), .B(n10947), .ZN(n10960) );
  NAND2_X1 U7989 ( .A1(n10963), .A2(n6803), .ZN(n6801) );
  NAND2_X1 U7990 ( .A1(n10960), .A2(P3_REG1_REG_3__SCAN_IN), .ZN(n6802) );
  NAND2_X1 U7991 ( .A1(n10940), .A2(n10939), .ZN(n6769) );
  OR2_X1 U7992 ( .A1(n10969), .A2(n10979), .ZN(n6895) );
  OAI21_X1 U7993 ( .B1(n11064), .B2(n7661), .A(n7659), .ZN(n10969) );
  NAND2_X1 U7994 ( .A1(n7657), .A2(n7656), .ZN(n10971) );
  NAND2_X1 U7995 ( .A1(n11064), .A2(n7659), .ZN(n7657) );
  AOI21_X1 U7996 ( .B1(n7659), .B2(n7661), .A(n11109), .ZN(n7656) );
  NAND2_X1 U7997 ( .A1(n6893), .A2(n10971), .ZN(n11099) );
  INV_X1 U7998 ( .A(n6894), .ZN(n6893) );
  NAND2_X1 U7999 ( .A1(n11048), .A2(n11047), .ZN(n6892) );
  INV_X1 U8000 ( .A(n7401), .ZN(n11048) );
  NAND2_X1 U8001 ( .A1(n11038), .A2(n11037), .ZN(n11193) );
  AND2_X1 U8002 ( .A1(n11041), .A2(n7078), .ZN(n7071) );
  INV_X1 U8003 ( .A(n11203), .ZN(n7073) );
  AOI21_X1 U8004 ( .B1(n11076), .B2(n11075), .A(n11074), .ZN(n11104) );
  OAI21_X1 U8005 ( .B1(n11585), .B2(n11584), .A(n11583), .ZN(n11611) );
  OAI21_X1 U8006 ( .B1(n11597), .B2(n6795), .A(n6793), .ZN(n12971) );
  INV_X1 U8007 ( .A(n6794), .ZN(n6793) );
  OAI21_X1 U8008 ( .B1(n11596), .B2(n6795), .A(n12087), .ZN(n6794) );
  OAI21_X1 U8009 ( .B1(n7404), .B2(n12983), .A(n12982), .ZN(n12992) );
  INV_X1 U8010 ( .A(n6898), .ZN(n6897) );
  OR2_X1 U8011 ( .A1(n12983), .A2(n7638), .ZN(n6896) );
  OR2_X1 U8012 ( .A1(n13030), .A2(n6715), .ZN(n7095) );
  NAND2_X1 U8013 ( .A1(n13055), .A2(n7684), .ZN(n7682) );
  AOI22_X1 U8014 ( .A1(n13086), .A2(n13085), .B1(P3_REG1_REG_16__SCAN_IN), 
        .B2(n13084), .ZN(n13102) );
  OR2_X1 U8015 ( .A1(n13095), .A2(n13096), .ZN(n7488) );
  NAND2_X1 U8016 ( .A1(n13169), .A2(n13340), .ZN(n7348) );
  INV_X1 U8017 ( .A(n13167), .ZN(n8610) );
  AND4_X1 U8018 ( .A1(n8508), .A2(n8507), .A3(n8506), .A4(n8505), .ZN(n13196)
         );
  NAND2_X1 U8019 ( .A1(n6994), .A2(n7000), .ZN(n7418) );
  AND2_X1 U8020 ( .A1(n7005), .A2(n7001), .ZN(n7000) );
  AOI21_X1 U8021 ( .B1(n6850), .B2(n13223), .A(n6849), .ZN(n6848) );
  INV_X1 U8022 ( .A(n12466), .ZN(n6849) );
  INV_X1 U8023 ( .A(n12441), .ZN(n8608) );
  NAND2_X1 U8024 ( .A1(n6544), .A2(n7003), .ZN(n6997) );
  NAND2_X1 U8025 ( .A1(n13243), .A2(n6999), .ZN(n6998) );
  NOR2_X1 U8026 ( .A1(n7004), .A2(n7002), .ZN(n6999) );
  NAND2_X1 U8027 ( .A1(n7761), .A2(n7759), .ZN(n13224) );
  AND2_X1 U8028 ( .A1(n7760), .A2(n12467), .ZN(n7759) );
  NAND2_X1 U8029 ( .A1(n8454), .A2(n12896), .ZN(n8475) );
  NAND2_X1 U8030 ( .A1(n6660), .A2(n12560), .ZN(n7777) );
  NAND2_X1 U8031 ( .A1(n6587), .A2(n8597), .ZN(n7780) );
  OR2_X1 U8032 ( .A1(n8232), .A2(P3_REG3_REG_8__SCAN_IN), .ZN(n8269) );
  NAND2_X1 U8033 ( .A1(n12423), .A2(n10615), .ZN(n7313) );
  INV_X1 U8034 ( .A(P3_REG3_REG_7__SCAN_IN), .ZN(n8230) );
  AND3_X1 U8035 ( .A1(n8248), .A2(n8247), .A3(n8246), .ZN(n11674) );
  NAND2_X1 U8036 ( .A1(n8211), .A2(n8210), .ZN(n12340) );
  NAND2_X1 U8037 ( .A1(n13182), .A2(n6582), .ZN(n13172) );
  AOI21_X1 U8038 ( .B1(n7766), .B2(n7764), .A(n7763), .ZN(n7762) );
  INV_X1 U8039 ( .A(n12471), .ZN(n7763) );
  INV_X1 U8040 ( .A(n8605), .ZN(n7764) );
  INV_X1 U8041 ( .A(n7766), .ZN(n7765) );
  AOI21_X1 U8042 ( .B1(n8605), .B2(n8606), .A(n7770), .ZN(n7769) );
  INV_X1 U8043 ( .A(n12472), .ZN(n7770) );
  AOI21_X1 U8044 ( .B1(n13281), .B2(n8466), .A(n8423), .ZN(n13266) );
  NAND2_X1 U8045 ( .A1(n8426), .A2(n6606), .ZN(n13264) );
  AND3_X1 U8046 ( .A1(n6862), .A2(n13258), .A3(n6861), .ZN(n8605) );
  OR2_X1 U8047 ( .A1(n8606), .A2(n13257), .ZN(n6862) );
  NAND2_X1 U8048 ( .A1(n8417), .A2(n8416), .ZN(n13384) );
  NAND2_X1 U8049 ( .A1(n13301), .A2(n8399), .ZN(n6991) );
  AOI21_X1 U8050 ( .B1(n6991), .B2(n6993), .A(n6989), .ZN(n6988) );
  INV_X1 U8051 ( .A(n6991), .ZN(n6990) );
  INV_X1 U8052 ( .A(n13312), .ZN(n8382) );
  NAND2_X1 U8053 ( .A1(n13318), .A2(n12480), .ZN(n13308) );
  AND2_X1 U8054 ( .A1(n12480), .A2(n12486), .ZN(n13325) );
  AOI21_X1 U8055 ( .B1(n7873), .B2(n7875), .A(n6631), .ZN(n7871) );
  INV_X1 U8056 ( .A(n8325), .ZN(n7875) );
  NAND2_X1 U8057 ( .A1(n8599), .A2(n12567), .ZN(n12217) );
  AND2_X1 U8058 ( .A1(n12479), .A2(n12484), .ZN(n12454) );
  INV_X1 U8059 ( .A(n13340), .ZN(n13267) );
  AOI21_X1 U8060 ( .B1(n11539), .B2(n8276), .A(n11787), .ZN(n7876) );
  OR2_X1 U8061 ( .A1(n11540), .A2(n11539), .ZN(n11542) );
  AND2_X1 U8062 ( .A1(n12561), .A2(n12560), .ZN(n11787) );
  NAND2_X1 U8063 ( .A1(n8596), .A2(n12545), .ZN(n11538) );
  AND2_X1 U8064 ( .A1(n12626), .A2(n10734), .ZN(n13340) );
  NAND2_X1 U8065 ( .A1(n7349), .A2(n13519), .ZN(n10621) );
  NAND2_X1 U8066 ( .A1(n7815), .A2(n7817), .ZN(n8127) );
  AOI21_X1 U8067 ( .B1(n8123), .B2(n7819), .A(n7818), .ZN(n7817) );
  NAND2_X1 U8068 ( .A1(n8499), .A2(n7816), .ZN(n7815) );
  INV_X1 U8069 ( .A(n8121), .ZN(n7819) );
  NAND2_X1 U8070 ( .A1(n8127), .A2(n8126), .ZN(n8529) );
  XNOR2_X1 U8071 ( .A(n7232), .B(P3_IR_REG_25__SCAN_IN), .ZN(n8579) );
  NAND2_X1 U8072 ( .A1(n8559), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7232) );
  NOR2_X1 U8073 ( .A1(n8552), .A2(P3_IR_REG_18__SCAN_IN), .ZN(n7218) );
  NAND2_X1 U8074 ( .A1(n8111), .A2(n8110), .ZN(n8451) );
  OR2_X1 U8075 ( .A1(n8542), .A2(P3_IR_REG_21__SCAN_IN), .ZN(n8576) );
  NAND2_X1 U8076 ( .A1(n8099), .A2(n6860), .ZN(n6859) );
  INV_X1 U8077 ( .A(n8097), .ZN(n6860) );
  NAND2_X1 U8078 ( .A1(n8098), .A2(n6541), .ZN(n6858) );
  NAND2_X1 U8079 ( .A1(n8367), .A2(n8099), .ZN(n8101) );
  AND2_X1 U8080 ( .A1(n8373), .A2(n8387), .ZN(n13088) );
  NAND2_X1 U8081 ( .A1(n7821), .A2(n7824), .ZN(n8340) );
  INV_X1 U8082 ( .A(n7825), .ZN(n7824) );
  OAI21_X1 U8083 ( .B1(n8089), .B2(n6581), .A(n8091), .ZN(n7825) );
  NAND2_X1 U8084 ( .A1(n8088), .A2(n8087), .ZN(n8311) );
  AOI21_X1 U8085 ( .B1(n7848), .B2(n6548), .A(n6654), .ZN(n7847) );
  NAND2_X1 U8086 ( .A1(n8264), .A2(n7848), .ZN(n6856) );
  OR2_X1 U8087 ( .A1(n8279), .A2(P3_IR_REG_9__SCAN_IN), .ZN(n8295) );
  AOI21_X1 U8088 ( .B1(n6588), .B2(n7830), .A(n7827), .ZN(n7826) );
  NOR2_X1 U8089 ( .A1(n10638), .A2(P2_DATAO_REG_7__SCAN_IN), .ZN(n7827) );
  XNOR2_X1 U8090 ( .A(n10636), .B(P1_DATAO_REG_7__SCAN_IN), .ZN(n8240) );
  INV_X1 U8091 ( .A(n7834), .ZN(n7833) );
  AOI21_X1 U8092 ( .B1(n7834), .B2(n7832), .A(n7831), .ZN(n7830) );
  INV_X1 U8093 ( .A(n8082), .ZN(n7831) );
  INV_X1 U8094 ( .A(n8171), .ZN(n7832) );
  XNOR2_X1 U8095 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(P2_DATAO_REG_5__SCAN_IN), 
        .ZN(n8171) );
  OAI21_X1 U8096 ( .B1(n8159), .B2(n8077), .A(n8076), .ZN(n8146) );
  NOR2_X1 U8097 ( .A1(n7633), .A2(n6936), .ZN(n6935) );
  INV_X1 U8098 ( .A(n11710), .ZN(n6936) );
  NOR2_X1 U8099 ( .A1(n7633), .A2(n11715), .ZN(n6933) );
  AND2_X1 U8100 ( .A1(n13580), .A2(n12671), .ZN(n12672) );
  INV_X1 U8101 ( .A(n6931), .ZN(n13565) );
  OAI21_X1 U8102 ( .B1(n7635), .B2(n6930), .A(n6928), .ZN(n6931) );
  INV_X1 U8103 ( .A(n6929), .ZN(n6928) );
  OAI21_X1 U8104 ( .B1(n13555), .B2(n6930), .A(n6644), .ZN(n6929) );
  OAI22_X1 U8105 ( .A1(n7628), .A2(n13598), .B1(n12655), .B2(n12656), .ZN(
        n7627) );
  NOR2_X1 U8106 ( .A1(n12681), .A2(n7612), .ZN(n7611) );
  INV_X1 U8107 ( .A(n12676), .ZN(n7612) );
  XNOR2_X1 U8108 ( .A(n14341), .B(n13615), .ZN(n12682) );
  AND2_X1 U8109 ( .A1(n13702), .A2(n6947), .ZN(n13630) );
  INV_X1 U8110 ( .A(n7627), .ZN(n7626) );
  OR2_X1 U8111 ( .A1(n13598), .A2(n7630), .ZN(n7629) );
  INV_X1 U8112 ( .A(n12651), .ZN(n7630) );
  NAND2_X1 U8113 ( .A1(n12184), .A2(n12183), .ZN(n12191) );
  NOR2_X1 U8114 ( .A1(n13670), .A2(n14261), .ZN(n13665) );
  XNOR2_X1 U8115 ( .A(n14351), .B(n13615), .ZN(n13664) );
  NAND2_X1 U8116 ( .A1(n10190), .A2(n7936), .ZN(n10142) );
  NOR2_X1 U8117 ( .A1(n10128), .A2(n7937), .ZN(n7936) );
  OR2_X1 U8118 ( .A1(n10230), .A2(n14180), .ZN(n7937) );
  NAND2_X1 U8119 ( .A1(n13816), .A2(n7568), .ZN(n10566) );
  OR2_X1 U8120 ( .A1(n10574), .A2(n10564), .ZN(n7568) );
  XNOR2_X1 U8121 ( .A(n6523), .B(P2_REG1_REG_2__SCAN_IN), .ZN(n10567) );
  NAND2_X1 U8122 ( .A1(n10691), .A2(n7566), .ZN(n15831) );
  NAND2_X1 U8123 ( .A1(n7567), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n7566) );
  INV_X1 U8124 ( .A(n6523), .ZN(n7567) );
  INV_X1 U8125 ( .A(n7565), .ZN(n6963) );
  NAND2_X1 U8126 ( .A1(n13904), .A2(n13903), .ZN(n13911) );
  INV_X1 U8127 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n13944) );
  NOR2_X1 U8128 ( .A1(n14401), .A2(n12384), .ZN(n7966) );
  NAND2_X1 U8129 ( .A1(n12385), .A2(n13962), .ZN(n12390) );
  AOI21_X2 U8130 ( .B1(n13968), .B2(n9550), .A(n9945), .ZN(n13614) );
  OR2_X1 U8131 ( .A1(n13972), .A2(n13614), .ZN(n12375) );
  OR2_X1 U8132 ( .A1(n9992), .A2(n9423), .ZN(n13959) );
  AND2_X1 U8133 ( .A1(n10009), .A2(n10008), .ZN(n13998) );
  AND2_X1 U8134 ( .A1(n7151), .A2(n6693), .ZN(n7642) );
  AOI21_X1 U8135 ( .B1(n7465), .B2(n7467), .A(n6627), .ZN(n7462) );
  INV_X1 U8136 ( .A(n6761), .ZN(n10031) );
  NAND2_X1 U8137 ( .A1(n10184), .A2(n6579), .ZN(n7808) );
  NAND2_X1 U8138 ( .A1(n14471), .A2(n7674), .ZN(n9904) );
  NAND2_X1 U8139 ( .A1(n7666), .A2(n10241), .ZN(n14057) );
  XNOR2_X1 U8140 ( .A(n14335), .B(n12686), .ZN(n14110) );
  NAND2_X1 U8141 ( .A1(n7477), .A2(n10173), .ZN(n14111) );
  NAND2_X1 U8142 ( .A1(n6741), .A2(n7479), .ZN(n7477) );
  NAND2_X1 U8143 ( .A1(n14111), .A2(n14110), .ZN(n14109) );
  NOR2_X1 U8144 ( .A1(n14351), .A2(n6882), .ZN(n6881) );
  NAND2_X1 U8145 ( .A1(n14156), .A2(n10230), .ZN(n10170) );
  AND2_X1 U8146 ( .A1(n6884), .A2(n6883), .ZN(n14163) );
  NOR2_X1 U8147 ( .A1(n14351), .A2(n14435), .ZN(n6883) );
  NAND2_X1 U8148 ( .A1(n6549), .A2(n6617), .ZN(n6808) );
  AND2_X1 U8149 ( .A1(n6609), .A2(n10226), .ZN(n12358) );
  AOI21_X1 U8150 ( .B1(n10164), .B2(n7474), .A(n6607), .ZN(n7473) );
  INV_X1 U8151 ( .A(n10163), .ZN(n7474) );
  INV_X1 U8152 ( .A(n10164), .ZN(n7475) );
  OR2_X1 U8153 ( .A1(n6619), .A2(n10165), .ZN(n14188) );
  AOI22_X1 U8154 ( .A1(n6658), .A2(n10222), .B1(n10221), .B2(n13801), .ZN(
        n10223) );
  NAND2_X1 U8155 ( .A1(n14239), .A2(n10162), .ZN(n14219) );
  INV_X1 U8156 ( .A(n10160), .ZN(n14271) );
  AND3_X1 U8157 ( .A1(n7960), .A2(n15901), .A3(n11564), .ZN(n12008) );
  XNOR2_X1 U8158 ( .A(n15901), .B(n13805), .ZN(n12000) );
  NAND2_X1 U8159 ( .A1(n11470), .A2(n11469), .ZN(n7437) );
  NAND2_X1 U8160 ( .A1(n7805), .A2(n7804), .ZN(n7803) );
  OR2_X1 U8161 ( .A1(n13809), .A2(n9522), .ZN(n11554) );
  NAND2_X1 U8162 ( .A1(n7677), .A2(n13815), .ZN(n7676) );
  INV_X1 U8163 ( .A(n10552), .ZN(n7677) );
  INV_X1 U8164 ( .A(n10578), .ZN(n7673) );
  INV_X1 U8165 ( .A(n14294), .ZN(n6821) );
  INV_X1 U8166 ( .A(n14396), .ZN(n14391) );
  NAND2_X1 U8167 ( .A1(n9492), .A2(n7959), .ZN(n7989) );
  AND2_X1 U8168 ( .A1(n7795), .A2(n7972), .ZN(n7440) );
  AND2_X1 U8169 ( .A1(n9500), .A2(n9501), .ZN(n6921) );
  XNOR2_X1 U8170 ( .A(n9670), .B(P2_IR_REG_10__SCAN_IN), .ZN(n11655) );
  OR2_X1 U8171 ( .A1(n9633), .A2(P2_IR_REG_8__SCAN_IN), .ZN(n9667) );
  NAND2_X1 U8172 ( .A1(n9569), .A2(n9568), .ZN(n9699) );
  AND2_X1 U8173 ( .A1(n14496), .A2(n7906), .ZN(n7902) );
  NAND2_X1 U8174 ( .A1(n7319), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n9090) );
  INV_X1 U8175 ( .A(n14570), .ZN(n7146) );
  AND2_X1 U8176 ( .A1(n10375), .A2(n14651), .ZN(n10376) );
  INV_X1 U8177 ( .A(n11962), .ZN(n14690) );
  AND4_X1 U8178 ( .A1(n8882), .A2(n8881), .A3(n8880), .A4(n8879), .ZN(n15466)
         );
  AND4_X1 U8179 ( .A1(n8841), .A2(n8840), .A3(n8839), .A4(n8838), .ZN(n12249)
         );
  AOI21_X1 U8180 ( .B1(n14976), .B2(P1_REG1_REG_1__SCAN_IN), .A(n14972), .ZN(
        n14984) );
  NOR2_X1 U8181 ( .A1(n14984), .A2(n14983), .ZN(n14982) );
  AOI21_X1 U8182 ( .B1(n14989), .B2(P1_REG1_REG_2__SCAN_IN), .A(n14982), .ZN(
        n10864) );
  NAND2_X1 U8183 ( .A1(n7241), .A2(n6623), .ZN(n7582) );
  NAND2_X1 U8184 ( .A1(n11984), .A2(n11980), .ZN(n7591) );
  NAND2_X1 U8185 ( .A1(n11477), .A2(n7590), .ZN(n7592) );
  NOR2_X1 U8186 ( .A1(n7588), .A2(n15730), .ZN(n7587) );
  NOR2_X1 U8187 ( .A1(n7590), .A2(n7589), .ZN(n7588) );
  INV_X1 U8188 ( .A(n7591), .ZN(n7589) );
  OR2_X1 U8189 ( .A1(n15036), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n7596) );
  NOR2_X1 U8190 ( .A1(n15061), .A2(n15060), .ZN(n15077) );
  INV_X1 U8191 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n15105) );
  NAND2_X1 U8192 ( .A1(n9197), .A2(n7124), .ZN(n15131) );
  AND2_X1 U8193 ( .A1(n6567), .A2(n7125), .ZN(n7124) );
  INV_X1 U8194 ( .A(n7707), .ZN(n7706) );
  NAND2_X1 U8195 ( .A1(n7311), .A2(n7709), .ZN(n7310) );
  OAI21_X1 U8196 ( .B1(n12735), .B2(n7708), .A(n15117), .ZN(n7707) );
  OR2_X1 U8197 ( .A1(n15160), .A2(n12754), .ZN(n10495) );
  NAND2_X1 U8198 ( .A1(n14467), .A2(n8743), .ZN(n10479) );
  NAND2_X1 U8199 ( .A1(n15205), .A2(n14805), .ZN(n15192) );
  XNOR2_X1 U8200 ( .A(n15214), .B(n15383), .ZN(n15217) );
  NAND2_X1 U8201 ( .A1(n15221), .A2(n6545), .ZN(n15205) );
  AND2_X1 U8202 ( .A1(n6530), .A2(n9023), .ZN(n7997) );
  OAI21_X1 U8203 ( .B1(n7284), .B2(n7068), .A(n7066), .ZN(n15266) );
  OAI21_X1 U8204 ( .B1(n9165), .B2(n7692), .A(n9167), .ZN(n7691) );
  INV_X1 U8205 ( .A(n15308), .ZN(n7692) );
  NOR2_X1 U8206 ( .A1(n15313), .A2(n15438), .ZN(n15278) );
  NAND2_X1 U8207 ( .A1(n14779), .A2(n14780), .ZN(n15289) );
  NAND2_X1 U8208 ( .A1(n8985), .A2(n7692), .ZN(n15305) );
  INV_X1 U8209 ( .A(n15307), .ZN(n8985) );
  XNOR2_X1 U8210 ( .A(n14772), .B(n15449), .ZN(n14941) );
  AND2_X2 U8211 ( .A1(n14768), .A2(n14771), .ZN(n14939) );
  NAND2_X1 U8212 ( .A1(n12263), .A2(n14766), .ZN(n12312) );
  NAND2_X1 U8213 ( .A1(n14939), .A2(n12312), .ZN(n12311) );
  INV_X1 U8214 ( .A(n15471), .ZN(n9195) );
  CLKBUF_X1 U8215 ( .A(n12313), .Z(n12314) );
  AOI21_X1 U8216 ( .B1(n8785), .B2(n8014), .A(n6616), .ZN(n8013) );
  INV_X1 U8217 ( .A(n8771), .ZN(n8014) );
  XNOR2_X1 U8218 ( .A(n14737), .B(n14618), .ZN(n14920) );
  AND2_X1 U8219 ( .A1(n8023), .A2(n9240), .ZN(n8022) );
  OR2_X1 U8220 ( .A1(n9199), .A2(n15820), .ZN(n8023) );
  INV_X1 U8221 ( .A(n15114), .ZN(n15348) );
  NAND2_X1 U8222 ( .A1(n6744), .A2(n15807), .ZN(n6743) );
  INV_X1 U8223 ( .A(n15382), .ZN(n6744) );
  AND2_X1 U8224 ( .A1(n9060), .A2(n9059), .ZN(n15401) );
  NAND2_X1 U8225 ( .A1(n12050), .A2(n8743), .ZN(n9068) );
  NAND2_X1 U8226 ( .A1(n8855), .A2(n8854), .ZN(n15490) );
  NOR2_X1 U8227 ( .A1(n10526), .A2(n9237), .ZN(n11211) );
  AND2_X1 U8228 ( .A1(n8025), .A2(n6826), .ZN(n6825) );
  NAND2_X1 U8229 ( .A1(n8644), .A2(n7092), .ZN(n7091) );
  AND2_X1 U8230 ( .A1(n8643), .A2(n8024), .ZN(n7092) );
  OR2_X1 U8231 ( .A1(n9209), .A2(n8645), .ZN(n7283) );
  AND2_X1 U8232 ( .A1(n7185), .A2(n9873), .ZN(n7183) );
  XNOR2_X1 U8233 ( .A(n9206), .B(n9205), .ZN(n10630) );
  OAI21_X1 U8234 ( .B1(n9204), .B2(n9203), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n9206) );
  OR2_X1 U8235 ( .A1(n7147), .A2(n8645), .ZN(n7017) );
  XNOR2_X1 U8236 ( .A(n9007), .B(n9006), .ZN(n11404) );
  XNOR2_X1 U8237 ( .A(n8884), .B(n8883), .ZN(n11247) );
  NAND2_X1 U8238 ( .A1(n8907), .A2(n8903), .ZN(n8884) );
  OAI21_X1 U8239 ( .B1(n8873), .B2(P1_IR_REG_11__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n8886) );
  NAND2_X1 U8240 ( .A1(n8907), .A2(n8872), .ZN(n11112) );
  OR2_X1 U8241 ( .A1(n8958), .A2(n8871), .ZN(n8872) );
  INV_X1 U8242 ( .A(n8756), .ZN(n8757) );
  OR2_X1 U8243 ( .A1(n8997), .A2(P1_IR_REG_5__SCAN_IN), .ZN(n8756) );
  NAND2_X1 U8244 ( .A1(n7445), .A2(n8754), .ZN(n7264) );
  INV_X1 U8245 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n7599) );
  NAND2_X1 U8246 ( .A1(P3_ADDR_REG_1__SCAN_IN), .A2(n7372), .ZN(n7371) );
  INV_X1 U8247 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n7372) );
  NAND2_X1 U8248 ( .A1(n15594), .A2(n15595), .ZN(n15598) );
  NAND2_X1 U8249 ( .A1(n15607), .A2(n15608), .ZN(n15611) );
  AOI21_X1 U8250 ( .B1(n7513), .B2(n7512), .A(n6726), .ZN(n15617) );
  INV_X1 U8251 ( .A(n15613), .ZN(n7512) );
  INV_X1 U8252 ( .A(n15678), .ZN(n7398) );
  OAI21_X1 U8253 ( .B1(n7510), .B2(n7033), .A(n7031), .ZN(n15620) );
  NAND2_X1 U8254 ( .A1(P3_ADDR_REG_13__SCAN_IN), .A2(n7032), .ZN(n7031) );
  INV_X1 U8255 ( .A(n15618), .ZN(n7033) );
  INV_X1 U8256 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n7032) );
  INV_X1 U8257 ( .A(n7721), .ZN(n7720) );
  NAND2_X1 U8258 ( .A1(n15627), .A2(n7508), .ZN(n15629) );
  NAND2_X1 U8259 ( .A1(P3_ADDR_REG_15__SCAN_IN), .A2(n7509), .ZN(n7508) );
  INV_X1 U8260 ( .A(n12831), .ZN(n7199) );
  NAND2_X1 U8261 ( .A1(n8474), .A2(n8473), .ZN(n13225) );
  NAND2_X1 U8262 ( .A1(n6739), .A2(n11088), .ZN(n11219) );
  AND2_X1 U8263 ( .A1(n8438), .A2(n8437), .ZN(n13247) );
  AND2_X1 U8264 ( .A1(n7738), .A2(n6697), .ZN(n7736) );
  AND2_X1 U8265 ( .A1(n7739), .A2(n12924), .ZN(n7738) );
  OAI21_X1 U8266 ( .B1(n12833), .B2(n7741), .A(n7740), .ZN(n7739) );
  NOR2_X1 U8267 ( .A1(n7745), .A2(n7746), .ZN(n7741) );
  NAND2_X1 U8268 ( .A1(n12833), .A2(n7744), .ZN(n7740) );
  NAND2_X1 U8269 ( .A1(n7743), .A2(n7744), .ZN(n7742) );
  INV_X1 U8270 ( .A(n12833), .ZN(n7743) );
  AOI21_X1 U8271 ( .B1(n13250), .B2(n8521), .A(n8448), .ZN(n13268) );
  NAND2_X1 U8272 ( .A1(n8332), .A2(n8331), .ZN(n12218) );
  AND2_X1 U8273 ( .A1(n10801), .A2(n10778), .ZN(n12929) );
  XNOR2_X1 U8274 ( .A(n12805), .B(n13170), .ZN(n12913) );
  NAND2_X1 U8275 ( .A1(n8501), .A2(n8500), .ZN(n12920) );
  OR2_X1 U8276 ( .A1(n12804), .A2(n13207), .ZN(n7337) );
  NAND2_X1 U8277 ( .A1(n11090), .A2(n12646), .ZN(n12934) );
  AND4_X1 U8278 ( .A1(n12403), .A2(n8547), .A3(n8546), .A4(n8545), .ZN(n12427)
         );
  INV_X1 U8279 ( .A(n13196), .ZN(n13170) );
  INV_X1 U8280 ( .A(n12897), .ZN(n13234) );
  INV_X1 U8281 ( .A(n13268), .ZN(n13233) );
  INV_X1 U8282 ( .A(n13266), .ZN(n13290) );
  INV_X1 U8283 ( .A(n12869), .ZN(n13303) );
  NAND2_X1 U8284 ( .A1(n8398), .A2(n8397), .ZN(n13313) );
  NAND4_X1 U8285 ( .A1(n8202), .A2(n8201), .A3(n8200), .A4(n8199), .ZN(n12953)
         );
  OR2_X1 U8286 ( .A1(n10942), .A2(n10941), .ZN(n11064) );
  AND2_X1 U8287 ( .A1(n8222), .A2(n8279), .ZN(n11574) );
  AND3_X1 U8288 ( .A1(n7488), .A2(n7487), .A3(n15914), .ZN(n13100) );
  NAND2_X1 U8289 ( .A1(n13095), .A2(n13096), .ZN(n7487) );
  OR2_X1 U8290 ( .A1(n13090), .A2(n7680), .ZN(n7679) );
  NAND2_X1 U8291 ( .A1(n7681), .A2(P3_REG2_REG_17__SCAN_IN), .ZN(n7680) );
  INV_X1 U8292 ( .A(n13141), .ZN(n15916) );
  NAND2_X1 U8293 ( .A1(n7353), .A2(n15915), .ZN(n6818) );
  OR2_X1 U8294 ( .A1(n13090), .A2(n13305), .ZN(n13108) );
  OAI21_X1 U8295 ( .B1(n13427), .B2(n13352), .A(n7415), .ZN(n7414) );
  NOR2_X1 U8296 ( .A1(n7417), .A2(n7416), .ZN(n7415) );
  INV_X1 U8297 ( .A(n8634), .ZN(n7417) );
  NOR2_X1 U8298 ( .A1(n13346), .A2(n13245), .ZN(n7412) );
  OAI21_X1 U8299 ( .B1(n13429), .B2(n13352), .A(n7098), .ZN(n7097) );
  INV_X1 U8300 ( .A(n13165), .ZN(n7098) );
  NAND2_X1 U8301 ( .A1(n8443), .A2(n8442), .ZN(n13251) );
  NAND2_X1 U8302 ( .A1(n8299), .A2(n8298), .ZN(n13411) );
  NAND2_X1 U8303 ( .A1(n15970), .A2(n8588), .ZN(n7314) );
  NAND2_X1 U8304 ( .A1(n8268), .A2(n8267), .ZN(n12551) );
  AND2_X1 U8305 ( .A1(n15973), .A2(n15960), .ZN(n13395) );
  INV_X1 U8306 ( .A(n13395), .ZN(n13403) );
  XNOR2_X1 U8307 ( .A(n12397), .B(n7786), .ZN(n13427) );
  INV_X1 U8308 ( .A(n12615), .ZN(n7786) );
  XNOR2_X1 U8309 ( .A(n7864), .B(n12615), .ZN(n7862) );
  NAND2_X1 U8310 ( .A1(n8526), .A2(n13169), .ZN(n7865) );
  INV_X1 U8311 ( .A(n7859), .ZN(n7858) );
  OAI21_X1 U8312 ( .B1(n8549), .B2(n7860), .A(n7863), .ZN(n7859) );
  NAND2_X1 U8313 ( .A1(n15961), .A2(n13424), .ZN(n7863) );
  NAND2_X1 U8314 ( .A1(n15963), .A2(n13245), .ZN(n7860) );
  XNOR2_X1 U8315 ( .A(n13151), .B(n13150), .ZN(n13429) );
  NAND2_X1 U8316 ( .A1(n13172), .A2(n8611), .ZN(n13151) );
  NOR2_X1 U8317 ( .A1(n6580), .A2(n13361), .ZN(n13434) );
  NAND2_X1 U8318 ( .A1(n8405), .A2(n8404), .ZN(n13469) );
  NAND2_X1 U8319 ( .A1(n8391), .A2(n8390), .ZN(n13477) );
  OR2_X1 U8320 ( .A1(n13416), .A2(n15961), .ZN(n13498) );
  INV_X1 U8321 ( .A(n13493), .ZN(n13480) );
  OR2_X1 U8322 ( .A1(n10897), .A2(n10921), .ZN(n8184) );
  OR2_X1 U8323 ( .A1(n15961), .A2(n15946), .ZN(n13493) );
  NAND2_X1 U8324 ( .A1(n9610), .A2(n9609), .ZN(n12026) );
  XNOR2_X1 U8325 ( .A(n13586), .B(n13587), .ZN(n13590) );
  NAND2_X1 U8326 ( .A1(n9892), .A2(n9891), .ZN(n14039) );
  NAND2_X1 U8327 ( .A1(n11877), .A2(n9628), .ZN(n9836) );
  NAND2_X1 U8328 ( .A1(n9750), .A2(n9749), .ZN(n14148) );
  NAND2_X1 U8329 ( .A1(n6937), .A2(n11715), .ZN(n11772) );
  NAND2_X1 U8330 ( .A1(n11713), .A2(n11710), .ZN(n6937) );
  OR2_X1 U8331 ( .A1(n11013), .A2(n11008), .ZN(n13736) );
  OAI21_X1 U8332 ( .B1(n10592), .B2(n9557), .A(n6791), .ZN(n9522) );
  INV_X1 U8333 ( .A(n6792), .ZN(n6791) );
  OAI22_X1 U8334 ( .A1(n9562), .A2(n10593), .B1(n6523), .B2(n10552), .ZN(n6792) );
  XNOR2_X1 U8335 ( .A(n11296), .B(n13615), .ZN(n11410) );
  AND3_X1 U8336 ( .A1(n10087), .A2(n10086), .A3(n10085), .ZN(n7516) );
  NAND2_X1 U8337 ( .A1(n9915), .A2(n9914), .ZN(n13787) );
  NAND2_X1 U8338 ( .A1(n9898), .A2(n9897), .ZN(n13788) );
  NAND2_X1 U8339 ( .A1(n9885), .A2(n9884), .ZN(n13789) );
  NAND2_X1 U8340 ( .A1(n7256), .A2(n7255), .ZN(n13820) );
  OR2_X1 U8341 ( .A1(n10574), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n7256) );
  NAND2_X1 U8342 ( .A1(n10574), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n7255) );
  NAND2_X1 U8343 ( .A1(n13865), .A2(n6618), .ZN(n10700) );
  NAND2_X1 U8344 ( .A1(n10878), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n7565) );
  NAND2_X1 U8345 ( .A1(n10700), .A2(n10699), .ZN(n10873) );
  INV_X1 U8346 ( .A(n13939), .ZN(n13941) );
  OAI21_X1 U8347 ( .B1(n13944), .B2(n15857), .A(n13943), .ZN(n7573) );
  NAND2_X1 U8348 ( .A1(n7967), .A2(n14261), .ZN(n13948) );
  OR2_X1 U8349 ( .A1(n12385), .A2(n12769), .ZN(n7965) );
  AND2_X1 U8350 ( .A1(n7962), .A2(n7961), .ZN(n7333) );
  OAI21_X1 U8351 ( .B1(n6822), .B2(n14127), .A(n14014), .ZN(n14293) );
  XNOR2_X1 U8352 ( .A(n7643), .B(n14013), .ZN(n6822) );
  AOI21_X1 U8353 ( .B1(n14017), .B2(n7644), .A(n7646), .ZN(n7643) );
  NAND2_X1 U8354 ( .A1(n7464), .A2(n7465), .ZN(n14004) );
  OR2_X1 U8355 ( .A1(n10184), .A2(n7467), .ZN(n7464) );
  OR2_X1 U8356 ( .A1(n14462), .A2(n7953), .ZN(n7954) );
  NAND2_X1 U8357 ( .A1(n12769), .A2(n14377), .ZN(n7297) );
  INV_X1 U8358 ( .A(n6868), .ZN(n6867) );
  NAND2_X1 U8359 ( .A1(n12769), .A2(n10276), .ZN(n7289) );
  NAND2_X1 U8360 ( .A1(n14460), .A2(n7674), .ZN(n9990) );
  NAND2_X1 U8361 ( .A1(n7229), .A2(n7228), .ZN(n7227) );
  INV_X1 U8362 ( .A(n14289), .ZN(n7228) );
  NAND2_X1 U8363 ( .A1(n11132), .A2(n15881), .ZN(n15906) );
  NAND2_X1 U8364 ( .A1(n6916), .A2(n6915), .ZN(n9503) );
  NOR2_X1 U8365 ( .A1(n6621), .A2(n6559), .ZN(n6915) );
  OAI21_X1 U8366 ( .B1(n14602), .B2(n7915), .A(n6653), .ZN(n10516) );
  AND2_X1 U8367 ( .A1(n7913), .A2(n7912), .ZN(n7911) );
  NAND2_X1 U8368 ( .A1(n10773), .A2(n8743), .ZN(n7442) );
  AND4_X1 U8369 ( .A1(n8897), .A2(n8896), .A3(n8895), .A4(n8894), .ZN(n14572)
         );
  OR2_X1 U8370 ( .A1(n15705), .A2(n6597), .ZN(n7136) );
  INV_X1 U8371 ( .A(n7918), .ZN(n7149) );
  NOR2_X2 U8372 ( .A1(n10525), .A2(n10520), .ZN(n15709) );
  AND3_X1 U8373 ( .A1(n8983), .A2(n8982), .A3(n8981), .ZN(n15434) );
  NAND2_X1 U8374 ( .A1(n11495), .A2(n8743), .ZN(n8942) );
  AND2_X1 U8375 ( .A1(n14690), .A2(n9194), .ZN(n14953) );
  INV_X1 U8376 ( .A(n15409), .ZN(n15428) );
  INV_X1 U8377 ( .A(n15435), .ZN(n15418) );
  INV_X1 U8378 ( .A(n15468), .ZN(n15449) );
  NOR2_X1 U8379 ( .A1(n15725), .A2(n15714), .ZN(n15745) );
  OAI21_X1 U8380 ( .B1(n15750), .B2(n15105), .A(n15104), .ZN(n7577) );
  OAI211_X1 U8381 ( .C1(n15128), .C2(n15124), .A(n15129), .B(n15123), .ZN(
        n7947) );
  OR2_X1 U8382 ( .A1(n15144), .A2(n15116), .ZN(n15124) );
  NAND2_X1 U8383 ( .A1(n15128), .A2(n15127), .ZN(n15129) );
  AOI21_X1 U8384 ( .B1(n12758), .B2(n15807), .A(n12757), .ZN(n15365) );
  NAND2_X1 U8385 ( .A1(n12756), .A2(n12755), .ZN(n12757) );
  NAND2_X1 U8386 ( .A1(n14962), .A2(n15798), .ZN(n12756) );
  INV_X1 U8387 ( .A(n15373), .ZN(n7127) );
  OAI21_X1 U8388 ( .B1(n15168), .B2(n15384), .A(n15167), .ZN(n15171) );
  NAND2_X1 U8389 ( .A1(n15246), .A2(n7704), .ZN(n15223) );
  AND2_X1 U8390 ( .A1(n15246), .A2(n9170), .ZN(n15224) );
  INV_X1 U8391 ( .A(n15281), .ZN(n15319) );
  NOR2_X1 U8392 ( .A1(n15286), .A2(n15465), .ZN(n15341) );
  NAND2_X1 U8393 ( .A1(n11387), .A2(n15178), .ZN(n15281) );
  NAND2_X1 U8394 ( .A1(n15312), .A2(n15470), .ZN(n15339) );
  AND2_X1 U8395 ( .A1(n15312), .A2(n15812), .ZN(n15290) );
  OR2_X1 U8396 ( .A1(n8022), .A2(n8027), .ZN(n8020) );
  NAND2_X1 U8397 ( .A1(n8022), .A2(n8019), .ZN(n8018) );
  NAND2_X1 U8398 ( .A1(n15820), .A2(n8021), .ZN(n8019) );
  INV_X1 U8399 ( .A(n8027), .ZN(n8021) );
  AND2_X1 U8400 ( .A1(n7994), .A2(n9191), .ZN(n7342) );
  NAND2_X1 U8401 ( .A1(n7118), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7952) );
  NOR2_X1 U8402 ( .A1(n15651), .A2(P2_ADDR_REG_9__SCAN_IN), .ZN(n7393) );
  XOR2_X1 U8403 ( .A(n15579), .B(n15578), .Z(n15656) );
  INV_X1 U8404 ( .A(n7043), .ZN(n15578) );
  OR2_X1 U8405 ( .A1(n15683), .A2(P2_ADDR_REG_13__SCAN_IN), .ZN(n7723) );
  NAND2_X1 U8406 ( .A1(n15683), .A2(P2_ADDR_REG_13__SCAN_IN), .ZN(n7721) );
  OAI21_X1 U8407 ( .B1(n7383), .B2(n7382), .A(n7380), .ZN(n15694) );
  NAND2_X1 U8408 ( .A1(n7386), .A2(n15692), .ZN(n7382) );
  OR2_X1 U8409 ( .A1(n15691), .A2(n7381), .ZN(n7380) );
  OR2_X1 U8410 ( .A1(n15691), .A2(n15690), .ZN(n7390) );
  NAND2_X1 U8411 ( .A1(n7054), .A2(n15635), .ZN(n7050) );
  MUX2_X1 U8412 ( .A(n12520), .B(n12519), .S(n12598), .Z(n12522) );
  NAND2_X1 U8413 ( .A1(n9856), .A2(n13808), .ZN(n7520) );
  AND2_X1 U8414 ( .A1(n7276), .A2(n7275), .ZN(n12577) );
  INV_X1 U8415 ( .A(n12568), .ZN(n7275) );
  OAI21_X1 U8416 ( .B1(n12559), .B2(n12558), .A(n12569), .ZN(n7276) );
  NAND2_X1 U8417 ( .A1(n6911), .A2(n6910), .ZN(n9625) );
  OR2_X1 U8418 ( .A1(n9606), .A2(n9607), .ZN(n6910) );
  NAND2_X1 U8419 ( .A1(n9592), .A2(n9596), .ZN(n6914) );
  NAND2_X1 U8420 ( .A1(n7366), .A2(n12626), .ZN(n7365) );
  INV_X1 U8421 ( .A(n12582), .ZN(n7366) );
  NAND2_X1 U8422 ( .A1(n14824), .A2(n15799), .ZN(n7016) );
  NAND2_X1 U8423 ( .A1(n14731), .A2(n7015), .ZN(n7014) );
  OR2_X1 U8424 ( .A1(n7564), .A2(n14727), .ZN(n7563) );
  NAND2_X1 U8425 ( .A1(n14730), .A2(n14732), .ZN(n7012) );
  INV_X1 U8426 ( .A(n9648), .ZN(n7531) );
  NAND2_X1 U8427 ( .A1(n14743), .A2(n14745), .ZN(n7558) );
  OAI21_X1 U8428 ( .B1(n14739), .B2(n7020), .A(n7018), .ZN(n7021) );
  NOR2_X1 U8429 ( .A1(n14738), .A2(n14741), .ZN(n7020) );
  NOR2_X1 U8430 ( .A1(n6562), .A2(n6642), .ZN(n7536) );
  NAND2_X1 U8431 ( .A1(n9715), .A2(n7983), .ZN(n7982) );
  NAND2_X1 U8432 ( .A1(n9715), .A2(n7985), .ZN(n7984) );
  NAND2_X1 U8433 ( .A1(n9696), .A2(n9695), .ZN(n7985) );
  INV_X1 U8434 ( .A(n12600), .ZN(n6766) );
  NAND2_X1 U8435 ( .A1(n7613), .A2(n9832), .ZN(n7617) );
  INV_X1 U8436 ( .A(n9831), .ZN(n7613) );
  INV_X1 U8437 ( .A(n7617), .ZN(n7622) );
  AND2_X1 U8438 ( .A1(n7620), .A2(n7618), .ZN(n6924) );
  OAI21_X1 U8439 ( .B1(n7618), .B2(n7620), .A(n7619), .ZN(n7615) );
  INV_X1 U8440 ( .A(n9844), .ZN(n7619) );
  INV_X1 U8441 ( .A(n14777), .ZN(n14778) );
  NAND2_X1 U8442 ( .A1(n14778), .A2(n7548), .ZN(n7547) );
  AND2_X1 U8443 ( .A1(n7549), .A2(n7552), .ZN(n7548) );
  NAND2_X1 U8444 ( .A1(n14778), .A2(n7552), .ZN(n7554) );
  NAND2_X1 U8445 ( .A1(n14778), .A2(n7549), .ZN(n7553) );
  AND3_X1 U8446 ( .A1(n14786), .A2(n14787), .A3(n14788), .ZN(n7546) );
  OR3_X1 U8447 ( .A1(n15289), .A2(n14785), .A3(n14784), .ZN(n14786) );
  NOR2_X1 U8448 ( .A1(n12446), .A2(n7878), .ZN(n12447) );
  NAND2_X1 U8449 ( .A1(n7526), .A2(n6569), .ZN(n7523) );
  NAND2_X1 U8450 ( .A1(n7602), .A2(n7978), .ZN(n7601) );
  NOR2_X1 U8451 ( .A1(n6575), .A2(P3_REG3_REG_25__SCAN_IN), .ZN(n8064) );
  NOR2_X1 U8452 ( .A1(n7845), .A2(n7842), .ZN(n7841) );
  INV_X1 U8453 ( .A(n8110), .ZN(n7842) );
  OR2_X1 U8454 ( .A1(n8450), .A2(n7846), .ZN(n7845) );
  INV_X1 U8455 ( .A(n8471), .ZN(n7846) );
  NAND2_X1 U8456 ( .A1(n7844), .A2(n8471), .ZN(n7843) );
  INV_X1 U8457 ( .A(n8112), .ZN(n7844) );
  INV_X1 U8458 ( .A(n8240), .ZN(n7829) );
  NAND2_X1 U8459 ( .A1(n7524), .A2(n7521), .ZN(n7525) );
  AND2_X1 U8460 ( .A1(n7523), .A2(n7522), .ZN(n7521) );
  INV_X1 U8461 ( .A(n9889), .ZN(n7522) );
  NAND2_X1 U8462 ( .A1(n9902), .A2(n9901), .ZN(n7981) );
  INV_X1 U8463 ( .A(n7674), .ZN(n7170) );
  AND2_X1 U8464 ( .A1(n9628), .A2(n10028), .ZN(n7167) );
  NOR2_X1 U8465 ( .A1(n7170), .A2(n7173), .ZN(n7162) );
  NOR2_X1 U8466 ( .A1(n10213), .A2(n7436), .ZN(n7435) );
  INV_X1 U8467 ( .A(n10211), .ZN(n7436) );
  AND2_X1 U8468 ( .A1(n10267), .A2(n15872), .ZN(n11006) );
  NOR2_X1 U8469 ( .A1(n7543), .A2(n7541), .ZN(n7540) );
  NOR2_X1 U8470 ( .A1(n15222), .A2(n15200), .ZN(n6841) );
  NAND2_X1 U8471 ( .A1(n7066), .A2(n7068), .ZN(n7065) );
  INV_X1 U8472 ( .A(n9168), .ZN(n7698) );
  INV_X1 U8473 ( .A(n14768), .ZN(n8010) );
  INV_X1 U8474 ( .A(n9971), .ZN(n7178) );
  NAND2_X1 U8475 ( .A1(n8990), .A2(n11055), .ZN(n9008) );
  NAND2_X1 U8476 ( .A1(n8967), .A2(n10892), .ZN(n8988) );
  NAND2_X1 U8477 ( .A1(n8929), .A2(n8928), .ZN(n8957) );
  AOI21_X1 U8478 ( .B1(n8826), .B2(n8829), .A(n8843), .ZN(n7606) );
  OAI21_X1 U8479 ( .B1(n10579), .B2(n10665), .A(n6872), .ZN(n6871) );
  NAND2_X1 U8480 ( .A1(n10579), .A2(P2_DATAO_REG_9__SCAN_IN), .ZN(n6872) );
  INV_X1 U8481 ( .A(n7447), .ZN(n7446) );
  OAI21_X1 U8482 ( .B1(n8750), .B2(n7448), .A(n8773), .ZN(n7447) );
  INV_X1 U8483 ( .A(n8754), .ZN(n7448) );
  OAI21_X1 U8484 ( .B1(n15592), .B2(P1_ADDR_REG_3__SCAN_IN), .A(n6645), .ZN(
        n7724) );
  NOR2_X1 U8485 ( .A1(n8475), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n8063) );
  INV_X1 U8486 ( .A(n12277), .ZN(n7734) );
  NAND2_X1 U8487 ( .A1(n12397), .A2(n12440), .ZN(n12438) );
  NOR2_X1 U8488 ( .A1(n12459), .A2(n13167), .ZN(n7839) );
  AND2_X1 U8489 ( .A1(n12617), .A2(n12413), .ZN(n12621) );
  NOR2_X1 U8490 ( .A1(n10925), .A2(n10954), .ZN(n7062) );
  AOI21_X1 U8491 ( .B1(n7660), .B2(n11062), .A(n6632), .ZN(n7659) );
  INV_X1 U8492 ( .A(n11063), .ZN(n7660) );
  NAND2_X1 U8493 ( .A1(n6895), .A2(P3_REG2_REG_5__SCAN_IN), .ZN(n6894) );
  INV_X1 U8494 ( .A(n12085), .ZN(n6795) );
  NAND2_X1 U8495 ( .A1(n7095), .A2(n7094), .ZN(n13048) );
  INV_X1 U8496 ( .A(n13046), .ZN(n7094) );
  NAND2_X1 U8497 ( .A1(n7488), .A2(n7486), .ZN(n7335) );
  XNOR2_X1 U8498 ( .A(n7335), .B(n7334), .ZN(n13114) );
  AND2_X1 U8499 ( .A1(n7300), .A2(n8064), .ZN(n8503) );
  INV_X1 U8500 ( .A(P3_REG3_REG_26__SCAN_IN), .ZN(n7300) );
  OAI21_X1 U8501 ( .B1(n13193), .B2(n7869), .A(n8511), .ZN(n7868) );
  AND2_X1 U8502 ( .A1(n12441), .A2(n13223), .ZN(n7005) );
  NOR2_X1 U8503 ( .A1(n6624), .A2(n7004), .ZN(n7001) );
  NOR2_X1 U8504 ( .A1(n7003), .A2(n6996), .ZN(n6995) );
  INV_X1 U8505 ( .A(n8439), .ZN(n6996) );
  INV_X1 U8506 ( .A(n6586), .ZN(n7003) );
  INV_X1 U8507 ( .A(n8449), .ZN(n7002) );
  AND2_X1 U8508 ( .A1(n7762), .A2(n12442), .ZN(n7757) );
  AND2_X1 U8509 ( .A1(n7112), .A2(n7111), .ZN(n7110) );
  AND2_X1 U8510 ( .A1(n8360), .A2(n7113), .ZN(n7112) );
  INV_X1 U8511 ( .A(P3_REG3_REG_16__SCAN_IN), .ZN(n7113) );
  INV_X1 U8512 ( .A(P3_REG3_REG_12__SCAN_IN), .ZN(n7116) );
  AND2_X1 U8513 ( .A1(n8284), .A2(n8300), .ZN(n7117) );
  NOR2_X1 U8514 ( .A1(n10796), .A2(n11190), .ZN(n10730) );
  OAI21_X1 U8515 ( .B1(n6582), .B2(n7773), .A(n12620), .ZN(n7772) );
  NOR2_X1 U8516 ( .A1(n13289), .A2(n8603), .ZN(n13257) );
  INV_X1 U8517 ( .A(n8351), .ZN(n6982) );
  AND2_X1 U8518 ( .A1(n12573), .A2(n7874), .ZN(n7873) );
  NAND2_X1 U8519 ( .A1(n12453), .A2(n8325), .ZN(n7874) );
  NOR2_X1 U8520 ( .A1(n8512), .A2(n8498), .ZN(n7816) );
  INV_X1 U8521 ( .A(n8124), .ZN(n7818) );
  NAND2_X1 U8522 ( .A1(n8131), .A2(n7370), .ZN(n7493) );
  NOR2_X1 U8523 ( .A1(n7494), .A2(n13504), .ZN(n7370) );
  NAND2_X1 U8524 ( .A1(n8113), .A2(n15547), .ZN(n8116) );
  NOR2_X1 U8525 ( .A1(n6581), .A2(n7823), .ZN(n7822) );
  INV_X1 U8526 ( .A(n8087), .ZN(n7823) );
  INV_X1 U8527 ( .A(n6592), .ZN(n6930) );
  AOI21_X1 U8528 ( .B1(n6947), .B2(n6945), .A(n13543), .ZN(n6944) );
  INV_X1 U8529 ( .A(n6947), .ZN(n6946) );
  NOR2_X1 U8530 ( .A1(n13935), .A2(n6723), .ZN(n13937) );
  INV_X1 U8531 ( .A(n7966), .ZN(n7964) );
  NAND2_X1 U8532 ( .A1(n14008), .A2(n6888), .ZN(n6887) );
  NAND2_X1 U8533 ( .A1(n7647), .A2(n10246), .ZN(n7645) );
  NOR2_X1 U8534 ( .A1(n7428), .A2(n7424), .ZN(n7423) );
  INV_X1 U8535 ( .A(n10241), .ZN(n7424) );
  AND2_X1 U8536 ( .A1(n14034), .A2(n7427), .ZN(n7426) );
  OR2_X1 U8537 ( .A1(n14056), .A2(n7428), .ZN(n7427) );
  AND2_X1 U8538 ( .A1(n7668), .A2(n14424), .ZN(n7973) );
  INV_X1 U8539 ( .A(n10236), .ZN(n7662) );
  NOR2_X1 U8540 ( .A1(n9786), .A2(n9767), .ZN(n6763) );
  NAND2_X1 U8541 ( .A1(n10199), .A2(n7969), .ZN(n7970) );
  NOR2_X1 U8542 ( .A1(n10210), .A2(n11930), .ZN(n7960) );
  INV_X1 U8543 ( .A(n11353), .ZN(n11002) );
  NAND2_X1 U8544 ( .A1(n6884), .A2(n10227), .ZN(n14176) );
  NAND2_X1 U8545 ( .A1(n7434), .A2(n10212), .ZN(n12001) );
  NAND4_X1 U8546 ( .A1(n6785), .A2(n10095), .A3(n7794), .A4(n9500), .ZN(n7793)
         );
  NOR2_X1 U8547 ( .A1(P2_IR_REG_25__SCAN_IN), .A2(P2_IR_REG_26__SCAN_IN), .ZN(
        n7972) );
  OR2_X1 U8548 ( .A1(n9699), .A2(P2_IR_REG_6__SCAN_IN), .ZN(n9629) );
  NOR2_X1 U8549 ( .A1(n8915), .A2(n8914), .ZN(n8943) );
  INV_X1 U8550 ( .A(n7896), .ZN(n7895) );
  AOI21_X1 U8551 ( .B1(n7896), .B2(n7894), .A(n7893), .ZN(n7892) );
  INV_X1 U8552 ( .A(n10355), .ZN(n7893) );
  NOR2_X1 U8553 ( .A1(n8978), .A2(n8977), .ZN(n7318) );
  MUX2_X1 U8554 ( .A(n14846), .B(n15114), .S(n14719), .Z(n14894) );
  NAND2_X1 U8555 ( .A1(n7306), .A2(n7305), .ZN(n14859) );
  NAND2_X1 U8556 ( .A1(n15344), .A2(n14719), .ZN(n7305) );
  OR2_X1 U8557 ( .A1(n15344), .A2(n7307), .ZN(n7306) );
  OR2_X1 U8558 ( .A1(n15119), .A2(n15118), .ZN(n15125) );
  NOR2_X1 U8559 ( .A1(n15379), .A2(n7126), .ZN(n7125) );
  NAND2_X1 U8560 ( .A1(n7127), .A2(n15187), .ZN(n7126) );
  AND2_X1 U8561 ( .A1(n12734), .A2(n15158), .ZN(n12735) );
  OR2_X1 U8562 ( .A1(n15148), .A2(n12733), .ZN(n12734) );
  INV_X1 U8563 ( .A(n6749), .ZN(n9105) );
  NOR2_X1 U8564 ( .A1(n15313), .A2(n7122), .ZN(n8033) );
  NAND2_X1 U8565 ( .A1(n8986), .A2(n15308), .ZN(n7251) );
  NAND2_X1 U8566 ( .A1(n8943), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n8978) );
  NOR2_X1 U8567 ( .A1(n8857), .A2(n8856), .ZN(n7321) );
  INV_X1 U8568 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n8811) );
  NAND2_X1 U8569 ( .A1(n11848), .A2(n8771), .ZN(n12148) );
  NAND2_X1 U8570 ( .A1(n8771), .A2(n8769), .ZN(n11850) );
  NOR2_X1 U8571 ( .A1(n7945), .A2(n14725), .ZN(n7944) );
  NAND2_X1 U8572 ( .A1(n14835), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n8666) );
  INV_X1 U8574 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n6826) );
  NAND2_X1 U8575 ( .A1(n9212), .A2(n8661), .ZN(n8026) );
  INV_X1 U8576 ( .A(n7920), .ZN(n7179) );
  NOR2_X1 U8577 ( .A1(P1_IR_REG_27__SCAN_IN), .A2(P1_IR_REG_26__SCAN_IN), .ZN(
        n8024) );
  OAI21_X1 U8578 ( .B1(n10004), .B2(n13522), .A(n10002), .ZN(n9985) );
  AOI21_X1 U8579 ( .B1(n7927), .B2(n7929), .A(n7925), .ZN(n7924) );
  INV_X1 U8580 ( .A(n9087), .ZN(n7925) );
  NAND2_X1 U8581 ( .A1(n9009), .A2(n7927), .ZN(n7187) );
  NAND2_X1 U8582 ( .A1(n7926), .A2(n9048), .ZN(n9081) );
  AND2_X1 U8583 ( .A1(n7900), .A2(n9361), .ZN(n7899) );
  NOR2_X1 U8584 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(P1_IR_REG_19__SCAN_IN), .ZN(
        n7900) );
  XNOR2_X1 U8585 ( .A(n9081), .B(n11752), .ZN(n9062) );
  NOR2_X1 U8586 ( .A1(n7308), .A2(P1_IR_REG_18__SCAN_IN), .ZN(n7147) );
  NAND2_X1 U8587 ( .A1(n8907), .A2(n6599), .ZN(n8904) );
  NAND2_X1 U8588 ( .A1(n8869), .A2(n10653), .ZN(n8903) );
  OR3_X1 U8589 ( .A1(n8852), .A2(P1_IR_REG_9__SCAN_IN), .A3(n8851), .ZN(n8873)
         );
  NAND2_X1 U8590 ( .A1(n8867), .A2(n8848), .ZN(n8865) );
  NAND2_X1 U8591 ( .A1(n6871), .A2(SI_9_), .ZN(n8829) );
  AND2_X1 U8592 ( .A1(n8827), .A2(n7454), .ZN(n7453) );
  INV_X1 U8593 ( .A(n8826), .ZN(n8827) );
  NAND2_X1 U8594 ( .A1(n8806), .A2(n8793), .ZN(n7454) );
  AOI21_X1 U8595 ( .B1(n8791), .B2(n7192), .A(n7191), .ZN(n7190) );
  INV_X1 U8596 ( .A(n8790), .ZN(n7192) );
  XNOR2_X1 U8597 ( .A(n6871), .B(SI_9_), .ZN(n8826) );
  INV_X1 U8598 ( .A(n8720), .ZN(n7154) );
  NAND2_X1 U8599 ( .A1(n6533), .A2(n10591), .ZN(n8703) );
  OR2_X1 U8600 ( .A1(n6532), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n7938) );
  OAI21_X1 U8601 ( .B1(n10580), .B2(n10575), .A(n7458), .ZN(n8700) );
  NAND2_X1 U8602 ( .A1(n6533), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n7458) );
  INV_X1 U8603 ( .A(P1_RD_REG_SCAN_IN), .ZN(n8133) );
  INV_X1 U8604 ( .A(P2_RD_REG_SCAN_IN), .ZN(n8135) );
  XNOR2_X1 U8605 ( .A(P3_ADDR_REG_1__SCAN_IN), .B(P1_ADDR_REG_1__SCAN_IN), 
        .ZN(n15585) );
  XNOR2_X1 U8606 ( .A(n7724), .B(n7501), .ZN(n15580) );
  OAI211_X1 U8607 ( .C1(n15596), .C2(n7036), .A(n7035), .B(n6713), .ZN(n7504)
         );
  NAND2_X1 U8608 ( .A1(n7038), .A2(n7037), .ZN(n7036) );
  XNOR2_X1 U8609 ( .A(n11759), .B(n15933), .ZN(n11216) );
  NOR2_X1 U8610 ( .A1(n12831), .A2(n7747), .ZN(n7746) );
  INV_X1 U8611 ( .A(n12913), .ZN(n7747) );
  NAND2_X1 U8612 ( .A1(n7235), .A2(n7234), .ZN(n10789) );
  NAND2_X1 U8613 ( .A1(n12832), .A2(n12496), .ZN(n7234) );
  NAND2_X1 U8614 ( .A1(n12119), .A2(n12118), .ZN(n12170) );
  AND2_X1 U8615 ( .A1(n12793), .A2(n12813), .ZN(n7267) );
  INV_X1 U8616 ( .A(n7350), .ZN(n7732) );
  NAND2_X1 U8617 ( .A1(n11453), .A2(n11454), .ZN(n11800) );
  INV_X1 U8618 ( .A(n12778), .ZN(n7728) );
  AND4_X1 U8619 ( .A1(n12403), .A2(n12402), .A3(n12401), .A4(n12400), .ZN(
        n13144) );
  AND4_X1 U8620 ( .A1(n8229), .A2(n8228), .A3(n8227), .A4(n8226), .ZN(n11795)
         );
  XNOR2_X1 U8621 ( .A(n8207), .B(n8206), .ZN(n10944) );
  OR2_X1 U8622 ( .A1(n10902), .A2(n10901), .ZN(n10905) );
  NAND2_X1 U8623 ( .A1(n12962), .A2(n10932), .ZN(n7061) );
  NAND2_X1 U8624 ( .A1(n6894), .A2(n10971), .ZN(n6774) );
  NAND2_X1 U8625 ( .A1(n6800), .A2(n6799), .ZN(n10964) );
  AOI21_X1 U8626 ( .B1(n6798), .B2(n11069), .A(n6550), .ZN(n6799) );
  NOR2_X1 U8627 ( .A1(n6797), .A2(n6803), .ZN(n6796) );
  NAND2_X1 U8628 ( .A1(n7077), .A2(n6552), .ZN(n11043) );
  NAND2_X1 U8629 ( .A1(n11104), .A2(n7078), .ZN(n7077) );
  NAND2_X1 U8630 ( .A1(n7655), .A2(P3_REG2_REG_7__SCAN_IN), .ZN(n11197) );
  NAND2_X1 U8631 ( .A1(n7075), .A2(n7074), .ZN(n7069) );
  OAI21_X1 U8632 ( .B1(n11191), .B2(n6790), .A(n6787), .ZN(n11576) );
  INV_X1 U8633 ( .A(n11194), .ZN(n6790) );
  NAND2_X1 U8634 ( .A1(n7655), .A2(n6583), .ZN(n7408) );
  AOI21_X1 U8635 ( .B1(n7655), .B2(n6612), .A(n7407), .ZN(n7406) );
  NOR2_X1 U8636 ( .A1(n6553), .A2(n11578), .ZN(n7407) );
  NOR2_X1 U8637 ( .A1(n7649), .A2(n12975), .ZN(n7648) );
  NOR2_X1 U8638 ( .A1(n12094), .A2(n12093), .ZN(n12096) );
  XNOR2_X1 U8639 ( .A(n13048), .B(n7093), .ZN(n13050) );
  NAND2_X1 U8640 ( .A1(n13050), .A2(n13049), .ZN(n13066) );
  NAND2_X1 U8641 ( .A1(n6810), .A2(n6809), .ZN(n13062) );
  INV_X1 U8642 ( .A(n6811), .ZN(n6810) );
  OAI21_X1 U8643 ( .B1(n6814), .B2(n13039), .A(n13043), .ZN(n6811) );
  NAND2_X1 U8644 ( .A1(n6890), .A2(n7682), .ZN(n13077) );
  OAI21_X1 U8645 ( .B1(n13067), .B2(n7093), .A(n13066), .ZN(n13094) );
  INV_X1 U8646 ( .A(n13048), .ZN(n13067) );
  OAI21_X1 U8647 ( .B1(n13120), .B2(n7498), .A(n15914), .ZN(n7497) );
  AND2_X1 U8648 ( .A1(n13114), .A2(n13115), .ZN(n7498) );
  AOI22_X1 U8649 ( .A1(n13104), .A2(P3_REG1_REG_17__SCAN_IN), .B1(n13112), 
        .B2(n13103), .ZN(n13134) );
  INV_X1 U8650 ( .A(n7335), .ZN(n13121) );
  NOR2_X1 U8651 ( .A1(n13114), .A2(n13115), .ZN(n13120) );
  AND4_X1 U8652 ( .A1(n8525), .A2(n8524), .A3(n8523), .A4(n8522), .ZN(n13181)
         );
  NOR2_X1 U8653 ( .A1(n8444), .A2(P3_REG3_REG_21__SCAN_IN), .ZN(n8454) );
  OR2_X1 U8654 ( .A1(n8431), .A2(P3_REG3_REG_20__SCAN_IN), .ZN(n8444) );
  NAND2_X1 U8655 ( .A1(n8419), .A2(n8418), .ZN(n8431) );
  AND2_X1 U8656 ( .A1(n8361), .A2(n7108), .ZN(n8419) );
  AND2_X1 U8657 ( .A1(n7110), .A2(n7109), .ZN(n7108) );
  INV_X1 U8658 ( .A(P3_REG3_REG_18__SCAN_IN), .ZN(n7109) );
  NAND2_X1 U8659 ( .A1(n8361), .A2(n7110), .ZN(n8406) );
  NAND2_X1 U8660 ( .A1(n8361), .A2(n8360), .ZN(n8377) );
  NAND2_X1 U8661 ( .A1(n8361), .A2(n7112), .ZN(n8392) );
  AND2_X1 U8662 ( .A1(n8347), .A2(n8346), .ZN(n8361) );
  AND2_X1 U8663 ( .A1(n8285), .A2(n7114), .ZN(n8347) );
  AND2_X1 U8664 ( .A1(n6703), .A2(n7115), .ZN(n7114) );
  INV_X1 U8665 ( .A(P3_REG3_REG_13__SCAN_IN), .ZN(n7115) );
  NAND2_X1 U8666 ( .A1(n8285), .A2(n6703), .ZN(n8335) );
  INV_X1 U8667 ( .A(P3_REG3_REG_11__SCAN_IN), .ZN(n8300) );
  NAND2_X1 U8668 ( .A1(n8285), .A2(n7117), .ZN(n8319) );
  AND2_X1 U8669 ( .A1(n8285), .A2(n8284), .ZN(n8301) );
  NOR2_X1 U8670 ( .A1(n8269), .A2(P3_REG3_REG_9__SCAN_IN), .ZN(n8285) );
  AND2_X1 U8671 ( .A1(n12350), .A2(n8230), .ZN(n7103) );
  AND2_X1 U8672 ( .A1(n8062), .A2(n7105), .ZN(n7102) );
  AND2_X1 U8673 ( .A1(n7106), .A2(n7104), .ZN(n8249) );
  AND2_X1 U8674 ( .A1(n7107), .A2(n7105), .ZN(n7104) );
  NAND2_X1 U8675 ( .A1(n7106), .A2(n7107), .ZN(n8250) );
  OR2_X1 U8676 ( .A1(n12952), .A2(n15933), .ZN(n12512) );
  NAND2_X1 U8677 ( .A1(n12350), .A2(n8062), .ZN(n9440) );
  NAND2_X2 U8678 ( .A1(n12504), .A2(n12509), .ZN(n12445) );
  INV_X1 U8679 ( .A(n10730), .ZN(n12494) );
  NAND2_X1 U8680 ( .A1(n12412), .A2(n12411), .ZN(n13147) );
  NAND2_X1 U8681 ( .A1(n8426), .A2(n8425), .ZN(n13262) );
  INV_X1 U8682 ( .A(n12443), .ZN(n13311) );
  NAND2_X1 U8683 ( .A1(n11949), .A2(n12566), .ZN(n12059) );
  NAND2_X1 U8684 ( .A1(n8595), .A2(n12538), .ZN(n11401) );
  AND2_X1 U8685 ( .A1(n12546), .A2(n12545), .ZN(n12450) );
  INV_X1 U8686 ( .A(n8214), .ZN(n8374) );
  AND3_X1 U8687 ( .A1(n10704), .A2(n10707), .A3(n10703), .ZN(n10801) );
  NAND2_X1 U8688 ( .A1(n12408), .A2(n12407), .ZN(n12416) );
  NAND2_X1 U8689 ( .A1(n8529), .A2(n8528), .ZN(n12406) );
  NOR2_X1 U8690 ( .A1(n8312), .A2(P3_IR_REG_27__SCAN_IN), .ZN(n7784) );
  INV_X1 U8691 ( .A(P3_IR_REG_28__SCAN_IN), .ZN(n8129) );
  OAI21_X1 U8692 ( .B1(n8462), .B2(n14473), .A(n8116), .ZN(n8487) );
  NAND2_X1 U8693 ( .A1(n7330), .A2(n7329), .ZN(n8540) );
  INV_X1 U8694 ( .A(n8553), .ZN(n7330) );
  INV_X1 U8695 ( .A(n7853), .ZN(n7852) );
  AOI21_X1 U8696 ( .B1(n7851), .B2(n7853), .A(n7850), .ZN(n7849) );
  NOR2_X1 U8697 ( .A1(n8400), .A2(n6706), .ZN(n7853) );
  OR2_X1 U8698 ( .A1(n8313), .A2(P3_IR_REG_6__SCAN_IN), .ZN(n8237) );
  INV_X1 U8699 ( .A(P3_IR_REG_5__SCAN_IN), .ZN(n8215) );
  XNOR2_X1 U8700 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(P2_DATAO_REG_4__SCAN_IN), 
        .ZN(n8145) );
  NAND2_X1 U8701 ( .A1(n7812), .A2(n8074), .ZN(n7811) );
  NAND2_X1 U8702 ( .A1(n11409), .A2(n11408), .ZN(n6927) );
  OR2_X1 U8703 ( .A1(n11415), .A2(n11414), .ZN(n11416) );
  XNOR2_X1 U8704 ( .A(n9522), .B(n11422), .ZN(n11414) );
  AND2_X1 U8705 ( .A1(n13561), .A2(n13560), .ZN(n13619) );
  OAI21_X1 U8706 ( .B1(n13586), .B2(n7636), .A(n6643), .ZN(n7635) );
  NAND2_X1 U8707 ( .A1(n13548), .A2(n7637), .ZN(n7636) );
  NAND2_X1 U8708 ( .A1(n13652), .A2(n13588), .ZN(n7637) );
  XNOR2_X1 U8709 ( .A(n11506), .B(n11422), .ZN(n11714) );
  NAND2_X1 U8710 ( .A1(n12651), .A2(n12189), .ZN(n12190) );
  NAND2_X1 U8711 ( .A1(n6760), .A2(n6705), .ZN(n9719) );
  INV_X1 U8712 ( .A(n9704), .ZN(n6760) );
  AND2_X1 U8713 ( .A1(n11007), .A2(n10102), .ZN(n13770) );
  AND2_X1 U8714 ( .A1(n11007), .A2(n10103), .ZN(n13769) );
  NAND2_X1 U8715 ( .A1(n11413), .A2(n11412), .ZN(n11409) );
  NAND2_X1 U8716 ( .A1(n13585), .A2(n12676), .ZN(n13666) );
  NOR2_X1 U8717 ( .A1(n10077), .A2(n7196), .ZN(n10086) );
  NOR4_X1 U8718 ( .A1(n10076), .A2(n10135), .A3(n6647), .A4(n10075), .ZN(
        n10077) );
  NAND2_X1 U8719 ( .A1(n7292), .A2(n7291), .ZN(n7290) );
  AOI21_X1 U8720 ( .B1(n9919), .B2(n9918), .A(n9920), .ZN(n7519) );
  NOR2_X1 U8721 ( .A1(n10134), .A2(n7647), .ZN(n7934) );
  INV_X1 U8722 ( .A(n10142), .ZN(n7935) );
  AND3_X1 U8723 ( .A1(n9827), .A2(n9826), .A3(n9825), .ZN(n12686) );
  AND4_X1 U8724 ( .A1(n9774), .A2(n9773), .A3(n9772), .A4(n9771), .ZN(n13670)
         );
  AND4_X1 U8725 ( .A1(n9681), .A2(n9680), .A3(n9679), .A4(n9678), .ZN(n13731)
         );
  AND4_X1 U8726 ( .A1(n9659), .A2(n9658), .A3(n9657), .A4(n9656), .ZN(n10220)
         );
  NAND2_X1 U8727 ( .A1(n10566), .A2(n10567), .ZN(n10691) );
  NAND2_X1 U8728 ( .A1(n15831), .A2(n15832), .ZN(n15829) );
  NAND2_X1 U8729 ( .A1(n11171), .A2(n11170), .ZN(n6964) );
  AOI21_X1 U8730 ( .B1(P2_REG1_REG_10__SCAN_IN), .B2(n11655), .A(n11654), .ZN(
        n11657) );
  NOR2_X1 U8731 ( .A1(n11657), .A2(n11656), .ZN(n11823) );
  INV_X1 U8732 ( .A(n11652), .ZN(n7253) );
  AOI21_X1 U8733 ( .B1(n6956), .B2(n6540), .A(n6955), .ZN(n13884) );
  INV_X1 U8734 ( .A(n6957), .ZN(n6955) );
  INV_X1 U8735 ( .A(n12304), .ZN(n6956) );
  AOI21_X1 U8736 ( .B1(n6540), .B2(n6960), .A(n12306), .ZN(n6957) );
  NAND2_X1 U8737 ( .A1(n12304), .A2(n6959), .ZN(n6958) );
  NOR2_X1 U8738 ( .A1(n13884), .A2(n7572), .ZN(n13902) );
  AND2_X1 U8739 ( .A1(n13885), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n7572) );
  NAND2_X1 U8740 ( .A1(n6954), .A2(n13931), .ZN(n6953) );
  INV_X1 U8741 ( .A(n13937), .ZN(n6954) );
  AND3_X1 U8742 ( .A1(n6953), .A2(n6952), .A3(P2_REG1_REG_18__SCAN_IN), .ZN(
        n15859) );
  OR2_X1 U8743 ( .A1(n13934), .A2(n13933), .ZN(n6757) );
  NAND2_X1 U8744 ( .A1(n12385), .A2(n7963), .ZN(n7962) );
  NOR2_X1 U8745 ( .A1(n7964), .A2(n13945), .ZN(n7963) );
  NAND2_X1 U8746 ( .A1(n7964), .A2(n13945), .ZN(n7961) );
  NOR2_X1 U8747 ( .A1(n12376), .A2(n14127), .ZN(n7430) );
  NOR2_X1 U8748 ( .A1(n6551), .A2(n12381), .ZN(n7431) );
  NAND3_X1 U8749 ( .A1(n12390), .A2(n7356), .A3(n14261), .ZN(n13958) );
  OR2_X1 U8750 ( .A1(n12385), .A2(n13962), .ZN(n7356) );
  AND2_X1 U8751 ( .A1(n13959), .A2(n9942), .ZN(n13968) );
  INV_X1 U8752 ( .A(n6875), .ZN(n6874) );
  NAND2_X1 U8753 ( .A1(n14017), .A2(n6877), .ZN(n6876) );
  NAND2_X1 U8754 ( .A1(n7355), .A2(n6886), .ZN(n13997) );
  INV_X1 U8755 ( .A(n6887), .ZN(n6886) );
  OR2_X1 U8756 ( .A1(n9908), .A2(n9907), .ZN(n10029) );
  INV_X1 U8757 ( .A(n10246), .ZN(n7646) );
  NAND2_X1 U8758 ( .A1(n7355), .A2(n14008), .ZN(n14006) );
  AOI21_X1 U8759 ( .B1(n7806), .B2(n7466), .A(n6641), .ZN(n7465) );
  INV_X1 U8760 ( .A(n6579), .ZN(n7466) );
  NOR2_X1 U8761 ( .A1(n14070), .A2(n14417), .ZN(n14050) );
  OR2_X1 U8762 ( .A1(n9862), .A2(n9861), .ZN(n9878) );
  NAND2_X1 U8763 ( .A1(n7668), .A2(n13791), .ZN(n7667) );
  NAND2_X1 U8764 ( .A1(n7665), .A2(n10237), .ZN(n7663) );
  NAND2_X1 U8765 ( .A1(n6762), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n9862) );
  INV_X1 U8766 ( .A(n10177), .ZN(n7797) );
  NOR2_X1 U8767 ( .A1(n14335), .A2(n14341), .ZN(n7974) );
  AND2_X1 U8768 ( .A1(n14114), .A2(n14424), .ZN(n14084) );
  INV_X1 U8769 ( .A(n6762), .ZN(n9838) );
  NAND2_X1 U8770 ( .A1(n6763), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n9753) );
  NAND2_X1 U8771 ( .A1(n9735), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n9821) );
  INV_X1 U8772 ( .A(n9753), .ZN(n9735) );
  NAND2_X1 U8773 ( .A1(n10201), .A2(n14131), .ZN(n14129) );
  INV_X1 U8774 ( .A(n14146), .ZN(n10201) );
  INV_X1 U8775 ( .A(n6763), .ZN(n9769) );
  INV_X1 U8776 ( .A(n10230), .ZN(n14159) );
  NAND2_X1 U8777 ( .A1(n6806), .A2(n10226), .ZN(n6805) );
  NAND2_X1 U8778 ( .A1(n6808), .A2(n6609), .ZN(n6806) );
  XNOR2_X1 U8779 ( .A(n14435), .B(n10119), .ZN(n14180) );
  OR2_X1 U8780 ( .A1(n9784), .A2(n9783), .ZN(n9786) );
  NAND2_X1 U8781 ( .A1(n6759), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n9784) );
  INV_X1 U8782 ( .A(n9719), .ZN(n6759) );
  NAND2_X1 U8783 ( .A1(n10200), .A2(n13712), .ZN(n14175) );
  AOI21_X1 U8784 ( .B1(n7470), .B2(n7475), .A(n6619), .ZN(n7468) );
  NOR2_X1 U8785 ( .A1(n10165), .A2(n7471), .ZN(n7470) );
  NOR2_X1 U8786 ( .A1(n7970), .A2(n14443), .ZN(n14208) );
  NAND2_X1 U8787 ( .A1(n9674), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n9704) );
  INV_X1 U8788 ( .A(n9676), .ZN(n9674) );
  NAND2_X1 U8789 ( .A1(n9636), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n9653) );
  INV_X1 U8790 ( .A(n9638), .ZN(n9636) );
  INV_X1 U8791 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n9652) );
  OR2_X1 U8792 ( .A1(n9653), .A2(n9652), .ZN(n9676) );
  NAND2_X1 U8793 ( .A1(n10199), .A2(n10198), .ZN(n14247) );
  NAND2_X1 U8794 ( .A1(n10218), .A2(n10217), .ZN(n14268) );
  NAND2_X1 U8795 ( .A1(n12024), .A2(n14393), .ZN(n14260) );
  NAND2_X1 U8796 ( .A1(n9615), .A2(n9614), .ZN(n9638) );
  AND2_X1 U8797 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_REG3_REG_7__SCAN_IN), 
        .ZN(n9614) );
  INV_X1 U8798 ( .A(n9613), .ZN(n9615) );
  NAND2_X1 U8799 ( .A1(n7960), .A2(n11564), .ZN(n12010) );
  NAND2_X1 U8800 ( .A1(n9573), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n9613) );
  INV_X1 U8801 ( .A(n9575), .ZN(n9573) );
  NAND2_X1 U8802 ( .A1(n11564), .A2(n11506), .ZN(n11931) );
  NAND2_X1 U8803 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n9575) );
  OR2_X1 U8804 ( .A1(n11252), .A2(n9522), .ZN(n11565) );
  NOR2_X1 U8805 ( .A1(n13955), .A2(n7485), .ZN(n7484) );
  OR2_X1 U8806 ( .A1(n12382), .A2(n13954), .ZN(n7485) );
  NAND2_X1 U8807 ( .A1(n11126), .A2(n11964), .ZN(n14307) );
  NAND2_X1 U8808 ( .A1(n7425), .A2(n10243), .ZN(n14035) );
  NAND2_X1 U8809 ( .A1(n14057), .A2(n14056), .ZN(n7425) );
  AND2_X1 U8810 ( .A1(n7968), .A2(n9701), .ZN(n14368) );
  NAND2_X1 U8811 ( .A1(n11112), .A2(n9628), .ZN(n7968) );
  INV_X1 U8812 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n6949) );
  AND2_X1 U8813 ( .A1(n14451), .A2(P2_IR_REG_19__SCAN_IN), .ZN(n6917) );
  INV_X1 U8814 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n6922) );
  AND2_X1 U8815 ( .A1(n6542), .A2(n9500), .ZN(n10096) );
  INV_X1 U8816 ( .A(n6785), .ZN(n9698) );
  INV_X2 U8817 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n9568) );
  CLKBUF_X1 U8818 ( .A(n9542), .Z(n9543) );
  NAND2_X1 U8819 ( .A1(n6532), .A2(n6625), .ZN(n9491) );
  INV_X1 U8820 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n9488) );
  NAND2_X1 U8821 ( .A1(n6532), .A2(SI_0_), .ZN(n9489) );
  INV_X1 U8822 ( .A(n15139), .ZN(n15352) );
  INV_X1 U8823 ( .A(n10514), .ZN(n7913) );
  NAND2_X1 U8824 ( .A1(n7914), .A2(n7910), .ZN(n7907) );
  INV_X1 U8825 ( .A(n8943), .ZN(n8945) );
  AND2_X1 U8826 ( .A1(n7897), .A2(n10345), .ZN(n7896) );
  INV_X1 U8827 ( .A(n14548), .ZN(n7897) );
  NAND2_X1 U8828 ( .A1(n14478), .A2(n14477), .ZN(n7898) );
  INV_X1 U8829 ( .A(n7318), .ZN(n9001) );
  INV_X1 U8830 ( .A(n7319), .ZN(n9069) );
  OR2_X1 U8831 ( .A1(n8892), .A2(n8891), .ZN(n8915) );
  NAND2_X1 U8832 ( .A1(n6753), .A2(n6752), .ZN(n6751) );
  XNOR2_X1 U8833 ( .A(n10293), .B(n14529), .ZN(n10297) );
  NAND2_X1 U8834 ( .A1(n10434), .A2(n10433), .ZN(n14664) );
  OR2_X1 U8835 ( .A1(n14823), .A2(n10295), .ZN(n10496) );
  NAND2_X1 U8837 ( .A1(n7882), .A2(n7880), .ZN(n14585) );
  AND2_X1 U8838 ( .A1(n7881), .A2(n10405), .ZN(n7880) );
  OAI21_X1 U8839 ( .B1(n14655), .B2(n7145), .A(n7142), .ZN(n7882) );
  NAND2_X1 U8840 ( .A1(n14819), .A2(n14821), .ZN(n7027) );
  NOR2_X1 U8841 ( .A1(n14886), .A2(n14888), .ZN(n14912) );
  AOI22_X1 U8842 ( .A1(n14891), .A2(n14890), .B1(n14889), .B2(n14888), .ZN(
        n14909) );
  OR4_X1 U8843 ( .A1(n14945), .A2(n15262), .A3(n15271), .A4(n14944), .ZN(
        n14946) );
  AND2_X1 U8844 ( .A1(n10510), .A2(n10509), .ZN(n14867) );
  AND2_X1 U8845 ( .A1(n15078), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n6764) );
  INV_X1 U8846 ( .A(n12746), .ZN(n6833) );
  INV_X1 U8847 ( .A(n15142), .ZN(n6830) );
  INV_X1 U8848 ( .A(n6832), .ZN(n6831) );
  OAI21_X1 U8849 ( .B1(n8041), .B2(n6833), .A(n15119), .ZN(n6832) );
  AND2_X1 U8850 ( .A1(n10532), .A2(n15132), .ZN(n14535) );
  NAND2_X1 U8851 ( .A1(n12747), .A2(n12746), .ZN(n12748) );
  OAI21_X1 U8852 ( .B1(n12720), .B2(n6833), .A(n6831), .ZN(n15143) );
  NAND2_X1 U8853 ( .A1(n14961), .A2(n15801), .ZN(n12755) );
  AND2_X1 U8854 ( .A1(n15142), .A2(n12745), .ZN(n15119) );
  NAND2_X1 U8855 ( .A1(n15139), .A2(n7942), .ZN(n12745) );
  NAND2_X1 U8856 ( .A1(n15159), .A2(n14866), .ZN(n12759) );
  NAND2_X1 U8857 ( .A1(n10504), .A2(n10503), .ZN(n14868) );
  XNOR2_X1 U8858 ( .A(n15373), .B(n14823), .ZN(n15158) );
  AND2_X1 U8859 ( .A1(n9184), .A2(n10488), .ZN(n15174) );
  NAND2_X1 U8860 ( .A1(n9122), .A2(n9121), .ZN(n15168) );
  NAND2_X1 U8861 ( .A1(n15201), .A2(n15200), .ZN(n15199) );
  AND2_X1 U8862 ( .A1(n7949), .A2(n7120), .ZN(n15208) );
  AND3_X1 U8863 ( .A1(n6531), .A2(n7121), .A3(n15214), .ZN(n7120) );
  INV_X1 U8864 ( .A(n7122), .ZN(n7121) );
  NOR2_X1 U8865 ( .A1(n15222), .A2(n7705), .ZN(n7704) );
  INV_X1 U8866 ( .A(n9170), .ZN(n7705) );
  NAND2_X1 U8867 ( .A1(n7949), .A2(n8033), .ZN(n15225) );
  NAND2_X1 U8868 ( .A1(n8033), .A2(n7951), .ZN(n15238) );
  AND2_X1 U8869 ( .A1(n8033), .A2(n15421), .ZN(n15251) );
  NOR2_X1 U8870 ( .A1(n15326), .A2(n15325), .ZN(n15328) );
  NAND2_X1 U8871 ( .A1(n7249), .A2(n7248), .ZN(n15326) );
  INV_X1 U8872 ( .A(n12332), .ZN(n7249) );
  AND2_X1 U8873 ( .A1(n14766), .A2(n14758), .ZN(n14937) );
  INV_X1 U8874 ( .A(n14937), .ZN(n12266) );
  NAND2_X1 U8875 ( .A1(n6747), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n8857) );
  INV_X1 U8876 ( .A(n8836), .ZN(n6747) );
  INV_X1 U8877 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n8856) );
  INV_X1 U8878 ( .A(n7321), .ZN(n8877) );
  AND4_X1 U8879 ( .A1(n15805), .A2(n7358), .A3(n11909), .A4(n7119), .ZN(n12203) );
  AND2_X1 U8880 ( .A1(n12203), .A2(n14753), .ZN(n12272) );
  NAND2_X1 U8881 ( .A1(n11909), .A2(n15805), .ZN(n12254) );
  OR2_X1 U8882 ( .A1(n8812), .A2(n8811), .ZN(n8814) );
  NAND2_X1 U8883 ( .A1(n6748), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n8836) );
  INV_X1 U8884 ( .A(n8814), .ZN(n6748) );
  AND4_X1 U8885 ( .A1(n8805), .A2(n8804), .A3(n8803), .A4(n8802), .ZN(n14513)
         );
  INV_X1 U8886 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n9414) );
  OR2_X1 U8887 ( .A1(n8779), .A2(n9414), .ZN(n8812) );
  NAND2_X1 U8888 ( .A1(n8761), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n8779) );
  INV_X1 U8889 ( .A(n8762), .ZN(n8761) );
  CLKBUF_X1 U8890 ( .A(n11853), .Z(n11854) );
  NAND2_X1 U8891 ( .A1(n8728), .A2(n6838), .ZN(n6837) );
  NAND2_X1 U8892 ( .A1(n8029), .A2(n8770), .ZN(n11848) );
  AND4_X1 U8893 ( .A1(n8784), .A2(n8783), .A3(n8782), .A4(n8781), .ZN(n14550)
         );
  NAND2_X1 U8894 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .ZN(n8732) );
  NAND2_X1 U8895 ( .A1(n8730), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n8762) );
  INV_X1 U8896 ( .A(n8732), .ZN(n8730) );
  NAND2_X1 U8897 ( .A1(n11281), .A2(n8728), .ZN(n11742) );
  NAND2_X1 U8898 ( .A1(n11512), .A2(n11283), .ZN(n11733) );
  CLKBUF_X1 U8899 ( .A(n11279), .Z(n11280) );
  NAND2_X1 U8900 ( .A1(n7361), .A2(n14699), .ZN(n11646) );
  INV_X1 U8901 ( .A(n11387), .ZN(n15135) );
  OR2_X1 U8902 ( .A1(n14834), .A2(n11692), .ZN(n8690) );
  CLKBUF_X1 U8903 ( .A(n11372), .Z(n11373) );
  NAND2_X1 U8904 ( .A1(n7995), .A2(n15807), .ZN(n7994) );
  XNOR2_X1 U8905 ( .A(n7996), .B(n9174), .ZN(n7995) );
  NAND2_X1 U8906 ( .A1(n9113), .A2(n12705), .ZN(n7996) );
  NAND2_X1 U8907 ( .A1(n7239), .A2(n7238), .ZN(n7237) );
  AND2_X1 U8908 ( .A1(n9964), .A2(n9963), .ZN(n9965) );
  NOR2_X1 U8909 ( .A1(n9959), .A2(n9958), .ZN(n7238) );
  XNOR2_X1 U8910 ( .A(n10052), .B(n10051), .ZN(n14842) );
  XNOR2_X1 U8911 ( .A(n9972), .B(n9971), .ZN(n14861) );
  NAND2_X1 U8912 ( .A1(n7174), .A2(n9952), .ZN(n9972) );
  NAND2_X1 U8913 ( .A1(n7180), .A2(n7175), .ZN(n7174) );
  NOR2_X1 U8914 ( .A1(n7179), .A2(n9950), .ZN(n7175) );
  NAND2_X1 U8915 ( .A1(n7180), .A2(n7920), .ZN(n9951) );
  INV_X1 U8916 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n8641) );
  XNOR2_X1 U8917 ( .A(n10004), .B(n10003), .ZN(n14464) );
  NAND2_X1 U8918 ( .A1(n7163), .A2(n10028), .ZN(n7172) );
  NAND2_X1 U8919 ( .A1(n7168), .A2(n10028), .ZN(n7165) );
  XNOR2_X1 U8920 ( .A(n9062), .B(n9083), .ZN(n11961) );
  AND2_X1 U8921 ( .A1(n8975), .A2(n8993), .ZN(n15059) );
  INV_X1 U8922 ( .A(n8938), .ZN(n8939) );
  NAND2_X1 U8923 ( .A1(n7155), .A2(n8720), .ZN(n8740) );
  XNOR2_X1 U8924 ( .A(n8718), .B(SI_3_), .ZN(n8717) );
  AND2_X1 U8925 ( .A1(n7940), .A2(n15717), .ZN(n8704) );
  AND2_X1 U8926 ( .A1(n7374), .A2(P3_ADDR_REG_0__SCAN_IN), .ZN(n15587) );
  INV_X1 U8927 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n7374) );
  XNOR2_X1 U8928 ( .A(n15561), .B(P3_ADDR_REG_3__SCAN_IN), .ZN(n15592) );
  XNOR2_X1 U8929 ( .A(n15580), .B(n15562), .ZN(n15582) );
  OAI21_X1 U8930 ( .B1(n15976), .B2(P2_ADDR_REG_5__SCAN_IN), .A(n6604), .ZN(
        n7395) );
  OAI211_X1 U8931 ( .C1(n15612), .C2(n7042), .A(n7040), .B(n7044), .ZN(n15614)
         );
  NAND2_X1 U8932 ( .A1(P3_ADDR_REG_10__SCAN_IN), .A2(n7045), .ZN(n7044) );
  OR2_X1 U8933 ( .A1(n15572), .A2(P1_ADDR_REG_9__SCAN_IN), .ZN(n7042) );
  INV_X1 U8934 ( .A(n15673), .ZN(n7714) );
  NAND2_X1 U8935 ( .A1(n15576), .A2(P1_ADDR_REG_12__SCAN_IN), .ZN(n7511) );
  NAND2_X1 U8936 ( .A1(n7384), .A2(n7387), .ZN(n7344) );
  NAND2_X1 U8937 ( .A1(n7386), .A2(n15697), .ZN(n7385) );
  NAND2_X1 U8938 ( .A1(n7375), .A2(n7388), .ZN(n7377) );
  XNOR2_X1 U8939 ( .A(n15638), .B(P3_ADDR_REG_17__SCAN_IN), .ZN(n15633) );
  INV_X1 U8940 ( .A(n7506), .ZN(n15636) );
  NAND2_X1 U8941 ( .A1(n7726), .A2(n7729), .ZN(n12779) );
  NAND2_X1 U8942 ( .A1(n7725), .A2(n6584), .ZN(n7726) );
  XNOR2_X1 U8943 ( .A(n11216), .B(n12952), .ZN(n11087) );
  INV_X1 U8944 ( .A(n7204), .ZN(n12822) );
  AND2_X1 U8945 ( .A1(n8460), .A2(n8459), .ZN(n13246) );
  AOI21_X1 U8946 ( .B1(n12170), .B2(n12121), .A(n7350), .ZN(n12235) );
  AND4_X1 U8947 ( .A1(n8470), .A2(n8469), .A3(n8468), .A4(n8467), .ZN(n13220)
         );
  INV_X1 U8948 ( .A(n13440), .ZN(n12851) );
  AND2_X1 U8949 ( .A1(n7207), .A2(n7206), .ZN(n7205) );
  NAND2_X1 U8950 ( .A1(n7212), .A2(n7213), .ZN(n7207) );
  NAND2_X1 U8951 ( .A1(n8464), .A2(n8463), .ZN(n13212) );
  AND2_X1 U8952 ( .A1(n11219), .A2(n11218), .ZN(n11224) );
  INV_X1 U8953 ( .A(n12889), .ZN(n7201) );
  INV_X1 U8954 ( .A(n7202), .ZN(n12888) );
  AND2_X1 U8955 ( .A1(n7731), .A2(n7730), .ZN(n12278) );
  INV_X1 U8956 ( .A(n7733), .ZN(n7730) );
  NAND2_X1 U8957 ( .A1(n7725), .A2(n7732), .ZN(n7731) );
  CLKBUF_X1 U8958 ( .A(n11088), .Z(n11085) );
  INV_X1 U8959 ( .A(n13207), .ZN(n13180) );
  NAND2_X1 U8960 ( .A1(n10733), .A2(n10732), .ZN(n12937) );
  NOR2_X1 U8961 ( .A1(n10895), .A2(n10718), .ZN(n12642) );
  XNOR2_X1 U8962 ( .A(n6758), .B(n13128), .ZN(n12635) );
  INV_X1 U8963 ( .A(n13157), .ZN(n12939) );
  INV_X1 U8964 ( .A(n13220), .ZN(n12941) );
  INV_X1 U8965 ( .A(n13246), .ZN(n12942) );
  NAND2_X1 U8966 ( .A1(n12398), .A2(P3_REG1_REG_6__SCAN_IN), .ZN(n6975) );
  INV_X1 U8967 ( .A(P3_ADDR_REG_0__SCAN_IN), .ZN(n15926) );
  AND2_X1 U8968 ( .A1(n10917), .A2(n10916), .ZN(n15913) );
  NAND2_X1 U8969 ( .A1(n10906), .A2(n10907), .ZN(n10940) );
  NAND2_X1 U8970 ( .A1(n6802), .A2(n10963), .ZN(n11068) );
  OAI211_X1 U8971 ( .C1(n10960), .C2(n6798), .A(n6801), .B(n11069), .ZN(n11067) );
  NAND2_X1 U8972 ( .A1(n7658), .A2(n11062), .ZN(n11066) );
  NAND2_X1 U8973 ( .A1(n11064), .A2(n11063), .ZN(n7658) );
  NAND2_X1 U8974 ( .A1(n6895), .A2(n10971), .ZN(n11097) );
  NAND2_X1 U8975 ( .A1(n7654), .A2(n11197), .ZN(n11051) );
  OR2_X1 U8976 ( .A1(n7655), .A2(P3_REG2_REG_7__SCAN_IN), .ZN(n7654) );
  XNOR2_X1 U8977 ( .A(n11193), .B(n11047), .ZN(n11191) );
  OAI211_X1 U8978 ( .C1(n7072), .C2(n7075), .A(n7070), .B(n6601), .ZN(n11585)
         );
  NAND2_X1 U8979 ( .A1(n6786), .A2(n11194), .ZN(n11572) );
  NAND2_X1 U8980 ( .A1(n11191), .A2(P3_REG1_REG_7__SCAN_IN), .ZN(n6786) );
  AOI21_X1 U8981 ( .B1(n11579), .B2(n11578), .A(n11598), .ZN(n11580) );
  AND3_X1 U8982 ( .A1(n6729), .A2(n7408), .A3(n6553), .ZN(n11579) );
  NAND2_X1 U8983 ( .A1(n11580), .A2(P3_REG2_REG_9__SCAN_IN), .ZN(n11601) );
  INV_X1 U8984 ( .A(n7651), .ZN(n12088) );
  OAI21_X1 U8985 ( .B1(n11580), .B2(n11598), .A(n6772), .ZN(n7651) );
  NAND2_X1 U8986 ( .A1(n11597), .A2(n11596), .ZN(n12086) );
  NOR2_X1 U8987 ( .A1(n12983), .A2(n7403), .ZN(n12984) );
  INV_X1 U8988 ( .A(n7404), .ZN(n7403) );
  NAND2_X1 U8989 ( .A1(n13018), .A2(n6781), .ZN(n12994) );
  NAND2_X1 U8990 ( .A1(n12992), .A2(n6782), .ZN(n6781) );
  NOR2_X1 U8991 ( .A1(n12994), .A2(n12995), .ZN(n13021) );
  AND2_X1 U8992 ( .A1(n6815), .A2(n6814), .ZN(n13040) );
  INV_X1 U8993 ( .A(n7095), .ZN(n13047) );
  XNOR2_X1 U8994 ( .A(n13062), .B(n7093), .ZN(n13041) );
  NAND2_X1 U8995 ( .A1(n13041), .A2(P3_REG1_REG_15__SCAN_IN), .ZN(n13064) );
  AOI21_X1 U8996 ( .B1(n13171), .B2(n13336), .A(n7346), .ZN(n13360) );
  NAND2_X1 U8997 ( .A1(n7348), .A2(n7347), .ZN(n7346) );
  NAND2_X1 U8998 ( .A1(n13170), .A2(n13339), .ZN(n7347) );
  OAI21_X1 U8999 ( .B1(n6633), .B2(n8610), .A(n13172), .ZN(n13359) );
  NAND2_X1 U9000 ( .A1(n6845), .A2(n6848), .ZN(n13199) );
  OR2_X1 U9001 ( .A1(n13224), .A2(n6851), .ZN(n6845) );
  NAND2_X1 U9002 ( .A1(n6852), .A2(n6850), .ZN(n13210) );
  AND2_X1 U9003 ( .A1(n6852), .A2(n12596), .ZN(n13211) );
  NAND2_X1 U9004 ( .A1(n13224), .A2(n13219), .ZN(n6852) );
  NAND2_X1 U9005 ( .A1(n8430), .A2(n8429), .ZN(n13381) );
  NAND2_X1 U9006 ( .A1(n7872), .A2(n8325), .ZN(n12214) );
  NAND2_X1 U9007 ( .A1(n12061), .A2(n12060), .ZN(n7872) );
  NAND2_X1 U9008 ( .A1(n7774), .A2(n7777), .ZN(n11950) );
  NAND2_X1 U9009 ( .A1(n11538), .A2(n7778), .ZN(n7774) );
  INV_X1 U9010 ( .A(n13310), .ZN(n13348) );
  INV_X1 U9011 ( .A(P3_REG3_REG_3__SCAN_IN), .ZN(n12350) );
  XNOR2_X1 U9012 ( .A(n7878), .B(n10794), .ZN(n10795) );
  INV_X1 U9013 ( .A(n13321), .ZN(n13345) );
  XNOR2_X1 U9014 ( .A(n7878), .B(n12494), .ZN(n11368) );
  AND2_X1 U9015 ( .A1(n12425), .A2(n12424), .ZN(n13419) );
  INV_X1 U9016 ( .A(n13147), .ZN(n13422) );
  NAND2_X1 U9017 ( .A1(n6855), .A2(n6853), .ZN(n13433) );
  AND2_X1 U9018 ( .A1(n13360), .A2(n6854), .ZN(n6853) );
  NAND2_X1 U9019 ( .A1(n13359), .A2(n13407), .ZN(n6855) );
  NAND2_X1 U9020 ( .A1(n13358), .A2(n15960), .ZN(n6854) );
  NAND2_X1 U9021 ( .A1(n8453), .A2(n8452), .ZN(n13451) );
  NAND2_X1 U9022 ( .A1(n13243), .A2(n8449), .ZN(n7006) );
  OR2_X1 U9023 ( .A1(n13254), .A2(n7765), .ZN(n7758) );
  NAND2_X1 U9024 ( .A1(n7767), .A2(n7769), .ZN(n13241) );
  NAND2_X1 U9025 ( .A1(n13296), .A2(n8605), .ZN(n7767) );
  NAND2_X1 U9026 ( .A1(n7768), .A2(n8605), .ZN(n13259) );
  OR2_X1 U9027 ( .A1(n13254), .A2(n8606), .ZN(n7768) );
  OAI21_X1 U9028 ( .B1(n8384), .B2(n6990), .A(n6988), .ZN(n13288) );
  NAND2_X1 U9029 ( .A1(n6987), .A2(n6991), .ZN(n8035) );
  NAND2_X1 U9030 ( .A1(n8384), .A2(n8383), .ZN(n13302) );
  NAND2_X1 U9031 ( .A1(n8376), .A2(n8375), .ZN(n13481) );
  NAND2_X1 U9032 ( .A1(n8359), .A2(n8358), .ZN(n13491) );
  NAND2_X1 U9033 ( .A1(n6983), .A2(n8351), .ZN(n13326) );
  NAND2_X1 U9034 ( .A1(n13335), .A2(n13334), .ZN(n6983) );
  NAND2_X1 U9035 ( .A1(n8345), .A2(n8344), .ZN(n13494) );
  NAND2_X1 U9036 ( .A1(n7781), .A2(n12484), .ZN(n13333) );
  NAND2_X1 U9037 ( .A1(n11542), .A2(n8276), .ZN(n11790) );
  OAI21_X1 U9038 ( .B1(n11538), .B2(n6587), .A(n8597), .ZN(n11788) );
  AND2_X1 U9039 ( .A1(n8564), .A2(n8563), .ZN(n10709) );
  OR2_X1 U9040 ( .A1(n10621), .A2(P3_D_REG_1__SCAN_IN), .ZN(n8564) );
  NAND2_X1 U9041 ( .A1(n13503), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7783) );
  XNOR2_X1 U9042 ( .A(n12406), .B(n12404), .ZN(n13509) );
  NAND2_X1 U9043 ( .A1(n8128), .A2(n8529), .ZN(n13513) );
  NAND2_X1 U9044 ( .A1(n7820), .A2(n8121), .ZN(n8513) );
  XNOR2_X1 U9045 ( .A(n8560), .B(P3_IR_REG_26__SCAN_IN), .ZN(n13519) );
  OAI21_X1 U9046 ( .B1(n8559), .B2(P3_IR_REG_25__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n8560) );
  XNOR2_X1 U9047 ( .A(n8499), .B(n8498), .ZN(n13520) );
  NAND2_X1 U9048 ( .A1(n7219), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8556) );
  OAI21_X1 U9049 ( .B1(n8451), .B2(n8450), .A(n8112), .ZN(n8472) );
  NAND2_X1 U9050 ( .A1(n8576), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8543) );
  NAND2_X1 U9051 ( .A1(n6858), .A2(n6857), .ZN(n8402) );
  AOI21_X1 U9052 ( .B1(n6541), .B2(n8366), .A(n6706), .ZN(n6857) );
  NAND2_X1 U9053 ( .A1(n8101), .A2(n8100), .ZN(n8386) );
  INV_X1 U9054 ( .A(SI_16_), .ZN(n10892) );
  INV_X1 U9055 ( .A(SI_14_), .ZN(n10662) );
  INV_X1 U9056 ( .A(SI_13_), .ZN(n10660) );
  NAND2_X1 U9057 ( .A1(n8311), .A2(n8089), .ZN(n8327) );
  INV_X1 U9058 ( .A(SI_11_), .ZN(n10633) );
  NAND2_X1 U9059 ( .A1(n6856), .A2(n7847), .ZN(n8294) );
  XNOR2_X1 U9060 ( .A(n8281), .B(n8280), .ZN(n12089) );
  OAI21_X1 U9061 ( .B1(n8264), .B2(n6548), .A(n8085), .ZN(n8278) );
  OAI21_X1 U9062 ( .B1(n8172), .B2(n7833), .A(n7830), .ZN(n8241) );
  NAND2_X1 U9063 ( .A1(n7836), .A2(n8080), .ZN(n8244) );
  NAND2_X1 U9064 ( .A1(n8172), .A2(n8171), .ZN(n7836) );
  NAND2_X1 U9065 ( .A1(n7814), .A2(n8073), .ZN(n8205) );
  NAND2_X1 U9066 ( .A1(n8182), .A2(n8181), .ZN(n7814) );
  NAND2_X1 U9067 ( .A1(n6783), .A2(n6817), .ZN(n6816) );
  INV_X1 U9068 ( .A(P3_IR_REG_31__SCAN_IN), .ZN(n6817) );
  NAND2_X1 U9069 ( .A1(n6933), .A2(n11779), .ZN(n6932) );
  OR2_X1 U9070 ( .A1(n13565), .A2(n13564), .ZN(n7309) );
  NAND2_X1 U9071 ( .A1(n13703), .A2(n12672), .ZN(n13585) );
  NAND2_X1 U9072 ( .A1(n12652), .A2(n12651), .ZN(n13599) );
  NAND2_X1 U9073 ( .A1(n13565), .A2(n13564), .ZN(n13629) );
  NAND2_X1 U9074 ( .A1(n10655), .A2(n9628), .ZN(n7483) );
  NAND2_X1 U9075 ( .A1(n13702), .A2(n13538), .ZN(n13631) );
  NAND2_X1 U9076 ( .A1(n12661), .A2(n12660), .ZN(n13640) );
  NAND2_X1 U9077 ( .A1(n7635), .A2(n13555), .ZN(n13750) );
  NAND2_X1 U9078 ( .A1(n6939), .A2(n7608), .ZN(n13684) );
  AOI21_X1 U9079 ( .B1(n7611), .B2(n7609), .A(n12680), .ZN(n7608) );
  NAND2_X1 U9080 ( .A1(n13651), .A2(n6594), .ZN(n13687) );
  XNOR2_X1 U9081 ( .A(n11709), .B(n11714), .ZN(n11430) );
  NAND2_X1 U9082 ( .A1(n7632), .A2(n7631), .ZN(n12652) );
  INV_X1 U9083 ( .A(n12190), .ZN(n7631) );
  INV_X1 U9084 ( .A(n12191), .ZN(n7632) );
  NAND2_X1 U9085 ( .A1(n13534), .A2(n13696), .ZN(n13702) );
  AND2_X1 U9086 ( .A1(n12697), .A2(n12693), .ZN(n12694) );
  NAND2_X1 U9087 ( .A1(n13704), .A2(n13705), .ZN(n13703) );
  AND2_X1 U9088 ( .A1(n11016), .A2(n11015), .ZN(n13773) );
  NAND2_X1 U9089 ( .A1(n7626), .A2(n7623), .ZN(n13729) );
  NAND2_X1 U9090 ( .A1(n7624), .A2(n12191), .ZN(n7623) );
  INV_X1 U9091 ( .A(n7629), .ZN(n7624) );
  NAND2_X1 U9092 ( .A1(n11772), .A2(n11771), .ZN(n11777) );
  NAND2_X1 U9093 ( .A1(n11772), .A2(n6938), .ZN(n11894) );
  AND2_X1 U9094 ( .A1(n11779), .A2(n11771), .ZN(n6938) );
  INV_X1 U9095 ( .A(n13775), .ZN(n13756) );
  AND2_X1 U9096 ( .A1(n11012), .A2(n14250), .ZN(n13749) );
  AND2_X1 U9097 ( .A1(n13750), .A2(n6592), .ZN(n13761) );
  INV_X1 U9098 ( .A(n13736), .ZN(n13766) );
  INV_X1 U9099 ( .A(n13751), .ZN(n13765) );
  INV_X1 U9100 ( .A(n13749), .ZN(n13777) );
  OR2_X1 U9101 ( .A1(n13983), .A2(n9535), .ZN(n9997) );
  NAND2_X1 U9102 ( .A1(n10015), .A2(n10014), .ZN(n13785) );
  OAI21_X1 U9103 ( .B1(n14010), .B2(n9535), .A(n10037), .ZN(n13786) );
  INV_X1 U9104 ( .A(n10220), .ZN(n13802) );
  NAND2_X1 U9105 ( .A1(n9549), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n7672) );
  NAND4_X1 U9106 ( .A1(n9487), .A2(n9486), .A3(n9485), .A4(n9484), .ZN(n13812)
         );
  NAND2_X1 U9107 ( .A1(n13818), .A2(n13817), .ZN(n13816) );
  NAND2_X1 U9108 ( .A1(n15839), .A2(n15838), .ZN(n15837) );
  NAND2_X1 U9109 ( .A1(n13828), .A2(n13829), .ZN(n13827) );
  NAND2_X1 U9110 ( .A1(n15829), .A2(n6950), .ZN(n13828) );
  OR2_X1 U9111 ( .A1(n10693), .A2(n10694), .ZN(n6950) );
  NAND2_X1 U9112 ( .A1(n13840), .A2(n13841), .ZN(n13839) );
  NAND2_X1 U9113 ( .A1(n13827), .A2(n7571), .ZN(n13840) );
  OR2_X1 U9114 ( .A1(n13830), .A2(n10695), .ZN(n7571) );
  NAND2_X1 U9115 ( .A1(n10676), .A2(n10675), .ZN(n13860) );
  NAND2_X1 U9116 ( .A1(n13839), .A2(n7570), .ZN(n13856) );
  OR2_X1 U9117 ( .A1(n13842), .A2(n10696), .ZN(n7570) );
  NAND2_X1 U9118 ( .A1(n13856), .A2(n13855), .ZN(n13854) );
  NAND2_X1 U9119 ( .A1(n10682), .A2(n10681), .ZN(n13876) );
  AND2_X1 U9120 ( .A1(n6965), .A2(n6964), .ZN(n11173) );
  OR2_X1 U9121 ( .A1(n11181), .A2(n11180), .ZN(n11649) );
  AND2_X1 U9122 ( .A1(n6965), .A2(n6962), .ZN(n11654) );
  AND2_X1 U9123 ( .A1(n11172), .A2(n6964), .ZN(n6962) );
  NOR2_X1 U9124 ( .A1(n11823), .A2(n7569), .ZN(n11824) );
  AND2_X1 U9125 ( .A1(n11826), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n7569) );
  NAND2_X1 U9126 ( .A1(n11824), .A2(n11825), .ZN(n12304) );
  AND2_X1 U9127 ( .A1(n12297), .A2(n12296), .ZN(n15853) );
  NAND2_X1 U9128 ( .A1(n15853), .A2(n15852), .ZN(n15851) );
  XNOR2_X1 U9129 ( .A(n13902), .B(n13893), .ZN(n13886) );
  OAI211_X1 U9130 ( .C1(n13923), .C2(n13921), .A(n13920), .B(n13919), .ZN(
        n13927) );
  AND2_X1 U9131 ( .A1(n13898), .A2(n13897), .ZN(n13923) );
  NAND2_X1 U9132 ( .A1(n13911), .A2(n6725), .ZN(n13913) );
  AND2_X1 U9133 ( .A1(n13913), .A2(n13912), .ZN(n13935) );
  NAND2_X1 U9134 ( .A1(n12385), .A2(n7966), .ZN(n13949) );
  AND2_X1 U9135 ( .A1(n13972), .A2(n13783), .ZN(n13954) );
  NAND2_X1 U9136 ( .A1(n7808), .A2(n7806), .ZN(n14021) );
  NAND2_X1 U9137 ( .A1(n7808), .A2(n10185), .ZN(n14019) );
  INV_X1 U9138 ( .A(n14299), .ZN(n14028) );
  NAND2_X1 U9139 ( .A1(n10184), .A2(n10183), .ZN(n14032) );
  INV_X1 U9140 ( .A(n14325), .ZN(n7668) );
  OAI21_X1 U9141 ( .B1(n14091), .B2(n10237), .A(n10236), .ZN(n14081) );
  NAND2_X1 U9142 ( .A1(n14109), .A2(n10175), .ZN(n14095) );
  NAND2_X1 U9143 ( .A1(n6741), .A2(n10172), .ZN(n14121) );
  NAND2_X1 U9144 ( .A1(n10170), .A2(n10169), .ZN(n14144) );
  NAND2_X1 U9145 ( .A1(n11495), .A2(n9628), .ZN(n7603) );
  NAND2_X1 U9146 ( .A1(n6807), .A2(n6808), .ZN(n12357) );
  NAND2_X1 U9147 ( .A1(n7472), .A2(n7473), .ZN(n14184) );
  OR2_X1 U9148 ( .A1(n14221), .A2(n7475), .ZN(n7472) );
  NAND2_X1 U9149 ( .A1(n14221), .A2(n10163), .ZN(n14203) );
  OR2_X1 U9150 ( .A1(n11330), .A2(n11354), .ZN(n14267) );
  NAND2_X1 U9151 ( .A1(n10159), .A2(n10158), .ZN(n14259) );
  NAND2_X1 U9152 ( .A1(n10624), .A2(n7674), .ZN(n6873) );
  NAND2_X1 U9153 ( .A1(n7437), .A2(n10211), .ZN(n11924) );
  OR2_X1 U9154 ( .A1(n11018), .A2(n15884), .ZN(n14250) );
  NAND2_X1 U9155 ( .A1(n14231), .A2(n11329), .ZN(n14251) );
  OAI21_X1 U9156 ( .B1(n6728), .B2(n11462), .A(n11463), .ZN(n11466) );
  INV_X1 U9157 ( .A(n7671), .ZN(n7670) );
  NAND2_X1 U9158 ( .A1(n7674), .A2(n7673), .ZN(n7669) );
  OAI21_X1 U9159 ( .B1(n9562), .B2(n10573), .A(n7676), .ZN(n7671) );
  INV_X1 U9160 ( .A(n14251), .ZN(n14265) );
  INV_X1 U9161 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n7296) );
  INV_X1 U9162 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n7288) );
  NOR2_X1 U9163 ( .A1(n14293), .A2(n6819), .ZN(n14296) );
  NAND2_X1 U9164 ( .A1(n6821), .A2(n6820), .ZN(n6819) );
  NAND2_X1 U9165 ( .A1(n7352), .A2(n14387), .ZN(n6820) );
  INV_X1 U9166 ( .A(n14148), .ZN(n14431) );
  NOR2_X1 U9167 ( .A1(n15884), .A2(n15872), .ZN(n15879) );
  AND2_X1 U9168 ( .A1(n11021), .A2(n10114), .ZN(n15882) );
  NAND2_X1 U9169 ( .A1(n10273), .A2(n10272), .ZN(n15881) );
  NAND2_X1 U9170 ( .A1(n7988), .A2(n7987), .ZN(n7986) );
  INV_X1 U9171 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n7987) );
  INV_X1 U9172 ( .A(n7989), .ZN(n7988) );
  NAND2_X1 U9173 ( .A1(n9493), .A2(n6564), .ZN(n7790) );
  INV_X1 U9174 ( .A(n10140), .ZN(n12052) );
  NAND2_X1 U9175 ( .A1(n6542), .A2(n6921), .ZN(n9816) );
  INV_X1 U9176 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n11757) );
  INV_X1 U9177 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n11407) );
  INV_X1 U9178 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n11292) );
  INV_X1 U9179 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n11449) );
  INV_X1 U9180 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n11248) );
  INV_X1 U9181 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n10838) );
  INV_X1 U9182 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n10656) );
  INV_X1 U9183 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n10638) );
  INV_X1 U9184 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n10625) );
  INV_X1 U9185 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n10591) );
  INV_X1 U9186 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n10593) );
  INV_X1 U9187 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n9521) );
  INV_X1 U9188 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n10573) );
  NAND2_X1 U9189 ( .A1(n9512), .A2(n14451), .ZN(n6966) );
  NAND2_X1 U9190 ( .A1(n7886), .A2(n10397), .ZN(n14486) );
  NAND2_X1 U9191 ( .A1(n14632), .A2(n14631), .ZN(n7886) );
  INV_X1 U9192 ( .A(n15383), .ZN(n15402) );
  AND2_X1 U9193 ( .A1(n7901), .A2(n7906), .ZN(n14495) );
  AND2_X1 U9194 ( .A1(n7891), .A2(n7889), .ZN(n14519) );
  NAND2_X1 U9195 ( .A1(n10442), .A2(n7891), .ZN(n14520) );
  AOI21_X1 U9196 ( .B1(n7914), .B2(n7910), .A(n7909), .ZN(n7908) );
  INV_X1 U9197 ( .A(n7912), .ZN(n7909) );
  NAND2_X1 U9198 ( .A1(n7898), .A2(n10345), .ZN(n14547) );
  OR2_X1 U9199 ( .A1(n10858), .A2(n10287), .ZN(n10288) );
  NAND2_X1 U9200 ( .A1(n14654), .A2(n10381), .ZN(n14571) );
  AND2_X1 U9201 ( .A1(n10318), .A2(n6597), .ZN(n7137) );
  NAND2_X1 U9202 ( .A1(n7134), .A2(n7133), .ZN(n11546) );
  AND4_X1 U9203 ( .A1(n8818), .A2(n8817), .A3(n8816), .A4(n8815), .ZN(n14618)
         );
  AND4_X1 U9204 ( .A1(n8920), .A2(n8919), .A3(n8918), .A4(n8917), .ZN(n15468)
         );
  NAND2_X1 U9205 ( .A1(n14835), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n7537) );
  NAND2_X1 U9206 ( .A1(n8778), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n7538) );
  AND3_X1 U9207 ( .A1(n9005), .A2(n9004), .A3(n9003), .ZN(n15311) );
  OR2_X1 U9208 ( .A1(n14606), .A2(n15467), .ZN(n14680) );
  INV_X1 U9209 ( .A(n14676), .ZN(n14684) );
  INV_X1 U9210 ( .A(n15709), .ZN(n14686) );
  INV_X1 U9211 ( .A(n14867), .ZN(n14962) );
  NAND2_X1 U9212 ( .A1(n9127), .A2(n9126), .ZN(n15384) );
  OR2_X1 U9213 ( .A1(n14498), .A2(n12754), .ZN(n9112) );
  NAND2_X1 U9214 ( .A1(n9076), .A2(n9075), .ZN(n15240) );
  OR2_X1 U9215 ( .A1(n15227), .A2(n12754), .ZN(n9076) );
  INV_X1 U9216 ( .A(n15401), .ZN(n15419) );
  INV_X1 U9217 ( .A(n14513), .ZN(n15800) );
  INV_X1 U9218 ( .A(n14550), .ZN(n15799) );
  OR2_X1 U9219 ( .A1(n10820), .A2(n10821), .ZN(n7584) );
  NAND2_X1 U9220 ( .A1(n10819), .A2(n7242), .ZN(n10820) );
  NAND2_X1 U9221 ( .A1(n7243), .A2(n10747), .ZN(n7242) );
  NAND2_X1 U9222 ( .A1(n7582), .A2(n6556), .ZN(n11146) );
  AND2_X1 U9223 ( .A1(n7584), .A2(n7583), .ZN(n10842) );
  NAND2_X1 U9224 ( .A1(n11477), .A2(n7593), .ZN(n11479) );
  AND2_X1 U9225 ( .A1(n7592), .A2(n7591), .ZN(n15731) );
  AOI21_X1 U9226 ( .B1(n7587), .B2(n7589), .A(n6712), .ZN(n7585) );
  INV_X1 U9227 ( .A(n15743), .ZN(n7595) );
  AND2_X1 U9228 ( .A1(n10741), .A2(n10632), .ZN(n15722) );
  NAND2_X1 U9229 ( .A1(n7359), .A2(n15447), .ZN(n15345) );
  INV_X1 U9230 ( .A(n14868), .ZN(n14866) );
  OAI21_X1 U9231 ( .B1(n14823), .B2(n12723), .A(n12722), .ZN(n12724) );
  NAND2_X1 U9232 ( .A1(n15139), .A2(n15801), .ZN(n12722) );
  INV_X1 U9233 ( .A(n15194), .ZN(n15386) );
  NAND2_X1 U9234 ( .A1(n15221), .A2(n9077), .ZN(n15207) );
  INV_X1 U9235 ( .A(n7336), .ZN(n9169) );
  NAND2_X1 U9236 ( .A1(n15268), .A2(n9023), .ZN(n15261) );
  INV_X1 U9237 ( .A(n15252), .ZN(n15421) );
  NAND2_X1 U9238 ( .A1(n7695), .A2(n9168), .ZN(n15250) );
  NAND2_X1 U9239 ( .A1(n15266), .A2(n15271), .ZN(n7695) );
  AND2_X1 U9240 ( .A1(n9041), .A2(n9040), .ZN(n15409) );
  AND2_X1 U9241 ( .A1(n9020), .A2(n9019), .ZN(n15435) );
  OAI21_X1 U9242 ( .B1(n7284), .B2(n7692), .A(n7690), .ZN(n15288) );
  NAND2_X1 U9243 ( .A1(n15305), .A2(n8986), .ZN(n15287) );
  NAND2_X1 U9244 ( .A1(n15302), .A2(n15308), .ZN(n15303) );
  NAND2_X1 U9245 ( .A1(n12314), .A2(n9160), .ZN(n12331) );
  CLKBUF_X1 U9246 ( .A(n12328), .Z(n12329) );
  NAND2_X1 U9247 ( .A1(n12311), .A2(n14768), .ZN(n12327) );
  NAND2_X1 U9248 ( .A1(n11247), .A2(n8743), .ZN(n8889) );
  NAND2_X1 U9249 ( .A1(n11112), .A2(n8743), .ZN(n8875) );
  NAND2_X1 U9250 ( .A1(n15497), .A2(n8842), .ZN(n12209) );
  OR2_X1 U9251 ( .A1(n12112), .A2(n14932), .ZN(n15497) );
  NAND2_X1 U9252 ( .A1(n11383), .A2(n11382), .ZN(n15294) );
  INV_X1 U9253 ( .A(n14699), .ZN(n14708) );
  INV_X1 U9254 ( .A(n15294), .ZN(n15331) );
  INV_X1 U9255 ( .A(n15339), .ZN(n15291) );
  NAND2_X1 U9256 ( .A1(n15345), .A2(n7246), .ZN(n15503) );
  INV_X1 U9257 ( .A(n7247), .ZN(n7246) );
  OAI21_X1 U9258 ( .B1(n7360), .B2(n15804), .A(n15346), .ZN(n7247) );
  INV_X1 U9259 ( .A(n15357), .ZN(n7948) );
  NAND2_X1 U9260 ( .A1(n7947), .A2(n15812), .ZN(n6735) );
  NAND2_X1 U9261 ( .A1(n6745), .A2(n6742), .ZN(n15509) );
  AND2_X1 U9262 ( .A1(n15381), .A2(n6743), .ZN(n6742) );
  NAND2_X1 U9263 ( .A1(n15380), .A2(n15812), .ZN(n6745) );
  CLKBUF_X1 U9264 ( .A(n9190), .Z(n15533) );
  XNOR2_X1 U9265 ( .A(n9213), .B(n9212), .ZN(n15542) );
  NAND2_X1 U9266 ( .A1(n7282), .A2(n7281), .ZN(n9210) );
  NAND2_X1 U9267 ( .A1(n9208), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7281) );
  XNOR2_X1 U9268 ( .A(n9101), .B(n9100), .ZN(n12166) );
  XNOR2_X1 U9269 ( .A(n9088), .B(P2_DATAO_REG_22__SCAN_IN), .ZN(n15551) );
  INV_X1 U9270 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n11405) );
  INV_X1 U9271 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n11294) );
  INV_X1 U9272 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n11447) );
  INV_X1 U9273 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n10836) );
  INV_X1 U9274 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n10776) );
  INV_X1 U9275 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n10667) );
  INV_X1 U9276 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n10659) );
  INV_X1 U9277 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n10636) );
  INV_X1 U9278 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n10627) );
  MUX2_X1 U9279 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8755), .S(
        P1_IR_REG_6__SCAN_IN), .Z(n8758) );
  INV_X1 U9280 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n10618) );
  INV_X1 U9281 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n10576) );
  NOR2_X1 U9282 ( .A1(n8673), .A2(n8645), .ZN(n7598) );
  NAND2_X1 U9283 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), .ZN(
        n8672) );
  AOI21_X1 U9284 ( .B1(n15646), .B2(n15591), .A(n15643), .ZN(n15982) );
  XNOR2_X1 U9285 ( .A(n15597), .B(n15598), .ZN(n15976) );
  XNOR2_X1 U9286 ( .A(n7395), .B(P2_ADDR_REG_6__SCAN_IN), .ZN(n15649) );
  INV_X1 U9287 ( .A(n7034), .ZN(n15600) );
  OAI21_X1 U9288 ( .B1(n15596), .B2(P1_ADDR_REG_5__SCAN_IN), .A(n7039), .ZN(
        n7034) );
  INV_X1 U9289 ( .A(n15566), .ZN(n7039) );
  XNOR2_X1 U9290 ( .A(n15605), .B(n15604), .ZN(n15980) );
  OR2_X1 U9291 ( .A1(n15655), .A2(n7716), .ZN(n7715) );
  NAND2_X1 U9292 ( .A1(n7378), .A2(n7376), .ZN(n7389) );
  AND2_X1 U9293 ( .A1(n7385), .A2(n7377), .ZN(n7376) );
  NAND2_X1 U9294 ( .A1(n7344), .A2(n7343), .ZN(n7378) );
  INV_X1 U9295 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n7052) );
  AND2_X1 U9296 ( .A1(n12810), .A2(n6661), .ZN(n7265) );
  NAND2_X1 U9297 ( .A1(n7738), .A2(n7742), .ZN(n7737) );
  NOR2_X1 U9298 ( .A1(n13100), .A2(n13099), .ZN(n6899) );
  NAND2_X1 U9299 ( .A1(n6778), .A2(n15916), .ZN(n6777) );
  NAND2_X1 U9300 ( .A1(n7679), .A2(n6554), .ZN(n6778) );
  NAND2_X1 U9301 ( .A1(n8549), .A2(n13350), .ZN(n7410) );
  INV_X1 U9302 ( .A(n7414), .ZN(n7413) );
  NAND2_X1 U9303 ( .A1(n6650), .A2(n7096), .ZN(P3_U3205) );
  INV_X1 U9304 ( .A(n7097), .ZN(n7096) );
  NAND2_X1 U9305 ( .A1(n7315), .A2(n7314), .ZN(n8622) );
  OAI21_X1 U9306 ( .B1(n13427), .B2(n13406), .A(n8619), .ZN(n8620) );
  NAND2_X1 U9307 ( .A1(n7278), .A2(n7277), .ZN(P3_U3487) );
  INV_X1 U9308 ( .A(n13357), .ZN(n7278) );
  INV_X1 U9309 ( .A(n13356), .ZN(n7277) );
  NOR2_X1 U9310 ( .A1(n7261), .A2(n7260), .ZN(n7259) );
  NOR2_X1 U9311 ( .A1(n15973), .A2(n13363), .ZN(n7260) );
  NOR2_X1 U9312 ( .A1(n13436), .A2(n13403), .ZN(n7261) );
  OR2_X1 U9313 ( .A1(n8549), .A2(n15961), .ZN(n7861) );
  NAND2_X1 U9314 ( .A1(n7280), .A2(n7279), .ZN(P3_U3455) );
  INV_X1 U9315 ( .A(n13432), .ZN(n7280) );
  INV_X1 U9316 ( .A(n13431), .ZN(n7279) );
  NAND2_X1 U9317 ( .A1(n6970), .A2(n6968), .ZN(P3_U3453) );
  NOR2_X1 U9318 ( .A1(n6708), .A2(n6969), .ZN(n6968) );
  OR2_X1 U9319 ( .A1(n13434), .A2(n15961), .ZN(n6970) );
  NOR2_X1 U9320 ( .A1(n15963), .A2(n13435), .ZN(n6969) );
  NOR2_X1 U9321 ( .A1(n10139), .A2(n10117), .ZN(n6902) );
  NAND2_X1 U9322 ( .A1(n7514), .A2(n6560), .ZN(n6903) );
  NAND2_X1 U9323 ( .A1(n10873), .A2(n7565), .ZN(n10876) );
  INV_X1 U9324 ( .A(n7573), .ZN(n6754) );
  NAND2_X1 U9325 ( .A1(n7574), .A2(n11354), .ZN(n6756) );
  AOI21_X1 U9326 ( .B1(n12768), .B2(n15912), .A(n7294), .ZN(n12393) );
  NAND2_X1 U9327 ( .A1(n7297), .A2(n7295), .ZN(n7294) );
  OR2_X1 U9328 ( .A1(n15912), .A2(n7296), .ZN(n7295) );
  OR2_X1 U9329 ( .A1(n15912), .A2(n9977), .ZN(n7687) );
  OR2_X1 U9330 ( .A1(n15912), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n7787) );
  NAND2_X1 U9331 ( .A1(n14405), .A2(n14377), .ZN(n7325) );
  NAND2_X1 U9332 ( .A1(n13995), .A2(n14377), .ZN(n7225) );
  AOI21_X1 U9333 ( .B1(n12768), .B2(n15908), .A(n7286), .ZN(n12770) );
  NAND2_X1 U9334 ( .A1(n7289), .A2(n7287), .ZN(n7286) );
  OR2_X1 U9335 ( .A1(n15908), .A2(n7288), .ZN(n7287) );
  INV_X1 U9336 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n7157) );
  AOI21_X1 U9337 ( .B1(n13972), .B2(n10276), .A(n10275), .ZN(n10277) );
  NAND2_X1 U9338 ( .A1(n14405), .A2(n10276), .ZN(n7327) );
  NAND2_X1 U9339 ( .A1(n13995), .A2(n10276), .ZN(n7224) );
  INV_X1 U9340 ( .A(n7302), .ZN(n7301) );
  OAI21_X1 U9341 ( .B1(n7127), .B2(n14676), .A(n14675), .ZN(n7302) );
  AOI22_X1 U9342 ( .A1(n14952), .A2(n14953), .B1(n14954), .B2(n14955), .ZN(
        n14960) );
  INV_X1 U9343 ( .A(n7577), .ZN(n7576) );
  INV_X1 U9344 ( .A(n7947), .ZN(n8031) );
  NAND2_X1 U9345 ( .A1(n15820), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n7456) );
  NAND2_X1 U9346 ( .A1(n15506), .A2(n15822), .ZN(n7457) );
  NAND2_X1 U9347 ( .A1(n8020), .A2(n8018), .ZN(n8017) );
  NAND2_X1 U9348 ( .A1(n7245), .A2(n7244), .ZN(P1_U3527) );
  NAND2_X1 U9349 ( .A1(n15813), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n7244) );
  NAND2_X1 U9350 ( .A1(n15503), .A2(n15815), .ZN(n7245) );
  NAND2_X1 U9351 ( .A1(n15813), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n7699) );
  NAND2_X1 U9352 ( .A1(n15506), .A2(n15815), .ZN(n7700) );
  NAND2_X1 U9353 ( .A1(n7084), .A2(n7083), .ZN(P1_U3520) );
  NAND2_X1 U9354 ( .A1(n15813), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n7083) );
  OAI21_X1 U9355 ( .B1(n15183), .B2(n9198), .A(n15815), .ZN(n7084) );
  INV_X1 U9356 ( .A(n15615), .ZN(n15677) );
  INV_X1 U9357 ( .A(n7397), .ZN(n15676) );
  NAND2_X1 U9358 ( .A1(n15682), .A2(n15683), .ZN(n15681) );
  NAND2_X1 U9359 ( .A1(n7722), .A2(n7721), .ZN(n15686) );
  AND2_X1 U9360 ( .A1(n7722), .A2(n6670), .ZN(n15685) );
  INV_X1 U9361 ( .A(n7390), .ZN(n15689) );
  INV_X1 U9362 ( .A(n7379), .ZN(n15696) );
  OAI21_X1 U9363 ( .B1(n7383), .B2(P2_ADDR_REG_15__SCAN_IN), .A(n7390), .ZN(
        n7379) );
  NAND2_X1 U9364 ( .A1(n7048), .A2(n7711), .ZN(n7047) );
  NAND2_X1 U9365 ( .A1(n7053), .A2(n7052), .ZN(n7051) );
  INV_X2 U9366 ( .A(n9504), .ZN(n9856) );
  INV_X2 U9367 ( .A(n9856), .ZN(n9947) );
  AND4_X2 U9368 ( .A1(n8996), .A2(n9208), .A3(n8995), .A4(n8641), .ZN(n6537)
         );
  NAND2_X1 U9369 ( .A1(n7355), .A2(n6593), .ZN(n6538) );
  XNOR2_X1 U9370 ( .A(n15133), .B(n15114), .ZN(n6539) );
  OAI21_X1 U9371 ( .B1(n7404), .B2(n6896), .A(n6897), .ZN(n13018) );
  NAND2_X1 U9372 ( .A1(n15849), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n6540) );
  AND2_X1 U9373 ( .A1(n7854), .A2(n6859), .ZN(n6541) );
  AND2_X1 U9374 ( .A1(n7795), .A2(n6785), .ZN(n6542) );
  NAND2_X2 U9375 ( .A1(n9782), .A2(n9781), .ZN(n14435) );
  NAND2_X2 U9376 ( .A1(n7250), .A2(n8976), .ZN(n15444) );
  INV_X2 U9377 ( .A(n9550), .ZN(n9535) );
  BUF_X1 U9378 ( .A(n8197), .Z(n8534) );
  INV_X1 U9379 ( .A(n14945), .ZN(n7703) );
  OR2_X1 U9380 ( .A1(n14824), .A2(n15795), .ZN(n6543) );
  OR2_X1 U9381 ( .A1(n13451), .A2(n12942), .ZN(n6544) );
  NAND2_X1 U9382 ( .A1(n8842), .A2(n7441), .ZN(n14932) );
  AND2_X1 U9383 ( .A1(n9098), .A2(n9077), .ZN(n6545) );
  NOR2_X1 U9384 ( .A1(n10094), .A2(n10093), .ZN(n6546) );
  NAND2_X1 U9385 ( .A1(n13494), .A2(n13327), .ZN(n6547) );
  NAND2_X1 U9386 ( .A1(n7439), .A2(n7438), .ZN(n14186) );
  AND2_X1 U9387 ( .A1(n10665), .A2(P2_DATAO_REG_9__SCAN_IN), .ZN(n6548) );
  OR2_X1 U9388 ( .A1(n14197), .A2(n10225), .ZN(n6549) );
  INV_X1 U9389 ( .A(n10970), .ZN(n7402) );
  INV_X1 U9390 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n9492) );
  NAND2_X1 U9391 ( .A1(n7406), .A2(n6598), .ZN(n11598) );
  AND2_X1 U9392 ( .A1(n10976), .A2(P3_REG1_REG_4__SCAN_IN), .ZN(n6550) );
  XNOR2_X1 U9393 ( .A(n15626), .B(n15625), .ZN(n15690) );
  AND4_X1 U9394 ( .A1(n12382), .A2(n12394), .A3(n14270), .A4(n13783), .ZN(
        n6551) );
  INV_X1 U9395 ( .A(n6851), .ZN(n6850) );
  NAND2_X1 U9396 ( .A1(n8608), .A2(n12596), .ZN(n6851) );
  OR2_X1 U9397 ( .A1(n7079), .A2(n10983), .ZN(n6552) );
  NAND2_X1 U9398 ( .A1(n11577), .A2(P3_REG2_REG_8__SCAN_IN), .ZN(n6553) );
  AND2_X1 U9399 ( .A1(n9197), .A2(n7125), .ZN(n15159) );
  INV_X1 U9400 ( .A(n13808), .ZN(n7805) );
  OR2_X1 U9401 ( .A1(n13107), .A2(n13106), .ZN(n6554) );
  XNOR2_X1 U9402 ( .A(n13993), .B(n13989), .ZN(n6555) );
  OR2_X1 U9403 ( .A1(n10841), .A2(n7583), .ZN(n6556) );
  NAND2_X1 U9404 ( .A1(n13255), .A2(n12474), .ZN(n13289) );
  INV_X1 U9405 ( .A(n13289), .ZN(n6989) );
  AND2_X1 U9406 ( .A1(n9174), .A2(n15144), .ZN(n6557) );
  AND2_X1 U9407 ( .A1(n6640), .A2(n15916), .ZN(n6558) );
  AND2_X1 U9408 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(n6922), .ZN(n6559) );
  INV_X1 U9409 ( .A(n7928), .ZN(n7927) );
  OAI21_X1 U9410 ( .B1(n7930), .B2(n7929), .A(n9080), .ZN(n7928) );
  AND2_X1 U9411 ( .A1(n6546), .A2(n6733), .ZN(n6560) );
  INV_X1 U9412 ( .A(n7128), .ZN(n15172) );
  NOR2_X1 U9413 ( .A1(n15173), .A2(n15379), .ZN(n7128) );
  AND2_X1 U9414 ( .A1(n13491), .A2(n12858), .ZN(n6561) );
  OR2_X1 U9415 ( .A1(n9810), .A2(n9794), .ZN(n6562) );
  AND2_X1 U9416 ( .A1(n9607), .A2(n9606), .ZN(n6563) );
  AND2_X1 U9417 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_27__SCAN_IN), .ZN(
        n6564) );
  INV_X1 U9418 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n10108) );
  INV_X1 U9419 ( .A(n8526), .ZN(n13428) );
  OAI21_X1 U9420 ( .B1(n13513), .B2(n8488), .A(n8138), .ZN(n8526) );
  INV_X1 U9421 ( .A(n11674), .ZN(n6977) );
  INV_X1 U9422 ( .A(n7915), .ZN(n7914) );
  NAND2_X1 U9423 ( .A1(n14580), .A2(n7917), .ZN(n7915) );
  AND2_X1 U9424 ( .A1(n7649), .A2(n12975), .ZN(n12983) );
  AND2_X1 U9425 ( .A1(n13715), .A2(n13717), .ZN(n6565) );
  AND2_X1 U9426 ( .A1(n9634), .A2(n9667), .ZN(n10878) );
  OR2_X1 U9427 ( .A1(n7733), .A2(n6724), .ZN(n6566) );
  AND2_X1 U9428 ( .A1(n14866), .A2(n7942), .ZN(n6567) );
  INV_X1 U9429 ( .A(n9193), .ZN(n9194) );
  XOR2_X1 U9430 ( .A(n14401), .B(n12380), .Z(n6568) );
  NAND2_X1 U9431 ( .A1(n8609), .A2(n12608), .ZN(n13185) );
  AND2_X1 U9432 ( .A1(n9871), .A2(n9870), .ZN(n6569) );
  INV_X1 U9433 ( .A(n8806), .ZN(n8791) );
  XNOR2_X1 U9434 ( .A(n8792), .B(SI_8_), .ZN(n8806) );
  NOR2_X1 U9435 ( .A1(n10877), .A2(n6963), .ZN(n6570) );
  AND2_X1 U9436 ( .A1(n9928), .A2(n7922), .ZN(n6571) );
  INV_X1 U9437 ( .A(n15495), .ZN(n7119) );
  INV_X1 U9438 ( .A(n13995), .ZN(n6888) );
  INV_X1 U9439 ( .A(n6960), .ZN(n6959) );
  NAND2_X1 U9440 ( .A1(n6702), .A2(n6961), .ZN(n6960) );
  AND2_X1 U9441 ( .A1(n7843), .A2(n6722), .ZN(n6572) );
  AND2_X1 U9442 ( .A1(n7944), .A2(n11512), .ZN(n6573) );
  AND2_X2 U9443 ( .A1(n10806), .A2(n10805), .ZN(n15961) );
  INV_X1 U9444 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n6920) );
  OR2_X1 U9445 ( .A1(n10092), .A2(n9856), .ZN(n6574) );
  BUF_X1 U9446 ( .A(n8693), .Z(n14839) );
  INV_X2 U9447 ( .A(n10296), .ZN(n10303) );
  NAND2_X1 U9448 ( .A1(n7299), .A2(n8063), .ZN(n6575) );
  NAND2_X1 U9449 ( .A1(n14664), .A2(n14663), .ZN(n7891) );
  INV_X1 U9450 ( .A(n9440), .ZN(n7106) );
  INV_X1 U9451 ( .A(n13803), .ZN(n7482) );
  XNOR2_X1 U9452 ( .A(n7783), .B(n8057), .ZN(n8061) );
  AND4_X2 U9453 ( .A1(n8055), .A2(n8551), .A3(n8550), .A4(n8554), .ZN(n6576)
         );
  INV_X1 U9454 ( .A(n7675), .ZN(n11296) );
  NAND2_X1 U9455 ( .A1(n7670), .A2(n7669), .ZN(n7675) );
  INV_X1 U9456 ( .A(n15222), .ZN(n9171) );
  INV_X1 U9457 ( .A(n14097), .ZN(n14424) );
  AND2_X1 U9458 ( .A1(n6998), .A2(n6997), .ZN(n6577) );
  OAI211_X1 U9459 ( .C1(n7171), .C2(n7170), .A(n7169), .B(n7166), .ZN(n14295)
         );
  NAND2_X1 U9460 ( .A1(n9169), .A2(n14945), .ZN(n15246) );
  NAND2_X1 U9461 ( .A1(n13251), .A2(n13233), .ZN(n6578) );
  INV_X1 U9462 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n8662) );
  NOR2_X1 U9463 ( .A1(n10186), .A2(n7809), .ZN(n6579) );
  AND2_X1 U9464 ( .A1(n13362), .A2(n13407), .ZN(n6580) );
  NAND2_X1 U9465 ( .A1(n8326), .A2(n8090), .ZN(n6581) );
  AND2_X1 U9466 ( .A1(n8610), .A2(n8609), .ZN(n6582) );
  INV_X1 U9467 ( .A(n10295), .ZN(n10469) );
  INV_X1 U9468 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n9361) );
  INV_X1 U9469 ( .A(n7647), .ZN(n7644) );
  INV_X1 U9470 ( .A(n14018), .ZN(n7647) );
  AND2_X1 U9471 ( .A1(n7409), .A2(P3_REG2_REG_7__SCAN_IN), .ZN(n6583) );
  AND2_X1 U9472 ( .A1(n7732), .A2(n7734), .ZN(n6584) );
  NAND2_X1 U9473 ( .A1(n13264), .A2(n8439), .ZN(n13243) );
  AND2_X1 U9474 ( .A1(n7939), .A2(n7940), .ZN(n8707) );
  OR2_X1 U9475 ( .A1(n15568), .A2(n11195), .ZN(n6585) );
  AND2_X1 U9476 ( .A1(n8461), .A2(n6578), .ZN(n6586) );
  NOR2_X1 U9477 ( .A1(n12551), .A2(n12947), .ZN(n6587) );
  AND2_X1 U9478 ( .A1(n7833), .A2(n7829), .ZN(n6588) );
  XNOR2_X1 U9479 ( .A(n12384), .B(n10136), .ZN(n12382) );
  INV_X1 U9480 ( .A(n12382), .ZN(n13956) );
  NOR2_X1 U9481 ( .A1(n13995), .A2(n13785), .ZN(n6589) );
  XNOR2_X1 U9482 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(P1_DATAO_REG_1__SCAN_IN), 
        .ZN(n8182) );
  AND3_X1 U9483 ( .A1(n9511), .A2(n9510), .A3(n9509), .ZN(n6590) );
  OAI21_X1 U9484 ( .B1(n14654), .B2(n7146), .A(n7144), .ZN(n14632) );
  AND2_X1 U9485 ( .A1(n7429), .A2(n7431), .ZN(n6591) );
  NAND2_X1 U9486 ( .A1(n10253), .A2(n10190), .ZN(n7240) );
  NAND2_X1 U9487 ( .A1(n9967), .A2(n9966), .ZN(n12769) );
  INV_X1 U9488 ( .A(n13972), .ZN(n12394) );
  OAI211_X1 U9489 ( .C1(n10102), .C2(n7953), .A(n7955), .B(n7954), .ZN(n11360)
         );
  INV_X1 U9490 ( .A(n11360), .ZN(n10196) );
  OR2_X1 U9491 ( .A1(n13225), .A2(n12897), .ZN(n12596) );
  NAND3_X1 U9492 ( .A1(n6967), .A2(n9540), .A3(n6966), .ZN(n10574) );
  AND2_X1 U9493 ( .A1(n13556), .A2(n13763), .ZN(n6592) );
  XNOR2_X1 U9494 ( .A(n13995), .B(n13785), .ZN(n13993) );
  NAND2_X1 U9495 ( .A1(n7758), .A2(n7762), .ZN(n13231) );
  NOR2_X1 U9496 ( .A1(n6887), .A2(n14405), .ZN(n6593) );
  INV_X1 U9497 ( .A(n14772), .ZN(n7248) );
  OR2_X1 U9498 ( .A1(n13586), .A2(n13652), .ZN(n6594) );
  XNOR2_X1 U9499 ( .A(n9128), .B(P1_IR_REG_21__SCAN_IN), .ZN(n9193) );
  NAND2_X1 U9500 ( .A1(n8061), .A2(n13510), .ZN(n8139) );
  AND2_X1 U9501 ( .A1(n12382), .A2(n14270), .ZN(n6595) );
  OR2_X1 U9502 ( .A1(n13251), .A2(n13268), .ZN(n6596) );
  NAND2_X1 U9503 ( .A1(n7284), .A2(n9165), .ZN(n15302) );
  AND2_X1 U9504 ( .A1(n10320), .A2(n10319), .ZN(n6597) );
  OR3_X1 U9505 ( .A1(n6689), .A2(n11196), .A3(n11578), .ZN(n6598) );
  XNOR2_X1 U9506 ( .A(n8556), .B(P3_IR_REG_24__SCAN_IN), .ZN(n8561) );
  AND3_X1 U9507 ( .A1(n8928), .A2(n10662), .A3(n8903), .ZN(n6599) );
  NAND2_X1 U9508 ( .A1(n14863), .A2(n14862), .ZN(n15350) );
  INV_X1 U9509 ( .A(n15350), .ZN(n7941) );
  NAND2_X1 U9510 ( .A1(n8649), .A2(n15525), .ZN(n15532) );
  OR2_X1 U9511 ( .A1(n15611), .A2(n15610), .ZN(n6600) );
  OR2_X1 U9512 ( .A1(n10476), .A2(n10477), .ZN(n7919) );
  INV_X1 U9513 ( .A(n7919), .ZN(n7910) );
  OR2_X1 U9514 ( .A1(n11203), .A2(n11204), .ZN(n6601) );
  AND2_X1 U9515 ( .A1(n7847), .A2(n8086), .ZN(n6602) );
  AND2_X1 U9516 ( .A1(n12596), .A2(n12597), .ZN(n13219) );
  INV_X1 U9517 ( .A(n13219), .ZN(n13223) );
  AND2_X1 U9518 ( .A1(n6593), .A2(n12394), .ZN(n6603) );
  OR2_X1 U9519 ( .A1(n15598), .A2(n15597), .ZN(n6604) );
  INV_X1 U9520 ( .A(n15670), .ZN(n7711) );
  AND2_X1 U9521 ( .A1(n10201), .A2(n7974), .ZN(n14114) );
  OR2_X1 U9522 ( .A1(n9089), .A2(n14994), .ZN(n6605) );
  INV_X1 U9523 ( .A(n7745), .ZN(n7744) );
  OAI22_X1 U9524 ( .A1(n12831), .A2(n7749), .B1(n12940), .B2(n12830), .ZN(
        n7745) );
  AND2_X1 U9525 ( .A1(n8604), .A2(n8425), .ZN(n6606) );
  INV_X1 U9526 ( .A(n8611), .ZN(n7773) );
  AND2_X1 U9527 ( .A1(n14443), .A2(n13800), .ZN(n6607) );
  INV_X1 U9528 ( .A(n12521), .ZN(n11303) );
  AND2_X1 U9529 ( .A1(n14414), .A2(n7971), .ZN(n6608) );
  NOR2_X1 U9530 ( .A1(n10922), .A2(n10921), .ZN(n10925) );
  INV_X1 U9531 ( .A(n10983), .ZN(n7080) );
  NAND2_X1 U9532 ( .A1(n14362), .A2(n13576), .ZN(n6609) );
  AND2_X1 U9533 ( .A1(n13153), .A2(n7839), .ZN(n6610) );
  NAND2_X1 U9534 ( .A1(n14865), .A2(n14871), .ZN(n6611) );
  AND2_X1 U9535 ( .A1(n6583), .A2(n11594), .ZN(n6612) );
  INV_X1 U9536 ( .A(n7594), .ZN(n7593) );
  NOR2_X1 U9537 ( .A1(n14771), .A2(n14719), .ZN(n6613) );
  AND2_X1 U9538 ( .A1(n13451), .A2(n13246), .ZN(n12469) );
  INV_X1 U9539 ( .A(P3_IR_REG_20__SCAN_IN), .ZN(n7332) );
  NAND2_X1 U9540 ( .A1(n6953), .A2(n6952), .ZN(n6614) );
  INV_X1 U9541 ( .A(n8497), .ZN(n7869) );
  OR2_X1 U9542 ( .A1(n12635), .A2(n12634), .ZN(n6615) );
  INV_X1 U9543 ( .A(n7779), .ZN(n7778) );
  NAND2_X1 U9544 ( .A1(n8597), .A2(n12560), .ZN(n7779) );
  AND2_X1 U9545 ( .A1(n14733), .A2(n14550), .ZN(n6616) );
  INV_X1 U9546 ( .A(n6993), .ZN(n6992) );
  NAND2_X1 U9547 ( .A1(n8399), .A2(n8383), .ZN(n6993) );
  NAND2_X1 U9548 ( .A1(n14187), .A2(n10224), .ZN(n6617) );
  INV_X1 U9549 ( .A(n7751), .ZN(n7750) );
  NOR2_X1 U9550 ( .A1(n12781), .A2(n12858), .ZN(n7751) );
  INV_X1 U9551 ( .A(n9832), .ZN(n7621) );
  OR2_X1 U9552 ( .A1(n13868), .A2(n10698), .ZN(n6618) );
  NOR2_X1 U9553 ( .A1(n14197), .A2(n13799), .ZN(n6619) );
  INV_X1 U9554 ( .A(n14823), .ZN(n14963) );
  INV_X1 U9555 ( .A(n12384), .ZN(n13962) );
  NAND2_X1 U9556 ( .A1(n9974), .A2(n9973), .ZN(n12384) );
  AND2_X1 U9557 ( .A1(n11849), .A2(n14725), .ZN(n6620) );
  AND2_X1 U9558 ( .A1(n6918), .A2(n6917), .ZN(n6621) );
  NAND2_X1 U9559 ( .A1(n11148), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n6622) );
  NOR2_X1 U9560 ( .A1(n10841), .A2(n10821), .ZN(n6623) );
  NAND2_X1 U9561 ( .A1(n8792), .A2(SI_8_), .ZN(n8793) );
  INV_X1 U9562 ( .A(n8793), .ZN(n7191) );
  INV_X1 U9563 ( .A(n7709), .ZN(n7708) );
  AND2_X1 U9564 ( .A1(n7710), .A2(n12737), .ZN(n7709) );
  AND2_X1 U9565 ( .A1(n6586), .A2(n7002), .ZN(n6624) );
  INV_X1 U9566 ( .A(n7542), .ZN(n7541) );
  NAND2_X1 U9567 ( .A1(n14810), .A2(n14809), .ZN(n7542) );
  AND2_X1 U9568 ( .A1(SI_0_), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n6625) );
  AND2_X1 U9569 ( .A1(n8741), .A2(SI_4_), .ZN(n6626) );
  NOR2_X1 U9570 ( .A1(n14295), .A2(n13786), .ZN(n6627) );
  NOR2_X1 U9571 ( .A1(n15438), .A2(n15274), .ZN(n6628) );
  NOR2_X1 U9572 ( .A1(n7226), .A2(n15428), .ZN(n6629) );
  NOR2_X1 U9573 ( .A1(n15405), .A2(n15240), .ZN(n6630) );
  NOR2_X1 U9574 ( .A1(n12218), .A2(n12238), .ZN(n6631) );
  AND2_X1 U9575 ( .A1(n10976), .A2(P3_REG2_REG_4__SCAN_IN), .ZN(n6632) );
  INV_X1 U9576 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n7959) );
  INV_X1 U9577 ( .A(n11600), .ZN(n7652) );
  INV_X1 U9578 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n8800) );
  AND2_X1 U9579 ( .A1(n13182), .A2(n8609), .ZN(n6633) );
  AND2_X1 U9580 ( .A1(n15438), .A2(n15274), .ZN(n6634) );
  INV_X1 U9581 ( .A(n7145), .ZN(n7144) );
  OAI21_X1 U9582 ( .B1(n7146), .B2(n10381), .A(n10389), .ZN(n7145) );
  NAND2_X1 U9583 ( .A1(n12785), .A2(n13303), .ZN(n7351) );
  AND2_X1 U9584 ( .A1(n14912), .A2(n14914), .ZN(n6635) );
  INV_X1 U9585 ( .A(n8986), .ZN(n8004) );
  INV_X1 U9586 ( .A(n7749), .ZN(n7748) );
  NAND2_X1 U9587 ( .A1(n13196), .A2(n12805), .ZN(n7749) );
  AND2_X1 U9588 ( .A1(n8774), .A2(SI_6_), .ZN(n6636) );
  AND2_X1 U9589 ( .A1(n7545), .A2(n7542), .ZN(n6637) );
  AND2_X1 U9590 ( .A1(n8845), .A2(SI_10_), .ZN(n6638) );
  AND2_X1 U9591 ( .A1(n11805), .A2(n12948), .ZN(n6639) );
  AND2_X1 U9592 ( .A1(n13107), .A2(n13106), .ZN(n6640) );
  AND2_X1 U9593 ( .A1(n14299), .A2(n13787), .ZN(n6641) );
  NAND2_X1 U9594 ( .A1(n9795), .A2(n7982), .ZN(n6642) );
  AND2_X1 U9595 ( .A1(n13550), .A2(n13549), .ZN(n6643) );
  NAND2_X1 U9596 ( .A1(n13559), .A2(n13558), .ZN(n6644) );
  NAND2_X1 U9597 ( .A1(P3_ADDR_REG_3__SCAN_IN), .A2(n15561), .ZN(n6645) );
  INV_X1 U9598 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n9512) );
  AND2_X1 U9599 ( .A1(n12464), .A2(n12463), .ZN(n13198) );
  INV_X1 U9600 ( .A(P3_IR_REG_18__SCAN_IN), .ZN(n7857) );
  OR2_X1 U9601 ( .A1(n14320), .A2(n10240), .ZN(n6646) );
  AND2_X1 U9602 ( .A1(n9949), .A2(n9948), .ZN(n6647) );
  AND2_X1 U9603 ( .A1(n12708), .A2(n6840), .ZN(n6648) );
  AND2_X1 U9604 ( .A1(n8253), .A2(n6976), .ZN(n6649) );
  AND2_X1 U9605 ( .A1(n13162), .A2(n13161), .ZN(n6650) );
  INV_X1 U9606 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n10589) );
  NAND2_X1 U9607 ( .A1(n12122), .A2(n12216), .ZN(n6651) );
  AND2_X1 U9609 ( .A1(n7911), .A2(n7907), .ZN(n6653) );
  AND2_X1 U9610 ( .A1(n10774), .A2(P2_DATAO_REG_10__SCAN_IN), .ZN(n6654) );
  NAND2_X1 U9611 ( .A1(n15368), .A2(n15367), .ZN(n6655) );
  NAND2_X1 U9612 ( .A1(n12776), .A2(n12777), .ZN(n6656) );
  INV_X1 U9613 ( .A(n8003), .ZN(n8002) );
  NAND2_X1 U9614 ( .A1(n7251), .A2(n14779), .ZN(n8003) );
  OR2_X1 U9615 ( .A1(n11036), .A2(n11442), .ZN(n6657) );
  AND2_X1 U9616 ( .A1(n10219), .A2(n14223), .ZN(n6658) );
  INV_X1 U9617 ( .A(n10397), .ZN(n7887) );
  AND2_X1 U9618 ( .A1(n13286), .A2(n12475), .ZN(n13301) );
  NAND2_X1 U9619 ( .A1(n12375), .A2(n10118), .ZN(n10189) );
  AND2_X1 U9620 ( .A1(n6658), .A2(n6878), .ZN(n6659) );
  NAND2_X1 U9621 ( .A1(n7780), .A2(n11787), .ZN(n6660) );
  INV_X1 U9622 ( .A(n14730), .ZN(n7015) );
  INV_X1 U9623 ( .A(n6544), .ZN(n7004) );
  INV_X1 U9624 ( .A(n15214), .ZN(n15395) );
  INV_X1 U9625 ( .A(n9872), .ZN(n7526) );
  INV_X1 U9626 ( .A(n7480), .ZN(n7479) );
  OR2_X1 U9627 ( .A1(n10174), .A2(n7481), .ZN(n7480) );
  INV_X1 U9628 ( .A(P3_ADDR_REG_1__SCAN_IN), .ZN(n15557) );
  NAND2_X1 U9629 ( .A1(n14857), .A2(n14856), .ZN(n15344) );
  INV_X1 U9630 ( .A(n15344), .ZN(n7360) );
  OR2_X1 U9631 ( .A1(n13175), .A2(n12937), .ZN(n6661) );
  NAND2_X1 U9632 ( .A1(n12744), .A2(n12743), .ZN(n15361) );
  INV_X1 U9633 ( .A(n15361), .ZN(n7942) );
  INV_X1 U9634 ( .A(n8604), .ZN(n6861) );
  INV_X1 U9635 ( .A(n14776), .ZN(n7552) );
  XNOR2_X1 U9636 ( .A(n14671), .B(n14670), .ZN(n6662) );
  INV_X1 U9637 ( .A(n6834), .ZN(n11212) );
  INV_X1 U9638 ( .A(n14934), .ZN(n7455) );
  NAND2_X2 U9639 ( .A1(n8889), .A2(n8888), .ZN(n15471) );
  INV_X1 U9640 ( .A(n13993), .ZN(n7420) );
  AND2_X1 U9641 ( .A1(n7830), .A2(n7829), .ZN(n6663) );
  AND2_X1 U9642 ( .A1(n6584), .A2(n12778), .ZN(n6664) );
  OR2_X1 U9643 ( .A1(n14341), .A2(n13794), .ZN(n10173) );
  OR2_X1 U9644 ( .A1(n14948), .A2(n6736), .ZN(n6665) );
  AND2_X1 U9645 ( .A1(n7924), .A2(n7186), .ZN(n6666) );
  AND2_X1 U9646 ( .A1(n7006), .A2(n6578), .ZN(n6667) );
  AND2_X1 U9647 ( .A1(n7135), .A2(n11548), .ZN(n6668) );
  INV_X1 U9648 ( .A(n15405), .ZN(n7950) );
  INV_X1 U9649 ( .A(n15901), .ZN(n12009) );
  AND2_X1 U9650 ( .A1(n9598), .A2(n6873), .ZN(n15901) );
  INV_X1 U9651 ( .A(n14476), .ZN(n7953) );
  AND2_X1 U9652 ( .A1(n8590), .A2(n12510), .ZN(n6669) );
  NOR2_X1 U9653 ( .A1(n15687), .A2(n7720), .ZN(n6670) );
  AND2_X1 U9654 ( .A1(n7918), .A2(n10502), .ZN(n6671) );
  NOR2_X1 U9655 ( .A1(n10144), .A2(n10143), .ZN(n6672) );
  AND2_X1 U9656 ( .A1(n7497), .A2(n7499), .ZN(n6673) );
  AND2_X1 U9657 ( .A1(n7100), .A2(n8611), .ZN(n6674) );
  XNOR2_X1 U9658 ( .A(n15344), .B(n15106), .ZN(n14899) );
  INV_X1 U9659 ( .A(n8786), .ZN(n8787) );
  XNOR2_X1 U9660 ( .A(n8789), .B(SI_7_), .ZN(n8786) );
  AND2_X1 U9661 ( .A1(n9547), .A2(n7520), .ZN(n6675) );
  AND2_X1 U9662 ( .A1(n12746), .A2(n12711), .ZN(n14947) );
  INV_X1 U9663 ( .A(n14947), .ZN(n7710) );
  NAND2_X1 U9664 ( .A1(n14792), .A2(n14791), .ZN(n6676) );
  AND2_X1 U9665 ( .A1(n8608), .A2(n6766), .ZN(n6677) );
  NAND2_X1 U9666 ( .A1(n11415), .A2(n11414), .ZN(n6678) );
  AND2_X1 U9667 ( .A1(n10188), .A2(n10129), .ZN(n13980) );
  INV_X1 U9668 ( .A(n13980), .ZN(n7933) );
  AND2_X1 U9669 ( .A1(n15259), .A2(n9042), .ZN(n6679) );
  AND2_X1 U9670 ( .A1(n14790), .A2(n14789), .ZN(n6680) );
  AND2_X1 U9671 ( .A1(n12606), .A2(n12605), .ZN(n6681) );
  AND2_X1 U9672 ( .A1(n10072), .A2(n7293), .ZN(n6682) );
  OR2_X1 U9673 ( .A1(n14790), .A2(n14789), .ZN(n6683) );
  AND2_X1 U9674 ( .A1(n6556), .A2(n6622), .ZN(n6684) );
  OR2_X1 U9675 ( .A1(n14743), .A2(n14745), .ZN(n6685) );
  AND2_X1 U9676 ( .A1(n8022), .A2(n8021), .ZN(n6686) );
  AND2_X1 U9677 ( .A1(n9161), .A2(n9160), .ZN(n6687) );
  AND2_X1 U9678 ( .A1(n6567), .A2(n7941), .ZN(n6688) );
  NAND2_X1 U9679 ( .A1(n7401), .A2(n11192), .ZN(n6689) );
  AND2_X1 U9680 ( .A1(n12787), .A2(n13290), .ZN(n6690) );
  INV_X1 U9681 ( .A(n7544), .ZN(n7543) );
  NOR2_X1 U9682 ( .A1(n14810), .A2(n14809), .ZN(n7544) );
  INV_X1 U9683 ( .A(n7078), .ZN(n7074) );
  AND2_X1 U9684 ( .A1(n7080), .A2(n11102), .ZN(n7078) );
  AND2_X1 U9685 ( .A1(n13956), .A2(n7430), .ZN(n6691) );
  NAND2_X1 U9686 ( .A1(n10776), .A2(P1_DATAO_REG_10__SCAN_IN), .ZN(n6692) );
  NAND2_X1 U9687 ( .A1(n7352), .A2(n13752), .ZN(n6693) );
  AND2_X1 U9688 ( .A1(n6918), .A2(P2_IR_REG_19__SCAN_IN), .ZN(n6694) );
  AND2_X1 U9689 ( .A1(n14451), .A2(n7959), .ZN(n6695) );
  AND2_X1 U9690 ( .A1(n6646), .A2(n7667), .ZN(n6696) );
  NAND2_X1 U9691 ( .A1(n12833), .A2(n7746), .ZN(n6697) );
  INV_X1 U9692 ( .A(P3_IR_REG_29__SCAN_IN), .ZN(n7782) );
  INV_X1 U9693 ( .A(P3_IR_REG_27__SCAN_IN), .ZN(n7494) );
  INV_X1 U9694 ( .A(n6885), .ZN(n10203) );
  NAND2_X1 U9695 ( .A1(n7973), .A2(n14114), .ZN(n6885) );
  NAND2_X1 U9696 ( .A1(n10090), .A2(n10089), .ZN(n6698) );
  OR2_X1 U9697 ( .A1(n7526), .A2(n6569), .ZN(n6699) );
  INV_X1 U9698 ( .A(n14813), .ZN(n7545) );
  AND4_X1 U9699 ( .A1(n8737), .A2(n8736), .A3(n8735), .A4(n8734), .ZN(n11849)
         );
  AND2_X1 U9700 ( .A1(SI_0_), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n6700) );
  INV_X1 U9702 ( .A(P3_IR_REG_19__SCAN_IN), .ZN(n7329) );
  AND2_X1 U9703 ( .A1(n7972), .A2(n7959), .ZN(n6701) );
  NAND3_X1 U9705 ( .A1(n7419), .A2(n7856), .A3(n8176), .ZN(n11438) );
  INV_X1 U9706 ( .A(n13696), .ZN(n6945) );
  AND2_X1 U9708 ( .A1(n12008), .A2(n12071), .ZN(n12024) );
  NAND2_X1 U9709 ( .A1(n10107), .A2(n10108), .ZN(n10104) );
  INV_X1 U9710 ( .A(n7331), .ZN(n12632) );
  NAND2_X1 U9711 ( .A1(n13128), .A2(n11753), .ZN(n7331) );
  INV_X1 U9712 ( .A(n13352), .ZN(n13324) );
  OR2_X1 U9713 ( .A1(n12305), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n6702) );
  INV_X1 U9714 ( .A(n7308), .ZN(n9029) );
  AND2_X1 U9715 ( .A1(n7117), .A2(n7116), .ZN(n6703) );
  OAI21_X1 U9716 ( .B1(n13335), .B2(n6980), .A(n6978), .ZN(n13312) );
  NAND2_X1 U9717 ( .A1(n8593), .A2(n8592), .ZN(n11300) );
  AND2_X1 U9718 ( .A1(n9971), .A2(n7176), .ZN(n6704) );
  INV_X1 U9719 ( .A(P3_ADDR_REG_4__SCAN_IN), .ZN(n15562) );
  INV_X1 U9720 ( .A(n10028), .ZN(n7173) );
  AND3_X1 U9721 ( .A1(n7977), .A2(n7975), .A3(n7976), .ZN(n10095) );
  NAND2_X1 U9722 ( .A1(n7357), .A2(n7795), .ZN(n7653) );
  XNOR2_X1 U9723 ( .A(n15612), .B(P1_ADDR_REG_9__SCAN_IN), .ZN(n15651) );
  AND2_X1 U9724 ( .A1(P2_REG3_REG_11__SCAN_IN), .A2(P2_REG3_REG_12__SCAN_IN), 
        .ZN(n6705) );
  INV_X1 U9725 ( .A(n7686), .ZN(n7685) );
  NOR2_X1 U9726 ( .A1(n13054), .A2(n7093), .ZN(n7686) );
  AND2_X1 U9727 ( .A1(n11407), .A2(P2_DATAO_REG_17__SCAN_IN), .ZN(n6706) );
  AND2_X1 U9728 ( .A1(n7898), .A2(n7896), .ZN(n6707) );
  NOR2_X1 U9729 ( .A1(n13436), .A2(n13493), .ZN(n6708) );
  NOR2_X1 U9730 ( .A1(n13469), .A2(n13303), .ZN(n6709) );
  NOR2_X1 U9731 ( .A1(n10053), .A2(n14470), .ZN(n6710) );
  OR2_X1 U9732 ( .A1(n13969), .A2(n14250), .ZN(n6711) );
  NOR2_X1 U9733 ( .A1(n15732), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n6712) );
  INV_X1 U9734 ( .A(n12932), .ZN(n13328) );
  AND3_X1 U9735 ( .A1(n8381), .A2(n8380), .A3(n8379), .ZN(n12932) );
  INV_X1 U9736 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n10665) );
  NAND2_X1 U9737 ( .A1(n15567), .A2(P3_ADDR_REG_6__SCAN_IN), .ZN(n6713) );
  AND2_X1 U9738 ( .A1(n7394), .A2(n7391), .ZN(n6714) );
  OR2_X1 U9739 ( .A1(n13032), .A2(n13029), .ZN(n6715) );
  AND2_X1 U9740 ( .A1(n6547), .A2(n12484), .ZN(n6716) );
  AND2_X1 U9741 ( .A1(n7439), .A2(n10223), .ZN(n6717) );
  OR2_X1 U9742 ( .A1(n14008), .A2(n13749), .ZN(n6718) );
  OR2_X1 U9743 ( .A1(n7686), .A2(n13330), .ZN(n6719) );
  AND2_X1 U9744 ( .A1(n12789), .A2(n13276), .ZN(n6720) );
  NOR2_X1 U9745 ( .A1(n12998), .A2(n12993), .ZN(n7638) );
  AND2_X1 U9746 ( .A1(n6958), .A2(n6540), .ZN(n6721) );
  INV_X1 U9747 ( .A(n7130), .ZN(n15447) );
  NAND2_X1 U9748 ( .A1(n14689), .A2(n9140), .ZN(n15807) );
  INV_X1 U9749 ( .A(n15973), .ZN(n15970) );
  NAND2_X1 U9750 ( .A1(n8799), .A2(n8798), .ZN(n14742) );
  INV_X1 U9751 ( .A(n14742), .ZN(n7358) );
  NAND2_X1 U9752 ( .A1(n10194), .A2(n14164), .ZN(n11003) );
  OR2_X1 U9753 ( .A1(n11282), .A2(n14926), .ZN(n11281) );
  AOI21_X1 U9754 ( .B1(n11599), .B2(n6773), .A(n11600), .ZN(n6772) );
  OR2_X1 U9755 ( .A1(n12164), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n6722) );
  NAND3_X1 U9756 ( .A1(n8254), .A2(n6649), .A3(n6975), .ZN(n12950) );
  INV_X1 U9757 ( .A(n12950), .ZN(n6974) );
  INV_X1 U9758 ( .A(n13334), .ZN(n6979) );
  INV_X1 U9759 ( .A(n12922), .ZN(n12924) );
  AND2_X1 U9760 ( .A1(n13936), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n6723) );
  INV_X1 U9761 ( .A(n11645), .ZN(n7361) );
  AND2_X1 U9762 ( .A1(n12123), .A2(n12238), .ZN(n6724) );
  OR2_X1 U9763 ( .A1(n13916), .A2(n14347), .ZN(n6725) );
  NAND2_X1 U9764 ( .A1(n6839), .A2(n14698), .ZN(n11282) );
  AND2_X1 U9765 ( .A1(n15574), .A2(P1_ADDR_REG_11__SCAN_IN), .ZN(n6726) );
  AND2_X1 U9766 ( .A1(n6729), .A2(n7408), .ZN(n6727) );
  NAND2_X1 U9767 ( .A1(n11962), .A2(n14688), .ZN(n7131) );
  INV_X1 U9768 ( .A(n7131), .ZN(n7129) );
  AND2_X1 U9769 ( .A1(n11465), .A2(n11464), .ZN(n6728) );
  INV_X1 U9770 ( .A(SI_22_), .ZN(n7186) );
  OR2_X1 U9771 ( .A1(n6689), .A2(n11196), .ZN(n6729) );
  AND2_X1 U9772 ( .A1(n7061), .A2(n7489), .ZN(n6730) );
  INV_X1 U9773 ( .A(n11771), .ZN(n7633) );
  INV_X1 U9774 ( .A(n7076), .ZN(n7075) );
  NAND2_X1 U9775 ( .A1(n6552), .A2(n11039), .ZN(n7076) );
  AND2_X1 U9776 ( .A1(n6774), .A2(n7402), .ZN(n6731) );
  OR2_X1 U9777 ( .A1(n15820), .A2(n8021), .ZN(n6732) );
  INV_X1 U9778 ( .A(P3_REG3_REG_17__SCAN_IN), .ZN(n7111) );
  INV_X1 U9779 ( .A(P3_REG1_REG_7__SCAN_IN), .ZN(n6789) );
  INV_X1 U9780 ( .A(n11062), .ZN(n7661) );
  INV_X1 U9781 ( .A(n15103), .ZN(n15178) );
  INV_X1 U9782 ( .A(n10822), .ZN(n7243) );
  INV_X1 U9783 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n8995) );
  AND2_X1 U9784 ( .A1(n10101), .A2(n10100), .ZN(n6733) );
  NAND2_X1 U9785 ( .A1(n9503), .A2(n9502), .ZN(n14164) );
  NAND4_X1 U9786 ( .A1(n6984), .A2(n8052), .A3(n6576), .A4(n7231), .ZN(n13503)
         );
  INV_X1 U9787 ( .A(n7388), .ZN(n7387) );
  NOR2_X1 U9788 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P2_ADDR_REG_15__SCAN_IN), 
        .ZN(n7388) );
  INV_X1 U9789 ( .A(n13106), .ZN(n7681) );
  AND2_X1 U9790 ( .A1(n15622), .A2(P1_ADDR_REG_14__SCAN_IN), .ZN(n6734) );
  INV_X1 U9791 ( .A(P3_REG1_REG_1__SCAN_IN), .ZN(n7495) );
  INV_X1 U9792 ( .A(P3_REG3_REG_24__SCAN_IN), .ZN(n7299) );
  INV_X1 U9793 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n7509) );
  INV_X1 U9794 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n7501) );
  INV_X1 U9795 ( .A(P3_REG1_REG_3__SCAN_IN), .ZN(n6803) );
  INV_X1 U9796 ( .A(P3_REG2_REG_1__SCAN_IN), .ZN(n7088) );
  INV_X1 U9797 ( .A(P3_REG2_REG_9__SCAN_IN), .ZN(n6773) );
  OAI22_X1 U9798 ( .A1(n13134), .A2(n13133), .B1(n13132), .B2(n13388), .ZN(
        n13137) );
  AOI21_X1 U9799 ( .B1(n15922), .B2(n13132), .A(n13117), .ZN(n7499) );
  INV_X1 U9800 ( .A(n13132), .ZN(n7334) );
  INV_X1 U9801 ( .A(n13063), .ZN(n7093) );
  NOR2_X1 U9802 ( .A1(n13045), .A2(n13063), .ZN(n7684) );
  NOR2_X1 U9803 ( .A1(n13027), .A2(n7638), .ZN(n6782) );
  OAI21_X1 U9804 ( .B1(n12982), .B2(n7638), .A(n13027), .ZN(n6898) );
  NOR2_X1 U9805 ( .A1(n13350), .A2(n8629), .ZN(n7416) );
  NAND2_X1 U9806 ( .A1(n13089), .A2(n13112), .ZN(n13107) );
  XNOR2_X1 U9807 ( .A(n13102), .B(n13112), .ZN(n13104) );
  NAND2_X1 U9808 ( .A1(n13113), .A2(n13112), .ZN(n7486) );
  NAND3_X1 U9809 ( .A1(n6735), .A2(n15358), .A3(n7948), .ZN(n15505) );
  NAND4_X1 U9810 ( .A1(n15170), .A2(n14899), .A3(n6557), .A4(n6539), .ZN(n6736) );
  NAND2_X1 U9811 ( .A1(n7889), .A2(n8032), .ZN(n7888) );
  NAND2_X1 U9812 ( .A1(n6737), .A2(n8610), .ZN(n12613) );
  NAND2_X1 U9813 ( .A1(n7271), .A2(n12607), .ZN(n6737) );
  INV_X1 U9814 ( .A(n8080), .ZN(n7835) );
  NAND2_X2 U9815 ( .A1(n13515), .A2(n13111), .ZN(n10897) );
  NAND2_X2 U9816 ( .A1(n7490), .A2(n7493), .ZN(n13111) );
  AND2_X1 U9817 ( .A1(n11087), .A2(n11086), .ZN(n6739) );
  INV_X1 U9818 ( .A(n12903), .ZN(n6740) );
  NAND2_X1 U9819 ( .A1(n6818), .A2(n6673), .ZN(n6780) );
  NAND2_X1 U9820 ( .A1(n6779), .A2(n6777), .ZN(P3_U3200) );
  NAND2_X1 U9821 ( .A1(n7266), .A2(n12802), .ZN(n12846) );
  NOR2_X1 U9822 ( .A1(n12887), .A2(n6720), .ZN(n12840) );
  NAND2_X1 U9823 ( .A1(n8487), .A2(n8486), .ZN(n8485) );
  NAND2_X1 U9824 ( .A1(n8079), .A2(n8078), .ZN(n8172) );
  NAND2_X1 U9825 ( .A1(n8111), .A2(n7841), .ZN(n7840) );
  NAND2_X1 U9826 ( .A1(n12625), .A2(n12624), .ZN(n7274) );
  AOI21_X1 U9827 ( .B1(n12867), .B2(n12863), .A(n12865), .ZN(n12904) );
  OAI21_X1 U9828 ( .B1(n8428), .B2(n8107), .A(n8106), .ZN(n8441) );
  XNOR2_X1 U9829 ( .A(n7200), .B(n7199), .ZN(n7198) );
  NAND2_X1 U9830 ( .A1(n8056), .A2(n7857), .ZN(n8553) );
  OAI21_X1 U9831 ( .B1(n7198), .B2(n12922), .A(n7265), .ZN(P3_U3154) );
  NAND2_X1 U9832 ( .A1(n7208), .A2(n7205), .ZN(n12867) );
  OAI21_X1 U9833 ( .B1(n11970), .B2(n11803), .A(n11802), .ZN(n7268) );
  INV_X1 U9834 ( .A(n14287), .ZN(n7326) );
  INV_X1 U9835 ( .A(n14404), .ZN(n7328) );
  NAND2_X1 U9836 ( .A1(n7461), .A2(n10159), .ZN(n14257) );
  OAI21_X2 U9837 ( .B1(n12356), .B2(n10167), .A(n10166), .ZN(n14181) );
  NAND2_X1 U9838 ( .A1(n7463), .A2(n7462), .ZN(n13992) );
  INV_X1 U9839 ( .A(n10175), .ZN(n7800) );
  NAND2_X1 U9840 ( .A1(n7476), .A2(n7796), .ZN(n14063) );
  NAND2_X1 U9841 ( .A1(n12316), .A2(n12315), .ZN(n12313) );
  NOR2_X1 U9842 ( .A1(n14288), .A2(n7227), .ZN(n14406) );
  NAND2_X1 U9843 ( .A1(n14290), .A2(n14396), .ZN(n7229) );
  NAND2_X1 U9844 ( .A1(n15985), .A2(n15986), .ZN(n15589) );
  XNOR2_X1 U9845 ( .A(n15588), .B(P2_ADDR_REG_1__SCAN_IN), .ZN(n15985) );
  INV_X1 U9846 ( .A(n15691), .ZN(n7343) );
  XNOR2_X1 U9847 ( .A(n7056), .B(n15663), .ZN(n15662) );
  NAND2_X1 U9848 ( .A1(n15975), .A2(n15974), .ZN(n15594) );
  OAI21_X2 U9849 ( .B1(n7394), .B2(n7393), .A(n7392), .ZN(n15657) );
  OAI21_X1 U9850 ( .B1(n14827), .B2(n14826), .A(n14825), .ZN(n14828) );
  NAND3_X1 U9852 ( .A1(n9116), .A2(n9114), .A3(n9115), .ZN(n9120) );
  INV_X1 U9853 ( .A(n7691), .ZN(n7690) );
  XNOR2_X1 U9854 ( .A(n10315), .B(n10314), .ZN(n15705) );
  AOI21_X2 U9855 ( .B1(n14579), .B2(n14580), .A(n7149), .ZN(n7148) );
  NAND2_X1 U9856 ( .A1(n7283), .A2(P1_IR_REG_24__SCAN_IN), .ZN(n7282) );
  NAND2_X1 U9857 ( .A1(n7138), .A2(n11547), .ZN(n11623) );
  NAND4_X1 U9858 ( .A1(n6746), .A2(n14545), .A3(n14544), .A4(n14546), .ZN(
        P1_U3220) );
  NAND3_X1 U9859 ( .A1(n14534), .A2(n14542), .A3(n15709), .ZN(n6746) );
  NAND2_X1 U9860 ( .A1(n10489), .A2(n10531), .ZN(n15160) );
  NAND2_X1 U9861 ( .A1(n7840), .A2(n6572), .ZN(n8114) );
  NAND2_X1 U9862 ( .A1(n7318), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n9014) );
  NAND2_X1 U9863 ( .A1(n7321), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n8892) );
  INV_X1 U9864 ( .A(n8073), .ZN(n7812) );
  INV_X1 U9865 ( .A(n7320), .ZN(n10488) );
  NAND2_X1 U9866 ( .A1(n6750), .A2(n12396), .ZN(P2_U3527) );
  NAND2_X1 U9867 ( .A1(n6864), .A2(n7787), .ZN(n6750) );
  NOR2_X1 U9868 ( .A1(n15910), .A2(n6867), .ZN(n6866) );
  NAND2_X1 U9869 ( .A1(n7254), .A2(n7253), .ZN(n11832) );
  OR2_X1 U9870 ( .A1(n13942), .A2(n11354), .ZN(n6755) );
  NAND2_X1 U9871 ( .A1(n13820), .A2(n13821), .ZN(n13819) );
  NAND2_X1 U9872 ( .A1(n10680), .A2(n10679), .ZN(n13874) );
  NAND2_X1 U9873 ( .A1(n11179), .A2(n11178), .ZN(n11181) );
  NAND2_X1 U9874 ( .A1(n10673), .A2(n10672), .ZN(n13845) );
  NAND2_X1 U9875 ( .A1(n11832), .A2(n11830), .ZN(n11828) );
  INV_X1 U9876 ( .A(n11653), .ZN(n7254) );
  NAND3_X1 U9877 ( .A1(n6756), .A2(n6755), .A3(n6754), .ZN(P2_U3233) );
  NAND2_X1 U9878 ( .A1(n12200), .A2(n9158), .ZN(n12267) );
  XNOR2_X1 U9879 ( .A(n8671), .B(n8670), .ZN(n10578) );
  NAND2_X1 U9880 ( .A1(n8340), .A2(n8093), .ZN(n8095) );
  NAND2_X1 U9881 ( .A1(n8116), .A2(n8115), .ZN(n8462) );
  INV_X1 U9882 ( .A(n8114), .ZN(n8113) );
  OAI21_X2 U9883 ( .B1(n8101), .B2(n7852), .A(n7849), .ZN(n8413) );
  NAND3_X1 U9884 ( .A1(n7837), .A2(n12630), .A3(n12628), .ZN(n6758) );
  NAND2_X1 U9885 ( .A1(n13973), .A2(n14396), .ZN(n7789) );
  NAND2_X1 U9886 ( .A1(n6682), .A2(n10073), .ZN(n10071) );
  NAND2_X1 U9887 ( .A1(n7788), .A2(n15908), .ZN(n10278) );
  NAND2_X1 U9888 ( .A1(n7469), .A2(n7468), .ZN(n12356) );
  NAND2_X1 U9889 ( .A1(n7579), .A2(n15178), .ZN(n7578) );
  INV_X1 U9890 ( .A(n10820), .ZN(n7241) );
  NOR2_X1 U9891 ( .A1(n15005), .A2(n15004), .ZN(n15003) );
  AND2_X1 U9892 ( .A1(n12586), .A2(n12585), .ZN(n12589) );
  NAND2_X1 U9893 ( .A1(n12633), .A2(n6615), .ZN(n12638) );
  NAND2_X1 U9894 ( .A1(n12581), .A2(n7365), .ZN(n7364) );
  NAND2_X1 U9895 ( .A1(n6767), .A2(n6677), .ZN(n7368) );
  NAND2_X1 U9896 ( .A1(n12601), .A2(n12602), .ZN(n6767) );
  INV_X1 U9897 ( .A(n10442), .ZN(n7890) );
  XNOR2_X1 U9898 ( .A(n7148), .B(n6662), .ZN(n14672) );
  NAND3_X1 U9899 ( .A1(n7801), .A2(n7802), .A3(n10150), .ZN(n11922) );
  AOI21_X2 U9900 ( .B1(n14270), .B2(n14024), .A(n14023), .ZN(n14301) );
  NAND2_X2 U9901 ( .A1(n14219), .A2(n14218), .ZN(n14221) );
  XNOR2_X1 U9902 ( .A(n6768), .B(n14164), .ZN(n10138) );
  NAND3_X1 U9903 ( .A1(n10137), .A2(n13956), .A3(n14013), .ZN(n6768) );
  NAND2_X1 U9904 ( .A1(n7188), .A2(n7190), .ZN(n8828) );
  NOR2_X1 U9905 ( .A1(n8806), .A2(n8786), .ZN(n7189) );
  NAND4_X1 U9906 ( .A1(n7934), .A2(n7935), .A3(n7933), .A4(n6568), .ZN(n7932)
         );
  NAND2_X1 U9907 ( .A1(n6769), .A2(n10961), .ZN(n11063) );
  NAND3_X1 U9908 ( .A1(n6771), .A2(n7650), .A3(n6770), .ZN(n7649) );
  OAI211_X2 U9909 ( .C1(n8183), .C2(n6783), .A(n6816), .B(n10902), .ZN(n10921)
         );
  INV_X2 U9910 ( .A(P3_IR_REG_0__SCAN_IN), .ZN(n15919) );
  NOR2_X1 U9911 ( .A1(n6784), .A2(n9698), .ZN(n7527) );
  NAND2_X1 U9912 ( .A1(n7262), .A2(n9500), .ZN(n6784) );
  XNOR2_X1 U9913 ( .A(n12971), .B(n12100), .ZN(n12970) );
  NAND2_X1 U9914 ( .A1(n10960), .A2(n6796), .ZN(n6800) );
  INV_X1 U9915 ( .A(n10963), .ZN(n6798) );
  OAI22_X2 U9916 ( .A1(n14170), .A2(n14180), .B1(n13797), .B2(n10227), .ZN(
        n14160) );
  NAND4_X1 U9917 ( .A1(n7439), .A2(n7438), .A3(n6549), .A4(n10226), .ZN(n6804)
         );
  NAND3_X1 U9918 ( .A1(n7439), .A2(n7438), .A3(n6549), .ZN(n6807) );
  NAND2_X1 U9919 ( .A1(n13017), .A2(n6812), .ZN(n6809) );
  NAND2_X1 U9920 ( .A1(n13017), .A2(P3_REG1_REG_13__SCAN_IN), .ZN(n6815) );
  NAND2_X1 U9921 ( .A1(n13016), .A2(n13027), .ZN(n6814) );
  AOI21_X2 U9922 ( .B1(n10910), .B2(n12955), .A(n10911), .ZN(n12959) );
  NAND2_X1 U9923 ( .A1(n6537), .A2(n8642), .ZN(n6827) );
  NAND4_X1 U9924 ( .A1(n8642), .A2(n6823), .A3(n8938), .A4(n8643), .ZN(n8647)
         );
  AND2_X1 U9925 ( .A1(n6537), .A2(n8025), .ZN(n6823) );
  NOR2_X2 U9926 ( .A1(n6824), .A2(n6827), .ZN(n8646) );
  NAND3_X1 U9927 ( .A1(n8938), .A2(n8643), .A3(n6825), .ZN(n6824) );
  OR2_X2 U9928 ( .A1(n8646), .A2(n8645), .ZN(n7150) );
  INV_X2 U9929 ( .A(n8997), .ZN(n8643) );
  AND3_X4 U9930 ( .A1(n7555), .A2(n7556), .A3(n7557), .ZN(n8938) );
  NAND2_X1 U9931 ( .A1(n14835), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n8734) );
  AND2_X4 U9932 ( .A1(n12389), .A2(n8650), .ZN(n14835) );
  NAND2_X1 U9933 ( .A1(n12720), .A2(n6831), .ZN(n6828) );
  NAND2_X1 U9934 ( .A1(n6828), .A2(n6829), .ZN(n15145) );
  NAND2_X1 U9935 ( .A1(n12720), .A2(n8041), .ZN(n12747) );
  NAND4_X1 U9936 ( .A1(n8028), .A2(n8656), .A3(n8657), .A4(n11497), .ZN(n6834)
         );
  NAND3_X1 U9937 ( .A1(n11517), .A2(n14924), .A3(n8728), .ZN(n6836) );
  NAND2_X1 U9938 ( .A1(n11517), .A2(n14924), .ZN(n6839) );
  NAND3_X1 U9939 ( .A1(n7999), .A2(n6837), .A3(n6836), .ZN(n8749) );
  OAI21_X2 U9940 ( .B1(n15220), .B2(n6842), .A(n6648), .ZN(n6843) );
  NAND2_X2 U9941 ( .A1(n6843), .A2(n12709), .ZN(n15166) );
  NAND3_X1 U9942 ( .A1(n7998), .A2(n6844), .A3(n14934), .ZN(n12208) );
  NAND2_X1 U9943 ( .A1(n13224), .A2(n6848), .ZN(n6847) );
  NAND2_X1 U9944 ( .A1(n8098), .A2(n8097), .ZN(n8367) );
  XNOR2_X1 U9945 ( .A(n6863), .B(n8717), .ZN(n10590) );
  NAND2_X1 U9946 ( .A1(n8702), .A2(n8701), .ZN(n6863) );
  NAND2_X1 U9947 ( .A1(n6870), .A2(n13622), .ZN(n13970) );
  NAND3_X1 U9948 ( .A1(n7789), .A2(n6866), .A3(n6870), .ZN(n6864) );
  NAND3_X1 U9949 ( .A1(n7789), .A2(n6868), .A3(n6870), .ZN(n7788) );
  NAND2_X2 U9950 ( .A1(n7263), .A2(n10245), .ZN(n14017) );
  NAND2_X1 U9951 ( .A1(n10227), .A2(n14431), .ZN(n6882) );
  NAND2_X1 U9952 ( .A1(n6884), .A2(n6881), .ZN(n14146) );
  NAND3_X1 U9953 ( .A1(n7973), .A2(n10202), .A3(n14114), .ZN(n14070) );
  NAND2_X1 U9954 ( .A1(n13077), .A2(n13075), .ZN(n13073) );
  NAND2_X1 U9955 ( .A1(n6889), .A2(n13063), .ZN(n13075) );
  NAND2_X1 U9956 ( .A1(n13055), .A2(n13054), .ZN(n6889) );
  NAND2_X1 U9957 ( .A1(n7400), .A2(n7399), .ZN(n13055) );
  NOR2_X1 U9958 ( .A1(n6891), .A2(n6719), .ZN(n6890) );
  INV_X1 U9959 ( .A(n7683), .ZN(n6891) );
  OAI211_X1 U9960 ( .C1(n13101), .C2(n13118), .A(n6900), .B(n6899), .ZN(
        P3_U3199) );
  NAND2_X1 U9961 ( .A1(n6901), .A2(n15916), .ZN(n6900) );
  OAI21_X1 U9962 ( .B1(n13091), .B2(P3_REG2_REG_17__SCAN_IN), .A(n13108), .ZN(
        n6901) );
  NAND3_X1 U9963 ( .A1(n6904), .A2(n6903), .A3(n6902), .ZN(P2_U3328) );
  NAND2_X1 U9964 ( .A1(n7514), .A2(n6546), .ZN(n6905) );
  NAND2_X1 U9965 ( .A1(n6905), .A2(n6672), .ZN(n6904) );
  AOI21_X1 U9966 ( .B1(n9890), .B2(n9889), .A(n9888), .ZN(n6907) );
  NOR2_X4 U9967 ( .A1(n9542), .A2(n9472), .ZN(n7795) );
  NAND2_X1 U9968 ( .A1(n6909), .A2(n6908), .ZN(n9542) );
  NAND3_X1 U9969 ( .A1(n6914), .A2(n6913), .A3(n6912), .ZN(n6911) );
  NAND2_X1 U9970 ( .A1(n6694), .A2(n6542), .ZN(n6916) );
  NAND2_X1 U9971 ( .A1(n7535), .A2(n9815), .ZN(n6926) );
  NAND3_X1 U9972 ( .A1(n11416), .A2(n6528), .A3(n6927), .ZN(n11417) );
  NAND2_X1 U9973 ( .A1(n11422), .A2(n10196), .ZN(n11412) );
  INV_X4 U9974 ( .A(n11422), .ZN(n13615) );
  AND2_X2 U9975 ( .A1(n11003), .A2(n11002), .ZN(n11422) );
  NAND3_X1 U9976 ( .A1(n6934), .A2(n6932), .A3(n11893), .ZN(n11896) );
  NAND3_X1 U9977 ( .A1(n11713), .A2(n11779), .A3(n6935), .ZN(n6934) );
  NAND2_X1 U9978 ( .A1(n13704), .A2(n6940), .ZN(n6939) );
  NAND2_X1 U9979 ( .A1(n12666), .A2(n13639), .ZN(n13704) );
  NAND2_X1 U9980 ( .A1(n13684), .A2(n12685), .ZN(n13738) );
  NAND2_X1 U9981 ( .A1(n13534), .A2(n6944), .ZN(n6943) );
  NAND2_X1 U9982 ( .A1(n7527), .A2(n7795), .ZN(n9502) );
  INV_X1 U9983 ( .A(n6953), .ZN(n6951) );
  NAND2_X1 U9984 ( .A1(n13937), .A2(n15870), .ZN(n6952) );
  NAND2_X1 U9985 ( .A1(n12304), .A2(n6702), .ZN(n15845) );
  INV_X1 U9986 ( .A(n6958), .ZN(n15844) );
  INV_X1 U9987 ( .A(n15846), .ZN(n6961) );
  NAND2_X1 U9988 ( .A1(n10873), .A2(n6570), .ZN(n6965) );
  INV_X1 U9989 ( .A(n6965), .ZN(n11169) );
  MUX2_X1 U9990 ( .A(n10564), .B(P2_REG1_REG_1__SCAN_IN), .S(n10574), .Z(
        n13818) );
  NAND3_X1 U9991 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .A3(
        P2_IR_REG_31__SCAN_IN), .ZN(n6967) );
  NAND4_X1 U9992 ( .A1(n7231), .A2(n8216), .A3(n8052), .A4(n6576), .ZN(n8058)
         );
  NAND2_X1 U9993 ( .A1(n8384), .A2(n6988), .ZN(n6986) );
  NAND2_X1 U9994 ( .A1(n13264), .A2(n6995), .ZN(n6994) );
  NAND3_X1 U9995 ( .A1(n7009), .A2(n7008), .A3(n14799), .ZN(n7007) );
  NAND2_X1 U9996 ( .A1(n6680), .A2(n6530), .ZN(n7008) );
  NAND3_X1 U9997 ( .A1(n7550), .A2(n7010), .A3(n7551), .ZN(n7009) );
  AND2_X1 U9998 ( .A1(n6530), .A2(n6683), .ZN(n7010) );
  NAND3_X1 U9999 ( .A1(n7013), .A2(n7012), .A3(n7011), .ZN(n7559) );
  NAND3_X1 U10000 ( .A1(n6543), .A2(n7016), .A3(n14735), .ZN(n7011) );
  NAND3_X1 U10001 ( .A1(n7561), .A2(n7563), .A3(n7014), .ZN(n7013) );
  XNOR2_X2 U10002 ( .A(n7017), .B(P1_IR_REG_19__SCAN_IN), .ZN(n15103) );
  NAND2_X1 U10003 ( .A1(n7354), .A2(n7544), .ZN(n7026) );
  NAND3_X1 U10004 ( .A1(n7023), .A2(n7022), .A3(n7027), .ZN(n14822) );
  NAND3_X1 U10005 ( .A1(n7025), .A2(n14811), .A3(n7024), .ZN(n7022) );
  NAND3_X1 U10006 ( .A1(n7025), .A2(n7029), .A3(n7024), .ZN(n7023) );
  INV_X1 U10007 ( .A(n7028), .ZN(n7025) );
  OAI21_X1 U10008 ( .B1(n7539), .B2(n14813), .A(n7026), .ZN(n7028) );
  MUX2_X1 U10009 ( .A(n11885), .B(n11849), .S(n14719), .Z(n14728) );
  AND2_X2 U10010 ( .A1(n14833), .A2(n14692), .ZN(n14719) );
  INV_X1 U10011 ( .A(n7502), .ZN(n15568) );
  XNOR2_X1 U10012 ( .A(n7502), .B(P3_ADDR_REG_8__SCAN_IN), .ZN(n15609) );
  NAND2_X1 U10013 ( .A1(n15566), .A2(n7038), .ZN(n7035) );
  XNOR2_X2 U10014 ( .A(n15565), .B(n15564), .ZN(n15596) );
  NAND2_X1 U10015 ( .A1(n15585), .A2(n15587), .ZN(n7373) );
  NAND2_X1 U10016 ( .A1(n15571), .A2(n7041), .ZN(n7040) );
  INV_X1 U10017 ( .A(n15614), .ZN(n7513) );
  OAI21_X1 U10018 ( .B1(n15612), .B2(P1_ADDR_REG_9__SCAN_IN), .A(n7505), .ZN(
        n7043) );
  INV_X1 U10019 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n7046) );
  OAI211_X1 U10020 ( .C1(n15670), .C2(n7051), .A(n7049), .B(n7047), .ZN(
        SUB_1596_U4) );
  INV_X1 U10021 ( .A(n7050), .ZN(n7048) );
  NAND3_X1 U10022 ( .A1(n15670), .A2(n7051), .A3(n7050), .ZN(n7049) );
  NAND2_X1 U10023 ( .A1(n15635), .A2(n15634), .ZN(n7056) );
  INV_X1 U10024 ( .A(n15663), .ZN(n7053) );
  AOI21_X1 U10025 ( .B1(n15663), .B2(P2_ADDR_REG_18__SCAN_IN), .A(n7055), .ZN(
        n7054) );
  INV_X1 U10026 ( .A(n15634), .ZN(n7055) );
  AND4_X2 U10027 ( .A1(n8850), .A2(n8637), .A3(n8830), .A4(n7057), .ZN(n7555)
         );
  NAND2_X1 U10028 ( .A1(n8757), .A2(n7057), .ZN(n8794) );
  NAND2_X1 U10029 ( .A1(n12963), .A2(n15917), .ZN(n12962) );
  OAI21_X1 U10030 ( .B1(n7489), .B2(n10954), .A(n10953), .ZN(n7059) );
  NAND2_X1 U10031 ( .A1(n7063), .A2(n7064), .ZN(n7693) );
  NAND2_X1 U10032 ( .A1(n9166), .A2(n7066), .ZN(n7063) );
  OAI211_X1 U10033 ( .C1(n7076), .C2(n11104), .A(n11041), .B(n7069), .ZN(
        n11205) );
  NAND3_X1 U10034 ( .A1(n11104), .A2(n7073), .A3(n7071), .ZN(n7070) );
  NAND2_X1 U10035 ( .A1(n7073), .A2(n11041), .ZN(n7072) );
  OAI21_X1 U10036 ( .B1(n11104), .B2(n11103), .A(n11102), .ZN(n11106) );
  AOI21_X1 U10037 ( .B1(n11102), .B2(n11103), .A(n10981), .ZN(n7079) );
  NAND2_X1 U10038 ( .A1(n12313), .A2(n6687), .ZN(n12328) );
  NAND3_X1 U10039 ( .A1(n7087), .A2(n7086), .A3(n7085), .ZN(n10923) );
  NAND3_X1 U10040 ( .A1(n7490), .A2(n7493), .A3(n7088), .ZN(n7087) );
  AND2_X2 U10041 ( .A1(n7089), .A2(n8052), .ZN(n8056) );
  NAND3_X1 U10042 ( .A1(n7089), .A2(n8052), .A3(n7218), .ZN(n7219) );
  NAND3_X1 U10043 ( .A1(n7784), .A2(n7089), .A3(n6576), .ZN(n8132) );
  NAND2_X2 U10044 ( .A1(n9190), .A2(n15536), .ZN(n9089) );
  NAND2_X1 U10045 ( .A1(n13197), .A2(n7100), .ZN(n13182) );
  NAND2_X1 U10046 ( .A1(n7099), .A2(n7771), .ZN(n8612) );
  NAND2_X1 U10047 ( .A1(n13197), .A2(n6674), .ZN(n7099) );
  NAND2_X1 U10048 ( .A1(n13197), .A2(n12463), .ZN(n13184) );
  NAND3_X1 U10049 ( .A1(n7103), .A2(n7102), .A3(n7107), .ZN(n8232) );
  NAND4_X1 U10050 ( .A1(n8642), .A2(n8643), .A3(n6652), .A4(n6537), .ZN(n7118)
         );
  NAND2_X1 U10051 ( .A1(n8644), .A2(n8643), .ZN(n9211) );
  AND3_X2 U10052 ( .A1(n8642), .A2(n8938), .A3(n6537), .ZN(n8644) );
  NAND3_X1 U10053 ( .A1(n15805), .A2(n7358), .A3(n11909), .ZN(n12255) );
  NAND2_X1 U10054 ( .A1(n9197), .A2(n15187), .ZN(n15173) );
  NAND2_X2 U10055 ( .A1(n9194), .A2(n7129), .ZN(n7130) );
  NAND2_X1 U10056 ( .A1(n7132), .A2(n7137), .ZN(n11547) );
  OR2_X1 U10057 ( .A1(n15706), .A2(n15705), .ZN(n7132) );
  OR2_X1 U10058 ( .A1(n10318), .A2(n6597), .ZN(n7135) );
  AOI21_X1 U10059 ( .B1(n15705), .B2(n10318), .A(n6597), .ZN(n7133) );
  NAND2_X1 U10060 ( .A1(n15706), .A2(n10318), .ZN(n7134) );
  OAI21_X1 U10061 ( .B1(n15706), .B2(n7136), .A(n6668), .ZN(n7138) );
  NAND2_X1 U10062 ( .A1(n7139), .A2(n10434), .ZN(n7141) );
  NAND2_X1 U10063 ( .A1(n7147), .A2(n9030), .ZN(n9139) );
  INV_X2 U10064 ( .A(n8692), .ZN(n8980) );
  XNOR2_X2 U10065 ( .A(n7150), .B(P1_IR_REG_30__SCAN_IN), .ZN(n8654) );
  NAND3_X1 U10066 ( .A1(n7645), .A2(n14013), .A3(n7646), .ZN(n7151) );
  NAND2_X1 U10067 ( .A1(n7152), .A2(n14017), .ZN(n7421) );
  NAND2_X1 U10068 ( .A1(n7158), .A2(n7156), .ZN(P2_U3496) );
  OR2_X1 U10069 ( .A1(n15908), .A2(n7157), .ZN(n7156) );
  NAND2_X1 U10070 ( .A1(n12388), .A2(n15908), .ZN(n7158) );
  INV_X1 U10071 ( .A(n13965), .ZN(n7159) );
  INV_X1 U10072 ( .A(n7161), .ZN(n7160) );
  NAND2_X1 U10073 ( .A1(n10025), .A2(n7164), .ZN(n7171) );
  NAND3_X1 U10074 ( .A1(n7171), .A2(n7172), .A3(n7165), .ZN(n14467) );
  NAND2_X1 U10075 ( .A1(n9009), .A2(n7181), .ZN(n7182) );
  NAND2_X1 U10076 ( .A1(n7187), .A2(n7924), .ZN(n9099) );
  NAND2_X1 U10077 ( .A1(n7187), .A2(n6666), .ZN(n7184) );
  NAND3_X1 U10078 ( .A1(n7184), .A2(n7185), .A3(n7182), .ZN(n9874) );
  NAND3_X1 U10079 ( .A1(n7184), .A2(n7183), .A3(n7182), .ZN(n9116) );
  NAND2_X1 U10080 ( .A1(n8788), .A2(n8787), .ZN(n7193) );
  NAND2_X1 U10081 ( .A1(n8788), .A2(n7189), .ZN(n7188) );
  NAND2_X1 U10082 ( .A1(n10078), .A2(n7194), .ZN(n7197) );
  OAI211_X1 U10083 ( .C1(n13945), .C2(n9947), .A(n7195), .B(n6574), .ZN(n7194)
         );
  NAND2_X1 U10084 ( .A1(n13945), .A2(n10092), .ZN(n7195) );
  OAI21_X1 U10085 ( .B1(n7290), .B2(n10071), .A(n7197), .ZN(n7196) );
  AND2_X2 U10086 ( .A1(n7202), .A2(n7201), .ZN(n12887) );
  OR2_X2 U10087 ( .A1(n12821), .A2(n6690), .ZN(n7202) );
  NAND2_X1 U10088 ( .A1(n12927), .A2(n7209), .ZN(n7208) );
  NAND2_X1 U10089 ( .A1(n12927), .A2(n12926), .ZN(n12925) );
  NAND2_X1 U10090 ( .A1(n12925), .A2(n7750), .ZN(n12856) );
  INV_X2 U10091 ( .A(n11759), .ZN(n12832) );
  INV_X1 U10092 ( .A(n7219), .ZN(n8555) );
  AOI21_X1 U10093 ( .B1(n12172), .B2(n6664), .A(n7727), .ZN(n12927) );
  INV_X1 U10094 ( .A(n11759), .ZN(n12791) );
  NAND2_X1 U10095 ( .A1(n11869), .A2(n11868), .ZN(n12119) );
  AND2_X1 U10096 ( .A1(n11451), .A2(n11222), .ZN(n11223) );
  INV_X1 U10097 ( .A(n14911), .ZN(n7304) );
  NAND2_X1 U10098 ( .A1(n7223), .A2(n10233), .ZN(n14106) );
  NAND3_X1 U10099 ( .A1(n7220), .A2(n13975), .A3(n13974), .ZN(P2_U3237) );
  OAI21_X1 U10100 ( .B1(n13970), .B2(n7221), .A(n14231), .ZN(n7220) );
  NAND2_X1 U10101 ( .A1(n7222), .A2(n6711), .ZN(n7221) );
  NAND2_X1 U10102 ( .A1(n13971), .A2(n14164), .ZN(n7222) );
  NAND2_X1 U10103 ( .A1(n12846), .A2(n12847), .ZN(n12803) );
  NAND3_X1 U10104 ( .A1(n14160), .A2(n14159), .A3(n10231), .ZN(n7223) );
  NAND2_X1 U10105 ( .A1(n7422), .A2(n7426), .ZN(n7263) );
  NAND2_X1 U10106 ( .A1(n14408), .A2(n7224), .ZN(P2_U3493) );
  NAND2_X1 U10107 ( .A1(n14292), .A2(n7225), .ZN(P2_U3525) );
  NAND2_X1 U10109 ( .A1(n10789), .A2(n10787), .ZN(n10993) );
  NAND2_X1 U10110 ( .A1(n10784), .A2(n11759), .ZN(n7235) );
  NAND2_X1 U10111 ( .A1(n12840), .A2(n12839), .ZN(n12838) );
  NAND2_X1 U10112 ( .A1(n12895), .A2(n7267), .ZN(n7266) );
  NAND2_X1 U10113 ( .A1(n15247), .A2(n7704), .ZN(n7236) );
  INV_X1 U10114 ( .A(n10048), .ZN(n7239) );
  INV_X1 U10115 ( .A(n7240), .ZN(n12377) );
  NAND2_X1 U10116 ( .A1(n7240), .A2(n6691), .ZN(n7429) );
  NAND2_X2 U10117 ( .A1(n8675), .A2(n8674), .ZN(n10752) );
  NAND2_X1 U10118 ( .A1(n7586), .A2(n7585), .ZN(n11981) );
  OAI22_X1 U10119 ( .A1(n15102), .A2(n15097), .B1(n15098), .B2(n15099), .ZN(
        n7579) );
  OAI211_X1 U10120 ( .C1(n7580), .C2(n15178), .A(n7578), .B(n7576), .ZN(
        P1_U3262) );
  NAND2_X1 U10121 ( .A1(n12373), .A2(n12372), .ZN(n12374) );
  XNOR2_X1 U10122 ( .A(n15110), .B(n7360), .ZN(n7359) );
  NAND2_X1 U10123 ( .A1(n13981), .A2(n13980), .ZN(n13979) );
  INV_X1 U10124 ( .A(n7806), .ZN(n7467) );
  INV_X4 U10125 ( .A(n8697), .ZN(n8743) );
  NAND2_X1 U10126 ( .A1(n8933), .A2(n8932), .ZN(n8937) );
  NAND2_X1 U10127 ( .A1(n11291), .A2(n8743), .ZN(n7250) );
  NOR2_X1 U10128 ( .A1(n13934), .A2(n7252), .ZN(n15865) );
  AND2_X1 U10129 ( .A1(n13930), .A2(n13931), .ZN(n7252) );
  INV_X2 U10130 ( .A(n10897), .ZN(n8415) );
  INV_X1 U10131 ( .A(n8132), .ZN(n7492) );
  OAI21_X1 U10132 ( .B1(n13434), .B2(n15970), .A(n7259), .ZN(P3_U3485) );
  NAND2_X1 U10133 ( .A1(n12042), .A2(n12041), .ZN(n12182) );
  NAND2_X1 U10134 ( .A1(n8039), .A2(n11416), .ZN(n7323) );
  XNOR2_X2 U10135 ( .A(n15284), .B(n15435), .ZN(n15271) );
  NAND2_X1 U10136 ( .A1(n9009), .A2(n7930), .ZN(n7926) );
  INV_X1 U10137 ( .A(n12438), .ZN(n12435) );
  NAND2_X1 U10138 ( .A1(n12247), .A2(n9156), .ZN(n12105) );
  NAND2_X1 U10139 ( .A1(n12147), .A2(n9154), .ZN(n11905) );
  XNOR2_X1 U10140 ( .A(n7264), .B(n8772), .ZN(n10624) );
  XNOR2_X2 U10141 ( .A(n7952), .B(n8662), .ZN(n15536) );
  NAND2_X1 U10142 ( .A1(n15153), .A2(n12737), .ZN(n12764) );
  XNOR2_X1 U10143 ( .A(n12764), .B(n14947), .ZN(n15366) );
  NAND2_X1 U10144 ( .A1(n9164), .A2(n9163), .ZN(n9166) );
  NAND2_X1 U10145 ( .A1(n7326), .A2(n7325), .ZN(P2_U3526) );
  NAND2_X1 U10146 ( .A1(n7328), .A2(n7327), .ZN(P2_U3494) );
  AOI21_X1 U10147 ( .B1(n11806), .B2(n7268), .A(n6639), .ZN(n11807) );
  NAND2_X1 U10148 ( .A1(n7753), .A2(n11808), .ZN(n11869) );
  NAND2_X1 U10149 ( .A1(n7269), .A2(n12580), .ZN(n12581) );
  NAND2_X1 U10150 ( .A1(n12578), .A2(n12579), .ZN(n7269) );
  NAND2_X1 U10151 ( .A1(n7364), .A2(n7362), .ZN(n12586) );
  NAND2_X1 U10152 ( .A1(n7340), .A2(n7338), .ZN(n12623) );
  NAND2_X1 U10153 ( .A1(n12604), .A2(n6681), .ZN(n7271) );
  NAND2_X1 U10154 ( .A1(n11438), .A2(n8257), .ZN(n8262) );
  NAND2_X1 U10155 ( .A1(n13192), .A2(n13193), .ZN(n13191) );
  NAND2_X1 U10156 ( .A1(n10329), .A2(n11621), .ZN(n11842) );
  NAND2_X1 U10157 ( .A1(n14562), .A2(n7904), .ZN(n7903) );
  NAND2_X2 U10158 ( .A1(n14603), .A2(n14604), .ZN(n14602) );
  OAI21_X2 U10159 ( .B1(n14503), .B2(n10377), .A(n10376), .ZN(n14654) );
  NOR2_X2 U10160 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_3__SCAN_IN), .ZN(
        n7939) );
  XNOR2_X1 U10161 ( .A(n8828), .B(n8826), .ZN(n10664) );
  NAND2_X1 U10162 ( .A1(n13687), .A2(n13686), .ZN(n13685) );
  NAND2_X1 U10163 ( .A1(n7626), .A2(n7629), .ZN(n7625) );
  OAI21_X1 U10164 ( .B1(n14807), .B2(n14808), .A(n14806), .ZN(n14811) );
  CLKBUF_X3 U10165 ( .A(n12832), .Z(n7285) );
  INV_X1 U10166 ( .A(n8006), .ZN(n8005) );
  NOR2_X1 U10167 ( .A1(n7540), .A2(n14815), .ZN(n7539) );
  NAND2_X1 U10168 ( .A1(n10067), .A2(n10068), .ZN(n10072) );
  NAND2_X1 U10169 ( .A1(n12388), .A2(n15912), .ZN(n7688) );
  NAND2_X1 U10170 ( .A1(n12621), .A2(n6610), .ZN(n7838) );
  NAND2_X1 U10171 ( .A1(n10308), .A2(n10307), .ZN(n15706) );
  NAND2_X1 U10172 ( .A1(n8196), .A2(n8195), .ZN(n11341) );
  NAND2_X1 U10173 ( .A1(n7303), .A2(n7301), .ZN(P1_U3240) );
  NAND2_X1 U10174 ( .A1(n14672), .A2(n15709), .ZN(n7303) );
  OAI21_X2 U10175 ( .B1(n14478), .B2(n7895), .A(n7892), .ZN(n14503) );
  NAND3_X1 U10176 ( .A1(n14901), .A2(n14860), .A3(n14900), .ZN(n14911) );
  NAND2_X1 U10177 ( .A1(n7903), .A2(n7902), .ZN(n14494) );
  NAND2_X1 U10178 ( .A1(n13191), .A2(n8497), .ZN(n13178) );
  INV_X1 U10180 ( .A(n7793), .ZN(n7357) );
  NAND3_X1 U10181 ( .A1(n13629), .A2(n7309), .A3(n13766), .ZN(n13571) );
  NAND2_X1 U10182 ( .A1(n7706), .A2(n7310), .ZN(n12765) );
  INV_X1 U10183 ( .A(n12736), .ZN(n7311) );
  INV_X1 U10184 ( .A(n7611), .ZN(n7610) );
  NAND2_X1 U10185 ( .A1(n7457), .A2(n7456), .ZN(P1_U3556) );
  NAND2_X1 U10186 ( .A1(n7700), .A2(n7699), .ZN(P1_U3524) );
  NAND3_X1 U10187 ( .A1(n7701), .A2(n15364), .A3(n15365), .ZN(n15506) );
  NAND2_X1 U10188 ( .A1(n8415), .A2(n11192), .ZN(n7312) );
  NAND2_X2 U10189 ( .A1(n12538), .A2(n12537), .ZN(n11760) );
  NAND2_X1 U10190 ( .A1(n7688), .A2(n7687), .ZN(P2_U3528) );
  NAND2_X1 U10191 ( .A1(n13739), .A2(n12694), .ZN(n13699) );
  NAND2_X1 U10192 ( .A1(n7386), .A2(n7375), .ZN(n7381) );
  OAI21_X1 U10193 ( .B1(n15617), .B2(n15616), .A(n7511), .ZN(n7510) );
  NOR2_X2 U10194 ( .A1(n9183), .A2(n9182), .ZN(n7320) );
  NAND3_X1 U10195 ( .A1(n7322), .A2(n6718), .A3(n13662), .ZN(P2_U3197) );
  OAI21_X1 U10196 ( .B1(n13656), .B2(n13657), .A(n13750), .ZN(n7322) );
  XNOR2_X1 U10197 ( .A(n12791), .B(n11339), .ZN(n11083) );
  NAND2_X1 U10198 ( .A1(n14025), .A2(n14028), .ZN(n14005) );
  NAND2_X1 U10199 ( .A1(n7965), .A2(n7333), .ZN(n7967) );
  NAND2_X1 U10200 ( .A1(n11265), .A2(n6669), .ZN(n8593) );
  NAND2_X1 U10201 ( .A1(n8589), .A2(n12504), .ZN(n11265) );
  NAND2_X1 U10202 ( .A1(n7781), .A2(n6716), .ZN(n8601) );
  INV_X1 U10203 ( .A(n9845), .ZN(n7618) );
  NAND2_X1 U10204 ( .A1(n7524), .A2(n7523), .ZN(n9890) );
  OAI21_X1 U10205 ( .B1(n7519), .B2(n7518), .A(n10088), .ZN(n7517) );
  INV_X1 U10206 ( .A(n12672), .ZN(n7609) );
  AOI21_X2 U10207 ( .B1(n13992), .B2(n10187), .A(n6589), .ZN(n13981) );
  NOR2_X1 U10208 ( .A1(n12096), .A2(n12095), .ZN(n12978) );
  NAND2_X1 U10209 ( .A1(n13173), .A2(n8521), .ZN(n8523) );
  NAND2_X1 U10210 ( .A1(n8519), .A2(n8520), .ZN(n13173) );
  INV_X1 U10211 ( .A(n8063), .ZN(n8476) );
  INV_X1 U10212 ( .A(n8064), .ZN(n8502) );
  NAND2_X2 U10213 ( .A1(n12803), .A2(n7337), .ZN(n12912) );
  NAND4_X1 U10214 ( .A1(n12613), .A2(n13153), .A3(n12612), .A4(n12614), .ZN(
        n7340) );
  NOR2_X1 U10215 ( .A1(n13120), .A2(n7341), .ZN(n13125) );
  AND2_X1 U10216 ( .A1(n13121), .A2(n13132), .ZN(n7341) );
  NAND2_X1 U10217 ( .A1(n12208), .A2(n8864), .ZN(n12264) );
  NAND2_X1 U10218 ( .A1(n8751), .A2(n8750), .ZN(n7445) );
  NAND2_X1 U10219 ( .A1(n8029), .A2(n8012), .ZN(n8011) );
  INV_X1 U10220 ( .A(n15270), .ZN(n9022) );
  OAI21_X1 U10221 ( .B1(n13940), .B2(n15860), .A(n7575), .ZN(n7574) );
  NAND2_X1 U10222 ( .A1(n15560), .A2(n15559), .ZN(n15561) );
  OAI21_X1 U10223 ( .B1(n15606), .B2(P1_ADDR_REG_7__SCAN_IN), .A(n7503), .ZN(
        n7502) );
  NOR2_X1 U10224 ( .A1(n10925), .A2(n10924), .ZN(n12963) );
  OR2_X1 U10225 ( .A1(n9666), .A2(n9665), .ZN(n9697) );
  NOR2_X1 U10226 ( .A1(n9919), .A2(n9918), .ZN(n7518) );
  NAND2_X1 U10227 ( .A1(n7534), .A2(n7530), .ZN(n9664) );
  XNOR2_X2 U10228 ( .A(n7345), .B(n9499), .ZN(n12056) );
  OAI21_X2 U10229 ( .B1(n9498), .B2(P2_IR_REG_21__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n7345) );
  NAND2_X1 U10230 ( .A1(n7993), .A2(n6675), .ZN(n7992) );
  NAND2_X1 U10231 ( .A1(n7991), .A2(n7990), .ZN(n9582) );
  NAND3_X1 U10232 ( .A1(n7600), .A2(n7601), .A3(n6699), .ZN(n7524) );
  NAND2_X1 U10233 ( .A1(n8309), .A2(n8308), .ZN(n12061) );
  NAND2_X1 U10234 ( .A1(n7877), .A2(n7876), .ZN(n11789) );
  NAND2_X1 U10235 ( .A1(n8558), .A2(n13529), .ZN(n7349) );
  NAND2_X1 U10236 ( .A1(n12838), .A2(n12812), .ZN(n12895) );
  NAND2_X1 U10237 ( .A1(n11452), .A2(n11451), .ZN(n11453) );
  OAI21_X1 U10238 ( .B1(n12171), .B2(n12120), .A(n12232), .ZN(n7350) );
  OAI21_X1 U10239 ( .B1(n10621), .B2(P3_D_REG_0__SCAN_IN), .A(n8562), .ZN(
        n10782) );
  NAND2_X2 U10240 ( .A1(n7605), .A2(n7604), .ZN(n8866) );
  NAND2_X1 U10241 ( .A1(n7634), .A2(n6700), .ZN(n8669) );
  AOI21_X2 U10242 ( .B1(n13978), .B2(n14270), .A(n13977), .ZN(n14285) );
  OAI21_X1 U10243 ( .B1(n8958), .B2(n8957), .A(n8956), .ZN(n8966) );
  NAND2_X1 U10244 ( .A1(n7515), .A2(n6698), .ZN(n7514) );
  NAND2_X1 U10245 ( .A1(n7418), .A2(n8484), .ZN(n13192) );
  NAND2_X1 U10246 ( .A1(n13168), .A2(n13167), .ZN(n13166) );
  XNOR2_X1 U10247 ( .A(n10309), .B(n15700), .ZN(n14924) );
  XNOR2_X1 U10248 ( .A(n13134), .B(n13133), .ZN(n7353) );
  NAND2_X1 U10249 ( .A1(n8828), .A2(n7606), .ZN(n7605) );
  NOR2_X1 U10250 ( .A1(n7492), .A2(n7491), .ZN(n7490) );
  NAND4_X1 U10251 ( .A1(n14207), .A2(n10199), .A3(n7969), .A4(n14368), .ZN(
        n12360) );
  NOR2_X1 U10252 ( .A1(n13002), .A2(n7496), .ZN(n13030) );
  NAND2_X1 U10253 ( .A1(n9152), .A2(n11850), .ZN(n11853) );
  NAND2_X1 U10254 ( .A1(n7938), .A2(n8703), .ZN(n8718) );
  NOR2_X2 U10255 ( .A1(n7946), .A2(n14733), .ZN(n11909) );
  NAND2_X1 U10256 ( .A1(n7368), .A2(n7367), .ZN(n12604) );
  NAND2_X1 U10257 ( .A1(n7369), .A2(n12593), .ZN(n12595) );
  NAND3_X1 U10258 ( .A1(n12591), .A2(n13240), .A3(n12592), .ZN(n7369) );
  OAI21_X1 U10259 ( .B1(n9697), .B2(n7984), .A(n7536), .ZN(n7535) );
  NAND2_X1 U10260 ( .A1(n7517), .A2(n7516), .ZN(n7515) );
  AND2_X2 U10261 ( .A1(n15691), .A2(n15690), .ZN(n7383) );
  NAND2_X1 U10262 ( .A1(n7375), .A2(n15697), .ZN(n7384) );
  INV_X1 U10263 ( .A(n15690), .ZN(n7375) );
  INV_X1 U10264 ( .A(n15695), .ZN(n7386) );
  INV_X1 U10265 ( .A(n7394), .ZN(n15652) );
  INV_X1 U10266 ( .A(n15651), .ZN(n7391) );
  NAND2_X1 U10267 ( .A1(n15651), .A2(P2_ADDR_REG_9__SCAN_IN), .ZN(n7392) );
  INV_X1 U10268 ( .A(n7395), .ZN(n15601) );
  NAND2_X1 U10269 ( .A1(n15649), .A2(n15648), .ZN(n15603) );
  NAND3_X1 U10270 ( .A1(n7400), .A2(n7399), .A3(n13063), .ZN(n7683) );
  NOR2_X1 U10271 ( .A1(n12983), .A2(n7648), .ZN(n12090) );
  INV_X1 U10272 ( .A(n11196), .ZN(n7409) );
  NAND2_X1 U10273 ( .A1(n7862), .A2(n7412), .ZN(n7411) );
  NAND3_X1 U10274 ( .A1(n7411), .A2(n7413), .A3(n7410), .ZN(P3_U3204) );
  NAND3_X1 U10275 ( .A1(n12340), .A2(n12521), .A3(n11301), .ZN(n7419) );
  NAND2_X2 U10276 ( .A1(n10897), .A2(n6533), .ZN(n8214) );
  NAND2_X1 U10277 ( .A1(n7666), .A2(n7423), .ZN(n7422) );
  NAND2_X1 U10278 ( .A1(n7437), .A2(n7435), .ZN(n7434) );
  AND2_X1 U10279 ( .A1(n14204), .A2(n10223), .ZN(n7438) );
  NAND2_X1 U10280 ( .A1(n15495), .A2(n12249), .ZN(n7441) );
  NAND2_X1 U10281 ( .A1(n8751), .A2(n7446), .ZN(n7444) );
  NAND2_X1 U10282 ( .A1(n8807), .A2(n7453), .ZN(n7452) );
  NAND3_X1 U10283 ( .A1(n7452), .A2(n8829), .A3(n7451), .ZN(n8844) );
  NAND2_X1 U10284 ( .A1(n8137), .A2(n8136), .ZN(n7459) );
  NAND2_X1 U10285 ( .A1(n8134), .A2(P3_ADDR_REG_19__SCAN_IN), .ZN(n7460) );
  XNOR2_X1 U10286 ( .A(n8700), .B(n8679), .ZN(n8698) );
  NAND2_X1 U10287 ( .A1(n10184), .A2(n7465), .ZN(n7463) );
  NAND2_X1 U10288 ( .A1(n14221), .A2(n7470), .ZN(n7469) );
  OAI211_X1 U10289 ( .C1(n14142), .C2(n10131), .A(n7798), .B(n7478), .ZN(n7476) );
  NAND2_X2 U10290 ( .A1(n13979), .A2(n10188), .ZN(n13955) );
  INV_X1 U10291 ( .A(n7724), .ZN(n15563) );
  XNOR2_X1 U10292 ( .A(n7504), .B(P3_ADDR_REG_7__SCAN_IN), .ZN(n15606) );
  INV_X1 U10293 ( .A(n15571), .ZN(n7505) );
  NAND2_X1 U10294 ( .A1(n9502), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9496) );
  NAND3_X1 U10295 ( .A1(n7529), .A2(n7528), .A3(n9647), .ZN(n7534) );
  NAND2_X1 U10296 ( .A1(n9626), .A2(n9648), .ZN(n7528) );
  NAND2_X1 U10297 ( .A1(n9627), .A2(n9648), .ZN(n7529) );
  NAND3_X1 U10298 ( .A1(n7533), .A2(n7532), .A3(n7531), .ZN(n7530) );
  OAI211_X1 U10299 ( .C1(n6613), .C2(n14770), .A(n7547), .B(n7546), .ZN(n7550)
         );
  NAND4_X1 U10300 ( .A1(n7553), .A2(n7546), .A3(n7554), .A4(n7547), .ZN(n7551)
         );
  NAND2_X1 U10301 ( .A1(n7559), .A2(n7560), .ZN(n14739) );
  NAND3_X1 U10302 ( .A1(n14724), .A2(n14723), .A3(n7562), .ZN(n7561) );
  INV_X1 U10303 ( .A(n7584), .ZN(n10839) );
  NAND2_X1 U10304 ( .A1(n10843), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n7583) );
  NAND2_X1 U10305 ( .A1(n11477), .A2(n7587), .ZN(n7586) );
  INV_X1 U10306 ( .A(n7592), .ZN(n11979) );
  NOR2_X1 U10307 ( .A1(n11482), .A2(n11478), .ZN(n7594) );
  XNOR2_X2 U10308 ( .A(n7598), .B(P1_IR_REG_2__SCAN_IN), .ZN(n14994) );
  OR2_X1 U10309 ( .A1(n7979), .A2(n9858), .ZN(n7600) );
  NAND2_X1 U10310 ( .A1(n14351), .A2(n9947), .ZN(n9777) );
  INV_X1 U10311 ( .A(n7615), .ZN(n7614) );
  NAND2_X1 U10312 ( .A1(n12190), .A2(n12651), .ZN(n7628) );
  OAI211_X1 U10313 ( .C1(n12191), .C2(n7627), .A(n7625), .B(n13728), .ZN(
        n12661) );
  INV_X1 U10314 ( .A(n6533), .ZN(n7634) );
  NAND2_X1 U10315 ( .A1(n8669), .A2(n9491), .ZN(n8682) );
  NAND2_X1 U10316 ( .A1(n11063), .A2(n7639), .ZN(n10942) );
  NAND2_X1 U10317 ( .A1(n7640), .A2(n10940), .ZN(n7639) );
  INV_X1 U10318 ( .A(n7653), .ZN(n10107) );
  NOR2_X1 U10319 ( .A1(n10239), .A2(n7662), .ZN(n7665) );
  NAND3_X1 U10320 ( .A1(n7664), .A2(n7663), .A3(n7667), .ZN(n14067) );
  NAND3_X1 U10321 ( .A1(n7664), .A2(n7663), .A3(n6696), .ZN(n7666) );
  XNOR2_X2 U10322 ( .A(n13810), .B(n7675), .ZN(n11138) );
  NAND2_X2 U10323 ( .A1(n6590), .A2(n7672), .ZN(n13810) );
  INV_X2 U10324 ( .A(n9557), .ZN(n7674) );
  INV_X1 U10325 ( .A(n11138), .ZN(n10148) );
  XNOR2_X1 U10326 ( .A(n7678), .B(n13123), .ZN(n13142) );
  NAND3_X1 U10327 ( .A1(n7679), .A2(n6554), .A3(n13119), .ZN(n7678) );
  NAND3_X1 U10328 ( .A1(n7683), .A2(n7685), .A3(n7682), .ZN(n13056) );
  NAND3_X1 U10329 ( .A1(n15360), .A2(n15812), .A3(n15359), .ZN(n7701) );
  NAND2_X1 U10330 ( .A1(n8685), .A2(n8684), .ZN(n8699) );
  NAND2_X1 U10331 ( .A1(n12248), .A2(n14933), .ZN(n12247) );
  NAND2_X1 U10332 ( .A1(n15216), .A2(n15217), .ZN(n9173) );
  NAND2_X1 U10333 ( .A1(n12201), .A2(n7455), .ZN(n12200) );
  OR2_X1 U10334 ( .A1(n8697), .A2(n10578), .ZN(n8677) );
  NAND2_X1 U10335 ( .A1(n10209), .A2(n10208), .ZN(n11470) );
  NAND2_X2 U10336 ( .A1(n9089), .A2(n10579), .ZN(n8697) );
  NOR2_X1 U10337 ( .A1(n7792), .A2(n6695), .ZN(n7791) );
  XNOR2_X1 U10338 ( .A(n9495), .B(P2_IR_REG_21__SCAN_IN), .ZN(n10056) );
  INV_X1 U10339 ( .A(n13738), .ZN(n12692) );
  INV_X1 U10340 ( .A(n7715), .ZN(n15674) );
  NAND2_X1 U10341 ( .A1(n7712), .A2(n15671), .ZN(n15615) );
  NAND2_X1 U10342 ( .A1(n7715), .A2(n7714), .ZN(n15671) );
  INV_X1 U10343 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n7713) );
  AOI21_X1 U10344 ( .B1(n15657), .B2(n15656), .A(P2_ADDR_REG_10__SCAN_IN), 
        .ZN(n7716) );
  NOR2_X1 U10345 ( .A1(n15657), .A2(n15656), .ZN(n15655) );
  AND2_X2 U10346 ( .A1(n7717), .A2(n7718), .ZN(n15691) );
  NAND2_X1 U10347 ( .A1(n8056), .A2(n6576), .ZN(n8131) );
  CLKBUF_X1 U10348 ( .A(n12172), .Z(n7725) );
  NAND2_X1 U10349 ( .A1(n6566), .A2(n7734), .ZN(n7729) );
  OAI21_X1 U10350 ( .B1(n7350), .B2(n12121), .A(n6651), .ZN(n7733) );
  NAND2_X1 U10351 ( .A1(n12912), .A2(n7736), .ZN(n7735) );
  OAI211_X1 U10352 ( .C1(n12912), .C2(n7737), .A(n12837), .B(n7735), .ZN(
        P3_U3160) );
  NAND2_X1 U10353 ( .A1(n11219), .A2(n7752), .ZN(n11452) );
  AND2_X1 U10354 ( .A1(n11223), .A2(n11218), .ZN(n7752) );
  AND2_X1 U10355 ( .A1(n11807), .A2(n11809), .ZN(n7753) );
  NAND2_X1 U10356 ( .A1(n11808), .A2(n11807), .ZN(n11811) );
  NAND2_X1 U10357 ( .A1(n12521), .A2(n12523), .ZN(n7754) );
  NAND3_X1 U10358 ( .A1(n7755), .A2(n12448), .A3(n7754), .ZN(n11437) );
  NAND3_X1 U10359 ( .A1(n8593), .A2(n8592), .A3(n12523), .ZN(n7755) );
  NAND2_X1 U10360 ( .A1(n7756), .A2(n12523), .ZN(n11435) );
  NAND2_X1 U10361 ( .A1(n11300), .A2(n11303), .ZN(n7756) );
  NAND2_X1 U10362 ( .A1(n13254), .A2(n7757), .ZN(n7761) );
  NAND3_X1 U10363 ( .A1(n7762), .A2(n7765), .A3(n12442), .ZN(n7760) );
  NAND3_X1 U10364 ( .A1(n11465), .A2(n11464), .A3(n11463), .ZN(n7801) );
  OAI21_X1 U10365 ( .B1(n10147), .B2(n11554), .A(n7803), .ZN(n11462) );
  INV_X1 U10366 ( .A(n15890), .ZN(n7804) );
  NAND3_X1 U10367 ( .A1(n8181), .A2(n8074), .A3(n8182), .ZN(n7813) );
  NAND3_X1 U10368 ( .A1(n7813), .A2(n8075), .A3(n7811), .ZN(n8159) );
  NAND2_X1 U10369 ( .A1(n8499), .A2(n8120), .ZN(n7820) );
  NAND2_X1 U10370 ( .A1(n8088), .A2(n7822), .ZN(n7821) );
  NAND2_X1 U10371 ( .A1(n8172), .A2(n6663), .ZN(n7828) );
  NAND3_X1 U10372 ( .A1(n11301), .A2(n12521), .A3(n11302), .ZN(n7856) );
  OR2_X1 U10373 ( .A1(n8056), .A2(n13504), .ZN(n8403) );
  OAI21_X1 U10374 ( .B1(n7862), .B2(n7861), .A(n7858), .ZN(n13425) );
  NAND2_X1 U10375 ( .A1(n13155), .A2(n7865), .ZN(n7864) );
  NAND2_X1 U10376 ( .A1(n12061), .A2(n7873), .ZN(n7870) );
  NAND2_X1 U10377 ( .A1(n7870), .A2(n7871), .ZN(n13335) );
  NAND2_X1 U10378 ( .A1(n11540), .A2(n8276), .ZN(n7877) );
  NAND2_X1 U10379 ( .A1(n10784), .A2(n10794), .ZN(n8196) );
  CLKBUF_X1 U10380 ( .A(n10784), .Z(n7878) );
  NAND3_X1 U10381 ( .A1(n7878), .A2(n12494), .A3(n7285), .ZN(n10788) );
  INV_X1 U10382 ( .A(n7233), .ZN(n13122) );
  NAND3_X1 U10383 ( .A1(n7884), .A2(n14487), .A3(n7887), .ZN(n7881) );
  AND2_X1 U10384 ( .A1(n9029), .A2(n7899), .ZN(n9130) );
  CLKBUF_X1 U10385 ( .A(n7903), .Z(n7901) );
  NAND2_X1 U10386 ( .A1(n14562), .A2(n10466), .ZN(n14643) );
  INV_X1 U10387 ( .A(n7901), .ZN(n14642) );
  INV_X1 U10388 ( .A(n14644), .ZN(n7905) );
  NAND2_X1 U10389 ( .A1(n10467), .A2(n10468), .ZN(n7906) );
  OAI21_X1 U10390 ( .B1(n14602), .B2(n7915), .A(n7908), .ZN(n10515) );
  NAND2_X1 U10391 ( .A1(n10485), .A2(n10484), .ZN(n7918) );
  OAI21_X2 U10392 ( .B1(n8866), .B2(n8865), .A(n8867), .ZN(n8958) );
  MUX2_X1 U10393 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(P2_DATAO_REG_8__SCAN_IN), 
        .S(n10579), .Z(n8792) );
  MUX2_X1 U10394 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(P2_DATAO_REG_10__SCAN_IN), 
        .S(n10579), .Z(n8845) );
  MUX2_X1 U10395 ( .A(n11248), .B(n11250), .S(n10579), .Z(n8902) );
  MUX2_X1 U10396 ( .A(n11145), .B(n8868), .S(n10579), .Z(n8869) );
  MUX2_X1 U10397 ( .A(n10838), .B(n10836), .S(n10579), .Z(n8846) );
  MUX2_X1 U10398 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(P2_DATAO_REG_15__SCAN_IN), 
        .S(n10579), .Z(n8934) );
  MUX2_X1 U10399 ( .A(n11449), .B(n11447), .S(n10579), .Z(n8959) );
  MUX2_X1 U10400 ( .A(n11292), .B(n11294), .S(n10579), .Z(n8967) );
  MUX2_X1 U10401 ( .A(n11407), .B(n11405), .S(n10579), .Z(n8990) );
  MUX2_X1 U10402 ( .A(n11757), .B(n11755), .S(n10579), .Z(n9043) );
  MUX2_X1 U10403 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(P2_DATAO_REG_19__SCAN_IN), 
        .S(n10579), .Z(n9046) );
  MUX2_X1 U10404 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(P2_DATAO_REG_20__SCAN_IN), 
        .S(n10579), .Z(n9082) );
  MUX2_X1 U10405 ( .A(n14473), .B(n15547), .S(n10579), .Z(n9923) );
  NAND3_X1 U10406 ( .A1(n7943), .A2(n11512), .A3(n7944), .ZN(n7946) );
  INV_X1 U10407 ( .A(n7946), .ZN(n12146) );
  NAND2_X1 U10408 ( .A1(n7792), .A2(n9492), .ZN(n7956) );
  NAND3_X1 U10409 ( .A1(n10102), .A2(n14462), .A3(P2_IR_REG_0__SCAN_IN), .ZN(
        n7955) );
  OAI211_X2 U10410 ( .C1(P2_IR_REG_31__SCAN_IN), .C2(P2_IR_REG_28__SCAN_IN), 
        .A(n7957), .B(n7956), .ZN(n10102) );
  INV_X1 U10411 ( .A(n7970), .ZN(n14233) );
  NOR2_X2 U10412 ( .A1(n9493), .A2(n7986), .ZN(n14449) );
  OAI21_X1 U10413 ( .B1(n9531), .B2(n9534), .A(n7992), .ZN(n7990) );
  OR2_X1 U10414 ( .A1(n7993), .A2(n6675), .ZN(n7991) );
  INV_X1 U10415 ( .A(n9548), .ZN(n7993) );
  NAND2_X2 U10416 ( .A1(n9022), .A2(n9021), .ZN(n15268) );
  NAND2_X1 U10417 ( .A1(n8007), .A2(n8005), .ZN(n8923) );
  NAND2_X1 U10418 ( .A1(n12263), .A2(n8008), .ZN(n8007) );
  NAND2_X1 U10419 ( .A1(n9200), .A2(n6686), .ZN(n8016) );
  OAI211_X1 U10420 ( .C1(n9200), .C2(n6732), .A(n8016), .B(n8017), .ZN(
        P1_U3552) );
  NAND2_X1 U10421 ( .A1(n9196), .A2(n9195), .ZN(n12332) );
  INV_X1 U10422 ( .A(n12320), .ZN(n9196) );
  NAND2_X1 U10423 ( .A1(n8146), .A2(n8145), .ZN(n8079) );
  NAND2_X1 U10424 ( .A1(n8058), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8059) );
  NAND2_X1 U10425 ( .A1(n15551), .A2(n9089), .ZN(n15214) );
  NAND2_X1 U10426 ( .A1(n13955), .A2(n12368), .ZN(n12373) );
  NAND2_X1 U10427 ( .A1(n9552), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n9511) );
  NAND2_X1 U10428 ( .A1(n8382), .A2(n8036), .ZN(n8384) );
  INV_X1 U10429 ( .A(n9483), .ZN(n14455) );
  OAI211_X2 U10430 ( .C1(n8488), .C2(n10581), .A(n8209), .B(n8208), .ZN(n11339) );
  NAND2_X1 U10431 ( .A1(n11789), .A2(n8292), .ZN(n11947) );
  OR2_X1 U10432 ( .A1(n14268), .A2(n10160), .ZN(n14269) );
  NAND2_X1 U10433 ( .A1(n13430), .A2(n13350), .ZN(n13162) );
  CLKBUF_X1 U10434 ( .A(n14156), .Z(n14157) );
  AND2_X2 U10435 ( .A1(n10897), .A2(n10579), .ZN(n8203) );
  INV_X1 U10436 ( .A(n12360), .ZN(n10200) );
  XNOR2_X1 U10437 ( .A(n15145), .B(n15144), .ZN(n15349) );
  INV_X1 U10438 ( .A(n15155), .ZN(n15156) );
  INV_X4 U10439 ( .A(n10295), .ZN(n14525) );
  AND2_X1 U10440 ( .A1(n10909), .A2(n7233), .ZN(n15915) );
  AND2_X2 U10441 ( .A1(n8749), .A2(n8748), .ZN(n8029) );
  NAND2_X2 U10442 ( .A1(n8654), .A2(n15532), .ZN(n14834) );
  INV_X1 U10443 ( .A(n8654), .ZN(n12389) );
  INV_X1 U10444 ( .A(n9482), .ZN(n12771) );
  NAND2_X1 U10445 ( .A1(n9482), .A2(n14455), .ZN(n9523) );
  INV_X1 U10446 ( .A(n10189), .ZN(n10190) );
  OR2_X1 U10447 ( .A1(n9470), .A2(n9469), .ZN(n8027) );
  NAND2_X1 U10448 ( .A1(n8631), .A2(n13321), .ZN(n13350) );
  AND2_X2 U10449 ( .A1(n11211), .A2(n11378), .ZN(n15822) );
  AND2_X1 U10450 ( .A1(n8653), .A2(n8652), .ZN(n8028) );
  INV_X1 U10451 ( .A(n14430), .ZN(n10276) );
  NOR2_X1 U10452 ( .A1(n9591), .A2(n9590), .ZN(n8030) );
  XNOR2_X1 U10453 ( .A(n13955), .B(n10190), .ZN(n13973) );
  INV_X1 U10454 ( .A(n15384), .ZN(n14812) );
  NAND2_X1 U10455 ( .A1(n14559), .A2(n10455), .ZN(n8032) );
  INV_X1 U10456 ( .A(n14797), .ZN(n14792) );
  NAND2_X2 U10457 ( .A1(n14706), .A2(n10549), .ZN(n10290) );
  AND2_X1 U10458 ( .A1(n8988), .A2(n8969), .ZN(n8034) );
  OR2_X1 U10459 ( .A1(n13481), .A2(n13328), .ZN(n8036) );
  INV_X1 U10460 ( .A(n12565), .ZN(n8598) );
  INV_X1 U10461 ( .A(n14386), .ZN(n10198) );
  NAND2_X2 U10462 ( .A1(n11330), .A2(n14250), .ZN(n14231) );
  INV_X1 U10463 ( .A(n14231), .ZN(n14210) );
  INV_X2 U10464 ( .A(n15906), .ZN(n15908) );
  INV_X1 U10465 ( .A(n14164), .ZN(n11354) );
  NOR4_X1 U10466 ( .A1(n14946), .A2(n15200), .A3(n9171), .A4(n15217), .ZN(
        n8037) );
  INV_X1 U10467 ( .A(n12596), .ZN(n8607) );
  AND2_X1 U10468 ( .A1(n15151), .A2(n15150), .ZN(n8038) );
  AND3_X1 U10469 ( .A1(n11413), .A2(n11412), .A3(n11411), .ZN(n8039) );
  OR2_X1 U10470 ( .A1(n9518), .A2(n9517), .ZN(n8040) );
  AND3_X1 U10471 ( .A1(n14947), .A2(n12719), .A3(n12718), .ZN(n8041) );
  INV_X1 U10472 ( .A(n11850), .ZN(n8770) );
  NAND2_X1 U10473 ( .A1(n13810), .A2(n9856), .ZN(n9514) );
  AOI21_X1 U10474 ( .B1(n9518), .B2(n9517), .A(n9515), .ZN(n9516) );
  AOI21_X1 U10475 ( .B1(n9664), .B2(n9663), .A(n9662), .ZN(n9666) );
  AND2_X1 U10476 ( .A1(n9762), .A2(n9761), .ZN(n9806) );
  AND2_X1 U10477 ( .A1(n14937), .A2(n14754), .ZN(n14755) );
  INV_X1 U10478 ( .A(n14798), .ZN(n14791) );
  NAND2_X1 U10479 ( .A1(n14970), .A2(n7945), .ZN(n9148) );
  INV_X1 U10480 ( .A(n10045), .ZN(n10041) );
  AND2_X1 U10481 ( .A1(n11735), .A2(n9148), .ZN(n9149) );
  INV_X1 U10482 ( .A(n14820), .ZN(n14821) );
  NAND2_X1 U10483 ( .A1(n11279), .A2(n9149), .ZN(n9151) );
  INV_X1 U10484 ( .A(n12445), .ZN(n12501) );
  AND2_X1 U10485 ( .A1(n10046), .A2(n10043), .ZN(n10088) );
  INV_X1 U10486 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n9478) );
  NOR2_X1 U10487 ( .A1(P3_IR_REG_17__SCAN_IN), .A2(P3_IR_REG_5__SCAN_IN), .ZN(
        n8051) );
  INV_X1 U10488 ( .A(P3_IR_REG_6__SCAN_IN), .ZN(n8043) );
  INV_X1 U10489 ( .A(n14320), .ZN(n10202) );
  NAND2_X1 U10490 ( .A1(n8927), .A2(n8926), .ZN(n8929) );
  NAND2_X1 U10491 ( .A1(n12637), .A2(n12632), .ZN(n12633) );
  INV_X1 U10492 ( .A(P3_IR_REG_24__SCAN_IN), .ZN(n8554) );
  OR2_X1 U10493 ( .A1(n14039), .A2(n13788), .ZN(n10185) );
  INV_X1 U10494 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n8891) );
  INV_X1 U10495 ( .A(n15122), .ZN(n15123) );
  INV_X1 U10496 ( .A(n15217), .ZN(n9098) );
  INV_X1 U10497 ( .A(n15271), .ZN(n9021) );
  INV_X1 U10498 ( .A(n14941), .ZN(n9161) );
  OAI211_X1 U10499 ( .C1(n7941), .C2(n15804), .A(n15356), .B(n15355), .ZN(
        n15357) );
  NOR2_X1 U10500 ( .A1(n14969), .A2(n14725), .ZN(n11851) );
  AOI21_X1 U10501 ( .B1(n8955), .B2(n8954), .A(n8953), .ZN(n8956) );
  INV_X1 U10502 ( .A(n8772), .ZN(n8773) );
  OAI21_X1 U10503 ( .B1(n12800), .B2(n12811), .A(n12799), .ZN(n12801) );
  INV_X1 U10504 ( .A(n11812), .ZN(n11809) );
  INV_X1 U10505 ( .A(P3_REG3_REG_10__SCAN_IN), .ZN(n8284) );
  INV_X1 U10506 ( .A(P3_REG3_REG_4__SCAN_IN), .ZN(n8062) );
  INV_X1 U10507 ( .A(n12454), .ZN(n12573) );
  NAND2_X1 U10508 ( .A1(n10116), .A2(n11354), .ZN(n10143) );
  INV_X1 U10509 ( .A(n14145), .ZN(n10171) );
  AND2_X1 U10510 ( .A1(n14269), .A2(n14222), .ZN(n14244) );
  NAND2_X1 U10511 ( .A1(n13812), .A2(n10196), .ZN(n10122) );
  OR2_X1 U10512 ( .A1(n10474), .A2(n10473), .ZN(n10475) );
  INV_X1 U10513 ( .A(n14503), .ZN(n14650) );
  INV_X1 U10514 ( .A(n8693), .ZN(n8778) );
  AND2_X1 U10515 ( .A1(n15363), .A2(n15362), .ZN(n15364) );
  AOI21_X1 U10516 ( .B1(n8964), .B2(n8963), .A(n8962), .ZN(n8965) );
  INV_X1 U10517 ( .A(P3_ADDR_REG_19__SCAN_IN), .ZN(n8136) );
  INV_X1 U10518 ( .A(n13169), .ZN(n12807) );
  INV_X1 U10519 ( .A(n12929), .ZN(n12917) );
  INV_X1 U10520 ( .A(n15914), .ZN(n13116) );
  NAND2_X1 U10521 ( .A1(n13346), .A2(P3_REG2_REG_28__SCAN_IN), .ZN(n13161) );
  AND2_X1 U10522 ( .A1(n12587), .A2(n13258), .ZN(n13279) );
  INV_X1 U10523 ( .A(n8594), .ZN(n12448) );
  OR2_X1 U10524 ( .A1(n10548), .A2(n10712), .ZN(n10895) );
  AND2_X1 U10525 ( .A1(n12583), .A2(n12580), .ZN(n12443) );
  AND2_X1 U10526 ( .A1(n12571), .A2(n12567), .ZN(n12453) );
  AND2_X1 U10527 ( .A1(n10591), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n8077) );
  AND2_X1 U10528 ( .A1(n10191), .A2(n10140), .ZN(n11007) );
  INV_X1 U10529 ( .A(n13773), .ZN(n13759) );
  AND2_X2 U10530 ( .A1(n12771), .A2(n9483), .ZN(n9550) );
  INV_X1 U10531 ( .A(n12769), .ZN(n13945) );
  INV_X1 U10532 ( .A(n13770), .ZN(n13743) );
  AND2_X1 U10533 ( .A1(n14187), .A2(n10121), .ZN(n14204) );
  NAND2_X1 U10534 ( .A1(n14854), .A2(n9628), .ZN(n9967) );
  INV_X1 U10535 ( .A(n14270), .ZN(n14127) );
  AND2_X1 U10536 ( .A1(n14468), .A2(n10265), .ZN(n10266) );
  INV_X1 U10537 ( .A(n15212), .ZN(n15392) );
  INV_X1 U10538 ( .A(n15240), .ZN(n15410) );
  OR2_X1 U10539 ( .A1(n14606), .A2(n12723), .ZN(n14681) );
  NAND2_X1 U10540 ( .A1(n14884), .A2(n14882), .ZN(n14883) );
  INV_X1 U10541 ( .A(n15798), .ZN(n12723) );
  INV_X1 U10542 ( .A(n10526), .ZN(n14956) );
  AND2_X1 U10543 ( .A1(n15550), .A2(n15542), .ZN(n10643) );
  INV_X1 U10544 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n9208) );
  AND2_X1 U10545 ( .A1(n9008), .A2(n8992), .ZN(n9006) );
  AND2_X1 U10546 ( .A1(n10721), .A2(n10720), .ZN(n11090) );
  INV_X1 U10547 ( .A(n12937), .ZN(n12919) );
  AND2_X1 U10548 ( .A1(n8483), .A2(n8482), .ZN(n12897) );
  INV_X1 U10549 ( .A(n13129), .ZN(n15922) );
  INV_X1 U10550 ( .A(n13265), .ZN(n13339) );
  AND2_X1 U10551 ( .A1(n8632), .A2(n11366), .ZN(n13310) );
  AND2_X1 U10552 ( .A1(n8582), .A2(n8581), .ZN(n8628) );
  INV_X1 U10553 ( .A(n12453), .ZN(n12060) );
  INV_X1 U10554 ( .A(n15946), .ZN(n15960) );
  NAND2_X1 U10555 ( .A1(n15957), .A2(n15956), .ZN(n13407) );
  NAND2_X1 U10556 ( .A1(n8618), .A2(n12490), .ZN(n15946) );
  INV_X1 U10557 ( .A(P3_IR_REG_10__SCAN_IN), .ZN(n8280) );
  NAND2_X1 U10558 ( .A1(n11426), .A2(P2_STATE_REG_SCAN_IN), .ZN(n13775) );
  INV_X1 U10559 ( .A(n15871), .ZN(n15850) );
  INV_X1 U10560 ( .A(n15860), .ZN(n15830) );
  OR2_X1 U10561 ( .A1(n10131), .A2(n10174), .ZN(n14124) );
  INV_X1 U10562 ( .A(n14256), .ZN(n14278) );
  INV_X1 U10563 ( .A(n14267), .ZN(n14253) );
  AND2_X1 U10564 ( .A1(n11324), .A2(n10271), .ZN(n11132) );
  NOR2_X1 U10565 ( .A1(n14466), .A2(n10266), .ZN(n15872) );
  OR2_X1 U10566 ( .A1(n10628), .A2(n11382), .ZN(n10741) );
  NOR2_X1 U10567 ( .A1(n15725), .A2(n10742), .ZN(n15742) );
  AND2_X1 U10568 ( .A1(n10631), .A2(n10742), .ZN(n15798) );
  AND2_X1 U10569 ( .A1(n11380), .A2(n14956), .ZN(n11387) );
  AOI21_X1 U10570 ( .B1(n9239), .B2(n9238), .A(n10643), .ZN(n11378) );
  INV_X1 U10571 ( .A(n15701), .ZN(n15804) );
  INV_X1 U10572 ( .A(n15807), .ZN(n15465) );
  INV_X1 U10573 ( .A(n15812), .ZN(n15492) );
  NAND2_X1 U10574 ( .A1(n11381), .A2(n11386), .ZN(n15701) );
  INV_X1 U10575 ( .A(n9239), .ZN(n10639) );
  INV_X1 U10576 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n8722) );
  INV_X1 U10577 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n15581) );
  INV_X1 U10578 ( .A(n15671), .ZN(n15672) );
  AND2_X1 U10579 ( .A1(n8580), .A2(n13519), .ZN(n10712) );
  NAND2_X1 U10580 ( .A1(n10729), .A2(n10728), .ZN(n12922) );
  INV_X1 U10581 ( .A(n13181), .ZN(n12940) );
  INV_X1 U10582 ( .A(n13247), .ZN(n13276) );
  INV_X1 U10583 ( .A(n15913), .ZN(n15925) );
  INV_X1 U10584 ( .A(n15915), .ZN(n13118) );
  OR2_X1 U10585 ( .A1(n10908), .A2(n10900), .ZN(n13141) );
  NAND2_X1 U10586 ( .A1(n13350), .A2(n8630), .ZN(n13352) );
  NAND2_X1 U10587 ( .A1(n10732), .A2(n10731), .ZN(n13321) );
  AND2_X2 U10588 ( .A1(n8628), .A2(n8587), .ZN(n15973) );
  INV_X1 U10589 ( .A(n12920), .ZN(n13436) );
  NAND2_X1 U10590 ( .A1(n10621), .A2(n10722), .ZN(n10622) );
  INV_X1 U10591 ( .A(n10548), .ZN(n10722) );
  INV_X1 U10592 ( .A(SI_17_), .ZN(n11055) );
  INV_X1 U10593 ( .A(SI_12_), .ZN(n10653) );
  NAND2_X1 U10594 ( .A1(n9997), .A2(n9996), .ZN(n13784) );
  OR2_X1 U10595 ( .A1(n10565), .A2(n12378), .ZN(n15860) );
  INV_X1 U10596 ( .A(n14231), .ZN(n14275) );
  NAND2_X1 U10597 ( .A1(n14231), .A2(n11326), .ZN(n14256) );
  AND2_X2 U10598 ( .A1(n11132), .A2(n11131), .ZN(n15912) );
  INV_X1 U10599 ( .A(n15912), .ZN(n15910) );
  INV_X1 U10600 ( .A(n14039), .ZN(n14414) );
  OR2_X1 U10601 ( .A1(n14384), .A2(n14383), .ZN(n14445) );
  INV_X1 U10602 ( .A(n15879), .ZN(n15877) );
  INV_X1 U10603 ( .A(n15882), .ZN(n15884) );
  INV_X1 U10604 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n11145) );
  AND2_X1 U10605 ( .A1(n10630), .A2(P1_STATE_REG_SCAN_IN), .ZN(n10640) );
  NAND2_X1 U10606 ( .A1(n10524), .A2(P1_STATE_REG_SCAN_IN), .ZN(n15713) );
  INV_X1 U10607 ( .A(n15413), .ZN(n15236) );
  OR2_X1 U10608 ( .A1(n15699), .A2(n15804), .ZN(n14676) );
  OAI21_X1 U10609 ( .B1(n15132), .B2(n12754), .A(n12753), .ZN(n14961) );
  INV_X1 U10610 ( .A(n14816), .ZN(n14964) );
  INV_X1 U10611 ( .A(n15311), .ZN(n15274) );
  INV_X1 U10612 ( .A(n15742), .ZN(n15068) );
  INV_X1 U10613 ( .A(n15745), .ZN(n15097) );
  INV_X1 U10614 ( .A(n15722), .ZN(n15750) );
  INV_X1 U10615 ( .A(n15341), .ZN(n15301) );
  INV_X1 U10616 ( .A(n15290), .ZN(n15343) );
  INV_X1 U10617 ( .A(n15822), .ZN(n15820) );
  INV_X1 U10618 ( .A(n15815), .ZN(n15813) );
  AND2_X2 U10619 ( .A1(n11211), .A2(n11210), .ZN(n15815) );
  INV_X1 U10620 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n11755) );
  INV_X1 U10621 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n11250) );
  XNOR2_X1 U10622 ( .A(n15582), .B(n15581), .ZN(n15975) );
  AND2_X2 U10623 ( .A1(n10722), .A2(n10712), .ZN(P3_U3897) );
  AND2_X1 U10624 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10553), .ZN(P2_U3947) );
  NOR2_X1 U10625 ( .A1(P3_IR_REG_8__SCAN_IN), .A2(P3_IR_REG_7__SCAN_IN), .ZN(
        n8045) );
  NAND4_X1 U10626 ( .A1(n8045), .A2(n8044), .A3(n8043), .A4(n8280), .ZN(n8312)
         );
  INV_X1 U10627 ( .A(P3_IR_REG_25__SCAN_IN), .ZN(n8054) );
  INV_X1 U10628 ( .A(P3_IR_REG_30__SCAN_IN), .ZN(n8057) );
  NAND2_X1 U10629 ( .A1(n8517), .A2(P3_REG0_REG_28__SCAN_IN), .ZN(n8072) );
  AND2_X2 U10630 ( .A1(n8061), .A2(n8060), .ZN(n8197) );
  NAND2_X1 U10631 ( .A1(n12398), .A2(P3_REG1_REG_28__SCAN_IN), .ZN(n8071) );
  INV_X1 U10632 ( .A(n8061), .ZN(n8068) );
  INV_X1 U10633 ( .A(P3_REG3_REG_27__SCAN_IN), .ZN(n12806) );
  INV_X1 U10634 ( .A(P3_REG3_REG_14__SCAN_IN), .ZN(n8346) );
  INV_X1 U10635 ( .A(P3_REG3_REG_15__SCAN_IN), .ZN(n8360) );
  INV_X1 U10636 ( .A(P3_REG3_REG_19__SCAN_IN), .ZN(n8418) );
  INV_X1 U10637 ( .A(P3_REG3_REG_22__SCAN_IN), .ZN(n12896) );
  NAND2_X1 U10638 ( .A1(n12806), .A2(n8503), .ZN(n8520) );
  INV_X1 U10639 ( .A(n8520), .ZN(n8066) );
  INV_X1 U10640 ( .A(P3_REG3_REG_28__SCAN_IN), .ZN(n8065) );
  NAND2_X1 U10641 ( .A1(n8520), .A2(P3_REG3_REG_28__SCAN_IN), .ZN(n8067) );
  NAND2_X1 U10642 ( .A1(n8633), .A2(n8067), .ZN(n13163) );
  NAND2_X1 U10643 ( .A1(n8466), .A2(n13163), .ZN(n8070) );
  NAND2_X2 U10644 ( .A1(n8068), .A2(n13510), .ZN(n8287) );
  NAND2_X1 U10645 ( .A1(n8492), .A2(P3_REG2_REG_28__SCAN_IN), .ZN(n8069) );
  NAND4_X1 U10646 ( .A1(n8072), .A2(n8071), .A3(n8070), .A4(n8069), .ZN(n13169) );
  NAND2_X1 U10647 ( .A1(n9488), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n8192) );
  NAND2_X1 U10648 ( .A1(n10573), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n8073) );
  INV_X1 U10649 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n10575) );
  NAND2_X1 U10650 ( .A1(n10575), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n8074) );
  NAND2_X1 U10651 ( .A1(n10593), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n8075) );
  NAND2_X1 U10652 ( .A1(n10576), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n8076) );
  NAND2_X1 U10653 ( .A1(n10589), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n8078) );
  NAND2_X1 U10654 ( .A1(n10618), .A2(P1_DATAO_REG_5__SCAN_IN), .ZN(n8080) );
  NAND2_X1 U10655 ( .A1(n10627), .A2(P1_DATAO_REG_6__SCAN_IN), .ZN(n8081) );
  NAND2_X1 U10656 ( .A1(n8082), .A2(n8081), .ZN(n8243) );
  NAND2_X1 U10657 ( .A1(n10656), .A2(P2_DATAO_REG_8__SCAN_IN), .ZN(n8083) );
  NAND2_X1 U10658 ( .A1(n10667), .A2(P1_DATAO_REG_9__SCAN_IN), .ZN(n8085) );
  INV_X1 U10659 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n10774) );
  NAND2_X1 U10660 ( .A1(n10838), .A2(P2_DATAO_REG_11__SCAN_IN), .ZN(n8086) );
  NAND2_X1 U10661 ( .A1(n10836), .A2(P1_DATAO_REG_11__SCAN_IN), .ZN(n8087) );
  XNOR2_X1 U10662 ( .A(n8868), .B(P1_DATAO_REG_12__SCAN_IN), .ZN(n8310) );
  INV_X1 U10663 ( .A(n8310), .ZN(n8089) );
  NAND2_X1 U10664 ( .A1(n8868), .A2(P1_DATAO_REG_12__SCAN_IN), .ZN(n8326) );
  NAND2_X1 U10665 ( .A1(n11250), .A2(P1_DATAO_REG_13__SCAN_IN), .ZN(n8090) );
  NAND2_X1 U10666 ( .A1(n11248), .A2(P2_DATAO_REG_13__SCAN_IN), .ZN(n8091) );
  NAND2_X1 U10667 ( .A1(n11449), .A2(P2_DATAO_REG_14__SCAN_IN), .ZN(n8094) );
  NAND2_X1 U10668 ( .A1(n11447), .A2(P1_DATAO_REG_14__SCAN_IN), .ZN(n8092) );
  NAND2_X1 U10669 ( .A1(n8094), .A2(n8092), .ZN(n8339) );
  INV_X1 U10670 ( .A(n8339), .ZN(n8093) );
  INV_X1 U10671 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n8096) );
  XNOR2_X1 U10672 ( .A(n8096), .B(P1_DATAO_REG_15__SCAN_IN), .ZN(n8352) );
  NAND2_X1 U10673 ( .A1(n8096), .A2(P1_DATAO_REG_15__SCAN_IN), .ZN(n8097) );
  XNOR2_X1 U10674 ( .A(n11294), .B(P1_DATAO_REG_16__SCAN_IN), .ZN(n8366) );
  INV_X1 U10675 ( .A(n8366), .ZN(n8099) );
  NAND2_X1 U10676 ( .A1(n11294), .A2(P1_DATAO_REG_16__SCAN_IN), .ZN(n8100) );
  AND2_X1 U10677 ( .A1(n11405), .A2(P1_DATAO_REG_17__SCAN_IN), .ZN(n8102) );
  NAND2_X1 U10678 ( .A1(n11755), .A2(P1_DATAO_REG_18__SCAN_IN), .ZN(n8104) );
  NAND2_X1 U10679 ( .A1(n11757), .A2(P2_DATAO_REG_18__SCAN_IN), .ZN(n8103) );
  NAND2_X1 U10680 ( .A1(n8104), .A2(n8103), .ZN(n8400) );
  INV_X1 U10681 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n11880) );
  XNOR2_X1 U10682 ( .A(n11880), .B(P2_DATAO_REG_19__SCAN_IN), .ZN(n8412) );
  INV_X1 U10683 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n11878) );
  INV_X1 U10684 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n11963) );
  NAND2_X1 U10685 ( .A1(n11963), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n8106) );
  INV_X1 U10686 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n11966) );
  NAND2_X1 U10687 ( .A1(n11966), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n8105) );
  AND2_X1 U10688 ( .A1(n8106), .A2(n8105), .ZN(n8427) );
  INV_X1 U10689 ( .A(n8427), .ZN(n8107) );
  INV_X1 U10690 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n12051) );
  NAND2_X1 U10691 ( .A1(n12051), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n8110) );
  INV_X1 U10692 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n12054) );
  NAND2_X1 U10693 ( .A1(n12054), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n8108) );
  NAND2_X1 U10694 ( .A1(n8110), .A2(n8108), .ZN(n8440) );
  INV_X1 U10695 ( .A(n8440), .ZN(n8109) );
  INV_X1 U10696 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n12058) );
  XNOR2_X1 U10697 ( .A(n12058), .B(P2_DATAO_REG_22__SCAN_IN), .ZN(n8450) );
  NAND2_X1 U10698 ( .A1(n12058), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n8112) );
  XNOR2_X1 U10699 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(P2_DATAO_REG_23__SCAN_IN), 
        .ZN(n8471) );
  INV_X1 U10700 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n12164) );
  INV_X1 U10701 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n15547) );
  NAND2_X1 U10702 ( .A1(n8114), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n8115) );
  INV_X1 U10703 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n14473) );
  INV_X1 U10704 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n15545) );
  NAND2_X1 U10705 ( .A1(n15545), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n8118) );
  INV_X1 U10706 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n14470) );
  NAND2_X1 U10707 ( .A1(n14470), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n8117) );
  AND2_X1 U10708 ( .A1(n8118), .A2(n8117), .ZN(n8486) );
  INV_X1 U10709 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n15540) );
  NAND2_X1 U10710 ( .A1(n15540), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n8121) );
  INV_X1 U10711 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n14465) );
  NAND2_X1 U10712 ( .A1(n14465), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n8119) );
  NAND2_X1 U10713 ( .A1(n8121), .A2(n8119), .ZN(n8498) );
  INV_X1 U10714 ( .A(n8498), .ZN(n8120) );
  INV_X1 U10715 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n15538) );
  NAND2_X1 U10716 ( .A1(n15538), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n8124) );
  INV_X1 U10717 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n14463) );
  NAND2_X1 U10718 ( .A1(n14463), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n8122) );
  NAND2_X1 U10719 ( .A1(n8124), .A2(n8122), .ZN(n8512) );
  INV_X1 U10720 ( .A(n8512), .ZN(n8123) );
  INV_X1 U10721 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n15535) );
  NAND2_X1 U10722 ( .A1(n15535), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n8528) );
  INV_X1 U10723 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n9938) );
  NAND2_X1 U10724 ( .A1(n9938), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n8125) );
  AND2_X1 U10725 ( .A1(n8528), .A2(n8125), .ZN(n8126) );
  OR2_X1 U10726 ( .A1(n8127), .A2(n8126), .ZN(n8128) );
  NAND2_X1 U10727 ( .A1(n8132), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8130) );
  NAND3_X1 U10728 ( .A1(n15105), .A2(n13944), .A3(n8133), .ZN(n8134) );
  NAND3_X1 U10729 ( .A1(n8135), .A2(P2_ADDR_REG_19__SCAN_IN), .A3(
        P1_ADDR_REG_19__SCAN_IN), .ZN(n8137) );
  NAND2_X1 U10730 ( .A1(n12410), .A2(SI_28_), .ZN(n8138) );
  NAND2_X1 U10731 ( .A1(n8534), .A2(P3_REG1_REG_4__SCAN_IN), .ZN(n8144) );
  NAND2_X1 U10732 ( .A1(n8517), .A2(P3_REG0_REG_4__SCAN_IN), .ZN(n8143) );
  NAND2_X1 U10733 ( .A1(P3_REG3_REG_4__SCAN_IN), .A2(P3_REG3_REG_3__SCAN_IN), 
        .ZN(n8140) );
  NAND2_X1 U10734 ( .A1(n9440), .A2(n8140), .ZN(n11272) );
  NAND2_X1 U10735 ( .A1(n8521), .A2(n11272), .ZN(n8142) );
  INV_X2 U10736 ( .A(n8287), .ZN(n12399) );
  NAND2_X1 U10737 ( .A1(n12399), .A2(P3_REG2_REG_4__SCAN_IN), .ZN(n8141) );
  XNOR2_X1 U10738 ( .A(n8146), .B(n8145), .ZN(n10605) );
  NAND2_X1 U10739 ( .A1(n8203), .A2(n10605), .ZN(n8153) );
  INV_X1 U10740 ( .A(n10902), .ZN(n8147) );
  NAND2_X1 U10741 ( .A1(n8147), .A2(n8206), .ZN(n8160) );
  OAI21_X1 U10742 ( .B1(n8160), .B2(P3_IR_REG_3__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n8148) );
  MUX2_X1 U10743 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8148), .S(
        P3_IR_REG_4__SCAN_IN), .Z(n8151) );
  INV_X1 U10744 ( .A(n8216), .ZN(n8150) );
  NAND2_X1 U10745 ( .A1(n8415), .A2(n10976), .ZN(n8152) );
  OAI211_X1 U10746 ( .C1(n8214), .C2(SI_4_), .A(n8153), .B(n8152), .ZN(n15939)
         );
  OR2_X1 U10747 ( .A1(n12344), .A2(n15939), .ZN(n12518) );
  NAND2_X1 U10748 ( .A1(n12344), .A2(n15939), .ZN(n8590) );
  NAND2_X1 U10749 ( .A1(n12398), .A2(P3_REG1_REG_3__SCAN_IN), .ZN(n8157) );
  NAND2_X1 U10750 ( .A1(n8466), .A2(n12350), .ZN(n8156) );
  NAND2_X1 U10751 ( .A1(n12399), .A2(P3_REG2_REG_3__SCAN_IN), .ZN(n8155) );
  NAND2_X1 U10752 ( .A1(n8517), .A2(P3_REG0_REG_3__SCAN_IN), .ZN(n8154) );
  XNOR2_X1 U10753 ( .A(n10591), .B(P2_DATAO_REG_3__SCAN_IN), .ZN(n8158) );
  XNOR2_X1 U10754 ( .A(n8159), .B(n8158), .ZN(n10609) );
  NAND2_X1 U10755 ( .A1(n8203), .A2(n10609), .ZN(n8164) );
  NAND2_X1 U10756 ( .A1(n8160), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8162) );
  INV_X1 U10757 ( .A(P3_IR_REG_3__SCAN_IN), .ZN(n8161) );
  XNOR2_X2 U10758 ( .A(n8162), .B(n8161), .ZN(n10961) );
  NAND2_X1 U10759 ( .A1(n8415), .A2(n10961), .ZN(n8163) );
  OAI211_X1 U10760 ( .C1(n8214), .C2(SI_3_), .A(n8164), .B(n8163), .ZN(n15933)
         );
  INV_X1 U10761 ( .A(n15933), .ZN(n12351) );
  AND2_X1 U10762 ( .A1(n12952), .A2(n12351), .ZN(n11267) );
  INV_X1 U10763 ( .A(n15939), .ZN(n11273) );
  AND2_X1 U10764 ( .A1(n12344), .A2(n11273), .ZN(n8165) );
  NAND2_X1 U10765 ( .A1(n12952), .A2(n15933), .ZN(n12510) );
  NAND2_X1 U10766 ( .A1(n12512), .A2(n12510), .ZN(n12446) );
  NAND2_X1 U10767 ( .A1(n12446), .A2(n12511), .ZN(n11302) );
  NAND2_X1 U10768 ( .A1(n8517), .A2(P3_REG0_REG_5__SCAN_IN), .ZN(n8170) );
  NAND2_X1 U10769 ( .A1(n12398), .A2(P3_REG1_REG_5__SCAN_IN), .ZN(n8169) );
  NAND2_X1 U10770 ( .A1(n9440), .A2(P3_REG3_REG_5__SCAN_IN), .ZN(n8166) );
  NAND2_X1 U10771 ( .A1(n8250), .A2(n8166), .ZN(n11450) );
  NAND2_X1 U10772 ( .A1(n8521), .A2(n11450), .ZN(n8168) );
  NAND2_X1 U10773 ( .A1(n8492), .A2(P3_REG2_REG_5__SCAN_IN), .ZN(n8167) );
  NAND4_X1 U10774 ( .A1(n8170), .A2(n8169), .A3(n8168), .A4(n8167), .ZN(n12951) );
  XNOR2_X1 U10775 ( .A(n8172), .B(n8171), .ZN(n10607) );
  NAND2_X1 U10776 ( .A1(n8203), .A2(n10607), .ZN(n8175) );
  INV_X1 U10777 ( .A(P3_IR_REG_31__SCAN_IN), .ZN(n13504) );
  OR2_X1 U10778 ( .A1(n8216), .A2(n13504), .ZN(n8173) );
  XNOR2_X1 U10779 ( .A(n8173), .B(n8215), .ZN(n10979) );
  NAND2_X1 U10780 ( .A1(n8415), .A2(n10979), .ZN(n8174) );
  OAI211_X1 U10781 ( .C1(n8214), .C2(SI_5_), .A(n8175), .B(n8174), .ZN(n15947)
         );
  OR2_X1 U10782 ( .A1(n12951), .A2(n15947), .ZN(n12523) );
  NAND2_X1 U10783 ( .A1(n12951), .A2(n15947), .ZN(n12527) );
  NAND2_X1 U10784 ( .A1(n12523), .A2(n12527), .ZN(n12521) );
  INV_X1 U10785 ( .A(n12951), .ZN(n11670) );
  NAND2_X1 U10786 ( .A1(n11670), .A2(n15947), .ZN(n8176) );
  NAND2_X1 U10787 ( .A1(n8521), .A2(P3_REG3_REG_1__SCAN_IN), .ZN(n8180) );
  NAND2_X1 U10788 ( .A1(n8197), .A2(P3_REG1_REG_1__SCAN_IN), .ZN(n8179) );
  NAND2_X1 U10789 ( .A1(n12399), .A2(P3_REG2_REG_1__SCAN_IN), .ZN(n8178) );
  NAND2_X1 U10790 ( .A1(n8517), .A2(P3_REG0_REG_1__SCAN_IN), .ZN(n8177) );
  NAND2_X1 U10791 ( .A1(n8374), .A2(SI_1_), .ZN(n8186) );
  XNOR2_X1 U10792 ( .A(n8182), .B(n8181), .ZN(n10596) );
  NAND2_X1 U10793 ( .A1(n8203), .A2(n10596), .ZN(n8185) );
  NAND2_X1 U10794 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(P3_IR_REG_0__SCAN_IN), 
        .ZN(n8183) );
  OR2_X1 U10795 ( .A1(n12954), .A2(n11310), .ZN(n12496) );
  NAND2_X1 U10796 ( .A1(n8492), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n8190) );
  NAND2_X1 U10797 ( .A1(n8521), .A2(P3_REG3_REG_0__SCAN_IN), .ZN(n8189) );
  NAND2_X1 U10798 ( .A1(n8197), .A2(P3_REG1_REG_0__SCAN_IN), .ZN(n8188) );
  NAND2_X1 U10799 ( .A1(n8517), .A2(P3_REG0_REG_0__SCAN_IN), .ZN(n8187) );
  INV_X1 U10800 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n8658) );
  NAND2_X1 U10801 ( .A1(n8658), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n8191) );
  AND2_X1 U10802 ( .A1(n8192), .A2(n8191), .ZN(n8193) );
  OAI21_X1 U10803 ( .B1(n6533), .B2(n8193), .A(n9489), .ZN(n13530) );
  INV_X1 U10804 ( .A(n13530), .ZN(n8194) );
  MUX2_X1 U10805 ( .A(n15919), .B(n8194), .S(n10897), .Z(n11190) );
  INV_X1 U10806 ( .A(n11190), .ZN(n10814) );
  NAND2_X1 U10807 ( .A1(n10796), .A2(n10814), .ZN(n10794) );
  INV_X1 U10808 ( .A(n12954), .ZN(n11343) );
  NAND2_X1 U10809 ( .A1(n11343), .A2(n11310), .ZN(n8195) );
  NAND2_X1 U10810 ( .A1(n8534), .A2(P3_REG1_REG_2__SCAN_IN), .ZN(n8202) );
  NAND2_X1 U10811 ( .A1(n8198), .A2(P3_REG3_REG_2__SCAN_IN), .ZN(n8201) );
  NAND2_X1 U10812 ( .A1(n12399), .A2(P3_REG2_REG_2__SCAN_IN), .ZN(n8200) );
  NAND2_X1 U10813 ( .A1(n8517), .A2(P3_REG0_REG_2__SCAN_IN), .ZN(n8199) );
  INV_X1 U10814 ( .A(n8203), .ZN(n8488) );
  XNOR2_X1 U10815 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(P2_DATAO_REG_2__SCAN_IN), 
        .ZN(n8204) );
  XNOR2_X1 U10816 ( .A(n8205), .B(n8204), .ZN(n10581) );
  INV_X1 U10817 ( .A(SI_2_), .ZN(n8679) );
  NAND2_X1 U10818 ( .A1(n8374), .A2(n8679), .ZN(n8209) );
  NAND2_X1 U10819 ( .A1(n10902), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8207) );
  NAND2_X1 U10820 ( .A1(n8415), .A2(n7298), .ZN(n8208) );
  NAND2_X1 U10821 ( .A1(n12953), .A2(n11339), .ZN(n12509) );
  NAND2_X1 U10822 ( .A1(n11341), .A2(n12445), .ZN(n8211) );
  INV_X1 U10823 ( .A(n12953), .ZN(n11089) );
  NAND2_X1 U10824 ( .A1(n11089), .A2(n11339), .ZN(n8210) );
  XNOR2_X1 U10825 ( .A(n10656), .B(P2_DATAO_REG_8__SCAN_IN), .ZN(n8212) );
  XNOR2_X1 U10826 ( .A(n8213), .B(n8212), .ZN(n10599) );
  INV_X2 U10827 ( .A(n8488), .ZN(n8514) );
  NAND2_X1 U10828 ( .A1(n10599), .A2(n8514), .ZN(n8224) );
  NAND2_X1 U10829 ( .A1(n8216), .A2(n8215), .ZN(n8313) );
  INV_X1 U10830 ( .A(n8237), .ZN(n8217) );
  INV_X1 U10831 ( .A(P3_IR_REG_7__SCAN_IN), .ZN(n8238) );
  NAND2_X1 U10832 ( .A1(n8217), .A2(n8238), .ZN(n8219) );
  NAND2_X1 U10833 ( .A1(n8219), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8218) );
  MUX2_X1 U10834 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8218), .S(
        P3_IR_REG_8__SCAN_IN), .Z(n8222) );
  INV_X1 U10835 ( .A(n8219), .ZN(n8221) );
  INV_X1 U10836 ( .A(P3_IR_REG_8__SCAN_IN), .ZN(n8220) );
  NAND2_X1 U10837 ( .A1(n8221), .A2(n8220), .ZN(n8279) );
  AOI22_X1 U10838 ( .A1(n12423), .A2(SI_8_), .B1(n8415), .B2(n11574), .ZN(
        n8223) );
  NAND2_X1 U10839 ( .A1(n8517), .A2(P3_REG0_REG_8__SCAN_IN), .ZN(n8229) );
  NAND2_X1 U10840 ( .A1(n8534), .A2(P3_REG1_REG_8__SCAN_IN), .ZN(n8228) );
  NAND2_X1 U10841 ( .A1(n8232), .A2(P3_REG3_REG_8__SCAN_IN), .ZN(n8225) );
  NAND2_X1 U10842 ( .A1(n8269), .A2(n8225), .ZN(n11975) );
  NAND2_X1 U10843 ( .A1(n8466), .A2(n11975), .ZN(n8227) );
  NAND2_X1 U10844 ( .A1(n8492), .A2(P3_REG2_REG_8__SCAN_IN), .ZN(n8226) );
  OR2_X1 U10845 ( .A1(n11974), .A2(n11795), .ZN(n12546) );
  NAND2_X1 U10846 ( .A1(n11974), .A2(n11795), .ZN(n12545) );
  NAND2_X1 U10847 ( .A1(n12398), .A2(P3_REG1_REG_7__SCAN_IN), .ZN(n8236) );
  NAND2_X1 U10848 ( .A1(n8492), .A2(P3_REG2_REG_7__SCAN_IN), .ZN(n8235) );
  OR2_X1 U10849 ( .A1(n8249), .A2(n8230), .ZN(n8231) );
  NAND2_X1 U10850 ( .A1(n8232), .A2(n8231), .ZN(n11764) );
  NAND2_X1 U10851 ( .A1(n8521), .A2(n11764), .ZN(n8234) );
  NAND2_X1 U10852 ( .A1(n8517), .A2(P3_REG0_REG_7__SCAN_IN), .ZN(n8233) );
  INV_X1 U10853 ( .A(SI_7_), .ZN(n10615) );
  NAND2_X1 U10854 ( .A1(n8237), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8239) );
  XNOR2_X1 U10855 ( .A(n8239), .B(n8238), .ZN(n11192) );
  XNOR2_X1 U10856 ( .A(n8241), .B(n8240), .ZN(n10616) );
  NAND2_X1 U10857 ( .A1(n10616), .A2(n12422), .ZN(n8242) );
  OR2_X2 U10858 ( .A1(n12949), .A2(n11761), .ZN(n12538) );
  NAND2_X1 U10859 ( .A1(n12949), .A2(n11761), .ZN(n12537) );
  XNOR2_X1 U10860 ( .A(n8244), .B(n8243), .ZN(n10612) );
  NAND2_X1 U10861 ( .A1(n8514), .A2(n10612), .ZN(n8248) );
  NAND2_X1 U10862 ( .A1(n12410), .A2(SI_6_), .ZN(n8247) );
  NAND2_X1 U10863 ( .A1(n8313), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8245) );
  XNOR2_X1 U10864 ( .A(n8245), .B(P3_IR_REG_6__SCAN_IN), .ZN(n11036) );
  NAND2_X1 U10865 ( .A1(n8415), .A2(n11036), .ZN(n8246) );
  NAND2_X1 U10866 ( .A1(n8517), .A2(P3_REG0_REG_6__SCAN_IN), .ZN(n8254) );
  INV_X1 U10867 ( .A(n8249), .ZN(n8252) );
  NAND2_X1 U10868 ( .A1(n8250), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n8251) );
  NAND2_X1 U10869 ( .A1(n8252), .A2(n8251), .ZN(n11668) );
  NAND2_X1 U10870 ( .A1(n12399), .A2(P3_REG2_REG_6__SCAN_IN), .ZN(n8253) );
  AND2_X1 U10871 ( .A1(n6977), .A2(n12950), .ZN(n11697) );
  NAND2_X1 U10872 ( .A1(n11760), .A2(n11697), .ZN(n8256) );
  INV_X1 U10873 ( .A(n11761), .ZN(n13413) );
  NAND2_X1 U10874 ( .A1(n13413), .A2(n12949), .ZN(n8255) );
  NAND2_X1 U10875 ( .A1(n8256), .A2(n8255), .ZN(n8258) );
  NOR2_X1 U10876 ( .A1(n12450), .A2(n8258), .ZN(n8257) );
  AND2_X1 U10877 ( .A1(n8594), .A2(n11760), .ZN(n11394) );
  NOR2_X1 U10878 ( .A1(n12450), .A2(n11394), .ZN(n8260) );
  INV_X1 U10879 ( .A(n8258), .ZN(n11395) );
  INV_X1 U10880 ( .A(n11795), .ZN(n12948) );
  NOR2_X1 U10881 ( .A1(n12948), .A2(n11974), .ZN(n8259) );
  AOI21_X1 U10882 ( .B1(n8260), .B2(n11395), .A(n8259), .ZN(n8261) );
  NAND2_X1 U10883 ( .A1(n8262), .A2(n8261), .ZN(n11540) );
  XNOR2_X1 U10884 ( .A(n10665), .B(P2_DATAO_REG_9__SCAN_IN), .ZN(n8263) );
  XNOR2_X1 U10885 ( .A(n8264), .B(n8263), .ZN(n10611) );
  NAND2_X1 U10886 ( .A1(n10611), .A2(n12422), .ZN(n8268) );
  INV_X1 U10887 ( .A(SI_9_), .ZN(n10610) );
  NAND2_X1 U10888 ( .A1(n8279), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8266) );
  INV_X1 U10889 ( .A(P3_IR_REG_9__SCAN_IN), .ZN(n8265) );
  XNOR2_X1 U10890 ( .A(n8266), .B(n8265), .ZN(n11594) );
  AOI22_X1 U10891 ( .A1(n12423), .A2(n10610), .B1(n8415), .B2(n11594), .ZN(
        n8267) );
  NAND2_X1 U10892 ( .A1(n8517), .A2(P3_REG0_REG_9__SCAN_IN), .ZN(n8275) );
  NAND2_X1 U10893 ( .A1(n12398), .A2(P3_REG1_REG_9__SCAN_IN), .ZN(n8274) );
  INV_X1 U10894 ( .A(n8285), .ZN(n8271) );
  NAND2_X1 U10895 ( .A1(n8269), .A2(P3_REG3_REG_9__SCAN_IN), .ZN(n8270) );
  NAND2_X1 U10896 ( .A1(n8271), .A2(n8270), .ZN(n11817) );
  NAND2_X1 U10897 ( .A1(n8521), .A2(n11817), .ZN(n8273) );
  NAND2_X1 U10898 ( .A1(n12399), .A2(P3_REG2_REG_9__SCAN_IN), .ZN(n8272) );
  NAND4_X1 U10899 ( .A1(n8275), .A2(n8274), .A3(n8273), .A4(n8272), .ZN(n12947) );
  XNOR2_X1 U10900 ( .A(n12551), .B(n12947), .ZN(n12550) );
  INV_X1 U10901 ( .A(n12550), .ZN(n11539) );
  INV_X1 U10902 ( .A(n12947), .ZN(n12552) );
  OR2_X1 U10903 ( .A1(n12551), .A2(n12552), .ZN(n8276) );
  XNOR2_X1 U10904 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(P2_DATAO_REG_10__SCAN_IN), 
        .ZN(n8277) );
  XNOR2_X1 U10905 ( .A(n8278), .B(n8277), .ZN(n10603) );
  NAND2_X1 U10906 ( .A1(n10603), .A2(n12422), .ZN(n8283) );
  INV_X1 U10907 ( .A(SI_10_), .ZN(n10602) );
  NAND2_X1 U10908 ( .A1(n8295), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8281) );
  AOI22_X1 U10909 ( .A1(n12423), .A2(n10602), .B1(n8415), .B2(n12089), .ZN(
        n8282) );
  NAND2_X1 U10910 ( .A1(n8283), .A2(n8282), .ZN(n11954) );
  NAND2_X1 U10911 ( .A1(n8517), .A2(P3_REG0_REG_10__SCAN_IN), .ZN(n8291) );
  NAND2_X1 U10912 ( .A1(n12398), .A2(P3_REG1_REG_10__SCAN_IN), .ZN(n8290) );
  NOR2_X1 U10913 ( .A1(n8285), .A2(n8284), .ZN(n8286) );
  OR2_X1 U10914 ( .A1(n8301), .A2(n8286), .ZN(n11958) );
  NAND2_X1 U10915 ( .A1(n8466), .A2(n11958), .ZN(n8289) );
  NAND2_X1 U10916 ( .A1(n8492), .A2(P3_REG2_REG_10__SCAN_IN), .ZN(n8288) );
  NAND4_X1 U10917 ( .A1(n8291), .A2(n8290), .A3(n8289), .A4(n8288), .ZN(n12946) );
  OR2_X1 U10918 ( .A1(n11954), .A2(n12946), .ZN(n12561) );
  NAND2_X1 U10919 ( .A1(n11954), .A2(n12946), .ZN(n12560) );
  INV_X1 U10920 ( .A(n11787), .ZN(n12558) );
  INV_X1 U10921 ( .A(n12946), .ZN(n11866) );
  OR2_X1 U10922 ( .A1(n11954), .A2(n11866), .ZN(n8292) );
  XNOR2_X1 U10923 ( .A(n10838), .B(P2_DATAO_REG_11__SCAN_IN), .ZN(n8293) );
  XNOR2_X1 U10924 ( .A(n8294), .B(n8293), .ZN(n10634) );
  NAND2_X1 U10925 ( .A1(n10634), .A2(n12422), .ZN(n8299) );
  OAI21_X1 U10926 ( .B1(n8295), .B2(P3_IR_REG_10__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n8297) );
  INV_X1 U10927 ( .A(P3_IR_REG_11__SCAN_IN), .ZN(n8296) );
  XNOR2_X1 U10928 ( .A(n8297), .B(n8296), .ZN(n12975) );
  AOI22_X1 U10929 ( .A1(n8415), .A2(n12975), .B1(n12410), .B2(n10633), .ZN(
        n8298) );
  NAND2_X1 U10930 ( .A1(n8517), .A2(P3_REG0_REG_11__SCAN_IN), .ZN(n8306) );
  NAND2_X1 U10931 ( .A1(n8534), .A2(P3_REG1_REG_11__SCAN_IN), .ZN(n8305) );
  OR2_X1 U10932 ( .A1(n8301), .A2(n8300), .ZN(n8302) );
  NAND2_X1 U10933 ( .A1(n8319), .A2(n8302), .ZN(n12178) );
  NAND2_X1 U10934 ( .A1(n8466), .A2(n12178), .ZN(n8304) );
  NAND2_X1 U10935 ( .A1(n8492), .A2(P3_REG2_REG_11__SCAN_IN), .ZN(n8303) );
  NAND4_X1 U10936 ( .A1(n8306), .A2(n8305), .A3(n8304), .A4(n8303), .ZN(n12945) );
  INV_X1 U10937 ( .A(n12945), .ZN(n12120) );
  NAND2_X1 U10938 ( .A1(n13411), .A2(n12120), .ZN(n8307) );
  NAND2_X1 U10939 ( .A1(n11947), .A2(n8307), .ZN(n8309) );
  OR2_X1 U10940 ( .A1(n13411), .A2(n12120), .ZN(n8308) );
  XNOR2_X1 U10941 ( .A(n8311), .B(n8310), .ZN(n10652) );
  NAND2_X1 U10942 ( .A1(n10652), .A2(n8514), .ZN(n8318) );
  OR2_X1 U10943 ( .A1(n8313), .A2(n8312), .ZN(n8370) );
  NAND2_X1 U10944 ( .A1(n8370), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8314) );
  MUX2_X1 U10945 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8314), .S(
        P3_IR_REG_12__SCAN_IN), .Z(n8316) );
  NOR2_X1 U10946 ( .A1(n8370), .A2(P3_IR_REG_12__SCAN_IN), .ZN(n8342) );
  INV_X1 U10947 ( .A(n8342), .ZN(n8315) );
  NAND2_X1 U10948 ( .A1(n8316), .A2(n8315), .ZN(n13008) );
  INV_X1 U10949 ( .A(n13008), .ZN(n12998) );
  AOI22_X1 U10950 ( .A1(n12423), .A2(SI_12_), .B1(n8415), .B2(n12998), .ZN(
        n8317) );
  NAND2_X1 U10951 ( .A1(n8318), .A2(n8317), .ZN(n12116) );
  NAND2_X1 U10952 ( .A1(n8517), .A2(P3_REG0_REG_12__SCAN_IN), .ZN(n8324) );
  NAND2_X1 U10953 ( .A1(n12398), .A2(P3_REG1_REG_12__SCAN_IN), .ZN(n8323) );
  NAND2_X1 U10954 ( .A1(n8319), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n8320) );
  NAND2_X1 U10955 ( .A1(n8335), .A2(n8320), .ZN(n12240) );
  NAND2_X1 U10956 ( .A1(n8521), .A2(n12240), .ZN(n8322) );
  NAND2_X1 U10957 ( .A1(n8492), .A2(P3_REG2_REG_12__SCAN_IN), .ZN(n8321) );
  OR2_X1 U10958 ( .A1(n12116), .A2(n12216), .ZN(n12571) );
  NAND2_X1 U10959 ( .A1(n12116), .A2(n12216), .ZN(n12567) );
  INV_X1 U10960 ( .A(n12216), .ZN(n12944) );
  NAND2_X1 U10961 ( .A1(n12116), .A2(n12944), .ZN(n8325) );
  NAND2_X1 U10962 ( .A1(n8327), .A2(n8326), .ZN(n8329) );
  XNOR2_X1 U10963 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(P2_DATAO_REG_13__SCAN_IN), 
        .ZN(n8328) );
  XNOR2_X1 U10964 ( .A(n8329), .B(n8328), .ZN(n10661) );
  NAND2_X1 U10965 ( .A1(n10661), .A2(n12422), .ZN(n8332) );
  OR2_X1 U10966 ( .A1(n8342), .A2(n13504), .ZN(n8330) );
  INV_X1 U10967 ( .A(P3_IR_REG_13__SCAN_IN), .ZN(n8341) );
  XNOR2_X1 U10968 ( .A(n8330), .B(n8341), .ZN(n13027) );
  AOI22_X1 U10969 ( .A1(n12423), .A2(n10660), .B1(n8415), .B2(n13027), .ZN(
        n8331) );
  INV_X1 U10970 ( .A(P3_REG2_REG_13__SCAN_IN), .ZN(n12995) );
  NAND2_X1 U10971 ( .A1(n8517), .A2(P3_REG0_REG_13__SCAN_IN), .ZN(n8334) );
  NAND2_X1 U10972 ( .A1(n12398), .A2(P3_REG1_REG_13__SCAN_IN), .ZN(n8333) );
  AND2_X1 U10973 ( .A1(n8334), .A2(n8333), .ZN(n8338) );
  AND2_X1 U10974 ( .A1(n8335), .A2(P3_REG3_REG_13__SCAN_IN), .ZN(n8336) );
  OR2_X1 U10975 ( .A1(n8336), .A2(n8347), .ZN(n12225) );
  NAND2_X1 U10976 ( .A1(n12225), .A2(n8466), .ZN(n8337) );
  OAI211_X1 U10977 ( .C1(n8287), .C2(n12995), .A(n8338), .B(n8337), .ZN(n13338) );
  NOR2_X1 U10978 ( .A1(n12218), .A2(n13338), .ZN(n8600) );
  INV_X1 U10979 ( .A(n8600), .ZN(n12479) );
  NAND2_X1 U10980 ( .A1(n12218), .A2(n13338), .ZN(n12484) );
  INV_X1 U10981 ( .A(n13338), .ZN(n12238) );
  XNOR2_X1 U10982 ( .A(n8340), .B(n8339), .ZN(n10663) );
  NAND2_X1 U10983 ( .A1(n10663), .A2(n12422), .ZN(n8345) );
  AND2_X1 U10984 ( .A1(n8342), .A2(n8341), .ZN(n8355) );
  OR2_X1 U10985 ( .A1(n8355), .A2(n13504), .ZN(n8343) );
  INV_X1 U10986 ( .A(P3_IR_REG_14__SCAN_IN), .ZN(n8354) );
  XNOR2_X1 U10987 ( .A(n8343), .B(n8354), .ZN(n13042) );
  AOI22_X1 U10988 ( .A1(n12423), .A2(n10662), .B1(n8415), .B2(n13042), .ZN(
        n8344) );
  INV_X1 U10989 ( .A(n8517), .ZN(n8480) );
  INV_X1 U10990 ( .A(P3_REG0_REG_14__SCAN_IN), .ZN(n13492) );
  NOR2_X1 U10991 ( .A1(n8347), .A2(n8346), .ZN(n8348) );
  OR2_X1 U10992 ( .A1(n8361), .A2(n8348), .ZN(n13344) );
  NAND2_X1 U10993 ( .A1(n13344), .A2(n8466), .ZN(n8350) );
  AOI22_X1 U10994 ( .A1(n8534), .A2(P3_REG1_REG_14__SCAN_IN), .B1(n8492), .B2(
        P3_REG2_REG_14__SCAN_IN), .ZN(n8349) );
  OAI211_X1 U10995 ( .C1(n8480), .C2(n13492), .A(n8350), .B(n8349), .ZN(n13327) );
  OR2_X1 U10996 ( .A1(n13494), .A2(n13327), .ZN(n12481) );
  NAND2_X1 U10997 ( .A1(n12481), .A2(n6547), .ZN(n13334) );
  INV_X1 U10998 ( .A(n13327), .ZN(n12777) );
  OR2_X1 U10999 ( .A1(n13494), .A2(n12777), .ZN(n8351) );
  XNOR2_X1 U11000 ( .A(n8353), .B(n8352), .ZN(n10739) );
  NAND2_X1 U11001 ( .A1(n10739), .A2(n8514), .ZN(n8359) );
  INV_X1 U11002 ( .A(SI_15_), .ZN(n10738) );
  NAND2_X1 U11003 ( .A1(n8355), .A2(n8354), .ZN(n8368) );
  NAND2_X1 U11004 ( .A1(n8368), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8357) );
  INV_X1 U11005 ( .A(P3_IR_REG_15__SCAN_IN), .ZN(n8356) );
  XNOR2_X1 U11006 ( .A(n8357), .B(n8356), .ZN(n13063) );
  AOI22_X1 U11007 ( .A1(n12423), .A2(n10738), .B1(n13063), .B2(n8415), .ZN(
        n8358) );
  INV_X1 U11008 ( .A(P3_REG2_REG_15__SCAN_IN), .ZN(n13330) );
  OR2_X1 U11009 ( .A1(n8361), .A2(n8360), .ZN(n8362) );
  NAND2_X1 U11010 ( .A1(n8377), .A2(n8362), .ZN(n13320) );
  NAND2_X1 U11011 ( .A1(n13320), .A2(n8521), .ZN(n8364) );
  AOI22_X1 U11012 ( .A1(n8517), .A2(P3_REG0_REG_15__SCAN_IN), .B1(n12398), 
        .B2(P3_REG1_REG_15__SCAN_IN), .ZN(n8363) );
  OAI211_X1 U11013 ( .C1(n8287), .C2(n13330), .A(n8364), .B(n8363), .ZN(n13341) );
  INV_X1 U11014 ( .A(n13341), .ZN(n12858) );
  NOR2_X1 U11015 ( .A1(n13491), .A2(n12858), .ZN(n8365) );
  XNOR2_X1 U11016 ( .A(n8367), .B(n8366), .ZN(n10891) );
  NAND2_X1 U11017 ( .A1(n10891), .A2(n12422), .ZN(n8376) );
  OAI21_X1 U11018 ( .B1(n8368), .B2(P3_IR_REG_15__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n8369) );
  MUX2_X1 U11019 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8369), .S(
        P3_IR_REG_16__SCAN_IN), .Z(n8373) );
  INV_X1 U11020 ( .A(n8370), .ZN(n8372) );
  NAND2_X1 U11021 ( .A1(n8372), .A2(n8371), .ZN(n8387) );
  AOI22_X1 U11022 ( .A1(n13088), .A2(n8415), .B1(n12410), .B2(SI_16_), .ZN(
        n8375) );
  NAND2_X1 U11023 ( .A1(n8377), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n8378) );
  NAND2_X1 U11024 ( .A1(n8392), .A2(n8378), .ZN(n13309) );
  NAND2_X1 U11025 ( .A1(n13309), .A2(n8521), .ZN(n8381) );
  AOI22_X1 U11026 ( .A1(n8517), .A2(P3_REG0_REG_16__SCAN_IN), .B1(n8534), .B2(
        P3_REG1_REG_16__SCAN_IN), .ZN(n8380) );
  NAND2_X1 U11027 ( .A1(n8492), .A2(P3_REG2_REG_16__SCAN_IN), .ZN(n8379) );
  NAND2_X1 U11028 ( .A1(n13481), .A2(n13328), .ZN(n8383) );
  XNOR2_X1 U11029 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(P2_DATAO_REG_17__SCAN_IN), 
        .ZN(n8385) );
  XNOR2_X1 U11030 ( .A(n8386), .B(n8385), .ZN(n11056) );
  NAND2_X1 U11031 ( .A1(n11056), .A2(n12422), .ZN(n8391) );
  NAND2_X1 U11032 ( .A1(n8387), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8389) );
  INV_X1 U11033 ( .A(P3_IR_REG_17__SCAN_IN), .ZN(n8388) );
  XNOR2_X1 U11034 ( .A(n8389), .B(n8388), .ZN(n13112) );
  AOI22_X1 U11035 ( .A1(n12423), .A2(n11055), .B1(n8415), .B2(n13112), .ZN(
        n8390) );
  NAND2_X1 U11036 ( .A1(n8392), .A2(P3_REG3_REG_17__SCAN_IN), .ZN(n8393) );
  NAND2_X1 U11037 ( .A1(n8406), .A2(n8393), .ZN(n13298) );
  NAND2_X1 U11038 ( .A1(n13298), .A2(n8466), .ZN(n8398) );
  INV_X1 U11039 ( .A(P3_REG0_REG_17__SCAN_IN), .ZN(n13474) );
  NAND2_X1 U11040 ( .A1(n12399), .A2(P3_REG2_REG_17__SCAN_IN), .ZN(n8395) );
  NAND2_X1 U11041 ( .A1(n8534), .A2(P3_REG1_REG_17__SCAN_IN), .ZN(n8394) );
  OAI211_X1 U11042 ( .C1(n8480), .C2(n13474), .A(n8395), .B(n8394), .ZN(n8396)
         );
  INV_X1 U11043 ( .A(n8396), .ZN(n8397) );
  NAND2_X1 U11044 ( .A1(n13477), .A2(n13313), .ZN(n12475) );
  INV_X1 U11045 ( .A(n13301), .ZN(n12584) );
  INV_X1 U11046 ( .A(n13313), .ZN(n12782) );
  OR2_X1 U11047 ( .A1(n13477), .A2(n12782), .ZN(n8399) );
  INV_X1 U11048 ( .A(n8400), .ZN(n8401) );
  XNOR2_X1 U11049 ( .A(n8402), .B(n8401), .ZN(n11276) );
  NAND2_X1 U11050 ( .A1(n11276), .A2(n8514), .ZN(n8405) );
  XNOR2_X1 U11051 ( .A(n8403), .B(P3_IR_REG_18__SCAN_IN), .ZN(n13132) );
  AOI22_X1 U11052 ( .A1(n12423), .A2(SI_18_), .B1(n8415), .B2(n13132), .ZN(
        n8404) );
  INV_X1 U11053 ( .A(n8419), .ZN(n8408) );
  NAND2_X1 U11054 ( .A1(n8406), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n8407) );
  NAND2_X1 U11055 ( .A1(n8408), .A2(n8407), .ZN(n13293) );
  INV_X1 U11056 ( .A(P3_REG0_REG_18__SCAN_IN), .ZN(n9432) );
  NAND2_X1 U11057 ( .A1(n12399), .A2(P3_REG2_REG_18__SCAN_IN), .ZN(n8410) );
  NAND2_X1 U11058 ( .A1(n12398), .A2(P3_REG1_REG_18__SCAN_IN), .ZN(n8409) );
  OAI211_X1 U11059 ( .C1(n8480), .C2(n9432), .A(n8410), .B(n8409), .ZN(n8411)
         );
  NAND2_X1 U11060 ( .A1(n13469), .A2(n12869), .ZN(n12474) );
  XNOR2_X1 U11061 ( .A(n8413), .B(n8412), .ZN(n11529) );
  NAND2_X1 U11062 ( .A1(n11529), .A2(n8514), .ZN(n8417) );
  AOI22_X1 U11063 ( .A1(n12423), .A2(SI_19_), .B1(n6525), .B2(n8415), .ZN(
        n8416) );
  OR2_X1 U11064 ( .A1(n8419), .A2(n8418), .ZN(n8420) );
  NAND2_X1 U11065 ( .A1(n8431), .A2(n8420), .ZN(n13281) );
  INV_X1 U11066 ( .A(P3_REG0_REG_19__SCAN_IN), .ZN(n9348) );
  NAND2_X1 U11067 ( .A1(n8492), .A2(P3_REG2_REG_19__SCAN_IN), .ZN(n8422) );
  NAND2_X1 U11068 ( .A1(n12398), .A2(P3_REG1_REG_19__SCAN_IN), .ZN(n8421) );
  OAI211_X1 U11069 ( .C1(n8480), .C2(n9348), .A(n8422), .B(n8421), .ZN(n8423)
         );
  NAND2_X1 U11070 ( .A1(n13384), .A2(n13290), .ZN(n8424) );
  OR2_X1 U11071 ( .A1(n13384), .A2(n13290), .ZN(n8425) );
  XNOR2_X1 U11072 ( .A(n8428), .B(n8427), .ZN(n11750) );
  NAND2_X1 U11073 ( .A1(n11750), .A2(n8514), .ZN(n8430) );
  NAND2_X1 U11074 ( .A1(n12410), .A2(SI_20_), .ZN(n8429) );
  NAND2_X1 U11075 ( .A1(n8431), .A2(P3_REG3_REG_20__SCAN_IN), .ZN(n8432) );
  NAND2_X1 U11076 ( .A1(n8444), .A2(n8432), .ZN(n13261) );
  NAND2_X1 U11077 ( .A1(n13261), .A2(n8466), .ZN(n8438) );
  INV_X1 U11078 ( .A(P3_REG2_REG_20__SCAN_IN), .ZN(n8435) );
  NAND2_X1 U11079 ( .A1(n8517), .A2(P3_REG0_REG_20__SCAN_IN), .ZN(n8434) );
  NAND2_X1 U11080 ( .A1(n8534), .A2(P3_REG1_REG_20__SCAN_IN), .ZN(n8433) );
  OAI211_X1 U11081 ( .C1(n8435), .C2(n8287), .A(n8434), .B(n8433), .ZN(n8436)
         );
  INV_X1 U11082 ( .A(n8436), .ZN(n8437) );
  NAND2_X1 U11083 ( .A1(n13381), .A2(n13247), .ZN(n12473) );
  NAND2_X1 U11084 ( .A1(n12472), .A2(n12473), .ZN(n8604) );
  NAND2_X1 U11085 ( .A1(n13381), .A2(n13276), .ZN(n8439) );
  XNOR2_X1 U11086 ( .A(n8441), .B(n8440), .ZN(n11881) );
  NAND2_X1 U11087 ( .A1(n11881), .A2(n12422), .ZN(n8443) );
  NAND2_X1 U11088 ( .A1(n12410), .A2(SI_21_), .ZN(n8442) );
  AND2_X1 U11089 ( .A1(n8444), .A2(P3_REG3_REG_21__SCAN_IN), .ZN(n8445) );
  OR2_X1 U11090 ( .A1(n8445), .A2(n8454), .ZN(n13250) );
  INV_X1 U11091 ( .A(P3_REG2_REG_21__SCAN_IN), .ZN(n13249) );
  NAND2_X1 U11092 ( .A1(n8517), .A2(P3_REG0_REG_21__SCAN_IN), .ZN(n8447) );
  NAND2_X1 U11093 ( .A1(n8197), .A2(P3_REG1_REG_21__SCAN_IN), .ZN(n8446) );
  OAI211_X1 U11094 ( .C1(n13249), .C2(n8287), .A(n8447), .B(n8446), .ZN(n8448)
         );
  OR2_X1 U11095 ( .A1(n13251), .A2(n13233), .ZN(n8449) );
  XNOR2_X1 U11096 ( .A(n8451), .B(n8450), .ZN(n11919) );
  NAND2_X1 U11097 ( .A1(n11919), .A2(n8514), .ZN(n8453) );
  NAND2_X1 U11098 ( .A1(n12410), .A2(SI_22_), .ZN(n8452) );
  OR2_X1 U11099 ( .A1(n8454), .A2(n12896), .ZN(n8455) );
  NAND2_X1 U11100 ( .A1(n8475), .A2(n8455), .ZN(n13237) );
  NAND2_X1 U11101 ( .A1(n13237), .A2(n8466), .ZN(n8460) );
  INV_X1 U11102 ( .A(P3_REG0_REG_22__SCAN_IN), .ZN(n13450) );
  NAND2_X1 U11103 ( .A1(n12399), .A2(P3_REG2_REG_22__SCAN_IN), .ZN(n8457) );
  NAND2_X1 U11104 ( .A1(n8534), .A2(P3_REG1_REG_22__SCAN_IN), .ZN(n8456) );
  OAI211_X1 U11105 ( .C1(n8480), .C2(n13450), .A(n8457), .B(n8456), .ZN(n8458)
         );
  INV_X1 U11106 ( .A(n8458), .ZN(n8459) );
  NAND2_X1 U11107 ( .A1(n13451), .A2(n12942), .ZN(n8461) );
  XNOR2_X1 U11108 ( .A(n8462), .B(P1_DATAO_REG_24__SCAN_IN), .ZN(n12292) );
  NAND2_X1 U11109 ( .A1(n12292), .A2(n8514), .ZN(n8464) );
  NAND2_X1 U11110 ( .A1(n12410), .A2(SI_24_), .ZN(n8463) );
  NAND2_X1 U11111 ( .A1(n12398), .A2(P3_REG1_REG_24__SCAN_IN), .ZN(n8470) );
  NAND2_X1 U11112 ( .A1(n12399), .A2(P3_REG2_REG_24__SCAN_IN), .ZN(n8469) );
  NAND2_X1 U11113 ( .A1(P3_REG3_REG_24__SCAN_IN), .A2(n8476), .ZN(n8465) );
  NAND2_X1 U11114 ( .A1(n8465), .A2(n6575), .ZN(n13213) );
  NAND2_X1 U11115 ( .A1(n8466), .A2(n13213), .ZN(n8468) );
  NAND2_X1 U11116 ( .A1(n8517), .A2(P3_REG0_REG_24__SCAN_IN), .ZN(n8467) );
  OR2_X1 U11117 ( .A1(n13212), .A2(n13220), .ZN(n12465) );
  NAND2_X1 U11118 ( .A1(n13212), .A2(n13220), .ZN(n12466) );
  NAND2_X1 U11119 ( .A1(n12465), .A2(n12466), .ZN(n12441) );
  XNOR2_X1 U11120 ( .A(n8472), .B(n8471), .ZN(n12082) );
  NAND2_X1 U11121 ( .A1(n12082), .A2(n8514), .ZN(n8474) );
  NAND2_X1 U11122 ( .A1(n12410), .A2(SI_23_), .ZN(n8473) );
  NAND2_X1 U11123 ( .A1(n8475), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n8477) );
  NAND2_X1 U11124 ( .A1(n8477), .A2(n8476), .ZN(n13226) );
  NAND2_X1 U11125 ( .A1(n13226), .A2(n8466), .ZN(n8483) );
  INV_X1 U11126 ( .A(P3_REG0_REG_23__SCAN_IN), .ZN(n13446) );
  NAND2_X1 U11127 ( .A1(n8492), .A2(P3_REG2_REG_23__SCAN_IN), .ZN(n8479) );
  NAND2_X1 U11128 ( .A1(n12398), .A2(P3_REG1_REG_23__SCAN_IN), .ZN(n8478) );
  OAI211_X1 U11129 ( .C1(n8480), .C2(n13446), .A(n8479), .B(n8478), .ZN(n8481)
         );
  INV_X1 U11130 ( .A(n8481), .ZN(n8482) );
  NAND2_X1 U11131 ( .A1(n13225), .A2(n12897), .ZN(n12597) );
  AND2_X1 U11132 ( .A1(n13225), .A2(n13234), .ZN(n13205) );
  AOI22_X1 U11133 ( .A1(n12441), .A2(n13205), .B1(n12941), .B2(n13212), .ZN(
        n8484) );
  OAI21_X1 U11134 ( .B1(n8487), .B2(n8486), .A(n8485), .ZN(n13526) );
  OR2_X1 U11135 ( .A1(n13526), .A2(n8488), .ZN(n8490) );
  NAND2_X1 U11136 ( .A1(n12410), .A2(SI_25_), .ZN(n8489) );
  NAND2_X1 U11137 ( .A1(n8197), .A2(P3_REG1_REG_25__SCAN_IN), .ZN(n8496) );
  NAND2_X1 U11138 ( .A1(n8517), .A2(P3_REG0_REG_25__SCAN_IN), .ZN(n8495) );
  NAND2_X1 U11139 ( .A1(P3_REG3_REG_25__SCAN_IN), .A2(n6575), .ZN(n8491) );
  NAND2_X1 U11140 ( .A1(n8491), .A2(n8502), .ZN(n13200) );
  NAND2_X1 U11141 ( .A1(n8521), .A2(n13200), .ZN(n8494) );
  NAND2_X1 U11142 ( .A1(n8492), .A2(P3_REG2_REG_25__SCAN_IN), .ZN(n8493) );
  NAND4_X1 U11143 ( .A1(n8496), .A2(n8495), .A3(n8494), .A4(n8493), .ZN(n13207) );
  NAND2_X1 U11144 ( .A1(n13440), .A2(n13207), .ZN(n12464) );
  NAND2_X1 U11145 ( .A1(n12851), .A2(n13180), .ZN(n12463) );
  INV_X1 U11146 ( .A(n13198), .ZN(n13193) );
  NAND2_X1 U11147 ( .A1(n12851), .A2(n13207), .ZN(n8497) );
  NAND2_X1 U11148 ( .A1(n13520), .A2(n12422), .ZN(n8501) );
  NAND2_X1 U11149 ( .A1(n12410), .A2(SI_26_), .ZN(n8500) );
  NAND2_X1 U11150 ( .A1(n8517), .A2(P3_REG0_REG_26__SCAN_IN), .ZN(n8508) );
  NAND2_X1 U11151 ( .A1(n8534), .A2(P3_REG1_REG_26__SCAN_IN), .ZN(n8507) );
  NAND2_X1 U11152 ( .A1(P3_REG3_REG_26__SCAN_IN), .A2(n8502), .ZN(n8504) );
  INV_X1 U11153 ( .A(n8503), .ZN(n8518) );
  NAND2_X1 U11154 ( .A1(n8504), .A2(n8518), .ZN(n13186) );
  NAND2_X1 U11155 ( .A1(n8466), .A2(n13186), .ZN(n8506) );
  NAND2_X1 U11156 ( .A1(n8492), .A2(P3_REG2_REG_26__SCAN_IN), .ZN(n8505) );
  OR2_X1 U11157 ( .A1(n12920), .A2(n13170), .ZN(n8511) );
  NAND2_X1 U11158 ( .A1(n12920), .A2(n13196), .ZN(n12608) );
  OR2_X1 U11159 ( .A1(n13185), .A2(n13436), .ZN(n8509) );
  INV_X1 U11160 ( .A(n8509), .ZN(n8510) );
  XNOR2_X1 U11161 ( .A(n8513), .B(n8512), .ZN(n13516) );
  NAND2_X1 U11162 ( .A1(n13516), .A2(n8514), .ZN(n8516) );
  NAND2_X1 U11163 ( .A1(n12410), .A2(SI_27_), .ZN(n8515) );
  NAND2_X1 U11164 ( .A1(n8517), .A2(P3_REG0_REG_27__SCAN_IN), .ZN(n8525) );
  NAND2_X1 U11165 ( .A1(n8197), .A2(P3_REG1_REG_27__SCAN_IN), .ZN(n8524) );
  NAND2_X1 U11166 ( .A1(P3_REG3_REG_27__SCAN_IN), .A2(n8518), .ZN(n8519) );
  NAND2_X1 U11167 ( .A1(n12399), .A2(P3_REG2_REG_27__SCAN_IN), .ZN(n8522) );
  NAND2_X1 U11168 ( .A1(n13358), .A2(n13181), .ZN(n8611) );
  NAND2_X1 U11169 ( .A1(n12611), .A2(n8611), .ZN(n13167) );
  NAND2_X1 U11170 ( .A1(n8526), .A2(n12807), .ZN(n12616) );
  NAND2_X1 U11171 ( .A1(n13428), .A2(n13169), .ZN(n12620) );
  OR2_X1 U11172 ( .A1(n13358), .A2(n12940), .ZN(n13152) );
  AND2_X1 U11173 ( .A1(n13150), .A2(n13152), .ZN(n8527) );
  NAND2_X1 U11174 ( .A1(n13166), .A2(n8527), .ZN(n13155) );
  INV_X1 U11175 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n15530) );
  NAND2_X1 U11176 ( .A1(n15530), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n12407) );
  INV_X1 U11177 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n14454) );
  NAND2_X1 U11178 ( .A1(n14454), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n8530) );
  NAND2_X1 U11179 ( .A1(n12407), .A2(n8530), .ZN(n12404) );
  NAND2_X1 U11180 ( .A1(n13509), .A2(n12422), .ZN(n8532) );
  NAND2_X1 U11181 ( .A1(n12410), .A2(SI_29_), .ZN(n8531) );
  INV_X1 U11182 ( .A(n8633), .ZN(n8533) );
  NAND2_X1 U11183 ( .A1(n8466), .A2(n8533), .ZN(n12403) );
  NAND2_X1 U11184 ( .A1(n8534), .A2(P3_REG1_REG_29__SCAN_IN), .ZN(n8537) );
  NAND2_X1 U11185 ( .A1(n12399), .A2(P3_REG2_REG_29__SCAN_IN), .ZN(n8536) );
  NAND2_X1 U11186 ( .A1(n8517), .A2(P3_REG0_REG_29__SCAN_IN), .ZN(n8535) );
  NAND2_X1 U11187 ( .A1(n8539), .A2(n7332), .ZN(n8542) );
  NAND2_X1 U11188 ( .A1(n8542), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8538) );
  NAND2_X1 U11189 ( .A1(n8540), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8541) );
  AND2_X1 U11190 ( .A1(n12493), .A2(n10705), .ZN(n12429) );
  INV_X1 U11191 ( .A(n12429), .ZN(n8544) );
  NAND2_X1 U11192 ( .A1(n12644), .A2(n6525), .ZN(n10706) );
  AND2_X4 U11193 ( .A1(n12644), .A2(n12493), .ZN(n12626) );
  INV_X1 U11194 ( .A(n13515), .ZN(n12641) );
  NAND2_X1 U11195 ( .A1(n12641), .A2(n13122), .ZN(n10900) );
  NAND2_X1 U11196 ( .A1(n10900), .A2(n10897), .ZN(n10734) );
  INV_X1 U11197 ( .A(n10734), .ZN(n10777) );
  NAND2_X1 U11198 ( .A1(n12626), .A2(n10777), .ZN(n13265) );
  NAND2_X1 U11199 ( .A1(n8517), .A2(P3_REG0_REG_30__SCAN_IN), .ZN(n8547) );
  NAND2_X1 U11200 ( .A1(n8197), .A2(P3_REG1_REG_30__SCAN_IN), .ZN(n8546) );
  NAND2_X1 U11201 ( .A1(n12399), .A2(P3_REG2_REG_30__SCAN_IN), .ZN(n8545) );
  NAND2_X1 U11202 ( .A1(n12641), .A2(P3_B_REG_SCAN_IN), .ZN(n8548) );
  NAND2_X1 U11203 ( .A1(n13340), .A2(n8548), .ZN(n13143) );
  OAI22_X1 U11204 ( .A1(n12807), .A2(n13265), .B1(n12427), .B2(n13143), .ZN(
        n8549) );
  INV_X1 U11205 ( .A(P3_REG1_REG_29__SCAN_IN), .ZN(n8588) );
  NAND3_X1 U11206 ( .A1(n8551), .A2(n8550), .A3(n7329), .ZN(n8552) );
  NAND2_X1 U11207 ( .A1(n8555), .A2(n8554), .ZN(n8559) );
  INV_X1 U11208 ( .A(n8579), .ZN(n13529) );
  INV_X1 U11209 ( .A(P3_B_REG_SCAN_IN), .ZN(n8557) );
  XNOR2_X1 U11210 ( .A(n8561), .B(n8557), .ZN(n8558) );
  OR2_X1 U11211 ( .A1(n13519), .A2(n8561), .ZN(n8562) );
  OR2_X1 U11212 ( .A1(n13519), .A2(n8579), .ZN(n8563) );
  XNOR2_X1 U11213 ( .A(n10707), .B(n10709), .ZN(n8582) );
  NOR2_X1 U11214 ( .A1(P3_D_REG_18__SCAN_IN), .A2(P3_D_REG_17__SCAN_IN), .ZN(
        n8568) );
  NOR4_X1 U11215 ( .A1(P3_D_REG_2__SCAN_IN), .A2(P3_D_REG_8__SCAN_IN), .A3(
        P3_D_REG_22__SCAN_IN), .A4(P3_D_REG_25__SCAN_IN), .ZN(n8567) );
  NOR4_X1 U11216 ( .A1(P3_D_REG_29__SCAN_IN), .A2(P3_D_REG_10__SCAN_IN), .A3(
        P3_D_REG_31__SCAN_IN), .A4(P3_D_REG_14__SCAN_IN), .ZN(n8566) );
  NOR4_X1 U11217 ( .A1(P3_D_REG_20__SCAN_IN), .A2(P3_D_REG_19__SCAN_IN), .A3(
        P3_D_REG_27__SCAN_IN), .A4(P3_D_REG_24__SCAN_IN), .ZN(n8565) );
  NAND4_X1 U11218 ( .A1(n8568), .A2(n8567), .A3(n8566), .A4(n8565), .ZN(n8574)
         );
  NOR4_X1 U11219 ( .A1(P3_D_REG_9__SCAN_IN), .A2(P3_D_REG_16__SCAN_IN), .A3(
        P3_D_REG_15__SCAN_IN), .A4(P3_D_REG_30__SCAN_IN), .ZN(n8572) );
  NOR4_X1 U11220 ( .A1(P3_D_REG_11__SCAN_IN), .A2(P3_D_REG_21__SCAN_IN), .A3(
        P3_D_REG_12__SCAN_IN), .A4(P3_D_REG_26__SCAN_IN), .ZN(n8571) );
  NOR4_X1 U11221 ( .A1(P3_D_REG_3__SCAN_IN), .A2(P3_D_REG_5__SCAN_IN), .A3(
        P3_D_REG_4__SCAN_IN), .A4(P3_D_REG_7__SCAN_IN), .ZN(n8570) );
  NOR4_X1 U11222 ( .A1(P3_D_REG_13__SCAN_IN), .A2(P3_D_REG_28__SCAN_IN), .A3(
        P3_D_REG_23__SCAN_IN), .A4(P3_D_REG_6__SCAN_IN), .ZN(n8569) );
  NAND4_X1 U11223 ( .A1(n8572), .A2(n8571), .A3(n8570), .A4(n8569), .ZN(n8573)
         );
  NOR2_X1 U11224 ( .A1(n8574), .A2(n8573), .ZN(n8575) );
  NOR2_X1 U11225 ( .A1(n10621), .A2(n8575), .ZN(n10708) );
  OAI21_X1 U11226 ( .B1(n8576), .B2(P3_IR_REG_22__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n8578) );
  INV_X1 U11227 ( .A(P3_IR_REG_23__SCAN_IN), .ZN(n8577) );
  XNOR2_X1 U11228 ( .A(n8578), .B(n8577), .ZN(n10896) );
  NAND2_X1 U11229 ( .A1(n10896), .A2(P3_STATE_REG_SCAN_IN), .ZN(n10548) );
  AND2_X1 U11230 ( .A1(n8579), .A2(n8561), .ZN(n8580) );
  NOR2_X1 U11231 ( .A1(n10708), .A2(n10895), .ZN(n8581) );
  OAI22_X1 U11232 ( .A1(n15946), .A2(n10705), .B1(n6525), .B2(n8618), .ZN(
        n8583) );
  AOI21_X1 U11233 ( .B1(n8583), .B2(n7331), .A(n12626), .ZN(n8586) );
  NAND3_X1 U11234 ( .A1(n12644), .A2(n10705), .A3(n13128), .ZN(n8584) );
  NAND2_X1 U11235 ( .A1(n12598), .A2(n8584), .ZN(n8624) );
  NAND2_X1 U11236 ( .A1(n12626), .A2(n7331), .ZN(n10714) );
  NAND2_X1 U11237 ( .A1(n8624), .A2(n10714), .ZN(n8623) );
  INV_X1 U11238 ( .A(n8623), .ZN(n8585) );
  MUX2_X1 U11239 ( .A(n8586), .B(n8585), .S(n10709), .Z(n8587) );
  NAND2_X1 U11240 ( .A1(n10730), .A2(n12495), .ZN(n10785) );
  NAND2_X1 U11241 ( .A1(n10785), .A2(n12496), .ZN(n11336) );
  NAND2_X1 U11242 ( .A1(n11336), .A2(n12501), .ZN(n8589) );
  INV_X1 U11243 ( .A(n8590), .ZN(n12520) );
  OAI21_X1 U11244 ( .B1(n12520), .B2(n12512), .A(n12518), .ZN(n8591) );
  INV_X1 U11245 ( .A(n8591), .ZN(n8592) );
  NAND2_X1 U11246 ( .A1(n11437), .A2(n12532), .ZN(n11696) );
  INV_X1 U11247 ( .A(n11760), .ZN(n12535) );
  NAND2_X1 U11248 ( .A1(n11696), .A2(n12535), .ZN(n8595) );
  NAND2_X1 U11249 ( .A1(n11401), .A2(n12450), .ZN(n8596) );
  NAND2_X1 U11250 ( .A1(n12551), .A2(n12947), .ZN(n8597) );
  XNOR2_X1 U11251 ( .A(n13411), .B(n12945), .ZN(n12565) );
  OR2_X1 U11252 ( .A1(n13411), .A2(n12945), .ZN(n12566) );
  NAND2_X1 U11253 ( .A1(n12059), .A2(n12453), .ZN(n8599) );
  NAND2_X1 U11254 ( .A1(n8601), .A2(n12481), .ZN(n13319) );
  OR2_X1 U11255 ( .A1(n13491), .A2(n13341), .ZN(n12480) );
  NAND2_X1 U11256 ( .A1(n13491), .A2(n13341), .ZN(n12486) );
  NAND2_X1 U11257 ( .A1(n13319), .A2(n13325), .ZN(n13318) );
  OR2_X1 U11258 ( .A1(n13481), .A2(n12932), .ZN(n12583) );
  NAND2_X1 U11259 ( .A1(n13481), .A2(n12932), .ZN(n12580) );
  NAND2_X1 U11260 ( .A1(n13308), .A2(n12443), .ZN(n8602) );
  NAND2_X1 U11261 ( .A1(n13297), .A2(n13301), .ZN(n13254) );
  NAND2_X1 U11262 ( .A1(n12587), .A2(n13255), .ZN(n8606) );
  INV_X1 U11263 ( .A(n13286), .ZN(n8603) );
  NAND2_X1 U11264 ( .A1(n13384), .A2(n13266), .ZN(n13258) );
  NAND2_X1 U11265 ( .A1(n13251), .A2(n13268), .ZN(n12471) );
  OR2_X1 U11266 ( .A1(n12493), .A2(n10705), .ZN(n8613) );
  XNOR2_X1 U11267 ( .A(n12644), .B(n8613), .ZN(n8615) );
  OR2_X1 U11268 ( .A1(n12493), .A2(n6525), .ZN(n8614) );
  NAND2_X1 U11269 ( .A1(n8615), .A2(n8614), .ZN(n10711) );
  NAND2_X1 U11270 ( .A1(n10711), .A2(n15946), .ZN(n10724) );
  MUX2_X1 U11271 ( .A(n10724), .B(n8618), .S(n10705), .Z(n8616) );
  INV_X1 U11272 ( .A(n8616), .ZN(n8617) );
  NAND2_X1 U11273 ( .A1(n8617), .A2(n13128), .ZN(n15957) );
  NAND2_X1 U11274 ( .A1(n11753), .A2(n6525), .ZN(n12636) );
  NAND2_X1 U11275 ( .A1(n8618), .A2(n10731), .ZN(n15956) );
  NAND2_X1 U11276 ( .A1(n15973), .A2(n13407), .ZN(n13406) );
  NAND2_X1 U11277 ( .A1(n13423), .A2(n13395), .ZN(n8619) );
  INV_X1 U11278 ( .A(n8620), .ZN(n8621) );
  NAND2_X1 U11279 ( .A1(n8622), .A2(n8621), .ZN(P3_U3488) );
  INV_X1 U11280 ( .A(P3_REG2_REG_29__SCAN_IN), .ZN(n8629) );
  INV_X1 U11281 ( .A(n10709), .ZN(n10704) );
  NAND2_X1 U11282 ( .A1(n8623), .A2(n10704), .ZN(n8626) );
  NAND2_X1 U11283 ( .A1(n10709), .A2(n8624), .ZN(n8625) );
  AND2_X1 U11284 ( .A1(n8626), .A2(n8625), .ZN(n8627) );
  NAND2_X1 U11285 ( .A1(n8628), .A2(n8627), .ZN(n8631) );
  NOR2_X1 U11286 ( .A1(n10895), .A2(n15946), .ZN(n10732) );
  NAND2_X1 U11287 ( .A1(n10731), .A2(n12493), .ZN(n11337) );
  NAND2_X1 U11288 ( .A1(n15957), .A2(n11337), .ZN(n8630) );
  INV_X1 U11289 ( .A(n8631), .ZN(n8632) );
  AND2_X1 U11290 ( .A1(n15960), .A2(n12636), .ZN(n11366) );
  NOR2_X1 U11291 ( .A1(n13321), .A2(n8633), .ZN(n13145) );
  AOI21_X1 U11292 ( .B1(n13423), .B2(n13310), .A(n13145), .ZN(n8634) );
  NOR2_X1 U11293 ( .A1(P1_IR_REG_12__SCAN_IN), .A2(P1_IR_REG_8__SCAN_IN), .ZN(
        n8636) );
  INV_X2 U11294 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n8850) );
  NOR2_X1 U11295 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(P1_IR_REG_19__SCAN_IN), 
        .ZN(n8640) );
  NOR2_X1 U11296 ( .A1(P1_IR_REG_21__SCAN_IN), .A2(P1_IR_REG_23__SCAN_IN), 
        .ZN(n8639) );
  NAND4_X1 U11297 ( .A1(n8640), .A2(n8639), .A3(n9361), .A4(n9201), .ZN(n9207)
         );
  NOR2_X2 U11298 ( .A1(P1_IR_REG_17__SCAN_IN), .A2(P1_IR_REG_16__SCAN_IN), 
        .ZN(n8996) );
  INV_X1 U11299 ( .A(n8646), .ZN(n15525) );
  NAND2_X1 U11300 ( .A1(n8647), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8648) );
  MUX2_X1 U11301 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8648), .S(
        P1_IR_REG_29__SCAN_IN), .Z(n8649) );
  NAND2_X1 U11302 ( .A1(n8980), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n8653) );
  INV_X1 U11303 ( .A(n15532), .ZN(n8650) );
  OR2_X2 U11304 ( .A1(n8654), .A2(n8650), .ZN(n8693) );
  INV_X1 U11305 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n8651) );
  OR2_X1 U11306 ( .A1(n8693), .A2(n8651), .ZN(n8652) );
  NAND2_X1 U11307 ( .A1(n14835), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n8657) );
  INV_X1 U11308 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n8655) );
  OR2_X1 U11309 ( .A1(n14834), .A2(n8655), .ZN(n8656) );
  INV_X1 U11310 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n15717) );
  INV_X1 U11311 ( .A(SI_0_), .ZN(n8659) );
  OAI21_X1 U11312 ( .B1(n6532), .B2(n8659), .A(n8658), .ZN(n8660) );
  NAND2_X1 U11313 ( .A1(n8669), .A2(n8660), .ZN(n15553) );
  MUX2_X1 U11314 ( .A(n15717), .B(n15553), .S(n9089), .Z(n11371) );
  INV_X1 U11315 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n10753) );
  OR2_X1 U11316 ( .A1(n14834), .A2(n10753), .ZN(n8668) );
  INV_X1 U11317 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n8663) );
  OR2_X1 U11318 ( .A1(n8693), .A2(n8663), .ZN(n8667) );
  INV_X1 U11319 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n8664) );
  NAND2_X1 U11320 ( .A1(n8980), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n8665) );
  NAND4_X1 U11321 ( .A1(n8666), .A2(n8667), .A3(n8668), .A4(n8665), .ZN(n10289) );
  INV_X1 U11322 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n10577) );
  OR2_X1 U11323 ( .A1(n6535), .A2(n10577), .ZN(n8678) );
  INV_X1 U11324 ( .A(SI_1_), .ZN(n10598) );
  XNOR2_X1 U11325 ( .A(n8682), .B(n10598), .ZN(n8671) );
  MUX2_X1 U11326 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(P1_DATAO_REG_1__SCAN_IN), 
        .S(n6532), .Z(n8670) );
  MUX2_X1 U11327 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8672), .S(
        P1_IR_REG_1__SCAN_IN), .Z(n8675) );
  INV_X1 U11328 ( .A(n8673), .ZN(n8674) );
  OR2_X1 U11329 ( .A1(n9089), .A2(n10752), .ZN(n8676) );
  AND3_X4 U11330 ( .A1(n8677), .A2(n8678), .A3(n8676), .ZN(n15783) );
  NAND2_X1 U11331 ( .A1(n10289), .A2(n15783), .ZN(n9141) );
  INV_X2 U11332 ( .A(n10289), .ZN(n10294) );
  NAND2_X1 U11333 ( .A1(n6533), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n8680) );
  OAI211_X1 U11334 ( .C1(n6532), .C2(n10577), .A(n8680), .B(n10598), .ZN(n8681) );
  NAND2_X1 U11335 ( .A1(n8682), .A2(n8681), .ZN(n8685) );
  NAND2_X1 U11336 ( .A1(n6533), .A2(n10573), .ZN(n8683) );
  OAI211_X1 U11337 ( .C1(P2_DATAO_REG_1__SCAN_IN), .C2(n6532), .A(n8683), .B(
        SI_1_), .ZN(n8684) );
  XNOR2_X1 U11338 ( .A(n8698), .B(n8699), .ZN(n10592) );
  INV_X1 U11339 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n11692) );
  NAND2_X1 U11340 ( .A1(n8778), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n8689) );
  INV_X1 U11341 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n8686) );
  INV_X1 U11342 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n14986) );
  OR2_X1 U11343 ( .A1(n8692), .A2(n14986), .ZN(n8687) );
  NAND2_X1 U11344 ( .A1(n11637), .A2(n14923), .ZN(n8691) );
  NAND2_X1 U11345 ( .A1(n14709), .A2(n14708), .ZN(n14693) );
  OR2_X1 U11347 ( .A1(n8692), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n8696) );
  INV_X1 U11348 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n8694) );
  INV_X1 U11349 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n11525) );
  OR2_X1 U11350 ( .A1(n14834), .A2(n11525), .ZN(n8695) );
  NAND2_X1 U11351 ( .A1(n8699), .A2(n8698), .ZN(n8702) );
  NAND2_X1 U11352 ( .A1(n8700), .A2(SI_2_), .ZN(n8701) );
  OR2_X1 U11353 ( .A1(n8724), .A2(n10576), .ZN(n8711) );
  NOR2_X1 U11354 ( .A1(n8704), .A2(n8645), .ZN(n8705) );
  MUX2_X1 U11355 ( .A(n8645), .B(n8705), .S(P1_IR_REG_3__SCAN_IN), .Z(n8706)
         );
  INV_X1 U11356 ( .A(n8706), .ZN(n8709) );
  INV_X1 U11357 ( .A(n8707), .ZN(n8708) );
  NAND2_X1 U11358 ( .A1(n8709), .A2(n8708), .ZN(n10872) );
  OR2_X1 U11359 ( .A1(n9089), .A2(n10872), .ZN(n8710) );
  INV_X4 U11360 ( .A(n8980), .ZN(n12754) );
  OAI21_X1 U11361 ( .B1(P1_REG3_REG_3__SCAN_IN), .B2(P1_REG3_REG_4__SCAN_IN), 
        .A(n8732), .ZN(n11724) );
  OR2_X1 U11362 ( .A1(n12754), .A2(n11724), .ZN(n8716) );
  NAND2_X1 U11363 ( .A1(n14835), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n8715) );
  INV_X1 U11364 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n10759) );
  OR2_X1 U11365 ( .A1(n14834), .A2(n10759), .ZN(n8714) );
  INV_X1 U11366 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n8712) );
  OR2_X1 U11367 ( .A1(n14839), .A2(n8712), .ZN(n8713) );
  INV_X1 U11368 ( .A(n8718), .ZN(n8719) );
  NAND2_X1 U11369 ( .A1(n8719), .A2(SI_3_), .ZN(n8720) );
  XNOR2_X1 U11370 ( .A(n8741), .B(SI_4_), .ZN(n8738) );
  XNOR2_X1 U11371 ( .A(n8740), .B(n8738), .ZN(n10588) );
  NAND2_X1 U11372 ( .A1(n8743), .A2(n10588), .ZN(n8727) );
  OR2_X1 U11373 ( .A1(n8707), .A2(n8645), .ZN(n8723) );
  XNOR2_X1 U11374 ( .A(n8723), .B(n8722), .ZN(n15010) );
  OR2_X1 U11375 ( .A1(n9089), .A2(n15010), .ZN(n8726) );
  OR2_X1 U11376 ( .A1(n8724), .A2(n10589), .ZN(n8725) );
  XNOR2_X1 U11377 ( .A(n14970), .B(n11283), .ZN(n14926) );
  NAND2_X1 U11378 ( .A1(n14970), .A2(n11283), .ZN(n8728) );
  NAND2_X1 U11379 ( .A1(n10533), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n8737) );
  INV_X1 U11380 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n8729) );
  OR2_X1 U11381 ( .A1(n14839), .A2(n8729), .ZN(n8736) );
  INV_X1 U11382 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n8731) );
  NAND2_X1 U11383 ( .A1(n8732), .A2(n8731), .ZN(n8733) );
  NAND2_X1 U11384 ( .A1(n8762), .A2(n8733), .ZN(n11884) );
  OR2_X1 U11385 ( .A1(n12754), .A2(n11884), .ZN(n8735) );
  INV_X1 U11386 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n10747) );
  INV_X1 U11387 ( .A(n8738), .ZN(n8739) );
  INV_X1 U11388 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n10620) );
  MUX2_X1 U11389 ( .A(n10618), .B(n10620), .S(n6533), .Z(n8752) );
  XNOR2_X1 U11390 ( .A(n8752), .B(SI_5_), .ZN(n8750) );
  INV_X1 U11391 ( .A(n8750), .ZN(n8742) );
  XNOR2_X1 U11392 ( .A(n8751), .B(n8742), .ZN(n10617) );
  NAND2_X1 U11393 ( .A1(n10617), .A2(n8743), .ZN(n8747) );
  INV_X2 U11394 ( .A(n8724), .ZN(n9031) );
  NAND2_X1 U11395 ( .A1(n8997), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8744) );
  MUX2_X1 U11396 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8744), .S(
        P1_IR_REG_5__SCAN_IN), .Z(n8745) );
  AND2_X1 U11397 ( .A1(n8745), .A2(n8756), .ZN(n10822) );
  AOI22_X1 U11398 ( .A1(n9031), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n10629), 
        .B2(n10822), .ZN(n8746) );
  INV_X1 U11399 ( .A(n14725), .ZN(n11885) );
  NAND2_X1 U11400 ( .A1(n14969), .A2(n11885), .ZN(n8748) );
  INV_X1 U11401 ( .A(n8752), .ZN(n8753) );
  NAND2_X1 U11402 ( .A1(n8753), .A2(SI_5_), .ZN(n8754) );
  MUX2_X1 U11403 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(P1_DATAO_REG_6__SCAN_IN), 
        .S(n6532), .Z(n8774) );
  NAND2_X1 U11404 ( .A1(n10624), .A2(n8743), .ZN(n8760) );
  NAND2_X1 U11405 ( .A1(n8756), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8755) );
  NAND2_X1 U11406 ( .A1(n8758), .A2(n8794), .ZN(n10832) );
  INV_X1 U11407 ( .A(n10832), .ZN(n10843) );
  AOI22_X1 U11408 ( .A1(n9031), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n10629), 
        .B2(n10843), .ZN(n8759) );
  INV_X1 U11409 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n11843) );
  NAND2_X1 U11410 ( .A1(n8762), .A2(n11843), .ZN(n8763) );
  NAND2_X1 U11411 ( .A1(n8779), .A2(n8763), .ZN(n11860) );
  OR2_X1 U11412 ( .A1(n12754), .A2(n11860), .ZN(n8768) );
  NAND2_X1 U11413 ( .A1(n14835), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n8767) );
  INV_X1 U11414 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n11859) );
  OR2_X1 U11415 ( .A1(n14834), .A2(n11859), .ZN(n8766) );
  INV_X1 U11416 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n8764) );
  OR2_X1 U11417 ( .A1(n14839), .A2(n8764), .ZN(n8765) );
  NAND4_X1 U11418 ( .A1(n8768), .A2(n8767), .A3(n8766), .A4(n8765), .ZN(n14968) );
  NAND2_X1 U11419 ( .A1(n7943), .A2(n14968), .ZN(n8769) );
  MUX2_X1 U11420 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(P1_DATAO_REG_7__SCAN_IN), 
        .S(n6532), .Z(n8789) );
  XNOR2_X1 U11421 ( .A(n8788), .B(n8786), .ZN(n10635) );
  NAND2_X1 U11422 ( .A1(n10635), .A2(n8743), .ZN(n8777) );
  NAND2_X1 U11423 ( .A1(n8794), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8775) );
  XNOR2_X1 U11424 ( .A(n8775), .B(P1_IR_REG_7__SCAN_IN), .ZN(n11148) );
  AOI22_X1 U11425 ( .A1(n9031), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n10629), 
        .B2(n11148), .ZN(n8776) );
  NAND2_X2 U11426 ( .A1(n8777), .A2(n8776), .ZN(n14733) );
  NAND2_X1 U11427 ( .A1(n10490), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n8784) );
  INV_X1 U11428 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n12158) );
  OR2_X1 U11429 ( .A1(n14834), .A2(n12158), .ZN(n8783) );
  NAND2_X1 U11430 ( .A1(n8779), .A2(n9414), .ZN(n8780) );
  NAND2_X1 U11431 ( .A1(n8812), .A2(n8780), .ZN(n14480) );
  OR2_X1 U11432 ( .A1(n12754), .A2(n14480), .ZN(n8782) );
  INV_X1 U11433 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n10840) );
  OR2_X1 U11434 ( .A1(n10536), .A2(n10840), .ZN(n8781) );
  OR2_X1 U11435 ( .A1(n14733), .A2(n14550), .ZN(n8785) );
  NAND2_X1 U11436 ( .A1(n8789), .A2(SI_7_), .ZN(n8790) );
  NAND2_X1 U11437 ( .A1(n10664), .A2(n8743), .ZN(n8799) );
  INV_X1 U11438 ( .A(n8794), .ZN(n8796) );
  NAND2_X1 U11439 ( .A1(n8796), .A2(n8795), .ZN(n8852) );
  NAND2_X1 U11440 ( .A1(n8852), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8808) );
  INV_X1 U11441 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n8849) );
  NAND2_X1 U11442 ( .A1(n8808), .A2(n8849), .ZN(n8797) );
  NAND2_X1 U11443 ( .A1(n8797), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8831) );
  XNOR2_X1 U11444 ( .A(n8831), .B(P1_IR_REG_9__SCAN_IN), .ZN(n11231) );
  AOI22_X1 U11445 ( .A1(n9031), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n11231), 
        .B2(n10629), .ZN(n8798) );
  NAND2_X1 U11446 ( .A1(n10490), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n8805) );
  INV_X1 U11447 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n12258) );
  OR2_X1 U11448 ( .A1(n10536), .A2(n12258), .ZN(n8804) );
  NAND2_X1 U11449 ( .A1(n8814), .A2(n8800), .ZN(n8801) );
  NAND2_X1 U11450 ( .A1(n8836), .A2(n8801), .ZN(n14617) );
  OR2_X1 U11451 ( .A1(n12754), .A2(n14617), .ZN(n8803) );
  INV_X1 U11452 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n11151) );
  OR2_X1 U11453 ( .A1(n14834), .A2(n11151), .ZN(n8802) );
  XNOR2_X1 U11454 ( .A(n8807), .B(n8806), .ZN(n10655) );
  NAND2_X1 U11455 ( .A1(n10655), .A2(n8743), .ZN(n8810) );
  XNOR2_X1 U11456 ( .A(n8808), .B(P1_IR_REG_8__SCAN_IN), .ZN(n15030) );
  AOI22_X1 U11457 ( .A1(n9031), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n10629), 
        .B2(n15030), .ZN(n8809) );
  NAND2_X2 U11458 ( .A1(n8810), .A2(n8809), .ZN(n14737) );
  NAND2_X1 U11459 ( .A1(n10490), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n8818) );
  INV_X1 U11460 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n11906) );
  OR2_X1 U11461 ( .A1(n14834), .A2(n11906), .ZN(n8817) );
  NAND2_X1 U11462 ( .A1(n8812), .A2(n8811), .ZN(n8813) );
  NAND2_X1 U11463 ( .A1(n8814), .A2(n8813), .ZN(n14549) );
  OR2_X1 U11464 ( .A1(n12754), .A2(n14549), .ZN(n8816) );
  INV_X1 U11465 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n11147) );
  OR2_X1 U11466 ( .A1(n10536), .A2(n11147), .ZN(n8815) );
  OR2_X1 U11467 ( .A1(n14737), .A2(n14618), .ZN(n12244) );
  OAI21_X1 U11468 ( .B1(n14742), .B2(n14513), .A(n12244), .ZN(n8819) );
  INV_X1 U11469 ( .A(n8819), .ZN(n8820) );
  NAND2_X1 U11470 ( .A1(n11912), .A2(n8820), .ZN(n8825) );
  NAND2_X1 U11471 ( .A1(n14737), .A2(n14618), .ZN(n8821) );
  NAND2_X1 U11472 ( .A1(n8821), .A2(n15800), .ZN(n8823) );
  INV_X1 U11473 ( .A(n14618), .ZN(n14967) );
  NOR2_X1 U11474 ( .A1(n14967), .A2(n15800), .ZN(n8822) );
  AOI22_X1 U11475 ( .A1(n14742), .A2(n8823), .B1(n8822), .B2(n14737), .ZN(
        n8824) );
  XNOR2_X1 U11476 ( .A(n8844), .B(n8843), .ZN(n10773) );
  NAND2_X1 U11477 ( .A1(n8831), .A2(n8830), .ZN(n8832) );
  NAND2_X1 U11478 ( .A1(n8832), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8833) );
  XNOR2_X1 U11479 ( .A(n8833), .B(P1_IR_REG_10__SCAN_IN), .ZN(n11239) );
  AOI22_X1 U11480 ( .A1(n11239), .A2(n10629), .B1(n9031), .B2(
        P2_DATAO_REG_10__SCAN_IN), .ZN(n8834) );
  NAND2_X1 U11481 ( .A1(n10490), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n8841) );
  INV_X1 U11482 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n8835) );
  OR2_X1 U11483 ( .A1(n14834), .A2(n8835), .ZN(n8840) );
  INV_X1 U11484 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n14511) );
  NAND2_X1 U11485 ( .A1(n8836), .A2(n14511), .ZN(n8837) );
  NAND2_X1 U11486 ( .A1(n8857), .A2(n8837), .ZN(n14512) );
  OR2_X1 U11487 ( .A1(n12754), .A2(n14512), .ZN(n8839) );
  INV_X1 U11488 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n11478) );
  OR2_X1 U11489 ( .A1(n10536), .A2(n11478), .ZN(n8838) );
  INV_X1 U11490 ( .A(n8846), .ZN(n8847) );
  NAND2_X1 U11491 ( .A1(n8847), .A2(SI_11_), .ZN(n8848) );
  XNOR2_X1 U11492 ( .A(n8866), .B(n8865), .ZN(n10835) );
  NAND2_X1 U11493 ( .A1(n10835), .A2(n8743), .ZN(n8855) );
  NAND2_X1 U11494 ( .A1(n8850), .A2(n8849), .ZN(n8851) );
  NAND2_X1 U11495 ( .A1(n8873), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8853) );
  XNOR2_X1 U11496 ( .A(n8853), .B(P1_IR_REG_11__SCAN_IN), .ZN(n11483) );
  AOI22_X1 U11497 ( .A1(n9031), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n10629), 
        .B2(n11483), .ZN(n8854) );
  NAND2_X1 U11498 ( .A1(n8857), .A2(n8856), .ZN(n8858) );
  NAND2_X1 U11499 ( .A1(n8877), .A2(n8858), .ZN(n14657) );
  OR2_X1 U11500 ( .A1(n12754), .A2(n14657), .ZN(n8863) );
  NAND2_X1 U11501 ( .A1(n14835), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n8862) );
  INV_X1 U11502 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n8859) );
  OR2_X1 U11503 ( .A1(n14839), .A2(n8859), .ZN(n8861) );
  INV_X1 U11504 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n12205) );
  OR2_X1 U11505 ( .A1(n14834), .A2(n12205), .ZN(n8860) );
  NAND4_X1 U11506 ( .A1(n8863), .A2(n8862), .A3(n8861), .A4(n8860), .ZN(n15478) );
  XNOR2_X1 U11507 ( .A(n15490), .B(n15478), .ZN(n14934) );
  INV_X1 U11508 ( .A(n15478), .ZN(n14574) );
  OR2_X1 U11509 ( .A1(n15490), .A2(n14574), .ZN(n8864) );
  INV_X1 U11510 ( .A(n8869), .ZN(n8870) );
  NAND2_X1 U11511 ( .A1(n8870), .A2(SI_12_), .ZN(n8925) );
  AND2_X1 U11512 ( .A1(n8903), .A2(n8925), .ZN(n8871) );
  XNOR2_X1 U11513 ( .A(n8886), .B(P1_IR_REG_12__SCAN_IN), .ZN(n15732) );
  AOI22_X1 U11514 ( .A1(n15732), .A2(n10629), .B1(n9031), .B2(
        P2_DATAO_REG_12__SCAN_IN), .ZN(n8874) );
  NAND2_X1 U11515 ( .A1(n10490), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n8882) );
  INV_X1 U11516 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n12268) );
  OR2_X1 U11517 ( .A1(n14834), .A2(n12268), .ZN(n8881) );
  INV_X1 U11518 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n8876) );
  NAND2_X1 U11519 ( .A1(n8877), .A2(n8876), .ZN(n8878) );
  NAND2_X1 U11520 ( .A1(n8892), .A2(n8878), .ZN(n14573) );
  OR2_X1 U11521 ( .A1(n12754), .A2(n14573), .ZN(n8880) );
  INV_X1 U11522 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n9451) );
  OR2_X1 U11523 ( .A1(n10536), .A2(n9451), .ZN(n8879) );
  NAND2_X1 U11524 ( .A1(n15480), .A2(n15466), .ZN(n14758) );
  XNOR2_X1 U11525 ( .A(n8902), .B(SI_13_), .ZN(n8883) );
  INV_X1 U11526 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n8885) );
  NAND2_X1 U11527 ( .A1(n8886), .A2(n8885), .ZN(n8887) );
  NAND2_X1 U11528 ( .A1(n8887), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8909) );
  XNOR2_X1 U11529 ( .A(n8909), .B(P1_IR_REG_13__SCAN_IN), .ZN(n12136) );
  AOI22_X1 U11530 ( .A1(n12136), .A2(n10629), .B1(n9031), .B2(
        P2_DATAO_REG_13__SCAN_IN), .ZN(n8888) );
  NAND2_X1 U11531 ( .A1(n10490), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n8897) );
  INV_X1 U11532 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n8890) );
  OR2_X1 U11533 ( .A1(n10536), .A2(n8890), .ZN(n8896) );
  NAND2_X1 U11534 ( .A1(n8892), .A2(n8891), .ZN(n8893) );
  NAND2_X1 U11535 ( .A1(n8915), .A2(n8893), .ZN(n14634) );
  OR2_X1 U11536 ( .A1(n12754), .A2(n14634), .ZN(n8895) );
  INV_X1 U11537 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n12317) );
  OR2_X1 U11538 ( .A1(n14834), .A2(n12317), .ZN(n8894) );
  NAND2_X1 U11539 ( .A1(n15471), .A2(n14572), .ZN(n14771) );
  INV_X1 U11540 ( .A(n8902), .ZN(n8898) );
  NAND2_X1 U11541 ( .A1(n8926), .A2(SI_14_), .ZN(n8906) );
  INV_X1 U11542 ( .A(n8906), .ZN(n8901) );
  OAI21_X1 U11543 ( .B1(SI_14_), .B2(n10660), .A(n8898), .ZN(n8900) );
  OAI21_X1 U11544 ( .B1(SI_13_), .B2(n10662), .A(n8902), .ZN(n8899) );
  AOI22_X1 U11545 ( .A1(n8901), .A2(n8927), .B1(n8900), .B2(n8899), .ZN(n8905)
         );
  NAND2_X1 U11546 ( .A1(n8902), .A2(n10660), .ZN(n8928) );
  NAND2_X1 U11547 ( .A1(n11446), .A2(n8743), .ZN(n8913) );
  INV_X1 U11548 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n8908) );
  NAND2_X1 U11549 ( .A1(n8909), .A2(n8908), .ZN(n8910) );
  NAND2_X1 U11550 ( .A1(n8910), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8911) );
  XNOR2_X1 U11551 ( .A(n8911), .B(P1_IR_REG_14__SCAN_IN), .ZN(n15036) );
  AOI22_X1 U11552 ( .A1(n15036), .A2(n10629), .B1(n9031), .B2(
        P2_DATAO_REG_14__SCAN_IN), .ZN(n8912) );
  NAND2_X1 U11553 ( .A1(n10490), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n8920) );
  INV_X1 U11554 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n15041) );
  OR2_X1 U11555 ( .A1(n14834), .A2(n15041), .ZN(n8919) );
  INV_X1 U11556 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n8914) );
  NAND2_X1 U11557 ( .A1(n8915), .A2(n8914), .ZN(n8916) );
  NAND2_X1 U11558 ( .A1(n8945), .A2(n8916), .ZN(n14489) );
  OR2_X1 U11559 ( .A1(n12754), .A2(n14489), .ZN(n8918) );
  INV_X1 U11560 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n12134) );
  OR2_X1 U11561 ( .A1(n10536), .A2(n12134), .ZN(n8917) );
  NAND2_X1 U11562 ( .A1(n14772), .A2(n15468), .ZN(n8921) );
  OR2_X1 U11563 ( .A1(n14772), .A2(n15468), .ZN(n8922) );
  NAND2_X1 U11564 ( .A1(n8923), .A2(n8922), .ZN(n15323) );
  NAND2_X1 U11565 ( .A1(n8924), .A2(n8959), .ZN(n8933) );
  NAND2_X1 U11566 ( .A1(n8926), .A2(n8925), .ZN(n8954) );
  INV_X1 U11567 ( .A(n8954), .ZN(n8930) );
  AOI21_X1 U11568 ( .B1(n8958), .B2(n8930), .A(n8957), .ZN(n8931) );
  NAND2_X1 U11569 ( .A1(n8934), .A2(SI_15_), .ZN(n8963) );
  INV_X1 U11570 ( .A(n8934), .ZN(n8935) );
  NAND2_X1 U11571 ( .A1(n8935), .A2(n10738), .ZN(n8961) );
  AND2_X1 U11572 ( .A1(n8963), .A2(n8961), .ZN(n8936) );
  OR2_X1 U11573 ( .A1(n8997), .A2(n8939), .ZN(n8970) );
  NAND2_X1 U11574 ( .A1(n8970), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8940) );
  XNOR2_X1 U11575 ( .A(n8940), .B(P1_IR_REG_15__SCAN_IN), .ZN(n15743) );
  AOI22_X1 U11576 ( .A1(n9031), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n10629), 
        .B2(n15743), .ZN(n8941) );
  INV_X1 U11577 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n8944) );
  NAND2_X1 U11578 ( .A1(n8945), .A2(n8944), .ZN(n8946) );
  NAND2_X1 U11579 ( .A1(n8978), .A2(n8946), .ZN(n15330) );
  OR2_X1 U11580 ( .A1(n15330), .A2(n12754), .ZN(n8950) );
  NAND2_X1 U11581 ( .A1(n10533), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n8949) );
  NAND2_X1 U11582 ( .A1(n10490), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n8948) );
  NAND2_X1 U11583 ( .A1(n14835), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n8947) );
  NAND4_X1 U11584 ( .A1(n8950), .A2(n8949), .A3(n8948), .A4(n8947), .ZN(n15458) );
  NAND2_X1 U11585 ( .A1(n15323), .A2(n15324), .ZN(n8952) );
  INV_X1 U11586 ( .A(n15458), .ZN(n15310) );
  OR2_X1 U11587 ( .A1(n15325), .A2(n15310), .ZN(n8951) );
  NAND2_X1 U11588 ( .A1(n8952), .A2(n8951), .ZN(n15307) );
  INV_X1 U11589 ( .A(n8957), .ZN(n8955) );
  OAI21_X1 U11590 ( .B1(n8959), .B2(n10662), .A(n8963), .ZN(n8953) );
  INV_X1 U11591 ( .A(n8959), .ZN(n8960) );
  NOR2_X1 U11592 ( .A1(n8960), .A2(SI_14_), .ZN(n8964) );
  INV_X1 U11593 ( .A(n8961), .ZN(n8962) );
  NAND2_X1 U11594 ( .A1(n8966), .A2(n8965), .ZN(n8987) );
  INV_X1 U11595 ( .A(n8967), .ZN(n8968) );
  NAND2_X1 U11596 ( .A1(n8968), .A2(SI_16_), .ZN(n8969) );
  XNOR2_X1 U11597 ( .A(n8987), .B(n8034), .ZN(n11291) );
  NOR2_X1 U11598 ( .A1(n8970), .A2(P1_IR_REG_15__SCAN_IN), .ZN(n8974) );
  INV_X1 U11599 ( .A(n8974), .ZN(n8971) );
  NAND2_X1 U11600 ( .A1(n8971), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8972) );
  MUX2_X1 U11601 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8972), .S(
        P1_IR_REG_16__SCAN_IN), .Z(n8975) );
  INV_X1 U11602 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n8973) );
  NAND2_X1 U11603 ( .A1(n8974), .A2(n8973), .ZN(n8993) );
  AOI22_X1 U11604 ( .A1(n9031), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n10629), 
        .B2(n15059), .ZN(n8976) );
  INV_X1 U11605 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n8977) );
  NAND2_X1 U11606 ( .A1(n8978), .A2(n8977), .ZN(n8979) );
  AND2_X1 U11607 ( .A1(n9001), .A2(n8979), .ZN(n15315) );
  NAND2_X1 U11608 ( .A1(n15315), .A2(n8980), .ZN(n8983) );
  AOI22_X1 U11609 ( .A1(n10490), .A2(P1_REG0_REG_16__SCAN_IN), .B1(n10533), 
        .B2(P1_REG2_REG_16__SCAN_IN), .ZN(n8982) );
  NAND2_X1 U11610 ( .A1(n14835), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n8981) );
  NAND2_X1 U11611 ( .A1(n15444), .A2(n15434), .ZN(n8986) );
  OR2_X1 U11612 ( .A1(n15444), .A2(n15434), .ZN(n8984) );
  NAND2_X1 U11613 ( .A1(n8987), .A2(n8034), .ZN(n8989) );
  INV_X1 U11614 ( .A(n8990), .ZN(n8991) );
  NAND2_X1 U11615 ( .A1(n8991), .A2(SI_17_), .ZN(n8992) );
  NAND2_X1 U11616 ( .A1(n11404), .A2(n8743), .ZN(n9000) );
  NAND2_X1 U11617 ( .A1(n8993), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8994) );
  MUX2_X1 U11618 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8994), .S(
        P1_IR_REG_17__SCAN_IN), .Z(n8998) );
  AND2_X1 U11619 ( .A1(n8998), .A2(n7308), .ZN(n15078) );
  AOI22_X1 U11620 ( .A1(n9031), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n10629), 
        .B2(n15078), .ZN(n8999) );
  INV_X1 U11621 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n9415) );
  NAND2_X1 U11622 ( .A1(n9001), .A2(n9415), .ZN(n9002) );
  NAND2_X1 U11623 ( .A1(n9014), .A2(n9002), .ZN(n15293) );
  OR2_X1 U11624 ( .A1(n15293), .A2(n12754), .ZN(n9005) );
  AOI22_X1 U11625 ( .A1(n10490), .A2(P1_REG0_REG_17__SCAN_IN), .B1(n10533), 
        .B2(P1_REG2_REG_17__SCAN_IN), .ZN(n9004) );
  NAND2_X1 U11626 ( .A1(n14835), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n9003) );
  NAND2_X1 U11627 ( .A1(n15438), .A2(n15311), .ZN(n14780) );
  NAND2_X2 U11628 ( .A1(n9007), .A2(n9006), .ZN(n9009) );
  XNOR2_X1 U11629 ( .A(n9024), .B(n9043), .ZN(n11754) );
  NAND2_X1 U11630 ( .A1(n11754), .A2(n8743), .ZN(n9012) );
  NAND2_X1 U11631 ( .A1(n7308), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9010) );
  XNOR2_X1 U11632 ( .A(n9010), .B(P1_IR_REG_18__SCAN_IN), .ZN(n15093) );
  AOI22_X1 U11633 ( .A1(n9031), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n10629), 
        .B2(n15093), .ZN(n9011) );
  NAND2_X2 U11634 ( .A1(n9012), .A2(n9011), .ZN(n15284) );
  INV_X1 U11635 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n9013) );
  NAND2_X1 U11636 ( .A1(n9014), .A2(n9013), .ZN(n9015) );
  NAND2_X1 U11637 ( .A1(n9035), .A2(n9015), .ZN(n15275) );
  OR2_X1 U11638 ( .A1(n15275), .A2(n12754), .ZN(n9020) );
  INV_X1 U11639 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n15080) );
  NAND2_X1 U11640 ( .A1(n10533), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n9017) );
  NAND2_X1 U11641 ( .A1(n10490), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n9016) );
  OAI211_X1 U11642 ( .C1(n15080), .C2(n10536), .A(n9017), .B(n9016), .ZN(n9018) );
  INV_X1 U11643 ( .A(n9018), .ZN(n9019) );
  OR2_X1 U11644 ( .A1(n15284), .A2(n15435), .ZN(n9023) );
  NAND2_X1 U11645 ( .A1(n9024), .A2(n9045), .ZN(n9026) );
  INV_X1 U11646 ( .A(SI_18_), .ZN(n11277) );
  OR2_X1 U11647 ( .A1(n9050), .A2(n11277), .ZN(n9025) );
  XNOR2_X1 U11648 ( .A(n9046), .B(SI_19_), .ZN(n9027) );
  INV_X1 U11649 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n9030) );
  AOI22_X1 U11650 ( .A1(n9031), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n15103), 
        .B2(n10629), .ZN(n9032) );
  INV_X1 U11651 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n9034) );
  OR2_X2 U11652 ( .A1(n9035), .A2(n9034), .ZN(n9053) );
  NAND2_X1 U11653 ( .A1(n9035), .A2(n9034), .ZN(n9036) );
  AND2_X1 U11654 ( .A1(n9053), .A2(n9036), .ZN(n15253) );
  NAND2_X1 U11655 ( .A1(n15253), .A2(n8980), .ZN(n9041) );
  INV_X1 U11656 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n15090) );
  NAND2_X1 U11657 ( .A1(n10533), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n9038) );
  NAND2_X1 U11658 ( .A1(n10490), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n9037) );
  OAI211_X1 U11659 ( .C1(n15090), .C2(n10536), .A(n9038), .B(n9037), .ZN(n9039) );
  INV_X1 U11660 ( .A(n9039), .ZN(n9040) );
  NAND2_X1 U11661 ( .A1(n15252), .A2(n15409), .ZN(n9042) );
  OAI22_X1 U11662 ( .A1(n9045), .A2(SI_18_), .B1(n9046), .B2(SI_19_), .ZN(
        n9049) );
  INV_X1 U11663 ( .A(SI_19_), .ZN(n11531) );
  OAI21_X1 U11664 ( .B1(n9043), .B2(n11277), .A(n11531), .ZN(n9047) );
  AND2_X1 U11665 ( .A1(SI_18_), .A2(SI_19_), .ZN(n9044) );
  AOI22_X1 U11666 ( .A1(n9047), .A2(n9046), .B1(n9045), .B2(n9044), .ZN(n9048)
         );
  INV_X1 U11667 ( .A(SI_20_), .ZN(n11752) );
  NAND2_X1 U11668 ( .A1(n11961), .A2(n8743), .ZN(n9052) );
  OR2_X1 U11669 ( .A1(n8724), .A2(n11963), .ZN(n9051) );
  INV_X1 U11670 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n14626) );
  NAND2_X1 U11671 ( .A1(n9053), .A2(n14626), .ZN(n9054) );
  AND2_X1 U11672 ( .A1(n9069), .A2(n9054), .ZN(n15239) );
  NAND2_X1 U11673 ( .A1(n15239), .A2(n8980), .ZN(n9060) );
  INV_X1 U11674 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n9057) );
  NAND2_X1 U11675 ( .A1(n10533), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n9056) );
  NAND2_X1 U11676 ( .A1(n10490), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n9055) );
  OAI211_X1 U11677 ( .C1(n9057), .C2(n10536), .A(n9056), .B(n9055), .ZN(n9058)
         );
  INV_X1 U11678 ( .A(n9058), .ZN(n9059) );
  XNOR2_X1 U11679 ( .A(n15413), .B(n15401), .ZN(n14945) );
  OR2_X1 U11680 ( .A1(n15413), .A2(n15401), .ZN(n9061) );
  NAND2_X1 U11681 ( .A1(n9062), .A2(n9082), .ZN(n9064) );
  NAND2_X1 U11682 ( .A1(n9081), .A2(SI_20_), .ZN(n9063) );
  NAND2_X1 U11683 ( .A1(n9064), .A2(n9063), .ZN(n9066) );
  MUX2_X1 U11684 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(P1_DATAO_REG_21__SCAN_IN), 
        .S(n6532), .Z(n9084) );
  XNOR2_X1 U11685 ( .A(n9084), .B(SI_21_), .ZN(n9065) );
  OR2_X1 U11686 ( .A1(n8724), .A2(n12051), .ZN(n9067) );
  INV_X1 U11687 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n14565) );
  NAND2_X1 U11688 ( .A1(n9069), .A2(n14565), .ZN(n9070) );
  NAND2_X1 U11689 ( .A1(n9090), .A2(n9070), .ZN(n15227) );
  INV_X1 U11690 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n9073) );
  NAND2_X1 U11691 ( .A1(n10533), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n9072) );
  NAND2_X1 U11692 ( .A1(n10490), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n9071) );
  OAI211_X1 U11693 ( .C1(n9073), .C2(n10536), .A(n9072), .B(n9071), .ZN(n9074)
         );
  INV_X1 U11694 ( .A(n9074), .ZN(n9075) );
  XNOR2_X1 U11695 ( .A(n15405), .B(n15240), .ZN(n15222) );
  OR2_X1 U11696 ( .A1(n15405), .A2(n15410), .ZN(n9077) );
  INV_X1 U11697 ( .A(n9084), .ZN(n9078) );
  INV_X1 U11698 ( .A(SI_21_), .ZN(n11882) );
  NAND2_X1 U11699 ( .A1(n9078), .A2(n11882), .ZN(n9085) );
  OAI21_X1 U11700 ( .B1(n9082), .B2(SI_20_), .A(n9085), .ZN(n9079) );
  INV_X1 U11701 ( .A(n9079), .ZN(n9080) );
  INV_X1 U11702 ( .A(n9082), .ZN(n9083) );
  NOR2_X1 U11703 ( .A1(n9083), .A2(n11752), .ZN(n9086) );
  AOI22_X1 U11704 ( .A1(n9086), .A2(n9085), .B1(n9084), .B2(SI_21_), .ZN(n9087) );
  OR2_X1 U11705 ( .A1(n9874), .A2(n6533), .ZN(n9088) );
  INV_X1 U11706 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n9428) );
  NAND2_X1 U11707 ( .A1(n9090), .A2(n9428), .ZN(n9091) );
  AND2_X1 U11708 ( .A1(n9105), .A2(n9091), .ZN(n15209) );
  NAND2_X1 U11709 ( .A1(n15209), .A2(n8980), .ZN(n9097) );
  INV_X1 U11710 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n9094) );
  NAND2_X1 U11711 ( .A1(n10490), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n9093) );
  NAND2_X1 U11712 ( .A1(n10533), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n9092) );
  OAI211_X1 U11713 ( .C1(n10536), .C2(n9094), .A(n9093), .B(n9092), .ZN(n9095)
         );
  INV_X1 U11714 ( .A(n9095), .ZN(n9096) );
  AND2_X1 U11715 ( .A1(n15395), .A2(n15402), .ZN(n12704) );
  INV_X1 U11716 ( .A(n12704), .ZN(n14805) );
  MUX2_X1 U11717 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(P1_DATAO_REG_22__SCAN_IN), 
        .S(n6532), .Z(n9873) );
  NAND2_X1 U11718 ( .A1(n9099), .A2(SI_22_), .ZN(n9115) );
  NAND2_X1 U11719 ( .A1(n9116), .A2(n9115), .ZN(n9101) );
  MUX2_X1 U11720 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(P1_DATAO_REG_23__SCAN_IN), 
        .S(n6533), .Z(n9117) );
  XNOR2_X1 U11721 ( .A(n9117), .B(SI_23_), .ZN(n9100) );
  NAND2_X1 U11722 ( .A1(n12166), .A2(n8743), .ZN(n9103) );
  OR2_X1 U11723 ( .A1(n8724), .A2(n12164), .ZN(n9102) );
  INV_X1 U11724 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n9104) );
  NAND2_X1 U11725 ( .A1(n9105), .A2(n9104), .ZN(n9106) );
  NAND2_X1 U11726 ( .A1(n9183), .A2(n9106), .ZN(n14498) );
  INV_X1 U11727 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n9109) );
  NAND2_X1 U11728 ( .A1(n10490), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n9108) );
  NAND2_X1 U11729 ( .A1(n10533), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n9107) );
  OAI211_X1 U11730 ( .C1(n10536), .C2(n9109), .A(n9108), .B(n9107), .ZN(n9110)
         );
  INV_X1 U11731 ( .A(n9110), .ZN(n9111) );
  NAND2_X2 U11732 ( .A1(n9112), .A2(n9111), .ZN(n15212) );
  NAND2_X1 U11733 ( .A1(n15194), .A2(n15212), .ZN(n12726) );
  AND2_X2 U11734 ( .A1(n12729), .A2(n12726), .ZN(n15200) );
  NAND2_X1 U11735 ( .A1(n15192), .A2(n15191), .ZN(n9113) );
  NAND2_X1 U11736 ( .A1(n15194), .A2(n15392), .ZN(n12705) );
  NAND2_X1 U11737 ( .A1(n9117), .A2(SI_23_), .ZN(n9114) );
  INV_X1 U11738 ( .A(n9117), .ZN(n9118) );
  INV_X1 U11739 ( .A(SI_23_), .ZN(n12084) );
  NAND2_X1 U11740 ( .A1(n9118), .A2(n12084), .ZN(n9119) );
  NAND2_X1 U11741 ( .A1(n14471), .A2(n8743), .ZN(n9122) );
  OR2_X1 U11742 ( .A1(n8724), .A2(n15547), .ZN(n9121) );
  XNOR2_X1 U11743 ( .A(n9183), .B(P1_REG3_REG_24__SCAN_IN), .ZN(n15185) );
  NAND2_X1 U11744 ( .A1(n15185), .A2(n8980), .ZN(n9127) );
  INV_X1 U11745 ( .A(P1_REG0_REG_24__SCAN_IN), .ZN(n9457) );
  NAND2_X1 U11746 ( .A1(n10533), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n9124) );
  NAND2_X1 U11747 ( .A1(n14835), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n9123) );
  OAI211_X1 U11748 ( .C1(n14839), .C2(n9457), .A(n9124), .B(n9123), .ZN(n9125)
         );
  INV_X1 U11749 ( .A(n9125), .ZN(n9126) );
  XNOR2_X1 U11750 ( .A(n15187), .B(n14812), .ZN(n9174) );
  INV_X1 U11751 ( .A(n9174), .ZN(n14949) );
  NAND2_X1 U11752 ( .A1(n9139), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9129) );
  MUX2_X1 U11753 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9129), .S(
        P1_IR_REG_20__SCAN_IN), .Z(n9131) );
  INV_X1 U11754 ( .A(n9130), .ZN(n9204) );
  NAND2_X1 U11755 ( .A1(n9193), .A2(n14690), .ZN(n14689) );
  INV_X1 U11756 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n9132) );
  INV_X1 U11757 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n9202) );
  NAND2_X1 U11758 ( .A1(n9132), .A2(n9202), .ZN(n9135) );
  INV_X1 U11759 ( .A(n9135), .ZN(n9133) );
  NAND2_X1 U11760 ( .A1(n9133), .A2(n9201), .ZN(n9138) );
  NAND3_X1 U11761 ( .A1(n9139), .A2(P1_IR_REG_31__SCAN_IN), .A3(
        P1_IR_REG_22__SCAN_IN), .ZN(n9137) );
  XNOR2_X1 U11762 ( .A(P1_IR_REG_31__SCAN_IN), .B(P1_IR_REG_22__SCAN_IN), .ZN(
        n9134) );
  OAI21_X1 U11763 ( .B1(n9135), .B2(n9201), .A(n9134), .ZN(n9136) );
  OAI211_X2 U11764 ( .C1(n9139), .C2(n9138), .A(n9137), .B(n9136), .ZN(n14688)
         );
  OR2_X1 U11765 ( .A1(n14688), .A2(n15178), .ZN(n9140) );
  NAND2_X1 U11766 ( .A1(n10283), .A2(n11497), .ZN(n11385) );
  NAND2_X1 U11768 ( .A1(n10294), .A2(n15783), .ZN(n11638) );
  NAND2_X1 U11769 ( .A1(n11384), .A2(n11638), .ZN(n9143) );
  INV_X1 U11770 ( .A(n14923), .ZN(n9142) );
  NAND2_X1 U11771 ( .A1(n9143), .A2(n9142), .ZN(n11518) );
  NAND2_X1 U11772 ( .A1(n11518), .A2(n9144), .ZN(n9146) );
  INV_X1 U11773 ( .A(n14924), .ZN(n9145) );
  NAND2_X1 U11774 ( .A1(n9146), .A2(n9145), .ZN(n11515) );
  INV_X1 U11775 ( .A(n6534), .ZN(n14701) );
  NAND2_X1 U11776 ( .A1(n14695), .A2(n14701), .ZN(n9147) );
  NAND2_X1 U11777 ( .A1(n11515), .A2(n9147), .ZN(n11279) );
  NAND2_X1 U11778 ( .A1(n14969), .A2(n14725), .ZN(n11735) );
  INV_X1 U11779 ( .A(n14970), .ZN(n11625) );
  NOR2_X1 U11780 ( .A1(n14970), .A2(n7945), .ZN(n11734) );
  AOI21_X1 U11781 ( .B1(n11734), .B2(n11735), .A(n11851), .ZN(n9150) );
  NAND2_X1 U11782 ( .A1(n9151), .A2(n9150), .ZN(n9152) );
  NAND2_X1 U11783 ( .A1(n7943), .A2(n14481), .ZN(n12149) );
  NAND2_X1 U11784 ( .A1(n11853), .A2(n12149), .ZN(n9153) );
  XNOR2_X1 U11785 ( .A(n14733), .B(n14550), .ZN(n12152) );
  NAND2_X1 U11786 ( .A1(n9153), .A2(n12152), .ZN(n12147) );
  OR2_X1 U11787 ( .A1(n14733), .A2(n15799), .ZN(n9154) );
  NAND2_X1 U11788 ( .A1(n11905), .A2(n14920), .ZN(n11904) );
  OR2_X1 U11789 ( .A1(n14737), .A2(n14967), .ZN(n9155) );
  NAND2_X1 U11790 ( .A1(n11904), .A2(n9155), .ZN(n12248) );
  OR2_X1 U11791 ( .A1(n14742), .A2(n15800), .ZN(n9156) );
  NAND2_X1 U11792 ( .A1(n12105), .A2(n14932), .ZN(n12104) );
  INV_X1 U11793 ( .A(n12249), .ZN(n14966) );
  OR2_X1 U11794 ( .A1(n15495), .A2(n14966), .ZN(n9157) );
  NAND2_X1 U11795 ( .A1(n12104), .A2(n9157), .ZN(n12201) );
  OR2_X1 U11796 ( .A1(n15490), .A2(n15478), .ZN(n9158) );
  NAND2_X1 U11797 ( .A1(n12267), .A2(n12266), .ZN(n12265) );
  INV_X1 U11798 ( .A(n15466), .ZN(n14965) );
  OR2_X1 U11799 ( .A1(n15480), .A2(n14965), .ZN(n9159) );
  NAND2_X1 U11800 ( .A1(n12265), .A2(n9159), .ZN(n12316) );
  INV_X1 U11801 ( .A(n14939), .ZN(n12315) );
  INV_X1 U11802 ( .A(n14572), .ZN(n15479) );
  OR2_X1 U11803 ( .A1(n15471), .A2(n15479), .ZN(n9160) );
  NAND2_X1 U11804 ( .A1(n14772), .A2(n15449), .ZN(n9162) );
  NAND2_X1 U11805 ( .A1(n12328), .A2(n9162), .ZN(n15322) );
  INV_X1 U11806 ( .A(n15322), .ZN(n9164) );
  INV_X1 U11807 ( .A(n15324), .ZN(n9163) );
  OR2_X1 U11808 ( .A1(n15325), .A2(n15458), .ZN(n9165) );
  INV_X1 U11809 ( .A(n15434), .ZN(n15450) );
  OR2_X1 U11810 ( .A1(n15444), .A2(n15450), .ZN(n9167) );
  OR2_X1 U11811 ( .A1(n15284), .A2(n15418), .ZN(n9168) );
  NAND2_X1 U11812 ( .A1(n15413), .A2(n15419), .ZN(n9170) );
  NAND2_X1 U11813 ( .A1(n15214), .A2(n15402), .ZN(n9172) );
  NAND2_X1 U11814 ( .A1(n15199), .A2(n12726), .ZN(n9175) );
  NAND2_X1 U11815 ( .A1(n9175), .A2(n9174), .ZN(n9177) );
  AND2_X1 U11816 ( .A1(n14949), .A2(n12726), .ZN(n9176) );
  NAND2_X1 U11817 ( .A1(n9177), .A2(n15167), .ZN(n9180) );
  INV_X1 U11818 ( .A(n14688), .ZN(n15552) );
  NAND2_X1 U11819 ( .A1(n14851), .A2(n15552), .ZN(n9179) );
  OR2_X1 U11820 ( .A1(n14688), .A2(n15103), .ZN(n9178) );
  AND2_X2 U11821 ( .A1(n9179), .A2(n14529), .ZN(n15812) );
  NAND2_X1 U11822 ( .A1(n9180), .A2(n15812), .ZN(n9192) );
  INV_X1 U11823 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n14607) );
  INV_X1 U11824 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n9181) );
  OAI21_X1 U11825 ( .B1(n9183), .B2(n14607), .A(n9181), .ZN(n9184) );
  NAND2_X1 U11826 ( .A1(P1_REG3_REG_24__SCAN_IN), .A2(P1_REG3_REG_25__SCAN_IN), 
        .ZN(n9182) );
  NAND2_X1 U11827 ( .A1(n15174), .A2(n8980), .ZN(n9189) );
  INV_X1 U11828 ( .A(P1_REG0_REG_25__SCAN_IN), .ZN(n9298) );
  NAND2_X1 U11829 ( .A1(n10533), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n9186) );
  NAND2_X1 U11830 ( .A1(n14835), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n9185) );
  OAI211_X1 U11831 ( .C1(n14839), .C2(n9298), .A(n9186), .B(n9185), .ZN(n9187)
         );
  INV_X1 U11832 ( .A(n9187), .ZN(n9188) );
  INV_X1 U11833 ( .A(n15533), .ZN(n10742) );
  OAI22_X1 U11834 ( .A1(n14816), .A2(n15467), .B1(n15392), .B2(n12723), .ZN(
        n14610) );
  INV_X1 U11835 ( .A(n14610), .ZN(n9191) );
  NAND2_X1 U11836 ( .A1(n14953), .A2(n14688), .ZN(n11386) );
  NAND2_X1 U11837 ( .A1(n15783), .A2(n11371), .ZN(n11645) );
  INV_X1 U11838 ( .A(n14733), .ZN(n15795) );
  INV_X1 U11839 ( .A(n14737), .ZN(n15805) );
  INV_X1 U11840 ( .A(n15490), .ZN(n14753) );
  INV_X1 U11841 ( .A(n15480), .ZN(n12271) );
  NAND2_X1 U11842 ( .A1(n12272), .A2(n12271), .ZN(n12320) );
  INV_X1 U11843 ( .A(n15444), .ZN(n15317) );
  NAND2_X1 U11844 ( .A1(n15328), .A2(n15317), .ZN(n15313) );
  AND2_X2 U11845 ( .A1(n15208), .A2(n15386), .ZN(n9197) );
  OAI211_X1 U11846 ( .C1(n9197), .C2(n15187), .A(n15447), .B(n15173), .ZN(
        n15184) );
  OAI21_X1 U11847 ( .B1(n15187), .B2(n15804), .A(n15184), .ZN(n9198) );
  INV_X1 U11848 ( .A(n9198), .ZN(n9199) );
  NAND2_X1 U11849 ( .A1(n15807), .A2(n10631), .ZN(n9219) );
  NAND2_X1 U11850 ( .A1(n9202), .A2(n9201), .ZN(n9203) );
  INV_X1 U11851 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n9205) );
  NAND2_X1 U11852 ( .A1(n9209), .A2(n9208), .ZN(n9214) );
  NAND2_X1 U11853 ( .A1(n9211), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9213) );
  NAND2_X1 U11854 ( .A1(n9214), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9215) );
  MUX2_X1 U11855 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9215), .S(
        P1_IR_REG_25__SCAN_IN), .Z(n9216) );
  AND2_X1 U11856 ( .A1(n9211), .A2(n9216), .ZN(n9220) );
  AND2_X1 U11857 ( .A1(n10630), .A2(n10549), .ZN(n9218) );
  NAND2_X1 U11858 ( .A1(n9219), .A2(n9218), .ZN(n10522) );
  INV_X1 U11859 ( .A(n9220), .ZN(n15543) );
  NAND3_X1 U11860 ( .A1(n15543), .A2(P1_B_REG_SCAN_IN), .A3(n15550), .ZN(n9224) );
  INV_X1 U11861 ( .A(n15550), .ZN(n9222) );
  INV_X1 U11862 ( .A(P1_B_REG_SCAN_IN), .ZN(n9221) );
  AOI21_X1 U11863 ( .B1(n9222), .B2(n9221), .A(n15542), .ZN(n9223) );
  INV_X1 U11864 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n9225) );
  NAND2_X1 U11865 ( .A1(n9239), .A2(n9225), .ZN(n9226) );
  NAND2_X1 U11866 ( .A1(n15543), .A2(n15542), .ZN(n10641) );
  NAND2_X1 U11867 ( .A1(n9226), .A2(n10641), .ZN(n10517) );
  NOR4_X1 U11868 ( .A1(P1_D_REG_7__SCAN_IN), .A2(P1_D_REG_8__SCAN_IN), .A3(
        P1_D_REG_9__SCAN_IN), .A4(P1_D_REG_10__SCAN_IN), .ZN(n9235) );
  NOR4_X1 U11869 ( .A1(P1_D_REG_18__SCAN_IN), .A2(P1_D_REG_3__SCAN_IN), .A3(
        P1_D_REG_4__SCAN_IN), .A4(P1_D_REG_5__SCAN_IN), .ZN(n9234) );
  INV_X1 U11870 ( .A(P1_D_REG_6__SCAN_IN), .ZN(n15776) );
  INV_X1 U11871 ( .A(P1_D_REG_2__SCAN_IN), .ZN(n15780) );
  INV_X1 U11872 ( .A(P1_D_REG_28__SCAN_IN), .ZN(n15754) );
  INV_X1 U11873 ( .A(P1_D_REG_13__SCAN_IN), .ZN(n15769) );
  NAND4_X1 U11874 ( .A1(n15776), .A2(n15780), .A3(n15754), .A4(n15769), .ZN(
        n9232) );
  NOR4_X1 U11875 ( .A1(P1_D_REG_16__SCAN_IN), .A2(P1_D_REG_17__SCAN_IN), .A3(
        P1_D_REG_19__SCAN_IN), .A4(P1_D_REG_20__SCAN_IN), .ZN(n9230) );
  NOR4_X1 U11876 ( .A1(P1_D_REG_14__SCAN_IN), .A2(P1_D_REG_11__SCAN_IN), .A3(
        P1_D_REG_12__SCAN_IN), .A4(P1_D_REG_15__SCAN_IN), .ZN(n9229) );
  NOR4_X1 U11877 ( .A1(P1_D_REG_25__SCAN_IN), .A2(P1_D_REG_26__SCAN_IN), .A3(
        P1_D_REG_27__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n9228) );
  NOR4_X1 U11878 ( .A1(P1_D_REG_21__SCAN_IN), .A2(P1_D_REG_22__SCAN_IN), .A3(
        P1_D_REG_23__SCAN_IN), .A4(P1_D_REG_24__SCAN_IN), .ZN(n9227) );
  NAND4_X1 U11879 ( .A1(n9230), .A2(n9229), .A3(n9228), .A4(n9227), .ZN(n9231)
         );
  NOR4_X1 U11880 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        n9232), .A4(n9231), .ZN(n9233) );
  AND3_X1 U11881 ( .A1(n9235), .A2(n9234), .A3(n9233), .ZN(n9236) );
  OR2_X1 U11882 ( .A1(n10639), .A2(n9236), .ZN(n10518) );
  NAND3_X1 U11883 ( .A1(n10517), .A2(n11381), .A3(n10518), .ZN(n9237) );
  INV_X1 U11884 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n9238) );
  NAND2_X1 U11885 ( .A1(n15820), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n9240) );
  INV_X1 U11886 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n15843) );
  AOI22_X1 U11887 ( .A1(n15843), .A2(keyinput100), .B1(keyinput77), .B2(n12205), .ZN(n9241) );
  OAI221_X1 U11888 ( .B1(n15843), .B2(keyinput100), .C1(n12205), .C2(
        keyinput77), .A(n9241), .ZN(n9293) );
  INV_X1 U11889 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n15624) );
  AOI22_X1 U11890 ( .A1(n15624), .A2(keyinput121), .B1(n9457), .B2(keyinput86), 
        .ZN(n9242) );
  OAI221_X1 U11891 ( .B1(n15624), .B2(keyinput121), .C1(n9457), .C2(keyinput86), .A(n9242), .ZN(n9247) );
  XNOR2_X1 U11892 ( .A(SI_6_), .B(keyinput62), .ZN(n9245) );
  NAND2_X1 U11893 ( .A1(n10097), .A2(keyinput64), .ZN(n9244) );
  XNOR2_X1 U11894 ( .A(keyinput23), .B(P2_D_REG_20__SCAN_IN), .ZN(n9243) );
  NAND3_X1 U11895 ( .A1(n9245), .A2(n9244), .A3(n9243), .ZN(n9246) );
  NOR2_X1 U11896 ( .A1(n9247), .A2(n9246), .ZN(n9281) );
  XNOR2_X1 U11897 ( .A(P3_B_REG_SCAN_IN), .B(keyinput81), .ZN(n9251) );
  XNOR2_X1 U11898 ( .A(P3_REG3_REG_6__SCAN_IN), .B(keyinput105), .ZN(n9250) );
  XNOR2_X1 U11899 ( .A(P1_IR_REG_26__SCAN_IN), .B(keyinput44), .ZN(n9249) );
  XNOR2_X1 U11900 ( .A(P1_IR_REG_7__SCAN_IN), .B(keyinput67), .ZN(n9248) );
  NAND4_X1 U11901 ( .A1(n9251), .A2(n9250), .A3(n9249), .A4(n9248), .ZN(n9257)
         );
  XNOR2_X1 U11902 ( .A(P1_IR_REG_30__SCAN_IN), .B(keyinput113), .ZN(n9255) );
  XNOR2_X1 U11903 ( .A(P1_REG1_REG_12__SCAN_IN), .B(keyinput111), .ZN(n9254)
         );
  XNOR2_X1 U11904 ( .A(P1_REG1_REG_0__SCAN_IN), .B(keyinput97), .ZN(n9253) );
  XNOR2_X1 U11905 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(keyinput99), .ZN(n9252)
         );
  NAND4_X1 U11906 ( .A1(n9255), .A2(n9254), .A3(n9253), .A4(n9252), .ZN(n9256)
         );
  NOR2_X1 U11907 ( .A1(n9257), .A2(n9256), .ZN(n9280) );
  XNOR2_X1 U11908 ( .A(P1_REG2_REG_20__SCAN_IN), .B(keyinput11), .ZN(n9261) );
  XNOR2_X1 U11909 ( .A(P1_REG3_REG_21__SCAN_IN), .B(keyinput16), .ZN(n9260) );
  XNOR2_X1 U11910 ( .A(P1_REG3_REG_26__SCAN_IN), .B(keyinput30), .ZN(n9259) );
  XNOR2_X1 U11911 ( .A(P2_IR_REG_17__SCAN_IN), .B(keyinput73), .ZN(n9258) );
  NAND4_X1 U11912 ( .A1(n9261), .A2(n9260), .A3(n9259), .A4(n9258), .ZN(n9267)
         );
  XNOR2_X1 U11913 ( .A(P2_IR_REG_15__SCAN_IN), .B(keyinput20), .ZN(n9265) );
  XNOR2_X1 U11914 ( .A(P2_D_REG_0__SCAN_IN), .B(keyinput88), .ZN(n9264) );
  XNOR2_X1 U11915 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(keyinput72), .ZN(n9263)
         );
  XNOR2_X1 U11916 ( .A(P2_REG1_REG_11__SCAN_IN), .B(keyinput58), .ZN(n9262) );
  NAND4_X1 U11917 ( .A1(n9265), .A2(n9264), .A3(n9263), .A4(n9262), .ZN(n9266)
         );
  NOR2_X1 U11918 ( .A1(n9267), .A2(n9266), .ZN(n9279) );
  XNOR2_X1 U11919 ( .A(P2_REG3_REG_10__SCAN_IN), .B(keyinput34), .ZN(n9271) );
  XNOR2_X1 U11920 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(keyinput74), .ZN(n9270)
         );
  XNOR2_X1 U11921 ( .A(P3_REG1_REG_30__SCAN_IN), .B(keyinput5), .ZN(n9269) );
  XNOR2_X1 U11922 ( .A(P3_IR_REG_6__SCAN_IN), .B(keyinput54), .ZN(n9268) );
  NAND4_X1 U11923 ( .A1(n9271), .A2(n9270), .A3(n9269), .A4(n9268), .ZN(n9277)
         );
  XNOR2_X1 U11924 ( .A(SI_2_), .B(keyinput109), .ZN(n9275) );
  XNOR2_X1 U11925 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(keyinput126), .ZN(n9274)
         );
  XNOR2_X1 U11926 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(keyinput107), .ZN(n9273)
         );
  XNOR2_X1 U11927 ( .A(P1_REG3_REG_7__SCAN_IN), .B(keyinput93), .ZN(n9272) );
  NAND4_X1 U11928 ( .A1(n9275), .A2(n9274), .A3(n9273), .A4(n9272), .ZN(n9276)
         );
  NOR2_X1 U11929 ( .A1(n9277), .A2(n9276), .ZN(n9278) );
  NAND4_X1 U11930 ( .A1(n9281), .A2(n9280), .A3(n9279), .A4(n9278), .ZN(n9292)
         );
  INV_X1 U11931 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n15697) );
  INV_X1 U11932 ( .A(P3_ADDR_REG_12__SCAN_IN), .ZN(n15576) );
  AOI22_X1 U11933 ( .A1(n15697), .A2(keyinput108), .B1(keyinput0), .B2(n15576), 
        .ZN(n9282) );
  OAI221_X1 U11934 ( .B1(n15697), .B2(keyinput108), .C1(n15576), .C2(keyinput0), .A(n9282), .ZN(n9291) );
  INV_X1 U11935 ( .A(P1_REG2_REG_26__SCAN_IN), .ZN(n9284) );
  AOI22_X1 U11936 ( .A1(n9284), .A2(keyinput10), .B1(keyinput101), .B2(n11525), 
        .ZN(n9283) );
  OAI221_X1 U11937 ( .B1(n9284), .B2(keyinput10), .C1(n11525), .C2(keyinput101), .A(n9283), .ZN(n9289) );
  INV_X1 U11938 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n15637) );
  INV_X1 U11939 ( .A(P3_REG0_REG_26__SCAN_IN), .ZN(n13435) );
  AOI22_X1 U11940 ( .A1(n15637), .A2(keyinput25), .B1(n13435), .B2(keyinput26), 
        .ZN(n9285) );
  OAI221_X1 U11941 ( .B1(n15637), .B2(keyinput25), .C1(n13435), .C2(keyinput26), .A(n9285), .ZN(n9288) );
  AOI22_X1 U11942 ( .A1(n13249), .A2(keyinput61), .B1(keyinput103), .B2(n15041), .ZN(n9286) );
  OAI221_X1 U11943 ( .B1(n13249), .B2(keyinput61), .C1(n15041), .C2(
        keyinput103), .A(n9286), .ZN(n9287) );
  OR3_X1 U11944 ( .A1(n9289), .A2(n9288), .A3(n9287), .ZN(n9290) );
  NOR4_X1 U11945 ( .A1(n9293), .A2(n9292), .A3(n9291), .A4(n9290), .ZN(n9321)
         );
  INV_X1 U11946 ( .A(P3_REG1_REG_5__SCAN_IN), .ZN(n15968) );
  INV_X1 U11947 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n9423) );
  AOI22_X1 U11948 ( .A1(n15968), .A2(keyinput79), .B1(keyinput127), .B2(n9423), 
        .ZN(n9294) );
  OAI221_X1 U11949 ( .B1(n15968), .B2(keyinput79), .C1(n9423), .C2(keyinput127), .A(n9294), .ZN(n9302) );
  INV_X1 U11950 ( .A(P3_REG0_REG_9__SCAN_IN), .ZN(n9296) );
  AOI22_X1 U11951 ( .A1(n9296), .A2(keyinput112), .B1(keyinput117), .B2(n9415), 
        .ZN(n9295) );
  OAI221_X1 U11952 ( .B1(n9296), .B2(keyinput112), .C1(n9415), .C2(keyinput117), .A(n9295), .ZN(n9301) );
  INV_X1 U11953 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n9299) );
  AOI22_X1 U11954 ( .A1(n9299), .A2(keyinput71), .B1(keyinput19), .B2(n9298), 
        .ZN(n9297) );
  OAI221_X1 U11955 ( .B1(n9299), .B2(keyinput71), .C1(n9298), .C2(keyinput19), 
        .A(n9297), .ZN(n9300) );
  NOR3_X1 U11956 ( .A1(n9302), .A2(n9301), .A3(n9300), .ZN(n9320) );
  INV_X1 U11957 ( .A(P2_D_REG_8__SCAN_IN), .ZN(n15876) );
  AOI22_X1 U11958 ( .A1(n15538), .A2(keyinput29), .B1(keyinput94), .B2(n15876), 
        .ZN(n9303) );
  OAI221_X1 U11959 ( .B1(n15538), .B2(keyinput29), .C1(n15876), .C2(keyinput94), .A(n9303), .ZN(n9306) );
  INV_X1 U11960 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n13659) );
  INV_X1 U11961 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n15632) );
  AOI22_X1 U11962 ( .A1(n13659), .A2(keyinput32), .B1(keyinput83), .B2(n15632), 
        .ZN(n9304) );
  OAI221_X1 U11963 ( .B1(n13659), .B2(keyinput32), .C1(n15632), .C2(keyinput83), .A(n9304), .ZN(n9305) );
  NOR2_X1 U11964 ( .A1(n9306), .A2(n9305), .ZN(n9319) );
  AOI22_X1 U11965 ( .A1(n12806), .A2(keyinput75), .B1(keyinput92), .B2(n11692), 
        .ZN(n9307) );
  OAI221_X1 U11966 ( .B1(n12806), .B2(keyinput75), .C1(n11692), .C2(keyinput92), .A(n9307), .ZN(n9312) );
  INV_X1 U11967 ( .A(P2_B_REG_SCAN_IN), .ZN(n10264) );
  AOI22_X1 U11968 ( .A1(n8435), .A2(keyinput123), .B1(keyinput57), .B2(n10264), 
        .ZN(n9308) );
  OAI221_X1 U11969 ( .B1(n8435), .B2(keyinput123), .C1(n10264), .C2(keyinput57), .A(n9308), .ZN(n9311) );
  AOI22_X1 U11970 ( .A1(n7111), .A2(keyinput52), .B1(keyinput66), .B2(n11757), 
        .ZN(n9309) );
  OAI221_X1 U11971 ( .B1(n7111), .B2(keyinput52), .C1(n11757), .C2(keyinput66), 
        .A(n9309), .ZN(n9310) );
  OR3_X1 U11972 ( .A1(n9312), .A2(n9311), .A3(n9310), .ZN(n9317) );
  INV_X1 U11973 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n13722) );
  AOI22_X1 U11974 ( .A1(n13722), .A2(keyinput102), .B1(keyinput28), .B2(n15562), .ZN(n9313) );
  OAI221_X1 U11975 ( .B1(n13722), .B2(keyinput102), .C1(n15562), .C2(
        keyinput28), .A(n9313), .ZN(n9316) );
  INV_X1 U11976 ( .A(P3_REG3_REG_0__SCAN_IN), .ZN(n10817) );
  AOI22_X1 U11977 ( .A1(n10817), .A2(keyinput89), .B1(keyinput49), .B2(n15754), 
        .ZN(n9314) );
  OAI221_X1 U11978 ( .B1(n10817), .B2(keyinput89), .C1(n15754), .C2(keyinput49), .A(n9314), .ZN(n9315) );
  NOR3_X1 U11979 ( .A1(n9317), .A2(n9316), .A3(n9315), .ZN(n9318) );
  NAND4_X1 U11980 ( .A1(n9321), .A2(n9320), .A3(n9319), .A4(n9318), .ZN(n9382)
         );
  INV_X1 U11981 ( .A(P3_REG1_REG_14__SCAN_IN), .ZN(n13402) );
  AOI22_X1 U11982 ( .A1(n12158), .A2(keyinput22), .B1(n13402), .B2(keyinput56), 
        .ZN(n9322) );
  OAI221_X1 U11983 ( .B1(n12158), .B2(keyinput22), .C1(n13402), .C2(keyinput56), .A(n9322), .ZN(n9330) );
  INV_X1 U11984 ( .A(P3_ADDR_REG_17__SCAN_IN), .ZN(n9324) );
  AOI22_X1 U11985 ( .A1(n9324), .A2(keyinput51), .B1(n8694), .B2(keyinput6), 
        .ZN(n9323) );
  OAI221_X1 U11986 ( .B1(n9324), .B2(keyinput51), .C1(n8694), .C2(keyinput6), 
        .A(n9323), .ZN(n9329) );
  INV_X1 U11987 ( .A(P3_REG2_REG_30__SCAN_IN), .ZN(n9421) );
  AOI22_X1 U11988 ( .A1(n10747), .A2(keyinput114), .B1(n9421), .B2(keyinput70), 
        .ZN(n9325) );
  OAI221_X1 U11989 ( .B1(n10747), .B2(keyinput114), .C1(n9421), .C2(keyinput70), .A(n9325), .ZN(n9328) );
  INV_X1 U11990 ( .A(P3_REG1_REG_18__SCAN_IN), .ZN(n13388) );
  AOI22_X1 U11991 ( .A1(n15556), .A2(keyinput95), .B1(n13388), .B2(keyinput35), 
        .ZN(n9326) );
  OAI221_X1 U11992 ( .B1(n15556), .B2(keyinput95), .C1(n13388), .C2(keyinput35), .A(n9326), .ZN(n9327) );
  NOR4_X1 U11993 ( .A1(n9330), .A2(n9329), .A3(n9328), .A4(n9327), .ZN(n9344)
         );
  INV_X1 U11994 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n12419) );
  INV_X1 U11995 ( .A(P3_D_REG_18__SCAN_IN), .ZN(n9332) );
  AOI22_X1 U11996 ( .A1(n12419), .A2(keyinput18), .B1(keyinput60), .B2(n9332), 
        .ZN(n9331) );
  OAI221_X1 U11997 ( .B1(n12419), .B2(keyinput18), .C1(n9332), .C2(keyinput60), 
        .A(n9331), .ZN(n9335) );
  INV_X1 U11998 ( .A(P3_DATAO_REG_4__SCAN_IN), .ZN(n10649) );
  INV_X1 U11999 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n9446) );
  AOI22_X1 U12000 ( .A1(n10649), .A2(keyinput45), .B1(n9446), .B2(keyinput69), 
        .ZN(n9333) );
  OAI221_X1 U12001 ( .B1(n10649), .B2(keyinput45), .C1(n9446), .C2(keyinput69), 
        .A(n9333), .ZN(n9334) );
  NOR2_X1 U12002 ( .A1(n9335), .A2(n9334), .ZN(n9343) );
  INV_X1 U12003 ( .A(P3_DATAO_REG_25__SCAN_IN), .ZN(n12018) );
  AOI22_X1 U12004 ( .A1(n7046), .A2(keyinput76), .B1(keyinput14), .B2(n12018), 
        .ZN(n9336) );
  OAI221_X1 U12005 ( .B1(n7046), .B2(keyinput76), .C1(n12018), .C2(keyinput14), 
        .A(n9336), .ZN(n9341) );
  INV_X1 U12006 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n12395) );
  INV_X1 U12007 ( .A(SI_30_), .ZN(n12649) );
  AOI22_X1 U12008 ( .A1(n12395), .A2(keyinput36), .B1(n12649), .B2(keyinput39), 
        .ZN(n9337) );
  OAI221_X1 U12009 ( .B1(n12395), .B2(keyinput36), .C1(n12649), .C2(keyinput39), .A(n9337), .ZN(n9340) );
  INV_X1 U12010 ( .A(P2_REG2_REG_30__SCAN_IN), .ZN(n9439) );
  AOI22_X1 U12011 ( .A1(n9439), .A2(keyinput41), .B1(n9432), .B2(keyinput31), 
        .ZN(n9338) );
  OAI221_X1 U12012 ( .B1(n9439), .B2(keyinput41), .C1(n9432), .C2(keyinput31), 
        .A(n9338), .ZN(n9339) );
  NOR3_X1 U12013 ( .A1(n9341), .A2(n9340), .A3(n9339), .ZN(n9342) );
  NAND3_X1 U12014 ( .A1(n9344), .A2(n9343), .A3(n9342), .ZN(n9381) );
  INV_X1 U12015 ( .A(P3_REG1_REG_4__SCAN_IN), .ZN(n15966) );
  INV_X1 U12016 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n9977) );
  AOI22_X1 U12017 ( .A1(n15966), .A2(keyinput47), .B1(keyinput21), .B2(n9977), 
        .ZN(n9345) );
  OAI221_X1 U12018 ( .B1(n15966), .B2(keyinput47), .C1(n9977), .C2(keyinput21), 
        .A(n9345), .ZN(n9356) );
  INV_X1 U12019 ( .A(P2_D_REG_22__SCAN_IN), .ZN(n15873) );
  AOI22_X1 U12020 ( .A1(n15873), .A2(keyinput104), .B1(n11292), .B2(keyinput53), .ZN(n9346) );
  OAI221_X1 U12021 ( .B1(n15873), .B2(keyinput104), .C1(n11292), .C2(
        keyinput53), .A(n9346), .ZN(n9355) );
  AOI22_X1 U12022 ( .A1(n8729), .A2(keyinput7), .B1(n9348), .B2(keyinput40), 
        .ZN(n9347) );
  OAI221_X1 U12023 ( .B1(n8729), .B2(keyinput7), .C1(n9348), .C2(keyinput40), 
        .A(n9347), .ZN(n9354) );
  XOR2_X1 U12024 ( .A(n8663), .B(keyinput119), .Z(n9352) );
  INV_X1 U12025 ( .A(P2_D_REG_2__SCAN_IN), .ZN(n15878) );
  XOR2_X1 U12026 ( .A(n15878), .B(keyinput13), .Z(n9351) );
  XNOR2_X1 U12027 ( .A(P3_REG3_REG_4__SCAN_IN), .B(keyinput3), .ZN(n9350) );
  XNOR2_X1 U12028 ( .A(P1_IR_REG_4__SCAN_IN), .B(keyinput15), .ZN(n9349) );
  NAND4_X1 U12029 ( .A1(n9352), .A2(n9351), .A3(n9350), .A4(n9349), .ZN(n9353)
         );
  NOR4_X1 U12030 ( .A1(n9356), .A2(n9355), .A3(n9354), .A4(n9353), .ZN(n9369)
         );
  XOR2_X1 U12031 ( .A(keyinput8), .B(n15776), .Z(n9368) );
  XOR2_X1 U12032 ( .A(P2_REG1_REG_2__SCAN_IN), .B(keyinput106), .Z(n9360) );
  XOR2_X1 U12033 ( .A(P3_REG3_REG_3__SCAN_IN), .B(keyinput91), .Z(n9359) );
  INV_X2 U12034 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n9471) );
  XNOR2_X1 U12035 ( .A(n9471), .B(keyinput63), .ZN(n9358) );
  XNOR2_X1 U12036 ( .A(n10836), .B(keyinput48), .ZN(n9357) );
  NOR4_X1 U12037 ( .A1(n9360), .A2(n9359), .A3(n9358), .A4(n9357), .ZN(n9367)
         );
  XOR2_X1 U12038 ( .A(P3_REG1_REG_27__SCAN_IN), .B(keyinput50), .Z(n9365) );
  XOR2_X1 U12039 ( .A(P1_REG3_REG_2__SCAN_IN), .B(keyinput17), .Z(n9364) );
  XNOR2_X1 U12040 ( .A(n9361), .B(keyinput24), .ZN(n9363) );
  XNOR2_X1 U12041 ( .A(n11248), .B(keyinput37), .ZN(n9362) );
  NOR4_X1 U12042 ( .A1(n9365), .A2(n9364), .A3(n9363), .A4(n9362), .ZN(n9366)
         );
  NAND4_X1 U12043 ( .A1(n9369), .A2(n9368), .A3(n9367), .A4(n9366), .ZN(n9380)
         );
  INV_X1 U12044 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n15586) );
  INV_X1 U12045 ( .A(P2_REG2_REG_31__SCAN_IN), .ZN(n9371) );
  AOI22_X1 U12046 ( .A1(n15586), .A2(keyinput46), .B1(n9371), .B2(keyinput38), 
        .ZN(n9370) );
  OAI221_X1 U12047 ( .B1(n15586), .B2(keyinput46), .C1(n9371), .C2(keyinput38), 
        .A(n9370), .ZN(n9378) );
  INV_X1 U12048 ( .A(P3_DATAO_REG_28__SCAN_IN), .ZN(n12285) );
  INV_X1 U12049 ( .A(P3_DATAO_REG_0__SCAN_IN), .ZN(n10651) );
  AOI22_X1 U12050 ( .A1(n12285), .A2(keyinput33), .B1(keyinput84), .B2(n10651), 
        .ZN(n9372) );
  OAI221_X1 U12051 ( .B1(n12285), .B2(keyinput33), .C1(n10651), .C2(keyinput84), .A(n9372), .ZN(n9377) );
  INV_X1 U12052 ( .A(P3_ADDR_REG_11__SCAN_IN), .ZN(n15574) );
  AOI22_X1 U12053 ( .A1(n15574), .A2(keyinput27), .B1(n8230), .B2(keyinput2), 
        .ZN(n9373) );
  OAI221_X1 U12054 ( .B1(n15574), .B2(keyinput27), .C1(n8230), .C2(keyinput2), 
        .A(n9373), .ZN(n9376) );
  INV_X1 U12055 ( .A(P3_REG1_REG_16__SCAN_IN), .ZN(n13394) );
  AOI22_X1 U12056 ( .A1(n6789), .A2(keyinput59), .B1(n13394), .B2(keyinput68), 
        .ZN(n9374) );
  OAI221_X1 U12057 ( .B1(n6789), .B2(keyinput59), .C1(n13394), .C2(keyinput68), 
        .A(n9374), .ZN(n9375) );
  OR4_X1 U12058 ( .A1(n9378), .A2(n9377), .A3(n9376), .A4(n9375), .ZN(n9379)
         );
  NOR4_X1 U12059 ( .A1(n9382), .A2(n9381), .A3(n9380), .A4(n9379), .ZN(n9413)
         );
  INV_X1 U12060 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n15907) );
  AOI22_X1 U12061 ( .A1(n15557), .A2(keyinput85), .B1(n15907), .B2(keyinput116), .ZN(n9383) );
  OAI221_X1 U12062 ( .B1(n15557), .B2(keyinput85), .C1(n15907), .C2(
        keyinput116), .A(n9383), .ZN(n9391) );
  INV_X1 U12063 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n15653) );
  AOI22_X1 U12064 ( .A1(n8850), .A2(keyinput43), .B1(keyinput118), .B2(n15653), 
        .ZN(n9384) );
  OAI221_X1 U12065 ( .B1(n8850), .B2(keyinput43), .C1(n15653), .C2(keyinput118), .A(n9384), .ZN(n9390) );
  INV_X1 U12066 ( .A(P1_D_REG_18__SCAN_IN), .ZN(n15764) );
  AOI22_X1 U12067 ( .A1(n15769), .A2(keyinput55), .B1(keyinput125), .B2(n15764), .ZN(n9385) );
  OAI221_X1 U12068 ( .B1(n15769), .B2(keyinput55), .C1(n15764), .C2(
        keyinput125), .A(n9385), .ZN(n9389) );
  INV_X1 U12069 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n9866) );
  INV_X1 U12070 ( .A(P3_REG0_REG_13__SCAN_IN), .ZN(n9387) );
  AOI22_X1 U12071 ( .A1(n9866), .A2(keyinput122), .B1(n9387), .B2(keyinput78), 
        .ZN(n9386) );
  OAI221_X1 U12072 ( .B1(n9866), .B2(keyinput122), .C1(n9387), .C2(keyinput78), 
        .A(n9386), .ZN(n9388) );
  NOR4_X1 U12073 ( .A1(n9391), .A2(n9390), .A3(n9389), .A4(n9388), .ZN(n9412)
         );
  INV_X1 U12074 ( .A(P2_D_REG_12__SCAN_IN), .ZN(n15875) );
  INV_X1 U12075 ( .A(P1_REG2_REG_29__SCAN_IN), .ZN(n15136) );
  AOI22_X1 U12076 ( .A1(n15875), .A2(keyinput9), .B1(keyinput90), .B2(n15136), 
        .ZN(n9392) );
  OAI221_X1 U12077 ( .B1(n15875), .B2(keyinput9), .C1(n15136), .C2(keyinput90), 
        .A(n9392), .ZN(n9400) );
  AOI22_X1 U12078 ( .A1(n9652), .A2(keyinput115), .B1(keyinput80), .B2(n11147), 
        .ZN(n9393) );
  OAI221_X1 U12079 ( .B1(n9652), .B2(keyinput115), .C1(n11147), .C2(keyinput80), .A(n9393), .ZN(n9399) );
  INV_X1 U12080 ( .A(P3_REG2_REG_27__SCAN_IN), .ZN(n9395) );
  INV_X1 U12081 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n10528) );
  AOI22_X1 U12082 ( .A1(n9395), .A2(keyinput124), .B1(keyinput98), .B2(n10528), 
        .ZN(n9394) );
  OAI221_X1 U12083 ( .B1(n9395), .B2(keyinput124), .C1(n10528), .C2(keyinput98), .A(n9394), .ZN(n9398) );
  INV_X1 U12084 ( .A(P3_REG1_REG_6__SCAN_IN), .ZN(n15971) );
  INV_X1 U12085 ( .A(SI_28_), .ZN(n13514) );
  AOI22_X1 U12086 ( .A1(n15971), .A2(keyinput120), .B1(n13514), .B2(keyinput96), .ZN(n9396) );
  OAI221_X1 U12087 ( .B1(n15971), .B2(keyinput120), .C1(n13514), .C2(
        keyinput96), .A(n9396), .ZN(n9397) );
  NOR4_X1 U12088 ( .A1(n9400), .A2(n9399), .A3(n9398), .A4(n9397), .ZN(n9411)
         );
  INV_X1 U12089 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n9402) );
  AOI22_X1 U12090 ( .A1(n9402), .A2(keyinput4), .B1(keyinput1), .B2(n8995), 
        .ZN(n9401) );
  OAI221_X1 U12091 ( .B1(n9402), .B2(keyinput4), .C1(n8995), .C2(keyinput1), 
        .A(n9401), .ZN(n9409) );
  INV_X1 U12092 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n10875) );
  AOI22_X1 U12093 ( .A1(n10875), .A2(keyinput110), .B1(P2_U3088), .B2(
        keyinput12), .ZN(n9403) );
  OAI221_X1 U12094 ( .B1(n10875), .B2(keyinput110), .C1(P2_U3088), .C2(
        keyinput12), .A(n9403), .ZN(n9408) );
  INV_X1 U12095 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n10507) );
  AOI22_X1 U12096 ( .A1(n10507), .A2(keyinput82), .B1(n9428), .B2(keyinput65), 
        .ZN(n9404) );
  OAI221_X1 U12097 ( .B1(n10507), .B2(keyinput82), .C1(n9428), .C2(keyinput65), 
        .A(n9404), .ZN(n9407) );
  INV_X1 U12098 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n9673) );
  AOI22_X1 U12099 ( .A1(n9673), .A2(keyinput87), .B1(keyinput42), .B2(n15780), 
        .ZN(n9405) );
  OAI221_X1 U12100 ( .B1(n9673), .B2(keyinput87), .C1(n15780), .C2(keyinput42), 
        .A(n9405), .ZN(n9406) );
  NOR4_X1 U12101 ( .A1(n9409), .A2(n9408), .A3(n9407), .A4(n9406), .ZN(n9410)
         );
  NAND4_X1 U12102 ( .A1(n9413), .A2(n9412), .A3(n9411), .A4(n9410), .ZN(n9470)
         );
  NOR4_X1 U12103 ( .A1(n9415), .A2(n9414), .A3(SI_28_), .A4(
        P1_IR_REG_18__SCAN_IN), .ZN(n9427) );
  NAND4_X1 U12104 ( .A1(P3_REG0_REG_19__SCAN_IN), .A2(P3_REG2_REG_20__SCAN_IN), 
        .A3(n10264), .A4(n8729), .ZN(n9418) );
  NAND4_X1 U12105 ( .A1(P3_REG3_REG_7__SCAN_IN), .A2(P2_REG2_REG_27__SCAN_IN), 
        .A3(P2_REG1_REG_8__SCAN_IN), .A4(P1_IR_REG_15__SCAN_IN), .ZN(n9417) );
  NAND2_X1 U12106 ( .A1(P2_DATAO_REG_31__SCAN_IN), .A2(n12419), .ZN(n9416) );
  NAND2_X1 U12107 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(P2_U3088), .ZN(n11174)
         );
  NOR4_X1 U12108 ( .A1(n9418), .A2(n9417), .A3(n9416), .A4(n11174), .ZN(n9425)
         );
  NOR4_X1 U12109 ( .A1(P2_REG0_REG_30__SCAN_IN), .A2(P1_IR_REG_30__SCAN_IN), 
        .A3(P1_REG0_REG_25__SCAN_IN), .A4(P1_REG1_REG_0__SCAN_IN), .ZN(n9420)
         );
  NOR4_X1 U12110 ( .A1(P2_DATAO_REG_13__SCAN_IN), .A2(P1_REG2_REG_26__SCAN_IN), 
        .A3(n15776), .A4(n11525), .ZN(n9419) );
  AND4_X1 U12111 ( .A1(P1_REG2_REG_7__SCAN_IN), .A2(n9421), .A3(n9420), .A4(
        n9419), .ZN(n9424) );
  NOR4_X1 U12112 ( .A1(P2_REG3_REG_25__SCAN_IN), .A2(P1_REG0_REG_3__SCAN_IN), 
        .A3(P2_ADDR_REG_17__SCAN_IN), .A4(P3_ADDR_REG_17__SCAN_IN), .ZN(n9422)
         );
  AND4_X1 U12113 ( .A1(n9425), .A2(n9424), .A3(n9423), .A4(n9422), .ZN(n9426)
         );
  NAND4_X1 U12114 ( .A1(n9427), .A2(P1_IR_REG_4__SCAN_IN), .A3(
        P2_D_REG_2__SCAN_IN), .A4(n9426), .ZN(n9430) );
  NAND4_X1 U12115 ( .A1(P1_D_REG_2__SCAN_IN), .A2(P2_REG1_REG_10__SCAN_IN), 
        .A3(P1_REG0_REG_27__SCAN_IN), .A4(n9428), .ZN(n9429) );
  NOR2_X1 U12116 ( .A1(n9430), .A2(n9429), .ZN(n9437) );
  NOR4_X1 U12117 ( .A1(P2_DATAO_REG_11__SCAN_IN), .A2(SI_2_), .A3(
        P1_DATAO_REG_13__SCAN_IN), .A4(P2_DATAO_REG_29__SCAN_IN), .ZN(n9436)
         );
  NOR4_X1 U12118 ( .A1(n10576), .A2(n9471), .A3(n10747), .A4(
        P1_REG3_REG_2__SCAN_IN), .ZN(n9435) );
  NAND4_X1 U12119 ( .A1(n13402), .A2(P3_REG3_REG_27__SCAN_IN), .A3(
        P3_REG1_REG_27__SCAN_IN), .A4(P3_REG0_REG_13__SCAN_IN), .ZN(n9433) );
  NAND2_X1 U12120 ( .A1(P3_REG1_REG_5__SCAN_IN), .A2(P3_REG0_REG_9__SCAN_IN), 
        .ZN(n9431) );
  NOR4_X1 U12121 ( .A1(n9433), .A2(n9432), .A3(n9431), .A4(
        P2_REG1_REG_2__SCAN_IN), .ZN(n9434) );
  NAND4_X1 U12122 ( .A1(n9437), .A2(n9436), .A3(n9435), .A4(n9434), .ZN(n9445)
         );
  NOR4_X1 U12123 ( .A1(P2_REG1_REG_21__SCAN_IN), .A2(P2_REG0_REG_6__SCAN_IN), 
        .A3(P1_IR_REG_10__SCAN_IN), .A4(n15764), .ZN(n9438) );
  NAND3_X1 U12124 ( .A1(P1_D_REG_13__SCAN_IN), .A2(P2_ADDR_REG_9__SCAN_IN), 
        .A3(n9438), .ZN(n9444) );
  NAND4_X1 U12125 ( .A1(P2_REG1_REG_11__SCAN_IN), .A2(P1_REG2_REG_14__SCAN_IN), 
        .A3(n13249), .A4(n13388), .ZN(n9443) );
  NAND4_X1 U12126 ( .A1(P2_IR_REG_15__SCAN_IN), .A2(P1_REG3_REG_21__SCAN_IN), 
        .A3(P1_ADDR_REG_9__SCAN_IN), .A4(P3_DATAO_REG_25__SCAN_IN), .ZN(n9441)
         );
  OR4_X1 U12127 ( .A1(n9441), .A2(n9440), .A3(n9439), .A4(P2_D_REG_20__SCAN_IN), .ZN(n9442) );
  NOR4_X1 U12128 ( .A1(n9445), .A2(n9444), .A3(n9443), .A4(n9442), .ZN(n9467)
         );
  INV_X1 U12129 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n15880) );
  NAND4_X1 U12130 ( .A1(P1_IR_REG_7__SCAN_IN), .A2(P3_DATAO_REG_4__SCAN_IN), 
        .A3(n13435), .A4(n15880), .ZN(n9450) );
  NAND4_X1 U12131 ( .A1(SI_6_), .A2(P1_REG2_REG_20__SCAN_IN), .A3(
        P1_REG2_REG_2__SCAN_IN), .A4(P1_ADDR_REG_17__SCAN_IN), .ZN(n9449) );
  NAND4_X1 U12132 ( .A1(P3_REG2_REG_27__SCAN_IN), .A2(P1_REG3_REG_28__SCAN_IN), 
        .A3(n15971), .A4(n11147), .ZN(n9448) );
  NAND4_X1 U12133 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(P2_D_REG_12__SCAN_IN), 
        .A3(n15136), .A4(n9446), .ZN(n9447) );
  NOR4_X1 U12134 ( .A1(n9450), .A2(n9449), .A3(n9448), .A4(n9447), .ZN(n9466)
         );
  NAND4_X1 U12135 ( .A1(P3_B_REG_SCAN_IN), .A2(P3_REG1_REG_4__SCAN_IN), .A3(
        P1_REG0_REG_1__SCAN_IN), .A4(n9977), .ZN(n9455) );
  NAND4_X1 U12136 ( .A1(P3_ADDR_REG_1__SCAN_IN), .A2(P3_ADDR_REG_2__SCAN_IN), 
        .A3(n15586), .A4(n15562), .ZN(n9454) );
  NAND4_X1 U12137 ( .A1(P3_REG1_REG_16__SCAN_IN), .A2(P2_REG2_REG_31__SCAN_IN), 
        .A3(P3_ADDR_REG_11__SCAN_IN), .A4(n6789), .ZN(n9453) );
  NAND4_X1 U12138 ( .A1(P3_IR_REG_6__SCAN_IN), .A2(P3_DATAO_REG_28__SCAN_IN), 
        .A3(n9451), .A4(n10651), .ZN(n9452) );
  NOR4_X1 U12139 ( .A1(n9455), .A2(n9454), .A3(n9453), .A4(n9452), .ZN(n9465)
         );
  NAND4_X1 U12140 ( .A1(P3_REG3_REG_0__SCAN_IN), .A2(P2_IR_REG_17__SCAN_IN), 
        .A3(P1_IR_REG_26__SCAN_IN), .A4(P1_D_REG_28__SCAN_IN), .ZN(n9456) );
  NOR3_X1 U12141 ( .A1(P3_REG1_REG_30__SCAN_IN), .A2(P3_D_REG_18__SCAN_IN), 
        .A3(n9456), .ZN(n9463) );
  NAND4_X1 U12142 ( .A1(P2_REG1_REG_28__SCAN_IN), .A2(P2_ADDR_REG_16__SCAN_IN), 
        .A3(n12649), .A4(n15576), .ZN(n9461) );
  NAND4_X1 U12143 ( .A1(P3_REG3_REG_6__SCAN_IN), .A2(P1_DATAO_REG_18__SCAN_IN), 
        .A3(P1_REG3_REG_26__SCAN_IN), .A4(n7111), .ZN(n9460) );
  NAND4_X1 U12144 ( .A1(P1_DATAO_REG_12__SCAN_IN), .A2(
        P1_DATAO_REG_16__SCAN_IN), .A3(P2_REG3_REG_22__SCAN_IN), .A4(n15873), 
        .ZN(n9459) );
  NAND4_X1 U12145 ( .A1(P1_REG2_REG_11__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .A3(n15843), .A4(n9457), .ZN(n9458) );
  NOR4_X1 U12146 ( .A1(n9461), .A2(n9460), .A3(n9459), .A4(n9458), .ZN(n9462)
         );
  AND4_X1 U12147 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n9463), .A3(n9462), .A4(
        n15538), .ZN(n9464) );
  NAND4_X1 U12148 ( .A1(n9467), .A2(n9466), .A3(n9465), .A4(n9464), .ZN(n9468)
         );
  AOI21_X1 U12149 ( .B1(n9468), .B2(n10097), .A(keyinput64), .ZN(n9469) );
  NAND3_X1 U12150 ( .A1(n9559), .A2(n9471), .A3(n9568), .ZN(n9472) );
  INV_X1 U12151 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n15886) );
  OR2_X1 U12152 ( .A1(n9523), .A2(n15886), .ZN(n9487) );
  NAND2_X1 U12153 ( .A1(n9599), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n9486) );
  NAND2_X1 U12154 ( .A1(n9552), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n9485) );
  NAND2_X1 U12155 ( .A1(n9550), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n9484) );
  NAND2_X1 U12156 ( .A1(n9489), .A2(n9488), .ZN(n9490) );
  AND2_X1 U12157 ( .A1(n9491), .A2(n9490), .ZN(n14476) );
  MUX2_X1 U12158 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9496), .S(
        P2_IR_REG_20__SCAN_IN), .Z(n9497) );
  AND2_X2 U12159 ( .A1(n10056), .A2(n11964), .ZN(n11353) );
  INV_X1 U12160 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n9499) );
  NAND2_X1 U12161 ( .A1(n11353), .A2(n12056), .ZN(n10193) );
  NOR2_X1 U12162 ( .A1(n10193), .A2(n14164), .ZN(n9504) );
  NAND2_X1 U12163 ( .A1(n10122), .A2(n6529), .ZN(n9508) );
  NAND2_X1 U12164 ( .A1(n11360), .A2(n11353), .ZN(n9505) );
  NAND3_X1 U12165 ( .A1(n13812), .A2(n9856), .A3(n9505), .ZN(n9506) );
  NAND3_X1 U12166 ( .A1(n9508), .A2(n9507), .A3(n9506), .ZN(n9518) );
  NAND2_X1 U12167 ( .A1(n9550), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n9510) );
  NAND2_X1 U12168 ( .A1(n9599), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n9509) );
  INV_X1 U12169 ( .A(n9523), .ZN(n9549) );
  INV_X1 U12170 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n15827) );
  NAND2_X1 U12171 ( .A1(n15827), .A2(n9512), .ZN(n9540) );
  NAND2_X1 U12172 ( .A1(n7675), .A2(n6529), .ZN(n9513) );
  NAND2_X1 U12173 ( .A1(n9514), .A2(n9513), .ZN(n9517) );
  AOI22_X1 U12174 ( .A1(n13810), .A2(n6529), .B1(n7675), .B2(n9856), .ZN(n9515) );
  INV_X1 U12175 ( .A(n9516), .ZN(n9519) );
  NAND2_X1 U12176 ( .A1(n9519), .A2(n8040), .ZN(n9533) );
  NAND2_X1 U12177 ( .A1(n9540), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9520) );
  NAND2_X1 U12178 ( .A1(n9522), .A2(n9856), .ZN(n9529) );
  NAND2_X1 U12179 ( .A1(n10032), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n9527) );
  NAND2_X1 U12180 ( .A1(n9550), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n9526) );
  NAND2_X1 U12181 ( .A1(n9552), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n9525) );
  INV_X2 U12182 ( .A(n9523), .ZN(n10058) );
  NAND2_X1 U12183 ( .A1(n10058), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n9524) );
  NAND2_X1 U12184 ( .A1(n13809), .A2(n9947), .ZN(n9528) );
  NAND2_X1 U12185 ( .A1(n9529), .A2(n9528), .ZN(n9532) );
  AOI22_X1 U12186 ( .A1(n13809), .A2(n9856), .B1(n9947), .B2(n9522), .ZN(n9530) );
  AOI21_X1 U12187 ( .B1(n9533), .B2(n9532), .A(n9530), .ZN(n9531) );
  NOR2_X1 U12188 ( .A1(n9533), .A2(n9532), .ZN(n9534) );
  NAND2_X1 U12189 ( .A1(n10032), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n9539) );
  OR2_X1 U12190 ( .A1(n9535), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n9538) );
  NAND2_X1 U12191 ( .A1(n9552), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n9537) );
  NAND2_X1 U12192 ( .A1(n10058), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n9536) );
  NAND4_X4 U12193 ( .A1(n9539), .A2(n9538), .A3(n9537), .A4(n9536), .ZN(n13808) );
  OAI21_X1 U12194 ( .B1(n9540), .B2(P2_IR_REG_2__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n9541) );
  MUX2_X1 U12195 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9541), .S(
        P2_IR_REG_3__SCAN_IN), .Z(n9544) );
  NAND2_X1 U12196 ( .A1(n9544), .A2(n9543), .ZN(n10693) );
  OR2_X1 U12197 ( .A1(n10590), .A2(n9557), .ZN(n9546) );
  OR2_X1 U12198 ( .A1(n9562), .A2(n10591), .ZN(n9545) );
  OAI211_X2 U12199 ( .C1(n10552), .C2(n10693), .A(n9546), .B(n9545), .ZN(
        n15890) );
  NAND2_X1 U12200 ( .A1(n15890), .A2(n9947), .ZN(n9547) );
  AOI22_X1 U12201 ( .A1(n13808), .A2(n9947), .B1(n15890), .B2(n9856), .ZN(
        n9548) );
  NAND2_X1 U12202 ( .A1(n9549), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n9556) );
  OAI21_X1 U12203 ( .B1(P2_REG3_REG_4__SCAN_IN), .B2(P2_REG3_REG_3__SCAN_IN), 
        .A(n9575), .ZN(n11505) );
  INV_X1 U12204 ( .A(n11505), .ZN(n9551) );
  NAND2_X1 U12205 ( .A1(n9550), .A2(n9551), .ZN(n9555) );
  NAND2_X1 U12206 ( .A1(n9599), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n9554) );
  NAND2_X1 U12207 ( .A1(n9552), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n9553) );
  NAND4_X1 U12208 ( .A1(n9556), .A2(n9555), .A3(n9554), .A4(n9553), .ZN(n13807) );
  INV_X2 U12209 ( .A(n9557), .ZN(n9628) );
  NAND2_X1 U12210 ( .A1(n9628), .A2(n10588), .ZN(n9565) );
  NAND2_X1 U12211 ( .A1(n9543), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9558) );
  MUX2_X1 U12212 ( .A(n9558), .B(P2_IR_REG_31__SCAN_IN), .S(n9559), .Z(n9561)
         );
  INV_X1 U12213 ( .A(n9543), .ZN(n9560) );
  NAND2_X1 U12214 ( .A1(n9560), .A2(n9559), .ZN(n9567) );
  OR2_X1 U12215 ( .A1(n10552), .A2(n13830), .ZN(n9564) );
  INV_X1 U12216 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n10595) );
  OR2_X1 U12217 ( .A1(n9562), .A2(n10595), .ZN(n9563) );
  INV_X1 U12218 ( .A(n11506), .ZN(n10210) );
  AOI22_X1 U12219 ( .A1(n13807), .A2(n9947), .B1(n10210), .B2(n9856), .ZN(
        n9583) );
  NAND2_X1 U12220 ( .A1(n9582), .A2(n9583), .ZN(n9594) );
  NAND2_X1 U12221 ( .A1(n9567), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9566) );
  MUX2_X1 U12222 ( .A(n9566), .B(P2_IR_REG_31__SCAN_IN), .S(n9568), .Z(n9570)
         );
  INV_X1 U12223 ( .A(n9567), .ZN(n9569) );
  NAND2_X1 U12224 ( .A1(n9570), .A2(n9699), .ZN(n13842) );
  INV_X1 U12225 ( .A(n13842), .ZN(n10677) );
  AOI22_X1 U12226 ( .A1(n9834), .A2(P1_DATAO_REG_5__SCAN_IN), .B1(n9833), .B2(
        n10677), .ZN(n9572) );
  NAND2_X1 U12227 ( .A1(n10617), .A2(n9628), .ZN(n9571) );
  NAND2_X1 U12228 ( .A1(n10058), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n9580) );
  INV_X1 U12229 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n9574) );
  NAND2_X1 U12230 ( .A1(n9575), .A2(n9574), .ZN(n9576) );
  NAND2_X1 U12231 ( .A1(n9613), .A2(n9576), .ZN(n11933) );
  OR2_X1 U12232 ( .A1(n9535), .A2(n11933), .ZN(n9579) );
  NAND2_X1 U12233 ( .A1(n9599), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n9578) );
  NAND2_X1 U12234 ( .A1(n9552), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n9577) );
  NAND2_X1 U12235 ( .A1(n13806), .A2(n6529), .ZN(n9581) );
  OAI21_X1 U12236 ( .B1(n10197), .B2(n6529), .A(n9581), .ZN(n9589) );
  AND2_X1 U12237 ( .A1(n9594), .A2(n9589), .ZN(n9592) );
  INV_X1 U12238 ( .A(n9582), .ZN(n9585) );
  INV_X1 U12239 ( .A(n9583), .ZN(n9584) );
  NAND2_X1 U12240 ( .A1(n9585), .A2(n9584), .ZN(n9588) );
  NAND2_X1 U12241 ( .A1(n13807), .A2(n10091), .ZN(n9586) );
  OAI21_X1 U12242 ( .B1(n11506), .B2(n10091), .A(n9586), .ZN(n9587) );
  NAND2_X1 U12243 ( .A1(n9588), .A2(n9587), .ZN(n9596) );
  INV_X1 U12244 ( .A(n9589), .ZN(n9591) );
  AOI22_X1 U12245 ( .A1(n13806), .A2(n10091), .B1(n6529), .B2(n11930), .ZN(
        n9593) );
  INV_X1 U12246 ( .A(n9593), .ZN(n9590) );
  AND2_X1 U12247 ( .A1(n9594), .A2(n9593), .ZN(n9595) );
  NAND2_X1 U12248 ( .A1(n9699), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9597) );
  XNOR2_X1 U12249 ( .A(n9597), .B(P2_IR_REG_6__SCAN_IN), .ZN(n13857) );
  AOI22_X1 U12250 ( .A1(n9834), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n9833), .B2(
        n13857), .ZN(n9598) );
  NAND2_X1 U12251 ( .A1(n12009), .A2(n10091), .ZN(n9605) );
  NAND2_X1 U12252 ( .A1(n9549), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n9603) );
  INV_X1 U12253 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n9612) );
  XNOR2_X1 U12254 ( .A(n9613), .B(n9612), .ZN(n12013) );
  OR2_X1 U12255 ( .A1(n9535), .A2(n12013), .ZN(n9602) );
  INV_X2 U12256 ( .A(n9599), .ZN(n9978) );
  INV_X4 U12257 ( .A(n9978), .ZN(n10032) );
  NAND2_X1 U12258 ( .A1(n10032), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n9601) );
  NAND2_X1 U12259 ( .A1(n9552), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n9600) );
  NAND4_X1 U12260 ( .A1(n9603), .A2(n9602), .A3(n9601), .A4(n9600), .ZN(n13805) );
  NAND2_X1 U12261 ( .A1(n13805), .A2(n9947), .ZN(n9604) );
  NAND2_X1 U12262 ( .A1(n9605), .A2(n9604), .ZN(n9607) );
  AOI22_X1 U12263 ( .A1(n6529), .A2(n12009), .B1(n13805), .B2(n9856), .ZN(
        n9606) );
  NAND2_X1 U12264 ( .A1(n10635), .A2(n9628), .ZN(n9610) );
  NAND2_X1 U12265 ( .A1(n9629), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9608) );
  XNOR2_X1 U12266 ( .A(n9608), .B(P2_IR_REG_7__SCAN_IN), .ZN(n13871) );
  AOI22_X1 U12267 ( .A1(n9834), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n9833), .B2(
        n13871), .ZN(n9609) );
  NAND2_X1 U12268 ( .A1(n12026), .A2(n9947), .ZN(n9622) );
  NAND2_X1 U12269 ( .A1(n10058), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n9620) );
  INV_X1 U12270 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n9611) );
  OAI21_X1 U12271 ( .B1(n9613), .B2(n9612), .A(n9611), .ZN(n9616) );
  NAND2_X1 U12272 ( .A1(n9616), .A2(n9638), .ZN(n12070) );
  OR2_X1 U12273 ( .A1(n9535), .A2(n12070), .ZN(n9619) );
  NAND2_X1 U12274 ( .A1(n10032), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n9618) );
  NAND2_X1 U12275 ( .A1(n9552), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n9617) );
  NAND4_X1 U12276 ( .A1(n9620), .A2(n9619), .A3(n9618), .A4(n9617), .ZN(n13804) );
  NAND2_X1 U12277 ( .A1(n13804), .A2(n10091), .ZN(n9621) );
  NAND2_X1 U12278 ( .A1(n9622), .A2(n9621), .ZN(n9624) );
  AOI22_X1 U12279 ( .A1(n12026), .A2(n10091), .B1(n6529), .B2(n13804), .ZN(
        n9623) );
  NOR2_X1 U12280 ( .A1(n9625), .A2(n9624), .ZN(n9626) );
  INV_X1 U12281 ( .A(n9629), .ZN(n9631) );
  INV_X1 U12282 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n9630) );
  NAND2_X1 U12283 ( .A1(n9631), .A2(n9630), .ZN(n9633) );
  NAND2_X1 U12284 ( .A1(n9633), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9632) );
  MUX2_X1 U12285 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9632), .S(
        P2_IR_REG_8__SCAN_IN), .Z(n9634) );
  AOI22_X1 U12286 ( .A1(n9834), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n9833), .B2(
        n10878), .ZN(n9635) );
  NAND2_X1 U12287 ( .A1(n14264), .A2(n10091), .ZN(n9645) );
  OR2_X1 U12288 ( .A1(n9978), .A2(n10875), .ZN(n9643) );
  INV_X1 U12289 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n9637) );
  NAND2_X1 U12290 ( .A1(n9638), .A2(n9637), .ZN(n9639) );
  NAND2_X1 U12291 ( .A1(n9653), .A2(n9639), .ZN(n12044) );
  OR2_X1 U12292 ( .A1(n9535), .A2(n12044), .ZN(n9642) );
  NAND2_X1 U12293 ( .A1(n10058), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n9641) );
  NAND2_X1 U12294 ( .A1(n9552), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n9640) );
  NAND4_X1 U12295 ( .A1(n9643), .A2(n9642), .A3(n9641), .A4(n9640), .ZN(n13803) );
  NAND2_X1 U12296 ( .A1(n13803), .A2(n9947), .ZN(n9644) );
  NAND2_X1 U12297 ( .A1(n9645), .A2(n9644), .ZN(n9648) );
  NAND2_X1 U12298 ( .A1(n14264), .A2(n9947), .ZN(n9646) );
  OAI21_X1 U12299 ( .B1(n7482), .B2(n6529), .A(n9646), .ZN(n9647) );
  NAND2_X1 U12300 ( .A1(n10664), .A2(n7674), .ZN(n9651) );
  NAND2_X1 U12301 ( .A1(n9667), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9649) );
  XNOR2_X1 U12302 ( .A(n9649), .B(P2_IR_REG_9__SCAN_IN), .ZN(n11177) );
  AOI22_X1 U12303 ( .A1(n9834), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n9833), .B2(
        n11177), .ZN(n9650) );
  NAND2_X1 U12304 ( .A1(n14386), .A2(n9947), .ZN(n9661) );
  NAND2_X1 U12305 ( .A1(n9552), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n9659) );
  INV_X1 U12306 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n11170) );
  OR2_X1 U12307 ( .A1(n9978), .A2(n11170), .ZN(n9658) );
  NAND2_X1 U12308 ( .A1(n9653), .A2(n9652), .ZN(n9654) );
  NAND2_X1 U12309 ( .A1(n9676), .A2(n9654), .ZN(n14249) );
  OR2_X1 U12310 ( .A1(n9535), .A2(n14249), .ZN(n9657) );
  INV_X1 U12311 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n9655) );
  OR2_X1 U12312 ( .A1(n9523), .A2(n9655), .ZN(n9656) );
  NAND2_X1 U12313 ( .A1(n13802), .A2(n10091), .ZN(n9660) );
  NAND2_X1 U12314 ( .A1(n9661), .A2(n9660), .ZN(n9663) );
  AOI22_X1 U12315 ( .A1(n14386), .A2(n10091), .B1(n9947), .B2(n13802), .ZN(
        n9662) );
  NOR2_X1 U12316 ( .A1(n9664), .A2(n9663), .ZN(n9665) );
  NAND2_X1 U12317 ( .A1(n10773), .A2(n9628), .ZN(n9672) );
  INV_X1 U12318 ( .A(n9667), .ZN(n9669) );
  INV_X1 U12319 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n9668) );
  NAND2_X1 U12320 ( .A1(n9669), .A2(n9668), .ZN(n9684) );
  NAND2_X1 U12321 ( .A1(n9684), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9670) );
  AOI22_X1 U12322 ( .A1(n9834), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n9833), 
        .B2(n11655), .ZN(n9671) );
  NAND2_X1 U12323 ( .A1(n14379), .A2(n10091), .ZN(n9683) );
  NAND2_X1 U12324 ( .A1(n10058), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n9681) );
  OR2_X1 U12325 ( .A1(n9978), .A2(n9673), .ZN(n9680) );
  INV_X1 U12326 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n9675) );
  NAND2_X1 U12327 ( .A1(n9676), .A2(n9675), .ZN(n9677) );
  NAND2_X1 U12328 ( .A1(n9704), .A2(n9677), .ZN(n14229) );
  OR2_X1 U12329 ( .A1(n9535), .A2(n14229), .ZN(n9679) );
  INV_X1 U12330 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n14230) );
  OR2_X1 U12331 ( .A1(n10035), .A2(n14230), .ZN(n9678) );
  INV_X1 U12332 ( .A(n13731), .ZN(n13801) );
  NAND2_X1 U12333 ( .A1(n13801), .A2(n9947), .ZN(n9682) );
  NAND2_X1 U12334 ( .A1(n9683), .A2(n9682), .ZN(n9696) );
  NAND2_X1 U12335 ( .A1(n10835), .A2(n9628), .ZN(n9687) );
  OAI21_X1 U12336 ( .B1(n9684), .B2(P2_IR_REG_10__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n9685) );
  XNOR2_X1 U12337 ( .A(n9685), .B(P2_IR_REG_11__SCAN_IN), .ZN(n11826) );
  AOI22_X1 U12338 ( .A1(n9834), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n11826), 
        .B2(n9833), .ZN(n9686) );
  NAND2_X1 U12339 ( .A1(n9549), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n9691) );
  INV_X1 U12340 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n9703) );
  XNOR2_X1 U12341 ( .A(n9704), .B(n9703), .ZN(n14212) );
  OR2_X1 U12342 ( .A1(n9535), .A2(n14212), .ZN(n9690) );
  NAND2_X1 U12343 ( .A1(n10032), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n9689) );
  NAND2_X1 U12344 ( .A1(n9552), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n9688) );
  NAND4_X1 U12345 ( .A1(n9691), .A2(n9690), .A3(n9689), .A4(n9688), .ZN(n13800) );
  AND2_X1 U12346 ( .A1(n13800), .A2(n10091), .ZN(n9692) );
  AOI21_X1 U12347 ( .B1(n14443), .B2(n6529), .A(n9692), .ZN(n9714) );
  NAND2_X1 U12348 ( .A1(n14443), .A2(n10091), .ZN(n9694) );
  NAND2_X1 U12349 ( .A1(n13800), .A2(n9947), .ZN(n9693) );
  NAND2_X1 U12350 ( .A1(n9694), .A2(n9693), .ZN(n9713) );
  AOI22_X1 U12351 ( .A1(n14379), .A2(n9947), .B1(n13801), .B2(n9856), .ZN(
        n9695) );
  OAI21_X1 U12352 ( .B1(n9699), .B2(n9698), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n9700) );
  XNOR2_X1 U12353 ( .A(n9700), .B(P2_IR_REG_12__SCAN_IN), .ZN(n12305) );
  AOI22_X1 U12354 ( .A1(n9834), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n9833), 
        .B2(n12305), .ZN(n9701) );
  NAND2_X1 U12355 ( .A1(n10032), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n9709) );
  INV_X1 U12356 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n9702) );
  OAI21_X1 U12357 ( .B1(n9704), .B2(n9703), .A(n9702), .ZN(n9705) );
  NAND2_X1 U12358 ( .A1(n9705), .A2(n9719), .ZN(n14194) );
  OR2_X1 U12359 ( .A1(n9535), .A2(n14194), .ZN(n9708) );
  NAND2_X1 U12360 ( .A1(n9549), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n9707) );
  NAND2_X1 U12361 ( .A1(n9552), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n9706) );
  NAND4_X1 U12362 ( .A1(n9709), .A2(n9708), .A3(n9707), .A4(n9706), .ZN(n13799) );
  AND2_X1 U12363 ( .A1(n13799), .A2(n10091), .ZN(n9710) );
  AOI21_X1 U12364 ( .B1(n14197), .B2(n6529), .A(n9710), .ZN(n9729) );
  NAND2_X1 U12365 ( .A1(n14197), .A2(n10091), .ZN(n9712) );
  NAND2_X1 U12366 ( .A1(n13799), .A2(n9947), .ZN(n9711) );
  NAND2_X1 U12367 ( .A1(n9712), .A2(n9711), .ZN(n9728) );
  AOI22_X1 U12368 ( .A1(n9729), .A2(n9728), .B1(n9714), .B2(n9713), .ZN(n9715)
         );
  NAND2_X1 U12369 ( .A1(n11247), .A2(n9628), .ZN(n9718) );
  OR2_X1 U12370 ( .A1(n6542), .A2(n14451), .ZN(n9716) );
  XNOR2_X1 U12371 ( .A(n9716), .B(P2_IR_REG_13__SCAN_IN), .ZN(n15849) );
  AOI22_X1 U12372 ( .A1(n9834), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n9833), 
        .B2(n15849), .ZN(n9717) );
  NAND2_X1 U12373 ( .A1(n9549), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n9724) );
  NAND2_X1 U12374 ( .A1(n9719), .A2(n15843), .ZN(n9720) );
  NAND2_X1 U12375 ( .A1(n9784), .A2(n9720), .ZN(n13706) );
  OR2_X1 U12376 ( .A1(n9535), .A2(n13706), .ZN(n9723) );
  NAND2_X1 U12377 ( .A1(n10032), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n9722) );
  NAND2_X1 U12378 ( .A1(n9552), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n9721) );
  NAND4_X1 U12379 ( .A1(n9724), .A2(n9723), .A3(n9722), .A4(n9721), .ZN(n13798) );
  AND2_X1 U12380 ( .A1(n13798), .A2(n6529), .ZN(n9725) );
  AOI21_X1 U12381 ( .B1(n14362), .B2(n10091), .A(n9725), .ZN(n9797) );
  NAND2_X1 U12382 ( .A1(n14362), .A2(n9947), .ZN(n9727) );
  NAND2_X1 U12383 ( .A1(n13798), .A2(n10091), .ZN(n9726) );
  NAND2_X1 U12384 ( .A1(n9727), .A2(n9726), .ZN(n9796) );
  INV_X1 U12385 ( .A(n9728), .ZN(n9731) );
  INV_X1 U12386 ( .A(n9729), .ZN(n9730) );
  AOI22_X1 U12387 ( .A1(n9797), .A2(n9796), .B1(n9731), .B2(n9730), .ZN(n9795)
         );
  NAND2_X1 U12388 ( .A1(n11404), .A2(n7674), .ZN(n9734) );
  OR2_X1 U12389 ( .A1(n10096), .A2(n14451), .ZN(n9732) );
  XNOR2_X1 U12390 ( .A(n9732), .B(P2_IR_REG_17__SCAN_IN), .ZN(n13936) );
  AOI22_X1 U12391 ( .A1(n9834), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n9833), 
        .B2(n13936), .ZN(n9733) );
  NAND2_X1 U12392 ( .A1(n10058), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n9741) );
  INV_X1 U12393 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n9783) );
  INV_X1 U12394 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n9767) );
  INV_X1 U12395 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n9736) );
  NAND2_X1 U12396 ( .A1(n9753), .A2(n9736), .ZN(n9737) );
  NAND2_X1 U12397 ( .A1(n9821), .A2(n9737), .ZN(n14132) );
  OR2_X1 U12398 ( .A1(n9535), .A2(n14132), .ZN(n9740) );
  NAND2_X1 U12399 ( .A1(n10032), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n9739) );
  NAND2_X1 U12400 ( .A1(n9552), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n9738) );
  NAND4_X1 U12401 ( .A1(n9741), .A2(n9740), .A3(n9739), .A4(n9738), .ZN(n13794) );
  AOI22_X1 U12402 ( .A1(n14341), .A2(n10091), .B1(n6529), .B2(n13794), .ZN(
        n9744) );
  NAND2_X1 U12403 ( .A1(n14341), .A2(n9947), .ZN(n9743) );
  NAND2_X1 U12404 ( .A1(n13794), .A2(n10091), .ZN(n9742) );
  NAND2_X1 U12405 ( .A1(n9743), .A2(n9742), .ZN(n9804) );
  NAND2_X1 U12406 ( .A1(n9744), .A2(n9804), .ZN(n9762) );
  NAND2_X1 U12407 ( .A1(n11291), .A2(n9628), .ZN(n9750) );
  INV_X1 U12408 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n9745) );
  NAND2_X1 U12409 ( .A1(n6542), .A2(n9745), .ZN(n9779) );
  OR2_X1 U12410 ( .A1(n9779), .A2(P2_IR_REG_14__SCAN_IN), .ZN(n9763) );
  OAI21_X1 U12411 ( .B1(n9763), .B2(P2_IR_REG_15__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n9746) );
  MUX2_X1 U12412 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9746), .S(
        P2_IR_REG_16__SCAN_IN), .Z(n9748) );
  INV_X1 U12413 ( .A(n10096), .ZN(n9747) );
  NAND2_X1 U12414 ( .A1(n9748), .A2(n9747), .ZN(n13916) );
  INV_X1 U12415 ( .A(n13916), .ZN(n13908) );
  AOI22_X1 U12416 ( .A1(n9834), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n9833), 
        .B2(n13908), .ZN(n9749) );
  NAND2_X1 U12417 ( .A1(n10058), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n9757) );
  INV_X1 U12418 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n9751) );
  NAND2_X1 U12419 ( .A1(n9769), .A2(n9751), .ZN(n9752) );
  NAND2_X1 U12420 ( .A1(n9753), .A2(n9752), .ZN(n14149) );
  OR2_X1 U12421 ( .A1(n9535), .A2(n14149), .ZN(n9756) );
  NAND2_X1 U12422 ( .A1(n10032), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n9755) );
  NAND2_X1 U12423 ( .A1(n9552), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n9754) );
  NAND4_X1 U12424 ( .A1(n9757), .A2(n9756), .A3(n9755), .A4(n9754), .ZN(n13795) );
  AND2_X1 U12425 ( .A1(n13795), .A2(n6529), .ZN(n9758) );
  AOI21_X1 U12426 ( .B1(n14148), .B2(n10091), .A(n9758), .ZN(n9801) );
  NAND2_X1 U12427 ( .A1(n14148), .A2(n9947), .ZN(n9760) );
  NAND2_X1 U12428 ( .A1(n13795), .A2(n10091), .ZN(n9759) );
  NAND2_X1 U12429 ( .A1(n9760), .A2(n9759), .ZN(n9800) );
  NAND2_X1 U12430 ( .A1(n9801), .A2(n9800), .ZN(n9761) );
  NAND2_X1 U12431 ( .A1(n9763), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9764) );
  XNOR2_X1 U12432 ( .A(n9764), .B(P2_IR_REG_15__SCAN_IN), .ZN(n13893) );
  AOI22_X1 U12433 ( .A1(n9834), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n9833), 
        .B2(n13893), .ZN(n9765) );
  NAND2_X1 U12434 ( .A1(n10058), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n9774) );
  INV_X1 U12435 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n9766) );
  OR2_X1 U12436 ( .A1(n9978), .A2(n9766), .ZN(n9773) );
  NAND2_X1 U12437 ( .A1(n9786), .A2(n9767), .ZN(n9768) );
  NAND2_X1 U12438 ( .A1(n9769), .A2(n9768), .ZN(n14166) );
  OR2_X1 U12439 ( .A1(n9535), .A2(n14166), .ZN(n9772) );
  INV_X1 U12440 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n9770) );
  OR2_X1 U12441 ( .A1(n10035), .A2(n9770), .ZN(n9771) );
  NOR2_X1 U12442 ( .A1(n13670), .A2(n9856), .ZN(n9775) );
  AOI21_X1 U12443 ( .B1(n14351), .B2(n10091), .A(n9775), .ZN(n9803) );
  INV_X1 U12444 ( .A(n13670), .ZN(n13796) );
  NAND2_X1 U12445 ( .A1(n13796), .A2(n10091), .ZN(n9776) );
  NAND2_X1 U12446 ( .A1(n9777), .A2(n9776), .ZN(n9802) );
  NAND2_X1 U12447 ( .A1(n9803), .A2(n9802), .ZN(n9778) );
  NAND2_X1 U12448 ( .A1(n9806), .A2(n9778), .ZN(n9810) );
  NAND2_X1 U12449 ( .A1(n11446), .A2(n7674), .ZN(n9782) );
  NAND2_X1 U12450 ( .A1(n9779), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9780) );
  XNOR2_X1 U12451 ( .A(n9780), .B(P2_IR_REG_14__SCAN_IN), .ZN(n13885) );
  AOI22_X1 U12452 ( .A1(n9834), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n9833), 
        .B2(n13885), .ZN(n9781) );
  NAND2_X1 U12453 ( .A1(n10032), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n9790) );
  NAND2_X1 U12454 ( .A1(n9784), .A2(n9783), .ZN(n9785) );
  NAND2_X1 U12455 ( .A1(n9786), .A2(n9785), .ZN(n14173) );
  OR2_X1 U12456 ( .A1(n9535), .A2(n14173), .ZN(n9789) );
  NAND2_X1 U12457 ( .A1(n10058), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n9788) );
  NAND2_X1 U12458 ( .A1(n9552), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n9787) );
  NAND4_X1 U12459 ( .A1(n9790), .A2(n9789), .A3(n9788), .A4(n9787), .ZN(n13797) );
  AND2_X1 U12460 ( .A1(n13797), .A2(n9947), .ZN(n9791) );
  AOI21_X1 U12461 ( .B1(n14435), .B2(n10091), .A(n9791), .ZN(n9809) );
  NAND2_X1 U12462 ( .A1(n14435), .A2(n9947), .ZN(n9793) );
  NAND2_X1 U12463 ( .A1(n13797), .A2(n10091), .ZN(n9792) );
  NAND2_X1 U12464 ( .A1(n9793), .A2(n9792), .ZN(n9808) );
  AND2_X1 U12465 ( .A1(n9809), .A2(n9808), .ZN(n9794) );
  INV_X1 U12466 ( .A(n9796), .ZN(n9799) );
  INV_X1 U12467 ( .A(n9797), .ZN(n9798) );
  NAND2_X1 U12468 ( .A1(n9799), .A2(n9798), .ZN(n9813) );
  OAI22_X1 U12469 ( .A1(n9803), .A2(n9802), .B1(n9801), .B2(n9800), .ZN(n9807)
         );
  INV_X1 U12470 ( .A(n9804), .ZN(n9805) );
  AOI22_X1 U12471 ( .A1(n9807), .A2(n9806), .B1(n9805), .B2(n10173), .ZN(n9812) );
  OR3_X1 U12472 ( .A1(n9810), .A2(n9809), .A3(n9808), .ZN(n9811) );
  OAI211_X1 U12473 ( .C1(n6562), .C2(n9813), .A(n9812), .B(n9811), .ZN(n9814)
         );
  INV_X1 U12474 ( .A(n9814), .ZN(n9815) );
  NAND2_X1 U12475 ( .A1(n11754), .A2(n9628), .ZN(n9819) );
  NAND2_X1 U12476 ( .A1(n9816), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9817) );
  XNOR2_X1 U12477 ( .A(n9817), .B(n6920), .ZN(n15870) );
  INV_X1 U12478 ( .A(n15870), .ZN(n13931) );
  AOI22_X1 U12479 ( .A1(n9834), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n9833), 
        .B2(n13931), .ZN(n9818) );
  NAND2_X2 U12480 ( .A1(n9819), .A2(n9818), .ZN(n14335) );
  NAND2_X1 U12481 ( .A1(n14335), .A2(n10091), .ZN(n9829) );
  INV_X1 U12482 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n9820) );
  NAND2_X1 U12483 ( .A1(n9821), .A2(n9820), .ZN(n9822) );
  AND2_X1 U12484 ( .A1(n9838), .A2(n9822), .ZN(n14115) );
  NAND2_X1 U12485 ( .A1(n14115), .A2(n9550), .ZN(n9827) );
  NAND2_X1 U12486 ( .A1(n10058), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n9824) );
  NAND2_X1 U12487 ( .A1(n10032), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n9823) );
  AND2_X1 U12488 ( .A1(n9824), .A2(n9823), .ZN(n9826) );
  NAND2_X1 U12489 ( .A1(n9552), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n9825) );
  OR2_X1 U12490 ( .A1(n12686), .A2(n9856), .ZN(n9828) );
  NAND2_X1 U12491 ( .A1(n9829), .A2(n9828), .ZN(n9832) );
  NAND2_X1 U12492 ( .A1(n14335), .A2(n9947), .ZN(n9830) );
  OAI21_X1 U12493 ( .B1(n12686), .B2(n6529), .A(n9830), .ZN(n9831) );
  AOI22_X1 U12494 ( .A1(n9834), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n11354), 
        .B2(n9833), .ZN(n9835) );
  NAND2_X1 U12495 ( .A1(n14097), .A2(n9947), .ZN(n9843) );
  INV_X1 U12496 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n14099) );
  INV_X1 U12497 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n9837) );
  NAND2_X1 U12498 ( .A1(n9838), .A2(n9837), .ZN(n9839) );
  NAND2_X1 U12499 ( .A1(n9862), .A2(n9839), .ZN(n14098) );
  OR2_X1 U12500 ( .A1(n14098), .A2(n9535), .ZN(n9841) );
  AOI22_X1 U12501 ( .A1(n10058), .A2(P2_REG0_REG_19__SCAN_IN), .B1(n10032), 
        .B2(P2_REG1_REG_19__SCAN_IN), .ZN(n9840) );
  OAI211_X1 U12502 ( .C1(n10035), .C2(n14099), .A(n9841), .B(n9840), .ZN(
        n13792) );
  NAND2_X1 U12503 ( .A1(n13792), .A2(n10091), .ZN(n9842) );
  NAND2_X1 U12504 ( .A1(n9843), .A2(n9842), .ZN(n9845) );
  AOI22_X1 U12505 ( .A1(n14097), .A2(n10091), .B1(n6529), .B2(n13792), .ZN(
        n9844) );
  NAND2_X1 U12506 ( .A1(n11961), .A2(n9628), .ZN(n9847) );
  OR2_X1 U12507 ( .A1(n10053), .A2(n11966), .ZN(n9846) );
  NAND2_X1 U12508 ( .A1(n14325), .A2(n10091), .ZN(n9855) );
  XNOR2_X1 U12509 ( .A(n9862), .B(P2_REG3_REG_20__SCAN_IN), .ZN(n14086) );
  NAND2_X1 U12510 ( .A1(n14086), .A2(n9550), .ZN(n9853) );
  INV_X1 U12511 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n9850) );
  NAND2_X1 U12512 ( .A1(n10058), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n9849) );
  NAND2_X1 U12513 ( .A1(n10032), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n9848) );
  OAI211_X1 U12514 ( .C1(n9850), .C2(n10035), .A(n9849), .B(n9848), .ZN(n9851)
         );
  INV_X1 U12515 ( .A(n9851), .ZN(n9852) );
  NAND2_X1 U12516 ( .A1(n9853), .A2(n9852), .ZN(n13791) );
  NAND2_X1 U12517 ( .A1(n13791), .A2(n9947), .ZN(n9854) );
  NAND2_X1 U12518 ( .A1(n9855), .A2(n9854), .ZN(n9858) );
  AOI22_X1 U12519 ( .A1(n14325), .A2(n9947), .B1(n13791), .B2(n9856), .ZN(
        n9857) );
  NAND2_X1 U12520 ( .A1(n12050), .A2(n7674), .ZN(n9860) );
  OR2_X1 U12521 ( .A1(n10053), .A2(n12054), .ZN(n9859) );
  NAND2_X1 U12522 ( .A1(n14320), .A2(n9947), .ZN(n9871) );
  INV_X1 U12523 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n13693) );
  INV_X1 U12524 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n13634) );
  OAI21_X1 U12525 ( .B1(n9862), .B2(n13693), .A(n13634), .ZN(n9863) );
  NAND2_X1 U12526 ( .A1(P2_REG3_REG_20__SCAN_IN), .A2(P2_REG3_REG_21__SCAN_IN), 
        .ZN(n9861) );
  AND2_X1 U12527 ( .A1(n9863), .A2(n9878), .ZN(n14072) );
  NAND2_X1 U12528 ( .A1(n14072), .A2(n9550), .ZN(n9869) );
  NAND2_X1 U12529 ( .A1(n10058), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n9865) );
  NAND2_X1 U12530 ( .A1(n9552), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n9864) );
  OAI211_X1 U12531 ( .C1(n9978), .C2(n9866), .A(n9865), .B(n9864), .ZN(n9867)
         );
  INV_X1 U12532 ( .A(n9867), .ZN(n9868) );
  NAND2_X1 U12533 ( .A1(n9869), .A2(n9868), .ZN(n13790) );
  NAND2_X1 U12534 ( .A1(n13790), .A2(n10091), .ZN(n9870) );
  AOI22_X1 U12535 ( .A1(n14320), .A2(n10091), .B1(n6529), .B2(n13790), .ZN(
        n9872) );
  XNOR2_X1 U12536 ( .A(n9874), .B(n9873), .ZN(n12055) );
  NAND2_X1 U12537 ( .A1(n12055), .A2(n9628), .ZN(n9876) );
  OR2_X1 U12538 ( .A1(n10053), .A2(n12058), .ZN(n9875) );
  NAND2_X1 U12539 ( .A1(n14417), .A2(n10091), .ZN(n9887) );
  NAND2_X1 U12540 ( .A1(n9878), .A2(n13722), .ZN(n9879) );
  NAND2_X1 U12541 ( .A1(n9908), .A2(n9879), .ZN(n14052) );
  OR2_X1 U12542 ( .A1(n14052), .A2(n9535), .ZN(n9885) );
  INV_X1 U12543 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n9882) );
  NAND2_X1 U12544 ( .A1(n9549), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n9881) );
  NAND2_X1 U12545 ( .A1(n9599), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n9880) );
  OAI211_X1 U12546 ( .C1(n9882), .C2(n10035), .A(n9881), .B(n9880), .ZN(n9883)
         );
  INV_X1 U12547 ( .A(n9883), .ZN(n9884) );
  NAND2_X1 U12548 ( .A1(n13789), .A2(n9947), .ZN(n9886) );
  NAND2_X1 U12549 ( .A1(n9887), .A2(n9886), .ZN(n9889) );
  AOI22_X1 U12550 ( .A1(n14417), .A2(n9947), .B1(n13789), .B2(n10091), .ZN(
        n9888) );
  NAND2_X1 U12551 ( .A1(n12166), .A2(n7674), .ZN(n9892) );
  INV_X1 U12552 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n12169) );
  OR2_X1 U12553 ( .A1(n10053), .A2(n12169), .ZN(n9891) );
  NAND2_X1 U12554 ( .A1(n14039), .A2(n9947), .ZN(n9900) );
  XNOR2_X1 U12555 ( .A(n9908), .B(P2_REG3_REG_23__SCAN_IN), .ZN(n14033) );
  NAND2_X1 U12556 ( .A1(n14033), .A2(n9550), .ZN(n9898) );
  INV_X1 U12557 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n9895) );
  NAND2_X1 U12558 ( .A1(n10058), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n9894) );
  NAND2_X1 U12559 ( .A1(n10032), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n9893) );
  OAI211_X1 U12560 ( .C1(n9895), .C2(n10035), .A(n9894), .B(n9893), .ZN(n9896)
         );
  INV_X1 U12561 ( .A(n9896), .ZN(n9897) );
  NAND2_X1 U12562 ( .A1(n13788), .A2(n10091), .ZN(n9899) );
  NAND2_X1 U12563 ( .A1(n9900), .A2(n9899), .ZN(n9902) );
  AOI22_X1 U12564 ( .A1(n14039), .A2(n10091), .B1(n6529), .B2(n13788), .ZN(
        n9901) );
  OR2_X1 U12565 ( .A1(n10053), .A2(n14473), .ZN(n9903) );
  NAND2_X1 U12566 ( .A1(n7324), .A2(n10091), .ZN(n9917) );
  INV_X1 U12567 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n9906) );
  INV_X1 U12568 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n9905) );
  OAI21_X1 U12569 ( .B1(n9908), .B2(n9906), .A(n9905), .ZN(n9909) );
  NAND2_X1 U12570 ( .A1(P2_REG3_REG_24__SCAN_IN), .A2(P2_REG3_REG_23__SCAN_IN), 
        .ZN(n9907) );
  NAND2_X1 U12571 ( .A1(n9909), .A2(n10029), .ZN(n13688) );
  OR2_X1 U12572 ( .A1(n13688), .A2(n9535), .ZN(n9915) );
  INV_X1 U12573 ( .A(P2_REG2_REG_24__SCAN_IN), .ZN(n9912) );
  NAND2_X1 U12574 ( .A1(n10032), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n9911) );
  NAND2_X1 U12575 ( .A1(n10058), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n9910) );
  OAI211_X1 U12576 ( .C1(n9912), .C2(n10035), .A(n9911), .B(n9910), .ZN(n9913)
         );
  INV_X1 U12577 ( .A(n9913), .ZN(n9914) );
  NAND2_X1 U12578 ( .A1(n13787), .A2(n9947), .ZN(n9916) );
  NAND2_X1 U12579 ( .A1(n9917), .A2(n9916), .ZN(n9918) );
  AOI22_X1 U12580 ( .A1(n7324), .A2(n9947), .B1(n13787), .B2(n10091), .ZN(
        n9920) );
  INV_X1 U12581 ( .A(SI_24_), .ZN(n12294) );
  MUX2_X1 U12582 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(P1_DATAO_REG_25__SCAN_IN), 
        .S(n6533), .Z(n9924) );
  NAND2_X1 U12583 ( .A1(n9924), .A2(SI_25_), .ZN(n10027) );
  OAI21_X1 U12584 ( .B1(n9923), .B2(n12294), .A(n10027), .ZN(n9921) );
  INV_X1 U12585 ( .A(n9921), .ZN(n9922) );
  INV_X1 U12586 ( .A(n9923), .ZN(n10020) );
  NOR2_X1 U12587 ( .A1(n10020), .A2(SI_24_), .ZN(n9927) );
  INV_X1 U12588 ( .A(n9924), .ZN(n9925) );
  INV_X1 U12589 ( .A(SI_25_), .ZN(n13527) );
  NAND2_X1 U12590 ( .A1(n9925), .A2(n13527), .ZN(n10026) );
  INV_X1 U12591 ( .A(n10026), .ZN(n9926) );
  AOI21_X1 U12592 ( .B1(n9927), .B2(n10027), .A(n9926), .ZN(n9928) );
  MUX2_X1 U12593 ( .A(n15540), .B(n14465), .S(n6532), .Z(n10002) );
  INV_X1 U12594 ( .A(n10002), .ZN(n9930) );
  MUX2_X1 U12595 ( .A(n15538), .B(n14463), .S(n6533), .Z(n9986) );
  INV_X1 U12596 ( .A(n9986), .ZN(n9931) );
  OAI22_X1 U12597 ( .A1(n9930), .A2(SI_26_), .B1(n9931), .B2(SI_27_), .ZN(
        n9934) );
  INV_X1 U12598 ( .A(SI_26_), .ZN(n13522) );
  INV_X1 U12599 ( .A(SI_27_), .ZN(n13517) );
  OAI21_X1 U12600 ( .B1(n10002), .B2(n13522), .A(n13517), .ZN(n9932) );
  AND2_X1 U12601 ( .A1(SI_26_), .A2(SI_27_), .ZN(n9929) );
  AOI22_X1 U12602 ( .A1(n9932), .A2(n9931), .B1(n9930), .B2(n9929), .ZN(n9933)
         );
  MUX2_X1 U12603 ( .A(n15535), .B(n9938), .S(n6533), .Z(n9935) );
  NAND2_X1 U12604 ( .A1(n9935), .A2(n13514), .ZN(n9952) );
  INV_X1 U12605 ( .A(n9935), .ZN(n9936) );
  NAND2_X1 U12606 ( .A1(n9936), .A2(SI_28_), .ZN(n9937) );
  NAND2_X1 U12607 ( .A1(n9952), .A2(n9937), .ZN(n9950) );
  NAND2_X1 U12608 ( .A1(n14456), .A2(n7674), .ZN(n9940) );
  OR2_X1 U12609 ( .A1(n10053), .A2(n9938), .ZN(n9939) );
  INV_X1 U12610 ( .A(n10009), .ZN(n9941) );
  NAND2_X1 U12611 ( .A1(n9941), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n9992) );
  NAND2_X1 U12612 ( .A1(n9992), .A2(n9423), .ZN(n9942) );
  NAND2_X1 U12613 ( .A1(n9552), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n9944) );
  NAND2_X1 U12614 ( .A1(n10058), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n9943) );
  OAI211_X1 U12615 ( .C1(n9978), .C2(n12395), .A(n9944), .B(n9943), .ZN(n9945)
         );
  NOR2_X1 U12616 ( .A1(n13614), .A2(n9856), .ZN(n9946) );
  AOI21_X1 U12617 ( .B1(n13972), .B2(n10091), .A(n9946), .ZN(n10074) );
  NAND2_X1 U12618 ( .A1(n13972), .A2(n9947), .ZN(n9949) );
  OR2_X1 U12619 ( .A1(n13614), .A2(n9947), .ZN(n9948) );
  MUX2_X1 U12620 ( .A(n15530), .B(n14454), .S(n6532), .Z(n9955) );
  XNOR2_X1 U12621 ( .A(n9955), .B(SI_29_), .ZN(n9971) );
  INV_X1 U12622 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n14843) );
  INV_X1 U12623 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n12774) );
  MUX2_X1 U12624 ( .A(n14843), .B(n12774), .S(n6532), .Z(n9954) );
  NOR2_X1 U12625 ( .A1(n9954), .A2(n12649), .ZN(n9958) );
  MUX2_X1 U12626 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n6533), .Z(n9953) );
  XNOR2_X1 U12627 ( .A(n9953), .B(SI_31_), .ZN(n9959) );
  NAND2_X1 U12628 ( .A1(n9954), .A2(n12649), .ZN(n10049) );
  INV_X1 U12629 ( .A(SI_29_), .ZN(n13512) );
  NAND2_X1 U12630 ( .A1(n9955), .A2(n13512), .ZN(n10047) );
  NAND2_X1 U12631 ( .A1(n10049), .A2(n10047), .ZN(n9960) );
  INV_X1 U12632 ( .A(n9959), .ZN(n9956) );
  NOR2_X1 U12633 ( .A1(n9960), .A2(n9956), .ZN(n9957) );
  INV_X1 U12634 ( .A(n9958), .ZN(n10050) );
  XNOR2_X1 U12635 ( .A(n9959), .B(n10050), .ZN(n9962) );
  NOR2_X1 U12636 ( .A1(n9960), .A2(n9959), .ZN(n9961) );
  OR2_X1 U12637 ( .A1(n9962), .A2(n9961), .ZN(n9963) );
  OR2_X1 U12638 ( .A1(n10053), .A2(n12419), .ZN(n9966) );
  NAND2_X1 U12639 ( .A1(n9599), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n9970) );
  NAND2_X1 U12640 ( .A1(n9552), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n9969) );
  NAND2_X1 U12641 ( .A1(n10058), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n9968) );
  NAND3_X1 U12642 ( .A1(n9970), .A2(n9969), .A3(n9968), .ZN(n13781) );
  XNOR2_X1 U12643 ( .A(n12769), .B(n13781), .ZN(n10073) );
  NAND2_X1 U12644 ( .A1(n14861), .A2(n9628), .ZN(n9974) );
  OR2_X1 U12645 ( .A1(n10053), .A2(n14454), .ZN(n9973) );
  NAND2_X1 U12646 ( .A1(n10058), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n9976) );
  NAND2_X1 U12647 ( .A1(n9552), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n9975) );
  OAI211_X1 U12648 ( .C1(n9978), .C2(n9977), .A(n9976), .B(n9975), .ZN(n9979)
         );
  INV_X1 U12649 ( .A(n9979), .ZN(n9980) );
  OAI21_X1 U12650 ( .B1(n13959), .B2(n9535), .A(n9980), .ZN(n13782) );
  AND2_X1 U12651 ( .A1(n13782), .A2(n10091), .ZN(n9981) );
  AOI21_X1 U12652 ( .B1(n12384), .B2(n6529), .A(n9981), .ZN(n10068) );
  NAND2_X1 U12653 ( .A1(n12384), .A2(n10091), .ZN(n9983) );
  NAND2_X1 U12654 ( .A1(n13782), .A2(n9947), .ZN(n9982) );
  NAND2_X1 U12655 ( .A1(n9983), .A2(n9982), .ZN(n10067) );
  NAND2_X1 U12656 ( .A1(n10004), .A2(n13522), .ZN(n9984) );
  NAND2_X1 U12657 ( .A1(n9985), .A2(n9984), .ZN(n9988) );
  XNOR2_X1 U12658 ( .A(n9986), .B(SI_27_), .ZN(n9987) );
  OR2_X1 U12659 ( .A1(n10053), .A2(n14463), .ZN(n9989) );
  INV_X1 U12660 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n13568) );
  NAND2_X1 U12661 ( .A1(n10009), .A2(n13568), .ZN(n9991) );
  NAND2_X1 U12662 ( .A1(n9992), .A2(n9991), .ZN(n13983) );
  NAND2_X1 U12663 ( .A1(n10058), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n9994) );
  NAND2_X1 U12664 ( .A1(n9599), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n9993) );
  OAI211_X1 U12665 ( .C1(n9402), .C2(n10035), .A(n9994), .B(n9993), .ZN(n9995)
         );
  INV_X1 U12666 ( .A(n9995), .ZN(n9996) );
  AND2_X1 U12667 ( .A1(n13784), .A2(n10091), .ZN(n9998) );
  AOI21_X1 U12668 ( .B1(n14405), .B2(n6529), .A(n9998), .ZN(n10070) );
  NAND2_X1 U12669 ( .A1(n14405), .A2(n10091), .ZN(n10000) );
  NAND2_X1 U12670 ( .A1(n13784), .A2(n9947), .ZN(n9999) );
  NAND2_X1 U12671 ( .A1(n10000), .A2(n9999), .ZN(n10069) );
  AND2_X1 U12672 ( .A1(n10070), .A2(n10069), .ZN(n10001) );
  XNOR2_X1 U12673 ( .A(n10002), .B(SI_26_), .ZN(n10003) );
  NAND2_X1 U12674 ( .A1(n14464), .A2(n9628), .ZN(n10006) );
  OR2_X1 U12675 ( .A1(n10053), .A2(n14465), .ZN(n10005) );
  INV_X1 U12676 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n10007) );
  NAND2_X1 U12677 ( .A1(n10031), .A2(n10007), .ZN(n10008) );
  NAND2_X1 U12678 ( .A1(n13998), .A2(n9550), .ZN(n10015) );
  INV_X1 U12679 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n10012) );
  NAND2_X1 U12680 ( .A1(n10058), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n10011) );
  NAND2_X1 U12681 ( .A1(n10032), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n10010) );
  OAI211_X1 U12682 ( .C1(n10012), .C2(n10035), .A(n10011), .B(n10010), .ZN(
        n10013) );
  INV_X1 U12683 ( .A(n10013), .ZN(n10014) );
  AND2_X1 U12684 ( .A1(n13785), .A2(n10091), .ZN(n10016) );
  AOI21_X1 U12685 ( .B1(n13995), .B2(n6529), .A(n10016), .ZN(n10081) );
  NAND2_X1 U12686 ( .A1(n13995), .A2(n10091), .ZN(n10018) );
  NAND2_X1 U12687 ( .A1(n13785), .A2(n6529), .ZN(n10017) );
  NAND2_X1 U12688 ( .A1(n10018), .A2(n10017), .ZN(n10080) );
  AND2_X1 U12689 ( .A1(n10081), .A2(n10080), .ZN(n10019) );
  NAND2_X1 U12690 ( .A1(n10021), .A2(n10020), .ZN(n10025) );
  INV_X1 U12691 ( .A(n10022), .ZN(n10023) );
  NAND2_X1 U12692 ( .A1(n10023), .A2(SI_24_), .ZN(n10024) );
  NAND2_X1 U12693 ( .A1(n10027), .A2(n10026), .ZN(n10028) );
  NAND2_X1 U12694 ( .A1(n7352), .A2(n6529), .ZN(n10039) );
  NAND2_X1 U12695 ( .A1(n10029), .A2(n13659), .ZN(n10030) );
  NAND2_X1 U12696 ( .A1(n10031), .A2(n10030), .ZN(n14010) );
  INV_X1 U12697 ( .A(P2_REG2_REG_25__SCAN_IN), .ZN(n14009) );
  NAND2_X1 U12698 ( .A1(n10058), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n10034) );
  NAND2_X1 U12699 ( .A1(n10032), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n10033) );
  OAI211_X1 U12700 ( .C1(n14009), .C2(n10035), .A(n10034), .B(n10033), .ZN(
        n10036) );
  INV_X1 U12701 ( .A(n10036), .ZN(n10037) );
  NAND2_X1 U12702 ( .A1(n13786), .A2(n10091), .ZN(n10038) );
  NAND2_X1 U12703 ( .A1(n10039), .A2(n10038), .ZN(n10044) );
  INV_X1 U12704 ( .A(n10044), .ZN(n10042) );
  AND2_X1 U12705 ( .A1(n13786), .A2(n9947), .ZN(n10040) );
  AOI21_X1 U12706 ( .B1(n7352), .B2(n10091), .A(n10040), .ZN(n10045) );
  NAND2_X1 U12707 ( .A1(n10042), .A2(n10041), .ZN(n10043) );
  NAND3_X1 U12708 ( .A1(n10046), .A2(n10045), .A3(n10044), .ZN(n10087) );
  INV_X1 U12709 ( .A(n13781), .ZN(n10092) );
  NAND2_X1 U12710 ( .A1(n10048), .A2(n10047), .ZN(n10052) );
  AND2_X1 U12711 ( .A1(n10050), .A2(n10049), .ZN(n10051) );
  NAND2_X1 U12712 ( .A1(n14842), .A2(n9628), .ZN(n10055) );
  OR2_X1 U12713 ( .A1(n10053), .A2(n12774), .ZN(n10054) );
  INV_X1 U12714 ( .A(n12056), .ZN(n10191) );
  NAND2_X1 U12715 ( .A1(n11354), .A2(n10191), .ZN(n10252) );
  INV_X1 U12716 ( .A(n10252), .ZN(n10057) );
  NAND2_X1 U12717 ( .A1(n14164), .A2(n11964), .ZN(n11014) );
  NAND2_X1 U12718 ( .A1(n11014), .A2(n10140), .ZN(n10268) );
  AOI21_X1 U12719 ( .B1(n10057), .B2(n11964), .A(n10268), .ZN(n10063) );
  NAND2_X1 U12720 ( .A1(n13781), .A2(n10091), .ZN(n10062) );
  NAND2_X1 U12721 ( .A1(n10032), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n10061) );
  NAND2_X1 U12722 ( .A1(n9552), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n10060) );
  NAND2_X1 U12723 ( .A1(n10058), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n10059) );
  AND3_X1 U12724 ( .A1(n10061), .A2(n10060), .A3(n10059), .ZN(n12380) );
  AOI21_X1 U12725 ( .B1(n10063), .B2(n10062), .A(n12380), .ZN(n10064) );
  AOI21_X1 U12726 ( .B1(n14401), .B2(n6529), .A(n10064), .ZN(n10090) );
  NAND2_X1 U12727 ( .A1(n14401), .A2(n10091), .ZN(n10066) );
  OR2_X1 U12728 ( .A1(n12380), .A2(n9856), .ZN(n10065) );
  NAND2_X1 U12729 ( .A1(n10066), .A2(n10065), .ZN(n10089) );
  OAI22_X1 U12730 ( .A1(n10090), .A2(n10089), .B1(n10068), .B2(n10067), .ZN(
        n10078) );
  INV_X1 U12731 ( .A(n10072), .ZN(n10076) );
  INV_X1 U12732 ( .A(n10073), .ZN(n10135) );
  INV_X1 U12733 ( .A(n10074), .ZN(n10075) );
  INV_X1 U12734 ( .A(n10079), .ZN(n10084) );
  INV_X1 U12735 ( .A(n10080), .ZN(n10083) );
  INV_X1 U12736 ( .A(n10081), .ZN(n10082) );
  NAND3_X1 U12737 ( .A1(n10084), .A2(n10083), .A3(n10082), .ZN(n10085) );
  NOR3_X1 U12738 ( .A1(n13945), .A2(n6529), .A3(n13781), .ZN(n10094) );
  NOR3_X1 U12739 ( .A1(n12769), .A2(n10092), .A3(n10091), .ZN(n10093) );
  NAND2_X1 U12740 ( .A1(n10096), .A2(n10095), .ZN(n10111) );
  NAND2_X1 U12741 ( .A1(n10111), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n10098) );
  XNOR2_X1 U12742 ( .A(n10098), .B(n10097), .ZN(n11021) );
  OR2_X1 U12743 ( .A1(n11021), .A2(P2_U3088), .ZN(n12167) );
  INV_X1 U12744 ( .A(n12167), .ZN(n10116) );
  OAI21_X1 U12745 ( .B1(n10140), .B2(n11964), .A(n10116), .ZN(n10099) );
  INV_X1 U12746 ( .A(n10099), .ZN(n10101) );
  NAND2_X1 U12747 ( .A1(n10193), .A2(n11354), .ZN(n10100) );
  INV_X1 U12748 ( .A(n10102), .ZN(n10103) );
  INV_X1 U12749 ( .A(n13769), .ZN(n13741) );
  NAND2_X1 U12750 ( .A1(n10104), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n10105) );
  MUX2_X1 U12751 ( .A(P2_IR_REG_31__SCAN_IN), .B(n10105), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n10106) );
  NAND2_X1 U12752 ( .A1(n10106), .A2(n9493), .ZN(n14466) );
  NAND2_X1 U12753 ( .A1(n7653), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n10109) );
  MUX2_X1 U12754 ( .A(n10109), .B(P2_IR_REG_31__SCAN_IN), .S(n10108), .Z(
        n10110) );
  NAND2_X1 U12755 ( .A1(n10110), .A2(n10104), .ZN(n14468) );
  OAI21_X1 U12756 ( .B1(n10111), .B2(P2_IR_REG_23__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n10112) );
  MUX2_X1 U12757 ( .A(P2_IR_REG_31__SCAN_IN), .B(n10112), .S(
        P2_IR_REG_24__SCAN_IN), .Z(n10113) );
  NAND2_X1 U12758 ( .A1(n10113), .A2(n7653), .ZN(n14475) );
  NOR3_X1 U12759 ( .A1(n14466), .A2(n14468), .A3(n14475), .ZN(n10547) );
  INV_X1 U12760 ( .A(n10547), .ZN(n11020) );
  AND2_X1 U12761 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n11020), .ZN(n10114) );
  NOR4_X1 U12762 ( .A1(n13741), .A2(n14462), .A3(n15884), .A4(n11014), .ZN(
        n10115) );
  AOI211_X1 U12763 ( .C1(n10116), .C2(n12056), .A(n10264), .B(n10115), .ZN(
        n10117) );
  NAND2_X1 U12764 ( .A1(n13972), .A2(n13614), .ZN(n10118) );
  INV_X1 U12765 ( .A(n13797), .ZN(n10119) );
  INV_X1 U12766 ( .A(n13798), .ZN(n13576) );
  OR2_X1 U12767 ( .A1(n14362), .A2(n13576), .ZN(n10226) );
  INV_X1 U12768 ( .A(n13800), .ZN(n10120) );
  NAND2_X1 U12769 ( .A1(n14443), .A2(n10120), .ZN(n14187) );
  OR2_X1 U12770 ( .A1(n14443), .A2(n10120), .ZN(n10121) );
  AND2_X1 U12771 ( .A1(n14197), .A2(n13799), .ZN(n10165) );
  INV_X1 U12772 ( .A(n10122), .ZN(n10123) );
  NOR2_X1 U12773 ( .A1(n13812), .A2(n10196), .ZN(n11137) );
  OR2_X1 U12774 ( .A1(n10123), .A2(n11137), .ZN(n11352) );
  NOR2_X1 U12775 ( .A1(n11352), .A2(n11964), .ZN(n10124) );
  XNOR2_X1 U12776 ( .A(n13809), .B(n9522), .ZN(n11251) );
  XNOR2_X1 U12777 ( .A(n13808), .B(n15890), .ZN(n11557) );
  NAND4_X1 U12778 ( .A1(n10124), .A2(n11138), .A3(n11251), .A4(n11557), .ZN(
        n10125) );
  XNOR2_X1 U12779 ( .A(n13806), .B(n10197), .ZN(n11923) );
  NOR4_X1 U12780 ( .A1(n10125), .A2(n11463), .A3(n12000), .A4(n11923), .ZN(
        n10126) );
  XNOR2_X1 U12781 ( .A(n14386), .B(n10220), .ZN(n14240) );
  INV_X1 U12782 ( .A(n14240), .ZN(n14243) );
  AND4_X1 U12783 ( .A1(n14188), .A2(n10126), .A3(n14243), .A4(n14271), .ZN(
        n10127) );
  XNOR2_X1 U12784 ( .A(n14379), .B(n13731), .ZN(n14218) );
  INV_X1 U12785 ( .A(n14218), .ZN(n14224) );
  NAND4_X1 U12786 ( .A1(n12358), .A2(n14204), .A3(n10127), .A4(n14224), .ZN(
        n10128) );
  NAND2_X1 U12787 ( .A1(n14405), .A2(n13784), .ZN(n10188) );
  NAND2_X1 U12788 ( .A1(n14320), .A2(n13790), .ZN(n10178) );
  OR2_X1 U12789 ( .A1(n14320), .A2(n13790), .ZN(n10130) );
  NAND2_X1 U12790 ( .A1(n10178), .A2(n10130), .ZN(n14066) );
  OR2_X1 U12791 ( .A1(n14097), .A2(n13792), .ZN(n10177) );
  NAND2_X1 U12792 ( .A1(n14097), .A2(n13792), .ZN(n10176) );
  NAND2_X1 U12793 ( .A1(n10177), .A2(n10176), .ZN(n14094) );
  XNOR2_X1 U12794 ( .A(n14148), .B(n13795), .ZN(n14145) );
  XNOR2_X1 U12795 ( .A(n12026), .B(n13804), .ZN(n12020) );
  INV_X1 U12796 ( .A(n10173), .ZN(n10131) );
  AND2_X1 U12797 ( .A1(n14341), .A2(n13794), .ZN(n10174) );
  AND4_X1 U12798 ( .A1(n14094), .A2(n14145), .A3(n12020), .A4(n14124), .ZN(
        n10132) );
  INV_X1 U12799 ( .A(n14110), .ZN(n14105) );
  XNOR2_X1 U12800 ( .A(n14325), .B(n13791), .ZN(n14080) );
  AND4_X1 U12801 ( .A1(n14066), .A2(n10132), .A3(n14105), .A4(n14080), .ZN(
        n10133) );
  XNOR2_X1 U12802 ( .A(n14417), .B(n13789), .ZN(n14056) );
  XNOR2_X1 U12803 ( .A(n14039), .B(n13788), .ZN(n14034) );
  NAND4_X1 U12804 ( .A1(n10133), .A2(n13993), .A3(n14056), .A4(n14034), .ZN(
        n10134) );
  INV_X1 U12805 ( .A(n13782), .ZN(n10136) );
  AND2_X1 U12806 ( .A1(n11354), .A2(n11964), .ZN(n10195) );
  NOR4_X1 U12807 ( .A1(n10138), .A2(n10140), .A3(n10195), .A4(n12167), .ZN(
        n10139) );
  INV_X1 U12808 ( .A(n11964), .ZN(n11010) );
  NAND2_X1 U12809 ( .A1(n10140), .A2(n11010), .ZN(n10251) );
  OAI21_X1 U12810 ( .B1(n12056), .B2(n11010), .A(n10251), .ZN(n10141) );
  AOI21_X1 U12811 ( .B1(n10142), .B2(n12052), .A(n10141), .ZN(n10144) );
  INV_X1 U12812 ( .A(n10147), .ZN(n10146) );
  NAND2_X1 U12813 ( .A1(n13809), .A2(n9522), .ZN(n10145) );
  AND2_X1 U12814 ( .A1(n10146), .A2(n10145), .ZN(n11465) );
  NAND2_X1 U12815 ( .A1(n13812), .A2(n11360), .ZN(n11121) );
  NAND2_X1 U12816 ( .A1(n10148), .A2(n11121), .ZN(n11134) );
  OR2_X1 U12817 ( .A1(n13810), .A2(n7675), .ZN(n10149) );
  NAND2_X1 U12818 ( .A1(n11134), .A2(n10149), .ZN(n11464) );
  INV_X1 U12819 ( .A(n13807), .ZN(n11711) );
  NAND2_X1 U12820 ( .A1(n11711), .A2(n11506), .ZN(n10150) );
  AOI22_X1 U12821 ( .A1(n12009), .A2(n13805), .B1(n13806), .B2(n11930), .ZN(
        n10151) );
  NAND2_X1 U12822 ( .A1(n11922), .A2(n10151), .ZN(n10156) );
  INV_X1 U12823 ( .A(n13806), .ZN(n10152) );
  NAND2_X1 U12824 ( .A1(n10152), .A2(n10197), .ZN(n11996) );
  NAND2_X1 U12825 ( .A1(n11996), .A2(n13805), .ZN(n10154) );
  NOR2_X1 U12826 ( .A1(n13806), .A2(n13805), .ZN(n10153) );
  AOI22_X1 U12827 ( .A1(n10154), .A2(n15901), .B1(n10153), .B2(n10197), .ZN(
        n10155) );
  NAND2_X1 U12828 ( .A1(n10156), .A2(n10155), .ZN(n12019) );
  NAND2_X1 U12829 ( .A1(n12026), .A2(n13804), .ZN(n10157) );
  NAND2_X1 U12830 ( .A1(n12019), .A2(n10157), .ZN(n10159) );
  OR2_X1 U12831 ( .A1(n12026), .A2(n13804), .ZN(n10158) );
  NAND2_X1 U12832 ( .A1(n14264), .A2(n13803), .ZN(n10161) );
  NAND2_X1 U12833 ( .A1(n14386), .A2(n13802), .ZN(n10162) );
  NAND2_X1 U12834 ( .A1(n14379), .A2(n13801), .ZN(n10163) );
  OR2_X1 U12835 ( .A1(n14443), .A2(n13800), .ZN(n10164) );
  NOR2_X1 U12836 ( .A1(n14362), .A2(n13798), .ZN(n10167) );
  NAND2_X1 U12837 ( .A1(n14362), .A2(n13798), .ZN(n10166) );
  AND2_X1 U12838 ( .A1(n14435), .A2(n13797), .ZN(n10168) );
  OAI22_X1 U12839 ( .A1(n14181), .A2(n10168), .B1(n14435), .B2(n13797), .ZN(
        n14156) );
  OR2_X1 U12840 ( .A1(n14351), .A2(n13796), .ZN(n10169) );
  NAND2_X1 U12841 ( .A1(n14148), .A2(n13795), .ZN(n10172) );
  INV_X1 U12842 ( .A(n12686), .ZN(n13793) );
  OR2_X1 U12843 ( .A1(n14335), .A2(n13793), .ZN(n10175) );
  NAND2_X1 U12844 ( .A1(n14325), .A2(n13791), .ZN(n14064) );
  NAND3_X1 U12845 ( .A1(n14063), .A2(n10178), .A3(n14064), .ZN(n14047) );
  OAI21_X1 U12846 ( .B1(n14325), .B2(n13791), .A(n13790), .ZN(n10180) );
  NOR2_X1 U12847 ( .A1(n13790), .A2(n13791), .ZN(n10179) );
  AOI22_X1 U12848 ( .A1(n10202), .A2(n10180), .B1(n7668), .B2(n10179), .ZN(
        n14046) );
  INV_X1 U12849 ( .A(n14056), .ZN(n10181) );
  AND2_X1 U12850 ( .A1(n14046), .A2(n10181), .ZN(n10182) );
  NAND2_X1 U12851 ( .A1(n14417), .A2(n13789), .ZN(n10183) );
  AND2_X1 U12852 ( .A1(n14039), .A2(n13788), .ZN(n10186) );
  NAND2_X1 U12853 ( .A1(n7352), .A2(n13786), .ZN(n13991) );
  AND2_X1 U12854 ( .A1(n7420), .A2(n13991), .ZN(n10187) );
  NAND2_X1 U12855 ( .A1(n10191), .A2(n11002), .ZN(n10192) );
  NAND2_X1 U12856 ( .A1(n10193), .A2(n10192), .ZN(n10194) );
  NAND2_X1 U12857 ( .A1(n10195), .A2(n12056), .ZN(n14303) );
  NAND2_X1 U12858 ( .A1(n11003), .A2(n14303), .ZN(n14396) );
  NAND2_X1 U12859 ( .A1(n11296), .A2(n10196), .ZN(n11252) );
  INV_X1 U12860 ( .A(n12026), .ZN(n12071) );
  INV_X1 U12861 ( .A(n14264), .ZN(n14393) );
  INV_X1 U12862 ( .A(n14443), .ZN(n14207) );
  AOI211_X1 U12863 ( .C1(n13972), .C2(n6538), .A(n15891), .B(n12385), .ZN(
        n13971) );
  NAND2_X1 U12864 ( .A1(n11138), .A2(n11137), .ZN(n10205) );
  OR2_X1 U12865 ( .A1(n13810), .A2(n11296), .ZN(n10204) );
  NAND2_X1 U12866 ( .A1(n10205), .A2(n10204), .ZN(n11255) );
  NAND2_X1 U12867 ( .A1(n11255), .A2(n11251), .ZN(n10207) );
  INV_X1 U12868 ( .A(n9522), .ZN(n11684) );
  OR2_X1 U12869 ( .A1(n13809), .A2(n11684), .ZN(n10206) );
  NAND2_X1 U12870 ( .A1(n10207), .A2(n10206), .ZN(n11558) );
  NAND2_X1 U12871 ( .A1(n11558), .A2(n11557), .ZN(n10209) );
  NAND2_X1 U12872 ( .A1(n7805), .A2(n15890), .ZN(n10208) );
  INV_X1 U12873 ( .A(n11463), .ZN(n11469) );
  NAND2_X1 U12874 ( .A1(n11711), .A2(n10210), .ZN(n10211) );
  NOR2_X1 U12875 ( .A1(n13806), .A2(n10197), .ZN(n10213) );
  NAND2_X1 U12876 ( .A1(n13806), .A2(n10197), .ZN(n10212) );
  INV_X1 U12877 ( .A(n13805), .ZN(n11899) );
  NAND2_X1 U12878 ( .A1(n11899), .A2(n12009), .ZN(n10214) );
  INV_X1 U12879 ( .A(n13804), .ZN(n10216) );
  OR2_X1 U12880 ( .A1(n10216), .A2(n12026), .ZN(n10215) );
  NAND2_X1 U12881 ( .A1(n12021), .A2(n10215), .ZN(n10218) );
  NAND2_X1 U12882 ( .A1(n12026), .A2(n10216), .ZN(n10217) );
  NAND2_X1 U12883 ( .A1(n14379), .A2(n13731), .ZN(n10219) );
  NAND2_X1 U12884 ( .A1(n14386), .A2(n10220), .ZN(n14223) );
  OR2_X1 U12885 ( .A1(n14264), .A2(n7482), .ZN(n14222) );
  OAI21_X1 U12886 ( .B1(n14386), .B2(n10220), .A(n14222), .ZN(n10222) );
  INV_X1 U12887 ( .A(n14379), .ZN(n10221) );
  INV_X1 U12888 ( .A(n13799), .ZN(n10225) );
  NAND2_X1 U12889 ( .A1(n14197), .A2(n10225), .ZN(n10224) );
  INV_X1 U12890 ( .A(n14435), .ZN(n10227) );
  INV_X1 U12891 ( .A(n13794), .ZN(n13742) );
  OR2_X1 U12892 ( .A1(n14341), .A2(n13742), .ZN(n10229) );
  INV_X1 U12893 ( .A(n13795), .ZN(n10228) );
  OR2_X1 U12894 ( .A1(n14148), .A2(n10228), .ZN(n14123) );
  AND2_X1 U12895 ( .A1(n10229), .A2(n14123), .ZN(n10231) );
  NAND2_X1 U12896 ( .A1(n14351), .A2(n13670), .ZN(n14122) );
  OAI21_X1 U12897 ( .B1(n14431), .B2(n13795), .A(n14122), .ZN(n10232) );
  AOI22_X1 U12898 ( .A1(n10232), .A2(n10231), .B1(n13742), .B2(n14341), .ZN(
        n10233) );
  AND2_X1 U12899 ( .A1(n14335), .A2(n12686), .ZN(n10235) );
  OR2_X1 U12900 ( .A1(n14335), .A2(n12686), .ZN(n10234) );
  INV_X1 U12901 ( .A(n13792), .ZN(n13744) );
  NOR2_X1 U12902 ( .A1(n14097), .A2(n13744), .ZN(n10237) );
  NAND2_X1 U12903 ( .A1(n14097), .A2(n13744), .ZN(n10236) );
  INV_X1 U12904 ( .A(n13791), .ZN(n10238) );
  AND2_X1 U12905 ( .A1(n14325), .A2(n10238), .ZN(n10239) );
  INV_X1 U12906 ( .A(n13790), .ZN(n10240) );
  NAND2_X1 U12907 ( .A1(n14320), .A2(n10240), .ZN(n10241) );
  INV_X1 U12908 ( .A(n13789), .ZN(n10242) );
  NAND2_X1 U12909 ( .A1(n14417), .A2(n10242), .ZN(n10243) );
  INV_X1 U12910 ( .A(n13788), .ZN(n10244) );
  NAND2_X1 U12911 ( .A1(n14039), .A2(n10244), .ZN(n10245) );
  INV_X1 U12912 ( .A(n13787), .ZN(n13649) );
  NAND2_X1 U12913 ( .A1(n14299), .A2(n13649), .ZN(n10246) );
  INV_X1 U12914 ( .A(n13786), .ZN(n13752) );
  INV_X1 U12915 ( .A(n13785), .ZN(n10247) );
  NAND2_X1 U12916 ( .A1(n13995), .A2(n10247), .ZN(n10248) );
  INV_X1 U12917 ( .A(n13784), .ZN(n10249) );
  AND2_X1 U12918 ( .A1(n14405), .A2(n10249), .ZN(n10250) );
  OAI21_X1 U12919 ( .B1(n10253), .B2(n10190), .A(n14270), .ZN(n10254) );
  AOI22_X1 U12920 ( .A1(n13782), .A2(n13770), .B1(n13784), .B2(n13769), .ZN(
        n13622) );
  NOR4_X1 U12921 ( .A1(P2_D_REG_12__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .A3(
        P2_D_REG_4__SCAN_IN), .A4(P2_D_REG_5__SCAN_IN), .ZN(n10263) );
  INV_X1 U12922 ( .A(P2_D_REG_20__SCAN_IN), .ZN(n15874) );
  NAND4_X1 U12923 ( .A1(n15876), .A2(n15873), .A3(n15874), .A4(n15878), .ZN(
        n10260) );
  NOR4_X1 U12924 ( .A1(P2_D_REG_16__SCAN_IN), .A2(P2_D_REG_17__SCAN_IN), .A3(
        P2_D_REG_18__SCAN_IN), .A4(P2_D_REG_19__SCAN_IN), .ZN(n10258) );
  NOR4_X1 U12925 ( .A1(P2_D_REG_14__SCAN_IN), .A2(P2_D_REG_11__SCAN_IN), .A3(
        P2_D_REG_13__SCAN_IN), .A4(P2_D_REG_15__SCAN_IN), .ZN(n10257) );
  NOR4_X1 U12926 ( .A1(P2_D_REG_26__SCAN_IN), .A2(P2_D_REG_27__SCAN_IN), .A3(
        P2_D_REG_28__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n10256) );
  NOR4_X1 U12927 ( .A1(P2_D_REG_21__SCAN_IN), .A2(P2_D_REG_23__SCAN_IN), .A3(
        P2_D_REG_24__SCAN_IN), .A4(P2_D_REG_25__SCAN_IN), .ZN(n10255) );
  NAND4_X1 U12928 ( .A1(n10258), .A2(n10257), .A3(n10256), .A4(n10255), .ZN(
        n10259) );
  NOR4_X1 U12929 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        n10260), .A4(n10259), .ZN(n10262) );
  NOR4_X1 U12930 ( .A1(P2_D_REG_6__SCAN_IN), .A2(P2_D_REG_7__SCAN_IN), .A3(
        P2_D_REG_9__SCAN_IN), .A4(P2_D_REG_10__SCAN_IN), .ZN(n10261) );
  NAND3_X1 U12931 ( .A1(n10263), .A2(n10262), .A3(n10261), .ZN(n10267) );
  XOR2_X1 U12932 ( .A(n14475), .B(n10264), .Z(n10265) );
  NOR2_X1 U12933 ( .A1(n10268), .A2(n12056), .ZN(n11023) );
  NOR2_X1 U12934 ( .A1(n11006), .A2(n11023), .ZN(n11324) );
  INV_X1 U12935 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n15885) );
  NAND2_X1 U12936 ( .A1(n15872), .A2(n15885), .ZN(n10270) );
  NAND2_X1 U12937 ( .A1(n14466), .A2(n14468), .ZN(n10269) );
  NAND2_X1 U12938 ( .A1(n10270), .A2(n10269), .ZN(n11321) );
  AND2_X1 U12939 ( .A1(n11321), .A2(n15882), .ZN(n15883) );
  NAND2_X1 U12940 ( .A1(n14261), .A2(n11354), .ZN(n11018) );
  AND2_X1 U12941 ( .A1(n15883), .A2(n11018), .ZN(n10271) );
  NAND2_X1 U12942 ( .A1(n15872), .A2(n15880), .ZN(n10273) );
  NAND2_X1 U12943 ( .A1(n14475), .A2(n14466), .ZN(n10272) );
  NAND2_X1 U12944 ( .A1(n15908), .A2(n14387), .ZN(n14430) );
  INV_X1 U12945 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n10274) );
  NOR2_X1 U12946 ( .A1(n15908), .A2(n10274), .ZN(n10275) );
  NAND2_X1 U12947 ( .A1(n10278), .A2(n10277), .ZN(P2_U3495) );
  INV_X1 U12948 ( .A(n10290), .ZN(n10279) );
  OAI22_X1 U12949 ( .A1(n15187), .A2(n10295), .B1(n14812), .B2(n10303), .ZN(
        n10477) );
  OAI22_X1 U12950 ( .A1(n15187), .A2(n10290), .B1(n14812), .B2(n10295), .ZN(
        n10280) );
  XNOR2_X1 U12951 ( .A(n10280), .B(n14529), .ZN(n10476) );
  OAI22_X1 U12952 ( .A1(n15214), .A2(n10295), .B1(n15402), .B2(n10303), .ZN(
        n10468) );
  OAI22_X1 U12953 ( .A1(n15214), .A2(n10290), .B1(n15402), .B2(n10295), .ZN(
        n10281) );
  XNOR2_X1 U12954 ( .A(n10281), .B(n14529), .ZN(n10467) );
  OAI22_X1 U12955 ( .A1(n10295), .A2(n11371), .B1(n15717), .B2(n10549), .ZN(
        n10282) );
  AOI21_X1 U12956 ( .B1(n10283), .B2(n10296), .A(n10282), .ZN(n10859) );
  NAND2_X1 U12957 ( .A1(n10283), .A2(n10469), .ZN(n10286) );
  INV_X1 U12958 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n10743) );
  OAI22_X1 U12959 ( .A1(n10290), .A2(n11371), .B1(n10743), .B2(n10549), .ZN(
        n10284) );
  INV_X1 U12960 ( .A(n10284), .ZN(n10285) );
  NAND2_X1 U12961 ( .A1(n10286), .A2(n10285), .ZN(n10858) );
  NAND2_X1 U12962 ( .A1(n10859), .A2(n10858), .ZN(n10857) );
  NAND2_X1 U12963 ( .A1(n10857), .A2(n10288), .ZN(n11163) );
  NAND2_X1 U12964 ( .A1(n10855), .A2(n10469), .ZN(n10292) );
  OR2_X1 U12965 ( .A1(n10290), .A2(n15783), .ZN(n10291) );
  NAND2_X1 U12966 ( .A1(n10292), .A2(n10291), .ZN(n10293) );
  INV_X1 U12967 ( .A(n10294), .ZN(n10855) );
  AOI22_X1 U12968 ( .A1(n10855), .A2(n10296), .B1(n11166), .B2(n14525), .ZN(
        n10298) );
  XNOR2_X1 U12969 ( .A(n10297), .B(n10298), .ZN(n11162) );
  NAND2_X1 U12970 ( .A1(n11163), .A2(n11162), .ZN(n10301) );
  INV_X1 U12971 ( .A(n10297), .ZN(n10299) );
  NAND2_X1 U12972 ( .A1(n10299), .A2(n10298), .ZN(n10300) );
  NAND2_X1 U12973 ( .A1(n10301), .A2(n10300), .ZN(n11314) );
  OAI22_X1 U12974 ( .A1(n14709), .A2(n10295), .B1(n14699), .B2(n10290), .ZN(
        n10302) );
  XNOR2_X1 U12975 ( .A(n10302), .B(n10287), .ZN(n10306) );
  OAI22_X1 U12976 ( .A1(n14709), .A2(n10303), .B1(n14699), .B2(n10295), .ZN(
        n10304) );
  XNOR2_X1 U12977 ( .A(n10306), .B(n10304), .ZN(n11315) );
  NAND2_X1 U12978 ( .A1(n11314), .A2(n11315), .ZN(n10308) );
  INV_X1 U12979 ( .A(n10304), .ZN(n10305) );
  NAND2_X1 U12980 ( .A1(n10306), .A2(n10305), .ZN(n10307) );
  NAND2_X1 U12981 ( .A1(n14531), .A2(n6534), .ZN(n10311) );
  NAND2_X1 U12982 ( .A1(n10309), .A2(n14525), .ZN(n10310) );
  NAND2_X1 U12983 ( .A1(n10311), .A2(n10310), .ZN(n10312) );
  XNOR2_X1 U12984 ( .A(n10312), .B(n10287), .ZN(n10314) );
  AND2_X1 U12985 ( .A1(n6534), .A2(n10469), .ZN(n10313) );
  INV_X1 U12986 ( .A(n10314), .ZN(n10317) );
  INV_X1 U12987 ( .A(n10315), .ZN(n10316) );
  NAND2_X1 U12988 ( .A1(n10317), .A2(n10316), .ZN(n10318) );
  NAND2_X1 U12989 ( .A1(n14970), .A2(n14526), .ZN(n10320) );
  OR2_X1 U12990 ( .A1(n11283), .A2(n10295), .ZN(n10319) );
  NAND2_X1 U12991 ( .A1(n14970), .A2(n14525), .ZN(n10322) );
  OR2_X1 U12992 ( .A1(n11283), .A2(n10290), .ZN(n10321) );
  NAND2_X1 U12993 ( .A1(n10322), .A2(n10321), .ZN(n10323) );
  XNOR2_X1 U12994 ( .A(n10323), .B(n10287), .ZN(n11548) );
  OAI22_X1 U12995 ( .A1(n11849), .A2(n10295), .B1(n11885), .B2(n10290), .ZN(
        n10324) );
  XNOR2_X1 U12996 ( .A(n10324), .B(n14529), .ZN(n10325) );
  OAI22_X1 U12997 ( .A1(n11849), .A2(n10303), .B1(n11885), .B2(n10295), .ZN(
        n10326) );
  NAND2_X1 U12998 ( .A1(n10325), .A2(n10326), .ZN(n11620) );
  NAND2_X1 U12999 ( .A1(n11623), .A2(n11620), .ZN(n10329) );
  INV_X1 U13000 ( .A(n10325), .ZN(n10328) );
  INV_X1 U13001 ( .A(n10326), .ZN(n10327) );
  NAND2_X1 U13002 ( .A1(n10328), .A2(n10327), .ZN(n11621) );
  OR2_X1 U13003 ( .A1(n7943), .A2(n10295), .ZN(n10331) );
  NAND2_X1 U13004 ( .A1(n14968), .A2(n14526), .ZN(n10330) );
  AND2_X1 U13005 ( .A1(n10331), .A2(n10330), .ZN(n10335) );
  NAND2_X1 U13006 ( .A1(n11842), .A2(n10335), .ZN(n10334) );
  NAND2_X1 U13007 ( .A1(n14968), .A2(n14525), .ZN(n10332) );
  OAI21_X1 U13008 ( .B1(n7943), .B2(n10290), .A(n10332), .ZN(n10333) );
  XNOR2_X1 U13009 ( .A(n10333), .B(n14529), .ZN(n11840) );
  NAND2_X1 U13010 ( .A1(n10334), .A2(n11840), .ZN(n10338) );
  INV_X1 U13011 ( .A(n11842), .ZN(n10336) );
  INV_X1 U13012 ( .A(n10335), .ZN(n11839) );
  NAND2_X1 U13013 ( .A1(n10336), .A2(n11839), .ZN(n10337) );
  NAND2_X1 U13014 ( .A1(n14733), .A2(n14531), .ZN(n10340) );
  NAND2_X1 U13015 ( .A1(n15799), .A2(n10469), .ZN(n10339) );
  NAND2_X1 U13016 ( .A1(n10340), .A2(n10339), .ZN(n10341) );
  XNOR2_X1 U13017 ( .A(n10341), .B(n14529), .ZN(n10342) );
  AOI22_X1 U13018 ( .A1(n14733), .A2(n10469), .B1(n15799), .B2(n14526), .ZN(
        n10343) );
  XNOR2_X1 U13019 ( .A(n10342), .B(n10343), .ZN(n14477) );
  INV_X1 U13020 ( .A(n10342), .ZN(n10344) );
  OR2_X1 U13021 ( .A1(n10344), .A2(n10343), .ZN(n10345) );
  NAND2_X1 U13022 ( .A1(n14737), .A2(n14531), .ZN(n10347) );
  NAND2_X1 U13023 ( .A1(n14967), .A2(n14525), .ZN(n10346) );
  NAND2_X1 U13024 ( .A1(n10347), .A2(n10346), .ZN(n10348) );
  XNOR2_X1 U13025 ( .A(n10348), .B(n10287), .ZN(n10350) );
  NOR2_X1 U13026 ( .A1(n14618), .A2(n10303), .ZN(n10349) );
  AOI21_X1 U13027 ( .B1(n14737), .B2(n14525), .A(n10349), .ZN(n10351) );
  NAND2_X1 U13028 ( .A1(n10350), .A2(n10351), .ZN(n10355) );
  INV_X1 U13029 ( .A(n10350), .ZN(n10353) );
  INV_X1 U13030 ( .A(n10351), .ZN(n10352) );
  NAND2_X1 U13031 ( .A1(n10353), .A2(n10352), .ZN(n10354) );
  NAND2_X1 U13032 ( .A1(n10355), .A2(n10354), .ZN(n14548) );
  NAND2_X1 U13033 ( .A1(n15495), .A2(n14531), .ZN(n10357) );
  NAND2_X1 U13034 ( .A1(n14966), .A2(n14525), .ZN(n10356) );
  NAND2_X1 U13035 ( .A1(n10357), .A2(n10356), .ZN(n10358) );
  XNOR2_X1 U13036 ( .A(n10358), .B(n10287), .ZN(n10367) );
  NOR2_X1 U13037 ( .A1(n12249), .A2(n10303), .ZN(n10359) );
  AOI21_X1 U13038 ( .B1(n15495), .B2(n14525), .A(n10359), .ZN(n10368) );
  NAND2_X1 U13039 ( .A1(n10367), .A2(n10368), .ZN(n14508) );
  NAND2_X1 U13040 ( .A1(n14742), .A2(n14531), .ZN(n10361) );
  NAND2_X1 U13041 ( .A1(n15800), .A2(n10469), .ZN(n10360) );
  NAND2_X1 U13042 ( .A1(n10361), .A2(n10360), .ZN(n10362) );
  XNOR2_X1 U13043 ( .A(n10362), .B(n10287), .ZN(n14615) );
  NOR2_X1 U13044 ( .A1(n14513), .A2(n10303), .ZN(n10363) );
  AOI21_X1 U13045 ( .B1(n14742), .B2(n14525), .A(n10363), .ZN(n10365) );
  NAND2_X1 U13046 ( .A1(n14615), .A2(n10365), .ZN(n10364) );
  NAND2_X1 U13047 ( .A1(n14508), .A2(n10364), .ZN(n10377) );
  INV_X1 U13048 ( .A(n10377), .ZN(n14648) );
  INV_X1 U13049 ( .A(n14615), .ZN(n10366) );
  INV_X1 U13050 ( .A(n10365), .ZN(n14504) );
  AND2_X1 U13051 ( .A1(n10366), .A2(n14504), .ZN(n14649) );
  INV_X1 U13052 ( .A(n10367), .ZN(n10370) );
  INV_X1 U13053 ( .A(n10368), .ZN(n10369) );
  AND2_X1 U13054 ( .A1(n10370), .A2(n10369), .ZN(n14507) );
  AOI21_X1 U13055 ( .B1(n14648), .B2(n14649), .A(n14507), .ZN(n10375) );
  NAND2_X1 U13056 ( .A1(n15490), .A2(n14531), .ZN(n10372) );
  NAND2_X1 U13057 ( .A1(n15478), .A2(n14525), .ZN(n10371) );
  NAND2_X1 U13058 ( .A1(n10372), .A2(n10371), .ZN(n10373) );
  XNOR2_X1 U13059 ( .A(n10373), .B(n14529), .ZN(n10378) );
  AND2_X1 U13060 ( .A1(n15478), .A2(n14526), .ZN(n10374) );
  AOI21_X1 U13061 ( .B1(n15490), .B2(n14525), .A(n10374), .ZN(n10379) );
  XNOR2_X1 U13062 ( .A(n10378), .B(n10379), .ZN(n14651) );
  INV_X1 U13063 ( .A(n10378), .ZN(n10380) );
  NAND2_X1 U13064 ( .A1(n10380), .A2(n10379), .ZN(n10381) );
  NAND2_X1 U13065 ( .A1(n15480), .A2(n14531), .ZN(n10383) );
  NAND2_X1 U13066 ( .A1(n14965), .A2(n14525), .ZN(n10382) );
  NAND2_X1 U13067 ( .A1(n10383), .A2(n10382), .ZN(n10384) );
  XNOR2_X1 U13068 ( .A(n10384), .B(n14529), .ZN(n10386) );
  NOR2_X1 U13069 ( .A1(n15466), .A2(n10303), .ZN(n10385) );
  AOI21_X1 U13070 ( .B1(n15480), .B2(n14525), .A(n10385), .ZN(n10387) );
  XNOR2_X1 U13071 ( .A(n10386), .B(n10387), .ZN(n14570) );
  INV_X1 U13072 ( .A(n10386), .ZN(n10388) );
  NAND2_X1 U13073 ( .A1(n10388), .A2(n10387), .ZN(n10389) );
  NAND2_X1 U13074 ( .A1(n15471), .A2(n14531), .ZN(n10391) );
  NAND2_X1 U13075 ( .A1(n15479), .A2(n14525), .ZN(n10390) );
  NAND2_X1 U13076 ( .A1(n10391), .A2(n10390), .ZN(n10392) );
  XNOR2_X1 U13077 ( .A(n10392), .B(n14529), .ZN(n10394) );
  NOR2_X1 U13078 ( .A1(n14572), .A2(n10303), .ZN(n10393) );
  AOI21_X1 U13079 ( .B1(n15471), .B2(n14525), .A(n10393), .ZN(n10395) );
  XNOR2_X1 U13080 ( .A(n10394), .B(n10395), .ZN(n14631) );
  INV_X1 U13081 ( .A(n10394), .ZN(n10396) );
  NAND2_X1 U13082 ( .A1(n10396), .A2(n10395), .ZN(n10397) );
  NAND2_X1 U13083 ( .A1(n14772), .A2(n14531), .ZN(n10399) );
  NAND2_X1 U13084 ( .A1(n15449), .A2(n14525), .ZN(n10398) );
  NAND2_X1 U13085 ( .A1(n10399), .A2(n10398), .ZN(n10400) );
  XNOR2_X1 U13086 ( .A(n10400), .B(n14529), .ZN(n10402) );
  NOR2_X1 U13087 ( .A1(n15468), .A2(n10303), .ZN(n10401) );
  AOI21_X1 U13088 ( .B1(n14772), .B2(n14525), .A(n10401), .ZN(n10403) );
  XNOR2_X1 U13089 ( .A(n10402), .B(n10403), .ZN(n14487) );
  INV_X1 U13090 ( .A(n10402), .ZN(n10404) );
  NAND2_X1 U13091 ( .A1(n10404), .A2(n10403), .ZN(n10405) );
  NAND2_X1 U13092 ( .A1(n15325), .A2(n14531), .ZN(n10407) );
  NAND2_X1 U13093 ( .A1(n15458), .A2(n14525), .ZN(n10406) );
  NAND2_X1 U13094 ( .A1(n10407), .A2(n10406), .ZN(n10408) );
  XNOR2_X1 U13095 ( .A(n10408), .B(n14529), .ZN(n10417) );
  NAND2_X1 U13096 ( .A1(n15325), .A2(n14525), .ZN(n10410) );
  NAND2_X1 U13097 ( .A1(n15458), .A2(n14526), .ZN(n10409) );
  NAND2_X1 U13098 ( .A1(n10410), .A2(n10409), .ZN(n14678) );
  NAND2_X1 U13099 ( .A1(n15444), .A2(n14531), .ZN(n10412) );
  OR2_X1 U13100 ( .A1(n15434), .A2(n10295), .ZN(n10411) );
  NAND2_X1 U13101 ( .A1(n10412), .A2(n10411), .ZN(n10413) );
  XNOR2_X1 U13102 ( .A(n10413), .B(n14529), .ZN(n14588) );
  NAND2_X1 U13103 ( .A1(n15444), .A2(n14525), .ZN(n10415) );
  OR2_X1 U13104 ( .A1(n15434), .A2(n10303), .ZN(n10414) );
  NAND2_X1 U13105 ( .A1(n10415), .A2(n10414), .ZN(n10421) );
  AND2_X1 U13106 ( .A1(n14588), .A2(n10421), .ZN(n10418) );
  AOI21_X1 U13107 ( .B1(n10417), .B2(n14678), .A(n10418), .ZN(n10416) );
  NAND2_X1 U13108 ( .A1(n14585), .A2(n10416), .ZN(n10425) );
  INV_X1 U13109 ( .A(n10417), .ZN(n14586) );
  INV_X1 U13110 ( .A(n10418), .ZN(n10420) );
  INV_X1 U13111 ( .A(n14678), .ZN(n10419) );
  AND2_X1 U13112 ( .A1(n10420), .A2(n10419), .ZN(n10423) );
  INV_X1 U13113 ( .A(n10421), .ZN(n14587) );
  INV_X1 U13114 ( .A(n14588), .ZN(n10422) );
  AOI22_X1 U13115 ( .A1(n14586), .A2(n10423), .B1(n14587), .B2(n10422), .ZN(
        n10424) );
  NAND2_X1 U13116 ( .A1(n10425), .A2(n10424), .ZN(n14596) );
  NAND2_X1 U13117 ( .A1(n15438), .A2(n14531), .ZN(n10427) );
  NAND2_X1 U13118 ( .A1(n15274), .A2(n14525), .ZN(n10426) );
  NAND2_X1 U13119 ( .A1(n10427), .A2(n10426), .ZN(n10428) );
  XNOR2_X1 U13120 ( .A(n10428), .B(n14529), .ZN(n10430) );
  NOR2_X1 U13121 ( .A1(n15311), .A2(n10303), .ZN(n10429) );
  AOI21_X1 U13122 ( .B1(n15438), .B2(n14525), .A(n10429), .ZN(n10431) );
  XNOR2_X1 U13123 ( .A(n10430), .B(n10431), .ZN(n14597) );
  NAND2_X1 U13124 ( .A1(n14596), .A2(n14597), .ZN(n10434) );
  INV_X1 U13125 ( .A(n10430), .ZN(n10432) );
  NAND2_X1 U13126 ( .A1(n10432), .A2(n10431), .ZN(n10433) );
  NAND2_X1 U13127 ( .A1(n15284), .A2(n14531), .ZN(n10436) );
  NAND2_X1 U13128 ( .A1(n15418), .A2(n14525), .ZN(n10435) );
  NAND2_X1 U13129 ( .A1(n10436), .A2(n10435), .ZN(n10437) );
  XNOR2_X1 U13130 ( .A(n10437), .B(n14529), .ZN(n10439) );
  NOR2_X1 U13131 ( .A1(n15435), .A2(n10303), .ZN(n10438) );
  AOI21_X1 U13132 ( .B1(n15284), .B2(n14525), .A(n10438), .ZN(n10440) );
  XNOR2_X1 U13133 ( .A(n10439), .B(n10440), .ZN(n14663) );
  INV_X1 U13134 ( .A(n10439), .ZN(n10441) );
  NAND2_X1 U13135 ( .A1(n10441), .A2(n10440), .ZN(n10442) );
  NAND2_X1 U13136 ( .A1(n15252), .A2(n14531), .ZN(n10444) );
  NAND2_X1 U13137 ( .A1(n15428), .A2(n14525), .ZN(n10443) );
  NAND2_X1 U13138 ( .A1(n10444), .A2(n10443), .ZN(n10445) );
  XNOR2_X1 U13139 ( .A(n10445), .B(n10287), .ZN(n10457) );
  NOR2_X1 U13140 ( .A1(n15409), .A2(n10303), .ZN(n10446) );
  AOI21_X1 U13141 ( .B1(n7226), .B2(n14525), .A(n10446), .ZN(n10458) );
  XNOR2_X1 U13142 ( .A(n10457), .B(n10458), .ZN(n14521) );
  NAND2_X1 U13143 ( .A1(n15413), .A2(n14531), .ZN(n10448) );
  NAND2_X1 U13144 ( .A1(n15419), .A2(n14525), .ZN(n10447) );
  NAND2_X1 U13145 ( .A1(n10448), .A2(n10447), .ZN(n10449) );
  XNOR2_X1 U13146 ( .A(n10449), .B(n10287), .ZN(n14559) );
  NOR2_X1 U13147 ( .A1(n15401), .A2(n10303), .ZN(n10450) );
  AOI21_X1 U13148 ( .B1(n15413), .B2(n14525), .A(n10450), .ZN(n10455) );
  NAND2_X1 U13149 ( .A1(n15405), .A2(n14531), .ZN(n10452) );
  NAND2_X1 U13150 ( .A1(n15240), .A2(n10469), .ZN(n10451) );
  NAND2_X1 U13151 ( .A1(n10452), .A2(n10451), .ZN(n10453) );
  XNOR2_X1 U13152 ( .A(n10453), .B(n14529), .ZN(n10465) );
  AND2_X1 U13153 ( .A1(n15240), .A2(n14526), .ZN(n10454) );
  AOI21_X1 U13154 ( .B1(n15405), .B2(n10469), .A(n10454), .ZN(n10463) );
  XNOR2_X1 U13155 ( .A(n10465), .B(n10463), .ZN(n14560) );
  INV_X1 U13156 ( .A(n14559), .ZN(n10456) );
  INV_X1 U13157 ( .A(n10455), .ZN(n14558) );
  NAND2_X1 U13158 ( .A1(n10456), .A2(n14558), .ZN(n14561) );
  INV_X1 U13159 ( .A(n10457), .ZN(n10460) );
  INV_X1 U13160 ( .A(n10458), .ZN(n10459) );
  AND2_X1 U13161 ( .A1(n10460), .A2(n10459), .ZN(n14555) );
  NAND2_X1 U13162 ( .A1(n8032), .A2(n14555), .ZN(n10461) );
  AND3_X1 U13163 ( .A1(n14560), .A2(n14561), .A3(n10461), .ZN(n10462) );
  INV_X1 U13164 ( .A(n10463), .ZN(n10464) );
  OR2_X1 U13165 ( .A1(n10465), .A2(n10464), .ZN(n10466) );
  XNOR2_X1 U13166 ( .A(n10467), .B(n10468), .ZN(n14644) );
  OAI22_X1 U13167 ( .A1(n15386), .A2(n10295), .B1(n15392), .B2(n10303), .ZN(
        n10473) );
  NAND2_X1 U13168 ( .A1(n15194), .A2(n14531), .ZN(n10471) );
  NAND2_X1 U13169 ( .A1(n15212), .A2(n10469), .ZN(n10470) );
  NAND2_X1 U13170 ( .A1(n10471), .A2(n10470), .ZN(n10472) );
  XNOR2_X1 U13171 ( .A(n10472), .B(n14529), .ZN(n10474) );
  XOR2_X1 U13172 ( .A(n10473), .B(n10474), .Z(n14496) );
  NAND2_X1 U13173 ( .A1(n14494), .A2(n10475), .ZN(n14603) );
  XOR2_X1 U13174 ( .A(n10477), .B(n10476), .Z(n14604) );
  OR2_X1 U13175 ( .A1(n8724), .A2(n15545), .ZN(n10478) );
  NAND2_X1 U13176 ( .A1(n15379), .A2(n14531), .ZN(n10481) );
  NAND2_X1 U13177 ( .A1(n14964), .A2(n14525), .ZN(n10480) );
  NAND2_X1 U13178 ( .A1(n10481), .A2(n10480), .ZN(n10482) );
  XNOR2_X1 U13179 ( .A(n10482), .B(n14529), .ZN(n10483) );
  AOI22_X1 U13180 ( .A1(n15379), .A2(n14525), .B1(n14526), .B2(n14964), .ZN(
        n10484) );
  XNOR2_X1 U13181 ( .A(n10483), .B(n10484), .ZN(n14580) );
  INV_X1 U13182 ( .A(n10483), .ZN(n10485) );
  NAND2_X1 U13183 ( .A1(n14464), .A2(n8743), .ZN(n10487) );
  OR2_X1 U13184 ( .A1(n8724), .A2(n15540), .ZN(n10486) );
  NAND2_X1 U13185 ( .A1(n15373), .A2(n14531), .ZN(n10497) );
  INV_X1 U13186 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n14673) );
  NAND2_X1 U13187 ( .A1(n10488), .A2(n14673), .ZN(n10489) );
  NAND2_X1 U13188 ( .A1(n10490), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n10492) );
  NAND2_X1 U13189 ( .A1(n14835), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n10491) );
  OAI211_X1 U13190 ( .C1(n14834), .C2(n9284), .A(n10492), .B(n10491), .ZN(
        n10493) );
  INV_X1 U13191 ( .A(n10493), .ZN(n10494) );
  NAND2_X1 U13192 ( .A1(n10497), .A2(n10496), .ZN(n10498) );
  XNOR2_X1 U13193 ( .A(n10498), .B(n10287), .ZN(n14671) );
  NOR2_X1 U13194 ( .A1(n14823), .A2(n10303), .ZN(n10499) );
  AOI21_X1 U13195 ( .B1(n15373), .B2(n14525), .A(n10499), .ZN(n14670) );
  NAND2_X1 U13196 ( .A1(n14671), .A2(n14670), .ZN(n10502) );
  INV_X1 U13197 ( .A(n14671), .ZN(n10501) );
  INV_X1 U13198 ( .A(n14670), .ZN(n10500) );
  NAND2_X1 U13199 ( .A1(n14460), .A2(n8743), .ZN(n10504) );
  OR2_X1 U13200 ( .A1(n8724), .A2(n15538), .ZN(n10503) );
  XNOR2_X1 U13201 ( .A(n10531), .B(P1_REG3_REG_27__SCAN_IN), .ZN(n12738) );
  NAND2_X1 U13202 ( .A1(n12738), .A2(n8980), .ZN(n10510) );
  NAND2_X1 U13203 ( .A1(n10533), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n10506) );
  NAND2_X1 U13204 ( .A1(n14835), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n10505) );
  OAI211_X1 U13205 ( .C1(n14839), .C2(n10507), .A(n10506), .B(n10505), .ZN(
        n10508) );
  INV_X1 U13206 ( .A(n10508), .ZN(n10509) );
  OAI22_X1 U13207 ( .A1(n14866), .A2(n10290), .B1(n14867), .B2(n10295), .ZN(
        n10511) );
  XNOR2_X1 U13208 ( .A(n10511), .B(n14529), .ZN(n10513) );
  OAI22_X1 U13209 ( .A1(n14866), .A2(n10295), .B1(n14867), .B2(n10303), .ZN(
        n10512) );
  NOR2_X1 U13210 ( .A1(n10513), .A2(n10512), .ZN(n14543) );
  AOI21_X1 U13211 ( .B1(n10513), .B2(n10512), .A(n14543), .ZN(n10514) );
  NAND2_X1 U13212 ( .A1(n10515), .A2(n10514), .ZN(n14541) );
  NAND2_X1 U13213 ( .A1(n14541), .A2(n10516), .ZN(n10521) );
  INV_X1 U13214 ( .A(n10517), .ZN(n10519) );
  NAND2_X1 U13215 ( .A1(n10519), .A2(n10518), .ZN(n11379) );
  INV_X1 U13216 ( .A(n11378), .ZN(n11210) );
  AND2_X1 U13217 ( .A1(n10640), .A2(n10549), .ZN(n11382) );
  INV_X1 U13218 ( .A(n10631), .ZN(n14850) );
  NAND3_X1 U13219 ( .A1(n15804), .A2(n11382), .A3(n14850), .ZN(n10520) );
  NAND2_X1 U13220 ( .A1(n10521), .A2(n15709), .ZN(n10546) );
  NAND2_X1 U13221 ( .A1(n14868), .A2(n15701), .ZN(n15367) );
  NAND2_X1 U13222 ( .A1(n10525), .A2(n11381), .ZN(n10856) );
  NAND2_X1 U13223 ( .A1(n10856), .A2(n11382), .ZN(n15699) );
  INV_X1 U13224 ( .A(n10522), .ZN(n10523) );
  NAND2_X1 U13225 ( .A1(n10856), .A2(n10523), .ZN(n10524) );
  INV_X1 U13226 ( .A(n15713), .ZN(n14639) );
  INV_X1 U13227 ( .A(n10525), .ZN(n10527) );
  NAND2_X1 U13228 ( .A1(n10527), .A2(n14956), .ZN(n14606) );
  INV_X1 U13229 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n10529) );
  OAI22_X1 U13230 ( .A1(n14823), .A2(n14681), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n10529), .ZN(n10542) );
  OAI21_X1 U13231 ( .B1(n10531), .B2(n10529), .A(n10528), .ZN(n10532) );
  NAND2_X1 U13232 ( .A1(P1_REG3_REG_27__SCAN_IN), .A2(P1_REG3_REG_28__SCAN_IN), 
        .ZN(n10530) );
  NAND2_X1 U13233 ( .A1(n14535), .A2(n8980), .ZN(n10540) );
  INV_X1 U13234 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n10537) );
  NAND2_X1 U13235 ( .A1(n10533), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n10535) );
  NAND2_X1 U13236 ( .A1(n10490), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n10534) );
  OAI211_X1 U13237 ( .C1(n10537), .C2(n10536), .A(n10535), .B(n10534), .ZN(
        n10538) );
  INV_X1 U13238 ( .A(n10538), .ZN(n10539) );
  NOR2_X1 U13239 ( .A1(n15352), .A2(n14680), .ZN(n10541) );
  AOI211_X1 U13240 ( .C1(n12738), .C2(n14639), .A(n10542), .B(n10541), .ZN(
        n10543) );
  OAI21_X1 U13241 ( .B1(n15367), .B2(n15699), .A(n10543), .ZN(n10544) );
  INV_X1 U13242 ( .A(n10544), .ZN(n10545) );
  NAND2_X1 U13243 ( .A1(n10546), .A2(n10545), .ZN(P1_U3214) );
  AND2_X1 U13244 ( .A1(n11021), .A2(n10547), .ZN(n10553) );
  INV_X1 U13245 ( .A(n10549), .ZN(n10550) );
  AND2_X2 U13246 ( .A1(n10640), .A2(n10550), .ZN(P1_U4016) );
  INV_X1 U13247 ( .A(P2_ADDR_REG_2__SCAN_IN), .ZN(n15646) );
  NAND2_X1 U13248 ( .A1(n11007), .A2(n11021), .ZN(n10551) );
  NAND2_X1 U13249 ( .A1(n10552), .A2(n10551), .ZN(n10555) );
  INV_X1 U13250 ( .A(n10553), .ZN(n10554) );
  NAND2_X1 U13251 ( .A1(n10555), .A2(n10554), .ZN(n10563) );
  OR2_X1 U13252 ( .A1(n10563), .A2(P2_U3088), .ZN(n15857) );
  NOR2_X1 U13253 ( .A1(n15646), .A2(n15857), .ZN(n10572) );
  NOR2_X1 U13254 ( .A1(n10102), .A2(P2_U3088), .ZN(n14457) );
  NAND2_X1 U13255 ( .A1(n10563), .A2(n14457), .ZN(n10565) );
  INV_X1 U13256 ( .A(n10565), .ZN(n10556) );
  INV_X1 U13257 ( .A(n14462), .ZN(n12378) );
  INV_X1 U13258 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n11328) );
  AND2_X1 U13259 ( .A1(P2_REG2_REG_0__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), 
        .ZN(n13821) );
  INV_X1 U13260 ( .A(n10574), .ZN(n13815) );
  NAND2_X1 U13261 ( .A1(n13815), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n10560) );
  NAND2_X1 U13262 ( .A1(n13819), .A2(n10560), .ZN(n10558) );
  INV_X1 U13263 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n10669) );
  MUX2_X1 U13264 ( .A(n10669), .B(P2_REG2_REG_2__SCAN_IN), .S(n10692), .Z(
        n10557) );
  NAND2_X1 U13265 ( .A1(n10558), .A2(n10557), .ZN(n10671) );
  MUX2_X1 U13266 ( .A(P2_REG2_REG_2__SCAN_IN), .B(n10669), .S(n6523), .Z(
        n10559) );
  NAND3_X1 U13267 ( .A1(n13819), .A2(n10560), .A3(n10559), .ZN(n10561) );
  AND3_X1 U13268 ( .A1(n15866), .A2(n10671), .A3(n10561), .ZN(n10571) );
  AND2_X1 U13269 ( .A1(n10102), .A2(P2_STATE_REG_SCAN_IN), .ZN(n10562) );
  NAND2_X1 U13270 ( .A1(n10563), .A2(n10562), .ZN(n15871) );
  INV_X1 U13271 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n10564) );
  OAI211_X1 U13272 ( .C1(n10567), .C2(n10566), .A(n15830), .B(n10691), .ZN(
        n10569) );
  NAND2_X1 U13273 ( .A1(P2_U3088), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n10568) );
  OAI211_X1 U13274 ( .C1(n15871), .C2(n6523), .A(n10569), .B(n10568), .ZN(
        n10570) );
  OR3_X1 U13275 ( .A1(n10572), .A2(n10571), .A3(n10570), .ZN(P2_U3216) );
  NAND2_X1 U13276 ( .A1(n6533), .A2(P2_U3088), .ZN(n14474) );
  AND2_X1 U13277 ( .A1(n10579), .A2(P2_U3088), .ZN(n14458) );
  INV_X2 U13278 ( .A(n14458), .ZN(n14472) );
  OAI222_X1 U13279 ( .A1(n10574), .A2(P2_U3088), .B1(n14474), .B2(n10578), 
        .C1(n10573), .C2(n14472), .ZN(P2_U3326) );
  NAND2_X1 U13280 ( .A1(n6532), .A2(P1_U3086), .ZN(n15539) );
  AND2_X1 U13281 ( .A1(n10579), .A2(P1_U3086), .ZN(n12162) );
  OAI222_X1 U13282 ( .A1(n15539), .A2(n10575), .B1(n15549), .B2(n10592), .C1(
        P1_U3086), .C2(n14994), .ZN(P1_U3353) );
  INV_X2 U13283 ( .A(n12162), .ZN(n15549) );
  OAI222_X1 U13284 ( .A1(n15539), .A2(n10576), .B1(n15549), .B2(n10590), .C1(
        P1_U3086), .C2(n10872), .ZN(P1_U3352) );
  INV_X1 U13285 ( .A(n15539), .ZN(n15527) );
  INV_X1 U13286 ( .A(n15527), .ZN(n15546) );
  OAI222_X1 U13287 ( .A1(n10752), .A2(P1_U3086), .B1(n15549), .B2(n10578), 
        .C1(n10577), .C2(n15546), .ZN(P1_U3354) );
  AND2_X1 U13288 ( .A1(n10579), .A2(P3_U3151), .ZN(n12081) );
  INV_X1 U13289 ( .A(n7298), .ZN(n10927) );
  NAND2_X1 U13290 ( .A1(n6532), .A2(P3_U3151), .ZN(n13528) );
  INV_X1 U13291 ( .A(n13528), .ZN(n13506) );
  AOI222_X1 U13292 ( .A1(n10581), .A2(n12081), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n10927), .C1(SI_2_), .C2(n13506), .ZN(n10582) );
  INV_X1 U13293 ( .A(n10582), .ZN(P3_U3293) );
  INV_X1 U13294 ( .A(P3_D_REG_1__SCAN_IN), .ZN(n10584) );
  NAND2_X1 U13295 ( .A1(n10709), .A2(n10722), .ZN(n10583) );
  OAI21_X1 U13296 ( .B1(n10722), .B2(n10584), .A(n10583), .ZN(P3_U3377) );
  INV_X1 U13297 ( .A(P3_D_REG_0__SCAN_IN), .ZN(n10587) );
  INV_X1 U13298 ( .A(n10707), .ZN(n10585) );
  NAND2_X1 U13299 ( .A1(n10585), .A2(n10722), .ZN(n10586) );
  OAI21_X1 U13300 ( .B1(n10722), .B2(n10587), .A(n10586), .ZN(P3_U3376) );
  INV_X1 U13301 ( .A(n10588), .ZN(n10594) );
  OAI222_X1 U13302 ( .A1(n15539), .A2(n10589), .B1(n15549), .B2(n10594), .C1(
        P1_U3086), .C2(n15010), .ZN(P1_U3351) );
  INV_X1 U13303 ( .A(n14474), .ZN(n12165) );
  INV_X1 U13304 ( .A(n12165), .ZN(n14461) );
  OAI222_X1 U13305 ( .A1(n14472), .A2(n10591), .B1(n14461), .B2(n10590), .C1(
        P2_U3088), .C2(n10693), .ZN(P2_U3324) );
  OAI222_X1 U13306 ( .A1(n14472), .A2(n10593), .B1(n14461), .B2(n10592), .C1(
        P2_U3088), .C2(n6523), .ZN(P2_U3325) );
  OAI222_X1 U13307 ( .A1(n14472), .A2(n10595), .B1(n14461), .B2(n10594), .C1(
        P2_U3088), .C2(n13830), .ZN(P2_U3323) );
  INV_X1 U13308 ( .A(n13506), .ZN(n13521) );
  INV_X1 U13309 ( .A(n10596), .ZN(n10597) );
  OAI222_X1 U13310 ( .A1(P3_U3151), .A2(n10921), .B1(n13521), .B2(n10598), 
        .C1(n13524), .C2(n10597), .ZN(P3_U3294) );
  INV_X2 U13311 ( .A(n12081), .ZN(n13524) );
  INV_X1 U13312 ( .A(n10599), .ZN(n10601) );
  INV_X1 U13313 ( .A(SI_8_), .ZN(n10600) );
  INV_X1 U13314 ( .A(n11574), .ZN(n11577) );
  OAI222_X1 U13315 ( .A1(n13524), .A2(n10601), .B1(n13521), .B2(n10600), .C1(
        n11577), .C2(P3_U3151), .ZN(P3_U3287) );
  OAI222_X1 U13316 ( .A1(n13524), .A2(n10603), .B1(n13521), .B2(n10602), .C1(
        n12089), .C2(P3_U3151), .ZN(P3_U3285) );
  INV_X1 U13317 ( .A(SI_4_), .ZN(n10604) );
  OAI222_X1 U13318 ( .A1(n13524), .A2(n10605), .B1(n13521), .B2(n10604), .C1(
        n10976), .C2(P3_U3151), .ZN(P3_U3291) );
  INV_X1 U13319 ( .A(SI_5_), .ZN(n10606) );
  OAI222_X1 U13320 ( .A1(n13524), .A2(n10607), .B1(n13521), .B2(n10606), .C1(
        n10979), .C2(P3_U3151), .ZN(P3_U3290) );
  INV_X1 U13321 ( .A(SI_3_), .ZN(n10608) );
  OAI222_X1 U13322 ( .A1(n10961), .A2(P3_U3151), .B1(n13524), .B2(n10609), 
        .C1(n10608), .C2(n13521), .ZN(P3_U3292) );
  OAI222_X1 U13323 ( .A1(n11594), .A2(P3_U3151), .B1(n13524), .B2(n10611), 
        .C1(n10610), .C2(n13521), .ZN(P3_U3286) );
  INV_X1 U13324 ( .A(n11036), .ZN(n11046) );
  INV_X1 U13325 ( .A(n10612), .ZN(n10614) );
  INV_X1 U13326 ( .A(SI_6_), .ZN(n10613) );
  OAI222_X1 U13327 ( .A1(n11046), .A2(P3_U3151), .B1(n13524), .B2(n10614), 
        .C1(n10613), .C2(n13521), .ZN(P3_U3289) );
  OAI222_X1 U13328 ( .A1(n11192), .A2(P3_U3151), .B1(n13524), .B2(n10616), 
        .C1(n10615), .C2(n13521), .ZN(P3_U3288) );
  INV_X1 U13329 ( .A(n10617), .ZN(n10619) );
  OAI222_X1 U13330 ( .A1(n15539), .A2(n10618), .B1(n15549), .B2(n10619), .C1(
        P1_U3086), .C2(n7243), .ZN(P1_U3350) );
  OAI222_X1 U13331 ( .A1(n14472), .A2(n10620), .B1(n14461), .B2(n10619), .C1(
        P2_U3088), .C2(n13842), .ZN(P2_U3322) );
  AND2_X1 U13332 ( .A1(n10622), .A2(P3_D_REG_11__SCAN_IN), .ZN(P3_U3254) );
  AND2_X1 U13333 ( .A1(n10622), .A2(P3_D_REG_27__SCAN_IN), .ZN(P3_U3238) );
  AND2_X1 U13334 ( .A1(n10622), .A2(P3_D_REG_25__SCAN_IN), .ZN(P3_U3240) );
  AND2_X1 U13335 ( .A1(n10622), .A2(P3_D_REG_10__SCAN_IN), .ZN(P3_U3255) );
  AND2_X1 U13336 ( .A1(n10622), .A2(P3_D_REG_28__SCAN_IN), .ZN(P3_U3237) );
  AND2_X1 U13337 ( .A1(n10622), .A2(P3_D_REG_7__SCAN_IN), .ZN(P3_U3258) );
  AND2_X1 U13338 ( .A1(n10622), .A2(P3_D_REG_8__SCAN_IN), .ZN(P3_U3257) );
  AND2_X1 U13339 ( .A1(n10622), .A2(P3_D_REG_9__SCAN_IN), .ZN(P3_U3256) );
  AND2_X1 U13340 ( .A1(n10622), .A2(P3_D_REG_5__SCAN_IN), .ZN(P3_U3260) );
  AND2_X1 U13341 ( .A1(n10622), .A2(P3_D_REG_15__SCAN_IN), .ZN(P3_U3250) );
  AND2_X1 U13342 ( .A1(n10622), .A2(P3_D_REG_12__SCAN_IN), .ZN(P3_U3253) );
  AND2_X1 U13343 ( .A1(n10622), .A2(P3_D_REG_13__SCAN_IN), .ZN(P3_U3252) );
  AND2_X1 U13344 ( .A1(n10622), .A2(P3_D_REG_14__SCAN_IN), .ZN(P3_U3251) );
  AND2_X1 U13345 ( .A1(n10622), .A2(P3_D_REG_22__SCAN_IN), .ZN(P3_U3243) );
  AND2_X1 U13346 ( .A1(n10622), .A2(P3_D_REG_6__SCAN_IN), .ZN(P3_U3259) );
  AND2_X1 U13347 ( .A1(n10622), .A2(P3_D_REG_24__SCAN_IN), .ZN(P3_U3241) );
  AND2_X1 U13348 ( .A1(n10622), .A2(P3_D_REG_3__SCAN_IN), .ZN(P3_U3262) );
  AND2_X1 U13349 ( .A1(n10622), .A2(P3_D_REG_26__SCAN_IN), .ZN(P3_U3239) );
  AND2_X1 U13350 ( .A1(n10622), .A2(P3_D_REG_17__SCAN_IN), .ZN(P3_U3248) );
  AND2_X1 U13351 ( .A1(n10622), .A2(P3_D_REG_31__SCAN_IN), .ZN(P3_U3234) );
  AND2_X1 U13352 ( .A1(n10622), .A2(P3_D_REG_29__SCAN_IN), .ZN(P3_U3236) );
  AND2_X1 U13353 ( .A1(n10622), .A2(P3_D_REG_30__SCAN_IN), .ZN(P3_U3235) );
  AND2_X1 U13354 ( .A1(n10622), .A2(P3_D_REG_2__SCAN_IN), .ZN(P3_U3263) );
  AND2_X1 U13355 ( .A1(n10622), .A2(P3_D_REG_21__SCAN_IN), .ZN(P3_U3244) );
  AND2_X1 U13356 ( .A1(n10622), .A2(P3_D_REG_16__SCAN_IN), .ZN(P3_U3249) );
  AND2_X1 U13357 ( .A1(n10622), .A2(P3_D_REG_20__SCAN_IN), .ZN(P3_U3245) );
  AND2_X1 U13358 ( .A1(n10622), .A2(P3_D_REG_19__SCAN_IN), .ZN(P3_U3246) );
  AND2_X1 U13359 ( .A1(n10622), .A2(P3_D_REG_23__SCAN_IN), .ZN(P3_U3242) );
  AND2_X1 U13360 ( .A1(n10622), .A2(P3_D_REG_4__SCAN_IN), .ZN(P3_U3261) );
  INV_X1 U13361 ( .A(n10622), .ZN(n10623) );
  NOR2_X1 U13362 ( .A1(n10623), .A2(n9332), .ZN(P3_U3247) );
  INV_X1 U13363 ( .A(n10624), .ZN(n10626) );
  INV_X1 U13364 ( .A(n13857), .ZN(n13851) );
  OAI222_X1 U13365 ( .A1(n14472), .A2(n10625), .B1(n14461), .B2(n10626), .C1(
        P2_U3088), .C2(n13851), .ZN(P2_U3321) );
  OAI222_X1 U13366 ( .A1(n15539), .A2(n10627), .B1(n15549), .B2(n10626), .C1(
        P1_U3086), .C2(n10832), .ZN(P1_U3349) );
  OR2_X1 U13367 ( .A1(n10630), .A2(P1_U3086), .ZN(n14959) );
  INV_X1 U13368 ( .A(n14959), .ZN(n10628) );
  AOI21_X1 U13369 ( .B1(n10631), .B2(n10630), .A(n10629), .ZN(n10740) );
  INV_X1 U13370 ( .A(n10740), .ZN(n10632) );
  NOR2_X1 U13371 ( .A1(n15722), .A2(P1_U4016), .ZN(P1_U3085) );
  OAI222_X1 U13372 ( .A1(n12975), .A2(P3_U3151), .B1(n13524), .B2(n10634), 
        .C1(n10633), .C2(n13521), .ZN(P3_U3284) );
  INV_X1 U13373 ( .A(n10635), .ZN(n10637) );
  INV_X1 U13374 ( .A(n11148), .ZN(n10851) );
  OAI222_X1 U13375 ( .A1(n15546), .A2(n10636), .B1(n15549), .B2(n10637), .C1(
        P1_U3086), .C2(n10851), .ZN(P1_U3348) );
  INV_X1 U13376 ( .A(n13871), .ZN(n13868) );
  OAI222_X1 U13377 ( .A1(n14472), .A2(n10638), .B1(n14461), .B2(n10637), .C1(
        P2_U3088), .C2(n13868), .ZN(P2_U3320) );
  AND2_X2 U13378 ( .A1(n11382), .A2(n10639), .ZN(n15781) );
  INV_X1 U13379 ( .A(n10640), .ZN(n10645) );
  OAI22_X1 U13380 ( .A1(n15781), .A2(P1_D_REG_1__SCAN_IN), .B1(n10645), .B2(
        n10641), .ZN(n10642) );
  INV_X1 U13381 ( .A(n10642), .ZN(P1_U3446) );
  INV_X1 U13382 ( .A(n10643), .ZN(n10644) );
  OAI22_X1 U13383 ( .A1(n15781), .A2(P1_D_REG_0__SCAN_IN), .B1(n10645), .B2(
        n10644), .ZN(n10646) );
  INV_X1 U13384 ( .A(n10646), .ZN(P1_U3445) );
  INV_X2 U13385 ( .A(P2_U3947), .ZN(n13811) );
  NAND2_X1 U13386 ( .A1(P2_DATAO_REG_30__SCAN_IN), .A2(n13811), .ZN(n10647) );
  OAI21_X1 U13387 ( .B1(n12380), .B2(n13811), .A(n10647), .ZN(P2_U3561) );
  NAND2_X1 U13388 ( .A1(P3_U3897), .A2(n12344), .ZN(n10648) );
  OAI21_X1 U13389 ( .B1(P3_U3897), .B2(n10649), .A(n10648), .ZN(P3_U3495) );
  NAND2_X1 U13390 ( .A1(P3_U3897), .A2(n10796), .ZN(n10650) );
  OAI21_X1 U13391 ( .B1(P3_U3897), .B2(n10651), .A(n10650), .ZN(P3_U3491) );
  INV_X1 U13392 ( .A(n10652), .ZN(n10654) );
  OAI222_X1 U13393 ( .A1(n13524), .A2(n10654), .B1(n13521), .B2(n10653), .C1(
        n13008), .C2(P3_U3151), .ZN(P3_U3283) );
  INV_X1 U13394 ( .A(n10655), .ZN(n10658) );
  INV_X1 U13395 ( .A(n10878), .ZN(n10874) );
  OAI222_X1 U13396 ( .A1(n14472), .A2(n10656), .B1(n14461), .B2(n10658), .C1(
        P2_U3088), .C2(n10874), .ZN(P2_U3319) );
  INV_X1 U13397 ( .A(n15030), .ZN(n10657) );
  OAI222_X1 U13398 ( .A1(n15539), .A2(n10659), .B1(n15549), .B2(n10658), .C1(
        P1_U3086), .C2(n10657), .ZN(P1_U3347) );
  OAI222_X1 U13399 ( .A1(n13524), .A2(n10661), .B1(n13521), .B2(n10660), .C1(
        n13027), .C2(P3_U3151), .ZN(P3_U3282) );
  OAI222_X1 U13400 ( .A1(n13524), .A2(n10663), .B1(n13521), .B2(n10662), .C1(
        n13042), .C2(P3_U3151), .ZN(P3_U3281) );
  INV_X1 U13401 ( .A(n10664), .ZN(n10666) );
  INV_X1 U13402 ( .A(n11177), .ZN(n11171) );
  OAI222_X1 U13403 ( .A1(n14472), .A2(n10665), .B1(n14461), .B2(n10666), .C1(
        P2_U3088), .C2(n11171), .ZN(P2_U3318) );
  INV_X1 U13404 ( .A(n11231), .ZN(n11236) );
  OAI222_X1 U13405 ( .A1(n15539), .A2(n10667), .B1(n15549), .B2(n10666), .C1(
        P1_U3086), .C2(n11236), .ZN(P1_U3346) );
  INV_X1 U13406 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n10668) );
  NAND2_X1 U13407 ( .A1(P2_U3088), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n12046) );
  OAI21_X1 U13408 ( .B1(n15857), .B2(n10668), .A(n12046), .ZN(n10690) );
  OR2_X1 U13409 ( .A1(n6523), .A2(n10669), .ZN(n10670) );
  NAND2_X1 U13410 ( .A1(n10671), .A2(n10670), .ZN(n15839) );
  INV_X1 U13411 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n11563) );
  MUX2_X1 U13412 ( .A(n11563), .B(P2_REG2_REG_3__SCAN_IN), .S(n10693), .Z(
        n15838) );
  INV_X1 U13413 ( .A(n10693), .ZN(n15836) );
  NAND2_X1 U13414 ( .A1(n15836), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n13832) );
  NAND2_X1 U13415 ( .A1(n15837), .A2(n13832), .ZN(n10673) );
  INV_X1 U13416 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n11504) );
  MUX2_X1 U13417 ( .A(n11504), .B(P2_REG2_REG_4__SCAN_IN), .S(n13830), .Z(
        n10672) );
  INV_X1 U13418 ( .A(n13830), .ZN(n10674) );
  NAND2_X1 U13419 ( .A1(n10674), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n13844) );
  NAND2_X1 U13420 ( .A1(n13845), .A2(n13844), .ZN(n10676) );
  INV_X1 U13421 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n11929) );
  MUX2_X1 U13422 ( .A(n11929), .B(P2_REG2_REG_5__SCAN_IN), .S(n13842), .Z(
        n10675) );
  NAND2_X1 U13423 ( .A1(n10677), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n13859) );
  NAND2_X1 U13424 ( .A1(n13860), .A2(n13859), .ZN(n10680) );
  INV_X1 U13425 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n10678) );
  MUX2_X1 U13426 ( .A(P2_REG2_REG_6__SCAN_IN), .B(n10678), .S(n13857), .Z(
        n10679) );
  NAND2_X1 U13427 ( .A1(n13857), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n13873) );
  NAND2_X1 U13428 ( .A1(n13874), .A2(n13873), .ZN(n10682) );
  INV_X1 U13429 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n12068) );
  MUX2_X1 U13430 ( .A(P2_REG2_REG_7__SCAN_IN), .B(n12068), .S(n13871), .Z(
        n10681) );
  NAND2_X1 U13431 ( .A1(n13871), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n10687) );
  NAND2_X1 U13432 ( .A1(n13876), .A2(n10687), .ZN(n10685) );
  INV_X1 U13433 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n10683) );
  MUX2_X1 U13434 ( .A(P2_REG2_REG_8__SCAN_IN), .B(n10683), .S(n10878), .Z(
        n10684) );
  NAND2_X1 U13435 ( .A1(n10685), .A2(n10684), .ZN(n10880) );
  MUX2_X1 U13436 ( .A(n10683), .B(P2_REG2_REG_8__SCAN_IN), .S(n10878), .Z(
        n10686) );
  NAND3_X1 U13437 ( .A1(n13876), .A2(n10687), .A3(n10686), .ZN(n10688) );
  AND3_X1 U13438 ( .A1(n10880), .A2(n15866), .A3(n10688), .ZN(n10689) );
  AOI211_X1 U13439 ( .C1(n15850), .C2(n10878), .A(n10690), .B(n10689), .ZN(
        n10702) );
  INV_X1 U13440 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n10698) );
  INV_X1 U13441 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n10697) );
  INV_X1 U13442 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n10696) );
  INV_X1 U13443 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n10695) );
  INV_X1 U13444 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n10694) );
  INV_X1 U13445 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n11261) );
  MUX2_X1 U13446 ( .A(n10694), .B(P2_REG1_REG_3__SCAN_IN), .S(n10693), .Z(
        n15832) );
  MUX2_X1 U13447 ( .A(n10695), .B(P2_REG1_REG_4__SCAN_IN), .S(n13830), .Z(
        n13829) );
  MUX2_X1 U13448 ( .A(n10696), .B(P2_REG1_REG_5__SCAN_IN), .S(n13842), .Z(
        n13841) );
  MUX2_X1 U13449 ( .A(P2_REG1_REG_6__SCAN_IN), .B(n10697), .S(n13857), .Z(
        n13855) );
  OAI21_X1 U13450 ( .B1(n10697), .B2(n13851), .A(n13854), .ZN(n13867) );
  MUX2_X1 U13451 ( .A(P2_REG1_REG_7__SCAN_IN), .B(n10698), .S(n13871), .Z(
        n13866) );
  NAND2_X1 U13452 ( .A1(n13867), .A2(n13866), .ZN(n13865) );
  XOR2_X1 U13453 ( .A(P2_REG1_REG_8__SCAN_IN), .B(n10878), .Z(n10699) );
  OAI211_X1 U13454 ( .C1(n10700), .C2(n10699), .A(n10873), .B(n15830), .ZN(
        n10701) );
  NAND2_X1 U13455 ( .A1(n10702), .A2(n10701), .ZN(P2_U3222) );
  INV_X1 U13456 ( .A(n10708), .ZN(n10703) );
  NAND2_X1 U13457 ( .A1(n12490), .A2(n10705), .ZN(n12634) );
  OR2_X1 U13458 ( .A1(n10706), .A2(n12634), .ZN(n10802) );
  NOR2_X1 U13459 ( .A1(n10708), .A2(n10707), .ZN(n10710) );
  AND2_X1 U13460 ( .A1(n10710), .A2(n10709), .ZN(n10803) );
  INV_X1 U13461 ( .A(n10711), .ZN(n10799) );
  OR2_X1 U13462 ( .A1(n10803), .A2(n10799), .ZN(n10716) );
  INV_X1 U13463 ( .A(n10712), .ZN(n10713) );
  AND2_X1 U13464 ( .A1(n10714), .A2(n10713), .ZN(n10715) );
  OAI211_X1 U13465 ( .C1(n10801), .C2(n10802), .A(n10716), .B(n10715), .ZN(
        n10717) );
  NAND2_X1 U13466 ( .A1(n10717), .A2(P3_STATE_REG_SCAN_IN), .ZN(n10721) );
  NAND2_X1 U13467 ( .A1(n12626), .A2(n12632), .ZN(n10718) );
  INV_X1 U13468 ( .A(n12642), .ZN(n10719) );
  OR2_X1 U13469 ( .A1(n10801), .A2(n10719), .ZN(n10720) );
  AND2_X1 U13470 ( .A1(n11090), .A2(n10722), .ZN(n11001) );
  INV_X1 U13471 ( .A(n10802), .ZN(n10723) );
  NAND2_X1 U13472 ( .A1(n10801), .A2(n10723), .ZN(n10727) );
  INV_X1 U13473 ( .A(n10724), .ZN(n10725) );
  NAND2_X1 U13474 ( .A1(n10803), .A2(n10725), .ZN(n10726) );
  NAND2_X1 U13475 ( .A1(n10727), .A2(n10726), .ZN(n10729) );
  INV_X1 U13476 ( .A(n10895), .ZN(n10728) );
  NAND2_X1 U13477 ( .A1(n10796), .A2(n11190), .ZN(n12491) );
  NAND2_X1 U13478 ( .A1(n12494), .A2(n12491), .ZN(n12444) );
  OR2_X1 U13479 ( .A1(n10803), .A2(n10731), .ZN(n10733) );
  AND2_X1 U13480 ( .A1(n12642), .A2(n10734), .ZN(n10735) );
  OAI22_X1 U13481 ( .A1(n12937), .A2(n11190), .B1(n12931), .B2(n11343), .ZN(
        n10736) );
  AOI21_X1 U13482 ( .B1(n12924), .B2(n12444), .A(n10736), .ZN(n10737) );
  OAI21_X1 U13483 ( .B1(n11001), .B2(n10817), .A(n10737), .ZN(P3_U3172) );
  OAI222_X1 U13484 ( .A1(n13063), .A2(P3_U3151), .B1(n13524), .B2(n10739), 
        .C1(n10738), .C2(n13521), .ZN(P3_U3280) );
  NAND2_X1 U13485 ( .A1(n10741), .A2(n10740), .ZN(n15725) );
  INV_X1 U13486 ( .A(n15010), .ZN(n15009) );
  INV_X1 U13487 ( .A(n10872), .ZN(n10745) );
  INV_X1 U13488 ( .A(n14994), .ZN(n14989) );
  INV_X1 U13489 ( .A(n10752), .ZN(n14976) );
  MUX2_X1 U13490 ( .A(P1_REG1_REG_1__SCAN_IN), .B(n8664), .S(n10752), .Z(
        n14973) );
  NOR3_X1 U13491 ( .A1(n14973), .A2(n15717), .A3(n10743), .ZN(n14972) );
  XOR2_X1 U13492 ( .A(P1_REG1_REG_2__SCAN_IN), .B(n14994), .Z(n14983) );
  INV_X1 U13493 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n10744) );
  MUX2_X1 U13494 ( .A(P1_REG1_REG_3__SCAN_IN), .B(n10744), .S(n10872), .Z(
        n10863) );
  NOR2_X1 U13495 ( .A1(n10864), .A2(n10863), .ZN(n10862) );
  AOI21_X1 U13496 ( .B1(n10745), .B2(P1_REG1_REG_3__SCAN_IN), .A(n10862), .ZN(
        n15005) );
  INV_X1 U13497 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n10746) );
  MUX2_X1 U13498 ( .A(P1_REG1_REG_4__SCAN_IN), .B(n10746), .S(n15010), .Z(
        n15004) );
  AOI21_X1 U13499 ( .B1(n15009), .B2(P1_REG1_REG_4__SCAN_IN), .A(n15003), .ZN(
        n10749) );
  MUX2_X1 U13500 ( .A(P1_REG1_REG_5__SCAN_IN), .B(n10747), .S(n10822), .Z(
        n10748) );
  NAND2_X1 U13501 ( .A1(n10749), .A2(n10748), .ZN(n10819) );
  OAI21_X1 U13502 ( .B1(n10749), .B2(n10748), .A(n10819), .ZN(n10769) );
  INV_X1 U13503 ( .A(n15536), .ZN(n15714) );
  INV_X1 U13504 ( .A(n15725), .ZN(n10751) );
  NOR2_X1 U13505 ( .A1(n15533), .A2(n15536), .ZN(n10750) );
  NAND2_X1 U13506 ( .A1(n10751), .A2(n10750), .ZN(n15099) );
  INV_X1 U13507 ( .A(n15099), .ZN(n15746) );
  MUX2_X1 U13508 ( .A(n11525), .B(P1_REG2_REG_3__SCAN_IN), .S(n10872), .Z(
        n10758) );
  MUX2_X1 U13509 ( .A(n10753), .B(P1_REG2_REG_1__SCAN_IN), .S(n10752), .Z(
        n14977) );
  AND2_X1 U13510 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n10754) );
  NAND2_X1 U13511 ( .A1(n14977), .A2(n10754), .ZN(n14997) );
  NAND2_X1 U13512 ( .A1(n14976), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n14995) );
  NAND2_X1 U13513 ( .A1(n14997), .A2(n14995), .ZN(n10756) );
  MUX2_X1 U13514 ( .A(n11692), .B(P1_REG2_REG_2__SCAN_IN), .S(n14994), .Z(
        n10755) );
  NAND2_X1 U13515 ( .A1(n10756), .A2(n10755), .ZN(n14999) );
  NAND2_X1 U13516 ( .A1(n14989), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n10865) );
  NAND2_X1 U13517 ( .A1(n14999), .A2(n10865), .ZN(n10757) );
  NAND2_X1 U13518 ( .A1(n10758), .A2(n10757), .ZN(n15013) );
  OR2_X1 U13519 ( .A1(n10872), .A2(n11525), .ZN(n15012) );
  NAND2_X1 U13520 ( .A1(n15013), .A2(n15012), .ZN(n10761) );
  MUX2_X1 U13521 ( .A(n10759), .B(P1_REG2_REG_4__SCAN_IN), .S(n15010), .Z(
        n10760) );
  NAND2_X1 U13522 ( .A1(n10761), .A2(n10760), .ZN(n15015) );
  NAND2_X1 U13523 ( .A1(n15009), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n10766) );
  NAND2_X1 U13524 ( .A1(n15015), .A2(n10766), .ZN(n10764) );
  INV_X1 U13525 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n10762) );
  MUX2_X1 U13526 ( .A(P1_REG2_REG_5__SCAN_IN), .B(n10762), .S(n10822), .Z(
        n10763) );
  NAND2_X1 U13527 ( .A1(n10764), .A2(n10763), .ZN(n10827) );
  MUX2_X1 U13528 ( .A(n10762), .B(P1_REG2_REG_5__SCAN_IN), .S(n10822), .Z(
        n10765) );
  NAND3_X1 U13529 ( .A1(n15015), .A2(n10766), .A3(n10765), .ZN(n10767) );
  AND3_X1 U13530 ( .A1(n15746), .A2(n10827), .A3(n10767), .ZN(n10768) );
  AOI21_X1 U13531 ( .B1(n10769), .B2(n15745), .A(n10768), .ZN(n10772) );
  NAND2_X1 U13532 ( .A1(P1_U3086), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n11624) );
  INV_X1 U13533 ( .A(n11624), .ZN(n10770) );
  AOI21_X1 U13534 ( .B1(n15722), .B2(P1_ADDR_REG_5__SCAN_IN), .A(n10770), .ZN(
        n10771) );
  OAI211_X1 U13535 ( .C1(n7243), .C2(n15068), .A(n10772), .B(n10771), .ZN(
        P1_U3248) );
  INV_X1 U13536 ( .A(n10773), .ZN(n10775) );
  INV_X1 U13537 ( .A(n11655), .ZN(n11175) );
  OAI222_X1 U13538 ( .A1(n14472), .A2(n10774), .B1(n14461), .B2(n10775), .C1(
        P2_U3088), .C2(n11175), .ZN(P2_U3317) );
  INV_X1 U13539 ( .A(n11239), .ZN(n11482) );
  OAI222_X1 U13540 ( .A1(n15539), .A2(n10776), .B1(n15549), .B2(n10775), .C1(
        P1_U3086), .C2(n11482), .ZN(P1_U3345) );
  INV_X1 U13541 ( .A(P3_REG3_REG_1__SCAN_IN), .ZN(n10793) );
  INV_X1 U13542 ( .A(n11310), .ZN(n11365) );
  AND2_X1 U13543 ( .A1(n12642), .A2(n10777), .ZN(n10778) );
  INV_X1 U13544 ( .A(n10796), .ZN(n10779) );
  OAI22_X1 U13545 ( .A1(n12917), .A2(n10779), .B1(n11089), .B2(n12931), .ZN(
        n10780) );
  AOI21_X1 U13546 ( .B1(n12919), .B2(n11365), .A(n10780), .ZN(n10792) );
  OAI21_X1 U13547 ( .B1(n10782), .B2(n12634), .A(n10781), .ZN(n10783) );
  INV_X2 U13548 ( .A(n10783), .ZN(n11759) );
  INV_X1 U13549 ( .A(n10794), .ZN(n10786) );
  OAI21_X1 U13550 ( .B1(n10786), .B2(n12832), .A(n10785), .ZN(n10787) );
  OAI211_X1 U13551 ( .C1(n10789), .C2(n10794), .A(n10993), .B(n10788), .ZN(
        n10790) );
  NAND2_X1 U13552 ( .A1(n10790), .A2(n12924), .ZN(n10791) );
  OAI211_X1 U13553 ( .C1(n11001), .C2(n10793), .A(n10792), .B(n10791), .ZN(
        P3_U3162) );
  NAND2_X1 U13554 ( .A1(n10795), .A2(n13336), .ZN(n10798) );
  AOI22_X1 U13555 ( .A1(n13339), .A2(n10796), .B1(n12953), .B2(n13340), .ZN(
        n10797) );
  NAND2_X1 U13556 ( .A1(n10798), .A2(n10797), .ZN(n11364) );
  AOI21_X1 U13557 ( .B1(n13407), .B2(n11368), .A(n11364), .ZN(n11313) );
  NOR2_X1 U13558 ( .A1(n10799), .A2(n10895), .ZN(n10800) );
  NAND2_X1 U13559 ( .A1(n10801), .A2(n10800), .ZN(n10806) );
  NOR2_X1 U13560 ( .A1(n10895), .A2(n10802), .ZN(n10804) );
  OAI21_X1 U13561 ( .B1(n12642), .B2(n10804), .A(n10803), .ZN(n10805) );
  INV_X2 U13562 ( .A(n15961), .ZN(n15963) );
  INV_X1 U13563 ( .A(P3_REG0_REG_1__SCAN_IN), .ZN(n10807) );
  OAI22_X1 U13564 ( .A1(n11310), .A2(n13493), .B1(n15963), .B2(n10807), .ZN(
        n10808) );
  INV_X1 U13565 ( .A(n10808), .ZN(n10809) );
  OAI21_X1 U13566 ( .B1(n11313), .B2(n15961), .A(n10809), .ZN(P3_U3393) );
  AND2_X1 U13567 ( .A1(n12598), .A2(n15946), .ZN(n10811) );
  AND2_X1 U13568 ( .A1(n12954), .A2(n13340), .ZN(n10810) );
  AOI21_X1 U13569 ( .B1(n12444), .B2(n10811), .A(n10810), .ZN(n11187) );
  INV_X1 U13570 ( .A(P3_REG0_REG_0__SCAN_IN), .ZN(n10812) );
  MUX2_X1 U13571 ( .A(n11187), .B(n10812), .S(n15961), .Z(n10813) );
  OAI21_X1 U13572 ( .B1(n11190), .B2(n13493), .A(n10813), .ZN(P3_U3390) );
  INV_X1 U13573 ( .A(P3_REG2_REG_0__SCAN_IN), .ZN(n10901) );
  MUX2_X1 U13574 ( .A(n10901), .B(n11187), .S(n13350), .Z(n10816) );
  NAND2_X1 U13575 ( .A1(n13310), .A2(n10814), .ZN(n10815) );
  OAI211_X1 U13576 ( .C1(n10817), .C2(n13321), .A(n10816), .B(n10815), .ZN(
        P3_U3233) );
  INV_X1 U13577 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n10818) );
  MUX2_X1 U13578 ( .A(P1_REG1_REG_6__SCAN_IN), .B(n10818), .S(n10832), .Z(
        n10821) );
  AOI211_X1 U13579 ( .C1(n10821), .C2(n10820), .A(n15097), .B(n10839), .ZN(
        n10834) );
  NAND2_X1 U13580 ( .A1(n10822), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n10826) );
  NAND2_X1 U13581 ( .A1(n10827), .A2(n10826), .ZN(n10824) );
  MUX2_X1 U13582 ( .A(n11859), .B(P1_REG2_REG_6__SCAN_IN), .S(n10832), .Z(
        n10823) );
  NAND2_X1 U13583 ( .A1(n10824), .A2(n10823), .ZN(n10848) );
  MUX2_X1 U13584 ( .A(P1_REG2_REG_6__SCAN_IN), .B(n11859), .S(n10832), .Z(
        n10825) );
  NAND3_X1 U13585 ( .A1(n10827), .A2(n10826), .A3(n10825), .ZN(n10828) );
  NAND3_X1 U13586 ( .A1(n15746), .A2(n10848), .A3(n10828), .ZN(n10831) );
  AND2_X1 U13587 ( .A1(P1_U3086), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n10829) );
  AOI21_X1 U13588 ( .B1(n15722), .B2(P1_ADDR_REG_6__SCAN_IN), .A(n10829), .ZN(
        n10830) );
  OAI211_X1 U13589 ( .C1(n15068), .C2(n10832), .A(n10831), .B(n10830), .ZN(
        n10833) );
  OR2_X1 U13590 ( .A1(n10834), .A2(n10833), .ZN(P1_U3249) );
  INV_X1 U13591 ( .A(n10835), .ZN(n10837) );
  INV_X1 U13592 ( .A(n11483), .ZN(n11984) );
  OAI222_X1 U13593 ( .A1(n15539), .A2(n10836), .B1(n15549), .B2(n10837), .C1(
        P1_U3086), .C2(n11984), .ZN(P1_U3344) );
  INV_X1 U13594 ( .A(n11826), .ZN(n11659) );
  OAI222_X1 U13595 ( .A1(n14472), .A2(n10838), .B1(n14461), .B2(n10837), .C1(
        P2_U3088), .C2(n11659), .ZN(P2_U3316) );
  MUX2_X1 U13596 ( .A(n10840), .B(P1_REG1_REG_7__SCAN_IN), .S(n11148), .Z(
        n10841) );
  AOI211_X1 U13597 ( .C1(n10842), .C2(n10841), .A(n15097), .B(n11146), .ZN(
        n10854) );
  NAND2_X1 U13598 ( .A1(n10843), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n10847) );
  NAND2_X1 U13599 ( .A1(n10848), .A2(n10847), .ZN(n10845) );
  MUX2_X1 U13600 ( .A(P1_REG2_REG_7__SCAN_IN), .B(n12158), .S(n11148), .Z(
        n10844) );
  NAND2_X1 U13601 ( .A1(n10845), .A2(n10844), .ZN(n15027) );
  MUX2_X1 U13602 ( .A(n12158), .B(P1_REG2_REG_7__SCAN_IN), .S(n11148), .Z(
        n10846) );
  NAND3_X1 U13603 ( .A1(n10848), .A2(n10847), .A3(n10846), .ZN(n10849) );
  AND3_X1 U13604 ( .A1(n15746), .A2(n15027), .A3(n10849), .ZN(n10853) );
  NAND2_X1 U13605 ( .A1(P1_U3086), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n14479) );
  NAND2_X1 U13606 ( .A1(n15722), .A2(P1_ADDR_REG_7__SCAN_IN), .ZN(n10850) );
  OAI211_X1 U13607 ( .C1(n15068), .C2(n10851), .A(n14479), .B(n10850), .ZN(
        n10852) );
  OR3_X1 U13608 ( .A1(n10854), .A2(n10853), .A3(n10852), .ZN(P1_U3250) );
  INV_X1 U13609 ( .A(n14680), .ZN(n14667) );
  NAND2_X1 U13610 ( .A1(n10856), .A2(n14956), .ZN(n11316) );
  AOI22_X1 U13611 ( .A1(n14667), .A2(n10855), .B1(P1_REG3_REG_0__SCAN_IN), 
        .B2(n11316), .ZN(n10861) );
  OAI21_X1 U13612 ( .B1(n10859), .B2(n10858), .A(n10857), .ZN(n14990) );
  NAND2_X1 U13613 ( .A1(n14990), .A2(n15709), .ZN(n10860) );
  OAI211_X1 U13614 ( .C1(n14676), .C2(n11371), .A(n10861), .B(n10860), .ZN(
        P1_U3232) );
  AOI211_X1 U13615 ( .C1(n10864), .C2(n10863), .A(n10862), .B(n15097), .ZN(
        n10869) );
  MUX2_X1 U13616 ( .A(P1_REG2_REG_3__SCAN_IN), .B(n11525), .S(n10872), .Z(
        n10866) );
  NAND3_X1 U13617 ( .A1(n10866), .A2(n14999), .A3(n10865), .ZN(n10867) );
  AND3_X1 U13618 ( .A1(n15746), .A2(n15013), .A3(n10867), .ZN(n10868) );
  NOR2_X1 U13619 ( .A1(n10869), .A2(n10868), .ZN(n10871) );
  AND2_X1 U13620 ( .A1(P1_U3086), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n15702) );
  AOI21_X1 U13621 ( .B1(n15722), .B2(P1_ADDR_REG_3__SCAN_IN), .A(n15702), .ZN(
        n10870) );
  OAI211_X1 U13622 ( .C1(n10872), .C2(n15068), .A(n10871), .B(n10870), .ZN(
        P1_U3246) );
  XNOR2_X1 U13623 ( .A(n11177), .B(P2_REG1_REG_9__SCAN_IN), .ZN(n10877) );
  AOI21_X1 U13624 ( .B1(n10877), .B2(n10876), .A(n11169), .ZN(n10890) );
  NAND2_X1 U13625 ( .A1(n10878), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n10879) );
  NAND2_X1 U13626 ( .A1(n10880), .A2(n10879), .ZN(n10883) );
  INV_X1 U13627 ( .A(n10883), .ZN(n10885) );
  INV_X1 U13628 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n10881) );
  MUX2_X1 U13629 ( .A(P2_REG2_REG_9__SCAN_IN), .B(n10881), .S(n11177), .Z(
        n10884) );
  MUX2_X1 U13630 ( .A(n10881), .B(P2_REG2_REG_9__SCAN_IN), .S(n11177), .Z(
        n10882) );
  OAI21_X1 U13631 ( .B1(n10885), .B2(n10884), .A(n11179), .ZN(n10888) );
  INV_X1 U13632 ( .A(n15857), .ZN(n15864) );
  NOR2_X1 U13633 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9652), .ZN(n12194) );
  AOI21_X1 U13634 ( .B1(n15864), .B2(P2_ADDR_REG_9__SCAN_IN), .A(n12194), .ZN(
        n10886) );
  OAI21_X1 U13635 ( .B1(n11171), .B2(n15871), .A(n10886), .ZN(n10887) );
  AOI21_X1 U13636 ( .B1(n10888), .B2(n15866), .A(n10887), .ZN(n10889) );
  OAI21_X1 U13637 ( .B1(n10890), .B2(n15860), .A(n10889), .ZN(P2_U3223) );
  INV_X1 U13638 ( .A(n10891), .ZN(n10893) );
  INV_X1 U13639 ( .A(n13088), .ZN(n13084) );
  OAI222_X1 U13640 ( .A1(n13524), .A2(n10893), .B1(n13521), .B2(n10892), .C1(
        n13084), .C2(P3_U3151), .ZN(P3_U3279) );
  INV_X1 U13641 ( .A(n10896), .ZN(n10894) );
  NAND2_X1 U13642 ( .A1(n10894), .A2(P3_STATE_REG_SCAN_IN), .ZN(n12646) );
  NAND2_X1 U13643 ( .A1(n10895), .A2(n12646), .ZN(n10917) );
  NAND2_X1 U13644 ( .A1(n12626), .A2(n10896), .ZN(n10898) );
  NAND2_X1 U13645 ( .A1(n10898), .A2(n10897), .ZN(n10916) );
  INV_X1 U13646 ( .A(n10916), .ZN(n10899) );
  NAND2_X1 U13647 ( .A1(n10917), .A2(n10899), .ZN(n10908) );
  INV_X1 U13648 ( .A(P3_U3897), .ZN(n12943) );
  MUX2_X1 U13649 ( .A(n10908), .B(n12943), .S(n12641), .Z(n13129) );
  INV_X1 U13650 ( .A(P3_REG2_REG_2__SCAN_IN), .ZN(n11349) );
  XNOR2_X1 U13651 ( .A(n7298), .B(n11349), .ZN(n10907) );
  AND2_X1 U13652 ( .A1(n15919), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n10903) );
  OAI21_X1 U13653 ( .B1(n10921), .B2(n10903), .A(n10905), .ZN(n10904) );
  INV_X1 U13654 ( .A(n10904), .ZN(n12957) );
  NAND2_X1 U13655 ( .A1(n12957), .A2(P3_REG2_REG_1__SCAN_IN), .ZN(n12956) );
  NAND2_X1 U13656 ( .A1(n12956), .A2(n10905), .ZN(n10906) );
  OAI21_X1 U13657 ( .B1(n10907), .B2(n10906), .A(n10940), .ZN(n10937) );
  INV_X1 U13658 ( .A(n10908), .ZN(n10909) );
  INV_X1 U13659 ( .A(P3_REG1_REG_2__SCAN_IN), .ZN(n10926) );
  MUX2_X1 U13660 ( .A(P3_REG1_REG_2__SCAN_IN), .B(n10926), .S(n10944), .Z(
        n10914) );
  NAND2_X1 U13661 ( .A1(P3_REG1_REG_0__SCAN_IN), .A2(n15919), .ZN(n10910) );
  INV_X1 U13662 ( .A(P3_REG1_REG_0__SCAN_IN), .ZN(n11188) );
  NOR3_X1 U13663 ( .A1(n11188), .A2(P3_IR_REG_1__SCAN_IN), .A3(
        P3_IR_REG_0__SCAN_IN), .ZN(n10911) );
  NAND2_X1 U13664 ( .A1(n12959), .A2(P3_REG1_REG_1__SCAN_IN), .ZN(n12958) );
  INV_X1 U13665 ( .A(n10911), .ZN(n10912) );
  NAND2_X1 U13666 ( .A1(n12958), .A2(n10912), .ZN(n10913) );
  NAND2_X1 U13667 ( .A1(n10913), .A2(n10914), .ZN(n10946) );
  OAI21_X1 U13668 ( .B1(n10914), .B2(n10913), .A(n10946), .ZN(n10915) );
  NAND2_X1 U13669 ( .A1(n15915), .A2(n10915), .ZN(n10920) );
  INV_X1 U13670 ( .A(P3_REG3_REG_2__SCAN_IN), .ZN(n11340) );
  NOR2_X1 U13671 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11340), .ZN(n10918) );
  AOI21_X1 U13672 ( .B1(n15913), .B2(P3_ADDR_REG_2__SCAN_IN), .A(n10918), .ZN(
        n10919) );
  NAND2_X1 U13673 ( .A1(n10920), .A2(n10919), .ZN(n10936) );
  NOR2_X1 U13674 ( .A1(n10923), .A2(n12955), .ZN(n10924) );
  MUX2_X1 U13675 ( .A(P3_REG2_REG_0__SCAN_IN), .B(P3_REG1_REG_0__SCAN_IN), .S(
        n6527), .Z(n15918) );
  NOR2_X1 U13676 ( .A1(n15918), .A2(n15919), .ZN(n15917) );
  INV_X1 U13677 ( .A(n10925), .ZN(n10932) );
  MUX2_X1 U13678 ( .A(n11349), .B(n10926), .S(n6527), .Z(n10928) );
  NAND2_X1 U13679 ( .A1(n10928), .A2(n10927), .ZN(n10951) );
  INV_X1 U13680 ( .A(n10928), .ZN(n10929) );
  NAND2_X1 U13681 ( .A1(n10929), .A2(n7298), .ZN(n10930) );
  NAND2_X1 U13682 ( .A1(n10951), .A2(n10930), .ZN(n10931) );
  INV_X1 U13683 ( .A(n6730), .ZN(n10934) );
  NAND3_X1 U13684 ( .A1(n12962), .A2(n10932), .A3(n10931), .ZN(n10933) );
  AND2_X1 U13685 ( .A1(P3_U3897), .A2(n13515), .ZN(n15914) );
  AOI21_X1 U13686 ( .B1(n10934), .B2(n10933), .A(n13116), .ZN(n10935) );
  AOI211_X1 U13687 ( .C1(n15916), .C2(n10937), .A(n10936), .B(n10935), .ZN(
        n10938) );
  OAI21_X1 U13688 ( .B1(n7298), .B2(n13129), .A(n10938), .ZN(P3_U3184) );
  NAND2_X1 U13689 ( .A1(n7298), .A2(P3_REG2_REG_2__SCAN_IN), .ZN(n10939) );
  INV_X1 U13690 ( .A(P3_REG2_REG_3__SCAN_IN), .ZN(n10941) );
  NAND2_X1 U13691 ( .A1(n10942), .A2(n10941), .ZN(n10943) );
  NAND2_X1 U13692 ( .A1(n11064), .A2(n10943), .ZN(n10958) );
  NAND2_X1 U13693 ( .A1(n7298), .A2(P3_REG1_REG_2__SCAN_IN), .ZN(n10945) );
  INV_X1 U13694 ( .A(n10961), .ZN(n10947) );
  XNOR2_X1 U13695 ( .A(n10960), .B(P3_REG1_REG_3__SCAN_IN), .ZN(n10948) );
  NAND2_X1 U13696 ( .A1(n15915), .A2(n10948), .ZN(n10950) );
  AOI22_X1 U13697 ( .A1(n15913), .A2(P3_ADDR_REG_3__SCAN_IN), .B1(
        P3_REG3_REG_3__SCAN_IN), .B2(P3_U3151), .ZN(n10949) );
  NAND2_X1 U13698 ( .A1(n10950), .A2(n10949), .ZN(n10957) );
  INV_X1 U13699 ( .A(n10951), .ZN(n10954) );
  MUX2_X1 U13700 ( .A(P3_REG2_REG_3__SCAN_IN), .B(P3_REG1_REG_3__SCAN_IN), .S(
        n7233), .Z(n10952) );
  NOR2_X1 U13701 ( .A1(n10952), .A2(n10961), .ZN(n10975) );
  AOI21_X1 U13702 ( .B1(n10952), .B2(n10961), .A(n10975), .ZN(n10953) );
  OR3_X1 U13703 ( .A1(n6730), .A2(n10954), .A3(n10953), .ZN(n10955) );
  AOI21_X1 U13704 ( .B1(n11076), .B2(n10955), .A(n13116), .ZN(n10956) );
  AOI211_X1 U13705 ( .C1(n15916), .C2(n10958), .A(n10957), .B(n10956), .ZN(
        n10959) );
  OAI21_X1 U13706 ( .B1(n10961), .B2(n13129), .A(n10959), .ZN(P3_U3185) );
  MUX2_X1 U13707 ( .A(n15971), .B(P3_REG1_REG_6__SCAN_IN), .S(n11036), .Z(
        n10968) );
  NAND2_X1 U13708 ( .A1(n10962), .A2(n10961), .ZN(n10963) );
  MUX2_X1 U13709 ( .A(P3_REG1_REG_4__SCAN_IN), .B(n15966), .S(n10976), .Z(
        n11069) );
  INV_X1 U13710 ( .A(n10979), .ZN(n11109) );
  XNOR2_X1 U13711 ( .A(n10964), .B(n11109), .ZN(n11096) );
  NAND2_X1 U13712 ( .A1(n11096), .A2(P3_REG1_REG_5__SCAN_IN), .ZN(n10966) );
  NAND2_X1 U13713 ( .A1(n10964), .A2(n10979), .ZN(n10965) );
  NAND2_X1 U13714 ( .A1(n10966), .A2(n10965), .ZN(n10967) );
  NAND2_X1 U13715 ( .A1(n10967), .A2(n10968), .ZN(n11038) );
  OAI21_X1 U13716 ( .B1(n10968), .B2(n10967), .A(n11038), .ZN(n10989) );
  INV_X1 U13717 ( .A(P3_REG2_REG_4__SCAN_IN), .ZN(n11271) );
  XNOR2_X1 U13718 ( .A(n10976), .B(n11271), .ZN(n11062) );
  INV_X1 U13719 ( .A(P3_REG2_REG_5__SCAN_IN), .ZN(n11306) );
  INV_X1 U13720 ( .A(P3_REG2_REG_6__SCAN_IN), .ZN(n11442) );
  XNOR2_X1 U13721 ( .A(n11036), .B(n11442), .ZN(n10970) );
  AND3_X1 U13722 ( .A1(n11099), .A2(n10970), .A3(n10971), .ZN(n10972) );
  OAI21_X1 U13723 ( .B1(n10972), .B2(n6731), .A(n15916), .ZN(n10974) );
  AND2_X1 U13724 ( .A1(P3_U3151), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n11676) );
  AOI21_X1 U13725 ( .B1(n15913), .B2(P3_ADDR_REG_6__SCAN_IN), .A(n11676), .ZN(
        n10973) );
  OAI211_X1 U13726 ( .C1(n13129), .C2(n11046), .A(n10974), .B(n10973), .ZN(
        n10988) );
  INV_X1 U13727 ( .A(n10975), .ZN(n11075) );
  MUX2_X1 U13728 ( .A(n11271), .B(n15966), .S(n7233), .Z(n10977) );
  INV_X1 U13729 ( .A(n10976), .ZN(n11081) );
  NAND2_X1 U13730 ( .A1(n10977), .A2(n11081), .ZN(n10978) );
  OAI21_X1 U13731 ( .B1(n10977), .B2(n11081), .A(n10978), .ZN(n11074) );
  INV_X1 U13732 ( .A(n10978), .ZN(n11103) );
  MUX2_X1 U13733 ( .A(P3_REG2_REG_5__SCAN_IN), .B(P3_REG1_REG_5__SCAN_IN), .S(
        n6527), .Z(n10980) );
  NOR2_X1 U13734 ( .A1(n10980), .A2(n10979), .ZN(n10981) );
  AOI21_X1 U13735 ( .B1(n10980), .B2(n10979), .A(n10981), .ZN(n11102) );
  INV_X1 U13736 ( .A(n10981), .ZN(n10984) );
  MUX2_X1 U13737 ( .A(n11442), .B(n15971), .S(n6527), .Z(n10982) );
  NAND2_X1 U13738 ( .A1(n10982), .A2(n11036), .ZN(n11039) );
  OAI21_X1 U13739 ( .B1(n10982), .B2(n11036), .A(n11039), .ZN(n10983) );
  INV_X1 U13740 ( .A(n11043), .ZN(n10986) );
  NAND3_X1 U13741 ( .A1(n11106), .A2(n10984), .A3(n10983), .ZN(n10985) );
  AOI21_X1 U13742 ( .B1(n10986), .B2(n10985), .A(n13116), .ZN(n10987) );
  AOI211_X1 U13743 ( .C1(n15915), .C2(n10989), .A(n10988), .B(n10987), .ZN(
        n10990) );
  INV_X1 U13744 ( .A(n10990), .ZN(P3_U3188) );
  XNOR2_X1 U13745 ( .A(n11083), .B(n11089), .ZN(n10995) );
  XNOR2_X1 U13746 ( .A(n12832), .B(n11365), .ZN(n10991) );
  NAND2_X1 U13747 ( .A1(n10991), .A2(n11343), .ZN(n10992) );
  NAND2_X1 U13748 ( .A1(n10993), .A2(n10992), .ZN(n10994) );
  NAND2_X1 U13749 ( .A1(n10994), .A2(n10995), .ZN(n11088) );
  OAI21_X1 U13750 ( .B1(n10995), .B2(n10994), .A(n11085), .ZN(n10996) );
  NAND2_X1 U13751 ( .A1(n10996), .A2(n12924), .ZN(n11000) );
  INV_X1 U13752 ( .A(n11339), .ZN(n10998) );
  INV_X1 U13753 ( .A(n12952), .ZN(n11342) );
  OAI22_X1 U13754 ( .A1(n12917), .A2(n11343), .B1(n11342), .B2(n12931), .ZN(
        n10997) );
  AOI21_X1 U13755 ( .B1(n10998), .B2(n12919), .A(n10997), .ZN(n10999) );
  OAI211_X1 U13756 ( .C1(n11001), .C2(n11340), .A(n11000), .B(n10999), .ZN(
        P3_U3177) );
  AND2_X1 U13757 ( .A1(n13810), .A2(n14307), .ZN(n11408) );
  INV_X1 U13758 ( .A(n11408), .ZN(n11411) );
  INV_X1 U13759 ( .A(n6528), .ZN(n11004) );
  XNOR2_X1 U13760 ( .A(n11004), .B(n11408), .ZN(n11122) );
  OR2_X1 U13761 ( .A1(n11121), .A2(n14261), .ZN(n11413) );
  NOR2_X1 U13762 ( .A1(n11122), .A2(n11409), .ZN(n11114) );
  AOI21_X1 U13763 ( .B1(n6528), .B2(n11411), .A(n11114), .ZN(n11035) );
  OR2_X1 U13764 ( .A1(n15881), .A2(n11321), .ZN(n11005) );
  NOR2_X1 U13765 ( .A1(n11006), .A2(n11005), .ZN(n11017) );
  NAND2_X1 U13766 ( .A1(n11017), .A2(n15882), .ZN(n11013) );
  OR2_X1 U13767 ( .A1(n14387), .A2(n11007), .ZN(n11008) );
  NAND2_X1 U13768 ( .A1(n13809), .A2(n14307), .ZN(n11415) );
  XNOR2_X1 U13769 ( .A(n11415), .B(n11414), .ZN(n11030) );
  INV_X1 U13770 ( .A(n11030), .ZN(n11009) );
  NAND2_X1 U13771 ( .A1(n13766), .A2(n11009), .ZN(n11034) );
  AND2_X1 U13772 ( .A1(n11126), .A2(n11010), .ZN(n11329) );
  INV_X1 U13773 ( .A(n11329), .ZN(n11011) );
  OR2_X1 U13774 ( .A1(n11013), .A2(n11011), .ZN(n11012) );
  INV_X1 U13775 ( .A(n11013), .ZN(n11016) );
  INV_X1 U13776 ( .A(n11014), .ZN(n11015) );
  AOI22_X1 U13777 ( .A1(n13769), .A2(n13810), .B1(n13808), .B2(n13770), .ZN(
        n11256) );
  INV_X1 U13778 ( .A(n11017), .ZN(n11019) );
  NAND2_X1 U13779 ( .A1(n11019), .A2(n11018), .ZN(n11025) );
  NAND2_X1 U13780 ( .A1(n11021), .A2(n11020), .ZN(n11022) );
  NOR2_X1 U13781 ( .A1(n11023), .A2(n11022), .ZN(n11024) );
  NAND2_X1 U13782 ( .A1(n11025), .A2(n11024), .ZN(n11426) );
  NOR2_X1 U13783 ( .A1(n11426), .A2(P2_U3088), .ZN(n11118) );
  INV_X1 U13784 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n11026) );
  OAI22_X1 U13785 ( .A1(n13759), .A2(n11256), .B1(n11118), .B2(n11026), .ZN(
        n11027) );
  AOI21_X1 U13786 ( .B1(n9522), .B2(n13777), .A(n11027), .ZN(n11033) );
  NAND2_X1 U13787 ( .A1(n13766), .A2(n15891), .ZN(n13751) );
  INV_X1 U13788 ( .A(n13810), .ZN(n11028) );
  OAI22_X1 U13789 ( .A1(n13751), .A2(n11028), .B1(n6528), .B2(n13736), .ZN(
        n11031) );
  INV_X1 U13790 ( .A(n11114), .ZN(n11029) );
  NAND3_X1 U13791 ( .A1(n11031), .A2(n11030), .A3(n11029), .ZN(n11032) );
  OAI211_X1 U13792 ( .C1(n11035), .C2(n11034), .A(n11033), .B(n11032), .ZN(
        P2_U3209) );
  OR2_X1 U13793 ( .A1(n11036), .A2(n15971), .ZN(n11037) );
  INV_X1 U13794 ( .A(n11192), .ZN(n11047) );
  XOR2_X1 U13795 ( .A(n11191), .B(P3_REG1_REG_7__SCAN_IN), .Z(n11054) );
  INV_X1 U13796 ( .A(n11039), .ZN(n11042) );
  MUX2_X1 U13797 ( .A(P3_REG2_REG_7__SCAN_IN), .B(P3_REG1_REG_7__SCAN_IN), .S(
        n7233), .Z(n11040) );
  AOI21_X1 U13798 ( .B1(n11040), .B2(n11192), .A(n11201), .ZN(n11041) );
  INV_X1 U13799 ( .A(n11205), .ZN(n11045) );
  NOR3_X1 U13800 ( .A1(n11043), .A2(n11042), .A3(n11041), .ZN(n11044) );
  OAI21_X1 U13801 ( .B1(n11045), .B2(n11044), .A(n15914), .ZN(n11053) );
  NOR2_X1 U13802 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n8230), .ZN(n11763) );
  AOI21_X1 U13803 ( .B1(n15913), .B2(P3_ADDR_REG_7__SCAN_IN), .A(n11763), .ZN(
        n11049) );
  OAI21_X1 U13804 ( .B1(n13129), .B2(n11192), .A(n11049), .ZN(n11050) );
  AOI21_X1 U13805 ( .B1(n11051), .B2(n15916), .A(n11050), .ZN(n11052) );
  OAI211_X1 U13806 ( .C1(n11054), .C2(n13118), .A(n11053), .B(n11052), .ZN(
        P3_U3189) );
  OAI222_X1 U13807 ( .A1(n13524), .A2(n11056), .B1(n13521), .B2(n11055), .C1(
        n13112), .C2(P3_U3151), .ZN(P3_U3278) );
  AOI21_X1 U13808 ( .B1(n13766), .B2(n11413), .A(n13777), .ZN(n11061) );
  INV_X1 U13809 ( .A(n11118), .ZN(n11058) );
  NAND2_X1 U13810 ( .A1(n13810), .A2(n13770), .ZN(n11128) );
  INV_X1 U13811 ( .A(n11128), .ZN(n11057) );
  AOI22_X1 U13812 ( .A1(n11058), .A2(P2_REG3_REG_0__SCAN_IN), .B1(n13773), 
        .B2(n11057), .ZN(n11060) );
  NAND3_X1 U13813 ( .A1(n13765), .A2(n13812), .A3(n11121), .ZN(n11059) );
  OAI211_X1 U13814 ( .C1(n11061), .C2(n10196), .A(n11060), .B(n11059), .ZN(
        P2_U3204) );
  NAND3_X1 U13815 ( .A1(n11064), .A2(n7661), .A3(n11063), .ZN(n11065) );
  AND2_X1 U13816 ( .A1(n11066), .A2(n11065), .ZN(n11073) );
  OAI21_X1 U13817 ( .B1(n11069), .B2(n11068), .A(n11067), .ZN(n11070) );
  NAND2_X1 U13818 ( .A1(n15915), .A2(n11070), .ZN(n11072) );
  AND2_X1 U13819 ( .A1(P3_U3151), .A2(P3_REG3_REG_4__SCAN_IN), .ZN(n11227) );
  AOI21_X1 U13820 ( .B1(n15913), .B2(P3_ADDR_REG_4__SCAN_IN), .A(n11227), .ZN(
        n11071) );
  OAI211_X1 U13821 ( .C1(n11073), .C2(n13141), .A(n11072), .B(n11071), .ZN(
        n11080) );
  INV_X1 U13822 ( .A(n11104), .ZN(n11078) );
  NAND3_X1 U13823 ( .A1(n11076), .A2(n11075), .A3(n11074), .ZN(n11077) );
  AOI21_X1 U13824 ( .B1(n11078), .B2(n11077), .A(n13116), .ZN(n11079) );
  AOI211_X1 U13825 ( .C1(n15922), .C2(n11081), .A(n11080), .B(n11079), .ZN(
        n11082) );
  INV_X1 U13826 ( .A(n11082), .ZN(P3_U3186) );
  INV_X1 U13827 ( .A(n11083), .ZN(n11084) );
  NAND2_X1 U13828 ( .A1(n11084), .A2(n11089), .ZN(n11086) );
  AOI21_X1 U13829 ( .B1(n11085), .B2(n11086), .A(n11087), .ZN(n11095) );
  NAND2_X1 U13830 ( .A1(n11219), .A2(n12924), .ZN(n11094) );
  INV_X1 U13831 ( .A(n12344), .ZN(n11456) );
  OAI22_X1 U13832 ( .A1(n12917), .A2(n11089), .B1(n11456), .B2(n12931), .ZN(
        n11092) );
  MUX2_X1 U13833 ( .A(P3_U3151), .B(n12934), .S(n12350), .Z(n11091) );
  AOI211_X1 U13834 ( .C1(n12919), .C2(n12351), .A(n11092), .B(n11091), .ZN(
        n11093) );
  OAI21_X1 U13835 ( .B1(n11095), .B2(n11094), .A(n11093), .ZN(P3_U3158) );
  XOR2_X1 U13836 ( .A(n11096), .B(P3_REG1_REG_5__SCAN_IN), .Z(n11111) );
  NAND2_X1 U13837 ( .A1(n11097), .A2(n11306), .ZN(n11098) );
  AND2_X1 U13838 ( .A1(n11099), .A2(n11098), .ZN(n11101) );
  AND2_X1 U13839 ( .A1(P3_U3151), .A2(P3_REG3_REG_5__SCAN_IN), .ZN(n11458) );
  AOI21_X1 U13840 ( .B1(n15913), .B2(P3_ADDR_REG_5__SCAN_IN), .A(n11458), .ZN(
        n11100) );
  OAI21_X1 U13841 ( .B1(n11101), .B2(n13141), .A(n11100), .ZN(n11108) );
  OR3_X1 U13842 ( .A1(n11104), .A2(n11103), .A3(n11102), .ZN(n11105) );
  AOI21_X1 U13843 ( .B1(n11106), .B2(n11105), .A(n13116), .ZN(n11107) );
  AOI211_X1 U13844 ( .C1(n15922), .C2(n11109), .A(n11108), .B(n11107), .ZN(
        n11110) );
  OAI21_X1 U13845 ( .B1(n11111), .B2(n13118), .A(n11110), .ZN(P3_U3187) );
  INV_X1 U13846 ( .A(n11112), .ZN(n11144) );
  AOI22_X1 U13847 ( .A1(n15732), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(n15527), .ZN(n11113) );
  OAI21_X1 U13848 ( .B1(n11144), .B2(n15549), .A(n11113), .ZN(P1_U3343) );
  INV_X1 U13849 ( .A(n11412), .ZN(n11115) );
  AOI21_X1 U13850 ( .B1(n11122), .B2(n11115), .A(n11114), .ZN(n11125) );
  INV_X1 U13851 ( .A(n13812), .ZN(n11117) );
  INV_X1 U13852 ( .A(n13809), .ZN(n11116) );
  OAI22_X1 U13853 ( .A1(n11117), .A2(n13741), .B1(n11116), .B2(n13743), .ZN(
        n11139) );
  INV_X1 U13854 ( .A(n11139), .ZN(n11119) );
  INV_X1 U13855 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n13813) );
  OAI22_X1 U13856 ( .A1(n13759), .A2(n11119), .B1(n11118), .B2(n13813), .ZN(
        n11120) );
  AOI21_X1 U13857 ( .B1(n7675), .B2(n13777), .A(n11120), .ZN(n11124) );
  INV_X1 U13858 ( .A(n11121), .ZN(n11136) );
  NAND3_X1 U13859 ( .A1(n13765), .A2(n11136), .A3(n11122), .ZN(n11123) );
  OAI211_X1 U13860 ( .C1(n11125), .C2(n13736), .A(n11124), .B(n11123), .ZN(
        P2_U3194) );
  INV_X1 U13861 ( .A(n14303), .ZN(n15905) );
  INV_X1 U13862 ( .A(n11126), .ZN(n11127) );
  NOR2_X1 U13863 ( .A1(n10196), .A2(n11127), .ZN(n11130) );
  INV_X1 U13864 ( .A(n11003), .ZN(n14185) );
  OAI21_X1 U13865 ( .B1(n14185), .B2(n14270), .A(n11352), .ZN(n11129) );
  NAND2_X1 U13866 ( .A1(n11129), .A2(n11128), .ZN(n11359) );
  AOI211_X1 U13867 ( .C1(n15905), .C2(n11352), .A(n11130), .B(n11359), .ZN(
        n15887) );
  INV_X1 U13868 ( .A(n15881), .ZN(n11131) );
  NAND2_X1 U13869 ( .A1(n15910), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n11133) );
  OAI21_X1 U13870 ( .B1(n15887), .B2(n15910), .A(n11133), .ZN(P2_U3499) );
  INV_X1 U13871 ( .A(n11134), .ZN(n11135) );
  AOI21_X1 U13872 ( .B1(n11136), .B2(n11138), .A(n11135), .ZN(n11335) );
  XNOR2_X1 U13873 ( .A(n11138), .B(n11137), .ZN(n11140) );
  AOI21_X1 U13874 ( .B1(n11140), .B2(n14270), .A(n11139), .ZN(n11327) );
  OAI211_X1 U13875 ( .C1(n10196), .C2(n11296), .A(n14261), .B(n11252), .ZN(
        n11331) );
  OAI211_X1 U13876 ( .C1(n11335), .C2(n14391), .A(n11327), .B(n11331), .ZN(
        n11298) );
  NAND2_X1 U13877 ( .A1(n15912), .A2(n14387), .ZN(n14349) );
  OAI22_X1 U13878 ( .A1(n14349), .A2(n11296), .B1(n15912), .B2(n10564), .ZN(
        n11141) );
  AOI21_X1 U13879 ( .B1(n11298), .B2(n15912), .A(n11141), .ZN(n11142) );
  INV_X1 U13880 ( .A(n11142), .ZN(P2_U3500) );
  INV_X1 U13881 ( .A(n12305), .ZN(n11143) );
  OAI222_X1 U13882 ( .A1(n14472), .A2(n11145), .B1(n14461), .B2(n11144), .C1(
        P2_U3088), .C2(n11143), .ZN(P2_U3315) );
  MUX2_X1 U13883 ( .A(P1_REG1_REG_8__SCAN_IN), .B(n11147), .S(n15030), .Z(
        n15021) );
  NAND2_X1 U13884 ( .A1(n15022), .A2(n15021), .ZN(n15020) );
  OAI21_X1 U13885 ( .B1(P1_REG1_REG_8__SCAN_IN), .B2(n15030), .A(n15020), .ZN(
        n11238) );
  XNOR2_X1 U13886 ( .A(n11231), .B(n12258), .ZN(n11237) );
  XNOR2_X1 U13887 ( .A(n11238), .B(n11237), .ZN(n11160) );
  NAND2_X1 U13888 ( .A1(n11148), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n15026) );
  NAND2_X1 U13889 ( .A1(n15027), .A2(n15026), .ZN(n11150) );
  MUX2_X1 U13890 ( .A(P1_REG2_REG_8__SCAN_IN), .B(n11906), .S(n15030), .Z(
        n11149) );
  NAND2_X1 U13891 ( .A1(n11150), .A2(n11149), .ZN(n15029) );
  NAND2_X1 U13892 ( .A1(n15030), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n11155) );
  NAND2_X1 U13893 ( .A1(n15029), .A2(n11155), .ZN(n11153) );
  MUX2_X1 U13894 ( .A(P1_REG2_REG_9__SCAN_IN), .B(n11151), .S(n11231), .Z(
        n11152) );
  NAND2_X1 U13895 ( .A1(n11153), .A2(n11152), .ZN(n11234) );
  MUX2_X1 U13896 ( .A(n11151), .B(P1_REG2_REG_9__SCAN_IN), .S(n11231), .Z(
        n11154) );
  NAND3_X1 U13897 ( .A1(n15029), .A2(n11155), .A3(n11154), .ZN(n11156) );
  NAND3_X1 U13898 ( .A1(n15746), .A2(n11234), .A3(n11156), .ZN(n11158) );
  AND2_X1 U13899 ( .A1(P1_U3086), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n14620) );
  AOI21_X1 U13900 ( .B1(n15722), .B2(P1_ADDR_REG_9__SCAN_IN), .A(n14620), .ZN(
        n11157) );
  OAI211_X1 U13901 ( .C1(n15068), .C2(n11236), .A(n11158), .B(n11157), .ZN(
        n11159) );
  AOI21_X1 U13902 ( .B1(n11160), .B2(n15745), .A(n11159), .ZN(n11161) );
  INV_X1 U13903 ( .A(n11161), .ZN(P1_U3252) );
  XOR2_X1 U13904 ( .A(n11163), .B(n11162), .Z(n11168) );
  INV_X1 U13905 ( .A(n10283), .ZN(n11377) );
  INV_X1 U13906 ( .A(n14709), .ZN(n14971) );
  AOI22_X1 U13907 ( .A1(n14667), .A2(n14971), .B1(P1_REG3_REG_1__SCAN_IN), 
        .B2(n11316), .ZN(n11164) );
  OAI21_X1 U13908 ( .B1(n11377), .B2(n14681), .A(n11164), .ZN(n11165) );
  AOI21_X1 U13909 ( .B1(n14684), .B2(n11166), .A(n11165), .ZN(n11167) );
  OAI21_X1 U13910 ( .B1(n11168), .B2(n14686), .A(n11167), .ZN(P1_U3222) );
  XOR2_X1 U13911 ( .A(P2_REG1_REG_10__SCAN_IN), .B(n11655), .Z(n11172) );
  OAI21_X1 U13912 ( .B1(n11173), .B2(n11172), .A(n15830), .ZN(n11186) );
  INV_X1 U13913 ( .A(n11174), .ZN(n13601) );
  NOR2_X1 U13914 ( .A1(n15871), .A2(n11175), .ZN(n11176) );
  AOI211_X1 U13915 ( .C1(n15864), .C2(P2_ADDR_REG_10__SCAN_IN), .A(n13601), 
        .B(n11176), .ZN(n11185) );
  OR2_X1 U13916 ( .A1(n11177), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n11178) );
  INV_X1 U13917 ( .A(n11181), .ZN(n11183) );
  MUX2_X1 U13918 ( .A(P2_REG2_REG_10__SCAN_IN), .B(n14230), .S(n11655), .Z(
        n11182) );
  MUX2_X1 U13919 ( .A(n14230), .B(P2_REG2_REG_10__SCAN_IN), .S(n11655), .Z(
        n11180) );
  OAI211_X1 U13920 ( .C1(n11183), .C2(n11182), .A(n15866), .B(n11649), .ZN(
        n11184) );
  OAI211_X1 U13921 ( .C1(n11186), .C2(n11654), .A(n11185), .B(n11184), .ZN(
        P2_U3224) );
  MUX2_X1 U13922 ( .A(n11188), .B(n11187), .S(n15973), .Z(n11189) );
  OAI21_X1 U13923 ( .B1(n13403), .B2(n11190), .A(n11189), .ZN(P3_U3459) );
  XNOR2_X1 U13924 ( .A(n11574), .B(P3_REG1_REG_8__SCAN_IN), .ZN(n11571) );
  NAND2_X1 U13925 ( .A1(n11193), .A2(n11192), .ZN(n11194) );
  XOR2_X1 U13926 ( .A(n11571), .B(n11572), .Z(n11209) );
  INV_X1 U13927 ( .A(P3_ADDR_REG_8__SCAN_IN), .ZN(n11195) );
  NAND2_X1 U13928 ( .A1(P3_U3151), .A2(P3_REG3_REG_8__SCAN_IN), .ZN(n11971) );
  OAI21_X1 U13929 ( .B1(n15925), .B2(n11195), .A(n11971), .ZN(n11200) );
  INV_X1 U13930 ( .A(P3_REG2_REG_8__SCAN_IN), .ZN(n11534) );
  XNOR2_X1 U13931 ( .A(n11574), .B(n11534), .ZN(n11196) );
  NAND3_X1 U13932 ( .A1(n11197), .A2(n11196), .A3(n6689), .ZN(n11198) );
  AOI21_X1 U13933 ( .B1(n6727), .B2(n11198), .A(n13141), .ZN(n11199) );
  AOI211_X1 U13934 ( .C1(n15922), .C2(n11574), .A(n11200), .B(n11199), .ZN(
        n11208) );
  INV_X1 U13935 ( .A(n11201), .ZN(n11204) );
  INV_X1 U13936 ( .A(P3_REG1_REG_8__SCAN_IN), .ZN(n11573) );
  MUX2_X1 U13937 ( .A(n11534), .B(n11573), .S(n6527), .Z(n11202) );
  NAND2_X1 U13938 ( .A1(n11202), .A2(n11574), .ZN(n11581) );
  OAI21_X1 U13939 ( .B1(n11202), .B2(n11574), .A(n11581), .ZN(n11203) );
  AND3_X1 U13940 ( .A1(n11205), .A2(n11204), .A3(n11203), .ZN(n11206) );
  OAI21_X1 U13941 ( .B1(n11585), .B2(n11206), .A(n15914), .ZN(n11207) );
  OAI211_X1 U13942 ( .C1(n11209), .C2(n13118), .A(n11208), .B(n11207), .ZN(
        P3_U3190) );
  AND2_X1 U13943 ( .A1(n10283), .A2(n11371), .ZN(n14707) );
  OR2_X1 U13944 ( .A1(n14707), .A2(n11212), .ZN(n14921) );
  NAND2_X1 U13945 ( .A1(n15492), .A2(n15465), .ZN(n11213) );
  AOI22_X1 U13946 ( .A1(n14921), .A2(n11213), .B1(n15801), .B2(n10855), .ZN(
        n11500) );
  NAND3_X1 U13947 ( .A1(n11497), .A2(n9194), .A3(n14688), .ZN(n11214) );
  NAND2_X1 U13948 ( .A1(n11500), .A2(n11214), .ZN(n15502) );
  NAND2_X1 U13949 ( .A1(n15502), .A2(n15815), .ZN(n11215) );
  OAI21_X1 U13950 ( .B1(n15815), .B2(n8651), .A(n11215), .ZN(P1_U3459) );
  INV_X1 U13951 ( .A(n11272), .ZN(n11230) );
  INV_X1 U13952 ( .A(n12934), .ZN(n11679) );
  INV_X1 U13953 ( .A(n11216), .ZN(n11217) );
  NAND2_X1 U13954 ( .A1(n11217), .A2(n12952), .ZN(n11218) );
  XNOR2_X1 U13955 ( .A(n12832), .B(n11273), .ZN(n11220) );
  NAND2_X1 U13956 ( .A1(n11220), .A2(n11456), .ZN(n11451) );
  INV_X1 U13957 ( .A(n11220), .ZN(n11221) );
  NAND2_X1 U13958 ( .A1(n11221), .A2(n12344), .ZN(n11222) );
  OAI21_X1 U13959 ( .B1(n11224), .B2(n11223), .A(n11452), .ZN(n11225) );
  NAND2_X1 U13960 ( .A1(n11225), .A2(n12924), .ZN(n11229) );
  OAI22_X1 U13961 ( .A1(n12937), .A2(n15939), .B1(n12931), .B2(n11670), .ZN(
        n11226) );
  AOI211_X1 U13962 ( .C1(n12929), .C2(n12952), .A(n11227), .B(n11226), .ZN(
        n11228) );
  OAI211_X1 U13963 ( .C1(n11230), .C2(n11679), .A(n11229), .B(n11228), .ZN(
        P3_U3170) );
  NAND2_X1 U13964 ( .A1(n11231), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n11233) );
  MUX2_X1 U13965 ( .A(n8835), .B(P1_REG2_REG_10__SCAN_IN), .S(n11239), .Z(
        n11232) );
  AOI21_X1 U13966 ( .B1(n11234), .B2(n11233), .A(n11232), .ZN(n11486) );
  NAND3_X1 U13967 ( .A1(n11234), .A2(n11233), .A3(n11232), .ZN(n11235) );
  NAND2_X1 U13968 ( .A1(n15746), .A2(n11235), .ZN(n11246) );
  XOR2_X1 U13969 ( .A(P1_REG1_REG_10__SCAN_IN), .B(n11239), .Z(n11240) );
  OAI211_X1 U13970 ( .C1(n11241), .C2(n11240), .A(n11477), .B(n15745), .ZN(
        n11245) );
  AND2_X1 U13971 ( .A1(P1_U3086), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n11243) );
  NOR2_X1 U13972 ( .A1(n15068), .A2(n11482), .ZN(n11242) );
  AOI211_X1 U13973 ( .C1(n15722), .C2(P1_ADDR_REG_10__SCAN_IN), .A(n11243), 
        .B(n11242), .ZN(n11244) );
  OAI211_X1 U13974 ( .C1(n11486), .C2(n11246), .A(n11245), .B(n11244), .ZN(
        P1_U3253) );
  INV_X1 U13975 ( .A(n11247), .ZN(n11249) );
  INV_X1 U13976 ( .A(n15849), .ZN(n12299) );
  OAI222_X1 U13977 ( .A1(n14472), .A2(n11248), .B1(n14474), .B2(n11249), .C1(
        n12299), .C2(P2_U3088), .ZN(P2_U3314) );
  INV_X1 U13978 ( .A(n12136), .ZN(n11992) );
  OAI222_X1 U13979 ( .A1(n15539), .A2(n11250), .B1(n15549), .B2(n11249), .C1(
        n11992), .C2(P1_U3086), .ZN(P1_U3342) );
  INV_X1 U13980 ( .A(n11251), .ZN(n11254) );
  NAND2_X1 U13981 ( .A1(n11464), .A2(n11254), .ZN(n11555) );
  OAI21_X1 U13982 ( .B1(n11464), .B2(n11254), .A(n11555), .ZN(n11682) );
  AOI21_X1 U13983 ( .B1(n11252), .B2(n9522), .A(n15891), .ZN(n11253) );
  AND2_X1 U13984 ( .A1(n11565), .A2(n11253), .ZN(n11683) );
  XNOR2_X1 U13985 ( .A(n11255), .B(n11254), .ZN(n11257) );
  OAI21_X1 U13986 ( .B1(n11257), .B2(n14127), .A(n11256), .ZN(n11681) );
  AOI211_X1 U13987 ( .C1(n14396), .C2(n11682), .A(n11683), .B(n11681), .ZN(
        n11264) );
  INV_X1 U13988 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n11258) );
  OAI22_X1 U13989 ( .A1(n14430), .A2(n11684), .B1(n15908), .B2(n11258), .ZN(
        n11259) );
  INV_X1 U13990 ( .A(n11259), .ZN(n11260) );
  OAI21_X1 U13991 ( .B1(n11264), .B2(n15906), .A(n11260), .ZN(P2_U3436) );
  OAI22_X1 U13992 ( .A1(n14349), .A2(n11684), .B1(n15912), .B2(n11261), .ZN(
        n11262) );
  INV_X1 U13993 ( .A(n11262), .ZN(n11263) );
  OAI21_X1 U13994 ( .B1(n11264), .B2(n15910), .A(n11263), .ZN(P2_U3501) );
  INV_X1 U13995 ( .A(n12446), .ZN(n12347) );
  NAND2_X1 U13996 ( .A1(n11265), .A2(n12347), .ZN(n12349) );
  NAND2_X1 U13997 ( .A1(n12349), .A2(n12512), .ZN(n11266) );
  XNOR2_X1 U13998 ( .A(n11266), .B(n12511), .ZN(n15940) );
  NOR2_X1 U13999 ( .A1(n12340), .A2(n12347), .ZN(n12343) );
  NOR2_X1 U14000 ( .A1(n12343), .A2(n11267), .ZN(n11268) );
  XNOR2_X1 U14001 ( .A(n11268), .B(n12511), .ZN(n11270) );
  OAI22_X1 U14002 ( .A1(n11342), .A2(n13265), .B1(n11670), .B2(n13267), .ZN(
        n11269) );
  AOI21_X1 U14003 ( .B1(n11270), .B2(n13336), .A(n11269), .ZN(n15941) );
  MUX2_X1 U14004 ( .A(n11271), .B(n15941), .S(n13350), .Z(n11275) );
  AOI22_X1 U14005 ( .A1(n13310), .A2(n11273), .B1(n13345), .B2(n11272), .ZN(
        n11274) );
  OAI211_X1 U14006 ( .C1(n13352), .C2(n15940), .A(n11275), .B(n11274), .ZN(
        P3_U3229) );
  INV_X1 U14007 ( .A(n11276), .ZN(n11278) );
  OAI222_X1 U14008 ( .A1(n13524), .A2(n11278), .B1(n13521), .B2(n11277), .C1(
        n7334), .C2(P3_U3151), .ZN(P3_U3277) );
  NAND2_X1 U14009 ( .A1(n11280), .A2(n14926), .ZN(n11738) );
  OAI21_X1 U14010 ( .B1(n11280), .B2(n14926), .A(n11738), .ZN(n11721) );
  NAND2_X1 U14011 ( .A1(n11282), .A2(n14926), .ZN(n11729) );
  NAND3_X1 U14012 ( .A1(n11281), .A2(n15807), .A3(n11729), .ZN(n11286) );
  AOI22_X1 U14013 ( .A1(n14969), .A2(n15801), .B1(n15798), .B2(n10309), .ZN(
        n11285) );
  OAI211_X1 U14014 ( .C1(n11512), .C2(n11283), .A(n15447), .B(n11733), .ZN(
        n11722) );
  NAND2_X1 U14015 ( .A1(n7945), .A2(n15701), .ZN(n11284) );
  NAND4_X1 U14016 ( .A1(n11286), .A2(n11285), .A3(n11722), .A4(n11284), .ZN(
        n11287) );
  AOI21_X1 U14017 ( .B1(n15812), .B2(n11721), .A(n11287), .ZN(n11290) );
  NAND2_X1 U14018 ( .A1(n15820), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n11288) );
  OAI21_X1 U14019 ( .B1(n11290), .B2(n15820), .A(n11288), .ZN(P1_U3532) );
  OR2_X1 U14020 ( .A1(n15815), .A2(n8712), .ZN(n11289) );
  OAI21_X1 U14021 ( .B1(n11290), .B2(n15813), .A(n11289), .ZN(P1_U3471) );
  INV_X1 U14022 ( .A(n11291), .ZN(n11293) );
  OAI222_X1 U14023 ( .A1(n14472), .A2(n11292), .B1(n14474), .B2(n11293), .C1(
        n13916), .C2(P2_U3088), .ZN(P2_U3311) );
  INV_X1 U14024 ( .A(n15059), .ZN(n15053) );
  OAI222_X1 U14025 ( .A1(n15546), .A2(n11294), .B1(n15549), .B2(n11293), .C1(
        n15053), .C2(P1_U3086), .ZN(P1_U3339) );
  INV_X1 U14026 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n11295) );
  OAI22_X1 U14027 ( .A1(n14430), .A2(n11296), .B1(n15908), .B2(n11295), .ZN(
        n11297) );
  AOI21_X1 U14028 ( .B1(n11298), .B2(n15908), .A(n11297), .ZN(n11299) );
  INV_X1 U14029 ( .A(n11299), .ZN(P2_U3433) );
  XNOR2_X1 U14030 ( .A(n11300), .B(n12521), .ZN(n15948) );
  OAI21_X1 U14031 ( .B1(n12340), .B2(n11302), .A(n11301), .ZN(n11304) );
  XNOR2_X1 U14032 ( .A(n11304), .B(n11303), .ZN(n11305) );
  AOI222_X1 U14033 ( .A1(n13336), .A2(n11305), .B1(n12950), .B2(n13340), .C1(
        n12344), .C2(n13339), .ZN(n15949) );
  MUX2_X1 U14034 ( .A(n11306), .B(n15949), .S(n13350), .Z(n11309) );
  INV_X1 U14035 ( .A(n15947), .ZN(n11307) );
  AOI22_X1 U14036 ( .A1(n13310), .A2(n11307), .B1(n13345), .B2(n11450), .ZN(
        n11308) );
  OAI211_X1 U14037 ( .C1(n13352), .C2(n15948), .A(n11309), .B(n11308), .ZN(
        P3_U3228) );
  OAI22_X1 U14038 ( .A1(n13403), .A2(n11310), .B1(n15973), .B2(n7495), .ZN(
        n11311) );
  INV_X1 U14039 ( .A(n11311), .ZN(n11312) );
  OAI21_X1 U14040 ( .B1(n11313), .B2(n15970), .A(n11312), .ZN(P3_U3460) );
  XOR2_X1 U14041 ( .A(n11315), .B(n11314), .Z(n11320) );
  INV_X1 U14042 ( .A(n14681), .ZN(n14591) );
  AOI22_X1 U14043 ( .A1(n14591), .A2(n10855), .B1(P1_REG3_REG_2__SCAN_IN), 
        .B2(n11316), .ZN(n11317) );
  OAI21_X1 U14044 ( .B1(n14695), .B2(n14680), .A(n11317), .ZN(n11318) );
  AOI21_X1 U14045 ( .B1(n14684), .B2(n14708), .A(n11318), .ZN(n11319) );
  OAI21_X1 U14046 ( .B1(n11320), .B2(n14686), .A(n11319), .ZN(P1_U3237) );
  INV_X1 U14047 ( .A(n11321), .ZN(n11322) );
  AND3_X1 U14048 ( .A1(n11322), .A2(n15882), .A3(n15881), .ZN(n11323) );
  NAND2_X1 U14049 ( .A1(n11324), .A2(n11323), .ZN(n11330) );
  NAND2_X1 U14050 ( .A1(n11003), .A2(n14164), .ZN(n11325) );
  AND2_X1 U14051 ( .A1(n13615), .A2(n11325), .ZN(n11326) );
  MUX2_X1 U14052 ( .A(n11328), .B(n11327), .S(n14231), .Z(n11334) );
  OAI22_X1 U14053 ( .A1(n14267), .A2(n11331), .B1(n13813), .B2(n14250), .ZN(
        n11332) );
  AOI21_X1 U14054 ( .B1(n14265), .B2(n7675), .A(n11332), .ZN(n11333) );
  OAI211_X1 U14055 ( .C1(n14256), .C2(n11335), .A(n11334), .B(n11333), .ZN(
        P2_U3264) );
  XNOR2_X1 U14056 ( .A(n12445), .B(n11336), .ZN(n15927) );
  INV_X1 U14057 ( .A(n11337), .ZN(n11338) );
  NAND2_X1 U14058 ( .A1(n13350), .A2(n11338), .ZN(n11351) );
  NOR2_X1 U14059 ( .A1(n11339), .A2(n15946), .ZN(n15929) );
  NOR2_X1 U14060 ( .A1(n13321), .A2(n11340), .ZN(n11347) );
  XNOR2_X1 U14061 ( .A(n11341), .B(n12445), .ZN(n11345) );
  OAI22_X1 U14062 ( .A1(n11343), .A2(n13265), .B1(n11342), .B2(n13267), .ZN(
        n11344) );
  AOI21_X1 U14063 ( .B1(n11345), .B2(n13336), .A(n11344), .ZN(n11346) );
  OAI21_X1 U14064 ( .B1(n15927), .B2(n15957), .A(n11346), .ZN(n15928) );
  AOI211_X1 U14065 ( .C1(n15929), .C2(n12636), .A(n11347), .B(n15928), .ZN(
        n11348) );
  MUX2_X1 U14066 ( .A(n11349), .B(n11348), .S(n13350), .Z(n11350) );
  OAI21_X1 U14067 ( .B1(n15927), .B2(n11351), .A(n11350), .ZN(P3_U3231) );
  INV_X1 U14068 ( .A(n11352), .ZN(n11363) );
  NAND2_X1 U14069 ( .A1(n11354), .A2(n11353), .ZN(n11355) );
  OR2_X1 U14070 ( .A1(n14210), .A2(n11355), .ZN(n14200) );
  INV_X1 U14071 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n11357) );
  INV_X1 U14072 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n11356) );
  OAI22_X1 U14073 ( .A1(n14231), .A2(n11357), .B1(n11356), .B2(n14250), .ZN(
        n11358) );
  AOI21_X1 U14074 ( .B1(n14231), .B2(n11359), .A(n11358), .ZN(n11362) );
  NAND2_X1 U14075 ( .A1(n14253), .A2(n14261), .ZN(n14041) );
  INV_X1 U14076 ( .A(n14041), .ZN(n11566) );
  OAI21_X1 U14077 ( .B1(n11566), .B2(n14265), .A(n11360), .ZN(n11361) );
  OAI211_X1 U14078 ( .C1(n11363), .C2(n14200), .A(n11362), .B(n11361), .ZN(
        P2_U3265) );
  AOI21_X1 U14079 ( .B1(n11366), .B2(n11365), .A(n11364), .ZN(n11367) );
  INV_X2 U14080 ( .A(n13350), .ZN(n13346) );
  MUX2_X1 U14081 ( .A(n11367), .B(n7088), .S(n13346), .Z(n11370) );
  AOI22_X1 U14082 ( .A1(n13324), .A2(n11368), .B1(P3_REG3_REG_1__SCAN_IN), 
        .B2(n13345), .ZN(n11369) );
  NAND2_X1 U14083 ( .A1(n11370), .A2(n11369), .ZN(P3_U3232) );
  OAI21_X1 U14084 ( .B1(n15783), .B2(n11371), .A(n11645), .ZN(n11388) );
  XNOR2_X1 U14085 ( .A(n10294), .B(n11388), .ZN(n11375) );
  INV_X1 U14086 ( .A(n11373), .ZN(n11374) );
  MUX2_X1 U14087 ( .A(n11375), .B(n11374), .S(n10283), .Z(n11376) );
  OAI222_X1 U14088 ( .A1(n15467), .A2(n14709), .B1(n12723), .B2(n11377), .C1(
        n11376), .C2(n15465), .ZN(n15784) );
  INV_X1 U14089 ( .A(n15784), .ZN(n11393) );
  NOR2_X1 U14090 ( .A1(n11379), .A2(n11378), .ZN(n11380) );
  INV_X1 U14091 ( .A(n11381), .ZN(n11383) );
  OAI21_X1 U14092 ( .B1(n11373), .B2(n11385), .A(n11384), .ZN(n15786) );
  INV_X1 U14093 ( .A(n11386), .ZN(n15470) );
  AOI22_X1 U14094 ( .A1(n15286), .A2(P1_REG2_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(n15331), .ZN(n11390) );
  OR2_X1 U14095 ( .A1(n11388), .A2(n7130), .ZN(n15782) );
  OR2_X1 U14096 ( .A1(n15281), .A2(n15782), .ZN(n11389) );
  OAI211_X1 U14097 ( .C1(n15783), .C2(n15339), .A(n11390), .B(n11389), .ZN(
        n11391) );
  AOI21_X1 U14098 ( .B1(n15290), .B2(n15786), .A(n11391), .ZN(n11392) );
  OAI21_X1 U14099 ( .B1(n11393), .B2(n15286), .A(n11392), .ZN(P1_U3292) );
  INV_X1 U14100 ( .A(n11394), .ZN(n11396) );
  OAI21_X1 U14101 ( .B1(n11438), .B2(n11396), .A(n11395), .ZN(n11397) );
  XNOR2_X1 U14102 ( .A(n11397), .B(n12450), .ZN(n11398) );
  NAND2_X1 U14103 ( .A1(n11398), .A2(n13336), .ZN(n11400) );
  AOI22_X1 U14104 ( .A1(n13340), .A2(n12947), .B1(n12949), .B2(n13339), .ZN(
        n11399) );
  AND2_X1 U14105 ( .A1(n11400), .A2(n11399), .ZN(n11533) );
  XNOR2_X1 U14106 ( .A(n11401), .B(n12450), .ZN(n11532) );
  INV_X1 U14107 ( .A(n13407), .ZN(n13416) );
  INV_X1 U14108 ( .A(n13498), .ZN(n13485) );
  NAND2_X1 U14109 ( .A1(n11532), .A2(n13485), .ZN(n11403) );
  AOI22_X1 U14110 ( .A1(n13480), .A2(n11974), .B1(n15961), .B2(
        P3_REG0_REG_8__SCAN_IN), .ZN(n11402) );
  OAI211_X1 U14111 ( .C1(n15961), .C2(n11533), .A(n11403), .B(n11402), .ZN(
        P3_U3414) );
  INV_X1 U14112 ( .A(n11404), .ZN(n11406) );
  INV_X1 U14113 ( .A(n15078), .ZN(n15074) );
  OAI222_X1 U14114 ( .A1(n15546), .A2(n11405), .B1(n15549), .B2(n11406), .C1(
        n15074), .C2(P1_U3086), .ZN(P1_U3338) );
  INV_X1 U14115 ( .A(n13936), .ZN(n13928) );
  OAI222_X1 U14116 ( .A1(n14472), .A2(n11407), .B1(n14474), .B2(n11406), .C1(
        n13928), .C2(P2_U3088), .ZN(P2_U3310) );
  AND2_X1 U14117 ( .A1(n13808), .A2(n14307), .ZN(n11418) );
  XNOR2_X1 U14118 ( .A(n15890), .B(n13615), .ZN(n11419) );
  NAND2_X1 U14119 ( .A1(n11418), .A2(n11419), .ZN(n11423) );
  INV_X1 U14120 ( .A(n11418), .ZN(n11420) );
  INV_X1 U14121 ( .A(n11419), .ZN(n11429) );
  NAND2_X1 U14122 ( .A1(n11420), .A2(n11429), .ZN(n11421) );
  AND2_X1 U14123 ( .A1(n11423), .A2(n11421), .ZN(n13607) );
  NAND2_X1 U14124 ( .A1(n13807), .A2(n15891), .ZN(n11709) );
  NAND3_X1 U14125 ( .A1(n13606), .A2(n11430), .A3(n11423), .ZN(n11713) );
  OAI21_X1 U14126 ( .B1(n13606), .B2(n11430), .A(n11713), .ZN(n11433) );
  NAND2_X1 U14127 ( .A1(n13806), .A2(n13770), .ZN(n11425) );
  NAND2_X1 U14128 ( .A1(n13808), .A2(n13769), .ZN(n11424) );
  NAND2_X1 U14129 ( .A1(n11425), .A2(n11424), .ZN(n11471) );
  AOI22_X1 U14130 ( .A1(n13773), .A2(n11471), .B1(P2_REG3_REG_4__SCAN_IN), 
        .B2(P2_U3088), .ZN(n11428) );
  OR2_X1 U14131 ( .A1(n13775), .A2(n11505), .ZN(n11427) );
  OAI211_X1 U14132 ( .C1(n11506), .C2(n13749), .A(n11428), .B(n11427), .ZN(
        n11432) );
  NOR4_X1 U14133 ( .A1(n13751), .A2(n11430), .A3(n7805), .A4(n11429), .ZN(
        n11431) );
  AOI211_X1 U14134 ( .C1(n11433), .C2(n13766), .A(n11432), .B(n11431), .ZN(
        n11434) );
  INV_X1 U14135 ( .A(n11434), .ZN(P2_U3202) );
  OR2_X1 U14136 ( .A1(n11435), .A2(n12448), .ZN(n11436) );
  AND2_X1 U14137 ( .A1(n11437), .A2(n11436), .ZN(n15955) );
  OR2_X1 U14138 ( .A1(n11438), .A2(n12448), .ZN(n11699) );
  NAND2_X1 U14139 ( .A1(n11438), .A2(n12448), .ZN(n11439) );
  NAND3_X1 U14140 ( .A1(n11699), .A2(n13336), .A3(n11439), .ZN(n11441) );
  AOI22_X1 U14141 ( .A1(n13340), .A2(n12949), .B1(n12951), .B2(n13339), .ZN(
        n11440) );
  NAND2_X1 U14142 ( .A1(n11441), .A2(n11440), .ZN(n15959) );
  INV_X1 U14143 ( .A(n15959), .ZN(n11443) );
  MUX2_X1 U14144 ( .A(n11443), .B(n11442), .S(n13346), .Z(n11445) );
  AOI22_X1 U14145 ( .A1(n13310), .A2(n6977), .B1(n13345), .B2(n11668), .ZN(
        n11444) );
  OAI211_X1 U14146 ( .C1(n13352), .C2(n15955), .A(n11445), .B(n11444), .ZN(
        P3_U3227) );
  INV_X1 U14147 ( .A(n11446), .ZN(n11448) );
  INV_X1 U14148 ( .A(n15036), .ZN(n15042) );
  OAI222_X1 U14149 ( .A1(n15546), .A2(n11447), .B1(n15549), .B2(n11448), .C1(
        P1_U3086), .C2(n15042), .ZN(P1_U3341) );
  INV_X1 U14150 ( .A(n13885), .ZN(n12302) );
  OAI222_X1 U14151 ( .A1(n14472), .A2(n11449), .B1(n14474), .B2(n11448), .C1(
        P2_U3088), .C2(n12302), .ZN(P2_U3313) );
  INV_X1 U14152 ( .A(n11450), .ZN(n11461) );
  XNOR2_X1 U14153 ( .A(n12832), .B(n15947), .ZN(n11669) );
  XNOR2_X1 U14154 ( .A(n11669), .B(n11670), .ZN(n11454) );
  OAI21_X1 U14155 ( .B1(n11454), .B2(n11453), .A(n11800), .ZN(n11455) );
  NAND2_X1 U14156 ( .A1(n11455), .A2(n12924), .ZN(n11460) );
  INV_X1 U14157 ( .A(n12931), .ZN(n12914) );
  OAI22_X1 U14158 ( .A1(n12917), .A2(n11456), .B1(n15947), .B2(n12937), .ZN(
        n11457) );
  AOI211_X1 U14159 ( .C1(n12914), .C2(n12950), .A(n11458), .B(n11457), .ZN(
        n11459) );
  OAI211_X1 U14160 ( .C1(n11461), .C2(n11679), .A(n11460), .B(n11459), .ZN(
        P3_U3167) );
  AOI211_X1 U14161 ( .C1(n11465), .C2(n11464), .A(n11463), .B(n11462), .ZN(
        n11468) );
  INV_X1 U14162 ( .A(n11466), .ZN(n11467) );
  NOR2_X1 U14163 ( .A1(n11468), .A2(n11467), .ZN(n11511) );
  XNOR2_X1 U14164 ( .A(n11470), .B(n11469), .ZN(n11472) );
  AOI21_X1 U14165 ( .B1(n11472), .B2(n14270), .A(n11471), .ZN(n11503) );
  OR2_X1 U14166 ( .A1(n11564), .A2(n11506), .ZN(n11473) );
  AND3_X1 U14167 ( .A1(n11931), .A2(n11473), .A3(n14261), .ZN(n11508) );
  INV_X1 U14168 ( .A(n11508), .ZN(n11474) );
  OAI211_X1 U14169 ( .C1(n14391), .C2(n11511), .A(n11503), .B(n11474), .ZN(
        n11493) );
  OAI22_X1 U14170 ( .A1(n14349), .A2(n11506), .B1(n15912), .B2(n10695), .ZN(
        n11475) );
  AOI21_X1 U14171 ( .B1(n11493), .B2(n15912), .A(n11475), .ZN(n11476) );
  INV_X1 U14172 ( .A(n11476), .ZN(P2_U3503) );
  XNOR2_X1 U14173 ( .A(n11483), .B(P1_REG1_REG_11__SCAN_IN), .ZN(n11480) );
  AOI21_X1 U14174 ( .B1(n11480), .B2(n11479), .A(n11979), .ZN(n11490) );
  AND2_X1 U14175 ( .A1(P1_U3086), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n14659) );
  NOR2_X1 U14176 ( .A1(n15068), .A2(n11984), .ZN(n11481) );
  AOI211_X1 U14177 ( .C1(n15722), .C2(P1_ADDR_REG_11__SCAN_IN), .A(n14659), 
        .B(n11481), .ZN(n11489) );
  NOR2_X1 U14178 ( .A1(n11482), .A2(n8835), .ZN(n11485) );
  MUX2_X1 U14179 ( .A(P1_REG2_REG_11__SCAN_IN), .B(n12205), .S(n11483), .Z(
        n11484) );
  OAI21_X1 U14180 ( .B1(n11486), .B2(n11485), .A(n11484), .ZN(n11983) );
  OR3_X1 U14181 ( .A1(n11486), .A2(n11485), .A3(n11484), .ZN(n11487) );
  NAND3_X1 U14182 ( .A1(n11983), .A2(n15746), .A3(n11487), .ZN(n11488) );
  OAI211_X1 U14183 ( .C1(n11490), .C2(n15097), .A(n11489), .B(n11488), .ZN(
        P1_U3254) );
  INV_X1 U14184 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n11491) );
  OAI22_X1 U14185 ( .A1(n14430), .A2(n11506), .B1(n15908), .B2(n11491), .ZN(
        n11492) );
  AOI21_X1 U14186 ( .B1(n11493), .B2(n15908), .A(n11492), .ZN(n11494) );
  INV_X1 U14187 ( .A(n11494), .ZN(P2_U3442) );
  INV_X1 U14188 ( .A(n11495), .ZN(n11569) );
  AOI22_X1 U14189 ( .A1(n15743), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_15__SCAN_IN), .B2(n15527), .ZN(n11496) );
  OAI21_X1 U14190 ( .B1(n11569), .B2(n15549), .A(n11496), .ZN(P1_U3340) );
  NOR2_X1 U14191 ( .A1(n15281), .A2(n7130), .ZN(n15329) );
  OAI21_X1 U14192 ( .B1(n15329), .B2(n15291), .A(n11497), .ZN(n11499) );
  AOI22_X1 U14193 ( .A1(n15286), .A2(P1_REG2_REG_0__SCAN_IN), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(n15331), .ZN(n11498) );
  OAI211_X1 U14194 ( .C1(n15286), .C2(n11500), .A(n11499), .B(n11498), .ZN(
        P1_U3293) );
  INV_X1 U14195 ( .A(n13406), .ZN(n13398) );
  AOI22_X1 U14196 ( .A1(n11532), .A2(n13398), .B1(n13395), .B2(n11974), .ZN(
        n11502) );
  MUX2_X1 U14197 ( .A(n11533), .B(n11573), .S(n15970), .Z(n11501) );
  NAND2_X1 U14198 ( .A1(n11502), .A2(n11501), .ZN(P3_U3467) );
  MUX2_X1 U14199 ( .A(n11504), .B(n11503), .S(n14231), .Z(n11510) );
  OAI22_X1 U14200 ( .A1(n14251), .A2(n11506), .B1(n11505), .B2(n14250), .ZN(
        n11507) );
  AOI21_X1 U14201 ( .B1(n14253), .B2(n11508), .A(n11507), .ZN(n11509) );
  OAI211_X1 U14202 ( .C1(n14256), .C2(n11511), .A(n11510), .B(n11509), .ZN(
        P2_U3261) );
  INV_X1 U14203 ( .A(n11646), .ZN(n11514) );
  INV_X1 U14204 ( .A(n11512), .ZN(n11513) );
  OAI211_X1 U14205 ( .C1(n14701), .C2(n11514), .A(n11513), .B(n15447), .ZN(
        n15788) );
  INV_X1 U14206 ( .A(n11515), .ZN(n11524) );
  NAND2_X1 U14207 ( .A1(n14970), .A2(n15801), .ZN(n11516) );
  OAI21_X1 U14208 ( .B1(n14709), .B2(n12723), .A(n11516), .ZN(n15707) );
  NOR2_X1 U14209 ( .A1(n11517), .A2(n15465), .ZN(n11522) );
  INV_X1 U14210 ( .A(n11517), .ZN(n11520) );
  NAND3_X1 U14211 ( .A1(n11518), .A2(n15812), .A3(n9144), .ZN(n11519) );
  OAI21_X1 U14212 ( .B1(n11520), .B2(n15465), .A(n11519), .ZN(n11521) );
  MUX2_X1 U14213 ( .A(n11522), .B(n11521), .S(n14924), .Z(n11523) );
  AOI211_X1 U14214 ( .C1(n11524), .C2(n15812), .A(n15707), .B(n11523), .ZN(
        n15789) );
  MUX2_X1 U14215 ( .A(n11525), .B(n15789), .S(n15312), .Z(n11528) );
  INV_X1 U14216 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n11526) );
  AOI22_X1 U14217 ( .A1(n15291), .A2(n6534), .B1(n15331), .B2(n11526), .ZN(
        n11527) );
  OAI211_X1 U14218 ( .C1(n15281), .C2(n15788), .A(n11528), .B(n11527), .ZN(
        P1_U3290) );
  INV_X1 U14219 ( .A(n11529), .ZN(n11530) );
  OAI222_X1 U14220 ( .A1(P3_U3151), .A2(n13128), .B1(n13528), .B2(n11531), 
        .C1(n13524), .C2(n11530), .ZN(P3_U3276) );
  INV_X1 U14221 ( .A(n11532), .ZN(n11537) );
  AOI22_X1 U14222 ( .A1(n13310), .A2(n11974), .B1(n13345), .B2(n11975), .ZN(
        n11536) );
  MUX2_X1 U14223 ( .A(n11534), .B(n11533), .S(n13350), .Z(n11535) );
  OAI211_X1 U14224 ( .C1(n11537), .C2(n13352), .A(n11536), .B(n11535), .ZN(
        P3_U3225) );
  XNOR2_X1 U14225 ( .A(n11538), .B(n11539), .ZN(n11630) );
  NAND2_X1 U14226 ( .A1(n11540), .A2(n11539), .ZN(n11541) );
  NAND3_X1 U14227 ( .A1(n11542), .A2(n13336), .A3(n11541), .ZN(n11544) );
  AOI22_X1 U14228 ( .A1(n12948), .A2(n13339), .B1(n13340), .B2(n12946), .ZN(
        n11543) );
  NAND2_X1 U14229 ( .A1(n11544), .A2(n11543), .ZN(n11632) );
  AOI21_X1 U14230 ( .B1(n11630), .B2(n13407), .A(n11632), .ZN(n11820) );
  INV_X1 U14231 ( .A(n12551), .ZN(n11631) );
  AOI22_X1 U14232 ( .A1(n13480), .A2(n11631), .B1(P3_REG0_REG_9__SCAN_IN), 
        .B2(n15961), .ZN(n11545) );
  OAI21_X1 U14233 ( .B1(n11820), .B2(n15961), .A(n11545), .ZN(P3_U3417) );
  NAND2_X1 U14234 ( .A1(n11547), .A2(n11546), .ZN(n11549) );
  XNOR2_X1 U14235 ( .A(n11549), .B(n11548), .ZN(n11553) );
  NAND2_X1 U14236 ( .A1(P1_U3086), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n15007) );
  OAI21_X1 U14237 ( .B1(n14680), .B2(n11849), .A(n15007), .ZN(n11551) );
  OAI22_X1 U14238 ( .A1(n14695), .A2(n14681), .B1(n15713), .B2(n11724), .ZN(
        n11550) );
  AOI211_X1 U14239 ( .C1(n14684), .C2(n7945), .A(n11551), .B(n11550), .ZN(
        n11552) );
  OAI21_X1 U14240 ( .B1(n11553), .B2(n14686), .A(n11552), .ZN(P1_U3230) );
  NAND2_X1 U14241 ( .A1(n11555), .A2(n11554), .ZN(n11556) );
  XNOR2_X1 U14242 ( .A(n11556), .B(n11557), .ZN(n15888) );
  INV_X1 U14243 ( .A(n14250), .ZN(n14263) );
  INV_X1 U14244 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n11561) );
  AOI22_X1 U14245 ( .A1(n13769), .A2(n13809), .B1(n13807), .B2(n13770), .ZN(
        n13609) );
  XNOR2_X1 U14246 ( .A(n11558), .B(n11557), .ZN(n11559) );
  NAND2_X1 U14247 ( .A1(n11559), .A2(n14270), .ZN(n11560) );
  OAI211_X1 U14248 ( .C1(n15888), .C2(n11003), .A(n13609), .B(n11560), .ZN(
        n15893) );
  AOI21_X1 U14249 ( .B1(n14263), .B2(n11561), .A(n15893), .ZN(n11562) );
  MUX2_X1 U14250 ( .A(n11563), .B(n11562), .S(n14231), .Z(n11568) );
  AOI21_X1 U14251 ( .B1(n15890), .B2(n11565), .A(n11564), .ZN(n15889) );
  AOI22_X1 U14252 ( .A1(n11566), .A2(n15889), .B1(n14265), .B2(n15890), .ZN(
        n11567) );
  OAI211_X1 U14253 ( .C1(n15888), .C2(n14200), .A(n11568), .B(n11567), .ZN(
        P2_U3262) );
  INV_X1 U14254 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n11570) );
  INV_X1 U14255 ( .A(n13893), .ZN(n13901) );
  OAI222_X1 U14256 ( .A1(n14472), .A2(n11570), .B1(n14474), .B2(n11569), .C1(
        n13901), .C2(P2_U3088), .ZN(P2_U3312) );
  OR2_X1 U14257 ( .A1(n11574), .A2(n11573), .ZN(n11575) );
  INV_X1 U14258 ( .A(n11594), .ZN(n11578) );
  XNOR2_X1 U14259 ( .A(n11595), .B(n11578), .ZN(n11593) );
  INV_X1 U14260 ( .A(P3_REG1_REG_9__SCAN_IN), .ZN(n11821) );
  XNOR2_X1 U14261 ( .A(n11593), .B(n11821), .ZN(n11592) );
  OAI21_X1 U14262 ( .B1(P3_REG2_REG_9__SCAN_IN), .B2(n11580), .A(n11601), .ZN(
        n11590) );
  INV_X1 U14263 ( .A(n11581), .ZN(n11584) );
  MUX2_X1 U14264 ( .A(P3_REG2_REG_9__SCAN_IN), .B(P3_REG1_REG_9__SCAN_IN), .S(
        n7233), .Z(n11582) );
  NOR2_X1 U14265 ( .A1(n11582), .A2(n11594), .ZN(n11603) );
  AOI21_X1 U14266 ( .B1(n11582), .B2(n11594), .A(n11603), .ZN(n11583) );
  OR3_X1 U14267 ( .A1(n11585), .A2(n11584), .A3(n11583), .ZN(n11586) );
  AOI21_X1 U14268 ( .B1(n11611), .B2(n11586), .A(n13116), .ZN(n11589) );
  NAND2_X1 U14269 ( .A1(P3_U3151), .A2(P3_REG3_REG_9__SCAN_IN), .ZN(n11813) );
  NAND2_X1 U14270 ( .A1(n15913), .A2(P3_ADDR_REG_9__SCAN_IN), .ZN(n11587) );
  OAI211_X1 U14271 ( .C1(n13129), .C2(n11594), .A(n11813), .B(n11587), .ZN(
        n11588) );
  AOI211_X1 U14272 ( .C1(n11590), .C2(n15916), .A(n11589), .B(n11588), .ZN(
        n11591) );
  OAI21_X1 U14273 ( .B1(n11592), .B2(n13118), .A(n11591), .ZN(P3_U3191) );
  INV_X1 U14274 ( .A(P3_REG1_REG_10__SCAN_IN), .ZN(n11604) );
  XNOR2_X1 U14275 ( .A(n12089), .B(n11604), .ZN(n12085) );
  NAND2_X1 U14276 ( .A1(n11593), .A2(P3_REG1_REG_9__SCAN_IN), .ZN(n11597) );
  NAND2_X1 U14277 ( .A1(n11595), .A2(n11594), .ZN(n11596) );
  XOR2_X1 U14278 ( .A(n12086), .B(n12085), .Z(n11619) );
  INV_X1 U14279 ( .A(n11598), .ZN(n11599) );
  XNOR2_X1 U14280 ( .A(n12089), .B(P3_REG2_REG_10__SCAN_IN), .ZN(n11600) );
  AND3_X1 U14281 ( .A1(n11601), .A2(n11600), .A3(n11599), .ZN(n11602) );
  OAI21_X1 U14282 ( .B1(n12088), .B2(n11602), .A(n15916), .ZN(n11618) );
  INV_X1 U14283 ( .A(n12089), .ZN(n11616) );
  INV_X1 U14284 ( .A(P3_ADDR_REG_10__SCAN_IN), .ZN(n15573) );
  NAND2_X1 U14285 ( .A1(P3_U3151), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n11872)
         );
  OAI21_X1 U14286 ( .B1(n15925), .B2(n15573), .A(n11872), .ZN(n11615) );
  INV_X1 U14287 ( .A(n11603), .ZN(n11610) );
  INV_X1 U14288 ( .A(P3_REG2_REG_10__SCAN_IN), .ZN(n11605) );
  MUX2_X1 U14289 ( .A(n11605), .B(n11604), .S(n6527), .Z(n11606) );
  NAND2_X1 U14290 ( .A1(n11606), .A2(n11616), .ZN(n12092) );
  INV_X1 U14291 ( .A(n11606), .ZN(n11607) );
  NAND2_X1 U14292 ( .A1(n11607), .A2(n12089), .ZN(n11608) );
  NAND2_X1 U14293 ( .A1(n12092), .A2(n11608), .ZN(n11609) );
  AOI21_X1 U14294 ( .B1(n11611), .B2(n11610), .A(n11609), .ZN(n12094) );
  INV_X1 U14295 ( .A(n12094), .ZN(n11613) );
  NAND3_X1 U14296 ( .A1(n11611), .A2(n11610), .A3(n11609), .ZN(n11612) );
  AOI21_X1 U14297 ( .B1(n11613), .B2(n11612), .A(n13116), .ZN(n11614) );
  AOI211_X1 U14298 ( .C1(n15922), .C2(n11616), .A(n11615), .B(n11614), .ZN(
        n11617) );
  OAI211_X1 U14299 ( .C1(n11619), .C2(n13118), .A(n11618), .B(n11617), .ZN(
        P3_U3192) );
  NAND2_X1 U14300 ( .A1(n11621), .A2(n11620), .ZN(n11622) );
  XNOR2_X1 U14301 ( .A(n11623), .B(n11622), .ZN(n11629) );
  OAI21_X1 U14302 ( .B1(n14680), .B2(n14481), .A(n11624), .ZN(n11627) );
  OAI22_X1 U14303 ( .A1(n11625), .A2(n14681), .B1(n15713), .B2(n11884), .ZN(
        n11626) );
  AOI211_X1 U14304 ( .C1(n14684), .C2(n14725), .A(n11627), .B(n11626), .ZN(
        n11628) );
  OAI21_X1 U14305 ( .B1(n11629), .B2(n14686), .A(n11628), .ZN(P1_U3227) );
  INV_X1 U14306 ( .A(n11630), .ZN(n11636) );
  AOI22_X1 U14307 ( .A1(n13310), .A2(n11631), .B1(n13345), .B2(n11817), .ZN(
        n11635) );
  INV_X1 U14308 ( .A(n11632), .ZN(n11633) );
  MUX2_X1 U14309 ( .A(n11633), .B(n6773), .S(n13346), .Z(n11634) );
  OAI211_X1 U14310 ( .C1(n11636), .C2(n13352), .A(n11635), .B(n11634), .ZN(
        P3_U3224) );
  INV_X1 U14311 ( .A(n11518), .ZN(n11644) );
  OAI22_X1 U14312 ( .A1(n10294), .A2(n12723), .B1(n14695), .B2(n15467), .ZN(
        n11643) );
  NOR2_X1 U14313 ( .A1(n11637), .A2(n15465), .ZN(n11641) );
  INV_X1 U14314 ( .A(n11637), .ZN(n14694) );
  NAND3_X1 U14315 ( .A1(n11384), .A2(n15812), .A3(n11638), .ZN(n11639) );
  OAI21_X1 U14316 ( .B1(n14694), .B2(n15465), .A(n11639), .ZN(n11640) );
  MUX2_X1 U14317 ( .A(n11641), .B(n11640), .S(n14923), .Z(n11642) );
  AOI211_X1 U14318 ( .C1(n11644), .C2(n15812), .A(n11643), .B(n11642), .ZN(
        n11691) );
  OAI211_X1 U14319 ( .C1(n7361), .C2(n14699), .A(n15447), .B(n11646), .ZN(
        n11695) );
  OAI211_X1 U14320 ( .C1(n14699), .C2(n15804), .A(n11691), .B(n11695), .ZN(
        n11665) );
  NAND2_X1 U14321 ( .A1(n11665), .A2(n15822), .ZN(n11647) );
  OAI21_X1 U14322 ( .B1(n15822), .B2(n8686), .A(n11647), .ZN(P1_U3530) );
  NAND2_X1 U14323 ( .A1(n11655), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n11648) );
  NAND2_X1 U14324 ( .A1(n11649), .A2(n11648), .ZN(n11653) );
  INV_X1 U14325 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n11650) );
  MUX2_X1 U14326 ( .A(n11650), .B(P2_REG2_REG_11__SCAN_IN), .S(n11826), .Z(
        n11652) );
  INV_X1 U14327 ( .A(n11832), .ZN(n11651) );
  AOI21_X1 U14328 ( .B1(n11653), .B2(n11652), .A(n11651), .ZN(n11664) );
  INV_X1 U14329 ( .A(n15866), .ZN(n15823) );
  XNOR2_X1 U14330 ( .A(n11826), .B(P2_REG1_REG_11__SCAN_IN), .ZN(n11656) );
  AOI211_X1 U14331 ( .C1(n11657), .C2(n11656), .A(n15860), .B(n11823), .ZN(
        n11658) );
  INV_X1 U14332 ( .A(n11658), .ZN(n11663) );
  NOR2_X1 U14333 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9703), .ZN(n11661) );
  NOR2_X1 U14334 ( .A1(n15871), .A2(n11659), .ZN(n11660) );
  AOI211_X1 U14335 ( .C1(n15864), .C2(P2_ADDR_REG_11__SCAN_IN), .A(n11661), 
        .B(n11660), .ZN(n11662) );
  OAI211_X1 U14336 ( .C1(n11664), .C2(n15823), .A(n11663), .B(n11662), .ZN(
        P2_U3225) );
  INV_X1 U14337 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n11667) );
  NAND2_X1 U14338 ( .A1(n11665), .A2(n15815), .ZN(n11666) );
  OAI21_X1 U14339 ( .B1(n15815), .B2(n11667), .A(n11666), .ZN(P1_U3465) );
  INV_X1 U14340 ( .A(n11668), .ZN(n11680) );
  INV_X1 U14341 ( .A(n11669), .ZN(n11671) );
  NAND2_X1 U14342 ( .A1(n11671), .A2(n11670), .ZN(n11796) );
  AND2_X1 U14343 ( .A1(n11800), .A2(n11796), .ZN(n11673) );
  XNOR2_X1 U14344 ( .A(n12832), .B(n11674), .ZN(n11797) );
  XOR2_X1 U14345 ( .A(n12950), .B(n11797), .Z(n11672) );
  NAND2_X1 U14346 ( .A1(n11673), .A2(n11672), .ZN(n11758) );
  OAI211_X1 U14347 ( .C1(n11673), .C2(n11672), .A(n11758), .B(n12924), .ZN(
        n11678) );
  INV_X1 U14348 ( .A(n12949), .ZN(n11801) );
  OAI22_X1 U14349 ( .A1(n12937), .A2(n11674), .B1(n12931), .B2(n11801), .ZN(
        n11675) );
  AOI211_X1 U14350 ( .C1(n12929), .C2(n12951), .A(n11676), .B(n11675), .ZN(
        n11677) );
  OAI211_X1 U14351 ( .C1(n11680), .C2(n11679), .A(n11678), .B(n11677), .ZN(
        P3_U3179) );
  INV_X1 U14352 ( .A(n11681), .ZN(n11690) );
  NAND2_X1 U14353 ( .A1(n11682), .A2(n14278), .ZN(n11688) );
  AOI22_X1 U14354 ( .A1(n14253), .A2(n11683), .B1(P2_REG3_REG_2__SCAN_IN), 
        .B2(n14263), .ZN(n11687) );
  OR2_X1 U14355 ( .A1(n14251), .A2(n11684), .ZN(n11686) );
  NAND2_X1 U14356 ( .A1(n14275), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n11685) );
  AND4_X1 U14357 ( .A1(n11688), .A2(n11687), .A3(n11686), .A4(n11685), .ZN(
        n11689) );
  OAI21_X1 U14358 ( .B1(n11690), .B2(n14275), .A(n11689), .ZN(P2_U3263) );
  MUX2_X1 U14359 ( .A(n11692), .B(n11691), .S(n15312), .Z(n11694) );
  AOI22_X1 U14360 ( .A1(n15291), .A2(n14708), .B1(P1_REG3_REG_2__SCAN_IN), 
        .B2(n15331), .ZN(n11693) );
  OAI211_X1 U14361 ( .C1(n15281), .C2(n11695), .A(n11694), .B(n11693), .ZN(
        P1_U3291) );
  XNOR2_X1 U14362 ( .A(n11696), .B(n11760), .ZN(n13415) );
  INV_X1 U14363 ( .A(n11697), .ZN(n11698) );
  NAND2_X1 U14364 ( .A1(n11699), .A2(n11698), .ZN(n11700) );
  XNOR2_X1 U14365 ( .A(n11700), .B(n12535), .ZN(n11701) );
  NAND2_X1 U14366 ( .A1(n11701), .A2(n13336), .ZN(n11703) );
  AOI22_X1 U14367 ( .A1(n12948), .A2(n13340), .B1(n13339), .B2(n12950), .ZN(
        n11702) );
  NAND2_X1 U14368 ( .A1(n11703), .A2(n11702), .ZN(n13412) );
  INV_X1 U14369 ( .A(n13412), .ZN(n11705) );
  INV_X1 U14370 ( .A(P3_REG2_REG_7__SCAN_IN), .ZN(n11704) );
  MUX2_X1 U14371 ( .A(n11705), .B(n11704), .S(n13346), .Z(n11707) );
  AOI22_X1 U14372 ( .A1(n13310), .A2(n13413), .B1(n13345), .B2(n11764), .ZN(
        n11706) );
  OAI211_X1 U14373 ( .C1(n13352), .C2(n13415), .A(n11707), .B(n11706), .ZN(
        P3_U3226) );
  INV_X1 U14374 ( .A(n11714), .ZN(n11708) );
  NAND2_X1 U14375 ( .A1(n11709), .A2(n11708), .ZN(n11710) );
  XNOR2_X1 U14376 ( .A(n11930), .B(n13615), .ZN(n11768) );
  NAND2_X1 U14377 ( .A1(n13806), .A2(n15891), .ZN(n11770) );
  XNOR2_X1 U14378 ( .A(n11768), .B(n11770), .ZN(n11715) );
  OAI22_X1 U14379 ( .A1(n11899), .A2(n13743), .B1(n11711), .B2(n13741), .ZN(
        n11927) );
  NAND2_X1 U14380 ( .A1(n13773), .A2(n11927), .ZN(n11712) );
  NAND2_X1 U14381 ( .A1(P2_REG3_REG_5__SCAN_IN), .A2(P2_U3088), .ZN(n13837) );
  OAI211_X1 U14382 ( .C1(n13775), .C2(n11933), .A(n11712), .B(n13837), .ZN(
        n11719) );
  INV_X1 U14383 ( .A(n11713), .ZN(n11717) );
  AOI22_X1 U14384 ( .A1(n13765), .A2(n13807), .B1(n13766), .B2(n11714), .ZN(
        n11716) );
  NOR3_X1 U14385 ( .A1(n11717), .A2(n11716), .A3(n11715), .ZN(n11718) );
  AOI211_X1 U14386 ( .C1(n11930), .C2(n13777), .A(n11719), .B(n11718), .ZN(
        n11720) );
  OAI21_X1 U14387 ( .B1(n11772), .B2(n13736), .A(n11720), .ZN(P2_U3199) );
  INV_X1 U14388 ( .A(n11721), .ZN(n11732) );
  NOR2_X1 U14389 ( .A1(n11722), .A2(n15103), .ZN(n11723) );
  MUX2_X1 U14390 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n11723), .S(n15312), .Z(
        n11728) );
  NOR2_X1 U14391 ( .A1(n15286), .A2(n12723), .ZN(n15336) );
  INV_X1 U14392 ( .A(n15336), .ZN(n15255) );
  NOR2_X1 U14393 ( .A1(n15286), .A2(n15467), .ZN(n15257) );
  INV_X1 U14394 ( .A(n11724), .ZN(n11725) );
  AOI22_X1 U14395 ( .A1(n15257), .A2(n14969), .B1(n11725), .B2(n15331), .ZN(
        n11726) );
  OAI21_X1 U14396 ( .B1(n14695), .B2(n15255), .A(n11726), .ZN(n11727) );
  AOI211_X1 U14397 ( .C1(n15291), .C2(n7945), .A(n11728), .B(n11727), .ZN(
        n11731) );
  NAND3_X1 U14398 ( .A1(n11281), .A2(n11729), .A3(n15341), .ZN(n11730) );
  OAI211_X1 U14399 ( .C1(n11732), .C2(n15343), .A(n11731), .B(n11730), .ZN(
        P1_U3289) );
  AOI211_X1 U14400 ( .C1(n14725), .C2(n11733), .A(n7130), .B(n6573), .ZN(
        n11889) );
  INV_X1 U14401 ( .A(n11734), .ZN(n11737) );
  INV_X1 U14402 ( .A(n11735), .ZN(n11736) );
  OR2_X1 U14403 ( .A1(n11736), .A2(n11851), .ZN(n14922) );
  AOI21_X1 U14404 ( .B1(n11738), .B2(n11737), .A(n14922), .ZN(n11852) );
  NAND2_X1 U14405 ( .A1(n11852), .A2(n15812), .ZN(n11746) );
  AOI22_X1 U14406 ( .A1(n15798), .A2(n14970), .B1(n14968), .B2(n15801), .ZN(
        n11745) );
  NAND3_X1 U14407 ( .A1(n11738), .A2(n15812), .A3(n11737), .ZN(n11739) );
  OAI21_X1 U14408 ( .B1(n11742), .B2(n15465), .A(n11739), .ZN(n11740) );
  NAND2_X1 U14409 ( .A1(n11740), .A2(n14922), .ZN(n11744) );
  INV_X1 U14410 ( .A(n14922), .ZN(n11741) );
  NAND3_X1 U14411 ( .A1(n11742), .A2(n11741), .A3(n15807), .ZN(n11743) );
  NAND4_X1 U14412 ( .A1(n11746), .A2(n11745), .A3(n11744), .A4(n11743), .ZN(
        n11886) );
  NAND2_X1 U14413 ( .A1(n15820), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n11747) );
  OAI21_X1 U14414 ( .B1(n11749), .B2(n15820), .A(n11747), .ZN(P1_U3533) );
  NAND2_X1 U14415 ( .A1(n15813), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n11748) );
  OAI21_X1 U14416 ( .B1(n11749), .B2(n15813), .A(n11748), .ZN(P1_U3474) );
  INV_X1 U14417 ( .A(n11750), .ZN(n11751) );
  OAI222_X1 U14418 ( .A1(P3_U3151), .A2(n11753), .B1(n13521), .B2(n11752), 
        .C1(n13524), .C2(n11751), .ZN(P3_U3275) );
  INV_X1 U14419 ( .A(n11754), .ZN(n11756) );
  INV_X1 U14420 ( .A(n15093), .ZN(n15086) );
  OAI222_X1 U14421 ( .A1(n15546), .A2(n11755), .B1(n15549), .B2(n11756), .C1(
        n15086), .C2(P1_U3086), .ZN(P1_U3337) );
  OAI222_X1 U14422 ( .A1(n14472), .A2(n11757), .B1(n14474), .B2(n11756), .C1(
        n15870), .C2(P2_U3088), .ZN(P2_U3309) );
  NAND2_X1 U14423 ( .A1(n11797), .A2(n12950), .ZN(n11803) );
  NAND2_X1 U14424 ( .A1(n11758), .A2(n11803), .ZN(n11968) );
  XNOR2_X1 U14425 ( .A(n11968), .B(n11802), .ZN(n11767) );
  OAI22_X1 U14426 ( .A1(n12917), .A2(n6974), .B1(n12937), .B2(n11761), .ZN(
        n11762) );
  AOI211_X1 U14427 ( .C1(n12914), .C2(n12948), .A(n11763), .B(n11762), .ZN(
        n11766) );
  NAND2_X1 U14428 ( .A1(n12934), .A2(n11764), .ZN(n11765) );
  OAI211_X1 U14429 ( .C1(n11767), .C2(n12922), .A(n11766), .B(n11765), .ZN(
        P3_U3153) );
  INV_X1 U14430 ( .A(n11768), .ZN(n11769) );
  NAND2_X1 U14431 ( .A1(n11770), .A2(n11769), .ZN(n11771) );
  XNOR2_X1 U14432 ( .A(n12009), .B(n13615), .ZN(n11773) );
  AND2_X1 U14433 ( .A1(n13805), .A2(n15891), .ZN(n11774) );
  NAND2_X1 U14434 ( .A1(n11773), .A2(n11774), .ZN(n11893) );
  INV_X1 U14435 ( .A(n11773), .ZN(n11892) );
  INV_X1 U14436 ( .A(n11774), .ZN(n11775) );
  NAND2_X1 U14437 ( .A1(n11892), .A2(n11775), .ZN(n11776) );
  NAND2_X1 U14438 ( .A1(n11893), .A2(n11776), .ZN(n11778) );
  AOI21_X1 U14439 ( .B1(n11777), .B2(n11778), .A(n13736), .ZN(n11780) );
  INV_X1 U14440 ( .A(n11778), .ZN(n11779) );
  NAND2_X1 U14441 ( .A1(n11780), .A2(n11894), .ZN(n11786) );
  INV_X1 U14442 ( .A(n12013), .ZN(n11784) );
  NAND2_X1 U14443 ( .A1(n13804), .A2(n13770), .ZN(n11782) );
  NAND2_X1 U14444 ( .A1(n13806), .A2(n13769), .ZN(n11781) );
  AND2_X1 U14445 ( .A1(n11782), .A2(n11781), .ZN(n12005) );
  NAND2_X1 U14446 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_U3088), .ZN(n13850) );
  OAI21_X1 U14447 ( .B1(n13759), .B2(n12005), .A(n13850), .ZN(n11783) );
  AOI21_X1 U14448 ( .B1(n11784), .B2(n13756), .A(n11783), .ZN(n11785) );
  OAI211_X1 U14449 ( .C1(n15901), .C2(n13749), .A(n11786), .B(n11785), .ZN(
        P2_U3211) );
  XNOR2_X1 U14450 ( .A(n11788), .B(n11787), .ZN(n11960) );
  INV_X1 U14451 ( .A(n11954), .ZN(n11917) );
  AOI22_X1 U14452 ( .A1(n13480), .A2(n11917), .B1(P3_REG0_REG_10__SCAN_IN), 
        .B2(n15961), .ZN(n11794) );
  OAI211_X1 U14453 ( .C1(n11790), .C2(n12558), .A(n11789), .B(n13336), .ZN(
        n11792) );
  AOI22_X1 U14454 ( .A1(n13339), .A2(n12947), .B1(n12945), .B2(n13340), .ZN(
        n11791) );
  NAND2_X1 U14455 ( .A1(n11792), .A2(n11791), .ZN(n11955) );
  NAND2_X1 U14456 ( .A1(n11955), .A2(n15963), .ZN(n11793) );
  OAI211_X1 U14457 ( .C1(n11960), .C2(n13498), .A(n11794), .B(n11793), .ZN(
        P3_U3420) );
  XNOR2_X1 U14458 ( .A(n12551), .B(n7285), .ZN(n11864) );
  XNOR2_X1 U14459 ( .A(n11864), .B(n12947), .ZN(n11812) );
  XNOR2_X1 U14460 ( .A(n12791), .B(n11974), .ZN(n11804) );
  XNOR2_X1 U14461 ( .A(n11804), .B(n11795), .ZN(n11970) );
  OAI211_X1 U14462 ( .C1(n11797), .C2(n12950), .A(n11796), .B(n11802), .ZN(
        n11798) );
  NOR2_X1 U14463 ( .A1(n11970), .A2(n11798), .ZN(n11799) );
  NAND2_X1 U14464 ( .A1(n11800), .A2(n11799), .ZN(n11808) );
  INV_X1 U14465 ( .A(n11802), .ZN(n11967) );
  OAI21_X1 U14466 ( .B1(n11970), .B2(n11801), .A(n11967), .ZN(n11806) );
  INV_X1 U14467 ( .A(n11804), .ZN(n11805) );
  INV_X1 U14468 ( .A(n11869), .ZN(n11810) );
  AOI21_X1 U14469 ( .B1(n11812), .B2(n11811), .A(n11810), .ZN(n11819) );
  OAI21_X1 U14470 ( .B1(n12931), .B2(n11866), .A(n11813), .ZN(n11814) );
  AOI21_X1 U14471 ( .B1(n12929), .B2(n12948), .A(n11814), .ZN(n11815) );
  OAI21_X1 U14472 ( .B1(n12551), .B2(n12937), .A(n11815), .ZN(n11816) );
  AOI21_X1 U14473 ( .B1(n11817), .B2(n12934), .A(n11816), .ZN(n11818) );
  OAI21_X1 U14474 ( .B1(n11819), .B2(n12922), .A(n11818), .ZN(P3_U3171) );
  MUX2_X1 U14475 ( .A(n11821), .B(n11820), .S(n15973), .Z(n11822) );
  OAI21_X1 U14476 ( .B1(n13403), .B2(n12551), .A(n11822), .ZN(P3_U3468) );
  XOR2_X1 U14477 ( .A(P2_REG1_REG_12__SCAN_IN), .B(n12305), .Z(n11825) );
  OAI21_X1 U14478 ( .B1(n11825), .B2(n11824), .A(n12304), .ZN(n11837) );
  OR2_X1 U14479 ( .A1(n11826), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n11830) );
  INV_X1 U14480 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n11827) );
  MUX2_X1 U14481 ( .A(P2_REG2_REG_12__SCAN_IN), .B(n11827), .S(n12305), .Z(
        n11829) );
  NAND2_X1 U14482 ( .A1(n11828), .A2(n11829), .ZN(n12297) );
  INV_X1 U14483 ( .A(n11829), .ZN(n11831) );
  NAND3_X1 U14484 ( .A1(n11832), .A2(n11831), .A3(n11830), .ZN(n11833) );
  AOI21_X1 U14485 ( .B1(n12297), .B2(n11833), .A(n15823), .ZN(n11836) );
  INV_X1 U14486 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n15679) );
  NAND2_X1 U14487 ( .A1(n15850), .A2(n12305), .ZN(n11834) );
  NAND2_X1 U14488 ( .A1(P2_U3088), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n13644)
         );
  OAI211_X1 U14489 ( .C1(n15679), .C2(n15857), .A(n11834), .B(n13644), .ZN(
        n11835) );
  AOI211_X1 U14490 ( .C1(n11837), .C2(n15830), .A(n11836), .B(n11835), .ZN(
        n11838) );
  INV_X1 U14491 ( .A(n11838), .ZN(P2_U3226) );
  XNOR2_X1 U14492 ( .A(n11840), .B(n11839), .ZN(n11841) );
  XNOR2_X1 U14493 ( .A(n11842), .B(n11841), .ZN(n11847) );
  OAI22_X1 U14494 ( .A1(n14681), .A2(n11849), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n11843), .ZN(n11845) );
  OAI22_X1 U14495 ( .A1(n14550), .A2(n14680), .B1(n15713), .B2(n11860), .ZN(
        n11844) );
  AOI211_X1 U14496 ( .C1(n14684), .C2(n14729), .A(n11845), .B(n11844), .ZN(
        n11846) );
  OAI21_X1 U14497 ( .B1(n11847), .B2(n14686), .A(n11846), .ZN(P1_U3239) );
  OAI211_X1 U14498 ( .C1(n7943), .C2(n6573), .A(n7946), .B(n15447), .ZN(n15790) );
  OAI21_X1 U14499 ( .B1(n8029), .B2(n8770), .A(n11848), .ZN(n11858) );
  OAI22_X1 U14500 ( .A1(n14550), .A2(n15467), .B1(n11849), .B2(n12723), .ZN(
        n11857) );
  OR3_X1 U14501 ( .A1(n11852), .A2(n11851), .A3(n11850), .ZN(n11855) );
  AOI21_X1 U14502 ( .B1(n11855), .B2(n11854), .A(n15492), .ZN(n11856) );
  AOI211_X1 U14503 ( .C1(n15807), .C2(n11858), .A(n11857), .B(n11856), .ZN(
        n15791) );
  MUX2_X1 U14504 ( .A(n11859), .B(n15791), .S(n15312), .Z(n11863) );
  INV_X1 U14505 ( .A(n11860), .ZN(n11861) );
  AOI22_X1 U14506 ( .A1(n15291), .A2(n14729), .B1(n11861), .B2(n15331), .ZN(
        n11862) );
  OAI211_X1 U14507 ( .C1(n15281), .C2(n15790), .A(n11863), .B(n11862), .ZN(
        P1_U3287) );
  INV_X1 U14508 ( .A(n11864), .ZN(n11865) );
  NAND2_X1 U14509 ( .A1(n11865), .A2(n12552), .ZN(n11867) );
  AND2_X1 U14510 ( .A1(n11869), .A2(n11867), .ZN(n11871) );
  XNOR2_X1 U14511 ( .A(n11954), .B(n7285), .ZN(n12117) );
  XNOR2_X1 U14512 ( .A(n12117), .B(n11866), .ZN(n11870) );
  AND2_X1 U14513 ( .A1(n11870), .A2(n11867), .ZN(n11868) );
  OAI211_X1 U14514 ( .C1(n11871), .C2(n11870), .A(n12924), .B(n12119), .ZN(
        n11876) );
  NAND2_X1 U14515 ( .A1(n12929), .A2(n12947), .ZN(n11873) );
  OAI211_X1 U14516 ( .C1(n12120), .C2(n12931), .A(n11873), .B(n11872), .ZN(
        n11874) );
  AOI21_X1 U14517 ( .B1(n12934), .B2(n11958), .A(n11874), .ZN(n11875) );
  OAI211_X1 U14518 ( .C1(n12937), .C2(n11954), .A(n11876), .B(n11875), .ZN(
        P3_U3157) );
  INV_X1 U14519 ( .A(n11877), .ZN(n11879) );
  OAI222_X1 U14520 ( .A1(n15546), .A2(n11878), .B1(n15549), .B2(n11879), .C1(
        P1_U3086), .C2(n15178), .ZN(P1_U3336) );
  OAI222_X1 U14521 ( .A1(n14472), .A2(n11880), .B1(n14474), .B2(n11879), .C1(
        n14164), .C2(P2_U3088), .ZN(P2_U3308) );
  INV_X1 U14522 ( .A(n11881), .ZN(n11883) );
  OAI222_X1 U14523 ( .A1(n12490), .A2(P3_U3151), .B1(n13524), .B2(n11883), 
        .C1(n11882), .C2(n13521), .ZN(P3_U3274) );
  OAI22_X1 U14524 ( .A1(n15339), .A2(n11885), .B1(n15294), .B2(n11884), .ZN(
        n11888) );
  MUX2_X1 U14525 ( .A(P1_REG2_REG_5__SCAN_IN), .B(n11886), .S(n15312), .Z(
        n11887) );
  AOI211_X1 U14526 ( .C1(n15319), .C2(n11889), .A(n11888), .B(n11887), .ZN(
        n11890) );
  INV_X1 U14527 ( .A(n11890), .ZN(P1_U3288) );
  XNOR2_X1 U14528 ( .A(n12026), .B(n13615), .ZN(n12040) );
  NAND2_X1 U14529 ( .A1(n13804), .A2(n15891), .ZN(n12038) );
  XNOR2_X1 U14530 ( .A(n12040), .B(n12038), .ZN(n11895) );
  INV_X1 U14531 ( .A(n11895), .ZN(n11891) );
  AOI21_X1 U14532 ( .B1(n11894), .B2(n11891), .A(n13736), .ZN(n11898) );
  NOR3_X1 U14533 ( .A1(n13751), .A2(n11899), .A3(n11892), .ZN(n11897) );
  NAND2_X1 U14534 ( .A1(n11896), .A2(n11895), .ZN(n12042) );
  OAI21_X1 U14535 ( .B1(n11898), .B2(n11897), .A(n12042), .ZN(n11903) );
  OAI22_X1 U14536 ( .A1(n11899), .A2(n13741), .B1(n7482), .B2(n13743), .ZN(
        n12022) );
  AOI22_X1 U14537 ( .A1(n13773), .A2(n12022), .B1(P2_REG3_REG_7__SCAN_IN), 
        .B2(P2_U3088), .ZN(n11900) );
  OAI21_X1 U14538 ( .B1(n12070), .B2(n13775), .A(n11900), .ZN(n11901) );
  AOI21_X1 U14539 ( .B1(n12026), .B2(n13777), .A(n11901), .ZN(n11902) );
  NAND2_X1 U14540 ( .A1(n11903), .A2(n11902), .ZN(P2_U3185) );
  OAI21_X1 U14541 ( .B1(n11905), .B2(n14920), .A(n11904), .ZN(n15811) );
  INV_X1 U14542 ( .A(n15811), .ZN(n11915) );
  INV_X1 U14543 ( .A(n15257), .ZN(n15334) );
  OAI22_X1 U14544 ( .A1(n15312), .A2(n11906), .B1(n14549), .B2(n15294), .ZN(
        n11907) );
  AOI21_X1 U14545 ( .B1(n15336), .B2(n15799), .A(n11907), .ZN(n11908) );
  OAI21_X1 U14546 ( .B1(n14513), .B2(n15334), .A(n11908), .ZN(n11911) );
  OAI211_X1 U14547 ( .C1(n11909), .C2(n15805), .A(n15447), .B(n12254), .ZN(
        n15803) );
  NOR2_X1 U14548 ( .A1(n15803), .A2(n15281), .ZN(n11910) );
  AOI211_X1 U14549 ( .C1(n15291), .C2(n14737), .A(n11911), .B(n11910), .ZN(
        n11914) );
  OR2_X1 U14550 ( .A1(n11912), .A2(n14920), .ZN(n15808) );
  NAND2_X1 U14551 ( .A1(n11912), .A2(n14920), .ZN(n15806) );
  NAND3_X1 U14552 ( .A1(n15808), .A2(n15806), .A3(n15341), .ZN(n11913) );
  OAI211_X1 U14553 ( .C1(n11915), .C2(n15343), .A(n11914), .B(n11913), .ZN(
        P1_U3285) );
  MUX2_X1 U14554 ( .A(P3_REG1_REG_10__SCAN_IN), .B(n11955), .S(n15973), .Z(
        n11916) );
  AOI21_X1 U14555 ( .B1(n13395), .B2(n11917), .A(n11916), .ZN(n11918) );
  OAI21_X1 U14556 ( .B1(n11960), .B2(n13406), .A(n11918), .ZN(P3_U3469) );
  INV_X1 U14557 ( .A(n11919), .ZN(n11921) );
  OAI22_X1 U14558 ( .A1(n12644), .A2(P3_U3151), .B1(SI_22_), .B2(n13521), .ZN(
        n11920) );
  AOI21_X1 U14559 ( .B1(n11921), .B2(n12081), .A(n11920), .ZN(P3_U3273) );
  NAND2_X1 U14560 ( .A1(n11922), .A2(n11923), .ZN(n11997) );
  OAI21_X1 U14561 ( .B1(n11922), .B2(n11923), .A(n11997), .ZN(n11928) );
  INV_X1 U14562 ( .A(n11928), .ZN(n11940) );
  XNOR2_X1 U14563 ( .A(n11924), .B(n11923), .ZN(n11925) );
  NOR2_X1 U14564 ( .A1(n11925), .A2(n14127), .ZN(n11926) );
  AOI211_X1 U14565 ( .C1(n14185), .C2(n11928), .A(n11927), .B(n11926), .ZN(
        n11939) );
  MUX2_X1 U14566 ( .A(n11929), .B(n11939), .S(n14231), .Z(n11936) );
  AOI21_X1 U14567 ( .B1(n11931), .B2(n11930), .A(n15891), .ZN(n11932) );
  AND2_X1 U14568 ( .A1(n11932), .A2(n12010), .ZN(n11937) );
  OAI22_X1 U14569 ( .A1(n14251), .A2(n10197), .B1(n14250), .B2(n11933), .ZN(
        n11934) );
  AOI21_X1 U14570 ( .B1(n14253), .B2(n11937), .A(n11934), .ZN(n11935) );
  OAI211_X1 U14571 ( .C1(n11940), .C2(n14200), .A(n11936), .B(n11935), .ZN(
        P2_U3260) );
  INV_X1 U14572 ( .A(n11937), .ZN(n11938) );
  OAI211_X1 U14573 ( .C1(n11940), .C2(n14303), .A(n11939), .B(n11938), .ZN(
        n11945) );
  OAI22_X1 U14574 ( .A1(n14349), .A2(n10197), .B1(n15912), .B2(n10696), .ZN(
        n11941) );
  AOI21_X1 U14575 ( .B1(n11945), .B2(n15912), .A(n11941), .ZN(n11942) );
  INV_X1 U14576 ( .A(n11942), .ZN(P2_U3504) );
  INV_X1 U14577 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n11943) );
  OAI22_X1 U14578 ( .A1(n14430), .A2(n10197), .B1(n15908), .B2(n11943), .ZN(
        n11944) );
  AOI21_X1 U14579 ( .B1(n11945), .B2(n15908), .A(n11944), .ZN(n11946) );
  INV_X1 U14580 ( .A(n11946), .ZN(P2_U3445) );
  XNOR2_X1 U14581 ( .A(n11947), .B(n8598), .ZN(n11948) );
  AOI222_X1 U14582 ( .A1(n13336), .A2(n11948), .B1(n12944), .B2(n13340), .C1(
        n12946), .C2(n13339), .ZN(n13409) );
  OAI21_X1 U14583 ( .B1(n11950), .B2(n8598), .A(n11949), .ZN(n13408) );
  AOI22_X1 U14584 ( .A1(n13346), .A2(P3_REG2_REG_11__SCAN_IN), .B1(n13345), 
        .B2(n12178), .ZN(n11951) );
  OAI21_X1 U14585 ( .B1(n13348), .B2(n13411), .A(n11951), .ZN(n11952) );
  AOI21_X1 U14586 ( .B1(n13408), .B2(n13324), .A(n11952), .ZN(n11953) );
  OAI21_X1 U14587 ( .B1(n13346), .B2(n13409), .A(n11953), .ZN(P3_U3222) );
  NOR2_X1 U14588 ( .A1(n13348), .A2(n11954), .ZN(n11957) );
  MUX2_X1 U14589 ( .A(n11955), .B(P3_REG2_REG_10__SCAN_IN), .S(n13346), .Z(
        n11956) );
  AOI211_X1 U14590 ( .C1(n13345), .C2(n11958), .A(n11957), .B(n11956), .ZN(
        n11959) );
  OAI21_X1 U14591 ( .B1(n11960), .B2(n13352), .A(n11959), .ZN(P3_U3223) );
  INV_X1 U14592 ( .A(n11961), .ZN(n11965) );
  OAI222_X1 U14593 ( .A1(n15546), .A2(n11963), .B1(n15549), .B2(n11965), .C1(
        P1_U3086), .C2(n11962), .ZN(P1_U3335) );
  OAI222_X1 U14594 ( .A1(n14472), .A2(n11966), .B1(n14474), .B2(n11965), .C1(
        n11964), .C2(P2_U3088), .ZN(P2_U3307) );
  MUX2_X1 U14595 ( .A(n11968), .B(n12949), .S(n11967), .Z(n11969) );
  XOR2_X1 U14596 ( .A(n11970), .B(n11969), .Z(n11978) );
  NAND2_X1 U14597 ( .A1(n12929), .A2(n12949), .ZN(n11972) );
  OAI211_X1 U14598 ( .C1(n12552), .C2(n12931), .A(n11972), .B(n11971), .ZN(
        n11973) );
  AOI21_X1 U14599 ( .B1(n12919), .B2(n11974), .A(n11973), .ZN(n11977) );
  NAND2_X1 U14600 ( .A1(n12934), .A2(n11975), .ZN(n11976) );
  OAI211_X1 U14601 ( .C1(n11978), .C2(n12922), .A(n11977), .B(n11976), .ZN(
        P3_U3161) );
  XNOR2_X1 U14602 ( .A(n12136), .B(P1_REG1_REG_13__SCAN_IN), .ZN(n11982) );
  INV_X1 U14603 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n11980) );
  XNOR2_X1 U14604 ( .A(n15732), .B(P1_REG1_REG_12__SCAN_IN), .ZN(n15730) );
  NOR2_X1 U14605 ( .A1(n11981), .A2(n11982), .ZN(n12135) );
  AOI211_X1 U14606 ( .C1(n11982), .C2(n11981), .A(n15097), .B(n12135), .ZN(
        n11995) );
  OAI21_X1 U14607 ( .B1(n12205), .B2(n11984), .A(n11983), .ZN(n15726) );
  MUX2_X1 U14608 ( .A(P1_REG2_REG_12__SCAN_IN), .B(n12268), .S(n15732), .Z(
        n15729) );
  INV_X1 U14609 ( .A(n15729), .ZN(n11985) );
  NOR2_X1 U14610 ( .A1(n15726), .A2(n11985), .ZN(n11989) );
  INV_X1 U14611 ( .A(n11989), .ZN(n15727) );
  OR2_X1 U14612 ( .A1(n15732), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n11987) );
  MUX2_X1 U14613 ( .A(P1_REG2_REG_13__SCAN_IN), .B(n12317), .S(n12136), .Z(
        n11986) );
  AOI21_X1 U14614 ( .B1(n15727), .B2(n11987), .A(n11986), .ZN(n11990) );
  NAND2_X1 U14615 ( .A1(n12136), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n12131) );
  OAI211_X1 U14616 ( .C1(n12136), .C2(P1_REG2_REG_13__SCAN_IN), .A(n12131), 
        .B(n11987), .ZN(n11988) );
  NOR2_X1 U14617 ( .A1(n11989), .A2(n11988), .ZN(n12133) );
  NOR3_X1 U14618 ( .A1(n11990), .A2(n12133), .A3(n15099), .ZN(n11994) );
  NAND2_X1 U14619 ( .A1(P1_U3086), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n14633)
         );
  NAND2_X1 U14620 ( .A1(n15722), .A2(P1_ADDR_REG_13__SCAN_IN), .ZN(n11991) );
  OAI211_X1 U14621 ( .C1(n15068), .C2(n11992), .A(n14633), .B(n11991), .ZN(
        n11993) );
  OR3_X1 U14622 ( .A1(n11995), .A2(n11994), .A3(n11993), .ZN(P1_U3256) );
  NAND2_X1 U14623 ( .A1(n11997), .A2(n11996), .ZN(n11999) );
  INV_X1 U14624 ( .A(n12000), .ZN(n11998) );
  XNOR2_X1 U14625 ( .A(n11999), .B(n11998), .ZN(n15897) );
  NAND2_X1 U14626 ( .A1(n12001), .A2(n12000), .ZN(n12002) );
  NAND2_X1 U14627 ( .A1(n12003), .A2(n12002), .ZN(n12004) );
  NAND2_X1 U14628 ( .A1(n12004), .A2(n14270), .ZN(n12006) );
  OAI211_X1 U14629 ( .C1(n15897), .C2(n11003), .A(n12006), .B(n12005), .ZN(
        n15902) );
  MUX2_X1 U14630 ( .A(n15902), .B(P2_REG2_REG_6__SCAN_IN), .S(n14210), .Z(
        n12007) );
  INV_X1 U14631 ( .A(n12007), .ZN(n12016) );
  NAND2_X1 U14632 ( .A1(n12010), .A2(n12009), .ZN(n12011) );
  NAND2_X1 U14633 ( .A1(n12011), .A2(n14261), .ZN(n12012) );
  NOR2_X1 U14634 ( .A1(n12008), .A2(n12012), .ZN(n15898) );
  OAI22_X1 U14635 ( .A1(n14251), .A2(n15901), .B1(n14250), .B2(n12013), .ZN(
        n12014) );
  AOI21_X1 U14636 ( .B1(n15898), .B2(n14253), .A(n12014), .ZN(n12015) );
  OAI211_X1 U14637 ( .C1(n15897), .C2(n14200), .A(n12016), .B(n12015), .ZN(
        P2_U3259) );
  NAND2_X1 U14638 ( .A1(P3_U3897), .A2(n13207), .ZN(n12017) );
  OAI21_X1 U14639 ( .B1(P3_U3897), .B2(n12018), .A(n12017), .ZN(P3_U3516) );
  XNOR2_X1 U14640 ( .A(n12019), .B(n12020), .ZN(n12076) );
  XNOR2_X1 U14641 ( .A(n12021), .B(n12020), .ZN(n12023) );
  AOI21_X1 U14642 ( .B1(n12023), .B2(n14270), .A(n12022), .ZN(n12069) );
  INV_X1 U14643 ( .A(n12008), .ZN(n12025) );
  AOI211_X1 U14644 ( .C1(n12026), .C2(n12025), .A(n15891), .B(n12024), .ZN(
        n12073) );
  INV_X1 U14645 ( .A(n12073), .ZN(n12027) );
  OAI211_X1 U14646 ( .C1(n14391), .C2(n12076), .A(n12069), .B(n12027), .ZN(
        n12032) );
  OAI22_X1 U14647 ( .A1(n14349), .A2(n12071), .B1(n15912), .B2(n10698), .ZN(
        n12028) );
  AOI21_X1 U14648 ( .B1(n12032), .B2(n15912), .A(n12028), .ZN(n12029) );
  INV_X1 U14649 ( .A(n12029), .ZN(P2_U3506) );
  INV_X1 U14650 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n12030) );
  OAI22_X1 U14651 ( .A1(n14430), .A2(n12071), .B1(n15908), .B2(n12030), .ZN(
        n12031) );
  AOI21_X1 U14652 ( .B1(n12032), .B2(n15908), .A(n12031), .ZN(n12033) );
  INV_X1 U14653 ( .A(n12033), .ZN(P2_U3451) );
  XNOR2_X1 U14654 ( .A(n14264), .B(n11422), .ZN(n12034) );
  NAND2_X1 U14655 ( .A1(n13803), .A2(n15891), .ZN(n12035) );
  NAND2_X1 U14656 ( .A1(n12034), .A2(n12035), .ZN(n12181) );
  INV_X1 U14657 ( .A(n12034), .ZN(n12037) );
  INV_X1 U14658 ( .A(n12035), .ZN(n12036) );
  NAND2_X1 U14659 ( .A1(n12037), .A2(n12036), .ZN(n12183) );
  NAND2_X1 U14660 ( .A1(n12181), .A2(n12183), .ZN(n12043) );
  INV_X1 U14661 ( .A(n12038), .ZN(n12039) );
  NAND2_X1 U14662 ( .A1(n12040), .A2(n12039), .ZN(n12041) );
  XOR2_X1 U14663 ( .A(n12043), .B(n12182), .Z(n12049) );
  AOI22_X1 U14664 ( .A1(n13802), .A2(n13770), .B1(n13769), .B2(n13804), .ZN(
        n14273) );
  INV_X1 U14665 ( .A(n12044), .ZN(n14262) );
  NAND2_X1 U14666 ( .A1(n13756), .A2(n14262), .ZN(n12045) );
  OAI211_X1 U14667 ( .C1(n13759), .C2(n14273), .A(n12046), .B(n12045), .ZN(
        n12047) );
  AOI21_X1 U14668 ( .B1(n14264), .B2(n13777), .A(n12047), .ZN(n12048) );
  OAI21_X1 U14669 ( .B1(n12049), .B2(n13736), .A(n12048), .ZN(P2_U3193) );
  INV_X1 U14670 ( .A(n12050), .ZN(n12053) );
  OAI222_X1 U14671 ( .A1(n15546), .A2(n12051), .B1(n15549), .B2(n12053), .C1(
        P1_U3086), .C2(n9194), .ZN(P1_U3334) );
  OAI222_X1 U14672 ( .A1(n14472), .A2(n12054), .B1(n14474), .B2(n12053), .C1(
        n12052), .C2(P2_U3088), .ZN(P2_U3306) );
  INV_X1 U14673 ( .A(n12055), .ZN(n12057) );
  OAI222_X1 U14674 ( .A1(n14472), .A2(n12058), .B1(n14474), .B2(n12057), .C1(
        n12056), .C2(P2_U3088), .ZN(P2_U3305) );
  XNOR2_X1 U14675 ( .A(n12059), .B(n12060), .ZN(n12080) );
  XNOR2_X1 U14676 ( .A(n12061), .B(n12060), .ZN(n12062) );
  INV_X1 U14677 ( .A(n13336), .ZN(n13245) );
  OAI222_X1 U14678 ( .A1(n13265), .A2(n12120), .B1(n13267), .B2(n12238), .C1(
        n12062), .C2(n13245), .ZN(n12077) );
  INV_X1 U14679 ( .A(n12116), .ZN(n12243) );
  INV_X1 U14680 ( .A(P3_REG1_REG_12__SCAN_IN), .ZN(n12969) );
  OAI22_X1 U14681 ( .A1(n12243), .A2(n13403), .B1(n15973), .B2(n12969), .ZN(
        n12063) );
  AOI21_X1 U14682 ( .B1(n12077), .B2(n15973), .A(n12063), .ZN(n12064) );
  OAI21_X1 U14683 ( .B1(n12080), .B2(n13406), .A(n12064), .ZN(P3_U3471) );
  AOI22_X1 U14684 ( .A1(n13346), .A2(P3_REG2_REG_12__SCAN_IN), .B1(n13345), 
        .B2(n12240), .ZN(n12065) );
  OAI21_X1 U14685 ( .B1(n12243), .B2(n13348), .A(n12065), .ZN(n12066) );
  AOI21_X1 U14686 ( .B1(n12077), .B2(n13350), .A(n12066), .ZN(n12067) );
  OAI21_X1 U14687 ( .B1(n12080), .B2(n13352), .A(n12067), .ZN(P3_U3221) );
  MUX2_X1 U14688 ( .A(n12069), .B(n12068), .S(n14275), .Z(n12075) );
  OAI22_X1 U14689 ( .A1(n14251), .A2(n12071), .B1(n12070), .B2(n14250), .ZN(
        n12072) );
  AOI21_X1 U14690 ( .B1(n12073), .B2(n14253), .A(n12072), .ZN(n12074) );
  OAI211_X1 U14691 ( .C1(n14256), .C2(n12076), .A(n12075), .B(n12074), .ZN(
        P2_U3258) );
  AOI22_X1 U14692 ( .A1(n12116), .A2(n13480), .B1(P3_REG0_REG_12__SCAN_IN), 
        .B2(n15961), .ZN(n12079) );
  NAND2_X1 U14693 ( .A1(n12077), .A2(n15963), .ZN(n12078) );
  OAI211_X1 U14694 ( .C1(n12080), .C2(n13498), .A(n12079), .B(n12078), .ZN(
        P3_U3426) );
  NAND2_X1 U14695 ( .A1(n12082), .A2(n12081), .ZN(n12083) );
  OAI211_X1 U14696 ( .C1(n12084), .C2(n13521), .A(n12083), .B(n12646), .ZN(
        P3_U3272) );
  NAND2_X1 U14697 ( .A1(n12089), .A2(P3_REG1_REG_10__SCAN_IN), .ZN(n12087) );
  INV_X1 U14698 ( .A(n12975), .ZN(n12100) );
  XOR2_X1 U14699 ( .A(n12970), .B(P3_REG1_REG_11__SCAN_IN), .Z(n12103) );
  NOR2_X1 U14700 ( .A1(n12090), .A2(P3_REG2_REG_11__SCAN_IN), .ZN(n12091) );
  OAI21_X1 U14701 ( .B1(n12091), .B2(n12984), .A(n15916), .ZN(n12102) );
  NAND2_X1 U14702 ( .A1(P3_U3151), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n12174)
         );
  OAI21_X1 U14703 ( .B1(n15925), .B2(n15574), .A(n12174), .ZN(n12099) );
  INV_X1 U14704 ( .A(n12092), .ZN(n12093) );
  MUX2_X1 U14705 ( .A(P3_REG2_REG_11__SCAN_IN), .B(P3_REG1_REG_11__SCAN_IN), 
        .S(n7233), .Z(n12974) );
  XNOR2_X1 U14706 ( .A(n12975), .B(n12974), .ZN(n12095) );
  AOI21_X1 U14707 ( .B1(n12096), .B2(n12095), .A(n12978), .ZN(n12097) );
  NOR2_X1 U14708 ( .A1(n12097), .A2(n13116), .ZN(n12098) );
  AOI211_X1 U14709 ( .C1(n15922), .C2(n12100), .A(n12099), .B(n12098), .ZN(
        n12101) );
  OAI211_X1 U14710 ( .C1(n12103), .C2(n13118), .A(n12102), .B(n12101), .ZN(
        P3_U3193) );
  OAI21_X1 U14711 ( .B1(n12105), .B2(n14932), .A(n12104), .ZN(n15494) );
  XNOR2_X1 U14712 ( .A(n12255), .B(n7119), .ZN(n12107) );
  AND2_X1 U14713 ( .A1(n15478), .A2(n15801), .ZN(n12106) );
  AOI21_X1 U14714 ( .B1(n12107), .B2(n15447), .A(n12106), .ZN(n15500) );
  NAND2_X1 U14715 ( .A1(n15286), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n12108) );
  OAI21_X1 U14716 ( .B1(n15294), .B2(n14512), .A(n12108), .ZN(n12109) );
  AOI21_X1 U14717 ( .B1(n15336), .B2(n15800), .A(n12109), .ZN(n12111) );
  NAND2_X1 U14718 ( .A1(n15495), .A2(n15291), .ZN(n12110) );
  OAI211_X1 U14719 ( .C1(n15500), .C2(n15281), .A(n12111), .B(n12110), .ZN(
        n12114) );
  NAND2_X1 U14720 ( .A1(n12112), .A2(n14932), .ZN(n15496) );
  AND3_X1 U14721 ( .A1(n15497), .A2(n15341), .A3(n15496), .ZN(n12113) );
  AOI211_X1 U14722 ( .C1(n15290), .C2(n15494), .A(n12114), .B(n12113), .ZN(
        n12115) );
  INV_X1 U14723 ( .A(n12115), .ZN(P1_U3283) );
  XNOR2_X1 U14724 ( .A(n12116), .B(n12832), .ZN(n12122) );
  NAND2_X1 U14725 ( .A1(n12117), .A2(n12946), .ZN(n12118) );
  XNOR2_X1 U14726 ( .A(n13411), .B(n12792), .ZN(n12171) );
  NAND2_X1 U14727 ( .A1(n12171), .A2(n12120), .ZN(n12121) );
  XNOR2_X1 U14728 ( .A(n12122), .B(n12944), .ZN(n12232) );
  XNOR2_X1 U14729 ( .A(n12218), .B(n7285), .ZN(n12124) );
  INV_X1 U14730 ( .A(n12124), .ZN(n12123) );
  AND2_X1 U14731 ( .A1(n12124), .A2(n13338), .ZN(n12277) );
  NOR2_X1 U14732 ( .A1(n6724), .A2(n12277), .ZN(n12125) );
  XNOR2_X1 U14733 ( .A(n12278), .B(n12125), .ZN(n12130) );
  NAND2_X1 U14734 ( .A1(n12929), .A2(n12944), .ZN(n12126) );
  NAND2_X1 U14735 ( .A1(P3_U3151), .A2(P3_REG3_REG_13__SCAN_IN), .ZN(n12996)
         );
  OAI211_X1 U14736 ( .C1(n12777), .C2(n12931), .A(n12126), .B(n12996), .ZN(
        n12128) );
  NOR2_X1 U14737 ( .A1(n12218), .A2(n12937), .ZN(n12127) );
  AOI211_X1 U14738 ( .C1(n12225), .C2(n12934), .A(n12128), .B(n12127), .ZN(
        n12129) );
  OAI21_X1 U14739 ( .B1(n12130), .B2(n12922), .A(n12129), .ZN(P3_U3174) );
  INV_X1 U14740 ( .A(n12131), .ZN(n12132) );
  XNOR2_X1 U14741 ( .A(n15036), .B(P1_REG2_REG_14__SCAN_IN), .ZN(n15043) );
  XNOR2_X1 U14742 ( .A(n15044), .B(n15043), .ZN(n12144) );
  XNOR2_X1 U14743 ( .A(n15036), .B(n12134), .ZN(n12138) );
  OAI21_X1 U14744 ( .B1(n12138), .B2(n12137), .A(n15035), .ZN(n12139) );
  NAND2_X1 U14745 ( .A1(n12139), .A2(n15745), .ZN(n12143) );
  INV_X1 U14746 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n12140) );
  NAND2_X1 U14747 ( .A1(P1_U3086), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n14488)
         );
  OAI21_X1 U14748 ( .B1(n15750), .B2(n12140), .A(n14488), .ZN(n12141) );
  AOI21_X1 U14749 ( .B1(n15036), .B2(n15742), .A(n12141), .ZN(n12142) );
  OAI211_X1 U14750 ( .C1(n12144), .C2(n15099), .A(n12143), .B(n12142), .ZN(
        P1_U3257) );
  INV_X1 U14751 ( .A(n11909), .ZN(n12145) );
  OAI211_X1 U14752 ( .C1(n15795), .C2(n12146), .A(n12145), .B(n15447), .ZN(
        n15793) );
  INV_X1 U14753 ( .A(n12147), .ZN(n12157) );
  OAI22_X1 U14754 ( .A1(n14481), .A2(n12723), .B1(n14618), .B2(n15467), .ZN(
        n12156) );
  NOR2_X1 U14755 ( .A1(n12148), .A2(n15465), .ZN(n12154) );
  INV_X1 U14756 ( .A(n12148), .ZN(n12151) );
  NAND3_X1 U14757 ( .A1(n11854), .A2(n15812), .A3(n12149), .ZN(n12150) );
  OAI21_X1 U14758 ( .B1(n12151), .B2(n15465), .A(n12150), .ZN(n12153) );
  INV_X1 U14759 ( .A(n12152), .ZN(n14928) );
  MUX2_X1 U14760 ( .A(n12154), .B(n12153), .S(n14928), .Z(n12155) );
  AOI211_X1 U14761 ( .C1(n12157), .C2(n15812), .A(n12156), .B(n12155), .ZN(
        n15794) );
  MUX2_X1 U14762 ( .A(n12158), .B(n15794), .S(n15312), .Z(n12161) );
  INV_X1 U14763 ( .A(n14480), .ZN(n12159) );
  AOI22_X1 U14764 ( .A1(n15291), .A2(n14733), .B1(n15331), .B2(n12159), .ZN(
        n12160) );
  OAI211_X1 U14765 ( .C1(n15281), .C2(n15793), .A(n12161), .B(n12160), .ZN(
        P1_U3286) );
  NAND2_X1 U14766 ( .A1(n12166), .A2(n12162), .ZN(n12163) );
  OAI211_X1 U14767 ( .C1(n12164), .C2(n15539), .A(n12163), .B(n14959), .ZN(
        P1_U3332) );
  NAND2_X1 U14768 ( .A1(n12166), .A2(n12165), .ZN(n12168) );
  OAI211_X1 U14769 ( .C1(n12169), .C2(n14472), .A(n12168), .B(n12167), .ZN(
        P2_U3304) );
  INV_X1 U14770 ( .A(n12170), .ZN(n12172) );
  NAND2_X1 U14771 ( .A1(n7725), .A2(n12171), .ZN(n12231) );
  OAI21_X1 U14772 ( .B1(n7725), .B2(n12171), .A(n12231), .ZN(n12173) );
  NOR2_X1 U14773 ( .A1(n12173), .A2(n12945), .ZN(n12234) );
  AOI21_X1 U14774 ( .B1(n12945), .B2(n12173), .A(n12234), .ZN(n12180) );
  NAND2_X1 U14775 ( .A1(n12929), .A2(n12946), .ZN(n12175) );
  OAI211_X1 U14776 ( .C1(n12216), .C2(n12931), .A(n12175), .B(n12174), .ZN(
        n12177) );
  NOR2_X1 U14777 ( .A1(n13411), .A2(n12937), .ZN(n12176) );
  AOI211_X1 U14778 ( .C1(n12178), .C2(n12934), .A(n12177), .B(n12176), .ZN(
        n12179) );
  OAI21_X1 U14779 ( .B1(n12180), .B2(n12922), .A(n12179), .ZN(P3_U3176) );
  NAND2_X1 U14780 ( .A1(n12182), .A2(n12181), .ZN(n12184) );
  XNOR2_X1 U14781 ( .A(n14386), .B(n11422), .ZN(n12185) );
  NAND2_X1 U14782 ( .A1(n13802), .A2(n15891), .ZN(n12186) );
  NAND2_X1 U14783 ( .A1(n12185), .A2(n12186), .ZN(n12651) );
  INV_X1 U14784 ( .A(n12185), .ZN(n12188) );
  INV_X1 U14785 ( .A(n12186), .ZN(n12187) );
  NAND2_X1 U14786 ( .A1(n12188), .A2(n12187), .ZN(n12189) );
  NAND2_X1 U14787 ( .A1(n12191), .A2(n12190), .ZN(n12192) );
  AOI21_X1 U14788 ( .B1(n12652), .B2(n12192), .A(n13736), .ZN(n12198) );
  NAND2_X1 U14789 ( .A1(n13777), .A2(n14386), .ZN(n12196) );
  NAND2_X1 U14790 ( .A1(n13803), .A2(n13769), .ZN(n12193) );
  OAI21_X1 U14791 ( .B1(n13731), .B2(n13743), .A(n12193), .ZN(n14245) );
  AOI21_X1 U14792 ( .B1(n13773), .B2(n14245), .A(n12194), .ZN(n12195) );
  OAI211_X1 U14793 ( .C1(n13775), .C2(n14249), .A(n12196), .B(n12195), .ZN(
        n12197) );
  OR2_X1 U14794 ( .A1(n12198), .A2(n12197), .ZN(P2_U3203) );
  NAND2_X1 U14795 ( .A1(n12943), .A2(P3_DATAO_REG_30__SCAN_IN), .ZN(n12199) );
  OAI21_X1 U14796 ( .B1(n12943), .B2(n12427), .A(n12199), .ZN(P3_U3521) );
  OAI21_X1 U14797 ( .B1(n12201), .B2(n7455), .A(n12200), .ZN(n12202) );
  INV_X1 U14798 ( .A(n12202), .ZN(n15493) );
  INV_X1 U14799 ( .A(n12203), .ZN(n12204) );
  AOI211_X1 U14800 ( .C1(n15490), .C2(n12204), .A(n7130), .B(n12272), .ZN(
        n15489) );
  NOR2_X1 U14801 ( .A1(n14753), .A2(n15339), .ZN(n12207) );
  OAI22_X1 U14802 ( .A1(n15312), .A2(n12205), .B1(n14657), .B2(n15294), .ZN(
        n12206) );
  AOI211_X1 U14803 ( .C1(n15489), .C2(n15319), .A(n12207), .B(n12206), .ZN(
        n12213) );
  OAI211_X1 U14804 ( .C1(n12209), .C2(n14934), .A(n12208), .B(n15807), .ZN(
        n12211) );
  OAI22_X1 U14805 ( .A1(n12249), .A2(n12723), .B1(n15466), .B2(n15467), .ZN(
        n14660) );
  INV_X1 U14806 ( .A(n14660), .ZN(n12210) );
  NAND2_X1 U14807 ( .A1(n12211), .A2(n12210), .ZN(n15488) );
  NAND2_X1 U14808 ( .A1(n15488), .A2(n15312), .ZN(n12212) );
  OAI211_X1 U14809 ( .C1(n15493), .C2(n15343), .A(n12213), .B(n12212), .ZN(
        P1_U3282) );
  XNOR2_X1 U14810 ( .A(n12214), .B(n12573), .ZN(n12215) );
  OAI222_X1 U14811 ( .A1(n13267), .A2(n12777), .B1(n13265), .B2(n12216), .C1(
        n12215), .C2(n13245), .ZN(n12224) );
  INV_X1 U14812 ( .A(n12224), .ZN(n12223) );
  XNOR2_X1 U14813 ( .A(n12217), .B(n12454), .ZN(n12227) );
  NAND2_X1 U14814 ( .A1(n12227), .A2(n13485), .ZN(n12220) );
  INV_X1 U14815 ( .A(n12218), .ZN(n12226) );
  AOI22_X1 U14816 ( .A1(n12226), .A2(n13480), .B1(P3_REG0_REG_13__SCAN_IN), 
        .B2(n15961), .ZN(n12219) );
  OAI211_X1 U14817 ( .C1(n15961), .C2(n12223), .A(n12220), .B(n12219), .ZN(
        P3_U3429) );
  NAND2_X1 U14818 ( .A1(n12227), .A2(n13398), .ZN(n12222) );
  AOI22_X1 U14819 ( .A1(n12226), .A2(n13395), .B1(P3_REG1_REG_13__SCAN_IN), 
        .B2(n15970), .ZN(n12221) );
  OAI211_X1 U14820 ( .C1(n12223), .C2(n15970), .A(n12222), .B(n12221), .ZN(
        P3_U3472) );
  AOI21_X1 U14821 ( .B1(n13345), .B2(n12225), .A(n12224), .ZN(n12230) );
  AOI22_X1 U14822 ( .A1(n12226), .A2(n13310), .B1(P3_REG2_REG_13__SCAN_IN), 
        .B2(n13346), .ZN(n12229) );
  NAND2_X1 U14823 ( .A1(n12227), .A2(n13324), .ZN(n12228) );
  OAI211_X1 U14824 ( .C1(n12230), .C2(n13346), .A(n12229), .B(n12228), .ZN(
        P3_U3220) );
  INV_X1 U14825 ( .A(n12231), .ZN(n12233) );
  NOR3_X1 U14826 ( .A1(n12234), .A2(n12233), .A3(n12232), .ZN(n12236) );
  OAI21_X1 U14827 ( .B1(n12236), .B2(n12235), .A(n12924), .ZN(n12242) );
  NAND2_X1 U14828 ( .A1(n12929), .A2(n12945), .ZN(n12237) );
  NAND2_X1 U14829 ( .A1(P3_U3151), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n12979)
         );
  OAI211_X1 U14830 ( .C1(n12238), .C2(n12931), .A(n12237), .B(n12979), .ZN(
        n12239) );
  AOI21_X1 U14831 ( .B1(n12934), .B2(n12240), .A(n12239), .ZN(n12241) );
  OAI211_X1 U14832 ( .C1(n12243), .C2(n12937), .A(n12242), .B(n12241), .ZN(
        P3_U3164) );
  NAND2_X1 U14833 ( .A1(n15808), .A2(n12244), .ZN(n12245) );
  XNOR2_X1 U14834 ( .A(n12245), .B(n14933), .ZN(n12246) );
  NAND2_X1 U14835 ( .A1(n12246), .A2(n15807), .ZN(n12253) );
  OAI21_X1 U14836 ( .B1(n14933), .B2(n12248), .A(n12247), .ZN(n12251) );
  OAI22_X1 U14837 ( .A1(n14618), .A2(n12723), .B1(n12249), .B2(n15467), .ZN(
        n12250) );
  AOI21_X1 U14838 ( .B1(n12251), .B2(n15812), .A(n12250), .ZN(n12252) );
  NAND2_X1 U14839 ( .A1(n12253), .A2(n12252), .ZN(n12286) );
  AOI21_X1 U14840 ( .B1(n12254), .B2(n14742), .A(n7130), .ZN(n12256) );
  NAND2_X1 U14841 ( .A1(n12256), .A2(n12255), .ZN(n12291) );
  OAI21_X1 U14842 ( .B1(n7358), .B2(n15804), .A(n12291), .ZN(n12257) );
  NOR2_X1 U14843 ( .A1(n12286), .A2(n12257), .ZN(n12260) );
  MUX2_X1 U14844 ( .A(n12258), .B(n12260), .S(n15822), .Z(n12259) );
  INV_X1 U14845 ( .A(n12259), .ZN(P1_U3537) );
  INV_X1 U14846 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n12261) );
  MUX2_X1 U14847 ( .A(n12261), .B(n12260), .S(n15815), .Z(n12262) );
  INV_X1 U14848 ( .A(n12262), .ZN(P1_U3486) );
  OAI211_X1 U14849 ( .C1(n12264), .C2(n14937), .A(n15807), .B(n12263), .ZN(
        n15484) );
  OAI21_X1 U14850 ( .B1(n12267), .B2(n12266), .A(n12265), .ZN(n15486) );
  NAND2_X1 U14851 ( .A1(n15486), .A2(n15290), .ZN(n12276) );
  OAI22_X1 U14852 ( .A1(n15312), .A2(n12268), .B1(n14573), .B2(n15294), .ZN(
        n12269) );
  AOI21_X1 U14853 ( .B1(n15257), .B2(n15479), .A(n12269), .ZN(n12270) );
  OAI21_X1 U14854 ( .B1(n14574), .B2(n15255), .A(n12270), .ZN(n12274) );
  OAI211_X1 U14855 ( .C1(n12272), .C2(n12271), .A(n15447), .B(n12320), .ZN(
        n15482) );
  NOR2_X1 U14856 ( .A1(n15482), .A2(n15281), .ZN(n12273) );
  AOI211_X1 U14857 ( .C1(n15291), .C2(n15480), .A(n12274), .B(n12273), .ZN(
        n12275) );
  OAI211_X1 U14858 ( .C1(n15286), .C2(n15484), .A(n12276), .B(n12275), .ZN(
        P1_U3281) );
  XNOR2_X1 U14859 ( .A(n13494), .B(n7285), .ZN(n12775) );
  XNOR2_X1 U14860 ( .A(n12775), .B(n12777), .ZN(n12778) );
  XOR2_X1 U14861 ( .A(n12778), .B(n12779), .Z(n12283) );
  NAND2_X1 U14862 ( .A1(n12929), .A2(n13338), .ZN(n12279) );
  NAND2_X1 U14863 ( .A1(P3_U3151), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n13024)
         );
  OAI211_X1 U14864 ( .C1(n12858), .C2(n12931), .A(n12279), .B(n13024), .ZN(
        n12281) );
  NOR2_X1 U14865 ( .A1(n13494), .A2(n12937), .ZN(n12280) );
  AOI211_X1 U14866 ( .C1(n13344), .C2(n12934), .A(n12281), .B(n12280), .ZN(
        n12282) );
  OAI21_X1 U14867 ( .B1(n12283), .B2(n12922), .A(n12282), .ZN(P3_U3155) );
  NAND2_X1 U14868 ( .A1(P3_U3897), .A2(n13169), .ZN(n12284) );
  OAI21_X1 U14869 ( .B1(P3_U3897), .B2(n12285), .A(n12284), .ZN(P3_U3519) );
  MUX2_X1 U14870 ( .A(n12286), .B(P1_REG2_REG_9__SCAN_IN), .S(n15286), .Z(
        n12287) );
  INV_X1 U14871 ( .A(n12287), .ZN(n12290) );
  INV_X1 U14872 ( .A(n14617), .ZN(n12288) );
  AOI22_X1 U14873 ( .A1(n14742), .A2(n15291), .B1(n15331), .B2(n12288), .ZN(
        n12289) );
  OAI211_X1 U14874 ( .C1(n12291), .C2(n15281), .A(n12290), .B(n12289), .ZN(
        P1_U3284) );
  INV_X1 U14875 ( .A(n8561), .ZN(n12295) );
  INV_X1 U14876 ( .A(n12292), .ZN(n12293) );
  OAI222_X1 U14877 ( .A1(n12295), .A2(P3_U3151), .B1(n13521), .B2(n12294), 
        .C1(n13524), .C2(n12293), .ZN(P3_U3271) );
  OR2_X1 U14878 ( .A1(n12305), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n12296) );
  INV_X1 U14879 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n12298) );
  NAND2_X1 U14880 ( .A1(n12299), .A2(n12298), .ZN(n12300) );
  NAND2_X1 U14881 ( .A1(n15849), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n12301) );
  AND2_X1 U14882 ( .A1(n12300), .A2(n12301), .ZN(n15852) );
  NAND2_X1 U14883 ( .A1(n15851), .A2(n12301), .ZN(n13881) );
  XNOR2_X1 U14884 ( .A(n13880), .B(P2_REG2_REG_14__SCAN_IN), .ZN(n12310) );
  INV_X1 U14885 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n12303) );
  NAND2_X1 U14886 ( .A1(P2_U3088), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n13574)
         );
  OAI21_X1 U14887 ( .B1(n15857), .B2(n12303), .A(n13574), .ZN(n12308) );
  XNOR2_X1 U14888 ( .A(n15849), .B(P2_REG1_REG_13__SCAN_IN), .ZN(n15846) );
  XNOR2_X1 U14889 ( .A(n13885), .B(P2_REG1_REG_14__SCAN_IN), .ZN(n12306) );
  AOI211_X1 U14890 ( .C1(n6721), .C2(n12306), .A(n15860), .B(n13884), .ZN(
        n12307) );
  AOI211_X1 U14891 ( .C1(n15850), .C2(n13885), .A(n12308), .B(n12307), .ZN(
        n12309) );
  OAI21_X1 U14892 ( .B1(n12310), .B2(n15823), .A(n12309), .ZN(P2_U3228) );
  OAI211_X1 U14893 ( .C1(n12312), .C2(n14939), .A(n15807), .B(n12311), .ZN(
        n15473) );
  OAI21_X1 U14894 ( .B1(n12316), .B2(n12315), .A(n12314), .ZN(n15476) );
  NAND2_X1 U14895 ( .A1(n15476), .A2(n15290), .ZN(n12326) );
  OAI22_X1 U14896 ( .A1(n15312), .A2(n12317), .B1(n14634), .B2(n15294), .ZN(
        n12318) );
  AOI21_X1 U14897 ( .B1(n15336), .B2(n14965), .A(n12318), .ZN(n12319) );
  OAI21_X1 U14898 ( .B1(n15468), .B2(n15334), .A(n12319), .ZN(n12324) );
  NAND2_X1 U14899 ( .A1(n12320), .A2(n15471), .ZN(n12321) );
  NAND2_X1 U14900 ( .A1(n12332), .A2(n12321), .ZN(n15474) );
  INV_X1 U14901 ( .A(n15329), .ZN(n12322) );
  NOR2_X1 U14902 ( .A1(n15474), .A2(n12322), .ZN(n12323) );
  AOI211_X1 U14903 ( .C1(n15291), .C2(n15471), .A(n12324), .B(n12323), .ZN(
        n12325) );
  OAI211_X1 U14904 ( .C1(n15286), .C2(n15473), .A(n12326), .B(n12325), .ZN(
        P1_U3280) );
  XNOR2_X1 U14905 ( .A(n12327), .B(n14941), .ZN(n15464) );
  INV_X1 U14906 ( .A(n12329), .ZN(n12330) );
  AOI21_X1 U14907 ( .B1(n14941), .B2(n12331), .A(n12330), .ZN(n15462) );
  AOI21_X1 U14908 ( .B1(n12332), .B2(n14772), .A(n7130), .ZN(n12333) );
  NAND2_X1 U14909 ( .A1(n12333), .A2(n15326), .ZN(n15460) );
  OAI22_X1 U14910 ( .A1(n15312), .A2(n15041), .B1(n14489), .B2(n15294), .ZN(
        n12334) );
  AOI21_X1 U14911 ( .B1(n15257), .B2(n15458), .A(n12334), .ZN(n12335) );
  OAI21_X1 U14912 ( .B1(n14572), .B2(n15255), .A(n12335), .ZN(n12336) );
  AOI21_X1 U14913 ( .B1(n14772), .B2(n15291), .A(n12336), .ZN(n12337) );
  OAI21_X1 U14914 ( .B1(n15460), .B2(n15281), .A(n12337), .ZN(n12338) );
  AOI21_X1 U14915 ( .B1(n15462), .B2(n15290), .A(n12338), .ZN(n12339) );
  OAI21_X1 U14916 ( .B1(n15301), .B2(n15464), .A(n12339), .ZN(P1_U3279) );
  NAND2_X1 U14917 ( .A1(n12340), .A2(n12347), .ZN(n12341) );
  NAND2_X1 U14918 ( .A1(n12341), .A2(n13336), .ZN(n12342) );
  OR2_X1 U14919 ( .A1(n12343), .A2(n12342), .ZN(n12346) );
  AOI22_X1 U14920 ( .A1(n13340), .A2(n12344), .B1(n12953), .B2(n13339), .ZN(
        n12345) );
  NAND2_X1 U14921 ( .A1(n12346), .A2(n12345), .ZN(n15936) );
  MUX2_X1 U14922 ( .A(n15936), .B(P3_REG2_REG_3__SCAN_IN), .S(n13346), .Z(
        n12355) );
  OR2_X1 U14923 ( .A1(n11265), .A2(n12347), .ZN(n12348) );
  NAND2_X1 U14924 ( .A1(n12349), .A2(n12348), .ZN(n15937) );
  NAND2_X1 U14925 ( .A1(n15937), .A2(n13324), .ZN(n12353) );
  AOI22_X1 U14926 ( .A1(n13310), .A2(n12351), .B1(n13345), .B2(n12350), .ZN(
        n12352) );
  NAND2_X1 U14927 ( .A1(n12353), .A2(n12352), .ZN(n12354) );
  OR2_X1 U14928 ( .A1(n12355), .A2(n12354), .ZN(P3_U3230) );
  XNOR2_X1 U14929 ( .A(n12356), .B(n12358), .ZN(n14364) );
  XOR2_X1 U14930 ( .A(n12358), .B(n12357), .Z(n12359) );
  AOI22_X1 U14931 ( .A1(n13769), .A2(n13799), .B1(n13797), .B2(n13770), .ZN(
        n13707) );
  OAI21_X1 U14932 ( .B1(n12359), .B2(n14127), .A(n13707), .ZN(n14360) );
  AOI21_X1 U14933 ( .B1(n12360), .B2(n14362), .A(n15891), .ZN(n12361) );
  AND2_X1 U14934 ( .A1(n12361), .A2(n14175), .ZN(n14361) );
  NAND2_X1 U14935 ( .A1(n14361), .A2(n14253), .ZN(n12365) );
  NAND2_X1 U14936 ( .A1(n14210), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n12362) );
  OAI21_X1 U14937 ( .B1(n14250), .B2(n13706), .A(n12362), .ZN(n12363) );
  AOI21_X1 U14938 ( .B1(n14362), .B2(n14265), .A(n12363), .ZN(n12364) );
  NAND2_X1 U14939 ( .A1(n12365), .A2(n12364), .ZN(n12366) );
  AOI21_X1 U14940 ( .B1(n14360), .B2(n14231), .A(n12366), .ZN(n12367) );
  OAI21_X1 U14941 ( .B1(n14364), .B2(n14256), .A(n12367), .ZN(P2_U3252) );
  INV_X1 U14942 ( .A(n13614), .ZN(n13783) );
  NOR2_X1 U14943 ( .A1(n13956), .A2(n10190), .ZN(n12368) );
  INV_X1 U14944 ( .A(n13954), .ZN(n12370) );
  NAND3_X1 U14945 ( .A1(n13956), .A2(n10190), .A3(n12370), .ZN(n12369) );
  OAI211_X1 U14946 ( .C1(n13956), .C2(n12370), .A(n12369), .B(n14396), .ZN(
        n12371) );
  INV_X1 U14947 ( .A(n12371), .ZN(n12372) );
  INV_X1 U14948 ( .A(n12375), .ZN(n12376) );
  NAND2_X1 U14949 ( .A1(n12378), .A2(P2_B_REG_SCAN_IN), .ZN(n12379) );
  NAND2_X1 U14950 ( .A1(n13770), .A2(n12379), .ZN(n12391) );
  OAI22_X1 U14951 ( .A1(n13614), .A2(n13741), .B1(n12380), .B2(n12391), .ZN(
        n12381) );
  INV_X1 U14952 ( .A(n14387), .ZN(n15900) );
  OAI21_X1 U14953 ( .B1(n13962), .B2(n15900), .A(n13958), .ZN(n12386) );
  INV_X1 U14954 ( .A(n12386), .ZN(n12387) );
  INV_X1 U14955 ( .A(n14842), .ZN(n12772) );
  OAI222_X1 U14956 ( .A1(n15539), .A2(n14843), .B1(P1_U3086), .B2(n12389), 
        .C1(n15549), .C2(n12772), .ZN(P1_U3325) );
  INV_X1 U14957 ( .A(n14349), .ZN(n14377) );
  INV_X1 U14958 ( .A(n12391), .ZN(n12392) );
  NAND2_X1 U14959 ( .A1(n13781), .A2(n12392), .ZN(n14280) );
  NAND2_X1 U14960 ( .A1(n13948), .A2(n14280), .ZN(n12768) );
  INV_X1 U14961 ( .A(n12393), .ZN(P2_U3530) );
  OR2_X1 U14962 ( .A1(n12394), .A2(n14349), .ZN(n12396) );
  OR2_X1 U14963 ( .A1(n13423), .A2(n13157), .ZN(n12440) );
  NAND2_X1 U14964 ( .A1(n8517), .A2(P3_REG0_REG_31__SCAN_IN), .ZN(n12402) );
  NAND2_X1 U14965 ( .A1(n12398), .A2(P3_REG1_REG_31__SCAN_IN), .ZN(n12401) );
  NAND2_X1 U14966 ( .A1(n12399), .A2(P3_REG2_REG_31__SCAN_IN), .ZN(n12400) );
  INV_X1 U14967 ( .A(n12404), .ZN(n12405) );
  NAND2_X1 U14968 ( .A1(n12406), .A2(n12405), .ZN(n12408) );
  XNOR2_X1 U14969 ( .A(n12774), .B(P2_DATAO_REG_30__SCAN_IN), .ZN(n12409) );
  XNOR2_X1 U14970 ( .A(n12416), .B(n12409), .ZN(n12648) );
  NAND2_X1 U14971 ( .A1(n12648), .A2(n12422), .ZN(n12412) );
  NAND2_X1 U14972 ( .A1(n12410), .A2(SI_30_), .ZN(n12411) );
  NAND2_X1 U14973 ( .A1(n13147), .A2(n12427), .ZN(n12617) );
  NAND2_X1 U14974 ( .A1(n13423), .A2(n13157), .ZN(n12413) );
  INV_X1 U14975 ( .A(n12621), .ZN(n12414) );
  AOI211_X1 U14976 ( .C1(n13144), .C2(n13147), .A(n6525), .B(n12414), .ZN(
        n12426) );
  NAND2_X1 U14977 ( .A1(n12774), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n12415) );
  NAND2_X1 U14978 ( .A1(n12416), .A2(n12415), .ZN(n12418) );
  NAND2_X1 U14979 ( .A1(n14843), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n12417) );
  NAND2_X1 U14980 ( .A1(n12418), .A2(n12417), .ZN(n12421) );
  XNOR2_X1 U14981 ( .A(n12419), .B(P2_DATAO_REG_31__SCAN_IN), .ZN(n12420) );
  XNOR2_X1 U14982 ( .A(n12421), .B(n12420), .ZN(n13502) );
  NAND2_X1 U14983 ( .A1(n13502), .A2(n12422), .ZN(n12425) );
  NAND2_X1 U14984 ( .A1(n12423), .A2(SI_31_), .ZN(n12424) );
  NAND2_X1 U14985 ( .A1(n12426), .A2(n12630), .ZN(n12434) );
  NOR2_X1 U14986 ( .A1(n13147), .A2(n12427), .ZN(n12439) );
  NOR2_X1 U14987 ( .A1(n12439), .A2(n13144), .ZN(n12436) );
  INV_X1 U14988 ( .A(n12436), .ZN(n12428) );
  NAND3_X1 U14989 ( .A1(n12428), .A2(n13128), .A3(n12460), .ZN(n12432) );
  INV_X1 U14990 ( .A(n13144), .ZN(n12938) );
  OAI211_X1 U14991 ( .C1(n12938), .C2(n13147), .A(n13419), .B(n6525), .ZN(
        n12430) );
  AND2_X1 U14992 ( .A1(n12430), .A2(n12429), .ZN(n12431) );
  OAI21_X1 U14993 ( .B1(n12436), .B2(n13419), .A(n6525), .ZN(n12437) );
  AOI21_X1 U14994 ( .B1(n12621), .B2(n12438), .A(n12437), .ZN(n12639) );
  INV_X1 U14995 ( .A(n12439), .ZN(n12624) );
  NAND2_X1 U14996 ( .A1(n12624), .A2(n12440), .ZN(n12462) );
  INV_X1 U14997 ( .A(n13185), .ZN(n12606) );
  INV_X1 U14998 ( .A(n12469), .ZN(n12442) );
  NAND2_X1 U14999 ( .A1(n12467), .A2(n12442), .ZN(n13232) );
  XNOR2_X1 U15000 ( .A(n13251), .B(n13268), .ZN(n13242) );
  INV_X1 U15001 ( .A(n13325), .ZN(n12487) );
  OR2_X1 U15002 ( .A1(n12487), .A2(n13334), .ZN(n12485) );
  NOR4_X1 U15003 ( .A1(n12445), .A2(n12511), .A3(n12521), .A4(n12444), .ZN(
        n12449) );
  NAND4_X1 U15004 ( .A1(n12449), .A2(n12535), .A3(n12448), .A4(n12447), .ZN(
        n12451) );
  INV_X1 U15005 ( .A(n12450), .ZN(n12541) );
  NOR4_X1 U15006 ( .A1(n12451), .A2(n12558), .A3(n12541), .A4(n12550), .ZN(
        n12452) );
  NAND4_X1 U15007 ( .A1(n12454), .A2(n8598), .A3(n12453), .A4(n12452), .ZN(
        n12455) );
  NOR4_X1 U15008 ( .A1(n12584), .A2(n13311), .A3(n12485), .A4(n12455), .ZN(
        n12456) );
  NAND4_X1 U15009 ( .A1(n6861), .A2(n6989), .A3(n13279), .A4(n12456), .ZN(
        n12457) );
  NOR4_X1 U15010 ( .A1(n13223), .A2(n13232), .A3(n13242), .A4(n12457), .ZN(
        n12458) );
  NAND4_X1 U15011 ( .A1(n12606), .A2(n8608), .A3(n13198), .A4(n12458), .ZN(
        n12459) );
  NAND2_X1 U15012 ( .A1(n12460), .A2(n13144), .ZN(n12628) );
  INV_X1 U15013 ( .A(n12462), .ZN(n12619) );
  NAND3_X1 U15014 ( .A1(n13358), .A2(n12626), .A3(n13181), .ZN(n12614) );
  MUX2_X1 U15015 ( .A(n12464), .B(n12463), .S(n12598), .Z(n12605) );
  MUX2_X1 U15016 ( .A(n12466), .B(n12465), .S(n12598), .Z(n12603) );
  INV_X1 U15017 ( .A(n12467), .ZN(n12468) );
  MUX2_X1 U15018 ( .A(n12469), .B(n12468), .S(n12598), .Z(n12470) );
  NOR2_X1 U15019 ( .A1(n13223), .A2(n12470), .ZN(n12602) );
  MUX2_X1 U15020 ( .A(n6596), .B(n12471), .S(n12626), .Z(n12593) );
  INV_X1 U15021 ( .A(n13242), .ZN(n13240) );
  MUX2_X1 U15022 ( .A(n12473), .B(n12472), .S(n12626), .Z(n12592) );
  OAI211_X1 U15023 ( .C1(n13289), .C2(n13286), .A(n12474), .B(n13258), .ZN(
        n12478) );
  INV_X1 U15024 ( .A(n12474), .ZN(n12476) );
  OAI211_X1 U15025 ( .C1(n12476), .C2(n12475), .A(n12587), .B(n13255), .ZN(
        n12477) );
  MUX2_X1 U15026 ( .A(n12478), .B(n12477), .S(n12626), .Z(n12590) );
  INV_X1 U15027 ( .A(n12485), .ZN(n12575) );
  OAI21_X1 U15028 ( .B1(n12573), .B2(n12567), .A(n12479), .ZN(n12483) );
  OAI211_X1 U15029 ( .C1(n12487), .C2(n12481), .A(n12580), .B(n12480), .ZN(
        n12482) );
  AOI21_X1 U15030 ( .B1(n12575), .B2(n12483), .A(n12482), .ZN(n12582) );
  NOR2_X1 U15031 ( .A1(n12485), .A2(n12484), .ZN(n12489) );
  OAI211_X1 U15032 ( .C1(n12487), .C2(n6547), .A(n12583), .B(n12486), .ZN(
        n12488) );
  OAI21_X1 U15033 ( .B1(n12489), .B2(n12488), .A(n12598), .ZN(n12579) );
  AOI21_X1 U15034 ( .B1(n12495), .B2(n12644), .A(n12490), .ZN(n12492) );
  MUX2_X1 U15035 ( .A(n12626), .B(n12492), .S(n12491), .Z(n12503) );
  OAI21_X1 U15036 ( .B1(n12494), .B2(n12493), .A(n12496), .ZN(n12502) );
  INV_X1 U15037 ( .A(n12495), .ZN(n12498) );
  INV_X1 U15038 ( .A(n12496), .ZN(n12497) );
  MUX2_X1 U15039 ( .A(n12498), .B(n12497), .S(n12626), .Z(n12499) );
  INV_X1 U15040 ( .A(n12499), .ZN(n12500) );
  OAI211_X1 U15041 ( .C1(n12503), .C2(n12502), .A(n12501), .B(n12500), .ZN(
        n12508) );
  NAND2_X1 U15042 ( .A1(n12512), .A2(n12504), .ZN(n12505) );
  NAND2_X1 U15043 ( .A1(n12505), .A2(n12598), .ZN(n12507) );
  INV_X1 U15044 ( .A(n12510), .ZN(n12506) );
  AOI21_X1 U15045 ( .B1(n12508), .B2(n12507), .A(n12506), .ZN(n12517) );
  AOI21_X1 U15046 ( .B1(n12510), .B2(n12509), .A(n12598), .ZN(n12516) );
  INV_X1 U15047 ( .A(n12511), .ZN(n12515) );
  INV_X1 U15048 ( .A(n12512), .ZN(n12513) );
  NAND2_X1 U15049 ( .A1(n12513), .A2(n12626), .ZN(n12514) );
  OAI211_X1 U15050 ( .C1(n12517), .C2(n12516), .A(n12515), .B(n12514), .ZN(
        n12526) );
  INV_X1 U15051 ( .A(n12518), .ZN(n12519) );
  NOR2_X1 U15052 ( .A1(n12522), .A2(n12521), .ZN(n12525) );
  AOI21_X1 U15053 ( .B1(n12532), .B2(n12523), .A(n12598), .ZN(n12524) );
  AOI21_X1 U15054 ( .B1(n12526), .B2(n12525), .A(n12524), .ZN(n12531) );
  INV_X1 U15055 ( .A(n12528), .ZN(n12530) );
  AND2_X1 U15056 ( .A1(n12528), .A2(n12527), .ZN(n12529) );
  OAI22_X1 U15057 ( .A1(n12531), .A2(n12530), .B1(n12626), .B2(n12529), .ZN(
        n12536) );
  INV_X1 U15058 ( .A(n12532), .ZN(n12533) );
  NAND2_X1 U15059 ( .A1(n12533), .A2(n12598), .ZN(n12534) );
  NAND3_X1 U15060 ( .A1(n12536), .A2(n12535), .A3(n12534), .ZN(n12544) );
  INV_X1 U15061 ( .A(n12537), .ZN(n12540) );
  INV_X1 U15062 ( .A(n12538), .ZN(n12539) );
  MUX2_X1 U15063 ( .A(n12540), .B(n12539), .S(n12626), .Z(n12542) );
  NOR2_X1 U15064 ( .A1(n12542), .A2(n12541), .ZN(n12543) );
  NAND2_X1 U15065 ( .A1(n12544), .A2(n12543), .ZN(n12557) );
  INV_X1 U15066 ( .A(n12545), .ZN(n12548) );
  INV_X1 U15067 ( .A(n12546), .ZN(n12547) );
  MUX2_X1 U15068 ( .A(n12548), .B(n12547), .S(n12626), .Z(n12549) );
  NOR2_X1 U15069 ( .A1(n12550), .A2(n12549), .ZN(n12556) );
  AND2_X1 U15070 ( .A1(n12551), .A2(n12598), .ZN(n12554) );
  NOR2_X1 U15071 ( .A1(n12551), .A2(n12598), .ZN(n12553) );
  MUX2_X1 U15072 ( .A(n12554), .B(n12553), .S(n12552), .Z(n12555) );
  AOI21_X1 U15073 ( .B1(n12557), .B2(n12556), .A(n12555), .ZN(n12559) );
  INV_X1 U15074 ( .A(n12560), .ZN(n12563) );
  INV_X1 U15075 ( .A(n12561), .ZN(n12562) );
  MUX2_X1 U15076 ( .A(n12563), .B(n12562), .S(n12626), .Z(n12564) );
  NOR2_X1 U15077 ( .A1(n12565), .A2(n12564), .ZN(n12569) );
  AOI21_X1 U15078 ( .B1(n12567), .B2(n12566), .A(n12626), .ZN(n12568) );
  INV_X1 U15079 ( .A(n12571), .ZN(n12576) );
  NAND2_X1 U15080 ( .A1(n13411), .A2(n12945), .ZN(n12570) );
  AOI21_X1 U15081 ( .B1(n12571), .B2(n12570), .A(n12598), .ZN(n12572) );
  NOR2_X1 U15082 ( .A1(n12573), .A2(n12572), .ZN(n12574) );
  OAI211_X1 U15083 ( .C1(n12577), .C2(n12576), .A(n12575), .B(n12574), .ZN(
        n12578) );
  NOR2_X1 U15084 ( .A1(n13289), .A2(n12584), .ZN(n12585) );
  MUX2_X1 U15085 ( .A(n13258), .B(n12587), .S(n12598), .Z(n12588) );
  OAI211_X1 U15086 ( .C1(n12590), .C2(n12589), .A(n6861), .B(n12588), .ZN(
        n12591) );
  INV_X1 U15087 ( .A(n13232), .ZN(n12594) );
  NAND2_X1 U15088 ( .A1(n12595), .A2(n12594), .ZN(n12601) );
  INV_X1 U15089 ( .A(n12597), .ZN(n12599) );
  MUX2_X1 U15090 ( .A(n8607), .B(n12599), .S(n12598), .Z(n12600) );
  OR3_X1 U15091 ( .A1(n12920), .A2(n12626), .A3(n13196), .ZN(n12607) );
  INV_X1 U15092 ( .A(n12608), .ZN(n12609) );
  NAND2_X1 U15093 ( .A1(n12611), .A2(n12609), .ZN(n12610) );
  MUX2_X1 U15094 ( .A(n12611), .B(n12610), .S(n12626), .Z(n12612) );
  INV_X1 U15095 ( .A(n12617), .ZN(n12618) );
  AOI21_X1 U15096 ( .B1(n12619), .B2(n12623), .A(n12618), .ZN(n12627) );
  INV_X1 U15097 ( .A(n12620), .ZN(n12622) );
  OAI21_X1 U15098 ( .B1(n12623), .B2(n12622), .A(n12621), .ZN(n12625) );
  INV_X1 U15099 ( .A(n12628), .ZN(n12629) );
  NAND3_X1 U15100 ( .A1(n12642), .A2(n12641), .A3(n6527), .ZN(n12643) );
  OAI211_X1 U15101 ( .C1(n12644), .C2(n12646), .A(n12643), .B(P3_B_REG_SCAN_IN), .ZN(n12645) );
  OAI21_X1 U15102 ( .B1(n12647), .B2(n12646), .A(n12645), .ZN(P3_U3296) );
  INV_X1 U15103 ( .A(n12648), .ZN(n12650) );
  OAI222_X1 U15104 ( .A1(n13524), .A2(n12650), .B1(n8061), .B2(P3_U3151), .C1(
        n12649), .C2(n13521), .ZN(P3_U3265) );
  XNOR2_X1 U15105 ( .A(n14379), .B(n13615), .ZN(n12653) );
  NOR2_X1 U15106 ( .A1(n13731), .A2(n14261), .ZN(n12654) );
  XNOR2_X1 U15107 ( .A(n12653), .B(n12654), .ZN(n13598) );
  INV_X1 U15108 ( .A(n12653), .ZN(n12656) );
  INV_X1 U15109 ( .A(n12654), .ZN(n12655) );
  XNOR2_X1 U15110 ( .A(n14443), .B(n13615), .ZN(n12659) );
  NAND2_X1 U15111 ( .A1(n13800), .A2(n15891), .ZN(n12657) );
  XNOR2_X1 U15112 ( .A(n12659), .B(n12657), .ZN(n13728) );
  INV_X1 U15113 ( .A(n12657), .ZN(n12658) );
  NAND2_X1 U15114 ( .A1(n12659), .A2(n12658), .ZN(n12660) );
  XNOR2_X1 U15115 ( .A(n14197), .B(n11422), .ZN(n12662) );
  NAND2_X1 U15116 ( .A1(n13799), .A2(n15891), .ZN(n12663) );
  NAND2_X1 U15117 ( .A1(n12662), .A2(n12663), .ZN(n13638) );
  NAND2_X1 U15118 ( .A1(n13640), .A2(n13638), .ZN(n12666) );
  INV_X1 U15119 ( .A(n12662), .ZN(n12665) );
  INV_X1 U15120 ( .A(n12663), .ZN(n12664) );
  NAND2_X1 U15121 ( .A1(n12665), .A2(n12664), .ZN(n13639) );
  XNOR2_X1 U15122 ( .A(n14362), .B(n13615), .ZN(n12667) );
  AND2_X1 U15123 ( .A1(n13798), .A2(n14307), .ZN(n12668) );
  NAND2_X1 U15124 ( .A1(n12667), .A2(n12668), .ZN(n12671) );
  INV_X1 U15125 ( .A(n12667), .ZN(n13577) );
  INV_X1 U15126 ( .A(n12668), .ZN(n12669) );
  NAND2_X1 U15127 ( .A1(n13577), .A2(n12669), .ZN(n12670) );
  AND2_X1 U15128 ( .A1(n12671), .A2(n12670), .ZN(n13705) );
  XNOR2_X1 U15129 ( .A(n14435), .B(n13615), .ZN(n12673) );
  NAND2_X1 U15130 ( .A1(n13797), .A2(n15891), .ZN(n12674) );
  XNOR2_X1 U15131 ( .A(n12673), .B(n12674), .ZN(n13580) );
  INV_X1 U15132 ( .A(n12673), .ZN(n12675) );
  NAND2_X1 U15133 ( .A1(n12675), .A2(n12674), .ZN(n12676) );
  AND2_X1 U15134 ( .A1(n13795), .A2(n14307), .ZN(n13663) );
  XNOR2_X1 U15135 ( .A(n14148), .B(n13615), .ZN(n13675) );
  OAI22_X1 U15136 ( .A1(n13664), .A2(n13665), .B1(n13663), .B2(n13675), .ZN(
        n12681) );
  AOI21_X1 U15137 ( .B1(n13664), .B2(n13665), .A(n13663), .ZN(n12679) );
  INV_X1 U15138 ( .A(n13675), .ZN(n12678) );
  NAND3_X1 U15139 ( .A1(n13664), .A2(n13665), .A3(n13663), .ZN(n12677) );
  NAND2_X1 U15140 ( .A1(n13794), .A2(n15891), .ZN(n12683) );
  XNOR2_X1 U15141 ( .A(n12682), .B(n12683), .ZN(n13676) );
  OAI211_X1 U15142 ( .C1(n12679), .C2(n12678), .A(n12677), .B(n13676), .ZN(
        n12680) );
  INV_X1 U15143 ( .A(n12682), .ZN(n12684) );
  NAND2_X1 U15144 ( .A1(n12684), .A2(n12683), .ZN(n12685) );
  XNOR2_X1 U15145 ( .A(n14335), .B(n13615), .ZN(n12695) );
  NOR2_X1 U15146 ( .A1(n12686), .A2(n14261), .ZN(n12687) );
  NAND2_X1 U15147 ( .A1(n12695), .A2(n12687), .ZN(n12693) );
  INV_X1 U15148 ( .A(n12695), .ZN(n12689) );
  INV_X1 U15149 ( .A(n12687), .ZN(n12688) );
  NAND2_X1 U15150 ( .A1(n12689), .A2(n12688), .ZN(n12690) );
  NAND2_X1 U15151 ( .A1(n12693), .A2(n12690), .ZN(n13737) );
  INV_X1 U15152 ( .A(n13737), .ZN(n12691) );
  XNOR2_X1 U15153 ( .A(n14097), .B(n13615), .ZN(n13531) );
  NAND2_X1 U15154 ( .A1(n13792), .A2(n15891), .ZN(n13532) );
  XNOR2_X1 U15155 ( .A(n13531), .B(n13532), .ZN(n12697) );
  NAND3_X1 U15156 ( .A1(n12695), .A2(n13765), .A3(n13793), .ZN(n12696) );
  OAI21_X1 U15157 ( .B1(n13739), .B2(n13736), .A(n12696), .ZN(n12699) );
  INV_X1 U15158 ( .A(n12697), .ZN(n12698) );
  NAND2_X1 U15159 ( .A1(n12699), .A2(n12698), .ZN(n12703) );
  NOR2_X1 U15160 ( .A1(n13775), .A2(n14098), .ZN(n12701) );
  AOI22_X1 U15161 ( .A1(n13791), .A2(n13770), .B1(n13793), .B2(n13769), .ZN(
        n14092) );
  NAND2_X1 U15162 ( .A1(P2_U3088), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n13943)
         );
  OAI21_X1 U15163 ( .B1(n14092), .B2(n13759), .A(n13943), .ZN(n12700) );
  AOI211_X1 U15164 ( .C1(n14097), .C2(n13777), .A(n12701), .B(n12700), .ZN(
        n12702) );
  OAI211_X1 U15165 ( .C1(n13699), .C2(n13736), .A(n12703), .B(n12702), .ZN(
        P2_U3191) );
  NAND2_X1 U15166 ( .A1(n15191), .A2(n12704), .ZN(n12706) );
  OAI211_X1 U15167 ( .C1(n15187), .C2(n15384), .A(n12706), .B(n12705), .ZN(
        n12707) );
  INV_X1 U15168 ( .A(n12707), .ZN(n12708) );
  NAND2_X1 U15169 ( .A1(n15187), .A2(n15384), .ZN(n12709) );
  XNOR2_X1 U15170 ( .A(n15379), .B(n14816), .ZN(n14951) );
  NAND2_X1 U15171 ( .A1(n15379), .A2(n14816), .ZN(n12713) );
  OAI21_X2 U15172 ( .B1(n15166), .B2(n14951), .A(n12713), .ZN(n15157) );
  OR2_X2 U15173 ( .A1(n15157), .A2(n15158), .ZN(n15155) );
  NAND2_X1 U15174 ( .A1(n7127), .A2(n14963), .ZN(n12710) );
  NAND2_X1 U15175 ( .A1(n15155), .A2(n12710), .ZN(n12712) );
  NAND2_X1 U15176 ( .A1(n14868), .A2(n14867), .ZN(n12746) );
  OR2_X1 U15177 ( .A1(n14868), .A2(n14867), .ZN(n12711) );
  NAND2_X1 U15178 ( .A1(n12712), .A2(n7710), .ZN(n12721) );
  INV_X1 U15179 ( .A(n12713), .ZN(n12714) );
  NAND2_X1 U15180 ( .A1(n15166), .A2(n12716), .ZN(n12720) );
  OAI21_X1 U15181 ( .B1(n15379), .B2(n14816), .A(n14823), .ZN(n12717) );
  NAND2_X1 U15182 ( .A1(n12717), .A2(n7127), .ZN(n12719) );
  OR3_X1 U15183 ( .A1(n15379), .A2(n14823), .A3(n14816), .ZN(n12718) );
  NAND2_X1 U15184 ( .A1(n12721), .A2(n12747), .ZN(n12725) );
  AOI21_X2 U15185 ( .B1(n12725), .B2(n15807), .A(n12724), .ZN(n15369) );
  NAND2_X1 U15186 ( .A1(n15379), .A2(n14964), .ZN(n15151) );
  INV_X1 U15187 ( .A(n12726), .ZN(n12727) );
  AOI21_X1 U15188 ( .B1(n15168), .B2(n15384), .A(n12727), .ZN(n15150) );
  NAND2_X1 U15189 ( .A1(n12729), .A2(n15384), .ZN(n12731) );
  INV_X1 U15190 ( .A(n12729), .ZN(n12730) );
  AOI22_X1 U15191 ( .A1(n15187), .A2(n12731), .B1(n12730), .B2(n14812), .ZN(
        n12732) );
  INV_X1 U15192 ( .A(n15151), .ZN(n12733) );
  NAND2_X1 U15193 ( .A1(n15373), .A2(n14963), .ZN(n12737) );
  OAI211_X1 U15194 ( .C1(n15159), .C2(n14866), .A(n12759), .B(n15447), .ZN(
        n15368) );
  NOR2_X1 U15195 ( .A1(n15368), .A2(n15281), .ZN(n12741) );
  AOI22_X1 U15196 ( .A1(n12738), .A2(n15331), .B1(P1_REG2_REG_27__SCAN_IN), 
        .B2(n15286), .ZN(n12739) );
  OAI21_X1 U15197 ( .B1(n14866), .B2(n15339), .A(n12739), .ZN(n12740) );
  AOI211_X1 U15198 ( .C1(n15366), .C2(n15290), .A(n12741), .B(n12740), .ZN(
        n12742) );
  OAI21_X1 U15199 ( .B1(n15369), .B2(n15286), .A(n12742), .ZN(P1_U3266) );
  NAND2_X1 U15200 ( .A1(n14456), .A2(n8743), .ZN(n12744) );
  OR2_X1 U15201 ( .A1(n8724), .A2(n15535), .ZN(n12743) );
  NAND2_X1 U15202 ( .A1(n15361), .A2(n15352), .ZN(n15142) );
  OAI21_X1 U15203 ( .B1(n15119), .B2(n12748), .A(n15143), .ZN(n12758) );
  INV_X1 U15204 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n12751) );
  NAND2_X1 U15205 ( .A1(n14835), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n12750) );
  OR2_X1 U15206 ( .A1(n14834), .A2(n15136), .ZN(n12749) );
  OAI211_X1 U15207 ( .C1(n14839), .C2(n12751), .A(n12750), .B(n12749), .ZN(
        n12752) );
  INV_X1 U15208 ( .A(n12752), .ZN(n12753) );
  AOI21_X1 U15209 ( .B1(n12759), .B2(n15361), .A(n7130), .ZN(n12760) );
  NAND2_X1 U15210 ( .A1(n12760), .A2(n15131), .ZN(n15363) );
  AOI22_X1 U15211 ( .A1(n14535), .A2(n15331), .B1(P1_REG2_REG_28__SCAN_IN), 
        .B2(n15286), .ZN(n12762) );
  NAND2_X1 U15212 ( .A1(n15361), .A2(n15291), .ZN(n12761) );
  OAI211_X1 U15213 ( .C1(n15363), .C2(n15281), .A(n12762), .B(n12761), .ZN(
        n12763) );
  INV_X1 U15214 ( .A(n12763), .ZN(n12767) );
  OR2_X1 U15215 ( .A1(n14868), .A2(n14962), .ZN(n15117) );
  NAND2_X1 U15216 ( .A1(n12765), .A2(n15119), .ZN(n15359) );
  NAND3_X1 U15217 ( .A1(n15360), .A2(n15359), .A3(n15290), .ZN(n12766) );
  OAI211_X1 U15218 ( .C1(n15365), .C2(n15286), .A(n12767), .B(n12766), .ZN(
        P1_U3265) );
  INV_X1 U15219 ( .A(n12770), .ZN(P2_U3498) );
  INV_X1 U15220 ( .A(n12771), .ZN(n12773) );
  OAI222_X1 U15221 ( .A1(n14472), .A2(n12774), .B1(P2_U3088), .B2(n12773), 
        .C1(n14474), .C2(n12772), .ZN(P2_U3297) );
  INV_X1 U15222 ( .A(n13358), .ZN(n13175) );
  XNOR2_X1 U15223 ( .A(n13440), .B(n7285), .ZN(n12804) );
  XNOR2_X1 U15224 ( .A(n13381), .B(n7285), .ZN(n12788) );
  INV_X1 U15225 ( .A(n12788), .ZN(n12789) );
  XNOR2_X1 U15226 ( .A(n13384), .B(n7285), .ZN(n12786) );
  INV_X1 U15227 ( .A(n12786), .ZN(n12787) );
  XNOR2_X1 U15228 ( .A(n13469), .B(n7285), .ZN(n12784) );
  INV_X1 U15229 ( .A(n12784), .ZN(n12785) );
  XNOR2_X1 U15230 ( .A(n13491), .B(n7285), .ZN(n12780) );
  INV_X1 U15231 ( .A(n12780), .ZN(n12781) );
  INV_X1 U15232 ( .A(n12775), .ZN(n12776) );
  XNOR2_X1 U15233 ( .A(n12780), .B(n12858), .ZN(n12926) );
  XOR2_X1 U15234 ( .A(n7285), .B(n13481), .Z(n12854) );
  XNOR2_X1 U15235 ( .A(n13477), .B(n12792), .ZN(n12783) );
  NAND2_X1 U15236 ( .A1(n12783), .A2(n12782), .ZN(n12863) );
  NOR2_X1 U15237 ( .A1(n12783), .A2(n12782), .ZN(n12865) );
  XNOR2_X1 U15238 ( .A(n12784), .B(n12869), .ZN(n12905) );
  XNOR2_X1 U15239 ( .A(n12786), .B(n13266), .ZN(n12823) );
  XNOR2_X1 U15240 ( .A(n12788), .B(n13247), .ZN(n12889) );
  XNOR2_X1 U15241 ( .A(n13251), .B(n7285), .ZN(n12790) );
  XNOR2_X1 U15242 ( .A(n12790), .B(n13233), .ZN(n12839) );
  NAND2_X1 U15243 ( .A1(n12790), .A2(n13268), .ZN(n12812) );
  XNOR2_X1 U15244 ( .A(n13451), .B(n12792), .ZN(n12893) );
  NAND2_X1 U15245 ( .A1(n12893), .A2(n12942), .ZN(n12813) );
  XOR2_X1 U15246 ( .A(n7285), .B(n13212), .Z(n12877) );
  XNOR2_X1 U15247 ( .A(n13225), .B(n12792), .ZN(n12875) );
  AOI22_X1 U15248 ( .A1(n12877), .A2(n12941), .B1(n12875), .B2(n13234), .ZN(
        n12793) );
  INV_X1 U15249 ( .A(n12793), .ZN(n12800) );
  INV_X1 U15250 ( .A(n12893), .ZN(n12794) );
  NAND2_X1 U15251 ( .A1(n12794), .A2(n13246), .ZN(n12811) );
  INV_X1 U15252 ( .A(n12877), .ZN(n12798) );
  OAI21_X1 U15253 ( .B1(n12875), .B2(n13234), .A(n12941), .ZN(n12797) );
  NOR2_X1 U15254 ( .A1(n13234), .A2(n12941), .ZN(n12796) );
  INV_X1 U15255 ( .A(n12875), .ZN(n12795) );
  AOI22_X1 U15256 ( .A1(n12798), .A2(n12797), .B1(n12796), .B2(n12795), .ZN(
        n12799) );
  INV_X1 U15257 ( .A(n12801), .ZN(n12802) );
  XNOR2_X1 U15258 ( .A(n12804), .B(n13180), .ZN(n12847) );
  XNOR2_X1 U15259 ( .A(n12920), .B(n7285), .ZN(n12805) );
  XNOR2_X1 U15260 ( .A(n13358), .B(n7285), .ZN(n12829) );
  OAI22_X1 U15261 ( .A1(n12931), .A2(n12807), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n12806), .ZN(n12809) );
  NOR2_X1 U15262 ( .A1(n12917), .A2(n13196), .ZN(n12808) );
  AOI211_X1 U15263 ( .C1(n13173), .C2(n12934), .A(n12809), .B(n12808), .ZN(
        n12810) );
  NAND3_X1 U15264 ( .A1(n12838), .A2(n12812), .A3(n12811), .ZN(n12814) );
  NAND2_X1 U15265 ( .A1(n12814), .A2(n12813), .ZN(n12874) );
  XNOR2_X1 U15266 ( .A(n12874), .B(n12875), .ZN(n12876) );
  XNOR2_X1 U15267 ( .A(n12876), .B(n12897), .ZN(n12820) );
  INV_X1 U15268 ( .A(P3_REG3_REG_23__SCAN_IN), .ZN(n12815) );
  OAI22_X1 U15269 ( .A1(n12931), .A2(n13220), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n12815), .ZN(n12817) );
  NOR2_X1 U15270 ( .A1(n13246), .A2(n12917), .ZN(n12816) );
  AOI211_X1 U15271 ( .C1(n13226), .C2(n12934), .A(n12817), .B(n12816), .ZN(
        n12819) );
  NAND2_X1 U15272 ( .A1(n13225), .A2(n12919), .ZN(n12818) );
  OAI211_X1 U15273 ( .C1(n12820), .C2(n12922), .A(n12819), .B(n12818), .ZN(
        P3_U3156) );
  INV_X1 U15274 ( .A(n13384), .ZN(n13283) );
  AOI211_X1 U15275 ( .C1(n12823), .C2(n12822), .A(n12922), .B(n12821), .ZN(
        n12824) );
  INV_X1 U15276 ( .A(n12824), .ZN(n12828) );
  NAND2_X1 U15277 ( .A1(n13303), .A2(n12929), .ZN(n12825) );
  NAND2_X1 U15278 ( .A1(P3_U3151), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n13127)
         );
  OAI211_X1 U15279 ( .C1(n13247), .C2(n12931), .A(n12825), .B(n13127), .ZN(
        n12826) );
  AOI21_X1 U15280 ( .B1(n13281), .B2(n12934), .A(n12826), .ZN(n12827) );
  OAI211_X1 U15281 ( .C1(n13283), .C2(n12937), .A(n12828), .B(n12827), .ZN(
        P3_U3159) );
  INV_X1 U15282 ( .A(n12829), .ZN(n12830) );
  XNOR2_X1 U15283 ( .A(n13150), .B(n7285), .ZN(n12833) );
  AOI22_X1 U15284 ( .A1(n12929), .A2(n12940), .B1(P3_REG3_REG_28__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12834) );
  OAI21_X1 U15285 ( .B1(n13157), .B2(n12931), .A(n12834), .ZN(n12836) );
  NOR2_X1 U15286 ( .A1(n13428), .A2(n12937), .ZN(n12835) );
  AOI211_X1 U15287 ( .C1(n13163), .C2(n12934), .A(n12836), .B(n12835), .ZN(
        n12837) );
  INV_X1 U15288 ( .A(n13251), .ZN(n13456) );
  OAI21_X1 U15289 ( .B1(n12840), .B2(n12839), .A(n12838), .ZN(n12841) );
  NAND2_X1 U15290 ( .A1(n12841), .A2(n12924), .ZN(n12845) );
  AOI22_X1 U15291 ( .A1(n13276), .A2(n12929), .B1(P3_REG3_REG_21__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12842) );
  OAI21_X1 U15292 ( .B1(n13246), .B2(n12931), .A(n12842), .ZN(n12843) );
  AOI21_X1 U15293 ( .B1(n13250), .B2(n12934), .A(n12843), .ZN(n12844) );
  OAI211_X1 U15294 ( .C1(n13456), .C2(n12937), .A(n12845), .B(n12844), .ZN(
        P3_U3163) );
  XOR2_X1 U15295 ( .A(n12847), .B(n12846), .Z(n12853) );
  NAND2_X1 U15296 ( .A1(n12934), .A2(n13200), .ZN(n12849) );
  AOI22_X1 U15297 ( .A1(n12914), .A2(n13170), .B1(P3_REG3_REG_25__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12848) );
  OAI211_X1 U15298 ( .C1(n13220), .C2(n12917), .A(n12849), .B(n12848), .ZN(
        n12850) );
  AOI21_X1 U15299 ( .B1(n12851), .B2(n12919), .A(n12850), .ZN(n12852) );
  OAI21_X1 U15300 ( .B1(n12853), .B2(n12922), .A(n12852), .ZN(P3_U3165) );
  XNOR2_X1 U15301 ( .A(n12854), .B(n12932), .ZN(n12855) );
  XNOR2_X1 U15302 ( .A(n12856), .B(n12855), .ZN(n12862) );
  NAND2_X1 U15303 ( .A1(n12914), .A2(n13313), .ZN(n12857) );
  NAND2_X1 U15304 ( .A1(P3_U3151), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n13072)
         );
  OAI211_X1 U15305 ( .C1(n12917), .C2(n12858), .A(n12857), .B(n13072), .ZN(
        n12859) );
  AOI21_X1 U15306 ( .B1(n12934), .B2(n13309), .A(n12859), .ZN(n12861) );
  NAND2_X1 U15307 ( .A1(n13481), .A2(n12919), .ZN(n12860) );
  OAI211_X1 U15308 ( .C1(n12862), .C2(n12922), .A(n12861), .B(n12860), .ZN(
        P3_U3166) );
  INV_X1 U15309 ( .A(n12863), .ZN(n12864) );
  NOR2_X1 U15310 ( .A1(n12865), .A2(n12864), .ZN(n12866) );
  XNOR2_X1 U15311 ( .A(n12867), .B(n12866), .ZN(n12873) );
  NOR2_X1 U15312 ( .A1(n7111), .A2(P3_STATE_REG_SCAN_IN), .ZN(n13097) );
  AOI21_X1 U15313 ( .B1(n13328), .B2(n12929), .A(n13097), .ZN(n12868) );
  OAI21_X1 U15314 ( .B1(n12869), .B2(n12931), .A(n12868), .ZN(n12871) );
  NOR2_X1 U15315 ( .A1(n13477), .A2(n12937), .ZN(n12870) );
  AOI211_X1 U15316 ( .C1(n13298), .C2(n12934), .A(n12871), .B(n12870), .ZN(
        n12872) );
  OAI21_X1 U15317 ( .B1(n12873), .B2(n12922), .A(n12872), .ZN(P3_U3168) );
  OAI22_X1 U15318 ( .A1(n12876), .A2(n13234), .B1(n12875), .B2(n12874), .ZN(
        n12879) );
  XNOR2_X1 U15319 ( .A(n12877), .B(n12941), .ZN(n12878) );
  XNOR2_X1 U15320 ( .A(n12879), .B(n12878), .ZN(n12884) );
  OAI22_X1 U15321 ( .A1(n12931), .A2(n13180), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n7299), .ZN(n12881) );
  NOR2_X1 U15322 ( .A1(n12897), .A2(n12917), .ZN(n12880) );
  AOI211_X1 U15323 ( .C1(n13213), .C2(n12934), .A(n12881), .B(n12880), .ZN(
        n12883) );
  NAND2_X1 U15324 ( .A1(n13212), .A2(n12919), .ZN(n12882) );
  OAI211_X1 U15325 ( .C1(n12884), .C2(n12922), .A(n12883), .B(n12882), .ZN(
        P3_U3169) );
  AOI22_X1 U15326 ( .A1(n13290), .A2(n12929), .B1(P3_REG3_REG_20__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12886) );
  NAND2_X1 U15327 ( .A1(n12934), .A2(n13261), .ZN(n12885) );
  OAI211_X1 U15328 ( .C1(n13268), .C2(n12931), .A(n12886), .B(n12885), .ZN(
        n12891) );
  AOI211_X1 U15329 ( .C1(n12889), .C2(n12888), .A(n12922), .B(n12887), .ZN(
        n12890) );
  AOI211_X1 U15330 ( .C1(n12919), .C2(n13381), .A(n12891), .B(n12890), .ZN(
        n12892) );
  INV_X1 U15331 ( .A(n12892), .ZN(P3_U3173) );
  XNOR2_X1 U15332 ( .A(n12893), .B(n12942), .ZN(n12894) );
  XNOR2_X1 U15333 ( .A(n12895), .B(n12894), .ZN(n12902) );
  OAI22_X1 U15334 ( .A1(n13268), .A2(n12917), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n12896), .ZN(n12899) );
  NOR2_X1 U15335 ( .A1(n12897), .A2(n12931), .ZN(n12898) );
  AOI211_X1 U15336 ( .C1(n13237), .C2(n12934), .A(n12899), .B(n12898), .ZN(
        n12901) );
  NAND2_X1 U15337 ( .A1(n13451), .A2(n12919), .ZN(n12900) );
  OAI211_X1 U15338 ( .C1(n12902), .C2(n12922), .A(n12901), .B(n12900), .ZN(
        P3_U3175) );
  INV_X1 U15339 ( .A(n13469), .ZN(n12911) );
  AOI211_X1 U15340 ( .C1(n12905), .C2(n12904), .A(n12922), .B(n12903), .ZN(
        n12906) );
  INV_X1 U15341 ( .A(n12906), .ZN(n12910) );
  NAND2_X1 U15342 ( .A1(n13313), .A2(n12929), .ZN(n12907) );
  NAND2_X1 U15343 ( .A1(P3_U3151), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n13109)
         );
  OAI211_X1 U15344 ( .C1(n13266), .C2(n12931), .A(n12907), .B(n13109), .ZN(
        n12908) );
  AOI21_X1 U15345 ( .B1(n13293), .B2(n12934), .A(n12908), .ZN(n12909) );
  OAI211_X1 U15346 ( .C1(n12911), .C2(n12937), .A(n12910), .B(n12909), .ZN(
        P3_U3178) );
  XOR2_X1 U15347 ( .A(n12913), .B(n12912), .Z(n12923) );
  NAND2_X1 U15348 ( .A1(n12934), .A2(n13186), .ZN(n12916) );
  AOI22_X1 U15349 ( .A1(n12914), .A2(n12940), .B1(P3_REG3_REG_26__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12915) );
  OAI211_X1 U15350 ( .C1(n13180), .C2(n12917), .A(n12916), .B(n12915), .ZN(
        n12918) );
  AOI21_X1 U15351 ( .B1(n12920), .B2(n12919), .A(n12918), .ZN(n12921) );
  OAI21_X1 U15352 ( .B1(n12923), .B2(n12922), .A(n12921), .ZN(P3_U3180) );
  OAI211_X1 U15353 ( .C1(n12927), .C2(n12926), .A(n12925), .B(n12924), .ZN(
        n12936) );
  AND2_X1 U15354 ( .A1(P3_U3151), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n13051) );
  AOI21_X1 U15355 ( .B1(n12929), .B2(n13327), .A(n13051), .ZN(n12930) );
  OAI21_X1 U15356 ( .B1(n12932), .B2(n12931), .A(n12930), .ZN(n12933) );
  AOI21_X1 U15357 ( .B1(n12934), .B2(n13320), .A(n12933), .ZN(n12935) );
  OAI211_X1 U15358 ( .C1(n12937), .C2(n13491), .A(n12936), .B(n12935), .ZN(
        P3_U3181) );
  MUX2_X1 U15359 ( .A(P3_DATAO_REG_31__SCAN_IN), .B(n12938), .S(P3_U3897), .Z(
        P3_U3522) );
  MUX2_X1 U15360 ( .A(P3_DATAO_REG_29__SCAN_IN), .B(n12939), .S(P3_U3897), .Z(
        P3_U3520) );
  MUX2_X1 U15361 ( .A(P3_DATAO_REG_27__SCAN_IN), .B(n12940), .S(P3_U3897), .Z(
        P3_U3518) );
  MUX2_X1 U15362 ( .A(P3_DATAO_REG_26__SCAN_IN), .B(n13170), .S(P3_U3897), .Z(
        P3_U3517) );
  MUX2_X1 U15363 ( .A(P3_DATAO_REG_24__SCAN_IN), .B(n12941), .S(P3_U3897), .Z(
        P3_U3515) );
  MUX2_X1 U15364 ( .A(P3_DATAO_REG_23__SCAN_IN), .B(n13234), .S(P3_U3897), .Z(
        P3_U3514) );
  MUX2_X1 U15365 ( .A(P3_DATAO_REG_22__SCAN_IN), .B(n12942), .S(P3_U3897), .Z(
        P3_U3513) );
  MUX2_X1 U15366 ( .A(P3_DATAO_REG_21__SCAN_IN), .B(n13233), .S(P3_U3897), .Z(
        P3_U3512) );
  MUX2_X1 U15367 ( .A(P3_DATAO_REG_20__SCAN_IN), .B(n13276), .S(P3_U3897), .Z(
        P3_U3511) );
  MUX2_X1 U15368 ( .A(n13290), .B(P3_DATAO_REG_19__SCAN_IN), .S(n12943), .Z(
        P3_U3510) );
  MUX2_X1 U15369 ( .A(P3_DATAO_REG_18__SCAN_IN), .B(n13303), .S(P3_U3897), .Z(
        P3_U3509) );
  MUX2_X1 U15370 ( .A(n13313), .B(P3_DATAO_REG_17__SCAN_IN), .S(n12943), .Z(
        P3_U3508) );
  MUX2_X1 U15371 ( .A(P3_DATAO_REG_16__SCAN_IN), .B(n13328), .S(P3_U3897), .Z(
        P3_U3507) );
  MUX2_X1 U15372 ( .A(n13341), .B(P3_DATAO_REG_15__SCAN_IN), .S(n12943), .Z(
        P3_U3506) );
  MUX2_X1 U15373 ( .A(P3_DATAO_REG_14__SCAN_IN), .B(n13327), .S(P3_U3897), .Z(
        P3_U3505) );
  MUX2_X1 U15374 ( .A(P3_DATAO_REG_13__SCAN_IN), .B(n13338), .S(P3_U3897), .Z(
        P3_U3504) );
  MUX2_X1 U15375 ( .A(P3_DATAO_REG_12__SCAN_IN), .B(n12944), .S(P3_U3897), .Z(
        P3_U3503) );
  MUX2_X1 U15376 ( .A(P3_DATAO_REG_11__SCAN_IN), .B(n12945), .S(P3_U3897), .Z(
        P3_U3502) );
  MUX2_X1 U15377 ( .A(P3_DATAO_REG_10__SCAN_IN), .B(n12946), .S(P3_U3897), .Z(
        P3_U3501) );
  MUX2_X1 U15378 ( .A(P3_DATAO_REG_9__SCAN_IN), .B(n12947), .S(P3_U3897), .Z(
        P3_U3500) );
  MUX2_X1 U15379 ( .A(P3_DATAO_REG_8__SCAN_IN), .B(n12948), .S(P3_U3897), .Z(
        P3_U3499) );
  MUX2_X1 U15380 ( .A(P3_DATAO_REG_7__SCAN_IN), .B(n12949), .S(P3_U3897), .Z(
        P3_U3498) );
  MUX2_X1 U15381 ( .A(P3_DATAO_REG_6__SCAN_IN), .B(n12950), .S(P3_U3897), .Z(
        P3_U3497) );
  MUX2_X1 U15382 ( .A(P3_DATAO_REG_5__SCAN_IN), .B(n12951), .S(P3_U3897), .Z(
        P3_U3496) );
  MUX2_X1 U15383 ( .A(P3_DATAO_REG_3__SCAN_IN), .B(n12952), .S(P3_U3897), .Z(
        P3_U3494) );
  MUX2_X1 U15384 ( .A(P3_DATAO_REG_2__SCAN_IN), .B(n12953), .S(P3_U3897), .Z(
        P3_U3493) );
  MUX2_X1 U15385 ( .A(P3_DATAO_REG_1__SCAN_IN), .B(n12954), .S(P3_U3897), .Z(
        P3_U3492) );
  NAND2_X1 U15386 ( .A1(n15922), .A2(n12955), .ZN(n12968) );
  OAI21_X1 U15387 ( .B1(P3_REG2_REG_1__SCAN_IN), .B2(n12957), .A(n12956), .ZN(
        n12961) );
  OAI21_X1 U15388 ( .B1(P3_REG1_REG_1__SCAN_IN), .B2(n12959), .A(n12958), .ZN(
        n12960) );
  AOI22_X1 U15389 ( .A1(n15916), .A2(n12961), .B1(n15915), .B2(n12960), .ZN(
        n12967) );
  OAI21_X1 U15390 ( .B1(n12963), .B2(n15917), .A(n12962), .ZN(n12964) );
  AOI22_X1 U15391 ( .A1(n15914), .A2(n12964), .B1(P3_REG3_REG_1__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12966) );
  NAND2_X1 U15392 ( .A1(n15913), .A2(P3_ADDR_REG_1__SCAN_IN), .ZN(n12965) );
  NAND4_X1 U15393 ( .A1(n12968), .A2(n12967), .A3(n12966), .A4(n12965), .ZN(
        P3_U3183) );
  XNOR2_X1 U15394 ( .A(n13008), .B(n12969), .ZN(n13009) );
  NAND2_X1 U15395 ( .A1(n12970), .A2(P3_REG1_REG_11__SCAN_IN), .ZN(n12973) );
  NAND2_X1 U15396 ( .A1(n12971), .A2(n12975), .ZN(n12972) );
  XOR2_X1 U15397 ( .A(n13009), .B(n13010), .Z(n12991) );
  NOR2_X1 U15398 ( .A1(n12975), .A2(n12974), .ZN(n12977) );
  MUX2_X1 U15399 ( .A(P3_REG2_REG_12__SCAN_IN), .B(P3_REG1_REG_12__SCAN_IN), 
        .S(n7233), .Z(n12997) );
  XNOR2_X1 U15400 ( .A(n12997), .B(n13008), .ZN(n12976) );
  NOR2_X1 U15401 ( .A1(n13002), .A2(n13116), .ZN(n12989) );
  OAI21_X1 U15402 ( .B1(n12978), .B2(n12977), .A(n12976), .ZN(n12988) );
  INV_X1 U15403 ( .A(n12979), .ZN(n12980) );
  AOI21_X1 U15404 ( .B1(n15913), .B2(P3_ADDR_REG_12__SCAN_IN), .A(n12980), 
        .ZN(n12981) );
  OAI21_X1 U15405 ( .B1(n13129), .B2(n13008), .A(n12981), .ZN(n12987) );
  INV_X1 U15406 ( .A(P3_REG2_REG_12__SCAN_IN), .ZN(n12993) );
  XNOR2_X1 U15407 ( .A(n13008), .B(n12993), .ZN(n12982) );
  OR3_X1 U15408 ( .A1(n12984), .A2(n12983), .A3(n12982), .ZN(n12985) );
  AOI21_X1 U15409 ( .B1(n12992), .B2(n12985), .A(n13141), .ZN(n12986) );
  AOI211_X1 U15410 ( .C1(n12989), .C2(n12988), .A(n12987), .B(n12986), .ZN(
        n12990) );
  OAI21_X1 U15411 ( .B1(n12991), .B2(n13118), .A(n12990), .ZN(P3_U3194) );
  AOI21_X1 U15412 ( .B1(n12995), .B2(n12994), .A(n13021), .ZN(n13014) );
  INV_X1 U15413 ( .A(n13027), .ZN(n13007) );
  INV_X1 U15414 ( .A(P3_ADDR_REG_13__SCAN_IN), .ZN(n15577) );
  OAI21_X1 U15415 ( .B1(n15925), .B2(n15577), .A(n12996), .ZN(n13006) );
  INV_X1 U15416 ( .A(n12997), .ZN(n12999) );
  NOR2_X1 U15417 ( .A1(n12999), .A2(n12998), .ZN(n13001) );
  MUX2_X1 U15418 ( .A(P3_REG2_REG_13__SCAN_IN), .B(P3_REG1_REG_13__SCAN_IN), 
        .S(n7233), .Z(n13028) );
  XNOR2_X1 U15419 ( .A(n13028), .B(n13027), .ZN(n13000) );
  INV_X1 U15420 ( .A(n13030), .ZN(n13004) );
  OAI21_X1 U15421 ( .B1(n13002), .B2(n13001), .A(n13000), .ZN(n13003) );
  AOI21_X1 U15422 ( .B1(n13004), .B2(n13003), .A(n13116), .ZN(n13005) );
  AOI211_X1 U15423 ( .C1(n15922), .C2(n13007), .A(n13006), .B(n13005), .ZN(
        n13013) );
  XNOR2_X1 U15424 ( .A(n13017), .B(P3_REG1_REG_13__SCAN_IN), .ZN(n13011) );
  NAND2_X1 U15425 ( .A1(n13011), .A2(n15915), .ZN(n13012) );
  OAI211_X1 U15426 ( .C1(n13014), .C2(n13141), .A(n13013), .B(n13012), .ZN(
        P3_U3195) );
  XNOR2_X1 U15427 ( .A(n13042), .B(P3_REG1_REG_14__SCAN_IN), .ZN(n13039) );
  INV_X1 U15428 ( .A(n13015), .ZN(n13016) );
  XOR2_X1 U15429 ( .A(n13039), .B(n13040), .Z(n13038) );
  INV_X1 U15430 ( .A(n13018), .ZN(n13020) );
  INV_X1 U15431 ( .A(P3_REG2_REG_14__SCAN_IN), .ZN(n13019) );
  XNOR2_X1 U15432 ( .A(n13042), .B(n13019), .ZN(n13025) );
  INV_X1 U15433 ( .A(n13055), .ZN(n13023) );
  NOR3_X1 U15434 ( .A1(n13021), .A2(n13020), .A3(n13025), .ZN(n13022) );
  OAI21_X1 U15435 ( .B1(n13023), .B2(n13022), .A(n15916), .ZN(n13037) );
  INV_X1 U15436 ( .A(n13042), .ZN(n13035) );
  INV_X1 U15437 ( .A(P3_ADDR_REG_14__SCAN_IN), .ZN(n15622) );
  OAI21_X1 U15438 ( .B1(n15925), .B2(n15622), .A(n13024), .ZN(n13034) );
  INV_X1 U15439 ( .A(n13025), .ZN(n13026) );
  MUX2_X1 U15440 ( .A(n13039), .B(n13026), .S(n13122), .Z(n13032) );
  NOR2_X1 U15441 ( .A1(n13028), .A2(n13027), .ZN(n13029) );
  OR2_X1 U15442 ( .A1(n13030), .A2(n13029), .ZN(n13031) );
  AOI211_X1 U15443 ( .C1(n13032), .C2(n13031), .A(n13116), .B(n13047), .ZN(
        n13033) );
  AOI211_X1 U15444 ( .C1(n15922), .C2(n13035), .A(n13034), .B(n13033), .ZN(
        n13036) );
  OAI211_X1 U15445 ( .C1(n13038), .C2(n13118), .A(n13037), .B(n13036), .ZN(
        P3_U3196) );
  NAND2_X1 U15446 ( .A1(n13042), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n13043) );
  OAI21_X1 U15447 ( .B1(n13041), .B2(P3_REG1_REG_15__SCAN_IN), .A(n13064), 
        .ZN(n13060) );
  NAND2_X1 U15448 ( .A1(n13042), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n13054) );
  INV_X1 U15449 ( .A(n13054), .ZN(n13045) );
  INV_X1 U15450 ( .A(n13043), .ZN(n13044) );
  MUX2_X1 U15451 ( .A(n13045), .B(n13044), .S(n7233), .Z(n13046) );
  MUX2_X1 U15452 ( .A(P3_REG2_REG_15__SCAN_IN), .B(P3_REG1_REG_15__SCAN_IN), 
        .S(n7233), .Z(n13049) );
  OAI211_X1 U15453 ( .C1(n13050), .C2(n13049), .A(n13066), .B(n15914), .ZN(
        n13053) );
  AOI21_X1 U15454 ( .B1(n15913), .B2(P3_ADDR_REG_15__SCAN_IN), .A(n13051), 
        .ZN(n13052) );
  OAI211_X1 U15455 ( .C1(n13129), .C2(n13063), .A(n13053), .B(n13052), .ZN(
        n13059) );
  NAND2_X1 U15456 ( .A1(n13056), .A2(n13330), .ZN(n13057) );
  AOI21_X1 U15457 ( .B1(n13077), .B2(n13057), .A(n13141), .ZN(n13058) );
  AOI211_X1 U15458 ( .C1(n15915), .C2(n13060), .A(n13059), .B(n13058), .ZN(
        n13061) );
  INV_X1 U15459 ( .A(n13061), .ZN(P3_U3197) );
  XNOR2_X1 U15460 ( .A(n13088), .B(P3_REG1_REG_16__SCAN_IN), .ZN(n13085) );
  NAND2_X1 U15461 ( .A1(n13063), .A2(n13062), .ZN(n13065) );
  NAND2_X1 U15462 ( .A1(n13065), .A2(n13064), .ZN(n13086) );
  XOR2_X1 U15463 ( .A(n13085), .B(n13086), .Z(n13083) );
  INV_X1 U15464 ( .A(P3_REG2_REG_16__SCAN_IN), .ZN(n13315) );
  MUX2_X1 U15465 ( .A(n13315), .B(n13394), .S(n6527), .Z(n13068) );
  NOR2_X1 U15466 ( .A1(n13088), .A2(n13068), .ZN(n13093) );
  INV_X1 U15467 ( .A(n13093), .ZN(n13069) );
  NAND2_X1 U15468 ( .A1(n13088), .A2(n13068), .ZN(n13092) );
  NAND2_X1 U15469 ( .A1(n13069), .A2(n13092), .ZN(n13070) );
  XNOR2_X1 U15470 ( .A(n13094), .B(n13070), .ZN(n13081) );
  NAND2_X1 U15471 ( .A1(n15913), .A2(P3_ADDR_REG_16__SCAN_IN), .ZN(n13071) );
  OAI211_X1 U15472 ( .C1(n13129), .C2(n13084), .A(n13072), .B(n13071), .ZN(
        n13080) );
  XNOR2_X1 U15473 ( .A(n13088), .B(P3_REG2_REG_16__SCAN_IN), .ZN(n13074) );
  NAND2_X1 U15474 ( .A1(n13073), .A2(n13074), .ZN(n13087) );
  INV_X1 U15475 ( .A(n13074), .ZN(n13076) );
  NAND3_X1 U15476 ( .A1(n13077), .A2(n13076), .A3(n13075), .ZN(n13078) );
  AOI21_X1 U15477 ( .B1(n13087), .B2(n13078), .A(n13141), .ZN(n13079) );
  AOI211_X1 U15478 ( .C1(n15914), .C2(n13081), .A(n13080), .B(n13079), .ZN(
        n13082) );
  OAI21_X1 U15479 ( .B1(n13118), .B2(n13083), .A(n13082), .ZN(P3_U3198) );
  XOR2_X1 U15480 ( .A(P3_REG1_REG_17__SCAN_IN), .B(n13104), .Z(n13101) );
  OAI21_X1 U15481 ( .B1(n13088), .B2(n13315), .A(n13087), .ZN(n13089) );
  OAI21_X1 U15482 ( .B1(n13089), .B2(n13112), .A(n13107), .ZN(n13090) );
  INV_X1 U15483 ( .A(n13090), .ZN(n13091) );
  INV_X1 U15484 ( .A(P3_REG2_REG_17__SCAN_IN), .ZN(n13305) );
  MUX2_X1 U15485 ( .A(P3_REG2_REG_17__SCAN_IN), .B(P3_REG1_REG_17__SCAN_IN), 
        .S(n7233), .Z(n13113) );
  XNOR2_X1 U15486 ( .A(n13113), .B(n13112), .ZN(n13096) );
  AOI21_X1 U15487 ( .B1(n15913), .B2(P3_ADDR_REG_17__SCAN_IN), .A(n13097), 
        .ZN(n13098) );
  OAI21_X1 U15488 ( .B1(n13129), .B2(n13112), .A(n13098), .ZN(n13099) );
  XOR2_X1 U15489 ( .A(P3_REG1_REG_18__SCAN_IN), .B(n13132), .Z(n13133) );
  INV_X1 U15490 ( .A(n13102), .ZN(n13103) );
  INV_X1 U15491 ( .A(P3_REG2_REG_18__SCAN_IN), .ZN(n13292) );
  OR2_X1 U15492 ( .A1(n13132), .A2(n13292), .ZN(n13119) );
  NAND2_X1 U15493 ( .A1(n13132), .A2(n13292), .ZN(n13105) );
  NAND2_X1 U15494 ( .A1(n13119), .A2(n13105), .ZN(n13106) );
  INV_X1 U15495 ( .A(P3_ADDR_REG_18__SCAN_IN), .ZN(n13110) );
  OAI21_X1 U15496 ( .B1(n15925), .B2(n13110), .A(n13109), .ZN(n13117) );
  MUX2_X1 U15497 ( .A(P3_REG2_REG_18__SCAN_IN), .B(P3_REG1_REG_18__SCAN_IN), 
        .S(n7233), .Z(n13115) );
  XNOR2_X1 U15498 ( .A(n13128), .B(P3_REG2_REG_19__SCAN_IN), .ZN(n13123) );
  XNOR2_X1 U15499 ( .A(n13128), .B(P3_REG1_REG_19__SCAN_IN), .ZN(n13135) );
  MUX2_X1 U15500 ( .A(n13135), .B(n13123), .S(n13122), .Z(n13124) );
  XNOR2_X1 U15501 ( .A(n13125), .B(n13124), .ZN(n13131) );
  NAND2_X1 U15502 ( .A1(n15913), .A2(P3_ADDR_REG_19__SCAN_IN), .ZN(n13126) );
  OAI211_X1 U15503 ( .C1(n13129), .C2(n13128), .A(n13127), .B(n13126), .ZN(
        n13130) );
  AOI21_X1 U15504 ( .B1(n13131), .B2(n15914), .A(n13130), .ZN(n13140) );
  INV_X1 U15505 ( .A(n13135), .ZN(n13136) );
  XNOR2_X1 U15506 ( .A(n13137), .B(n13136), .ZN(n13138) );
  NAND2_X1 U15507 ( .A1(n13138), .A2(n15915), .ZN(n13139) );
  OAI211_X1 U15508 ( .C1(n13142), .C2(n13141), .A(n13140), .B(n13139), .ZN(
        P3_U3201) );
  NOR2_X1 U15509 ( .A1(n13144), .A2(n13143), .ZN(n13417) );
  AOI21_X1 U15510 ( .B1(n13350), .B2(n13417), .A(n13145), .ZN(n13149) );
  NAND2_X1 U15511 ( .A1(n13346), .A2(P3_REG2_REG_31__SCAN_IN), .ZN(n13146) );
  OAI211_X1 U15512 ( .C1(n13419), .C2(n13348), .A(n13149), .B(n13146), .ZN(
        P3_U3202) );
  NAND2_X1 U15513 ( .A1(n13346), .A2(P3_REG2_REG_30__SCAN_IN), .ZN(n13148) );
  OAI211_X1 U15514 ( .C1(n13422), .C2(n13348), .A(n13149), .B(n13148), .ZN(
        P3_U3203) );
  NAND2_X1 U15515 ( .A1(n13166), .A2(n13152), .ZN(n13154) );
  NAND2_X1 U15516 ( .A1(n13154), .A2(n13153), .ZN(n13156) );
  NAND3_X1 U15517 ( .A1(n13156), .A2(n13336), .A3(n13155), .ZN(n13160) );
  OAI22_X1 U15518 ( .A1(n13181), .A2(n13265), .B1(n13157), .B2(n13267), .ZN(
        n13158) );
  INV_X1 U15519 ( .A(n13158), .ZN(n13159) );
  NAND2_X1 U15520 ( .A1(n13160), .A2(n13159), .ZN(n13430) );
  INV_X1 U15521 ( .A(n13163), .ZN(n13164) );
  OAI22_X1 U15522 ( .A1(n13428), .A2(n13348), .B1(n13164), .B2(n13321), .ZN(
        n13165) );
  OAI21_X1 U15523 ( .B1(n13168), .B2(n13167), .A(n13166), .ZN(n13171) );
  AOI22_X1 U15524 ( .A1(n13346), .A2(P3_REG2_REG_27__SCAN_IN), .B1(n13345), 
        .B2(n13173), .ZN(n13174) );
  OAI21_X1 U15525 ( .B1(n13175), .B2(n13348), .A(n13174), .ZN(n13176) );
  AOI21_X1 U15526 ( .B1(n13359), .B2(n13324), .A(n13176), .ZN(n13177) );
  OAI21_X1 U15527 ( .B1(n13360), .B2(n13346), .A(n13177), .ZN(P3_U3206) );
  XNOR2_X1 U15528 ( .A(n13178), .B(n13185), .ZN(n13179) );
  INV_X1 U15529 ( .A(n13361), .ZN(n13190) );
  INV_X1 U15530 ( .A(n13182), .ZN(n13183) );
  AOI21_X1 U15531 ( .B1(n13185), .B2(n13184), .A(n13183), .ZN(n13362) );
  AOI22_X1 U15532 ( .A1(n13346), .A2(P3_REG2_REG_26__SCAN_IN), .B1(n13345), 
        .B2(n13186), .ZN(n13187) );
  OAI21_X1 U15533 ( .B1(n13436), .B2(n13348), .A(n13187), .ZN(n13188) );
  AOI21_X1 U15534 ( .B1(n13362), .B2(n13324), .A(n13188), .ZN(n13189) );
  OAI21_X1 U15535 ( .B1(n13346), .B2(n13190), .A(n13189), .ZN(P3_U3207) );
  OAI211_X1 U15536 ( .C1(n13193), .C2(n13192), .A(n13191), .B(n13336), .ZN(
        n13195) );
  OR2_X1 U15537 ( .A1(n13220), .A2(n13265), .ZN(n13194) );
  OAI211_X1 U15538 ( .C1(n13196), .C2(n13267), .A(n13195), .B(n13194), .ZN(
        n13364) );
  INV_X1 U15539 ( .A(n13364), .ZN(n13204) );
  OAI21_X1 U15540 ( .B1(n13199), .B2(n13198), .A(n13197), .ZN(n13365) );
  AOI22_X1 U15541 ( .A1(n13346), .A2(P3_REG2_REG_25__SCAN_IN), .B1(n13345), 
        .B2(n13200), .ZN(n13201) );
  OAI21_X1 U15542 ( .B1(n13440), .B2(n13348), .A(n13201), .ZN(n13202) );
  AOI21_X1 U15543 ( .B1(n13365), .B2(n13324), .A(n13202), .ZN(n13203) );
  OAI21_X1 U15544 ( .B1(n13346), .B2(n13204), .A(n13203), .ZN(P3_U3208) );
  NOR2_X1 U15545 ( .A1(n6577), .A2(n13219), .ZN(n13218) );
  NOR2_X1 U15546 ( .A1(n13218), .A2(n13205), .ZN(n13206) );
  XNOR2_X1 U15547 ( .A(n13206), .B(n8608), .ZN(n13209) );
  AOI22_X1 U15548 ( .A1(n13234), .A2(n13339), .B1(n13340), .B2(n13207), .ZN(
        n13208) );
  OAI21_X1 U15549 ( .B1(n13209), .B2(n13245), .A(n13208), .ZN(n13368) );
  INV_X1 U15550 ( .A(n13368), .ZN(n13217) );
  OAI21_X1 U15551 ( .B1(n13211), .B2(n8608), .A(n13210), .ZN(n13369) );
  INV_X1 U15552 ( .A(n13212), .ZN(n13444) );
  AOI22_X1 U15553 ( .A1(n13346), .A2(P3_REG2_REG_24__SCAN_IN), .B1(n13345), 
        .B2(n13213), .ZN(n13214) );
  OAI21_X1 U15554 ( .B1(n13444), .B2(n13348), .A(n13214), .ZN(n13215) );
  AOI21_X1 U15555 ( .B1(n13369), .B2(n13324), .A(n13215), .ZN(n13216) );
  OAI21_X1 U15556 ( .B1(n13217), .B2(n13346), .A(n13216), .ZN(P3_U3209) );
  AOI211_X1 U15557 ( .C1(n13219), .C2(n6577), .A(n13245), .B(n13218), .ZN(
        n13222) );
  OAI22_X1 U15558 ( .A1(n13246), .A2(n13265), .B1(n13220), .B2(n13267), .ZN(
        n13221) );
  OR2_X1 U15559 ( .A1(n13222), .A2(n13221), .ZN(n13372) );
  INV_X1 U15560 ( .A(n13372), .ZN(n13230) );
  XNOR2_X1 U15561 ( .A(n13224), .B(n13223), .ZN(n13373) );
  INV_X1 U15562 ( .A(n13225), .ZN(n13448) );
  AOI22_X1 U15563 ( .A1(n13226), .A2(n13345), .B1(n13346), .B2(
        P3_REG2_REG_23__SCAN_IN), .ZN(n13227) );
  OAI21_X1 U15564 ( .B1(n13448), .B2(n13348), .A(n13227), .ZN(n13228) );
  AOI21_X1 U15565 ( .B1(n13373), .B2(n13324), .A(n13228), .ZN(n13229) );
  OAI21_X1 U15566 ( .B1(n13230), .B2(n13346), .A(n13229), .ZN(P3_U3210) );
  XNOR2_X1 U15567 ( .A(n13231), .B(n13232), .ZN(n13454) );
  INV_X1 U15568 ( .A(P3_REG2_REG_22__SCAN_IN), .ZN(n13236) );
  XNOR2_X1 U15569 ( .A(n6667), .B(n13232), .ZN(n13235) );
  AOI222_X1 U15570 ( .A1(n13336), .A2(n13235), .B1(n13234), .B2(n13340), .C1(
        n13233), .C2(n13339), .ZN(n13449) );
  MUX2_X1 U15571 ( .A(n13236), .B(n13449), .S(n13350), .Z(n13239) );
  AOI22_X1 U15572 ( .A1(n13451), .A2(n13310), .B1(n13345), .B2(n13237), .ZN(
        n13238) );
  OAI211_X1 U15573 ( .C1(n13454), .C2(n13352), .A(n13239), .B(n13238), .ZN(
        P3_U3211) );
  XNOR2_X1 U15574 ( .A(n13241), .B(n13240), .ZN(n13457) );
  XNOR2_X1 U15575 ( .A(n13243), .B(n13242), .ZN(n13244) );
  OAI222_X1 U15576 ( .A1(n13265), .A2(n13247), .B1(n13267), .B2(n13246), .C1(
        n13245), .C2(n13244), .ZN(n13455) );
  INV_X1 U15577 ( .A(n13455), .ZN(n13248) );
  MUX2_X1 U15578 ( .A(n13249), .B(n13248), .S(n13350), .Z(n13253) );
  AOI22_X1 U15579 ( .A1(n13251), .A2(n13310), .B1(n13345), .B2(n13250), .ZN(
        n13252) );
  OAI211_X1 U15580 ( .C1(n13457), .C2(n13352), .A(n13253), .B(n13252), .ZN(
        P3_U3212) );
  INV_X1 U15581 ( .A(n13255), .ZN(n13256) );
  AOI21_X1 U15582 ( .B1(n13296), .B2(n13257), .A(n13256), .ZN(n13280) );
  NAND2_X1 U15583 ( .A1(n13280), .A2(n13279), .ZN(n13278) );
  AND2_X1 U15584 ( .A1(n13278), .A2(n13258), .ZN(n13260) );
  OAI21_X1 U15585 ( .B1(n13260), .B2(n6861), .A(n13259), .ZN(n13461) );
  AOI22_X1 U15586 ( .A1(n13381), .A2(n13310), .B1(n13345), .B2(n13261), .ZN(
        n13274) );
  NAND2_X1 U15587 ( .A1(n13262), .A2(n6861), .ZN(n13263) );
  NAND3_X1 U15588 ( .A1(n13264), .A2(n13336), .A3(n13263), .ZN(n13271) );
  OAI22_X1 U15589 ( .A1(n13268), .A2(n13267), .B1(n13266), .B2(n13265), .ZN(
        n13269) );
  INV_X1 U15590 ( .A(n13269), .ZN(n13270) );
  NAND2_X1 U15591 ( .A1(n13271), .A2(n13270), .ZN(n13462) );
  MUX2_X1 U15592 ( .A(n13462), .B(P3_REG2_REG_20__SCAN_IN), .S(n13346), .Z(
        n13272) );
  INV_X1 U15593 ( .A(n13272), .ZN(n13273) );
  OAI211_X1 U15594 ( .C1(n13461), .C2(n13352), .A(n13274), .B(n13273), .ZN(
        P3_U3213) );
  XOR2_X1 U15595 ( .A(n13275), .B(n13279), .Z(n13277) );
  AOI222_X1 U15596 ( .A1(n13336), .A2(n13277), .B1(n13276), .B2(n13340), .C1(
        n13303), .C2(n13339), .ZN(n13386) );
  OAI21_X1 U15597 ( .B1(n13280), .B2(n13279), .A(n13278), .ZN(n13385) );
  AOI22_X1 U15598 ( .A1(n13345), .A2(n13281), .B1(n13346), .B2(
        P3_REG2_REG_19__SCAN_IN), .ZN(n13282) );
  OAI21_X1 U15599 ( .B1(n13283), .B2(n13348), .A(n13282), .ZN(n13284) );
  AOI21_X1 U15600 ( .B1(n13385), .B2(n13324), .A(n13284), .ZN(n13285) );
  OAI21_X1 U15601 ( .B1(n13346), .B2(n13386), .A(n13285), .ZN(P3_U3214) );
  NAND2_X1 U15602 ( .A1(n13296), .A2(n13286), .ZN(n13287) );
  XNOR2_X1 U15603 ( .A(n13287), .B(n13289), .ZN(n13471) );
  OAI21_X1 U15604 ( .B1(n8035), .B2(n13289), .A(n13288), .ZN(n13291) );
  AOI222_X1 U15605 ( .A1(n13336), .A2(n13291), .B1(n13313), .B2(n13339), .C1(
        n13290), .C2(n13340), .ZN(n13466) );
  MUX2_X1 U15606 ( .A(n13292), .B(n13466), .S(n13350), .Z(n13295) );
  AOI22_X1 U15607 ( .A1(n13469), .A2(n13310), .B1(n13345), .B2(n13293), .ZN(
        n13294) );
  OAI211_X1 U15608 ( .C1(n13471), .C2(n13352), .A(n13295), .B(n13294), .ZN(
        P3_U3215) );
  OAI21_X1 U15609 ( .B1(n13297), .B2(n13301), .A(n13296), .ZN(n13472) );
  INV_X1 U15610 ( .A(n13298), .ZN(n13299) );
  OAI22_X1 U15611 ( .A1(n13477), .A2(n13348), .B1(n13299), .B2(n13321), .ZN(
        n13300) );
  AOI21_X1 U15612 ( .B1(n13472), .B2(n13324), .A(n13300), .ZN(n13307) );
  XNOR2_X1 U15613 ( .A(n13302), .B(n13301), .ZN(n13304) );
  AOI222_X1 U15614 ( .A1(n13336), .A2(n13304), .B1(n13303), .B2(n13340), .C1(
        n13328), .C2(n13339), .ZN(n13473) );
  MUX2_X1 U15615 ( .A(n13305), .B(n13473), .S(n13350), .Z(n13306) );
  NAND2_X1 U15616 ( .A1(n13307), .A2(n13306), .ZN(P3_U3216) );
  XNOR2_X1 U15617 ( .A(n13308), .B(n13311), .ZN(n13484) );
  AOI22_X1 U15618 ( .A1(n13481), .A2(n13310), .B1(n13345), .B2(n13309), .ZN(
        n13317) );
  XNOR2_X1 U15619 ( .A(n13312), .B(n13311), .ZN(n13314) );
  AOI222_X1 U15620 ( .A1(n13336), .A2(n13314), .B1(n13313), .B2(n13340), .C1(
        n13341), .C2(n13339), .ZN(n13478) );
  MUX2_X1 U15621 ( .A(n13315), .B(n13478), .S(n13350), .Z(n13316) );
  OAI211_X1 U15622 ( .C1(n13484), .C2(n13352), .A(n13317), .B(n13316), .ZN(
        P3_U3217) );
  OAI21_X1 U15623 ( .B1(n13319), .B2(n13325), .A(n13318), .ZN(n13486) );
  INV_X1 U15624 ( .A(n13320), .ZN(n13322) );
  OAI22_X1 U15625 ( .A1(n13491), .A2(n13348), .B1(n13322), .B2(n13321), .ZN(
        n13323) );
  AOI21_X1 U15626 ( .B1(n13486), .B2(n13324), .A(n13323), .ZN(n13332) );
  XNOR2_X1 U15627 ( .A(n13326), .B(n13325), .ZN(n13329) );
  AOI222_X1 U15628 ( .A1(n13336), .A2(n13329), .B1(n13328), .B2(n13340), .C1(
        n13327), .C2(n13339), .ZN(n13487) );
  MUX2_X1 U15629 ( .A(n13330), .B(n13487), .S(n13350), .Z(n13331) );
  NAND2_X1 U15630 ( .A1(n13332), .A2(n13331), .ZN(P3_U3218) );
  XOR2_X1 U15631 ( .A(n13334), .B(n13333), .Z(n13499) );
  XNOR2_X1 U15632 ( .A(n13335), .B(n6979), .ZN(n13337) );
  NAND2_X1 U15633 ( .A1(n13337), .A2(n13336), .ZN(n13343) );
  AOI22_X1 U15634 ( .A1(n13341), .A2(n13340), .B1(n13339), .B2(n13338), .ZN(
        n13342) );
  NAND2_X1 U15635 ( .A1(n13343), .A2(n13342), .ZN(n13496) );
  AOI22_X1 U15636 ( .A1(n13346), .A2(P3_REG2_REG_14__SCAN_IN), .B1(n13345), 
        .B2(n13344), .ZN(n13347) );
  OAI21_X1 U15637 ( .B1(n13494), .B2(n13348), .A(n13347), .ZN(n13349) );
  AOI21_X1 U15638 ( .B1(n13496), .B2(n13350), .A(n13349), .ZN(n13351) );
  OAI21_X1 U15639 ( .B1(n13499), .B2(n13352), .A(n13351), .ZN(P3_U3219) );
  NAND2_X1 U15640 ( .A1(n15973), .A2(n13417), .ZN(n13354) );
  NAND2_X1 U15641 ( .A1(n15970), .A2(P3_REG1_REG_31__SCAN_IN), .ZN(n13353) );
  OAI211_X1 U15642 ( .C1(n13419), .C2(n13403), .A(n13354), .B(n13353), .ZN(
        P3_U3490) );
  NAND2_X1 U15643 ( .A1(n15970), .A2(P3_REG1_REG_30__SCAN_IN), .ZN(n13355) );
  OAI211_X1 U15644 ( .C1(n13422), .C2(n13403), .A(n13355), .B(n13354), .ZN(
        P3_U3489) );
  OAI22_X1 U15645 ( .A1(n13429), .A2(n13406), .B1(n13428), .B2(n13403), .ZN(
        n13357) );
  MUX2_X1 U15646 ( .A(P3_REG1_REG_28__SCAN_IN), .B(n13430), .S(n15973), .Z(
        n13356) );
  MUX2_X1 U15647 ( .A(P3_REG1_REG_27__SCAN_IN), .B(n13433), .S(n15973), .Z(
        P3_U3486) );
  INV_X1 U15648 ( .A(P3_REG1_REG_26__SCAN_IN), .ZN(n13363) );
  INV_X1 U15649 ( .A(P3_REG1_REG_25__SCAN_IN), .ZN(n13366) );
  AOI21_X1 U15650 ( .B1(n13365), .B2(n13407), .A(n13364), .ZN(n13437) );
  MUX2_X1 U15651 ( .A(n13366), .B(n13437), .S(n15973), .Z(n13367) );
  OAI21_X1 U15652 ( .B1(n13440), .B2(n13403), .A(n13367), .ZN(P3_U3484) );
  INV_X1 U15653 ( .A(P3_REG1_REG_24__SCAN_IN), .ZN(n13370) );
  AOI21_X1 U15654 ( .B1(n13407), .B2(n13369), .A(n13368), .ZN(n13441) );
  MUX2_X1 U15655 ( .A(n13370), .B(n13441), .S(n15973), .Z(n13371) );
  OAI21_X1 U15656 ( .B1(n13444), .B2(n13403), .A(n13371), .ZN(P3_U3483) );
  INV_X1 U15657 ( .A(P3_REG1_REG_23__SCAN_IN), .ZN(n13374) );
  AOI21_X1 U15658 ( .B1(n13407), .B2(n13373), .A(n13372), .ZN(n13445) );
  MUX2_X1 U15659 ( .A(n13374), .B(n13445), .S(n15973), .Z(n13375) );
  OAI21_X1 U15660 ( .B1(n13448), .B2(n13403), .A(n13375), .ZN(P3_U3482) );
  INV_X1 U15661 ( .A(P3_REG1_REG_22__SCAN_IN), .ZN(n13376) );
  MUX2_X1 U15662 ( .A(n13376), .B(n13449), .S(n15973), .Z(n13378) );
  NAND2_X1 U15663 ( .A1(n13451), .A2(n13395), .ZN(n13377) );
  OAI211_X1 U15664 ( .C1(n13406), .C2(n13454), .A(n13378), .B(n13377), .ZN(
        P3_U3481) );
  MUX2_X1 U15665 ( .A(n13455), .B(P3_REG1_REG_21__SCAN_IN), .S(n15970), .Z(
        n13380) );
  OAI22_X1 U15666 ( .A1(n13457), .A2(n13406), .B1(n13456), .B2(n13403), .ZN(
        n13379) );
  OR2_X1 U15667 ( .A1(n13380), .A2(n13379), .ZN(P3_U3480) );
  INV_X1 U15668 ( .A(n13381), .ZN(n13460) );
  OAI22_X1 U15669 ( .A1(n13461), .A2(n13406), .B1(n13460), .B2(n13403), .ZN(
        n13383) );
  MUX2_X1 U15670 ( .A(n13462), .B(P3_REG1_REG_20__SCAN_IN), .S(n15970), .Z(
        n13382) );
  OR2_X1 U15671 ( .A1(n13383), .A2(n13382), .ZN(P3_U3479) );
  AOI22_X1 U15672 ( .A1(n13385), .A2(n13407), .B1(n15960), .B2(n13384), .ZN(
        n13387) );
  NAND2_X1 U15673 ( .A1(n13387), .A2(n13386), .ZN(n13465) );
  MUX2_X1 U15674 ( .A(P3_REG1_REG_19__SCAN_IN), .B(n13465), .S(n15973), .Z(
        P3_U3478) );
  MUX2_X1 U15675 ( .A(n13388), .B(n13466), .S(n15973), .Z(n13390) );
  NAND2_X1 U15676 ( .A1(n13469), .A2(n13395), .ZN(n13389) );
  OAI211_X1 U15677 ( .C1(n13471), .C2(n13406), .A(n13390), .B(n13389), .ZN(
        P3_U3477) );
  NAND2_X1 U15678 ( .A1(n13472), .A2(n13398), .ZN(n13393) );
  INV_X1 U15679 ( .A(P3_REG1_REG_17__SCAN_IN), .ZN(n13391) );
  MUX2_X1 U15680 ( .A(n13391), .B(n13473), .S(n15973), .Z(n13392) );
  OAI211_X1 U15681 ( .C1(n13403), .C2(n13477), .A(n13393), .B(n13392), .ZN(
        P3_U3476) );
  MUX2_X1 U15682 ( .A(n13394), .B(n13478), .S(n15973), .Z(n13397) );
  NAND2_X1 U15683 ( .A1(n13481), .A2(n13395), .ZN(n13396) );
  OAI211_X1 U15684 ( .C1(n13484), .C2(n13406), .A(n13397), .B(n13396), .ZN(
        P3_U3475) );
  NAND2_X1 U15685 ( .A1(n13486), .A2(n13398), .ZN(n13401) );
  INV_X1 U15686 ( .A(P3_REG1_REG_15__SCAN_IN), .ZN(n13399) );
  MUX2_X1 U15687 ( .A(n13399), .B(n13487), .S(n15973), .Z(n13400) );
  OAI211_X1 U15688 ( .C1(n13403), .C2(n13491), .A(n13401), .B(n13400), .ZN(
        P3_U3474) );
  OAI22_X1 U15689 ( .A1(n13494), .A2(n13403), .B1(n15973), .B2(n13402), .ZN(
        n13404) );
  AOI21_X1 U15690 ( .B1(n13496), .B2(n15973), .A(n13404), .ZN(n13405) );
  OAI21_X1 U15691 ( .B1(n13499), .B2(n13406), .A(n13405), .ZN(P3_U3473) );
  NAND2_X1 U15692 ( .A1(n13408), .A2(n13407), .ZN(n13410) );
  OAI211_X1 U15693 ( .C1(n15946), .C2(n13411), .A(n13410), .B(n13409), .ZN(
        n13500) );
  MUX2_X1 U15694 ( .A(P3_REG1_REG_11__SCAN_IN), .B(n13500), .S(n15973), .Z(
        P3_U3470) );
  AOI21_X1 U15695 ( .B1(n13413), .B2(n15960), .A(n13412), .ZN(n13414) );
  OAI21_X1 U15696 ( .B1(n13416), .B2(n13415), .A(n13414), .ZN(n13501) );
  MUX2_X1 U15697 ( .A(P3_REG1_REG_7__SCAN_IN), .B(n13501), .S(n15973), .Z(
        P3_U3466) );
  NAND2_X1 U15698 ( .A1(n15963), .A2(n13417), .ZN(n13420) );
  NAND2_X1 U15699 ( .A1(n15961), .A2(P3_REG0_REG_31__SCAN_IN), .ZN(n13418) );
  OAI211_X1 U15700 ( .C1(n13419), .C2(n13493), .A(n13420), .B(n13418), .ZN(
        P3_U3458) );
  NAND2_X1 U15701 ( .A1(n15961), .A2(P3_REG0_REG_30__SCAN_IN), .ZN(n13421) );
  OAI211_X1 U15702 ( .C1(n13422), .C2(n13493), .A(n13421), .B(n13420), .ZN(
        P3_U3457) );
  NAND2_X1 U15703 ( .A1(n13423), .A2(n13480), .ZN(n13426) );
  INV_X1 U15704 ( .A(P3_REG0_REG_29__SCAN_IN), .ZN(n13424) );
  OAI211_X1 U15705 ( .C1(n13427), .C2(n13498), .A(n13426), .B(n13425), .ZN(
        P3_U3456) );
  OAI22_X1 U15706 ( .A1(n13429), .A2(n13498), .B1(n13428), .B2(n13493), .ZN(
        n13432) );
  MUX2_X1 U15707 ( .A(n13430), .B(P3_REG0_REG_28__SCAN_IN), .S(n15961), .Z(
        n13431) );
  MUX2_X1 U15708 ( .A(P3_REG0_REG_27__SCAN_IN), .B(n13433), .S(n15963), .Z(
        P3_U3454) );
  INV_X1 U15709 ( .A(P3_REG0_REG_25__SCAN_IN), .ZN(n13438) );
  MUX2_X1 U15710 ( .A(n13438), .B(n13437), .S(n15963), .Z(n13439) );
  OAI21_X1 U15711 ( .B1(n13440), .B2(n13493), .A(n13439), .ZN(P3_U3452) );
  INV_X1 U15712 ( .A(P3_REG0_REG_24__SCAN_IN), .ZN(n13442) );
  MUX2_X1 U15713 ( .A(n13442), .B(n13441), .S(n15963), .Z(n13443) );
  OAI21_X1 U15714 ( .B1(n13444), .B2(n13493), .A(n13443), .ZN(P3_U3451) );
  MUX2_X1 U15715 ( .A(n13446), .B(n13445), .S(n15963), .Z(n13447) );
  OAI21_X1 U15716 ( .B1(n13448), .B2(n13493), .A(n13447), .ZN(P3_U3450) );
  MUX2_X1 U15717 ( .A(n13450), .B(n13449), .S(n15963), .Z(n13453) );
  NAND2_X1 U15718 ( .A1(n13451), .A2(n13480), .ZN(n13452) );
  OAI211_X1 U15719 ( .C1(n13454), .C2(n13498), .A(n13453), .B(n13452), .ZN(
        P3_U3449) );
  MUX2_X1 U15720 ( .A(n13455), .B(P3_REG0_REG_21__SCAN_IN), .S(n15961), .Z(
        n13459) );
  OAI22_X1 U15721 ( .A1(n13457), .A2(n13498), .B1(n13456), .B2(n13493), .ZN(
        n13458) );
  OR2_X1 U15722 ( .A1(n13459), .A2(n13458), .ZN(P3_U3448) );
  OAI22_X1 U15723 ( .A1(n13461), .A2(n13498), .B1(n13460), .B2(n13493), .ZN(
        n13464) );
  MUX2_X1 U15724 ( .A(n13462), .B(P3_REG0_REG_20__SCAN_IN), .S(n15961), .Z(
        n13463) );
  OR2_X1 U15725 ( .A1(n13464), .A2(n13463), .ZN(P3_U3447) );
  MUX2_X1 U15726 ( .A(P3_REG0_REG_19__SCAN_IN), .B(n13465), .S(n15963), .Z(
        P3_U3446) );
  INV_X1 U15727 ( .A(n13466), .ZN(n13467) );
  MUX2_X1 U15728 ( .A(P3_REG0_REG_18__SCAN_IN), .B(n13467), .S(n15963), .Z(
        n13468) );
  AOI21_X1 U15729 ( .B1(n13480), .B2(n13469), .A(n13468), .ZN(n13470) );
  OAI21_X1 U15730 ( .B1(n13498), .B2(n13471), .A(n13470), .ZN(P3_U3444) );
  NAND2_X1 U15731 ( .A1(n13472), .A2(n13485), .ZN(n13476) );
  MUX2_X1 U15732 ( .A(n13474), .B(n13473), .S(n15963), .Z(n13475) );
  OAI211_X1 U15733 ( .C1(n13493), .C2(n13477), .A(n13476), .B(n13475), .ZN(
        P3_U3441) );
  INV_X1 U15734 ( .A(P3_REG0_REG_16__SCAN_IN), .ZN(n13479) );
  MUX2_X1 U15735 ( .A(n13479), .B(n13478), .S(n15963), .Z(n13483) );
  NAND2_X1 U15736 ( .A1(n13481), .A2(n13480), .ZN(n13482) );
  OAI211_X1 U15737 ( .C1(n13484), .C2(n13498), .A(n13483), .B(n13482), .ZN(
        P3_U3438) );
  NAND2_X1 U15738 ( .A1(n13486), .A2(n13485), .ZN(n13490) );
  INV_X1 U15739 ( .A(P3_REG0_REG_15__SCAN_IN), .ZN(n13488) );
  MUX2_X1 U15740 ( .A(n13488), .B(n13487), .S(n15963), .Z(n13489) );
  OAI211_X1 U15741 ( .C1(n13493), .C2(n13491), .A(n13490), .B(n13489), .ZN(
        P3_U3435) );
  OAI22_X1 U15742 ( .A1(n13494), .A2(n13493), .B1(n13492), .B2(n15963), .ZN(
        n13495) );
  AOI21_X1 U15743 ( .B1(n13496), .B2(n15963), .A(n13495), .ZN(n13497) );
  OAI21_X1 U15744 ( .B1(n13499), .B2(n13498), .A(n13497), .ZN(P3_U3432) );
  MUX2_X1 U15745 ( .A(P3_REG0_REG_11__SCAN_IN), .B(n13500), .S(n15963), .Z(
        P3_U3423) );
  MUX2_X1 U15746 ( .A(n13501), .B(P3_REG0_REG_7__SCAN_IN), .S(n15961), .Z(
        P3_U3411) );
  INV_X1 U15747 ( .A(n13502), .ZN(n13508) );
  NOR4_X1 U15748 ( .A1(n13503), .A2(P3_IR_REG_30__SCAN_IN), .A3(P3_U3151), 
        .A4(n13504), .ZN(n13505) );
  AOI21_X1 U15749 ( .B1(n13506), .B2(SI_31_), .A(n13505), .ZN(n13507) );
  OAI21_X1 U15750 ( .B1(n13508), .B2(n13524), .A(n13507), .ZN(P3_U3264) );
  INV_X1 U15751 ( .A(n13509), .ZN(n13511) );
  OAI222_X1 U15752 ( .A1(n13528), .A2(n13512), .B1(n13524), .B2(n13511), .C1(
        P3_U3151), .C2(n13510), .ZN(P3_U3266) );
  OAI222_X1 U15753 ( .A1(P3_U3151), .A2(n13515), .B1(n13528), .B2(n13514), 
        .C1(n13524), .C2(n13513), .ZN(P3_U3267) );
  INV_X1 U15754 ( .A(n13516), .ZN(n13518) );
  OAI222_X1 U15755 ( .A1(n13111), .A2(P3_U3151), .B1(n13524), .B2(n13518), 
        .C1(n13517), .C2(n13528), .ZN(P3_U3268) );
  INV_X1 U15756 ( .A(n13519), .ZN(n13525) );
  INV_X1 U15757 ( .A(n13520), .ZN(n13523) );
  OAI222_X1 U15758 ( .A1(P3_U3151), .A2(n13525), .B1(n13524), .B2(n13523), 
        .C1(n13522), .C2(n13521), .ZN(P3_U3269) );
  OAI222_X1 U15759 ( .A1(n13529), .A2(P3_U3151), .B1(n13528), .B2(n13527), 
        .C1(n13524), .C2(n13526), .ZN(P3_U3270) );
  MUX2_X1 U15760 ( .A(n13530), .B(P3_IR_REG_0__SCAN_IN), .S(
        P3_STATE_REG_SCAN_IN), .Z(P3_U3295) );
  INV_X1 U15761 ( .A(n14405), .ZN(n13572) );
  XNOR2_X1 U15762 ( .A(n14039), .B(n11422), .ZN(n13652) );
  NAND2_X1 U15763 ( .A1(n13788), .A2(n15891), .ZN(n13588) );
  XNOR2_X1 U15764 ( .A(n7324), .B(n13615), .ZN(n13544) );
  AND2_X1 U15765 ( .A1(n13787), .A2(n14307), .ZN(n13545) );
  NOR2_X1 U15766 ( .A1(n13544), .A2(n13545), .ZN(n13654) );
  INV_X1 U15767 ( .A(n13531), .ZN(n13697) );
  NAND2_X1 U15768 ( .A1(n13697), .A2(n13532), .ZN(n13533) );
  NAND2_X1 U15769 ( .A1(n13699), .A2(n13533), .ZN(n13534) );
  XNOR2_X1 U15770 ( .A(n14325), .B(n13615), .ZN(n13535) );
  NAND2_X1 U15771 ( .A1(n13791), .A2(n15891), .ZN(n13536) );
  XNOR2_X1 U15772 ( .A(n13535), .B(n13536), .ZN(n13696) );
  INV_X1 U15773 ( .A(n13535), .ZN(n13537) );
  NAND2_X1 U15774 ( .A1(n13537), .A2(n13536), .ZN(n13538) );
  XNOR2_X1 U15775 ( .A(n14320), .B(n11422), .ZN(n13539) );
  NAND2_X1 U15776 ( .A1(n13790), .A2(n15891), .ZN(n13540) );
  XNOR2_X1 U15777 ( .A(n13539), .B(n13540), .ZN(n13632) );
  XNOR2_X1 U15778 ( .A(n14417), .B(n11422), .ZN(n13715) );
  NAND2_X1 U15779 ( .A1(n13789), .A2(n15891), .ZN(n13717) );
  INV_X1 U15780 ( .A(n13539), .ZN(n13542) );
  INV_X1 U15781 ( .A(n13540), .ZN(n13541) );
  NAND2_X1 U15782 ( .A1(n13542), .A2(n13541), .ZN(n13713) );
  OAI21_X1 U15783 ( .B1(n13715), .B2(n13717), .A(n13713), .ZN(n13543) );
  INV_X1 U15784 ( .A(n13544), .ZN(n13650) );
  INV_X1 U15785 ( .A(n13545), .ZN(n13546) );
  NOR2_X1 U15786 ( .A1(n13650), .A2(n13546), .ZN(n13653) );
  INV_X1 U15787 ( .A(n13654), .ZN(n13548) );
  NOR2_X1 U15788 ( .A1(n13652), .A2(n13588), .ZN(n13547) );
  NAND2_X1 U15789 ( .A1(n13548), .A2(n13547), .ZN(n13549) );
  XNOR2_X1 U15790 ( .A(n7352), .B(n13615), .ZN(n13551) );
  AND2_X1 U15791 ( .A1(n13786), .A2(n14307), .ZN(n13552) );
  NAND2_X1 U15792 ( .A1(n13551), .A2(n13552), .ZN(n13556) );
  INV_X1 U15793 ( .A(n13551), .ZN(n13753) );
  INV_X1 U15794 ( .A(n13552), .ZN(n13553) );
  NAND2_X1 U15795 ( .A1(n13753), .A2(n13553), .ZN(n13554) );
  NAND2_X1 U15796 ( .A1(n13556), .A2(n13554), .ZN(n13655) );
  INV_X1 U15797 ( .A(n13655), .ZN(n13555) );
  XNOR2_X1 U15798 ( .A(n13995), .B(n13615), .ZN(n13557) );
  NAND2_X1 U15799 ( .A1(n13785), .A2(n15891), .ZN(n13558) );
  XNOR2_X1 U15800 ( .A(n13557), .B(n13558), .ZN(n13763) );
  INV_X1 U15801 ( .A(n13557), .ZN(n13559) );
  XNOR2_X1 U15802 ( .A(n14405), .B(n13615), .ZN(n13561) );
  INV_X1 U15803 ( .A(n13561), .ZN(n13563) );
  AND2_X1 U15804 ( .A1(n13784), .A2(n14307), .ZN(n13560) );
  INV_X1 U15805 ( .A(n13560), .ZN(n13562) );
  AOI21_X1 U15806 ( .B1(n13563), .B2(n13562), .A(n13619), .ZN(n13564) );
  OR2_X1 U15807 ( .A1(n13614), .A2(n13743), .ZN(n13567) );
  NAND2_X1 U15808 ( .A1(n13785), .A2(n13769), .ZN(n13566) );
  NAND2_X1 U15809 ( .A1(n13567), .A2(n13566), .ZN(n13977) );
  OAI22_X1 U15810 ( .A1(n13983), .A2(n13775), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13568), .ZN(n13569) );
  AOI21_X1 U15811 ( .B1(n13977), .B2(n13773), .A(n13569), .ZN(n13570) );
  OAI211_X1 U15812 ( .C1(n13572), .C2(n13749), .A(n13571), .B(n13570), .ZN(
        P2_U3186) );
  NAND2_X1 U15813 ( .A1(n13798), .A2(n13769), .ZN(n13573) );
  OAI21_X1 U15814 ( .B1(n13670), .B2(n13743), .A(n13573), .ZN(n14171) );
  NAND2_X1 U15815 ( .A1(n13773), .A2(n14171), .ZN(n13575) );
  OAI211_X1 U15816 ( .C1(n13775), .C2(n14173), .A(n13575), .B(n13574), .ZN(
        n13583) );
  INV_X1 U15817 ( .A(n13703), .ZN(n13579) );
  NOR3_X1 U15818 ( .A1(n13577), .A2(n13576), .A3(n13751), .ZN(n13578) );
  AOI21_X1 U15819 ( .B1(n13579), .B2(n13766), .A(n13578), .ZN(n13581) );
  NOR2_X1 U15820 ( .A1(n13581), .A2(n13580), .ZN(n13582) );
  AOI211_X1 U15821 ( .C1(n14435), .C2(n13777), .A(n13583), .B(n13582), .ZN(
        n13584) );
  OAI21_X1 U15822 ( .B1(n13585), .B2(n13736), .A(n13584), .ZN(P2_U3187) );
  INV_X1 U15823 ( .A(n13652), .ZN(n13587) );
  AOI22_X1 U15824 ( .A1(n13590), .A2(n13766), .B1(n13765), .B2(n13788), .ZN(
        n13597) );
  INV_X1 U15825 ( .A(n13588), .ZN(n13589) );
  NAND2_X1 U15826 ( .A1(n13590), .A2(n13589), .ZN(n13651) );
  INV_X1 U15827 ( .A(n13651), .ZN(n13596) );
  NAND2_X1 U15828 ( .A1(n13787), .A2(n13770), .ZN(n13592) );
  NAND2_X1 U15829 ( .A1(n13789), .A2(n13769), .ZN(n13591) );
  AND2_X1 U15830 ( .A1(n13592), .A2(n13591), .ZN(n14304) );
  AOI22_X1 U15831 ( .A1(n13756), .A2(n14033), .B1(P2_REG3_REG_23__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13593) );
  OAI21_X1 U15832 ( .B1(n14304), .B2(n13759), .A(n13593), .ZN(n13594) );
  AOI21_X1 U15833 ( .B1(n14039), .B2(n13777), .A(n13594), .ZN(n13595) );
  OAI21_X1 U15834 ( .B1(n13597), .B2(n13596), .A(n13595), .ZN(P2_U3188) );
  XNOR2_X1 U15835 ( .A(n13599), .B(n13598), .ZN(n13605) );
  INV_X1 U15836 ( .A(n14229), .ZN(n13602) );
  AOI22_X1 U15837 ( .A1(n13802), .A2(n13769), .B1(n13770), .B2(n13800), .ZN(
        n14227) );
  NOR2_X1 U15838 ( .A1(n13759), .A2(n14227), .ZN(n13600) );
  AOI211_X1 U15839 ( .C1(n13756), .C2(n13602), .A(n13601), .B(n13600), .ZN(
        n13604) );
  NAND2_X1 U15840 ( .A1(n14379), .A2(n13777), .ZN(n13603) );
  OAI211_X1 U15841 ( .C1(n13605), .C2(n13736), .A(n13604), .B(n13603), .ZN(
        P2_U3189) );
  OAI211_X1 U15842 ( .C1(n13608), .C2(n13607), .A(n13606), .B(n13766), .ZN(
        n13613) );
  INV_X1 U15843 ( .A(n13609), .ZN(n13610) );
  AOI22_X1 U15844 ( .A1(n13777), .A2(n15890), .B1(n13773), .B2(n13610), .ZN(
        n13612) );
  MUX2_X1 U15845 ( .A(n13775), .B(P2_STATE_REG_SCAN_IN), .S(
        P2_REG3_REG_3__SCAN_IN), .Z(n13611) );
  NAND3_X1 U15846 ( .A1(n13613), .A2(n13612), .A3(n13611), .ZN(P2_U3190) );
  OR2_X1 U15847 ( .A1(n13614), .A2(n14261), .ZN(n13616) );
  XNOR2_X1 U15848 ( .A(n13616), .B(n13615), .ZN(n13617) );
  XNOR2_X1 U15849 ( .A(n13972), .B(n13617), .ZN(n13620) );
  INV_X1 U15850 ( .A(n13620), .ZN(n13618) );
  NAND2_X1 U15851 ( .A1(n13618), .A2(n13766), .ZN(n13628) );
  INV_X1 U15852 ( .A(n13619), .ZN(n13623) );
  NAND4_X1 U15853 ( .A1(n13629), .A2(n13766), .A3(n13623), .A4(n13620), .ZN(
        n13627) );
  AOI22_X1 U15854 ( .A1(n13968), .A2(n13756), .B1(P2_REG3_REG_28__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13621) );
  OAI21_X1 U15855 ( .B1(n13622), .B2(n13759), .A(n13621), .ZN(n13625) );
  NOR2_X1 U15856 ( .A1(n13623), .A2(n13628), .ZN(n13624) );
  AOI211_X1 U15857 ( .C1(n13972), .C2(n13777), .A(n13625), .B(n13624), .ZN(
        n13626) );
  OAI211_X1 U15858 ( .C1(n13629), .C2(n13628), .A(n13627), .B(n13626), .ZN(
        P2_U3192) );
  AOI211_X1 U15859 ( .C1(n13632), .C2(n13631), .A(n13736), .B(n13630), .ZN(
        n13633) );
  INV_X1 U15860 ( .A(n13633), .ZN(n13637) );
  AOI22_X1 U15861 ( .A1(n13789), .A2(n13770), .B1(n13769), .B2(n13791), .ZN(
        n14068) );
  OAI22_X1 U15862 ( .A1(n14068), .A2(n13759), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13634), .ZN(n13635) );
  AOI21_X1 U15863 ( .B1(n14072), .B2(n13756), .A(n13635), .ZN(n13636) );
  OAI211_X1 U15864 ( .C1(n10202), .C2(n13749), .A(n13637), .B(n13636), .ZN(
        P2_U3195) );
  NAND2_X1 U15865 ( .A1(n13639), .A2(n13638), .ZN(n13641) );
  XOR2_X1 U15866 ( .A(n13641), .B(n13640), .Z(n13648) );
  NOR2_X1 U15867 ( .A1(n13775), .A2(n14194), .ZN(n13646) );
  NAND2_X1 U15868 ( .A1(n13800), .A2(n13769), .ZN(n13643) );
  NAND2_X1 U15869 ( .A1(n13798), .A2(n13770), .ZN(n13642) );
  AND2_X1 U15870 ( .A1(n13643), .A2(n13642), .ZN(n14192) );
  OAI21_X1 U15871 ( .B1(n13759), .B2(n14192), .A(n13644), .ZN(n13645) );
  AOI211_X1 U15872 ( .C1(n14197), .C2(n13777), .A(n13646), .B(n13645), .ZN(
        n13647) );
  OAI21_X1 U15873 ( .B1(n13648), .B2(n13736), .A(n13647), .ZN(P2_U3196) );
  INV_X1 U15874 ( .A(n7352), .ZN(n14008) );
  NOR3_X1 U15875 ( .A1(n13650), .A2(n13649), .A3(n13751), .ZN(n13657) );
  NOR2_X1 U15876 ( .A1(n13654), .A2(n13653), .ZN(n13686) );
  AOI21_X1 U15877 ( .B1(n13685), .B2(n13655), .A(n13736), .ZN(n13656) );
  AND2_X1 U15878 ( .A1(n13787), .A2(n13769), .ZN(n13658) );
  AOI21_X1 U15879 ( .B1(n13785), .B2(n13770), .A(n13658), .ZN(n14014) );
  INV_X1 U15880 ( .A(n14014), .ZN(n13661) );
  OAI22_X1 U15881 ( .A1(n14010), .A2(n13775), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13659), .ZN(n13660) );
  AOI21_X1 U15882 ( .B1(n13661), .B2(n13773), .A(n13660), .ZN(n13662) );
  XNOR2_X1 U15883 ( .A(n13675), .B(n13663), .ZN(n13669) );
  INV_X1 U15884 ( .A(n13664), .ZN(n13667) );
  XNOR2_X1 U15885 ( .A(n13666), .B(n13664), .ZN(n13767) );
  NAND2_X1 U15886 ( .A1(n13767), .A2(n13665), .ZN(n13768) );
  OAI21_X1 U15887 ( .B1(n13667), .B2(n13666), .A(n13768), .ZN(n13668) );
  NOR2_X1 U15888 ( .A1(n13668), .A2(n13669), .ZN(n13678) );
  AOI21_X1 U15889 ( .B1(n13669), .B2(n13668), .A(n13678), .ZN(n13674) );
  OAI22_X1 U15890 ( .A1(n13742), .A2(n13743), .B1(n13670), .B2(n13741), .ZN(
        n14139) );
  NAND2_X1 U15891 ( .A1(n13773), .A2(n14139), .ZN(n13671) );
  NAND2_X1 U15892 ( .A1(P2_U3088), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n13899)
         );
  OAI211_X1 U15893 ( .C1(n13775), .C2(n14149), .A(n13671), .B(n13899), .ZN(
        n13672) );
  AOI21_X1 U15894 ( .B1(n14148), .B2(n13777), .A(n13672), .ZN(n13673) );
  OAI21_X1 U15895 ( .B1(n13674), .B2(n13736), .A(n13673), .ZN(P2_U3198) );
  AOI22_X1 U15896 ( .A1(n13675), .A2(n13766), .B1(n13765), .B2(n13795), .ZN(
        n13677) );
  OR3_X1 U15897 ( .A1(n13678), .A2(n13677), .A3(n13676), .ZN(n13683) );
  AOI22_X1 U15898 ( .A1(n13793), .A2(n13770), .B1(n13769), .B2(n13795), .ZN(
        n14126) );
  INV_X1 U15899 ( .A(n14126), .ZN(n13679) );
  AOI22_X1 U15900 ( .A1(n13679), .A2(n13773), .B1(P2_REG3_REG_17__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13680) );
  OAI21_X1 U15901 ( .B1(n14132), .B2(n13775), .A(n13680), .ZN(n13681) );
  AOI21_X1 U15902 ( .B1(n14341), .B2(n13777), .A(n13681), .ZN(n13682) );
  OAI211_X1 U15903 ( .C1(n13736), .C2(n13684), .A(n13683), .B(n13682), .ZN(
        P2_U3200) );
  OAI211_X1 U15904 ( .C1(n13687), .C2(n13686), .A(n13685), .B(n13766), .ZN(
        n13692) );
  AOI22_X1 U15905 ( .A1(n13786), .A2(n13770), .B1(n13769), .B2(n13788), .ZN(
        n14022) );
  INV_X1 U15906 ( .A(n13688), .ZN(n14026) );
  AOI22_X1 U15907 ( .A1(n14026), .A2(n13756), .B1(P2_REG3_REG_24__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13689) );
  OAI21_X1 U15908 ( .B1(n14022), .B2(n13759), .A(n13689), .ZN(n13690) );
  AOI21_X1 U15909 ( .B1(n7324), .B2(n13777), .A(n13690), .ZN(n13691) );
  NAND2_X1 U15910 ( .A1(n13692), .A2(n13691), .ZN(P2_U3201) );
  AOI22_X1 U15911 ( .A1(n13790), .A2(n13770), .B1(n13769), .B2(n13792), .ZN(
        n14082) );
  OAI22_X1 U15912 ( .A1(n14082), .A2(n13759), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13693), .ZN(n13695) );
  NOR2_X1 U15913 ( .A1(n7668), .A2(n13749), .ZN(n13694) );
  AOI211_X1 U15914 ( .C1(n13756), .C2(n14086), .A(n13695), .B(n13694), .ZN(
        n13701) );
  OAI22_X1 U15915 ( .A1(n13697), .A2(n13736), .B1(n13744), .B2(n13751), .ZN(
        n13698) );
  NAND3_X1 U15916 ( .A1(n13699), .A2(n6945), .A3(n13698), .ZN(n13700) );
  OAI211_X1 U15917 ( .C1(n13702), .C2(n13736), .A(n13701), .B(n13700), .ZN(
        P2_U3205) );
  INV_X1 U15918 ( .A(n14362), .ZN(n13712) );
  OAI211_X1 U15919 ( .C1(n13705), .C2(n13704), .A(n13703), .B(n13766), .ZN(
        n13711) );
  INV_X1 U15920 ( .A(n13706), .ZN(n13709) );
  OAI22_X1 U15921 ( .A1(n13759), .A2(n13707), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n15843), .ZN(n13708) );
  AOI21_X1 U15922 ( .B1(n13709), .B2(n13756), .A(n13708), .ZN(n13710) );
  OAI211_X1 U15923 ( .C1(n13712), .C2(n13749), .A(n13711), .B(n13710), .ZN(
        P2_U3206) );
  INV_X1 U15924 ( .A(n13713), .ZN(n13714) );
  OR2_X1 U15925 ( .A1(n13630), .A2(n13714), .ZN(n13716) );
  XNOR2_X1 U15926 ( .A(n13716), .B(n13715), .ZN(n13718) );
  NAND3_X1 U15927 ( .A1(n13718), .A2(n13766), .A3(n13717), .ZN(n13727) );
  INV_X1 U15928 ( .A(n13718), .ZN(n13719) );
  NAND3_X1 U15929 ( .A1(n13719), .A2(n13765), .A3(n13789), .ZN(n13726) );
  NAND2_X1 U15930 ( .A1(n13788), .A2(n13770), .ZN(n13721) );
  NAND2_X1 U15931 ( .A1(n13790), .A2(n13769), .ZN(n13720) );
  NAND2_X1 U15932 ( .A1(n13721), .A2(n13720), .ZN(n14058) );
  OAI22_X1 U15933 ( .A1(n13775), .A2(n14052), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13722), .ZN(n13723) );
  AOI21_X1 U15934 ( .B1(n14058), .B2(n13773), .A(n13723), .ZN(n13725) );
  NAND2_X1 U15935 ( .A1(n14417), .A2(n13777), .ZN(n13724) );
  NAND4_X1 U15936 ( .A1(n13727), .A2(n13726), .A3(n13725), .A4(n13724), .ZN(
        P2_U3207) );
  XNOR2_X1 U15937 ( .A(n13729), .B(n13728), .ZN(n13735) );
  NAND2_X1 U15938 ( .A1(n13799), .A2(n13770), .ZN(n13730) );
  OAI21_X1 U15939 ( .B1(n13731), .B2(n13741), .A(n13730), .ZN(n14205) );
  AOI22_X1 U15940 ( .A1(n13773), .A2(n14205), .B1(P2_U3088), .B2(
        P2_REG3_REG_11__SCAN_IN), .ZN(n13732) );
  OAI21_X1 U15941 ( .B1(n14212), .B2(n13775), .A(n13732), .ZN(n13733) );
  AOI21_X1 U15942 ( .B1(n14443), .B2(n13777), .A(n13733), .ZN(n13734) );
  OAI21_X1 U15943 ( .B1(n13735), .B2(n13736), .A(n13734), .ZN(P2_U3208) );
  INV_X1 U15944 ( .A(n14335), .ZN(n14118) );
  AOI21_X1 U15945 ( .B1(n13738), .B2(n13737), .A(n13736), .ZN(n13740) );
  NAND2_X1 U15946 ( .A1(n13740), .A2(n13739), .ZN(n13748) );
  OAI22_X1 U15947 ( .A1(n13744), .A2(n13743), .B1(n13742), .B2(n13741), .ZN(
        n14107) );
  INV_X1 U15948 ( .A(n14107), .ZN(n13745) );
  NAND2_X1 U15949 ( .A1(P2_U3088), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n15858)
         );
  OAI21_X1 U15950 ( .B1(n13745), .B2(n13759), .A(n15858), .ZN(n13746) );
  AOI21_X1 U15951 ( .B1(n14115), .B2(n13756), .A(n13746), .ZN(n13747) );
  OAI211_X1 U15952 ( .C1(n14118), .C2(n13749), .A(n13748), .B(n13747), .ZN(
        P2_U3210) );
  INV_X1 U15953 ( .A(n13750), .ZN(n13755) );
  NOR3_X1 U15954 ( .A1(n13753), .A2(n13752), .A3(n13751), .ZN(n13754) );
  AOI21_X1 U15955 ( .B1(n13755), .B2(n13766), .A(n13754), .ZN(n13764) );
  AOI22_X1 U15956 ( .A1(n13784), .A2(n13770), .B1(n13769), .B2(n13786), .ZN(
        n13990) );
  NAND2_X1 U15957 ( .A1(n13995), .A2(n13777), .ZN(n13758) );
  AOI22_X1 U15958 ( .A1(n13998), .A2(n13756), .B1(P2_REG3_REG_26__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13757) );
  OAI211_X1 U15959 ( .C1(n13990), .C2(n13759), .A(n13758), .B(n13757), .ZN(
        n13760) );
  AOI21_X1 U15960 ( .B1(n13761), .B2(n13766), .A(n13760), .ZN(n13762) );
  OAI21_X1 U15961 ( .B1(n13764), .B2(n13763), .A(n13762), .ZN(P2_U3212) );
  AOI22_X1 U15962 ( .A1(n13767), .A2(n13766), .B1(n13765), .B2(n13796), .ZN(
        n13780) );
  INV_X1 U15963 ( .A(n13768), .ZN(n13779) );
  NAND2_X1 U15964 ( .A1(n13797), .A2(n13769), .ZN(n13772) );
  NAND2_X1 U15965 ( .A1(n13795), .A2(n13770), .ZN(n13771) );
  NAND2_X1 U15966 ( .A1(n13772), .A2(n13771), .ZN(n14161) );
  AOI22_X1 U15967 ( .A1(n13773), .A2(n14161), .B1(P2_REG3_REG_15__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13774) );
  OAI21_X1 U15968 ( .B1(n14166), .B2(n13775), .A(n13774), .ZN(n13776) );
  AOI21_X1 U15969 ( .B1(n14351), .B2(n13777), .A(n13776), .ZN(n13778) );
  OAI21_X1 U15970 ( .B1(n13780), .B2(n13779), .A(n13778), .ZN(P2_U3213) );
  MUX2_X1 U15971 ( .A(n13781), .B(P2_DATAO_REG_31__SCAN_IN), .S(n13811), .Z(
        P2_U3562) );
  MUX2_X1 U15972 ( .A(n13782), .B(P2_DATAO_REG_29__SCAN_IN), .S(n13811), .Z(
        P2_U3560) );
  MUX2_X1 U15973 ( .A(n13783), .B(P2_DATAO_REG_28__SCAN_IN), .S(n13811), .Z(
        P2_U3559) );
  MUX2_X1 U15974 ( .A(n13784), .B(P2_DATAO_REG_27__SCAN_IN), .S(n13811), .Z(
        P2_U3558) );
  MUX2_X1 U15975 ( .A(n13785), .B(P2_DATAO_REG_26__SCAN_IN), .S(n13811), .Z(
        P2_U3557) );
  MUX2_X1 U15976 ( .A(n13786), .B(P2_DATAO_REG_25__SCAN_IN), .S(n13811), .Z(
        P2_U3556) );
  MUX2_X1 U15977 ( .A(n13787), .B(P2_DATAO_REG_24__SCAN_IN), .S(n13811), .Z(
        P2_U3555) );
  MUX2_X1 U15978 ( .A(n13788), .B(P2_DATAO_REG_23__SCAN_IN), .S(n13811), .Z(
        P2_U3554) );
  MUX2_X1 U15979 ( .A(n13789), .B(P2_DATAO_REG_22__SCAN_IN), .S(n13811), .Z(
        P2_U3553) );
  MUX2_X1 U15980 ( .A(n13790), .B(P2_DATAO_REG_21__SCAN_IN), .S(n13811), .Z(
        P2_U3552) );
  MUX2_X1 U15981 ( .A(n13791), .B(P2_DATAO_REG_20__SCAN_IN), .S(n13811), .Z(
        P2_U3551) );
  MUX2_X1 U15982 ( .A(n13792), .B(P2_DATAO_REG_19__SCAN_IN), .S(n13811), .Z(
        P2_U3550) );
  MUX2_X1 U15983 ( .A(n13793), .B(P2_DATAO_REG_18__SCAN_IN), .S(n13811), .Z(
        P2_U3549) );
  MUX2_X1 U15984 ( .A(n13794), .B(P2_DATAO_REG_17__SCAN_IN), .S(n13811), .Z(
        P2_U3548) );
  MUX2_X1 U15985 ( .A(n13795), .B(P2_DATAO_REG_16__SCAN_IN), .S(n13811), .Z(
        P2_U3547) );
  MUX2_X1 U15986 ( .A(n13796), .B(P2_DATAO_REG_15__SCAN_IN), .S(n13811), .Z(
        P2_U3546) );
  MUX2_X1 U15987 ( .A(n13797), .B(P2_DATAO_REG_14__SCAN_IN), .S(n13811), .Z(
        P2_U3545) );
  MUX2_X1 U15988 ( .A(n13798), .B(P2_DATAO_REG_13__SCAN_IN), .S(n13811), .Z(
        P2_U3544) );
  MUX2_X1 U15989 ( .A(n13799), .B(P2_DATAO_REG_12__SCAN_IN), .S(n13811), .Z(
        P2_U3543) );
  MUX2_X1 U15990 ( .A(n13800), .B(P2_DATAO_REG_11__SCAN_IN), .S(n13811), .Z(
        P2_U3542) );
  MUX2_X1 U15991 ( .A(n13801), .B(P2_DATAO_REG_10__SCAN_IN), .S(n13811), .Z(
        P2_U3541) );
  MUX2_X1 U15992 ( .A(n13802), .B(P2_DATAO_REG_9__SCAN_IN), .S(n13811), .Z(
        P2_U3540) );
  MUX2_X1 U15993 ( .A(n13803), .B(P2_DATAO_REG_8__SCAN_IN), .S(n13811), .Z(
        P2_U3539) );
  MUX2_X1 U15994 ( .A(n13804), .B(P2_DATAO_REG_7__SCAN_IN), .S(n13811), .Z(
        P2_U3538) );
  MUX2_X1 U15995 ( .A(n13805), .B(P2_DATAO_REG_6__SCAN_IN), .S(n13811), .Z(
        P2_U3537) );
  MUX2_X1 U15996 ( .A(n13806), .B(P2_DATAO_REG_5__SCAN_IN), .S(n13811), .Z(
        P2_U3536) );
  MUX2_X1 U15997 ( .A(n13807), .B(P2_DATAO_REG_4__SCAN_IN), .S(n13811), .Z(
        P2_U3535) );
  MUX2_X1 U15998 ( .A(n13808), .B(P2_DATAO_REG_3__SCAN_IN), .S(n13811), .Z(
        P2_U3534) );
  MUX2_X1 U15999 ( .A(n13809), .B(P2_DATAO_REG_2__SCAN_IN), .S(n13811), .Z(
        P2_U3533) );
  MUX2_X1 U16000 ( .A(n13810), .B(P2_DATAO_REG_1__SCAN_IN), .S(n13811), .Z(
        P2_U3532) );
  MUX2_X1 U16001 ( .A(n13812), .B(P2_DATAO_REG_0__SCAN_IN), .S(n13811), .Z(
        P2_U3531) );
  OAI22_X1 U16002 ( .A1(n15857), .A2(n15586), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13813), .ZN(n13814) );
  AOI21_X1 U16003 ( .B1(n13815), .B2(n15850), .A(n13814), .ZN(n13824) );
  AND2_X1 U16004 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), 
        .ZN(n13817) );
  OAI211_X1 U16005 ( .C1(n13818), .C2(n13817), .A(n15830), .B(n13816), .ZN(
        n13823) );
  OAI211_X1 U16006 ( .C1(n13821), .C2(n13820), .A(n15866), .B(n13819), .ZN(
        n13822) );
  NAND3_X1 U16007 ( .A1(n13824), .A2(n13823), .A3(n13822), .ZN(P2_U3215) );
  AND2_X1 U16008 ( .A1(P2_U3088), .A2(P2_REG3_REG_4__SCAN_IN), .ZN(n13826) );
  NOR2_X1 U16009 ( .A1(n15871), .A2(n13830), .ZN(n13825) );
  AOI211_X1 U16010 ( .C1(n15864), .C2(P2_ADDR_REG_4__SCAN_IN), .A(n13826), .B(
        n13825), .ZN(n13836) );
  OAI211_X1 U16011 ( .C1(n13829), .C2(n13828), .A(n15830), .B(n13827), .ZN(
        n13835) );
  MUX2_X1 U16012 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n11504), .S(n13830), .Z(
        n13831) );
  NAND3_X1 U16013 ( .A1(n15837), .A2(n13832), .A3(n13831), .ZN(n13833) );
  NAND3_X1 U16014 ( .A1(n15866), .A2(n13845), .A3(n13833), .ZN(n13834) );
  NAND3_X1 U16015 ( .A1(n13836), .A2(n13835), .A3(n13834), .ZN(P2_U3218) );
  OAI21_X1 U16016 ( .B1(n15871), .B2(n13842), .A(n13837), .ZN(n13838) );
  AOI21_X1 U16017 ( .B1(n15864), .B2(P2_ADDR_REG_5__SCAN_IN), .A(n13838), .ZN(
        n13849) );
  OAI211_X1 U16018 ( .C1(n13841), .C2(n13840), .A(n15830), .B(n13839), .ZN(
        n13848) );
  MUX2_X1 U16019 ( .A(P2_REG2_REG_5__SCAN_IN), .B(n11929), .S(n13842), .Z(
        n13843) );
  NAND3_X1 U16020 ( .A1(n13845), .A2(n13844), .A3(n13843), .ZN(n13846) );
  NAND3_X1 U16021 ( .A1(n15866), .A2(n13860), .A3(n13846), .ZN(n13847) );
  NAND3_X1 U16022 ( .A1(n13849), .A2(n13848), .A3(n13847), .ZN(P2_U3219) );
  INV_X1 U16023 ( .A(n13850), .ZN(n13853) );
  NOR2_X1 U16024 ( .A1(n15871), .A2(n13851), .ZN(n13852) );
  AOI211_X1 U16025 ( .C1(n15864), .C2(P2_ADDR_REG_6__SCAN_IN), .A(n13853), .B(
        n13852), .ZN(n13864) );
  OAI211_X1 U16026 ( .C1(n13856), .C2(n13855), .A(n13854), .B(n15830), .ZN(
        n13863) );
  MUX2_X1 U16027 ( .A(n10678), .B(P2_REG2_REG_6__SCAN_IN), .S(n13857), .Z(
        n13858) );
  NAND3_X1 U16028 ( .A1(n13860), .A2(n13859), .A3(n13858), .ZN(n13861) );
  NAND3_X1 U16029 ( .A1(n15866), .A2(n13874), .A3(n13861), .ZN(n13862) );
  NAND3_X1 U16030 ( .A1(n13864), .A2(n13863), .A3(n13862), .ZN(P2_U3220) );
  OAI211_X1 U16031 ( .C1(n13867), .C2(n13866), .A(n13865), .B(n15830), .ZN(
        n13879) );
  AND2_X1 U16032 ( .A1(P2_U3088), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n13870) );
  NOR2_X1 U16033 ( .A1(n15871), .A2(n13868), .ZN(n13869) );
  AOI211_X1 U16034 ( .C1(n15864), .C2(P2_ADDR_REG_7__SCAN_IN), .A(n13870), .B(
        n13869), .ZN(n13878) );
  MUX2_X1 U16035 ( .A(n12068), .B(P2_REG2_REG_7__SCAN_IN), .S(n13871), .Z(
        n13872) );
  NAND3_X1 U16036 ( .A1(n13874), .A2(n13873), .A3(n13872), .ZN(n13875) );
  NAND3_X1 U16037 ( .A1(n15866), .A2(n13876), .A3(n13875), .ZN(n13877) );
  NAND3_X1 U16038 ( .A1(n13879), .A2(n13878), .A3(n13877), .ZN(P2_U3221) );
  NAND2_X1 U16039 ( .A1(n13880), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n13883) );
  NAND2_X1 U16040 ( .A1(n13881), .A2(n13885), .ZN(n13882) );
  NAND2_X1 U16041 ( .A1(n13883), .A2(n13882), .ZN(n13894) );
  XNOR2_X1 U16042 ( .A(n13894), .B(n13901), .ZN(n13892) );
  XNOR2_X1 U16043 ( .A(n13892), .B(P2_REG2_REG_15__SCAN_IN), .ZN(n13891) );
  NAND2_X1 U16044 ( .A1(n13886), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n13900) );
  OAI211_X1 U16045 ( .C1(n13886), .C2(P2_REG1_REG_15__SCAN_IN), .A(n13900), 
        .B(n15830), .ZN(n13890) );
  AND2_X1 U16046 ( .A1(P2_U3088), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n13888) );
  NOR2_X1 U16047 ( .A1(n15871), .A2(n13901), .ZN(n13887) );
  AOI211_X1 U16048 ( .C1(n15864), .C2(P2_ADDR_REG_15__SCAN_IN), .A(n13888), 
        .B(n13887), .ZN(n13889) );
  OAI211_X1 U16049 ( .C1(n13891), .C2(n15823), .A(n13890), .B(n13889), .ZN(
        P2_U3229) );
  NAND2_X1 U16050 ( .A1(n13892), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n13896) );
  NAND2_X1 U16051 ( .A1(n13894), .A2(n13893), .ZN(n13895) );
  NAND2_X1 U16052 ( .A1(n13896), .A2(n13895), .ZN(n13898) );
  INV_X1 U16053 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n14150) );
  MUX2_X1 U16054 ( .A(n14150), .B(P2_REG2_REG_16__SCAN_IN), .S(n13916), .Z(
        n13897) );
  OAI21_X1 U16055 ( .B1(n13898), .B2(n13897), .A(n15866), .ZN(n13910) );
  OAI21_X1 U16056 ( .B1(n15857), .B2(n15697), .A(n13899), .ZN(n13907) );
  OAI21_X1 U16057 ( .B1(n13902), .B2(n13901), .A(n13900), .ZN(n13904) );
  XNOR2_X1 U16058 ( .A(n13916), .B(P2_REG1_REG_16__SCAN_IN), .ZN(n13903) );
  OAI211_X1 U16059 ( .C1(n13904), .C2(n13903), .A(n13911), .B(n15830), .ZN(
        n13905) );
  INV_X1 U16060 ( .A(n13905), .ZN(n13906) );
  AOI211_X1 U16061 ( .C1(n15850), .C2(n13908), .A(n13907), .B(n13906), .ZN(
        n13909) );
  OAI21_X1 U16062 ( .B1(n13923), .B2(n13910), .A(n13909), .ZN(P2_U3230) );
  INV_X1 U16063 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n14347) );
  XOR2_X1 U16064 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n13936), .Z(n13912) );
  OAI21_X1 U16065 ( .B1(n13913), .B2(n13912), .A(n15830), .ZN(n13926) );
  AND2_X1 U16066 ( .A1(P2_U3088), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n13915) );
  NOR2_X1 U16067 ( .A1(n15871), .A2(n13928), .ZN(n13914) );
  AOI211_X1 U16068 ( .C1(n15864), .C2(P2_ADDR_REG_17__SCAN_IN), .A(n13915), 
        .B(n13914), .ZN(n13925) );
  NOR2_X1 U16069 ( .A1(n13916), .A2(n14150), .ZN(n13921) );
  INV_X1 U16070 ( .A(n13921), .ZN(n13918) );
  NAND2_X1 U16071 ( .A1(n13928), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n13917) );
  OAI211_X1 U16072 ( .C1(P2_REG2_REG_17__SCAN_IN), .C2(n13928), .A(n13918), 
        .B(n13917), .ZN(n13922) );
  NAND2_X1 U16073 ( .A1(n13936), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n13920) );
  INV_X1 U16074 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n13929) );
  NAND2_X1 U16075 ( .A1(n13928), .A2(n13929), .ZN(n13919) );
  OAI211_X1 U16076 ( .C1(n13923), .C2(n13922), .A(n13927), .B(n15866), .ZN(
        n13924) );
  OAI211_X1 U16077 ( .C1(n13926), .C2(n13935), .A(n13925), .B(n13924), .ZN(
        P2_U3231) );
  OAI21_X1 U16078 ( .B1(n13929), .B2(n13928), .A(n13927), .ZN(n13930) );
  NOR2_X1 U16079 ( .A1(n13930), .A2(n13931), .ZN(n13934) );
  INV_X1 U16080 ( .A(n15865), .ZN(n13932) );
  NOR2_X1 U16081 ( .A1(n13932), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n13933) );
  XNOR2_X1 U16082 ( .A(n13938), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n13940) );
  AOI22_X1 U16083 ( .A1(n13941), .A2(n15866), .B1(n15830), .B2(n13940), .ZN(
        n13942) );
  NOR2_X1 U16084 ( .A1(n14210), .A2(n14280), .ZN(n13951) );
  NOR2_X1 U16085 ( .A1(n13945), .A2(n14251), .ZN(n13946) );
  AOI211_X1 U16086 ( .C1(P2_REG2_REG_31__SCAN_IN), .C2(n14210), .A(n13951), 
        .B(n13946), .ZN(n13947) );
  OAI21_X1 U16087 ( .B1(n13948), .B2(n14267), .A(n13947), .ZN(P2_U3234) );
  AOI21_X1 U16088 ( .B1(n12390), .B2(n14401), .A(n15891), .ZN(n13950) );
  NAND2_X1 U16089 ( .A1(n13950), .A2(n13949), .ZN(n14281) );
  AOI21_X1 U16090 ( .B1(n14275), .B2(P2_REG2_REG_30__SCAN_IN), .A(n13951), 
        .ZN(n13953) );
  NAND2_X1 U16091 ( .A1(n14401), .A2(n14265), .ZN(n13952) );
  OAI211_X1 U16092 ( .C1(n14281), .C2(n14267), .A(n13953), .B(n13952), .ZN(
        P2_U3235) );
  AOI21_X1 U16093 ( .B1(n13955), .B2(n10189), .A(n13954), .ZN(n13957) );
  XNOR2_X1 U16094 ( .A(n13957), .B(n13956), .ZN(n13967) );
  NOR2_X1 U16095 ( .A1(n13958), .A2(n14267), .ZN(n13964) );
  INV_X1 U16096 ( .A(n13959), .ZN(n13960) );
  AOI22_X1 U16097 ( .A1(n13960), .A2(n14263), .B1(P2_REG2_REG_29__SCAN_IN), 
        .B2(n14275), .ZN(n13961) );
  OAI21_X1 U16098 ( .B1(n13962), .B2(n14251), .A(n13961), .ZN(n13963) );
  AOI211_X1 U16099 ( .C1(n13965), .C2(n14231), .A(n13964), .B(n13963), .ZN(
        n13966) );
  OAI21_X1 U16100 ( .B1(n13967), .B2(n14256), .A(n13966), .ZN(P2_U3236) );
  INV_X1 U16101 ( .A(n13968), .ZN(n13969) );
  AOI22_X1 U16102 ( .A1(n13972), .A2(n14265), .B1(n14275), .B2(
        P2_REG2_REG_28__SCAN_IN), .ZN(n13975) );
  NAND2_X1 U16103 ( .A1(n13973), .A2(n14278), .ZN(n13974) );
  XNOR2_X1 U16104 ( .A(n13976), .B(n7933), .ZN(n13978) );
  OAI21_X1 U16105 ( .B1(n13981), .B2(n13980), .A(n13979), .ZN(n14286) );
  INV_X1 U16106 ( .A(n14286), .ZN(n13987) );
  AOI21_X1 U16107 ( .B1(n13997), .B2(n14405), .A(n15891), .ZN(n13982) );
  NAND2_X1 U16108 ( .A1(n6538), .A2(n13982), .ZN(n14284) );
  OAI22_X1 U16109 ( .A1(n13983), .A2(n14250), .B1(n9402), .B2(n14231), .ZN(
        n13984) );
  AOI21_X1 U16110 ( .B1(n14405), .B2(n14265), .A(n13984), .ZN(n13985) );
  OAI21_X1 U16111 ( .B1(n14284), .B2(n14267), .A(n13985), .ZN(n13986) );
  AOI21_X1 U16112 ( .B1(n13987), .B2(n14278), .A(n13986), .ZN(n13988) );
  OAI21_X1 U16113 ( .B1(n14285), .B2(n14210), .A(n13988), .ZN(P2_U3238) );
  INV_X1 U16114 ( .A(n14288), .ZN(n14003) );
  NAND2_X1 U16115 ( .A1(n13992), .A2(n13991), .ZN(n13994) );
  XNOR2_X1 U16116 ( .A(n13994), .B(n13993), .ZN(n14290) );
  AOI21_X1 U16117 ( .B1(n14006), .B2(n13995), .A(n15891), .ZN(n13996) );
  AND2_X1 U16118 ( .A1(n13997), .A2(n13996), .ZN(n14289) );
  NAND2_X1 U16119 ( .A1(n14289), .A2(n14253), .ZN(n14000) );
  AOI22_X1 U16120 ( .A1(n13998), .A2(n14263), .B1(P2_REG2_REG_26__SCAN_IN), 
        .B2(n14275), .ZN(n13999) );
  OAI211_X1 U16121 ( .C1(n6888), .C2(n14251), .A(n14000), .B(n13999), .ZN(
        n14001) );
  AOI21_X1 U16122 ( .B1(n14290), .B2(n14278), .A(n14001), .ZN(n14002) );
  OAI21_X1 U16123 ( .B1(n14003), .B2(n14275), .A(n14002), .ZN(P2_U3239) );
  XOR2_X1 U16124 ( .A(n14013), .B(n14004), .Z(n14297) );
  AOI21_X1 U16125 ( .B1(n14005), .B2(n7352), .A(n15891), .ZN(n14007) );
  AND2_X1 U16126 ( .A1(n14006), .A2(n14007), .ZN(n14294) );
  NOR2_X1 U16127 ( .A1(n14008), .A2(n14251), .ZN(n14012) );
  OAI22_X1 U16128 ( .A1(n14010), .A2(n14250), .B1(n14231), .B2(n14009), .ZN(
        n14011) );
  AOI211_X1 U16129 ( .C1(n14294), .C2(n14253), .A(n14012), .B(n14011), .ZN(
        n14016) );
  NAND2_X1 U16130 ( .A1(n14293), .A2(n14231), .ZN(n14015) );
  OAI211_X1 U16131 ( .C1(n14297), .C2(n14256), .A(n14016), .B(n14015), .ZN(
        P2_U3240) );
  XNOR2_X1 U16132 ( .A(n14017), .B(n7644), .ZN(n14024) );
  NAND2_X1 U16133 ( .A1(n14019), .A2(n14018), .ZN(n14020) );
  NAND2_X1 U16134 ( .A1(n14021), .A2(n14020), .ZN(n14302) );
  OAI21_X1 U16135 ( .B1(n14302), .B2(n11003), .A(n14022), .ZN(n14023) );
  INV_X1 U16136 ( .A(n14025), .ZN(n14038) );
  AOI211_X1 U16137 ( .C1(n7324), .C2(n14038), .A(n15891), .B(n7355), .ZN(
        n14298) );
  AOI22_X1 U16138 ( .A1(n14026), .A2(n14263), .B1(P2_REG2_REG_24__SCAN_IN), 
        .B2(n14275), .ZN(n14027) );
  OAI21_X1 U16139 ( .B1(n14028), .B2(n14251), .A(n14027), .ZN(n14030) );
  NOR2_X1 U16140 ( .A1(n14302), .A2(n14200), .ZN(n14029) );
  AOI211_X1 U16141 ( .C1(n14298), .C2(n14253), .A(n14030), .B(n14029), .ZN(
        n14031) );
  OAI21_X1 U16142 ( .B1(n14275), .B2(n14301), .A(n14031), .ZN(P2_U3241) );
  XNOR2_X1 U16143 ( .A(n14032), .B(n14034), .ZN(n14309) );
  INV_X1 U16144 ( .A(n14309), .ZN(n14045) );
  INV_X1 U16145 ( .A(n14033), .ZN(n14037) );
  XNOR2_X1 U16146 ( .A(n14035), .B(n14034), .ZN(n14036) );
  NAND2_X1 U16147 ( .A1(n14036), .A2(n14270), .ZN(n14305) );
  OAI211_X1 U16148 ( .C1(n14250), .C2(n14037), .A(n14305), .B(n14304), .ZN(
        n14043) );
  OAI21_X1 U16149 ( .B1(n14414), .B2(n14050), .A(n14038), .ZN(n14306) );
  AOI22_X1 U16150 ( .A1(n14039), .A2(n14265), .B1(n14275), .B2(
        P2_REG2_REG_23__SCAN_IN), .ZN(n14040) );
  OAI21_X1 U16151 ( .B1(n14306), .B2(n14041), .A(n14040), .ZN(n14042) );
  AOI21_X1 U16152 ( .B1(n14043), .B2(n14231), .A(n14042), .ZN(n14044) );
  OAI21_X1 U16153 ( .B1(n14045), .B2(n14256), .A(n14044), .ZN(P2_U3242) );
  NAND2_X1 U16154 ( .A1(n14047), .A2(n14046), .ZN(n14048) );
  XNOR2_X1 U16155 ( .A(n14048), .B(n10181), .ZN(n14312) );
  NAND2_X1 U16156 ( .A1(n14070), .A2(n14417), .ZN(n14049) );
  NAND2_X1 U16157 ( .A1(n14049), .A2(n14261), .ZN(n14051) );
  OR2_X1 U16158 ( .A1(n14051), .A2(n14050), .ZN(n14313) );
  INV_X1 U16159 ( .A(n14052), .ZN(n14053) );
  AOI22_X1 U16160 ( .A1(P2_REG2_REG_22__SCAN_IN), .A2(n14275), .B1(n14053), 
        .B2(n14263), .ZN(n14055) );
  NAND2_X1 U16161 ( .A1(n14417), .A2(n14265), .ZN(n14054) );
  OAI211_X1 U16162 ( .C1(n14313), .C2(n14267), .A(n14055), .B(n14054), .ZN(
        n14061) );
  XNOR2_X1 U16163 ( .A(n14057), .B(n14056), .ZN(n14059) );
  AOI21_X1 U16164 ( .B1(n14059), .B2(n14270), .A(n14058), .ZN(n14314) );
  NOR2_X1 U16165 ( .A1(n14314), .A2(n14275), .ZN(n14060) );
  AOI211_X1 U16166 ( .C1(n14312), .C2(n14278), .A(n14061), .B(n14060), .ZN(
        n14062) );
  INV_X1 U16167 ( .A(n14062), .ZN(P2_U3243) );
  OR2_X1 U16168 ( .A1(n14063), .A2(n14080), .ZN(n14077) );
  NAND2_X1 U16169 ( .A1(n14077), .A2(n14064), .ZN(n14065) );
  XOR2_X1 U16170 ( .A(n14065), .B(n14066), .Z(n14322) );
  XNOR2_X1 U16171 ( .A(n14067), .B(n14066), .ZN(n14069) );
  OAI21_X1 U16172 ( .B1(n14069), .B2(n14127), .A(n14068), .ZN(n14318) );
  INV_X1 U16173 ( .A(n14070), .ZN(n14071) );
  AOI211_X1 U16174 ( .C1(n14320), .C2(n6885), .A(n15891), .B(n14071), .ZN(
        n14319) );
  NAND2_X1 U16175 ( .A1(n14319), .A2(n14253), .ZN(n14074) );
  AOI22_X1 U16176 ( .A1(n14210), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n14072), 
        .B2(n14263), .ZN(n14073) );
  OAI211_X1 U16177 ( .C1(n10202), .C2(n14251), .A(n14074), .B(n14073), .ZN(
        n14075) );
  AOI21_X1 U16178 ( .B1(n14318), .B2(n14231), .A(n14075), .ZN(n14076) );
  OAI21_X1 U16179 ( .B1(n14322), .B2(n14256), .A(n14076), .ZN(P2_U3244) );
  INV_X1 U16180 ( .A(n14063), .ZN(n14079) );
  INV_X1 U16181 ( .A(n14080), .ZN(n14078) );
  OAI21_X1 U16182 ( .B1(n14079), .B2(n14078), .A(n14077), .ZN(n14327) );
  XOR2_X1 U16183 ( .A(n14081), .B(n14080), .Z(n14083) );
  OAI21_X1 U16184 ( .B1(n14083), .B2(n14127), .A(n14082), .ZN(n14323) );
  INV_X1 U16185 ( .A(n14084), .ZN(n14085) );
  AOI211_X1 U16186 ( .C1(n14325), .C2(n14085), .A(n15891), .B(n10203), .ZN(
        n14324) );
  NAND2_X1 U16187 ( .A1(n14324), .A2(n14253), .ZN(n14088) );
  AOI22_X1 U16188 ( .A1(n14210), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n14086), 
        .B2(n14263), .ZN(n14087) );
  OAI211_X1 U16189 ( .C1(n7668), .C2(n14251), .A(n14088), .B(n14087), .ZN(
        n14089) );
  AOI21_X1 U16190 ( .B1(n14323), .B2(n14231), .A(n14089), .ZN(n14090) );
  OAI21_X1 U16191 ( .B1(n14327), .B2(n14256), .A(n14090), .ZN(P2_U3245) );
  XNOR2_X1 U16192 ( .A(n14091), .B(n14094), .ZN(n14093) );
  OAI21_X1 U16193 ( .B1(n14093), .B2(n14127), .A(n14092), .ZN(n14328) );
  INV_X1 U16194 ( .A(n14328), .ZN(n14104) );
  XOR2_X1 U16195 ( .A(n14094), .B(n14095), .Z(n14330) );
  NAND2_X1 U16196 ( .A1(n14330), .A2(n14278), .ZN(n14103) );
  INV_X1 U16197 ( .A(n14114), .ZN(n14096) );
  AOI211_X1 U16198 ( .C1(n14097), .C2(n14096), .A(n15891), .B(n14084), .ZN(
        n14329) );
  NOR2_X1 U16199 ( .A1(n14424), .A2(n14251), .ZN(n14101) );
  OAI22_X1 U16200 ( .A1(n14231), .A2(n14099), .B1(n14098), .B2(n14250), .ZN(
        n14100) );
  AOI211_X1 U16201 ( .C1(n14329), .C2(n14253), .A(n14101), .B(n14100), .ZN(
        n14102) );
  OAI211_X1 U16202 ( .C1(n14275), .C2(n14104), .A(n14103), .B(n14102), .ZN(
        P2_U3246) );
  XNOR2_X1 U16203 ( .A(n14106), .B(n14105), .ZN(n14108) );
  AOI21_X1 U16204 ( .B1(n14108), .B2(n14270), .A(n14107), .ZN(n14337) );
  OAI21_X1 U16205 ( .B1(n14111), .B2(n14110), .A(n14109), .ZN(n14333) );
  NAND2_X1 U16206 ( .A1(n14129), .A2(n14335), .ZN(n14112) );
  NAND2_X1 U16207 ( .A1(n14112), .A2(n14261), .ZN(n14113) );
  NOR2_X1 U16208 ( .A1(n14114), .A2(n14113), .ZN(n14334) );
  NAND2_X1 U16209 ( .A1(n14334), .A2(n14253), .ZN(n14117) );
  AOI22_X1 U16210 ( .A1(n14210), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n14115), 
        .B2(n14263), .ZN(n14116) );
  OAI211_X1 U16211 ( .C1(n14118), .C2(n14251), .A(n14117), .B(n14116), .ZN(
        n14119) );
  AOI21_X1 U16212 ( .B1(n14333), .B2(n14278), .A(n14119), .ZN(n14120) );
  OAI21_X1 U16213 ( .B1(n14275), .B2(n14337), .A(n14120), .ZN(P2_U3247) );
  XOR2_X1 U16214 ( .A(n14124), .B(n14121), .Z(n14343) );
  NAND2_X1 U16215 ( .A1(n14160), .A2(n14159), .ZN(n14158) );
  AND2_X1 U16216 ( .A1(n14158), .A2(n14122), .ZN(n14138) );
  NAND2_X1 U16217 ( .A1(n14138), .A2(n14145), .ZN(n14137) );
  NAND2_X1 U16218 ( .A1(n14137), .A2(n14123), .ZN(n14125) );
  XNOR2_X1 U16219 ( .A(n14125), .B(n14124), .ZN(n14128) );
  OAI21_X1 U16220 ( .B1(n14128), .B2(n14127), .A(n14126), .ZN(n14339) );
  NAND2_X1 U16221 ( .A1(n14339), .A2(n14231), .ZN(n14136) );
  INV_X1 U16222 ( .A(n14129), .ZN(n14130) );
  AOI211_X1 U16223 ( .C1(n14341), .C2(n14146), .A(n15891), .B(n14130), .ZN(
        n14340) );
  INV_X1 U16224 ( .A(n14341), .ZN(n14131) );
  NOR2_X1 U16225 ( .A1(n14131), .A2(n14251), .ZN(n14134) );
  OAI22_X1 U16226 ( .A1(n14231), .A2(n13929), .B1(n14132), .B2(n14250), .ZN(
        n14133) );
  AOI211_X1 U16227 ( .C1(n14340), .C2(n14253), .A(n14134), .B(n14133), .ZN(
        n14135) );
  OAI211_X1 U16228 ( .C1(n14343), .C2(n14256), .A(n14136), .B(n14135), .ZN(
        P2_U3248) );
  OAI211_X1 U16229 ( .C1(n14138), .C2(n14145), .A(n14137), .B(n14270), .ZN(
        n14141) );
  INV_X1 U16230 ( .A(n14139), .ZN(n14140) );
  NAND2_X1 U16231 ( .A1(n14141), .A2(n14140), .ZN(n14344) );
  INV_X1 U16232 ( .A(n14344), .ZN(n14155) );
  INV_X1 U16233 ( .A(n6741), .ZN(n14143) );
  AOI21_X1 U16234 ( .B1(n14145), .B2(n14144), .A(n14143), .ZN(n14346) );
  NAND2_X1 U16235 ( .A1(n14346), .A2(n14278), .ZN(n14154) );
  INV_X1 U16236 ( .A(n14163), .ZN(n14147) );
  AOI211_X1 U16237 ( .C1(n14148), .C2(n14147), .A(n15891), .B(n10201), .ZN(
        n14345) );
  NOR2_X1 U16238 ( .A1(n14431), .A2(n14251), .ZN(n14152) );
  OAI22_X1 U16239 ( .A1(n14231), .A2(n14150), .B1(n14149), .B2(n14250), .ZN(
        n14151) );
  AOI211_X1 U16240 ( .C1(n14345), .C2(n14253), .A(n14152), .B(n14151), .ZN(
        n14153) );
  OAI211_X1 U16241 ( .C1(n14155), .C2(n14210), .A(n14154), .B(n14153), .ZN(
        P2_U3249) );
  XNOR2_X1 U16242 ( .A(n14157), .B(n14159), .ZN(n14354) );
  OAI21_X1 U16243 ( .B1(n14160), .B2(n14159), .A(n14158), .ZN(n14162) );
  AOI21_X1 U16244 ( .B1(n14162), .B2(n14270), .A(n14161), .ZN(n14353) );
  AOI211_X1 U16245 ( .C1(n14351), .C2(n14176), .A(n15891), .B(n14163), .ZN(
        n14350) );
  NAND2_X1 U16246 ( .A1(n14350), .A2(n14164), .ZN(n14165) );
  OAI211_X1 U16247 ( .C1(n14250), .C2(n14166), .A(n14353), .B(n14165), .ZN(
        n14167) );
  NAND2_X1 U16248 ( .A1(n14167), .A2(n14231), .ZN(n14169) );
  AOI22_X1 U16249 ( .A1(n14351), .A2(n14265), .B1(P2_REG2_REG_15__SCAN_IN), 
        .B2(n14210), .ZN(n14168) );
  OAI211_X1 U16250 ( .C1(n14354), .C2(n14256), .A(n14169), .B(n14168), .ZN(
        P2_U3250) );
  XNOR2_X1 U16251 ( .A(n14170), .B(n14180), .ZN(n14172) );
  AOI21_X1 U16252 ( .B1(n14172), .B2(n14270), .A(n14171), .ZN(n14356) );
  INV_X1 U16253 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n14174) );
  OAI22_X1 U16254 ( .A1(n14231), .A2(n14174), .B1(n14173), .B2(n14250), .ZN(
        n14179) );
  AOI21_X1 U16255 ( .B1(n14175), .B2(n14435), .A(n15891), .ZN(n14177) );
  NAND2_X1 U16256 ( .A1(n14177), .A2(n14176), .ZN(n14355) );
  NOR2_X1 U16257 ( .A1(n14355), .A2(n14267), .ZN(n14178) );
  AOI211_X1 U16258 ( .C1(n14265), .C2(n14435), .A(n14179), .B(n14178), .ZN(
        n14183) );
  XNOR2_X1 U16259 ( .A(n14181), .B(n14180), .ZN(n14357) );
  OR2_X1 U16260 ( .A1(n14357), .A2(n14256), .ZN(n14182) );
  OAI211_X1 U16261 ( .C1(n14356), .C2(n14210), .A(n14183), .B(n14182), .ZN(
        P2_U3251) );
  XNOR2_X1 U16262 ( .A(n14184), .B(n14188), .ZN(n14365) );
  INV_X1 U16263 ( .A(n14365), .ZN(n14201) );
  NAND2_X1 U16264 ( .A1(n14365), .A2(n14185), .ZN(n14193) );
  NAND2_X1 U16265 ( .A1(n14186), .A2(n14187), .ZN(n14189) );
  XNOR2_X1 U16266 ( .A(n14189), .B(n14188), .ZN(n14190) );
  NAND2_X1 U16267 ( .A1(n14190), .A2(n14270), .ZN(n14191) );
  NAND3_X1 U16268 ( .A1(n14193), .A2(n14192), .A3(n14191), .ZN(n14370) );
  NAND2_X1 U16269 ( .A1(n14370), .A2(n14231), .ZN(n14199) );
  OAI22_X1 U16270 ( .A1(n14231), .A2(n11827), .B1(n14194), .B2(n14250), .ZN(
        n14196) );
  OAI211_X1 U16271 ( .C1(n14208), .C2(n14368), .A(n14261), .B(n12360), .ZN(
        n14366) );
  NOR2_X1 U16272 ( .A1(n14366), .A2(n14267), .ZN(n14195) );
  AOI211_X1 U16273 ( .C1(n14265), .C2(n14197), .A(n14196), .B(n14195), .ZN(
        n14198) );
  OAI211_X1 U16274 ( .C1(n14201), .C2(n14200), .A(n14199), .B(n14198), .ZN(
        P2_U3253) );
  INV_X1 U16275 ( .A(n14204), .ZN(n14202) );
  XNOR2_X1 U16276 ( .A(n14203), .B(n14202), .ZN(n14375) );
  OAI21_X1 U16277 ( .B1(n6717), .B2(n14204), .A(n14186), .ZN(n14206) );
  AOI21_X1 U16278 ( .B1(n14206), .B2(n14270), .A(n14205), .ZN(n14374) );
  INV_X1 U16279 ( .A(n14374), .ZN(n14216) );
  OAI21_X1 U16280 ( .B1(n14233), .B2(n14207), .A(n14261), .ZN(n14209) );
  OR2_X1 U16281 ( .A1(n14209), .A2(n14208), .ZN(n14373) );
  NAND2_X1 U16282 ( .A1(n14210), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n14211) );
  OAI21_X1 U16283 ( .B1(n14250), .B2(n14212), .A(n14211), .ZN(n14213) );
  AOI21_X1 U16284 ( .B1(n14443), .B2(n14265), .A(n14213), .ZN(n14214) );
  OAI21_X1 U16285 ( .B1(n14373), .B2(n14267), .A(n14214), .ZN(n14215) );
  AOI21_X1 U16286 ( .B1(n14216), .B2(n14231), .A(n14215), .ZN(n14217) );
  OAI21_X1 U16287 ( .B1(n14256), .B2(n14375), .A(n14217), .ZN(P2_U3254) );
  OR2_X1 U16288 ( .A1(n14219), .A2(n14218), .ZN(n14220) );
  NAND2_X1 U16289 ( .A1(n14221), .A2(n14220), .ZN(n14382) );
  NAND2_X1 U16290 ( .A1(n14244), .A2(n14243), .ZN(n14242) );
  NAND2_X1 U16291 ( .A1(n14242), .A2(n14223), .ZN(n14225) );
  XNOR2_X1 U16292 ( .A(n14225), .B(n14224), .ZN(n14226) );
  NAND2_X1 U16293 ( .A1(n14226), .A2(n14270), .ZN(n14228) );
  NAND2_X1 U16294 ( .A1(n14228), .A2(n14227), .ZN(n14384) );
  NAND2_X1 U16295 ( .A1(n14384), .A2(n14231), .ZN(n14238) );
  OAI22_X1 U16296 ( .A1(n14231), .A2(n14230), .B1(n14229), .B2(n14250), .ZN(
        n14236) );
  NAND2_X1 U16297 ( .A1(n14247), .A2(n14379), .ZN(n14232) );
  NAND2_X1 U16298 ( .A1(n14232), .A2(n14261), .ZN(n14234) );
  OR2_X1 U16299 ( .A1(n14234), .A2(n14233), .ZN(n14381) );
  NOR2_X1 U16300 ( .A1(n14381), .A2(n14267), .ZN(n14235) );
  AOI211_X1 U16301 ( .C1(n14265), .C2(n14379), .A(n14236), .B(n14235), .ZN(
        n14237) );
  OAI211_X1 U16302 ( .C1(n14256), .C2(n14382), .A(n14238), .B(n14237), .ZN(
        P2_U3255) );
  OAI21_X1 U16303 ( .B1(n14241), .B2(n14240), .A(n14239), .ZN(n14390) );
  OAI21_X1 U16304 ( .B1(n14244), .B2(n14243), .A(n14242), .ZN(n14246) );
  AOI21_X1 U16305 ( .B1(n14246), .B2(n14270), .A(n14245), .ZN(n14389) );
  MUX2_X1 U16306 ( .A(n14389), .B(n10881), .S(n14275), .Z(n14255) );
  INV_X1 U16307 ( .A(n14247), .ZN(n14248) );
  AOI211_X1 U16308 ( .C1(n14386), .C2(n14260), .A(n15891), .B(n14248), .ZN(
        n14385) );
  OAI22_X1 U16309 ( .A1(n10198), .A2(n14251), .B1(n14250), .B2(n14249), .ZN(
        n14252) );
  AOI21_X1 U16310 ( .B1(n14385), .B2(n14253), .A(n14252), .ZN(n14254) );
  OAI211_X1 U16311 ( .C1(n14256), .C2(n14390), .A(n14255), .B(n14254), .ZN(
        P2_U3256) );
  INV_X1 U16312 ( .A(n14257), .ZN(n14258) );
  AOI21_X1 U16313 ( .B1(n14271), .B2(n14259), .A(n14258), .ZN(n14397) );
  OAI211_X1 U16314 ( .C1(n12024), .C2(n14393), .A(n14261), .B(n14260), .ZN(
        n14392) );
  AOI22_X1 U16315 ( .A1(n14265), .A2(n14264), .B1(n14263), .B2(n14262), .ZN(
        n14266) );
  OAI21_X1 U16316 ( .B1(n14392), .B2(n14267), .A(n14266), .ZN(n14277) );
  INV_X1 U16317 ( .A(n14268), .ZN(n14272) );
  OAI211_X1 U16318 ( .C1(n14272), .C2(n14271), .A(n14270), .B(n14269), .ZN(
        n14274) );
  NAND2_X1 U16319 ( .A1(n14274), .A2(n14273), .ZN(n14394) );
  MUX2_X1 U16320 ( .A(n14394), .B(P2_REG2_REG_8__SCAN_IN), .S(n14275), .Z(
        n14276) );
  AOI211_X1 U16321 ( .C1(n14397), .C2(n14278), .A(n14277), .B(n14276), .ZN(
        n14279) );
  INV_X1 U16322 ( .A(n14279), .ZN(P2_U3257) );
  NAND2_X1 U16323 ( .A1(n14281), .A2(n14280), .ZN(n14399) );
  MUX2_X1 U16324 ( .A(n14399), .B(P2_REG1_REG_30__SCAN_IN), .S(n15910), .Z(
        n14282) );
  AOI21_X1 U16325 ( .B1(n14377), .B2(n14401), .A(n14282), .ZN(n14283) );
  INV_X1 U16326 ( .A(n14283), .ZN(P2_U3529) );
  OAI211_X1 U16327 ( .C1(n14286), .C2(n14391), .A(n14285), .B(n14284), .ZN(
        n14403) );
  MUX2_X1 U16328 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n14403), .S(n15912), .Z(
        n14287) );
  INV_X1 U16329 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n14291) );
  MUX2_X1 U16330 ( .A(n14291), .B(n14406), .S(n15912), .Z(n14292) );
  OAI21_X1 U16331 ( .B1(n14391), .B2(n14297), .A(n14296), .ZN(n14409) );
  MUX2_X1 U16332 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n14409), .S(n15912), .Z(
        P2_U3524) );
  AOI21_X1 U16333 ( .B1(n14387), .B2(n7324), .A(n14298), .ZN(n14300) );
  OAI211_X1 U16334 ( .C1(n14303), .C2(n14302), .A(n14301), .B(n14300), .ZN(
        n14410) );
  MUX2_X1 U16335 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n14410), .S(n15912), .Z(
        P2_U3523) );
  INV_X1 U16336 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n14310) );
  OAI211_X1 U16337 ( .C1(n14307), .C2(n14306), .A(n14305), .B(n14304), .ZN(
        n14308) );
  AOI21_X1 U16338 ( .B1(n14396), .B2(n14309), .A(n14308), .ZN(n14411) );
  MUX2_X1 U16339 ( .A(n14310), .B(n14411), .S(n15912), .Z(n14311) );
  OAI21_X1 U16340 ( .B1(n14414), .B2(n14349), .A(n14311), .ZN(P2_U3522) );
  NAND2_X1 U16341 ( .A1(n14312), .A2(n14396), .ZN(n14315) );
  NAND3_X1 U16342 ( .A1(n14315), .A2(n14314), .A3(n14313), .ZN(n14415) );
  MUX2_X1 U16343 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n14415), .S(n15912), .Z(
        n14316) );
  AOI21_X1 U16344 ( .B1(n14377), .B2(n14417), .A(n14316), .ZN(n14317) );
  INV_X1 U16345 ( .A(n14317), .ZN(P2_U3521) );
  AOI211_X1 U16346 ( .C1(n14387), .C2(n14320), .A(n14319), .B(n14318), .ZN(
        n14321) );
  OAI21_X1 U16347 ( .B1(n14322), .B2(n14391), .A(n14321), .ZN(n14419) );
  MUX2_X1 U16348 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n14419), .S(n15912), .Z(
        P2_U3520) );
  AOI211_X1 U16349 ( .C1(n14387), .C2(n14325), .A(n14324), .B(n14323), .ZN(
        n14326) );
  OAI21_X1 U16350 ( .B1(n14391), .B2(n14327), .A(n14326), .ZN(n14420) );
  MUX2_X1 U16351 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n14420), .S(n15912), .Z(
        P2_U3519) );
  INV_X1 U16352 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n14331) );
  AOI211_X1 U16353 ( .C1(n14330), .C2(n14396), .A(n14329), .B(n14328), .ZN(
        n14421) );
  MUX2_X1 U16354 ( .A(n14331), .B(n14421), .S(n15912), .Z(n14332) );
  OAI21_X1 U16355 ( .B1(n14424), .B2(n14349), .A(n14332), .ZN(P2_U3518) );
  INV_X1 U16356 ( .A(n14333), .ZN(n14338) );
  AOI21_X1 U16357 ( .B1(n14387), .B2(n14335), .A(n14334), .ZN(n14336) );
  OAI211_X1 U16358 ( .C1(n14338), .C2(n14391), .A(n14337), .B(n14336), .ZN(
        n14425) );
  MUX2_X1 U16359 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n14425), .S(n15912), .Z(
        P2_U3517) );
  AOI211_X1 U16360 ( .C1(n14387), .C2(n14341), .A(n14340), .B(n14339), .ZN(
        n14342) );
  OAI21_X1 U16361 ( .B1(n14391), .B2(n14343), .A(n14342), .ZN(n14426) );
  MUX2_X1 U16362 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n14426), .S(n15912), .Z(
        P2_U3516) );
  AOI211_X1 U16363 ( .C1(n14346), .C2(n14396), .A(n14345), .B(n14344), .ZN(
        n14427) );
  MUX2_X1 U16364 ( .A(n14347), .B(n14427), .S(n15912), .Z(n14348) );
  OAI21_X1 U16365 ( .B1(n14431), .B2(n14349), .A(n14348), .ZN(P2_U3515) );
  AOI21_X1 U16366 ( .B1(n14387), .B2(n14351), .A(n14350), .ZN(n14352) );
  OAI211_X1 U16367 ( .C1(n14391), .C2(n14354), .A(n14353), .B(n14352), .ZN(
        n14432) );
  MUX2_X1 U16368 ( .A(P2_REG1_REG_15__SCAN_IN), .B(n14432), .S(n15912), .Z(
        P2_U3514) );
  OAI211_X1 U16369 ( .C1(n14391), .C2(n14357), .A(n14356), .B(n14355), .ZN(
        n14433) );
  MUX2_X1 U16370 ( .A(P2_REG1_REG_14__SCAN_IN), .B(n14433), .S(n15912), .Z(
        n14358) );
  AOI21_X1 U16371 ( .B1(n14377), .B2(n14435), .A(n14358), .ZN(n14359) );
  INV_X1 U16372 ( .A(n14359), .ZN(P2_U3513) );
  AOI211_X1 U16373 ( .C1(n14387), .C2(n14362), .A(n14361), .B(n14360), .ZN(
        n14363) );
  OAI21_X1 U16374 ( .B1(n14391), .B2(n14364), .A(n14363), .ZN(n14437) );
  MUX2_X1 U16375 ( .A(P2_REG1_REG_13__SCAN_IN), .B(n14437), .S(n15912), .Z(
        P2_U3512) );
  INV_X1 U16376 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n14371) );
  NAND2_X1 U16377 ( .A1(n14365), .A2(n15905), .ZN(n14367) );
  OAI211_X1 U16378 ( .C1(n14368), .C2(n15900), .A(n14367), .B(n14366), .ZN(
        n14369) );
  NOR2_X1 U16379 ( .A1(n14370), .A2(n14369), .ZN(n14438) );
  MUX2_X1 U16380 ( .A(n14371), .B(n14438), .S(n15912), .Z(n14372) );
  INV_X1 U16381 ( .A(n14372), .ZN(P2_U3511) );
  OAI211_X1 U16382 ( .C1(n14391), .C2(n14375), .A(n14374), .B(n14373), .ZN(
        n14441) );
  MUX2_X1 U16383 ( .A(P2_REG1_REG_11__SCAN_IN), .B(n14441), .S(n15912), .Z(
        n14376) );
  AOI21_X1 U16384 ( .B1(n14377), .B2(n14443), .A(n14376), .ZN(n14378) );
  INV_X1 U16385 ( .A(n14378), .ZN(P2_U3510) );
  NAND2_X1 U16386 ( .A1(n14379), .A2(n14387), .ZN(n14380) );
  OAI211_X1 U16387 ( .C1(n14382), .C2(n14391), .A(n14381), .B(n14380), .ZN(
        n14383) );
  MUX2_X1 U16388 ( .A(n14445), .B(P2_REG1_REG_10__SCAN_IN), .S(n15910), .Z(
        P2_U3509) );
  AOI21_X1 U16389 ( .B1(n14387), .B2(n14386), .A(n14385), .ZN(n14388) );
  OAI211_X1 U16390 ( .C1(n14391), .C2(n14390), .A(n14389), .B(n14388), .ZN(
        n14446) );
  MUX2_X1 U16391 ( .A(n14446), .B(P2_REG1_REG_9__SCAN_IN), .S(n15910), .Z(
        P2_U3508) );
  OAI21_X1 U16392 ( .B1(n14393), .B2(n15900), .A(n14392), .ZN(n14395) );
  AOI211_X1 U16393 ( .C1(n14397), .C2(n14396), .A(n14395), .B(n14394), .ZN(
        n14448) );
  NAND2_X1 U16394 ( .A1(n15910), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n14398) );
  OAI21_X1 U16395 ( .B1(n14448), .B2(n15910), .A(n14398), .ZN(P2_U3507) );
  MUX2_X1 U16396 ( .A(P2_REG0_REG_30__SCAN_IN), .B(n14399), .S(n15908), .Z(
        n14400) );
  AOI21_X1 U16397 ( .B1(n10276), .B2(n14401), .A(n14400), .ZN(n14402) );
  INV_X1 U16398 ( .A(n14402), .ZN(P2_U3497) );
  MUX2_X1 U16399 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n14403), .S(n15908), .Z(
        n14404) );
  INV_X1 U16400 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n14407) );
  MUX2_X1 U16401 ( .A(n14407), .B(n14406), .S(n15908), .Z(n14408) );
  MUX2_X1 U16402 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n14409), .S(n15908), .Z(
        P2_U3492) );
  MUX2_X1 U16403 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n14410), .S(n15908), .Z(
        P2_U3491) );
  INV_X1 U16404 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n14412) );
  MUX2_X1 U16405 ( .A(n14412), .B(n14411), .S(n15908), .Z(n14413) );
  OAI21_X1 U16406 ( .B1(n14414), .B2(n14430), .A(n14413), .ZN(P2_U3490) );
  MUX2_X1 U16407 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n14415), .S(n15908), .Z(
        n14416) );
  AOI21_X1 U16408 ( .B1(n10276), .B2(n14417), .A(n14416), .ZN(n14418) );
  INV_X1 U16409 ( .A(n14418), .ZN(P2_U3489) );
  MUX2_X1 U16410 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n14419), .S(n15908), .Z(
        P2_U3488) );
  MUX2_X1 U16411 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n14420), .S(n15908), .Z(
        P2_U3487) );
  INV_X1 U16412 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n14422) );
  MUX2_X1 U16413 ( .A(n14422), .B(n14421), .S(n15908), .Z(n14423) );
  OAI21_X1 U16414 ( .B1(n14424), .B2(n14430), .A(n14423), .ZN(P2_U3486) );
  MUX2_X1 U16415 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n14425), .S(n15908), .Z(
        P2_U3484) );
  MUX2_X1 U16416 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n14426), .S(n15908), .Z(
        P2_U3481) );
  INV_X1 U16417 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n14428) );
  MUX2_X1 U16418 ( .A(n14428), .B(n14427), .S(n15908), .Z(n14429) );
  OAI21_X1 U16419 ( .B1(n14431), .B2(n14430), .A(n14429), .ZN(P2_U3478) );
  MUX2_X1 U16420 ( .A(P2_REG0_REG_15__SCAN_IN), .B(n14432), .S(n15908), .Z(
        P2_U3475) );
  MUX2_X1 U16421 ( .A(P2_REG0_REG_14__SCAN_IN), .B(n14433), .S(n15908), .Z(
        n14434) );
  AOI21_X1 U16422 ( .B1(n10276), .B2(n14435), .A(n14434), .ZN(n14436) );
  INV_X1 U16423 ( .A(n14436), .ZN(P2_U3472) );
  MUX2_X1 U16424 ( .A(P2_REG0_REG_13__SCAN_IN), .B(n14437), .S(n15908), .Z(
        P2_U3469) );
  INV_X1 U16425 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n14439) );
  MUX2_X1 U16426 ( .A(n14439), .B(n14438), .S(n15908), .Z(n14440) );
  INV_X1 U16427 ( .A(n14440), .ZN(P2_U3466) );
  MUX2_X1 U16428 ( .A(P2_REG0_REG_11__SCAN_IN), .B(n14441), .S(n15908), .Z(
        n14442) );
  AOI21_X1 U16429 ( .B1(n10276), .B2(n14443), .A(n14442), .ZN(n14444) );
  INV_X1 U16430 ( .A(n14444), .ZN(P2_U3463) );
  MUX2_X1 U16431 ( .A(n14445), .B(P2_REG0_REG_10__SCAN_IN), .S(n15906), .Z(
        P2_U3460) );
  MUX2_X1 U16432 ( .A(P2_REG0_REG_9__SCAN_IN), .B(n14446), .S(n15908), .Z(
        P2_U3457) );
  NAND2_X1 U16433 ( .A1(n15906), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n14447) );
  OAI21_X1 U16434 ( .B1(n14448), .B2(n15906), .A(n14447), .ZN(P2_U3454) );
  INV_X1 U16435 ( .A(n14854), .ZN(n15529) );
  INV_X1 U16436 ( .A(n14449), .ZN(n14450) );
  NOR4_X1 U16437 ( .A1(n14450), .A2(P2_IR_REG_30__SCAN_IN), .A3(n14451), .A4(
        P2_U3088), .ZN(n14452) );
  AOI21_X1 U16438 ( .B1(n14458), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n14452), 
        .ZN(n14453) );
  OAI21_X1 U16439 ( .B1(n15529), .B2(n14461), .A(n14453), .ZN(P2_U3296) );
  INV_X1 U16440 ( .A(n14861), .ZN(n15531) );
  OAI222_X1 U16441 ( .A1(n14461), .A2(n15531), .B1(P2_U3088), .B2(n14455), 
        .C1(n14454), .C2(n14472), .ZN(P2_U3298) );
  INV_X1 U16442 ( .A(n14456), .ZN(n15534) );
  AOI21_X1 U16443 ( .B1(n14458), .B2(P1_DATAO_REG_28__SCAN_IN), .A(n14457), 
        .ZN(n14459) );
  OAI21_X1 U16444 ( .B1(n15534), .B2(n14461), .A(n14459), .ZN(P2_U3299) );
  INV_X1 U16445 ( .A(n14460), .ZN(n15537) );
  OAI222_X1 U16446 ( .A1(n14472), .A2(n14463), .B1(P2_U3088), .B2(n14462), 
        .C1(n14461), .C2(n15537), .ZN(P2_U3300) );
  INV_X1 U16447 ( .A(n14464), .ZN(n15541) );
  OAI222_X1 U16448 ( .A1(P2_U3088), .A2(n14466), .B1(n14474), .B2(n15541), 
        .C1(n14465), .C2(n14472), .ZN(P2_U3301) );
  INV_X1 U16449 ( .A(n14467), .ZN(n15544) );
  OAI222_X1 U16450 ( .A1(n14472), .A2(n14470), .B1(n14474), .B2(n15544), .C1(
        P2_U3088), .C2(n14468), .ZN(P2_U3302) );
  INV_X1 U16451 ( .A(n14471), .ZN(n15548) );
  OAI222_X1 U16452 ( .A1(P2_U3088), .A2(n14475), .B1(n14474), .B2(n15548), 
        .C1(n14473), .C2(n14472), .ZN(P2_U3303) );
  MUX2_X1 U16453 ( .A(n14476), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3327) );
  XNOR2_X1 U16454 ( .A(n14478), .B(n14477), .ZN(n14485) );
  OAI21_X1 U16455 ( .B1(n14680), .B2(n14618), .A(n14479), .ZN(n14483) );
  OAI22_X1 U16456 ( .A1(n14481), .A2(n14681), .B1(n15713), .B2(n14480), .ZN(
        n14482) );
  AOI211_X1 U16457 ( .C1(n14684), .C2(n14733), .A(n14483), .B(n14482), .ZN(
        n14484) );
  OAI21_X1 U16458 ( .B1(n14485), .B2(n14686), .A(n14484), .ZN(P1_U3213) );
  XOR2_X1 U16459 ( .A(n14487), .B(n14486), .Z(n14493) );
  OAI21_X1 U16460 ( .B1(n14681), .B2(n14572), .A(n14488), .ZN(n14491) );
  OAI22_X1 U16461 ( .A1(n15310), .A2(n14680), .B1(n15713), .B2(n14489), .ZN(
        n14490) );
  AOI211_X1 U16462 ( .C1(n14772), .C2(n14684), .A(n14491), .B(n14490), .ZN(
        n14492) );
  OAI21_X1 U16463 ( .B1(n14493), .B2(n14686), .A(n14492), .ZN(P1_U3215) );
  OAI21_X1 U16464 ( .B1(n14496), .B2(n14495), .A(n14494), .ZN(n14497) );
  NAND2_X1 U16465 ( .A1(n14497), .A2(n15709), .ZN(n14502) );
  INV_X1 U16466 ( .A(n14498), .ZN(n15195) );
  AOI22_X1 U16467 ( .A1(n15195), .A2(n14639), .B1(P1_REG3_REG_23__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14499) );
  OAI21_X1 U16468 ( .B1(n15402), .B2(n14681), .A(n14499), .ZN(n14500) );
  AOI21_X1 U16469 ( .B1(n14667), .B2(n15384), .A(n14500), .ZN(n14501) );
  OAI211_X1 U16470 ( .C1(n15386), .C2(n14676), .A(n14502), .B(n14501), .ZN(
        P1_U3216) );
  NOR2_X1 U16471 ( .A1(n14650), .A2(n14504), .ZN(n14505) );
  AOI21_X1 U16472 ( .B1(n14650), .B2(n14504), .A(n14505), .ZN(n14614) );
  NAND2_X1 U16473 ( .A1(n14614), .A2(n14615), .ZN(n14613) );
  INV_X1 U16474 ( .A(n14505), .ZN(n14506) );
  NAND2_X1 U16475 ( .A1(n14613), .A2(n14506), .ZN(n14510) );
  INV_X1 U16476 ( .A(n14507), .ZN(n14652) );
  NAND2_X1 U16477 ( .A1(n14652), .A2(n14508), .ZN(n14509) );
  XNOR2_X1 U16478 ( .A(n14510), .B(n14509), .ZN(n14517) );
  OAI22_X1 U16479 ( .A1(n14680), .A2(n14574), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14511), .ZN(n14515) );
  OAI22_X1 U16480 ( .A1(n14513), .A2(n14681), .B1(n15713), .B2(n14512), .ZN(
        n14514) );
  AOI211_X1 U16481 ( .C1(n15495), .C2(n14684), .A(n14515), .B(n14514), .ZN(
        n14516) );
  OAI21_X1 U16482 ( .B1(n14517), .B2(n14686), .A(n14516), .ZN(P1_U3217) );
  AOI22_X1 U16483 ( .A1(n15419), .A2(n14667), .B1(n14639), .B2(n15253), .ZN(
        n14518) );
  NAND2_X1 U16484 ( .A1(P1_U3086), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n15104)
         );
  OAI211_X1 U16485 ( .C1(n15435), .C2(n14681), .A(n14518), .B(n15104), .ZN(
        n14523) );
  INV_X1 U16486 ( .A(n14519), .ZN(n14557) );
  AOI211_X1 U16487 ( .C1(n14521), .C2(n14520), .A(n14686), .B(n14519), .ZN(
        n14522) );
  AOI211_X1 U16488 ( .C1(n14684), .C2(n7226), .A(n14523), .B(n14522), .ZN(
        n14524) );
  INV_X1 U16489 ( .A(n14524), .ZN(P1_U3219) );
  INV_X1 U16490 ( .A(n14541), .ZN(n14534) );
  NAND2_X1 U16491 ( .A1(n15361), .A2(n14525), .ZN(n14528) );
  NAND2_X1 U16492 ( .A1(n15139), .A2(n14526), .ZN(n14527) );
  NAND2_X1 U16493 ( .A1(n14528), .A2(n14527), .ZN(n14530) );
  XNOR2_X1 U16494 ( .A(n14530), .B(n14529), .ZN(n14533) );
  AOI22_X1 U16495 ( .A1(n15361), .A2(n14531), .B1(n14525), .B2(n15139), .ZN(
        n14532) );
  XNOR2_X1 U16496 ( .A(n14533), .B(n14532), .ZN(n14542) );
  AOI22_X1 U16497 ( .A1(n14535), .A2(n14639), .B1(P1_REG3_REG_28__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14537) );
  NAND2_X1 U16498 ( .A1(n14961), .A2(n14667), .ZN(n14536) );
  OAI211_X1 U16499 ( .C1(n14867), .C2(n14681), .A(n14537), .B(n14536), .ZN(
        n14538) );
  AOI21_X1 U16500 ( .B1(n15361), .B2(n14684), .A(n14538), .ZN(n14546) );
  INV_X1 U16501 ( .A(n14543), .ZN(n14540) );
  INV_X1 U16502 ( .A(n14542), .ZN(n14539) );
  NAND4_X1 U16503 ( .A1(n14541), .A2(n15709), .A3(n14540), .A4(n14539), .ZN(
        n14545) );
  NAND3_X1 U16504 ( .A1(n14543), .A2(n15709), .A3(n14542), .ZN(n14544) );
  AOI21_X1 U16505 ( .B1(n14548), .B2(n14547), .A(n6707), .ZN(n14554) );
  AND2_X1 U16506 ( .A1(P1_U3086), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n15024) );
  OAI22_X1 U16507 ( .A1(n14550), .A2(n14681), .B1(n15713), .B2(n14549), .ZN(
        n14551) );
  AOI211_X1 U16508 ( .C1(n14667), .C2(n15800), .A(n15024), .B(n14551), .ZN(
        n14553) );
  NAND2_X1 U16509 ( .A1(n14684), .A2(n14737), .ZN(n14552) );
  OAI211_X1 U16510 ( .C1(n14554), .C2(n14686), .A(n14553), .B(n14552), .ZN(
        P1_U3221) );
  INV_X1 U16511 ( .A(n14555), .ZN(n14556) );
  NAND2_X1 U16512 ( .A1(n14557), .A2(n14556), .ZN(n14625) );
  XNOR2_X1 U16513 ( .A(n14559), .B(n14558), .ZN(n14624) );
  NAND2_X1 U16514 ( .A1(n14625), .A2(n14624), .ZN(n14623) );
  AOI21_X1 U16515 ( .B1(n14623), .B2(n14561), .A(n14560), .ZN(n14564) );
  INV_X1 U16516 ( .A(n14562), .ZN(n14563) );
  OAI21_X1 U16517 ( .B1(n14564), .B2(n14563), .A(n15709), .ZN(n14569) );
  NOR2_X1 U16518 ( .A1(n15227), .A2(n15713), .ZN(n14567) );
  OAI22_X1 U16519 ( .A1(n15401), .A2(n14681), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14565), .ZN(n14566) );
  AOI211_X1 U16520 ( .C1(n14667), .C2(n15383), .A(n14567), .B(n14566), .ZN(
        n14568) );
  OAI211_X1 U16521 ( .C1(n7950), .C2(n14676), .A(n14569), .B(n14568), .ZN(
        P1_U3223) );
  XOR2_X1 U16522 ( .A(n14571), .B(n14570), .Z(n14578) );
  NAND2_X1 U16523 ( .A1(P1_U3086), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n15735)
         );
  OAI21_X1 U16524 ( .B1(n14680), .B2(n14572), .A(n15735), .ZN(n14576) );
  OAI22_X1 U16525 ( .A1(n14574), .A2(n14681), .B1(n15713), .B2(n14573), .ZN(
        n14575) );
  AOI211_X1 U16526 ( .C1(n15480), .C2(n14684), .A(n14576), .B(n14575), .ZN(
        n14577) );
  OAI21_X1 U16527 ( .B1(n14578), .B2(n14686), .A(n14577), .ZN(P1_U3224) );
  XOR2_X1 U16528 ( .A(n14580), .B(n14579), .Z(n14584) );
  OAI22_X1 U16529 ( .A1(n14823), .A2(n15467), .B1(n14812), .B2(n12723), .ZN(
        n15378) );
  INV_X1 U16530 ( .A(n15378), .ZN(n15175) );
  AOI22_X1 U16531 ( .A1(n15174), .A2(n14639), .B1(P1_REG3_REG_25__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14581) );
  OAI21_X1 U16532 ( .B1(n15175), .B2(n14606), .A(n14581), .ZN(n14582) );
  AOI21_X1 U16533 ( .B1(n15379), .B2(n14684), .A(n14582), .ZN(n14583) );
  OAI21_X1 U16534 ( .B1(n14584), .B2(n14686), .A(n14583), .ZN(P1_U3225) );
  XNOR2_X1 U16535 ( .A(n14585), .B(n14586), .ZN(n14679) );
  NOR2_X1 U16536 ( .A1(n14679), .A2(n14678), .ZN(n14677) );
  AOI21_X1 U16537 ( .B1(n14586), .B2(n14585), .A(n14677), .ZN(n14590) );
  XNOR2_X1 U16538 ( .A(n14588), .B(n14587), .ZN(n14589) );
  XNOR2_X1 U16539 ( .A(n14590), .B(n14589), .ZN(n14595) );
  AOI22_X1 U16540 ( .A1(n15315), .A2(n14639), .B1(n14591), .B2(n15458), .ZN(
        n14592) );
  NAND2_X1 U16541 ( .A1(P1_U3086), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n15052)
         );
  OAI211_X1 U16542 ( .C1(n15311), .C2(n14680), .A(n14592), .B(n15052), .ZN(
        n14593) );
  AOI21_X1 U16543 ( .B1(n15444), .B2(n14684), .A(n14593), .ZN(n14594) );
  OAI21_X1 U16544 ( .B1(n14595), .B2(n14686), .A(n14594), .ZN(P1_U3226) );
  XOR2_X1 U16545 ( .A(n14596), .B(n14597), .Z(n14601) );
  NAND2_X1 U16546 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n15063)
         );
  OAI21_X1 U16547 ( .B1(n14681), .B2(n15434), .A(n15063), .ZN(n14599) );
  OAI22_X1 U16548 ( .A1(n15435), .A2(n14680), .B1(n15713), .B2(n15293), .ZN(
        n14598) );
  AOI211_X1 U16549 ( .C1(n15438), .C2(n14684), .A(n14599), .B(n14598), .ZN(
        n14600) );
  OAI21_X1 U16550 ( .B1(n14601), .B2(n14686), .A(n14600), .ZN(P1_U3228) );
  OAI21_X1 U16551 ( .B1(n14604), .B2(n14603), .A(n14602), .ZN(n14605) );
  NAND2_X1 U16552 ( .A1(n14605), .A2(n15709), .ZN(n14612) );
  INV_X1 U16553 ( .A(n14606), .ZN(n15708) );
  INV_X1 U16554 ( .A(n15185), .ZN(n14608) );
  OAI22_X1 U16555 ( .A1(n14608), .A2(n15713), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14607), .ZN(n14609) );
  AOI21_X1 U16556 ( .B1(n14610), .B2(n15708), .A(n14609), .ZN(n14611) );
  OAI211_X1 U16557 ( .C1(n15187), .C2(n14676), .A(n14612), .B(n14611), .ZN(
        P1_U3229) );
  OAI21_X1 U16558 ( .B1(n14615), .B2(n14614), .A(n14613), .ZN(n14616) );
  NAND2_X1 U16559 ( .A1(n14616), .A2(n15709), .ZN(n14622) );
  OAI22_X1 U16560 ( .A1(n14618), .A2(n14681), .B1(n15713), .B2(n14617), .ZN(
        n14619) );
  AOI211_X1 U16561 ( .C1(n14667), .C2(n14966), .A(n14620), .B(n14619), .ZN(
        n14621) );
  OAI211_X1 U16562 ( .C1(n7358), .C2(n14676), .A(n14622), .B(n14621), .ZN(
        P1_U3231) );
  OAI211_X1 U16563 ( .C1(n14625), .C2(n14624), .A(n14623), .B(n15709), .ZN(
        n14630) );
  OAI22_X1 U16564 ( .A1(n15409), .A2(n14681), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14626), .ZN(n14628) );
  NOR2_X1 U16565 ( .A1(n15410), .A2(n14680), .ZN(n14627) );
  AOI211_X1 U16566 ( .C1(n14639), .C2(n15239), .A(n14628), .B(n14627), .ZN(
        n14629) );
  OAI211_X1 U16567 ( .C1(n15236), .C2(n14676), .A(n14630), .B(n14629), .ZN(
        P1_U3233) );
  XOR2_X1 U16568 ( .A(n14632), .B(n14631), .Z(n14638) );
  OAI21_X1 U16569 ( .B1(n14681), .B2(n15466), .A(n14633), .ZN(n14636) );
  OAI22_X1 U16570 ( .A1(n15468), .A2(n14680), .B1(n15713), .B2(n14634), .ZN(
        n14635) );
  AOI211_X1 U16571 ( .C1(n15471), .C2(n14684), .A(n14636), .B(n14635), .ZN(
        n14637) );
  OAI21_X1 U16572 ( .B1(n14638), .B2(n14686), .A(n14637), .ZN(P1_U3234) );
  NAND2_X1 U16573 ( .A1(n15212), .A2(n14667), .ZN(n14641) );
  AOI22_X1 U16574 ( .A1(n15209), .A2(n14639), .B1(P1_REG3_REG_22__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14640) );
  OAI211_X1 U16575 ( .C1(n15410), .C2(n14681), .A(n14641), .B(n14640), .ZN(
        n14646) );
  AOI211_X1 U16576 ( .C1(n14644), .C2(n14643), .A(n14686), .B(n14642), .ZN(
        n14645) );
  AOI211_X1 U16577 ( .C1(n14684), .C2(n15395), .A(n14646), .B(n14645), .ZN(
        n14647) );
  INV_X1 U16578 ( .A(n14647), .ZN(P1_U3235) );
  OAI21_X1 U16579 ( .B1(n14650), .B2(n14649), .A(n14648), .ZN(n14653) );
  AOI21_X1 U16580 ( .B1(n14653), .B2(n14652), .A(n14651), .ZN(n14656) );
  INV_X1 U16581 ( .A(n14654), .ZN(n14655) );
  OAI21_X1 U16582 ( .B1(n14656), .B2(n14655), .A(n15709), .ZN(n14662) );
  NOR2_X1 U16583 ( .A1(n15713), .A2(n14657), .ZN(n14658) );
  AOI211_X1 U16584 ( .C1(n15708), .C2(n14660), .A(n14659), .B(n14658), .ZN(
        n14661) );
  OAI211_X1 U16585 ( .C1(n14753), .C2(n14676), .A(n14662), .B(n14661), .ZN(
        P1_U3236) );
  NAND2_X1 U16586 ( .A1(n15284), .A2(n15701), .ZN(n15429) );
  XNOR2_X1 U16587 ( .A(n14664), .B(n14663), .ZN(n14665) );
  NAND2_X1 U16588 ( .A1(n14665), .A2(n15709), .ZN(n14669) );
  AND2_X1 U16589 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n15070) );
  OAI22_X1 U16590 ( .A1(n15311), .A2(n14681), .B1(n15713), .B2(n15275), .ZN(
        n14666) );
  AOI211_X1 U16591 ( .C1(n14667), .C2(n15428), .A(n15070), .B(n14666), .ZN(
        n14668) );
  OAI211_X1 U16592 ( .C1(n15429), .C2(n15699), .A(n14669), .B(n14668), .ZN(
        P1_U3238) );
  OAI22_X1 U16593 ( .A1(n14867), .A2(n15467), .B1(n14816), .B2(n12723), .ZN(
        n15372) );
  OAI22_X1 U16594 ( .A1(n15160), .A2(n15713), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14673), .ZN(n14674) );
  AOI21_X1 U16595 ( .B1(n15372), .B2(n15708), .A(n14674), .ZN(n14675) );
  AOI21_X1 U16596 ( .B1(n14679), .B2(n14678), .A(n14677), .ZN(n14687) );
  NAND2_X1 U16597 ( .A1(P1_U3086), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n15748)
         );
  OAI21_X1 U16598 ( .B1(n14680), .B2(n15434), .A(n15748), .ZN(n14683) );
  OAI22_X1 U16599 ( .A1(n15468), .A2(n14681), .B1(n15713), .B2(n15330), .ZN(
        n14682) );
  AOI211_X1 U16600 ( .C1(n15325), .C2(n14684), .A(n14683), .B(n14682), .ZN(
        n14685) );
  OAI21_X1 U16601 ( .B1(n14687), .B2(n14686), .A(n14685), .ZN(P1_U3241) );
  XNOR2_X1 U16602 ( .A(n15103), .B(n14688), .ZN(n14691) );
  NAND2_X1 U16603 ( .A1(n14691), .A2(n9194), .ZN(n14848) );
  NAND2_X1 U16604 ( .A1(n14848), .A2(n14689), .ZN(n14833) );
  NAND2_X1 U16605 ( .A1(n14691), .A2(n14690), .ZN(n14692) );
  MUX2_X1 U16606 ( .A(n15168), .B(n15384), .S(n14824), .Z(n14814) );
  INV_X1 U16607 ( .A(n14814), .ZN(n14815) );
  NAND4_X1 U16608 ( .A1(n14694), .A2(n14719), .A3(n14698), .A4(n14693), .ZN(
        n14717) );
  NAND3_X1 U16609 ( .A1(n14695), .A2(n6534), .A3(n14864), .ZN(n14697) );
  NAND3_X1 U16610 ( .A1(n10309), .A2(n14701), .A3(n14719), .ZN(n14696) );
  AND2_X1 U16611 ( .A1(n14697), .A2(n14696), .ZN(n14716) );
  NAND3_X1 U16612 ( .A1(n14698), .A2(n14971), .A3(n14719), .ZN(n14700) );
  NAND2_X1 U16613 ( .A1(n14700), .A2(n14699), .ZN(n14704) );
  NAND2_X1 U16614 ( .A1(n10309), .A2(n14701), .ZN(n14711) );
  NAND3_X1 U16615 ( .A1(n14711), .A2(n14709), .A3(n14864), .ZN(n14702) );
  NAND2_X1 U16616 ( .A1(n14702), .A2(n14708), .ZN(n14703) );
  NAND2_X1 U16617 ( .A1(n14704), .A2(n14703), .ZN(n14715) );
  OAI211_X1 U16618 ( .C1(n14707), .C2(n14706), .A(n6834), .B(n14705), .ZN(
        n14713) );
  OAI211_X1 U16619 ( .C1(n14709), .C2(n14708), .A(n14864), .B(n9141), .ZN(
        n14710) );
  INV_X1 U16620 ( .A(n14710), .ZN(n14712) );
  NAND3_X1 U16621 ( .A1(n14713), .A2(n14712), .A3(n14711), .ZN(n14714) );
  NAND4_X1 U16622 ( .A1(n14717), .A2(n14716), .A3(n14715), .A4(n14714), .ZN(
        n14722) );
  MUX2_X1 U16623 ( .A(n14970), .B(n7945), .S(n14719), .Z(n14718) );
  INV_X1 U16624 ( .A(n14718), .ZN(n14721) );
  MUX2_X1 U16625 ( .A(n14970), .B(n7945), .S(n14864), .Z(n14720) );
  OAI21_X1 U16626 ( .B1(n14722), .B2(n14721), .A(n14720), .ZN(n14724) );
  NAND2_X1 U16627 ( .A1(n14722), .A2(n14721), .ZN(n14723) );
  MUX2_X1 U16628 ( .A(n14725), .B(n14969), .S(n14864), .Z(n14726) );
  MUX2_X1 U16629 ( .A(n14968), .B(n14729), .S(n14719), .Z(n14731) );
  MUX2_X1 U16630 ( .A(n14968), .B(n14729), .S(n14864), .Z(n14730) );
  INV_X1 U16631 ( .A(n14731), .ZN(n14732) );
  MUX2_X1 U16632 ( .A(n15799), .B(n14733), .S(n14864), .Z(n14735) );
  INV_X1 U16633 ( .A(n14735), .ZN(n14736) );
  MUX2_X1 U16634 ( .A(n14967), .B(n14737), .S(n14719), .Z(n14740) );
  MUX2_X1 U16635 ( .A(n14967), .B(n14737), .S(n14824), .Z(n14738) );
  INV_X1 U16636 ( .A(n14740), .ZN(n14741) );
  MUX2_X1 U16637 ( .A(n15800), .B(n14742), .S(n14824), .Z(n14744) );
  MUX2_X1 U16638 ( .A(n15800), .B(n14742), .S(n14719), .Z(n14743) );
  INV_X1 U16639 ( .A(n14744), .ZN(n14745) );
  MUX2_X1 U16640 ( .A(n14966), .B(n15495), .S(n14719), .Z(n14749) );
  NAND2_X1 U16641 ( .A1(n14748), .A2(n14749), .ZN(n14747) );
  MUX2_X1 U16642 ( .A(n14966), .B(n15495), .S(n14824), .Z(n14746) );
  NAND2_X1 U16643 ( .A1(n14747), .A2(n14746), .ZN(n14757) );
  INV_X1 U16644 ( .A(n14748), .ZN(n14751) );
  INV_X1 U16645 ( .A(n14749), .ZN(n14750) );
  NAND2_X1 U16646 ( .A1(n14751), .A2(n14750), .ZN(n14756) );
  MUX2_X1 U16647 ( .A(n15478), .B(n15490), .S(n14824), .Z(n14760) );
  NAND2_X1 U16648 ( .A1(n15478), .A2(n14864), .ZN(n14752) );
  OAI211_X1 U16649 ( .C1(n14753), .C2(n14864), .A(n14760), .B(n14752), .ZN(
        n14754) );
  NAND3_X1 U16650 ( .A1(n14757), .A2(n14756), .A3(n14755), .ZN(n14765) );
  NAND2_X1 U16651 ( .A1(n14771), .A2(n14758), .ZN(n14759) );
  NAND2_X1 U16652 ( .A1(n14759), .A2(n14719), .ZN(n14764) );
  INV_X1 U16653 ( .A(n14760), .ZN(n14762) );
  MUX2_X1 U16654 ( .A(n15478), .B(n15490), .S(n14719), .Z(n14761) );
  NAND3_X1 U16655 ( .A1(n14937), .A2(n14762), .A3(n14761), .ZN(n14763) );
  NAND3_X1 U16656 ( .A1(n14765), .A2(n14764), .A3(n14763), .ZN(n14769) );
  AOI21_X1 U16657 ( .B1(n14768), .B2(n14766), .A(n14719), .ZN(n14767) );
  AOI21_X1 U16658 ( .B1(n14769), .B2(n14768), .A(n14767), .ZN(n14770) );
  MUX2_X1 U16659 ( .A(n15449), .B(n14772), .S(n14824), .Z(n14776) );
  MUX2_X1 U16660 ( .A(n7248), .B(n15468), .S(n14824), .Z(n14775) );
  INV_X1 U16661 ( .A(n15325), .ZN(n15453) );
  MUX2_X1 U16662 ( .A(n15458), .B(n15325), .S(n14719), .Z(n14781) );
  MUX2_X1 U16663 ( .A(n15450), .B(n15444), .S(n14824), .Z(n14785) );
  NOR2_X1 U16664 ( .A1(n15434), .A2(n14719), .ZN(n14773) );
  AOI21_X1 U16665 ( .B1(n15444), .B2(n14719), .A(n14773), .ZN(n14784) );
  AND2_X1 U16666 ( .A1(n14785), .A2(n14784), .ZN(n14774) );
  OAI21_X1 U16667 ( .B1(n14782), .B2(n14781), .A(n14783), .ZN(n14777) );
  MUX2_X1 U16668 ( .A(n14780), .B(n14779), .S(n14824), .Z(n14788) );
  NAND3_X1 U16669 ( .A1(n14783), .A2(n14782), .A3(n14781), .ZN(n14787) );
  INV_X1 U16670 ( .A(n15284), .ZN(n15280) );
  MUX2_X1 U16671 ( .A(n15418), .B(n15284), .S(n14719), .Z(n14789) );
  MUX2_X1 U16672 ( .A(n15401), .B(n15236), .S(n14864), .Z(n14797) );
  MUX2_X1 U16673 ( .A(n15419), .B(n15413), .S(n14719), .Z(n14798) );
  NOR2_X1 U16674 ( .A1(n15252), .A2(n14719), .ZN(n14794) );
  NOR2_X1 U16675 ( .A1(n15421), .A2(n14864), .ZN(n14793) );
  MUX2_X1 U16676 ( .A(n14794), .B(n14793), .S(n15409), .Z(n14795) );
  MUX2_X1 U16677 ( .A(n15410), .B(n7950), .S(n14824), .Z(n14802) );
  NAND2_X1 U16678 ( .A1(n15214), .A2(n15383), .ZN(n14804) );
  MUX2_X1 U16679 ( .A(n14804), .B(n14805), .S(n14864), .Z(n14800) );
  OAI21_X1 U16680 ( .B1(n14803), .B2(n14802), .A(n14800), .ZN(n14808) );
  MUX2_X1 U16681 ( .A(n15240), .B(n15405), .S(n14719), .Z(n14801) );
  AOI21_X1 U16682 ( .B1(n14803), .B2(n14802), .A(n14801), .ZN(n14807) );
  MUX2_X1 U16683 ( .A(n14805), .B(n14804), .S(n14864), .Z(n14806) );
  MUX2_X1 U16684 ( .A(n15392), .B(n15386), .S(n14864), .Z(n14810) );
  MUX2_X1 U16685 ( .A(n15194), .B(n15212), .S(n14864), .Z(n14809) );
  MUX2_X1 U16686 ( .A(n14812), .B(n15187), .S(n14864), .Z(n14813) );
  MUX2_X1 U16687 ( .A(n14964), .B(n15379), .S(n14864), .Z(n14820) );
  INV_X1 U16688 ( .A(n15379), .ZN(n14817) );
  MUX2_X1 U16689 ( .A(n14817), .B(n14816), .S(n14864), .Z(n14818) );
  INV_X1 U16690 ( .A(n14818), .ZN(n14819) );
  INV_X1 U16691 ( .A(n14822), .ZN(n14827) );
  MUX2_X1 U16692 ( .A(n7127), .B(n14823), .S(n14864), .Z(n14826) );
  INV_X1 U16693 ( .A(n14826), .ZN(n14829) );
  MUX2_X1 U16694 ( .A(n14963), .B(n15373), .S(n14824), .Z(n14825) );
  OAI21_X1 U16695 ( .B1(n14822), .B2(n14829), .A(n14828), .ZN(n14884) );
  INV_X1 U16696 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n14832) );
  NAND2_X1 U16697 ( .A1(n14835), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n14831) );
  INV_X1 U16698 ( .A(P1_REG2_REG_31__SCAN_IN), .ZN(n15107) );
  OR2_X1 U16699 ( .A1(n14834), .A2(n15107), .ZN(n14830) );
  OAI211_X1 U16700 ( .C1(n14839), .C2(n14832), .A(n14831), .B(n14830), .ZN(
        n15106) );
  INV_X1 U16701 ( .A(n14833), .ZN(n14840) );
  INV_X1 U16702 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n14838) );
  INV_X1 U16703 ( .A(P1_REG2_REG_30__SCAN_IN), .ZN(n15111) );
  OR2_X1 U16704 ( .A1(n14834), .A2(n15111), .ZN(n14837) );
  NAND2_X1 U16705 ( .A1(n14835), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n14836) );
  OAI211_X1 U16706 ( .C1(n14839), .C2(n14838), .A(n14837), .B(n14836), .ZN(
        n15133) );
  OAI21_X1 U16707 ( .B1(n15106), .B2(n14840), .A(n15133), .ZN(n14841) );
  INV_X1 U16708 ( .A(n14841), .ZN(n14846) );
  NAND2_X1 U16709 ( .A1(n14842), .A2(n8743), .ZN(n14845) );
  OR2_X1 U16710 ( .A1(n8724), .A2(n14843), .ZN(n14844) );
  NAND2_X1 U16711 ( .A1(n15106), .A2(n14719), .ZN(n14858) );
  INV_X1 U16712 ( .A(n15133), .ZN(n14847) );
  AOI21_X1 U16713 ( .B1(n14848), .B2(n14858), .A(n14847), .ZN(n14849) );
  AOI21_X1 U16714 ( .B1(n15114), .B2(n14824), .A(n14849), .ZN(n14895) );
  OR2_X1 U16715 ( .A1(n14894), .A2(n14895), .ZN(n14860) );
  NAND2_X1 U16716 ( .A1(n14850), .A2(n7131), .ZN(n14853) );
  NAND2_X1 U16717 ( .A1(n14851), .A2(n15103), .ZN(n14852) );
  AND2_X1 U16718 ( .A1(n14853), .A2(n14852), .ZN(n14900) );
  NAND2_X1 U16719 ( .A1(n14854), .A2(n8743), .ZN(n14857) );
  INV_X1 U16720 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n14855) );
  OR2_X1 U16721 ( .A1(n8724), .A2(n14855), .ZN(n14856) );
  NAND2_X1 U16722 ( .A1(n14859), .A2(n14858), .ZN(n14901) );
  NAND2_X1 U16723 ( .A1(n14861), .A2(n8743), .ZN(n14863) );
  OR2_X1 U16724 ( .A1(n8724), .A2(n15530), .ZN(n14862) );
  MUX2_X1 U16725 ( .A(n14961), .B(n15350), .S(n14719), .Z(n14872) );
  INV_X1 U16726 ( .A(n14872), .ZN(n14865) );
  MUX2_X1 U16727 ( .A(n14961), .B(n15350), .S(n14864), .Z(n14871) );
  MUX2_X1 U16728 ( .A(n15352), .B(n7942), .S(n14719), .Z(n14875) );
  MUX2_X1 U16729 ( .A(n15139), .B(n15361), .S(n14864), .Z(n14874) );
  AND2_X1 U16730 ( .A1(n14875), .A2(n14874), .ZN(n14888) );
  MUX2_X1 U16731 ( .A(n14867), .B(n14866), .S(n14719), .Z(n14879) );
  MUX2_X1 U16732 ( .A(n14962), .B(n14868), .S(n14824), .Z(n14878) );
  NAND2_X1 U16733 ( .A1(n14879), .A2(n14878), .ZN(n14914) );
  NAND2_X1 U16734 ( .A1(n14894), .A2(n14895), .ZN(n14870) );
  INV_X1 U16735 ( .A(n14900), .ZN(n14896) );
  AND2_X1 U16736 ( .A1(n14899), .A2(n14896), .ZN(n14869) );
  NAND2_X1 U16737 ( .A1(n14870), .A2(n14869), .ZN(n14892) );
  INV_X1 U16738 ( .A(n14871), .ZN(n14873) );
  AND2_X1 U16739 ( .A1(n14873), .A2(n14872), .ZN(n14885) );
  INV_X1 U16740 ( .A(n14874), .ZN(n14877) );
  INV_X1 U16741 ( .A(n14875), .ZN(n14876) );
  AND2_X1 U16742 ( .A1(n14877), .A2(n14876), .ZN(n14890) );
  INV_X1 U16743 ( .A(n14878), .ZN(n14881) );
  INV_X1 U16744 ( .A(n14879), .ZN(n14880) );
  NAND2_X1 U16745 ( .A1(n14881), .A2(n14880), .ZN(n14916) );
  NAND2_X1 U16746 ( .A1(n14913), .A2(n14916), .ZN(n14882) );
  OAI21_X1 U16747 ( .B1(n14884), .B2(n6635), .A(n14883), .ZN(n14955) );
  INV_X1 U16748 ( .A(n14885), .ZN(n14910) );
  INV_X1 U16749 ( .A(n14886), .ZN(n14891) );
  INV_X1 U16750 ( .A(n14887), .ZN(n14889) );
  NOR2_X1 U16751 ( .A1(n14892), .A2(n6611), .ZN(n14907) );
  INV_X1 U16752 ( .A(n14901), .ZN(n14893) );
  AOI21_X1 U16753 ( .B1(n14893), .B2(n14896), .A(n14953), .ZN(n14905) );
  NAND4_X1 U16754 ( .A1(n14901), .A2(n14895), .A3(n14900), .A4(n14894), .ZN(
        n14904) );
  INV_X1 U16755 ( .A(n14894), .ZN(n14898) );
  INV_X1 U16756 ( .A(n14895), .ZN(n14897) );
  NAND4_X1 U16757 ( .A1(n14898), .A2(n14897), .A3(n14896), .A4(n14899), .ZN(
        n14903) );
  INV_X1 U16758 ( .A(n14899), .ZN(n14950) );
  NAND3_X1 U16759 ( .A1(n14901), .A2(n14900), .A3(n14950), .ZN(n14902) );
  NAND4_X1 U16760 ( .A1(n14905), .A2(n14904), .A3(n14903), .A4(n14902), .ZN(
        n14906) );
  NOR2_X1 U16761 ( .A1(n14907), .A2(n14906), .ZN(n14908) );
  OAI211_X1 U16762 ( .C1(n14911), .C2(n14910), .A(n14909), .B(n14908), .ZN(
        n14919) );
  INV_X1 U16763 ( .A(n14912), .ZN(n14917) );
  INV_X1 U16764 ( .A(n14913), .ZN(n14915) );
  OAI22_X1 U16765 ( .A1(n14917), .A2(n14916), .B1(n14915), .B2(n14914), .ZN(
        n14918) );
  NOR2_X1 U16766 ( .A1(n14919), .A2(n14918), .ZN(n14954) );
  INV_X1 U16767 ( .A(n15289), .ZN(n14943) );
  INV_X1 U16768 ( .A(n14920), .ZN(n14930) );
  NOR2_X1 U16769 ( .A1(n14921), .A2(n11373), .ZN(n14925) );
  NAND4_X1 U16770 ( .A1(n14925), .A2(n14924), .A3(n14923), .A4(n14922), .ZN(
        n14927) );
  NOR2_X1 U16771 ( .A1(n14927), .A2(n14926), .ZN(n14929) );
  NAND4_X1 U16772 ( .A1(n14930), .A2(n8770), .A3(n14929), .A4(n14928), .ZN(
        n14931) );
  NOR2_X1 U16773 ( .A1(n14932), .A2(n14931), .ZN(n14936) );
  INV_X1 U16774 ( .A(n14933), .ZN(n14935) );
  AND4_X1 U16775 ( .A1(n14937), .A2(n14936), .A3(n14935), .A4(n14934), .ZN(
        n14938) );
  NAND2_X1 U16776 ( .A1(n14939), .A2(n14938), .ZN(n14940) );
  NOR2_X1 U16777 ( .A1(n14940), .A2(n15308), .ZN(n14942) );
  NAND4_X1 U16778 ( .A1(n15324), .A2(n14943), .A3(n14942), .A4(n14941), .ZN(
        n14944) );
  INV_X1 U16779 ( .A(n15158), .ZN(n15152) );
  NAND4_X1 U16780 ( .A1(n8037), .A2(n15119), .A3(n14947), .A4(n15152), .ZN(
        n14948) );
  INV_X1 U16781 ( .A(n14951), .ZN(n15170) );
  XNOR2_X1 U16782 ( .A(n6665), .B(n15103), .ZN(n14952) );
  NAND3_X1 U16783 ( .A1(n14956), .A2(n15714), .A3(n15798), .ZN(n14957) );
  OAI211_X1 U16784 ( .C1(n15552), .C2(n14959), .A(n14957), .B(P1_B_REG_SCAN_IN), .ZN(n14958) );
  OAI21_X1 U16785 ( .B1(n14960), .B2(n14959), .A(n14958), .ZN(P1_U3242) );
  MUX2_X1 U16786 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(n15106), .S(P1_U4016), .Z(
        P1_U3591) );
  MUX2_X1 U16787 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n15133), .S(P1_U4016), .Z(
        P1_U3590) );
  MUX2_X1 U16788 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n14961), .S(P1_U4016), .Z(
        P1_U3589) );
  MUX2_X1 U16789 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n15139), .S(P1_U4016), .Z(
        P1_U3588) );
  MUX2_X1 U16790 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n14962), .S(P1_U4016), .Z(
        P1_U3587) );
  MUX2_X1 U16791 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n14963), .S(P1_U4016), .Z(
        P1_U3586) );
  MUX2_X1 U16792 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n14964), .S(P1_U4016), .Z(
        P1_U3585) );
  MUX2_X1 U16793 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n15384), .S(P1_U4016), .Z(
        P1_U3584) );
  MUX2_X1 U16794 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n15212), .S(P1_U4016), .Z(
        P1_U3583) );
  MUX2_X1 U16795 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n15383), .S(P1_U4016), .Z(
        P1_U3582) );
  MUX2_X1 U16796 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n15240), .S(P1_U4016), .Z(
        P1_U3581) );
  MUX2_X1 U16797 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n15419), .S(P1_U4016), .Z(
        P1_U3580) );
  MUX2_X1 U16798 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n15428), .S(P1_U4016), .Z(
        P1_U3579) );
  MUX2_X1 U16799 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n15418), .S(P1_U4016), .Z(
        P1_U3578) );
  MUX2_X1 U16800 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n15274), .S(P1_U4016), .Z(
        P1_U3577) );
  MUX2_X1 U16801 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n15450), .S(P1_U4016), .Z(
        P1_U3576) );
  MUX2_X1 U16802 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n15458), .S(P1_U4016), .Z(
        P1_U3575) );
  MUX2_X1 U16803 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n15449), .S(P1_U4016), .Z(
        P1_U3574) );
  MUX2_X1 U16804 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n15479), .S(P1_U4016), .Z(
        P1_U3573) );
  MUX2_X1 U16805 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n14965), .S(P1_U4016), .Z(
        P1_U3572) );
  MUX2_X1 U16806 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n15478), .S(P1_U4016), .Z(
        P1_U3571) );
  MUX2_X1 U16807 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n14966), .S(P1_U4016), .Z(
        P1_U3570) );
  MUX2_X1 U16808 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n15800), .S(P1_U4016), .Z(
        P1_U3569) );
  MUX2_X1 U16809 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n14967), .S(P1_U4016), .Z(
        P1_U3568) );
  MUX2_X1 U16810 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n15799), .S(P1_U4016), .Z(
        P1_U3567) );
  MUX2_X1 U16811 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n14968), .S(P1_U4016), .Z(
        P1_U3566) );
  MUX2_X1 U16812 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n14969), .S(P1_U4016), .Z(
        P1_U3565) );
  MUX2_X1 U16813 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n14970), .S(P1_U4016), .Z(
        P1_U3564) );
  MUX2_X1 U16814 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n10309), .S(P1_U4016), .Z(
        P1_U3563) );
  MUX2_X1 U16815 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n14971), .S(P1_U4016), .Z(
        P1_U3562) );
  MUX2_X1 U16816 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n10855), .S(P1_U4016), .Z(
        P1_U3561) );
  MUX2_X1 U16817 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(n10283), .S(P1_U4016), .Z(
        P1_U3560) );
  NAND2_X1 U16818 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), 
        .ZN(n14974) );
  AOI211_X1 U16819 ( .C1(n14974), .C2(n14973), .A(n14972), .B(n15097), .ZN(
        n14975) );
  INV_X1 U16820 ( .A(n14975), .ZN(n14981) );
  AOI22_X1 U16821 ( .A1(n15722), .A2(P1_ADDR_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(P1_U3086), .ZN(n14980) );
  NAND2_X1 U16822 ( .A1(n15742), .A2(n14976), .ZN(n14979) );
  NAND2_X1 U16823 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n14991) );
  OAI211_X1 U16824 ( .C1(n10754), .C2(n14977), .A(n15746), .B(n14997), .ZN(
        n14978) );
  NAND4_X1 U16825 ( .A1(n14981), .A2(n14980), .A3(n14979), .A4(n14978), .ZN(
        P1_U3244) );
  AOI211_X1 U16826 ( .C1(n14984), .C2(n14983), .A(n14982), .B(n15097), .ZN(
        n14985) );
  INV_X1 U16827 ( .A(n14985), .ZN(n15002) );
  INV_X1 U16828 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n14987) );
  OAI22_X1 U16829 ( .A1(n15750), .A2(n14987), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14986), .ZN(n14988) );
  AOI21_X1 U16830 ( .B1(n14989), .B2(n15742), .A(n14988), .ZN(n15001) );
  MUX2_X1 U16831 ( .A(n14991), .B(n14990), .S(n15536), .Z(n14993) );
  NOR2_X1 U16832 ( .A1(n15536), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n14992) );
  OR2_X1 U16833 ( .A1(n15533), .A2(n14992), .ZN(n15715) );
  NAND2_X1 U16834 ( .A1(n15715), .A2(n15717), .ZN(n15720) );
  OAI211_X1 U16835 ( .C1(n14993), .C2(n15533), .A(P1_U4016), .B(n15720), .ZN(
        n15017) );
  MUX2_X1 U16836 ( .A(P1_REG2_REG_2__SCAN_IN), .B(n11692), .S(n14994), .Z(
        n14996) );
  NAND3_X1 U16837 ( .A1(n14997), .A2(n14996), .A3(n14995), .ZN(n14998) );
  NAND3_X1 U16838 ( .A1(n15746), .A2(n14999), .A3(n14998), .ZN(n15000) );
  NAND4_X1 U16839 ( .A1(n15002), .A2(n15001), .A3(n15017), .A4(n15000), .ZN(
        P1_U3245) );
  AOI211_X1 U16840 ( .C1(n15005), .C2(n15004), .A(n15097), .B(n15003), .ZN(
        n15006) );
  INV_X1 U16841 ( .A(n15006), .ZN(n15019) );
  OAI21_X1 U16842 ( .B1(n15750), .B2(n7501), .A(n15007), .ZN(n15008) );
  AOI21_X1 U16843 ( .B1(n15009), .B2(n15742), .A(n15008), .ZN(n15018) );
  MUX2_X1 U16844 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n10759), .S(n15010), .Z(
        n15011) );
  NAND3_X1 U16845 ( .A1(n15013), .A2(n15012), .A3(n15011), .ZN(n15014) );
  NAND3_X1 U16846 ( .A1(n15746), .A2(n15015), .A3(n15014), .ZN(n15016) );
  NAND4_X1 U16847 ( .A1(n15019), .A2(n15018), .A3(n15017), .A4(n15016), .ZN(
        P1_U3247) );
  OAI21_X1 U16848 ( .B1(n15022), .B2(n15021), .A(n15020), .ZN(n15023) );
  NAND2_X1 U16849 ( .A1(n15023), .A2(n15745), .ZN(n15034) );
  AOI21_X1 U16850 ( .B1(n15722), .B2(P1_ADDR_REG_8__SCAN_IN), .A(n15024), .ZN(
        n15033) );
  MUX2_X1 U16851 ( .A(n11906), .B(P1_REG2_REG_8__SCAN_IN), .S(n15030), .Z(
        n15025) );
  NAND3_X1 U16852 ( .A1(n15027), .A2(n15026), .A3(n15025), .ZN(n15028) );
  NAND3_X1 U16853 ( .A1(n15746), .A2(n15029), .A3(n15028), .ZN(n15032) );
  NAND2_X1 U16854 ( .A1(n15742), .A2(n15030), .ZN(n15031) );
  NAND4_X1 U16855 ( .A1(n15034), .A2(n15033), .A3(n15032), .A4(n15031), .ZN(
        P1_U3251) );
  XNOR2_X1 U16856 ( .A(n15059), .B(P1_REG1_REG_16__SCAN_IN), .ZN(n15040) );
  INV_X1 U16857 ( .A(n15037), .ZN(n15038) );
  NOR2_X1 U16858 ( .A1(n15039), .A2(n15040), .ZN(n15058) );
  AOI211_X1 U16859 ( .C1(n15040), .C2(n15039), .A(n15097), .B(n15058), .ZN(
        n15056) );
  OAI22_X1 U16860 ( .A1(n15044), .A2(n15043), .B1(n15042), .B2(n15041), .ZN(
        n15045) );
  AOI21_X1 U16861 ( .B1(n15743), .B2(n15045), .A(n15046), .ZN(n15740) );
  INV_X1 U16862 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n15739) );
  NAND2_X1 U16863 ( .A1(n15740), .A2(n15739), .ZN(n15738) );
  INV_X1 U16864 ( .A(n15046), .ZN(n15047) );
  NAND2_X1 U16865 ( .A1(n15738), .A2(n15047), .ZN(n15050) );
  INV_X1 U16866 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n15048) );
  MUX2_X1 U16867 ( .A(n15048), .B(P1_REG2_REG_16__SCAN_IN), .S(n15059), .Z(
        n15049) );
  NOR2_X1 U16868 ( .A1(n15050), .A2(n15049), .ZN(n15057) );
  AOI211_X1 U16869 ( .C1(n15050), .C2(n15049), .A(n15099), .B(n15057), .ZN(
        n15055) );
  NAND2_X1 U16870 ( .A1(n15722), .A2(P1_ADDR_REG_16__SCAN_IN), .ZN(n15051) );
  OAI211_X1 U16871 ( .C1(n15068), .C2(n15053), .A(n15052), .B(n15051), .ZN(
        n15054) );
  OR3_X1 U16872 ( .A1(n15056), .A2(n15055), .A3(n15054), .ZN(P1_U3259) );
  AOI21_X1 U16873 ( .B1(n15059), .B2(P1_REG2_REG_16__SCAN_IN), .A(n15057), 
        .ZN(n15071) );
  INV_X1 U16874 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n15075) );
  MUX2_X1 U16875 ( .A(n15075), .B(P1_REG2_REG_17__SCAN_IN), .S(n15078), .Z(
        n15072) );
  XNOR2_X1 U16876 ( .A(n15071), .B(n15072), .ZN(n15067) );
  AOI21_X1 U16877 ( .B1(P1_REG1_REG_16__SCAN_IN), .B2(n15059), .A(n15058), 
        .ZN(n15061) );
  XNOR2_X1 U16878 ( .A(n15078), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n15060) );
  AOI211_X1 U16879 ( .C1(n15061), .C2(n15060), .A(n15097), .B(n15077), .ZN(
        n15062) );
  INV_X1 U16880 ( .A(n15062), .ZN(n15066) );
  OAI21_X1 U16881 ( .B1(n15750), .B2(n15637), .A(n15063), .ZN(n15064) );
  AOI21_X1 U16882 ( .B1(n15078), .B2(n15742), .A(n15064), .ZN(n15065) );
  OAI211_X1 U16883 ( .C1(n15099), .C2(n15067), .A(n15066), .B(n15065), .ZN(
        P1_U3260) );
  NOR2_X1 U16884 ( .A1(n15068), .A2(n15086), .ZN(n15069) );
  AOI211_X1 U16885 ( .C1(n15722), .C2(P1_ADDR_REG_18__SCAN_IN), .A(n15070), 
        .B(n15069), .ZN(n15085) );
  OR2_X1 U16886 ( .A1(n15072), .A2(n15071), .ZN(n15073) );
  OAI21_X1 U16887 ( .B1(n15075), .B2(n15074), .A(n15073), .ZN(n15092) );
  XNOR2_X1 U16888 ( .A(n15086), .B(n15092), .ZN(n15076) );
  NAND2_X1 U16889 ( .A1(P1_REG2_REG_18__SCAN_IN), .A2(n15076), .ZN(n15094) );
  OAI211_X1 U16890 ( .C1(P1_REG2_REG_18__SCAN_IN), .C2(n15076), .A(n15746), 
        .B(n15094), .ZN(n15084) );
  XNOR2_X1 U16891 ( .A(n15086), .B(n15087), .ZN(n15079) );
  INV_X1 U16892 ( .A(n15079), .ZN(n15082) );
  NOR2_X1 U16893 ( .A1(n15080), .A2(n15079), .ZN(n15089) );
  INV_X1 U16894 ( .A(n15089), .ZN(n15081) );
  OAI211_X1 U16895 ( .C1(P1_REG1_REG_18__SCAN_IN), .C2(n15082), .A(n15745), 
        .B(n15081), .ZN(n15083) );
  NAND3_X1 U16896 ( .A1(n15085), .A2(n15084), .A3(n15083), .ZN(P1_U3261) );
  NOR2_X1 U16897 ( .A1(n15087), .A2(n15086), .ZN(n15088) );
  NOR2_X1 U16898 ( .A1(n15089), .A2(n15088), .ZN(n15091) );
  XNOR2_X1 U16899 ( .A(n15091), .B(n15090), .ZN(n15102) );
  NAND2_X1 U16900 ( .A1(n15093), .A2(n15092), .ZN(n15095) );
  NAND2_X1 U16901 ( .A1(n15095), .A2(n15094), .ZN(n15096) );
  XNOR2_X1 U16902 ( .A(P1_REG2_REG_19__SCAN_IN), .B(n15096), .ZN(n15098) );
  INV_X1 U16903 ( .A(n15098), .ZN(n15100) );
  NOR2_X1 U16904 ( .A1(n15100), .A2(n15099), .ZN(n15101) );
  NAND2_X1 U16905 ( .A1(n15130), .A2(n15348), .ZN(n15110) );
  AOI21_X1 U16906 ( .B1(n15714), .B2(P1_B_REG_SCAN_IN), .A(n15467), .ZN(n15134) );
  NAND2_X1 U16907 ( .A1(n15134), .A2(n15106), .ZN(n15346) );
  NOR2_X1 U16908 ( .A1(n15286), .A2(n15346), .ZN(n15113) );
  NOR2_X1 U16909 ( .A1(n15312), .A2(n15107), .ZN(n15108) );
  AOI211_X1 U16910 ( .C1(n15344), .C2(n15291), .A(n15113), .B(n15108), .ZN(
        n15109) );
  OAI21_X1 U16911 ( .B1(n15345), .B2(n15281), .A(n15109), .ZN(P1_U3263) );
  OAI211_X1 U16912 ( .C1(n15130), .C2(n15348), .A(n15447), .B(n15110), .ZN(
        n15347) );
  NOR2_X1 U16913 ( .A1(n15312), .A2(n15111), .ZN(n15112) );
  AOI211_X1 U16914 ( .C1(n15114), .C2(n15291), .A(n15113), .B(n15112), .ZN(
        n15115) );
  OAI21_X1 U16915 ( .B1(n15347), .B2(n15281), .A(n15115), .ZN(P1_U3264) );
  AND2_X1 U16916 ( .A1(n15361), .A2(n15139), .ZN(n15116) );
  INV_X1 U16917 ( .A(n15116), .ZN(n15121) );
  INV_X1 U16918 ( .A(n15117), .ZN(n15118) );
  AOI21_X1 U16919 ( .B1(n15125), .B2(n15121), .A(n15144), .ZN(n15120) );
  AOI21_X1 U16920 ( .B1(n15144), .B2(n15121), .A(n15120), .ZN(n15122) );
  INV_X1 U16921 ( .A(n15144), .ZN(n15126) );
  NOR2_X1 U16922 ( .A1(n15126), .A2(n15125), .ZN(n15127) );
  AOI211_X1 U16923 ( .C1(n15350), .C2(n15131), .A(n7130), .B(n15130), .ZN(
        n15354) );
  NOR2_X1 U16924 ( .A1(n15132), .A2(n15294), .ZN(n15138) );
  NAND2_X1 U16925 ( .A1(n15134), .A2(n15133), .ZN(n15351) );
  OAI22_X1 U16926 ( .A1(n15312), .A2(n15136), .B1(n15351), .B2(n15135), .ZN(
        n15137) );
  AOI211_X1 U16927 ( .C1(n15139), .C2(n15336), .A(n15138), .B(n15137), .ZN(
        n15140) );
  OAI21_X1 U16928 ( .B1(n7941), .B2(n15339), .A(n15140), .ZN(n15141) );
  AOI21_X1 U16929 ( .B1(n15354), .B2(n15319), .A(n15141), .ZN(n15147) );
  NAND2_X1 U16930 ( .A1(n15349), .A2(n15341), .ZN(n15146) );
  OAI211_X1 U16931 ( .C1(n8031), .C2(n15343), .A(n15147), .B(n15146), .ZN(
        P1_U3356) );
  INV_X1 U16932 ( .A(n15148), .ZN(n15149) );
  AOI21_X1 U16933 ( .B1(n12728), .B2(n15150), .A(n15149), .ZN(n15169) );
  NAND2_X1 U16934 ( .A1(n15152), .A2(n15151), .ZN(n15154) );
  OAI21_X1 U16935 ( .B1(n15169), .B2(n15154), .A(n15153), .ZN(n15376) );
  AOI21_X1 U16936 ( .B1(n15158), .B2(n15157), .A(n15156), .ZN(n15370) );
  NAND2_X1 U16937 ( .A1(n15370), .A2(n15341), .ZN(n15165) );
  AOI211_X1 U16938 ( .C1(n15373), .C2(n15172), .A(n7130), .B(n15159), .ZN(
        n15371) );
  OAI22_X1 U16939 ( .A1(n15160), .A2(n15294), .B1(n9284), .B2(n15312), .ZN(
        n15161) );
  AOI21_X1 U16940 ( .B1(n15372), .B2(n15312), .A(n15161), .ZN(n15162) );
  OAI21_X1 U16941 ( .B1(n7127), .B2(n15339), .A(n15162), .ZN(n15163) );
  AOI21_X1 U16942 ( .B1(n15371), .B2(n15319), .A(n15163), .ZN(n15164) );
  OAI211_X1 U16943 ( .C1(n15376), .C2(n15343), .A(n15165), .B(n15164), .ZN(
        P1_U3267) );
  XNOR2_X1 U16944 ( .A(n15166), .B(n15170), .ZN(n15382) );
  AOI211_X1 U16945 ( .C1(n15379), .C2(n15173), .A(n7130), .B(n7128), .ZN(
        n15377) );
  INV_X1 U16946 ( .A(n15174), .ZN(n15176) );
  OAI21_X1 U16947 ( .B1(n15176), .B2(n15294), .A(n15175), .ZN(n15177) );
  AOI21_X1 U16948 ( .B1(n15377), .B2(n15178), .A(n15177), .ZN(n15180) );
  AOI22_X1 U16949 ( .A1(n15379), .A2(n15291), .B1(n15286), .B2(
        P1_REG2_REG_25__SCAN_IN), .ZN(n15179) );
  OAI21_X1 U16950 ( .B1(n15180), .B2(n15286), .A(n15179), .ZN(n15181) );
  AOI21_X1 U16951 ( .B1(n15380), .B2(n15290), .A(n15181), .ZN(n15182) );
  OAI21_X1 U16952 ( .B1(n15301), .B2(n15382), .A(n15182), .ZN(P1_U3268) );
  NOR2_X1 U16953 ( .A1(n15184), .A2(n15281), .ZN(n15189) );
  AOI22_X1 U16954 ( .A1(n15185), .A2(n15331), .B1(P1_REG2_REG_24__SCAN_IN), 
        .B2(n15286), .ZN(n15186) );
  OAI21_X1 U16955 ( .B1(n15187), .B2(n15339), .A(n15186), .ZN(n15188) );
  AOI211_X1 U16956 ( .C1(n15183), .C2(n15312), .A(n15189), .B(n15188), .ZN(
        n15190) );
  INV_X1 U16957 ( .A(n15190), .ZN(P1_U3269) );
  XNOR2_X1 U16958 ( .A(n15192), .B(n15191), .ZN(n15193) );
  NAND2_X1 U16959 ( .A1(n15193), .A2(n15807), .ZN(n15389) );
  XNOR2_X1 U16960 ( .A(n15208), .B(n15194), .ZN(n15388) );
  AOI22_X1 U16961 ( .A1(n15195), .A2(n15331), .B1(P1_REG2_REG_23__SCAN_IN), 
        .B2(n15286), .ZN(n15196) );
  OAI21_X1 U16962 ( .B1(n15402), .B2(n15255), .A(n15196), .ZN(n15197) );
  AOI21_X1 U16963 ( .B1(n15257), .B2(n15384), .A(n15197), .ZN(n15198) );
  OAI21_X1 U16964 ( .B1(n15386), .B2(n15339), .A(n15198), .ZN(n15203) );
  INV_X1 U16965 ( .A(n12728), .ZN(n15201) );
  OAI21_X1 U16966 ( .B1(n15201), .B2(n15200), .A(n15199), .ZN(n15391) );
  NOR2_X1 U16967 ( .A1(n15391), .A2(n15343), .ZN(n15202) );
  AOI211_X1 U16968 ( .C1(n15388), .C2(n15329), .A(n15203), .B(n15202), .ZN(
        n15204) );
  OAI21_X1 U16969 ( .B1(n15286), .B2(n15389), .A(n15204), .ZN(P1_U3270) );
  INV_X1 U16970 ( .A(n15205), .ZN(n15206) );
  AOI21_X1 U16971 ( .B1(n15217), .B2(n15207), .A(n15206), .ZN(n15399) );
  AOI211_X1 U16972 ( .C1(n15395), .C2(n15225), .A(n7130), .B(n15208), .ZN(
        n15393) );
  AOI22_X1 U16973 ( .A1(n15209), .A2(n15331), .B1(P1_REG2_REG_22__SCAN_IN), 
        .B2(n15286), .ZN(n15210) );
  OAI21_X1 U16974 ( .B1(n15410), .B2(n15255), .A(n15210), .ZN(n15211) );
  AOI21_X1 U16975 ( .B1(n15257), .B2(n15212), .A(n15211), .ZN(n15213) );
  OAI21_X1 U16976 ( .B1(n15214), .B2(n15339), .A(n15213), .ZN(n15215) );
  AOI21_X1 U16977 ( .B1(n15393), .B2(n15319), .A(n15215), .ZN(n15219) );
  XNOR2_X1 U16978 ( .A(n15216), .B(n15217), .ZN(n15396) );
  NAND2_X1 U16979 ( .A1(n15396), .A2(n15290), .ZN(n15218) );
  OAI211_X1 U16980 ( .C1(n15399), .C2(n15301), .A(n15219), .B(n15218), .ZN(
        P1_U3271) );
  OAI21_X1 U16981 ( .B1(n15220), .B2(n15222), .A(n15221), .ZN(n15408) );
  OAI21_X1 U16982 ( .B1(n15224), .B2(n9171), .A(n15223), .ZN(n15400) );
  NAND2_X1 U16983 ( .A1(n15400), .A2(n15290), .ZN(n15234) );
  AOI21_X1 U16984 ( .B1(n15238), .B2(n15405), .A(n7130), .ZN(n15226) );
  AND2_X1 U16985 ( .A1(n15226), .A2(n15225), .ZN(n15403) );
  INV_X1 U16986 ( .A(n15227), .ZN(n15228) );
  AOI22_X1 U16987 ( .A1(n15228), .A2(n15331), .B1(P1_REG2_REG_21__SCAN_IN), 
        .B2(n15286), .ZN(n15229) );
  OAI21_X1 U16988 ( .B1(n15401), .B2(n15255), .A(n15229), .ZN(n15230) );
  AOI21_X1 U16989 ( .B1(n15257), .B2(n15383), .A(n15230), .ZN(n15231) );
  OAI21_X1 U16990 ( .B1(n7950), .B2(n15339), .A(n15231), .ZN(n15232) );
  AOI21_X1 U16991 ( .B1(n15403), .B2(n15319), .A(n15232), .ZN(n15233) );
  OAI211_X1 U16992 ( .C1(n15408), .C2(n15301), .A(n15234), .B(n15233), .ZN(
        P1_U3272) );
  OAI21_X1 U16993 ( .B1(n6679), .B2(n7703), .A(n15235), .ZN(n15417) );
  OR2_X1 U16994 ( .A1(n15251), .A2(n15236), .ZN(n15237) );
  AND3_X1 U16995 ( .A1(n15238), .A2(n15237), .A3(n15447), .ZN(n15411) );
  NAND2_X1 U16996 ( .A1(n15413), .A2(n15291), .ZN(n15244) );
  AOI22_X1 U16997 ( .A1(n15239), .A2(n15331), .B1(P1_REG2_REG_20__SCAN_IN), 
        .B2(n15286), .ZN(n15243) );
  NAND2_X1 U16998 ( .A1(n15240), .A2(n15257), .ZN(n15242) );
  NAND2_X1 U16999 ( .A1(n15428), .A2(n15336), .ZN(n15241) );
  NAND4_X1 U17000 ( .A1(n15244), .A2(n15243), .A3(n15242), .A4(n15241), .ZN(
        n15245) );
  AOI21_X1 U17001 ( .B1(n15411), .B2(n15319), .A(n15245), .ZN(n15249) );
  NAND2_X1 U17002 ( .A1(n7336), .A2(n7703), .ZN(n15414) );
  NAND3_X1 U17003 ( .A1(n15246), .A2(n15414), .A3(n15290), .ZN(n15248) );
  OAI211_X1 U17004 ( .C1(n15417), .C2(n15301), .A(n15249), .B(n15248), .ZN(
        P1_U3273) );
  XOR2_X1 U17005 ( .A(n15262), .B(n15250), .Z(n15427) );
  INV_X1 U17006 ( .A(n8033), .ZN(n15279) );
  AOI21_X1 U17007 ( .B1(n7226), .B2(n15279), .A(n15251), .ZN(n15425) );
  AOI22_X1 U17008 ( .A1(n15253), .A2(n15331), .B1(n15286), .B2(
        P1_REG2_REG_19__SCAN_IN), .ZN(n15254) );
  OAI21_X1 U17009 ( .B1(n15255), .B2(n15435), .A(n15254), .ZN(n15256) );
  AOI21_X1 U17010 ( .B1(n15257), .B2(n15419), .A(n15256), .ZN(n15258) );
  OAI21_X1 U17011 ( .B1(n15421), .B2(n15339), .A(n15258), .ZN(n15264) );
  INV_X1 U17012 ( .A(n15259), .ZN(n15260) );
  AOI21_X1 U17013 ( .B1(n15262), .B2(n15261), .A(n15260), .ZN(n15422) );
  NOR2_X1 U17014 ( .A1(n15422), .A2(n15301), .ZN(n15263) );
  AOI211_X1 U17015 ( .C1(n15425), .C2(n15329), .A(n15264), .B(n15263), .ZN(
        n15265) );
  OAI21_X1 U17016 ( .B1(n15343), .B2(n15427), .A(n15265), .ZN(P1_U3274) );
  XOR2_X1 U17017 ( .A(n15266), .B(n15271), .Z(n15267) );
  NOR2_X1 U17018 ( .A1(n15267), .A2(n15492), .ZN(n15273) );
  INV_X1 U17019 ( .A(n15268), .ZN(n15269) );
  AOI211_X1 U17020 ( .C1(n15271), .C2(n15270), .A(n15465), .B(n15269), .ZN(
        n15272) );
  INV_X1 U17021 ( .A(n15275), .ZN(n15276) );
  AOI22_X1 U17022 ( .A1(n15286), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n15276), 
        .B2(n15331), .ZN(n15277) );
  OAI21_X1 U17023 ( .B1(n15334), .B2(n15409), .A(n15277), .ZN(n15283) );
  OAI211_X1 U17024 ( .C1(n15280), .C2(n15278), .A(n15279), .B(n15447), .ZN(
        n15430) );
  NOR2_X1 U17025 ( .A1(n15430), .A2(n15281), .ZN(n15282) );
  AOI211_X1 U17026 ( .C1(n15291), .C2(n15284), .A(n15283), .B(n15282), .ZN(
        n15285) );
  OAI21_X1 U17027 ( .B1(n15432), .B2(n15286), .A(n15285), .ZN(P1_U3275) );
  XNOR2_X1 U17028 ( .A(n15289), .B(n15287), .ZN(n15441) );
  XNOR2_X1 U17029 ( .A(n15289), .B(n15288), .ZN(n15433) );
  NAND2_X1 U17030 ( .A1(n15433), .A2(n15290), .ZN(n15300) );
  AOI211_X1 U17031 ( .C1(n15438), .C2(n15313), .A(n7130), .B(n15278), .ZN(
        n15436) );
  NAND2_X1 U17032 ( .A1(n15438), .A2(n15291), .ZN(n15297) );
  NAND2_X1 U17033 ( .A1(n15286), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n15292) );
  OAI21_X1 U17034 ( .B1(n15294), .B2(n15293), .A(n15292), .ZN(n15295) );
  AOI21_X1 U17035 ( .B1(n15336), .B2(n15450), .A(n15295), .ZN(n15296) );
  OAI211_X1 U17036 ( .C1(n15435), .C2(n15334), .A(n15297), .B(n15296), .ZN(
        n15298) );
  AOI21_X1 U17037 ( .B1(n15436), .B2(n15319), .A(n15298), .ZN(n15299) );
  OAI211_X1 U17038 ( .C1(n15441), .C2(n15301), .A(n15300), .B(n15299), .ZN(
        P1_U3276) );
  OAI21_X1 U17039 ( .B1(n15302), .B2(n15308), .A(n15303), .ZN(n15304) );
  INV_X1 U17040 ( .A(n15304), .ZN(n15446) );
  INV_X1 U17041 ( .A(n15305), .ZN(n15306) );
  AOI21_X1 U17042 ( .B1(n15308), .B2(n15307), .A(n15306), .ZN(n15309) );
  OAI222_X1 U17043 ( .A1(n15467), .A2(n15311), .B1(n12723), .B2(n15310), .C1(
        n15309), .C2(n15465), .ZN(n15442) );
  NAND2_X1 U17044 ( .A1(n15442), .A2(n15312), .ZN(n15321) );
  INV_X1 U17045 ( .A(n15328), .ZN(n15314) );
  AOI211_X1 U17046 ( .C1(n15444), .C2(n15314), .A(n7130), .B(n6531), .ZN(
        n15443) );
  AOI22_X1 U17047 ( .A1(n15286), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n15315), 
        .B2(n15331), .ZN(n15316) );
  OAI21_X1 U17048 ( .B1(n15317), .B2(n15339), .A(n15316), .ZN(n15318) );
  AOI21_X1 U17049 ( .B1(n15443), .B2(n15319), .A(n15318), .ZN(n15320) );
  OAI211_X1 U17050 ( .C1(n15446), .C2(n15343), .A(n15321), .B(n15320), .ZN(
        P1_U3277) );
  XOR2_X1 U17051 ( .A(n15322), .B(n15324), .Z(n15457) );
  XOR2_X1 U17052 ( .A(n15323), .B(n15324), .Z(n15455) );
  AND2_X1 U17053 ( .A1(n15326), .A2(n15325), .ZN(n15327) );
  NOR2_X1 U17054 ( .A1(n15328), .A2(n15327), .ZN(n15448) );
  NAND2_X1 U17055 ( .A1(n15448), .A2(n15329), .ZN(n15338) );
  INV_X1 U17056 ( .A(n15330), .ZN(n15332) );
  AOI22_X1 U17057 ( .A1(n15286), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n15332), 
        .B2(n15331), .ZN(n15333) );
  OAI21_X1 U17058 ( .B1(n15334), .B2(n15434), .A(n15333), .ZN(n15335) );
  AOI21_X1 U17059 ( .B1(n15336), .B2(n15449), .A(n15335), .ZN(n15337) );
  OAI211_X1 U17060 ( .C1(n15453), .C2(n15339), .A(n15338), .B(n15337), .ZN(
        n15340) );
  AOI21_X1 U17061 ( .B1(n15455), .B2(n15341), .A(n15340), .ZN(n15342) );
  OAI21_X1 U17062 ( .B1(n15457), .B2(n15343), .A(n15342), .ZN(P1_U3278) );
  MUX2_X1 U17063 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n15503), .S(n15822), .Z(
        P1_U3559) );
  OAI211_X1 U17064 ( .C1(n15804), .C2(n15348), .A(n15347), .B(n15346), .ZN(
        n15504) );
  MUX2_X1 U17065 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n15504), .S(n15822), .Z(
        P1_U3558) );
  NAND2_X1 U17066 ( .A1(n15349), .A2(n15807), .ZN(n15358) );
  OAI21_X1 U17067 ( .B1(n15352), .B2(n12723), .A(n15351), .ZN(n15353) );
  INV_X1 U17068 ( .A(n15353), .ZN(n15356) );
  INV_X1 U17069 ( .A(n15354), .ZN(n15355) );
  MUX2_X1 U17070 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n15505), .S(n15822), .Z(
        P1_U3557) );
  NAND2_X1 U17071 ( .A1(n15361), .A2(n15701), .ZN(n15362) );
  NAND2_X1 U17072 ( .A1(n15369), .A2(n8042), .ZN(n15507) );
  MUX2_X1 U17073 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n15507), .S(n15822), .Z(
        P1_U3555) );
  NAND2_X1 U17074 ( .A1(n15370), .A2(n15807), .ZN(n15375) );
  AOI211_X1 U17075 ( .C1(n15373), .C2(n15701), .A(n15372), .B(n15371), .ZN(
        n15374) );
  OAI211_X1 U17076 ( .C1(n15492), .C2(n15376), .A(n15375), .B(n15374), .ZN(
        n15508) );
  MUX2_X1 U17077 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n15508), .S(n15822), .Z(
        P1_U3554) );
  AOI211_X1 U17078 ( .C1(n15379), .C2(n15701), .A(n15378), .B(n15377), .ZN(
        n15381) );
  MUX2_X1 U17079 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n15509), .S(n15822), .Z(
        P1_U3553) );
  AOI22_X1 U17080 ( .A1(n15384), .A2(n15801), .B1(n15798), .B2(n15383), .ZN(
        n15385) );
  OAI21_X1 U17081 ( .B1(n15386), .B2(n15804), .A(n15385), .ZN(n15387) );
  AOI21_X1 U17082 ( .B1(n15388), .B2(n15447), .A(n15387), .ZN(n15390) );
  OAI211_X1 U17083 ( .C1(n15391), .C2(n15492), .A(n15390), .B(n15389), .ZN(
        n15510) );
  MUX2_X1 U17084 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n15510), .S(n15822), .Z(
        P1_U3551) );
  OAI22_X1 U17085 ( .A1(n15392), .A2(n15467), .B1(n15410), .B2(n12723), .ZN(
        n15394) );
  AOI211_X1 U17086 ( .C1(n15395), .C2(n15701), .A(n15394), .B(n15393), .ZN(
        n15398) );
  NAND2_X1 U17087 ( .A1(n15396), .A2(n15812), .ZN(n15397) );
  OAI211_X1 U17088 ( .C1(n15399), .C2(n15465), .A(n15398), .B(n15397), .ZN(
        n15511) );
  MUX2_X1 U17089 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n15511), .S(n15822), .Z(
        P1_U3550) );
  NAND2_X1 U17090 ( .A1(n15400), .A2(n15812), .ZN(n15407) );
  OAI22_X1 U17091 ( .A1(n15402), .A2(n15467), .B1(n15401), .B2(n12723), .ZN(
        n15404) );
  AOI211_X1 U17092 ( .C1(n15405), .C2(n15701), .A(n15404), .B(n15403), .ZN(
        n15406) );
  OAI211_X1 U17093 ( .C1(n15465), .C2(n15408), .A(n15407), .B(n15406), .ZN(
        n15512) );
  MUX2_X1 U17094 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n15512), .S(n15822), .Z(
        P1_U3549) );
  OAI22_X1 U17095 ( .A1(n15410), .A2(n15467), .B1(n15409), .B2(n12723), .ZN(
        n15412) );
  AOI211_X1 U17096 ( .C1(n15413), .C2(n15701), .A(n15412), .B(n15411), .ZN(
        n15416) );
  NAND3_X1 U17097 ( .A1(n15246), .A2(n15414), .A3(n15812), .ZN(n15415) );
  OAI211_X1 U17098 ( .C1(n15417), .C2(n15465), .A(n15416), .B(n15415), .ZN(
        n15513) );
  MUX2_X1 U17099 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n15513), .S(n15822), .Z(
        P1_U3548) );
  AOI22_X1 U17100 ( .A1(n15419), .A2(n15801), .B1(n15798), .B2(n15418), .ZN(
        n15420) );
  OAI21_X1 U17101 ( .B1(n15421), .B2(n15804), .A(n15420), .ZN(n15424) );
  NOR2_X1 U17102 ( .A1(n15422), .A2(n15465), .ZN(n15423) );
  AOI211_X1 U17103 ( .C1(n15447), .C2(n15425), .A(n15424), .B(n15423), .ZN(
        n15426) );
  OAI21_X1 U17104 ( .B1(n15492), .B2(n15427), .A(n15426), .ZN(n15514) );
  MUX2_X1 U17105 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n15514), .S(n15822), .Z(
        P1_U3547) );
  NAND2_X1 U17106 ( .A1(n15428), .A2(n15801), .ZN(n15431) );
  NAND4_X1 U17107 ( .A1(n15432), .A2(n15431), .A3(n15430), .A4(n15429), .ZN(
        n15515) );
  MUX2_X1 U17108 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n15515), .S(n15822), .Z(
        P1_U3546) );
  NAND2_X1 U17109 ( .A1(n15433), .A2(n15812), .ZN(n15440) );
  OAI22_X1 U17110 ( .A1(n15435), .A2(n15467), .B1(n15434), .B2(n12723), .ZN(
        n15437) );
  AOI211_X1 U17111 ( .C1(n15438), .C2(n15701), .A(n15437), .B(n15436), .ZN(
        n15439) );
  OAI211_X1 U17112 ( .C1(n15465), .C2(n15441), .A(n15440), .B(n15439), .ZN(
        n15516) );
  MUX2_X1 U17113 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n15516), .S(n15822), .Z(
        P1_U3545) );
  AOI211_X1 U17114 ( .C1(n15444), .C2(n15701), .A(n15443), .B(n15442), .ZN(
        n15445) );
  OAI21_X1 U17115 ( .B1(n15446), .B2(n15492), .A(n15445), .ZN(n15517) );
  MUX2_X1 U17116 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n15517), .S(n15822), .Z(
        P1_U3544) );
  NAND2_X1 U17117 ( .A1(n15448), .A2(n15447), .ZN(n15452) );
  AOI22_X1 U17118 ( .A1(n15450), .A2(n15801), .B1(n15798), .B2(n15449), .ZN(
        n15451) );
  OAI211_X1 U17119 ( .C1(n15453), .C2(n15804), .A(n15452), .B(n15451), .ZN(
        n15454) );
  AOI21_X1 U17120 ( .B1(n15455), .B2(n15807), .A(n15454), .ZN(n15456) );
  OAI21_X1 U17121 ( .B1(n15457), .B2(n15492), .A(n15456), .ZN(n15518) );
  MUX2_X1 U17122 ( .A(P1_REG1_REG_15__SCAN_IN), .B(n15518), .S(n15822), .Z(
        P1_U3543) );
  AOI22_X1 U17123 ( .A1(n15479), .A2(n15798), .B1(n15801), .B2(n15458), .ZN(
        n15459) );
  OAI211_X1 U17124 ( .C1(n7248), .C2(n15804), .A(n15460), .B(n15459), .ZN(
        n15461) );
  AOI21_X1 U17125 ( .B1(n15462), .B2(n15812), .A(n15461), .ZN(n15463) );
  OAI21_X1 U17126 ( .B1(n15465), .B2(n15464), .A(n15463), .ZN(n15519) );
  MUX2_X1 U17127 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n15519), .S(n15822), .Z(
        P1_U3542) );
  OAI22_X1 U17128 ( .A1(n15468), .A2(n15467), .B1(n15466), .B2(n12723), .ZN(
        n15469) );
  AOI21_X1 U17129 ( .B1(n15471), .B2(n15470), .A(n15469), .ZN(n15472) );
  OAI211_X1 U17130 ( .C1(n7130), .C2(n15474), .A(n15473), .B(n15472), .ZN(
        n15475) );
  AOI21_X1 U17131 ( .B1(n15812), .B2(n15476), .A(n15475), .ZN(n15477) );
  INV_X1 U17132 ( .A(n15477), .ZN(n15520) );
  MUX2_X1 U17133 ( .A(P1_REG1_REG_13__SCAN_IN), .B(n15520), .S(n15822), .Z(
        P1_U3541) );
  AOI22_X1 U17134 ( .A1(n15479), .A2(n15801), .B1(n15798), .B2(n15478), .ZN(
        n15483) );
  NAND2_X1 U17135 ( .A1(n15480), .A2(n15701), .ZN(n15481) );
  NAND4_X1 U17136 ( .A1(n15484), .A2(n15483), .A3(n15482), .A4(n15481), .ZN(
        n15485) );
  AOI21_X1 U17137 ( .B1(n15812), .B2(n15486), .A(n15485), .ZN(n15487) );
  INV_X1 U17138 ( .A(n15487), .ZN(n15521) );
  MUX2_X1 U17139 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n15521), .S(n15822), .Z(
        P1_U3540) );
  AOI211_X1 U17140 ( .C1(n15490), .C2(n15701), .A(n15489), .B(n15488), .ZN(
        n15491) );
  OAI21_X1 U17141 ( .B1(n15493), .B2(n15492), .A(n15491), .ZN(n15522) );
  MUX2_X1 U17142 ( .A(P1_REG1_REG_11__SCAN_IN), .B(n15522), .S(n15822), .Z(
        P1_U3539) );
  NAND2_X1 U17143 ( .A1(n15494), .A2(n15812), .ZN(n15501) );
  AOI22_X1 U17144 ( .A1(n15495), .A2(n15701), .B1(n15798), .B2(n15800), .ZN(
        n15499) );
  NAND3_X1 U17145 ( .A1(n15497), .A2(n15496), .A3(n15807), .ZN(n15498) );
  NAND4_X1 U17146 ( .A1(n15501), .A2(n15500), .A3(n15499), .A4(n15498), .ZN(
        n15523) );
  MUX2_X1 U17147 ( .A(n15523), .B(P1_REG1_REG_10__SCAN_IN), .S(n15820), .Z(
        P1_U3538) );
  MUX2_X1 U17148 ( .A(P1_REG1_REG_0__SCAN_IN), .B(n15502), .S(n15822), .Z(
        P1_U3528) );
  MUX2_X1 U17149 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n15504), .S(n15815), .Z(
        P1_U3526) );
  MUX2_X1 U17150 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n15505), .S(n15815), .Z(
        P1_U3525) );
  MUX2_X1 U17151 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n15507), .S(n15815), .Z(
        P1_U3523) );
  MUX2_X1 U17152 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n15508), .S(n15815), .Z(
        P1_U3522) );
  MUX2_X1 U17153 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n15509), .S(n15815), .Z(
        P1_U3521) );
  MUX2_X1 U17154 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n15510), .S(n15815), .Z(
        P1_U3519) );
  MUX2_X1 U17155 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n15511), .S(n15815), .Z(
        P1_U3518) );
  MUX2_X1 U17156 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n15512), .S(n15815), .Z(
        P1_U3517) );
  MUX2_X1 U17157 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n15513), .S(n15815), .Z(
        P1_U3516) );
  MUX2_X1 U17158 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n15514), .S(n15815), .Z(
        P1_U3515) );
  MUX2_X1 U17159 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n15515), .S(n15815), .Z(
        P1_U3513) );
  MUX2_X1 U17160 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n15516), .S(n15815), .Z(
        P1_U3510) );
  MUX2_X1 U17161 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n15517), .S(n15815), .Z(
        P1_U3507) );
  MUX2_X1 U17162 ( .A(P1_REG0_REG_15__SCAN_IN), .B(n15518), .S(n15815), .Z(
        P1_U3504) );
  MUX2_X1 U17163 ( .A(P1_REG0_REG_14__SCAN_IN), .B(n15519), .S(n15815), .Z(
        P1_U3501) );
  MUX2_X1 U17164 ( .A(P1_REG0_REG_13__SCAN_IN), .B(n15520), .S(n15815), .Z(
        P1_U3498) );
  MUX2_X1 U17165 ( .A(P1_REG0_REG_12__SCAN_IN), .B(n15521), .S(n15815), .Z(
        P1_U3495) );
  MUX2_X1 U17166 ( .A(P1_REG0_REG_11__SCAN_IN), .B(n15522), .S(n15815), .Z(
        P1_U3492) );
  MUX2_X1 U17167 ( .A(n15523), .B(P1_REG0_REG_10__SCAN_IN), .S(n15813), .Z(
        P1_U3489) );
  NOR4_X1 U17168 ( .A1(n15525), .A2(P1_IR_REG_30__SCAN_IN), .A3(n8645), .A4(
        P1_U3086), .ZN(n15526) );
  AOI21_X1 U17169 ( .B1(n15527), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n15526), 
        .ZN(n15528) );
  OAI21_X1 U17170 ( .B1(n15529), .B2(n15549), .A(n15528), .ZN(P1_U3324) );
  OAI222_X1 U17171 ( .A1(P1_U3086), .A2(n15532), .B1(n15549), .B2(n15531), 
        .C1(n15530), .C2(n15539), .ZN(P1_U3326) );
  OAI222_X1 U17172 ( .A1(n15546), .A2(n15535), .B1(n15549), .B2(n15534), .C1(
        P1_U3086), .C2(n15533), .ZN(P1_U3327) );
  OAI222_X1 U17173 ( .A1(n15546), .A2(n15538), .B1(n15549), .B2(n15537), .C1(
        n15536), .C2(P1_U3086), .ZN(P1_U3328) );
  OAI222_X1 U17174 ( .A1(P1_U3086), .A2(n15542), .B1(n15549), .B2(n15541), 
        .C1(n15540), .C2(n15539), .ZN(P1_U3329) );
  OAI222_X1 U17175 ( .A1(n15546), .A2(n15545), .B1(n15549), .B2(n15544), .C1(
        P1_U3086), .C2(n15543), .ZN(P1_U3330) );
  OAI222_X1 U17176 ( .A1(P1_U3086), .A2(n15550), .B1(n15549), .B2(n15548), 
        .C1(n15547), .C2(n15546), .ZN(P1_U3331) );
  MUX2_X1 U17177 ( .A(n15552), .B(n15551), .S(P1_U3086), .Z(P1_U3333) );
  INV_X1 U17178 ( .A(n15553), .ZN(n15554) );
  MUX2_X1 U17179 ( .A(n15554), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  INV_X1 U17180 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n15692) );
  XNOR2_X1 U17181 ( .A(n15622), .B(P1_ADDR_REG_14__SCAN_IN), .ZN(n15621) );
  NAND2_X1 U17182 ( .A1(P1_ADDR_REG_11__SCAN_IN), .A2(n15574), .ZN(n15555) );
  OAI21_X1 U17183 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(n15574), .A(n15555), 
        .ZN(n15613) );
  NAND2_X1 U17184 ( .A1(n15584), .A2(n15583), .ZN(n15560) );
  INV_X1 U17185 ( .A(n15558), .ZN(n15559) );
  INV_X1 U17186 ( .A(P3_ADDR_REG_5__SCAN_IN), .ZN(n15564) );
  NOR2_X1 U17187 ( .A1(n15565), .A2(n15564), .ZN(n15566) );
  XOR2_X1 U17188 ( .A(P1_ADDR_REG_6__SCAN_IN), .B(P3_ADDR_REG_6__SCAN_IN), .Z(
        n15599) );
  INV_X1 U17189 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n15567) );
  INV_X1 U17190 ( .A(P3_ADDR_REG_9__SCAN_IN), .ZN(n15570) );
  NOR2_X1 U17191 ( .A1(n15569), .A2(n15570), .ZN(n15571) );
  AND2_X1 U17192 ( .A1(n15573), .A2(P1_ADDR_REG_10__SCAN_IN), .ZN(n15572) );
  NAND2_X1 U17193 ( .A1(P1_ADDR_REG_12__SCAN_IN), .A2(n15576), .ZN(n15575) );
  OAI21_X1 U17194 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(n15576), .A(n15575), 
        .ZN(n15616) );
  XNOR2_X1 U17195 ( .A(P3_ADDR_REG_13__SCAN_IN), .B(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n15618) );
  XOR2_X1 U17196 ( .A(n15621), .B(n15620), .Z(n15687) );
  INV_X1 U17197 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n15658) );
  XNOR2_X1 U17198 ( .A(P3_ADDR_REG_10__SCAN_IN), .B(P1_ADDR_REG_10__SCAN_IN), 
        .ZN(n15579) );
  NAND2_X1 U17199 ( .A1(P2_ADDR_REG_4__SCAN_IN), .A2(n15582), .ZN(n15595) );
  XNOR2_X1 U17200 ( .A(n15584), .B(n15583), .ZN(n15644) );
  XOR2_X1 U17201 ( .A(n15585), .B(n15587), .Z(n15588) );
  OR2_X1 U17202 ( .A1(n15586), .A2(n15588), .ZN(n15590) );
  AOI21_X1 U17203 ( .B1(P1_ADDR_REG_0__SCAN_IN), .B2(n15926), .A(n15587), .ZN(
        n15978) );
  INV_X1 U17204 ( .A(P2_ADDR_REG_0__SCAN_IN), .ZN(n15977) );
  NOR2_X1 U17205 ( .A1(n15978), .A2(n15977), .ZN(n15986) );
  NAND2_X1 U17206 ( .A1(n15590), .A2(n15589), .ZN(n15645) );
  NAND2_X1 U17207 ( .A1(n15644), .A2(n15645), .ZN(n15591) );
  NOR2_X1 U17208 ( .A1(n15644), .A2(n15645), .ZN(n15643) );
  XNOR2_X1 U17209 ( .A(P1_ADDR_REG_3__SCAN_IN), .B(n15592), .ZN(n15983) );
  NOR2_X1 U17210 ( .A1(n15982), .A2(n15983), .ZN(n15593) );
  INV_X1 U17211 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n15842) );
  NAND2_X1 U17212 ( .A1(n15982), .A2(n15983), .ZN(n15981) );
  OAI21_X1 U17213 ( .B1(n15593), .B2(n15842), .A(n15981), .ZN(n15974) );
  XNOR2_X1 U17214 ( .A(P1_ADDR_REG_5__SCAN_IN), .B(n15596), .ZN(n15597) );
  XNOR2_X1 U17215 ( .A(n15600), .B(n15599), .ZN(n15648) );
  NAND2_X1 U17216 ( .A1(n15601), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n15602) );
  NAND2_X1 U17217 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(n15605), .ZN(n15608) );
  INV_X1 U17218 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n15604) );
  XNOR2_X1 U17219 ( .A(P1_ADDR_REG_7__SCAN_IN), .B(n15606), .ZN(n15979) );
  NAND2_X1 U17220 ( .A1(n15980), .A2(n15979), .ZN(n15607) );
  XNOR2_X1 U17221 ( .A(P1_ADDR_REG_8__SCAN_IN), .B(n15609), .ZN(n15610) );
  XOR2_X1 U17222 ( .A(n15614), .B(n15613), .Z(n15673) );
  XOR2_X1 U17223 ( .A(n15617), .B(n15616), .Z(n15678) );
  XNOR2_X1 U17224 ( .A(n15619), .B(n15618), .ZN(n15683) );
  INV_X1 U17225 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n15856) );
  INV_X1 U17226 ( .A(P3_ADDR_REG_15__SCAN_IN), .ZN(n15628) );
  NOR2_X1 U17227 ( .A1(P1_ADDR_REG_15__SCAN_IN), .A2(n15628), .ZN(n15623) );
  AOI21_X1 U17228 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(n15628), .A(n15623), 
        .ZN(n15625) );
  INV_X1 U17229 ( .A(P3_ADDR_REG_16__SCAN_IN), .ZN(n15631) );
  AOI22_X1 U17230 ( .A1(P1_ADDR_REG_16__SCAN_IN), .A2(n15631), .B1(
        P3_ADDR_REG_16__SCAN_IN), .B2(n15624), .ZN(n15630) );
  NAND2_X1 U17231 ( .A1(n15626), .A2(n15625), .ZN(n15627) );
  XNOR2_X1 U17232 ( .A(n15630), .B(n15629), .ZN(n15695) );
  XNOR2_X1 U17233 ( .A(n15632), .B(n15633), .ZN(n15660) );
  NAND2_X1 U17234 ( .A1(n15661), .A2(n15660), .ZN(n15635) );
  NAND2_X1 U17235 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(n15633), .ZN(n15634) );
  XNOR2_X1 U17236 ( .A(P3_ADDR_REG_18__SCAN_IN), .B(P1_ADDR_REG_18__SCAN_IN), 
        .ZN(n15665) );
  NAND2_X1 U17237 ( .A1(n15637), .A2(n15636), .ZN(n15640) );
  NAND2_X1 U17238 ( .A1(P3_ADDR_REG_17__SCAN_IN), .A2(n15638), .ZN(n15639) );
  NAND2_X1 U17239 ( .A1(n15640), .A2(n15639), .ZN(n15664) );
  XNOR2_X1 U17240 ( .A(n15665), .B(n15664), .ZN(n15663) );
  XNOR2_X1 U17241 ( .A(P2_ADDR_REG_18__SCAN_IN), .B(n15662), .ZN(SUB_1596_U62)
         );
  AOI21_X1 U17242 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(
        P3_WR_REG_SCAN_IN), .ZN(n15641) );
  OAI21_X1 U17243 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(n15641), 
        .ZN(U28) );
  AOI21_X1 U17244 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(
        P3_RD_REG_SCAN_IN), .ZN(n15642) );
  OAI21_X1 U17245 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(n15642), 
        .ZN(U29) );
  AOI21_X1 U17246 ( .B1(n15645), .B2(n15644), .A(n15643), .ZN(n15647) );
  XNOR2_X1 U17247 ( .A(n15647), .B(n15646), .ZN(SUB_1596_U61) );
  XOR2_X1 U17248 ( .A(n15649), .B(n15648), .Z(SUB_1596_U57) );
  XNOR2_X1 U17249 ( .A(P2_ADDR_REG_8__SCAN_IN), .B(n15650), .ZN(SUB_1596_U55)
         );
  AOI21_X1 U17250 ( .B1(n15652), .B2(n15651), .A(n6714), .ZN(n15654) );
  XNOR2_X1 U17251 ( .A(n15654), .B(n15653), .ZN(SUB_1596_U54) );
  AOI21_X1 U17252 ( .B1(n15657), .B2(n15656), .A(n15655), .ZN(n15659) );
  XNOR2_X1 U17253 ( .A(n15659), .B(n15658), .ZN(SUB_1596_U70) );
  XOR2_X1 U17254 ( .A(n15661), .B(n15660), .Z(SUB_1596_U63) );
  NAND2_X1 U17255 ( .A1(n15665), .A2(n15664), .ZN(n15666) );
  OAI21_X1 U17256 ( .B1(n13110), .B2(P1_ADDR_REG_18__SCAN_IN), .A(n15666), 
        .ZN(n15669) );
  XNOR2_X1 U17257 ( .A(P2_ADDR_REG_19__SCAN_IN), .B(P1_ADDR_REG_19__SCAN_IN), 
        .ZN(n15667) );
  XNOR2_X1 U17258 ( .A(n15667), .B(P3_ADDR_REG_19__SCAN_IN), .ZN(n15668) );
  XNOR2_X1 U17259 ( .A(n15669), .B(n15668), .ZN(n15670) );
  AOI21_X1 U17260 ( .B1(n15674), .B2(n15673), .A(n15672), .ZN(n15675) );
  XNOR2_X1 U17261 ( .A(n15675), .B(n7713), .ZN(SUB_1596_U69) );
  AOI21_X1 U17262 ( .B1(n15678), .B2(n15677), .A(n15676), .ZN(n15680) );
  XNOR2_X1 U17263 ( .A(n15680), .B(n15679), .ZN(SUB_1596_U68) );
  OAI21_X1 U17264 ( .B1(n15683), .B2(n15682), .A(n15681), .ZN(n15684) );
  XNOR2_X1 U17265 ( .A(n15684), .B(P2_ADDR_REG_13__SCAN_IN), .ZN(SUB_1596_U67)
         );
  AOI21_X1 U17266 ( .B1(n15687), .B2(n15686), .A(n15685), .ZN(n15688) );
  XNOR2_X1 U17267 ( .A(n15688), .B(n12303), .ZN(SUB_1596_U66) );
  AOI21_X1 U17268 ( .B1(n15691), .B2(n15690), .A(n15689), .ZN(n15693) );
  XNOR2_X1 U17269 ( .A(n15693), .B(n15692), .ZN(SUB_1596_U65) );
  AOI21_X1 U17270 ( .B1(n15696), .B2(n15695), .A(n15694), .ZN(n15698) );
  XNOR2_X1 U17271 ( .A(n15698), .B(n15697), .ZN(SUB_1596_U64) );
  INV_X1 U17272 ( .A(n15699), .ZN(n15704) );
  NAND2_X1 U17273 ( .A1(n15701), .A2(n6534), .ZN(n15787) );
  INV_X1 U17274 ( .A(n15787), .ZN(n15703) );
  AOI21_X1 U17275 ( .B1(n15704), .B2(n15703), .A(n15702), .ZN(n15712) );
  XOR2_X1 U17276 ( .A(n15706), .B(n15705), .Z(n15710) );
  AOI22_X1 U17277 ( .A1(n15710), .A2(n15709), .B1(n15708), .B2(n15707), .ZN(
        n15711) );
  OAI211_X1 U17278 ( .C1(P1_REG3_REG_3__SCAN_IN), .C2(n15713), .A(n15712), .B(
        n15711), .ZN(P1_U3218) );
  NOR2_X1 U17279 ( .A1(n15714), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n15716) );
  OR2_X1 U17280 ( .A1(n15715), .A2(n15716), .ZN(n15719) );
  INV_X1 U17281 ( .A(n15716), .ZN(n15718) );
  MUX2_X1 U17282 ( .A(n15719), .B(n15718), .S(n15717), .Z(n15721) );
  NAND2_X1 U17283 ( .A1(n15721), .A2(n15720), .ZN(n15724) );
  AOI22_X1 U17284 ( .A1(n15722), .A2(P1_ADDR_REG_0__SCAN_IN), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(P1_U3086), .ZN(n15723) );
  OAI21_X1 U17285 ( .B1(n15725), .B2(n15724), .A(n15723), .ZN(P1_U3243) );
  INV_X1 U17286 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n15737) );
  INV_X1 U17287 ( .A(n15726), .ZN(n15728) );
  OAI21_X1 U17288 ( .B1(n15729), .B2(n15728), .A(n15727), .ZN(n15734) );
  XNOR2_X1 U17289 ( .A(n15731), .B(n15730), .ZN(n15733) );
  AOI222_X1 U17290 ( .A1(n15734), .A2(n15746), .B1(n15745), .B2(n15733), .C1(
        n15732), .C2(n15742), .ZN(n15736) );
  OAI211_X1 U17291 ( .C1(n15737), .C2(n15750), .A(n15736), .B(n15735), .ZN(
        P1_U3255) );
  OAI21_X1 U17292 ( .B1(n15740), .B2(n15739), .A(n15738), .ZN(n15747) );
  XNOR2_X1 U17293 ( .A(n15741), .B(P1_REG1_REG_15__SCAN_IN), .ZN(n15744) );
  AOI222_X1 U17294 ( .A1(n15747), .A2(n15746), .B1(n15745), .B2(n15744), .C1(
        n15743), .C2(n15742), .ZN(n15749) );
  OAI211_X1 U17295 ( .C1(n7509), .C2(n15750), .A(n15749), .B(n15748), .ZN(
        P1_U3258) );
  INV_X1 U17296 ( .A(P1_D_REG_31__SCAN_IN), .ZN(n15751) );
  NOR2_X1 U17297 ( .A1(n15781), .A2(n15751), .ZN(P1_U3294) );
  INV_X1 U17298 ( .A(P1_D_REG_30__SCAN_IN), .ZN(n15752) );
  NOR2_X1 U17299 ( .A1(n15781), .A2(n15752), .ZN(P1_U3295) );
  INV_X1 U17300 ( .A(P1_D_REG_29__SCAN_IN), .ZN(n15753) );
  NOR2_X1 U17301 ( .A1(n15781), .A2(n15753), .ZN(P1_U3296) );
  NOR2_X1 U17302 ( .A1(n15781), .A2(n15754), .ZN(P1_U3297) );
  INV_X1 U17303 ( .A(P1_D_REG_27__SCAN_IN), .ZN(n15755) );
  NOR2_X1 U17304 ( .A1(n15781), .A2(n15755), .ZN(P1_U3298) );
  INV_X1 U17305 ( .A(P1_D_REG_26__SCAN_IN), .ZN(n15756) );
  NOR2_X1 U17306 ( .A1(n15781), .A2(n15756), .ZN(P1_U3299) );
  INV_X1 U17307 ( .A(P1_D_REG_25__SCAN_IN), .ZN(n15757) );
  NOR2_X1 U17308 ( .A1(n15781), .A2(n15757), .ZN(P1_U3300) );
  INV_X1 U17309 ( .A(P1_D_REG_24__SCAN_IN), .ZN(n15758) );
  NOR2_X1 U17310 ( .A1(n15781), .A2(n15758), .ZN(P1_U3301) );
  INV_X1 U17311 ( .A(P1_D_REG_23__SCAN_IN), .ZN(n15759) );
  NOR2_X1 U17312 ( .A1(n15781), .A2(n15759), .ZN(P1_U3302) );
  INV_X1 U17313 ( .A(P1_D_REG_22__SCAN_IN), .ZN(n15760) );
  NOR2_X1 U17314 ( .A1(n15781), .A2(n15760), .ZN(P1_U3303) );
  INV_X1 U17315 ( .A(P1_D_REG_21__SCAN_IN), .ZN(n15761) );
  NOR2_X1 U17316 ( .A1(n15781), .A2(n15761), .ZN(P1_U3304) );
  INV_X1 U17317 ( .A(P1_D_REG_20__SCAN_IN), .ZN(n15762) );
  NOR2_X1 U17318 ( .A1(n15781), .A2(n15762), .ZN(P1_U3305) );
  INV_X1 U17319 ( .A(P1_D_REG_19__SCAN_IN), .ZN(n15763) );
  NOR2_X1 U17320 ( .A1(n15781), .A2(n15763), .ZN(P1_U3306) );
  NOR2_X1 U17321 ( .A1(n15781), .A2(n15764), .ZN(P1_U3307) );
  INV_X1 U17322 ( .A(P1_D_REG_17__SCAN_IN), .ZN(n15765) );
  NOR2_X1 U17323 ( .A1(n15781), .A2(n15765), .ZN(P1_U3308) );
  INV_X1 U17324 ( .A(P1_D_REG_16__SCAN_IN), .ZN(n15766) );
  NOR2_X1 U17325 ( .A1(n15781), .A2(n15766), .ZN(P1_U3309) );
  INV_X1 U17326 ( .A(P1_D_REG_15__SCAN_IN), .ZN(n15767) );
  NOR2_X1 U17327 ( .A1(n15781), .A2(n15767), .ZN(P1_U3310) );
  INV_X1 U17328 ( .A(P1_D_REG_14__SCAN_IN), .ZN(n15768) );
  NOR2_X1 U17329 ( .A1(n15781), .A2(n15768), .ZN(P1_U3311) );
  NOR2_X1 U17330 ( .A1(n15781), .A2(n15769), .ZN(P1_U3312) );
  INV_X1 U17331 ( .A(P1_D_REG_12__SCAN_IN), .ZN(n15770) );
  NOR2_X1 U17332 ( .A1(n15781), .A2(n15770), .ZN(P1_U3313) );
  INV_X1 U17333 ( .A(P1_D_REG_11__SCAN_IN), .ZN(n15771) );
  NOR2_X1 U17334 ( .A1(n15781), .A2(n15771), .ZN(P1_U3314) );
  INV_X1 U17335 ( .A(P1_D_REG_10__SCAN_IN), .ZN(n15772) );
  NOR2_X1 U17336 ( .A1(n15781), .A2(n15772), .ZN(P1_U3315) );
  INV_X1 U17337 ( .A(P1_D_REG_9__SCAN_IN), .ZN(n15773) );
  NOR2_X1 U17338 ( .A1(n15781), .A2(n15773), .ZN(P1_U3316) );
  INV_X1 U17339 ( .A(P1_D_REG_8__SCAN_IN), .ZN(n15774) );
  NOR2_X1 U17340 ( .A1(n15781), .A2(n15774), .ZN(P1_U3317) );
  INV_X1 U17341 ( .A(P1_D_REG_7__SCAN_IN), .ZN(n15775) );
  NOR2_X1 U17342 ( .A1(n15781), .A2(n15775), .ZN(P1_U3318) );
  NOR2_X1 U17343 ( .A1(n15781), .A2(n15776), .ZN(P1_U3319) );
  INV_X1 U17344 ( .A(P1_D_REG_5__SCAN_IN), .ZN(n15777) );
  NOR2_X1 U17345 ( .A1(n15781), .A2(n15777), .ZN(P1_U3320) );
  INV_X1 U17346 ( .A(P1_D_REG_4__SCAN_IN), .ZN(n15778) );
  NOR2_X1 U17347 ( .A1(n15781), .A2(n15778), .ZN(P1_U3321) );
  INV_X1 U17348 ( .A(P1_D_REG_3__SCAN_IN), .ZN(n15779) );
  NOR2_X1 U17349 ( .A1(n15781), .A2(n15779), .ZN(P1_U3322) );
  NOR2_X1 U17350 ( .A1(n15781), .A2(n15780), .ZN(P1_U3323) );
  OAI21_X1 U17351 ( .B1(n15783), .B2(n15804), .A(n15782), .ZN(n15785) );
  AOI211_X1 U17352 ( .C1(n15812), .C2(n15786), .A(n15785), .B(n15784), .ZN(
        n15816) );
  AOI22_X1 U17353 ( .A1(n15815), .A2(n15816), .B1(n8663), .B2(n15813), .ZN(
        P1_U3462) );
  AND3_X1 U17354 ( .A1(n15789), .A2(n15788), .A3(n15787), .ZN(n15817) );
  AOI22_X1 U17355 ( .A1(n15815), .A2(n15817), .B1(n8694), .B2(n15813), .ZN(
        P1_U3468) );
  OAI211_X1 U17356 ( .C1(n7943), .C2(n15804), .A(n15791), .B(n15790), .ZN(
        n15792) );
  INV_X1 U17357 ( .A(n15792), .ZN(n15818) );
  AOI22_X1 U17358 ( .A1(n15815), .A2(n15818), .B1(n8764), .B2(n15813), .ZN(
        P1_U3477) );
  OAI211_X1 U17359 ( .C1(n15795), .C2(n15804), .A(n15794), .B(n15793), .ZN(
        n15796) );
  INV_X1 U17360 ( .A(n15796), .ZN(n15819) );
  INV_X1 U17361 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n15797) );
  AOI22_X1 U17362 ( .A1(n15815), .A2(n15819), .B1(n15797), .B2(n15813), .ZN(
        P1_U3480) );
  AOI22_X1 U17363 ( .A1(n15801), .A2(n15800), .B1(n15799), .B2(n15798), .ZN(
        n15802) );
  OAI211_X1 U17364 ( .C1(n15805), .C2(n15804), .A(n15803), .B(n15802), .ZN(
        n15810) );
  AND3_X1 U17365 ( .A1(n15808), .A2(n15807), .A3(n15806), .ZN(n15809) );
  AOI211_X1 U17366 ( .C1(n15812), .C2(n15811), .A(n15810), .B(n15809), .ZN(
        n15821) );
  INV_X1 U17367 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n15814) );
  AOI22_X1 U17368 ( .A1(n15815), .A2(n15821), .B1(n15814), .B2(n15813), .ZN(
        P1_U3483) );
  AOI22_X1 U17369 ( .A1(n15822), .A2(n15816), .B1(n8664), .B2(n15820), .ZN(
        P1_U3529) );
  AOI22_X1 U17370 ( .A1(n15822), .A2(n15817), .B1(n10744), .B2(n15820), .ZN(
        P1_U3531) );
  AOI22_X1 U17371 ( .A1(n15822), .A2(n15818), .B1(n10818), .B2(n15820), .ZN(
        P1_U3534) );
  AOI22_X1 U17372 ( .A1(n15822), .A2(n15819), .B1(n10840), .B2(n15820), .ZN(
        P1_U3535) );
  AOI22_X1 U17373 ( .A1(n15822), .A2(n15821), .B1(n11147), .B2(n15820), .ZN(
        P1_U3536) );
  NOR2_X1 U17374 ( .A1(n15864), .A2(P2_U3947), .ZN(P2_U3087) );
  AOI22_X1 U17375 ( .A1(P2_REG1_REG_0__SCAN_IN), .A2(n15830), .B1(n15866), 
        .B2(P2_REG2_REG_0__SCAN_IN), .ZN(n15828) );
  OAI22_X1 U17376 ( .A1(n15823), .A2(P2_REG2_REG_0__SCAN_IN), .B1(
        P2_REG1_REG_0__SCAN_IN), .B2(n15860), .ZN(n15824) );
  NOR2_X1 U17377 ( .A1(n15850), .A2(n15824), .ZN(n15826) );
  AOI22_X1 U17378 ( .A1(n15864), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3088), .ZN(n15825) );
  OAI221_X1 U17379 ( .B1(P2_IR_REG_0__SCAN_IN), .B2(n15828), .C1(n15827), .C2(
        n15826), .A(n15825), .ZN(P2_U3214) );
  AND2_X1 U17380 ( .A1(P2_U3088), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n15835) );
  OAI211_X1 U17381 ( .C1(n15832), .C2(n15831), .A(n15830), .B(n15829), .ZN(
        n15833) );
  INV_X1 U17382 ( .A(n15833), .ZN(n15834) );
  AOI211_X1 U17383 ( .C1(n15850), .C2(n15836), .A(n15835), .B(n15834), .ZN(
        n15841) );
  OAI211_X1 U17384 ( .C1(n15839), .C2(n15838), .A(n15866), .B(n15837), .ZN(
        n15840) );
  OAI211_X1 U17385 ( .C1(n15857), .C2(n15842), .A(n15841), .B(n15840), .ZN(
        P2_U3217) );
  NOR2_X1 U17386 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n15843), .ZN(n15848) );
  AOI211_X1 U17387 ( .C1(n15846), .C2(n15845), .A(n15860), .B(n15844), .ZN(
        n15847) );
  AOI211_X1 U17388 ( .C1(n15850), .C2(n15849), .A(n15848), .B(n15847), .ZN(
        n15855) );
  OAI211_X1 U17389 ( .C1(n15853), .C2(n15852), .A(n15851), .B(n15866), .ZN(
        n15854) );
  OAI211_X1 U17390 ( .C1(n15857), .C2(n15856), .A(n15855), .B(n15854), .ZN(
        P2_U3227) );
  INV_X1 U17391 ( .A(n15858), .ZN(n15863) );
  INV_X1 U17392 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n15861) );
  AOI211_X1 U17393 ( .C1(n15861), .C2(n6614), .A(n15860), .B(n15859), .ZN(
        n15862) );
  AOI211_X1 U17394 ( .C1(P2_ADDR_REG_18__SCAN_IN), .C2(n15864), .A(n15863), 
        .B(n15862), .ZN(n15869) );
  XOR2_X1 U17395 ( .A(P2_REG2_REG_18__SCAN_IN), .B(n15865), .Z(n15867) );
  NAND2_X1 U17396 ( .A1(n15867), .A2(n15866), .ZN(n15868) );
  OAI211_X1 U17397 ( .C1(n15871), .C2(n15870), .A(n15869), .B(n15868), .ZN(
        P2_U3232) );
  AND2_X1 U17398 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n15877), .ZN(P2_U3266) );
  AND2_X1 U17399 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n15877), .ZN(P2_U3267) );
  AND2_X1 U17400 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n15877), .ZN(P2_U3268) );
  AND2_X1 U17401 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n15877), .ZN(P2_U3269) );
  AND2_X1 U17402 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n15877), .ZN(P2_U3270) );
  AND2_X1 U17403 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n15877), .ZN(P2_U3271) );
  AND2_X1 U17404 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n15877), .ZN(P2_U3272) );
  AND2_X1 U17405 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n15877), .ZN(P2_U3273) );
  AND2_X1 U17406 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n15877), .ZN(P2_U3274) );
  NOR2_X1 U17407 ( .A1(n15879), .A2(n15873), .ZN(P2_U3275) );
  AND2_X1 U17408 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n15877), .ZN(P2_U3276) );
  NOR2_X1 U17409 ( .A1(n15879), .A2(n15874), .ZN(P2_U3277) );
  AND2_X1 U17410 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n15877), .ZN(P2_U3278) );
  AND2_X1 U17411 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n15877), .ZN(P2_U3279) );
  AND2_X1 U17412 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n15877), .ZN(P2_U3280) );
  AND2_X1 U17413 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n15877), .ZN(P2_U3281) );
  AND2_X1 U17414 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n15877), .ZN(P2_U3282) );
  AND2_X1 U17415 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n15877), .ZN(P2_U3283) );
  AND2_X1 U17416 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n15877), .ZN(P2_U3284) );
  NOR2_X1 U17417 ( .A1(n15879), .A2(n15875), .ZN(P2_U3285) );
  AND2_X1 U17418 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n15877), .ZN(P2_U3286) );
  AND2_X1 U17419 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n15877), .ZN(P2_U3287) );
  AND2_X1 U17420 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n15877), .ZN(P2_U3288) );
  NOR2_X1 U17421 ( .A1(n15879), .A2(n15876), .ZN(P2_U3289) );
  AND2_X1 U17422 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n15877), .ZN(P2_U3290) );
  AND2_X1 U17423 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n15877), .ZN(P2_U3291) );
  AND2_X1 U17424 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n15877), .ZN(P2_U3292) );
  AND2_X1 U17425 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n15877), .ZN(P2_U3293) );
  AND2_X1 U17426 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n15877), .ZN(P2_U3294) );
  NOR2_X1 U17427 ( .A1(n15879), .A2(n15878), .ZN(P2_U3295) );
  AOI22_X1 U17428 ( .A1(n15882), .A2(n15881), .B1(n15880), .B2(n15884), .ZN(
        P2_U3416) );
  AOI21_X1 U17429 ( .B1(n15885), .B2(n15884), .A(n15883), .ZN(P2_U3417) );
  AOI22_X1 U17430 ( .A1(n15908), .A2(n15887), .B1(n15886), .B2(n15906), .ZN(
        P2_U3430) );
  INV_X1 U17431 ( .A(n15888), .ZN(n15895) );
  INV_X1 U17432 ( .A(n15889), .ZN(n15892) );
  OAI22_X1 U17433 ( .A1(n15892), .A2(n15891), .B1(n7804), .B2(n15900), .ZN(
        n15894) );
  AOI211_X1 U17434 ( .C1(n15905), .C2(n15895), .A(n15894), .B(n15893), .ZN(
        n15909) );
  INV_X1 U17435 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n15896) );
  AOI22_X1 U17436 ( .A1(n15908), .A2(n15909), .B1(n15896), .B2(n15906), .ZN(
        P2_U3439) );
  INV_X1 U17437 ( .A(n15897), .ZN(n15904) );
  INV_X1 U17438 ( .A(n15898), .ZN(n15899) );
  OAI21_X1 U17439 ( .B1(n15901), .B2(n15900), .A(n15899), .ZN(n15903) );
  AOI211_X1 U17440 ( .C1(n15905), .C2(n15904), .A(n15903), .B(n15902), .ZN(
        n15911) );
  AOI22_X1 U17441 ( .A1(n15908), .A2(n15911), .B1(n15907), .B2(n15906), .ZN(
        P2_U3448) );
  AOI22_X1 U17442 ( .A1(n15912), .A2(n15909), .B1(n10694), .B2(n15910), .ZN(
        P2_U3502) );
  AOI22_X1 U17443 ( .A1(n15912), .A2(n15911), .B1(n10697), .B2(n15910), .ZN(
        P2_U3505) );
  NOR2_X1 U17444 ( .A1(P3_U3897), .A2(n15913), .ZN(P3_U3150) );
  NOR3_X1 U17445 ( .A1(n15916), .A2(n15915), .A3(n15914), .ZN(n15921) );
  AOI21_X1 U17446 ( .B1(n15919), .B2(n15918), .A(n15917), .ZN(n15920) );
  OR2_X1 U17447 ( .A1(n15921), .A2(n15920), .ZN(n15924) );
  AOI22_X1 U17448 ( .A1(n15922), .A2(P3_IR_REG_0__SCAN_IN), .B1(
        P3_REG3_REG_0__SCAN_IN), .B2(P3_U3151), .ZN(n15923) );
  OAI211_X1 U17449 ( .C1(n15926), .C2(n15925), .A(n15924), .B(n15923), .ZN(
        P3_U3182) );
  INV_X1 U17450 ( .A(n15927), .ZN(n15931) );
  INV_X1 U17451 ( .A(n15956), .ZN(n15930) );
  AOI211_X1 U17452 ( .C1(n15931), .C2(n15930), .A(n15929), .B(n15928), .ZN(
        n15964) );
  INV_X1 U17453 ( .A(P3_REG0_REG_2__SCAN_IN), .ZN(n15932) );
  AOI22_X1 U17454 ( .A1(n15963), .A2(n15964), .B1(n15932), .B2(n15961), .ZN(
        P3_U3396) );
  INV_X1 U17455 ( .A(n15957), .ZN(n15953) );
  INV_X1 U17456 ( .A(n15937), .ZN(n15934) );
  OAI22_X1 U17457 ( .A1(n15934), .A2(n15956), .B1(n15933), .B2(n15946), .ZN(
        n15935) );
  AOI211_X1 U17458 ( .C1(n15953), .C2(n15937), .A(n15936), .B(n15935), .ZN(
        n15965) );
  INV_X1 U17459 ( .A(P3_REG0_REG_3__SCAN_IN), .ZN(n15938) );
  AOI22_X1 U17460 ( .A1(n15963), .A2(n15965), .B1(n15938), .B2(n15961), .ZN(
        P3_U3399) );
  INV_X1 U17461 ( .A(n15940), .ZN(n15944) );
  OAI22_X1 U17462 ( .A1(n15940), .A2(n15956), .B1(n15939), .B2(n15946), .ZN(
        n15943) );
  INV_X1 U17463 ( .A(n15941), .ZN(n15942) );
  AOI211_X1 U17464 ( .C1(n15953), .C2(n15944), .A(n15943), .B(n15942), .ZN(
        n15967) );
  INV_X1 U17465 ( .A(P3_REG0_REG_4__SCAN_IN), .ZN(n15945) );
  AOI22_X1 U17466 ( .A1(n15963), .A2(n15967), .B1(n15945), .B2(n15961), .ZN(
        P3_U3402) );
  INV_X1 U17467 ( .A(n15948), .ZN(n15952) );
  OAI22_X1 U17468 ( .A1(n15948), .A2(n15956), .B1(n15947), .B2(n15946), .ZN(
        n15951) );
  INV_X1 U17469 ( .A(n15949), .ZN(n15950) );
  AOI211_X1 U17470 ( .C1(n15953), .C2(n15952), .A(n15951), .B(n15950), .ZN(
        n15969) );
  INV_X1 U17471 ( .A(P3_REG0_REG_5__SCAN_IN), .ZN(n15954) );
  AOI22_X1 U17472 ( .A1(n15963), .A2(n15969), .B1(n15954), .B2(n15961), .ZN(
        P3_U3405) );
  AOI21_X1 U17473 ( .B1(n15957), .B2(n15956), .A(n15955), .ZN(n15958) );
  AOI211_X1 U17474 ( .C1(n15960), .C2(n6977), .A(n15959), .B(n15958), .ZN(
        n15972) );
  INV_X1 U17475 ( .A(P3_REG0_REG_6__SCAN_IN), .ZN(n15962) );
  AOI22_X1 U17476 ( .A1(n15963), .A2(n15972), .B1(n15962), .B2(n15961), .ZN(
        P3_U3408) );
  AOI22_X1 U17477 ( .A1(n15973), .A2(n15964), .B1(n10926), .B2(n15970), .ZN(
        P3_U3461) );
  AOI22_X1 U17478 ( .A1(n15973), .A2(n15965), .B1(n6803), .B2(n15970), .ZN(
        P3_U3462) );
  AOI22_X1 U17479 ( .A1(n15973), .A2(n15967), .B1(n15966), .B2(n15970), .ZN(
        P3_U3463) );
  AOI22_X1 U17480 ( .A1(n15973), .A2(n15969), .B1(n15968), .B2(n15970), .ZN(
        P3_U3464) );
  AOI22_X1 U17481 ( .A1(n15973), .A2(n15972), .B1(n15971), .B2(n15970), .ZN(
        P3_U3465) );
  XOR2_X1 U17482 ( .A(n15975), .B(n15974), .Z(SUB_1596_U59) );
  XNOR2_X1 U17483 ( .A(n15976), .B(P2_ADDR_REG_5__SCAN_IN), .ZN(SUB_1596_U58)
         );
  AOI21_X1 U17484 ( .B1(n15978), .B2(n15977), .A(n15986), .ZN(SUB_1596_U53) );
  XOR2_X1 U17485 ( .A(n15980), .B(n15979), .Z(SUB_1596_U56) );
  OAI21_X1 U17486 ( .B1(n15983), .B2(n15982), .A(n15981), .ZN(n15984) );
  XNOR2_X1 U17487 ( .A(n15984), .B(P2_ADDR_REG_3__SCAN_IN), .ZN(SUB_1596_U60)
         );
  XOR2_X1 U17488 ( .A(n15986), .B(n15985), .Z(SUB_1596_U5) );
  NAND2_X1 U9707 ( .A1(n8825), .A2(n8824), .ZN(n12112) );
  NAND2_X1 U10179 ( .A1(n8011), .A2(n8013), .ZN(n11912) );
  NAND2_X2 U9704 ( .A1(n12264), .A2(n14937), .ZN(n12263) );
  NAND2_X1 U11346 ( .A1(n8691), .A2(n14693), .ZN(n11517) );
  AND4_X2 U9608 ( .A1(n7555), .A2(n7556), .A3(n7557), .A4(n9212), .ZN(n6652)
         );
  NAND2_X2 U11767 ( .A1(n11372), .A2(n11385), .ZN(n11384) );
  INV_X2 U9701 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n9212) );
  NAND2_X1 U8573 ( .A1(n14705), .A2(n9141), .ZN(n11372) );
  AND2_X2 U7540 ( .A1(n8636), .A2(n8635), .ZN(n7556) );
  INV_X1 U7348 ( .A(n14729), .ZN(n7943) );
  INV_X2 U7380 ( .A(n14307), .ZN(n14261) );
  INV_X2 U7289 ( .A(n14719), .ZN(n14864) );
  NOR2_X1 U7304 ( .A1(P1_IR_REG_27__SCAN_IN), .A2(n8026), .ZN(n8025) );
  NOR2_X1 U7309 ( .A1(P1_IR_REG_14__SCAN_IN), .A2(P1_IR_REG_13__SCAN_IN), .ZN(
        n8635) );
  NAND2_X1 U7343 ( .A1(n11166), .A2(n10294), .ZN(n14705) );
  CLKBUF_X1 U7346 ( .A(n12461), .Z(n6525) );
  CLKBUF_X2 U7349 ( .A(n9562), .Z(n10053) );
  CLKBUF_X1 U7350 ( .A(n10296), .Z(n14526) );
  CLKBUF_X2 U7351 ( .A(n13111), .Z(n6527) );
  CLKBUF_X2 U7353 ( .A(n8198), .Z(n8466) );
  CLKBUF_X2 U7373 ( .A(n13111), .Z(n7233) );
  CLKBUF_X1 U7376 ( .A(n14295), .Z(n7352) );
  CLKBUF_X1 U7377 ( .A(n8778), .Z(n10490) );
  CLKBUF_X2 U7390 ( .A(n11410), .Z(n6528) );
  CLKBUF_X1 U7514 ( .A(n15252), .Z(n7226) );
  OR2_X1 U7531 ( .A1(n12765), .A2(n15119), .ZN(n15360) );
  CLKBUF_X1 U7535 ( .A(n10944), .Z(n7298) );
  INV_X1 U7547 ( .A(n15168), .ZN(n15187) );
  NAND3_X1 U7920 ( .A1(n8028), .A2(n8657), .A3(n8656), .ZN(n10283) );
endmodule

