

module b22_C_gen_AntiSAT_k_128_5 ( P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN, 
        P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN, 
        P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN, 
        P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN, 
        P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN, 
        P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN, 
        P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN, 
        P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN, 
        P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN, 
        P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN, P3_REG3_REG_0__SCAN_IN, 
        P3_REG3_REG_20__SCAN_IN, P3_REG3_REG_13__SCAN_IN, 
        P3_REG3_REG_22__SCAN_IN, P3_REG3_REG_11__SCAN_IN, 
        P3_REG3_REG_2__SCAN_IN, P3_REG3_REG_18__SCAN_IN, 
        P3_REG3_REG_6__SCAN_IN, P3_REG3_REG_26__SCAN_IN, 
        P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_ADDR_REG_0__SCAN_IN, 
        P3_ADDR_REG_1__SCAN_IN, P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN, 
        P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN, P3_ADDR_REG_6__SCAN_IN, 
        P3_ADDR_REG_7__SCAN_IN, P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, 
        P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, 
        P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, 
        P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, 
        P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, 
        P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, 
        P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, 
        P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, 
        P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, 
        P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, 
        P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, 
        P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, 
        P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, 
        P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, 
        P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, 
        P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, 
        P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, 
        P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, 
        P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, 
        P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, 
        P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, 
        P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, 
        P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, 
        P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, 
        P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, 
        P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, 
        P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN, 
        P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN, 
        P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN, 
        P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN, 
        P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN, 
        P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN, 
        P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN, 
        P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN, 
        P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN, 
        P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN, 
        P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN, 
        P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN, 
        P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN, 
        P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN, 
        P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN, 
        P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN, 
        P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN, 
        P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_4__SCAN_IN, 
        P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_17__SCAN_IN, 
        P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_16__SCAN_IN, 
        P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_12__SCAN_IN, 
        P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_1__SCAN_IN, 
        P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_28__SCAN_IN, 
        P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_3__SCAN_IN, 
        P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_23__SCAN_IN, 
        P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_27__SCAN_IN, 
        P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN, P2_RD_REG_SCAN_IN, 
        P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN, P3_IR_REG_1__SCAN_IN, 
        P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN, P3_IR_REG_4__SCAN_IN, 
        P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN, P3_IR_REG_7__SCAN_IN, 
        P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN, P3_IR_REG_10__SCAN_IN, 
        P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN, P3_IR_REG_13__SCAN_IN, 
        P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN, P3_IR_REG_16__SCAN_IN, 
        P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN, P3_IR_REG_19__SCAN_IN, 
        P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN, P3_IR_REG_22__SCAN_IN, 
        P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN, P3_IR_REG_25__SCAN_IN, 
        P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN, P3_IR_REG_28__SCAN_IN, 
        P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN, P3_IR_REG_31__SCAN_IN, 
        P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN, P3_D_REG_2__SCAN_IN, 
        P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN, P3_D_REG_5__SCAN_IN, 
        P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN, P3_D_REG_8__SCAN_IN, 
        P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN, P3_D_REG_11__SCAN_IN, 
        P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN, P3_D_REG_14__SCAN_IN, 
        P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN, P3_D_REG_17__SCAN_IN, 
        P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN, P3_D_REG_20__SCAN_IN, 
        P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN, P3_D_REG_23__SCAN_IN, 
        P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN, P3_D_REG_26__SCAN_IN, 
        P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN, P3_D_REG_29__SCAN_IN, 
        P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN, P3_REG0_REG_0__SCAN_IN, 
        P3_REG0_REG_1__SCAN_IN, P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN, 
        P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN, P3_REG0_REG_6__SCAN_IN, 
        P3_REG0_REG_7__SCAN_IN, P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN, 
        P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN, 
        P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN, 
        P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN, 
        P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN, 
        P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN, 
        P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN, 
        P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN, 
        P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN, 
        P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN, 
        P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN, 
        P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN, 
        P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN, P3_REG1_REG_2__SCAN_IN, 
        P3_REG1_REG_3__SCAN_IN, P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN, 
        P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN, P3_REG1_REG_8__SCAN_IN, 
        P3_REG1_REG_9__SCAN_IN, P3_REG1_REG_10__SCAN_IN, 
        P3_REG1_REG_11__SCAN_IN, P3_REG1_REG_12__SCAN_IN, 
        P3_REG1_REG_13__SCAN_IN, P3_REG1_REG_14__SCAN_IN, 
        P3_REG1_REG_15__SCAN_IN, P3_REG1_REG_16__SCAN_IN, 
        P3_REG1_REG_17__SCAN_IN, P3_REG1_REG_18__SCAN_IN, 
        P3_REG1_REG_19__SCAN_IN, P3_REG1_REG_20__SCAN_IN, 
        P3_REG1_REG_21__SCAN_IN, P3_REG1_REG_22__SCAN_IN, 
        P3_REG1_REG_23__SCAN_IN, P3_REG1_REG_24__SCAN_IN, 
        P3_REG1_REG_25__SCAN_IN, P3_REG1_REG_26__SCAN_IN, 
        P3_REG1_REG_27__SCAN_IN, P3_REG1_REG_28__SCAN_IN, 
        P3_REG1_REG_29__SCAN_IN, P3_REG1_REG_30__SCAN_IN, 
        P3_REG1_REG_31__SCAN_IN, P3_REG2_REG_0__SCAN_IN, 
        P3_REG2_REG_1__SCAN_IN, P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN, 
        P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN, P3_REG2_REG_6__SCAN_IN, 
        P3_REG2_REG_7__SCAN_IN, P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN, 
        P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN, 
        P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN, 
        P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN, 
        P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN, 
        P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN, 
        P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN, 
        P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN, 
        P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN, 
        P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN, 
        P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN, 
        P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN, 
        P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN, 
        P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN, 
        P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN, 
        P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN, 
        P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, keyinput_f0, 
        keyinput_f1, keyinput_f2, keyinput_f3, keyinput_f4, keyinput_f5, 
        keyinput_f6, keyinput_f7, keyinput_f8, keyinput_f9, keyinput_f10, 
        keyinput_f11, keyinput_f12, keyinput_f13, keyinput_f14, keyinput_f15, 
        keyinput_f16, keyinput_f17, keyinput_f18, keyinput_f19, keyinput_f20, 
        keyinput_f21, keyinput_f22, keyinput_f23, keyinput_f24, keyinput_f25, 
        keyinput_f26, keyinput_f27, keyinput_f28, keyinput_f29, keyinput_f30, 
        keyinput_f31, keyinput_f32, keyinput_f33, keyinput_f34, keyinput_f35, 
        keyinput_f36, keyinput_f37, keyinput_f38, keyinput_f39, keyinput_f40, 
        keyinput_f41, keyinput_f42, keyinput_f43, keyinput_f44, keyinput_f45, 
        keyinput_f46, keyinput_f47, keyinput_f48, keyinput_f49, keyinput_f50, 
        keyinput_f51, keyinput_f52, keyinput_f53, keyinput_f54, keyinput_f55, 
        keyinput_f56, keyinput_f57, keyinput_f58, keyinput_f59, keyinput_f60, 
        keyinput_f61, keyinput_f62, keyinput_f63, keyinput_g0, keyinput_g1, 
        keyinput_g2, keyinput_g3, keyinput_g4, keyinput_g5, keyinput_g6, 
        keyinput_g7, keyinput_g8, keyinput_g9, keyinput_g10, keyinput_g11, 
        keyinput_g12, keyinput_g13, keyinput_g14, keyinput_g15, keyinput_g16, 
        keyinput_g17, keyinput_g18, keyinput_g19, keyinput_g20, keyinput_g21, 
        keyinput_g22, keyinput_g23, keyinput_g24, keyinput_g25, keyinput_g26, 
        keyinput_g27, keyinput_g28, keyinput_g29, keyinput_g30, keyinput_g31, 
        keyinput_g32, keyinput_g33, keyinput_g34, keyinput_g35, keyinput_g36, 
        keyinput_g37, keyinput_g38, keyinput_g39, keyinput_g40, keyinput_g41, 
        keyinput_g42, keyinput_g43, keyinput_g44, keyinput_g45, keyinput_g46, 
        keyinput_g47, keyinput_g48, keyinput_g49, keyinput_g50, keyinput_g51, 
        keyinput_g52, keyinput_g53, keyinput_g54, keyinput_g55, keyinput_g56, 
        keyinput_g57, keyinput_g58, keyinput_g59, keyinput_g60, keyinput_g61, 
        keyinput_g62, keyinput_g63, SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, 
        SUB_1596_U64, SUB_1596_U65, SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, 
        SUB_1596_U69, SUB_1596_U70, SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, 
        SUB_1596_U57, SUB_1596_U58, SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, 
        SUB_1596_U5, SUB_1596_U53, U29, U28, P1_U3355, P1_U3354, P1_U3353, 
        P1_U3352, P1_U3351, P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, 
        P1_U3345, P1_U3344, P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, 
        P1_U3338, P1_U3337, P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, 
        P1_U3331, P1_U3330, P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, 
        P1_U3324, P1_U3445, P1_U3446, P1_U3323, P1_U3322, P1_U3321, P1_U3320, 
        P1_U3319, P1_U3318, P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, 
        P1_U3312, P1_U3311, P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, 
        P1_U3305, P1_U3304, P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, 
        P1_U3298, P1_U3297, P1_U3296, P1_U3295, P1_U3294, P1_U3459, P1_U3462, 
        P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483, 
        P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504, 
        P1_U3507, P1_U3510, P1_U3513, P1_U3515, P1_U3516, P1_U3517, P1_U3518, 
        P1_U3519, P1_U3520, P1_U3521, P1_U3522, P1_U3523, P1_U3524, P1_U3525, 
        P1_U3526, P1_U3527, P1_U3528, P1_U3529, P1_U3530, P1_U3531, P1_U3532, 
        P1_U3533, P1_U3534, P1_U3535, P1_U3536, P1_U3537, P1_U3538, P1_U3539, 
        P1_U3540, P1_U3541, P1_U3542, P1_U3543, P1_U3544, P1_U3545, P1_U3546, 
        P1_U3547, P1_U3548, P1_U3549, P1_U3550, P1_U3551, P1_U3552, P1_U3553, 
        P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3293, 
        P1_U3292, P1_U3291, P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, 
        P1_U3285, P1_U3284, P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, 
        P1_U3278, P1_U3277, P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, 
        P1_U3271, P1_U3270, P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, 
        P1_U3356, P1_U3264, P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, 
        P1_U3258, P1_U3257, P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, 
        P1_U3251, P1_U3250, P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, 
        P1_U3244, P1_U3243, P1_U3560, P1_U3561, P1_U3562, P1_U3563, P1_U3564, 
        P1_U3565, P1_U3566, P1_U3567, P1_U3568, P1_U3569, P1_U3570, P1_U3571, 
        P1_U3572, P1_U3573, P1_U3574, P1_U3575, P1_U3576, P1_U3577, P1_U3578, 
        P1_U3579, P1_U3580, P1_U3581, P1_U3582, P1_U3583, P1_U3584, P1_U3585, 
        P1_U3586, P1_U3587, P1_U3588, P1_U3589, P1_U3590, P1_U3591, P1_U3242, 
        P1_U3241, P1_U3240, P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, 
        P1_U3234, P1_U3233, P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, 
        P1_U3227, P1_U3226, P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, 
        P1_U3220, P1_U3219, P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, 
        P1_U3213, P1_U3086, P1_U3085, P1_U4016, P2_U3327, P2_U3326, P2_U3325, 
        P2_U3324, P2_U3323, P2_U3322, P2_U3321, P2_U3320, P2_U3319, P2_U3318, 
        P2_U3317, P2_U3316, P2_U3315, P2_U3314, P2_U3313, P2_U3312, P2_U3311, 
        P2_U3310, P2_U3309, P2_U3308, P2_U3307, P2_U3306, P2_U3305, P2_U3304, 
        P2_U3303, P2_U3302, P2_U3301, P2_U3300, P2_U3299, P2_U3298, P2_U3297, 
        P2_U3296, P2_U3416, P2_U3417, P2_U3295, P2_U3294, P2_U3293, P2_U3292, 
        P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, 
        P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, 
        P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, 
        P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3430, P2_U3433, 
        P2_U3436, P2_U3439, P2_U3442, P2_U3445, P2_U3448, P2_U3451, P2_U3454, 
        P2_U3457, P2_U3460, P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, 
        P2_U3478, P2_U3481, P2_U3484, P2_U3486, P2_U3487, P2_U3488, P2_U3489, 
        P2_U3490, P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, 
        P2_U3497, P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, 
        P2_U3504, P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, 
        P2_U3511, P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, 
        P2_U3518, P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, 
        P2_U3525, P2_U3526, P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3265, 
        P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258, 
        P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251, 
        P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244, 
        P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, 
        P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, 
        P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, 
        P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, 
        P2_U3215, P2_U3214, P2_U3531, P2_U3532, P2_U3533, P2_U3534, P2_U3535, 
        P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540, P2_U3541, P2_U3542, 
        P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547, P2_U3548, P2_U3549, 
        P2_U3550, P2_U3551, P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, 
        P2_U3557, P2_U3558, P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3328, 
        P2_U3213, P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3208, P2_U3207, 
        P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, 
        P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, 
        P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, 
        P2_U3185, P2_U3088, P2_U3087, P2_U3947, P3_U3295, P3_U3294, P3_U3293, 
        P3_U3292, P3_U3291, P3_U3290, P3_U3289, P3_U3288, P3_U3287, P3_U3286, 
        P3_U3285, P3_U3284, P3_U3283, P3_U3282, P3_U3281, P3_U3280, P3_U3279, 
        P3_U3278, P3_U3277, P3_U3276, P3_U3275, P3_U3274, P3_U3273, P3_U3272, 
        P3_U3271, P3_U3270, P3_U3269, P3_U3268, P3_U3267, P3_U3266, P3_U3265, 
        P3_U3264, P3_U3376, P3_U3377, P3_U3263, P3_U3262, P3_U3261, P3_U3260, 
        P3_U3259, P3_U3258, P3_U3257, P3_U3256, P3_U3255, P3_U3254, P3_U3253, 
        P3_U3252, P3_U3251, P3_U3250, P3_U3249, P3_U3248, P3_U3247, P3_U3246, 
        P3_U3245, P3_U3244, P3_U3243, P3_U3242, P3_U3241, P3_U3240, P3_U3239, 
        P3_U3238, P3_U3237, P3_U3236, P3_U3235, P3_U3234, P3_U3390, P3_U3393, 
        P3_U3396, P3_U3399, P3_U3402, P3_U3405, P3_U3408, P3_U3411, P3_U3414, 
        P3_U3417, P3_U3420, P3_U3423, P3_U3426, P3_U3429, P3_U3432, P3_U3435, 
        P3_U3438, P3_U3441, P3_U3444, P3_U3446, P3_U3447, P3_U3448, P3_U3449, 
        P3_U3450, P3_U3451, P3_U3452, P3_U3453, P3_U3454, P3_U3455, P3_U3456, 
        P3_U3457, P3_U3458, P3_U3459, P3_U3460, P3_U3461, P3_U3462, P3_U3463, 
        P3_U3464, P3_U3465, P3_U3466, P3_U3467, P3_U3468, P3_U3469, P3_U3470, 
        P3_U3471, P3_U3472, P3_U3473, P3_U3474, P3_U3475, P3_U3476, P3_U3477, 
        P3_U3478, P3_U3479, P3_U3480, P3_U3481, P3_U3482, P3_U3483, P3_U3484, 
        P3_U3485, P3_U3486, P3_U3487, P3_U3488, P3_U3489, P3_U3490, P3_U3233, 
        P3_U3232, P3_U3231, P3_U3230, P3_U3229, P3_U3228, P3_U3227, P3_U3226, 
        P3_U3225, P3_U3224, P3_U3223, P3_U3222, P3_U3221, P3_U3220, P3_U3219, 
        P3_U3218, P3_U3217, P3_U3216, P3_U3215, P3_U3214, P3_U3213, P3_U3212, 
        P3_U3211, P3_U3210, P3_U3209, P3_U3208, P3_U3207, P3_U3206, P3_U3205, 
        P3_U3204, P3_U3203, P3_U3202, P3_U3201, P3_U3200, P3_U3199, P3_U3198, 
        P3_U3197, P3_U3196, P3_U3195, P3_U3194, P3_U3193, P3_U3192, P3_U3191, 
        P3_U3190, P3_U3189, P3_U3188, P3_U3187, P3_U3186, P3_U3185, P3_U3184, 
        P3_U3183, P3_U3182, P3_U3491, P3_U3492, P3_U3493, P3_U3494, P3_U3495, 
        P3_U3496, P3_U3497, P3_U3498, P3_U3499, P3_U3500, P3_U3501, P3_U3502, 
        P3_U3503, P3_U3504, P3_U3505, P3_U3506, P3_U3507, P3_U3508, P3_U3509, 
        P3_U3510, P3_U3511, P3_U3512, P3_U3513, P3_U3514, P3_U3515, P3_U3516, 
        P3_U3517, P3_U3518, P3_U3519, P3_U3520, P3_U3521, P3_U3522, P3_U3296, 
        P3_U3181, P3_U3180, P3_U3179, P3_U3178, P3_U3177, P3_U3176, P3_U3175, 
        P3_U3174, P3_U3173, P3_U3172, P3_U3171, P3_U3170, P3_U3169, P3_U3168, 
        P3_U3167, P3_U3166, P3_U3165, P3_U3164, P3_U3163, P3_U3162, P3_U3161, 
        P3_U3160, P3_U3159, P3_U3158, P3_U3157, P3_U3156, P3_U3155, P3_U3154, 
        P3_U3153, P3_U3151, P3_U3150, P3_U3897 );
  input P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN,
         P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN,
         P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN,
         P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN,
         P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN,
         P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN,
         P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN,
         P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN,
         P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN,
         P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN,
         P3_REG3_REG_0__SCAN_IN, P3_REG3_REG_20__SCAN_IN,
         P3_REG3_REG_13__SCAN_IN, P3_REG3_REG_22__SCAN_IN,
         P3_REG3_REG_11__SCAN_IN, P3_REG3_REG_2__SCAN_IN,
         P3_REG3_REG_18__SCAN_IN, P3_REG3_REG_6__SCAN_IN,
         P3_REG3_REG_26__SCAN_IN, P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN,
         P3_DATAO_REG_31__SCAN_IN, P3_DATAO_REG_30__SCAN_IN,
         P3_DATAO_REG_29__SCAN_IN, P3_DATAO_REG_28__SCAN_IN,
         P3_DATAO_REG_27__SCAN_IN, P3_DATAO_REG_26__SCAN_IN,
         P3_DATAO_REG_25__SCAN_IN, P3_DATAO_REG_24__SCAN_IN,
         P3_DATAO_REG_23__SCAN_IN, P3_DATAO_REG_22__SCAN_IN,
         P3_DATAO_REG_21__SCAN_IN, P3_DATAO_REG_20__SCAN_IN,
         P3_DATAO_REG_19__SCAN_IN, P3_DATAO_REG_18__SCAN_IN,
         P3_DATAO_REG_17__SCAN_IN, P3_DATAO_REG_16__SCAN_IN,
         P3_DATAO_REG_15__SCAN_IN, P3_DATAO_REG_14__SCAN_IN,
         P3_DATAO_REG_13__SCAN_IN, P3_DATAO_REG_12__SCAN_IN,
         P3_DATAO_REG_11__SCAN_IN, P3_DATAO_REG_10__SCAN_IN,
         P3_DATAO_REG_9__SCAN_IN, P3_DATAO_REG_8__SCAN_IN,
         P3_DATAO_REG_7__SCAN_IN, P3_DATAO_REG_6__SCAN_IN,
         P3_DATAO_REG_5__SCAN_IN, P3_DATAO_REG_4__SCAN_IN,
         P3_DATAO_REG_3__SCAN_IN, P3_DATAO_REG_2__SCAN_IN,
         P3_DATAO_REG_1__SCAN_IN, P3_DATAO_REG_0__SCAN_IN,
         P3_ADDR_REG_0__SCAN_IN, P3_ADDR_REG_1__SCAN_IN,
         P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN,
         P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN,
         P3_ADDR_REG_6__SCAN_IN, P3_ADDR_REG_7__SCAN_IN,
         P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, P1_IR_REG_0__SCAN_IN,
         P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN,
         P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN,
         P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN,
         P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN,
         P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN,
         P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN,
         P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN,
         P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN,
         P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN,
         P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN,
         P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN,
         P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN,
         P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN,
         P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN,
         P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN,
         P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN,
         P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN,
         P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN,
         P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN,
         P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN,
         P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN,
         P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN,
         P2_RD_REG_SCAN_IN, P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN,
         P3_IR_REG_1__SCAN_IN, P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN,
         P3_IR_REG_4__SCAN_IN, P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN,
         P3_IR_REG_7__SCAN_IN, P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN,
         P3_IR_REG_10__SCAN_IN, P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN,
         P3_IR_REG_13__SCAN_IN, P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN,
         P3_IR_REG_16__SCAN_IN, P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN,
         P3_IR_REG_19__SCAN_IN, P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN,
         P3_IR_REG_22__SCAN_IN, P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN,
         P3_IR_REG_25__SCAN_IN, P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN,
         P3_IR_REG_28__SCAN_IN, P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN,
         P3_IR_REG_31__SCAN_IN, P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN,
         P3_D_REG_2__SCAN_IN, P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN,
         P3_D_REG_5__SCAN_IN, P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN,
         P3_D_REG_8__SCAN_IN, P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN,
         P3_D_REG_11__SCAN_IN, P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN,
         P3_D_REG_14__SCAN_IN, P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN,
         P3_D_REG_17__SCAN_IN, P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN,
         P3_D_REG_20__SCAN_IN, P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN,
         P3_D_REG_23__SCAN_IN, P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN,
         P3_D_REG_26__SCAN_IN, P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN,
         P3_D_REG_29__SCAN_IN, P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN,
         P3_REG0_REG_0__SCAN_IN, P3_REG0_REG_1__SCAN_IN,
         P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN,
         P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN,
         P3_REG0_REG_6__SCAN_IN, P3_REG0_REG_7__SCAN_IN,
         P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN,
         P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN,
         P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN,
         P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN,
         P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN,
         P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN,
         P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN,
         P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN,
         P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN,
         P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN,
         P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN,
         P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN,
         P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN,
         P3_REG1_REG_2__SCAN_IN, P3_REG1_REG_3__SCAN_IN,
         P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN,
         P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN,
         P3_REG1_REG_8__SCAN_IN, P3_REG1_REG_9__SCAN_IN,
         P3_REG1_REG_10__SCAN_IN, P3_REG1_REG_11__SCAN_IN,
         P3_REG1_REG_12__SCAN_IN, P3_REG1_REG_13__SCAN_IN,
         P3_REG1_REG_14__SCAN_IN, P3_REG1_REG_15__SCAN_IN,
         P3_REG1_REG_16__SCAN_IN, P3_REG1_REG_17__SCAN_IN,
         P3_REG1_REG_18__SCAN_IN, P3_REG1_REG_19__SCAN_IN,
         P3_REG1_REG_20__SCAN_IN, P3_REG1_REG_21__SCAN_IN,
         P3_REG1_REG_22__SCAN_IN, P3_REG1_REG_23__SCAN_IN,
         P3_REG1_REG_24__SCAN_IN, P3_REG1_REG_25__SCAN_IN,
         P3_REG1_REG_26__SCAN_IN, P3_REG1_REG_27__SCAN_IN,
         P3_REG1_REG_28__SCAN_IN, P3_REG1_REG_29__SCAN_IN,
         P3_REG1_REG_30__SCAN_IN, P3_REG1_REG_31__SCAN_IN,
         P3_REG2_REG_0__SCAN_IN, P3_REG2_REG_1__SCAN_IN,
         P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN,
         P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN,
         P3_REG2_REG_6__SCAN_IN, P3_REG2_REG_7__SCAN_IN,
         P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN,
         P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN,
         P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN,
         P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN,
         P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN,
         P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN,
         P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN,
         P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN,
         P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN,
         P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN,
         P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN,
         P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN,
         P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN,
         P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN,
         P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN,
         P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN,
         P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, keyinput_f0,
         keyinput_f1, keyinput_f2, keyinput_f3, keyinput_f4, keyinput_f5,
         keyinput_f6, keyinput_f7, keyinput_f8, keyinput_f9, keyinput_f10,
         keyinput_f11, keyinput_f12, keyinput_f13, keyinput_f14, keyinput_f15,
         keyinput_f16, keyinput_f17, keyinput_f18, keyinput_f19, keyinput_f20,
         keyinput_f21, keyinput_f22, keyinput_f23, keyinput_f24, keyinput_f25,
         keyinput_f26, keyinput_f27, keyinput_f28, keyinput_f29, keyinput_f30,
         keyinput_f31, keyinput_f32, keyinput_f33, keyinput_f34, keyinput_f35,
         keyinput_f36, keyinput_f37, keyinput_f38, keyinput_f39, keyinput_f40,
         keyinput_f41, keyinput_f42, keyinput_f43, keyinput_f44, keyinput_f45,
         keyinput_f46, keyinput_f47, keyinput_f48, keyinput_f49, keyinput_f50,
         keyinput_f51, keyinput_f52, keyinput_f53, keyinput_f54, keyinput_f55,
         keyinput_f56, keyinput_f57, keyinput_f58, keyinput_f59, keyinput_f60,
         keyinput_f61, keyinput_f62, keyinput_f63, keyinput_g0, keyinput_g1,
         keyinput_g2, keyinput_g3, keyinput_g4, keyinput_g5, keyinput_g6,
         keyinput_g7, keyinput_g8, keyinput_g9, keyinput_g10, keyinput_g11,
         keyinput_g12, keyinput_g13, keyinput_g14, keyinput_g15, keyinput_g16,
         keyinput_g17, keyinput_g18, keyinput_g19, keyinput_g20, keyinput_g21,
         keyinput_g22, keyinput_g23, keyinput_g24, keyinput_g25, keyinput_g26,
         keyinput_g27, keyinput_g28, keyinput_g29, keyinput_g30, keyinput_g31,
         keyinput_g32, keyinput_g33, keyinput_g34, keyinput_g35, keyinput_g36,
         keyinput_g37, keyinput_g38, keyinput_g39, keyinput_g40, keyinput_g41,
         keyinput_g42, keyinput_g43, keyinput_g44, keyinput_g45, keyinput_g46,
         keyinput_g47, keyinput_g48, keyinput_g49, keyinput_g50, keyinput_g51,
         keyinput_g52, keyinput_g53, keyinput_g54, keyinput_g55, keyinput_g56,
         keyinput_g57, keyinput_g58, keyinput_g59, keyinput_g60, keyinput_g61,
         keyinput_g62, keyinput_g63;
  output SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65,
         SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70,
         SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58,
         SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53,
         U29, U28, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350,
         P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343,
         P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336,
         P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329,
         P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446,
         P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317,
         P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310,
         P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303,
         P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296,
         P1_U3295, P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471,
         P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492,
         P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556,
         P1_U3557, P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290,
         P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283,
         P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276,
         P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269,
         P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263,
         P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256,
         P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249,
         P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588,
         P1_U3589, P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239,
         P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232,
         P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085,
         P1_U4016, P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322,
         P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315,
         P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308,
         P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301,
         P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417,
         P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289,
         P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282,
         P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275,
         P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268,
         P2_U3267, P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442,
         P2_U3445, P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463,
         P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484,
         P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492,
         P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499,
         P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506,
         P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513,
         P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520,
         P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527,
         P2_U3528, P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262,
         P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255,
         P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248,
         P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241,
         P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234,
         P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227,
         P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220,
         P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531,
         P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538,
         P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545,
         P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552,
         P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559,
         P2_U3560, P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204,
         P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197,
         P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190,
         P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087,
         P2_U3947, P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290,
         P3_U3289, P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283,
         P3_U3282, P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276,
         P3_U3275, P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269,
         P3_U3268, P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377,
         P3_U3263, P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257,
         P3_U3256, P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250,
         P3_U3249, P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243,
         P3_U3242, P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236,
         P3_U3235, P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402,
         P3_U3405, P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423,
         P3_U3426, P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444,
         P3_U3446, P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452,
         P3_U3453, P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459,
         P3_U3460, P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466,
         P3_U3467, P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473,
         P3_U3474, P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480,
         P3_U3481, P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487,
         P3_U3488, P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230,
         P3_U3229, P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223,
         P3_U3222, P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216,
         P3_U3215, P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209,
         P3_U3208, P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202,
         P3_U3201, P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195,
         P3_U3194, P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188,
         P3_U3187, P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491,
         P3_U3492, P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498,
         P3_U3499, P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505,
         P3_U3506, P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512,
         P3_U3513, P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519,
         P3_U3520, P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179,
         P3_U3178, P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172,
         P3_U3171, P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165,
         P3_U3164, P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158,
         P3_U3157, P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150,
         P3_U3897;
  wire   n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476,
         n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486,
         n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496,
         n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506,
         n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516,
         n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526,
         n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536,
         n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546,
         n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556,
         n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566,
         n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576,
         n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586,
         n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596,
         n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606,
         n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616,
         n6617, n6618, n6619, n6620, n6622, n6623, n6624, n6625, n6626, n6627,
         n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637,
         n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647,
         n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657,
         n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667,
         n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677,
         n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687,
         n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697,
         n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707,
         n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717,
         n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727,
         n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737,
         n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747,
         n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757,
         n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767,
         n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777,
         n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787,
         n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797,
         n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807,
         n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817,
         n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827,
         n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837,
         n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847,
         n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857,
         n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867,
         n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877,
         n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887,
         n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897,
         n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907,
         n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917,
         n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927,
         n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937,
         n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947,
         n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957,
         n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967,
         n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977,
         n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987,
         n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997,
         n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007,
         n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017,
         n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027,
         n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037,
         n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047,
         n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057,
         n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067,
         n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077,
         n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087,
         n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097,
         n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107,
         n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117,
         n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127,
         n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137,
         n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147,
         n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157,
         n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167,
         n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177,
         n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187,
         n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197,
         n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207,
         n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217,
         n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227,
         n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237,
         n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247,
         n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257,
         n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267,
         n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277,
         n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287,
         n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297,
         n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307,
         n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317,
         n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327,
         n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337,
         n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347,
         n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357,
         n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367,
         n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377,
         n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387,
         n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397,
         n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407,
         n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417,
         n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427,
         n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437,
         n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447,
         n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457,
         n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467,
         n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477,
         n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487,
         n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497,
         n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507,
         n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517,
         n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527,
         n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537,
         n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547,
         n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557,
         n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567,
         n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577,
         n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587,
         n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597,
         n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607,
         n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617,
         n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627,
         n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637,
         n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647,
         n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657,
         n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667,
         n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677,
         n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687,
         n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697,
         n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707,
         n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717,
         n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727,
         n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737,
         n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747,
         n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757,
         n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767,
         n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777,
         n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787,
         n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797,
         n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807,
         n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817,
         n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827,
         n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837,
         n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847,
         n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857,
         n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867,
         n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877,
         n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887,
         n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897,
         n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907,
         n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917,
         n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927,
         n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937,
         n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947,
         n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957,
         n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967,
         n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977,
         n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987,
         n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997,
         n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007,
         n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017,
         n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027,
         n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037,
         n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047,
         n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057,
         n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067,
         n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077,
         n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087,
         n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097,
         n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107,
         n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117,
         n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127,
         n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137,
         n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147,
         n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157,
         n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167,
         n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177,
         n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187,
         n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197,
         n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207,
         n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217,
         n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227,
         n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237,
         n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247,
         n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257,
         n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267,
         n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277,
         n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287,
         n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297,
         n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307,
         n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317,
         n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327,
         n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337,
         n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347,
         n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357,
         n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367,
         n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377,
         n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387,
         n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397,
         n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407,
         n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417,
         n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427,
         n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437,
         n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447,
         n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457,
         n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467,
         n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477,
         n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487,
         n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497,
         n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507,
         n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517,
         n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527,
         n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537,
         n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547,
         n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557,
         n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567,
         n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577,
         n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587,
         n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597,
         n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607,
         n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617,
         n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627,
         n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637,
         n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647,
         n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657,
         n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667,
         n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677,
         n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687,
         n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697,
         n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707,
         n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717,
         n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727,
         n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737,
         n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747,
         n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757,
         n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767,
         n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777,
         n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787,
         n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797,
         n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807,
         n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817,
         n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827,
         n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837,
         n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847,
         n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857,
         n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867,
         n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877,
         n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887,
         n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897,
         n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907,
         n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917,
         n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927,
         n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937,
         n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947,
         n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957,
         n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967,
         n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977,
         n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987,
         n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997,
         n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007,
         n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017,
         n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027,
         n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037,
         n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047,
         n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057,
         n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067,
         n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077,
         n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087,
         n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097,
         n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107,
         n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117,
         n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127,
         n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137,
         n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147,
         n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157,
         n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167,
         n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177,
         n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187,
         n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197,
         n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207,
         n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217,
         n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227,
         n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237,
         n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247,
         n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257,
         n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267,
         n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277,
         n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287,
         n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297,
         n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307,
         n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317,
         n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327,
         n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337,
         n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347,
         n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357,
         n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367,
         n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377,
         n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387,
         n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397,
         n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407,
         n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417,
         n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427,
         n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437,
         n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447,
         n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457,
         n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467,
         n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477,
         n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487,
         n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497,
         n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507,
         n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517,
         n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527,
         n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537,
         n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547,
         n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557,
         n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567,
         n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577,
         n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587,
         n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597,
         n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607,
         n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617,
         n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627,
         n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637,
         n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647,
         n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657,
         n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667,
         n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677,
         n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687,
         n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697,
         n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707,
         n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717,
         n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727,
         n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737,
         n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747,
         n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757,
         n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767,
         n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777,
         n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787,
         n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797,
         n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807,
         n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817,
         n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827,
         n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837,
         n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847,
         n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857,
         n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867,
         n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877,
         n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887,
         n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897,
         n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907,
         n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917,
         n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927,
         n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937,
         n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947,
         n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957,
         n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967,
         n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977,
         n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987,
         n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997,
         n9998, n9999, n10000, n10001, n10002, n10003, n10004, n10005, n10006,
         n10007, n10008, n10009, n10010, n10011, n10012, n10013, n10014,
         n10015, n10016, n10017, n10018, n10019, n10020, n10021, n10022,
         n10023, n10024, n10025, n10026, n10027, n10028, n10029, n10030,
         n10031, n10032, n10033, n10034, n10035, n10036, n10037, n10038,
         n10039, n10040, n10041, n10042, n10043, n10044, n10045, n10046,
         n10047, n10048, n10049, n10050, n10051, n10052, n10053, n10054,
         n10055, n10056, n10057, n10058, n10059, n10060, n10061, n10062,
         n10063, n10064, n10065, n10066, n10067, n10068, n10069, n10070,
         n10071, n10072, n10073, n10074, n10075, n10076, n10077, n10078,
         n10079, n10080, n10081, n10082, n10083, n10084, n10085, n10086,
         n10087, n10088, n10089, n10090, n10091, n10092, n10093, n10094,
         n10095, n10096, n10097, n10098, n10099, n10100, n10101, n10102,
         n10103, n10104, n10105, n10106, n10107, n10108, n10109, n10110,
         n10111, n10112, n10113, n10114, n10115, n10116, n10117, n10118,
         n10119, n10120, n10121, n10122, n10123, n10124, n10125, n10126,
         n10127, n10128, n10129, n10130, n10131, n10132, n10133, n10134,
         n10135, n10136, n10137, n10138, n10139, n10140, n10141, n10142,
         n10143, n10144, n10145, n10146, n10147, n10148, n10149, n10150,
         n10151, n10152, n10153, n10154, n10155, n10156, n10157, n10158,
         n10159, n10160, n10161, n10162, n10163, n10164, n10165, n10166,
         n10167, n10168, n10169, n10170, n10171, n10172, n10173, n10174,
         n10175, n10176, n10177, n10178, n10179, n10180, n10181, n10182,
         n10183, n10184, n10185, n10186, n10187, n10188, n10189, n10190,
         n10191, n10192, n10193, n10194, n10195, n10196, n10197, n10198,
         n10199, n10200, n10201, n10202, n10203, n10204, n10205, n10206,
         n10207, n10208, n10209, n10210, n10211, n10212, n10213, n10214,
         n10215, n10216, n10217, n10218, n10219, n10220, n10221, n10222,
         n10223, n10224, n10225, n10226, n10227, n10228, n10229, n10230,
         n10231, n10232, n10233, n10234, n10235, n10236, n10237, n10238,
         n10239, n10240, n10241, n10242, n10243, n10244, n10245, n10246,
         n10247, n10248, n10249, n10250, n10251, n10252, n10253, n10254,
         n10255, n10256, n10257, n10258, n10259, n10260, n10261, n10262,
         n10263, n10264, n10265, n10266, n10267, n10268, n10269, n10270,
         n10271, n10272, n10273, n10274, n10275, n10276, n10277, n10278,
         n10279, n10280, n10281, n10282, n10283, n10284, n10285, n10286,
         n10287, n10288, n10289, n10290, n10291, n10292, n10293, n10294,
         n10295, n10296, n10297, n10298, n10299, n10300, n10301, n10302,
         n10303, n10304, n10305, n10306, n10307, n10308, n10309, n10310,
         n10311, n10312, n10313, n10314, n10315, n10316, n10317, n10318,
         n10319, n10320, n10321, n10322, n10323, n10324, n10325, n10326,
         n10327, n10328, n10329, n10330, n10331, n10332, n10333, n10334,
         n10335, n10336, n10337, n10338, n10339, n10340, n10341, n10342,
         n10343, n10344, n10345, n10346, n10347, n10348, n10349, n10350,
         n10351, n10352, n10353, n10354, n10355, n10356, n10357, n10358,
         n10359, n10360, n10361, n10362, n10363, n10364, n10365, n10366,
         n10367, n10368, n10369, n10370, n10371, n10372, n10373, n10374,
         n10375, n10376, n10377, n10378, n10379, n10380, n10381, n10382,
         n10383, n10384, n10385, n10386, n10387, n10388, n10389, n10390,
         n10391, n10392, n10393, n10394, n10395, n10396, n10397, n10398,
         n10399, n10400, n10401, n10402, n10403, n10404, n10405, n10406,
         n10407, n10408, n10409, n10410, n10411, n10412, n10413, n10414,
         n10415, n10416, n10417, n10418, n10419, n10420, n10421, n10422,
         n10423, n10424, n10425, n10426, n10427, n10428, n10429, n10430,
         n10431, n10432, n10433, n10434, n10435, n10436, n10437, n10438,
         n10439, n10440, n10441, n10442, n10443, n10444, n10445, n10446,
         n10447, n10448, n10449, n10450, n10451, n10452, n10453, n10454,
         n10455, n10456, n10457, n10458, n10459, n10460, n10461, n10462,
         n10463, n10464, n10465, n10466, n10467, n10468, n10469, n10470,
         n10471, n10472, n10473, n10474, n10475, n10476, n10477, n10478,
         n10479, n10480, n10481, n10482, n10483, n10484, n10485, n10486,
         n10487, n10488, n10489, n10490, n10491, n10492, n10493, n10494,
         n10495, n10496, n10497, n10498, n10499, n10500, n10501, n10502,
         n10503, n10504, n10505, n10506, n10507, n10508, n10509, n10510,
         n10511, n10512, n10513, n10514, n10515, n10516, n10517, n10518,
         n10519, n10520, n10521, n10522, n10523, n10524, n10525, n10526,
         n10527, n10528, n10529, n10530, n10531, n10532, n10533, n10534,
         n10535, n10536, n10537, n10538, n10539, n10540, n10541, n10542,
         n10543, n10544, n10545, n10546, n10547, n10548, n10549, n10550,
         n10551, n10552, n10553, n10554, n10555, n10556, n10557, n10558,
         n10559, n10560, n10561, n10562, n10563, n10564, n10565, n10566,
         n10567, n10568, n10569, n10570, n10571, n10572, n10573, n10574,
         n10575, n10576, n10577, n10578, n10579, n10580, n10581, n10582,
         n10583, n10584, n10585, n10586, n10587, n10588, n10589, n10590,
         n10591, n10592, n10593, n10594, n10595, n10596, n10597, n10598,
         n10599, n10600, n10601, n10602, n10603, n10604, n10605, n10606,
         n10607, n10608, n10609, n10610, n10611, n10612, n10613, n10614,
         n10615, n10616, n10617, n10618, n10619, n10620, n10621, n10622,
         n10623, n10624, n10625, n10626, n10627, n10628, n10629, n10630,
         n10631, n10632, n10633, n10634, n10635, n10636, n10637, n10638,
         n10639, n10640, n10641, n10642, n10643, n10644, n10645, n10646,
         n10647, n10648, n10649, n10650, n10651, n10652, n10653, n10654,
         n10655, n10656, n10657, n10658, n10659, n10660, n10661, n10662,
         n10663, n10664, n10665, n10666, n10667, n10668, n10669, n10670,
         n10671, n10672, n10673, n10674, n10675, n10676, n10677, n10678,
         n10679, n10680, n10681, n10682, n10683, n10684, n10685, n10686,
         n10687, n10688, n10689, n10690, n10691, n10692, n10693, n10694,
         n10695, n10696, n10697, n10698, n10699, n10700, n10701, n10702,
         n10703, n10704, n10705, n10706, n10707, n10708, n10709, n10710,
         n10711, n10712, n10713, n10714, n10715, n10716, n10717, n10718,
         n10719, n10720, n10721, n10722, n10723, n10724, n10725, n10726,
         n10727, n10728, n10729, n10730, n10731, n10732, n10733, n10734,
         n10735, n10736, n10737, n10738, n10739, n10740, n10741, n10742,
         n10743, n10744, n10745, n10746, n10747, n10748, n10749, n10750,
         n10751, n10752, n10753, n10754, n10755, n10756, n10757, n10758,
         n10759, n10760, n10761, n10762, n10763, n10764, n10765, n10766,
         n10767, n10768, n10769, n10770, n10771, n10772, n10773, n10774,
         n10775, n10776, n10777, n10778, n10779, n10780, n10781, n10782,
         n10783, n10784, n10785, n10786, n10787, n10788, n10789, n10790,
         n10791, n10792, n10793, n10794, n10795, n10796, n10797, n10798,
         n10799, n10800, n10801, n10802, n10803, n10804, n10805, n10806,
         n10807, n10808, n10809, n10810, n10811, n10812, n10813, n10814,
         n10815, n10816, n10817, n10818, n10819, n10820, n10821, n10822,
         n10823, n10824, n10825, n10826, n10827, n10828, n10829, n10830,
         n10831, n10832, n10833, n10834, n10835, n10836, n10837, n10838,
         n10839, n10840, n10841, n10842, n10843, n10844, n10845, n10846,
         n10847, n10848, n10849, n10850, n10851, n10852, n10853, n10854,
         n10855, n10856, n10857, n10858, n10859, n10860, n10861, n10862,
         n10863, n10864, n10865, n10866, n10867, n10868, n10869, n10870,
         n10871, n10872, n10873, n10874, n10875, n10876, n10877, n10878,
         n10879, n10880, n10881, n10882, n10883, n10884, n10885, n10886,
         n10887, n10888, n10889, n10890, n10891, n10892, n10893, n10894,
         n10895, n10896, n10897, n10898, n10899, n10900, n10901, n10902,
         n10903, n10904, n10905, n10906, n10907, n10908, n10909, n10910,
         n10911, n10912, n10913, n10914, n10915, n10916, n10917, n10918,
         n10919, n10920, n10921, n10922, n10923, n10924, n10925, n10926,
         n10927, n10928, n10929, n10930, n10931, n10932, n10933, n10934,
         n10935, n10936, n10937, n10938, n10939, n10940, n10941, n10942,
         n10943, n10944, n10945, n10946, n10947, n10948, n10949, n10950,
         n10951, n10952, n10953, n10954, n10955, n10956, n10957, n10958,
         n10959, n10960, n10961, n10962, n10963, n10964, n10965, n10966,
         n10967, n10968, n10969, n10970, n10971, n10972, n10973, n10974,
         n10975, n10976, n10977, n10978, n10979, n10980, n10981, n10982,
         n10983, n10984, n10985, n10986, n10987, n10988, n10989, n10990,
         n10991, n10992, n10993, n10994, n10995, n10996, n10997, n10998,
         n10999, n11000, n11001, n11002, n11003, n11004, n11005, n11006,
         n11007, n11008, n11009, n11010, n11011, n11012, n11013, n11014,
         n11015, n11016, n11017, n11018, n11019, n11020, n11021, n11022,
         n11023, n11024, n11025, n11026, n11027, n11028, n11029, n11030,
         n11031, n11032, n11033, n11034, n11035, n11036, n11037, n11038,
         n11039, n11040, n11041, n11042, n11043, n11044, n11045, n11046,
         n11047, n11048, n11049, n11050, n11051, n11052, n11053, n11054,
         n11055, n11056, n11057, n11058, n11059, n11060, n11061, n11062,
         n11063, n11064, n11065, n11066, n11067, n11068, n11069, n11070,
         n11071, n11072, n11073, n11074, n11075, n11076, n11077, n11078,
         n11079, n11080, n11081, n11082, n11083, n11084, n11085, n11086,
         n11087, n11088, n11089, n11090, n11091, n11092, n11093, n11094,
         n11095, n11096, n11097, n11098, n11099, n11100, n11101, n11102,
         n11103, n11104, n11105, n11106, n11107, n11108, n11109, n11110,
         n11111, n11112, n11113, n11114, n11115, n11116, n11117, n11118,
         n11119, n11120, n11121, n11122, n11123, n11124, n11125, n11126,
         n11127, n11128, n11129, n11130, n11131, n11132, n11133, n11134,
         n11135, n11136, n11137, n11138, n11139, n11140, n11141, n11142,
         n11143, n11144, n11145, n11146, n11147, n11148, n11149, n11150,
         n11151, n11152, n11153, n11154, n11155, n11156, n11157, n11158,
         n11159, n11160, n11161, n11162, n11163, n11164, n11165, n11166,
         n11167, n11168, n11169, n11170, n11171, n11172, n11173, n11174,
         n11175, n11176, n11177, n11178, n11179, n11180, n11181, n11182,
         n11183, n11184, n11185, n11186, n11187, n11188, n11189, n11190,
         n11191, n11192, n11193, n11194, n11195, n11196, n11197, n11198,
         n11199, n11200, n11201, n11202, n11203, n11204, n11205, n11206,
         n11207, n11208, n11209, n11210, n11211, n11212, n11213, n11214,
         n11215, n11216, n11217, n11218, n11219, n11220, n11221, n11222,
         n11223, n11224, n11225, n11226, n11227, n11228, n11229, n11230,
         n11231, n11232, n11233, n11234, n11235, n11236, n11237, n11238,
         n11239, n11240, n11241, n11242, n11243, n11244, n11245, n11246,
         n11247, n11248, n11249, n11250, n11251, n11252, n11253, n11254,
         n11255, n11256, n11257, n11258, n11259, n11260, n11261, n11262,
         n11263, n11264, n11265, n11266, n11267, n11268, n11269, n11270,
         n11271, n11272, n11273, n11274, n11275, n11276, n11277, n11278,
         n11279, n11280, n11281, n11282, n11283, n11284, n11285, n11286,
         n11287, n11288, n11289, n11290, n11291, n11292, n11293, n11294,
         n11295, n11296, n11297, n11298, n11299, n11300, n11301, n11302,
         n11303, n11304, n11305, n11306, n11307, n11308, n11309, n11310,
         n11311, n11312, n11313, n11314, n11315, n11316, n11317, n11318,
         n11319, n11320, n11321, n11322, n11323, n11324, n11325, n11326,
         n11327, n11328, n11329, n11330, n11331, n11332, n11333, n11334,
         n11335, n11336, n11337, n11338, n11339, n11340, n11341, n11342,
         n11343, n11344, n11345, n11346, n11347, n11348, n11349, n11350,
         n11351, n11352, n11353, n11354, n11355, n11356, n11357, n11358,
         n11359, n11360, n11361, n11362, n11363, n11364, n11365, n11366,
         n11367, n11368, n11369, n11370, n11371, n11372, n11373, n11374,
         n11375, n11376, n11377, n11378, n11379, n11380, n11381, n11382,
         n11383, n11384, n11385, n11386, n11387, n11388, n11389, n11390,
         n11391, n11392, n11393, n11394, n11395, n11396, n11397, n11398,
         n11399, n11400, n11401, n11402, n11403, n11404, n11405, n11406,
         n11407, n11408, n11409, n11410, n11411, n11412, n11413, n11414,
         n11415, n11416, n11417, n11418, n11419, n11420, n11421, n11422,
         n11423, n11424, n11425, n11426, n11427, n11428, n11429, n11430,
         n11431, n11432, n11433, n11434, n11435, n11436, n11437, n11438,
         n11439, n11440, n11441, n11442, n11443, n11444, n11445, n11446,
         n11447, n11448, n11449, n11450, n11451, n11452, n11453, n11454,
         n11455, n11456, n11457, n11458, n11459, n11460, n11461, n11462,
         n11463, n11464, n11465, n11466, n11467, n11468, n11469, n11470,
         n11471, n11472, n11473, n11474, n11475, n11476, n11477, n11478,
         n11479, n11480, n11481, n11482, n11483, n11484, n11485, n11486,
         n11487, n11488, n11489, n11490, n11491, n11492, n11493, n11494,
         n11495, n11496, n11497, n11498, n11499, n11500, n11501, n11502,
         n11503, n11504, n11505, n11506, n11507, n11508, n11509, n11510,
         n11511, n11512, n11513, n11514, n11515, n11516, n11517, n11518,
         n11519, n11520, n11521, n11522, n11523, n11524, n11525, n11526,
         n11527, n11528, n11529, n11530, n11531, n11532, n11533, n11534,
         n11535, n11536, n11537, n11538, n11539, n11540, n11541, n11542,
         n11543, n11544, n11545, n11546, n11547, n11548, n11549, n11550,
         n11551, n11552, n11553, n11554, n11555, n11556, n11557, n11558,
         n11559, n11560, n11561, n11562, n11563, n11564, n11565, n11566,
         n11567, n11568, n11569, n11570, n11571, n11572, n11573, n11574,
         n11575, n11576, n11577, n11578, n11579, n11580, n11581, n11582,
         n11583, n11584, n11585, n11586, n11587, n11588, n11589, n11590,
         n11591, n11592, n11593, n11594, n11595, n11596, n11597, n11598,
         n11599, n11600, n11601, n11602, n11603, n11604, n11605, n11606,
         n11607, n11608, n11609, n11610, n11611, n11612, n11613, n11614,
         n11615, n11616, n11617, n11618, n11619, n11620, n11621, n11622,
         n11623, n11624, n11625, n11626, n11627, n11628, n11629, n11630,
         n11631, n11632, n11633, n11634, n11635, n11636, n11637, n11638,
         n11639, n11640, n11641, n11642, n11643, n11644, n11645, n11646,
         n11647, n11648, n11649, n11650, n11651, n11652, n11653, n11654,
         n11655, n11656, n11657, n11658, n11659, n11660, n11661, n11662,
         n11663, n11664, n11665, n11666, n11667, n11669, n11670, n11671,
         n11672, n11673, n11674, n11675, n11676, n11677, n11678, n11679,
         n11680, n11681, n11682, n11683, n11684, n11685, n11686, n11687,
         n11688, n11689, n11690, n11691, n11692, n11693, n11694, n11695,
         n11696, n11697, n11698, n11699, n11700, n11701, n11702, n11703,
         n11704, n11705, n11706, n11707, n11708, n11709, n11710, n11711,
         n11712, n11713, n11714, n11715, n11716, n11717, n11718, n11719,
         n11720, n11721, n11722, n11723, n11724, n11725, n11726, n11727,
         n11728, n11729, n11730, n11731, n11732, n11733, n11734, n11735,
         n11736, n11737, n11738, n11739, n11740, n11741, n11742, n11743,
         n11744, n11745, n11746, n11747, n11748, n11749, n11750, n11751,
         n11752, n11753, n11754, n11755, n11756, n11757, n11758, n11759,
         n11760, n11761, n11762, n11763, n11764, n11765, n11766, n11767,
         n11768, n11769, n11770, n11771, n11772, n11773, n11774, n11775,
         n11776, n11777, n11778, n11779, n11780, n11781, n11782, n11783,
         n11784, n11785, n11786, n11787, n11788, n11789, n11790, n11791,
         n11792, n11793, n11794, n11795, n11796, n11797, n11798, n11799,
         n11800, n11801, n11802, n11803, n11804, n11805, n11806, n11807,
         n11808, n11809, n11810, n11811, n11812, n11813, n11814, n11815,
         n11816, n11817, n11818, n11819, n11820, n11821, n11822, n11823,
         n11824, n11825, n11826, n11827, n11828, n11829, n11830, n11831,
         n11832, n11833, n11834, n11835, n11836, n11837, n11838, n11839,
         n11840, n11841, n11842, n11843, n11844, n11845, n11846, n11847,
         n11848, n11849, n11850, n11851, n11852, n11853, n11854, n11855,
         n11856, n11857, n11858, n11859, n11860, n11861, n11862, n11863,
         n11864, n11865, n11866, n11867, n11868, n11869, n11870, n11871,
         n11872, n11873, n11874, n11875, n11876, n11877, n11878, n11879,
         n11880, n11881, n11882, n11883, n11884, n11885, n11886, n11887,
         n11888, n11889, n11890, n11891, n11892, n11893, n11894, n11895,
         n11896, n11897, n11898, n11899, n11900, n11901, n11902, n11903,
         n11904, n11905, n11906, n11907, n11908, n11909, n11910, n11911,
         n11912, n11913, n11914, n11915, n11916, n11917, n11918, n11919,
         n11920, n11921, n11922, n11923, n11924, n11925, n11926, n11927,
         n11928, n11929, n11930, n11931, n11932, n11933, n11934, n11935,
         n11936, n11937, n11938, n11939, n11940, n11941, n11942, n11943,
         n11944, n11945, n11946, n11947, n11948, n11949, n11950, n11951,
         n11952, n11953, n11954, n11955, n11956, n11957, n11958, n11959,
         n11960, n11961, n11962, n11963, n11964, n11965, n11966, n11967,
         n11968, n11969, n11970, n11971, n11972, n11973, n11974, n11975,
         n11976, n11977, n11978, n11979, n11980, n11981, n11982, n11983,
         n11984, n11985, n11986, n11987, n11988, n11989, n11990, n11991,
         n11992, n11993, n11994, n11995, n11996, n11997, n11998, n11999,
         n12000, n12001, n12002, n12003, n12004, n12005, n12006, n12007,
         n12008, n12009, n12010, n12011, n12012, n12013, n12014, n12015,
         n12016, n12017, n12018, n12019, n12020, n12021, n12022, n12023,
         n12024, n12025, n12026, n12027, n12028, n12029, n12030, n12031,
         n12032, n12033, n12034, n12035, n12036, n12037, n12038, n12039,
         n12040, n12041, n12042, n12043, n12044, n12045, n12046, n12047,
         n12048, n12049, n12050, n12051, n12052, n12053, n12054, n12055,
         n12056, n12057, n12058, n12059, n12060, n12061, n12062, n12063,
         n12064, n12065, n12066, n12067, n12068, n12069, n12070, n12071,
         n12072, n12073, n12074, n12075, n12076, n12077, n12078, n12079,
         n12080, n12081, n12082, n12083, n12084, n12085, n12086, n12087,
         n12088, n12089, n12090, n12091, n12092, n12093, n12094, n12095,
         n12096, n12097, n12098, n12099, n12100, n12101, n12102, n12103,
         n12104, n12105, n12106, n12107, n12108, n12109, n12110, n12111,
         n12112, n12113, n12114, n12115, n12116, n12117, n12118, n12119,
         n12120, n12121, n12122, n12123, n12124, n12125, n12126, n12127,
         n12128, n12129, n12130, n12131, n12132, n12133, n12134, n12135,
         n12136, n12137, n12138, n12139, n12140, n12141, n12142, n12143,
         n12144, n12145, n12146, n12147, n12148, n12150, n12151, n12152,
         n12153, n12154, n12155, n12156, n12157, n12158, n12159, n12160,
         n12161, n12162, n12163, n12164, n12165, n12166, n12167, n12168,
         n12169, n12170, n12171, n12172, n12173, n12174, n12175, n12176,
         n12177, n12178, n12179, n12180, n12181, n12182, n12183, n12184,
         n12185, n12186, n12187, n12188, n12189, n12190, n12191, n12192,
         n12193, n12194, n12195, n12196, n12197, n12198, n12199, n12200,
         n12201, n12202, n12203, n12204, n12205, n12206, n12207, n12208,
         n12209, n12210, n12211, n12212, n12213, n12214, n12215, n12216,
         n12217, n12218, n12219, n12220, n12221, n12222, n12223, n12224,
         n12225, n12226, n12227, n12228, n12229, n12230, n12231, n12232,
         n12233, n12234, n12235, n12236, n12237, n12238, n12239, n12240,
         n12241, n12242, n12243, n12244, n12245, n12246, n12247, n12248,
         n12249, n12250, n12251, n12252, n12253, n12254, n12255, n12256,
         n12257, n12258, n12259, n12260, n12261, n12262, n12263, n12264,
         n12265, n12266, n12267, n12268, n12269, n12270, n12271, n12272,
         n12273, n12274, n12275, n12276, n12277, n12278, n12279, n12280,
         n12281, n12282, n12283, n12284, n12285, n12286, n12287, n12288,
         n12289, n12290, n12291, n12292, n12293, n12294, n12295, n12296,
         n12297, n12298, n12299, n12300, n12301, n12302, n12303, n12304,
         n12305, n12306, n12307, n12308, n12309, n12310, n12311, n12312,
         n12313, n12314, n12315, n12316, n12317, n12318, n12319, n12320,
         n12321, n12322, n12323, n12324, n12325, n12326, n12327, n12328,
         n12329, n12330, n12331, n12332, n12333, n12334, n12335, n12336,
         n12337, n12338, n12339, n12340, n12341, n12342, n12343, n12344,
         n12345, n12346, n12347, n12348, n12349, n12350, n12351, n12352,
         n12353, n12354, n12355, n12356, n12357, n12358, n12359, n12360,
         n12361, n12362, n12363, n12364, n12365, n12366, n12367, n12368,
         n12369, n12370, n12371, n12372, n12373, n12374, n12375, n12376,
         n12377, n12378, n12379, n12380, n12381, n12382, n12383, n12384,
         n12385, n12386, n12387, n12388, n12389, n12390, n12391, n12392,
         n12393, n12394, n12395, n12396, n12397, n12398, n12399, n12400,
         n12401, n12402, n12403, n12404, n12405, n12406, n12407, n12408,
         n12409, n12410, n12411, n12412, n12413, n12414, n12415, n12416,
         n12417, n12418, n12419, n12420, n12421, n12422, n12423, n12424,
         n12425, n12426, n12427, n12428, n12429, n12430, n12431, n12432,
         n12433, n12434, n12435, n12436, n12437, n12438, n12439, n12440,
         n12441, n12442, n12443, n12444, n12445, n12446, n12447, n12448,
         n12449, n12450, n12451, n12452, n12453, n12454, n12455, n12456,
         n12457, n12458, n12459, n12460, n12461, n12462, n12463, n12464,
         n12465, n12466, n12467, n12468, n12469, n12470, n12471, n12472,
         n12473, n12474, n12475, n12476, n12477, n12478, n12479, n12480,
         n12481, n12482, n12483, n12484, n12485, n12486, n12487, n12488,
         n12489, n12490, n12491, n12492, n12493, n12494, n12495, n12496,
         n12497, n12498, n12499, n12500, n12501, n12502, n12503, n12504,
         n12505, n12506, n12507, n12508, n12509, n12510, n12511, n12512,
         n12513, n12514, n12515, n12516, n12517, n12518, n12519, n12520,
         n12521, n12522, n12523, n12524, n12525, n12526, n12527, n12528,
         n12529, n12530, n12531, n12532, n12533, n12534, n12535, n12536,
         n12537, n12538, n12539, n12540, n12541, n12542, n12543, n12544,
         n12545, n12546, n12547, n12548, n12549, n12550, n12551, n12552,
         n12553, n12554, n12555, n12556, n12557, n12558, n12559, n12560,
         n12561, n12562, n12563, n12564, n12565, n12566, n12567, n12568,
         n12569, n12570, n12571, n12572, n12573, n12574, n12575, n12576,
         n12577, n12578, n12579, n12580, n12581, n12582, n12583, n12584,
         n12585, n12586, n12587, n12588, n12589, n12590, n12591, n12592,
         n12593, n12594, n12595, n12596, n12597, n12598, n12599, n12600,
         n12601, n12602, n12603, n12604, n12605, n12606, n12607, n12608,
         n12609, n12610, n12611, n12612, n12613, n12614, n12615, n12616,
         n12617, n12618, n12619, n12620, n12621, n12622, n12623, n12624,
         n12625, n12626, n12627, n12628, n12629, n12630, n12631, n12632,
         n12633, n12634, n12635, n12636, n12637, n12638, n12639, n12640,
         n12641, n12642, n12643, n12644, n12645, n12646, n12647, n12648,
         n12649, n12650, n12651, n12652, n12653, n12654, n12655, n12656,
         n12657, n12658, n12659, n12660, n12661, n12662, n12663, n12664,
         n12665, n12666, n12667, n12668, n12669, n12670, n12671, n12672,
         n12673, n12674, n12675, n12676, n12677, n12678, n12679, n12680,
         n12681, n12682, n12683, n12684, n12685, n12686, n12687, n12688,
         n12689, n12690, n12691, n12692, n12693, n12694, n12695, n12696,
         n12697, n12698, n12699, n12700, n12701, n12702, n12703, n12704,
         n12705, n12706, n12707, n12708, n12709, n12710, n12711, n12712,
         n12713, n12714, n12715, n12716, n12717, n12718, n12719, n12720,
         n12721, n12722, n12723, n12724, n12725, n12726, n12727, n12728,
         n12729, n12730, n12731, n12732, n12733, n12734, n12735, n12736,
         n12737, n12738, n12739, n12740, n12741, n12742, n12743, n12744,
         n12745, n12746, n12747, n12748, n12749, n12750, n12751, n12752,
         n12753, n12754, n12755, n12756, n12757, n12758, n12759, n12760,
         n12761, n12762, n12763, n12764, n12765, n12766, n12767, n12768,
         n12769, n12770, n12771, n12772, n12773, n12774, n12775, n12776,
         n12777, n12778, n12779, n12780, n12781, n12782, n12783, n12784,
         n12785, n12786, n12787, n12788, n12789, n12790, n12791, n12792,
         n12793, n12794, n12795, n12796, n12797, n12798, n12799, n12800,
         n12801, n12802, n12803, n12804, n12805, n12806, n12807, n12808,
         n12809, n12810, n12811, n12812, n12813, n12814, n12815, n12816,
         n12817, n12818, n12819, n12820, n12821, n12822, n12823, n12824,
         n12825, n12826, n12827, n12828, n12829, n12830, n12831, n12832,
         n12833, n12834, n12835, n12836, n12837, n12838, n12839, n12840,
         n12841, n12842, n12843, n12844, n12845, n12846, n12847, n12848,
         n12849, n12850, n12851, n12852, n12853, n12854, n12855, n12856,
         n12857, n12858, n12859, n12860, n12861, n12862, n12863, n12864,
         n12865, n12866, n12867, n12868, n12869, n12870, n12871, n12872,
         n12873, n12874, n12875, n12876, n12877, n12878, n12879, n12880,
         n12881, n12882, n12883, n12884, n12885, n12886, n12887, n12888,
         n12889, n12890, n12891, n12892, n12893, n12894, n12895, n12896,
         n12897, n12898, n12899, n12900, n12901, n12902, n12903, n12904,
         n12905, n12906, n12907, n12908, n12909, n12910, n12911, n12912,
         n12913, n12914, n12915, n12916, n12917, n12918, n12919, n12920,
         n12921, n12922, n12923, n12924, n12925, n12926, n12927, n12928,
         n12929, n12930, n12931, n12932, n12933, n12934, n12935, n12936,
         n12937, n12938, n12939, n12940, n12941, n12942, n12943, n12944,
         n12945, n12946, n12947, n12948, n12949, n12950, n12951, n12952,
         n12953, n12954, n12955, n12956, n12957, n12958, n12959, n12960,
         n12961, n12962, n12963, n12964, n12965, n12966, n12967, n12968,
         n12969, n12970, n12971, n12972, n12973, n12974, n12975, n12976,
         n12977, n12978, n12979, n12980, n12981, n12982, n12983, n12984,
         n12985, n12986, n12987, n12988, n12989, n12990, n12991, n12992,
         n12993, n12994, n12995, n12996, n12997, n12998, n12999, n13000,
         n13001, n13002, n13003, n13004, n13005, n13006, n13007, n13008,
         n13009, n13010, n13011, n13012, n13013, n13014, n13015, n13016,
         n13017, n13018, n13019, n13020, n13021, n13022, n13023, n13024,
         n13025, n13026, n13027, n13028, n13029, n13030, n13031, n13032,
         n13033, n13034, n13035, n13036, n13037, n13038, n13039, n13040,
         n13041, n13042, n13043, n13044, n13045, n13046, n13047, n13048,
         n13049, n13050, n13051, n13052, n13053, n13054, n13055, n13056,
         n13057, n13058, n13059, n13060, n13061, n13062, n13063, n13064,
         n13065, n13066, n13067, n13068, n13069, n13070, n13071, n13072,
         n13073, n13074, n13075, n13076, n13077, n13078, n13079, n13080,
         n13081, n13082, n13083, n13084, n13085, n13086, n13087, n13088,
         n13089, n13090, n13091, n13092, n13093, n13094, n13095, n13096,
         n13097, n13098, n13099, n13100, n13101, n13102, n13103, n13104,
         n13105, n13106, n13107, n13108, n13109, n13110, n13111, n13112,
         n13113, n13114, n13115, n13116, n13117, n13118, n13119, n13120,
         n13121, n13122, n13123, n13124, n13125, n13126, n13127, n13128,
         n13129, n13130, n13131, n13132, n13133, n13134, n13135, n13136,
         n13137, n13138, n13139, n13140, n13141, n13142, n13143, n13144,
         n13145, n13146, n13147, n13148, n13149, n13150, n13151, n13152,
         n13153, n13154, n13155, n13156, n13157, n13158, n13159, n13160,
         n13161, n13162, n13163, n13164, n13165, n13166, n13167, n13168,
         n13169, n13170, n13171, n13172, n13173, n13174, n13175, n13176,
         n13177, n13178, n13179, n13180, n13181, n13182, n13183, n13184,
         n13185, n13186, n13187, n13188, n13189, n13190, n13191, n13192,
         n13193, n13194, n13195, n13196, n13197, n13198, n13199, n13200,
         n13201, n13202, n13203, n13204, n13205, n13206, n13207, n13208,
         n13209, n13210, n13211, n13212, n13213, n13214, n13215, n13216,
         n13217, n13218, n13219, n13220, n13221, n13222, n13223, n13224,
         n13225, n13226, n13227, n13228, n13229, n13230, n13231, n13232,
         n13233, n13234, n13235, n13236, n13237, n13238, n13239, n13240,
         n13241, n13242, n13243, n13244, n13245, n13246, n13247, n13248,
         n13249, n13250, n13251, n13252, n13253, n13254, n13255, n13256,
         n13257, n13258, n13259, n13260, n13261, n13262, n13263, n13264,
         n13265, n13266, n13267, n13268, n13269, n13270, n13271, n13272,
         n13273, n13274, n13275, n13276, n13277, n13278, n13279, n13280,
         n13281, n13282, n13283, n13284, n13285, n13286, n13287, n13288,
         n13289, n13290, n13291, n13292, n13293, n13294, n13295, n13296,
         n13297, n13298, n13299, n13300, n13301, n13302, n13303, n13304,
         n13305, n13306, n13307, n13308, n13309, n13310, n13311, n13312,
         n13313, n13314, n13315, n13316, n13317, n13318, n13319, n13320,
         n13321, n13322, n13323, n13324, n13325, n13326, n13327, n13328,
         n13329, n13330, n13331, n13332, n13333, n13334, n13335, n13336,
         n13337, n13338, n13339, n13340, n13341, n13342, n13343, n13344,
         n13345, n13346, n13347, n13348, n13349, n13350, n13351, n13352,
         n13353, n13354, n13355, n13356, n13357, n13358, n13359, n13360,
         n13361, n13362, n13363, n13364, n13365, n13366, n13367, n13368,
         n13369, n13370, n13371, n13372, n13373, n13374, n13375, n13376,
         n13377, n13378, n13379, n13380, n13381, n13382, n13383, n13384,
         n13385, n13386, n13387, n13388, n13389, n13390, n13391, n13392,
         n13393, n13394, n13395, n13396, n13397, n13398, n13399, n13400,
         n13401, n13402, n13403, n13404, n13405, n13406, n13407, n13408,
         n13409, n13410, n13411, n13412, n13413, n13414, n13415, n13416,
         n13417, n13418, n13419, n13420, n13421, n13422, n13423, n13424,
         n13425, n13426, n13427, n13428, n13429, n13430, n13431, n13432,
         n13433, n13434, n13435, n13436, n13437, n13438, n13439, n13440,
         n13441, n13442, n13443, n13444, n13445, n13446, n13447, n13448,
         n13449, n13450, n13451, n13452, n13453, n13454, n13455, n13456,
         n13457, n13458, n13459, n13460, n13461, n13462, n13463, n13464,
         n13465, n13466, n13467, n13468, n13469, n13470, n13471, n13472,
         n13473, n13474, n13475, n13476, n13477, n13478, n13479, n13480,
         n13481, n13482, n13483, n13484, n13485, n13486, n13487, n13488,
         n13489, n13490, n13491, n13492, n13493, n13494, n13495, n13496,
         n13497, n13498, n13499, n13500, n13501, n13502, n13503, n13504,
         n13505, n13506, n13507, n13508, n13509, n13510, n13511, n13512,
         n13513, n13514, n13515, n13516, n13517, n13518, n13519, n13520,
         n13521, n13522, n13523, n13524, n13525, n13526, n13527, n13528,
         n13529, n13530, n13531, n13532, n13533, n13534, n13535, n13536,
         n13537, n13538, n13539, n13540, n13541, n13542, n13543, n13544,
         n13545, n13546, n13547, n13548, n13549, n13550, n13551, n13552,
         n13553, n13554, n13555, n13556, n13557, n13558, n13559, n13560,
         n13561, n13562, n13563, n13564, n13565, n13566, n13567, n13568,
         n13569, n13570, n13571, n13572, n13573, n13574, n13575, n13576,
         n13577, n13578, n13579, n13580, n13581, n13582, n13583, n13584,
         n13585, n13586, n13587, n13588, n13589, n13590, n13591, n13592,
         n13593, n13594, n13595, n13596, n13597, n13598, n13599, n13600,
         n13601, n13602, n13603, n13604, n13605, n13606, n13607, n13608,
         n13609, n13610, n13611, n13612, n13613, n13614, n13615, n13616,
         n13617, n13618, n13619, n13620, n13621, n13622, n13623, n13624,
         n13625, n13626, n13627, n13628, n13629, n13630, n13631, n13632,
         n13633, n13634, n13635, n13636, n13637, n13638, n13639, n13640,
         n13641, n13642, n13643, n13644, n13645, n13646, n13647, n13648,
         n13649, n13650, n13651, n13652, n13653, n13654, n13655, n13656,
         n13657, n13658, n13659, n13660, n13661, n13662, n13663, n13664,
         n13665, n13666, n13667, n13668, n13669, n13670, n13671, n13672,
         n13673, n13674, n13675, n13676, n13677, n13678, n13679, n13680,
         n13681, n13682, n13683, n13684, n13685, n13686, n13687, n13688,
         n13689, n13690, n13691, n13692, n13693, n13694, n13695, n13696,
         n13697, n13698, n13699, n13700, n13701, n13702, n13703, n13704,
         n13705, n13706, n13707, n13708, n13709, n13710, n13711, n13712,
         n13713, n13714, n13715, n13716, n13717, n13718, n13719, n13720,
         n13721, n13722, n13723, n13724, n13725, n13726, n13727, n13728,
         n13729, n13730, n13731, n13732, n13733, n13734, n13735, n13736,
         n13737, n13738, n13739, n13740, n13741, n13742, n13743, n13744,
         n13745, n13746, n13747, n13748, n13749, n13750, n13751, n13752,
         n13753, n13754, n13755, n13756, n13757, n13758, n13759, n13760,
         n13761, n13762, n13763, n13764, n13765, n13766, n13767, n13768,
         n13769, n13770, n13771, n13772, n13773, n13774, n13775, n13776,
         n13777, n13778, n13779, n13780, n13781, n13782, n13783, n13784,
         n13785, n13786, n13787, n13788, n13789, n13790, n13791, n13792,
         n13793, n13794, n13795, n13796, n13797, n13798, n13799, n13800,
         n13801, n13802, n13803, n13804, n13805, n13806, n13807, n13808,
         n13809, n13810, n13811, n13812, n13813, n13814, n13815, n13816,
         n13817, n13818, n13819, n13820, n13821, n13822, n13823, n13824,
         n13825, n13826, n13827, n13828, n13829, n13830, n13831, n13832,
         n13833, n13834, n13835, n13836, n13837, n13838, n13839, n13840,
         n13841, n13842, n13843, n13844, n13845, n13846, n13847, n13848,
         n13849, n13850, n13851, n13852, n13853, n13854, n13855, n13856,
         n13857, n13858, n13859, n13860, n13861, n13862, n13863, n13864,
         n13865, n13866, n13867, n13868, n13869, n13870, n13871, n13872,
         n13873, n13874, n13875, n13876, n13877, n13878, n13879, n13880,
         n13881, n13882, n13883, n13884, n13885, n13886, n13887, n13888,
         n13889, n13890, n13891, n13892, n13893, n13894, n13895, n13896,
         n13897, n13898, n13899, n13900, n13901, n13902, n13903, n13904,
         n13905, n13906, n13907, n13908, n13909, n13910, n13911, n13912,
         n13913, n13914, n13915, n13916, n13917, n13918, n13919, n13920,
         n13921, n13922, n13923, n13924, n13925, n13926, n13927, n13928,
         n13929, n13930, n13931, n13932, n13933, n13934, n13935, n13936,
         n13937, n13938, n13939, n13940, n13941, n13942, n13943, n13944,
         n13945, n13946, n13947, n13948, n13949, n13950, n13951, n13952,
         n13953, n13954, n13955, n13956, n13957, n13958, n13959, n13960,
         n13961, n13962, n13963, n13964, n13965, n13966, n13967, n13968,
         n13969, n13970, n13971, n13972, n13973, n13974, n13975, n13976,
         n13977, n13978, n13979, n13980, n13981, n13982, n13983, n13984,
         n13985, n13986, n13987, n13988, n13989, n13990, n13991, n13992,
         n13993, n13994, n13995, n13996, n13997, n13998, n13999, n14000,
         n14001, n14002, n14003, n14004, n14005, n14006, n14007, n14008,
         n14009, n14010, n14011, n14012, n14013, n14014, n14015, n14016,
         n14017, n14018, n14019, n14020, n14021, n14022, n14023, n14024,
         n14025, n14026, n14027, n14028, n14029, n14030, n14031, n14032,
         n14033, n14034, n14035, n14036, n14037, n14038, n14039, n14040,
         n14041, n14042, n14043, n14044, n14045, n14046, n14047, n14048,
         n14049, n14050, n14051, n14052, n14053, n14054, n14055, n14056,
         n14057, n14058, n14059, n14060, n14061, n14062, n14063, n14064,
         n14065, n14066, n14067, n14068, n14069, n14070, n14071, n14072,
         n14073, n14074, n14075, n14076, n14077, n14078, n14079, n14080,
         n14081, n14082, n14083, n14084, n14085, n14086, n14087, n14088,
         n14089, n14090, n14091, n14092, n14093, n14094, n14095, n14096,
         n14097, n14098, n14099, n14100, n14101, n14102, n14103, n14104,
         n14105, n14106, n14107, n14108, n14109, n14110, n14111, n14112,
         n14113, n14114, n14115, n14116, n14117, n14118, n14119, n14120,
         n14121, n14122, n14123, n14124, n14125, n14126, n14127, n14128,
         n14129, n14130, n14131, n14132, n14133, n14134, n14135, n14136,
         n14137, n14138, n14139, n14140, n14141, n14142, n14143, n14144,
         n14145, n14146, n14147, n14148, n14149, n14150, n14151, n14152,
         n14153, n14154, n14155, n14156, n14157, n14158, n14159, n14160,
         n14161, n14162, n14163, n14164, n14165, n14166, n14167, n14168,
         n14169, n14170, n14171, n14172, n14173, n14174, n14175, n14176,
         n14177, n14178, n14179, n14180, n14181, n14182, n14183, n14184,
         n14185, n14186, n14187, n14188, n14189, n14190, n14191, n14192,
         n14193, n14194, n14195, n14196, n14197, n14198, n14199, n14200,
         n14201, n14202, n14203, n14204, n14205, n14206, n14207, n14208,
         n14209, n14210, n14211, n14212, n14213, n14214, n14215, n14216,
         n14217, n14218, n14219, n14220, n14221, n14222, n14223, n14224,
         n14225, n14226, n14227, n14228, n14229, n14230, n14231, n14232,
         n14233, n14234, n14235, n14236, n14237, n14238, n14239, n14240,
         n14241, n14242, n14243, n14244, n14245, n14246, n14247, n14248,
         n14249, n14250, n14251, n14252, n14253, n14254, n14255, n14256,
         n14257, n14258, n14259, n14260, n14261, n14262, n14263, n14264,
         n14265, n14266, n14267, n14268, n14269, n14270, n14271, n14272,
         n14273, n14274, n14275, n14276, n14277, n14278, n14279, n14280,
         n14281, n14282, n14283, n14284, n14285, n14286, n14287, n14288,
         n14289, n14290, n14291, n14292, n14293, n14294, n14295, n14296,
         n14297, n14298, n14299, n14300, n14301, n14302, n14303, n14304,
         n14305, n14306, n14307, n14308, n14309, n14310, n14311, n14312,
         n14313, n14314, n14315, n14316, n14317, n14318, n14319, n14320,
         n14321, n14322, n14323, n14324, n14325, n14326, n14327, n14328,
         n14329, n14330, n14331, n14332, n14333, n14334, n14335, n14336,
         n14337, n14338, n14339, n14340, n14341, n14342, n14343, n14344,
         n14345, n14346, n14347, n14348, n14349, n14350, n14351, n14352,
         n14353, n14354, n14355, n14356, n14357, n14358, n14359, n14360,
         n14361, n14362, n14363, n14364, n14365, n14366, n14367, n14368,
         n14369, n14370, n14371, n14372, n14373, n14374, n14375, n14376,
         n14377, n14378, n14379, n14380, n14381, n14382, n14383, n14384,
         n14385, n14386, n14387, n14388, n14389, n14390, n14391, n14392,
         n14393, n14394, n14395, n14396, n14397, n14398, n14399, n14400,
         n14401, n14402, n14403, n14404, n14405, n14406, n14407, n14408,
         n14409, n14410, n14411, n14412, n14413, n14414, n14415, n14416,
         n14417, n14418, n14419, n14420, n14421, n14422, n14423, n14424,
         n14425, n14426, n14427, n14428, n14429, n14430, n14431, n14432,
         n14433, n14434, n14435, n14436, n14437, n14438, n14439, n14440,
         n14441, n14442, n14443, n14444, n14445, n14446, n14447, n14448,
         n14449, n14450, n14451, n14452, n14453, n14454, n14455, n14456,
         n14457, n14458, n14459, n14460, n14461, n14462, n14463, n14464,
         n14465, n14466, n14467, n14468, n14469, n14470, n14471, n14472,
         n14473, n14474, n14475, n14476, n14477, n14478, n14479, n14480,
         n14481, n14482, n14483, n14484, n14485, n14486, n14487, n14488,
         n14489, n14490, n14491, n14492, n14493, n14494, n14495, n14496,
         n14497, n14498, n14499, n14500, n14501, n14502, n14503, n14504,
         n14505, n14506, n14507, n14508, n14509, n14510, n14511, n14512,
         n14513, n14514, n14515, n14516, n14517, n14518, n14519, n14520,
         n14521, n14522, n14523, n14524, n14525, n14526, n14527, n14528,
         n14529, n14530, n14531, n14532, n14533, n14534, n14535, n14536,
         n14537, n14538, n14539, n14540, n14541, n14542, n14543, n14544,
         n14545, n14546, n14547, n14548, n14549, n14550, n14551, n14552,
         n14553, n14554, n14555, n14556, n14557, n14558, n14559, n14560,
         n14561, n14562, n14563, n14564, n14565, n14566, n14567, n14568,
         n14569, n14570, n14571, n14572, n14573, n14574, n14575, n14576,
         n14577, n14578, n14579, n14580, n14581, n14582, n14583, n14584,
         n14585, n14586, n14587, n14588, n14589, n14590, n14591, n14592,
         n14593, n14594, n14595, n14596, n14597, n14598, n14599, n14600,
         n14601, n14602, n14603, n14604, n14605, n14606, n14607, n14608,
         n14609, n14610, n14611, n14612, n14613, n14614, n14615, n14616,
         n14617, n14618, n14619, n14620, n14621, n14622, n14623, n14624,
         n14625, n14626, n14627, n14628, n14629, n14630, n14631, n14632,
         n14633, n14634, n14635, n14636, n14637, n14638, n14639, n14640,
         n14641, n14642, n14643, n14644, n14645, n14646, n14647, n14648,
         n14649, n14650, n14651, n14652, n14653, n14654, n14655, n14656,
         n14657, n14658, n14659, n14660, n14661, n14662, n14663, n14664,
         n14665, n14666, n14667, n14668, n14669, n14670, n14671, n14672,
         n14673, n14674, n14675, n14676, n14677, n14678, n14679, n14680,
         n14681, n14682, n14683, n14684, n14685, n14686, n14687, n14688,
         n14689, n14690, n14691, n14692, n14693, n14694, n14695, n14696,
         n14697, n14698, n14699, n14700, n14701, n14702, n14703, n14704,
         n14705, n14706, n14707, n14708, n14709, n14710, n14711, n14712,
         n14713, n14714, n14715, n14716, n14717, n14718, n14719, n14720,
         n14721, n14722, n14723, n14724, n14725, n14726, n14727, n14728,
         n14729, n14730, n14731, n14732, n14733, n14734, n14735, n14736,
         n14737, n14738, n14739, n14740, n14741, n14742, n14743, n14744,
         n14745, n14746, n14747, n14748, n14749, n14750, n14751, n14752,
         n14753, n14754, n14755, n14756, n14757, n14758, n14759, n14760,
         n14761, n14762, n14763, n14764, n14765, n14766, n14767, n14768,
         n14769, n14770, n14771, n14772, n14773, n14774, n14775, n14776,
         n14777, n14778, n14779, n14780, n14781, n14782, n14783, n14784,
         n14785, n14786, n14787, n14788, n14789, n14790, n14791, n14792,
         n14793, n14794, n14795, n14796, n14797, n14798, n14799, n14800,
         n14801, n14802, n14803, n14804, n14805, n14806, n14807, n14808,
         n14809, n14810, n14811, n14812, n14813, n14814, n14815, n14816,
         n14817, n14818, n14819, n14820, n14821, n14822, n14823, n14824,
         n14825, n14826, n14827, n14828, n14829, n14830, n14831, n14832,
         n14833, n14834, n14835, n14836, n14837, n14838, n14839, n14840,
         n14841, n14842, n14843, n14844, n14845, n14846, n14847, n14848,
         n14849, n14850, n14851, n14852, n14853, n14854, n14855, n14856,
         n14857, n14858, n14859, n14860, n14861, n14862, n14863, n14864,
         n14865, n14866, n14867, n14868, n14869, n14870, n14871, n14872,
         n14873, n14874, n14875, n14876, n14877, n14878, n14879, n14880,
         n14881, n14882, n14883, n14884, n14885, n14886, n14887, n14888,
         n14889, n14890, n14891, n14892, n14893, n14894, n14895, n14896,
         n14897, n14898, n14899, n14900, n14901, n14902, n14903, n14904,
         n14905, n14906, n14907, n14908, n14909, n14910, n14911, n14912,
         n14913, n14914, n14915, n14916, n14917, n14918, n14919, n14920,
         n14921, n14922, n14923, n14924, n14925, n14926, n14927, n14928,
         n14929, n14930, n14931, n14932, n14933, n14934, n14935, n14936,
         n14937, n14938, n14939, n14940, n14941, n14942, n14943, n14944,
         n14945, n14947, n14948, n14949, n14950, n14951, n14952, n14953,
         n14954, n14955, n14956, n14957, n14958, n14959, n14960, n14961,
         n14962, n14963, n14964, n14965, n14966, n14967, n14968, n14969,
         n14970, n14971, n14972, n14973, n14974, n14975, n14976, n14977,
         n14978, n14979, n14980, n14981, n14982, n14983, n14984, n14985,
         n14986, n14987, n14988, n14989, n14990, n14991, n14992, n14993,
         n14994, n14995, n14996, n14997, n14998, n14999, n15000, n15001,
         n15002, n15003, n15004, n15005, n15006, n15007, n15008, n15009,
         n15010, n15011, n15012, n15013, n15014, n15015, n15016, n15017,
         n15018, n15019, n15020, n15021, n15022, n15023, n15024, n15025,
         n15026, n15027, n15028, n15029, n15030, n15031, n15032, n15033,
         n15034, n15035, n15036, n15037, n15038, n15039, n15040, n15041,
         n15042, n15043, n15044, n15045, n15046, n15047, n15048, n15049,
         n15050, n15051, n15052, n15053, n15054, n15055, n15056, n15057,
         n15058, n15059, n15060, n15061, n15062, n15063, n15064, n15065,
         n15066, n15067, n15068, n15069, n15070, n15071, n15072, n15073,
         n15074, n15075, n15076, n15077, n15078, n15079, n15080, n15081,
         n15082, n15083, n15084, n15085, n15086, n15087, n15088, n15089,
         n15090, n15091, n15092, n15093, n15094, n15095, n15096, n15097,
         n15098, n15099, n15100, n15101, n15102, n15103, n15104, n15105,
         n15106, n15107, n15108, n15109, n15110, n15111, n15112, n15113,
         n15114, n15115, n15116, n15117, n15118, n15119, n15120, n15121,
         n15122, n15123, n15124, n15125, n15126, n15127, n15128, n15129,
         n15130, n15131, n15132, n15133, n15134, n15135, n15136, n15137,
         n15138, n15139, n15140, n15141, n15142, n15143, n15144, n15145,
         n15146, n15147, n15148, n15149, n15150, n15151, n15152, n15153,
         n15154, n15155, n15156, n15157, n15158, n15159, n15160, n15161,
         n15162, n15163, n15164, n15165, n15166, n15167, n15168, n15169,
         n15170, n15171, n15172, n15173, n15174, n15175, n15176, n15177,
         n15178, n15179, n15180, n15181, n15182, n15183, n15184, n15185,
         n15186, n15187, n15188, n15189, n15190, n15191, n15192, n15193,
         n15194, n15195, n15196, n15197, n15198, n15199, n15200, n15201,
         n15202, n15203, n15204, n15205, n15206, n15207, n15208;

  INV_X4 U7215 ( .A(P3_STATE_REG_SCAN_IN), .ZN(P3_U3151) );
  NAND2_X1 U7216 ( .A1(n11576), .A2(n11575), .ZN(n14216) );
  XNOR2_X1 U7217 ( .A(n8659), .B(SI_24_), .ZN(n8635) );
  INV_X1 U7218 ( .A(n9355), .ZN(n12273) );
  NAND2_X1 U7219 ( .A1(n9412), .A2(n9324), .ZN(n12223) );
  CLKBUF_X1 U7220 ( .A(n6973), .Z(n6482) );
  CLKBUF_X2 U7221 ( .A(n11797), .Z(n6483) );
  NAND2_X1 U7222 ( .A1(n8089), .A2(n8088), .ZN(n13270) );
  CLKBUF_X1 U7223 ( .A(n8049), .Z(n8746) );
  INV_X1 U7224 ( .A(n8056), .ZN(n9640) );
  INV_X1 U7225 ( .A(n8066), .ZN(n8667) );
  AND2_X2 U7226 ( .A1(n11647), .A2(n11667), .ZN(n7454) );
  NAND2_X2 U7227 ( .A1(n9350), .A2(n9349), .ZN(n14187) );
  AND2_X1 U7228 ( .A1(n9328), .A2(n9327), .ZN(n10452) );
  CLKBUF_X2 U7229 ( .A(n8069), .Z(n8780) );
  INV_X2 U7230 ( .A(n6483), .ZN(n11980) );
  XNOR2_X1 U7231 ( .A(n10092), .B(n15069), .ZN(n15058) );
  XNOR2_X1 U7233 ( .A(n13729), .B(n13304), .ZN(n13565) );
  NAND2_X1 U7234 ( .A1(n8056), .A2(n9434), .ZN(n8066) );
  NAND2_X1 U7235 ( .A1(n13534), .A2(n13526), .ZN(n13515) );
  INV_X1 U7236 ( .A(n9342), .ZN(n12303) );
  INV_X2 U7237 ( .A(n12223), .ZN(n10746) );
  AND2_X1 U7238 ( .A1(n9329), .A2(n9327), .ZN(n10474) );
  INV_X1 U7239 ( .A(n10088), .ZN(n10111) );
  INV_X1 U7240 ( .A(n12754), .ZN(n13003) );
  INV_X1 U7241 ( .A(n12671), .ZN(n12689) );
  AND3_X1 U7242 ( .A1(n7435), .A2(n7352), .A3(n7434), .ZN(n15125) );
  INV_X1 U7243 ( .A(n8050), .ZN(n8768) );
  NAND2_X2 U7244 ( .A1(n8821), .A2(n8820), .ZN(n8056) );
  NAND2_X1 U7245 ( .A1(n8516), .A2(n8515), .ZN(n13752) );
  NAND2_X1 U7246 ( .A1(n8254), .A2(n7980), .ZN(n8009) );
  NAND2_X2 U7247 ( .A1(n11554), .A2(n11553), .ZN(n14226) );
  OR2_X1 U7248 ( .A1(n14089), .A2(n14221), .ZN(n14071) );
  INV_X1 U7249 ( .A(n14149), .ZN(n12035) );
  INV_X1 U7250 ( .A(n12273), .ZN(n11452) );
  NOR2_X2 U7251 ( .A1(n14071), .A2(n14216), .ZN(n11693) );
  INV_X2 U7252 ( .A(n14493), .ZN(n7114) );
  OAI21_X1 U7253 ( .B1(n8084), .B2(P2_DATAO_REG_1__SCAN_IN), .A(n8031), .ZN(
        n8063) );
  XNOR2_X1 U7254 ( .A(n10261), .B(n10269), .ZN(n10154) );
  XNOR2_X1 U7255 ( .A(n7385), .B(P3_IR_REG_30__SCAN_IN), .ZN(n7391) );
  OAI21_X1 U7256 ( .B1(n8056), .B2(n8008), .A(n8007), .ZN(n10216) );
  AOI21_X1 U7257 ( .B1(n13706), .B2(n14986), .A(n13705), .ZN(n13707) );
  INV_X1 U7258 ( .A(n9377), .ZN(n9420) );
  BUF_X1 U7259 ( .A(n14176), .Z(n6473) );
  INV_X2 U7260 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n10128) );
  NAND2_X1 U7261 ( .A1(n14728), .A2(n13995), .ZN(n6467) );
  INV_X1 U7262 ( .A(n11792), .ZN(n11797) );
  OR2_X2 U7263 ( .A1(n11786), .A2(n11787), .ZN(n6584) );
  AOI21_X2 U7264 ( .B1(n11690), .B2(n14701), .A(n11689), .ZN(n14214) );
  NOR2_X2 U7265 ( .A1(n10062), .A2(n15021), .ZN(n15020) );
  NAND2_X2 U7266 ( .A1(n8179), .A2(n8178), .ZN(n8209) );
  INV_X1 U7267 ( .A(n9174), .ZN(n6468) );
  INV_X1 U7268 ( .A(n6468), .ZN(n6469) );
  NOR2_X2 U7269 ( .A1(n10799), .A2(n14987), .ZN(n6677) );
  NAND2_X2 U7270 ( .A1(n10877), .A2(n7874), .ZN(n10892) );
  NAND2_X2 U7271 ( .A1(n10938), .A2(n10937), .ZN(n14478) );
  CLKBUF_X1 U7272 ( .A(n14012), .Z(n6470) );
  XNOR2_X1 U7273 ( .A(n9373), .B(P1_IR_REG_2__SCAN_IN), .ZN(n14012) );
  MUX2_X2 U7274 ( .A(n14728), .B(n13995), .S(n6476), .Z(n11786) );
  OR2_X2 U7275 ( .A1(n14728), .A2(n13995), .ZN(n9755) );
  NOR2_X1 U7276 ( .A1(n14728), .A2(n10396), .ZN(n10399) );
  NAND2_X1 U7277 ( .A1(n7916), .A2(n7915), .ZN(n6471) );
  NAND2_X1 U7278 ( .A1(n7916), .A2(n7915), .ZN(n6472) );
  NAND2_X1 U7279 ( .A1(n7916), .A2(n7915), .ZN(n7450) );
  NAND2_X2 U7280 ( .A1(n14724), .A2(n11972), .ZN(n14493) );
  AOI21_X2 U7281 ( .B1(n9525), .B2(n7930), .A(n6570), .ZN(n13239) );
  INV_X4 U7282 ( .A(n7471), .ZN(n12515) );
  OR3_X2 U7283 ( .A1(n12542), .A2(n12541), .A3(n12893), .ZN(n12720) );
  OAI211_X1 U7284 ( .C1(n9435), .C2(n9371), .A(n9345), .B(n6907), .ZN(n14176)
         );
  CLKBUF_X1 U7285 ( .A(n10474), .Z(n6474) );
  BUF_X4 U7286 ( .A(n10474), .Z(n6475) );
  XNOR2_X2 U7287 ( .A(n7990), .B(n7989), .ZN(n11662) );
  NAND2_X2 U7288 ( .A1(n7988), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7990) );
  XNOR2_X2 U7289 ( .A(n14226), .B(n12275), .ZN(n14082) );
  INV_X1 U7290 ( .A(n12763), .ZN(n15112) );
  MUX2_X1 U7291 ( .A(n11978), .B(n11979), .S(n11963), .Z(n6476) );
  MUX2_X2 U7292 ( .A(n11978), .B(n11979), .S(n11963), .Z(n11792) );
  OAI211_X4 U7293 ( .C1(n9343), .C2(n7074), .A(n9344), .B(n7073), .ZN(n9582)
         );
  OAI21_X2 U7294 ( .B1(n9795), .B2(n9962), .A(n9785), .ZN(n9786) );
  NAND2_X2 U7295 ( .A1(n7430), .A2(n7429), .ZN(n9795) );
  AND2_X2 U7296 ( .A1(n11951), .A2(n6676), .ZN(n11953) );
  AND2_X2 U7297 ( .A1(n6747), .A2(n8101), .ZN(n8254) );
  AOI21_X2 U7298 ( .B1(n12872), .B2(n15167), .A(n12867), .ZN(n8898) );
  OAI21_X2 U7299 ( .B1(n8879), .B2(n15115), .A(n8878), .ZN(n12867) );
  AOI21_X2 U7300 ( .B1(P3_ADDR_REG_12__SCAN_IN), .B2(n14586), .A(n8915), .ZN(
        n8928) );
  XNOR2_X2 U7301 ( .A(n11734), .B(n11325), .ZN(n11327) );
  AND2_X2 U7302 ( .A1(n7184), .A2(n7183), .ZN(n10092) );
  OAI22_X2 U7303 ( .A1(n13543), .A2(n13547), .B1(n6955), .B2(n13378), .ZN(
        n13531) );
  AOI21_X2 U7304 ( .B1(n13566), .B2(n13561), .A(n12116), .ZN(n13543) );
  OAI21_X2 U7305 ( .B1(n10353), .B2(n10352), .A(n11718), .ZN(n10354) );
  XNOR2_X2 U7306 ( .A(n12088), .B(n12086), .ZN(n13261) );
  NAND2_X2 U7307 ( .A1(n7671), .A2(n7670), .ZN(n13167) );
  NAND2_X2 U7308 ( .A1(n8617), .A2(n8616), .ZN(n13729) );
  NOR2_X2 U7309 ( .A1(n14351), .A2(n14353), .ZN(n14352) );
  AOI21_X1 U7310 ( .B1(P3_REG2_REG_10__SCAN_IN), .B2(n11021), .A(n11020), .ZN(
        n11138) );
  XNOR2_X2 U7311 ( .A(n10694), .B(n10714), .ZN(n15080) );
  AOI21_X1 U7312 ( .B1(n11634), .B2(n14701), .A(n11633), .ZN(n11635) );
  AOI211_X1 U7313 ( .C1(n13701), .C2(n13669), .A(n12147), .B(n12146), .ZN(
        n12148) );
  NAND2_X1 U7314 ( .A1(n14078), .A2(n14077), .ZN(n14076) );
  NAND2_X1 U7315 ( .A1(n11749), .A2(n11752), .ZN(n12066) );
  NOR2_X1 U7316 ( .A1(n12768), .A2(n13067), .ZN(n12787) );
  INV_X1 U7317 ( .A(n12761), .ZN(n10876) );
  NAND2_X2 U7318 ( .A1(n15112), .A2(n7868), .ZN(n12563) );
  NAND2_X1 U7319 ( .A1(n7441), .A2(n6522), .ZN(n12763) );
  INV_X1 U7320 ( .A(n15135), .ZN(n7868) );
  INV_X1 U7321 ( .A(n15107), .ZN(n15130) );
  INV_X2 U7322 ( .A(n7454), .ZN(n7471) );
  CLKBUF_X3 U7323 ( .A(n10036), .Z(n6485) );
  CLKBUF_X2 U7324 ( .A(n12163), .Z(n12159) );
  CLKBUF_X2 U7326 ( .A(n8667), .Z(n8761) );
  NOR2_X2 U7327 ( .A1(n12547), .A2(n10288), .ZN(n12727) );
  NAND2_X1 U7328 ( .A1(n6472), .A2(n9434), .ZN(n7462) );
  XNOR2_X1 U7329 ( .A(n7298), .B(P1_IR_REG_30__SCAN_IN), .ZN(n9329) );
  AND2_X2 U7330 ( .A1(n8021), .A2(n10871), .ZN(n9832) );
  NAND2_X1 U7331 ( .A1(n9438), .A2(P3_U3151), .ZN(n13247) );
  NAND2_X1 U7332 ( .A1(n9308), .A2(n9311), .ZN(n9325) );
  CLKBUF_X1 U7333 ( .A(n7667), .Z(n7668) );
  INV_X1 U7334 ( .A(P2_RD_REG_SCAN_IN), .ZN(n14305) );
  INV_X1 U7335 ( .A(n6705), .ZN(n14218) );
  OAI21_X1 U7336 ( .B1(n14219), .B2(n11636), .A(n11635), .ZN(n6705) );
  OR2_X1 U7337 ( .A1(n8887), .A2(n8886), .ZN(n12887) );
  AND2_X1 U7338 ( .A1(n7919), .A2(n7918), .ZN(n12882) );
  NAND2_X1 U7339 ( .A1(n13875), .A2(n12284), .ZN(n13952) );
  AND2_X1 U7340 ( .A1(n8892), .A2(n8893), .ZN(n6852) );
  NAND2_X1 U7341 ( .A1(n8863), .A2(n12679), .ZN(n12505) );
  NAND2_X1 U7342 ( .A1(n6741), .A2(n6517), .ZN(n11631) );
  OR2_X1 U7343 ( .A1(n14208), .A2(n14721), .ZN(n6507) );
  XNOR2_X1 U7344 ( .A(n11601), .B(n6889), .ZN(n14208) );
  NOR2_X1 U7345 ( .A1(n7907), .A2(n12685), .ZN(n8869) );
  AND2_X1 U7346 ( .A1(n13508), .A2(n13507), .ZN(n13708) );
  NAND2_X1 U7347 ( .A1(n7262), .A2(n7261), .ZN(n14067) );
  NOR2_X1 U7348 ( .A1(n13713), .A2(n13712), .ZN(n13714) );
  NAND2_X1 U7349 ( .A1(n6756), .A2(n7148), .ZN(n13503) );
  NAND2_X1 U7350 ( .A1(n6894), .A2(n6893), .ZN(n11694) );
  AOI21_X1 U7351 ( .B1(n6963), .B2(n6966), .A(n12677), .ZN(n6961) );
  OR2_X1 U7352 ( .A1(n13335), .A2(n12089), .ZN(n13297) );
  OR2_X1 U7353 ( .A1(n8880), .A2(n11677), .ZN(n12687) );
  NOR2_X1 U7354 ( .A1(n11610), .A2(n7265), .ZN(n7264) );
  OR2_X1 U7355 ( .A1(n14082), .A2(n7267), .ZN(n7263) );
  NOR2_X1 U7356 ( .A1(n12449), .A2(n12751), .ZN(n12448) );
  NAND2_X1 U7357 ( .A1(n7840), .A2(n7839), .ZN(n7954) );
  NAND2_X1 U7358 ( .A1(n8764), .A2(n8763), .ZN(n13706) );
  NAND2_X1 U7359 ( .A1(n8641), .A2(n8640), .ZN(n13724) );
  NAND2_X1 U7360 ( .A1(n7828), .A2(n7827), .ZN(n12535) );
  NAND2_X1 U7361 ( .A1(n8669), .A2(n8668), .ZN(n13719) );
  NAND2_X1 U7362 ( .A1(n12066), .A2(n12065), .ZN(n12081) );
  INV_X1 U7363 ( .A(n12667), .ZN(n6977) );
  OR2_X1 U7364 ( .A1(n14157), .A2(n14165), .ZN(n14155) );
  OAI21_X1 U7365 ( .B1(n7837), .B2(n7836), .A(n7835), .ZN(n8865) );
  OR2_X1 U7366 ( .A1(n11262), .A2(n11261), .ZN(n14487) );
  NAND2_X1 U7367 ( .A1(n7894), .A2(n7893), .ZN(n12997) );
  XNOR2_X1 U7368 ( .A(n8635), .B(n8660), .ZN(n11543) );
  NAND2_X1 U7369 ( .A1(n13275), .A2(n6523), .ZN(n13277) );
  NAND2_X1 U7370 ( .A1(n8596), .A2(n8595), .ZN(n13735) );
  NOR2_X1 U7371 ( .A1(n7195), .A2(n7192), .ZN(n14389) );
  NAND2_X1 U7372 ( .A1(n8568), .A2(n8567), .ZN(n13740) );
  OAI21_X1 U7373 ( .B1(n7800), .B2(P2_DATAO_REG_24__SCAN_IN), .A(n7799), .ZN(
        n7811) );
  NOR2_X1 U7374 ( .A1(n14373), .A2(n14372), .ZN(n14374) );
  NAND2_X1 U7375 ( .A1(n8594), .A2(n8593), .ZN(n8612) );
  NAND2_X1 U7376 ( .A1(n6811), .A2(n7750), .ZN(n12545) );
  NAND2_X1 U7377 ( .A1(n6729), .A2(n7237), .ZN(n11183) );
  OR2_X1 U7378 ( .A1(n7787), .A2(n11396), .ZN(n7799) );
  NAND2_X1 U7379 ( .A1(n6952), .A2(n6951), .ZN(n13662) );
  NAND2_X1 U7380 ( .A1(n11360), .A2(n11361), .ZN(n11359) );
  INV_X1 U7381 ( .A(n13672), .ZN(n6952) );
  NAND2_X1 U7382 ( .A1(n12327), .A2(n9215), .ZN(n12492) );
  OAI21_X1 U7383 ( .B1(n11288), .B2(n6552), .A(n6503), .ZN(n6719) );
  NAND2_X1 U7384 ( .A1(n6662), .A2(n6556), .ZN(n11734) );
  NAND2_X1 U7385 ( .A1(n11432), .A2(n11431), .ZN(n11899) );
  NAND2_X1 U7386 ( .A1(n8467), .A2(n8466), .ZN(n13763) );
  NAND2_X1 U7387 ( .A1(n6720), .A2(n6536), .ZN(n11288) );
  XNOR2_X1 U7388 ( .A(n6897), .B(n8486), .ZN(n11428) );
  NAND2_X1 U7389 ( .A1(n8513), .A2(SI_20_), .ZN(n8539) );
  OR2_X1 U7390 ( .A1(n11016), .A2(n11015), .ZN(n14513) );
  NAND2_X1 U7391 ( .A1(n8364), .A2(n8363), .ZN(n13767) );
  XNOR2_X1 U7392 ( .A(n14027), .B(n11164), .ZN(n11407) );
  OAI21_X1 U7393 ( .B1(n8482), .B2(n8503), .A(n8483), .ZN(n6897) );
  AND2_X1 U7394 ( .A1(n14603), .A2(n7078), .ZN(n14027) );
  INV_X1 U7395 ( .A(n11632), .ZN(n11633) );
  AND2_X1 U7396 ( .A1(n13110), .A2(n12603), .ZN(n13090) );
  NAND2_X1 U7397 ( .A1(n11182), .A2(n11181), .ZN(n14498) );
  OAI21_X1 U7398 ( .B1(n8461), .B2(n6932), .A(n6931), .ZN(n8511) );
  NAND2_X1 U7399 ( .A1(n8377), .A2(n8376), .ZN(n13772) );
  NAND2_X1 U7400 ( .A1(n6994), .A2(n6545), .ZN(n10840) );
  NAND2_X1 U7401 ( .A1(n6900), .A2(n8356), .ZN(n8461) );
  AOI21_X1 U7402 ( .B1(P3_ADDR_REG_11__SCAN_IN), .B2(n14574), .A(n8914), .ZN(
        n8976) );
  NAND2_X1 U7403 ( .A1(n8397), .A2(n8396), .ZN(n13780) );
  NAND2_X1 U7404 ( .A1(n10988), .A2(n10987), .ZN(n14442) );
  OAI21_X1 U7405 ( .B1(n7628), .B2(n7046), .A(n7044), .ZN(n7647) );
  NAND2_X1 U7406 ( .A1(n10945), .A2(n10944), .ZN(n11849) );
  NAND2_X1 U7407 ( .A1(n10941), .A2(n10940), .ZN(n14477) );
  NAND2_X1 U7408 ( .A1(n8288), .A2(n8287), .ZN(n10854) );
  OAI21_X1 U7409 ( .B1(n8325), .B2(n6492), .A(n6938), .ZN(n8347) );
  NAND2_X1 U7410 ( .A1(n10570), .A2(n10569), .ZN(n14778) );
  NOR2_X1 U7411 ( .A1(n10266), .A2(n10265), .ZN(n10693) );
  AND2_X1 U7412 ( .A1(n12595), .A2(n12594), .ZN(n12707) );
  NAND2_X1 U7413 ( .A1(n13267), .A2(n10043), .ZN(n11716) );
  NAND2_X1 U7414 ( .A1(n6715), .A2(n8211), .ZN(n8231) );
  OAI21_X2 U7415 ( .B1(n9819), .B2(n10141), .A(n13607), .ZN(n9820) );
  INV_X2 U7416 ( .A(n13606), .ZN(n13671) );
  NAND2_X1 U7417 ( .A1(n12703), .A2(n10412), .ZN(n15114) );
  AND2_X1 U7418 ( .A1(n7207), .A2(n7206), .ZN(n10152) );
  INV_X1 U7419 ( .A(n9888), .ZN(n10669) );
  OR2_X1 U7420 ( .A1(n15057), .A2(n10094), .ZN(n7207) );
  NOR2_X1 U7421 ( .A1(n8906), .A2(n8907), .ZN(n8952) );
  NAND2_X1 U7422 ( .A1(n6916), .A2(n8154), .ZN(n8176) );
  NOR2_X1 U7423 ( .A1(n8946), .A2(P1_ADDR_REG_5__SCAN_IN), .ZN(n8906) );
  NAND4_X1 U7424 ( .A1(n7418), .A2(n7417), .A3(n7416), .A4(n7415), .ZN(n12766)
         );
  INV_X1 U7425 ( .A(n15125), .ZN(n10416) );
  OAI211_X1 U7426 ( .C1(n7448), .C2(n14313), .A(n7410), .B(n6972), .ZN(n15107)
         );
  NAND2_X1 U7427 ( .A1(n7453), .A2(n7452), .ZN(n15135) );
  NAND2_X1 U7428 ( .A1(n6675), .A2(n8138), .ZN(n8152) );
  AND2_X2 U7429 ( .A1(n9166), .A2(n9165), .ZN(n9178) );
  AND4_X1 U7430 ( .A1(n9333), .A2(n9332), .A3(n9331), .A4(n9330), .ZN(n9892)
         );
  AND3_X1 U7431 ( .A1(n9348), .A2(n9347), .A3(n9346), .ZN(n9350) );
  AND4_X1 U7432 ( .A1(n9363), .A2(n9362), .A3(n9361), .A4(n9360), .ZN(n11775)
         );
  AND2_X1 U7433 ( .A1(n7391), .A2(n7390), .ZN(n7437) );
  BUF_X2 U7434 ( .A(n11954), .Z(n11526) );
  OR2_X1 U7435 ( .A1(n15046), .A2(n15045), .ZN(n7184) );
  INV_X1 U7436 ( .A(n6477), .ZN(n6478) );
  INV_X1 U7437 ( .A(n6477), .ZN(n6479) );
  NAND4_X1 U7438 ( .A1(n8055), .A2(n8054), .A3(n8053), .A4(n8052), .ZN(n8841)
         );
  CLKBUF_X3 U7439 ( .A(n6564), .Z(n11960) );
  INV_X2 U7440 ( .A(n10036), .ZN(n12098) );
  NAND2_X2 U7441 ( .A1(n14988), .A2(n13680), .ZN(n12163) );
  INV_X1 U7442 ( .A(n9329), .ZN(n9328) );
  INV_X2 U7443 ( .A(n8075), .ZN(n8767) );
  XNOR2_X1 U7444 ( .A(n6818), .B(P3_ADDR_REG_4__SCAN_IN), .ZN(n8930) );
  CLKBUF_X1 U7445 ( .A(n8050), .Z(n8750) );
  OAI21_X1 U7446 ( .B1(n8230), .B2(n6888), .A(n8251), .ZN(n6887) );
  CLKBUF_X1 U7447 ( .A(n8075), .Z(n8694) );
  NAND2_X1 U7448 ( .A1(n7387), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7388) );
  OAI21_X1 U7449 ( .B1(n8942), .B2(P1_ADDR_REG_3__SCAN_IN), .A(n6493), .ZN(
        n6818) );
  AND2_X1 U7450 ( .A1(n7992), .A2(n7991), .ZN(n8075) );
  NAND2_X1 U7451 ( .A1(n14287), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7298) );
  NAND2_X1 U7452 ( .A1(n11705), .A2(n7991), .ZN(n8050) );
  INV_X1 U7453 ( .A(n9327), .ZN(n14294) );
  CLKBUF_X3 U7454 ( .A(n7916), .Z(n12836) );
  NOR2_X1 U7455 ( .A1(n10108), .A2(n7351), .ZN(n10089) );
  INV_X1 U7456 ( .A(n13490), .ZN(n13680) );
  XNOR2_X1 U7457 ( .A(n9326), .B(P1_IR_REG_29__SCAN_IN), .ZN(n9327) );
  NAND2_X1 U7458 ( .A1(n9340), .A2(n9339), .ZN(n14149) );
  CLKBUF_X2 U7459 ( .A(n8021), .Z(n14938) );
  AND2_X1 U7460 ( .A1(n11705), .A2(n11662), .ZN(n8049) );
  AND2_X1 U7461 ( .A1(n7992), .A2(n11662), .ZN(n8095) );
  INV_X2 U7462 ( .A(n13813), .ZN(n13822) );
  MUX2_X1 U7463 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9338), .S(
        P1_IR_REG_19__SCAN_IN), .Z(n9340) );
  NAND2_X1 U7464 ( .A1(n9325), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6659) );
  OAI21_X1 U7465 ( .B1(n9325), .B2(P1_IR_REG_28__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n9326) );
  NAND2_X1 U7466 ( .A1(n8803), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8017) );
  XNOR2_X1 U7467 ( .A(n7987), .B(n7986), .ZN(n11705) );
  MUX2_X1 U7468 ( .A(P2_IR_REG_31__SCAN_IN), .B(n7999), .S(
        P2_IR_REG_27__SCAN_IN), .Z(n8002) );
  AND2_X1 U7469 ( .A1(n7691), .A2(n7723), .ZN(n7851) );
  CLKBUF_X1 U7470 ( .A(n9302), .Z(n6668) );
  NOR3_X1 U7471 ( .A1(n7668), .A2(P3_IR_REG_26__SCAN_IN), .A3(n6982), .ZN(
        n6981) );
  AND2_X1 U7472 ( .A1(n7687), .A2(n7378), .ZN(n7691) );
  AND3_X1 U7473 ( .A1(n7477), .A2(n7377), .A3(n6605), .ZN(n6842) );
  INV_X4 U7474 ( .A(n8084), .ZN(n11519) );
  AND2_X1 U7475 ( .A1(n9284), .A2(n9336), .ZN(n9294) );
  AND3_X1 U7476 ( .A1(n9279), .A2(n9278), .A3(n9277), .ZN(n9281) );
  AND2_X1 U7477 ( .A1(n7381), .A2(n7378), .ZN(n7345) );
  AND2_X1 U7478 ( .A1(n9283), .A2(n9282), .ZN(n9336) );
  AND2_X1 U7479 ( .A1(n9274), .A2(n9569), .ZN(n9279) );
  AND4_X1 U7480 ( .A1(n7371), .A2(n7370), .A3(n7369), .A4(n7368), .ZN(n7377)
         );
  AND4_X1 U7481 ( .A1(n7375), .A2(n7476), .A3(n7374), .A4(n7373), .ZN(n7376)
         );
  NAND2_X1 U7482 ( .A1(n7383), .A2(n6983), .ZN(n6982) );
  AND2_X1 U7483 ( .A1(n8057), .A2(n7975), .ZN(n8101) );
  AND4_X1 U7484 ( .A1(n7380), .A2(n7379), .A3(n7854), .A4(n7850), .ZN(n7381)
         );
  AND4_X1 U7485 ( .A1(n7974), .A2(n7973), .A3(n7972), .A4(n7971), .ZN(n6747)
         );
  NOR2_X1 U7486 ( .A1(P1_IR_REG_16__SCAN_IN), .A2(P1_IR_REG_15__SCAN_IN), .ZN(
        n9282) );
  NOR2_X1 U7487 ( .A1(P1_IR_REG_18__SCAN_IN), .A2(P1_IR_REG_17__SCAN_IN), .ZN(
        n9283) );
  INV_X1 U7488 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n9286) );
  NOR2_X1 U7489 ( .A1(P3_IR_REG_10__SCAN_IN), .A2(P3_IR_REG_14__SCAN_IN), .ZN(
        n7369) );
  NOR2_X1 U7490 ( .A1(P3_IR_REG_13__SCAN_IN), .A2(P3_IR_REG_15__SCAN_IN), .ZN(
        n7370) );
  NOR2_X1 U7491 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(P1_IR_REG_9__SCAN_IN), .ZN(
        n9569) );
  NOR2_X1 U7492 ( .A1(P3_IR_REG_8__SCAN_IN), .A2(P3_IR_REG_7__SCAN_IN), .ZN(
        n7368) );
  INV_X4 U7493 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3088) );
  NOR3_X1 U7494 ( .A1(P1_IR_REG_11__SCAN_IN), .A2(P1_IR_REG_5__SCAN_IN), .A3(
        P1_IR_REG_4__SCAN_IN), .ZN(n9277) );
  INV_X1 U7495 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n9309) );
  NOR2_X1 U7496 ( .A1(P3_IR_REG_21__SCAN_IN), .A2(P3_IR_REG_23__SCAN_IN), .ZN(
        n7379) );
  NOR2_X1 U7497 ( .A1(P2_IR_REG_4__SCAN_IN), .A2(P2_IR_REG_3__SCAN_IN), .ZN(
        n7973) );
  INV_X4 U7498 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  NOR2_X2 U7499 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n9372) );
  NOR2_X1 U7500 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n8057) );
  NOR2_X1 U7501 ( .A1(P2_IR_REG_7__SCAN_IN), .A2(P2_IR_REG_9__SCAN_IN), .ZN(
        n7972) );
  BUF_X1 U7502 ( .A(P1_IR_REG_0__SCAN_IN), .Z(n14299) );
  INV_X1 U7503 ( .A(n11521), .ZN(n11429) );
  AND2_X1 U7504 ( .A1(n14298), .A2(n11521), .ZN(n14247) );
  NOR2_X1 U7505 ( .A1(n11022), .A2(n11023), .ZN(n11140) );
  NOR2_X2 U7506 ( .A1(n11316), .A2(n13767), .ZN(n6954) );
  INV_X1 U7507 ( .A(n8060), .ZN(n8068) );
  NOR3_X2 U7508 ( .A1(n9836), .A2(n9835), .A3(n9837), .ZN(n9931) );
  INV_X1 U7509 ( .A(n11429), .ZN(n6477) );
  INV_X4 U7510 ( .A(n7468), .ZN(n7423) );
  NOR2_X1 U7511 ( .A1(n10012), .A2(n10216), .ZN(n10013) );
  NOR2_X2 U7512 ( .A1(n10354), .A2(n10355), .ZN(n10596) );
  AOI22_X2 U7513 ( .A1(n9374), .A2(P2_DATAO_REG_2__SCAN_IN), .B1(n11429), .B2(
        n6470), .ZN(n9375) );
  CLKBUF_X1 U7514 ( .A(n9506), .Z(n6484) );
  XNOR2_X1 U7515 ( .A(n9312), .B(n9311), .ZN(n9506) );
  AND2_X1 U7516 ( .A1(n11007), .A2(n6508), .ZN(n11243) );
  NOR2_X2 U7517 ( .A1(n14480), .A2(n11849), .ZN(n11007) );
  AOI21_X2 U7518 ( .B1(P1_REG2_REG_16__SCAN_IN), .B2(n14625), .A(n14620), .ZN(
        n14635) );
  NOR2_X2 U7519 ( .A1(n11363), .A2(n13780), .ZN(n11366) );
  OR2_X2 U7520 ( .A1(n11277), .A2(n13784), .ZN(n11363) );
  XNOR2_X2 U7521 ( .A(n7998), .B(n7997), .ZN(n8821) );
  OR2_X1 U7522 ( .A1(n8026), .A2(n8117), .ZN(n6657) );
  NAND2_X1 U7523 ( .A1(n12889), .A2(n7904), .ZN(n7326) );
  INV_X1 U7524 ( .A(n6982), .ZN(n6841) );
  NOR2_X1 U7525 ( .A1(n11613), .A2(n14209), .ZN(n6901) );
  NAND2_X1 U7526 ( .A1(n14164), .A2(n11605), .ZN(n14141) );
  INV_X1 U7527 ( .A(n12762), .ZN(n10363) );
  INV_X1 U7528 ( .A(n10660), .ZN(n9182) );
  NAND2_X1 U7529 ( .A1(n9386), .A2(n9408), .ZN(n6772) );
  NAND2_X1 U7530 ( .A1(n14130), .A2(n6898), .ZN(n14112) );
  NOR2_X1 U7531 ( .A1(n14102), .A2(n6899), .ZN(n6898) );
  INV_X1 U7532 ( .A(n11542), .ZN(n6899) );
  NAND2_X1 U7533 ( .A1(n8073), .A2(n6529), .ZN(n7212) );
  NAND2_X1 U7534 ( .A1(n8541), .A2(SI_21_), .ZN(n8563) );
  INV_X1 U7535 ( .A(n7437), .ZN(n7455) );
  INV_X1 U7536 ( .A(n11667), .ZN(n7390) );
  NAND2_X1 U7537 ( .A1(n11024), .A2(n6872), .ZN(n11145) );
  OR2_X1 U7538 ( .A1(n11025), .A2(n13178), .ZN(n6872) );
  OR2_X1 U7539 ( .A1(n12480), .A2(n9266), .ZN(n12540) );
  OR2_X1 U7540 ( .A1(n13134), .A2(n12450), .ZN(n12669) );
  NAND2_X1 U7541 ( .A1(n12764), .A2(n15125), .ZN(n12557) );
  NOR2_X1 U7542 ( .A1(n7327), .A2(n7325), .ZN(n7324) );
  INV_X1 U7543 ( .A(n7905), .ZN(n7325) );
  INV_X1 U7544 ( .A(n12541), .ZN(n7327) );
  INV_X1 U7545 ( .A(P3_IR_REG_24__SCAN_IN), .ZN(n7382) );
  NAND2_X1 U7546 ( .A1(n7060), .A2(n7058), .ZN(n7786) );
  AOI21_X1 U7547 ( .B1(n7053), .B2(n7056), .A(n6796), .ZN(n6795) );
  INV_X1 U7548 ( .A(n7705), .ZN(n6796) );
  NAND2_X1 U7549 ( .A1(n7610), .A2(n7609), .ZN(n6809) );
  INV_X1 U7550 ( .A(n7051), .ZN(n7050) );
  OAI21_X1 U7551 ( .B1(n7566), .B2(n7052), .A(n7594), .ZN(n7051) );
  OR2_X1 U7552 ( .A1(n7569), .A2(P3_IR_REG_9__SCAN_IN), .ZN(n7604) );
  OR2_X1 U7553 ( .A1(n7547), .A2(P3_IR_REG_8__SCAN_IN), .ZN(n7569) );
  INV_X1 U7554 ( .A(n6803), .ZN(n6802) );
  OAI21_X1 U7555 ( .B1(n7481), .B2(n6804), .A(n7495), .ZN(n6803) );
  XNOR2_X1 U7556 ( .A(n13694), .B(n13372), .ZN(n8827) );
  INV_X1 U7557 ( .A(n13376), .ZN(n12143) );
  NAND2_X1 U7558 ( .A1(n10852), .A2(n10851), .ZN(n6755) );
  INV_X1 U7559 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n7985) );
  NAND2_X1 U7560 ( .A1(n6590), .A2(n12227), .ZN(n6783) );
  INV_X1 U7561 ( .A(n10942), .ZN(n7287) );
  NOR2_X1 U7562 ( .A1(n12006), .A2(n7260), .ZN(n7259) );
  INV_X1 U7563 ( .A(n10567), .ZN(n7260) );
  NAND2_X1 U7564 ( .A1(n14096), .A2(n6895), .ZN(n6894) );
  NOR2_X1 U7565 ( .A1(n7295), .A2(n6896), .ZN(n6895) );
  INV_X1 U7566 ( .A(n11562), .ZN(n6896) );
  INV_X1 U7567 ( .A(n7244), .ZN(n7243) );
  OAI21_X1 U7568 ( .B1(n11434), .B2(n6745), .A(n6743), .ZN(n7242) );
  OAI21_X1 U7569 ( .B1(n12019), .B2(n7245), .A(n14165), .ZN(n7244) );
  NAND2_X1 U7570 ( .A1(n10980), .A2(n10979), .ZN(n11053) );
  INV_X1 U7571 ( .A(n13988), .ZN(n11109) );
  NAND2_X1 U7572 ( .A1(n8708), .A2(n8707), .ZN(n8760) );
  OR2_X1 U7573 ( .A1(n8705), .A2(n8704), .ZN(n8708) );
  NAND2_X1 U7574 ( .A1(n8564), .A2(n8563), .ZN(n8592) );
  INV_X1 U7575 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n9284) );
  AOI22_X1 U7576 ( .A1(P3_ADDR_REG_15__SCAN_IN), .A2(n8980), .B1(n8981), .B2(
        n8919), .ZN(n8983) );
  AND2_X1 U7577 ( .A1(n6488), .A2(n6528), .ZN(n7034) );
  AND4_X1 U7578 ( .A1(n7660), .A2(n7659), .A3(n7658), .A4(n7657), .ZN(n12332)
         );
  INV_X1 U7579 ( .A(n10096), .ZN(n7206) );
  INV_X1 U7580 ( .A(n12817), .ZN(n7179) );
  OAI21_X1 U7581 ( .B1(n14373), .B2(n7198), .A(n7196), .ZN(n7195) );
  NAND2_X1 U7582 ( .A1(n12848), .A2(n7199), .ZN(n7198) );
  NOR2_X1 U7583 ( .A1(n7197), .A2(n7201), .ZN(n7196) );
  NOR2_X1 U7584 ( .A1(n14379), .A2(n7202), .ZN(n7201) );
  NAND2_X1 U7585 ( .A1(n14373), .A2(n7194), .ZN(n7193) );
  INV_X1 U7586 ( .A(n7200), .ZN(n7194) );
  OAI21_X1 U7587 ( .B1(n6813), .B2(n6583), .A(n6812), .ZN(n12933) );
  INV_X1 U7588 ( .A(n6515), .ZN(n6812) );
  INV_X1 U7589 ( .A(n12947), .ZN(n6813) );
  INV_X1 U7590 ( .A(n13103), .ZN(n15115) );
  NAND2_X1 U7591 ( .A1(n12887), .A2(n6850), .ZN(n6846) );
  OR2_X1 U7592 ( .A1(n15120), .A2(n15161), .ZN(n6850) );
  INV_X1 U7593 ( .A(n7448), .ZN(n12520) );
  NAND2_X1 U7594 ( .A1(n13242), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7385) );
  NAND2_X1 U7595 ( .A1(n6793), .A2(n6795), .ZN(n7718) );
  OR2_X1 U7596 ( .A1(n7665), .A2(n6797), .ZN(n6793) );
  AND2_X1 U7597 ( .A1(n7703), .A2(n7686), .ZN(n7701) );
  NAND2_X1 U7598 ( .A1(n6809), .A2(n10982), .ZN(n7627) );
  AND2_X1 U7599 ( .A1(n6991), .A2(n6592), .ZN(n6989) );
  AND2_X1 U7600 ( .A1(n14939), .A2(n14938), .ZN(n9824) );
  INV_X1 U7601 ( .A(n13694), .ZN(n6945) );
  INV_X1 U7602 ( .A(n8745), .ZN(n8765) );
  NAND2_X1 U7603 ( .A1(n8689), .A2(n8688), .ZN(n13711) );
  NAND2_X1 U7604 ( .A1(n6955), .A2(n7152), .ZN(n7151) );
  NOR2_X1 U7605 ( .A1(n13564), .A2(n12141), .ZN(n13548) );
  AND2_X1 U7606 ( .A1(n13729), .A2(n13379), .ZN(n12141) );
  NAND2_X1 U7607 ( .A1(n13548), .A2(n13547), .ZN(n13546) );
  INV_X1 U7608 ( .A(n12117), .ZN(n13547) );
  AND2_X1 U7609 ( .A1(n13729), .A2(n13304), .ZN(n12116) );
  OR2_X1 U7610 ( .A1(n11126), .A2(n7178), .ZN(n7170) );
  AND2_X1 U7611 ( .A1(n11730), .A2(n11123), .ZN(n11126) );
  INV_X1 U7612 ( .A(n11398), .ZN(n9800) );
  NAND2_X1 U7613 ( .A1(n9383), .A2(n9385), .ZN(n9386) );
  OR2_X1 U7614 ( .A1(n14462), .A2(n14461), .ZN(n6780) );
  NAND2_X1 U7615 ( .A1(n10646), .A2(n10645), .ZN(n6767) );
  NAND2_X1 U7616 ( .A1(n6777), .A2(n6776), .ZN(n12176) );
  AOI21_X1 U7617 ( .B1(n6778), .B2(n14461), .A(n6588), .ZN(n6776) );
  NAND2_X1 U7618 ( .A1(n14096), .A2(n11562), .ZN(n14078) );
  NAND2_X1 U7619 ( .A1(n14137), .A2(n14142), .ZN(n7292) );
  NAND2_X1 U7620 ( .A1(n6693), .A2(n6546), .ZN(n11427) );
  NAND2_X1 U7621 ( .A1(n6691), .A2(n6690), .ZN(n6693) );
  AND2_X1 U7622 ( .A1(n6692), .A2(n6598), .ZN(n6690) );
  AOI21_X1 U7623 ( .B1(n11015), .B2(n7241), .A(n7240), .ZN(n7239) );
  INV_X1 U7624 ( .A(n10995), .ZN(n7241) );
  INV_X1 U7625 ( .A(n11862), .ZN(n7240) );
  NAND2_X1 U7626 ( .A1(n6746), .A2(n10564), .ZN(n14672) );
  NAND2_X1 U7627 ( .A1(n10562), .A2(n11960), .ZN(n6746) );
  XNOR2_X1 U7628 ( .A(n14672), .B(n11109), .ZN(n14664) );
  AND2_X1 U7629 ( .A1(n6903), .A2(n6902), .ZN(n14206) );
  AOI21_X1 U7630 ( .B1(n9723), .B2(n8974), .A(n14541), .ZN(n8978) );
  NAND2_X1 U7631 ( .A1(n6837), .A2(n14908), .ZN(n6836) );
  INV_X1 U7632 ( .A(n14555), .ZN(n6837) );
  OR2_X1 U7633 ( .A1(n8923), .A2(n8922), .ZN(n8988) );
  NAND2_X1 U7634 ( .A1(n6822), .A2(n14927), .ZN(n7087) );
  AND2_X1 U7635 ( .A1(n14560), .A2(n6821), .ZN(n6820) );
  INV_X1 U7636 ( .A(n14341), .ZN(n6821) );
  NAND2_X1 U7637 ( .A1(n7727), .A2(n7726), .ZN(n12991) );
  NAND2_X1 U7638 ( .A1(n10657), .A2(n9185), .ZN(n10754) );
  NAND2_X1 U7639 ( .A1(n6944), .A2(n13694), .ZN(n6943) );
  INV_X1 U7640 ( .A(n6946), .ZN(n6944) );
  NAND2_X1 U7641 ( .A1(n11535), .A2(n11534), .ZN(n14239) );
  OR2_X1 U7642 ( .A1(n14545), .A2(P2_ADDR_REG_12__SCAN_IN), .ZN(n6825) );
  XOR2_X1 U7643 ( .A(n8988), .B(n8989), .Z(n14302) );
  NAND2_X1 U7644 ( .A1(n11786), .A2(n6467), .ZN(n7300) );
  OAI21_X1 U7645 ( .B1(n10143), .B2(n8117), .A(n8072), .ZN(n8073) );
  INV_X1 U7646 ( .A(n8092), .ZN(n6673) );
  OAI21_X1 U7647 ( .B1(n8206), .B2(n7346), .A(n8205), .ZN(n8226) );
  OR2_X1 U7648 ( .A1(n8204), .A2(n8203), .ZN(n8205) );
  NOR2_X1 U7649 ( .A1(n8249), .A2(n6544), .ZN(n7226) );
  NOR2_X1 U7650 ( .A1(n11869), .A2(n6561), .ZN(n7315) );
  NOR2_X1 U7651 ( .A1(n12011), .A2(n7317), .ZN(n7316) );
  NOR2_X1 U7652 ( .A1(n11860), .A2(n11861), .ZN(n7317) );
  NAND2_X1 U7653 ( .A1(n6656), .A2(n6655), .ZN(n6654) );
  INV_X1 U7654 ( .A(n6601), .ZN(n7217) );
  INV_X1 U7655 ( .A(n6602), .ZN(n7214) );
  NAND2_X1 U7656 ( .A1(n11928), .A2(n7306), .ZN(n7305) );
  INV_X1 U7657 ( .A(n11927), .ZN(n7306) );
  MUX2_X1 U7658 ( .A(n14121), .B(n14233), .S(n11980), .Z(n11927) );
  NOR2_X1 U7659 ( .A1(n12916), .A2(n6979), .ZN(n6978) );
  INV_X1 U7660 ( .A(n12669), .ZN(n6979) );
  AOI21_X1 U7661 ( .B1(n7720), .B2(n7043), .A(n7042), .ZN(n7041) );
  INV_X1 U7662 ( .A(n7733), .ZN(n7042) );
  INV_X1 U7663 ( .A(n7717), .ZN(n7043) );
  NAND2_X1 U7664 ( .A1(n6928), .A2(n6926), .ZN(n8512) );
  AOI21_X1 U7665 ( .B1(n6929), .B2(n6932), .A(n6927), .ZN(n6926) );
  NOR2_X1 U7666 ( .A1(n8510), .A2(n6930), .ZN(n6929) );
  NAND2_X1 U7667 ( .A1(n8350), .A2(n9639), .ZN(n8353) );
  NAND2_X1 U7668 ( .A1(n8325), .A2(n6487), .ZN(n6891) );
  INV_X1 U7669 ( .A(n8326), .ZN(n8329) );
  INV_X1 U7670 ( .A(n8233), .ZN(n6888) );
  INV_X1 U7671 ( .A(n8930), .ZN(n7081) );
  INV_X1 U7672 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n7080) );
  AND2_X1 U7673 ( .A1(n7951), .A2(n7950), .ZN(n9249) );
  NAND2_X1 U7674 ( .A1(n10159), .A2(n6873), .ZN(n10272) );
  OR2_X1 U7675 ( .A1(n10160), .A2(n15184), .ZN(n6873) );
  NAND2_X1 U7676 ( .A1(n10698), .A2(n6874), .ZN(n10700) );
  OR2_X1 U7677 ( .A1(n10699), .A2(n15188), .ZN(n6874) );
  INV_X1 U7678 ( .A(n12827), .ZN(n7182) );
  AOI21_X1 U7679 ( .B1(n12833), .B2(n12848), .A(n14382), .ZN(n12834) );
  NAND2_X1 U7680 ( .A1(n12929), .A2(n6978), .ZN(n12911) );
  OR2_X1 U7681 ( .A1(n13145), .A2(n12990), .ZN(n12650) );
  OR2_X1 U7682 ( .A1(n14417), .A2(n13050), .ZN(n12617) );
  NAND2_X1 U7683 ( .A1(n7334), .A2(n12706), .ZN(n7332) );
  NOR2_X1 U7684 ( .A1(n12707), .A2(n7335), .ZN(n7334) );
  INV_X1 U7685 ( .A(n7875), .ZN(n7335) );
  NOR2_X1 U7686 ( .A1(n7772), .A2(n7065), .ZN(n7064) );
  INV_X1 U7687 ( .A(n7758), .ZN(n7065) );
  NAND2_X1 U7688 ( .A1(n7853), .A2(n7854), .ZN(n7857) );
  INV_X1 U7689 ( .A(P3_IR_REG_19__SCAN_IN), .ZN(n7850) );
  INV_X1 U7690 ( .A(P3_IR_REG_17__SCAN_IN), .ZN(n7378) );
  INV_X1 U7691 ( .A(n7684), .ZN(n7057) );
  INV_X1 U7692 ( .A(n7581), .ZN(n7052) );
  INV_X1 U7693 ( .A(n7483), .ZN(n6804) );
  OR2_X1 U7694 ( .A1(n7479), .A2(P3_IR_REG_5__SCAN_IN), .ZN(n7509) );
  OAI21_X1 U7695 ( .B1(n8655), .B2(n8654), .A(n6582), .ZN(n7229) );
  AND2_X1 U7696 ( .A1(n6495), .A2(n6604), .ZN(n6722) );
  NAND2_X1 U7697 ( .A1(n6587), .A2(n12135), .ZN(n7144) );
  OAI21_X1 U7698 ( .B1(n7168), .B2(n7171), .A(n7175), .ZN(n7165) );
  NAND2_X1 U7699 ( .A1(n7176), .A2(n13386), .ZN(n7175) );
  INV_X1 U7700 ( .A(n10860), .ZN(n7173) );
  INV_X1 U7701 ( .A(n7132), .ZN(n7131) );
  OAI21_X1 U7702 ( .B1(n10373), .B2(n7133), .A(n10328), .ZN(n7132) );
  NAND2_X1 U7703 ( .A1(n7122), .A2(n8835), .ZN(n9922) );
  OR2_X1 U7704 ( .A1(n13767), .A2(n13316), .ZN(n12112) );
  XNOR2_X1 U7705 ( .A(n8011), .B(P2_IR_REG_21__SCAN_IN), .ZN(n8021) );
  INV_X1 U7706 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n7971) );
  INV_X1 U7707 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n7975) );
  NAND2_X1 U7708 ( .A1(n12247), .A2(n7109), .ZN(n7108) );
  INV_X1 U7709 ( .A(n12244), .ZN(n7109) );
  NAND3_X1 U7710 ( .A1(n14448), .A2(n7348), .A3(n6784), .ZN(n6782) );
  AND2_X1 U7711 ( .A1(n6542), .A2(n12227), .ZN(n6784) );
  AND2_X1 U7712 ( .A1(P1_REG3_REG_21__SCAN_IN), .A2(n11476), .ZN(n11522) );
  INV_X1 U7713 ( .A(n11475), .ZN(n11476) );
  NOR2_X1 U7714 ( .A1(n14634), .A2(n6648), .ZN(n14031) );
  OAI21_X1 U7715 ( .B1(n14138), .B2(n7249), .A(n14131), .ZN(n7248) );
  OR2_X1 U7716 ( .A1(n12184), .A2(n12188), .ZN(n11867) );
  OAI21_X1 U7717 ( .B1(n10578), .B2(n6489), .A(n14664), .ZN(n7274) );
  AND2_X1 U7718 ( .A1(n7270), .A2(n6696), .ZN(n6695) );
  NOR2_X1 U7719 ( .A1(n6489), .A2(n7271), .ZN(n7270) );
  NAND2_X1 U7720 ( .A1(n14687), .A2(n6697), .ZN(n6696) );
  INV_X1 U7721 ( .A(n13992), .ZN(n10650) );
  NAND2_X1 U7722 ( .A1(n6467), .A2(n9755), .ZN(n11997) );
  INV_X1 U7723 ( .A(n14204), .ZN(n11613) );
  AOI21_X1 U7724 ( .B1(n7294), .B2(n12026), .A(n6566), .ZN(n7293) );
  AND2_X1 U7725 ( .A1(n12203), .A2(n11243), .ZN(n11387) );
  AND2_X1 U7726 ( .A1(n12004), .A2(n7253), .ZN(n7252) );
  NAND2_X1 U7727 ( .A1(n14687), .A2(n10497), .ZN(n7253) );
  INV_X1 U7728 ( .A(n11979), .ZN(n11965) );
  NAND2_X1 U7729 ( .A1(n8760), .A2(n6512), .ZN(n6917) );
  AOI21_X1 U7730 ( .B1(n6512), .B2(n6919), .A(n6651), .ZN(n6918) );
  INV_X1 U7731 ( .A(n6924), .ZN(n6919) );
  AOI21_X1 U7732 ( .B1(n6924), .B2(n6923), .A(n6641), .ZN(n6922) );
  INV_X1 U7733 ( .A(n6633), .ZN(n6923) );
  OAI21_X1 U7734 ( .B1(n8659), .B2(n6936), .A(n6934), .ZN(n8705) );
  AOI21_X1 U7735 ( .B1(n6937), .B2(n6935), .A(n6639), .ZN(n6934) );
  INV_X1 U7736 ( .A(n6937), .ZN(n6936) );
  INV_X1 U7737 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n9304) );
  NAND2_X1 U7738 ( .A1(n8545), .A2(n8544), .ZN(n8564) );
  OAI21_X2 U7739 ( .B1(n6714), .B2(n6716), .A(n6884), .ZN(n8275) );
  NAND2_X1 U7740 ( .A1(n6886), .A2(n6717), .ZN(n6716) );
  AOI21_X1 U7741 ( .B1(n6886), .B2(n6888), .A(n6578), .ZN(n6884) );
  NOR2_X1 U7742 ( .A1(n8209), .A2(n6718), .ZN(n6714) );
  OAI21_X1 U7743 ( .B1(n8965), .B2(n8964), .A(n7099), .ZN(n7098) );
  NAND2_X1 U7744 ( .A1(n10224), .A2(P3_ADDR_REG_9__SCAN_IN), .ZN(n7099) );
  NOR2_X1 U7745 ( .A1(n8973), .A2(n8972), .ZN(n8914) );
  AOI21_X1 U7746 ( .B1(n7016), .B2(n9244), .A(n6576), .ZN(n7013) );
  OR2_X1 U7747 ( .A1(n12483), .A2(n9244), .ZN(n7014) );
  INV_X1 U7748 ( .A(n9232), .ZN(n7039) );
  AND2_X1 U7749 ( .A1(n9245), .A2(n7017), .ZN(n7016) );
  OR2_X1 U7750 ( .A1(n12483), .A2(n9244), .ZN(n7017) );
  AND2_X1 U7751 ( .A1(n7740), .A2(n9134), .ZN(n7751) );
  NAND2_X1 U7752 ( .A1(n7751), .A2(n12367), .ZN(n7762) );
  NOR2_X1 U7753 ( .A1(n12490), .A2(n12332), .ZN(n7027) );
  INV_X1 U7754 ( .A(n12492), .ZN(n7030) );
  NOR2_X1 U7755 ( .A1(n12399), .A2(n7027), .ZN(n7026) );
  BUF_X1 U7756 ( .A(n9178), .Z(n9242) );
  INV_X1 U7757 ( .A(n12406), .ZN(n7021) );
  AOI21_X1 U7758 ( .B1(n7026), .B2(n7031), .A(n7023), .ZN(n7022) );
  INV_X1 U7759 ( .A(n12397), .ZN(n7023) );
  NAND2_X1 U7760 ( .A1(n7067), .A2(n12724), .ZN(n12694) );
  AND4_X1 U7761 ( .A1(n12519), .A2(n7914), .A3(n7913), .A4(n7912), .ZN(n11677)
         );
  AND4_X1 U7762 ( .A1(n7798), .A2(n7797), .A3(n7796), .A4(n7795), .ZN(n12389)
         );
  AND4_X1 U7763 ( .A1(n7782), .A2(n7781), .A3(n7780), .A4(n7779), .ZN(n12450)
         );
  NAND2_X1 U7764 ( .A1(n15042), .A2(n15043), .ZN(n15041) );
  XNOR2_X1 U7765 ( .A(n10080), .B(n15069), .ZN(n15067) );
  NAND2_X1 U7766 ( .A1(n15041), .A2(n6871), .ZN(n10080) );
  NAND2_X1 U7767 ( .A1(n15051), .A2(P3_REG1_REG_4__SCAN_IN), .ZN(n6871) );
  XNOR2_X1 U7768 ( .A(n10272), .B(n10269), .ZN(n10161) );
  NOR2_X1 U7769 ( .A1(n10160), .A2(n10095), .ZN(n7205) );
  NAND2_X1 U7770 ( .A1(n10276), .A2(n10277), .ZN(n10698) );
  NOR2_X1 U7771 ( .A1(n10699), .A2(n10264), .ZN(n6688) );
  XNOR2_X1 U7772 ( .A(n10700), .B(n10714), .ZN(n15096) );
  NAND2_X1 U7773 ( .A1(n11146), .A2(n11147), .ZN(n11148) );
  NAND2_X1 U7774 ( .A1(n11148), .A2(n11149), .ZN(n12769) );
  AND2_X1 U7775 ( .A1(n12773), .A2(P3_REG2_REG_12__SCAN_IN), .ZN(n7211) );
  INV_X1 U7776 ( .A(n12858), .ZN(n6882) );
  NAND2_X1 U7777 ( .A1(n7193), .A2(P3_REG2_REG_17__SCAN_IN), .ZN(n7192) );
  XNOR2_X1 U7778 ( .A(n12922), .B(n12389), .ZN(n12916) );
  NAND2_X1 U7779 ( .A1(n7898), .A2(n7329), .ZN(n7328) );
  NOR2_X1 U7780 ( .A1(n7900), .A2(n7330), .ZN(n7329) );
  INV_X1 U7781 ( .A(n7897), .ZN(n7330) );
  AND2_X1 U7782 ( .A1(n12669), .A2(n12661), .ZN(n12930) );
  AOI21_X1 U7783 ( .B1(n12545), .B2(n12752), .A(n6810), .ZN(n7899) );
  INV_X1 U7784 ( .A(n12961), .ZN(n6810) );
  INV_X1 U7785 ( .A(n12752), .ZN(n12973) );
  NAND2_X1 U7786 ( .A1(n7898), .A2(n7897), .ZN(n12972) );
  OR2_X1 U7787 ( .A1(n7681), .A2(n7680), .ZN(n7682) );
  AOI21_X1 U7788 ( .B1(n7340), .B2(n7339), .A(n6559), .ZN(n7338) );
  INV_X1 U7789 ( .A(n6519), .ZN(n7339) );
  OR2_X1 U7790 ( .A1(n13231), .A2(n13051), .ZN(n13024) );
  NAND2_X1 U7791 ( .A1(n7336), .A2(n7334), .ZN(n11077) );
  NAND2_X1 U7792 ( .A1(n10892), .A2(n10891), .ZN(n7336) );
  NAND2_X1 U7793 ( .A1(n11076), .A2(n12707), .ZN(n11075) );
  NAND2_X1 U7794 ( .A1(n6840), .A2(n12570), .ZN(n10519) );
  NAND2_X1 U7795 ( .A1(n7864), .A2(n7962), .ZN(n15120) );
  NOR2_X1 U7796 ( .A1(n9767), .A2(n15170), .ZN(n10028) );
  AND2_X1 U7797 ( .A1(n7917), .A2(n12689), .ZN(n13100) );
  OR2_X1 U7798 ( .A1(n8891), .A2(n15115), .ZN(n8892) );
  NAND2_X1 U7799 ( .A1(n7326), .A2(n7905), .ZN(n8890) );
  INV_X1 U7800 ( .A(n13007), .ZN(n6843) );
  OR2_X1 U7801 ( .A1(n7448), .A2(n9441), .ZN(n7434) );
  OR2_X1 U7802 ( .A1(n7462), .A2(n9442), .ZN(n7435) );
  INV_X1 U7803 ( .A(n13100), .ZN(n15111) );
  OR2_X1 U7804 ( .A1(n12739), .A2(n12547), .ZN(n15170) );
  AND2_X1 U7805 ( .A1(n7929), .A2(n7951), .ZN(n9525) );
  OAI22_X1 U7806 ( .A1(n11644), .A2(n11643), .B1(P2_DATAO_REG_29__SCAN_IN), 
        .B2(n11663), .ZN(n12509) );
  NOR2_X1 U7807 ( .A1(P3_IR_REG_27__SCAN_IN), .A2(P3_IR_REG_26__SCAN_IN), .ZN(
        n7323) );
  NAND2_X1 U7808 ( .A1(n7799), .A2(n7788), .ZN(n7800) );
  NAND2_X1 U7809 ( .A1(n7745), .A2(n7744), .ZN(n7748) );
  AND2_X1 U7810 ( .A1(n7851), .A2(n7850), .ZN(n7853) );
  OR2_X1 U7811 ( .A1(n7736), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n7745) );
  AND2_X1 U7812 ( .A1(n7717), .A2(n7704), .ZN(n7705) );
  AOI21_X1 U7813 ( .B1(n7055), .B2(n7057), .A(n7054), .ZN(n7053) );
  INV_X1 U7814 ( .A(n7703), .ZN(n7054) );
  AND2_X1 U7815 ( .A1(n7684), .A2(n7663), .ZN(n7664) );
  NAND2_X1 U7816 ( .A1(n7662), .A2(n7661), .ZN(n7665) );
  NAND2_X1 U7817 ( .A1(n7665), .A2(n7664), .ZN(n7685) );
  NAND2_X1 U7818 ( .A1(n7647), .A2(n7646), .ZN(n7662) );
  AND2_X1 U7819 ( .A1(n7644), .A2(n7629), .ZN(n7642) );
  NAND2_X1 U7820 ( .A1(n6808), .A2(P1_DATAO_REG_13__SCAN_IN), .ZN(n7628) );
  NOR2_X1 U7821 ( .A1(n7604), .A2(n7603), .ZN(n7614) );
  INV_X1 U7822 ( .A(P3_IR_REG_12__SCAN_IN), .ZN(n7613) );
  AND2_X1 U7823 ( .A1(n7581), .A2(n7565), .ZN(n7566) );
  NAND2_X1 U7824 ( .A1(n7564), .A2(n7563), .ZN(n7567) );
  NAND2_X1 U7825 ( .A1(n7567), .A2(n7566), .ZN(n7582) );
  AND2_X1 U7826 ( .A1(n7483), .A2(n7465), .ZN(n7481) );
  NAND2_X1 U7827 ( .A1(n7464), .A2(n7463), .ZN(n7482) );
  NAND2_X1 U7828 ( .A1(n7446), .A2(n7445), .ZN(n7464) );
  NAND2_X1 U7829 ( .A1(n6686), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n6685) );
  OR2_X1 U7830 ( .A1(n12157), .A2(n12156), .ZN(n7357) );
  NOR2_X1 U7831 ( .A1(n11215), .A2(n11216), .ZN(n7002) );
  INV_X1 U7832 ( .A(n13377), .ZN(n13305) );
  OR2_X1 U7833 ( .A1(n8598), .A2(n8597), .ZN(n8618) );
  AND2_X1 U7834 ( .A1(n11763), .A2(n10548), .ZN(n6998) );
  NOR2_X1 U7835 ( .A1(n11096), .A2(n7004), .ZN(n7003) );
  INV_X1 U7836 ( .A(n7005), .ZN(n7004) );
  NAND2_X1 U7837 ( .A1(n10840), .A2(n10839), .ZN(n11090) );
  NAND2_X1 U7838 ( .A1(n6530), .A2(n8827), .ZN(n8858) );
  AOI21_X1 U7839 ( .B1(P2_REG1_REG_14__SCAN_IN), .B2(n14889), .A(n14883), .ZN(
        n10927) );
  NOR2_X1 U7840 ( .A1(n13498), .A2(n13700), .ZN(n6946) );
  NAND2_X1 U7841 ( .A1(n6486), .A2(n6491), .ZN(n6711) );
  NAND2_X1 U7842 ( .A1(n6710), .A2(n6491), .ZN(n6709) );
  AND2_X1 U7843 ( .A1(n8765), .A2(n8693), .ZN(n13524) );
  NOR2_X1 U7844 ( .A1(n12136), .A2(n7147), .ZN(n7146) );
  INV_X1 U7845 ( .A(n13683), .ZN(n12133) );
  NAND2_X1 U7846 ( .A1(n12133), .A2(n12132), .ZN(n13681) );
  AND2_X1 U7847 ( .A1(n13636), .A2(n8831), .ZN(n13652) );
  NAND2_X1 U7848 ( .A1(n6721), .A2(n6495), .ZN(n13650) );
  NAND2_X1 U7849 ( .A1(n6954), .A2(n6953), .ZN(n13672) );
  AND2_X1 U7850 ( .A1(n7128), .A2(n11300), .ZN(n7127) );
  NAND2_X1 U7851 ( .A1(n11299), .A2(n7129), .ZN(n7128) );
  INV_X1 U7852 ( .A(n11298), .ZN(n7129) );
  NAND2_X1 U7853 ( .A1(n6757), .A2(n11299), .ZN(n7126) );
  INV_X1 U7854 ( .A(n6719), .ZN(n11360) );
  AOI21_X1 U7855 ( .B1(n6497), .B2(n7136), .A(n6586), .ZN(n7135) );
  NAND2_X1 U7856 ( .A1(n6497), .A2(n6754), .ZN(n6753) );
  AND2_X1 U7857 ( .A1(n11125), .A2(n7173), .ZN(n7171) );
  NAND2_X1 U7858 ( .A1(n6755), .A2(n10859), .ZN(n11121) );
  NOR2_X1 U7859 ( .A1(n14995), .A2(n13388), .ZN(n7178) );
  NAND2_X1 U7860 ( .A1(n7174), .A2(n7173), .ZN(n7172) );
  NOR2_X2 U7861 ( .A1(n10786), .A2(n10854), .ZN(n10864) );
  INV_X1 U7862 ( .A(n6751), .ZN(n6750) );
  OAI21_X1 U7863 ( .B1(n7131), .B2(n6752), .A(n11498), .ZN(n6751) );
  INV_X1 U7864 ( .A(n10618), .ZN(n6752) );
  NAND2_X1 U7865 ( .A1(n10370), .A2(n10320), .ZN(n7130) );
  INV_X1 U7866 ( .A(n10627), .ZN(n11498) );
  NAND2_X1 U7867 ( .A1(n7130), .A2(n7131), .ZN(n10619) );
  NAND2_X1 U7868 ( .A1(n7134), .A2(n10373), .ZN(n10368) );
  INV_X1 U7869 ( .A(n10370), .ZN(n7134) );
  XNOR2_X1 U7870 ( .A(n13395), .B(n13270), .ZN(n10179) );
  XNOR2_X1 U7871 ( .A(n8841), .B(n9953), .ZN(n9948) );
  AND2_X1 U7872 ( .A1(n9824), .A2(n8823), .ZN(n13640) );
  INV_X1 U7873 ( .A(n13657), .ZN(n13642) );
  AND2_X1 U7874 ( .A1(n14988), .A2(n13490), .ZN(n9912) );
  AND2_X1 U7875 ( .A1(n13711), .A2(n14986), .ZN(n13712) );
  AOI21_X1 U7876 ( .B1(n13546), .B2(n6499), .A(n12142), .ZN(n13523) );
  AND2_X1 U7877 ( .A1(n9797), .A2(n9800), .ZN(n14928) );
  AND2_X1 U7878 ( .A1(n9273), .A2(n9641), .ZN(n10046) );
  INV_X1 U7879 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n7221) );
  NAND4_X1 U7880 ( .A1(n8254), .A2(n7980), .A3(n7985), .A4(n6526), .ZN(n8814)
         );
  NAND2_X1 U7881 ( .A1(n8804), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8817) );
  OR2_X1 U7882 ( .A1(n8803), .A2(P2_IR_REG_22__SCAN_IN), .ZN(n8804) );
  AND2_X1 U7883 ( .A1(n13889), .A2(n12257), .ZN(n13837) );
  AND2_X1 U7884 ( .A1(n13826), .A2(n7105), .ZN(n7104) );
  OR2_X1 U7885 ( .A1(n13953), .A2(n12292), .ZN(n7105) );
  NAND2_X1 U7886 ( .A1(n6770), .A2(n6769), .ZN(n10644) );
  NAND2_X1 U7887 ( .A1(n6772), .A2(n10338), .ZN(n6770) );
  AOI21_X1 U7888 ( .B1(n13940), .B2(n6787), .A(n6786), .ZN(n11225) );
  AND2_X1 U7889 ( .A1(n7112), .A2(n6788), .ZN(n6787) );
  INV_X1 U7890 ( .A(n7110), .ZN(n6786) );
  NOR2_X1 U7891 ( .A1(n7117), .A2(n6548), .ZN(n7116) );
  NOR3_X1 U7892 ( .A1(n12220), .A2(n7119), .A3(n7118), .ZN(n7117) );
  NAND2_X1 U7893 ( .A1(n11437), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n11475) );
  OR2_X1 U7894 ( .A1(n12246), .A2(n12245), .ZN(n13833) );
  XNOR2_X1 U7895 ( .A(n9383), .B(n9384), .ZN(n13923) );
  NAND2_X1 U7896 ( .A1(n13922), .A2(n13923), .ZN(n13921) );
  NAND2_X1 U7897 ( .A1(n13952), .A2(n13953), .ZN(n13951) );
  NAND2_X1 U7898 ( .A1(n12183), .A2(n12182), .ZN(n12189) );
  OR2_X1 U7899 ( .A1(n12181), .A2(n12180), .ZN(n12182) );
  NAND2_X1 U7900 ( .A1(n6660), .A2(n7296), .ZN(n11951) );
  OR3_X1 U7901 ( .A1(n9387), .A2(n12150), .A3(n9389), .ZN(n9412) );
  OR2_X1 U7902 ( .A1(n9855), .A2(n9854), .ZN(n7076) );
  OR2_X1 U7903 ( .A1(n9979), .A2(n9978), .ZN(n7072) );
  AND2_X1 U7904 ( .A1(n7072), .A2(n7071), .ZN(n10229) );
  NAND2_X1 U7905 ( .A1(n10462), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n7071) );
  OR2_X1 U7906 ( .A1(n10229), .A2(n10228), .ZN(n7070) );
  NOR2_X1 U7907 ( .A1(n11403), .A2(n7077), .ZN(n14568) );
  AND2_X1 U7908 ( .A1(n11411), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n7077) );
  NOR2_X1 U7909 ( .A1(n14568), .A2(n14567), .ZN(n14566) );
  OR2_X1 U7910 ( .A1(n9611), .A2(P1_IR_REG_11__SCAN_IN), .ZN(n9612) );
  NOR2_X1 U7911 ( .A1(n14592), .A2(n6629), .ZN(n14608) );
  NAND2_X1 U7912 ( .A1(n14610), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n7078) );
  NAND2_X1 U7913 ( .A1(n14606), .A2(n6870), .ZN(n14035) );
  OR2_X1 U7914 ( .A1(n14610), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n6870) );
  OR2_X1 U7915 ( .A1(n14619), .A2(n14618), .ZN(n6861) );
  AND2_X1 U7916 ( .A1(n6861), .A2(n6860), .ZN(n14630) );
  NAND2_X1 U7917 ( .A1(n14625), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n6860) );
  OR2_X1 U7918 ( .A1(n14630), .A2(n14631), .ZN(n6859) );
  OR2_X1 U7919 ( .A1(n10310), .A2(P1_IR_REG_17__SCAN_IN), .ZN(n10679) );
  XNOR2_X1 U7920 ( .A(n14031), .B(n14043), .ZN(n14654) );
  NOR2_X1 U7921 ( .A1(n14654), .A2(n14653), .ZN(n14652) );
  NAND2_X1 U7922 ( .A1(n11971), .A2(n11970), .ZN(n12045) );
  INV_X1 U7923 ( .A(n6736), .ZN(n6732) );
  AOI21_X1 U7924 ( .B1(n6738), .B2(n6737), .A(n6560), .ZN(n6736) );
  INV_X1 U7925 ( .A(n6520), .ZN(n6737) );
  NAND2_X1 U7926 ( .A1(n6738), .A2(n6734), .ZN(n6733) );
  AND2_X1 U7927 ( .A1(n11612), .A2(n12026), .ZN(n6734) );
  NAND2_X1 U7928 ( .A1(n14088), .A2(n14093), .ZN(n14089) );
  NAND2_X1 U7929 ( .A1(n7268), .A2(n7263), .ZN(n7261) );
  NAND2_X1 U7930 ( .A1(n7250), .A2(n14138), .ZN(n14139) );
  NAND3_X1 U7931 ( .A1(n6498), .A2(n14162), .A3(n11387), .ZN(n14158) );
  NAND2_X1 U7932 ( .A1(n11490), .A2(n11491), .ZN(n7276) );
  INV_X1 U7933 ( .A(n11473), .ZN(n7246) );
  AOI21_X1 U7934 ( .B1(n7288), .B2(n7290), .A(n6569), .ZN(n6692) );
  NAND2_X1 U7935 ( .A1(n6626), .A2(n7288), .ZN(n6691) );
  INV_X1 U7936 ( .A(n12015), .ZN(n11261) );
  AOI21_X1 U7937 ( .B1(n7239), .B2(n12011), .A(n11167), .ZN(n7237) );
  NAND2_X1 U7938 ( .A1(n11054), .A2(n7239), .ZN(n6729) );
  NAND2_X1 U7939 ( .A1(n6626), .A2(n11167), .ZN(n11197) );
  INV_X1 U7940 ( .A(n6700), .ZN(n6699) );
  NAND2_X1 U7941 ( .A1(n11054), .A2(n10995), .ZN(n7238) );
  AND2_X1 U7942 ( .A1(n12008), .A2(n7286), .ZN(n7285) );
  OR2_X1 U7943 ( .A1(n14479), .A2(n7287), .ZN(n7286) );
  NAND2_X1 U7944 ( .A1(n6742), .A2(n7256), .ZN(n14473) );
  AND2_X1 U7945 ( .A1(n7255), .A2(n10958), .ZN(n6742) );
  NAND2_X1 U7946 ( .A1(n10566), .A2(n10565), .ZN(n14667) );
  NAND2_X1 U7947 ( .A1(n14682), .A2(n14687), .ZN(n10460) );
  NAND2_X1 U7948 ( .A1(n7254), .A2(n12002), .ZN(n14684) );
  INV_X1 U7949 ( .A(n14686), .ZN(n7254) );
  INV_X1 U7950 ( .A(n11779), .ZN(n9746) );
  NAND2_X1 U7951 ( .A1(n9668), .A2(n10400), .ZN(n14777) );
  AND2_X1 U7952 ( .A1(n9392), .A2(n9483), .ZN(n10394) );
  XNOR2_X1 U7953 ( .A(n8723), .B(n6647), .ZN(n11961) );
  NAND2_X1 U7954 ( .A1(n6920), .A2(n6922), .ZN(n8723) );
  NAND2_X1 U7955 ( .A1(n6921), .A2(n6924), .ZN(n6920) );
  INV_X1 U7956 ( .A(n8760), .ZN(n6921) );
  NOR2_X1 U7957 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_26__SCAN_IN), .ZN(
        n6774) );
  AND2_X1 U7958 ( .A1(n9288), .A2(n9292), .ZN(n7121) );
  INV_X1 U7959 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n9285) );
  OAI21_X1 U7960 ( .B1(n9519), .B2(P1_IR_REG_8__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n9571) );
  XNOR2_X1 U7961 ( .A(n8252), .B(n8250), .ZN(n10562) );
  NAND2_X1 U7962 ( .A1(n6885), .A2(n8233), .ZN(n8252) );
  NAND2_X1 U7963 ( .A1(n8231), .A2(n8230), .ZN(n6885) );
  OR2_X1 U7964 ( .A1(n9513), .A2(P1_IR_REG_7__SCAN_IN), .ZN(n9519) );
  INV_X1 U7965 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n7074) );
  NAND2_X1 U7966 ( .A1(n6814), .A2(n6616), .ZN(n7094) );
  INV_X1 U7967 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n8901) );
  XNOR2_X1 U7968 ( .A(n8930), .B(P1_ADDR_REG_4__SCAN_IN), .ZN(n8931) );
  INV_X1 U7969 ( .A(n6817), .ZN(n8950) );
  OAI21_X1 U7970 ( .B1(n15196), .B2(P2_ADDR_REG_5__SCAN_IN), .A(n6563), .ZN(
        n6817) );
  INV_X1 U7971 ( .A(n6826), .ZN(n8961) );
  OAI21_X1 U7972 ( .B1(n15201), .B2(n15200), .A(n6580), .ZN(n6826) );
  OAI21_X1 U7973 ( .B1(n8966), .B2(n14852), .A(n14324), .ZN(n8970) );
  NOR2_X1 U7974 ( .A1(n8927), .A2(n8926), .ZN(n8918) );
  OAI21_X1 U7975 ( .B1(n6836), .B2(n6834), .A(n8985), .ZN(n6833) );
  NAND2_X1 U7976 ( .A1(n7033), .A2(n7032), .ZN(n12328) );
  NAND2_X1 U7977 ( .A1(n6589), .A2(n6488), .ZN(n7032) );
  INV_X1 U7978 ( .A(n13099), .ZN(n12352) );
  NAND2_X1 U7979 ( .A1(n11042), .A2(n11041), .ZN(n11040) );
  OR2_X1 U7980 ( .A1(n9221), .A2(n13003), .ZN(n9222) );
  NAND2_X1 U7981 ( .A1(n7761), .A2(n7760), .ZN(n12954) );
  NAND2_X1 U7982 ( .A1(n7710), .A2(n7709), .ZN(n13004) );
  INV_X1 U7983 ( .A(n12500), .ZN(n12476) );
  OR2_X1 U7984 ( .A1(n9260), .A2(n9259), .ZN(n12497) );
  NAND2_X1 U7985 ( .A1(n7769), .A2(n7768), .ZN(n12751) );
  INV_X1 U7986 ( .A(n12332), .ZN(n13051) );
  AND2_X1 U7987 ( .A1(n7460), .A2(n7457), .ZN(n6661) );
  AND2_X1 U7988 ( .A1(n10122), .A2(n9775), .ZN(n9776) );
  NAND2_X1 U7989 ( .A1(n10082), .A2(n10083), .ZN(n10159) );
  NOR2_X1 U7990 ( .A1(n12765), .A2(n12737), .ZN(n15064) );
  INV_X1 U7991 ( .A(n12840), .ZN(n14394) );
  XNOR2_X1 U7992 ( .A(n12719), .B(n12505), .ZN(n12872) );
  NAND2_X1 U7993 ( .A1(n6962), .A2(n12539), .ZN(n8885) );
  NAND2_X1 U7994 ( .A1(n11666), .A2(n12520), .ZN(n7040) );
  NAND2_X1 U7995 ( .A1(n7694), .A2(n7693), .ZN(n13226) );
  AND2_X1 U7996 ( .A1(n6994), .A2(n6506), .ZN(n10769) );
  NAND2_X1 U7997 ( .A1(n8311), .A2(n8310), .ZN(n11730) );
  NOR2_X1 U7998 ( .A1(n13331), .A2(n13314), .ZN(n6992) );
  NAND2_X1 U7999 ( .A1(n6993), .A2(n6550), .ZN(n6991) );
  XNOR2_X1 U8000 ( .A(n11706), .B(n10347), .ZN(n10044) );
  NAND2_X1 U8001 ( .A1(n8838), .A2(n10216), .ZN(n10001) );
  NAND2_X1 U8002 ( .A1(n13277), .A2(n11748), .ZN(n11749) );
  OR2_X1 U8003 ( .A1(n11750), .A2(n11747), .ZN(n11748) );
  INV_X1 U8004 ( .A(n13392), .ZN(n11766) );
  NAND2_X1 U8005 ( .A1(n8577), .A2(n8576), .ZN(n13625) );
  NAND2_X1 U8006 ( .A1(n8719), .A2(n8718), .ZN(n13694) );
  NAND2_X1 U8007 ( .A1(n6712), .A2(n6486), .ZN(n13519) );
  NAND2_X1 U8008 ( .A1(n13531), .A2(n13538), .ZN(n6712) );
  INV_X1 U8009 ( .A(n13987), .ZN(n11234) );
  OAI22_X1 U8010 ( .A1(n11227), .A2(n11226), .B1(n11225), .B2(n11111), .ZN(
        n11339) );
  NAND2_X1 U8011 ( .A1(n6780), .A2(n6781), .ZN(n11351) );
  XNOR2_X1 U8012 ( .A(n11225), .B(n11111), .ZN(n11227) );
  NAND2_X1 U8013 ( .A1(n11566), .A2(n11565), .ZN(n14221) );
  XNOR2_X1 U8014 ( .A(n9582), .B(P1_REG2_REG_1__SCAN_IN), .ZN(n14002) );
  NOR2_X1 U8015 ( .A1(n14017), .A2(n6533), .ZN(n9585) );
  AND2_X1 U8016 ( .A1(n7070), .A2(n7069), .ZN(n10532) );
  NAND2_X1 U8017 ( .A1(n10563), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n7069) );
  INV_X1 U8018 ( .A(n14098), .ZN(n6689) );
  NAND2_X1 U8019 ( .A1(n14130), .A2(n11542), .ZN(n14114) );
  NAND2_X1 U8020 ( .A1(n14207), .A2(n14701), .ZN(n7230) );
  AND2_X1 U8021 ( .A1(n8970), .A2(n8969), .ZN(n14328) );
  NAND2_X1 U8022 ( .A1(n6823), .A2(n7089), .ZN(n14552) );
  NAND2_X1 U8023 ( .A1(n6825), .A2(n6824), .ZN(n6823) );
  AND2_X1 U8024 ( .A1(n7088), .A2(n6535), .ZN(n6824) );
  NOR2_X1 U8025 ( .A1(n14551), .A2(n14552), .ZN(n14550) );
  NAND2_X1 U8026 ( .A1(n8979), .A2(n14893), .ZN(n6828) );
  NAND2_X1 U8027 ( .A1(n8987), .A2(P2_ADDR_REG_18__SCAN_IN), .ZN(n6664) );
  AND2_X1 U8028 ( .A1(n14340), .A2(n7085), .ZN(n7082) );
  INV_X1 U8029 ( .A(n9755), .ZN(n11787) );
  NOR2_X1 U8030 ( .A1(n8041), .A2(n8040), .ZN(n8045) );
  AND2_X1 U8031 ( .A1(n8836), .A2(n8069), .ZN(n8041) );
  NAND2_X1 U8032 ( .A1(n11814), .A2(n11816), .ZN(n7311) );
  OR2_X1 U8033 ( .A1(n8172), .A2(n8173), .ZN(n7218) );
  INV_X1 U8034 ( .A(n11835), .ZN(n7303) );
  NAND2_X1 U8035 ( .A1(n11846), .A2(n11848), .ZN(n7302) );
  NAND2_X1 U8036 ( .A1(n7222), .A2(n7225), .ZN(n8268) );
  NAND2_X1 U8037 ( .A1(n8249), .A2(n6544), .ZN(n7225) );
  INV_X1 U8038 ( .A(n8268), .ZN(n6656) );
  INV_X1 U8039 ( .A(n8267), .ZN(n6655) );
  NOR2_X1 U8040 ( .A1(n6567), .A2(n7314), .ZN(n7312) );
  INV_X1 U8041 ( .A(n11868), .ZN(n7314) );
  NAND2_X1 U8042 ( .A1(n11909), .A2(n7319), .ZN(n7318) );
  NAND2_X1 U8043 ( .A1(n8502), .A2(n6601), .ZN(n6681) );
  NAND2_X1 U8044 ( .A1(n8562), .A2(n6602), .ZN(n6683) );
  NAND2_X1 U8045 ( .A1(n11929), .A2(n11927), .ZN(n7307) );
  NAND2_X1 U8046 ( .A1(n7227), .A2(n7228), .ZN(n8632) );
  NAND2_X1 U8047 ( .A1(n6525), .A2(n6500), .ZN(n7228) );
  NAND2_X1 U8048 ( .A1(n7322), .A2(n11938), .ZN(n7321) );
  INV_X1 U8049 ( .A(n6931), .ZN(n6930) );
  INV_X1 U8050 ( .A(n8509), .ZN(n6927) );
  INV_X1 U8051 ( .A(P3_IR_REG_25__SCAN_IN), .ZN(n7383) );
  INV_X1 U8052 ( .A(P3_IR_REG_16__SCAN_IN), .ZN(n6983) );
  INV_X1 U8053 ( .A(n7783), .ZN(n7059) );
  INV_X1 U8054 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n8416) );
  INV_X1 U8055 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n8337) );
  OR2_X1 U8056 ( .A1(n8338), .A2(n8337), .ZN(n8417) );
  NAND2_X1 U8057 ( .A1(n14216), .A2(n12309), .ZN(n6740) );
  INV_X1 U8058 ( .A(n10446), .ZN(n6697) );
  INV_X1 U8059 ( .A(n10459), .ZN(n7271) );
  AND2_X1 U8060 ( .A1(n6744), .A2(n11602), .ZN(n6743) );
  OR2_X1 U8061 ( .A1(n6518), .A2(n6745), .ZN(n6744) );
  INV_X1 U8062 ( .A(n11900), .ZN(n6745) );
  NOR2_X1 U8063 ( .A1(n11899), .A2(n14270), .ZN(n6915) );
  INV_X1 U8064 ( .A(n8665), .ZN(n6935) );
  NAND2_X1 U8065 ( .A1(n8460), .A2(SI_17_), .ZN(n6931) );
  NOR2_X1 U8066 ( .A1(n8460), .A2(SI_17_), .ZN(n6932) );
  AOI21_X1 U8067 ( .B1(n6492), .B2(n6487), .A(n6573), .ZN(n6892) );
  INV_X1 U8068 ( .A(n8211), .ZN(n6718) );
  INV_X1 U8069 ( .A(n6887), .ZN(n6886) );
  NAND2_X1 U8070 ( .A1(n8207), .A2(n8211), .ZN(n6717) );
  INV_X1 U8071 ( .A(P3_ADDR_REG_19__SCAN_IN), .ZN(n7401) );
  NOR2_X2 U8072 ( .A1(n12448), .A2(n9231), .ZN(n9233) );
  INV_X1 U8073 ( .A(n13087), .ZN(n9205) );
  NAND2_X1 U8074 ( .A1(n15051), .A2(P3_REG2_REG_4__SCAN_IN), .ZN(n7183) );
  INV_X1 U8075 ( .A(n14372), .ZN(n7199) );
  INV_X1 U8076 ( .A(n7203), .ZN(n7202) );
  NOR2_X1 U8077 ( .A1(n7200), .A2(n7199), .ZN(n7197) );
  NAND2_X1 U8078 ( .A1(n7202), .A2(n14379), .ZN(n7200) );
  NAND2_X1 U8079 ( .A1(n14367), .A2(n12847), .ZN(n12849) );
  AND2_X1 U8080 ( .A1(n12534), .A2(n6964), .ZN(n6963) );
  NAND2_X1 U8081 ( .A1(n6965), .A2(n12539), .ZN(n6964) );
  INV_X1 U8082 ( .A(n12540), .ZN(n6965) );
  INV_X1 U8083 ( .A(n12539), .ZN(n6966) );
  NAND2_X1 U8084 ( .A1(n6976), .A2(n12667), .ZN(n6975) );
  INV_X1 U8085 ( .A(n6978), .ZN(n6976) );
  NOR2_X1 U8086 ( .A1(P3_REG3_REG_22__SCAN_IN), .A2(n7762), .ZN(n7776) );
  OR2_X1 U8087 ( .A1(n12954), .A2(n7770), .ZN(n12660) );
  OR2_X1 U8088 ( .A1(n13226), .A2(n12756), .ZN(n12638) );
  INV_X1 U8089 ( .A(n7889), .ZN(n7341) );
  INV_X1 U8090 ( .A(n12595), .ZN(n6971) );
  INV_X1 U8091 ( .A(n6970), .ZN(n6969) );
  OAI21_X1 U8092 ( .B1(n12707), .B2(n6971), .A(n12599), .ZN(n6970) );
  AOI21_X1 U8093 ( .B1(n6511), .B2(n6797), .A(n6791), .ZN(n6790) );
  INV_X1 U8094 ( .A(n7041), .ZN(n6791) );
  NAND2_X1 U8095 ( .A1(n7735), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n7744) );
  INV_X1 U8096 ( .A(n7053), .ZN(n6797) );
  INV_X1 U8097 ( .A(P3_IR_REG_7__SCAN_IN), .ZN(n7529) );
  INV_X1 U8098 ( .A(n6713), .ZN(n6710) );
  AOI21_X1 U8099 ( .B1(n12118), .B2(n6486), .A(n13518), .ZN(n6713) );
  OR2_X1 U8100 ( .A1(n13706), .A2(n8828), .ZN(n12119) );
  OAI21_X1 U8101 ( .B1(n7146), .B2(n7144), .A(n12137), .ZN(n7143) );
  NAND2_X1 U8102 ( .A1(n8489), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n8518) );
  AND2_X1 U8103 ( .A1(n8378), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n8365) );
  NOR2_X1 U8104 ( .A1(n8417), .A2(n8416), .ZN(n8398) );
  AND2_X1 U8105 ( .A1(n8398), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n8378) );
  INV_X1 U8106 ( .A(n10859), .ZN(n6754) );
  INV_X1 U8107 ( .A(n6521), .ZN(n7136) );
  INV_X1 U8108 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n8258) );
  INV_X1 U8109 ( .A(n10372), .ZN(n7157) );
  NOR2_X1 U8110 ( .A1(n7157), .A2(n7158), .ZN(n7156) );
  INV_X1 U8111 ( .A(n6760), .ZN(n7158) );
  NAND2_X1 U8112 ( .A1(n8837), .A2(n9922), .ZN(n9915) );
  NAND2_X1 U8113 ( .A1(n6950), .A2(n10317), .ZN(n10381) );
  INV_X1 U8114 ( .A(n10323), .ZN(n6950) );
  OR2_X1 U8115 ( .A1(n8158), .A2(n8157), .ZN(n8181) );
  INV_X1 U8116 ( .A(n10747), .ZN(n7111) );
  INV_X1 U8117 ( .A(n12207), .ZN(n7118) );
  NAND2_X1 U8118 ( .A1(n11948), .A2(n7297), .ZN(n7296) );
  INV_X1 U8119 ( .A(n11609), .ZN(n7267) );
  NOR2_X1 U8120 ( .A1(n12184), .A2(n6913), .ZN(n6912) );
  INV_X1 U8121 ( .A(n6914), .ZN(n6913) );
  NOR2_X1 U8122 ( .A1(n14442), .A2(n11858), .ZN(n6914) );
  INV_X1 U8123 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n10571) );
  NAND2_X1 U8124 ( .A1(n11965), .A2(n11972), .ZN(n11781) );
  NAND2_X1 U8125 ( .A1(n11387), .A2(n6915), .ZN(n11485) );
  NAND2_X1 U8126 ( .A1(n11387), .A2(n12209), .ZN(n11435) );
  NAND2_X1 U8127 ( .A1(n14473), .A2(n10959), .ZN(n10961) );
  NAND2_X1 U8128 ( .A1(n6905), .A2(n6904), .ZN(n14711) );
  INV_X1 U8129 ( .A(n8741), .ZN(n6925) );
  XNOR2_X1 U8130 ( .A(n8355), .B(SI_16_), .ZN(n8374) );
  AND2_X1 U8131 ( .A1(n8353), .A2(n8352), .ZN(n8389) );
  NOR2_X1 U8132 ( .A1(n7353), .A2(n6554), .ZN(n6938) );
  XNOR2_X1 U8133 ( .A(n8330), .B(SI_12_), .ZN(n8326) );
  NAND2_X1 U8134 ( .A1(n8280), .A2(n8279), .ZN(n8328) );
  NAND2_X1 U8135 ( .A1(n8209), .A2(n8208), .ZN(n6715) );
  INV_X1 U8136 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n9468) );
  NOR2_X1 U8137 ( .A1(n9316), .A2(P1_IR_REG_4__SCAN_IN), .ZN(n9469) );
  XNOR2_X1 U8138 ( .A(n8137), .B(n6708), .ZN(n8135) );
  INV_X1 U8139 ( .A(SI_4_), .ZN(n6708) );
  XNOR2_X1 U8140 ( .A(n6816), .B(P1_ADDR_REG_1__SCAN_IN), .ZN(n8934) );
  INV_X1 U8141 ( .A(P3_ADDR_REG_1__SCAN_IN), .ZN(n6816) );
  AND2_X1 U8142 ( .A1(n7092), .A2(n7091), .ZN(n8903) );
  NAND2_X1 U8143 ( .A1(n8902), .A2(P3_ADDR_REG_2__SCAN_IN), .ZN(n7091) );
  INV_X1 U8144 ( .A(n8932), .ZN(n7093) );
  AND2_X1 U8145 ( .A1(n7079), .A2(n6593), .ZN(n8905) );
  XNOR2_X1 U8146 ( .A(n8905), .B(n15078), .ZN(n8946) );
  AND2_X1 U8147 ( .A1(n7097), .A2(n7096), .ZN(n8908) );
  NAND2_X1 U8148 ( .A1(n9607), .A2(P3_ADDR_REG_6__SCAN_IN), .ZN(n7096) );
  OR2_X1 U8149 ( .A1(n8952), .A2(n8951), .ZN(n7097) );
  OAI21_X1 U8150 ( .B1(P3_ADDR_REG_16__SCAN_IN), .B2(n14628), .A(n8920), .ZN(
        n8921) );
  INV_X1 U8151 ( .A(P3_REG3_REG_20__SCAN_IN), .ZN(n9134) );
  INV_X1 U8152 ( .A(n9208), .ZN(n7035) );
  OR2_X1 U8153 ( .A1(n7634), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n7654) );
  NOR2_X1 U8154 ( .A1(n7728), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n7740) );
  OR2_X1 U8155 ( .A1(n7711), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n7728) );
  INV_X1 U8156 ( .A(P3_REG3_REG_8__SCAN_IN), .ZN(n10279) );
  NOR2_X1 U8157 ( .A1(n7654), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n7672) );
  INV_X1 U8158 ( .A(P3_REG3_REG_16__SCAN_IN), .ZN(n12401) );
  AND2_X1 U8159 ( .A1(n7672), .A2(n12401), .ZN(n7695) );
  INV_X1 U8160 ( .A(n9203), .ZN(n7037) );
  XNOR2_X1 U8161 ( .A(n12954), .B(n11671), .ZN(n9228) );
  INV_X1 U8162 ( .A(SI_22_), .ZN(n8565) );
  NAND2_X1 U8163 ( .A1(n12349), .A2(n9203), .ZN(n12373) );
  OR2_X1 U8164 ( .A1(n7804), .A2(P3_REG3_REG_25__SCAN_IN), .ZN(n7817) );
  AND4_X1 U8165 ( .A1(n7639), .A2(n7638), .A3(n7637), .A4(n7636), .ZN(n12493)
         );
  NAND2_X1 U8166 ( .A1(n12514), .A2(P3_REG2_REG_2__SCAN_IN), .ZN(n7411) );
  INV_X1 U8167 ( .A(n7184), .ZN(n15044) );
  NAND2_X1 U8168 ( .A1(n15022), .A2(n10079), .ZN(n15042) );
  NAND2_X1 U8169 ( .A1(n10274), .A2(n10275), .ZN(n10276) );
  NAND2_X1 U8170 ( .A1(n15095), .A2(n10701), .ZN(n10702) );
  NAND2_X1 U8171 ( .A1(n10702), .A2(n10703), .ZN(n11024) );
  XNOR2_X1 U8172 ( .A(n11145), .B(n11139), .ZN(n11026) );
  NOR2_X1 U8173 ( .A1(n11032), .A2(n11031), .ZN(n11154) );
  NAND2_X1 U8174 ( .A1(n12769), .A2(n6628), .ZN(n12792) );
  NAND2_X1 U8175 ( .A1(n7182), .A2(n12818), .ZN(n7180) );
  NOR2_X1 U8176 ( .A1(n14348), .A2(n14349), .ZN(n14347) );
  NAND2_X1 U8177 ( .A1(n14345), .A2(n12846), .ZN(n14368) );
  NAND2_X1 U8178 ( .A1(n14368), .A2(n14369), .ZN(n14367) );
  XNOR2_X1 U8179 ( .A(n12849), .B(n14379), .ZN(n14381) );
  NAND2_X1 U8180 ( .A1(n12835), .A2(n6513), .ZN(n7187) );
  NAND2_X1 U8181 ( .A1(n7189), .A2(n12837), .ZN(n7188) );
  NAND2_X1 U8182 ( .A1(n14405), .A2(n6513), .ZN(n7189) );
  NOR2_X1 U8183 ( .A1(n14361), .A2(n7204), .ZN(n7203) );
  INV_X1 U8184 ( .A(n12542), .ZN(n12685) );
  NAND2_X1 U8185 ( .A1(n12911), .A2(n12667), .ZN(n12899) );
  NAND2_X1 U8186 ( .A1(n12929), .A2(n12669), .ZN(n12913) );
  OR2_X1 U8187 ( .A1(n12972), .A2(n12971), .ZN(n12975) );
  OR2_X1 U8188 ( .A1(n13004), .A2(n13018), .ZN(n12985) );
  NAND2_X1 U8189 ( .A1(n6959), .A2(n12638), .ZN(n13007) );
  NAND2_X1 U8190 ( .A1(n13012), .A2(n13013), .ZN(n6959) );
  INV_X1 U8191 ( .A(n13015), .ZN(n13013) );
  AND4_X1 U8192 ( .A1(n7677), .A2(n7676), .A3(n7675), .A4(n7674), .ZN(n13017)
         );
  AND2_X1 U8193 ( .A1(n13024), .A2(n12625), .ZN(n13038) );
  INV_X1 U8194 ( .A(n12617), .ZN(n6980) );
  OR2_X1 U8195 ( .A1(n7575), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n7588) );
  OR2_X1 U8196 ( .A1(n7557), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n7575) );
  INV_X1 U8197 ( .A(SI_11_), .ZN(n8279) );
  INV_X1 U8198 ( .A(n12606), .ZN(n7587) );
  AOI21_X1 U8199 ( .B1(n6969), .B2(n6971), .A(n6968), .ZN(n6967) );
  INV_X1 U8200 ( .A(n12598), .ZN(n6968) );
  NAND2_X1 U8201 ( .A1(n11076), .A2(n6969), .ZN(n6844) );
  INV_X1 U8202 ( .A(n13112), .ZN(n7573) );
  OAI21_X1 U8203 ( .B1(n10892), .B2(n7333), .A(n7331), .ZN(n11065) );
  INV_X1 U8204 ( .A(n7334), .ZN(n7333) );
  AND2_X1 U8205 ( .A1(n7332), .A2(n7877), .ZN(n7331) );
  INV_X1 U8206 ( .A(n12573), .ZN(n6839) );
  NAND2_X1 U8207 ( .A1(n7871), .A2(n7870), .ZN(n10683) );
  NAND2_X1 U8208 ( .A1(n12563), .A2(n12562), .ZN(n10727) );
  NAND2_X1 U8209 ( .A1(n7815), .A2(n7814), .ZN(n12480) );
  OR2_X1 U8210 ( .A1(n6481), .A2(n11202), .ZN(n7814) );
  NAND2_X1 U8211 ( .A1(n7803), .A2(n7802), .ZN(n12382) );
  NAND2_X1 U8212 ( .A1(n7775), .A2(n7774), .ZN(n13134) );
  OR2_X1 U8213 ( .A1(n6480), .A2(n10423), .ZN(n7750) );
  OR2_X1 U8214 ( .A1(n10422), .A2(n7448), .ZN(n6811) );
  INV_X1 U8215 ( .A(n6481), .ZN(n7725) );
  OR2_X1 U8216 ( .A1(n15120), .A2(n15161), .ZN(n15167) );
  INV_X1 U8217 ( .A(P3_IR_REG_23__SCAN_IN), .ZN(n7948) );
  OAI21_X1 U8218 ( .B1(n8865), .B2(n8864), .A(n8867), .ZN(n11644) );
  NAND2_X1 U8219 ( .A1(n7066), .A2(n7812), .ZN(n7824) );
  NAND2_X1 U8220 ( .A1(n7811), .A2(n7810), .ZN(n7066) );
  XNOR2_X1 U8221 ( .A(n7928), .B(P3_IR_REG_26__SCAN_IN), .ZN(n7951) );
  AOI21_X1 U8222 ( .B1(n7062), .B2(n7064), .A(n6642), .ZN(n7061) );
  INV_X1 U8223 ( .A(n7747), .ZN(n7062) );
  INV_X1 U8224 ( .A(n7064), .ZN(n7063) );
  INV_X1 U8225 ( .A(P3_IR_REG_18__SCAN_IN), .ZN(n7723) );
  INV_X1 U8226 ( .A(n7045), .ZN(n7044) );
  OAI21_X1 U8227 ( .B1(n7627), .B2(n7046), .A(n7644), .ZN(n7045) );
  INV_X1 U8228 ( .A(n7642), .ZN(n7046) );
  AND2_X1 U8229 ( .A1(n7661), .A2(n7645), .ZN(n7646) );
  OR2_X1 U8230 ( .A1(n7616), .A2(P3_IR_REG_13__SCAN_IN), .ZN(n7649) );
  OAI21_X1 U8231 ( .B1(n6809), .B2(n10982), .A(n7627), .ZN(n7611) );
  AOI21_X1 U8232 ( .B1(n7050), .B2(n7052), .A(n7049), .ZN(n7048) );
  INV_X1 U8233 ( .A(n7596), .ZN(n7049) );
  AND2_X1 U8234 ( .A1(n7609), .A2(n7597), .ZN(n7598) );
  XNOR2_X1 U8235 ( .A(n7570), .B(P3_IR_REG_10__SCAN_IN), .ZN(n11025) );
  AND2_X1 U8236 ( .A1(n7563), .A2(n7551), .ZN(n7552) );
  NAND2_X1 U8237 ( .A1(n7533), .A2(n7532), .ZN(n7536) );
  OR2_X1 U8238 ( .A1(n7517), .A2(n7516), .ZN(n7533) );
  AOI21_X1 U8239 ( .B1(n6802), .B2(n6804), .A(n6800), .ZN(n6799) );
  INV_X1 U8240 ( .A(n7497), .ZN(n6800) );
  INV_X1 U8241 ( .A(P3_IR_REG_2__SCAN_IN), .ZN(n6878) );
  NAND2_X1 U8242 ( .A1(n8004), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n7432) );
  INV_X1 U8243 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n8215) );
  NAND2_X2 U8244 ( .A1(n13654), .A2(n8023), .ZN(n10036) );
  OR2_X1 U8245 ( .A1(n8518), .A2(n8517), .ZN(n8551) );
  AND2_X1 U8246 ( .A1(n12097), .A2(n12095), .ZN(n13299) );
  INV_X1 U8247 ( .A(n13379), .ZN(n13304) );
  NAND2_X1 U8248 ( .A1(n13261), .A2(n12085), .ZN(n13298) );
  OR2_X1 U8249 ( .A1(n8618), .A2(n13340), .ZN(n8643) );
  NAND2_X1 U8250 ( .A1(n13289), .A2(n12077), .ZN(n13346) );
  OR2_X1 U8251 ( .A1(n8468), .A2(n13364), .ZN(n8491) );
  OR2_X1 U8252 ( .A1(n13334), .A2(n12083), .ZN(n13327) );
  OR2_X1 U8253 ( .A1(n11267), .A2(n6940), .ZN(n6939) );
  OR2_X1 U8254 ( .A1(n14938), .A2(n13490), .ZN(n6940) );
  AOI21_X1 U8255 ( .B1(n14863), .B2(P2_REG1_REG_10__SCAN_IN), .A(n14859), .ZN(
        n9741) );
  AOI21_X1 U8256 ( .B1(P2_REG1_REG_17__SCAN_IN), .B2(n13468), .A(n14909), .ZN(
        n13475) );
  NAND2_X1 U8257 ( .A1(n8725), .A2(n8724), .ZN(n13498) );
  NAND2_X1 U8258 ( .A1(n13506), .A2(n13505), .ZN(n13504) );
  INV_X1 U8259 ( .A(n7149), .ZN(n7148) );
  NAND2_X1 U8260 ( .A1(n13546), .A2(n6565), .ZN(n6756) );
  OAI21_X1 U8261 ( .B1(n13522), .B2(n7150), .A(n6504), .ZN(n7149) );
  NAND2_X1 U8262 ( .A1(n6956), .A2(n6955), .ZN(n13556) );
  INV_X1 U8263 ( .A(n13554), .ZN(n6956) );
  NOR2_X2 U8264 ( .A1(n13556), .A2(n13719), .ZN(n13534) );
  OR2_X1 U8265 ( .A1(n13590), .A2(n13380), .ZN(n7358) );
  INV_X1 U8266 ( .A(n8570), .ZN(n8569) );
  NAND2_X1 U8267 ( .A1(n13617), .A2(n13622), .ZN(n12139) );
  NAND2_X1 U8268 ( .A1(n6725), .A2(n6724), .ZN(n13595) );
  AND2_X1 U8269 ( .A1(n7159), .A2(n7162), .ZN(n6724) );
  NAND2_X1 U8270 ( .A1(n13747), .A2(n13597), .ZN(n7162) );
  OAI21_X1 U8271 ( .B1(n13683), .B2(n6759), .A(n7142), .ZN(n13617) );
  NAND2_X1 U8272 ( .A1(n12132), .A2(n7145), .ZN(n6759) );
  INV_X1 U8273 ( .A(n7143), .ZN(n7142) );
  INV_X1 U8274 ( .A(n7144), .ZN(n7145) );
  AOI21_X1 U8275 ( .B1(n13650), .B2(n13636), .A(n13637), .ZN(n13635) );
  AND2_X1 U8276 ( .A1(n6721), .A2(n6527), .ZN(n13651) );
  INV_X1 U8277 ( .A(n6954), .ZN(n13674) );
  AOI21_X1 U8278 ( .B1(n7123), .B2(n11361), .A(n6496), .ZN(n6758) );
  AOI22_X1 U8279 ( .A1(n11307), .A2(n11306), .B1(n13328), .B2(n13772), .ZN(
        n11308) );
  NAND2_X1 U8280 ( .A1(n11359), .A2(n11290), .ZN(n11307) );
  NAND2_X1 U8281 ( .A1(n7166), .A2(n7164), .ZN(n6720) );
  INV_X1 U8282 ( .A(n7165), .ZN(n7164) );
  NAND2_X1 U8283 ( .A1(n11130), .A2(n7176), .ZN(n11277) );
  NAND2_X1 U8284 ( .A1(n8289), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n8313) );
  INV_X1 U8285 ( .A(n8291), .ZN(n8289) );
  INV_X1 U8286 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n8312) );
  INV_X1 U8287 ( .A(n11730), .ZN(n11124) );
  OR2_X1 U8288 ( .A1(n8216), .A2(n8215), .ZN(n8240) );
  NAND2_X1 U8289 ( .A1(n6750), .A2(n6752), .ZN(n6748) );
  NAND2_X1 U8290 ( .A1(n7130), .A2(n6750), .ZN(n6749) );
  NOR2_X2 U8291 ( .A1(n10381), .A2(n10380), .ZN(n10382) );
  NAND2_X1 U8292 ( .A1(n10183), .A2(n10184), .ZN(n10374) );
  NAND2_X1 U8293 ( .A1(n9915), .A2(n10001), .ZN(n10002) );
  NAND2_X1 U8295 ( .A1(n8257), .A2(n8256), .ZN(n14987) );
  OAI22_X1 U8296 ( .A1(n8762), .A2(n9450), .B1(n8056), .B2(n8059), .ZN(n8060)
         );
  CLKBUF_X1 U8297 ( .A(n9920), .Z(n14937) );
  AND2_X1 U8298 ( .A1(n9815), .A2(n10141), .ZN(n14994) );
  INV_X1 U8299 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n8808) );
  NAND2_X1 U8300 ( .A1(n7008), .A2(n7007), .ZN(n8803) );
  NOR3_X1 U8301 ( .A1(P2_IR_REG_20__SCAN_IN), .A2(P2_IR_REG_21__SCAN_IN), .A3(
        n8010), .ZN(n7007) );
  OR2_X1 U8302 ( .A1(P2_IR_REG_18__SCAN_IN), .A2(P2_IR_REG_19__SCAN_IN), .ZN(
        n8010) );
  OR2_X1 U8303 ( .A1(n8411), .A2(P2_IR_REG_14__SCAN_IN), .ZN(n8391) );
  INV_X1 U8304 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n8156) );
  NAND2_X1 U8305 ( .A1(n10741), .A2(n6789), .ZN(n6788) );
  INV_X1 U8306 ( .A(n10742), .ZN(n6789) );
  NOR2_X1 U8307 ( .A1(n10963), .A2(n10962), .ZN(n10989) );
  INV_X1 U8308 ( .A(n10822), .ZN(n7113) );
  NOR2_X1 U8309 ( .A1(n9369), .A2(n9354), .ZN(n13858) );
  AND2_X1 U8310 ( .A1(n9353), .A2(n9352), .ZN(n9354) );
  OR2_X1 U8311 ( .A1(n11345), .A2(n11344), .ZN(n6781) );
  NOR2_X1 U8312 ( .A1(n11352), .A2(n6779), .ZN(n6778) );
  INV_X1 U8313 ( .A(n6781), .ZN(n6779) );
  INV_X1 U8314 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n10946) );
  OR2_X1 U8315 ( .A1(n10947), .A2(n10946), .ZN(n10963) );
  NAND2_X1 U8316 ( .A1(n7106), .A2(n7107), .ZN(n13870) );
  AND2_X1 U8317 ( .A1(n12268), .A2(n7108), .ZN(n7107) );
  AND2_X1 U8318 ( .A1(n12284), .A2(n12282), .ZN(n13871) );
  OR2_X1 U8319 ( .A1(n10997), .A2(n11419), .ZN(n11173) );
  NOR2_X1 U8320 ( .A1(n11173), .A2(n11172), .ZN(n11188) );
  AND2_X1 U8321 ( .A1(n13873), .A2(n12267), .ZN(n13890) );
  NAND2_X1 U8322 ( .A1(n13834), .A2(n12247), .ZN(n13838) );
  INV_X1 U8323 ( .A(n11556), .ZN(n11555) );
  AND2_X1 U8324 ( .A1(n11536), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n11546) );
  INV_X1 U8325 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n10475) );
  OR2_X1 U8326 ( .A1(n10476), .A2(n10475), .ZN(n10572) );
  OR2_X1 U8327 ( .A1(n10465), .A2(n10827), .ZN(n10476) );
  AND2_X1 U8328 ( .A1(n9368), .A2(n9367), .ZN(n9676) );
  AOI22_X1 U8329 ( .A1(n10746), .A2(n14725), .B1(n14299), .B2(n9366), .ZN(
        n9367) );
  NAND2_X1 U8330 ( .A1(n13996), .A2(n12301), .ZN(n9368) );
  NAND2_X1 U8331 ( .A1(n9676), .A2(n9675), .ZN(n9674) );
  NAND2_X1 U8332 ( .A1(n6524), .A2(n12244), .ZN(n13834) );
  AND2_X1 U8333 ( .A1(n13835), .A2(n12243), .ZN(n13912) );
  NOR2_X1 U8334 ( .A1(n10572), .A2(n10571), .ZN(n10582) );
  OR2_X1 U8335 ( .A1(n13930), .A2(n13931), .ZN(n13847) );
  AND2_X1 U8336 ( .A1(n12206), .A2(n12200), .ZN(n7119) );
  NOR2_X1 U8337 ( .A1(n6764), .A2(n6765), .ZN(n6762) );
  INV_X1 U8338 ( .A(n10647), .ZN(n6765) );
  AND2_X1 U8339 ( .A1(n11251), .A2(n11250), .ZN(n13851) );
  OR2_X1 U8340 ( .A1(n9585), .A2(n9584), .ZN(n6865) );
  NAND2_X1 U8341 ( .A1(n6865), .A2(n6864), .ZN(n6863) );
  NAND2_X1 U8342 ( .A1(n9601), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n6864) );
  AND2_X1 U8343 ( .A1(n7076), .A2(n7075), .ZN(n9622) );
  NAND2_X1 U8344 ( .A1(n9885), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n7075) );
  NOR2_X1 U8345 ( .A1(n9622), .A2(n9621), .ZN(n9620) );
  NAND2_X1 U8346 ( .A1(n14608), .A2(n14607), .ZN(n14606) );
  XNOR2_X1 U8347 ( .A(n14035), .B(n11164), .ZN(n11417) );
  NAND2_X1 U8348 ( .A1(n14042), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n6858) );
  NOR2_X1 U8349 ( .A1(n14652), .A2(n14032), .ZN(n14033) );
  NAND2_X1 U8350 ( .A1(n11693), .A2(n11692), .ZN(n11691) );
  NAND2_X1 U8351 ( .A1(n6735), .A2(n6738), .ZN(n11686) );
  NAND2_X1 U8352 ( .A1(n6741), .A2(n6520), .ZN(n6735) );
  INV_X1 U8353 ( .A(n7263), .ZN(n7266) );
  NAND2_X1 U8354 ( .A1(n14106), .A2(n11609), .ZN(n14083) );
  INV_X1 U8355 ( .A(n7248), .ZN(n7247) );
  NAND2_X1 U8356 ( .A1(n11608), .A2(n14102), .ZN(n14106) );
  NAND2_X1 U8357 ( .A1(n11513), .A2(n11512), .ZN(n14157) );
  NAND2_X1 U8358 ( .A1(n11468), .A2(n11900), .ZN(n11473) );
  NAND2_X1 U8359 ( .A1(n11434), .A2(n6518), .ZN(n11468) );
  AND2_X1 U8360 ( .A1(n11245), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n11378) );
  AND2_X1 U8361 ( .A1(n11188), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n11245) );
  AND2_X1 U8362 ( .A1(n11242), .A2(n11241), .ZN(n12203) );
  NAND2_X1 U8363 ( .A1(n11007), .A2(n6912), .ZN(n11187) );
  NAND2_X1 U8364 ( .A1(n11007), .A2(n11006), .ZN(n11050) );
  AOI21_X1 U8365 ( .B1(n7285), .B2(n7287), .A(n6568), .ZN(n7283) );
  AOI21_X1 U8366 ( .B1(n14664), .B2(n7259), .A(n6579), .ZN(n7257) );
  INV_X1 U8367 ( .A(n7259), .ZN(n7258) );
  INV_X1 U8368 ( .A(n7274), .ZN(n7273) );
  NOR2_X1 U8369 ( .A1(n14711), .A2(n13945), .ZN(n14694) );
  NAND2_X1 U8370 ( .A1(n14694), .A2(n14754), .ZN(n14693) );
  OR2_X1 U8371 ( .A1(n10471), .A2(n12035), .ZN(n11636) );
  NAND2_X1 U8372 ( .A1(n7269), .A2(n9889), .ZN(n10425) );
  NOR2_X1 U8373 ( .A1(n7233), .A2(n9751), .ZN(n7232) );
  NAND2_X1 U8374 ( .A1(n9756), .A2(n11999), .ZN(n7269) );
  NAND2_X1 U8375 ( .A1(n9656), .A2(n6906), .ZN(n10396) );
  INV_X1 U8376 ( .A(n14167), .ZN(n14455) );
  AND2_X1 U8377 ( .A1(n7293), .A2(n11593), .ZN(n6893) );
  NAND2_X1 U8378 ( .A1(n6894), .A2(n7293), .ZN(n11695) );
  NAND2_X1 U8379 ( .A1(n11603), .A2(n11602), .ZN(n14166) );
  NAND2_X1 U8380 ( .A1(n14684), .A2(n10497), .ZN(n10498) );
  NOR2_X1 U8381 ( .A1(n14297), .A2(n11965), .ZN(n14724) );
  INV_X1 U8382 ( .A(n14701), .ZN(n14780) );
  NAND2_X1 U8383 ( .A1(n6917), .A2(n6918), .ZN(n8716) );
  XNOR2_X1 U8384 ( .A(n8760), .B(n8759), .ZN(n11655) );
  XNOR2_X1 U8385 ( .A(n8705), .B(n8687), .ZN(n11664) );
  NAND2_X1 U8386 ( .A1(n8591), .A2(n8590), .ZN(n8594) );
  XNOR2_X1 U8387 ( .A(n9323), .B(P1_IR_REG_20__SCAN_IN), .ZN(n11978) );
  XNOR2_X1 U8388 ( .A(n8514), .B(n8538), .ZN(n11469) );
  AND2_X1 U8389 ( .A1(n9636), .A2(n9877), .ZN(n11416) );
  XNOR2_X1 U8390 ( .A(n6726), .B(n8326), .ZN(n10943) );
  OAI21_X1 U8391 ( .B1(n8325), .B2(n8327), .A(n8328), .ZN(n6726) );
  OR2_X1 U8392 ( .A1(n9476), .A2(P1_IR_REG_6__SCAN_IN), .ZN(n9513) );
  XNOR2_X1 U8393 ( .A(n8136), .B(n6707), .ZN(n9884) );
  INV_X1 U8394 ( .A(n8135), .ZN(n6707) );
  INV_X1 U8395 ( .A(P3_ADDR_REG_0__SCAN_IN), .ZN(n9959) );
  XNOR2_X1 U8396 ( .A(n8903), .B(n7090), .ZN(n8942) );
  NAND2_X1 U8397 ( .A1(n8944), .A2(n8945), .ZN(n8948) );
  XNOR2_X1 U8398 ( .A(n8946), .B(P1_ADDR_REG_5__SCAN_IN), .ZN(n8947) );
  NAND2_X1 U8399 ( .A1(n8953), .A2(n8954), .ZN(n8956) );
  XNOR2_X1 U8400 ( .A(n8908), .B(n7095), .ZN(n8955) );
  AND2_X1 U8401 ( .A1(n7101), .A2(n7100), .ZN(n8965) );
  NAND2_X1 U8402 ( .A1(n9975), .A2(P3_ADDR_REG_8__SCAN_IN), .ZN(n7100) );
  NOR2_X1 U8403 ( .A1(n8913), .A2(n8912), .ZN(n8973) );
  XOR2_X1 U8404 ( .A(n14646), .B(n8921), .Z(n8924) );
  AND2_X1 U8405 ( .A1(n7013), .A2(n7011), .ZN(n7010) );
  INV_X1 U8406 ( .A(n7016), .ZN(n7011) );
  NAND2_X1 U8407 ( .A1(n7013), .A2(n7015), .ZN(n7012) );
  OR2_X1 U8408 ( .A1(n9245), .A2(n9244), .ZN(n7015) );
  NAND2_X1 U8409 ( .A1(n7028), .A2(n7025), .ZN(n12398) );
  INV_X1 U8410 ( .A(n7027), .ZN(n7025) );
  NAND2_X1 U8411 ( .A1(n7030), .A2(n7029), .ZN(n7028) );
  NAND2_X1 U8412 ( .A1(n12492), .A2(n7026), .ZN(n7018) );
  NAND2_X1 U8413 ( .A1(n7790), .A2(n7789), .ZN(n12922) );
  AND4_X1 U8414 ( .A1(n7626), .A2(n7625), .A3(n7624), .A4(n7623), .ZN(n12437)
         );
  NAND2_X1 U8415 ( .A1(n7036), .A2(n9208), .ZN(n12440) );
  NAND2_X1 U8416 ( .A1(n12349), .A2(n6528), .ZN(n7036) );
  AND4_X2 U8417 ( .A1(n7427), .A2(n7426), .A3(n7425), .A4(n7424), .ZN(n15110)
         );
  NAND2_X1 U8418 ( .A1(n7022), .A2(n7021), .ZN(n7020) );
  NAND2_X1 U8419 ( .A1(n7038), .A2(n6557), .ZN(n10811) );
  NAND2_X1 U8420 ( .A1(n7038), .A2(n9187), .ZN(n10810) );
  NAND2_X1 U8421 ( .A1(n10028), .A2(n9248), .ZN(n12500) );
  AND2_X1 U8422 ( .A1(n9247), .A2(n12736), .ZN(n12502) );
  OR2_X1 U8423 ( .A1(n12696), .A2(n7349), .ZN(n12531) );
  NAND2_X1 U8424 ( .A1(n12728), .A2(n12727), .ZN(n12729) );
  NAND4_X1 U8425 ( .A1(n7834), .A2(n7833), .A3(n7832), .A4(n7831), .ZN(n12746)
         );
  OAI211_X1 U8426 ( .C1(n7471), .C2(n13208), .A(n7754), .B(n7753), .ZN(n12752)
         );
  OAI211_X1 U8427 ( .C1(n7471), .C2(n13211), .A(n7743), .B(n7742), .ZN(n12753)
         );
  INV_X1 U8428 ( .A(n12493), .ZN(n13063) );
  INV_X1 U8429 ( .A(n12437), .ZN(n13050) );
  NAND2_X1 U8430 ( .A1(n15066), .A2(n10081), .ZN(n10082) );
  INV_X1 U8431 ( .A(n15064), .ZN(n15090) );
  INV_X1 U8432 ( .A(n7207), .ZN(n10097) );
  OAI22_X1 U8433 ( .A1(n10158), .A2(n10157), .B1(n10156), .B2(n10155), .ZN(
        n10271) );
  NOR2_X1 U8434 ( .A1(n10262), .A2(n10263), .ZN(n10266) );
  NOR2_X1 U8435 ( .A1(n15080), .A2(n15081), .ZN(n15079) );
  OAI21_X1 U8436 ( .B1(n15080), .B2(n7209), .A(n7208), .ZN(n11020) );
  NAND2_X1 U8437 ( .A1(n7210), .A2(P3_REG2_REG_9__SCAN_IN), .ZN(n7209) );
  NAND2_X1 U8438 ( .A1(n10695), .A2(n7210), .ZN(n7208) );
  INV_X1 U8439 ( .A(n10697), .ZN(n7210) );
  XNOR2_X1 U8440 ( .A(n11138), .B(n11139), .ZN(n11022) );
  XNOR2_X1 U8441 ( .A(n12792), .B(n12802), .ZN(n12771) );
  NAND2_X1 U8442 ( .A1(n7193), .A2(n7191), .ZN(n14387) );
  INV_X1 U8443 ( .A(n7195), .ZN(n7191) );
  NAND2_X1 U8444 ( .A1(n7186), .A2(n6882), .ZN(n6881) );
  NAND2_X1 U8445 ( .A1(n14404), .A2(n6650), .ZN(n7186) );
  OR2_X1 U8446 ( .A1(n12854), .A2(n12853), .ZN(n6883) );
  OR2_X1 U8447 ( .A1(n12837), .A2(n14405), .ZN(n7190) );
  AND2_X1 U8448 ( .A1(n6543), .A2(n7328), .ZN(n12935) );
  AND2_X1 U8449 ( .A1(n12971), .A2(n12647), .ZN(n6974) );
  NAND2_X1 U8450 ( .A1(n7732), .A2(n12647), .ZN(n12981) );
  NAND2_X1 U8451 ( .A1(n7739), .A2(n7738), .ZN(n13145) );
  NAND2_X1 U8452 ( .A1(n7342), .A2(n7889), .ZN(n13028) );
  NAND2_X1 U8453 ( .A1(n7343), .A2(n6519), .ZN(n7342) );
  NAND2_X1 U8454 ( .A1(n11074), .A2(n11073), .ZN(n13113) );
  NAND2_X1 U8455 ( .A1(n11075), .A2(n12595), .ZN(n11063) );
  NAND2_X1 U8456 ( .A1(n7336), .A2(n7875), .ZN(n11079) );
  NAND2_X1 U8457 ( .A1(n10519), .A2(n12573), .ZN(n10685) );
  NAND2_X1 U8458 ( .A1(n6973), .A2(n10088), .ZN(n6972) );
  NAND2_X1 U8459 ( .A1(n10028), .A2(n12695), .ZN(n15108) );
  NAND2_X1 U8460 ( .A1(n12524), .A2(n12523), .ZN(n13186) );
  AND2_X1 U8461 ( .A1(n8892), .A2(n6848), .ZN(n6847) );
  AND2_X1 U8462 ( .A1(n8893), .A2(n15177), .ZN(n6848) );
  INV_X1 U8463 ( .A(n12535), .ZN(n12885) );
  INV_X1 U8464 ( .A(n12480), .ZN(n13193) );
  INV_X1 U8465 ( .A(n12545), .ZN(n13210) );
  NAND2_X1 U8466 ( .A1(n7653), .A2(n7652), .ZN(n13231) );
  NAND2_X1 U8467 ( .A1(n9766), .A2(P3_STATE_REG_SCAN_IN), .ZN(n13238) );
  INV_X1 U8468 ( .A(n7391), .ZN(n11647) );
  XNOR2_X1 U8469 ( .A(n11644), .B(n11642), .ZN(n11666) );
  INV_X1 U8470 ( .A(P3_IR_REG_28__SCAN_IN), .ZN(n7393) );
  NAND2_X1 U8471 ( .A1(n7923), .A2(n6514), .ZN(n10912) );
  MUX2_X1 U8472 ( .A(P3_IR_REG_31__SCAN_IN), .B(n7922), .S(
        P3_IR_REG_24__SCAN_IN), .Z(n7923) );
  NAND2_X1 U8473 ( .A1(n7345), .A2(n7687), .ZN(n7921) );
  INV_X1 U8474 ( .A(SI_24_), .ZN(n10910) );
  NAND2_X1 U8475 ( .A1(n7759), .A2(n7758), .ZN(n7773) );
  OR2_X1 U8476 ( .A1(n7853), .A2(n13241), .ZN(n7855) );
  INV_X1 U8477 ( .A(SI_19_), .ZN(n9992) );
  NAND2_X1 U8478 ( .A1(n7721), .A2(n7720), .ZN(n7734) );
  NAND2_X1 U8479 ( .A1(n7718), .A2(n7717), .ZN(n7721) );
  INV_X1 U8480 ( .A(SI_18_), .ZN(n9883) );
  NAND2_X1 U8481 ( .A1(n6794), .A2(n7053), .ZN(n7706) );
  NAND2_X1 U8482 ( .A1(n7665), .A2(n7055), .ZN(n6794) );
  NAND2_X1 U8483 ( .A1(n7685), .A2(n7684), .ZN(n7702) );
  INV_X1 U8484 ( .A(SI_15_), .ZN(n9639) );
  NAND2_X1 U8485 ( .A1(n7628), .A2(n7627), .ZN(n7643) );
  INV_X1 U8486 ( .A(SI_12_), .ZN(n9489) );
  XNOR2_X1 U8487 ( .A(n7605), .B(n7613), .ZN(n12773) );
  NAND2_X1 U8488 ( .A1(n7582), .A2(n7581), .ZN(n7595) );
  INV_X1 U8489 ( .A(n11025), .ZN(n11021) );
  NAND2_X1 U8490 ( .A1(n6801), .A2(n7483), .ZN(n7496) );
  NAND2_X1 U8491 ( .A1(n7482), .A2(n7481), .ZN(n6801) );
  NOR2_X1 U8492 ( .A1(n9434), .A2(P3_STATE_REG_SCAN_IN), .ZN(n14317) );
  NAND2_X1 U8493 ( .A1(n6687), .A2(n6685), .ZN(n7430) );
  NAND2_X1 U8494 ( .A1(n12158), .A2(n7357), .ZN(n13253) );
  NOR2_X1 U8495 ( .A1(n13252), .A2(n6987), .ZN(n6986) );
  INV_X1 U8496 ( .A(n7357), .ZN(n6987) );
  NAND2_X1 U8497 ( .A1(n7002), .A2(n7001), .ZN(n7000) );
  INV_X1 U8498 ( .A(n7003), .ZN(n7001) );
  NAND2_X1 U8499 ( .A1(n12066), .A2(n7006), .ZN(n13289) );
  AND2_X1 U8500 ( .A1(n13290), .A2(n12065), .ZN(n7006) );
  INV_X1 U8501 ( .A(n12081), .ZN(n13291) );
  NAND2_X1 U8502 ( .A1(n11092), .A2(n11725), .ZN(n11732) );
  AND2_X1 U8503 ( .A1(n10044), .A2(n10042), .ZN(n10043) );
  AND2_X1 U8504 ( .A1(n6998), .A2(n6997), .ZN(n6996) );
  INV_X1 U8505 ( .A(n10556), .ZN(n6997) );
  OR2_X1 U8506 ( .A1(n10556), .A2(n10551), .ZN(n6995) );
  NAND2_X1 U8507 ( .A1(n11762), .A2(n6998), .ZN(n11774) );
  NAND2_X1 U8508 ( .A1(n11732), .A2(n7005), .ZN(n11095) );
  AND2_X1 U8509 ( .A1(n13360), .A2(n6989), .ZN(n6988) );
  AND2_X1 U8510 ( .A1(n6990), .A2(n6989), .ZN(n13361) );
  OR2_X1 U8511 ( .A1(n13366), .A2(n13657), .ZN(n13351) );
  OR2_X1 U8512 ( .A1(n13366), .A2(n13655), .ZN(n13353) );
  NAND2_X1 U8513 ( .A1(n10049), .A2(P2_STATE_REG_SCAN_IN), .ZN(n13352) );
  NAND2_X1 U8514 ( .A1(n9823), .A2(n9816), .ZN(n13334) );
  INV_X1 U8515 ( .A(n13334), .ZN(n13359) );
  NOR2_X1 U8516 ( .A1(n8858), .A2(n6939), .ZN(n7367) );
  NOR2_X1 U8517 ( .A1(n8856), .A2(n11267), .ZN(n6670) );
  NAND2_X1 U8518 ( .A1(n8700), .A2(n8699), .ZN(n13376) );
  NAND2_X1 U8519 ( .A1(n8679), .A2(n8678), .ZN(n13377) );
  NAND4_X1 U8520 ( .A1(n8079), .A2(n8078), .A3(n8077), .A4(n8076), .ZN(n13395)
         );
  NAND2_X1 U8521 ( .A1(n8694), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n8052) );
  NOR2_X1 U8522 ( .A1(n14839), .A2(n14838), .ZN(n14841) );
  AOI21_X1 U8523 ( .B1(n14875), .B2(P2_REG1_REG_13__SCAN_IN), .A(n14870), .ZN(
        n14886) );
  NOR2_X1 U8524 ( .A1(n10928), .A2(n14894), .ZN(n10930) );
  OR2_X1 U8525 ( .A1(n9644), .A2(n11657), .ZN(n14884) );
  INV_X1 U8526 ( .A(n13711), .ZN(n13526) );
  NAND2_X1 U8527 ( .A1(n13546), .A2(n7151), .ZN(n13539) );
  OAI21_X1 U8528 ( .B1(n13650), .B2(n13637), .A(n7160), .ZN(n7163) );
  OAI211_X1 U8529 ( .C1(n7141), .C2(n12133), .A(n7140), .B(n12135), .ZN(n13630) );
  INV_X1 U8530 ( .A(n7146), .ZN(n7141) );
  NAND2_X1 U8531 ( .A1(n13684), .A2(n7146), .ZN(n7140) );
  NAND2_X1 U8532 ( .A1(n13681), .A2(n12134), .ZN(n13653) );
  NAND2_X1 U8533 ( .A1(n7126), .A2(n7127), .ZN(n11302) );
  NAND2_X1 U8534 ( .A1(n7126), .A2(n7123), .ZN(n13775) );
  NAND2_X1 U8535 ( .A1(n7363), .A2(n11298), .ZN(n11358) );
  NAND2_X1 U8536 ( .A1(n7167), .A2(n7169), .ZN(n11280) );
  NAND2_X1 U8537 ( .A1(n7174), .A2(n7171), .ZN(n7167) );
  NAND2_X1 U8538 ( .A1(n7138), .A2(n11122), .ZN(n11275) );
  NAND2_X1 U8539 ( .A1(n7139), .A2(n6521), .ZN(n7138) );
  INV_X1 U8540 ( .A(n11121), .ZN(n7139) );
  NAND2_X1 U8541 ( .A1(n7172), .A2(n7177), .ZN(n11127) );
  INV_X1 U8542 ( .A(n7178), .ZN(n7177) );
  NAND2_X1 U8543 ( .A1(n8237), .A2(n8236), .ZN(n10779) );
  OAI21_X1 U8544 ( .B1(n7130), .B2(n6752), .A(n6750), .ZN(n11501) );
  NAND2_X1 U8545 ( .A1(n10619), .A2(n10618), .ZN(n11499) );
  NAND2_X1 U8546 ( .A1(n10368), .A2(n10320), .ZN(n10321) );
  NAND2_X1 U8547 ( .A1(n13606), .A2(n10142), .ZN(n13688) );
  NAND2_X1 U8548 ( .A1(n14932), .A2(n9912), .ZN(n13607) );
  OR2_X1 U8549 ( .A1(n10138), .A2(n12163), .ZN(n11660) );
  INV_X1 U8550 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n8008) );
  NAND2_X1 U8551 ( .A1(n8056), .A2(n13824), .ZN(n8007) );
  INV_X1 U8552 ( .A(n13688), .ZN(n13553) );
  INV_X1 U8553 ( .A(n11660), .ZN(n13669) );
  NAND2_X1 U8554 ( .A1(n6949), .A2(n6947), .ZN(n13789) );
  NOR2_X1 U8555 ( .A1(n6541), .A2(n6948), .ZN(n6947) );
  INV_X1 U8556 ( .A(n13697), .ZN(n6948) );
  NAND2_X1 U8557 ( .A1(n6679), .A2(n15000), .ZN(n6678) );
  INV_X1 U8558 ( .A(n13703), .ZN(n6679) );
  INV_X1 U8559 ( .A(n13710), .ZN(n13718) );
  OAI21_X1 U8560 ( .B1(n13715), .B2(n14984), .A(n13714), .ZN(n13716) );
  NAND2_X1 U8561 ( .A1(n9799), .A2(n9798), .ZN(n14931) );
  AND2_X1 U8562 ( .A1(n10046), .A2(P2_STATE_REG_SCAN_IN), .ZN(n14932) );
  INV_X1 U8563 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n7986) );
  NAND2_X1 U8564 ( .A1(n13809), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7987) );
  INV_X1 U8565 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n7989) );
  INV_X1 U8566 ( .A(n8811), .ZN(n8812) );
  XNOR2_X1 U8567 ( .A(n8819), .B(n8818), .ZN(n13818) );
  INV_X1 U8568 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n8818) );
  INV_X1 U8569 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n11651) );
  INV_X1 U8570 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n10212) );
  INV_X1 U8571 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n10134) );
  INV_X1 U8572 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n9876) );
  INV_X1 U8573 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n9616) );
  INV_X1 U8574 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n9568) );
  INV_X1 U8575 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n9559) );
  INV_X1 U8576 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n9518) );
  INV_X1 U8577 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n9512) );
  INV_X1 U8578 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n9482) );
  AND2_X1 U8579 ( .A1(n8188), .A2(n8234), .ZN(n13444) );
  INV_X1 U8580 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n9451) );
  INV_X1 U8581 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n9448) );
  INV_X1 U8582 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n9452) );
  INV_X1 U8583 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n9446) );
  NAND2_X1 U8584 ( .A1(n10748), .A2(n10747), .ZN(n10823) );
  NAND2_X1 U8585 ( .A1(n13940), .A2(n6788), .ZN(n10748) );
  AND2_X1 U8586 ( .A1(n11580), .A2(n11596), .ZN(n13828) );
  NAND2_X1 U8587 ( .A1(n13825), .A2(n6768), .ZN(n13827) );
  OAI21_X1 U8588 ( .B1(n13952), .B2(n12292), .A(n7104), .ZN(n13825) );
  NAND2_X1 U8589 ( .A1(n13951), .A2(n6501), .ZN(n6768) );
  NAND2_X1 U8590 ( .A1(n12176), .A2(n12175), .ZN(n14441) );
  INV_X1 U8591 ( .A(n6772), .ZN(n6771) );
  NAND2_X1 U8592 ( .A1(n13921), .A2(n9386), .ZN(n9409) );
  AOI21_X1 U8593 ( .B1(n7104), .B2(n12292), .A(n12300), .ZN(n7103) );
  AND2_X1 U8594 ( .A1(n10823), .A2(n7112), .ZN(n11108) );
  NAND2_X1 U8595 ( .A1(n10823), .A2(n10822), .ZN(n10824) );
  AND2_X1 U8596 ( .A1(n11477), .A2(n11523), .ZN(n14160) );
  NAND2_X1 U8597 ( .A1(n6780), .A2(n6778), .ZN(n11458) );
  NAND2_X1 U8598 ( .A1(n14448), .A2(n7348), .ZN(n14449) );
  AND2_X1 U8599 ( .A1(n14449), .A2(n12200), .ZN(n13883) );
  INV_X1 U8600 ( .A(n12203), .ZN(n14489) );
  XNOR2_X1 U8601 ( .A(n10644), .B(n10645), .ZN(n10648) );
  NAND2_X1 U8602 ( .A1(n11458), .A2(n11457), .ZN(n11461) );
  AND2_X1 U8603 ( .A1(n11525), .A2(n11524), .ZN(n14148) );
  AOI21_X1 U8604 ( .B1(n11339), .B2(n11338), .A(n7355), .ZN(n14462) );
  NAND2_X1 U8605 ( .A1(n7115), .A2(n12207), .ZN(n13930) );
  NAND2_X1 U8606 ( .A1(n14449), .A2(n7119), .ZN(n7115) );
  NAND2_X1 U8607 ( .A1(n9407), .A2(n9406), .ZN(n13938) );
  AND2_X1 U8608 ( .A1(n13946), .A2(n14777), .ZN(n14463) );
  AND4_X1 U8609 ( .A1(n10994), .A2(n10993), .A3(n10992), .A4(n10991), .ZN(
        n13965) );
  XNOR2_X1 U8610 ( .A(n12189), .B(n12190), .ZN(n13962) );
  NAND2_X1 U8611 ( .A1(n13962), .A2(n13961), .ZN(n14448) );
  INV_X1 U8612 ( .A(n13938), .ZN(n14465) );
  AND2_X1 U8613 ( .A1(n11987), .A2(n6596), .ZN(n12053) );
  OR2_X1 U8614 ( .A1(n9412), .A2(n9306), .ZN(n13979) );
  INV_X1 U8615 ( .A(n11775), .ZN(n13996) );
  NOR2_X1 U8616 ( .A1(n9593), .A2(n6537), .ZN(n9855) );
  INV_X1 U8617 ( .A(n7076), .ZN(n9853) );
  INV_X1 U8618 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n9607) );
  NOR2_X1 U8619 ( .A1(n9689), .A2(n9688), .ZN(n9969) );
  NOR2_X1 U8620 ( .A1(n9686), .A2(n6867), .ZN(n9689) );
  NOR2_X1 U8621 ( .A1(n6869), .A2(n6868), .ZN(n6867) );
  NOR2_X1 U8622 ( .A1(n9969), .A2(n6866), .ZN(n9972) );
  AND2_X1 U8623 ( .A1(n10449), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n6866) );
  NAND2_X1 U8624 ( .A1(n9972), .A2(n9971), .ZN(n10219) );
  INV_X1 U8625 ( .A(n7072), .ZN(n10225) );
  INV_X1 U8626 ( .A(n7070), .ZN(n10528) );
  NOR2_X1 U8627 ( .A1(n11410), .A2(n6857), .ZN(n14565) );
  AND2_X1 U8628 ( .A1(n11411), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n6857) );
  NAND2_X1 U8629 ( .A1(n14565), .A2(n14564), .ZN(n14563) );
  NOR2_X1 U8630 ( .A1(n14566), .A2(n6623), .ZN(n14579) );
  NAND2_X1 U8631 ( .A1(n14579), .A2(n14580), .ZN(n14578) );
  NAND2_X1 U8632 ( .A1(n14563), .A2(n6855), .ZN(n14577) );
  NAND2_X1 U8633 ( .A1(n6856), .A2(n11412), .ZN(n6855) );
  NAND2_X1 U8634 ( .A1(n14577), .A2(n14576), .ZN(n14575) );
  NAND2_X1 U8635 ( .A1(n11407), .A2(n11406), .ZN(n14028) );
  INV_X1 U8636 ( .A(n6861), .ZN(n14617) );
  INV_X1 U8637 ( .A(n14638), .ZN(n14651) );
  INV_X1 U8638 ( .A(n6859), .ZN(n14629) );
  INV_X1 U8639 ( .A(n14642), .ZN(n14658) );
  INV_X1 U8640 ( .A(n12045), .ZN(n14197) );
  AOI21_X1 U8641 ( .B1(n11961), .B2(n11960), .A(n11959), .ZN(n14201) );
  AOI21_X1 U8642 ( .B1(n11661), .B2(n11960), .A(n11595), .ZN(n14204) );
  XNOR2_X1 U8643 ( .A(n7231), .B(n6889), .ZN(n14207) );
  NAND2_X1 U8644 ( .A1(n6732), .A2(n11612), .ZN(n6731) );
  NAND2_X1 U8645 ( .A1(n14076), .A2(n7294), .ZN(n11629) );
  NAND2_X1 U8646 ( .A1(n11630), .A2(n12027), .ZN(n6706) );
  NAND2_X1 U8647 ( .A1(n14076), .A2(n11574), .ZN(n11630) );
  NAND2_X1 U8648 ( .A1(n14139), .A2(n11606), .ZN(n14118) );
  AND2_X1 U8649 ( .A1(n12024), .A2(n11531), .ZN(n7291) );
  NAND2_X1 U8650 ( .A1(n7292), .A2(n11531), .ZN(n14132) );
  NAND2_X1 U8651 ( .A1(n7276), .A2(n11492), .ZN(n11494) );
  NAND2_X1 U8652 ( .A1(n6691), .A2(n6692), .ZN(n11372) );
  NAND2_X1 U8653 ( .A1(n11197), .A2(n11196), .ZN(n11239) );
  OAI21_X1 U8654 ( .B1(n11054), .B2(n12011), .A(n7239), .ZN(n11171) );
  NAND2_X1 U8655 ( .A1(n7238), .A2(n11015), .ZN(n11170) );
  NAND2_X1 U8656 ( .A1(n7284), .A2(n10942), .ZN(n11013) );
  NAND2_X1 U8657 ( .A1(n14478), .A2(n14479), .ZN(n7284) );
  NAND2_X1 U8658 ( .A1(n14667), .A2(n10567), .ZN(n10957) );
  AOI21_X1 U8659 ( .B1(n10579), .B2(n10578), .A(n6489), .ZN(n7272) );
  INV_X1 U8660 ( .A(n7281), .ZN(n10503) );
  AOI21_X1 U8661 ( .B1(n14698), .B2(n14700), .A(n7282), .ZN(n7281) );
  AND2_X1 U8662 ( .A1(n7235), .A2(n7234), .ZN(n7236) );
  INV_X1 U8663 ( .A(n9751), .ZN(n7234) );
  INV_X1 U8664 ( .A(n14188), .ZN(n14704) );
  OR2_X1 U8665 ( .A1(n11775), .A2(n14725), .ZN(n11776) );
  INV_X1 U8666 ( .A(n14174), .ZN(n14483) );
  OR2_X1 U8667 ( .A1(n14231), .A2(n14230), .ZN(n14279) );
  AND2_X2 U8668 ( .A1(n9704), .A2(n10395), .ZN(n14787) );
  NAND2_X1 U8669 ( .A1(n7299), .A2(n6547), .ZN(n14287) );
  INV_X1 U8670 ( .A(n9325), .ZN(n7299) );
  OAI21_X1 U8671 ( .B1(n9339), .B2(n9299), .A(n6631), .ZN(n6775) );
  NOR2_X1 U8672 ( .A1(n9308), .A2(n6774), .ZN(n6773) );
  XNOR2_X1 U8673 ( .A(n9290), .B(n9289), .ZN(n9387) );
  INV_X1 U8674 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n9289) );
  NAND2_X1 U8675 ( .A1(n7120), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9290) );
  XNOR2_X1 U8676 ( .A(n9293), .B(n9292), .ZN(n12150) );
  XNOR2_X1 U8677 ( .A(n9322), .B(n9286), .ZN(n11979) );
  INV_X1 U8678 ( .A(n11978), .ZN(n11972) );
  NAND2_X1 U8679 ( .A1(n9302), .A2(n9336), .ZN(n9337) );
  INV_X1 U8680 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n10312) );
  INV_X1 U8681 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n10210) );
  INV_X1 U8682 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n10132) );
  INV_X1 U8683 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n9881) );
  XNOR2_X1 U8684 ( .A(n9878), .B(P1_IR_REG_14__SCAN_IN), .ZN(n14610) );
  INV_X1 U8685 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n10982) );
  INV_X1 U8686 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n9613) );
  INV_X1 U8687 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n9574) );
  INV_X1 U8688 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n9524) );
  AND2_X1 U8689 ( .A1(n9521), .A2(n9560), .ZN(n10563) );
  INV_X1 U8690 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n9517) );
  INV_X1 U8691 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n9479) );
  INV_X1 U8692 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n9472) );
  INV_X1 U8693 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n9464) );
  OR2_X1 U8694 ( .A1(n9372), .A2(n10128), .ZN(n9373) );
  NAND2_X1 U8695 ( .A1(n10128), .A2(n7074), .ZN(n7073) );
  INV_X1 U8696 ( .A(n7094), .ZN(n8933) );
  XNOR2_X1 U8697 ( .A(n8948), .B(n8947), .ZN(n15196) );
  XNOR2_X1 U8698 ( .A(n8956), .B(P2_ADDR_REG_7__SCAN_IN), .ZN(n15201) );
  XNOR2_X1 U8699 ( .A(n8961), .B(n8960), .ZN(n14323) );
  NOR2_X1 U8700 ( .A1(n14329), .A2(n8971), .ZN(n14543) );
  OR2_X1 U8701 ( .A1(n8986), .A2(n8985), .ZN(n14560) );
  NAND2_X1 U8702 ( .A1(n6831), .A2(n6835), .ZN(n8986) );
  INV_X1 U8703 ( .A(n6833), .ZN(n6832) );
  NAND2_X1 U8704 ( .A1(n14558), .A2(n14560), .ZN(n14342) );
  NAND2_X1 U8705 ( .A1(n10360), .A2(n9181), .ZN(n10659) );
  NAND2_X1 U8706 ( .A1(n11040), .A2(n9196), .ZN(n12421) );
  OAI21_X1 U8707 ( .B1(n8898), .B2(n15190), .A(n6984), .ZN(P3_U3488) );
  NOR2_X1 U8708 ( .A1(n6627), .A2(n6985), .ZN(n6984) );
  NOR2_X1 U8709 ( .A1(n15193), .A2(n8899), .ZN(n6985) );
  INV_X1 U8710 ( .A(n6805), .ZN(P3_U3487) );
  AOI21_X1 U8711 ( .B1(n7969), .B2(n15193), .A(n6806), .ZN(n6805) );
  OAI21_X1 U8712 ( .B1(n7970), .B2(n13179), .A(n6807), .ZN(n6806) );
  NAND2_X1 U8713 ( .A1(n15190), .A2(P3_REG1_REG_28__SCAN_IN), .ZN(n6807) );
  AOI21_X1 U8714 ( .B1(n8880), .B2(n13185), .A(n8882), .ZN(n8883) );
  MUX2_X1 U8715 ( .A(n13492), .B(n13491), .S(n13490), .Z(n13495) );
  NAND2_X1 U8716 ( .A1(n6910), .A2(n6649), .ZN(P1_U3525) );
  NAND2_X1 U8717 ( .A1(n14275), .A2(n14787), .ZN(n6910) );
  INV_X1 U8718 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n6909) );
  NOR2_X1 U8719 ( .A1(n14548), .A2(n14547), .ZN(n14546) );
  AND2_X1 U8720 ( .A1(n6825), .A2(n6535), .ZN(n14548) );
  NOR2_X1 U8721 ( .A1(n14556), .A2(n14555), .ZN(n14554) );
  AND2_X1 U8722 ( .A1(n6827), .A2(n6828), .ZN(n14556) );
  NAND2_X1 U8723 ( .A1(n14301), .A2(n14302), .ZN(n7083) );
  XNOR2_X1 U8724 ( .A(n6663), .B(n9164), .ZN(SUB_1596_U4) );
  NAND2_X1 U8725 ( .A1(n7086), .A2(n6664), .ZN(n6663) );
  OR2_X1 U8726 ( .A1(n13537), .A2(n13377), .ZN(n6486) );
  AND2_X1 U8727 ( .A1(n6938), .A2(n6553), .ZN(n6487) );
  INV_X1 U8728 ( .A(n12011), .ZN(n11015) );
  AND2_X1 U8729 ( .A1(n13719), .A2(n13377), .ZN(n12142) );
  NAND2_X1 U8730 ( .A1(n9412), .A2(n11781), .ZN(n9342) );
  INV_X1 U8731 ( .A(n10091), .ZN(n15051) );
  NAND2_X1 U8732 ( .A1(n9211), .A2(n13050), .ZN(n6488) );
  NOR2_X1 U8733 ( .A1(n11826), .A2(n13989), .ZN(n6489) );
  INV_X1 U8734 ( .A(P3_IR_REG_31__SCAN_IN), .ZN(n13241) );
  OR2_X1 U8735 ( .A1(n9233), .A2(n9232), .ZN(n6490) );
  OR2_X1 U8736 ( .A1(n13526), .A2(n13376), .ZN(n6491) );
  INV_X2 U8737 ( .A(n7574), .ZN(n7522) );
  AND2_X2 U8738 ( .A1(n11647), .A2(n7390), .ZN(n7422) );
  AND2_X1 U8739 ( .A1(n14226), .A2(n12275), .ZN(n11610) );
  OR2_X1 U8740 ( .A1(n8327), .A2(n8329), .ZN(n6492) );
  OR2_X1 U8741 ( .A1(n8903), .A2(n7090), .ZN(n6493) );
  INV_X1 U8742 ( .A(n11807), .ZN(n6904) );
  OR2_X1 U8743 ( .A1(n13747), .A2(n13597), .ZN(n6494) );
  NAND2_X2 U8744 ( .A1(n7404), .A2(n7403), .ZN(n8084) );
  AND2_X1 U8745 ( .A1(n13652), .A2(n6527), .ZN(n6495) );
  INV_X1 U8746 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n8012) );
  AND2_X1 U8747 ( .A1(n13772), .A2(n13383), .ZN(n6496) );
  AND2_X1 U8748 ( .A1(n11122), .A2(n6534), .ZN(n6497) );
  AND2_X1 U8749 ( .A1(n6915), .A2(n13905), .ZN(n6498) );
  AND2_X1 U8750 ( .A1(n7151), .A2(n6574), .ZN(n6499) );
  AND2_X1 U8751 ( .A1(n8607), .A2(n8606), .ZN(n6500) );
  INV_X1 U8752 ( .A(n13724), .ZN(n6955) );
  INV_X1 U8753 ( .A(n12026), .ZN(n14077) );
  INV_X1 U8754 ( .A(n13331), .ZN(n6993) );
  NAND2_X1 U8755 ( .A1(n8414), .A2(n8413), .ZN(n13784) );
  NOR2_X1 U8756 ( .A1(n13826), .A2(n12292), .ZN(n6501) );
  AND2_X1 U8757 ( .A1(n6883), .A2(n6880), .ZN(n6502) );
  INV_X1 U8758 ( .A(n11196), .ZN(n7290) );
  NAND2_X1 U8759 ( .A1(n8548), .A2(n8547), .ZN(n13747) );
  OR2_X1 U8760 ( .A1(n13784), .A2(n11329), .ZN(n6503) );
  INV_X1 U8761 ( .A(n7289), .ZN(n7288) );
  OAI21_X1 U8762 ( .B1(n11167), .B2(n7290), .A(n11238), .ZN(n7289) );
  INV_X1 U8763 ( .A(n8562), .ZN(n7215) );
  OR2_X1 U8764 ( .A1(n13526), .A2(n12143), .ZN(n6504) );
  AND2_X1 U8765 ( .A1(n7985), .A2(n7221), .ZN(n6505) );
  AND2_X1 U8766 ( .A1(n6995), .A2(n6562), .ZN(n6506) );
  INV_X1 U8767 ( .A(n13518), .ZN(n13522) );
  AND2_X1 U8768 ( .A1(n6912), .A2(n6911), .ZN(n6508) );
  AND2_X1 U8769 ( .A1(n9197), .A2(n9196), .ZN(n6509) );
  AND2_X1 U8770 ( .A1(n7019), .A2(n6551), .ZN(n6510) );
  INV_X1 U8771 ( .A(n7124), .ZN(n7123) );
  NAND2_X1 U8772 ( .A1(n7127), .A2(n7125), .ZN(n7124) );
  AND2_X1 U8773 ( .A1(n6795), .A2(n7720), .ZN(n6511) );
  INV_X1 U8774 ( .A(n9915), .ZN(n9921) );
  AND2_X1 U8775 ( .A1(n6922), .A2(n6647), .ZN(n6512) );
  NAND2_X1 U8776 ( .A1(n12840), .A2(P3_REG2_REG_18__SCAN_IN), .ZN(n6513) );
  CLKBUF_X3 U8777 ( .A(n8095), .Z(n8747) );
  XNOR2_X1 U8778 ( .A(n13920), .B(n14168), .ZN(n14138) );
  INV_X1 U8779 ( .A(n10891), .ZN(n12706) );
  NAND2_X1 U8780 ( .A1(n7687), .A2(n7344), .ZN(n6514) );
  NOR2_X1 U8781 ( .A1(n12954), .A2(n12751), .ZN(n6515) );
  NAND4_X1 U8782 ( .A1(n8099), .A2(n8098), .A3(n8097), .A4(n8096), .ZN(n8833)
         );
  NAND2_X1 U8783 ( .A1(n15130), .A2(n10204), .ZN(n7436) );
  INV_X1 U8784 ( .A(n7384), .ZN(n7925) );
  XNOR2_X1 U8785 ( .A(n14233), .B(n14121), .ZN(n14102) );
  INV_X1 U8786 ( .A(n14102), .ZN(n7265) );
  INV_X1 U8787 ( .A(n12031), .ZN(n6889) );
  AND2_X1 U8788 ( .A1(n6863), .A2(n6862), .ZN(n6516) );
  OR2_X1 U8789 ( .A1(n14075), .A2(n14085), .ZN(n6517) );
  AND2_X1 U8790 ( .A1(n12020), .A2(n11433), .ZN(n6518) );
  XNOR2_X1 U8791 ( .A(n14216), .B(n14069), .ZN(n12027) );
  INV_X1 U8792 ( .A(n12027), .ZN(n6739) );
  OR2_X1 U8793 ( .A1(n13231), .A2(n12332), .ZN(n6519) );
  AND2_X1 U8794 ( .A1(n6517), .A2(n6740), .ZN(n6520) );
  NAND2_X1 U8795 ( .A1(n11730), .A2(n13387), .ZN(n6521) );
  AND3_X1 U8796 ( .A1(n7440), .A2(n7439), .A3(n7438), .ZN(n6522) );
  NOR2_X1 U8797 ( .A1(n13283), .A2(n11745), .ZN(n6523) );
  NAND2_X1 U8798 ( .A1(n6782), .A2(n6783), .ZN(n6524) );
  INV_X1 U8799 ( .A(P3_IR_REG_27__SCAN_IN), .ZN(n7396) );
  NAND2_X1 U8800 ( .A1(n8609), .A2(n8608), .ZN(n6525) );
  AND4_X1 U8801 ( .A1(n7984), .A2(n7983), .A3(n7982), .A4(n7981), .ZN(n6526)
         );
  AND2_X1 U8802 ( .A1(n11867), .A2(n11866), .ZN(n12014) );
  NAND2_X1 U8803 ( .A1(n13490), .A2(n11649), .ZN(n8022) );
  INV_X1 U8804 ( .A(n11610), .ZN(n7268) );
  OR2_X1 U8805 ( .A1(n13656), .A2(n13763), .ZN(n6527) );
  NOR2_X1 U8806 ( .A1(n9209), .A2(n7037), .ZN(n6528) );
  AND2_X1 U8807 ( .A1(n8071), .A2(n8070), .ZN(n6529) );
  AND4_X1 U8808 ( .A1(n8853), .A2(n8852), .A3(n12144), .A4(n12117), .ZN(n6530)
         );
  AND2_X1 U8809 ( .A1(n6785), .A2(n7116), .ZN(n6531) );
  AND2_X1 U8810 ( .A1(n6859), .A2(n6858), .ZN(n6532) );
  AND2_X1 U8811 ( .A1(n6470), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n6533) );
  NAND2_X1 U8812 ( .A1(n8336), .A2(n8335), .ZN(n11281) );
  INV_X1 U8813 ( .A(n11281), .ZN(n7176) );
  OR2_X1 U8814 ( .A1(n11281), .A2(n13386), .ZN(n6534) );
  OR2_X1 U8815 ( .A1(n8978), .A2(n8977), .ZN(n6535) );
  OR2_X1 U8816 ( .A1(n7176), .A2(n13386), .ZN(n6536) );
  AND2_X1 U8817 ( .A1(n9601), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n6537) );
  NAND2_X1 U8818 ( .A1(n7246), .A2(n12019), .ZN(n11603) );
  OR3_X1 U8819 ( .A1(P3_IR_REG_2__SCAN_IN), .A2(P3_IR_REG_1__SCAN_IN), .A3(
        P3_IR_REG_0__SCAN_IN), .ZN(n6538) );
  INV_X1 U8820 ( .A(n12024), .ZN(n14131) );
  INV_X1 U8821 ( .A(n11949), .ZN(n7297) );
  INV_X1 U8822 ( .A(n11910), .ZN(n7319) );
  INV_X1 U8823 ( .A(n12012), .ZN(n11238) );
  AND2_X1 U8824 ( .A1(n12573), .A2(n12563), .ZN(n6539) );
  AND2_X1 U8825 ( .A1(n12985), .A2(n12641), .ZN(n13000) );
  NAND2_X1 U8826 ( .A1(n13834), .A2(n13833), .ZN(n6540) );
  AND2_X1 U8827 ( .A1(n13694), .A2(n14986), .ZN(n6541) );
  NAND2_X1 U8828 ( .A1(n11586), .A2(n11585), .ZN(n14209) );
  NOR2_X1 U8829 ( .A1(n12220), .A2(n7118), .ZN(n6542) );
  XNOR2_X1 U8830 ( .A(n12535), .B(n12746), .ZN(n12534) );
  OR2_X1 U8831 ( .A1(n12933), .A2(n12930), .ZN(n6543) );
  AND2_X1 U8832 ( .A1(n8247), .A2(n8246), .ZN(n6544) );
  AND2_X1 U8833 ( .A1(n6506), .A2(n10768), .ZN(n6545) );
  OR2_X1 U8834 ( .A1(n12203), .A2(n12201), .ZN(n6546) );
  INV_X1 U8835 ( .A(n11939), .ZN(n7322) );
  INV_X1 U8836 ( .A(n7450), .ZN(n6973) );
  NOR2_X1 U8837 ( .A1(P1_IR_REG_28__SCAN_IN), .A2(P1_IR_REG_29__SCAN_IN), .ZN(
        n6547) );
  INV_X1 U8838 ( .A(n10320), .ZN(n7133) );
  INV_X1 U8839 ( .A(n13905), .ZN(n14256) );
  AND2_X1 U8840 ( .A1(n11472), .A2(n11471), .ZN(n13905) );
  INV_X1 U8841 ( .A(P3_ADDR_REG_3__SCAN_IN), .ZN(n7090) );
  NOR2_X1 U8842 ( .A1(n7350), .A2(n13846), .ZN(n6548) );
  AND2_X1 U8843 ( .A1(n14106), .A2(n7266), .ZN(n6549) );
  AND2_X1 U8844 ( .A1(n11375), .A2(n11374), .ZN(n12209) );
  INV_X1 U8845 ( .A(n12209), .ZN(n14270) );
  AND2_X1 U8846 ( .A1(n13329), .A2(n11740), .ZN(n6550) );
  INV_X1 U8847 ( .A(n6835), .ZN(n6834) );
  NAND2_X1 U8848 ( .A1(n14555), .A2(P2_ADDR_REG_15__SCAN_IN), .ZN(n6835) );
  OR2_X1 U8849 ( .A1(n9218), .A2(n13002), .ZN(n6551) );
  INV_X1 U8850 ( .A(n12184), .ZN(n14506) );
  NAND2_X1 U8851 ( .A1(n11166), .A2(n11165), .ZN(n12184) );
  INV_X1 U8852 ( .A(P3_IR_REG_29__SCAN_IN), .ZN(n6854) );
  AND2_X1 U8853 ( .A1(n13784), .A2(n11329), .ZN(n6552) );
  OR2_X1 U8854 ( .A1(n8346), .A2(SI_13_), .ZN(n6553) );
  AND2_X1 U8855 ( .A1(n8330), .A2(n9489), .ZN(n6554) );
  OR2_X1 U8856 ( .A1(n8632), .A2(n8631), .ZN(n6555) );
  NAND2_X1 U8857 ( .A1(n11323), .A2(n11322), .ZN(n6556) );
  AND2_X1 U8858 ( .A1(n9188), .A2(n9187), .ZN(n6557) );
  AND2_X1 U8859 ( .A1(n6852), .A2(n6849), .ZN(n6558) );
  INV_X1 U8860 ( .A(n7031), .ZN(n7029) );
  AND2_X1 U8861 ( .A1(n12490), .A2(n12332), .ZN(n7031) );
  NAND2_X1 U8862 ( .A1(n8744), .A2(n8743), .ZN(n13700) );
  AND2_X1 U8863 ( .A1(n13167), .A2(n12757), .ZN(n6559) );
  AND2_X1 U8864 ( .A1(n14209), .A2(n11611), .ZN(n6560) );
  INV_X1 U8865 ( .A(n7169), .ZN(n7168) );
  NAND2_X1 U8866 ( .A1(n7170), .A2(n11125), .ZN(n7169) );
  INV_X1 U8867 ( .A(n6958), .ZN(n13585) );
  AND2_X1 U8868 ( .A1(n11860), .A2(n11861), .ZN(n6561) );
  NAND2_X1 U8869 ( .A1(n10766), .A2(n10765), .ZN(n6562) );
  OR2_X1 U8870 ( .A1(n8948), .A2(n8947), .ZN(n6563) );
  AND2_X1 U8871 ( .A1(n11521), .A2(n11519), .ZN(n6564) );
  AND2_X1 U8872 ( .A1(n13518), .A2(n6499), .ZN(n6565) );
  NOR2_X1 U8873 ( .A1(n14216), .A2(n14069), .ZN(n6566) );
  INV_X1 U8874 ( .A(n7295), .ZN(n7294) );
  NAND2_X1 U8875 ( .A1(n6739), .A2(n11574), .ZN(n7295) );
  NOR2_X1 U8876 ( .A1(n11869), .A2(n7316), .ZN(n6567) );
  NOR2_X1 U8877 ( .A1(n11849), .A2(n14456), .ZN(n6568) );
  NOR2_X1 U8878 ( .A1(n14498), .A2(n13983), .ZN(n6569) );
  NOR2_X1 U8879 ( .A1(n7951), .A2(n7931), .ZN(n6570) );
  OR2_X1 U8880 ( .A1(n9229), .A2(n9228), .ZN(n6571) );
  OR2_X1 U8881 ( .A1(n6525), .A2(n6500), .ZN(n6572) );
  AND2_X1 U8882 ( .A1(n8346), .A2(SI_13_), .ZN(n6573) );
  NAND2_X1 U8883 ( .A1(n13537), .A2(n13305), .ZN(n6574) );
  AND2_X1 U8884 ( .A1(n7872), .A2(n7870), .ZN(n6575) );
  INV_X1 U8885 ( .A(n8009), .ZN(n7008) );
  NOR2_X1 U8886 ( .A1(n7014), .A2(n9245), .ZN(n6576) );
  AND2_X1 U8887 ( .A1(n12665), .A2(n6975), .ZN(n6577) );
  AND2_X1 U8888 ( .A1(n8253), .A2(SI_9_), .ZN(n6578) );
  NOR2_X1 U8889 ( .A1(n14778), .A2(n10956), .ZN(n6579) );
  OR2_X1 U8890 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(n8956), .ZN(n6580) );
  INV_X1 U8891 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n13808) );
  NAND2_X1 U8892 ( .A1(n13752), .A2(n13658), .ZN(n6581) );
  NAND2_X1 U8893 ( .A1(n8682), .A2(n8683), .ZN(n6582) );
  NAND2_X1 U8894 ( .A1(n11517), .A2(n11516), .ZN(n14252) );
  AND2_X1 U8895 ( .A1(n12954), .A2(n12751), .ZN(n6583) );
  INV_X1 U8896 ( .A(n12142), .ZN(n7150) );
  NOR2_X1 U8897 ( .A1(P2_IR_REG_28__SCAN_IN), .A2(P2_IR_REG_29__SCAN_IN), .ZN(
        n6585) );
  NOR2_X1 U8898 ( .A1(n7176), .A2(n11282), .ZN(n6586) );
  NAND2_X1 U8899 ( .A1(n13752), .A2(n13624), .ZN(n6587) );
  AOI21_X1 U8900 ( .B1(n7112), .B2(n7111), .A(n7365), .ZN(n7110) );
  INV_X1 U8901 ( .A(n11790), .ZN(n7233) );
  NAND2_X1 U8902 ( .A1(n11459), .A2(n11457), .ZN(n6588) );
  NAND2_X1 U8903 ( .A1(n6739), .A2(n6740), .ZN(n6738) );
  OR2_X1 U8904 ( .A1(n9210), .A2(n7035), .ZN(n6589) );
  NAND2_X1 U8905 ( .A1(n7116), .A2(n13902), .ZN(n6590) );
  INV_X1 U8906 ( .A(n11950), .ZN(n6676) );
  AND2_X1 U8907 ( .A1(n7002), .A2(n11725), .ZN(n6591) );
  OR2_X1 U8908 ( .A1(n11743), .A2(n11742), .ZN(n6592) );
  OR2_X1 U8909 ( .A1(n8904), .A2(n15056), .ZN(n6593) );
  AND2_X1 U8910 ( .A1(n6967), .A2(n7573), .ZN(n6594) );
  AND2_X1 U8911 ( .A1(n6892), .A2(n6890), .ZN(n6595) );
  NOR2_X1 U8912 ( .A1(n10825), .A2(n7113), .ZN(n7112) );
  INV_X1 U8913 ( .A(n11602), .ZN(n7245) );
  AND2_X1 U8914 ( .A1(n11993), .A2(n12039), .ZN(n6596) );
  AND2_X1 U8915 ( .A1(n7412), .A2(n7413), .ZN(n6597) );
  NAND2_X1 U8916 ( .A1(n12203), .A2(n12201), .ZN(n6598) );
  NOR2_X1 U8917 ( .A1(n14206), .A2(n14205), .ZN(n6599) );
  AND2_X1 U8918 ( .A1(n6945), .A2(n6946), .ZN(n6600) );
  INV_X1 U8919 ( .A(n11606), .ZN(n7249) );
  AND2_X1 U8920 ( .A1(n12650), .A2(n12651), .ZN(n12971) );
  NOR2_X1 U8921 ( .A1(n7890), .A2(n7341), .ZN(n7340) );
  AND2_X1 U8922 ( .A1(n8500), .A2(n8499), .ZN(n6601) );
  AND2_X1 U8923 ( .A1(n8560), .A2(n8559), .ZN(n6602) );
  AND2_X1 U8924 ( .A1(n9182), .A2(n9181), .ZN(n6603) );
  AND2_X1 U8925 ( .A1(n12115), .A2(n6494), .ZN(n6604) );
  AND2_X1 U8926 ( .A1(n7376), .A2(n6841), .ZN(n6605) );
  OR2_X1 U8927 ( .A1(n7297), .A2(n11948), .ZN(n6606) );
  OR2_X1 U8928 ( .A1(n7319), .A2(n11909), .ZN(n6607) );
  OR2_X1 U8929 ( .A1(n11837), .A2(n11835), .ZN(n6608) );
  OR2_X1 U8930 ( .A1(n11848), .A2(n11846), .ZN(n6609) );
  OR2_X1 U8931 ( .A1(n7219), .A2(n7220), .ZN(n6610) );
  INV_X1 U8932 ( .A(n10432), .ZN(n7282) );
  OR2_X1 U8933 ( .A1(n7322), .A2(n11938), .ZN(n6611) );
  INV_X1 U8934 ( .A(n7161), .ZN(n7160) );
  OAI21_X1 U8935 ( .B1(n13637), .B2(n13636), .A(n6581), .ZN(n7161) );
  OR2_X1 U8936 ( .A1(n8321), .A2(n8323), .ZN(n6612) );
  OR2_X1 U8937 ( .A1(n7303), .A2(n11836), .ZN(n6613) );
  OR2_X1 U8938 ( .A1(n8322), .A2(n8324), .ZN(n6614) );
  OR2_X1 U8939 ( .A1(n8854), .A2(n7367), .ZN(n6615) );
  NAND2_X1 U8940 ( .A1(n8901), .A2(P3_ADDR_REG_1__SCAN_IN), .ZN(n6616) );
  AND2_X1 U8941 ( .A1(n12247), .A2(n6783), .ZN(n6617) );
  INV_X1 U8942 ( .A(n12017), .ZN(n14165) );
  NAND2_X1 U8943 ( .A1(n7214), .A2(n7215), .ZN(n6618) );
  NAND2_X1 U8944 ( .A1(n7217), .A2(n8501), .ZN(n6619) );
  AND2_X1 U8945 ( .A1(n6585), .A2(n6505), .ZN(n6620) );
  INV_X1 U8946 ( .A(P3_IR_REG_1__SCAN_IN), .ZN(n6686) );
  INV_X1 U8947 ( .A(n6497), .ZN(n7137) );
  OR2_X1 U8948 ( .A1(n13495), .A2(n13494), .ZN(P2_U3233) );
  INV_X1 U8949 ( .A(n15089), .ZN(n10714) );
  NAND2_X1 U8950 ( .A1(n7040), .A2(n8868), .ZN(n8880) );
  NAND2_X1 U8951 ( .A1(n7018), .A2(n7022), .ZN(n12396) );
  INV_X1 U8952 ( .A(n13729), .ZN(n6957) );
  NAND2_X1 U8953 ( .A1(n11738), .A2(n11737), .ZN(n13311) );
  NAND2_X1 U8954 ( .A1(n6498), .A2(n11387), .ZN(n6622) );
  NAND2_X1 U8955 ( .A1(n7276), .A2(n7275), .ZN(n11513) );
  INV_X1 U8956 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n9450) );
  AND2_X1 U8957 ( .A1(n11413), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n6623) );
  AND2_X1 U8958 ( .A1(n11007), .A2(n6914), .ZN(n6624) );
  INV_X1 U8959 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n6868) );
  INV_X1 U8960 ( .A(n10160), .ZN(n10155) );
  INV_X1 U8961 ( .A(n10699), .ZN(n10709) );
  INV_X1 U8962 ( .A(n13684), .ZN(n12132) );
  NAND2_X2 U8963 ( .A1(n7391), .A2(n11667), .ZN(n7468) );
  NAND2_X1 U8964 ( .A1(n8558), .A2(n8557), .ZN(n13643) );
  NAND2_X1 U8965 ( .A1(n8650), .A2(n8649), .ZN(n13378) );
  INV_X1 U8966 ( .A(n13378), .ZN(n7152) );
  AND2_X1 U8967 ( .A1(n11732), .A2(n7003), .ZN(n6625) );
  AND2_X1 U8968 ( .A1(n14513), .A2(n11162), .ZN(n6626) );
  INV_X1 U8969 ( .A(n7056), .ZN(n7055) );
  OAI21_X1 U8970 ( .B1(n7664), .B2(n7057), .A(n7701), .ZN(n7056) );
  INV_X1 U8971 ( .A(n7026), .ZN(n7024) );
  AND2_X1 U8972 ( .A1(n8880), .A2(n8900), .ZN(n6627) );
  OR2_X1 U8973 ( .A1(n12770), .A2(n14426), .ZN(n6628) );
  AND2_X1 U8974 ( .A1(n11416), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n6629) );
  AND2_X1 U8975 ( .A1(n7733), .A2(n7719), .ZN(n7720) );
  AND2_X1 U8976 ( .A1(n6990), .A2(n6991), .ZN(n6630) );
  AND2_X1 U8977 ( .A1(P1_IR_REG_26__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), .ZN(
        n6631) );
  AND2_X1 U8978 ( .A1(n11434), .A2(n11433), .ZN(n6632) );
  INV_X1 U8979 ( .A(P3_IR_REG_0__SCAN_IN), .ZN(n6876) );
  INV_X1 U8980 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n9292) );
  NAND2_X1 U8981 ( .A1(n11762), .A2(n6996), .ZN(n6994) );
  OR2_X1 U8982 ( .A1(n8709), .A2(SI_28_), .ZN(n6633) );
  INV_X1 U8983 ( .A(n13763), .ZN(n6953) );
  AND2_X2 U8984 ( .A1(n10026), .A2(n7968), .ZN(n15193) );
  NOR2_X1 U8985 ( .A1(n11130), .A2(n10865), .ZN(n6634) );
  INV_X1 U8986 ( .A(SI_14_), .ZN(n6890) );
  NAND2_X1 U8987 ( .A1(n8488), .A2(n8487), .ZN(n13757) );
  INV_X1 U8988 ( .A(n13757), .ZN(n6951) );
  INV_X1 U8989 ( .A(n14498), .ZN(n6911) );
  NAND2_X1 U8990 ( .A1(n10460), .A2(n10459), .ZN(n10579) );
  NAND2_X1 U8991 ( .A1(n10447), .A2(n10446), .ZN(n14682) );
  INV_X1 U8992 ( .A(n7272), .ZN(n14663) );
  AOI21_X1 U8993 ( .B1(n8759), .B2(n6633), .A(n6925), .ZN(n6924) );
  OR2_X1 U8994 ( .A1(n10652), .A2(n10651), .ZN(n6635) );
  NAND2_X1 U8995 ( .A1(n6844), .A2(n6967), .ZN(n13111) );
  NOR2_X1 U8996 ( .A1(n15079), .A2(n10695), .ZN(n6636) );
  INV_X1 U8997 ( .A(P3_ADDR_REG_7__SCAN_IN), .ZN(n7095) );
  AND2_X1 U8998 ( .A1(n6771), .A2(n13921), .ZN(n6637) );
  AND2_X1 U8999 ( .A1(n6994), .A2(n6995), .ZN(n6638) );
  AND2_X1 U9000 ( .A1(n8686), .A2(n11202), .ZN(n6639) );
  NAND2_X1 U9001 ( .A1(n9303), .A2(n9295), .ZN(n6640) );
  AND2_X1 U9002 ( .A1(n8711), .A2(n11670), .ZN(n6641) );
  INV_X1 U9003 ( .A(SI_17_), .ZN(n9764) );
  AND2_X1 U9004 ( .A1(n11651), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n6642) );
  INV_X1 U9005 ( .A(n12802), .ZN(n12793) );
  AND2_X1 U9006 ( .A1(n6635), .A2(n10740), .ZN(n6643) );
  OR2_X1 U9007 ( .A1(n12818), .A2(n7182), .ZN(n6644) );
  INV_X1 U9008 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n9295) );
  AND2_X1 U9009 ( .A1(n8684), .A2(SI_26_), .ZN(n6645) );
  OR2_X1 U9010 ( .A1(n15101), .A2(n7190), .ZN(n6646) );
  INV_X1 U9011 ( .A(n11413), .ZN(n6856) );
  BUF_X1 U9012 ( .A(n8836), .Z(n13396) );
  INV_X1 U9013 ( .A(n8836), .ZN(n7122) );
  NAND2_X1 U9014 ( .A1(n8002), .A2(n8001), .ZN(n8820) );
  XOR2_X1 U9015 ( .A(n8712), .B(SI_30_), .Z(n6647) );
  INV_X1 U9016 ( .A(n14361), .ZN(n12842) );
  AND2_X1 U9017 ( .A1(n14042), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n6648) );
  OR2_X1 U9018 ( .A1(n14787), .A2(n6909), .ZN(n6649) );
  AND2_X1 U9019 ( .A1(n7188), .A2(n7187), .ZN(n6650) );
  INV_X1 U9020 ( .A(n6905), .ZN(n14710) );
  NOR2_X1 U9021 ( .A1(n9890), .A2(n11798), .ZN(n6905) );
  NOR2_X1 U9022 ( .A1(n8713), .A2(n12522), .ZN(n6651) );
  INV_X1 U9023 ( .A(n14988), .ZN(n14996) );
  INV_X1 U9024 ( .A(n10434), .ZN(n6869) );
  INV_X1 U9025 ( .A(n12825), .ZN(n12857) );
  INV_X1 U9026 ( .A(P3_REG2_REG_16__SCAN_IN), .ZN(n7204) );
  AND2_X1 U9027 ( .A1(n12837), .A2(n6513), .ZN(n6652) );
  INV_X1 U9028 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n8902) );
  INV_X1 U9029 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n7399) );
  INV_X1 U9030 ( .A(P1_RD_REG_SCAN_IN), .ZN(n7398) );
  AND2_X1 U9031 ( .A1(n9412), .A2(n9486), .ZN(n12057) );
  OR2_X1 U9032 ( .A1(n10253), .A2(n10299), .ZN(n10323) );
  XNOR2_X1 U9033 ( .A(n6485), .B(n10299), .ZN(n11706) );
  NAND2_X1 U9034 ( .A1(n6653), .A2(n7406), .ZN(n7409) );
  NAND2_X1 U9035 ( .A1(n7405), .A2(n7433), .ZN(n6653) );
  OR2_X1 U9036 ( .A1(n12693), .A2(n12692), .ZN(n7068) );
  INV_X1 U9037 ( .A(n7611), .ZN(n6808) );
  INV_X1 U9038 ( .A(n12694), .ZN(n12697) );
  NAND2_X1 U9039 ( .A1(n6792), .A2(n6790), .ZN(n7735) );
  NAND2_X1 U9040 ( .A1(n7599), .A2(n7598), .ZN(n7610) );
  NAND2_X1 U9041 ( .A1(n7786), .A2(n7785), .ZN(n7787) );
  NAND3_X1 U9042 ( .A1(n8535), .A2(n8536), .A3(n6618), .ZN(n6684) );
  OR2_X1 U9043 ( .A1(n8428), .A2(n8432), .ZN(n8459) );
  NAND2_X1 U9044 ( .A1(n8633), .A2(n6555), .ZN(n8655) );
  NAND2_X1 U9045 ( .A1(n8272), .A2(n6654), .ZN(n8303) );
  OAI22_X1 U9046 ( .A1(n7229), .A2(n8656), .B1(n8682), .B2(n8683), .ZN(n8783)
         );
  OR2_X2 U9047 ( .A1(n9920), .A2(n10976), .ZN(n8531) );
  XNOR2_X2 U9048 ( .A(n8019), .B(P2_IR_REG_19__SCAN_IN), .ZN(n13490) );
  OAI21_X1 U9049 ( .B1(n8149), .B2(n8148), .A(n6610), .ZN(n6680) );
  NAND2_X1 U9050 ( .A1(n6658), .A2(n6657), .ZN(n8046) );
  NAND2_X1 U9051 ( .A1(n7008), .A2(n8462), .ZN(n8018) );
  OAI21_X1 U9052 ( .B1(n8479), .B2(n8478), .A(n8477), .ZN(n8481) );
  AOI21_X1 U9053 ( .B1(n6671), .B2(n6670), .A(n6615), .ZN(n6669) );
  NAND3_X1 U9054 ( .A1(n8026), .A2(n8024), .A3(n8025), .ZN(n6658) );
  NAND2_X1 U9055 ( .A1(n10216), .A2(n9832), .ZN(n8014) );
  INV_X1 U9056 ( .A(n8859), .ZN(n6671) );
  OAI21_X1 U9057 ( .B1(n8147), .B2(n6680), .A(n7218), .ZN(n8204) );
  XNOR2_X2 U9058 ( .A(n6659), .B(n9309), .ZN(n9428) );
  NAND3_X1 U9059 ( .A1(n11947), .A2(n11946), .A3(n6606), .ZN(n6660) );
  OAI21_X1 U9060 ( .B1(n11906), .B2(n11905), .A(n11904), .ZN(n11908) );
  NAND2_X1 U9061 ( .A1(n6990), .A2(n6988), .ZN(n13275) );
  NOR2_X1 U9062 ( .A1(n10039), .A2(n7364), .ZN(n13269) );
  OAI21_X2 U9063 ( .B1(n8009), .B2(n8010), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n8013) );
  NAND2_X1 U9064 ( .A1(n11736), .A2(n11735), .ZN(n13313) );
  NAND2_X2 U9065 ( .A1(n7771), .A2(n12660), .ZN(n12931) );
  NAND2_X2 U9066 ( .A1(n12931), .A2(n12930), .ZN(n12929) );
  AOI211_X2 U9067 ( .C1(n12687), .C2(n12528), .A(n12722), .B(n12527), .ZN(
        n12532) );
  NAND2_X1 U9068 ( .A1(n7608), .A2(n12611), .ZN(n13071) );
  NAND2_X1 U9069 ( .A1(n12882), .A2(n7920), .ZN(n7969) );
  NAND3_X2 U9070 ( .A1(n7459), .A2(n7458), .A3(n6661), .ZN(n12762) );
  INV_X1 U9071 ( .A(n13270), .ZN(n10238) );
  NAND2_X1 U9072 ( .A1(n13631), .A2(n13621), .ZN(n13603) );
  NAND2_X1 U9073 ( .A1(n13349), .A2(n12082), .ZN(n12088) );
  OR2_X1 U9074 ( .A1(n8015), .A2(n13808), .ZN(n8011) );
  INV_X1 U9075 ( .A(n11324), .ZN(n6662) );
  INV_X1 U9076 ( .A(n9931), .ZN(n9938) );
  NAND2_X2 U9077 ( .A1(n12096), .A2(n13299), .ZN(n12101) );
  NAND2_X1 U9078 ( .A1(n11738), .A2(n6992), .ZN(n6990) );
  NAND2_X1 U9079 ( .A1(n7428), .A2(P3_IR_REG_1__SCAN_IN), .ZN(n6687) );
  NOR2_X1 U9080 ( .A1(n14374), .A2(n7203), .ZN(n12822) );
  XNOR2_X1 U9081 ( .A(n11649), .B(n9832), .ZN(n9833) );
  NOR2_X1 U9082 ( .A1(n9772), .A2(n9786), .ZN(n10086) );
  OAI21_X2 U9083 ( .B1(n10596), .B2(n10547), .A(n10595), .ZN(n11762) );
  OAI22_X1 U9084 ( .A1(n8928), .A2(n8917), .B1(P1_ADDR_REG_13__SCAN_IN), .B2(
        n8916), .ZN(n8926) );
  NAND2_X1 U9085 ( .A1(n7094), .A2(n7093), .ZN(n7092) );
  NAND2_X1 U9086 ( .A1(n7081), .A2(n7080), .ZN(n7079) );
  AOI21_X1 U9087 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(n12800), .A(n8918), .ZN(
        n8981) );
  INV_X1 U9088 ( .A(n7098), .ZN(n8911) );
  NOR2_X1 U9089 ( .A1(n8976), .A2(n8975), .ZN(n8915) );
  NOR2_X1 U9090 ( .A1(n8910), .A2(n8909), .ZN(n8958) );
  OR2_X1 U9091 ( .A1(n8958), .A2(n8957), .ZN(n7101) );
  NOR2_X1 U9092 ( .A1(n8968), .A2(n8967), .ZN(n8912) );
  XNOR2_X2 U9093 ( .A(n8058), .B(P2_IR_REG_2__SCAN_IN), .ZN(n14807) );
  NAND2_X1 U9094 ( .A1(n12328), .A2(n12329), .ZN(n12327) );
  NOR2_X4 U9095 ( .A1(P3_IR_REG_1__SCAN_IN), .A2(P3_IR_REG_0__SCAN_IN), .ZN(
        n10087) );
  NAND2_X1 U9096 ( .A1(n10362), .A2(n10361), .ZN(n10360) );
  AOI22_X1 U9097 ( .A1(n12469), .A2(n12470), .B1(n9220), .B2(n12755), .ZN(
        n12357) );
  INV_X4 U9098 ( .A(n9178), .ZN(n11671) );
  NAND2_X1 U9099 ( .A1(n6665), .A2(n6613), .ZN(n11840) );
  NAND3_X1 U9100 ( .A1(n11834), .A2(n11833), .A3(n6608), .ZN(n6665) );
  NAND2_X1 U9101 ( .A1(n6666), .A2(n7302), .ZN(n11852) );
  NAND3_X1 U9102 ( .A1(n11845), .A2(n11844), .A3(n6609), .ZN(n6666) );
  NAND2_X1 U9103 ( .A1(n9337), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9338) );
  NAND2_X1 U9104 ( .A1(n6667), .A2(n7318), .ZN(n11913) );
  NAND3_X1 U9105 ( .A1(n11908), .A2(n11907), .A3(n6607), .ZN(n6667) );
  OAI21_X2 U9106 ( .B1(n11894), .B2(n11893), .A(n11892), .ZN(n11895) );
  NAND2_X1 U9107 ( .A1(n11973), .A2(n12035), .ZN(n11777) );
  NAND2_X1 U9108 ( .A1(n11825), .A2(n11824), .ZN(n11829) );
  AOI21_X1 U9109 ( .B1(n12859), .B2(n15064), .A(n6881), .ZN(n6880) );
  NAND2_X1 U9111 ( .A1(n7309), .A2(n11815), .ZN(n7308) );
  NAND3_X1 U9112 ( .A1(n8860), .A2(n8855), .A3(n6669), .ZN(P2_U3328) );
  NAND2_X1 U9113 ( .A1(n6682), .A2(n6681), .ZN(n8530) );
  OAI21_X1 U9114 ( .B1(n8094), .B2(n8093), .A(n6672), .ZN(n8121) );
  NAND2_X1 U9115 ( .A1(n6674), .A2(n6673), .ZN(n6672) );
  NAND2_X1 U9116 ( .A1(n8094), .A2(n8093), .ZN(n6674) );
  XNOR2_X1 U9117 ( .A(n9178), .B(n15107), .ZN(n9175) );
  OAI21_X2 U9118 ( .B1(n12384), .B2(n12386), .A(n12385), .ZN(n12383) );
  NAND2_X2 U9119 ( .A1(n12383), .A2(n9241), .ZN(n12482) );
  OAI21_X1 U9120 ( .B1(n12357), .B2(n12356), .A(n9222), .ZN(n12431) );
  AOI21_X1 U9121 ( .B1(n10289), .B2(n10290), .A(n9177), .ZN(n10362) );
  NAND2_X1 U9122 ( .A1(n8136), .A2(n8135), .ZN(n6675) );
  NAND2_X1 U9123 ( .A1(n8373), .A2(n8374), .ZN(n6900) );
  NAND2_X1 U9124 ( .A1(n8084), .A2(n9437), .ZN(n8031) );
  NAND2_X1 U9125 ( .A1(n8349), .A2(n6933), .ZN(n8410) );
  OR2_X2 U9126 ( .A1(n13603), .A2(n13740), .ZN(n13601) );
  INV_X1 U9127 ( .A(n6677), .ZN(n10786) );
  NOR2_X4 U9128 ( .A1(n13515), .A2(n13706), .ZN(n13509) );
  AND2_X1 U9129 ( .A1(n10013), .A2(n10143), .ZN(n9951) );
  NAND2_X1 U9130 ( .A1(n6958), .A2(n6957), .ZN(n13554) );
  NAND3_X1 U9131 ( .A1(n13704), .A2(n13702), .A3(n6678), .ZN(n13791) );
  NAND2_X4 U9132 ( .A1(n8056), .A2(n11519), .ZN(n8762) );
  NOR2_X1 U9133 ( .A1(n8530), .A2(n8529), .ZN(n8528) );
  NAND2_X1 U9134 ( .A1(n6684), .A2(n6683), .ZN(n8584) );
  AOI21_X1 U9135 ( .B1(n8149), .B2(n8148), .A(n8146), .ZN(n8147) );
  NAND2_X1 U9136 ( .A1(n8303), .A2(n8304), .ZN(n8302) );
  NAND3_X1 U9137 ( .A1(n8481), .A2(n8480), .A3(n6619), .ZN(n6682) );
  NAND2_X1 U9138 ( .A1(n7216), .A2(n6612), .ZN(n8431) );
  NAND2_X1 U9139 ( .A1(n7213), .A2(n7212), .ZN(n8094) );
  NOR2_X1 U9140 ( .A1(n15058), .A2(n10072), .ZN(n15057) );
  NAND4_X1 U9141 ( .A1(n14408), .A2(n14410), .A3(n14409), .A4(n14411), .ZN(
        P3_U3200) );
  NOR2_X2 U9142 ( .A1(n10693), .A2(n6688), .ZN(n10694) );
  XNOR2_X1 U9143 ( .A(n12785), .B(n12802), .ZN(n12768) );
  NOR2_X2 U9144 ( .A1(n12823), .A2(n14389), .ZN(n14406) );
  NOR2_X1 U9145 ( .A1(n15020), .A2(n10090), .ZN(n15046) );
  NAND2_X2 U9146 ( .A1(n6689), .A2(n14082), .ZN(n14096) );
  OAI21_X1 U9147 ( .B1(n10447), .B2(n12002), .A(n6695), .ZN(n6694) );
  NAND2_X1 U9148 ( .A1(n6694), .A2(n7273), .ZN(n10581) );
  NAND2_X1 U9149 ( .A1(n6699), .A2(n6698), .ZN(n11016) );
  NAND2_X1 U9150 ( .A1(n14478), .A2(n6701), .ZN(n6698) );
  OAI21_X1 U9151 ( .B1(n7283), .B2(n6703), .A(n11014), .ZN(n6700) );
  NOR2_X1 U9152 ( .A1(n6704), .A2(n6703), .ZN(n6701) );
  NAND2_X1 U9153 ( .A1(n6702), .A2(n7283), .ZN(n11048) );
  NAND2_X1 U9154 ( .A1(n14478), .A2(n7285), .ZN(n6702) );
  INV_X1 U9155 ( .A(n12009), .ZN(n6703) );
  INV_X1 U9156 ( .A(n7285), .ZN(n6704) );
  AND2_X2 U9157 ( .A1(n9302), .A2(n9301), .ZN(n9308) );
  AND2_X2 U9158 ( .A1(n6706), .A2(n11629), .ZN(n14219) );
  OAI21_X1 U9159 ( .B1(n13531), .B2(n6711), .A(n6709), .ZN(n13506) );
  NAND2_X1 U9160 ( .A1(n13675), .A2(n12114), .ZN(n6723) );
  NAND2_X1 U9161 ( .A1(n6723), .A2(n6722), .ZN(n6725) );
  CLKBUF_X1 U9162 ( .A(n6723), .Z(n6721) );
  NOR2_X1 U9163 ( .A1(n13595), .A2(n13596), .ZN(n13593) );
  NAND2_X1 U9164 ( .A1(n6727), .A2(n11607), .ZN(n14103) );
  NAND2_X1 U9165 ( .A1(n6728), .A2(n7247), .ZN(n6727) );
  NAND2_X1 U9166 ( .A1(n14141), .A2(n11606), .ZN(n6728) );
  NAND2_X2 U9167 ( .A1(n11053), .A2(n6703), .ZN(n11054) );
  OR2_X2 U9168 ( .A1(n14067), .A2(n14077), .ZN(n6741) );
  INV_X1 U9169 ( .A(n6730), .ZN(n7231) );
  OAI21_X1 U9170 ( .B1(n14067), .B2(n6733), .A(n6731), .ZN(n6730) );
  AND2_X2 U9171 ( .A1(n8811), .A2(n6505), .ZN(n8000) );
  AND4_X2 U9172 ( .A1(n7980), .A2(n6526), .A3(n6747), .A4(n8101), .ZN(n8811)
         );
  AND4_X2 U9173 ( .A1(n7979), .A2(n7977), .A3(n7978), .A4(n7976), .ZN(n7980)
         );
  NAND3_X1 U9174 ( .A1(n6749), .A2(n10620), .A3(n6748), .ZN(n10621) );
  OAI211_X1 U9175 ( .C1(n7137), .C2(n6755), .A(n6753), .B(n7135), .ZN(n11297)
         );
  INV_X1 U9176 ( .A(n7363), .ZN(n6757) );
  OAI21_X1 U9177 ( .B1(n6757), .B2(n7124), .A(n6758), .ZN(n11313) );
  AND2_X1 U9178 ( .A1(n8834), .A2(n6760), .ZN(n10249) );
  NAND2_X1 U9179 ( .A1(n11710), .A2(n10299), .ZN(n6760) );
  NAND2_X1 U9180 ( .A1(n10247), .A2(n6760), .ZN(n10183) );
  OAI211_X1 U9181 ( .C1(n6767), .C2(n6764), .A(n6761), .B(n10740), .ZN(n13942)
         );
  NAND2_X1 U9182 ( .A1(n10648), .A2(n6762), .ZN(n6761) );
  NAND2_X1 U9183 ( .A1(n6763), .A2(n6767), .ZN(n6766) );
  NAND2_X1 U9184 ( .A1(n10648), .A2(n10647), .ZN(n6763) );
  INV_X1 U9185 ( .A(n6635), .ZN(n6764) );
  XNOR2_X1 U9186 ( .A(n6766), .B(n6643), .ZN(n10653) );
  NAND3_X1 U9187 ( .A1(n13922), .A2(n13923), .A3(n10338), .ZN(n6769) );
  NAND2_X1 U9188 ( .A1(n13856), .A2(n9370), .ZN(n13922) );
  NAND2_X1 U9189 ( .A1(n6775), .A2(n6773), .ZN(n9389) );
  NAND2_X1 U9190 ( .A1(n9302), .A2(n9294), .ZN(n9339) );
  NAND2_X1 U9191 ( .A1(n14462), .A2(n6778), .ZN(n6777) );
  NAND2_X1 U9192 ( .A1(n6782), .A2(n6617), .ZN(n7106) );
  NAND3_X1 U9193 ( .A1(n7348), .A2(n14448), .A3(n6542), .ZN(n6785) );
  NAND2_X1 U9194 ( .A1(n7665), .A2(n6511), .ZN(n6792) );
  NAND2_X1 U9195 ( .A1(n7482), .A2(n6802), .ZN(n6798) );
  NAND2_X1 U9196 ( .A1(n6798), .A2(n6799), .ZN(n7512) );
  INV_X1 U9197 ( .A(n8936), .ZN(n8935) );
  NAND2_X1 U9198 ( .A1(n6815), .A2(n8936), .ZN(n6814) );
  INV_X1 U9199 ( .A(n8934), .ZN(n6815) );
  INV_X1 U9200 ( .A(n6818), .ZN(n8904) );
  INV_X1 U9201 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n6819) );
  NAND2_X1 U9202 ( .A1(n6820), .A2(n14558), .ZN(n6822) );
  NAND2_X1 U9203 ( .A1(n14340), .A2(n7087), .ZN(n14301) );
  INV_X1 U9204 ( .A(n14550), .ZN(n6827) );
  NAND2_X1 U9205 ( .A1(n14550), .A2(n6835), .ZN(n6829) );
  NAND3_X1 U9206 ( .A1(n6827), .A2(n6828), .A3(n6836), .ZN(n6831) );
  NAND3_X1 U9207 ( .A1(n6832), .A2(n6830), .A3(n6829), .ZN(n14561) );
  NAND3_X1 U9208 ( .A1(n6835), .A2(n14893), .A3(n8979), .ZN(n6830) );
  AND2_X2 U9209 ( .A1(n12561), .A2(n7436), .ZN(n12556) );
  AND3_X1 U9210 ( .A1(n7411), .A2(n7414), .A3(n6597), .ZN(n10204) );
  NAND2_X1 U9211 ( .A1(n10726), .A2(n6539), .ZN(n6838) );
  OAI211_X1 U9212 ( .C1(n12570), .C2(n6839), .A(n12701), .B(n6838), .ZN(n7487)
         );
  NAND2_X1 U9213 ( .A1(n10726), .A2(n12563), .ZN(n6840) );
  NAND3_X1 U9214 ( .A1(n7477), .A2(n7377), .A3(n7376), .ZN(n7667) );
  AND2_X2 U9215 ( .A1(n7344), .A2(n6842), .ZN(n7384) );
  AND2_X2 U9216 ( .A1(n7372), .A2(n10087), .ZN(n7477) );
  NAND2_X2 U9217 ( .A1(n13147), .A2(n12650), .ZN(n12960) );
  NAND2_X2 U9218 ( .A1(n7732), .A2(n6974), .ZN(n13147) );
  NAND2_X2 U9219 ( .A1(n13158), .A2(n12637), .ZN(n7732) );
  NAND2_X2 U9220 ( .A1(n6843), .A2(n13000), .ZN(n13158) );
  NAND2_X1 U9221 ( .A1(n6844), .A2(n6594), .ZN(n13110) );
  NAND2_X1 U9222 ( .A1(n12887), .A2(n15120), .ZN(n6849) );
  NAND2_X1 U9223 ( .A1(n6847), .A2(n6846), .ZN(n6845) );
  AND2_X1 U9224 ( .A1(n6846), .A2(n6852), .ZN(n8896) );
  NAND2_X1 U9225 ( .A1(n6845), .A2(n6851), .ZN(n8897) );
  OR2_X1 U9226 ( .A1(n15177), .A2(P3_REG0_REG_27__SCAN_IN), .ZN(n6851) );
  OAI21_X2 U9227 ( .B1(n12892), .B2(n6966), .A(n6963), .ZN(n8884) );
  NAND2_X2 U9228 ( .A1(n6853), .A2(n12672), .ZN(n12892) );
  OAI21_X2 U9229 ( .B1(n12929), .B2(n6977), .A(n6577), .ZN(n6853) );
  XNOR2_X2 U9230 ( .A(n7388), .B(n6854), .ZN(n11667) );
  NAND2_X1 U9231 ( .A1(n9372), .A2(n9280), .ZN(n9313) );
  INV_X1 U9232 ( .A(n6865), .ZN(n9600) );
  INV_X1 U9233 ( .A(n6863), .ZN(n9852) );
  INV_X1 U9234 ( .A(n9851), .ZN(n6862) );
  OAI211_X1 U9235 ( .C1(P3_IR_REG_1__SCAN_IN), .C2(P3_IR_REG_0__SCAN_IN), .A(
        P3_IR_REG_2__SCAN_IN), .B(P3_IR_REG_31__SCAN_IN), .ZN(n6879) );
  NAND3_X1 U9236 ( .A1(n6879), .A2(n6877), .A3(n6875), .ZN(n10088) );
  NAND3_X1 U9237 ( .A1(n6878), .A2(n6686), .A3(n6876), .ZN(n6875) );
  OR2_X1 U9238 ( .A1(P3_IR_REG_2__SCAN_IN), .A2(P3_IR_REG_31__SCAN_IN), .ZN(
        n6877) );
  NAND3_X1 U9239 ( .A1(n6507), .A2(n7230), .A3(n6599), .ZN(n14275) );
  NAND2_X1 U9240 ( .A1(n6891), .A2(n6595), .ZN(n6933) );
  NAND2_X1 U9241 ( .A1(n6891), .A2(n6892), .ZN(n8348) );
  NAND2_X1 U9242 ( .A1(n14112), .A2(n11552), .ZN(n14098) );
  NAND2_X2 U9243 ( .A1(n7292), .A2(n7291), .ZN(n14130) );
  NAND2_X1 U9244 ( .A1(n11693), .A2(n6901), .ZN(n6902) );
  INV_X1 U9245 ( .A(n6902), .ZN(n14063) );
  AOI21_X1 U9246 ( .B1(n11691), .B2(n11613), .A(n14493), .ZN(n6903) );
  INV_X2 U9247 ( .A(n14176), .ZN(n6906) );
  NAND2_X1 U9248 ( .A1(n6564), .A2(n6908), .ZN(n6907) );
  INV_X1 U9249 ( .A(n9436), .ZN(n6908) );
  NAND2_X1 U9250 ( .A1(n8152), .A2(n8151), .ZN(n6916) );
  OAI21_X1 U9251 ( .B1(n8760), .B2(n8759), .A(n6633), .ZN(n8742) );
  NAND2_X1 U9252 ( .A1(n8461), .A2(n6929), .ZN(n6928) );
  OAI21_X2 U9253 ( .B1(n8410), .B2(n8409), .A(n6933), .ZN(n8390) );
  OAI21_X1 U9254 ( .B1(n8659), .B2(n8658), .A(n8665), .ZN(n8685) );
  AOI21_X1 U9255 ( .B1(n8658), .B2(n8665), .A(n6645), .ZN(n6937) );
  NAND2_X2 U9256 ( .A1(n8278), .A2(n8277), .ZN(n8325) );
  OR2_X2 U9257 ( .A1(n8000), .A2(n13808), .ZN(n7998) );
  AND2_X1 U9258 ( .A1(n13509), .A2(n6946), .ZN(n13496) );
  NAND2_X1 U9259 ( .A1(n13509), .A2(n12129), .ZN(n13497) );
  NAND3_X1 U9260 ( .A1(n6941), .A2(n6942), .A3(n6943), .ZN(n13695) );
  NAND4_X1 U9261 ( .A1(n6942), .A2(n6941), .A3(n6943), .A4(n14988), .ZN(n6949)
         );
  NAND2_X1 U9262 ( .A1(n13509), .A2(n6600), .ZN(n6941) );
  OR2_X1 U9263 ( .A1(n13509), .A2(n6945), .ZN(n6942) );
  AND2_X2 U9264 ( .A1(n11505), .A2(n14970), .ZN(n11507) );
  AND2_X2 U9265 ( .A1(n10382), .A2(n14962), .ZN(n11505) );
  AND2_X2 U9266 ( .A1(n10864), .A2(n11124), .ZN(n11130) );
  NOR2_X2 U9267 ( .A1(n13662), .A2(n13752), .ZN(n13631) );
  NOR2_X2 U9268 ( .A1(n13601), .A2(n13735), .ZN(n6958) );
  NAND2_X1 U9269 ( .A1(n6960), .A2(n6961), .ZN(n8863) );
  NAND2_X1 U9270 ( .A1(n12892), .A2(n6963), .ZN(n6960) );
  NAND2_X1 U9271 ( .A1(n12892), .A2(n12540), .ZN(n6962) );
  OAI21_X2 U9272 ( .B1(n13071), .B2(n6980), .A(n12618), .ZN(n13059) );
  NAND2_X1 U9273 ( .A1(n7344), .A2(n6981), .ZN(n7395) );
  NOR2_X2 U9274 ( .A1(n7667), .A2(P3_IR_REG_16__SCAN_IN), .ZN(n7687) );
  NAND2_X2 U9275 ( .A1(n6471), .A2(n11519), .ZN(n7448) );
  XNOR2_X2 U9276 ( .A(n7397), .B(n7396), .ZN(n7916) );
  NAND2_X1 U9277 ( .A1(n12158), .A2(n6986), .ZN(n13257) );
  NAND2_X2 U9278 ( .A1(n12101), .A2(n12100), .ZN(n12158) );
  NAND2_X1 U9279 ( .A1(n11092), .A2(n6591), .ZN(n6999) );
  NAND2_X1 U9280 ( .A1(n6999), .A2(n7000), .ZN(n11324) );
  OR2_X1 U9281 ( .A1(n11093), .A2(n11094), .ZN(n7005) );
  NOR3_X1 U9282 ( .A1(n8009), .A2(P2_IR_REG_20__SCAN_IN), .A3(n8010), .ZN(
        n8015) );
  NAND2_X1 U9283 ( .A1(n10351), .A2(n11707), .ZN(n11718) );
  AOI21_X1 U9284 ( .B1(n9938), .B2(n9933), .A(n9939), .ZN(n10039) );
  NAND2_X1 U9285 ( .A1(n13269), .A2(n13268), .ZN(n13267) );
  NAND2_X1 U9286 ( .A1(n8540), .A2(n8539), .ZN(n8545) );
  NAND2_X1 U9287 ( .A1(n8064), .A2(n7354), .ZN(n8105) );
  NAND2_X1 U9288 ( .A1(n12482), .A2(n7010), .ZN(n7009) );
  OAI211_X1 U9289 ( .C1(n12482), .C2(n7012), .A(n12502), .B(n7009), .ZN(n9271)
         );
  NAND2_X1 U9290 ( .A1(n12482), .A2(n12483), .ZN(n12481) );
  OAI21_X1 U9291 ( .B1(n12482), .B2(n9244), .A(n7016), .ZN(n11684) );
  OAI21_X1 U9292 ( .B1(n12492), .B2(n7020), .A(n6510), .ZN(n12469) );
  NAND3_X1 U9293 ( .A1(n7022), .A2(n7024), .A3(n7021), .ZN(n7019) );
  NAND2_X1 U9294 ( .A1(n12348), .A2(n7034), .ZN(n7033) );
  NAND2_X1 U9295 ( .A1(n10754), .A2(n10753), .ZN(n7038) );
  XNOR2_X1 U9296 ( .A(n9233), .B(n7039), .ZN(n12337) );
  NAND2_X1 U9297 ( .A1(n12337), .A2(n12450), .ZN(n12336) );
  AOI21_X2 U9298 ( .B1(n12336), .B2(n6490), .A(n12412), .ZN(n12384) );
  NAND2_X1 U9299 ( .A1(n11040), .A2(n6509), .ZN(n12344) );
  NAND2_X1 U9300 ( .A1(n10360), .A2(n6603), .ZN(n10657) );
  NAND2_X1 U9301 ( .A1(n7567), .A2(n7050), .ZN(n7047) );
  NAND2_X1 U9302 ( .A1(n7047), .A2(n7048), .ZN(n7599) );
  NAND2_X1 U9303 ( .A1(n7748), .A2(n7061), .ZN(n7060) );
  NAND2_X1 U9304 ( .A1(n7748), .A2(n7747), .ZN(n7759) );
  OAI21_X1 U9305 ( .B1(n7748), .B2(n7063), .A(n7061), .ZN(n7784) );
  AOI21_X1 U9306 ( .B1(n7061), .B2(n7063), .A(n7059), .ZN(n7058) );
  OAI21_X2 U9307 ( .B1(n7824), .B2(n7823), .A(n7825), .ZN(n7837) );
  NAND3_X1 U9308 ( .A1(n7068), .A2(n12690), .A3(n12691), .ZN(n7067) );
  INV_X1 U9309 ( .A(n14302), .ZN(n7085) );
  NAND2_X1 U9310 ( .A1(n7087), .A2(n7082), .ZN(n7086) );
  NAND2_X1 U9311 ( .A1(n7083), .A2(n7086), .ZN(n7084) );
  XNOR2_X1 U9312 ( .A(n7084), .B(P2_ADDR_REG_18__SCAN_IN), .ZN(SUB_1596_U62)
         );
  OR2_X1 U9313 ( .A1(n14547), .A2(P2_ADDR_REG_13__SCAN_IN), .ZN(n7088) );
  NAND2_X1 U9314 ( .A1(n14547), .A2(P2_ADDR_REG_13__SCAN_IN), .ZN(n7089) );
  NAND2_X1 U9315 ( .A1(n7102), .A2(n7103), .ZN(n12307) );
  NAND2_X1 U9316 ( .A1(n13952), .A2(n7104), .ZN(n7102) );
  INV_X2 U9317 ( .A(n12276), .ZN(n12301) );
  OR2_X4 U9318 ( .A1(n9342), .A2(n7114), .ZN(n12276) );
  AND2_X1 U9319 ( .A1(n9287), .A2(n9302), .ZN(n9303) );
  NAND3_X1 U9320 ( .A1(n9287), .A2(n7121), .A3(n6668), .ZN(n7120) );
  NAND3_X1 U9321 ( .A1(n9287), .A2(n6668), .A3(n9288), .ZN(n9291) );
  INV_X1 U9322 ( .A(n9303), .ZN(n9334) );
  NAND3_X1 U9323 ( .A1(n8820), .A2(n8822), .A3(n8037), .ZN(n8038) );
  INV_X1 U9324 ( .A(n8835), .ZN(n9834) );
  NAND4_X1 U9325 ( .A1(n8028), .A2(n8030), .A3(n8027), .A4(n8029), .ZN(n8836)
         );
  INV_X1 U9326 ( .A(n11301), .ZN(n7125) );
  INV_X1 U9327 ( .A(n12134), .ZN(n7147) );
  OAI21_X1 U9328 ( .B1(n10184), .B2(n7157), .A(n10371), .ZN(n7153) );
  NAND2_X1 U9329 ( .A1(n10247), .A2(n7156), .ZN(n7155) );
  INV_X1 U9330 ( .A(n7153), .ZN(n7154) );
  NAND2_X1 U9331 ( .A1(n7155), .A2(n7154), .ZN(n10376) );
  NAND2_X1 U9332 ( .A1(n7161), .A2(n6494), .ZN(n7159) );
  INV_X1 U9333 ( .A(n7163), .ZN(n13623) );
  INV_X1 U9334 ( .A(n10861), .ZN(n7174) );
  NAND2_X1 U9335 ( .A1(n10861), .A2(n7169), .ZN(n7166) );
  NAND2_X1 U9336 ( .A1(n7179), .A2(n12827), .ZN(n12819) );
  NAND2_X1 U9337 ( .A1(n12817), .A2(n12818), .ZN(n7181) );
  OAI211_X1 U9338 ( .C1(n12817), .C2(n6644), .A(n7181), .B(n7180), .ZN(n14351)
         );
  OAI211_X1 U9339 ( .C1(n14406), .C2(n6646), .A(n7185), .B(n6502), .ZN(
        P3_U3201) );
  NAND3_X1 U9340 ( .A1(n14406), .A2(n6652), .A3(n14404), .ZN(n7185) );
  NOR2_X1 U9341 ( .A1(n14406), .A2(n14405), .ZN(n14407) );
  NOR2_X2 U9342 ( .A1(n10152), .A2(n7205), .ZN(n10261) );
  NOR2_X2 U9343 ( .A1(n12787), .A2(n12786), .ZN(n12788) );
  NOR2_X2 U9344 ( .A1(n12767), .A2(n7211), .ZN(n12785) );
  OAI211_X1 U9345 ( .C1(n8073), .C2(n6529), .A(n8047), .B(n8048), .ZN(n7213)
         );
  NAND2_X1 U9346 ( .A1(n8584), .A2(n8585), .ZN(n8583) );
  NAND3_X1 U9347 ( .A1(n8308), .A2(n8307), .A3(n6614), .ZN(n7216) );
  INV_X1 U9348 ( .A(n8172), .ZN(n7219) );
  INV_X1 U9349 ( .A(n8173), .ZN(n7220) );
  NAND2_X1 U9350 ( .A1(n8811), .A2(n6620), .ZN(n13809) );
  NAND2_X1 U9351 ( .A1(n7224), .A2(n7223), .ZN(n7222) );
  INV_X1 U9352 ( .A(n8228), .ZN(n7223) );
  NOR2_X1 U9353 ( .A1(n8227), .A2(n7226), .ZN(n7224) );
  NAND3_X1 U9354 ( .A1(n8589), .A2(n8588), .A3(n6572), .ZN(n7227) );
  NAND2_X2 U9355 ( .A1(n9428), .A2(n9506), .ZN(n11521) );
  NAND2_X1 U9356 ( .A1(n11997), .A2(n10403), .ZN(n7235) );
  NAND2_X1 U9357 ( .A1(n7235), .A2(n7232), .ZN(n9901) );
  XNOR2_X1 U9358 ( .A(n7236), .B(n11788), .ZN(n10677) );
  NAND2_X1 U9359 ( .A1(n7242), .A2(n7243), .ZN(n14164) );
  INV_X1 U9360 ( .A(n14141), .ZN(n7250) );
  NAND2_X1 U9361 ( .A1(n14686), .A2(n10497), .ZN(n7251) );
  NAND2_X1 U9362 ( .A1(n7251), .A2(n7252), .ZN(n10561) );
  OAI21_X1 U9363 ( .B1(n10566), .B2(n7258), .A(n7257), .ZN(n14470) );
  NAND2_X1 U9364 ( .A1(n7257), .A2(n7258), .ZN(n7255) );
  NAND2_X1 U9365 ( .A1(n10566), .A2(n7257), .ZN(n7256) );
  NAND2_X1 U9366 ( .A1(n11608), .A2(n7264), .ZN(n7262) );
  OAI21_X1 U9367 ( .B1(n11999), .B2(n9756), .A(n7269), .ZN(n10675) );
  INV_X1 U9368 ( .A(n11997), .ZN(n10404) );
  AND2_X1 U9369 ( .A1(n11493), .A2(n11492), .ZN(n7275) );
  NAND2_X1 U9370 ( .A1(n10427), .A2(n10426), .ZN(n14698) );
  NAND2_X1 U9371 ( .A1(n7279), .A2(n7277), .ZN(n10447) );
  INV_X1 U9372 ( .A(n7278), .ZN(n7277) );
  OAI21_X1 U9373 ( .B1(n7282), .B2(n14700), .A(n10509), .ZN(n7278) );
  NAND2_X1 U9374 ( .A1(n7280), .A2(n10427), .ZN(n7279) );
  AND2_X1 U9375 ( .A1(n10426), .A2(n10432), .ZN(n7280) );
  NAND2_X1 U9376 ( .A1(n7301), .A2(n7300), .ZN(n11789) );
  NAND3_X1 U9377 ( .A1(n6584), .A2(n11784), .A3(n11785), .ZN(n7301) );
  NAND2_X1 U9378 ( .A1(n7304), .A2(n7307), .ZN(n11932) );
  NAND3_X1 U9379 ( .A1(n11926), .A2(n11925), .A3(n7305), .ZN(n7304) );
  NAND3_X1 U9380 ( .A1(n11813), .A2(n11812), .A3(n7308), .ZN(n7310) );
  INV_X1 U9381 ( .A(n11814), .ZN(n7309) );
  NAND2_X1 U9382 ( .A1(n7310), .A2(n7311), .ZN(n11820) );
  NAND3_X1 U9383 ( .A1(n11857), .A2(n11856), .A3(n7315), .ZN(n7313) );
  NAND2_X1 U9384 ( .A1(n7313), .A2(n7312), .ZN(n11876) );
  NAND2_X1 U9385 ( .A1(n7320), .A2(n7321), .ZN(n11942) );
  NAND3_X1 U9386 ( .A1(n11937), .A2(n6611), .A3(n11936), .ZN(n7320) );
  NAND2_X2 U9387 ( .A1(n12557), .A2(n12559), .ZN(n12703) );
  NAND2_X1 U9388 ( .A1(n15110), .A2(n10416), .ZN(n12559) );
  INV_X1 U9389 ( .A(n15110), .ZN(n12764) );
  NAND2_X1 U9390 ( .A1(n7384), .A2(n7323), .ZN(n7392) );
  NOR2_X2 U9391 ( .A1(n7392), .A2(P3_IR_REG_28__SCAN_IN), .ZN(n7386) );
  NAND2_X1 U9392 ( .A1(n7326), .A2(n7324), .ZN(n8888) );
  NAND3_X1 U9393 ( .A1(n6543), .A2(n7901), .A3(n7328), .ZN(n12917) );
  NAND2_X1 U9394 ( .A1(n10879), .A2(n7873), .ZN(n10877) );
  NAND2_X1 U9395 ( .A1(n6575), .A2(n7871), .ZN(n10879) );
  INV_X1 U9396 ( .A(n13037), .ZN(n7343) );
  NAND2_X1 U9397 ( .A1(n7337), .A2(n7338), .ZN(n13014) );
  NAND2_X1 U9398 ( .A1(n13037), .A2(n7340), .ZN(n7337) );
  AND2_X2 U9399 ( .A1(n7345), .A2(n7382), .ZN(n7344) );
  AND2_X1 U9400 ( .A1(n13838), .A2(n13837), .ZN(n13892) );
  INV_X1 U9401 ( .A(n7953), .ZN(n7956) );
  MUX2_X2 U9402 ( .A(n7969), .B(P3_REG0_REG_28__SCAN_IN), .S(n15175), .Z(n7953) );
  NAND2_X1 U9403 ( .A1(n15125), .A2(n15110), .ZN(n15113) );
  INV_X1 U9404 ( .A(n8121), .ZN(n8124) );
  AND2_X1 U9405 ( .A1(n8204), .A2(n8203), .ZN(n8206) );
  INV_X1 U9406 ( .A(n11662), .ZN(n7991) );
  NAND4_X2 U9407 ( .A1(n9381), .A2(n9380), .A3(n9379), .A4(n9378), .ZN(n13995)
         );
  CLKBUF_X1 U9408 ( .A(n13110), .Z(n13175) );
  NAND2_X1 U9409 ( .A1(n6474), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n9348) );
  OAI21_X1 U9410 ( .B1(n8859), .B2(n9817), .A(n7366), .ZN(n8860) );
  AOI22_X2 U9411 ( .A1(n8180), .A2(P1_DATAO_REG_3__SCAN_IN), .B1(n9640), .B2(
        n9728), .ZN(n8088) );
  NOR2_X1 U9412 ( .A1(n12532), .A2(n12531), .ZN(n12533) );
  AND2_X1 U9413 ( .A1(n8202), .A2(n8201), .ZN(n7346) );
  INV_X1 U9414 ( .A(n13275), .ZN(n13276) );
  OR2_X1 U9415 ( .A1(n12885), .A2(n13179), .ZN(n7347) );
  NAND2_X2 U9416 ( .A1(n10030), .A2(n15108), .ZN(n13106) );
  INV_X1 U9417 ( .A(n13179), .ZN(n8900) );
  AND2_X1 U9418 ( .A1(n14447), .A2(n14450), .ZN(n7348) );
  AND2_X1 U9419 ( .A1(n12721), .A2(n12530), .ZN(n7349) );
  AND2_X1 U9420 ( .A1(n12215), .A2(n12214), .ZN(n7350) );
  AND2_X1 U9421 ( .A1(n10088), .A2(P3_REG2_REG_2__SCAN_IN), .ZN(n7351) );
  NAND2_X1 U9422 ( .A1(n6973), .A2(n7431), .ZN(n7352) );
  NOR2_X1 U9423 ( .A1(n8329), .A2(n8328), .ZN(n7353) );
  OR2_X1 U9424 ( .A1(n8063), .A2(n9442), .ZN(n7354) );
  AND2_X1 U9425 ( .A1(n11337), .A2(n11336), .ZN(n7355) );
  OR2_X1 U9426 ( .A1(n12885), .A2(n13234), .ZN(n7356) );
  INV_X1 U9427 ( .A(n14296), .ZN(n11270) );
  INV_X1 U9428 ( .A(n11270), .ZN(n12152) );
  INV_X1 U9429 ( .A(n14379), .ZN(n12848) );
  INV_X1 U9430 ( .A(P3_REG3_REG_9__SCAN_IN), .ZN(n7540) );
  AND2_X2 U9431 ( .A1(n7952), .A2(n12736), .ZN(n15177) );
  INV_X1 U9432 ( .A(n15109), .ZN(n13098) );
  NAND2_X1 U9433 ( .A1(n11327), .A2(n11326), .ZN(n11736) );
  NAND2_X1 U9434 ( .A1(n15177), .A2(n15152), .ZN(n13234) );
  OR2_X1 U9435 ( .A1(n7450), .A2(n15035), .ZN(n7359) );
  INV_X1 U9436 ( .A(n10871), .ZN(n9817) );
  XNOR2_X1 U9437 ( .A(n7394), .B(n7393), .ZN(n7915) );
  NOR2_X1 U9438 ( .A1(n12545), .A2(n12752), .ZN(n7360) );
  AND2_X1 U9439 ( .A1(n9224), .A2(n12753), .ZN(n7361) );
  INV_X4 U9440 ( .A(n11519), .ZN(n9434) );
  AND2_X1 U9441 ( .A1(n13740), .A2(n13625), .ZN(n7362) );
  INV_X1 U9442 ( .A(n14706), .ZN(n14179) );
  AND2_X2 U9443 ( .A1(n11622), .A2(n14188), .ZN(n14706) );
  OR2_X1 U9444 ( .A1(n11297), .A2(n11296), .ZN(n7363) );
  AND2_X1 U9445 ( .A1(n10038), .A2(n10037), .ZN(n7364) );
  INV_X1 U9446 ( .A(n14088), .ZN(n14108) );
  NOR2_X1 U9447 ( .A1(n14119), .A2(n14233), .ZN(n14088) );
  AND2_X1 U9448 ( .A1(n11107), .A2(n11106), .ZN(n7365) );
  AND2_X2 U9449 ( .A1(n9984), .A2(n9914), .ZN(n15019) );
  INV_X1 U9450 ( .A(n14953), .ZN(n15002) );
  AND4_X1 U9451 ( .A1(n8858), .A2(n13490), .A3(n8857), .A4(n10976), .ZN(n7366)
         );
  NAND2_X1 U9452 ( .A1(n10138), .A2(n13607), .ZN(n13606) );
  INV_X1 U9453 ( .A(n13645), .ZN(n13594) );
  INV_X1 U9454 ( .A(n11224), .ZN(n11111) );
  NAND2_X1 U9455 ( .A1(n10216), .A2(n8023), .ZN(n8024) );
  AND2_X1 U9456 ( .A1(n8531), .A2(n10012), .ZN(n8040) );
  INV_X1 U9457 ( .A(n8122), .ZN(n8123) );
  INV_X1 U9458 ( .A(n8269), .ZN(n8270) );
  INV_X1 U9459 ( .A(n8532), .ZN(n8533) );
  OR2_X1 U9460 ( .A1(n13993), .A2(n10484), .ZN(n10485) );
  INV_X1 U9461 ( .A(n12721), .ZN(n12691) );
  INV_X1 U9462 ( .A(n13000), .ZN(n7893) );
  INV_X1 U9463 ( .A(P3_IR_REG_4__SCAN_IN), .ZN(n7476) );
  INV_X1 U9464 ( .A(n9724), .ZN(n8037) );
  INV_X1 U9465 ( .A(n8610), .ZN(n8611) );
  INV_X1 U9466 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n9280) );
  INV_X1 U9467 ( .A(n14344), .ZN(n12818) );
  INV_X1 U9468 ( .A(n12701), .ZN(n7872) );
  NOR2_X1 U9469 ( .A1(P3_IR_REG_2__SCAN_IN), .A2(P3_IR_REG_3__SCAN_IN), .ZN(
        n7372) );
  INV_X1 U9470 ( .A(n8551), .ZN(n8549) );
  INV_X1 U9471 ( .A(n8491), .ZN(n8489) );
  INV_X1 U9472 ( .A(n8240), .ZN(n8238) );
  NAND2_X1 U9473 ( .A1(n10337), .A2(n10336), .ZN(n10338) );
  INV_X1 U9474 ( .A(n11858), .ZN(n11006) );
  NOR2_X1 U9475 ( .A1(P1_ADDR_REG_7__SCAN_IN), .A2(n8955), .ZN(n8909) );
  INV_X1 U9476 ( .A(P3_REG3_REG_17__SCAN_IN), .ZN(n9125) );
  INV_X1 U9477 ( .A(P3_REG3_REG_13__SCAN_IN), .ZN(n7620) );
  OR2_X1 U9478 ( .A1(n7829), .A2(P3_REG3_REG_27__SCAN_IN), .ZN(n7843) );
  NAND2_X1 U9479 ( .A1(n7640), .A2(n12622), .ZN(n7641) );
  INV_X1 U9480 ( .A(n15140), .ZN(n10661) );
  OR2_X1 U9481 ( .A1(n14413), .A2(n13063), .ZN(n12621) );
  NAND2_X1 U9482 ( .A1(n12739), .A2(n12547), .ZN(n12671) );
  AND2_X1 U9483 ( .A1(n7451), .A2(n7359), .ZN(n7452) );
  AND2_X1 U9484 ( .A1(n10023), .A2(n10024), .ZN(n7958) );
  OR2_X1 U9485 ( .A1(n7857), .A2(P3_IR_REG_21__SCAN_IN), .ZN(n7947) );
  AND2_X1 U9486 ( .A1(n7596), .A2(n7583), .ZN(n7594) );
  NOR2_X1 U9487 ( .A1(n7509), .A2(P3_IR_REG_6__SCAN_IN), .ZN(n7530) );
  AND2_X1 U9488 ( .A1(n10848), .A2(n10838), .ZN(n10839) );
  AND2_X1 U9489 ( .A1(n8690), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n8745) );
  NAND2_X1 U9490 ( .A1(n8642), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n8672) );
  NAND2_X1 U9491 ( .A1(n8549), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n8570) );
  NAND2_X1 U9492 ( .A1(n8365), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n8468) );
  OR2_X1 U9493 ( .A1(n8259), .A2(n8258), .ZN(n8291) );
  NAND2_X1 U9494 ( .A1(n8569), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n8598) );
  OR2_X1 U9495 ( .A1(n8313), .A2(n8312), .ZN(n8338) );
  NAND2_X1 U9496 ( .A1(n8238), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n8259) );
  INV_X1 U9497 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n7997) );
  INV_X1 U9498 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n10962) );
  AND2_X1 U9499 ( .A1(n11522), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n11536) );
  OR2_X1 U9500 ( .A1(n13880), .A2(n13881), .ZN(n12206) );
  INV_X1 U9501 ( .A(n10452), .ZN(n10999) );
  NAND2_X1 U9502 ( .A1(n11692), .A2(n13975), .ZN(n11612) );
  INV_X1 U9503 ( .A(n12029), .ZN(n11593) );
  INV_X1 U9504 ( .A(n12019), .ZN(n11493) );
  INV_X1 U9505 ( .A(n11998), .ZN(n9657) );
  INV_X1 U9506 ( .A(n11007), .ZN(n11049) );
  NOR2_X1 U9507 ( .A1(n14673), .A2(n14672), .ZN(n14676) );
  OR2_X1 U9508 ( .A1(n14493), .A2(n14149), .ZN(n9668) );
  AND2_X1 U9509 ( .A1(n9304), .A2(n9295), .ZN(n9288) );
  NOR2_X1 U9510 ( .A1(n7503), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n7523) );
  AND2_X1 U9511 ( .A1(n7523), .A2(n10279), .ZN(n7541) );
  NOR2_X1 U9512 ( .A1(n7588), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n7621) );
  NAND2_X1 U9513 ( .A1(n7695), .A2(n9125), .ZN(n7711) );
  NAND2_X1 U9514 ( .A1(n7792), .A2(n7791), .ZN(n7804) );
  NAND2_X1 U9515 ( .A1(n7541), .A2(n7540), .ZN(n7557) );
  NAND2_X1 U9516 ( .A1(n7621), .A2(n7620), .ZN(n7634) );
  NAND2_X1 U9517 ( .A1(n9168), .A2(n9167), .ZN(n9173) );
  INV_X1 U9518 ( .A(n12496), .ZN(n12486) );
  INV_X1 U9519 ( .A(n9262), .ZN(n12735) );
  INV_X1 U9520 ( .A(n12773), .ZN(n12770) );
  AND2_X1 U9521 ( .A1(n12737), .A2(n12826), .ZN(n9783) );
  INV_X1 U9522 ( .A(n12971), .ZN(n12982) );
  INV_X1 U9523 ( .A(n12755), .ZN(n13018) );
  OR2_X1 U9524 ( .A1(n7488), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n7503) );
  INV_X1 U9525 ( .A(n10027), .ZN(n12695) );
  AOI21_X1 U9526 ( .B1(n12745), .B2(n13098), .A(n8877), .ZN(n8878) );
  OR2_X1 U9527 ( .A1(n6481), .A2(n10910), .ZN(n7789) );
  OR3_X1 U9528 ( .A1(n9783), .A2(n6482), .A3(n12671), .ZN(n15109) );
  OR2_X1 U9529 ( .A1(n13238), .A2(n9249), .ZN(n9767) );
  OAI21_X1 U9530 ( .B1(n7947), .B2(P3_IR_REG_22__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n7949) );
  OAI21_X1 U9531 ( .B1(n7735), .B2(P1_DATAO_REG_20__SCAN_IN), .A(n7744), .ZN(
        n7736) );
  AND2_X1 U9532 ( .A1(n7549), .A2(n7534), .ZN(n7535) );
  AND2_X1 U9533 ( .A1(n7497), .A2(n7484), .ZN(n7495) );
  OR2_X1 U9534 ( .A1(n11724), .A2(n11088), .ZN(n11089) );
  OR2_X1 U9535 ( .A1(n11734), .A2(n11733), .ZN(n11735) );
  INV_X1 U9536 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n13364) );
  OR2_X1 U9537 ( .A1(n10048), .A2(n10047), .ZN(n10049) );
  INV_X1 U9538 ( .A(n8826), .ZN(n8854) );
  OR2_X1 U9539 ( .A1(n8050), .A2(n8051), .ZN(n8054) );
  NOR2_X1 U9540 ( .A1(n13611), .A2(n7362), .ZN(n13584) );
  INV_X1 U9541 ( .A(n13380), .ZN(n13598) );
  NAND2_X1 U9542 ( .A1(n10002), .A2(n9916), .ZN(n9946) );
  INV_X1 U9543 ( .A(n12123), .ZN(n12124) );
  INV_X1 U9544 ( .A(n14994), .ZN(n14986) );
  OR2_X1 U9546 ( .A1(n9796), .A2(n13818), .ZN(n9797) );
  OR2_X1 U9547 ( .A1(n8285), .A2(P2_IR_REG_11__SCAN_IN), .ZN(n8332) );
  INV_X1 U9548 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n10827) );
  NAND2_X1 U9549 ( .A1(n10819), .A2(n10821), .ZN(n10822) );
  INV_X1 U9550 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n11172) );
  INV_X1 U9551 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n11419) );
  AND2_X1 U9552 ( .A1(n11378), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n11437) );
  INV_X1 U9553 ( .A(n14120), .ZN(n14168) );
  OR2_X1 U9554 ( .A1(n11975), .A2(n9586), .ZN(n14167) );
  OR2_X1 U9555 ( .A1(n11622), .A2(n12035), .ZN(n11701) );
  INV_X1 U9556 ( .A(n12001), .ZN(n10509) );
  INV_X1 U9557 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n9311) );
  AND2_X1 U9558 ( .A1(n12496), .A2(n13100), .ZN(n12471) );
  INV_X1 U9559 ( .A(n12474), .ZN(n12441) );
  AND4_X1 U9560 ( .A1(n12519), .A2(n12518), .A3(n12517), .A4(n12516), .ZN(
        n12861) );
  AND4_X1 U9561 ( .A1(n7809), .A2(n7808), .A3(n7807), .A4(n7806), .ZN(n12415)
         );
  AND4_X1 U9562 ( .A1(n7580), .A2(n7579), .A3(n7578), .A4(n7577), .ZN(n12464)
         );
  NOR2_X1 U9563 ( .A1(n11141), .A2(n11140), .ZN(n11144) );
  INV_X1 U9564 ( .A(n12853), .ZN(n15097) );
  AND2_X1 U9565 ( .A1(n9784), .A2(n9783), .ZN(n14404) );
  OR2_X1 U9566 ( .A1(n7944), .A2(n12733), .ZN(n13103) );
  INV_X1 U9567 ( .A(n11074), .ZN(n12926) );
  INV_X1 U9568 ( .A(n15108), .ZN(n13092) );
  AND3_X1 U9569 ( .A1(n7961), .A2(n7960), .A3(n7959), .ZN(n10026) );
  INV_X1 U9570 ( .A(n15170), .ZN(n15152) );
  INV_X1 U9571 ( .A(n15171), .ZN(n15161) );
  XNOR2_X1 U9572 ( .A(n7949), .B(n7948), .ZN(n9766) );
  XNOR2_X1 U9573 ( .A(n7852), .B(P3_IR_REG_22__SCAN_IN), .ZN(n12739) );
  AND2_X1 U9574 ( .A1(n7617), .A2(n7649), .ZN(n12802) );
  INV_X1 U9575 ( .A(n11519), .ZN(n9438) );
  INV_X1 U9576 ( .A(n13351), .ZN(n11753) );
  INV_X1 U9577 ( .A(n9819), .ZN(n9823) );
  NAND2_X1 U9578 ( .A1(n8801), .A2(n8800), .ZN(n8859) );
  OR2_X1 U9579 ( .A1(n12106), .A2(n8767), .ZN(n8679) );
  INV_X1 U9580 ( .A(n8746), .ZN(n8771) );
  INV_X1 U9581 ( .A(n14884), .ZN(n14913) );
  INV_X1 U9582 ( .A(n14890), .ZN(n14922) );
  INV_X1 U9583 ( .A(n14880), .ZN(n14918) );
  INV_X1 U9584 ( .A(n13611), .ZN(n13743) );
  INV_X1 U9585 ( .A(n12115), .ZN(n13637) );
  OR2_X1 U9586 ( .A1(n9925), .A2(n9924), .ZN(n13645) );
  INV_X1 U9587 ( .A(n13594), .ZN(n13677) );
  INV_X1 U9588 ( .A(n14931), .ZN(n9914) );
  AND2_X1 U9589 ( .A1(n13654), .A2(n14937), .ZN(n14984) );
  INV_X1 U9590 ( .A(n14984), .ZN(n15000) );
  AND2_X1 U9591 ( .A1(n14933), .A2(n9913), .ZN(n9984) );
  OR2_X1 U9592 ( .A1(n11394), .A2(n9800), .ZN(n9798) );
  XNOR2_X1 U9593 ( .A(n8810), .B(P2_IR_REG_24__SCAN_IN), .ZN(n11394) );
  AND2_X1 U9594 ( .A1(n8286), .A2(n8332), .ZN(n9866) );
  INV_X1 U9595 ( .A(n14466), .ZN(n13934) );
  AND2_X1 U9596 ( .A1(n9419), .A2(n12055), .ZN(n14466) );
  INV_X1 U9597 ( .A(n12312), .ZN(n13969) );
  AND4_X1 U9598 ( .A1(n11600), .A2(n11599), .A3(n11598), .A4(n11597), .ZN(
        n12311) );
  AND2_X1 U9599 ( .A1(n11444), .A2(n11443), .ZN(n14170) );
  AND2_X1 U9600 ( .A1(n11001), .A2(n11000), .ZN(n12188) );
  OR2_X1 U9601 ( .A1(n9587), .A2(n12056), .ZN(n14647) );
  INV_X1 U9602 ( .A(n14647), .ZN(n14633) );
  AND2_X1 U9603 ( .A1(n9579), .A2(n9578), .ZN(n14638) );
  NAND2_X1 U9604 ( .A1(n11688), .A2(n11687), .ZN(n11689) );
  NAND2_X1 U9605 ( .A1(n9411), .A2(n11958), .ZN(n14701) );
  NAND2_X1 U9606 ( .A1(n12057), .A2(n9696), .ZN(n14188) );
  INV_X1 U9607 ( .A(n11701), .ZN(n14713) );
  INV_X1 U9608 ( .A(n14708), .ZN(n14476) );
  INV_X1 U9609 ( .A(n10394), .ZN(n9671) );
  INV_X1 U9610 ( .A(n14777), .ZN(n14753) );
  AND2_X1 U9611 ( .A1(n11636), .A2(n14730), .ZN(n14721) );
  INV_X1 U9612 ( .A(n14721), .ZN(n14783) );
  AND3_X1 U9613 ( .A1(n9703), .A2(n9702), .A3(n9701), .ZN(n10395) );
  AND2_X1 U9614 ( .A1(n9782), .A2(n9781), .ZN(n15094) );
  INV_X1 U9615 ( .A(n9269), .ZN(n9270) );
  INV_X1 U9616 ( .A(n12502), .ZN(n12478) );
  AND4_X1 U9617 ( .A1(n12519), .A2(n8874), .A3(n8873), .A4(n8872), .ZN(n12529)
         );
  INV_X1 U9618 ( .A(n13017), .ZN(n12757) );
  OR2_X2 U9619 ( .A1(n9307), .A2(n13238), .ZN(n12765) );
  INV_X1 U9620 ( .A(P3_ADDR_REG_4__SCAN_IN), .ZN(n15056) );
  INV_X1 U9621 ( .A(n14404), .ZN(n15101) );
  NAND2_X1 U9622 ( .A1(n10031), .A2(n15105), .ZN(n13094) );
  INV_X1 U9623 ( .A(n13106), .ZN(n13116) );
  NAND2_X1 U9624 ( .A1(n13106), .A2(n15123), .ZN(n11074) );
  NAND2_X1 U9625 ( .A1(n15193), .A2(n15152), .ZN(n13179) );
  INV_X1 U9626 ( .A(n15193), .ZN(n15190) );
  INV_X1 U9627 ( .A(n12530), .ZN(n13184) );
  INV_X1 U9628 ( .A(n12382), .ZN(n13197) );
  INV_X1 U9629 ( .A(n15177), .ZN(n15175) );
  INV_X1 U9630 ( .A(SI_26_), .ZN(n11202) );
  INV_X1 U9631 ( .A(SI_20_), .ZN(n10287) );
  INV_X1 U9632 ( .A(SI_16_), .ZN(n9679) );
  INV_X1 U9633 ( .A(n11139), .ZN(n14320) );
  INV_X1 U9634 ( .A(n14317), .ZN(n13250) );
  INV_X1 U9635 ( .A(n14926), .ZN(n14800) );
  INV_X1 U9636 ( .A(n13747), .ZN(n13621) );
  INV_X1 U9637 ( .A(n9820), .ZN(n13371) );
  NAND2_X1 U9638 ( .A1(n8775), .A2(n8774), .ZN(n13375) );
  NAND2_X1 U9639 ( .A1(n8498), .A2(n8497), .ZN(n13641) );
  OR2_X1 U9640 ( .A1(n9644), .A2(n8820), .ZN(n14880) );
  OR2_X1 U9641 ( .A1(n9648), .A2(P2_U3088), .ZN(n14926) );
  AND2_X1 U9642 ( .A1(n10798), .A2(n10797), .ZN(n14991) );
  NAND2_X1 U9643 ( .A1(n13606), .A2(n10147), .ZN(n13649) );
  INV_X1 U9644 ( .A(n15019), .ZN(n15017) );
  NAND2_X1 U9645 ( .A1(n13718), .A2(n13717), .ZN(n13793) );
  AND3_X1 U9646 ( .A1(n14992), .A2(n14991), .A3(n14990), .ZN(n15016) );
  INV_X1 U9647 ( .A(n15002), .ZN(n15004) );
  AND2_X1 U9648 ( .A1(n9984), .A2(n14931), .ZN(n14953) );
  OR2_X1 U9649 ( .A1(n14934), .A2(n14928), .ZN(n14929) );
  INV_X1 U9650 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n9630) );
  INV_X1 U9651 ( .A(n14247), .ZN(n13920) );
  INV_X1 U9652 ( .A(n14463), .ZN(n13972) );
  NAND4_X1 U9653 ( .A1(n11584), .A2(n11583), .A3(n11582), .A4(n11581), .ZN(
        n14069) );
  INV_X1 U9654 ( .A(n14170), .ZN(n13978) );
  OR2_X1 U9655 ( .A1(n9587), .A2(n9586), .ZN(n14642) );
  NAND2_X1 U9656 ( .A1(n9505), .A2(n9503), .ZN(n14661) );
  OR2_X1 U9657 ( .A1(n14706), .A2(n10400), .ZN(n14708) );
  INV_X1 U9658 ( .A(n14179), .ZN(n14681) );
  OR2_X1 U9659 ( .A1(n14706), .A2(n10471), .ZN(n14174) );
  INV_X1 U9660 ( .A(n14799), .ZN(n14797) );
  AND2_X2 U9661 ( .A1(n9672), .A2(n9671), .ZN(n14799) );
  INV_X1 U9662 ( .A(n14787), .ZN(n14785) );
  AND2_X1 U9663 ( .A1(n9500), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9486) );
  OR2_X1 U9664 ( .A1(n10131), .A2(n10308), .ZN(n14036) );
  INV_X1 U9665 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n9564) );
  XNOR2_X1 U9666 ( .A(n8950), .B(n8949), .ZN(n14322) );
  INV_X1 U9667 ( .A(n14560), .ZN(n14559) );
  INV_X1 U9668 ( .A(n12765), .ZN(P3_U3897) );
  NAND2_X1 U9669 ( .A1(n7956), .A2(n7955), .ZN(P3_U3455) );
  AND2_X1 U9670 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9643), .ZN(P2_U3947) );
  INV_X2 U9671 ( .A(n13979), .ZN(P1_U4016) );
  NOR2_X1 U9672 ( .A1(P3_IR_REG_12__SCAN_IN), .A2(P3_IR_REG_11__SCAN_IN), .ZN(
        n7371) );
  INV_X1 U9673 ( .A(P3_IR_REG_5__SCAN_IN), .ZN(n7375) );
  INV_X1 U9674 ( .A(P3_IR_REG_9__SCAN_IN), .ZN(n7374) );
  INV_X1 U9675 ( .A(P3_IR_REG_6__SCAN_IN), .ZN(n7373) );
  NOR2_X1 U9676 ( .A1(P3_IR_REG_22__SCAN_IN), .A2(P3_IR_REG_18__SCAN_IN), .ZN(
        n7380) );
  INV_X2 U9677 ( .A(P3_IR_REG_20__SCAN_IN), .ZN(n7854) );
  NAND2_X1 U9678 ( .A1(n7386), .A2(n6854), .ZN(n13242) );
  INV_X1 U9679 ( .A(n7386), .ZN(n7387) );
  INV_X1 U9680 ( .A(P3_REG3_REG_2__SCAN_IN), .ZN(n7389) );
  OR2_X1 U9681 ( .A1(n7455), .A2(n7389), .ZN(n7414) );
  NAND2_X1 U9682 ( .A1(n7422), .A2(P3_REG1_REG_2__SCAN_IN), .ZN(n7413) );
  NAND2_X1 U9683 ( .A1(n7454), .A2(P3_REG0_REG_2__SCAN_IN), .ZN(n7412) );
  INV_X2 U9684 ( .A(n7468), .ZN(n12514) );
  NAND2_X1 U9685 ( .A1(n7392), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7394) );
  NAND2_X1 U9686 ( .A1(n7395), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7397) );
  NAND3_X1 U9687 ( .A1(n7399), .A2(n7398), .A3(P3_ADDR_REG_19__SCAN_IN), .ZN(
        n7400) );
  NAND2_X1 U9688 ( .A1(n7400), .A2(n14056), .ZN(n7404) );
  NAND3_X1 U9689 ( .A1(n7401), .A2(n14305), .A3(P2_ADDR_REG_19__SCAN_IN), .ZN(
        n7402) );
  NAND2_X1 U9690 ( .A1(n7402), .A2(P1_ADDR_REG_19__SCAN_IN), .ZN(n7403) );
  XNOR2_X1 U9691 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .ZN(n7433) );
  INV_X1 U9692 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n8004) );
  INV_X1 U9693 ( .A(n7432), .ZN(n7405) );
  INV_X1 U9694 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n9437) );
  NAND2_X1 U9695 ( .A1(n9437), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n7406) );
  NAND2_X1 U9696 ( .A1(n9450), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n7442) );
  INV_X1 U9697 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n9461) );
  NAND2_X1 U9698 ( .A1(n9461), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n7407) );
  AND2_X1 U9699 ( .A1(n7442), .A2(n7407), .ZN(n7408) );
  NAND2_X1 U9700 ( .A1(n7409), .A2(n7408), .ZN(n7443) );
  OAI21_X1 U9701 ( .B1(n7409), .B2(n7408), .A(n7443), .ZN(n14313) );
  OR2_X1 U9702 ( .A1(n7462), .A2(SI_2_), .ZN(n7410) );
  NAND4_X1 U9703 ( .A1(n7414), .A2(n7413), .A3(n7412), .A4(n7411), .ZN(n9174)
         );
  NAND2_X1 U9704 ( .A1(n9174), .A2(n15107), .ZN(n12561) );
  NAND2_X1 U9705 ( .A1(n7422), .A2(P3_REG1_REG_0__SCAN_IN), .ZN(n7418) );
  NAND2_X1 U9706 ( .A1(n7454), .A2(P3_REG0_REG_0__SCAN_IN), .ZN(n7417) );
  NAND2_X1 U9707 ( .A1(n7423), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n7416) );
  NAND2_X1 U9708 ( .A1(n7437), .A2(P3_REG3_REG_0__SCAN_IN), .ZN(n7415) );
  INV_X1 U9709 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n9356) );
  NAND2_X1 U9710 ( .A1(n9356), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n7419) );
  AND2_X1 U9711 ( .A1(n7432), .A2(n7419), .ZN(n7420) );
  NAND2_X1 U9712 ( .A1(n8084), .A2(SI_0_), .ZN(n8005) );
  OAI21_X1 U9713 ( .B1(n9434), .B2(n7420), .A(n8005), .ZN(n13251) );
  INV_X1 U9714 ( .A(n13251), .ZN(n7421) );
  MUX2_X1 U9715 ( .A(n6876), .B(n7421), .S(n7450), .Z(n10104) );
  NOR2_X2 U9716 ( .A1(n12766), .A2(n10104), .ZN(n12553) );
  NAND2_X1 U9717 ( .A1(n7454), .A2(P3_REG0_REG_1__SCAN_IN), .ZN(n7427) );
  NAND2_X1 U9718 ( .A1(n7422), .A2(P3_REG1_REG_1__SCAN_IN), .ZN(n7426) );
  NAND2_X1 U9719 ( .A1(n7423), .A2(P3_REG2_REG_1__SCAN_IN), .ZN(n7425) );
  NAND2_X1 U9720 ( .A1(n7437), .A2(P3_REG3_REG_1__SCAN_IN), .ZN(n7424) );
  INV_X1 U9721 ( .A(SI_1_), .ZN(n9442) );
  NAND2_X1 U9722 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(P3_IR_REG_0__SCAN_IN), .ZN(
        n7428) );
  INV_X1 U9723 ( .A(n10087), .ZN(n7429) );
  INV_X1 U9724 ( .A(n9795), .ZN(n7431) );
  XNOR2_X1 U9725 ( .A(n7433), .B(n7432), .ZN(n9441) );
  NAND2_X1 U9726 ( .A1(n12553), .A2(n12557), .ZN(n9171) );
  NAND2_X1 U9727 ( .A1(n9171), .A2(n12559), .ZN(n15104) );
  NAND2_X1 U9728 ( .A1(n12556), .A2(n15104), .ZN(n15103) );
  NAND2_X1 U9729 ( .A1(n15103), .A2(n7436), .ZN(n10724) );
  NAND2_X1 U9730 ( .A1(n12514), .A2(P3_REG2_REG_3__SCAN_IN), .ZN(n7441) );
  NAND2_X1 U9731 ( .A1(n7454), .A2(P3_REG0_REG_3__SCAN_IN), .ZN(n7440) );
  NAND2_X1 U9732 ( .A1(n7422), .A2(P3_REG1_REG_3__SCAN_IN), .ZN(n7439) );
  INV_X1 U9733 ( .A(P3_REG3_REG_3__SCAN_IN), .ZN(n9095) );
  NAND2_X1 U9734 ( .A1(n7437), .A2(n9095), .ZN(n7438) );
  OR2_X1 U9735 ( .A1(n6481), .A2(SI_3_), .ZN(n7453) );
  NAND2_X1 U9736 ( .A1(n7443), .A2(n7442), .ZN(n7446) );
  NAND2_X1 U9737 ( .A1(n9446), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n7463) );
  INV_X1 U9738 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n9467) );
  NAND2_X1 U9739 ( .A1(n9467), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n7444) );
  AND2_X1 U9740 ( .A1(n7463), .A2(n7444), .ZN(n7445) );
  OR2_X1 U9741 ( .A1(n7446), .A2(n7445), .ZN(n7447) );
  NAND2_X1 U9742 ( .A1(n7464), .A2(n7447), .ZN(n14310) );
  OR2_X1 U9743 ( .A1(n7448), .A2(n14310), .ZN(n7451) );
  NAND2_X1 U9744 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(n6538), .ZN(n7449) );
  XNOR2_X1 U9745 ( .A(n7449), .B(P3_IR_REG_3__SCAN_IN), .ZN(n15035) );
  NAND2_X1 U9746 ( .A1(n12763), .A2(n15135), .ZN(n12562) );
  INV_X1 U9747 ( .A(n10727), .ZN(n12705) );
  NAND2_X1 U9748 ( .A1(n10724), .A2(n12705), .ZN(n10726) );
  NAND2_X1 U9749 ( .A1(n7422), .A2(P3_REG1_REG_4__SCAN_IN), .ZN(n7460) );
  NAND2_X1 U9750 ( .A1(n12515), .A2(P3_REG0_REG_4__SCAN_IN), .ZN(n7459) );
  INV_X4 U9751 ( .A(n7455), .ZN(n7911) );
  AND2_X1 U9752 ( .A1(P3_REG3_REG_4__SCAN_IN), .A2(P3_REG3_REG_3__SCAN_IN), 
        .ZN(n7456) );
  NOR2_X1 U9753 ( .A1(P3_REG3_REG_3__SCAN_IN), .A2(P3_REG3_REG_4__SCAN_IN), 
        .ZN(n7469) );
  OR2_X1 U9754 ( .A1(n7456), .A2(n7469), .ZN(n10665) );
  NAND2_X1 U9755 ( .A1(n7911), .A2(n10665), .ZN(n7458) );
  NAND2_X1 U9756 ( .A1(n12514), .A2(P3_REG2_REG_4__SCAN_IN), .ZN(n7457) );
  OR2_X1 U9757 ( .A1(n7477), .A2(n13241), .ZN(n7461) );
  XNOR2_X1 U9758 ( .A(n7461), .B(P3_IR_REG_4__SCAN_IN), .ZN(n10091) );
  OR2_X1 U9759 ( .A1(n6481), .A2(SI_4_), .ZN(n7467) );
  NAND2_X1 U9760 ( .A1(n9452), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n7483) );
  INV_X1 U9761 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n9475) );
  NAND2_X1 U9762 ( .A1(n9475), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n7465) );
  XNOR2_X1 U9763 ( .A(n7482), .B(n7481), .ZN(n9497) );
  OR2_X1 U9764 ( .A1(n7448), .A2(n9497), .ZN(n7466) );
  OAI211_X1 U9765 ( .C1(n10091), .C2(n6472), .A(n7467), .B(n7466), .ZN(n15140)
         );
  NAND2_X1 U9766 ( .A1(n10363), .A2(n10661), .ZN(n12573) );
  NAND2_X1 U9767 ( .A1(n12762), .A2(n15140), .ZN(n12572) );
  NAND2_X1 U9768 ( .A1(n12573), .A2(n12572), .ZN(n12698) );
  INV_X1 U9769 ( .A(n12698), .ZN(n12570) );
  NAND2_X1 U9770 ( .A1(n7423), .A2(P3_REG2_REG_5__SCAN_IN), .ZN(n7475) );
  NAND2_X1 U9771 ( .A1(n7422), .A2(P3_REG1_REG_5__SCAN_IN), .ZN(n7474) );
  NAND2_X1 U9772 ( .A1(n7469), .A2(n9149), .ZN(n7488) );
  OR2_X1 U9773 ( .A1(n7469), .A2(n9149), .ZN(n7470) );
  NAND2_X1 U9774 ( .A1(n7488), .A2(n7470), .ZN(n10759) );
  NAND2_X1 U9775 ( .A1(n7911), .A2(n10759), .ZN(n7473) );
  NAND2_X1 U9776 ( .A1(n12515), .A2(P3_REG0_REG_5__SCAN_IN), .ZN(n7472) );
  NAND4_X1 U9777 ( .A1(n7475), .A2(n7474), .A3(n7473), .A4(n7472), .ZN(n12761)
         );
  NAND2_X1 U9778 ( .A1(n7477), .A2(n7476), .ZN(n7479) );
  NAND2_X1 U9779 ( .A1(n7479), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7478) );
  MUX2_X1 U9780 ( .A(P3_IR_REG_31__SCAN_IN), .B(n7478), .S(
        P3_IR_REG_5__SCAN_IN), .Z(n7480) );
  NAND2_X1 U9781 ( .A1(n7480), .A2(n7509), .ZN(n10093) );
  INV_X1 U9782 ( .A(n10093), .ZN(n15069) );
  OR2_X1 U9783 ( .A1(n6480), .A2(SI_5_), .ZN(n7486) );
  NAND2_X1 U9784 ( .A1(n9448), .A2(P2_DATAO_REG_5__SCAN_IN), .ZN(n7497) );
  NAND2_X1 U9785 ( .A1(n9464), .A2(P1_DATAO_REG_5__SCAN_IN), .ZN(n7484) );
  XNOR2_X1 U9786 ( .A(n7496), .B(n7495), .ZN(n9491) );
  OR2_X1 U9787 ( .A1(n7448), .A2(n9491), .ZN(n7485) );
  OAI211_X1 U9788 ( .C1(n15069), .C2(n7450), .A(n7486), .B(n7485), .ZN(n15146)
         );
  INV_X1 U9789 ( .A(n15146), .ZN(n10755) );
  NAND2_X1 U9790 ( .A1(n10876), .A2(n10755), .ZN(n12576) );
  NAND2_X1 U9791 ( .A1(n12761), .A2(n15146), .ZN(n12577) );
  AND2_X2 U9792 ( .A1(n12576), .A2(n12577), .ZN(n12701) );
  NAND2_X1 U9793 ( .A1(n7487), .A2(n12576), .ZN(n10875) );
  NAND2_X1 U9794 ( .A1(n7423), .A2(P3_REG2_REG_6__SCAN_IN), .ZN(n7493) );
  NAND2_X1 U9795 ( .A1(n7522), .A2(P3_REG1_REG_6__SCAN_IN), .ZN(n7492) );
  NAND2_X1 U9796 ( .A1(n7488), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n7489) );
  NAND2_X1 U9797 ( .A1(n7503), .A2(n7489), .ZN(n10884) );
  NAND2_X1 U9798 ( .A1(n7911), .A2(n10884), .ZN(n7491) );
  NAND2_X1 U9799 ( .A1(n12515), .A2(P3_REG0_REG_6__SCAN_IN), .ZN(n7490) );
  NAND4_X1 U9800 ( .A1(n7493), .A2(n7492), .A3(n7491), .A4(n7490), .ZN(n12760)
         );
  INV_X1 U9801 ( .A(n12760), .ZN(n7501) );
  NAND2_X1 U9802 ( .A1(n7509), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7494) );
  XNOR2_X1 U9803 ( .A(n7494), .B(P3_IR_REG_6__SCAN_IN), .ZN(n10160) );
  INV_X1 U9804 ( .A(SI_6_), .ZN(n9457) );
  OR2_X1 U9805 ( .A1(n6480), .A2(n9457), .ZN(n7500) );
  XNOR2_X1 U9806 ( .A(n9451), .B(P2_DATAO_REG_6__SCAN_IN), .ZN(n7498) );
  XNOR2_X1 U9807 ( .A(n7512), .B(n7498), .ZN(n9458) );
  OR2_X1 U9808 ( .A1(n7448), .A2(n9458), .ZN(n7499) );
  OAI211_X1 U9809 ( .C1(n10155), .C2(n6472), .A(n7500), .B(n7499), .ZN(n15151)
         );
  NAND2_X1 U9810 ( .A1(n7501), .A2(n15151), .ZN(n12584) );
  INV_X1 U9811 ( .A(n15151), .ZN(n7502) );
  NAND2_X1 U9812 ( .A1(n12760), .A2(n7502), .ZN(n12583) );
  NAND2_X1 U9813 ( .A1(n12584), .A2(n12583), .ZN(n12704) );
  INV_X1 U9814 ( .A(n12704), .ZN(n10874) );
  NAND2_X1 U9815 ( .A1(n10875), .A2(n10874), .ZN(n10873) );
  NAND2_X1 U9816 ( .A1(n10873), .A2(n12584), .ZN(n10888) );
  NAND2_X1 U9817 ( .A1(n7423), .A2(P3_REG2_REG_7__SCAN_IN), .ZN(n7508) );
  NAND2_X1 U9818 ( .A1(n7522), .A2(P3_REG1_REG_7__SCAN_IN), .ZN(n7507) );
  AND2_X1 U9819 ( .A1(n7503), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n7504) );
  OR2_X1 U9820 ( .A1(n7504), .A2(n7523), .ZN(n12322) );
  NAND2_X1 U9821 ( .A1(n7911), .A2(n12322), .ZN(n7506) );
  NAND2_X1 U9822 ( .A1(n12515), .A2(P3_REG0_REG_7__SCAN_IN), .ZN(n7505) );
  NAND4_X1 U9823 ( .A1(n7508), .A2(n7507), .A3(n7506), .A4(n7505), .ZN(n12759)
         );
  OR2_X1 U9824 ( .A1(n7530), .A2(n13241), .ZN(n7510) );
  XNOR2_X1 U9825 ( .A(n7510), .B(P3_IR_REG_7__SCAN_IN), .ZN(n10269) );
  OR2_X1 U9826 ( .A1(n6480), .A2(SI_7_), .ZN(n7520) );
  NAND2_X1 U9827 ( .A1(n9472), .A2(P1_DATAO_REG_6__SCAN_IN), .ZN(n7511) );
  NAND2_X1 U9828 ( .A1(n7512), .A2(n7511), .ZN(n7514) );
  NAND2_X1 U9829 ( .A1(n9451), .A2(P2_DATAO_REG_6__SCAN_IN), .ZN(n7513) );
  NAND2_X1 U9830 ( .A1(n7514), .A2(n7513), .ZN(n7517) );
  NAND2_X1 U9831 ( .A1(n9479), .A2(P1_DATAO_REG_7__SCAN_IN), .ZN(n7532) );
  NAND2_X1 U9832 ( .A1(n9482), .A2(P2_DATAO_REG_7__SCAN_IN), .ZN(n7515) );
  NAND2_X1 U9833 ( .A1(n7532), .A2(n7515), .ZN(n7516) );
  NAND2_X1 U9834 ( .A1(n7517), .A2(n7516), .ZN(n7518) );
  AND2_X1 U9835 ( .A1(n7533), .A2(n7518), .ZN(n9495) );
  OR2_X1 U9836 ( .A1(n7448), .A2(n9495), .ZN(n7519) );
  OAI211_X1 U9837 ( .C1(n10269), .C2(n7450), .A(n7520), .B(n7519), .ZN(n15157)
         );
  XNOR2_X1 U9838 ( .A(n12759), .B(n15157), .ZN(n10891) );
  NAND2_X1 U9839 ( .A1(n10888), .A2(n12706), .ZN(n10890) );
  INV_X1 U9840 ( .A(n12759), .ZN(n12587) );
  INV_X1 U9841 ( .A(n15157), .ZN(n12588) );
  NAND2_X1 U9842 ( .A1(n12587), .A2(n12588), .ZN(n7521) );
  NAND2_X1 U9843 ( .A1(n10890), .A2(n7521), .ZN(n11076) );
  INV_X1 U9844 ( .A(n7422), .ZN(n7574) );
  NAND2_X1 U9845 ( .A1(n7522), .A2(P3_REG1_REG_8__SCAN_IN), .ZN(n7528) );
  NAND2_X1 U9846 ( .A1(n7423), .A2(P3_REG2_REG_8__SCAN_IN), .ZN(n7527) );
  NOR2_X1 U9847 ( .A1(n7523), .A2(n10279), .ZN(n7524) );
  OR2_X1 U9848 ( .A1(n7541), .A2(n7524), .ZN(n11039) );
  NAND2_X1 U9849 ( .A1(n7911), .A2(n11039), .ZN(n7526) );
  NAND2_X1 U9850 ( .A1(n12515), .A2(P3_REG0_REG_8__SCAN_IN), .ZN(n7525) );
  NAND4_X1 U9851 ( .A1(n7528), .A2(n7527), .A3(n7526), .A4(n7525), .ZN(n12758)
         );
  INV_X1 U9852 ( .A(n12758), .ZN(n7876) );
  NAND2_X1 U9853 ( .A1(n7530), .A2(n7529), .ZN(n7547) );
  NAND2_X1 U9854 ( .A1(n7547), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7531) );
  XNOR2_X1 U9855 ( .A(n7531), .B(P3_IR_REG_8__SCAN_IN), .ZN(n10699) );
  NAND2_X1 U9856 ( .A1(n9517), .A2(P1_DATAO_REG_8__SCAN_IN), .ZN(n7549) );
  NAND2_X1 U9857 ( .A1(n9512), .A2(P2_DATAO_REG_8__SCAN_IN), .ZN(n7534) );
  NAND2_X1 U9858 ( .A1(n7536), .A2(n7535), .ZN(n7550) );
  OR2_X1 U9859 ( .A1(n7536), .A2(n7535), .ZN(n7537) );
  NAND2_X1 U9860 ( .A1(n7550), .A2(n7537), .ZN(n9439) );
  OR2_X1 U9861 ( .A1(n7448), .A2(n9439), .ZN(n7539) );
  INV_X1 U9862 ( .A(SI_8_), .ZN(n9440) );
  OR2_X1 U9863 ( .A1(n6481), .A2(n9440), .ZN(n7538) );
  OAI211_X1 U9864 ( .C1(n10709), .C2(n6472), .A(n7539), .B(n7538), .ZN(n11045)
         );
  NAND2_X1 U9865 ( .A1(n7876), .A2(n11045), .ZN(n12595) );
  INV_X1 U9866 ( .A(n11045), .ZN(n15163) );
  NAND2_X1 U9867 ( .A1(n12758), .A2(n15163), .ZN(n12594) );
  NAND2_X1 U9868 ( .A1(n12514), .A2(P3_REG2_REG_9__SCAN_IN), .ZN(n7546) );
  NAND2_X1 U9869 ( .A1(n7522), .A2(P3_REG1_REG_9__SCAN_IN), .ZN(n7545) );
  OR2_X1 U9870 ( .A1(n7541), .A2(n7540), .ZN(n7542) );
  NAND2_X1 U9871 ( .A1(n7557), .A2(n7542), .ZN(n12427) );
  NAND2_X1 U9872 ( .A1(n7911), .A2(n12427), .ZN(n7544) );
  NAND2_X1 U9873 ( .A1(n12515), .A2(P3_REG0_REG_9__SCAN_IN), .ZN(n7543) );
  NAND4_X1 U9874 ( .A1(n7546), .A2(n7545), .A3(n7544), .A4(n7543), .ZN(n13099)
         );
  NAND2_X1 U9875 ( .A1(n7569), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7548) );
  XNOR2_X1 U9876 ( .A(n7548), .B(n7374), .ZN(n15089) );
  NAND2_X1 U9877 ( .A1(n7550), .A2(n7549), .ZN(n7553) );
  NAND2_X1 U9878 ( .A1(n9524), .A2(P1_DATAO_REG_9__SCAN_IN), .ZN(n7563) );
  NAND2_X1 U9879 ( .A1(n9518), .A2(P2_DATAO_REG_9__SCAN_IN), .ZN(n7551) );
  NAND2_X1 U9880 ( .A1(n7553), .A2(n7552), .ZN(n7564) );
  OR2_X1 U9881 ( .A1(n7553), .A2(n7552), .ZN(n7554) );
  AND2_X1 U9882 ( .A1(n7564), .A2(n7554), .ZN(n9493) );
  OR2_X1 U9883 ( .A1(n7448), .A2(n9493), .ZN(n7556) );
  OR2_X1 U9884 ( .A1(n6481), .A2(SI_9_), .ZN(n7555) );
  OAI211_X1 U9885 ( .C1(n10714), .C2(n7450), .A(n7556), .B(n7555), .ZN(n15169)
         );
  NAND2_X1 U9886 ( .A1(n13099), .A2(n15169), .ZN(n12599) );
  INV_X1 U9887 ( .A(n15169), .ZN(n12423) );
  NAND2_X1 U9888 ( .A1(n12352), .A2(n12423), .ZN(n12598) );
  NAND2_X1 U9889 ( .A1(n7522), .A2(P3_REG1_REG_10__SCAN_IN), .ZN(n7562) );
  NAND2_X1 U9890 ( .A1(n12515), .A2(P3_REG0_REG_10__SCAN_IN), .ZN(n7561) );
  NAND2_X1 U9891 ( .A1(n7557), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n7558) );
  NAND2_X1 U9892 ( .A1(n7575), .A2(n7558), .ZN(n13104) );
  NAND2_X1 U9893 ( .A1(n7911), .A2(n13104), .ZN(n7560) );
  NAND2_X1 U9894 ( .A1(n7423), .A2(P3_REG2_REG_10__SCAN_IN), .ZN(n7559) );
  NAND4_X1 U9895 ( .A1(n7562), .A2(n7561), .A3(n7560), .A4(n7559), .ZN(n13086)
         );
  INV_X1 U9896 ( .A(n13086), .ZN(n12461) );
  NAND2_X1 U9897 ( .A1(n9564), .A2(P1_DATAO_REG_10__SCAN_IN), .ZN(n7581) );
  NAND2_X1 U9898 ( .A1(n9559), .A2(P2_DATAO_REG_10__SCAN_IN), .ZN(n7565) );
  OR2_X1 U9899 ( .A1(n7567), .A2(n7566), .ZN(n7568) );
  NAND2_X1 U9900 ( .A1(n7582), .A2(n7568), .ZN(n9443) );
  NAND2_X1 U9901 ( .A1(n9443), .A2(n12520), .ZN(n7572) );
  NAND2_X1 U9902 ( .A1(n7604), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7570) );
  OR2_X1 U9903 ( .A1(n6472), .A2(n11025), .ZN(n7571) );
  OAI211_X1 U9904 ( .C1(SI_10_), .C2(n6480), .A(n7572), .B(n7571), .ZN(n13233)
         );
  INV_X1 U9905 ( .A(n13233), .ZN(n13109) );
  NAND2_X1 U9906 ( .A1(n12461), .A2(n13109), .ZN(n12605) );
  NAND2_X1 U9907 ( .A1(n13086), .A2(n13233), .ZN(n12603) );
  NAND2_X1 U9908 ( .A1(n12605), .A2(n12603), .ZN(n13112) );
  NAND2_X1 U9909 ( .A1(n7522), .A2(P3_REG1_REG_11__SCAN_IN), .ZN(n7580) );
  NAND2_X1 U9910 ( .A1(n12515), .A2(P3_REG0_REG_11__SCAN_IN), .ZN(n7579) );
  NAND2_X1 U9911 ( .A1(n7575), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n7576) );
  NAND2_X1 U9912 ( .A1(n7588), .A2(n7576), .ZN(n13091) );
  NAND2_X1 U9913 ( .A1(n7911), .A2(n13091), .ZN(n7578) );
  NAND2_X1 U9914 ( .A1(n7423), .A2(P3_REG2_REG_11__SCAN_IN), .ZN(n7577) );
  NAND2_X1 U9915 ( .A1(n9574), .A2(P1_DATAO_REG_11__SCAN_IN), .ZN(n7596) );
  NAND2_X1 U9916 ( .A1(n9568), .A2(P2_DATAO_REG_11__SCAN_IN), .ZN(n7583) );
  XNOR2_X1 U9917 ( .A(n7595), .B(n7594), .ZN(n14315) );
  NAND2_X1 U9918 ( .A1(n14315), .A2(n12520), .ZN(n7586) );
  OAI21_X1 U9919 ( .B1(n7604), .B2(P3_IR_REG_10__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n7584) );
  XNOR2_X1 U9920 ( .A(n7584), .B(P3_IR_REG_11__SCAN_IN), .ZN(n11139) );
  AOI22_X1 U9921 ( .A1(n7725), .A2(n8279), .B1(n6482), .B2(n14320), .ZN(n7585)
         );
  NAND2_X1 U9922 ( .A1(n7586), .A2(n7585), .ZN(n14428) );
  INV_X1 U9923 ( .A(n14428), .ZN(n12467) );
  OR2_X1 U9924 ( .A1(n12464), .A2(n12467), .ZN(n12602) );
  NAND2_X1 U9925 ( .A1(n12467), .A2(n12464), .ZN(n12604) );
  NAND2_X1 U9926 ( .A1(n12602), .A2(n12604), .ZN(n12606) );
  NAND2_X1 U9927 ( .A1(n13090), .A2(n7587), .ZN(n13089) );
  NAND2_X1 U9928 ( .A1(n13089), .A2(n12604), .ZN(n13074) );
  NAND2_X1 U9929 ( .A1(n7522), .A2(P3_REG1_REG_12__SCAN_IN), .ZN(n7593) );
  NAND2_X1 U9930 ( .A1(n12514), .A2(P3_REG2_REG_12__SCAN_IN), .ZN(n7592) );
  AND2_X1 U9931 ( .A1(n7588), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n7589) );
  OR2_X1 U9932 ( .A1(n7589), .A2(n7621), .ZN(n13079) );
  NAND2_X1 U9933 ( .A1(n7911), .A2(n13079), .ZN(n7591) );
  NAND2_X1 U9934 ( .A1(n12515), .A2(P3_REG0_REG_12__SCAN_IN), .ZN(n7590) );
  NAND4_X1 U9935 ( .A1(n7593), .A2(n7592), .A3(n7591), .A4(n7590), .ZN(n13087)
         );
  NAND2_X1 U9936 ( .A1(n9613), .A2(P1_DATAO_REG_12__SCAN_IN), .ZN(n7609) );
  NAND2_X1 U9937 ( .A1(n9616), .A2(P2_DATAO_REG_12__SCAN_IN), .ZN(n7597) );
  OR2_X1 U9938 ( .A1(n7599), .A2(n7598), .ZN(n7600) );
  NAND2_X1 U9939 ( .A1(n7610), .A2(n7600), .ZN(n9490) );
  OR2_X1 U9940 ( .A1(n9490), .A2(n7448), .ZN(n7607) );
  INV_X1 U9941 ( .A(P3_IR_REG_10__SCAN_IN), .ZN(n7602) );
  INV_X1 U9942 ( .A(P3_IR_REG_11__SCAN_IN), .ZN(n7601) );
  NAND2_X1 U9943 ( .A1(n7602), .A2(n7601), .ZN(n7603) );
  OR2_X1 U9944 ( .A1(n7614), .A2(n13241), .ZN(n7605) );
  AOI22_X1 U9945 ( .A1(n7725), .A2(SI_12_), .B1(n6482), .B2(n12770), .ZN(n7606) );
  NAND2_X1 U9946 ( .A1(n7607), .A2(n7606), .ZN(n14425) );
  OR2_X1 U9947 ( .A1(n9205), .A2(n14425), .ZN(n12610) );
  NAND2_X1 U9948 ( .A1(n14425), .A2(n9205), .ZN(n12611) );
  NAND2_X1 U9949 ( .A1(n12610), .A2(n12611), .ZN(n13076) );
  INV_X1 U9950 ( .A(n13076), .ZN(n12711) );
  NAND2_X1 U9951 ( .A1(n13074), .A2(n12711), .ZN(n7608) );
  NAND2_X1 U9952 ( .A1(n7611), .A2(n9630), .ZN(n7612) );
  NAND2_X1 U9953 ( .A1(n7628), .A2(n7612), .ZN(n9565) );
  NAND2_X1 U9954 ( .A1(n9565), .A2(n12520), .ZN(n7619) );
  INV_X1 U9955 ( .A(SI_13_), .ZN(n9566) );
  NAND2_X1 U9956 ( .A1(n7614), .A2(n7613), .ZN(n7616) );
  NAND2_X1 U9957 ( .A1(n7616), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7615) );
  MUX2_X1 U9958 ( .A(P3_IR_REG_31__SCAN_IN), .B(n7615), .S(
        P3_IR_REG_13__SCAN_IN), .Z(n7617) );
  AOI22_X1 U9959 ( .A1(n7725), .A2(n9566), .B1(n6482), .B2(n12793), .ZN(n7618)
         );
  NAND2_X1 U9960 ( .A1(n7619), .A2(n7618), .ZN(n14417) );
  OR2_X1 U9961 ( .A1(n7621), .A2(n7620), .ZN(n7622) );
  NAND2_X1 U9962 ( .A1(n7634), .A2(n7622), .ZN(n13065) );
  NAND2_X1 U9963 ( .A1(n7911), .A2(n13065), .ZN(n7626) );
  NAND2_X1 U9964 ( .A1(n7522), .A2(P3_REG1_REG_13__SCAN_IN), .ZN(n7625) );
  NAND2_X1 U9965 ( .A1(n12515), .A2(P3_REG0_REG_13__SCAN_IN), .ZN(n7624) );
  NAND2_X1 U9966 ( .A1(n12514), .A2(P3_REG2_REG_13__SCAN_IN), .ZN(n7623) );
  NAND2_X1 U9967 ( .A1(n14417), .A2(n13050), .ZN(n12618) );
  INV_X1 U9968 ( .A(n13059), .ZN(n7640) );
  NAND2_X1 U9969 ( .A1(n9881), .A2(P1_DATAO_REG_14__SCAN_IN), .ZN(n7644) );
  NAND2_X1 U9970 ( .A1(n9876), .A2(P2_DATAO_REG_14__SCAN_IN), .ZN(n7629) );
  XNOR2_X1 U9971 ( .A(n7643), .B(n7642), .ZN(n9575) );
  NAND2_X1 U9972 ( .A1(n9575), .A2(n12520), .ZN(n7633) );
  NAND2_X1 U9973 ( .A1(n7649), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7631) );
  INV_X1 U9974 ( .A(P3_IR_REG_14__SCAN_IN), .ZN(n7630) );
  XNOR2_X1 U9975 ( .A(n7631), .B(n7630), .ZN(n12790) );
  AOI22_X1 U9976 ( .A1(n7725), .A2(n6890), .B1(n6482), .B2(n12790), .ZN(n7632)
         );
  NAND2_X1 U9977 ( .A1(n7633), .A2(n7632), .ZN(n14413) );
  NAND2_X1 U9978 ( .A1(n7423), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n7639) );
  NAND2_X1 U9979 ( .A1(n7522), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n7638) );
  NAND2_X1 U9980 ( .A1(n7634), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n7635) );
  NAND2_X1 U9981 ( .A1(n7654), .A2(n7635), .ZN(n13053) );
  NAND2_X1 U9982 ( .A1(n7911), .A2(n13053), .ZN(n7637) );
  NAND2_X1 U9983 ( .A1(n12515), .A2(P3_REG0_REG_14__SCAN_IN), .ZN(n7636) );
  NAND2_X1 U9984 ( .A1(n14413), .A2(n13063), .ZN(n12622) );
  NAND2_X1 U9985 ( .A1(n7641), .A2(n12621), .ZN(n13036) );
  NAND2_X1 U9986 ( .A1(n10132), .A2(P1_DATAO_REG_15__SCAN_IN), .ZN(n7661) );
  NAND2_X1 U9987 ( .A1(n10134), .A2(P2_DATAO_REG_15__SCAN_IN), .ZN(n7645) );
  OR2_X1 U9988 ( .A1(n7647), .A2(n7646), .ZN(n7648) );
  NAND2_X1 U9989 ( .A1(n7662), .A2(n7648), .ZN(n9638) );
  NAND2_X1 U9990 ( .A1(n9638), .A2(n12520), .ZN(n7653) );
  OAI21_X1 U9991 ( .B1(n7649), .B2(P3_IR_REG_14__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n7650) );
  XNOR2_X1 U9992 ( .A(n7650), .B(P3_IR_REG_15__SCAN_IN), .ZN(n14344) );
  OAI22_X1 U9993 ( .A1(n6480), .A2(SI_15_), .B1(n14344), .B2(n6472), .ZN(n7651) );
  INV_X1 U9994 ( .A(n7651), .ZN(n7652) );
  NAND2_X1 U9995 ( .A1(n7423), .A2(P3_REG2_REG_15__SCAN_IN), .ZN(n7660) );
  NAND2_X1 U9996 ( .A1(n7522), .A2(P3_REG1_REG_15__SCAN_IN), .ZN(n7659) );
  INV_X1 U9997 ( .A(n7672), .ZN(n7656) );
  NAND2_X1 U9998 ( .A1(n7654), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n7655) );
  NAND2_X1 U9999 ( .A1(n7656), .A2(n7655), .ZN(n13042) );
  NAND2_X1 U10000 ( .A1(n7911), .A2(n13042), .ZN(n7658) );
  NAND2_X1 U10001 ( .A1(n12515), .A2(P3_REG0_REG_15__SCAN_IN), .ZN(n7657) );
  NAND2_X1 U10002 ( .A1(n13231), .A2(n13051), .ZN(n12625) );
  NAND2_X1 U10003 ( .A1(n10210), .A2(P1_DATAO_REG_16__SCAN_IN), .ZN(n7684) );
  NAND2_X1 U10004 ( .A1(n10212), .A2(P2_DATAO_REG_16__SCAN_IN), .ZN(n7663) );
  OR2_X1 U10005 ( .A1(n7665), .A2(n7664), .ZN(n7666) );
  NAND2_X1 U10006 ( .A1(n7685), .A2(n7666), .ZN(n9680) );
  OR2_X1 U10007 ( .A1(n9680), .A2(n7448), .ZN(n7671) );
  NAND2_X1 U10008 ( .A1(n7668), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7669) );
  XNOR2_X1 U10009 ( .A(n7669), .B(P3_IR_REG_16__SCAN_IN), .ZN(n14361) );
  AOI22_X1 U10010 ( .A1(n7725), .A2(SI_16_), .B1(n6482), .B2(n14361), .ZN(
        n7670) );
  NAND2_X1 U10011 ( .A1(n12514), .A2(P3_REG2_REG_16__SCAN_IN), .ZN(n7677) );
  NAND2_X1 U10012 ( .A1(n7522), .A2(P3_REG1_REG_16__SCAN_IN), .ZN(n7676) );
  NOR2_X1 U10013 ( .A1(n7672), .A2(n12401), .ZN(n7673) );
  OR2_X1 U10014 ( .A1(n7695), .A2(n7673), .ZN(n13031) );
  NAND2_X1 U10015 ( .A1(n7911), .A2(n13031), .ZN(n7675) );
  NAND2_X1 U10016 ( .A1(n12515), .A2(P3_REG0_REG_16__SCAN_IN), .ZN(n7674) );
  NAND2_X1 U10017 ( .A1(n13167), .A2(n13017), .ZN(n12630) );
  INV_X1 U10018 ( .A(n12630), .ZN(n12627) );
  XNOR2_X1 U10019 ( .A(n13167), .B(n12757), .ZN(n13027) );
  OR2_X1 U10020 ( .A1(n12627), .A2(n13027), .ZN(n7679) );
  AND2_X1 U10021 ( .A1(n13038), .A2(n7679), .ZN(n7678) );
  NAND2_X1 U10022 ( .A1(n13036), .A2(n7678), .ZN(n7683) );
  INV_X1 U10023 ( .A(n7679), .ZN(n7681) );
  AND2_X1 U10024 ( .A1(n13024), .A2(n12630), .ZN(n7680) );
  NAND2_X1 U10025 ( .A1(n7683), .A2(n7682), .ZN(n13012) );
  NAND2_X1 U10026 ( .A1(n10312), .A2(P1_DATAO_REG_17__SCAN_IN), .ZN(n7703) );
  INV_X1 U10027 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n10314) );
  NAND2_X1 U10028 ( .A1(n10314), .A2(P2_DATAO_REG_17__SCAN_IN), .ZN(n7686) );
  XNOR2_X1 U10029 ( .A(n7702), .B(n7701), .ZN(n9765) );
  NAND2_X1 U10030 ( .A1(n9765), .A2(n12520), .ZN(n7694) );
  INV_X1 U10031 ( .A(n7687), .ZN(n7688) );
  NAND2_X1 U10032 ( .A1(n7688), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7689) );
  MUX2_X1 U10033 ( .A(P3_IR_REG_31__SCAN_IN), .B(n7689), .S(
        P3_IR_REG_17__SCAN_IN), .Z(n7690) );
  INV_X1 U10034 ( .A(n7690), .ZN(n7692) );
  NOR2_X1 U10035 ( .A1(n7692), .A2(n7691), .ZN(n14379) );
  AOI22_X1 U10036 ( .A1(n7725), .A2(n9764), .B1(n6482), .B2(n12848), .ZN(n7693) );
  NAND2_X1 U10037 ( .A1(n7522), .A2(P3_REG1_REG_17__SCAN_IN), .ZN(n7700) );
  NAND2_X1 U10038 ( .A1(n12514), .A2(P3_REG2_REG_17__SCAN_IN), .ZN(n7699) );
  OR2_X1 U10039 ( .A1(n7695), .A2(n9125), .ZN(n7696) );
  NAND2_X1 U10040 ( .A1(n7711), .A2(n7696), .ZN(n13019) );
  NAND2_X1 U10041 ( .A1(n7911), .A2(n13019), .ZN(n7698) );
  NAND2_X1 U10042 ( .A1(n12515), .A2(P3_REG0_REG_17__SCAN_IN), .ZN(n7697) );
  NAND4_X1 U10043 ( .A1(n7700), .A2(n7699), .A3(n7698), .A4(n7697), .ZN(n12756) );
  NAND2_X1 U10044 ( .A1(n13226), .A2(n12756), .ZN(n12634) );
  NAND2_X1 U10045 ( .A1(n12638), .A2(n12634), .ZN(n13015) );
  INV_X1 U10046 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n10682) );
  NAND2_X1 U10047 ( .A1(n10682), .A2(P1_DATAO_REG_18__SCAN_IN), .ZN(n7717) );
  INV_X1 U10048 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n10678) );
  NAND2_X1 U10049 ( .A1(n10678), .A2(P2_DATAO_REG_18__SCAN_IN), .ZN(n7704) );
  OR2_X1 U10050 ( .A1(n7706), .A2(n7705), .ZN(n7707) );
  NAND2_X1 U10051 ( .A1(n7718), .A2(n7707), .ZN(n9882) );
  OR2_X1 U10052 ( .A1(n9882), .A2(n7448), .ZN(n7710) );
  OR2_X1 U10053 ( .A1(n7691), .A2(n13241), .ZN(n7708) );
  XNOR2_X1 U10054 ( .A(n7708), .B(n7723), .ZN(n12840) );
  AOI22_X1 U10055 ( .A1(n7725), .A2(SI_18_), .B1(n6482), .B2(n14394), .ZN(
        n7709) );
  NAND2_X1 U10056 ( .A1(n7711), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n7712) );
  NAND2_X1 U10057 ( .A1(n7728), .A2(n7712), .ZN(n13005) );
  NAND2_X1 U10058 ( .A1(n13005), .A2(n7911), .ZN(n7716) );
  NAND2_X1 U10059 ( .A1(n7522), .A2(P3_REG1_REG_18__SCAN_IN), .ZN(n7715) );
  NAND2_X1 U10060 ( .A1(n12515), .A2(P3_REG0_REG_18__SCAN_IN), .ZN(n7714) );
  NAND2_X1 U10061 ( .A1(n7423), .A2(P3_REG2_REG_18__SCAN_IN), .ZN(n7713) );
  NAND4_X1 U10062 ( .A1(n7716), .A2(n7715), .A3(n7714), .A4(n7713), .ZN(n12755) );
  NAND2_X1 U10063 ( .A1(n13004), .A2(n13018), .ZN(n12641) );
  INV_X1 U10064 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n11654) );
  NAND2_X1 U10065 ( .A1(n11654), .A2(P1_DATAO_REG_19__SCAN_IN), .ZN(n7733) );
  INV_X1 U10066 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n10764) );
  NAND2_X1 U10067 ( .A1(n10764), .A2(P2_DATAO_REG_19__SCAN_IN), .ZN(n7719) );
  OR2_X1 U10068 ( .A1(n7721), .A2(n7720), .ZN(n7722) );
  NAND2_X1 U10069 ( .A1(n7734), .A2(n7722), .ZN(n9991) );
  OR2_X1 U10070 ( .A1(n9991), .A2(n7448), .ZN(n7727) );
  OR2_X1 U10071 ( .A1(n7851), .A2(n13241), .ZN(n7724) );
  XNOR2_X2 U10072 ( .A(n7724), .B(P3_IR_REG_19__SCAN_IN), .ZN(n12825) );
  AOI22_X1 U10073 ( .A1(n7725), .A2(SI_19_), .B1(n6482), .B2(n12825), .ZN(
        n7726) );
  INV_X1 U10074 ( .A(P3_REG0_REG_19__SCAN_IN), .ZN(n13216) );
  AND2_X1 U10075 ( .A1(n7728), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n7729) );
  OR2_X1 U10076 ( .A1(n7729), .A2(n7740), .ZN(n12992) );
  NAND2_X1 U10077 ( .A1(n12992), .A2(n7911), .ZN(n7731) );
  AOI22_X1 U10078 ( .A1(P3_REG2_REG_19__SCAN_IN), .A2(n12514), .B1(n7522), 
        .B2(P3_REG1_REG_19__SCAN_IN), .ZN(n7730) );
  OAI211_X1 U10079 ( .C1(n7471), .C2(n13216), .A(n7731), .B(n7730), .ZN(n12754) );
  OR2_X1 U10080 ( .A1(n12991), .A2(n13003), .ZN(n12646) );
  AND2_X1 U10081 ( .A1(n12646), .A2(n12985), .ZN(n12637) );
  NAND2_X1 U10082 ( .A1(n12991), .A2(n13003), .ZN(n12647) );
  NAND2_X1 U10083 ( .A1(n7736), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n7737) );
  NAND2_X1 U10084 ( .A1(n7745), .A2(n7737), .ZN(n10286) );
  OR2_X1 U10085 ( .A1(n10286), .A2(n7448), .ZN(n7739) );
  OR2_X1 U10086 ( .A1(n6481), .A2(n10287), .ZN(n7738) );
  INV_X1 U10087 ( .A(P3_REG0_REG_20__SCAN_IN), .ZN(n13211) );
  NOR2_X1 U10088 ( .A1(n7740), .A2(n9134), .ZN(n7741) );
  OR2_X1 U10089 ( .A1(n7751), .A2(n7741), .ZN(n12977) );
  NAND2_X1 U10090 ( .A1(n12977), .A2(n7911), .ZN(n7743) );
  AOI22_X1 U10091 ( .A1(n7423), .A2(P3_REG2_REG_20__SCAN_IN), .B1(n7522), .B2(
        P3_REG1_REG_20__SCAN_IN), .ZN(n7742) );
  INV_X1 U10092 ( .A(n12753), .ZN(n12990) );
  NAND2_X1 U10093 ( .A1(n13145), .A2(n12990), .ZN(n12651) );
  INV_X1 U10094 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n11515) );
  NAND2_X1 U10095 ( .A1(n11515), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n7758) );
  INV_X1 U10096 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n10977) );
  NAND2_X1 U10097 ( .A1(n10977), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n7746) );
  AND2_X1 U10098 ( .A1(n7758), .A2(n7746), .ZN(n7747) );
  OR2_X1 U10099 ( .A1(n7748), .A2(n7747), .ZN(n7749) );
  NAND2_X1 U10100 ( .A1(n7759), .A2(n7749), .ZN(n10422) );
  INV_X1 U10101 ( .A(SI_21_), .ZN(n10423) );
  INV_X1 U10102 ( .A(P3_REG0_REG_21__SCAN_IN), .ZN(n13208) );
  INV_X1 U10103 ( .A(P3_REG3_REG_21__SCAN_IN), .ZN(n12367) );
  OR2_X1 U10104 ( .A1(n7751), .A2(n12367), .ZN(n7752) );
  NAND2_X1 U10105 ( .A1(n7762), .A2(n7752), .ZN(n12966) );
  NAND2_X1 U10106 ( .A1(n12966), .A2(n7911), .ZN(n7754) );
  AOI22_X1 U10107 ( .A1(n12514), .A2(P3_REG2_REG_21__SCAN_IN), .B1(n7522), 
        .B2(P3_REG1_REG_21__SCAN_IN), .ZN(n7753) );
  NAND2_X1 U10108 ( .A1(n12545), .A2(n12973), .ZN(n7755) );
  NAND2_X1 U10109 ( .A1(n12960), .A2(n7755), .ZN(n7757) );
  OR2_X1 U10110 ( .A1(n12545), .A2(n12973), .ZN(n7756) );
  NAND2_X1 U10111 ( .A1(n7757), .A2(n7756), .ZN(n12945) );
  XNOR2_X1 U10112 ( .A(n11651), .B(P2_DATAO_REG_22__SCAN_IN), .ZN(n7772) );
  XNOR2_X1 U10113 ( .A(n7773), .B(n7772), .ZN(n10605) );
  NAND2_X1 U10114 ( .A1(n10605), .A2(n12520), .ZN(n7761) );
  OR2_X1 U10115 ( .A1(n6480), .A2(n8565), .ZN(n7760) );
  NAND2_X1 U10116 ( .A1(n7762), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n7763) );
  INV_X1 U10117 ( .A(n7776), .ZN(n7777) );
  NAND2_X1 U10118 ( .A1(n7763), .A2(n7777), .ZN(n12955) );
  NAND2_X1 U10119 ( .A1(n12955), .A2(n7911), .ZN(n7769) );
  INV_X1 U10120 ( .A(P3_REG2_REG_22__SCAN_IN), .ZN(n7766) );
  NAND2_X1 U10121 ( .A1(n12515), .A2(P3_REG0_REG_22__SCAN_IN), .ZN(n7765) );
  NAND2_X1 U10122 ( .A1(n7522), .A2(P3_REG1_REG_22__SCAN_IN), .ZN(n7764) );
  OAI211_X1 U10123 ( .C1(n7468), .C2(n7766), .A(n7765), .B(n7764), .ZN(n7767)
         );
  INV_X1 U10124 ( .A(n7767), .ZN(n7768) );
  INV_X1 U10125 ( .A(n12751), .ZN(n7770) );
  NAND2_X1 U10126 ( .A1(n12954), .A2(n7770), .ZN(n12658) );
  NAND2_X1 U10127 ( .A1(n12945), .A2(n12658), .ZN(n7771) );
  XNOR2_X1 U10128 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(P2_DATAO_REG_23__SCAN_IN), 
        .ZN(n7783) );
  XNOR2_X1 U10129 ( .A(n7784), .B(n7783), .ZN(n10762) );
  NAND2_X1 U10130 ( .A1(n10762), .A2(n12520), .ZN(n7775) );
  OR2_X1 U10131 ( .A1(n6481), .A2(n9113), .ZN(n7774) );
  NAND2_X1 U10132 ( .A1(n7423), .A2(P3_REG2_REG_23__SCAN_IN), .ZN(n7782) );
  NAND2_X1 U10133 ( .A1(n7522), .A2(P3_REG1_REG_23__SCAN_IN), .ZN(n7781) );
  INV_X1 U10134 ( .A(P3_REG3_REG_23__SCAN_IN), .ZN(n12340) );
  NAND2_X1 U10135 ( .A1(n12340), .A2(n7776), .ZN(n7793) );
  NAND2_X1 U10136 ( .A1(P3_REG3_REG_23__SCAN_IN), .A2(n7777), .ZN(n7778) );
  NAND2_X1 U10137 ( .A1(n7793), .A2(n7778), .ZN(n12940) );
  NAND2_X1 U10138 ( .A1(n7911), .A2(n12940), .ZN(n7780) );
  NAND2_X1 U10139 ( .A1(n12515), .A2(P3_REG0_REG_23__SCAN_IN), .ZN(n7779) );
  NAND2_X1 U10140 ( .A1(n13134), .A2(n12450), .ZN(n12661) );
  INV_X1 U10141 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n11269) );
  NAND2_X1 U10142 ( .A1(n11269), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n7785) );
  INV_X1 U10143 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n11396) );
  NAND2_X1 U10144 ( .A1(n7787), .A2(n11396), .ZN(n7788) );
  INV_X1 U10145 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n12153) );
  XNOR2_X1 U10146 ( .A(n7800), .B(n12153), .ZN(n10909) );
  NAND2_X1 U10147 ( .A1(n10909), .A2(n12520), .ZN(n7790) );
  NAND2_X1 U10148 ( .A1(n7423), .A2(P3_REG2_REG_24__SCAN_IN), .ZN(n7798) );
  NAND2_X1 U10149 ( .A1(n7522), .A2(P3_REG1_REG_24__SCAN_IN), .ZN(n7797) );
  INV_X1 U10150 ( .A(n7793), .ZN(n7792) );
  INV_X1 U10151 ( .A(P3_REG3_REG_24__SCAN_IN), .ZN(n7791) );
  NAND2_X1 U10152 ( .A1(n7793), .A2(P3_REG3_REG_24__SCAN_IN), .ZN(n7794) );
  NAND2_X1 U10153 ( .A1(n7804), .A2(n7794), .ZN(n12923) );
  NAND2_X1 U10154 ( .A1(n7911), .A2(n12923), .ZN(n7796) );
  NAND2_X1 U10155 ( .A1(n12515), .A2(P3_REG0_REG_24__SCAN_IN), .ZN(n7795) );
  NAND2_X1 U10156 ( .A1(n12922), .A2(n12389), .ZN(n12667) );
  INV_X1 U10157 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n13823) );
  XNOR2_X1 U10158 ( .A(n13823), .B(P2_DATAO_REG_25__SCAN_IN), .ZN(n7801) );
  XNOR2_X1 U10159 ( .A(n7811), .B(n7801), .ZN(n11102) );
  NAND2_X1 U10160 ( .A1(n11102), .A2(n12520), .ZN(n7803) );
  INV_X1 U10161 ( .A(SI_25_), .ZN(n11104) );
  OR2_X1 U10162 ( .A1(n6480), .A2(n11104), .ZN(n7802) );
  NAND2_X1 U10163 ( .A1(n12514), .A2(P3_REG2_REG_25__SCAN_IN), .ZN(n7809) );
  NAND2_X1 U10164 ( .A1(n7522), .A2(P3_REG1_REG_25__SCAN_IN), .ZN(n7808) );
  NAND2_X1 U10165 ( .A1(n7804), .A2(P3_REG3_REG_25__SCAN_IN), .ZN(n7805) );
  NAND2_X1 U10166 ( .A1(n7817), .A2(n7805), .ZN(n12906) );
  NAND2_X1 U10167 ( .A1(n7911), .A2(n12906), .ZN(n7807) );
  NAND2_X1 U10168 ( .A1(n12515), .A2(P3_REG0_REG_25__SCAN_IN), .ZN(n7806) );
  OR2_X1 U10169 ( .A1(n12382), .A2(n12415), .ZN(n12673) );
  NAND2_X1 U10170 ( .A1(n12382), .A2(n12415), .ZN(n12672) );
  NAND2_X1 U10171 ( .A1(n12673), .A2(n12672), .ZN(n12901) );
  INV_X1 U10172 ( .A(n12901), .ZN(n12665) );
  NAND2_X1 U10173 ( .A1(n13823), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n7810) );
  INV_X1 U10174 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n12318) );
  NAND2_X1 U10175 ( .A1(n12318), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n7812) );
  INV_X1 U10176 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n11397) );
  XNOR2_X1 U10177 ( .A(n11397), .B(P2_DATAO_REG_26__SCAN_IN), .ZN(n7813) );
  XNOR2_X1 U10178 ( .A(n7824), .B(n7813), .ZN(n11200) );
  NAND2_X1 U10179 ( .A1(n11200), .A2(n12520), .ZN(n7815) );
  NAND2_X1 U10180 ( .A1(n7522), .A2(P3_REG1_REG_26__SCAN_IN), .ZN(n7822) );
  NAND2_X1 U10181 ( .A1(n12514), .A2(P3_REG2_REG_26__SCAN_IN), .ZN(n7821) );
  INV_X1 U10182 ( .A(n7817), .ZN(n7816) );
  INV_X1 U10183 ( .A(P3_REG3_REG_26__SCAN_IN), .ZN(n12485) );
  NAND2_X1 U10184 ( .A1(n7816), .A2(n12485), .ZN(n7829) );
  NAND2_X1 U10185 ( .A1(n7817), .A2(P3_REG3_REG_26__SCAN_IN), .ZN(n7818) );
  NAND2_X1 U10186 ( .A1(n7829), .A2(n7818), .ZN(n12894) );
  NAND2_X1 U10187 ( .A1(n7911), .A2(n12894), .ZN(n7820) );
  NAND2_X1 U10188 ( .A1(n12515), .A2(P3_REG0_REG_26__SCAN_IN), .ZN(n7819) );
  NAND4_X1 U10189 ( .A1(n7822), .A2(n7821), .A3(n7820), .A4(n7819), .ZN(n12747) );
  INV_X1 U10190 ( .A(n12747), .ZN(n9266) );
  NAND2_X1 U10191 ( .A1(n12480), .A2(n9266), .ZN(n12539) );
  INV_X1 U10192 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n11564) );
  AND2_X1 U10193 ( .A1(n11564), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n7823) );
  NAND2_X1 U10194 ( .A1(n11397), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n7825) );
  XNOR2_X1 U10195 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(P2_DATAO_REG_27__SCAN_IN), 
        .ZN(n7826) );
  XNOR2_X1 U10196 ( .A(n7837), .B(n7826), .ZN(n11272) );
  NAND2_X1 U10197 ( .A1(n11272), .A2(n12520), .ZN(n7828) );
  INV_X1 U10198 ( .A(SI_27_), .ZN(n11273) );
  OR2_X1 U10199 ( .A1(n6480), .A2(n11273), .ZN(n7827) );
  NAND2_X1 U10200 ( .A1(n12514), .A2(P3_REG2_REG_27__SCAN_IN), .ZN(n7834) );
  NAND2_X1 U10201 ( .A1(n7522), .A2(P3_REG1_REG_27__SCAN_IN), .ZN(n7833) );
  NAND2_X1 U10202 ( .A1(n7829), .A2(P3_REG3_REG_27__SCAN_IN), .ZN(n7830) );
  NAND2_X1 U10203 ( .A1(n7843), .A2(n7830), .ZN(n12883) );
  NAND2_X1 U10204 ( .A1(n7911), .A2(n12883), .ZN(n7832) );
  NAND2_X1 U10205 ( .A1(n12515), .A2(P3_REG0_REG_27__SCAN_IN), .ZN(n7831) );
  INV_X1 U10206 ( .A(n12746), .ZN(n12536) );
  NAND2_X1 U10207 ( .A1(n12535), .A2(n12536), .ZN(n8861) );
  NAND2_X1 U10208 ( .A1(n8884), .A2(n8861), .ZN(n7849) );
  INV_X1 U10209 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n13817) );
  AND2_X1 U10210 ( .A1(n13817), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n7836) );
  INV_X1 U10211 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n11665) );
  NAND2_X1 U10212 ( .A1(n11665), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n7835) );
  INV_X1 U10213 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n8866) );
  XNOR2_X1 U10214 ( .A(n8866), .B(P2_DATAO_REG_28__SCAN_IN), .ZN(n7838) );
  XNOR2_X1 U10215 ( .A(n8865), .B(n7838), .ZN(n13246) );
  NAND2_X1 U10216 ( .A1(n13246), .A2(n12520), .ZN(n7840) );
  INV_X1 U10217 ( .A(SI_28_), .ZN(n13248) );
  OR2_X1 U10218 ( .A1(n6481), .A2(n13248), .ZN(n7839) );
  NAND2_X1 U10219 ( .A1(n7422), .A2(P3_REG1_REG_28__SCAN_IN), .ZN(n7848) );
  NAND2_X1 U10220 ( .A1(n12515), .A2(P3_REG0_REG_28__SCAN_IN), .ZN(n7847) );
  INV_X1 U10221 ( .A(n7843), .ZN(n7842) );
  INV_X1 U10222 ( .A(P3_REG3_REG_28__SCAN_IN), .ZN(n7841) );
  NAND2_X1 U10223 ( .A1(n7842), .A2(n7841), .ZN(n12862) );
  NAND2_X1 U10224 ( .A1(n7843), .A2(P3_REG3_REG_28__SCAN_IN), .ZN(n7844) );
  NAND2_X1 U10225 ( .A1(n12862), .A2(n7844), .ZN(n12875) );
  NAND2_X1 U10226 ( .A1(n7911), .A2(n12875), .ZN(n7846) );
  NAND2_X1 U10227 ( .A1(n12514), .A2(P3_REG2_REG_28__SCAN_IN), .ZN(n7845) );
  NAND4_X1 U10228 ( .A1(n7848), .A2(n7847), .A3(n7846), .A4(n7845), .ZN(n12745) );
  INV_X1 U10229 ( .A(n12745), .ZN(n8871) );
  OR2_X2 U10230 ( .A1(n7954), .A2(n8871), .ZN(n12679) );
  NAND2_X1 U10231 ( .A1(n7954), .A2(n8871), .ZN(n8862) );
  NAND2_X1 U10232 ( .A1(n12679), .A2(n8862), .ZN(n12542) );
  XNOR2_X1 U10233 ( .A(n7849), .B(n12685), .ZN(n12879) );
  NAND2_X1 U10234 ( .A1(n7947), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7852) );
  XNOR2_X2 U10235 ( .A(n7855), .B(n7854), .ZN(n10288) );
  NAND2_X1 U10236 ( .A1(n12739), .A2(n10288), .ZN(n7856) );
  NAND2_X1 U10237 ( .A1(n7856), .A2(n12825), .ZN(n7859) );
  NAND2_X1 U10238 ( .A1(n7857), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7858) );
  XNOR2_X2 U10239 ( .A(n7858), .B(P3_IR_REG_21__SCAN_IN), .ZN(n12547) );
  INV_X1 U10240 ( .A(n12547), .ZN(n12552) );
  NAND2_X1 U10241 ( .A1(n7859), .A2(n12552), .ZN(n7862) );
  INV_X1 U10242 ( .A(n10288), .ZN(n7964) );
  NOR2_X1 U10243 ( .A1(n12547), .A2(n7964), .ZN(n7860) );
  OR2_X1 U10244 ( .A1(n12739), .A2(n7860), .ZN(n7861) );
  NAND2_X1 U10245 ( .A1(n7862), .A2(n7861), .ZN(n9252) );
  NAND2_X1 U10246 ( .A1(n10288), .A2(n12857), .ZN(n9262) );
  NAND3_X1 U10247 ( .A1(n9252), .A2(n12735), .A3(n15170), .ZN(n7864) );
  NOR2_X1 U10248 ( .A1(n10288), .A2(n12825), .ZN(n7863) );
  NAND2_X1 U10249 ( .A1(n12739), .A2(n7863), .ZN(n7962) );
  NAND2_X1 U10250 ( .A1(n10288), .A2(n12825), .ZN(n10027) );
  OR2_X1 U10251 ( .A1(n12739), .A2(n10027), .ZN(n15171) );
  NAND2_X1 U10252 ( .A1(n12879), .A2(n15167), .ZN(n7920) );
  INV_X1 U10253 ( .A(n10104), .ZN(n10032) );
  NAND2_X1 U10254 ( .A1(n12766), .A2(n10032), .ZN(n10412) );
  NAND2_X1 U10255 ( .A1(n15114), .A2(n15113), .ZN(n7866) );
  INV_X1 U10256 ( .A(n12556), .ZN(n7865) );
  NAND2_X1 U10257 ( .A1(n7866), .A2(n7865), .ZN(n15117) );
  NAND2_X1 U10258 ( .A1(n10204), .A2(n15107), .ZN(n10728) );
  AND2_X1 U10259 ( .A1(n10727), .A2(n10728), .ZN(n7867) );
  NAND2_X1 U10260 ( .A1(n15117), .A2(n7867), .ZN(n10729) );
  NAND2_X1 U10261 ( .A1(n12763), .A2(n7868), .ZN(n7869) );
  NAND2_X1 U10262 ( .A1(n10729), .A2(n7869), .ZN(n10517) );
  NAND2_X1 U10263 ( .A1(n10517), .A2(n12698), .ZN(n7871) );
  NAND2_X1 U10264 ( .A1(n12762), .A2(n10661), .ZN(n7870) );
  NAND2_X1 U10265 ( .A1(n10876), .A2(n15146), .ZN(n10878) );
  AND2_X1 U10266 ( .A1(n12704), .A2(n10878), .ZN(n7873) );
  NAND2_X1 U10267 ( .A1(n12760), .A2(n15151), .ZN(n7874) );
  NAND2_X1 U10268 ( .A1(n12759), .A2(n12588), .ZN(n7875) );
  NAND2_X1 U10269 ( .A1(n12598), .A2(n12599), .ZN(n12593) );
  NAND2_X1 U10270 ( .A1(n7876), .A2(n15163), .ZN(n11064) );
  AND2_X1 U10271 ( .A1(n12593), .A2(n11064), .ZN(n7877) );
  NAND2_X1 U10272 ( .A1(n13099), .A2(n12423), .ZN(n7878) );
  NAND2_X1 U10273 ( .A1(n11065), .A2(n7878), .ZN(n13097) );
  NAND2_X1 U10274 ( .A1(n13097), .A2(n13112), .ZN(n7880) );
  NAND2_X1 U10275 ( .A1(n13086), .A2(n13109), .ZN(n7879) );
  NAND2_X1 U10276 ( .A1(n7880), .A2(n7879), .ZN(n13085) );
  NAND2_X1 U10277 ( .A1(n13085), .A2(n12606), .ZN(n7882) );
  OR2_X1 U10278 ( .A1(n12464), .A2(n14428), .ZN(n7881) );
  NAND2_X1 U10279 ( .A1(n7882), .A2(n7881), .ZN(n13075) );
  NAND2_X1 U10280 ( .A1(n13075), .A2(n13076), .ZN(n7884) );
  NAND2_X1 U10281 ( .A1(n14425), .A2(n13087), .ZN(n7883) );
  NAND2_X1 U10282 ( .A1(n7884), .A2(n7883), .ZN(n13062) );
  NAND2_X1 U10283 ( .A1(n12617), .A2(n12618), .ZN(n13070) );
  NAND2_X1 U10284 ( .A1(n13062), .A2(n13070), .ZN(n7886) );
  OR2_X1 U10285 ( .A1(n14417), .A2(n12437), .ZN(n7885) );
  NAND2_X1 U10286 ( .A1(n7886), .A2(n7885), .ZN(n13048) );
  NAND2_X1 U10287 ( .A1(n12621), .A2(n12622), .ZN(n13058) );
  NAND2_X1 U10288 ( .A1(n13048), .A2(n13058), .ZN(n7888) );
  OR2_X1 U10289 ( .A1(n14413), .A2(n12493), .ZN(n7887) );
  NAND2_X1 U10290 ( .A1(n7888), .A2(n7887), .ZN(n13037) );
  NAND2_X1 U10291 ( .A1(n13231), .A2(n12332), .ZN(n7889) );
  NOR2_X1 U10292 ( .A1(n13167), .A2(n12757), .ZN(n7890) );
  NAND2_X1 U10293 ( .A1(n13014), .A2(n13015), .ZN(n7892) );
  INV_X1 U10294 ( .A(n12756), .ZN(n13002) );
  OR2_X1 U10295 ( .A1(n13226), .A2(n13002), .ZN(n7891) );
  NAND2_X1 U10296 ( .A1(n7892), .A2(n7891), .ZN(n12999) );
  INV_X1 U10297 ( .A(n12999), .ZN(n7894) );
  OR2_X1 U10298 ( .A1(n13004), .A2(n12755), .ZN(n7895) );
  NAND2_X1 U10299 ( .A1(n12997), .A2(n7895), .ZN(n12987) );
  NAND2_X1 U10300 ( .A1(n12991), .A2(n12754), .ZN(n7896) );
  NAND2_X1 U10301 ( .A1(n12987), .A2(n7896), .ZN(n7898) );
  OR2_X1 U10302 ( .A1(n12991), .A2(n12754), .ZN(n7897) );
  OR2_X1 U10303 ( .A1(n12971), .A2(n7360), .ZN(n12946) );
  OR2_X1 U10304 ( .A1(n12946), .A2(n6515), .ZN(n12932) );
  OR2_X1 U10305 ( .A1(n12932), .A2(n12930), .ZN(n7900) );
  NAND2_X1 U10306 ( .A1(n13145), .A2(n12753), .ZN(n12961) );
  OR2_X1 U10307 ( .A1(n7360), .A2(n7899), .ZN(n12947) );
  INV_X1 U10308 ( .A(n12450), .ZN(n12750) );
  NAND2_X1 U10309 ( .A1(n13134), .A2(n12750), .ZN(n7901) );
  NAND2_X1 U10310 ( .A1(n12917), .A2(n12916), .ZN(n12915) );
  INV_X1 U10311 ( .A(n12389), .ZN(n12749) );
  NAND2_X1 U10312 ( .A1(n12922), .A2(n12749), .ZN(n7902) );
  NAND2_X1 U10313 ( .A1(n12915), .A2(n7902), .ZN(n12902) );
  NAND2_X1 U10314 ( .A1(n12902), .A2(n12901), .ZN(n12900) );
  INV_X1 U10315 ( .A(n12415), .ZN(n12748) );
  NAND2_X1 U10316 ( .A1(n12382), .A2(n12748), .ZN(n7903) );
  NAND2_X1 U10317 ( .A1(n12900), .A2(n7903), .ZN(n12889) );
  OR2_X1 U10318 ( .A1(n12480), .A2(n12747), .ZN(n7904) );
  NAND2_X1 U10319 ( .A1(n12480), .A2(n12747), .ZN(n7905) );
  OR2_X1 U10320 ( .A1(n12535), .A2(n12746), .ZN(n7906) );
  NAND2_X1 U10321 ( .A1(n8888), .A2(n7906), .ZN(n7907) );
  NAND2_X1 U10322 ( .A1(n7907), .A2(n12685), .ZN(n7908) );
  AND2_X1 U10323 ( .A1(n12739), .A2(n12825), .ZN(n7944) );
  AND2_X1 U10324 ( .A1(n7964), .A2(n12547), .ZN(n12733) );
  NAND2_X1 U10325 ( .A1(n7908), .A2(n13103), .ZN(n7909) );
  OR2_X1 U10326 ( .A1(n8869), .A2(n7909), .ZN(n7919) );
  INV_X1 U10327 ( .A(n12862), .ZN(n7910) );
  NAND2_X1 U10328 ( .A1(n7911), .A2(n7910), .ZN(n12519) );
  NAND2_X1 U10329 ( .A1(n12514), .A2(P3_REG2_REG_29__SCAN_IN), .ZN(n7914) );
  NAND2_X1 U10330 ( .A1(n7422), .A2(P3_REG1_REG_29__SCAN_IN), .ZN(n7913) );
  NAND2_X1 U10331 ( .A1(n7454), .A2(P3_REG0_REG_29__SCAN_IN), .ZN(n7912) );
  INV_X1 U10332 ( .A(n11677), .ZN(n12744) );
  INV_X1 U10333 ( .A(n7915), .ZN(n12737) );
  INV_X1 U10334 ( .A(n12836), .ZN(n12826) );
  OR2_X1 U10335 ( .A1(n6482), .A2(n9783), .ZN(n7917) );
  AOI22_X1 U10336 ( .A1(n12744), .A2(n13100), .B1(n13098), .B2(n12746), .ZN(
        n7918) );
  NAND2_X1 U10337 ( .A1(n7921), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7922) );
  XNOR2_X1 U10338 ( .A(n10912), .B(P3_B_REG_SCAN_IN), .ZN(n7927) );
  NAND2_X1 U10339 ( .A1(n6514), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7924) );
  MUX2_X1 U10340 ( .A(P3_IR_REG_31__SCAN_IN), .B(n7924), .S(
        P3_IR_REG_25__SCAN_IN), .Z(n7926) );
  NAND2_X1 U10341 ( .A1(n7926), .A2(n7925), .ZN(n11105) );
  NAND2_X1 U10342 ( .A1(n7927), .A2(n11105), .ZN(n7929) );
  NAND2_X1 U10343 ( .A1(n7925), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7928) );
  INV_X1 U10344 ( .A(P3_D_REG_0__SCAN_IN), .ZN(n7930) );
  INV_X1 U10345 ( .A(n10912), .ZN(n7931) );
  INV_X1 U10346 ( .A(n13239), .ZN(n10023) );
  INV_X1 U10347 ( .A(P3_D_REG_1__SCAN_IN), .ZN(n9455) );
  NAND2_X1 U10348 ( .A1(n9525), .A2(n9455), .ZN(n7933) );
  INV_X1 U10349 ( .A(n7951), .ZN(n11203) );
  NAND2_X1 U10350 ( .A1(n11203), .A2(n11105), .ZN(n7932) );
  NAND2_X1 U10351 ( .A1(n7933), .A2(n7932), .ZN(n10024) );
  NOR2_X1 U10352 ( .A1(P3_D_REG_17__SCAN_IN), .A2(P3_D_REG_22__SCAN_IN), .ZN(
        n7937) );
  NOR4_X1 U10353 ( .A1(P3_D_REG_2__SCAN_IN), .A2(P3_D_REG_8__SCAN_IN), .A3(
        P3_D_REG_25__SCAN_IN), .A4(P3_D_REG_20__SCAN_IN), .ZN(n7936) );
  NOR4_X1 U10354 ( .A1(P3_D_REG_29__SCAN_IN), .A2(P3_D_REG_10__SCAN_IN), .A3(
        P3_D_REG_31__SCAN_IN), .A4(P3_D_REG_14__SCAN_IN), .ZN(n7935) );
  NOR4_X1 U10355 ( .A1(P3_D_REG_19__SCAN_IN), .A2(P3_D_REG_18__SCAN_IN), .A3(
        P3_D_REG_27__SCAN_IN), .A4(P3_D_REG_24__SCAN_IN), .ZN(n7934) );
  NAND4_X1 U10356 ( .A1(n7937), .A2(n7936), .A3(n7935), .A4(n7934), .ZN(n7943)
         );
  NOR4_X1 U10357 ( .A1(P3_D_REG_9__SCAN_IN), .A2(P3_D_REG_16__SCAN_IN), .A3(
        P3_D_REG_15__SCAN_IN), .A4(P3_D_REG_30__SCAN_IN), .ZN(n7941) );
  NOR4_X1 U10358 ( .A1(P3_D_REG_11__SCAN_IN), .A2(P3_D_REG_21__SCAN_IN), .A3(
        P3_D_REG_12__SCAN_IN), .A4(P3_D_REG_26__SCAN_IN), .ZN(n7940) );
  NOR4_X1 U10359 ( .A1(P3_D_REG_3__SCAN_IN), .A2(P3_D_REG_5__SCAN_IN), .A3(
        P3_D_REG_4__SCAN_IN), .A4(P3_D_REG_7__SCAN_IN), .ZN(n7939) );
  NOR4_X1 U10360 ( .A1(P3_D_REG_13__SCAN_IN), .A2(P3_D_REG_28__SCAN_IN), .A3(
        P3_D_REG_23__SCAN_IN), .A4(P3_D_REG_6__SCAN_IN), .ZN(n7938) );
  NAND4_X1 U10361 ( .A1(n7941), .A2(n7940), .A3(n7939), .A4(n7938), .ZN(n7942)
         );
  OAI21_X1 U10362 ( .B1(n7943), .B2(n7942), .A(n9525), .ZN(n7959) );
  NAND2_X1 U10363 ( .A1(n7958), .A2(n7959), .ZN(n9261) );
  INV_X1 U10364 ( .A(n9252), .ZN(n7946) );
  INV_X1 U10365 ( .A(n10024), .ZN(n9453) );
  NAND3_X1 U10366 ( .A1(n9453), .A2(n13239), .A3(n7959), .ZN(n9253) );
  OR2_X1 U10367 ( .A1(n12671), .A2(n9262), .ZN(n9993) );
  NAND2_X1 U10368 ( .A1(n7944), .A2(n12727), .ZN(n9254) );
  AND2_X1 U10369 ( .A1(n9993), .A2(n9254), .ZN(n7945) );
  OAI22_X1 U10370 ( .A1(n9261), .A2(n7946), .B1(n9253), .B2(n7945), .ZN(n7952)
         );
  NOR2_X1 U10371 ( .A1(n11105), .A2(n10912), .ZN(n7950) );
  INV_X1 U10372 ( .A(n9767), .ZN(n12736) );
  INV_X1 U10373 ( .A(n13234), .ZN(n13185) );
  NAND2_X1 U10374 ( .A1(n7954), .A2(n13185), .ZN(n7955) );
  OR2_X1 U10375 ( .A1(n12671), .A2(n12735), .ZN(n9250) );
  INV_X1 U10376 ( .A(n9250), .ZN(n7957) );
  NOR2_X1 U10377 ( .A1(n9767), .A2(n7957), .ZN(n7961) );
  INV_X1 U10378 ( .A(n7958), .ZN(n7960) );
  AND2_X1 U10379 ( .A1(n12671), .A2(n7962), .ZN(n10022) );
  NAND2_X1 U10380 ( .A1(n12739), .A2(n12857), .ZN(n7963) );
  OAI21_X1 U10381 ( .B1(n15170), .B2(n7964), .A(n7963), .ZN(n7965) );
  NAND2_X1 U10382 ( .A1(n7965), .A2(n9262), .ZN(n7966) );
  NAND3_X1 U10383 ( .A1(n7966), .A2(n12671), .A3(n10024), .ZN(n7967) );
  OAI21_X1 U10384 ( .B1(n13239), .B2(n10022), .A(n7967), .ZN(n7968) );
  INV_X1 U10385 ( .A(n7954), .ZN(n7970) );
  NOR2_X1 U10386 ( .A1(P2_IR_REG_6__SCAN_IN), .A2(P2_IR_REG_5__SCAN_IN), .ZN(
        n7974) );
  NOR2_X1 U10387 ( .A1(P2_IR_REG_11__SCAN_IN), .A2(P2_IR_REG_10__SCAN_IN), 
        .ZN(n7979) );
  NOR2_X1 U10388 ( .A1(P2_IR_REG_12__SCAN_IN), .A2(P2_IR_REG_16__SCAN_IN), 
        .ZN(n7978) );
  NOR2_X1 U10389 ( .A1(P2_IR_REG_15__SCAN_IN), .A2(P2_IR_REG_17__SCAN_IN), 
        .ZN(n7977) );
  NOR2_X1 U10390 ( .A1(P2_IR_REG_14__SCAN_IN), .A2(P2_IR_REG_13__SCAN_IN), 
        .ZN(n7976) );
  NOR2_X1 U10391 ( .A1(P2_IR_REG_22__SCAN_IN), .A2(P2_IR_REG_23__SCAN_IN), 
        .ZN(n7984) );
  NOR2_X1 U10392 ( .A1(P2_IR_REG_20__SCAN_IN), .A2(P2_IR_REG_21__SCAN_IN), 
        .ZN(n7983) );
  NOR2_X1 U10393 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_18__SCAN_IN), 
        .ZN(n7982) );
  NOR2_X1 U10394 ( .A1(P2_IR_REG_24__SCAN_IN), .A2(P2_IR_REG_25__SCAN_IN), 
        .ZN(n7981) );
  NAND2_X1 U10395 ( .A1(n8000), .A2(n7997), .ZN(n7988) );
  INV_X1 U10396 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n9646) );
  OR2_X1 U10397 ( .A1(n8050), .A2(n9646), .ZN(n7996) );
  INV_X1 U10398 ( .A(n11705), .ZN(n7992) );
  NAND2_X1 U10399 ( .A1(n8075), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n7995) );
  NAND2_X1 U10400 ( .A1(n8095), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n7994) );
  NAND2_X1 U10401 ( .A1(n8049), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n7993) );
  NAND4_X1 U10402 ( .A1(n7996), .A2(n7995), .A3(n7994), .A4(n7993), .ZN(n8838)
         );
  NAND2_X1 U10403 ( .A1(n8814), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7999) );
  INV_X1 U10404 ( .A(n8000), .ZN(n8001) );
  INV_X1 U10405 ( .A(n8005), .ZN(n8003) );
  NAND2_X1 U10406 ( .A1(n8003), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n8033) );
  NAND2_X1 U10407 ( .A1(n8005), .A2(n8004), .ZN(n8006) );
  AND2_X1 U10408 ( .A1(n8033), .A2(n8006), .ZN(n13824) );
  XNOR2_X2 U10409 ( .A(n8013), .B(n8012), .ZN(n10871) );
  NAND2_X1 U10410 ( .A1(n8838), .A2(n8014), .ZN(n8026) );
  INV_X1 U10411 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n8016) );
  XNOR2_X2 U10412 ( .A(n8017), .B(n8016), .ZN(n11649) );
  NAND2_X1 U10413 ( .A1(n8018), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8019) );
  INV_X1 U10414 ( .A(n8022), .ZN(n8020) );
  NAND2_X1 U10415 ( .A1(n8020), .A2(n10871), .ZN(n9920) );
  INV_X1 U10416 ( .A(n14938), .ZN(n10976) );
  INV_X2 U10417 ( .A(n8531), .ZN(n8117) );
  NAND2_X1 U10418 ( .A1(n8022), .A2(n9832), .ZN(n8025) );
  INV_X1 U10419 ( .A(n9832), .ZN(n8023) );
  NAND2_X1 U10420 ( .A1(n8075), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n8030) );
  NAND2_X1 U10421 ( .A1(n8095), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n8029) );
  INV_X1 U10422 ( .A(n8050), .ZN(n8074) );
  NAND2_X1 U10423 ( .A1(n8074), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n8028) );
  NAND2_X1 U10424 ( .A1(n8049), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n8027) );
  AND2_X1 U10425 ( .A1(n8020), .A2(n9832), .ZN(n8069) );
  INV_X1 U10426 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n9435) );
  XNOR2_X1 U10427 ( .A(n8063), .B(SI_1_), .ZN(n8062) );
  AND2_X1 U10428 ( .A1(P2_DATAO_REG_0__SCAN_IN), .A2(SI_0_), .ZN(n8032) );
  NAND2_X1 U10429 ( .A1(n11519), .A2(n8032), .ZN(n9359) );
  NAND2_X1 U10430 ( .A1(n8033), .A2(n9359), .ZN(n8061) );
  XNOR2_X1 U10431 ( .A(n8062), .B(n8061), .ZN(n9436) );
  NOR2_X1 U10432 ( .A1(n9434), .A2(n9437), .ZN(n8034) );
  NAND2_X1 U10433 ( .A1(n8056), .A2(n8034), .ZN(n8039) );
  INV_X1 U10434 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n8036) );
  NAND2_X1 U10435 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), 
        .ZN(n8035) );
  XNOR2_X1 U10436 ( .A(n8036), .B(n8035), .ZN(n9724) );
  OAI211_X1 U10437 ( .C1(n8066), .C2(n9436), .A(n8039), .B(n8038), .ZN(n8835)
         );
  NAND2_X1 U10438 ( .A1(n8069), .A2(n10012), .ZN(n8043) );
  NAND2_X1 U10439 ( .A1(n13396), .A2(n8531), .ZN(n8042) );
  NAND2_X1 U10440 ( .A1(n8043), .A2(n8042), .ZN(n8044) );
  OAI21_X1 U10441 ( .B1(n8046), .B2(n8045), .A(n8044), .ZN(n8048) );
  NAND2_X1 U10442 ( .A1(n8046), .A2(n8045), .ZN(n8047) );
  NAND2_X1 U10443 ( .A1(n8049), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n8055) );
  INV_X1 U10444 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n8051) );
  NAND2_X1 U10445 ( .A1(n8747), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n8053) );
  NAND2_X1 U10446 ( .A1(n8841), .A2(n8531), .ZN(n8071) );
  OR2_X1 U10447 ( .A1(n8057), .A2(n13808), .ZN(n8058) );
  INV_X1 U10448 ( .A(n14807), .ZN(n8059) );
  NAND2_X1 U10449 ( .A1(n8062), .A2(n8061), .ZN(n8064) );
  INV_X1 U10450 ( .A(n8105), .ZN(n8065) );
  XNOR2_X1 U10451 ( .A(n8065), .B(SI_2_), .ZN(n8081) );
  MUX2_X1 U10452 ( .A(n9461), .B(n9450), .S(n8084), .Z(n8107) );
  XNOR2_X1 U10453 ( .A(n8081), .B(n8107), .ZN(n9449) );
  NAND2_X1 U10454 ( .A1(n9449), .A2(n8667), .ZN(n8067) );
  NAND2_X2 U10455 ( .A1(n8068), .A2(n8067), .ZN(n9953) );
  INV_X1 U10456 ( .A(n8069), .ZN(n8581) );
  NAND2_X1 U10457 ( .A1(n9953), .A2(n8069), .ZN(n8070) );
  INV_X2 U10458 ( .A(n9953), .ZN(n10143) );
  NAND2_X1 U10459 ( .A1(n8841), .A2(n8069), .ZN(n8072) );
  NAND2_X1 U10460 ( .A1(n8074), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n8079) );
  NAND2_X1 U10461 ( .A1(n8746), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n8078) );
  OR2_X1 U10462 ( .A1(n8767), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n8077) );
  NAND2_X1 U10463 ( .A1(n8747), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n8076) );
  NAND2_X1 U10464 ( .A1(n13395), .A2(n8069), .ZN(n8091) );
  INV_X1 U10465 ( .A(n8107), .ZN(n8080) );
  NAND2_X1 U10466 ( .A1(n8081), .A2(n8080), .ZN(n8083) );
  NAND2_X1 U10467 ( .A1(n8105), .A2(SI_2_), .ZN(n8082) );
  NAND2_X1 U10468 ( .A1(n8083), .A2(n8082), .ZN(n8086) );
  MUX2_X1 U10469 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(P1_DATAO_REG_3__SCAN_IN), 
        .S(n8084), .Z(n8108) );
  XNOR2_X1 U10470 ( .A(n8108), .B(SI_3_), .ZN(n8085) );
  XNOR2_X1 U10471 ( .A(n8086), .B(n8085), .ZN(n9445) );
  NAND2_X1 U10472 ( .A1(n9445), .A2(n8667), .ZN(n8089) );
  INV_X1 U10473 ( .A(n8762), .ZN(n8180) );
  OR2_X1 U10474 ( .A1(n8101), .A2(n13808), .ZN(n8087) );
  XNOR2_X1 U10475 ( .A(n8087), .B(P2_IR_REG_3__SCAN_IN), .ZN(n9728) );
  INV_X4 U10476 ( .A(n8117), .ZN(n8736) );
  NAND2_X1 U10477 ( .A1(n13270), .A2(n8736), .ZN(n8090) );
  NAND2_X1 U10478 ( .A1(n8091), .A2(n8090), .ZN(n8093) );
  AOI22_X1 U10479 ( .A1(n13395), .A2(n8736), .B1(n13270), .B2(n8069), .ZN(
        n8092) );
  NAND2_X1 U10480 ( .A1(n8768), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n8099) );
  NAND2_X1 U10481 ( .A1(n8747), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n8098) );
  NAND2_X1 U10482 ( .A1(n8746), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n8097) );
  NAND2_X1 U10483 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n8129) );
  OAI21_X1 U10484 ( .B1(P2_REG3_REG_4__SCAN_IN), .B2(P2_REG3_REG_3__SCAN_IN), 
        .A(n8129), .ZN(n10296) );
  OR2_X1 U10485 ( .A1(n8767), .A2(n10296), .ZN(n8096) );
  NAND2_X1 U10486 ( .A1(n8833), .A2(n8531), .ZN(n8116) );
  INV_X1 U10487 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n8100) );
  NAND2_X1 U10488 ( .A1(n8101), .A2(n8100), .ZN(n8158) );
  NAND2_X1 U10489 ( .A1(n8158), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8139) );
  XNOR2_X1 U10490 ( .A(n8139), .B(n8156), .ZN(n13421) );
  INV_X1 U10491 ( .A(n8108), .ZN(n8103) );
  INV_X1 U10492 ( .A(SI_3_), .ZN(n8102) );
  NAND2_X1 U10493 ( .A1(n8103), .A2(n8102), .ZN(n8109) );
  INV_X1 U10494 ( .A(SI_2_), .ZN(n8106) );
  NAND2_X1 U10495 ( .A1(n8107), .A2(n8106), .ZN(n8104) );
  NAND3_X1 U10496 ( .A1(n8105), .A2(n8109), .A3(n8104), .ZN(n8112) );
  NOR2_X1 U10497 ( .A1(n8107), .A2(n8106), .ZN(n8110) );
  AOI22_X1 U10498 ( .A1(n8110), .A2(n8109), .B1(n8108), .B2(SI_3_), .ZN(n8111)
         );
  NAND2_X1 U10499 ( .A1(n8112), .A2(n8111), .ZN(n8136) );
  MUX2_X1 U10500 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(P1_DATAO_REG_4__SCAN_IN), 
        .S(n8084), .Z(n8137) );
  NAND2_X1 U10501 ( .A1(n9884), .A2(n8667), .ZN(n8114) );
  OR2_X1 U10502 ( .A1(n8762), .A2(n9452), .ZN(n8113) );
  OAI211_X1 U10503 ( .C1(n8056), .C2(n13421), .A(n8114), .B(n8113), .ZN(n10299) );
  INV_X1 U10504 ( .A(n8581), .ZN(n8738) );
  NAND2_X1 U10505 ( .A1(n10299), .A2(n8738), .ZN(n8115) );
  NAND2_X1 U10506 ( .A1(n8116), .A2(n8115), .ZN(n8122) );
  NAND2_X1 U10507 ( .A1(n8121), .A2(n8122), .ZN(n8120) );
  AOI22_X1 U10508 ( .A1(n8833), .A2(n8780), .B1(n10299), .B2(n8736), .ZN(n8118) );
  INV_X1 U10509 ( .A(n8118), .ZN(n8119) );
  NAND2_X1 U10510 ( .A1(n8120), .A2(n8119), .ZN(n8126) );
  NAND2_X1 U10511 ( .A1(n8124), .A2(n8123), .ZN(n8125) );
  NAND2_X1 U10512 ( .A1(n8126), .A2(n8125), .ZN(n8149) );
  NAND2_X1 U10513 ( .A1(n8747), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n8134) );
  NAND2_X1 U10514 ( .A1(n8768), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n8133) );
  INV_X1 U10515 ( .A(n8129), .ZN(n8127) );
  NAND2_X1 U10516 ( .A1(n8127), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n8164) );
  INV_X1 U10517 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n8128) );
  NAND2_X1 U10518 ( .A1(n8129), .A2(n8128), .ZN(n8130) );
  NAND2_X1 U10519 ( .A1(n8164), .A2(n8130), .ZN(n11712) );
  OR2_X1 U10520 ( .A1(n8767), .A2(n11712), .ZN(n8132) );
  NAND2_X1 U10521 ( .A1(n8746), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n8131) );
  NAND4_X1 U10522 ( .A1(n8134), .A2(n8133), .A3(n8132), .A4(n8131), .ZN(n13394) );
  NAND2_X1 U10523 ( .A1(n13394), .A2(n8738), .ZN(n8145) );
  NAND2_X1 U10524 ( .A1(n8137), .A2(SI_4_), .ZN(n8138) );
  MUX2_X1 U10525 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(P1_DATAO_REG_5__SCAN_IN), 
        .S(n8084), .Z(n8153) );
  XNOR2_X1 U10526 ( .A(n8153), .B(SI_5_), .ZN(n8150) );
  XNOR2_X1 U10527 ( .A(n8152), .B(n8150), .ZN(n10428) );
  NAND2_X1 U10528 ( .A1(n10428), .A2(n8667), .ZN(n8143) );
  INV_X1 U10529 ( .A(n8762), .ZN(n8465) );
  NAND2_X1 U10530 ( .A1(n8139), .A2(n8156), .ZN(n8140) );
  NAND2_X1 U10531 ( .A1(n8140), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8141) );
  XNOR2_X1 U10532 ( .A(n8141), .B(P2_IR_REG_5__SCAN_IN), .ZN(n14819) );
  AOI22_X1 U10533 ( .A1(n8465), .A2(P1_DATAO_REG_5__SCAN_IN), .B1(n9640), .B2(
        n14819), .ZN(n8142) );
  NAND2_X1 U10534 ( .A1(n8143), .A2(n8142), .ZN(n14947) );
  NAND2_X1 U10535 ( .A1(n14947), .A2(n8736), .ZN(n8144) );
  NAND2_X1 U10536 ( .A1(n8145), .A2(n8144), .ZN(n8148) );
  AOI22_X1 U10537 ( .A1(n13394), .A2(n8736), .B1(n14947), .B2(n8738), .ZN(
        n8146) );
  INV_X1 U10538 ( .A(n8150), .ZN(n8151) );
  NAND2_X1 U10539 ( .A1(n8153), .A2(SI_5_), .ZN(n8154) );
  MUX2_X1 U10540 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(P1_DATAO_REG_6__SCAN_IN), 
        .S(n9434), .Z(n8177) );
  XNOR2_X1 U10541 ( .A(n8177), .B(SI_6_), .ZN(n8174) );
  XNOR2_X1 U10542 ( .A(n8176), .B(n8174), .ZN(n10433) );
  NAND2_X1 U10543 ( .A1(n10433), .A2(n8667), .ZN(n8161) );
  INV_X1 U10544 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n8155) );
  NAND2_X1 U10545 ( .A1(n8156), .A2(n8155), .ZN(n8157) );
  NAND2_X1 U10546 ( .A1(n8181), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8159) );
  XNOR2_X1 U10547 ( .A(n8159), .B(P2_IR_REG_6__SCAN_IN), .ZN(n9733) );
  AOI22_X1 U10548 ( .A1(n8465), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n9640), .B2(
        n9733), .ZN(n8160) );
  NAND2_X1 U10549 ( .A1(n8161), .A2(n8160), .ZN(n10380) );
  NAND2_X1 U10550 ( .A1(n10380), .A2(n8738), .ZN(n8171) );
  NAND2_X1 U10551 ( .A1(n8768), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n8169) );
  NAND2_X1 U10552 ( .A1(n8747), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n8168) );
  INV_X1 U10553 ( .A(n8164), .ZN(n8162) );
  NAND2_X1 U10554 ( .A1(n8162), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n8193) );
  INV_X1 U10555 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n8163) );
  NAND2_X1 U10556 ( .A1(n8164), .A2(n8163), .ZN(n8165) );
  NAND2_X1 U10557 ( .A1(n8193), .A2(n8165), .ZN(n10385) );
  OR2_X1 U10558 ( .A1(n8767), .A2(n10385), .ZN(n8167) );
  NAND2_X1 U10559 ( .A1(n8746), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n8166) );
  NAND4_X1 U10560 ( .A1(n8169), .A2(n8168), .A3(n8167), .A4(n8166), .ZN(n13393) );
  NAND2_X1 U10561 ( .A1(n13393), .A2(n8736), .ZN(n8170) );
  NAND2_X1 U10562 ( .A1(n8171), .A2(n8170), .ZN(n8173) );
  AOI22_X1 U10563 ( .A1(n10380), .A2(n8531), .B1(n8780), .B2(n13393), .ZN(
        n8172) );
  INV_X1 U10564 ( .A(n8174), .ZN(n8175) );
  NAND2_X1 U10565 ( .A1(n8176), .A2(n8175), .ZN(n8179) );
  NAND2_X1 U10566 ( .A1(n8177), .A2(SI_6_), .ZN(n8178) );
  MUX2_X1 U10567 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(P1_DATAO_REG_7__SCAN_IN), 
        .S(n9434), .Z(n8210) );
  XNOR2_X1 U10568 ( .A(n8210), .B(SI_7_), .ZN(n8207) );
  XNOR2_X1 U10569 ( .A(n8209), .B(n8207), .ZN(n10448) );
  NAND2_X1 U10570 ( .A1(n10448), .A2(n8667), .ZN(n8190) );
  INV_X1 U10571 ( .A(n8181), .ZN(n8183) );
  INV_X1 U10572 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n8182) );
  NAND2_X1 U10573 ( .A1(n8183), .A2(n8182), .ZN(n8185) );
  NAND2_X1 U10574 ( .A1(n8185), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8184) );
  MUX2_X1 U10575 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8184), .S(
        P2_IR_REG_7__SCAN_IN), .Z(n8188) );
  INV_X1 U10576 ( .A(n8185), .ZN(n8187) );
  INV_X1 U10577 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n8186) );
  NAND2_X1 U10578 ( .A1(n8187), .A2(n8186), .ZN(n8234) );
  AOI22_X1 U10579 ( .A1(n8465), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n9640), .B2(
        n13444), .ZN(n8189) );
  NAND2_X1 U10580 ( .A1(n8190), .A2(n8189), .ZN(n10624) );
  NAND2_X1 U10581 ( .A1(n10624), .A2(n8736), .ZN(n8200) );
  NAND2_X1 U10582 ( .A1(n8768), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n8198) );
  NAND2_X1 U10583 ( .A1(n8747), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n8197) );
  INV_X1 U10584 ( .A(n8193), .ZN(n8191) );
  NAND2_X1 U10585 ( .A1(n8191), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n8216) );
  INV_X1 U10586 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n8192) );
  NAND2_X1 U10587 ( .A1(n8193), .A2(n8192), .ZN(n8194) );
  NAND2_X1 U10588 ( .A1(n8216), .A2(n8194), .ZN(n10600) );
  OR2_X1 U10589 ( .A1(n8767), .A2(n10600), .ZN(n8196) );
  NAND2_X1 U10590 ( .A1(n8746), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n8195) );
  NAND4_X1 U10591 ( .A1(n8198), .A2(n8197), .A3(n8196), .A4(n8195), .ZN(n13392) );
  NAND2_X1 U10592 ( .A1(n13392), .A2(n8738), .ZN(n8199) );
  NAND2_X1 U10593 ( .A1(n8200), .A2(n8199), .ZN(n8203) );
  NAND2_X1 U10594 ( .A1(n10624), .A2(n8738), .ZN(n8202) );
  NAND2_X1 U10595 ( .A1(n13392), .A2(n8736), .ZN(n8201) );
  INV_X1 U10596 ( .A(n8207), .ZN(n8208) );
  NAND2_X1 U10597 ( .A1(n8210), .A2(SI_7_), .ZN(n8211) );
  MUX2_X1 U10598 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(P1_DATAO_REG_8__SCAN_IN), 
        .S(n9434), .Z(n8232) );
  XNOR2_X1 U10599 ( .A(n8232), .B(SI_8_), .ZN(n8229) );
  XNOR2_X1 U10600 ( .A(n8231), .B(n8229), .ZN(n10461) );
  NAND2_X1 U10601 ( .A1(n10461), .A2(n8667), .ZN(n8214) );
  NAND2_X1 U10602 ( .A1(n8234), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8212) );
  XNOR2_X1 U10603 ( .A(n8212), .B(P2_IR_REG_8__SCAN_IN), .ZN(n9736) );
  AOI22_X1 U10604 ( .A1(n8465), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n9640), .B2(
        n9736), .ZN(n8213) );
  NAND2_X1 U10605 ( .A1(n8214), .A2(n8213), .ZN(n11771) );
  NAND2_X1 U10606 ( .A1(n11771), .A2(n8738), .ZN(n8223) );
  NAND2_X1 U10607 ( .A1(n8768), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n8221) );
  NAND2_X1 U10608 ( .A1(n8747), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n8220) );
  NAND2_X1 U10609 ( .A1(n8216), .A2(n8215), .ZN(n8217) );
  NAND2_X1 U10610 ( .A1(n8240), .A2(n8217), .ZN(n11767) );
  OR2_X1 U10611 ( .A1(n8767), .A2(n11767), .ZN(n8219) );
  NAND2_X1 U10612 ( .A1(n8746), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n8218) );
  NAND4_X1 U10613 ( .A1(n8221), .A2(n8220), .A3(n8219), .A4(n8218), .ZN(n13391) );
  NAND2_X1 U10614 ( .A1(n13391), .A2(n8736), .ZN(n8222) );
  NAND2_X1 U10615 ( .A1(n8223), .A2(n8222), .ZN(n8225) );
  AOI22_X1 U10616 ( .A1(n11771), .A2(n8531), .B1(n8780), .B2(n13391), .ZN(
        n8224) );
  AOI21_X1 U10617 ( .B1(n8226), .B2(n8225), .A(n8224), .ZN(n8228) );
  NOR2_X1 U10618 ( .A1(n8226), .A2(n8225), .ZN(n8227) );
  INV_X1 U10619 ( .A(n8229), .ZN(n8230) );
  NAND2_X1 U10620 ( .A1(n8232), .A2(SI_8_), .ZN(n8233) );
  MUX2_X1 U10621 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(P1_DATAO_REG_9__SCAN_IN), 
        .S(n9434), .Z(n8253) );
  XNOR2_X1 U10622 ( .A(n8253), .B(SI_9_), .ZN(n8250) );
  NAND2_X1 U10623 ( .A1(n10562), .A2(n8761), .ZN(n8237) );
  OAI21_X1 U10624 ( .B1(n8234), .B2(P2_IR_REG_8__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n8235) );
  XNOR2_X1 U10625 ( .A(n8235), .B(P2_IR_REG_9__SCAN_IN), .ZN(n14846) );
  AOI22_X1 U10626 ( .A1(n8465), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n9640), .B2(
        n14846), .ZN(n8236) );
  NAND2_X1 U10627 ( .A1(n10779), .A2(n8736), .ZN(n8247) );
  INV_X1 U10628 ( .A(n8747), .ZN(n8728) );
  INV_X1 U10629 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n10634) );
  OR2_X1 U10630 ( .A1(n8728), .A2(n10634), .ZN(n8245) );
  OR2_X1 U10631 ( .A1(n8750), .A2(n15013), .ZN(n8244) );
  NAND2_X1 U10632 ( .A1(n8746), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n8243) );
  INV_X1 U10633 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n8239) );
  NAND2_X1 U10634 ( .A1(n8240), .A2(n8239), .ZN(n8241) );
  NAND2_X1 U10635 ( .A1(n8259), .A2(n8241), .ZN(n10633) );
  OR2_X1 U10636 ( .A1(n8767), .A2(n10633), .ZN(n8242) );
  NAND4_X1 U10637 ( .A1(n8245), .A2(n8244), .A3(n8243), .A4(n8242), .ZN(n13390) );
  NAND2_X1 U10638 ( .A1(n13390), .A2(n8738), .ZN(n8246) );
  INV_X1 U10639 ( .A(n13390), .ZN(n11768) );
  NAND2_X1 U10640 ( .A1(n10779), .A2(n8738), .ZN(n8248) );
  OAI21_X1 U10641 ( .B1(n11768), .B2(n8117), .A(n8248), .ZN(n8249) );
  INV_X1 U10642 ( .A(n8250), .ZN(n8251) );
  MUX2_X1 U10643 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(P1_DATAO_REG_10__SCAN_IN), 
        .S(n9434), .Z(n8276) );
  XNOR2_X1 U10644 ( .A(n8276), .B(SI_10_), .ZN(n8273) );
  XNOR2_X1 U10645 ( .A(n8275), .B(n8273), .ZN(n10568) );
  NAND2_X1 U10646 ( .A1(n10568), .A2(n8667), .ZN(n8257) );
  OR2_X1 U10647 ( .A1(n8254), .A2(n13808), .ZN(n8255) );
  XNOR2_X1 U10648 ( .A(n8255), .B(P2_IR_REG_10__SCAN_IN), .ZN(n14863) );
  AOI22_X1 U10649 ( .A1(n8465), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n9640), 
        .B2(n14863), .ZN(n8256) );
  NAND2_X1 U10650 ( .A1(n14987), .A2(n8780), .ZN(n8266) );
  NAND2_X1 U10651 ( .A1(n8095), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n8264) );
  NAND2_X1 U10652 ( .A1(n8768), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n8263) );
  NAND2_X1 U10653 ( .A1(n8259), .A2(n8258), .ZN(n8260) );
  NAND2_X1 U10654 ( .A1(n8291), .A2(n8260), .ZN(n10800) );
  OR2_X1 U10655 ( .A1(n8767), .A2(n10800), .ZN(n8262) );
  NAND2_X1 U10656 ( .A1(n8746), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n8261) );
  NAND4_X1 U10657 ( .A1(n8264), .A2(n8263), .A3(n8262), .A4(n8261), .ZN(n13389) );
  NAND2_X1 U10658 ( .A1(n13389), .A2(n8736), .ZN(n8265) );
  NAND2_X1 U10659 ( .A1(n8266), .A2(n8265), .ZN(n8267) );
  NAND2_X1 U10660 ( .A1(n8268), .A2(n8267), .ZN(n8271) );
  AOI22_X1 U10661 ( .A1(n14987), .A2(n8531), .B1(n8780), .B2(n13389), .ZN(
        n8269) );
  NAND2_X1 U10662 ( .A1(n8271), .A2(n8270), .ZN(n8272) );
  INV_X1 U10663 ( .A(n8273), .ZN(n8274) );
  NAND2_X1 U10664 ( .A1(n8275), .A2(n8274), .ZN(n8278) );
  NAND2_X1 U10665 ( .A1(n8276), .A2(SI_10_), .ZN(n8277) );
  MUX2_X1 U10666 ( .A(n9574), .B(n9568), .S(n9434), .Z(n8280) );
  INV_X1 U10667 ( .A(n8280), .ZN(n8281) );
  NAND2_X1 U10668 ( .A1(n8281), .A2(SI_11_), .ZN(n8282) );
  NAND2_X1 U10669 ( .A1(n8328), .A2(n8282), .ZN(n8327) );
  XNOR2_X1 U10670 ( .A(n8325), .B(n8327), .ZN(n10939) );
  NAND2_X1 U10671 ( .A1(n10939), .A2(n8667), .ZN(n8288) );
  INV_X1 U10672 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n8283) );
  NAND2_X1 U10673 ( .A1(n8254), .A2(n8283), .ZN(n8285) );
  NAND2_X1 U10674 ( .A1(n8285), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8284) );
  MUX2_X1 U10675 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8284), .S(
        P2_IR_REG_11__SCAN_IN), .Z(n8286) );
  AOI22_X1 U10676 ( .A1(n8180), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n9640), 
        .B2(n9866), .ZN(n8287) );
  NAND2_X1 U10677 ( .A1(n10854), .A2(n8736), .ZN(n8298) );
  NAND2_X1 U10678 ( .A1(n8768), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n8296) );
  INV_X1 U10679 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n10788) );
  OR2_X1 U10680 ( .A1(n8728), .A2(n10788), .ZN(n8295) );
  INV_X1 U10681 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n8290) );
  NAND2_X1 U10682 ( .A1(n8291), .A2(n8290), .ZN(n8292) );
  NAND2_X1 U10683 ( .A1(n8313), .A2(n8292), .ZN(n10843) );
  OR2_X1 U10684 ( .A1(n8767), .A2(n10843), .ZN(n8294) );
  NAND2_X1 U10685 ( .A1(n8746), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n8293) );
  NAND4_X1 U10686 ( .A1(n8296), .A2(n8295), .A3(n8294), .A4(n8293), .ZN(n13388) );
  NAND2_X1 U10687 ( .A1(n13388), .A2(n8069), .ZN(n8297) );
  NAND2_X1 U10688 ( .A1(n8298), .A2(n8297), .ZN(n8304) );
  NAND2_X1 U10689 ( .A1(n10854), .A2(n8738), .ZN(n8300) );
  NAND2_X1 U10690 ( .A1(n13388), .A2(n8736), .ZN(n8299) );
  NAND2_X1 U10691 ( .A1(n8300), .A2(n8299), .ZN(n8301) );
  NAND2_X1 U10692 ( .A1(n8302), .A2(n8301), .ZN(n8308) );
  INV_X1 U10693 ( .A(n8303), .ZN(n8306) );
  INV_X1 U10694 ( .A(n8304), .ZN(n8305) );
  NAND2_X1 U10695 ( .A1(n8306), .A2(n8305), .ZN(n8307) );
  MUX2_X1 U10696 ( .A(n9613), .B(n9616), .S(n9434), .Z(n8330) );
  NAND2_X1 U10697 ( .A1(n10943), .A2(n8761), .ZN(n8311) );
  NAND2_X1 U10698 ( .A1(n8332), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8309) );
  XNOR2_X1 U10699 ( .A(n8309), .B(P2_IR_REG_12__SCAN_IN), .ZN(n10925) );
  AOI22_X1 U10700 ( .A1(n8465), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n9640), 
        .B2(n10925), .ZN(n8310) );
  NAND2_X1 U10701 ( .A1(n11730), .A2(n8738), .ZN(n8320) );
  INV_X1 U10702 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n9867) );
  OR2_X1 U10703 ( .A1(n8750), .A2(n9867), .ZN(n8318) );
  NAND2_X1 U10704 ( .A1(n8746), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n8317) );
  NAND2_X1 U10705 ( .A1(n8313), .A2(n8312), .ZN(n8314) );
  NAND2_X1 U10706 ( .A1(n8338), .A2(n8314), .ZN(n11719) );
  OR2_X1 U10707 ( .A1(n8767), .A2(n11719), .ZN(n8316) );
  OR2_X1 U10708 ( .A1(n8728), .A2(n10866), .ZN(n8315) );
  NAND4_X1 U10709 ( .A1(n8318), .A2(n8317), .A3(n8316), .A4(n8315), .ZN(n13387) );
  NAND2_X1 U10710 ( .A1(n13387), .A2(n8736), .ZN(n8319) );
  NAND2_X1 U10711 ( .A1(n8320), .A2(n8319), .ZN(n8323) );
  AOI22_X1 U10712 ( .A1(n11730), .A2(n8531), .B1(n8780), .B2(n13387), .ZN(
        n8321) );
  INV_X1 U10713 ( .A(n8321), .ZN(n8322) );
  INV_X1 U10714 ( .A(n8323), .ZN(n8324) );
  MUX2_X1 U10715 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(P1_DATAO_REG_13__SCAN_IN), 
        .S(n9438), .Z(n8346) );
  XNOR2_X1 U10716 ( .A(n8346), .B(n9566), .ZN(n8331) );
  XNOR2_X1 U10717 ( .A(n8347), .B(n8331), .ZN(n10981) );
  NAND2_X1 U10718 ( .A1(n10981), .A2(n8761), .ZN(n8336) );
  NOR2_X1 U10719 ( .A1(n8332), .A2(P2_IR_REG_12__SCAN_IN), .ZN(n8359) );
  INV_X1 U10720 ( .A(n8359), .ZN(n8333) );
  NAND2_X1 U10721 ( .A1(n8333), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8334) );
  XNOR2_X1 U10722 ( .A(n8334), .B(P2_IR_REG_13__SCAN_IN), .ZN(n14875) );
  AOI22_X1 U10723 ( .A1(n8180), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n9640), 
        .B2(n14875), .ZN(n8335) );
  NAND2_X1 U10724 ( .A1(n11281), .A2(n8736), .ZN(n8345) );
  NAND2_X1 U10725 ( .A1(n8768), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n8343) );
  NAND2_X1 U10726 ( .A1(n8747), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n8342) );
  NAND2_X1 U10727 ( .A1(n8338), .A2(n8337), .ZN(n8339) );
  NAND2_X1 U10728 ( .A1(n8417), .A2(n8339), .ZN(n11097) );
  OR2_X1 U10729 ( .A1(n8767), .A2(n11097), .ZN(n8341) );
  NAND2_X1 U10730 ( .A1(n8746), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n8340) );
  NAND4_X1 U10731 ( .A1(n8343), .A2(n8342), .A3(n8341), .A4(n8340), .ZN(n13386) );
  NAND2_X1 U10732 ( .A1(n13386), .A2(n8780), .ZN(n8344) );
  NAND2_X1 U10733 ( .A1(n8345), .A2(n8344), .ZN(n8430) );
  NAND2_X1 U10734 ( .A1(n8348), .A2(SI_14_), .ZN(n8349) );
  MUX2_X1 U10735 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(P1_DATAO_REG_14__SCAN_IN), 
        .S(n9434), .Z(n8409) );
  MUX2_X1 U10736 ( .A(n10132), .B(n10134), .S(n9434), .Z(n8350) );
  INV_X1 U10737 ( .A(n8350), .ZN(n8351) );
  NAND2_X1 U10738 ( .A1(n8351), .A2(SI_15_), .ZN(n8352) );
  NAND2_X1 U10739 ( .A1(n8390), .A2(n8389), .ZN(n8354) );
  NAND2_X1 U10740 ( .A1(n8354), .A2(n8353), .ZN(n8373) );
  MUX2_X1 U10741 ( .A(n10210), .B(n10212), .S(n9438), .Z(n8355) );
  NAND2_X1 U10742 ( .A1(n8355), .A2(n9679), .ZN(n8356) );
  MUX2_X1 U10743 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(P1_DATAO_REG_17__SCAN_IN), 
        .S(n9438), .Z(n8460) );
  XNOR2_X1 U10744 ( .A(n8460), .B(n9764), .ZN(n8357) );
  XNOR2_X1 U10745 ( .A(n8461), .B(n8357), .ZN(n11240) );
  NAND2_X1 U10746 ( .A1(n11240), .A2(n8761), .ZN(n8364) );
  INV_X1 U10747 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n8358) );
  NAND2_X1 U10748 ( .A1(n8359), .A2(n8358), .ZN(n8411) );
  INV_X1 U10749 ( .A(n8391), .ZN(n8361) );
  INV_X1 U10750 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n8360) );
  NAND2_X1 U10751 ( .A1(n8361), .A2(n8360), .ZN(n8393) );
  OAI21_X1 U10752 ( .B1(n8393), .B2(P2_IR_REG_16__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n8362) );
  XNOR2_X1 U10753 ( .A(n8362), .B(P2_IR_REG_17__SCAN_IN), .ZN(n13468) );
  AOI22_X1 U10754 ( .A1(n13468), .A2(n9640), .B1(n8465), .B2(
        P1_DATAO_REG_17__SCAN_IN), .ZN(n8363) );
  INV_X1 U10755 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n8369) );
  INV_X1 U10756 ( .A(n8365), .ZN(n8381) );
  INV_X1 U10757 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n13323) );
  NAND2_X1 U10758 ( .A1(n8381), .A2(n13323), .ZN(n8366) );
  NAND2_X1 U10759 ( .A1(n8468), .A2(n8366), .ZN(n13324) );
  OR2_X1 U10760 ( .A1(n13324), .A2(n8767), .ZN(n8368) );
  AOI22_X1 U10761 ( .A1(n8768), .A2(P2_REG1_REG_17__SCAN_IN), .B1(n8747), .B2(
        P2_REG2_REG_17__SCAN_IN), .ZN(n8367) );
  OAI211_X1 U10762 ( .C1(n8771), .C2(n8369), .A(n8368), .B(n8367), .ZN(n13382)
         );
  AND2_X1 U10763 ( .A1(n13382), .A2(n8780), .ZN(n8370) );
  AOI21_X1 U10764 ( .B1(n13767), .B2(n8736), .A(n8370), .ZN(n8445) );
  NAND2_X1 U10765 ( .A1(n13767), .A2(n8780), .ZN(n8372) );
  NAND2_X1 U10766 ( .A1(n13382), .A2(n8736), .ZN(n8371) );
  NAND2_X1 U10767 ( .A1(n8372), .A2(n8371), .ZN(n8443) );
  NAND2_X1 U10768 ( .A1(n8445), .A2(n8443), .ZN(n8388) );
  XNOR2_X1 U10769 ( .A(n8373), .B(n8374), .ZN(n11180) );
  NAND2_X1 U10770 ( .A1(n11180), .A2(n8761), .ZN(n8377) );
  NAND2_X1 U10771 ( .A1(n8393), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8375) );
  XNOR2_X1 U10772 ( .A(n8375), .B(P2_IR_REG_16__SCAN_IN), .ZN(n13467) );
  AOI22_X1 U10773 ( .A1(n13467), .A2(n9640), .B1(n8465), .B2(
        P1_DATAO_REG_16__SCAN_IN), .ZN(n8376) );
  INV_X1 U10774 ( .A(n8378), .ZN(n8400) );
  INV_X1 U10775 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n8379) );
  NAND2_X1 U10776 ( .A1(n8400), .A2(n8379), .ZN(n8380) );
  NAND2_X1 U10777 ( .A1(n8381), .A2(n8380), .ZN(n13317) );
  AOI22_X1 U10778 ( .A1(n8768), .A2(P2_REG1_REG_16__SCAN_IN), .B1(n8747), .B2(
        P2_REG2_REG_16__SCAN_IN), .ZN(n8383) );
  NAND2_X1 U10779 ( .A1(n8746), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n8382) );
  OAI211_X1 U10780 ( .C1(n13317), .C2(n8767), .A(n8383), .B(n8382), .ZN(n13383) );
  AND2_X1 U10781 ( .A1(n13383), .A2(n8738), .ZN(n8384) );
  AOI21_X1 U10782 ( .B1(n13772), .B2(n8736), .A(n8384), .ZN(n8439) );
  NAND2_X1 U10783 ( .A1(n13772), .A2(n8780), .ZN(n8386) );
  NAND2_X1 U10784 ( .A1(n13383), .A2(n8736), .ZN(n8385) );
  NAND2_X1 U10785 ( .A1(n8386), .A2(n8385), .ZN(n8438) );
  NAND2_X1 U10786 ( .A1(n8439), .A2(n8438), .ZN(n8387) );
  NAND2_X1 U10787 ( .A1(n8388), .A2(n8387), .ZN(n8452) );
  XNOR2_X1 U10788 ( .A(n8390), .B(n8389), .ZN(n11163) );
  NAND2_X1 U10789 ( .A1(n11163), .A2(n8761), .ZN(n8397) );
  NAND2_X1 U10790 ( .A1(n8391), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8392) );
  MUX2_X1 U10791 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8392), .S(
        P2_IR_REG_15__SCAN_IN), .Z(n8394) );
  NAND2_X1 U10792 ( .A1(n8394), .A2(n8393), .ZN(n14904) );
  OAI22_X1 U10793 ( .A1(n8762), .A2(n10134), .B1(n14904), .B2(n8056), .ZN(
        n8395) );
  INV_X1 U10794 ( .A(n8395), .ZN(n8396) );
  INV_X1 U10795 ( .A(n8398), .ZN(n8419) );
  INV_X1 U10796 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n11328) );
  NAND2_X1 U10797 ( .A1(n8419), .A2(n11328), .ZN(n8399) );
  NAND2_X1 U10798 ( .A1(n8400), .A2(n8399), .ZN(n11368) );
  OR2_X1 U10799 ( .A1(n11368), .A2(n8767), .ZN(n8404) );
  INV_X1 U10800 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n14899) );
  OR2_X1 U10801 ( .A1(n8728), .A2(n14899), .ZN(n8403) );
  INV_X1 U10802 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n14895) );
  OR2_X1 U10803 ( .A1(n8750), .A2(n14895), .ZN(n8402) );
  NAND2_X1 U10804 ( .A1(n8746), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n8401) );
  NAND4_X1 U10805 ( .A1(n8404), .A2(n8403), .A3(n8402), .A4(n8401), .ZN(n13384) );
  AND2_X1 U10806 ( .A1(n13384), .A2(n8780), .ZN(n8405) );
  AOI21_X1 U10807 ( .B1(n13780), .B2(n8736), .A(n8405), .ZN(n8451) );
  NAND2_X1 U10808 ( .A1(n13780), .A2(n8738), .ZN(n8407) );
  NAND2_X1 U10809 ( .A1(n13384), .A2(n8736), .ZN(n8406) );
  NAND2_X1 U10810 ( .A1(n8407), .A2(n8406), .ZN(n8450) );
  AND2_X1 U10811 ( .A1(n8451), .A2(n8450), .ZN(n8408) );
  NOR2_X1 U10812 ( .A1(n8452), .A2(n8408), .ZN(n8433) );
  XNOR2_X1 U10813 ( .A(n8410), .B(n8409), .ZN(n10986) );
  NAND2_X1 U10814 ( .A1(n10986), .A2(n8761), .ZN(n8414) );
  NAND2_X1 U10815 ( .A1(n8411), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8412) );
  XNOR2_X1 U10816 ( .A(n8412), .B(P2_IR_REG_14__SCAN_IN), .ZN(n14889) );
  AOI22_X1 U10817 ( .A1(n8465), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n9640), 
        .B2(n14889), .ZN(n8413) );
  NAND2_X1 U10818 ( .A1(n8747), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n8423) );
  INV_X1 U10819 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n8415) );
  OR2_X1 U10820 ( .A1(n8750), .A2(n8415), .ZN(n8422) );
  NAND2_X1 U10821 ( .A1(n8417), .A2(n8416), .ZN(n8418) );
  NAND2_X1 U10822 ( .A1(n8419), .A2(n8418), .ZN(n11217) );
  OR2_X1 U10823 ( .A1(n8767), .A2(n11217), .ZN(n8421) );
  NAND2_X1 U10824 ( .A1(n8746), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n8420) );
  NAND4_X1 U10825 ( .A1(n8423), .A2(n8422), .A3(n8421), .A4(n8420), .ZN(n13385) );
  AND2_X1 U10826 ( .A1(n13385), .A2(n8780), .ZN(n8424) );
  AOI21_X1 U10827 ( .B1(n13784), .B2(n8736), .A(n8424), .ZN(n8435) );
  NAND2_X1 U10828 ( .A1(n13784), .A2(n8780), .ZN(n8426) );
  NAND2_X1 U10829 ( .A1(n13385), .A2(n8736), .ZN(n8425) );
  NAND2_X1 U10830 ( .A1(n8426), .A2(n8425), .ZN(n8434) );
  NAND2_X1 U10831 ( .A1(n8435), .A2(n8434), .ZN(n8427) );
  OAI211_X1 U10832 ( .C1(n8431), .C2(n8430), .A(n8433), .B(n8427), .ZN(n8428)
         );
  AOI22_X1 U10833 ( .A1(n11281), .A2(n8780), .B1(n13386), .B2(n8736), .ZN(
        n8429) );
  AOI21_X1 U10834 ( .B1(n8431), .B2(n8430), .A(n8429), .ZN(n8432) );
  INV_X1 U10835 ( .A(n8433), .ZN(n8456) );
  INV_X1 U10836 ( .A(n8434), .ZN(n8437) );
  INV_X1 U10837 ( .A(n8435), .ZN(n8436) );
  NAND2_X1 U10838 ( .A1(n8437), .A2(n8436), .ZN(n8455) );
  INV_X1 U10839 ( .A(n8438), .ZN(n8441) );
  INV_X1 U10840 ( .A(n8439), .ZN(n8440) );
  NAND2_X1 U10841 ( .A1(n8441), .A2(n8440), .ZN(n8444) );
  INV_X1 U10842 ( .A(n13767), .ZN(n8442) );
  INV_X1 U10843 ( .A(n13382), .ZN(n13316) );
  NAND3_X1 U10844 ( .A1(n8444), .A2(n8442), .A3(n13316), .ZN(n8449) );
  INV_X1 U10845 ( .A(n8443), .ZN(n8448) );
  INV_X1 U10846 ( .A(n8444), .ZN(n8447) );
  INV_X1 U10847 ( .A(n8445), .ZN(n8446) );
  AOI22_X1 U10848 ( .A1(n8449), .A2(n8448), .B1(n8447), .B2(n8446), .ZN(n8454)
         );
  OR3_X1 U10849 ( .A1(n8452), .A2(n8451), .A3(n8450), .ZN(n8453) );
  OAI211_X1 U10850 ( .C1(n8456), .C2(n8455), .A(n8454), .B(n8453), .ZN(n8457)
         );
  INV_X1 U10851 ( .A(n8457), .ZN(n8458) );
  NAND2_X1 U10852 ( .A1(n8459), .A2(n8458), .ZN(n8479) );
  XNOR2_X1 U10853 ( .A(n8511), .B(SI_18_), .ZN(n8482) );
  MUX2_X1 U10854 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(P1_DATAO_REG_18__SCAN_IN), 
        .S(n9438), .Z(n8504) );
  XNOR2_X1 U10855 ( .A(n8482), .B(n8504), .ZN(n11373) );
  NAND2_X1 U10856 ( .A1(n11373), .A2(n8761), .ZN(n8467) );
  NAND2_X1 U10857 ( .A1(n8009), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8463) );
  INV_X1 U10858 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n8462) );
  XNOR2_X1 U10859 ( .A(n8463), .B(n8462), .ZN(n13479) );
  INV_X1 U10860 ( .A(n13479), .ZN(n8464) );
  AOI22_X1 U10861 ( .A1(n8465), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n9640), 
        .B2(n8464), .ZN(n8466) );
  NAND2_X1 U10862 ( .A1(n8468), .A2(n13364), .ZN(n8469) );
  AND2_X1 U10863 ( .A1(n8491), .A2(n8469), .ZN(n13686) );
  NAND2_X1 U10864 ( .A1(n13686), .A2(n8694), .ZN(n8474) );
  INV_X1 U10865 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n13469) );
  NAND2_X1 U10866 ( .A1(n8747), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n8471) );
  NAND2_X1 U10867 ( .A1(n8746), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n8470) );
  OAI211_X1 U10868 ( .C1(n8750), .C2(n13469), .A(n8471), .B(n8470), .ZN(n8472)
         );
  INV_X1 U10869 ( .A(n8472), .ZN(n8473) );
  NAND2_X1 U10870 ( .A1(n8474), .A2(n8473), .ZN(n13381) );
  AND2_X1 U10871 ( .A1(n13381), .A2(n8736), .ZN(n8475) );
  AOI21_X1 U10872 ( .B1(n13763), .B2(n8780), .A(n8475), .ZN(n8478) );
  INV_X1 U10873 ( .A(n13381), .ZN(n13656) );
  NAND2_X1 U10874 ( .A1(n13763), .A2(n8736), .ZN(n8476) );
  OAI21_X1 U10875 ( .B1(n13656), .B2(n8581), .A(n8476), .ZN(n8477) );
  NAND2_X1 U10876 ( .A1(n8479), .A2(n8478), .ZN(n8480) );
  NAND2_X1 U10877 ( .A1(n8511), .A2(SI_18_), .ZN(n8483) );
  MUX2_X1 U10878 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(P1_DATAO_REG_19__SCAN_IN), 
        .S(n9434), .Z(n8484) );
  NAND2_X1 U10879 ( .A1(n8484), .A2(SI_19_), .ZN(n8507) );
  INV_X1 U10880 ( .A(n8484), .ZN(n8485) );
  NAND2_X1 U10881 ( .A1(n8485), .A2(n9992), .ZN(n8505) );
  NAND2_X1 U10882 ( .A1(n8507), .A2(n8505), .ZN(n8486) );
  NAND2_X1 U10883 ( .A1(n11428), .A2(n8667), .ZN(n8488) );
  AOI22_X1 U10884 ( .A1(n8180), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n13490), 
        .B2(n9640), .ZN(n8487) );
  NAND2_X1 U10885 ( .A1(n13757), .A2(n8736), .ZN(n8500) );
  INV_X1 U10886 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n8490) );
  NAND2_X1 U10887 ( .A1(n8491), .A2(n8490), .ZN(n8492) );
  NAND2_X1 U10888 ( .A1(n8518), .A2(n8492), .ZN(n13279) );
  OR2_X1 U10889 ( .A1(n13279), .A2(n8767), .ZN(n8498) );
  INV_X1 U10890 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n8495) );
  NAND2_X1 U10891 ( .A1(n8747), .A2(P2_REG2_REG_19__SCAN_IN), .ZN(n8494) );
  NAND2_X1 U10892 ( .A1(n8746), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n8493) );
  OAI211_X1 U10893 ( .C1(n8750), .C2(n8495), .A(n8494), .B(n8493), .ZN(n8496)
         );
  INV_X1 U10894 ( .A(n8496), .ZN(n8497) );
  NAND2_X1 U10895 ( .A1(n13641), .A2(n8780), .ZN(n8499) );
  AOI22_X1 U10896 ( .A1(n13757), .A2(n8780), .B1(n13641), .B2(n8736), .ZN(
        n8501) );
  INV_X1 U10897 ( .A(n8501), .ZN(n8502) );
  INV_X1 U10898 ( .A(n8504), .ZN(n8503) );
  OAI21_X1 U10899 ( .B1(n8503), .B2(n9883), .A(n8507), .ZN(n8510) );
  NOR2_X1 U10900 ( .A1(n8504), .A2(SI_18_), .ZN(n8508) );
  INV_X1 U10901 ( .A(n8505), .ZN(n8506) );
  AOI21_X1 U10902 ( .B1(n8508), .B2(n8507), .A(n8506), .ZN(n8509) );
  INV_X1 U10903 ( .A(n8512), .ZN(n8513) );
  NAND2_X1 U10904 ( .A1(n8512), .A2(n10287), .ZN(n8537) );
  NAND2_X1 U10905 ( .A1(n8539), .A2(n8537), .ZN(n8514) );
  MUX2_X1 U10906 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(P1_DATAO_REG_20__SCAN_IN), 
        .S(n9438), .Z(n8538) );
  NAND2_X1 U10907 ( .A1(n11469), .A2(n8761), .ZN(n8516) );
  INV_X1 U10908 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n10872) );
  OR2_X1 U10909 ( .A1(n8762), .A2(n10872), .ZN(n8515) );
  NAND2_X1 U10910 ( .A1(n13752), .A2(n8780), .ZN(n8527) );
  INV_X1 U10911 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n8517) );
  NAND2_X1 U10912 ( .A1(n8518), .A2(n8517), .ZN(n8519) );
  AND2_X1 U10913 ( .A1(n8551), .A2(n8519), .ZN(n13632) );
  NAND2_X1 U10914 ( .A1(n13632), .A2(n8694), .ZN(n8525) );
  INV_X1 U10915 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n8522) );
  NAND2_X1 U10916 ( .A1(n8768), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n8521) );
  NAND2_X1 U10917 ( .A1(n8747), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n8520) );
  OAI211_X1 U10918 ( .C1(n8771), .C2(n8522), .A(n8521), .B(n8520), .ZN(n8523)
         );
  INV_X1 U10919 ( .A(n8523), .ZN(n8524) );
  NAND2_X1 U10920 ( .A1(n8525), .A2(n8524), .ZN(n13624) );
  NAND2_X1 U10921 ( .A1(n13624), .A2(n8736), .ZN(n8526) );
  NAND2_X1 U10922 ( .A1(n8527), .A2(n8526), .ZN(n8529) );
  INV_X1 U10923 ( .A(n8528), .ZN(n8536) );
  NAND2_X1 U10924 ( .A1(n8530), .A2(n8529), .ZN(n8534) );
  AOI22_X1 U10925 ( .A1(n13752), .A2(n8531), .B1(n8780), .B2(n13624), .ZN(
        n8532) );
  NAND2_X1 U10926 ( .A1(n8534), .A2(n8533), .ZN(n8535) );
  NAND2_X1 U10927 ( .A1(n8538), .A2(n8537), .ZN(n8540) );
  INV_X1 U10928 ( .A(n8545), .ZN(n8542) );
  MUX2_X1 U10929 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(P1_DATAO_REG_21__SCAN_IN), 
        .S(n9434), .Z(n8541) );
  OAI21_X1 U10930 ( .B1(SI_21_), .B2(n8541), .A(n8563), .ZN(n8543) );
  NAND2_X1 U10931 ( .A1(n8542), .A2(n8543), .ZN(n8546) );
  INV_X1 U10932 ( .A(n8543), .ZN(n8544) );
  AND2_X1 U10933 ( .A1(n8546), .A2(n8564), .ZN(n11514) );
  NAND2_X1 U10934 ( .A1(n11514), .A2(n8761), .ZN(n8548) );
  OR2_X1 U10935 ( .A1(n8762), .A2(n10977), .ZN(n8547) );
  NAND2_X1 U10936 ( .A1(n13747), .A2(n8736), .ZN(n8560) );
  INV_X1 U10937 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n8550) );
  NAND2_X1 U10938 ( .A1(n8551), .A2(n8550), .ZN(n8552) );
  NAND2_X1 U10939 ( .A1(n8570), .A2(n8552), .ZN(n13618) );
  OR2_X1 U10940 ( .A1(n13618), .A2(n8767), .ZN(n8558) );
  INV_X1 U10941 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n8555) );
  NAND2_X1 U10942 ( .A1(n8747), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n8554) );
  NAND2_X1 U10943 ( .A1(n8768), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n8553) );
  OAI211_X1 U10944 ( .C1(n8555), .C2(n8771), .A(n8554), .B(n8553), .ZN(n8556)
         );
  INV_X1 U10945 ( .A(n8556), .ZN(n8557) );
  NAND2_X1 U10946 ( .A1(n13643), .A2(n8738), .ZN(n8559) );
  INV_X1 U10947 ( .A(n13643), .ZN(n13597) );
  NAND2_X1 U10948 ( .A1(n13747), .A2(n8780), .ZN(n8561) );
  OAI21_X1 U10949 ( .B1(n13597), .B2(n8117), .A(n8561), .ZN(n8562) );
  XNOR2_X2 U10950 ( .A(n8592), .B(n8565), .ZN(n8591) );
  MUX2_X1 U10951 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(P1_DATAO_REG_22__SCAN_IN), 
        .S(n9438), .Z(n8590) );
  INV_X1 U10952 ( .A(n8590), .ZN(n8566) );
  XNOR2_X1 U10953 ( .A(n8591), .B(n8566), .ZN(n11648) );
  NAND2_X1 U10954 ( .A1(n11648), .A2(n8761), .ZN(n8568) );
  OR2_X1 U10955 ( .A1(n8762), .A2(n11651), .ZN(n8567) );
  NAND2_X1 U10956 ( .A1(n13740), .A2(n8780), .ZN(n8579) );
  INV_X1 U10957 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n13350) );
  NAND2_X1 U10958 ( .A1(n8570), .A2(n13350), .ZN(n8571) );
  NAND2_X1 U10959 ( .A1(n8598), .A2(n8571), .ZN(n13608) );
  OR2_X1 U10960 ( .A1(n13608), .A2(n8767), .ZN(n8577) );
  INV_X1 U10961 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n8574) );
  NAND2_X1 U10962 ( .A1(n8747), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n8573) );
  NAND2_X1 U10963 ( .A1(n8768), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n8572) );
  OAI211_X1 U10964 ( .C1(n8574), .C2(n8771), .A(n8573), .B(n8572), .ZN(n8575)
         );
  INV_X1 U10965 ( .A(n8575), .ZN(n8576) );
  NAND2_X1 U10966 ( .A1(n13625), .A2(n8736), .ZN(n8578) );
  NAND2_X1 U10967 ( .A1(n8579), .A2(n8578), .ZN(n8585) );
  INV_X1 U10968 ( .A(n13625), .ZN(n13292) );
  NAND2_X1 U10969 ( .A1(n13740), .A2(n8736), .ZN(n8580) );
  OAI21_X1 U10970 ( .B1(n13292), .B2(n8581), .A(n8580), .ZN(n8582) );
  NAND2_X1 U10971 ( .A1(n8583), .A2(n8582), .ZN(n8589) );
  INV_X1 U10972 ( .A(n8584), .ZN(n8587) );
  INV_X1 U10973 ( .A(n8585), .ZN(n8586) );
  NAND2_X1 U10974 ( .A1(n8587), .A2(n8586), .ZN(n8588) );
  NAND2_X1 U10975 ( .A1(n8592), .A2(SI_22_), .ZN(n8593) );
  MUX2_X1 U10976 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(P1_DATAO_REG_23__SCAN_IN), 
        .S(n9438), .Z(n8613) );
  XNOR2_X1 U10977 ( .A(n8613), .B(SI_23_), .ZN(n8610) );
  XNOR2_X1 U10978 ( .A(n8612), .B(n8610), .ZN(n11532) );
  NAND2_X1 U10979 ( .A1(n11532), .A2(n8761), .ZN(n8596) );
  OR2_X1 U10980 ( .A1(n8762), .A2(n11269), .ZN(n8595) );
  NAND2_X1 U10981 ( .A1(n13735), .A2(n8736), .ZN(n8607) );
  INV_X1 U10982 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n8597) );
  NAND2_X1 U10983 ( .A1(n8598), .A2(n8597), .ZN(n8599) );
  NAND2_X1 U10984 ( .A1(n8618), .A2(n8599), .ZN(n13586) );
  OR2_X1 U10985 ( .A1(n13586), .A2(n8767), .ZN(n8605) );
  INV_X1 U10986 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n8602) );
  NAND2_X1 U10987 ( .A1(n8768), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n8601) );
  NAND2_X1 U10988 ( .A1(n8747), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n8600) );
  OAI211_X1 U10989 ( .C1(n8771), .C2(n8602), .A(n8601), .B(n8600), .ZN(n8603)
         );
  INV_X1 U10990 ( .A(n8603), .ZN(n8604) );
  NAND2_X1 U10991 ( .A1(n8605), .A2(n8604), .ZN(n13380) );
  NAND2_X1 U10992 ( .A1(n13380), .A2(n8780), .ZN(n8606) );
  NAND2_X1 U10993 ( .A1(n13735), .A2(n8738), .ZN(n8609) );
  NAND2_X1 U10994 ( .A1(n13380), .A2(n8736), .ZN(n8608) );
  NAND2_X1 U10995 ( .A1(n8612), .A2(n8611), .ZN(n8615) );
  NAND2_X1 U10996 ( .A1(n8613), .A2(SI_23_), .ZN(n8614) );
  NAND2_X2 U10997 ( .A1(n8615), .A2(n8614), .ZN(n8659) );
  MUX2_X1 U10998 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(P1_DATAO_REG_24__SCAN_IN), 
        .S(n9438), .Z(n8660) );
  NAND2_X1 U10999 ( .A1(n11543), .A2(n8761), .ZN(n8617) );
  OR2_X1 U11000 ( .A1(n8762), .A2(n11396), .ZN(n8616) );
  NAND2_X1 U11001 ( .A1(n13729), .A2(n8780), .ZN(n8627) );
  INV_X1 U11002 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n13340) );
  NAND2_X1 U11003 ( .A1(n8618), .A2(n13340), .ZN(n8619) );
  AND2_X1 U11004 ( .A1(n8643), .A2(n8619), .ZN(n13571) );
  NAND2_X1 U11005 ( .A1(n13571), .A2(n8694), .ZN(n8625) );
  INV_X1 U11006 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n8622) );
  NAND2_X1 U11007 ( .A1(n8095), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n8621) );
  NAND2_X1 U11008 ( .A1(n8768), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n8620) );
  OAI211_X1 U11009 ( .C1(n8622), .C2(n8771), .A(n8621), .B(n8620), .ZN(n8623)
         );
  INV_X1 U11010 ( .A(n8623), .ZN(n8624) );
  NAND2_X1 U11011 ( .A1(n8625), .A2(n8624), .ZN(n13379) );
  NAND2_X1 U11012 ( .A1(n13379), .A2(n8736), .ZN(n8626) );
  NAND2_X1 U11013 ( .A1(n8627), .A2(n8626), .ZN(n8631) );
  NAND2_X1 U11014 ( .A1(n8632), .A2(n8631), .ZN(n8630) );
  AOI22_X1 U11015 ( .A1(n13729), .A2(n8736), .B1(n8780), .B2(n13379), .ZN(
        n8628) );
  INV_X1 U11016 ( .A(n8628), .ZN(n8629) );
  NAND2_X1 U11017 ( .A1(n8630), .A2(n8629), .ZN(n8633) );
  INV_X1 U11018 ( .A(n8660), .ZN(n8657) );
  INV_X1 U11019 ( .A(n8659), .ZN(n8634) );
  OAI22_X1 U11020 ( .A1(n8635), .A2(n8657), .B1(n8634), .B2(n10910), .ZN(n8639) );
  MUX2_X1 U11021 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(P1_DATAO_REG_25__SCAN_IN), 
        .S(n9434), .Z(n8636) );
  NAND2_X1 U11022 ( .A1(n8636), .A2(SI_25_), .ZN(n8663) );
  INV_X1 U11023 ( .A(n8636), .ZN(n8637) );
  NAND2_X1 U11024 ( .A1(n8637), .A2(n11104), .ZN(n8661) );
  NAND2_X1 U11025 ( .A1(n8663), .A2(n8661), .ZN(n8638) );
  XNOR2_X1 U11026 ( .A(n8639), .B(n8638), .ZN(n12317) );
  NAND2_X1 U11027 ( .A1(n12317), .A2(n8761), .ZN(n8641) );
  OR2_X1 U11028 ( .A1(n8762), .A2(n13823), .ZN(n8640) );
  NAND2_X1 U11029 ( .A1(n13724), .A2(n8736), .ZN(n8652) );
  INV_X1 U11030 ( .A(n8643), .ZN(n8642) );
  INV_X1 U11031 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n13306) );
  NAND2_X1 U11032 ( .A1(n8643), .A2(n13306), .ZN(n8644) );
  NAND2_X1 U11033 ( .A1(n8672), .A2(n8644), .ZN(n13551) );
  OR2_X1 U11034 ( .A1(n13551), .A2(n8767), .ZN(n8650) );
  INV_X1 U11035 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n8647) );
  NAND2_X1 U11036 ( .A1(n8747), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n8646) );
  NAND2_X1 U11037 ( .A1(n8768), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n8645) );
  OAI211_X1 U11038 ( .C1(n8647), .C2(n8771), .A(n8646), .B(n8645), .ZN(n8648)
         );
  INV_X1 U11039 ( .A(n8648), .ZN(n8649) );
  NAND2_X1 U11040 ( .A1(n13378), .A2(n8780), .ZN(n8651) );
  NAND2_X1 U11041 ( .A1(n8652), .A2(n8651), .ZN(n8654) );
  AOI22_X1 U11042 ( .A1(n13724), .A2(n8780), .B1(n13378), .B2(n8736), .ZN(
        n8653) );
  AOI21_X1 U11043 ( .B1(n8655), .B2(n8654), .A(n8653), .ZN(n8656) );
  OAI21_X1 U11044 ( .B1(n10910), .B2(n8657), .A(n8663), .ZN(n8658) );
  NOR2_X1 U11045 ( .A1(n8660), .A2(SI_24_), .ZN(n8664) );
  INV_X1 U11046 ( .A(n8661), .ZN(n8662) );
  AOI21_X1 U11047 ( .B1(n8664), .B2(n8663), .A(n8662), .ZN(n8665) );
  MUX2_X1 U11048 ( .A(n11564), .B(n11397), .S(n9438), .Z(n8686) );
  XNOR2_X1 U11049 ( .A(n8686), .B(SI_26_), .ZN(n8666) );
  XNOR2_X1 U11050 ( .A(n8685), .B(n8666), .ZN(n11563) );
  NAND2_X1 U11051 ( .A1(n11563), .A2(n8667), .ZN(n8669) );
  OR2_X1 U11052 ( .A1(n8762), .A2(n11397), .ZN(n8668) );
  NAND2_X1 U11053 ( .A1(n13719), .A2(n8738), .ZN(n8681) );
  INV_X1 U11054 ( .A(n8672), .ZN(n8670) );
  NAND2_X1 U11055 ( .A1(n8670), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n8692) );
  INV_X1 U11056 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n8671) );
  NAND2_X1 U11057 ( .A1(n8672), .A2(n8671), .ZN(n8673) );
  NAND2_X1 U11058 ( .A1(n8692), .A2(n8673), .ZN(n12106) );
  INV_X1 U11059 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n8676) );
  NAND2_X1 U11060 ( .A1(n8747), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n8675) );
  NAND2_X1 U11061 ( .A1(n8768), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n8674) );
  OAI211_X1 U11062 ( .C1(n8676), .C2(n8771), .A(n8675), .B(n8674), .ZN(n8677)
         );
  INV_X1 U11063 ( .A(n8677), .ZN(n8678) );
  NAND2_X1 U11064 ( .A1(n13377), .A2(n8736), .ZN(n8680) );
  NAND2_X1 U11065 ( .A1(n8681), .A2(n8680), .ZN(n8683) );
  AOI22_X1 U11066 ( .A1(n13719), .A2(n8736), .B1(n8780), .B2(n13377), .ZN(
        n8682) );
  INV_X1 U11067 ( .A(n8686), .ZN(n8684) );
  MUX2_X1 U11068 ( .A(n11665), .B(n13817), .S(n9438), .Z(n8703) );
  XNOR2_X1 U11069 ( .A(n8703), .B(SI_27_), .ZN(n8687) );
  NAND2_X1 U11070 ( .A1(n11664), .A2(n8761), .ZN(n8689) );
  OR2_X1 U11071 ( .A1(n8762), .A2(n13817), .ZN(n8688) );
  NAND2_X1 U11072 ( .A1(n13711), .A2(n8736), .ZN(n8702) );
  INV_X1 U11073 ( .A(n8692), .ZN(n8690) );
  INV_X1 U11074 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n8691) );
  NAND2_X1 U11075 ( .A1(n8692), .A2(n8691), .ZN(n8693) );
  NAND2_X1 U11076 ( .A1(n13524), .A2(n8694), .ZN(n8700) );
  INV_X1 U11077 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n8697) );
  NAND2_X1 U11078 ( .A1(n8768), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n8696) );
  NAND2_X1 U11079 ( .A1(n8747), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n8695) );
  OAI211_X1 U11080 ( .C1(n8697), .C2(n8771), .A(n8696), .B(n8695), .ZN(n8698)
         );
  INV_X1 U11081 ( .A(n8698), .ZN(n8699) );
  NAND2_X1 U11082 ( .A1(n13376), .A2(n8738), .ZN(n8701) );
  NAND2_X1 U11083 ( .A1(n8702), .A2(n8701), .ZN(n8782) );
  INV_X1 U11084 ( .A(n8703), .ZN(n8706) );
  NOR2_X1 U11085 ( .A1(n8706), .A2(SI_27_), .ZN(n8704) );
  NAND2_X1 U11086 ( .A1(n8706), .A2(SI_27_), .ZN(n8707) );
  MUX2_X1 U11087 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(P1_DATAO_REG_28__SCAN_IN), 
        .S(n9438), .Z(n8709) );
  XNOR2_X1 U11088 ( .A(n8709), .B(SI_28_), .ZN(n8759) );
  MUX2_X1 U11089 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(P1_DATAO_REG_29__SCAN_IN), 
        .S(n9434), .Z(n8710) );
  INV_X1 U11090 ( .A(SI_29_), .ZN(n11670) );
  XNOR2_X1 U11091 ( .A(n8710), .B(n11670), .ZN(n8741) );
  INV_X1 U11092 ( .A(n8710), .ZN(n8711) );
  MUX2_X1 U11093 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(P1_DATAO_REG_30__SCAN_IN), 
        .S(n9434), .Z(n8712) );
  INV_X1 U11094 ( .A(n8712), .ZN(n8713) );
  INV_X1 U11095 ( .A(SI_30_), .ZN(n12522) );
  MUX2_X1 U11096 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n9438), .Z(n8714) );
  XNOR2_X1 U11097 ( .A(n8714), .B(SI_31_), .ZN(n8715) );
  XNOR2_X1 U11098 ( .A(n8716), .B(n8715), .ZN(n13807) );
  NAND2_X1 U11099 ( .A1(n13807), .A2(n8761), .ZN(n8719) );
  INV_X1 U11100 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n8717) );
  OR2_X1 U11101 ( .A1(n8762), .A2(n8717), .ZN(n8718) );
  INV_X1 U11102 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n8722) );
  NAND2_X1 U11103 ( .A1(n8747), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n8721) );
  NAND2_X1 U11104 ( .A1(n8768), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n8720) );
  OAI211_X1 U11105 ( .C1(n8771), .C2(n8722), .A(n8721), .B(n8720), .ZN(n13372)
         );
  NAND2_X1 U11106 ( .A1(n11961), .A2(n8761), .ZN(n8725) );
  INV_X1 U11107 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n12506) );
  OR2_X1 U11108 ( .A1(n8762), .A2(n12506), .ZN(n8724) );
  INV_X1 U11109 ( .A(n11649), .ZN(n14939) );
  AND2_X1 U11110 ( .A1(n14939), .A2(n13490), .ZN(n9925) );
  NAND2_X1 U11111 ( .A1(n10871), .A2(n13680), .ZN(n8824) );
  NAND2_X1 U11112 ( .A1(n14938), .A2(n8824), .ZN(n9827) );
  AOI21_X1 U11113 ( .B1(n9925), .B2(n10871), .A(n9827), .ZN(n8734) );
  NAND2_X1 U11114 ( .A1(n13372), .A2(n8736), .ZN(n8733) );
  INV_X1 U11115 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n8726) );
  OR2_X1 U11116 ( .A1(n8750), .A2(n8726), .ZN(n8732) );
  INV_X1 U11117 ( .A(P2_REG2_REG_30__SCAN_IN), .ZN(n8727) );
  OR2_X1 U11118 ( .A1(n8728), .A2(n8727), .ZN(n8731) );
  INV_X1 U11119 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n8729) );
  OR2_X1 U11120 ( .A1(n8771), .A2(n8729), .ZN(n8730) );
  AND3_X1 U11121 ( .A1(n8732), .A2(n8731), .A3(n8730), .ZN(n8737) );
  AOI21_X1 U11122 ( .B1(n8734), .B2(n8733), .A(n8737), .ZN(n8735) );
  AOI21_X1 U11123 ( .B1(n13498), .B2(n8780), .A(n8735), .ZN(n8792) );
  NAND2_X1 U11124 ( .A1(n13498), .A2(n8736), .ZN(n8740) );
  INV_X1 U11125 ( .A(n8737), .ZN(n13373) );
  NAND2_X1 U11126 ( .A1(n13373), .A2(n8738), .ZN(n8739) );
  NAND2_X1 U11127 ( .A1(n8740), .A2(n8739), .ZN(n8791) );
  XNOR2_X1 U11128 ( .A(n8742), .B(n8741), .ZN(n11661) );
  NAND2_X1 U11129 ( .A1(n11661), .A2(n8761), .ZN(n8744) );
  INV_X1 U11130 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n11663) );
  OR2_X1 U11131 ( .A1(n8762), .A2(n11663), .ZN(n8743) );
  NAND2_X1 U11132 ( .A1(n8745), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n12126) );
  OR2_X1 U11133 ( .A1(n12126), .A2(n8767), .ZN(n8754) );
  INV_X1 U11134 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n8751) );
  NAND2_X1 U11135 ( .A1(n8746), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n8749) );
  NAND2_X1 U11136 ( .A1(n8747), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n8748) );
  OAI211_X1 U11137 ( .C1(n8751), .C2(n8750), .A(n8749), .B(n8748), .ZN(n8752)
         );
  INV_X1 U11138 ( .A(n8752), .ZN(n8753) );
  NAND2_X1 U11139 ( .A1(n8754), .A2(n8753), .ZN(n13374) );
  AND2_X1 U11140 ( .A1(n13374), .A2(n8736), .ZN(n8755) );
  AOI21_X1 U11141 ( .B1(n13700), .B2(n8780), .A(n8755), .ZN(n8789) );
  NAND2_X1 U11142 ( .A1(n13700), .A2(n8736), .ZN(n8757) );
  NAND2_X1 U11143 ( .A1(n13374), .A2(n8069), .ZN(n8756) );
  NAND2_X1 U11144 ( .A1(n8757), .A2(n8756), .ZN(n8788) );
  OAI22_X1 U11145 ( .A1(n8792), .A2(n8791), .B1(n8789), .B2(n8788), .ZN(n8758)
         );
  NAND2_X1 U11146 ( .A1(n8827), .A2(n8758), .ZN(n8794) );
  NAND2_X1 U11147 ( .A1(n11655), .A2(n8761), .ZN(n8764) );
  OR2_X1 U11148 ( .A1(n8762), .A2(n8866), .ZN(n8763) );
  INV_X1 U11149 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n12168) );
  NAND2_X1 U11150 ( .A1(n8765), .A2(n12168), .ZN(n8766) );
  NAND2_X1 U11151 ( .A1(n12126), .A2(n8766), .ZN(n13511) );
  OR2_X1 U11152 ( .A1(n13511), .A2(n8767), .ZN(n8775) );
  INV_X1 U11153 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n8772) );
  NAND2_X1 U11154 ( .A1(n8095), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n8770) );
  NAND2_X1 U11155 ( .A1(n8768), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n8769) );
  OAI211_X1 U11156 ( .C1(n8772), .C2(n8771), .A(n8770), .B(n8769), .ZN(n8773)
         );
  INV_X1 U11157 ( .A(n8773), .ZN(n8774) );
  AND2_X1 U11158 ( .A1(n13375), .A2(n8780), .ZN(n8776) );
  AOI21_X1 U11159 ( .B1(n13706), .B2(n8736), .A(n8776), .ZN(n8785) );
  NAND2_X1 U11160 ( .A1(n13706), .A2(n8069), .ZN(n8778) );
  NAND2_X1 U11161 ( .A1(n13375), .A2(n8736), .ZN(n8777) );
  NAND2_X1 U11162 ( .A1(n8778), .A2(n8777), .ZN(n8784) );
  NAND2_X1 U11163 ( .A1(n8785), .A2(n8784), .ZN(n8779) );
  OAI211_X1 U11164 ( .C1(n8783), .C2(n8782), .A(n8794), .B(n8779), .ZN(n8797)
         );
  AOI22_X1 U11165 ( .A1(n13711), .A2(n8780), .B1(n13376), .B2(n8736), .ZN(
        n8781) );
  AOI21_X1 U11166 ( .B1(n8783), .B2(n8782), .A(n8781), .ZN(n8796) );
  INV_X1 U11167 ( .A(n8784), .ZN(n8787) );
  INV_X1 U11168 ( .A(n8785), .ZN(n8786) );
  AOI22_X1 U11169 ( .A1(n8789), .A2(n8788), .B1(n8787), .B2(n8786), .ZN(n8790)
         );
  NAND2_X1 U11170 ( .A1(n8827), .A2(n8790), .ZN(n8793) );
  AOI22_X1 U11171 ( .A1(n8794), .A2(n8793), .B1(n8792), .B2(n8791), .ZN(n8795)
         );
  OAI21_X1 U11172 ( .B1(n8797), .B2(n8796), .A(n8795), .ZN(n8801) );
  NAND2_X1 U11173 ( .A1(n13372), .A2(n8117), .ZN(n8799) );
  OR2_X1 U11174 ( .A1(n13372), .A2(n8780), .ZN(n8798) );
  MUX2_X1 U11175 ( .A(n8799), .B(n8798), .S(n13694), .Z(n8800) );
  MUX2_X1 U11176 ( .A(n14939), .B(n14938), .S(n9817), .Z(n8802) );
  INV_X1 U11177 ( .A(n8802), .ZN(n8806) );
  XNOR2_X1 U11178 ( .A(n8817), .B(n8808), .ZN(n9641) );
  INV_X1 U11179 ( .A(n9641), .ZN(n9272) );
  NAND2_X1 U11180 ( .A1(n9272), .A2(P2_STATE_REG_SCAN_IN), .ZN(n11267) );
  INV_X1 U11181 ( .A(n11267), .ZN(n8857) );
  NAND2_X1 U11182 ( .A1(n8857), .A2(n13490), .ZN(n8805) );
  NOR2_X1 U11183 ( .A1(n8806), .A2(n8805), .ZN(n8807) );
  NAND2_X1 U11184 ( .A1(n8859), .A2(n8807), .ZN(n8855) );
  NAND2_X1 U11185 ( .A1(n8817), .A2(n8808), .ZN(n8809) );
  NAND2_X1 U11186 ( .A1(n8809), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8810) );
  NAND2_X1 U11187 ( .A1(n8812), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8813) );
  MUX2_X1 U11188 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8813), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n8815) );
  NAND2_X1 U11189 ( .A1(n8815), .A2(n8814), .ZN(n11398) );
  OAI21_X1 U11190 ( .B1(P2_IR_REG_23__SCAN_IN), .B2(P2_IR_REG_24__SCAN_IN), 
        .A(P2_IR_REG_31__SCAN_IN), .ZN(n8816) );
  NAND2_X1 U11191 ( .A1(n8817), .A2(n8816), .ZN(n8819) );
  NAND3_X1 U11192 ( .A1(n11394), .A2(n9800), .A3(n13818), .ZN(n9273) );
  INV_X1 U11193 ( .A(n8820), .ZN(n11657) );
  INV_X1 U11195 ( .A(n8822), .ZN(n8823) );
  INV_X1 U11196 ( .A(n8824), .ZN(n9822) );
  NAND4_X1 U11197 ( .A1(n14932), .A2(n11657), .A3(n13640), .A4(n9822), .ZN(
        n8825) );
  OAI211_X1 U11198 ( .C1(n14939), .C2(n11267), .A(n8825), .B(P2_B_REG_SCAN_IN), 
        .ZN(n8826) );
  XNOR2_X1 U11199 ( .A(n13498), .B(n13373), .ZN(n8853) );
  INV_X1 U11200 ( .A(n13375), .ZN(n8828) );
  NAND2_X1 U11201 ( .A1(n13706), .A2(n8828), .ZN(n8829) );
  NAND2_X1 U11202 ( .A1(n12119), .A2(n8829), .ZN(n13502) );
  XNOR2_X1 U11203 ( .A(n13711), .B(n12143), .ZN(n13518) );
  XNOR2_X1 U11204 ( .A(n13719), .B(n13305), .ZN(n12118) );
  XNOR2_X1 U11205 ( .A(n13735), .B(n13598), .ZN(n13583) );
  XNOR2_X1 U11206 ( .A(n13740), .B(n13625), .ZN(n13612) );
  XNOR2_X1 U11207 ( .A(n13752), .B(n13624), .ZN(n12115) );
  INV_X1 U11208 ( .A(n13641), .ZN(n8830) );
  NAND2_X1 U11209 ( .A1(n13757), .A2(n8830), .ZN(n13636) );
  OR2_X1 U11210 ( .A1(n13757), .A2(n8830), .ZN(n8831) );
  AND2_X1 U11211 ( .A1(n12115), .A2(n13652), .ZN(n8849) );
  XNOR2_X1 U11212 ( .A(n13747), .B(n13643), .ZN(n13616) );
  INV_X1 U11213 ( .A(n13384), .ZN(n13318) );
  NAND2_X1 U11214 ( .A1(n13780), .A2(n13318), .ZN(n11290) );
  OR2_X1 U11215 ( .A1(n13780), .A2(n13318), .ZN(n8832) );
  NAND2_X1 U11216 ( .A1(n11290), .A2(n8832), .ZN(n11299) );
  INV_X1 U11217 ( .A(n13385), .ZN(n11329) );
  XNOR2_X1 U11218 ( .A(n13784), .B(n11329), .ZN(n11283) );
  INV_X1 U11219 ( .A(n13386), .ZN(n11282) );
  XNOR2_X1 U11220 ( .A(n11281), .B(n11282), .ZN(n11128) );
  INV_X1 U11221 ( .A(n13388), .ZN(n11723) );
  XNOR2_X1 U11222 ( .A(n10854), .B(n11723), .ZN(n10860) );
  INV_X1 U11223 ( .A(n13387), .ZN(n11123) );
  XNOR2_X1 U11224 ( .A(n11730), .B(n11123), .ZN(n10862) );
  XNOR2_X1 U11225 ( .A(n14987), .B(n13389), .ZN(n10794) );
  XNOR2_X1 U11226 ( .A(n10380), .B(n13393), .ZN(n10371) );
  INV_X1 U11227 ( .A(n8833), .ZN(n11710) );
  INV_X1 U11228 ( .A(n10299), .ZN(n10194) );
  NAND2_X1 U11229 ( .A1(n8833), .A2(n10194), .ZN(n8834) );
  NAND2_X1 U11230 ( .A1(n13396), .A2(n9834), .ZN(n8837) );
  OAI21_X1 U11231 ( .B1(n8838), .B2(n10216), .A(n10001), .ZN(n14936) );
  NAND4_X1 U11232 ( .A1(n10249), .A2(n9921), .A3(n9817), .A4(n14936), .ZN(
        n8840) );
  INV_X1 U11233 ( .A(n13394), .ZN(n10377) );
  NAND2_X1 U11234 ( .A1(n10377), .A2(n14947), .ZN(n10372) );
  INV_X1 U11235 ( .A(n14947), .ZN(n10317) );
  NAND2_X1 U11236 ( .A1(n10317), .A2(n13394), .ZN(n8839) );
  NAND2_X1 U11237 ( .A1(n10372), .A2(n8839), .ZN(n10196) );
  NOR2_X1 U11238 ( .A1(n8840), .A2(n10196), .ZN(n8842) );
  NAND4_X1 U11239 ( .A1(n10179), .A2(n10371), .A3(n8842), .A4(n9948), .ZN(
        n8843) );
  XNOR2_X1 U11240 ( .A(n10624), .B(n11766), .ZN(n10328) );
  NOR2_X1 U11241 ( .A1(n8843), .A2(n10328), .ZN(n8844) );
  XNOR2_X1 U11242 ( .A(n10779), .B(n13390), .ZN(n10777) );
  XNOR2_X1 U11243 ( .A(n11771), .B(n13391), .ZN(n10627) );
  NAND4_X1 U11244 ( .A1(n10794), .A2(n8844), .A3(n10777), .A4(n10627), .ZN(
        n8845) );
  OR4_X1 U11245 ( .A1(n11128), .A2(n10860), .A3(n10862), .A4(n8845), .ZN(n8846) );
  NOR3_X1 U11246 ( .A1(n11299), .A2(n11283), .A3(n8846), .ZN(n8847) );
  XNOR2_X1 U11247 ( .A(n13767), .B(n13382), .ZN(n11311) );
  XNOR2_X1 U11248 ( .A(n13772), .B(n13383), .ZN(n11301) );
  AND4_X1 U11249 ( .A1(n13616), .A2(n8847), .A3(n11311), .A4(n11301), .ZN(
        n8848) );
  XNOR2_X1 U11250 ( .A(n13763), .B(n13381), .ZN(n13684) );
  NAND4_X1 U11251 ( .A1(n13612), .A2(n8849), .A3(n8848), .A4(n13684), .ZN(
        n8850) );
  OR3_X1 U11252 ( .A1(n12118), .A2(n13583), .A3(n8850), .ZN(n8851) );
  NOR4_X1 U11253 ( .A1(n13502), .A2(n13518), .A3(n13565), .A4(n8851), .ZN(
        n8852) );
  XNOR2_X1 U11254 ( .A(n13700), .B(n13374), .ZN(n12144) );
  XNOR2_X1 U11255 ( .A(n13724), .B(n13378), .ZN(n12117) );
  NAND2_X1 U11256 ( .A1(n10976), .A2(n9817), .ZN(n9813) );
  AOI22_X1 U11257 ( .A1(n11649), .A2(n9832), .B1(n9813), .B2(n13680), .ZN(
        n8856) );
  NAND2_X1 U11258 ( .A1(n8862), .A2(n8861), .ZN(n12677) );
  NOR2_X1 U11259 ( .A1(n8866), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n8864) );
  NAND2_X1 U11260 ( .A1(n8866), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n8867) );
  XNOR2_X1 U11261 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(P2_DATAO_REG_29__SCAN_IN), 
        .ZN(n11642) );
  OR2_X1 U11262 ( .A1(n6480), .A2(n11670), .ZN(n8868) );
  NAND2_X1 U11263 ( .A1(n8880), .A2(n11677), .ZN(n12686) );
  NAND2_X1 U11264 ( .A1(n12687), .A2(n12686), .ZN(n12719) );
  AOI21_X1 U11265 ( .B1(n7954), .B2(n12745), .A(n8869), .ZN(n8870) );
  XOR2_X1 U11266 ( .A(n12719), .B(n8870), .Z(n8879) );
  NAND2_X1 U11267 ( .A1(n7423), .A2(P3_REG2_REG_30__SCAN_IN), .ZN(n8874) );
  NAND2_X1 U11268 ( .A1(n7522), .A2(P3_REG1_REG_30__SCAN_IN), .ZN(n8873) );
  NAND2_X1 U11269 ( .A1(n7454), .A2(P3_REG0_REG_30__SCAN_IN), .ZN(n8872) );
  INV_X1 U11270 ( .A(P3_B_REG_SCAN_IN), .ZN(n8875) );
  OR2_X1 U11271 ( .A1(n7915), .A2(n8875), .ZN(n8876) );
  NAND2_X1 U11272 ( .A1(n13100), .A2(n8876), .ZN(n12860) );
  NOR2_X1 U11273 ( .A1(n12529), .A2(n12860), .ZN(n8877) );
  INV_X1 U11274 ( .A(n8880), .ZN(n12870) );
  INV_X1 U11275 ( .A(P3_REG0_REG_29__SCAN_IN), .ZN(n8881) );
  NOR2_X1 U11276 ( .A1(n15177), .A2(n8881), .ZN(n8882) );
  OAI21_X1 U11277 ( .B1(n8898), .B2(n15175), .A(n8883), .ZN(P3_U3456) );
  INV_X1 U11278 ( .A(P3_REG1_REG_27__SCAN_IN), .ZN(n8894) );
  INV_X1 U11279 ( .A(n8884), .ZN(n8887) );
  NOR2_X1 U11280 ( .A1(n8885), .A2(n12534), .ZN(n8886) );
  AOI22_X1 U11281 ( .A1(n13098), .A2(n12747), .B1(n12745), .B2(n13100), .ZN(
        n8893) );
  INV_X1 U11282 ( .A(n8888), .ZN(n8889) );
  AOI21_X1 U11283 ( .B1(n12534), .B2(n8890), .A(n8889), .ZN(n8891) );
  MUX2_X1 U11284 ( .A(n8894), .B(n8896), .S(n15193), .Z(n8895) );
  NAND2_X1 U11285 ( .A1(n8895), .A2(n7347), .ZN(P3_U3486) );
  NAND2_X1 U11286 ( .A1(n8897), .A2(n7356), .ZN(P3_U3454) );
  INV_X1 U11287 ( .A(P3_REG1_REG_29__SCAN_IN), .ZN(n8899) );
  INV_X1 U11288 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n14628) );
  XOR2_X1 U11289 ( .A(P3_ADDR_REG_16__SCAN_IN), .B(n14628), .Z(n8984) );
  INV_X1 U11290 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n8980) );
  INV_X1 U11291 ( .A(P3_ADDR_REG_14__SCAN_IN), .ZN(n12800) );
  INV_X1 U11292 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n14616) );
  XNOR2_X1 U11293 ( .A(P3_ADDR_REG_14__SCAN_IN), .B(n14616), .ZN(n8927) );
  INV_X1 U11294 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n14586) );
  INV_X1 U11295 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n14574) );
  INV_X1 U11296 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n10224) );
  INV_X1 U11297 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n9975) );
  NOR2_X1 U11298 ( .A1(n9959), .A2(P1_ADDR_REG_0__SCAN_IN), .ZN(n8936) );
  XNOR2_X1 U11299 ( .A(n8902), .B(P3_ADDR_REG_2__SCAN_IN), .ZN(n8932) );
  INV_X1 U11300 ( .A(P3_ADDR_REG_5__SCAN_IN), .ZN(n15078) );
  NOR2_X1 U11301 ( .A1(n8905), .A2(n15078), .ZN(n8907) );
  XNOR2_X1 U11302 ( .A(n9607), .B(P3_ADDR_REG_6__SCAN_IN), .ZN(n8951) );
  NOR2_X1 U11303 ( .A1(n8908), .A2(n7095), .ZN(n8910) );
  XNOR2_X1 U11304 ( .A(n9975), .B(P3_ADDR_REG_8__SCAN_IN), .ZN(n8957) );
  XNOR2_X1 U11305 ( .A(n10224), .B(P3_ADDR_REG_9__SCAN_IN), .ZN(n8964) );
  NOR2_X1 U11306 ( .A1(P1_ADDR_REG_10__SCAN_IN), .A2(n8911), .ZN(n8913) );
  INV_X1 U11307 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n10538) );
  XOR2_X1 U11308 ( .A(n10538), .B(n8911), .Z(n8968) );
  INV_X1 U11309 ( .A(P3_ADDR_REG_10__SCAN_IN), .ZN(n8967) );
  XNOR2_X1 U11310 ( .A(n14574), .B(P3_ADDR_REG_11__SCAN_IN), .ZN(n8972) );
  XNOR2_X1 U11311 ( .A(n14586), .B(P3_ADDR_REG_12__SCAN_IN), .ZN(n8975) );
  INV_X1 U11312 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n14602) );
  NOR2_X1 U11313 ( .A1(P3_ADDR_REG_13__SCAN_IN), .A2(n14602), .ZN(n8917) );
  INV_X1 U11314 ( .A(P3_ADDR_REG_13__SCAN_IN), .ZN(n8916) );
  OR2_X1 U11315 ( .A1(n8980), .A2(P3_ADDR_REG_15__SCAN_IN), .ZN(n8919) );
  NAND2_X1 U11316 ( .A1(n8984), .A2(n8983), .ZN(n8920) );
  NOR2_X1 U11317 ( .A1(P1_ADDR_REG_17__SCAN_IN), .A2(n8921), .ZN(n8923) );
  INV_X1 U11318 ( .A(P3_ADDR_REG_17__SCAN_IN), .ZN(n8925) );
  INV_X1 U11319 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n14646) );
  NOR2_X1 U11320 ( .A1(n8925), .A2(n8924), .ZN(n8922) );
  INV_X1 U11321 ( .A(P3_ADDR_REG_18__SCAN_IN), .ZN(n8991) );
  XOR2_X1 U11322 ( .A(n8991), .B(P1_ADDR_REG_18__SCAN_IN), .Z(n8989) );
  XOR2_X1 U11323 ( .A(n8925), .B(n8924), .Z(n14341) );
  INV_X1 U11324 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n14562) );
  INV_X1 U11325 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n14908) );
  INV_X1 U11326 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n14893) );
  XOR2_X1 U11327 ( .A(n8927), .B(n8926), .Z(n14551) );
  INV_X1 U11328 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n14878) );
  XOR2_X1 U11329 ( .A(n14602), .B(P3_ADDR_REG_13__SCAN_IN), .Z(n8929) );
  XOR2_X1 U11330 ( .A(n8929), .B(n8928), .Z(n14547) );
  INV_X1 U11331 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n9723) );
  INV_X1 U11332 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n13447) );
  NAND2_X1 U11333 ( .A1(P2_ADDR_REG_4__SCAN_IN), .A2(n8931), .ZN(n8945) );
  XOR2_X1 U11334 ( .A(n8931), .B(P2_ADDR_REG_4__SCAN_IN), .Z(n15195) );
  INV_X1 U11335 ( .A(P2_ADDR_REG_2__SCAN_IN), .ZN(n8941) );
  XNOR2_X1 U11336 ( .A(n8933), .B(n8932), .ZN(n14307) );
  XNOR2_X1 U11337 ( .A(n8935), .B(n8934), .ZN(n8937) );
  NAND2_X1 U11338 ( .A1(P2_ADDR_REG_1__SCAN_IN), .A2(n8937), .ZN(n8939) );
  AOI21_X1 U11339 ( .B1(P1_ADDR_REG_0__SCAN_IN), .B2(n9959), .A(n8936), .ZN(
        n15199) );
  INV_X1 U11340 ( .A(P2_ADDR_REG_0__SCAN_IN), .ZN(n15198) );
  NOR2_X1 U11341 ( .A1(n15199), .A2(n15198), .ZN(n15208) );
  XOR2_X1 U11342 ( .A(n8937), .B(P2_ADDR_REG_1__SCAN_IN), .Z(n15207) );
  NAND2_X1 U11343 ( .A1(n15208), .A2(n15207), .ZN(n8938) );
  NAND2_X1 U11344 ( .A1(n8939), .A2(n8938), .ZN(n14308) );
  NAND2_X1 U11345 ( .A1(n14307), .A2(n14308), .ZN(n8940) );
  NOR2_X1 U11346 ( .A1(n14307), .A2(n14308), .ZN(n14306) );
  AOI21_X1 U11347 ( .B1(n8941), .B2(n8940), .A(n14306), .ZN(n15203) );
  XOR2_X1 U11348 ( .A(n6819), .B(n8942), .Z(n15204) );
  NOR2_X1 U11349 ( .A1(n15203), .A2(n15204), .ZN(n8943) );
  INV_X1 U11350 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n15205) );
  NAND2_X1 U11351 ( .A1(n15203), .A2(n15204), .ZN(n15202) );
  OAI21_X1 U11352 ( .B1(n8943), .B2(n15205), .A(n15202), .ZN(n15194) );
  NAND2_X1 U11353 ( .A1(n15195), .A2(n15194), .ZN(n8944) );
  NAND2_X1 U11354 ( .A1(n8950), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n8954) );
  INV_X1 U11355 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n8949) );
  XNOR2_X1 U11356 ( .A(n8952), .B(n8951), .ZN(n14321) );
  NAND2_X1 U11357 ( .A1(n14322), .A2(n14321), .ZN(n8953) );
  INV_X1 U11358 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n9692) );
  XOR2_X1 U11359 ( .A(n9692), .B(n8955), .Z(n15200) );
  XNOR2_X1 U11360 ( .A(n8958), .B(n8957), .ZN(n8959) );
  NAND2_X1 U11361 ( .A1(n8961), .A2(n8959), .ZN(n8963) );
  INV_X1 U11362 ( .A(n8959), .ZN(n8960) );
  NAND2_X1 U11363 ( .A1(n14323), .A2(P2_ADDR_REG_8__SCAN_IN), .ZN(n8962) );
  NAND2_X1 U11364 ( .A1(n8963), .A2(n8962), .ZN(n14326) );
  XNOR2_X1 U11365 ( .A(n8965), .B(n8964), .ZN(n14325) );
  NOR2_X1 U11366 ( .A1(n14326), .A2(n14325), .ZN(n8966) );
  INV_X1 U11367 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n14852) );
  NAND2_X1 U11368 ( .A1(n14326), .A2(n14325), .ZN(n14324) );
  XNOR2_X1 U11369 ( .A(n8968), .B(n8967), .ZN(n8969) );
  NOR2_X1 U11370 ( .A1(n8970), .A2(n8969), .ZN(n14329) );
  NOR2_X1 U11371 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(n14328), .ZN(n8971) );
  XNOR2_X1 U11372 ( .A(n8973), .B(n8972), .ZN(n14542) );
  NAND2_X1 U11373 ( .A1(n14543), .A2(n14542), .ZN(n8974) );
  NOR2_X1 U11374 ( .A1(n14543), .A2(n14542), .ZN(n14541) );
  XNOR2_X1 U11375 ( .A(n8976), .B(n8975), .ZN(n8977) );
  XNOR2_X1 U11376 ( .A(n8978), .B(n8977), .ZN(n14545) );
  NAND2_X1 U11377 ( .A1(n14551), .A2(n14552), .ZN(n8979) );
  XOR2_X1 U11378 ( .A(P3_ADDR_REG_15__SCAN_IN), .B(n8980), .Z(n8982) );
  XNOR2_X1 U11379 ( .A(n8982), .B(n8981), .ZN(n14555) );
  XOR2_X1 U11380 ( .A(n8984), .B(n8983), .Z(n8985) );
  NAND2_X1 U11381 ( .A1(n14562), .A2(n14561), .ZN(n14558) );
  NAND2_X1 U11382 ( .A1(n14341), .A2(n14342), .ZN(n14340) );
  NAND2_X1 U11383 ( .A1(n14302), .A2(n14301), .ZN(n8987) );
  NAND2_X1 U11384 ( .A1(n8989), .A2(n8988), .ZN(n8990) );
  OAI21_X1 U11385 ( .B1(n8991), .B2(P1_ADDR_REG_18__SCAN_IN), .A(n8990), .ZN(
        n8994) );
  XNOR2_X1 U11386 ( .A(P3_ADDR_REG_19__SCAN_IN), .B(P2_ADDR_REG_19__SCAN_IN), 
        .ZN(n8992) );
  INV_X1 U11387 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n14056) );
  XNOR2_X1 U11388 ( .A(n8992), .B(n14056), .ZN(n8993) );
  XNOR2_X1 U11389 ( .A(n8994), .B(n8993), .ZN(n9163) );
  INV_X1 U11390 ( .A(P3_REG3_REG_18__SCAN_IN), .ZN(n9074) );
  AOI22_X1 U11391 ( .A1(SI_17_), .A2(keyinput_f15), .B1(
        P3_REG3_REG_10__SCAN_IN), .B2(keyinput_f39), .ZN(n8995) );
  OAI221_X1 U11392 ( .B1(SI_17_), .B2(keyinput_f15), .C1(
        P3_REG3_REG_10__SCAN_IN), .C2(keyinput_f39), .A(n8995), .ZN(n9002) );
  AOI22_X1 U11393 ( .A1(SI_2_), .A2(keyinput_f30), .B1(SI_22_), .B2(
        keyinput_f10), .ZN(n8996) );
  OAI221_X1 U11394 ( .B1(SI_2_), .B2(keyinput_f30), .C1(SI_22_), .C2(
        keyinput_f10), .A(n8996), .ZN(n9001) );
  AOI22_X1 U11395 ( .A1(keyinput_f0), .A2(P3_WR_REG_SCAN_IN), .B1(SI_23_), 
        .B2(keyinput_f9), .ZN(n8997) );
  OAI221_X1 U11396 ( .B1(keyinput_f0), .B2(P3_WR_REG_SCAN_IN), .C1(SI_23_), 
        .C2(keyinput_f9), .A(n8997), .ZN(n9000) );
  AOI22_X1 U11397 ( .A1(SI_11_), .A2(keyinput_f21), .B1(
        P3_REG3_REG_19__SCAN_IN), .B2(keyinput_f41), .ZN(n8998) );
  OAI221_X1 U11398 ( .B1(SI_11_), .B2(keyinput_f21), .C1(
        P3_REG3_REG_19__SCAN_IN), .C2(keyinput_f41), .A(n8998), .ZN(n8999) );
  NOR4_X1 U11399 ( .A1(n9002), .A2(n9001), .A3(n9000), .A4(n8999), .ZN(n9030)
         );
  XNOR2_X1 U11400 ( .A(n7791), .B(keyinput_f51), .ZN(n9009) );
  AOI22_X1 U11401 ( .A1(P3_REG3_REG_15__SCAN_IN), .A2(keyinput_f63), .B1(
        P3_REG3_REG_25__SCAN_IN), .B2(keyinput_f47), .ZN(n9003) );
  OAI221_X1 U11402 ( .B1(P3_REG3_REG_15__SCAN_IN), .B2(keyinput_f63), .C1(
        P3_REG3_REG_25__SCAN_IN), .C2(keyinput_f47), .A(n9003), .ZN(n9008) );
  AOI22_X1 U11403 ( .A1(P3_REG3_REG_0__SCAN_IN), .A2(keyinput_f54), .B1(
        P3_REG3_REG_28__SCAN_IN), .B2(keyinput_f42), .ZN(n9004) );
  OAI221_X1 U11404 ( .B1(P3_REG3_REG_0__SCAN_IN), .B2(keyinput_f54), .C1(
        P3_REG3_REG_28__SCAN_IN), .C2(keyinput_f42), .A(n9004), .ZN(n9007) );
  AOI22_X1 U11405 ( .A1(SI_25_), .A2(keyinput_f7), .B1(SI_14_), .B2(
        keyinput_f18), .ZN(n9005) );
  OAI221_X1 U11406 ( .B1(SI_25_), .B2(keyinput_f7), .C1(SI_14_), .C2(
        keyinput_f18), .A(n9005), .ZN(n9006) );
  NOR4_X1 U11407 ( .A1(n9009), .A2(n9008), .A3(n9007), .A4(n9006), .ZN(n9029)
         );
  AOI22_X1 U11408 ( .A1(SI_3_), .A2(keyinput_f29), .B1(SI_12_), .B2(
        keyinput_f20), .ZN(n9010) );
  OAI221_X1 U11409 ( .B1(SI_3_), .B2(keyinput_f29), .C1(SI_12_), .C2(
        keyinput_f20), .A(n9010), .ZN(n9018) );
  INV_X1 U11410 ( .A(SI_10_), .ZN(n9444) );
  AOI22_X1 U11411 ( .A1(n9566), .A2(keyinput_f19), .B1(keyinput_f22), .B2(
        n9444), .ZN(n9011) );
  OAI221_X1 U11412 ( .B1(n9566), .B2(keyinput_f19), .C1(n9444), .C2(
        keyinput_f22), .A(n9011), .ZN(n9017) );
  AOI22_X1 U11413 ( .A1(SI_26_), .A2(keyinput_f6), .B1(P3_REG3_REG_20__SCAN_IN), .B2(keyinput_f55), .ZN(n9012) );
  OAI221_X1 U11414 ( .B1(SI_26_), .B2(keyinput_f6), .C1(
        P3_REG3_REG_20__SCAN_IN), .C2(keyinput_f55), .A(n9012), .ZN(n9016) );
  XNOR2_X1 U11415 ( .A(P3_REG3_REG_8__SCAN_IN), .B(keyinput_f43), .ZN(n9014)
         );
  XNOR2_X1 U11416 ( .A(SI_9_), .B(keyinput_f23), .ZN(n9013) );
  NAND2_X1 U11417 ( .A1(n9014), .A2(n9013), .ZN(n9015) );
  NOR4_X1 U11418 ( .A1(n9018), .A2(n9017), .A3(n9016), .A4(n9015), .ZN(n9028)
         );
  AOI22_X1 U11419 ( .A1(P3_REG3_REG_22__SCAN_IN), .A2(keyinput_f57), .B1(
        P3_REG3_REG_26__SCAN_IN), .B2(keyinput_f62), .ZN(n9019) );
  OAI221_X1 U11420 ( .B1(P3_REG3_REG_22__SCAN_IN), .B2(keyinput_f57), .C1(
        P3_REG3_REG_26__SCAN_IN), .C2(keyinput_f62), .A(n9019), .ZN(n9026) );
  AOI22_X1 U11421 ( .A1(SI_28_), .A2(keyinput_f4), .B1(P3_REG3_REG_3__SCAN_IN), 
        .B2(keyinput_f40), .ZN(n9020) );
  OAI221_X1 U11422 ( .B1(SI_28_), .B2(keyinput_f4), .C1(P3_REG3_REG_3__SCAN_IN), .C2(keyinput_f40), .A(n9020), .ZN(n9025) );
  AOI22_X1 U11423 ( .A1(P3_REG3_REG_5__SCAN_IN), .A2(keyinput_f49), .B1(
        P3_REG3_REG_12__SCAN_IN), .B2(keyinput_f46), .ZN(n9021) );
  OAI221_X1 U11424 ( .B1(P3_REG3_REG_5__SCAN_IN), .B2(keyinput_f49), .C1(
        P3_REG3_REG_12__SCAN_IN), .C2(keyinput_f46), .A(n9021), .ZN(n9024) );
  AOI22_X1 U11425 ( .A1(SI_30_), .A2(keyinput_f2), .B1(SI_15_), .B2(
        keyinput_f17), .ZN(n9022) );
  OAI221_X1 U11426 ( .B1(SI_30_), .B2(keyinput_f2), .C1(SI_15_), .C2(
        keyinput_f17), .A(n9022), .ZN(n9023) );
  NOR4_X1 U11427 ( .A1(n9026), .A2(n9025), .A3(n9024), .A4(n9023), .ZN(n9027)
         );
  NAND4_X1 U11428 ( .A1(n9030), .A2(n9029), .A3(n9028), .A4(n9027), .ZN(n9072)
         );
  INV_X1 U11429 ( .A(P3_REG3_REG_6__SCAN_IN), .ZN(n10084) );
  AOI22_X1 U11430 ( .A1(n9679), .A2(keyinput_f16), .B1(n10084), .B2(
        keyinput_f61), .ZN(n9031) );
  OAI221_X1 U11431 ( .B1(n9679), .B2(keyinput_f16), .C1(n10084), .C2(
        keyinput_f61), .A(n9031), .ZN(n9039) );
  XOR2_X1 U11432 ( .A(SI_4_), .B(keyinput_f28), .Z(n9038) );
  XNOR2_X1 U11433 ( .A(SI_1_), .B(keyinput_f31), .ZN(n9035) );
  XNOR2_X1 U11434 ( .A(SI_7_), .B(keyinput_f25), .ZN(n9034) );
  XNOR2_X1 U11435 ( .A(P3_REG3_REG_23__SCAN_IN), .B(keyinput_f38), .ZN(n9033)
         );
  XNOR2_X1 U11436 ( .A(SI_5_), .B(keyinput_f27), .ZN(n9032) );
  NAND4_X1 U11437 ( .A1(n9035), .A2(n9034), .A3(n9033), .A4(n9032), .ZN(n9037)
         );
  XNOR2_X1 U11438 ( .A(n9125), .B(keyinput_f50), .ZN(n9036) );
  NOR4_X1 U11439 ( .A1(n9039), .A2(n9038), .A3(n9037), .A4(n9036), .ZN(n9070)
         );
  AOI22_X1 U11440 ( .A1(n12401), .A2(keyinput_f48), .B1(n12367), .B2(
        keyinput_f45), .ZN(n9040) );
  OAI221_X1 U11441 ( .B1(n12401), .B2(keyinput_f48), .C1(n12367), .C2(
        keyinput_f45), .A(n9040), .ZN(n9048) );
  AOI22_X1 U11442 ( .A1(n7540), .A2(keyinput_f53), .B1(keyinput_f13), .B2(
        n9992), .ZN(n9041) );
  OAI221_X1 U11443 ( .B1(n7540), .B2(keyinput_f53), .C1(n9992), .C2(
        keyinput_f13), .A(n9041), .ZN(n9047) );
  AOI22_X1 U11444 ( .A1(n7389), .A2(keyinput_f59), .B1(n10910), .B2(
        keyinput_f8), .ZN(n9042) );
  OAI221_X1 U11445 ( .B1(n7389), .B2(keyinput_f59), .C1(n10910), .C2(
        keyinput_f8), .A(n9042), .ZN(n9046) );
  XNOR2_X1 U11446 ( .A(P3_STATE_REG_SCAN_IN), .B(keyinput_f34), .ZN(n9044) );
  XNOR2_X1 U11447 ( .A(SI_0_), .B(keyinput_f32), .ZN(n9043) );
  NAND2_X1 U11448 ( .A1(n9044), .A2(n9043), .ZN(n9045) );
  NOR4_X1 U11449 ( .A1(n9048), .A2(n9047), .A3(n9046), .A4(n9045), .ZN(n9069)
         );
  AOI22_X1 U11450 ( .A1(n10287), .A2(keyinput_f12), .B1(n7620), .B2(
        keyinput_f56), .ZN(n9049) );
  OAI221_X1 U11451 ( .B1(n10287), .B2(keyinput_f12), .C1(n7620), .C2(
        keyinput_f56), .A(n9049), .ZN(n9056) );
  INV_X1 U11452 ( .A(P3_REG3_REG_27__SCAN_IN), .ZN(n9137) );
  AOI22_X1 U11453 ( .A1(n9137), .A2(keyinput_f36), .B1(keyinput_f14), .B2(
        n9883), .ZN(n9050) );
  OAI221_X1 U11454 ( .B1(n9137), .B2(keyinput_f36), .C1(n9883), .C2(
        keyinput_f14), .A(n9050), .ZN(n9055) );
  INV_X1 U11455 ( .A(P3_RD_REG_SCAN_IN), .ZN(n14304) );
  AOI22_X1 U11456 ( .A1(n11273), .A2(keyinput_f5), .B1(keyinput_f33), .B2(
        n14304), .ZN(n9051) );
  OAI221_X1 U11457 ( .B1(n11273), .B2(keyinput_f5), .C1(n14304), .C2(
        keyinput_f33), .A(n9051), .ZN(n9054) );
  INV_X1 U11458 ( .A(P3_REG3_REG_4__SCAN_IN), .ZN(n9124) );
  INV_X1 U11459 ( .A(SI_31_), .ZN(n13245) );
  AOI22_X1 U11460 ( .A1(n9124), .A2(keyinput_f52), .B1(keyinput_f1), .B2(
        n13245), .ZN(n9052) );
  OAI221_X1 U11461 ( .B1(n9124), .B2(keyinput_f52), .C1(n13245), .C2(
        keyinput_f1), .A(n9052), .ZN(n9053) );
  NOR4_X1 U11462 ( .A1(n9056), .A2(n9055), .A3(n9054), .A4(n9053), .ZN(n9068)
         );
  INV_X1 U11463 ( .A(P3_REG3_REG_11__SCAN_IN), .ZN(n9147) );
  AOI22_X1 U11464 ( .A1(n10423), .A2(keyinput_f11), .B1(n9147), .B2(
        keyinput_f58), .ZN(n9057) );
  OAI221_X1 U11465 ( .B1(n10423), .B2(keyinput_f11), .C1(n9147), .C2(
        keyinput_f58), .A(n9057), .ZN(n9066) );
  INV_X1 U11466 ( .A(P3_REG3_REG_1__SCAN_IN), .ZN(n10417) );
  INV_X1 U11467 ( .A(P3_REG3_REG_14__SCAN_IN), .ZN(n9059) );
  AOI22_X1 U11468 ( .A1(n10417), .A2(keyinput_f44), .B1(n9059), .B2(
        keyinput_f37), .ZN(n9058) );
  OAI221_X1 U11469 ( .B1(n10417), .B2(keyinput_f44), .C1(n9059), .C2(
        keyinput_f37), .A(n9058), .ZN(n9065) );
  XNOR2_X1 U11470 ( .A(SI_29_), .B(keyinput_f3), .ZN(n9063) );
  XNOR2_X1 U11471 ( .A(SI_8_), .B(keyinput_f24), .ZN(n9062) );
  XNOR2_X1 U11472 ( .A(SI_6_), .B(keyinput_f26), .ZN(n9061) );
  XNOR2_X1 U11473 ( .A(keyinput_f35), .B(P3_REG3_REG_7__SCAN_IN), .ZN(n9060)
         );
  NAND4_X1 U11474 ( .A1(n9063), .A2(n9062), .A3(n9061), .A4(n9060), .ZN(n9064)
         );
  NOR3_X1 U11475 ( .A1(n9066), .A2(n9065), .A3(n9064), .ZN(n9067) );
  NAND4_X1 U11476 ( .A1(n9070), .A2(n9069), .A3(n9068), .A4(n9067), .ZN(n9071)
         );
  OAI22_X1 U11477 ( .A1(keyinput_f60), .A2(n9074), .B1(n9072), .B2(n9071), 
        .ZN(n9073) );
  AOI21_X1 U11478 ( .B1(keyinput_f60), .B2(n9074), .A(n9073), .ZN(n9161) );
  AOI22_X1 U11479 ( .A1(SI_20_), .A2(keyinput_g12), .B1(SI_11_), .B2(
        keyinput_g21), .ZN(n9075) );
  OAI221_X1 U11480 ( .B1(SI_20_), .B2(keyinput_g12), .C1(SI_11_), .C2(
        keyinput_g21), .A(n9075), .ZN(n9082) );
  AOI22_X1 U11481 ( .A1(SI_14_), .A2(keyinput_g18), .B1(SI_22_), .B2(
        keyinput_g10), .ZN(n9076) );
  OAI221_X1 U11482 ( .B1(SI_14_), .B2(keyinput_g18), .C1(SI_22_), .C2(
        keyinput_g10), .A(n9076), .ZN(n9081) );
  AOI22_X1 U11483 ( .A1(SI_5_), .A2(keyinput_g27), .B1(SI_29_), .B2(
        keyinput_g3), .ZN(n9077) );
  OAI221_X1 U11484 ( .B1(SI_5_), .B2(keyinput_g27), .C1(SI_29_), .C2(
        keyinput_g3), .A(n9077), .ZN(n9080) );
  AOI22_X1 U11485 ( .A1(P3_REG3_REG_22__SCAN_IN), .A2(keyinput_g57), .B1(
        P3_REG3_REG_26__SCAN_IN), .B2(keyinput_g62), .ZN(n9078) );
  OAI221_X1 U11486 ( .B1(P3_REG3_REG_22__SCAN_IN), .B2(keyinput_g57), .C1(
        P3_REG3_REG_26__SCAN_IN), .C2(keyinput_g62), .A(n9078), .ZN(n9079) );
  NOR4_X1 U11487 ( .A1(n9082), .A2(n9081), .A3(n9080), .A4(n9079), .ZN(n9111)
         );
  AOI22_X1 U11488 ( .A1(P3_RD_REG_SCAN_IN), .A2(keyinput_g33), .B1(SI_15_), 
        .B2(keyinput_g17), .ZN(n9083) );
  OAI221_X1 U11489 ( .B1(P3_RD_REG_SCAN_IN), .B2(keyinput_g33), .C1(SI_15_), 
        .C2(keyinput_g17), .A(n9083), .ZN(n9089) );
  INV_X1 U11490 ( .A(P3_REG3_REG_0__SCAN_IN), .ZN(n10107) );
  AOI22_X1 U11491 ( .A1(P3_STATE_REG_SCAN_IN), .A2(keyinput_g34), .B1(n10107), 
        .B2(keyinput_g54), .ZN(n9084) );
  OAI221_X1 U11492 ( .B1(P3_STATE_REG_SCAN_IN), .B2(keyinput_g34), .C1(n10107), 
        .C2(keyinput_g54), .A(n9084), .ZN(n9088) );
  AOI22_X1 U11493 ( .A1(P3_REG3_REG_14__SCAN_IN), .A2(keyinput_g37), .B1(
        P3_REG3_REG_15__SCAN_IN), .B2(keyinput_g63), .ZN(n9085) );
  OAI221_X1 U11494 ( .B1(P3_REG3_REG_14__SCAN_IN), .B2(keyinput_g37), .C1(
        P3_REG3_REG_15__SCAN_IN), .C2(keyinput_g63), .A(n9085), .ZN(n9087) );
  XNOR2_X1 U11495 ( .A(SI_4_), .B(keyinput_g28), .ZN(n9086) );
  NOR4_X1 U11496 ( .A1(n9089), .A2(n9088), .A3(n9087), .A4(n9086), .ZN(n9110)
         );
  AOI22_X1 U11497 ( .A1(SI_0_), .A2(keyinput_g32), .B1(P3_REG3_REG_12__SCAN_IN), .B2(keyinput_g46), .ZN(n9090) );
  OAI221_X1 U11498 ( .B1(SI_0_), .B2(keyinput_g32), .C1(
        P3_REG3_REG_12__SCAN_IN), .C2(keyinput_g46), .A(n9090), .ZN(n9099) );
  AOI22_X1 U11499 ( .A1(P3_REG3_REG_2__SCAN_IN), .A2(keyinput_g59), .B1(SI_17_), .B2(keyinput_g15), .ZN(n9091) );
  OAI221_X1 U11500 ( .B1(P3_REG3_REG_2__SCAN_IN), .B2(keyinput_g59), .C1(
        SI_17_), .C2(keyinput_g15), .A(n9091), .ZN(n9098) );
  INV_X1 U11501 ( .A(P3_WR_REG_SCAN_IN), .ZN(n9093) );
  AOI22_X1 U11502 ( .A1(n9093), .A2(keyinput_g0), .B1(n9444), .B2(keyinput_g22), .ZN(n9092) );
  OAI221_X1 U11503 ( .B1(n9093), .B2(keyinput_g0), .C1(n9444), .C2(
        keyinput_g22), .A(n9092), .ZN(n9097) );
  AOI22_X1 U11504 ( .A1(n9095), .A2(keyinput_g40), .B1(keyinput_g20), .B2(
        n9489), .ZN(n9094) );
  OAI221_X1 U11505 ( .B1(n9095), .B2(keyinput_g40), .C1(n9489), .C2(
        keyinput_g20), .A(n9094), .ZN(n9096) );
  NOR4_X1 U11506 ( .A1(n9099), .A2(n9098), .A3(n9097), .A4(n9096), .ZN(n9109)
         );
  AOI22_X1 U11507 ( .A1(SI_2_), .A2(keyinput_g30), .B1(P3_REG3_REG_28__SCAN_IN), .B2(keyinput_g42), .ZN(n9100) );
  OAI221_X1 U11508 ( .B1(SI_2_), .B2(keyinput_g30), .C1(
        P3_REG3_REG_28__SCAN_IN), .C2(keyinput_g42), .A(n9100), .ZN(n9107) );
  AOI22_X1 U11509 ( .A1(SI_8_), .A2(keyinput_g24), .B1(SI_13_), .B2(
        keyinput_g19), .ZN(n9101) );
  OAI221_X1 U11510 ( .B1(SI_8_), .B2(keyinput_g24), .C1(SI_13_), .C2(
        keyinput_g19), .A(n9101), .ZN(n9106) );
  AOI22_X1 U11511 ( .A1(SI_25_), .A2(keyinput_g7), .B1(SI_3_), .B2(
        keyinput_g29), .ZN(n9102) );
  OAI221_X1 U11512 ( .B1(SI_25_), .B2(keyinput_g7), .C1(SI_3_), .C2(
        keyinput_g29), .A(n9102), .ZN(n9105) );
  AOI22_X1 U11513 ( .A1(SI_9_), .A2(keyinput_g23), .B1(P3_REG3_REG_19__SCAN_IN), .B2(keyinput_g41), .ZN(n9103) );
  OAI221_X1 U11514 ( .B1(SI_9_), .B2(keyinput_g23), .C1(
        P3_REG3_REG_19__SCAN_IN), .C2(keyinput_g41), .A(n9103), .ZN(n9104) );
  NOR4_X1 U11515 ( .A1(n9107), .A2(n9106), .A3(n9105), .A4(n9104), .ZN(n9108)
         );
  NAND4_X1 U11516 ( .A1(n9111), .A2(n9110), .A3(n9109), .A4(n9108), .ZN(n9159)
         );
  INV_X1 U11517 ( .A(SI_23_), .ZN(n9113) );
  AOI22_X1 U11518 ( .A1(n9113), .A2(keyinput_g9), .B1(n12367), .B2(
        keyinput_g45), .ZN(n9112) );
  OAI221_X1 U11519 ( .B1(n9113), .B2(keyinput_g9), .C1(n12367), .C2(
        keyinput_g45), .A(n9112), .ZN(n9121) );
  AOI22_X1 U11520 ( .A1(n10279), .A2(keyinput_g43), .B1(keyinput_g44), .B2(
        n10417), .ZN(n9114) );
  OAI221_X1 U11521 ( .B1(n10279), .B2(keyinput_g43), .C1(n10417), .C2(
        keyinput_g44), .A(n9114), .ZN(n9120) );
  AOI22_X1 U11522 ( .A1(n11202), .A2(keyinput_g6), .B1(n12401), .B2(
        keyinput_g48), .ZN(n9115) );
  OAI221_X1 U11523 ( .B1(n11202), .B2(keyinput_g6), .C1(n12401), .C2(
        keyinput_g48), .A(n9115), .ZN(n9119) );
  XNOR2_X1 U11524 ( .A(SI_6_), .B(keyinput_g26), .ZN(n9117) );
  XNOR2_X1 U11525 ( .A(SI_19_), .B(keyinput_g13), .ZN(n9116) );
  NAND2_X1 U11526 ( .A1(n9117), .A2(n9116), .ZN(n9118) );
  NOR4_X1 U11527 ( .A1(n9121), .A2(n9120), .A3(n9119), .A4(n9118), .ZN(n9157)
         );
  AOI22_X1 U11528 ( .A1(n7620), .A2(keyinput_g56), .B1(n7791), .B2(
        keyinput_g51), .ZN(n9122) );
  OAI221_X1 U11529 ( .B1(n7620), .B2(keyinput_g56), .C1(n7791), .C2(
        keyinput_g51), .A(n9122), .ZN(n9132) );
  AOI22_X1 U11530 ( .A1(n9125), .A2(keyinput_g50), .B1(keyinput_g52), .B2(
        n9124), .ZN(n9123) );
  OAI221_X1 U11531 ( .B1(n9125), .B2(keyinput_g50), .C1(n9124), .C2(
        keyinput_g52), .A(n9123), .ZN(n9131) );
  INV_X1 U11532 ( .A(P3_REG3_REG_25__SCAN_IN), .ZN(n12392) );
  AOI22_X1 U11533 ( .A1(n10084), .A2(keyinput_g61), .B1(n12392), .B2(
        keyinput_g47), .ZN(n9126) );
  OAI221_X1 U11534 ( .B1(n10084), .B2(keyinput_g61), .C1(n12392), .C2(
        keyinput_g47), .A(n9126), .ZN(n9130) );
  XNOR2_X1 U11535 ( .A(SI_1_), .B(keyinput_g31), .ZN(n9128) );
  XNOR2_X1 U11536 ( .A(keyinput_g35), .B(P3_REG3_REG_7__SCAN_IN), .ZN(n9127)
         );
  NAND2_X1 U11537 ( .A1(n9128), .A2(n9127), .ZN(n9129) );
  NOR4_X1 U11538 ( .A1(n9132), .A2(n9131), .A3(n9130), .A4(n9129), .ZN(n9156)
         );
  AOI22_X1 U11539 ( .A1(n10910), .A2(keyinput_g8), .B1(n9134), .B2(
        keyinput_g55), .ZN(n9133) );
  OAI221_X1 U11540 ( .B1(n10910), .B2(keyinput_g8), .C1(n9134), .C2(
        keyinput_g55), .A(n9133), .ZN(n9143) );
  INV_X1 U11541 ( .A(P3_REG3_REG_10__SCAN_IN), .ZN(n10704) );
  AOI22_X1 U11542 ( .A1(n9883), .A2(keyinput_g14), .B1(n10704), .B2(
        keyinput_g39), .ZN(n9135) );
  OAI221_X1 U11543 ( .B1(n9883), .B2(keyinput_g14), .C1(n10704), .C2(
        keyinput_g39), .A(n9135), .ZN(n9142) );
  AOI22_X1 U11544 ( .A1(n9679), .A2(keyinput_g16), .B1(n9137), .B2(
        keyinput_g36), .ZN(n9136) );
  OAI221_X1 U11545 ( .B1(n9679), .B2(keyinput_g16), .C1(n9137), .C2(
        keyinput_g36), .A(n9136), .ZN(n9141) );
  XOR2_X1 U11546 ( .A(n7540), .B(keyinput_g53), .Z(n9139) );
  XNOR2_X1 U11547 ( .A(SI_7_), .B(keyinput_g25), .ZN(n9138) );
  NAND2_X1 U11548 ( .A1(n9139), .A2(n9138), .ZN(n9140) );
  NOR4_X1 U11549 ( .A1(n9143), .A2(n9142), .A3(n9141), .A4(n9140), .ZN(n9155)
         );
  AOI22_X1 U11550 ( .A1(n13248), .A2(keyinput_g4), .B1(keyinput_g2), .B2(
        n12522), .ZN(n9144) );
  OAI221_X1 U11551 ( .B1(n13248), .B2(keyinput_g4), .C1(n12522), .C2(
        keyinput_g2), .A(n9144), .ZN(n9153) );
  AOI22_X1 U11552 ( .A1(n13245), .A2(keyinput_g1), .B1(n10423), .B2(
        keyinput_g11), .ZN(n9145) );
  OAI221_X1 U11553 ( .B1(n13245), .B2(keyinput_g1), .C1(n10423), .C2(
        keyinput_g11), .A(n9145), .ZN(n9152) );
  AOI22_X1 U11554 ( .A1(n9147), .A2(keyinput_g58), .B1(keyinput_g5), .B2(
        n11273), .ZN(n9146) );
  OAI221_X1 U11555 ( .B1(n9147), .B2(keyinput_g58), .C1(n11273), .C2(
        keyinput_g5), .A(n9146), .ZN(n9151) );
  INV_X1 U11556 ( .A(P3_REG3_REG_5__SCAN_IN), .ZN(n9149) );
  AOI22_X1 U11557 ( .A1(n9149), .A2(keyinput_g49), .B1(n12340), .B2(
        keyinput_g38), .ZN(n9148) );
  OAI221_X1 U11558 ( .B1(n9149), .B2(keyinput_g49), .C1(n12340), .C2(
        keyinput_g38), .A(n9148), .ZN(n9150) );
  NOR4_X1 U11559 ( .A1(n9153), .A2(n9152), .A3(n9151), .A4(n9150), .ZN(n9154)
         );
  NAND4_X1 U11560 ( .A1(n9157), .A2(n9156), .A3(n9155), .A4(n9154), .ZN(n9158)
         );
  OAI22_X1 U11561 ( .A1(P3_REG3_REG_18__SCAN_IN), .A2(keyinput_g60), .B1(n9159), .B2(n9158), .ZN(n9160) );
  AOI211_X1 U11562 ( .C1(P3_REG3_REG_18__SCAN_IN), .C2(keyinput_g60), .A(n9161), .B(n9160), .ZN(n9162) );
  XNOR2_X1 U11563 ( .A(n9163), .B(n9162), .ZN(n9164) );
  NAND2_X1 U11564 ( .A1(n13239), .A2(n12727), .ZN(n9166) );
  OAI21_X1 U11565 ( .B1(n12547), .B2(n12857), .A(n10288), .ZN(n9165) );
  XNOR2_X1 U11566 ( .A(n12535), .B(n9242), .ZN(n11678) );
  NOR2_X1 U11567 ( .A1(n11678), .A2(n12746), .ZN(n11673) );
  AOI21_X1 U11568 ( .B1(n11678), .B2(n12746), .A(n11673), .ZN(n9245) );
  NAND2_X1 U11569 ( .A1(n12559), .A2(n11671), .ZN(n9168) );
  NAND2_X1 U11570 ( .A1(n15113), .A2(n9178), .ZN(n9167) );
  NAND3_X1 U11571 ( .A1(n12764), .A2(n9178), .A3(n10416), .ZN(n9169) );
  AND2_X1 U11572 ( .A1(n9173), .A2(n9169), .ZN(n10202) );
  NAND2_X1 U11573 ( .A1(n10412), .A2(n9178), .ZN(n9170) );
  NAND2_X1 U11574 ( .A1(n9171), .A2(n9170), .ZN(n9172) );
  NAND2_X1 U11575 ( .A1(n10202), .A2(n9172), .ZN(n10199) );
  NAND2_X1 U11576 ( .A1(n10199), .A2(n9173), .ZN(n10289) );
  XNOR2_X1 U11577 ( .A(n9175), .B(n6469), .ZN(n10290) );
  INV_X1 U11578 ( .A(n9175), .ZN(n9176) );
  NOR2_X1 U11579 ( .A1(n9176), .A2(n6469), .ZN(n9177) );
  XNOR2_X1 U11580 ( .A(n15135), .B(n9178), .ZN(n9179) );
  XNOR2_X1 U11581 ( .A(n9179), .B(n12763), .ZN(n10361) );
  INV_X1 U11582 ( .A(n9179), .ZN(n9180) );
  NAND2_X1 U11583 ( .A1(n9180), .A2(n12763), .ZN(n9181) );
  XNOR2_X1 U11584 ( .A(n15140), .B(n11671), .ZN(n9183) );
  XNOR2_X1 U11585 ( .A(n9183), .B(n12762), .ZN(n10660) );
  INV_X1 U11586 ( .A(n9183), .ZN(n9184) );
  NAND2_X1 U11587 ( .A1(n10363), .A2(n9184), .ZN(n9185) );
  XNOR2_X1 U11588 ( .A(n15146), .B(n9242), .ZN(n9186) );
  XNOR2_X1 U11589 ( .A(n9186), .B(n12761), .ZN(n10753) );
  NAND2_X1 U11590 ( .A1(n10876), .A2(n9186), .ZN(n9187) );
  XNOR2_X1 U11591 ( .A(n15151), .B(n9242), .ZN(n9189) );
  XNOR2_X1 U11592 ( .A(n9189), .B(n12760), .ZN(n10809) );
  INV_X1 U11593 ( .A(n10809), .ZN(n9188) );
  NAND2_X1 U11594 ( .A1(n9189), .A2(n12760), .ZN(n9190) );
  NAND2_X1 U11595 ( .A1(n10811), .A2(n9190), .ZN(n12321) );
  XNOR2_X1 U11596 ( .A(n15157), .B(n9242), .ZN(n9191) );
  XNOR2_X1 U11597 ( .A(n9191), .B(n12759), .ZN(n12320) );
  NAND2_X1 U11598 ( .A1(n12321), .A2(n12320), .ZN(n12319) );
  INV_X1 U11599 ( .A(n9191), .ZN(n9192) );
  NAND2_X1 U11600 ( .A1(n9192), .A2(n12759), .ZN(n9193) );
  NAND2_X1 U11601 ( .A1(n12319), .A2(n9193), .ZN(n11042) );
  XNOR2_X1 U11602 ( .A(n11045), .B(n11671), .ZN(n9194) );
  XNOR2_X1 U11603 ( .A(n9194), .B(n12758), .ZN(n11041) );
  INV_X1 U11604 ( .A(n9194), .ZN(n9195) );
  NAND2_X1 U11605 ( .A1(n9195), .A2(n12758), .ZN(n9196) );
  XNOR2_X1 U11606 ( .A(n15169), .B(n11671), .ZN(n9198) );
  XNOR2_X1 U11607 ( .A(n9198), .B(n13099), .ZN(n12422) );
  INV_X1 U11608 ( .A(n12422), .ZN(n9197) );
  XNOR2_X1 U11609 ( .A(n13233), .B(n11671), .ZN(n9202) );
  XNOR2_X1 U11610 ( .A(n9202), .B(n13086), .ZN(n12346) );
  INV_X1 U11611 ( .A(n12346), .ZN(n9200) );
  INV_X1 U11612 ( .A(n9198), .ZN(n9199) );
  NAND2_X1 U11613 ( .A1(n12352), .A2(n9199), .ZN(n12345) );
  AND2_X1 U11614 ( .A1(n9200), .A2(n12345), .ZN(n9201) );
  NAND2_X1 U11615 ( .A1(n12344), .A2(n9201), .ZN(n12348) );
  NAND2_X1 U11616 ( .A1(n9202), .A2(n13086), .ZN(n9203) );
  XNOR2_X1 U11617 ( .A(n14428), .B(n9242), .ZN(n12371) );
  XNOR2_X1 U11618 ( .A(n14425), .B(n9242), .ZN(n12374) );
  NAND2_X1 U11619 ( .A1(n12374), .A2(n13087), .ZN(n9207) );
  OAI21_X1 U11620 ( .B1(n12464), .B2(n12371), .A(n9207), .ZN(n9209) );
  AND2_X1 U11621 ( .A1(n12371), .A2(n12464), .ZN(n9206) );
  INV_X1 U11622 ( .A(n12374), .ZN(n9204) );
  AOI22_X1 U11623 ( .A1(n9207), .A2(n9206), .B1(n9205), .B2(n9204), .ZN(n9208)
         );
  XNOR2_X1 U11624 ( .A(n14417), .B(n9242), .ZN(n12438) );
  AND2_X1 U11625 ( .A1(n12438), .A2(n12437), .ZN(n9210) );
  INV_X1 U11626 ( .A(n12438), .ZN(n9211) );
  XNOR2_X1 U11627 ( .A(n14413), .B(n9242), .ZN(n9212) );
  NAND2_X1 U11628 ( .A1(n9212), .A2(n12493), .ZN(n9215) );
  INV_X1 U11629 ( .A(n9212), .ZN(n9213) );
  NAND2_X1 U11630 ( .A1(n9213), .A2(n13063), .ZN(n9214) );
  AND2_X1 U11631 ( .A1(n9215), .A2(n9214), .ZN(n12329) );
  XNOR2_X1 U11632 ( .A(n13231), .B(n9242), .ZN(n12490) );
  XNOR2_X1 U11633 ( .A(n13167), .B(n11671), .ZN(n9216) );
  NOR2_X1 U11634 ( .A1(n9216), .A2(n13017), .ZN(n12399) );
  NAND2_X1 U11635 ( .A1(n9216), .A2(n13017), .ZN(n12397) );
  XNOR2_X1 U11636 ( .A(n13226), .B(n11671), .ZN(n9217) );
  XNOR2_X1 U11637 ( .A(n9217), .B(n12756), .ZN(n12406) );
  INV_X1 U11638 ( .A(n9217), .ZN(n9218) );
  XNOR2_X1 U11639 ( .A(n13004), .B(n11671), .ZN(n9219) );
  XNOR2_X1 U11640 ( .A(n9219), .B(n12755), .ZN(n12470) );
  INV_X1 U11641 ( .A(n9219), .ZN(n9220) );
  XNOR2_X1 U11642 ( .A(n12991), .B(n11671), .ZN(n9221) );
  XOR2_X1 U11643 ( .A(n12754), .B(n9221), .Z(n12356) );
  XNOR2_X1 U11644 ( .A(n13145), .B(n11671), .ZN(n9223) );
  XNOR2_X1 U11645 ( .A(n9223), .B(n12753), .ZN(n12430) );
  INV_X1 U11646 ( .A(n9223), .ZN(n9224) );
  AOI21_X1 U11647 ( .B1(n12431), .B2(n12430), .A(n7361), .ZN(n12364) );
  XNOR2_X1 U11648 ( .A(n12545), .B(n9242), .ZN(n9225) );
  NOR2_X1 U11649 ( .A1(n9225), .A2(n12752), .ZN(n9226) );
  AOI21_X1 U11650 ( .B1(n9225), .B2(n12752), .A(n9226), .ZN(n12365) );
  NAND2_X1 U11651 ( .A1(n12364), .A2(n12365), .ZN(n12363) );
  INV_X1 U11652 ( .A(n9226), .ZN(n9227) );
  NAND2_X1 U11653 ( .A1(n12363), .A2(n9227), .ZN(n9229) );
  NAND2_X1 U11654 ( .A1(n9229), .A2(n9228), .ZN(n9230) );
  NAND2_X1 U11655 ( .A1(n6571), .A2(n9230), .ZN(n12449) );
  INV_X1 U11656 ( .A(n9230), .ZN(n9231) );
  XOR2_X1 U11657 ( .A(n11671), .B(n13134), .Z(n9232) );
  XNOR2_X1 U11658 ( .A(n12922), .B(n11671), .ZN(n9234) );
  NAND2_X1 U11659 ( .A1(n9234), .A2(n12389), .ZN(n9237) );
  INV_X1 U11660 ( .A(n9234), .ZN(n9235) );
  NAND2_X1 U11661 ( .A1(n9235), .A2(n12749), .ZN(n9236) );
  NAND2_X1 U11662 ( .A1(n9237), .A2(n9236), .ZN(n12412) );
  INV_X1 U11663 ( .A(n9237), .ZN(n12386) );
  XNOR2_X1 U11664 ( .A(n12382), .B(n11671), .ZN(n9238) );
  NAND2_X1 U11665 ( .A1(n9238), .A2(n12415), .ZN(n9241) );
  INV_X1 U11666 ( .A(n9238), .ZN(n9239) );
  NAND2_X1 U11667 ( .A1(n9239), .A2(n12748), .ZN(n9240) );
  AND2_X1 U11668 ( .A1(n9241), .A2(n9240), .ZN(n12385) );
  XNOR2_X1 U11669 ( .A(n12480), .B(n9242), .ZN(n9243) );
  NOR2_X1 U11670 ( .A1(n9243), .A2(n12747), .ZN(n9244) );
  AOI21_X1 U11671 ( .B1(n9243), .B2(n12747), .A(n9244), .ZN(n12483) );
  NAND2_X1 U11672 ( .A1(n9252), .A2(n15170), .ZN(n9246) );
  OAI22_X1 U11673 ( .A1(n9261), .A2(n9254), .B1(n9253), .B2(n9246), .ZN(n9247)
         );
  NAND2_X1 U11674 ( .A1(n9253), .A2(n10027), .ZN(n9248) );
  INV_X1 U11675 ( .A(n9249), .ZN(n9307) );
  NAND3_X1 U11676 ( .A1(n9250), .A2(n9307), .A3(n9766), .ZN(n9251) );
  AOI21_X1 U11677 ( .B1(n9253), .B2(n9252), .A(n9251), .ZN(n9257) );
  INV_X1 U11678 ( .A(n9254), .ZN(n9255) );
  NAND2_X1 U11679 ( .A1(n9261), .A2(n9255), .ZN(n9256) );
  AOI21_X1 U11680 ( .B1(n9257), .B2(n9256), .A(P3_U3151), .ZN(n9260) );
  NOR2_X1 U11681 ( .A1(n9767), .A2(n9993), .ZN(n9258) );
  AND2_X1 U11682 ( .A1(n9261), .A2(n9258), .ZN(n9259) );
  INV_X1 U11683 ( .A(n9261), .ZN(n9264) );
  NOR2_X1 U11684 ( .A1(n9767), .A2(n9262), .ZN(n9263) );
  AND2_X1 U11685 ( .A1(n9264), .A2(n9263), .ZN(n12496) );
  NAND2_X1 U11686 ( .A1(n12496), .A2(n13098), .ZN(n12474) );
  AOI22_X1 U11687 ( .A1(n12471), .A2(n12745), .B1(P3_REG3_REG_27__SCAN_IN), 
        .B2(P3_U3151), .ZN(n9265) );
  OAI21_X1 U11688 ( .B1(n9266), .B2(n12474), .A(n9265), .ZN(n9267) );
  AOI21_X1 U11689 ( .B1(n12883), .B2(n12497), .A(n9267), .ZN(n9268) );
  OAI21_X1 U11690 ( .B1(n12885), .B2(n12500), .A(n9268), .ZN(n9269) );
  NAND2_X1 U11691 ( .A1(n9271), .A2(n9270), .ZN(P3_U3154) );
  NOR2_X1 U11692 ( .A1(n9273), .A2(n9272), .ZN(n9643) );
  NOR2_X1 U11693 ( .A1(P1_IR_REG_6__SCAN_IN), .A2(P1_IR_REG_8__SCAN_IN), .ZN(
        n9274) );
  NOR2_X1 U11694 ( .A1(P1_IR_REG_12__SCAN_IN), .A2(P1_IR_REG_13__SCAN_IN), 
        .ZN(n9276) );
  NOR2_X1 U11695 ( .A1(P1_IR_REG_7__SCAN_IN), .A2(P1_IR_REG_14__SCAN_IN), .ZN(
        n9275) );
  AND2_X1 U11696 ( .A1(n9276), .A2(n9275), .ZN(n9278) );
  NOR2_X2 U11697 ( .A1(n9313), .A2(P1_IR_REG_3__SCAN_IN), .ZN(n9315) );
  AND2_X2 U11698 ( .A1(n9281), .A2(n9315), .ZN(n9302) );
  AND2_X2 U11699 ( .A1(n9294), .A2(n9285), .ZN(n9320) );
  AND2_X2 U11700 ( .A1(n9320), .A2(n9286), .ZN(n9287) );
  NAND2_X1 U11701 ( .A1(n9291), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9293) );
  NOR2_X1 U11702 ( .A1(P1_IR_REG_25__SCAN_IN), .A2(P1_IR_REG_24__SCAN_IN), 
        .ZN(n9297) );
  NOR2_X1 U11703 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(P1_IR_REG_23__SCAN_IN), 
        .ZN(n9296) );
  NAND4_X1 U11704 ( .A1(n9297), .A2(n9296), .A3(n9286), .A4(n9295), .ZN(n9299)
         );
  NOR2_X1 U11705 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P1_IR_REG_26__SCAN_IN), 
        .ZN(n9298) );
  NAND2_X1 U11706 ( .A1(n9336), .A2(n9298), .ZN(n9300) );
  NOR2_X1 U11707 ( .A1(n9300), .A2(n9299), .ZN(n9301) );
  INV_X1 U11708 ( .A(n9308), .ZN(n9310) );
  NAND2_X1 U11709 ( .A1(n6640), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9305) );
  XNOR2_X1 U11710 ( .A(n9305), .B(n9304), .ZN(n9500) );
  INV_X1 U11711 ( .A(n9486), .ZN(n9306) );
  NAND2_X1 U11712 ( .A1(n9310), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9312) );
  NAND2_X1 U11713 ( .A1(n9445), .A2(n11960), .ZN(n9319) );
  NAND2_X4 U11714 ( .A1(n11521), .A2(n9434), .ZN(n9371) );
  INV_X2 U11715 ( .A(n9371), .ZN(n11430) );
  NAND2_X1 U11716 ( .A1(n9313), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9314) );
  MUX2_X1 U11717 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9314), .S(
        P1_IR_REG_3__SCAN_IN), .Z(n9317) );
  INV_X1 U11718 ( .A(n9315), .ZN(n9316) );
  AND2_X1 U11719 ( .A1(n9317), .A2(n9316), .ZN(n9601) );
  AOI22_X1 U11720 ( .A1(n11430), .A2(P2_DATAO_REG_3__SCAN_IN), .B1(n6479), 
        .B2(n9601), .ZN(n9318) );
  NAND2_X1 U11721 ( .A1(n9319), .A2(n9318), .ZN(n9888) );
  NAND2_X1 U11722 ( .A1(n6668), .A2(n9320), .ZN(n9321) );
  NAND2_X1 U11723 ( .A1(n9321), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9322) );
  NAND2_X1 U11724 ( .A1(n9339), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9323) );
  INV_X1 U11725 ( .A(n11781), .ZN(n9324) );
  INV_X1 U11726 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n9422) );
  NAND2_X1 U11727 ( .A1(n6475), .A2(n9422), .ZN(n9333) );
  NAND2_X1 U11728 ( .A1(n10452), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n9332) );
  AND2_X2 U11729 ( .A1(n9328), .A2(n14294), .ZN(n11954) );
  NAND2_X1 U11730 ( .A1(n11954), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n9331) );
  AND2_X2 U11731 ( .A1(n9329), .A2(n14294), .ZN(n9377) );
  NAND2_X1 U11732 ( .A1(n9377), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n9330) );
  OAI22_X1 U11733 ( .A1(n10669), .A2(n9342), .B1(n12223), .B2(n9892), .ZN(
        n9341) );
  XNOR2_X2 U11734 ( .A(n9335), .B(P1_IR_REG_22__SCAN_IN), .ZN(n14297) );
  NAND2_X1 U11735 ( .A1(n14297), .A2(n14149), .ZN(n11778) );
  NAND2_X1 U11736 ( .A1(n11778), .A2(n11781), .ZN(n9355) );
  XNOR2_X1 U11737 ( .A(n9341), .B(n11452), .ZN(n10337) );
  OAI22_X1 U11738 ( .A1(n12276), .A2(n9892), .B1(n10669), .B2(n12223), .ZN(
        n10336) );
  XNOR2_X1 U11739 ( .A(n10337), .B(n10336), .ZN(n9410) );
  NAND2_X1 U11740 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(n14299), .ZN(n9343) );
  INV_X1 U11741 ( .A(n9372), .ZN(n9344) );
  OR2_X1 U11742 ( .A1(n11521), .A2(n9582), .ZN(n9345) );
  NAND2_X1 U11743 ( .A1(n11954), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n9347) );
  NAND2_X1 U11744 ( .A1(n9377), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n9346) );
  NAND2_X1 U11745 ( .A1(n10452), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n9349) );
  INV_X1 U11746 ( .A(n14187), .ZN(n9752) );
  OAI22_X1 U11747 ( .A1(n6906), .A2(n9342), .B1(n12223), .B2(n9752), .ZN(n9351) );
  XNOR2_X1 U11748 ( .A(n9351), .B(n11452), .ZN(n9353) );
  OAI22_X1 U11749 ( .A1(n12276), .A2(n9752), .B1(n6906), .B2(n12223), .ZN(
        n9352) );
  NOR2_X1 U11750 ( .A1(n9353), .A2(n9352), .ZN(n9369) );
  INV_X1 U11751 ( .A(SI_0_), .ZN(n9357) );
  OAI21_X1 U11752 ( .B1(n9438), .B2(n9357), .A(n9356), .ZN(n9358) );
  AND2_X1 U11753 ( .A1(n9359), .A2(n9358), .ZN(n14300) );
  MUX2_X1 U11754 ( .A(n14299), .B(n14300), .S(n11521), .Z(n14725) );
  INV_X1 U11755 ( .A(n14725), .ZN(n9656) );
  NAND2_X1 U11756 ( .A1(n6475), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n9363) );
  NAND2_X1 U11757 ( .A1(n10452), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n9362) );
  NAND2_X1 U11758 ( .A1(n11954), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n9361) );
  NAND2_X1 U11759 ( .A1(n9377), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n9360) );
  NAND2_X1 U11760 ( .A1(n10746), .A2(n13996), .ZN(n9365) );
  INV_X1 U11761 ( .A(n9412), .ZN(n9366) );
  NAND2_X1 U11762 ( .A1(n9366), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n9364) );
  OAI211_X1 U11763 ( .C1(n9342), .C2(n9656), .A(n9365), .B(n9364), .ZN(n9675)
         );
  OAI21_X1 U11764 ( .B1(n12273), .B2(n9675), .A(n9674), .ZN(n13857) );
  NAND2_X1 U11765 ( .A1(n13858), .A2(n13857), .ZN(n13856) );
  INV_X1 U11766 ( .A(n9369), .ZN(n9370) );
  NAND2_X1 U11767 ( .A1(n9449), .A2(n6564), .ZN(n9376) );
  INV_X1 U11768 ( .A(n9371), .ZN(n9374) );
  NAND2_X2 U11769 ( .A1(n9376), .A2(n9375), .ZN(n14728) );
  NAND2_X1 U11770 ( .A1(n6475), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n9381) );
  NAND2_X1 U11771 ( .A1(n10452), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n9380) );
  NAND2_X1 U11772 ( .A1(n11954), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n9379) );
  NAND2_X1 U11773 ( .A1(n9377), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n9378) );
  AOI22_X1 U11774 ( .A1(n12303), .A2(n14728), .B1(n10746), .B2(n13995), .ZN(
        n9382) );
  XNOR2_X1 U11775 ( .A(n9382), .B(n11452), .ZN(n9383) );
  INV_X1 U11776 ( .A(n13995), .ZN(n9750) );
  INV_X1 U11777 ( .A(n14728), .ZN(n10401) );
  OAI22_X1 U11778 ( .A1(n12276), .A2(n9750), .B1(n10401), .B2(n12223), .ZN(
        n9384) );
  INV_X1 U11779 ( .A(n9384), .ZN(n9385) );
  NAND2_X1 U11780 ( .A1(n9387), .A2(P1_B_REG_SCAN_IN), .ZN(n9388) );
  MUX2_X1 U11781 ( .A(P1_B_REG_SCAN_IN), .B(n9388), .S(n12150), .Z(n9390) );
  INV_X1 U11782 ( .A(n9389), .ZN(n9391) );
  NAND2_X1 U11783 ( .A1(n9390), .A2(n9391), .ZN(n9700) );
  OR2_X1 U11784 ( .A1(n9700), .A2(P1_D_REG_1__SCAN_IN), .ZN(n9392) );
  NAND2_X1 U11785 ( .A1(n9387), .A2(n9389), .ZN(n9483) );
  NOR4_X1 U11786 ( .A1(P1_D_REG_18__SCAN_IN), .A2(P1_D_REG_19__SCAN_IN), .A3(
        P1_D_REG_20__SCAN_IN), .A4(P1_D_REG_21__SCAN_IN), .ZN(n9396) );
  NOR4_X1 U11787 ( .A1(P1_D_REG_16__SCAN_IN), .A2(P1_D_REG_14__SCAN_IN), .A3(
        P1_D_REG_15__SCAN_IN), .A4(P1_D_REG_17__SCAN_IN), .ZN(n9395) );
  NOR4_X1 U11788 ( .A1(P1_D_REG_26__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n9394) );
  NOR4_X1 U11789 ( .A1(P1_D_REG_22__SCAN_IN), .A2(P1_D_REG_23__SCAN_IN), .A3(
        P1_D_REG_24__SCAN_IN), .A4(P1_D_REG_25__SCAN_IN), .ZN(n9393) );
  AND4_X1 U11790 ( .A1(n9396), .A2(n9395), .A3(n9394), .A4(n9393), .ZN(n9402)
         );
  NOR2_X1 U11791 ( .A1(P1_D_REG_2__SCAN_IN), .A2(P1_D_REG_3__SCAN_IN), .ZN(
        n9400) );
  NOR4_X1 U11792 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        P1_D_REG_4__SCAN_IN), .A4(P1_D_REG_5__SCAN_IN), .ZN(n9399) );
  NOR4_X1 U11793 ( .A1(P1_D_REG_10__SCAN_IN), .A2(P1_D_REG_11__SCAN_IN), .A3(
        P1_D_REG_12__SCAN_IN), .A4(P1_D_REG_13__SCAN_IN), .ZN(n9398) );
  NOR4_X1 U11794 ( .A1(P1_D_REG_6__SCAN_IN), .A2(P1_D_REG_7__SCAN_IN), .A3(
        P1_D_REG_8__SCAN_IN), .A4(P1_D_REG_9__SCAN_IN), .ZN(n9397) );
  AND4_X1 U11795 ( .A1(n9400), .A2(n9399), .A3(n9398), .A4(n9397), .ZN(n9401)
         );
  NAND2_X1 U11796 ( .A1(n9402), .A2(n9401), .ZN(n9698) );
  INV_X1 U11797 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n9488) );
  NOR2_X1 U11798 ( .A1(n9698), .A2(n9488), .ZN(n9403) );
  OR2_X1 U11799 ( .A1(n9700), .A2(n9403), .ZN(n9404) );
  NAND2_X1 U11800 ( .A1(n12150), .A2(n9389), .ZN(n9697) );
  AND2_X1 U11801 ( .A1(n9404), .A2(n9697), .ZN(n9670) );
  NAND2_X1 U11802 ( .A1(n10394), .A2(n9670), .ZN(n9417) );
  INV_X1 U11803 ( .A(n9417), .ZN(n9407) );
  NAND2_X1 U11804 ( .A1(n14724), .A2(n11978), .ZN(n10400) );
  NAND2_X1 U11805 ( .A1(n14297), .A2(n11965), .ZN(n11975) );
  INV_X1 U11806 ( .A(n11975), .ZN(n9501) );
  NOR2_X1 U11807 ( .A1(n14777), .A2(n9501), .ZN(n9405) );
  AND2_X1 U11808 ( .A1(n12057), .A2(n9405), .ZN(n9406) );
  INV_X1 U11809 ( .A(n9410), .ZN(n9408) );
  AOI211_X1 U11810 ( .C1(n9410), .C2(n9409), .A(n13938), .B(n6637), .ZN(n9433)
         );
  NAND2_X1 U11811 ( .A1(n9417), .A2(n9668), .ZN(n9413) );
  NAND2_X1 U11812 ( .A1(n14297), .A2(n12035), .ZN(n9411) );
  NAND2_X1 U11813 ( .A1(n11965), .A2(n11978), .ZN(n11958) );
  NAND2_X1 U11814 ( .A1(n14701), .A2(n9501), .ZN(n12055) );
  NAND3_X1 U11815 ( .A1(n9413), .A2(n9412), .A3(n12055), .ZN(n9414) );
  NAND2_X1 U11816 ( .A1(n9414), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9416) );
  INV_X1 U11817 ( .A(n9500), .ZN(n9415) );
  NAND2_X1 U11818 ( .A1(n9415), .A2(P1_STATE_REG_SCAN_IN), .ZN(n12060) );
  AND2_X1 U11819 ( .A1(n9416), .A2(n12060), .ZN(n14469) );
  INV_X1 U11820 ( .A(n14469), .ZN(n13955) );
  MUX2_X1 U11821 ( .A(n13955), .B(P1_U3086), .S(P1_REG3_REG_3__SCAN_IN), .Z(
        n9432) );
  INV_X1 U11822 ( .A(n12057), .ZN(n9499) );
  NOR2_X1 U11823 ( .A1(n9417), .A2(n9499), .ZN(n9419) );
  INV_X1 U11824 ( .A(n9419), .ZN(n9418) );
  INV_X1 U11825 ( .A(n9668), .ZN(n9696) );
  NAND2_X1 U11826 ( .A1(n9418), .A2(n14188), .ZN(n13946) );
  NAND2_X1 U11827 ( .A1(n10452), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n9427) );
  INV_X2 U11828 ( .A(n9420), .ZN(n11587) );
  NAND2_X1 U11829 ( .A1(n11587), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n9426) );
  INV_X1 U11830 ( .A(P1_REG3_REG_4__SCAN_IN), .ZN(n9421) );
  NAND2_X1 U11831 ( .A1(n9422), .A2(n9421), .ZN(n9423) );
  NAND2_X1 U11832 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n10439) );
  AND2_X1 U11833 ( .A1(n9423), .A2(n10439), .ZN(n10612) );
  NAND2_X1 U11834 ( .A1(n9893), .A2(n10612), .ZN(n9425) );
  NAND2_X1 U11835 ( .A1(n11526), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n9424) );
  NAND4_X1 U11836 ( .A1(n9427), .A2(n9426), .A3(n9425), .A4(n9424), .ZN(n13993) );
  INV_X1 U11837 ( .A(n9428), .ZN(n9586) );
  NAND2_X1 U11838 ( .A1(n13993), .A2(n14455), .ZN(n9430) );
  AND2_X2 U11839 ( .A1(n9501), .A2(n9586), .ZN(n14457) );
  NAND2_X1 U11840 ( .A1(n13995), .A2(n14457), .ZN(n9429) );
  AND2_X1 U11841 ( .A1(n9430), .A2(n9429), .ZN(n10668) );
  OAI22_X1 U11842 ( .A1(n13972), .A2(n10669), .B1(n13934), .B2(n10668), .ZN(
        n9431) );
  OR3_X1 U11843 ( .A1(n9433), .A2(n9432), .A3(n9431), .ZN(P1_U3218) );
  NAND2_X1 U11844 ( .A1(n9434), .A2(P1_U3086), .ZN(n14292) );
  NAND2_X1 U11845 ( .A1(n11519), .A2(P1_U3086), .ZN(n14296) );
  OAI222_X1 U11846 ( .A1(n14292), .A2(n9435), .B1(n12152), .B2(n9436), .C1(
        P1_U3086), .C2(n9582), .ZN(P1_U3354) );
  NOR2_X1 U11847 ( .A1(n9438), .A2(P2_STATE_REG_SCAN_IN), .ZN(n13813) );
  AND2_X1 U11848 ( .A1(n9438), .A2(P2_U3088), .ZN(n11266) );
  INV_X2 U11849 ( .A(n11266), .ZN(n13820) );
  OAI222_X1 U11850 ( .A1(n13822), .A2(n9437), .B1(n13820), .B2(n9436), .C1(
        P2_U3088), .C2(n9724), .ZN(P2_U3326) );
  OAI222_X1 U11851 ( .A1(P3_U3151), .A2(n10709), .B1(n13247), .B2(n9440), .C1(
        n13250), .C2(n9439), .ZN(P3_U3287) );
  OAI222_X1 U11852 ( .A1(P3_U3151), .A2(n9795), .B1(n13247), .B2(n9442), .C1(
        n13250), .C2(n9441), .ZN(P3_U3294) );
  OAI222_X1 U11853 ( .A1(P3_U3151), .A2(n11021), .B1(n13247), .B2(n9444), .C1(
        n13250), .C2(n9443), .ZN(P3_U3285) );
  INV_X1 U11854 ( .A(n9445), .ZN(n9466) );
  INV_X1 U11855 ( .A(n9728), .ZN(n13409) );
  OAI222_X1 U11856 ( .A1(n13822), .A2(n9446), .B1(n13820), .B2(n9466), .C1(
        P2_U3088), .C2(n13409), .ZN(P2_U3324) );
  INV_X1 U11857 ( .A(n10428), .ZN(n9463) );
  INV_X1 U11858 ( .A(n14819), .ZN(n9447) );
  OAI222_X1 U11859 ( .A1(n13822), .A2(n9448), .B1(n13820), .B2(n9463), .C1(
        P2_U3088), .C2(n9447), .ZN(P2_U3322) );
  INV_X1 U11860 ( .A(n9449), .ZN(n9460) );
  OAI222_X1 U11861 ( .A1(n13822), .A2(n9450), .B1(n13820), .B2(n9460), .C1(
        P2_U3088), .C2(n8059), .ZN(P2_U3325) );
  INV_X1 U11862 ( .A(n10433), .ZN(n9471) );
  INV_X1 U11863 ( .A(n9733), .ZN(n13433) );
  OAI222_X1 U11864 ( .A1(n13822), .A2(n9451), .B1(n13820), .B2(n9471), .C1(
        P2_U3088), .C2(n13433), .ZN(P2_U3321) );
  INV_X1 U11865 ( .A(n9884), .ZN(n9474) );
  OAI222_X1 U11866 ( .A1(n13822), .A2(n9452), .B1(n13820), .B2(n9474), .C1(
        P2_U3088), .C2(n13421), .ZN(P2_U3323) );
  INV_X1 U11867 ( .A(n13238), .ZN(n9456) );
  NAND2_X1 U11868 ( .A1(n9453), .A2(n9456), .ZN(n9454) );
  OAI21_X1 U11869 ( .B1(n9456), .B2(n9455), .A(n9454), .ZN(P3_U3377) );
  OAI222_X1 U11870 ( .A1(n10155), .A2(P3_U3151), .B1(n13250), .B2(n9458), .C1(
        n9457), .C2(n13247), .ZN(P3_U3289) );
  INV_X1 U11871 ( .A(n14292), .ZN(n14289) );
  INV_X1 U11872 ( .A(n14289), .ZN(n11652) );
  INV_X1 U11873 ( .A(n6470), .ZN(n9459) );
  OAI222_X1 U11874 ( .A1(n11652), .A2(n9461), .B1(n12152), .B2(n9460), .C1(
        P1_U3086), .C2(n9459), .ZN(P1_U3353) );
  OR2_X1 U11875 ( .A1(n9469), .A2(n10128), .ZN(n9462) );
  XNOR2_X1 U11876 ( .A(n9462), .B(P1_IR_REG_5__SCAN_IN), .ZN(n10429) );
  INV_X1 U11877 ( .A(n10429), .ZN(n9628) );
  OAI222_X1 U11878 ( .A1(n11652), .A2(n9464), .B1(n12152), .B2(n9463), .C1(
        P1_U3086), .C2(n9628), .ZN(P1_U3350) );
  INV_X1 U11879 ( .A(n9601), .ZN(n9465) );
  OAI222_X1 U11880 ( .A1(n11652), .A2(n9467), .B1(n14296), .B2(n9466), .C1(
        P1_U3086), .C2(n9465), .ZN(P1_U3352) );
  NAND2_X1 U11881 ( .A1(n9469), .A2(n9468), .ZN(n9476) );
  NAND2_X1 U11882 ( .A1(n9476), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9470) );
  XNOR2_X1 U11883 ( .A(n9470), .B(P1_IR_REG_6__SCAN_IN), .ZN(n10434) );
  OAI222_X1 U11884 ( .A1(n11652), .A2(n9472), .B1(n14296), .B2(n9471), .C1(
        P1_U3086), .C2(n6869), .ZN(P1_U3349) );
  NAND2_X1 U11885 ( .A1(n9316), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9473) );
  XNOR2_X1 U11886 ( .A(n9473), .B(P1_IR_REG_4__SCAN_IN), .ZN(n9885) );
  INV_X1 U11887 ( .A(n9885), .ZN(n9857) );
  OAI222_X1 U11888 ( .A1(n11652), .A2(n9475), .B1(n14296), .B2(n9474), .C1(
        P1_U3086), .C2(n9857), .ZN(P1_U3351) );
  INV_X1 U11889 ( .A(n10448), .ZN(n9481) );
  NAND2_X1 U11890 ( .A1(n9513), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9477) );
  XNOR2_X1 U11891 ( .A(n9477), .B(P1_IR_REG_7__SCAN_IN), .ZN(n10449) );
  INV_X1 U11892 ( .A(n10449), .ZN(n9478) );
  OAI222_X1 U11893 ( .A1(n11652), .A2(n9479), .B1(n14296), .B2(n9481), .C1(
        P1_U3086), .C2(n9478), .ZN(P1_U3348) );
  INV_X1 U11894 ( .A(n13444), .ZN(n9480) );
  OAI222_X1 U11895 ( .A1(n13822), .A2(n9482), .B1(n13820), .B2(n9481), .C1(
        P2_U3088), .C2(n9480), .ZN(P2_U3320) );
  NAND2_X1 U11896 ( .A1(n9700), .A2(n12057), .ZN(n14718) );
  INV_X1 U11897 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n9485) );
  INV_X1 U11898 ( .A(n9483), .ZN(n9484) );
  AOI22_X1 U11899 ( .A1(n14718), .A2(n9485), .B1(n9484), .B2(n9486), .ZN(
        P1_U3446) );
  INV_X1 U11900 ( .A(n9697), .ZN(n9487) );
  AOI22_X1 U11901 ( .A1(n14718), .A2(n9488), .B1(n9487), .B2(n9486), .ZN(
        P1_U3445) );
  OAI222_X1 U11902 ( .A1(n13250), .A2(n9490), .B1(n12773), .B2(P3_U3151), .C1(
        n9489), .C2(n13247), .ZN(P3_U3283) );
  INV_X1 U11903 ( .A(n13247), .ZN(n14316) );
  AOI222_X1 U11904 ( .A1(n9491), .A2(n14317), .B1(SI_5_), .B2(n14316), .C1(
        P3_STATE_REG_SCAN_IN), .C2(n15069), .ZN(n9492) );
  INV_X1 U11905 ( .A(n9492), .ZN(P3_U3290) );
  AOI222_X1 U11906 ( .A1(n9493), .A2(n14317), .B1(SI_9_), .B2(n14316), .C1(
        P3_STATE_REG_SCAN_IN), .C2(n10714), .ZN(n9494) );
  INV_X1 U11907 ( .A(n9494), .ZN(P3_U3286) );
  AOI222_X1 U11908 ( .A1(n9495), .A2(n14317), .B1(SI_7_), .B2(n14316), .C1(
        P3_STATE_REG_SCAN_IN), .C2(n10269), .ZN(n9496) );
  INV_X1 U11909 ( .A(n9496), .ZN(P3_U3288) );
  AOI222_X1 U11910 ( .A1(n9497), .A2(n14317), .B1(SI_4_), .B2(n14316), .C1(
        P3_STATE_REG_SCAN_IN), .C2(n10091), .ZN(n9498) );
  INV_X1 U11911 ( .A(n9498), .ZN(P3_U3291) );
  NAND2_X1 U11912 ( .A1(n9499), .A2(n12060), .ZN(n9505) );
  NAND2_X1 U11913 ( .A1(n9501), .A2(n9500), .ZN(n9502) );
  NAND2_X1 U11914 ( .A1(n9502), .A2(n11521), .ZN(n9503) );
  INV_X1 U11915 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n9511) );
  INV_X1 U11916 ( .A(n9503), .ZN(n9504) );
  NAND2_X1 U11917 ( .A1(n9505), .A2(n9504), .ZN(n9587) );
  INV_X1 U11918 ( .A(n9587), .ZN(n9579) );
  INV_X1 U11919 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n9507) );
  OAI21_X1 U11920 ( .B1(n6484), .B2(P1_REG2_REG_0__SCAN_IN), .A(n9586), .ZN(
        n9849) );
  AOI21_X1 U11921 ( .B1(n6484), .B2(n9507), .A(n9849), .ZN(n9508) );
  INV_X1 U11922 ( .A(n14299), .ZN(n9850) );
  XNOR2_X1 U11923 ( .A(n9508), .B(n9850), .ZN(n9509) );
  AOI22_X1 U11924 ( .A1(n9579), .A2(n9509), .B1(P1_REG3_REG_0__SCAN_IN), .B2(
        P1_U3086), .ZN(n9510) );
  OAI21_X1 U11925 ( .B1(n14661), .B2(n9511), .A(n9510), .ZN(P1_U3243) );
  INV_X1 U11926 ( .A(n10461), .ZN(n9516) );
  INV_X1 U11927 ( .A(n9736), .ZN(n14833) );
  OAI222_X1 U11928 ( .A1(n13822), .A2(n9512), .B1(n13820), .B2(n9516), .C1(
        P2_U3088), .C2(n14833), .ZN(P2_U3319) );
  NAND2_X1 U11929 ( .A1(n9519), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9514) );
  XNOR2_X1 U11930 ( .A(n9514), .B(P1_IR_REG_8__SCAN_IN), .ZN(n10462) );
  INV_X1 U11931 ( .A(n10462), .ZN(n9515) );
  OAI222_X1 U11932 ( .A1(n11652), .A2(n9517), .B1(n14296), .B2(n9516), .C1(
        P1_U3086), .C2(n9515), .ZN(P1_U3347) );
  INV_X1 U11933 ( .A(n14661), .ZN(n14003) );
  NOR2_X1 U11934 ( .A1(n14003), .A2(P1_U4016), .ZN(P1_U3085) );
  INV_X1 U11935 ( .A(n10562), .ZN(n9523) );
  INV_X1 U11936 ( .A(n14846), .ZN(n9738) );
  OAI222_X1 U11937 ( .A1(n13822), .A2(n9518), .B1(n13820), .B2(n9523), .C1(
        P2_U3088), .C2(n9738), .ZN(P2_U3318) );
  INV_X1 U11938 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n9520) );
  OR2_X1 U11939 ( .A1(n9571), .A2(n9520), .ZN(n9521) );
  NAND2_X1 U11940 ( .A1(n9571), .A2(n9520), .ZN(n9560) );
  INV_X1 U11941 ( .A(n10563), .ZN(n9522) );
  OAI222_X1 U11942 ( .A1(n11652), .A2(n9524), .B1(n14296), .B2(n9523), .C1(
        P1_U3086), .C2(n9522), .ZN(P1_U3346) );
  NOR2_X1 U11943 ( .A1(n13238), .A2(n9525), .ZN(n9527) );
  CLKBUF_X1 U11944 ( .A(n9527), .Z(n9557) );
  INV_X1 U11945 ( .A(P3_D_REG_17__SCAN_IN), .ZN(n9526) );
  NOR2_X1 U11946 ( .A1(n9557), .A2(n9526), .ZN(P3_U3248) );
  INV_X1 U11947 ( .A(P3_D_REG_3__SCAN_IN), .ZN(n9528) );
  NOR2_X1 U11948 ( .A1(n9557), .A2(n9528), .ZN(P3_U3262) );
  INV_X1 U11949 ( .A(P3_D_REG_26__SCAN_IN), .ZN(n9529) );
  NOR2_X1 U11950 ( .A1(n9527), .A2(n9529), .ZN(P3_U3239) );
  INV_X1 U11951 ( .A(P3_D_REG_24__SCAN_IN), .ZN(n9530) );
  NOR2_X1 U11952 ( .A1(n9527), .A2(n9530), .ZN(P3_U3241) );
  INV_X1 U11953 ( .A(P3_D_REG_2__SCAN_IN), .ZN(n9531) );
  NOR2_X1 U11954 ( .A1(n9557), .A2(n9531), .ZN(P3_U3263) );
  INV_X1 U11955 ( .A(P3_D_REG_20__SCAN_IN), .ZN(n9532) );
  NOR2_X1 U11956 ( .A1(n9527), .A2(n9532), .ZN(P3_U3245) );
  INV_X1 U11957 ( .A(P3_D_REG_25__SCAN_IN), .ZN(n9533) );
  NOR2_X1 U11958 ( .A1(n9527), .A2(n9533), .ZN(P3_U3240) );
  INV_X1 U11959 ( .A(P3_D_REG_18__SCAN_IN), .ZN(n9534) );
  NOR2_X1 U11960 ( .A1(n9557), .A2(n9534), .ZN(P3_U3247) );
  INV_X1 U11961 ( .A(P3_D_REG_11__SCAN_IN), .ZN(n9535) );
  NOR2_X1 U11962 ( .A1(n9557), .A2(n9535), .ZN(P3_U3254) );
  INV_X1 U11963 ( .A(P3_D_REG_31__SCAN_IN), .ZN(n9536) );
  NOR2_X1 U11964 ( .A1(n9527), .A2(n9536), .ZN(P3_U3234) );
  INV_X1 U11965 ( .A(P3_D_REG_21__SCAN_IN), .ZN(n9537) );
  NOR2_X1 U11966 ( .A1(n9527), .A2(n9537), .ZN(P3_U3244) );
  INV_X1 U11967 ( .A(P3_D_REG_29__SCAN_IN), .ZN(n9538) );
  NOR2_X1 U11968 ( .A1(n9527), .A2(n9538), .ZN(P3_U3236) );
  INV_X1 U11969 ( .A(P3_D_REG_28__SCAN_IN), .ZN(n9539) );
  NOR2_X1 U11970 ( .A1(n9527), .A2(n9539), .ZN(P3_U3237) );
  INV_X1 U11971 ( .A(P3_D_REG_27__SCAN_IN), .ZN(n9540) );
  NOR2_X1 U11972 ( .A1(n9527), .A2(n9540), .ZN(P3_U3238) );
  INV_X1 U11973 ( .A(P3_D_REG_5__SCAN_IN), .ZN(n9541) );
  NOR2_X1 U11974 ( .A1(n9527), .A2(n9541), .ZN(P3_U3260) );
  INV_X1 U11975 ( .A(P3_D_REG_10__SCAN_IN), .ZN(n9542) );
  NOR2_X1 U11976 ( .A1(n9557), .A2(n9542), .ZN(P3_U3255) );
  INV_X1 U11977 ( .A(P3_D_REG_9__SCAN_IN), .ZN(n9543) );
  NOR2_X1 U11978 ( .A1(n9557), .A2(n9543), .ZN(P3_U3256) );
  INV_X1 U11979 ( .A(P3_D_REG_23__SCAN_IN), .ZN(n9544) );
  NOR2_X1 U11980 ( .A1(n9527), .A2(n9544), .ZN(P3_U3242) );
  INV_X1 U11981 ( .A(P3_D_REG_4__SCAN_IN), .ZN(n9545) );
  NOR2_X1 U11982 ( .A1(n9557), .A2(n9545), .ZN(P3_U3261) );
  INV_X1 U11983 ( .A(P3_D_REG_6__SCAN_IN), .ZN(n9546) );
  NOR2_X1 U11984 ( .A1(n9557), .A2(n9546), .ZN(P3_U3259) );
  INV_X1 U11985 ( .A(P3_D_REG_30__SCAN_IN), .ZN(n9547) );
  NOR2_X1 U11986 ( .A1(n9557), .A2(n9547), .ZN(P3_U3235) );
  INV_X1 U11987 ( .A(P3_D_REG_22__SCAN_IN), .ZN(n9548) );
  NOR2_X1 U11988 ( .A1(n9557), .A2(n9548), .ZN(P3_U3243) );
  INV_X1 U11989 ( .A(P3_D_REG_19__SCAN_IN), .ZN(n9549) );
  NOR2_X1 U11990 ( .A1(n9557), .A2(n9549), .ZN(P3_U3246) );
  INV_X1 U11991 ( .A(P3_D_REG_14__SCAN_IN), .ZN(n9550) );
  NOR2_X1 U11992 ( .A1(n9557), .A2(n9550), .ZN(P3_U3251) );
  INV_X1 U11993 ( .A(P3_D_REG_13__SCAN_IN), .ZN(n9551) );
  NOR2_X1 U11994 ( .A1(n9557), .A2(n9551), .ZN(P3_U3252) );
  INV_X1 U11995 ( .A(P3_D_REG_12__SCAN_IN), .ZN(n9552) );
  NOR2_X1 U11996 ( .A1(n9557), .A2(n9552), .ZN(P3_U3253) );
  INV_X1 U11997 ( .A(P3_D_REG_7__SCAN_IN), .ZN(n9553) );
  NOR2_X1 U11998 ( .A1(n9557), .A2(n9553), .ZN(P3_U3258) );
  INV_X1 U11999 ( .A(P3_D_REG_16__SCAN_IN), .ZN(n9554) );
  NOR2_X1 U12000 ( .A1(n9557), .A2(n9554), .ZN(P3_U3249) );
  INV_X1 U12001 ( .A(P3_D_REG_8__SCAN_IN), .ZN(n9555) );
  NOR2_X1 U12002 ( .A1(n9557), .A2(n9555), .ZN(P3_U3257) );
  INV_X1 U12003 ( .A(P3_D_REG_15__SCAN_IN), .ZN(n9556) );
  NOR2_X1 U12004 ( .A1(n9557), .A2(n9556), .ZN(P3_U3250) );
  INV_X1 U12005 ( .A(n10568), .ZN(n9563) );
  INV_X1 U12006 ( .A(n14863), .ZN(n9558) );
  OAI222_X1 U12007 ( .A1(n13822), .A2(n9559), .B1(n13820), .B2(n9563), .C1(
        P2_U3088), .C2(n9558), .ZN(P2_U3317) );
  NAND2_X1 U12008 ( .A1(n9560), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9561) );
  XNOR2_X1 U12009 ( .A(n9561), .B(P1_IR_REG_10__SCAN_IN), .ZN(n11411) );
  INV_X1 U12010 ( .A(n11411), .ZN(n9562) );
  OAI222_X1 U12011 ( .A1(n11652), .A2(n9564), .B1(n12152), .B2(n9563), .C1(
        P1_U3086), .C2(n9562), .ZN(P1_U3345) );
  OAI222_X1 U12012 ( .A1(P3_U3151), .A2(n12793), .B1(n13247), .B2(n9566), .C1(
        n13250), .C2(n9565), .ZN(P3_U3282) );
  INV_X1 U12013 ( .A(n10939), .ZN(n9573) );
  INV_X1 U12014 ( .A(n9866), .ZN(n9567) );
  OAI222_X1 U12015 ( .A1(n13822), .A2(n9568), .B1(n13820), .B2(n9573), .C1(
        P2_U3088), .C2(n9567), .ZN(P2_U3316) );
  OR2_X1 U12016 ( .A1(n9569), .A2(n10128), .ZN(n9570) );
  NAND2_X1 U12017 ( .A1(n9571), .A2(n9570), .ZN(n9611) );
  INV_X1 U12018 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n9572) );
  XNOR2_X1 U12019 ( .A(n9611), .B(n9572), .ZN(n11413) );
  OAI222_X1 U12020 ( .A1(n9574), .A2(n14292), .B1(P1_U3086), .B2(n6856), .C1(
        n12152), .C2(n9573), .ZN(P1_U3344) );
  OAI222_X1 U12021 ( .A1(n12790), .A2(P3_U3151), .B1(n13250), .B2(n9575), .C1(
        n6890), .C2(n13247), .ZN(P3_U3281) );
  INV_X1 U12022 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n9576) );
  MUX2_X1 U12023 ( .A(P1_REG2_REG_2__SCAN_IN), .B(n9576), .S(n14012), .Z(
        n14016) );
  AND2_X1 U12024 ( .A1(n14299), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n14001) );
  NAND2_X1 U12025 ( .A1(n14002), .A2(n14001), .ZN(n14000) );
  INV_X1 U12026 ( .A(n9582), .ZN(n14004) );
  NAND2_X1 U12027 ( .A1(n14004), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n9577) );
  NAND2_X1 U12028 ( .A1(n14000), .A2(n9577), .ZN(n14015) );
  AND2_X1 U12029 ( .A1(n14016), .A2(n14015), .ZN(n14013) );
  AOI21_X1 U12030 ( .B1(n6470), .B2(P1_REG2_REG_2__SCAN_IN), .A(n14013), .ZN(
        n9581) );
  XNOR2_X1 U12031 ( .A(n9601), .B(P1_REG2_REG_3__SCAN_IN), .ZN(n9580) );
  NOR2_X1 U12032 ( .A1(n9581), .A2(n9580), .ZN(n9593) );
  NOR2_X1 U12033 ( .A1(n9428), .A2(n6484), .ZN(n9578) );
  AOI211_X1 U12034 ( .C1(n9581), .C2(n9580), .A(n9593), .B(n14651), .ZN(n9592)
         );
  INV_X1 U12035 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n14789) );
  MUX2_X1 U12036 ( .A(P1_REG1_REG_2__SCAN_IN), .B(n14789), .S(n6470), .Z(
        n14020) );
  XNOR2_X1 U12037 ( .A(n9582), .B(P1_REG1_REG_1__SCAN_IN), .ZN(n13999) );
  AND2_X1 U12038 ( .A1(n14299), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n13998) );
  NAND2_X1 U12039 ( .A1(n13999), .A2(n13998), .ZN(n13997) );
  NAND2_X1 U12040 ( .A1(n14004), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n9583) );
  NAND2_X1 U12041 ( .A1(n13997), .A2(n9583), .ZN(n14019) );
  AND2_X1 U12042 ( .A1(n14020), .A2(n14019), .ZN(n14017) );
  XNOR2_X1 U12043 ( .A(n9601), .B(P1_REG1_REG_3__SCAN_IN), .ZN(n9584) );
  INV_X1 U12044 ( .A(n6484), .ZN(n12056) );
  AOI211_X1 U12045 ( .C1(n9585), .C2(n9584), .A(n9600), .B(n14647), .ZN(n9591)
         );
  NAND2_X1 U12046 ( .A1(n14658), .A2(n9601), .ZN(n9589) );
  NAND2_X1 U12047 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_U3086), .ZN(n9588) );
  OAI211_X1 U12048 ( .C1(n6819), .C2(n14661), .A(n9589), .B(n9588), .ZN(n9590)
         );
  OR3_X1 U12049 ( .A1(n9592), .A2(n9591), .A3(n9590), .ZN(P1_U3246) );
  XNOR2_X1 U12050 ( .A(n9885), .B(P1_REG2_REG_4__SCAN_IN), .ZN(n9854) );
  INV_X1 U12051 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n9594) );
  MUX2_X1 U12052 ( .A(P1_REG2_REG_5__SCAN_IN), .B(n9594), .S(n10429), .Z(n9595) );
  INV_X1 U12053 ( .A(n9595), .ZN(n9621) );
  AOI21_X1 U12054 ( .B1(P1_REG2_REG_5__SCAN_IN), .B2(n10429), .A(n9620), .ZN(
        n9599) );
  INV_X1 U12055 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n9596) );
  MUX2_X1 U12056 ( .A(P1_REG2_REG_6__SCAN_IN), .B(n9596), .S(n10434), .Z(n9597) );
  INV_X1 U12057 ( .A(n9597), .ZN(n9598) );
  NOR2_X1 U12058 ( .A1(n9599), .A2(n9598), .ZN(n9681) );
  AOI211_X1 U12059 ( .C1(n9599), .C2(n9598), .A(n14651), .B(n9681), .ZN(n9610)
         );
  MUX2_X1 U12060 ( .A(n6868), .B(P1_REG1_REG_6__SCAN_IN), .S(n10434), .Z(n9604) );
  XNOR2_X1 U12061 ( .A(n9885), .B(P1_REG1_REG_4__SCAN_IN), .ZN(n9851) );
  AOI21_X1 U12062 ( .B1(n9885), .B2(P1_REG1_REG_4__SCAN_IN), .A(n6516), .ZN(
        n9619) );
  INV_X1 U12063 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n9602) );
  MUX2_X1 U12064 ( .A(P1_REG1_REG_5__SCAN_IN), .B(n9602), .S(n10429), .Z(n9618) );
  NAND2_X1 U12065 ( .A1(n9619), .A2(n9618), .ZN(n9617) );
  OAI21_X1 U12066 ( .B1(n10429), .B2(P1_REG1_REG_5__SCAN_IN), .A(n9617), .ZN(
        n9603) );
  NOR2_X1 U12067 ( .A1(n9603), .A2(n9604), .ZN(n9686) );
  AOI211_X1 U12068 ( .C1(n9604), .C2(n9603), .A(n14647), .B(n9686), .ZN(n9609)
         );
  NAND2_X1 U12069 ( .A1(n14658), .A2(n10434), .ZN(n9606) );
  NAND2_X1 U12070 ( .A1(P1_REG3_REG_6__SCAN_IN), .A2(P1_U3086), .ZN(n9605) );
  OAI211_X1 U12071 ( .C1(n9607), .C2(n14661), .A(n9606), .B(n9605), .ZN(n9608)
         );
  OR3_X1 U12072 ( .A1(n9610), .A2(n9609), .A3(n9608), .ZN(P1_U3249) );
  INV_X1 U12073 ( .A(n10943), .ZN(n9615) );
  NAND2_X1 U12074 ( .A1(n9612), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9632) );
  XNOR2_X1 U12075 ( .A(n9632), .B(P1_IR_REG_12__SCAN_IN), .ZN(n14582) );
  INV_X1 U12076 ( .A(n14582), .ZN(n11401) );
  OAI222_X1 U12077 ( .A1(n11652), .A2(n9613), .B1(n12152), .B2(n9615), .C1(
        n11401), .C2(P1_U3086), .ZN(P1_U3343) );
  INV_X1 U12078 ( .A(n10925), .ZN(n9614) );
  OAI222_X1 U12079 ( .A1(n13822), .A2(n9616), .B1(n13820), .B2(n9615), .C1(
        n9614), .C2(P2_U3088), .ZN(P2_U3315) );
  OAI21_X1 U12080 ( .B1(n9619), .B2(n9618), .A(n9617), .ZN(n9624) );
  AOI211_X1 U12081 ( .C1(n9622), .C2(n9621), .A(n9620), .B(n14651), .ZN(n9623)
         );
  AOI21_X1 U12082 ( .B1(n14633), .B2(n9624), .A(n9623), .ZN(n9627) );
  NAND2_X1 U12083 ( .A1(P1_U3086), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n10642) );
  INV_X1 U12084 ( .A(n10642), .ZN(n9625) );
  AOI21_X1 U12085 ( .B1(n14003), .B2(P1_ADDR_REG_5__SCAN_IN), .A(n9625), .ZN(
        n9626) );
  OAI211_X1 U12086 ( .C1(n9628), .C2(n14642), .A(n9627), .B(n9626), .ZN(
        P1_U3248) );
  INV_X1 U12087 ( .A(n10981), .ZN(n9637) );
  INV_X1 U12088 ( .A(n14875), .ZN(n9629) );
  OAI222_X1 U12089 ( .A1(n13822), .A2(n9630), .B1(n13820), .B2(n9637), .C1(
        n9629), .C2(P2_U3088), .ZN(P2_U3314) );
  INV_X1 U12090 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n9631) );
  AOI21_X1 U12091 ( .B1(n9632), .B2(n9631), .A(n10128), .ZN(n9633) );
  NAND2_X1 U12092 ( .A1(n9633), .A2(P1_IR_REG_13__SCAN_IN), .ZN(n9636) );
  INV_X1 U12093 ( .A(n9633), .ZN(n9635) );
  INV_X1 U12094 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n9634) );
  NAND2_X1 U12095 ( .A1(n9635), .A2(n9634), .ZN(n9877) );
  INV_X1 U12096 ( .A(n11416), .ZN(n14598) );
  OAI222_X1 U12097 ( .A1(n11652), .A2(n10982), .B1(n12152), .B2(n9637), .C1(
        n14598), .C2(P1_U3086), .ZN(P1_U3342) );
  OAI222_X1 U12098 ( .A1(P3_U3151), .A2(n12818), .B1(n13247), .B2(n9639), .C1(
        n13250), .C2(n9638), .ZN(P3_U3280) );
  AOI21_X1 U12099 ( .B1(n9824), .B2(n9641), .A(n9640), .ZN(n9642) );
  OR2_X1 U12100 ( .A1(n9643), .A2(n9642), .ZN(n9648) );
  NOR2_X1 U12101 ( .A1(n8822), .A2(P2_U3088), .ZN(n13812) );
  NAND2_X1 U12102 ( .A1(n9648), .A2(n13812), .ZN(n9644) );
  INV_X1 U12103 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n9645) );
  OAI22_X1 U12104 ( .A1(n9646), .A2(n14884), .B1(n14880), .B2(n9645), .ZN(
        n9651) );
  NAND2_X1 U12105 ( .A1(n14913), .A2(n9646), .ZN(n9649) );
  AND2_X1 U12106 ( .A1(n8822), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9647) );
  AND2_X1 U12107 ( .A1(n9648), .A2(n9647), .ZN(n14890) );
  OAI211_X1 U12108 ( .C1(P2_REG2_REG_0__SCAN_IN), .C2(n14880), .A(n9649), .B(
        n14922), .ZN(n9650) );
  MUX2_X1 U12109 ( .A(n9651), .B(n9650), .S(P2_IR_REG_0__SCAN_IN), .Z(n9652)
         );
  INV_X1 U12110 ( .A(n9652), .ZN(n9654) );
  NAND2_X1 U12111 ( .A1(P2_U3088), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n9653) );
  OAI211_X1 U12112 ( .C1(n15198), .C2(n14926), .A(n9654), .B(n9653), .ZN(
        P2_U3214) );
  INV_X1 U12113 ( .A(n14297), .ZN(n11973) );
  INV_X1 U12114 ( .A(n11777), .ZN(n9655) );
  NAND2_X1 U12115 ( .A1(n9655), .A2(n11972), .ZN(n14730) );
  INV_X1 U12116 ( .A(n14730), .ZN(n14759) );
  XNOR2_X2 U12117 ( .A(n14187), .B(n6473), .ZN(n11998) );
  OR2_X1 U12118 ( .A1(n11775), .A2(n9656), .ZN(n9658) );
  NAND2_X1 U12119 ( .A1(n9657), .A2(n9658), .ZN(n9754) );
  INV_X1 U12120 ( .A(n9658), .ZN(n9659) );
  NAND2_X1 U12121 ( .A1(n9659), .A2(n11998), .ZN(n9660) );
  NAND2_X1 U12122 ( .A1(n9754), .A2(n9660), .ZN(n14177) );
  NAND2_X1 U12123 ( .A1(n6473), .A2(n14725), .ZN(n9661) );
  AND2_X1 U12124 ( .A1(n10396), .A2(n9661), .ZN(n14180) );
  INV_X1 U12125 ( .A(n14180), .ZN(n9662) );
  OAI22_X1 U12126 ( .A1(n14753), .A2(n6906), .B1(n9662), .B2(n14493), .ZN(
        n9667) );
  XNOR2_X1 U12127 ( .A(n14180), .B(n14187), .ZN(n9663) );
  MUX2_X1 U12128 ( .A(n9663), .B(n11998), .S(n13996), .Z(n9666) );
  OAI21_X1 U12129 ( .B1(n11778), .B2(n11781), .A(n11452), .ZN(n10471) );
  INV_X1 U12130 ( .A(n11636), .ZN(n14743) );
  NAND2_X1 U12131 ( .A1(n14177), .A2(n14743), .ZN(n9665) );
  AOI22_X1 U12132 ( .A1(n13996), .A2(n14457), .B1(n14455), .B2(n13995), .ZN(
        n9664) );
  OAI211_X1 U12133 ( .C1(n14780), .C2(n9666), .A(n9665), .B(n9664), .ZN(n14178) );
  AOI211_X1 U12134 ( .C1(n14759), .C2(n14177), .A(n9667), .B(n14178), .ZN(
        n9705) );
  AND3_X1 U12135 ( .A1(n12057), .A2(n9668), .A3(n12055), .ZN(n9669) );
  AND2_X1 U12136 ( .A1(n9670), .A2(n9669), .ZN(n9672) );
  NAND2_X1 U12137 ( .A1(n14797), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n9673) );
  OAI21_X1 U12138 ( .B1(n9705), .B2(n14797), .A(n9673), .ZN(P1_U3529) );
  NAND2_X1 U12139 ( .A1(n14466), .A2(n14455), .ZN(n12312) );
  AOI22_X1 U12140 ( .A1(n13969), .A2(n14187), .B1(n14463), .B2(n14725), .ZN(
        n9678) );
  OAI21_X1 U12141 ( .B1(n9676), .B2(n9675), .A(n9674), .ZN(n9845) );
  NAND2_X1 U12142 ( .A1(n13946), .A2(n12055), .ZN(n13925) );
  AOI22_X1 U12143 ( .A1(n9845), .A2(n14465), .B1(P1_REG3_REG_0__SCAN_IN), .B2(
        n13925), .ZN(n9677) );
  NAND2_X1 U12144 ( .A1(n9678), .A2(n9677), .ZN(P1_U3232) );
  OAI222_X1 U12145 ( .A1(n13250), .A2(n9680), .B1(n12842), .B2(P3_U3151), .C1(
        n9679), .C2(n13247), .ZN(P3_U3279) );
  AOI21_X1 U12146 ( .B1(n10434), .B2(P1_REG2_REG_6__SCAN_IN), .A(n9681), .ZN(
        n9685) );
  INV_X1 U12147 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n9682) );
  MUX2_X1 U12148 ( .A(P1_REG2_REG_7__SCAN_IN), .B(n9682), .S(n10449), .Z(n9683) );
  INV_X1 U12149 ( .A(n9683), .ZN(n9684) );
  NOR2_X1 U12150 ( .A1(n9685), .A2(n9684), .ZN(n9976) );
  AOI211_X1 U12151 ( .C1(n9685), .C2(n9684), .A(n14651), .B(n9976), .ZN(n9695)
         );
  INV_X1 U12152 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n9687) );
  MUX2_X1 U12153 ( .A(n9687), .B(P1_REG1_REG_7__SCAN_IN), .S(n10449), .Z(n9688) );
  AOI211_X1 U12154 ( .C1(n9689), .C2(n9688), .A(n14647), .B(n9969), .ZN(n9694)
         );
  NAND2_X1 U12155 ( .A1(n14658), .A2(n10449), .ZN(n9691) );
  NAND2_X1 U12156 ( .A1(P1_REG3_REG_7__SCAN_IN), .A2(P1_U3086), .ZN(n9690) );
  OAI211_X1 U12157 ( .C1(n9692), .C2(n14661), .A(n9691), .B(n9690), .ZN(n9693)
         );
  OR3_X1 U12158 ( .A1(n9695), .A2(n9694), .A3(n9693), .ZN(P1_U3250) );
  NOR2_X1 U12159 ( .A1(n10394), .A2(n9696), .ZN(n9704) );
  OAI21_X1 U12160 ( .B1(n9700), .B2(P1_D_REG_0__SCAN_IN), .A(n9697), .ZN(n9703) );
  AND2_X1 U12161 ( .A1(n12057), .A2(n12055), .ZN(n9702) );
  INV_X1 U12162 ( .A(n9698), .ZN(n9699) );
  OR2_X1 U12163 ( .A1(n9700), .A2(n9699), .ZN(n9701) );
  INV_X1 U12164 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n9707) );
  OR2_X1 U12165 ( .A1(n9705), .A2(n14785), .ZN(n9706) );
  OAI21_X1 U12166 ( .B1(n14787), .B2(n9707), .A(n9706), .ZN(P1_U3462) );
  XNOR2_X1 U12167 ( .A(n9866), .B(n10788), .ZN(n9721) );
  INV_X1 U12168 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n10140) );
  MUX2_X1 U12169 ( .A(P2_REG2_REG_2__SCAN_IN), .B(n10140), .S(n14807), .Z(
        n14806) );
  XNOR2_X1 U12170 ( .A(n9724), .B(P2_REG2_REG_1__SCAN_IN), .ZN(n13403) );
  AND2_X1 U12171 ( .A1(P2_REG2_REG_0__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), 
        .ZN(n13402) );
  NAND2_X1 U12172 ( .A1(n13403), .A2(n13402), .ZN(n13401) );
  NAND2_X1 U12173 ( .A1(n8037), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n9708) );
  NAND2_X1 U12174 ( .A1(n13401), .A2(n9708), .ZN(n14805) );
  NAND2_X1 U12175 ( .A1(n14806), .A2(n14805), .ZN(n14804) );
  NAND2_X1 U12176 ( .A1(n14807), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n9709) );
  NAND2_X1 U12177 ( .A1(n14804), .A2(n9709), .ZN(n13412) );
  INV_X1 U12178 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n9710) );
  XNOR2_X1 U12179 ( .A(n9728), .B(n9710), .ZN(n13413) );
  NAND2_X1 U12180 ( .A1(n13412), .A2(n13413), .ZN(n13411) );
  NAND2_X1 U12181 ( .A1(n9728), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n9711) );
  NAND2_X1 U12182 ( .A1(n13411), .A2(n9711), .ZN(n13424) );
  INV_X1 U12183 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n10297) );
  MUX2_X1 U12184 ( .A(n10297), .B(P2_REG2_REG_4__SCAN_IN), .S(n13421), .Z(
        n13425) );
  NAND2_X1 U12185 ( .A1(n13424), .A2(n13425), .ZN(n13423) );
  OR2_X1 U12186 ( .A1(n13421), .A2(n10297), .ZN(n9712) );
  NAND2_X1 U12187 ( .A1(n13423), .A2(n9712), .ZN(n14814) );
  INV_X1 U12188 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n10188) );
  XNOR2_X1 U12189 ( .A(n14819), .B(n10188), .ZN(n14815) );
  NAND2_X1 U12190 ( .A1(n14814), .A2(n14815), .ZN(n14813) );
  NAND2_X1 U12191 ( .A1(n14819), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n9713) );
  NAND2_X1 U12192 ( .A1(n14813), .A2(n9713), .ZN(n13436) );
  INV_X1 U12193 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n9714) );
  MUX2_X1 U12194 ( .A(P2_REG2_REG_6__SCAN_IN), .B(n9714), .S(n9733), .Z(n13437) );
  NAND2_X1 U12195 ( .A1(n13436), .A2(n13437), .ZN(n13435) );
  NAND2_X1 U12196 ( .A1(n9733), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n9715) );
  NAND2_X1 U12197 ( .A1(n13435), .A2(n9715), .ZN(n13453) );
  INV_X1 U12198 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n10322) );
  XNOR2_X1 U12199 ( .A(n13444), .B(n10322), .ZN(n13454) );
  NAND2_X1 U12200 ( .A1(n13453), .A2(n13454), .ZN(n13452) );
  NAND2_X1 U12201 ( .A1(n13444), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n9716) );
  NAND2_X1 U12202 ( .A1(n13452), .A2(n9716), .ZN(n14826) );
  INV_X1 U12203 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n9717) );
  MUX2_X1 U12204 ( .A(P2_REG2_REG_8__SCAN_IN), .B(n9717), .S(n9736), .Z(n14827) );
  NAND2_X1 U12205 ( .A1(n14826), .A2(n14827), .ZN(n14825) );
  NAND2_X1 U12206 ( .A1(n9736), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n9718) );
  NAND2_X1 U12207 ( .A1(n14825), .A2(n9718), .ZN(n14843) );
  XNOR2_X1 U12208 ( .A(n14846), .B(P2_REG2_REG_9__SCAN_IN), .ZN(n14842) );
  NOR2_X1 U12209 ( .A1(n14843), .A2(n14842), .ZN(n14845) );
  AOI21_X1 U12210 ( .B1(n10634), .B2(n9738), .A(n14845), .ZN(n14854) );
  INV_X1 U12211 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n9719) );
  MUX2_X1 U12212 ( .A(P2_REG2_REG_10__SCAN_IN), .B(n9719), .S(n14863), .Z(
        n14853) );
  AND2_X1 U12213 ( .A1(n14854), .A2(n14853), .ZN(n14855) );
  AOI21_X1 U12214 ( .B1(n14863), .B2(P2_REG2_REG_10__SCAN_IN), .A(n14855), 
        .ZN(n9720) );
  NAND2_X1 U12215 ( .A1(n9720), .A2(n9721), .ZN(n9861) );
  OAI21_X1 U12216 ( .B1(n9721), .B2(n9720), .A(n9861), .ZN(n9744) );
  NAND2_X1 U12217 ( .A1(n14890), .A2(n9866), .ZN(n9722) );
  NAND2_X1 U12218 ( .A1(P2_REG3_REG_11__SCAN_IN), .A2(P2_U3088), .ZN(n10841)
         );
  OAI211_X1 U12219 ( .C1(n9723), .C2(n14926), .A(n9722), .B(n10841), .ZN(n9743) );
  MUX2_X1 U12220 ( .A(P2_REG1_REG_2__SCAN_IN), .B(n8051), .S(n14807), .Z(
        n14803) );
  XNOR2_X1 U12221 ( .A(n9724), .B(P2_REG1_REG_1__SCAN_IN), .ZN(n13400) );
  AND2_X1 U12222 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), 
        .ZN(n13399) );
  NAND2_X1 U12223 ( .A1(n13400), .A2(n13399), .ZN(n13398) );
  NAND2_X1 U12224 ( .A1(n8037), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n9725) );
  NAND2_X1 U12225 ( .A1(n13398), .A2(n9725), .ZN(n14802) );
  NAND2_X1 U12226 ( .A1(n14803), .A2(n14802), .ZN(n14801) );
  NAND2_X1 U12227 ( .A1(n14807), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n9726) );
  NAND2_X1 U12228 ( .A1(n14801), .A2(n9726), .ZN(n13415) );
  INV_X1 U12229 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n9727) );
  XNOR2_X1 U12230 ( .A(n9728), .B(n9727), .ZN(n13416) );
  NAND2_X1 U12231 ( .A1(n13415), .A2(n13416), .ZN(n13414) );
  NAND2_X1 U12232 ( .A1(n9728), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n9729) );
  NAND2_X1 U12233 ( .A1(n13414), .A2(n9729), .ZN(n13427) );
  INV_X1 U12234 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n10260) );
  MUX2_X1 U12235 ( .A(n10260), .B(P2_REG1_REG_4__SCAN_IN), .S(n13421), .Z(
        n13428) );
  NAND2_X1 U12236 ( .A1(n13427), .A2(n13428), .ZN(n13426) );
  OR2_X1 U12237 ( .A1(n13421), .A2(n10260), .ZN(n9730) );
  NAND2_X1 U12238 ( .A1(n13426), .A2(n9730), .ZN(n14817) );
  INV_X1 U12239 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n9731) );
  XNOR2_X1 U12240 ( .A(n14819), .B(n9731), .ZN(n14818) );
  NAND2_X1 U12241 ( .A1(n14817), .A2(n14818), .ZN(n14816) );
  NAND2_X1 U12242 ( .A1(n14819), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n9732) );
  NAND2_X1 U12243 ( .A1(n14816), .A2(n9732), .ZN(n13439) );
  INV_X1 U12244 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n15007) );
  MUX2_X1 U12245 ( .A(P2_REG1_REG_6__SCAN_IN), .B(n15007), .S(n9733), .Z(
        n13440) );
  NAND2_X1 U12246 ( .A1(n13439), .A2(n13440), .ZN(n13438) );
  NAND2_X1 U12247 ( .A1(n9733), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n9734) );
  NAND2_X1 U12248 ( .A1(n13438), .A2(n9734), .ZN(n13450) );
  INV_X1 U12249 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n15009) );
  MUX2_X1 U12250 ( .A(P2_REG1_REG_7__SCAN_IN), .B(n15009), .S(n13444), .Z(
        n13451) );
  NAND2_X1 U12251 ( .A1(n13450), .A2(n13451), .ZN(n13449) );
  NAND2_X1 U12252 ( .A1(n13444), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n9735) );
  NAND2_X1 U12253 ( .A1(n13449), .A2(n9735), .ZN(n14829) );
  INV_X1 U12254 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n15011) );
  MUX2_X1 U12255 ( .A(P2_REG1_REG_8__SCAN_IN), .B(n15011), .S(n9736), .Z(
        n14830) );
  NAND2_X1 U12256 ( .A1(n14829), .A2(n14830), .ZN(n14828) );
  NAND2_X1 U12257 ( .A1(n9736), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n9737) );
  NAND2_X1 U12258 ( .A1(n14828), .A2(n9737), .ZN(n14839) );
  INV_X1 U12259 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n15013) );
  MUX2_X1 U12260 ( .A(n15013), .B(P2_REG1_REG_9__SCAN_IN), .S(n14846), .Z(
        n14838) );
  AOI21_X1 U12261 ( .B1(n15013), .B2(n9738), .A(n14841), .ZN(n14858) );
  INV_X1 U12262 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n15015) );
  MUX2_X1 U12263 ( .A(P2_REG1_REG_10__SCAN_IN), .B(n15015), .S(n14863), .Z(
        n14857) );
  AND2_X1 U12264 ( .A1(n14858), .A2(n14857), .ZN(n14859) );
  INV_X1 U12265 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n9739) );
  MUX2_X1 U12266 ( .A(n9739), .B(P2_REG1_REG_11__SCAN_IN), .S(n9866), .Z(n9740) );
  NOR2_X1 U12267 ( .A1(n9741), .A2(n9740), .ZN(n9865) );
  AOI211_X1 U12268 ( .C1(n9741), .C2(n9740), .A(n14884), .B(n9865), .ZN(n9742)
         );
  AOI211_X1 U12269 ( .C1(n14918), .C2(n9744), .A(n9743), .B(n9742), .ZN(n9745)
         );
  INV_X1 U12270 ( .A(n9745), .ZN(P2_U3225) );
  INV_X1 U12271 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n9760) );
  NAND2_X1 U12272 ( .A1(n6906), .A2(n14187), .ZN(n9747) );
  NAND2_X1 U12273 ( .A1(n11775), .A2(n14725), .ZN(n11779) );
  NAND2_X1 U12274 ( .A1(n9747), .A2(n9746), .ZN(n9749) );
  NAND2_X1 U12275 ( .A1(n9752), .A2(n6473), .ZN(n9748) );
  NAND2_X1 U12276 ( .A1(n9749), .A2(n9748), .ZN(n10403) );
  AND2_X1 U12277 ( .A1(n9750), .A2(n14728), .ZN(n9751) );
  OR2_X1 U12278 ( .A1(n9888), .A2(n9892), .ZN(n11791) );
  NAND2_X1 U12279 ( .A1(n9888), .A2(n9892), .ZN(n11790) );
  AND2_X1 U12280 ( .A1(n11791), .A2(n11790), .ZN(n11788) );
  NAND2_X1 U12281 ( .A1(n9752), .A2(n6906), .ZN(n9753) );
  NAND2_X1 U12282 ( .A1(n9754), .A2(n9753), .ZN(n10391) );
  NAND2_X1 U12283 ( .A1(n10391), .A2(n10404), .ZN(n10393) );
  NAND2_X1 U12284 ( .A1(n10393), .A2(n9755), .ZN(n9756) );
  INV_X1 U12285 ( .A(n11788), .ZN(n11999) );
  NAND2_X1 U12286 ( .A1(n10669), .A2(n10399), .ZN(n9890) );
  OAI211_X1 U12287 ( .C1(n10669), .C2(n10399), .A(n7114), .B(n9890), .ZN(
        n10673) );
  OAI211_X1 U12288 ( .C1(n10669), .C2(n14753), .A(n10673), .B(n10668), .ZN(
        n9757) );
  AOI21_X1 U12289 ( .B1(n10675), .B2(n14783), .A(n9757), .ZN(n9758) );
  OAI21_X1 U12290 ( .B1(n14780), .B2(n10677), .A(n9758), .ZN(n9761) );
  NAND2_X1 U12291 ( .A1(n9761), .A2(n14799), .ZN(n9759) );
  OAI21_X1 U12292 ( .B1(n14799), .B2(n9760), .A(n9759), .ZN(P1_U3531) );
  INV_X1 U12293 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n9763) );
  NAND2_X1 U12294 ( .A1(n9761), .A2(n14787), .ZN(n9762) );
  OAI21_X1 U12295 ( .B1(n14787), .B2(n9763), .A(n9762), .ZN(P1_U3468) );
  OAI222_X1 U12296 ( .A1(n12848), .A2(P3_U3151), .B1(n13250), .B2(n9765), .C1(
        n9764), .C2(n13247), .ZN(P3_U3278) );
  INV_X1 U12297 ( .A(n9766), .ZN(n9768) );
  NAND2_X1 U12298 ( .A1(n9768), .A2(P3_STATE_REG_SCAN_IN), .ZN(n12741) );
  NAND2_X1 U12299 ( .A1(n9767), .A2(n12741), .ZN(n9781) );
  OR2_X1 U12300 ( .A1(n12671), .A2(n9768), .ZN(n9769) );
  AND2_X1 U12301 ( .A1(n7450), .A2(n9769), .ZN(n9780) );
  AND2_X1 U12302 ( .A1(n9781), .A2(n9780), .ZN(n9784) );
  INV_X1 U12303 ( .A(n9784), .ZN(n9770) );
  MUX2_X1 U12304 ( .A(n9770), .B(n12765), .S(n12737), .Z(n15088) );
  MUX2_X1 U12305 ( .A(n10035), .B(n9995), .S(n12836), .Z(n9963) );
  AND2_X1 U12306 ( .A1(n9963), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n9957) );
  INV_X1 U12307 ( .A(P3_REG2_REG_1__SCAN_IN), .ZN(n9772) );
  INV_X1 U12308 ( .A(P3_REG1_REG_1__SCAN_IN), .ZN(n9771) );
  MUX2_X1 U12309 ( .A(n9772), .B(n9771), .S(n7916), .Z(n9773) );
  NAND2_X1 U12310 ( .A1(n9773), .A2(n7431), .ZN(n10122) );
  INV_X1 U12311 ( .A(n9773), .ZN(n9774) );
  NAND2_X1 U12312 ( .A1(n9774), .A2(n9795), .ZN(n9775) );
  NAND2_X1 U12313 ( .A1(n9776), .A2(n9957), .ZN(n10124) );
  OAI21_X1 U12314 ( .B1(n9957), .B2(n9776), .A(n10124), .ZN(n9793) );
  NAND2_X1 U12315 ( .A1(n9784), .A2(n12836), .ZN(n12853) );
  INV_X1 U12316 ( .A(P3_REG1_REG_0__SCAN_IN), .ZN(n9995) );
  NOR2_X1 U12317 ( .A1(n9995), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n9958) );
  INV_X1 U12318 ( .A(n9958), .ZN(n10077) );
  NOR2_X1 U12319 ( .A1(P3_IR_REG_1__SCAN_IN), .A2(n10077), .ZN(n9777) );
  AOI21_X1 U12320 ( .B1(n7431), .B2(n10077), .A(n9777), .ZN(n9778) );
  NAND2_X1 U12321 ( .A1(P3_REG1_REG_1__SCAN_IN), .A2(n9778), .ZN(n10076) );
  OAI21_X1 U12322 ( .B1(n9778), .B2(P3_REG1_REG_1__SCAN_IN), .A(n10076), .ZN(
        n9779) );
  NAND2_X1 U12323 ( .A1(n15097), .A2(n9779), .ZN(n9791) );
  INV_X1 U12324 ( .A(n9780), .ZN(n9782) );
  AOI22_X1 U12325 ( .A1(n15094), .A2(P3_ADDR_REG_1__SCAN_IN), .B1(
        P3_REG3_REG_1__SCAN_IN), .B2(P3_U3151), .ZN(n9790) );
  INV_X1 U12326 ( .A(P3_REG2_REG_0__SCAN_IN), .ZN(n10035) );
  NOR2_X1 U12327 ( .A1(P3_IR_REG_0__SCAN_IN), .A2(n10035), .ZN(n9962) );
  NAND2_X1 U12328 ( .A1(n10087), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n9785) );
  AOI21_X1 U12329 ( .B1(n9786), .B2(n9772), .A(n10086), .ZN(n9787) );
  INV_X1 U12330 ( .A(n9787), .ZN(n9788) );
  NAND2_X1 U12331 ( .A1(n14404), .A2(n9788), .ZN(n9789) );
  NAND3_X1 U12332 ( .A1(n9791), .A2(n9790), .A3(n9789), .ZN(n9792) );
  AOI21_X1 U12333 ( .B1(n15064), .B2(n9793), .A(n9792), .ZN(n9794) );
  OAI21_X1 U12334 ( .B1(n9795), .B2(n15088), .A(n9794), .ZN(P3_U3183) );
  XNOR2_X1 U12335 ( .A(n11394), .B(P2_B_REG_SCAN_IN), .ZN(n9796) );
  INV_X1 U12336 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n14930) );
  NAND2_X1 U12337 ( .A1(n14928), .A2(n14930), .ZN(n9799) );
  INV_X1 U12338 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n14935) );
  NAND2_X1 U12339 ( .A1(n14928), .A2(n14935), .ZN(n9802) );
  OR2_X1 U12340 ( .A1(n13818), .A2(n9800), .ZN(n9801) );
  NAND2_X1 U12341 ( .A1(n9802), .A2(n9801), .ZN(n9909) );
  INV_X1 U12342 ( .A(n9909), .ZN(n10136) );
  NOR4_X1 U12343 ( .A1(P2_D_REG_6__SCAN_IN), .A2(P2_D_REG_7__SCAN_IN), .A3(
        P2_D_REG_8__SCAN_IN), .A4(P2_D_REG_9__SCAN_IN), .ZN(n9811) );
  OR4_X1 U12344 ( .A1(P2_D_REG_2__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .A3(
        P2_D_REG_4__SCAN_IN), .A4(P2_D_REG_5__SCAN_IN), .ZN(n9808) );
  NOR4_X1 U12345 ( .A1(P2_D_REG_18__SCAN_IN), .A2(P2_D_REG_19__SCAN_IN), .A3(
        P2_D_REG_20__SCAN_IN), .A4(P2_D_REG_21__SCAN_IN), .ZN(n9806) );
  NOR4_X1 U12346 ( .A1(P2_D_REG_16__SCAN_IN), .A2(P2_D_REG_14__SCAN_IN), .A3(
        P2_D_REG_15__SCAN_IN), .A4(P2_D_REG_17__SCAN_IN), .ZN(n9805) );
  NOR4_X1 U12347 ( .A1(P2_D_REG_26__SCAN_IN), .A2(P2_D_REG_27__SCAN_IN), .A3(
        P2_D_REG_28__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n9804) );
  NOR4_X1 U12348 ( .A1(P2_D_REG_22__SCAN_IN), .A2(P2_D_REG_23__SCAN_IN), .A3(
        P2_D_REG_24__SCAN_IN), .A4(P2_D_REG_25__SCAN_IN), .ZN(n9803) );
  NAND4_X1 U12349 ( .A1(n9806), .A2(n9805), .A3(n9804), .A4(n9803), .ZN(n9807)
         );
  NOR4_X1 U12350 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        n9808), .A4(n9807), .ZN(n9810) );
  NOR4_X1 U12351 ( .A1(P2_D_REG_10__SCAN_IN), .A2(P2_D_REG_11__SCAN_IN), .A3(
        P2_D_REG_12__SCAN_IN), .A4(P2_D_REG_13__SCAN_IN), .ZN(n9809) );
  NAND3_X1 U12352 ( .A1(n9811), .A2(n9810), .A3(n9809), .ZN(n9812) );
  NAND2_X1 U12353 ( .A1(n14928), .A2(n9812), .ZN(n9911) );
  NAND3_X1 U12354 ( .A1(n9914), .A2(n10136), .A3(n9911), .ZN(n9826) );
  INV_X1 U12355 ( .A(n14932), .ZN(n14934) );
  OR2_X1 U12356 ( .A1(n9826), .A2(n14934), .ZN(n9819) );
  OR2_X1 U12357 ( .A1(n8022), .A2(n14938), .ZN(n9815) );
  INV_X1 U12358 ( .A(n9813), .ZN(n9814) );
  NAND2_X1 U12359 ( .A1(n9814), .A2(n11649), .ZN(n10141) );
  NOR2_X1 U12360 ( .A1(n14986), .A2(n9824), .ZN(n9816) );
  NOR2_X1 U12361 ( .A1(n14938), .A2(n9817), .ZN(n9818) );
  AND2_X4 U12362 ( .A1(n11649), .A2(n9818), .ZN(n14988) );
  INV_X1 U12363 ( .A(n12163), .ZN(n12083) );
  NOR2_X1 U12364 ( .A1(n10001), .A2(n12083), .ZN(n9835) );
  INV_X1 U12365 ( .A(n9835), .ZN(n9821) );
  AOI21_X1 U12366 ( .B1(n13359), .B2(n9821), .A(n9820), .ZN(n9831) );
  INV_X1 U12367 ( .A(n10216), .ZN(n14940) );
  NAND2_X1 U12368 ( .A1(n9823), .A2(n9822), .ZN(n13366) );
  NAND2_X1 U12369 ( .A1(n9824), .A2(n8822), .ZN(n13657) );
  INV_X1 U12370 ( .A(n9912), .ZN(n9825) );
  NAND2_X1 U12371 ( .A1(n9826), .A2(n9825), .ZN(n9828) );
  OR2_X1 U12372 ( .A1(n11649), .A2(n9827), .ZN(n9910) );
  NAND2_X1 U12373 ( .A1(n9828), .A2(n9910), .ZN(n10048) );
  OR2_X1 U12374 ( .A1(n10048), .A2(n14934), .ZN(n9936) );
  AOI22_X1 U12375 ( .A1(n11753), .A2(n13396), .B1(P2_REG3_REG_0__SCAN_IN), 
        .B2(n9936), .ZN(n9830) );
  INV_X1 U12376 ( .A(n13327), .ZN(n13347) );
  NAND3_X1 U12377 ( .A1(n13347), .A2(n8838), .A3(n10001), .ZN(n9829) );
  OAI211_X1 U12378 ( .C1(n9831), .C2(n14940), .A(n9830), .B(n9829), .ZN(
        P2_U3204) );
  NAND2_X2 U12379 ( .A1(n9833), .A2(n13680), .ZN(n13654) );
  NOR2_X1 U12380 ( .A1(n10036), .A2(n10216), .ZN(n9837) );
  XNOR2_X2 U12381 ( .A(n10036), .B(n9834), .ZN(n9937) );
  NAND2_X1 U12382 ( .A1(n13396), .A2(n12163), .ZN(n9932) );
  XNOR2_X1 U12383 ( .A(n9937), .B(n9932), .ZN(n9836) );
  AOI21_X1 U12384 ( .B1(n9837), .B2(n9836), .A(n9931), .ZN(n9844) );
  INV_X1 U12385 ( .A(n8838), .ZN(n10008) );
  INV_X1 U12386 ( .A(n13640), .ZN(n13655) );
  INV_X1 U12387 ( .A(n8841), .ZN(n10007) );
  OAI22_X1 U12388 ( .A1(n10008), .A2(n13353), .B1(n13351), .B2(n10007), .ZN(
        n9842) );
  INV_X1 U12389 ( .A(n9836), .ZN(n9838) );
  NOR3_X1 U12390 ( .A1(n13327), .A2(n10001), .A3(n9838), .ZN(n9841) );
  INV_X1 U12391 ( .A(n9936), .ZN(n9839) );
  INV_X1 U12392 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n10169) );
  OAI22_X1 U12393 ( .A1(n13371), .A2(n9834), .B1(n9839), .B2(n10169), .ZN(
        n9840) );
  NOR3_X1 U12394 ( .A1(n9842), .A2(n9841), .A3(n9840), .ZN(n9843) );
  OAI21_X1 U12395 ( .B1(n9844), .B2(n13334), .A(n9843), .ZN(P2_U3194) );
  INV_X1 U12396 ( .A(n14001), .ZN(n9846) );
  MUX2_X1 U12397 ( .A(n9846), .B(n9845), .S(n6484), .Z(n9847) );
  NOR2_X1 U12398 ( .A1(n9847), .A2(n9428), .ZN(n9848) );
  AOI211_X1 U12399 ( .C1(n9850), .C2(n9849), .A(n13979), .B(n9848), .ZN(n14009) );
  AOI211_X1 U12400 ( .C1(n9852), .C2(n9851), .A(n6516), .B(n14647), .ZN(n9860)
         );
  AOI211_X1 U12401 ( .C1(n9855), .C2(n9854), .A(n9853), .B(n14651), .ZN(n9859)
         );
  AND2_X1 U12402 ( .A1(P1_U3086), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n10339) );
  AOI21_X1 U12403 ( .B1(n14003), .B2(P1_ADDR_REG_4__SCAN_IN), .A(n10339), .ZN(
        n9856) );
  OAI21_X1 U12404 ( .B1(n9857), .B2(n14642), .A(n9856), .ZN(n9858) );
  OR4_X1 U12405 ( .A1(n14009), .A2(n9860), .A3(n9859), .A4(n9858), .ZN(
        P1_U3247) );
  MUX2_X1 U12406 ( .A(P2_REG2_REG_12__SCAN_IN), .B(n10866), .S(n10925), .Z(
        n9863) );
  OAI21_X1 U12407 ( .B1(P2_REG2_REG_11__SCAN_IN), .B2(n9866), .A(n9861), .ZN(
        n9862) );
  NAND2_X1 U12408 ( .A1(n9862), .A2(n9863), .ZN(n10913) );
  OAI21_X1 U12409 ( .B1(n9863), .B2(n9862), .A(n10913), .ZN(n9864) );
  INV_X1 U12410 ( .A(n9864), .ZN(n9875) );
  AOI21_X1 U12411 ( .B1(n9866), .B2(P2_REG1_REG_11__SCAN_IN), .A(n9865), .ZN(
        n9869) );
  MUX2_X1 U12412 ( .A(P2_REG1_REG_12__SCAN_IN), .B(n9867), .S(n10925), .Z(
        n9868) );
  NAND2_X1 U12413 ( .A1(n9869), .A2(n9868), .ZN(n10924) );
  OAI21_X1 U12414 ( .B1(n9869), .B2(n9868), .A(n10924), .ZN(n9873) );
  INV_X1 U12415 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n9871) );
  NAND2_X1 U12416 ( .A1(n14890), .A2(n10925), .ZN(n9870) );
  NAND2_X1 U12417 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(P2_U3088), .ZN(n11721)
         );
  OAI211_X1 U12418 ( .C1(n14926), .C2(n9871), .A(n9870), .B(n11721), .ZN(n9872) );
  AOI21_X1 U12419 ( .B1(n9873), .B2(n14913), .A(n9872), .ZN(n9874) );
  OAI21_X1 U12420 ( .B1(n9875), .B2(n14880), .A(n9874), .ZN(P2_U3226) );
  INV_X1 U12421 ( .A(n10986), .ZN(n9880) );
  INV_X1 U12422 ( .A(n14889), .ZN(n10914) );
  OAI222_X1 U12423 ( .A1(n13822), .A2(n9876), .B1(n13820), .B2(n9880), .C1(
        n10914), .C2(P2_U3088), .ZN(P2_U3313) );
  NAND2_X1 U12424 ( .A1(n9877), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9878) );
  INV_X1 U12425 ( .A(n14610), .ZN(n9879) );
  OAI222_X1 U12426 ( .A1(n14292), .A2(n9881), .B1(n12152), .B2(n9880), .C1(
        n9879), .C2(P1_U3086), .ZN(P1_U3341) );
  OAI222_X1 U12427 ( .A1(P3_U3151), .A2(n12840), .B1(n13247), .B2(n9883), .C1(
        n13250), .C2(n9882), .ZN(P3_U3277) );
  INV_X1 U12428 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n9905) );
  NAND2_X1 U12429 ( .A1(n9884), .A2(n11960), .ZN(n9887) );
  AOI22_X1 U12430 ( .A1(n11430), .A2(P2_DATAO_REG_4__SCAN_IN), .B1(n6478), 
        .B2(n9885), .ZN(n9886) );
  NAND2_X1 U12431 ( .A1(n9887), .A2(n9886), .ZN(n11798) );
  XNOR2_X1 U12432 ( .A(n13993), .B(n11798), .ZN(n11996) );
  INV_X1 U12433 ( .A(n9892), .ZN(n13994) );
  OR2_X1 U12434 ( .A1(n13994), .A2(n9888), .ZN(n9889) );
  XOR2_X1 U12435 ( .A(n11996), .B(n10425), .Z(n10615) );
  AOI21_X1 U12436 ( .B1(n9890), .B2(n11798), .A(n14493), .ZN(n9891) );
  NAND2_X1 U12437 ( .A1(n9891), .A2(n14710), .ZN(n10608) );
  INV_X1 U12438 ( .A(n14457), .ZN(n14169) );
  OR2_X1 U12439 ( .A1(n9892), .A2(n14169), .ZN(n9899) );
  NAND2_X1 U12440 ( .A1(n11587), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n9897) );
  NAND2_X1 U12441 ( .A1(n10452), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n9896) );
  BUF_X1 U12442 ( .A(n6475), .Z(n9893) );
  XNOR2_X1 U12443 ( .A(n10439), .B(P1_REG3_REG_5__SCAN_IN), .ZN(n14705) );
  NAND2_X1 U12444 ( .A1(n9893), .A2(n14705), .ZN(n9895) );
  NAND2_X1 U12445 ( .A1(n11526), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n9894) );
  NAND4_X1 U12446 ( .A1(n9897), .A2(n9896), .A3(n9895), .A4(n9894), .ZN(n13992) );
  NAND2_X1 U12447 ( .A1(n13992), .A2(n14455), .ZN(n9898) );
  NAND2_X1 U12448 ( .A1(n9899), .A2(n9898), .ZN(n10610) );
  INV_X1 U12449 ( .A(n10610), .ZN(n9900) );
  OAI211_X1 U12450 ( .C1(n10484), .C2(n14753), .A(n10608), .B(n9900), .ZN(
        n9903) );
  NAND2_X1 U12451 ( .A1(n9901), .A2(n11791), .ZN(n10486) );
  XNOR2_X1 U12452 ( .A(n10486), .B(n11996), .ZN(n9902) );
  NOR2_X1 U12453 ( .A1(n9902), .A2(n14780), .ZN(n10609) );
  AOI211_X1 U12454 ( .C1(n10615), .C2(n14783), .A(n9903), .B(n10609), .ZN(
        n9906) );
  OR2_X1 U12455 ( .A1(n9906), .A2(n14797), .ZN(n9904) );
  OAI21_X1 U12456 ( .B1(n14799), .B2(n9905), .A(n9904), .ZN(P1_U3532) );
  INV_X1 U12457 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n9908) );
  OR2_X1 U12458 ( .A1(n9906), .A2(n14785), .ZN(n9907) );
  OAI21_X1 U12459 ( .B1(n14787), .B2(n9908), .A(n9907), .ZN(P1_U3471) );
  AND2_X1 U12460 ( .A1(n9909), .A2(n14932), .ZN(n14933) );
  NAND2_X1 U12461 ( .A1(n9911), .A2(n9910), .ZN(n10135) );
  NOR2_X1 U12462 ( .A1(n10135), .A2(n9912), .ZN(n9913) );
  INV_X1 U12463 ( .A(n9948), .ZN(n9945) );
  OR2_X1 U12464 ( .A1(n13396), .A2(n10012), .ZN(n9916) );
  NAND2_X1 U12465 ( .A1(n9945), .A2(n9946), .ZN(n9944) );
  OR2_X1 U12466 ( .A1(n8841), .A2(n9953), .ZN(n9917) );
  NAND2_X1 U12467 ( .A1(n9944), .A2(n9917), .ZN(n9919) );
  INV_X1 U12468 ( .A(n10179), .ZN(n9918) );
  NAND2_X1 U12469 ( .A1(n9919), .A2(n9918), .ZN(n10193) );
  OAI21_X1 U12470 ( .B1(n9919), .B2(n9918), .A(n10193), .ZN(n10240) );
  INV_X1 U12471 ( .A(n10240), .ZN(n9929) );
  NOR2_X1 U12472 ( .A1(n8838), .A2(n14940), .ZN(n10006) );
  NAND2_X1 U12473 ( .A1(n9921), .A2(n10006), .ZN(n10005) );
  NAND2_X1 U12474 ( .A1(n10005), .A2(n9922), .ZN(n9949) );
  NAND2_X1 U12475 ( .A1(n9949), .A2(n9948), .ZN(n9947) );
  OR2_X1 U12476 ( .A1(n8841), .A2(n10143), .ZN(n9923) );
  NAND2_X1 U12477 ( .A1(n9947), .A2(n9923), .ZN(n10180) );
  XNOR2_X1 U12478 ( .A(n10180), .B(n10179), .ZN(n9926) );
  AND2_X1 U12479 ( .A1(n14938), .A2(n9817), .ZN(n9924) );
  OAI22_X1 U12480 ( .A1(n10007), .A2(n13655), .B1(n11710), .B2(n13657), .ZN(
        n13271) );
  AOI21_X1 U12481 ( .B1(n9926), .B2(n13677), .A(n13271), .ZN(n10242) );
  NAND2_X1 U12482 ( .A1(n9951), .A2(n10238), .ZN(n10253) );
  OR2_X1 U12483 ( .A1(n9951), .A2(n10238), .ZN(n9927) );
  AND2_X1 U12484 ( .A1(n10253), .A2(n9927), .ZN(n10235) );
  AOI22_X1 U12485 ( .A1(n10235), .A2(n14988), .B1(n13270), .B2(n14986), .ZN(
        n9928) );
  OAI211_X1 U12486 ( .C1(n9929), .C2(n14984), .A(n10242), .B(n9928), .ZN(n9988) );
  NAND2_X1 U12487 ( .A1(n9988), .A2(n15019), .ZN(n9930) );
  OAI21_X1 U12488 ( .B1(n15019), .B2(n9727), .A(n9930), .ZN(P2_U3502) );
  NAND2_X1 U12489 ( .A1(n9937), .A2(n9932), .ZN(n9933) );
  XNOR2_X1 U12490 ( .A(n12098), .B(n9953), .ZN(n10038) );
  NAND2_X1 U12491 ( .A1(n8841), .A2(n12163), .ZN(n10037) );
  XNOR2_X1 U12492 ( .A(n10038), .B(n10037), .ZN(n9939) );
  INV_X1 U12493 ( .A(n10039), .ZN(n9943) );
  NOR2_X1 U12494 ( .A1(n13371), .A2(n10143), .ZN(n9935) );
  INV_X1 U12495 ( .A(n13395), .ZN(n10191) );
  OAI22_X1 U12496 ( .A1(n7122), .A2(n13353), .B1(n13351), .B2(n10191), .ZN(
        n9934) );
  AOI211_X1 U12497 ( .C1(P2_REG3_REG_2__SCAN_IN), .C2(n9936), .A(n9935), .B(
        n9934), .ZN(n9942) );
  OAI22_X1 U12498 ( .A1(n13327), .A2(n7122), .B1(n9937), .B2(n13334), .ZN(
        n9940) );
  NAND3_X1 U12499 ( .A1(n9940), .A2(n9939), .A3(n9938), .ZN(n9941) );
  OAI211_X1 U12500 ( .C1(n13334), .C2(n9943), .A(n9942), .B(n9941), .ZN(
        P2_U3209) );
  OAI21_X1 U12501 ( .B1(n9946), .B2(n9945), .A(n9944), .ZN(n10148) );
  INV_X1 U12502 ( .A(n10148), .ZN(n9955) );
  OAI21_X1 U12503 ( .B1(n9949), .B2(n9948), .A(n9947), .ZN(n9950) );
  AOI222_X1 U12504 ( .A1(n13677), .A2(n9950), .B1(n13395), .B2(n13642), .C1(
        n13396), .C2(n13640), .ZN(n10151) );
  INV_X1 U12505 ( .A(n10013), .ZN(n9952) );
  AOI21_X1 U12506 ( .B1(n9953), .B2(n9952), .A(n9951), .ZN(n10146) );
  AOI22_X1 U12507 ( .A1(n10146), .A2(n14988), .B1(n9953), .B2(n14986), .ZN(
        n9954) );
  OAI211_X1 U12508 ( .C1(n14984), .C2(n9955), .A(n10151), .B(n9954), .ZN(n9985) );
  NAND2_X1 U12509 ( .A1(n9985), .A2(n15019), .ZN(n9956) );
  OAI21_X1 U12510 ( .B1(n15019), .B2(n8051), .A(n9956), .ZN(P2_U3501) );
  NOR3_X1 U12511 ( .A1(n15097), .A2(n14404), .A3(n15064), .ZN(n9968) );
  INV_X1 U12512 ( .A(n9957), .ZN(n9967) );
  AND2_X1 U12513 ( .A1(n15097), .A2(n9958), .ZN(n9961) );
  INV_X1 U12514 ( .A(n15094), .ZN(n15077) );
  OAI22_X1 U12515 ( .A1(n15077), .A2(n9959), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n10107), .ZN(n9960) );
  AOI211_X1 U12516 ( .C1(n9962), .C2(n14404), .A(n9961), .B(n9960), .ZN(n9966)
         );
  OR2_X1 U12517 ( .A1(n15090), .A2(n9963), .ZN(n9964) );
  MUX2_X1 U12518 ( .A(n9964), .B(n15088), .S(P3_IR_REG_0__SCAN_IN), .Z(n9965)
         );
  OAI211_X1 U12519 ( .C1(n9968), .C2(n9967), .A(n9966), .B(n9965), .ZN(
        P3_U3182) );
  INV_X1 U12520 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n9970) );
  MUX2_X1 U12521 ( .A(P1_REG1_REG_8__SCAN_IN), .B(n9970), .S(n10462), .Z(n9971) );
  OAI21_X1 U12522 ( .B1(n9972), .B2(n9971), .A(n10219), .ZN(n9982) );
  NAND2_X1 U12523 ( .A1(n14658), .A2(n10462), .ZN(n9974) );
  NAND2_X1 U12524 ( .A1(P1_REG3_REG_8__SCAN_IN), .A2(P1_U3086), .ZN(n9973) );
  OAI211_X1 U12525 ( .C1(n9975), .C2(n14661), .A(n9974), .B(n9973), .ZN(n9981)
         );
  AOI21_X1 U12526 ( .B1(n10449), .B2(P1_REG2_REG_7__SCAN_IN), .A(n9976), .ZN(
        n9979) );
  INV_X1 U12527 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n9977) );
  MUX2_X1 U12528 ( .A(n9977), .B(P1_REG2_REG_8__SCAN_IN), .S(n10462), .Z(n9978) );
  AOI211_X1 U12529 ( .C1(n9979), .C2(n9978), .A(n14651), .B(n10225), .ZN(n9980) );
  AOI211_X1 U12530 ( .C1(n14633), .C2(n9982), .A(n9981), .B(n9980), .ZN(n9983)
         );
  INV_X1 U12531 ( .A(n9983), .ZN(P1_U3251) );
  INV_X1 U12532 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n9987) );
  NAND2_X1 U12533 ( .A1(n9985), .A2(n14953), .ZN(n9986) );
  OAI21_X1 U12534 ( .B1(n14953), .B2(n9987), .A(n9986), .ZN(P2_U3436) );
  INV_X1 U12535 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n9990) );
  NAND2_X1 U12536 ( .A1(n9988), .A2(n15004), .ZN(n9989) );
  OAI21_X1 U12537 ( .B1(n14953), .B2(n9990), .A(n9989), .ZN(P2_U3439) );
  OAI222_X1 U12538 ( .A1(P3_U3151), .A2(n12857), .B1(n13247), .B2(n9992), .C1(
        n13250), .C2(n9991), .ZN(P3_U3276) );
  AND2_X1 U12539 ( .A1(n12766), .A2(n10104), .ZN(n12546) );
  OR2_X1 U12540 ( .A1(n12546), .A2(n12553), .ZN(n12699) );
  NAND3_X1 U12541 ( .A1(n12699), .A2(n15170), .A3(n9993), .ZN(n9994) );
  OAI21_X1 U12542 ( .B1(n15110), .B2(n15111), .A(n9994), .ZN(n10029) );
  OAI22_X1 U12543 ( .A1(n13179), .A2(n10104), .B1(n15193), .B2(n9995), .ZN(
        n9996) );
  AOI21_X1 U12544 ( .B1(n10029), .B2(n15193), .A(n9996), .ZN(n9997) );
  INV_X1 U12545 ( .A(n9997), .ZN(P3_U3459) );
  INV_X1 U12546 ( .A(P3_REG0_REG_0__SCAN_IN), .ZN(n9998) );
  OAI22_X1 U12547 ( .A1(n13234), .A2(n10104), .B1(n15177), .B2(n9998), .ZN(
        n9999) );
  AOI21_X1 U12548 ( .B1(n10029), .B2(n15177), .A(n9999), .ZN(n10000) );
  INV_X1 U12549 ( .A(n10000), .ZN(P3_U3390) );
  INV_X1 U12550 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n10018) );
  INV_X1 U12551 ( .A(n10001), .ZN(n10004) );
  INV_X1 U12552 ( .A(n10002), .ZN(n10003) );
  AOI21_X1 U12553 ( .B1(n9921), .B2(n10004), .A(n10003), .ZN(n10175) );
  OAI21_X1 U12554 ( .B1(n9921), .B2(n10006), .A(n10005), .ZN(n10011) );
  OAI22_X1 U12555 ( .A1(n10008), .A2(n13655), .B1(n10007), .B2(n13657), .ZN(
        n10010) );
  NOR2_X1 U12556 ( .A1(n10175), .A2(n13654), .ZN(n10009) );
  AOI211_X1 U12557 ( .C1(n13645), .C2(n10011), .A(n10010), .B(n10009), .ZN(
        n10170) );
  AND2_X1 U12558 ( .A1(n10012), .A2(n10216), .ZN(n10014) );
  OR2_X1 U12559 ( .A1(n10014), .A2(n10013), .ZN(n10172) );
  OAI22_X1 U12560 ( .A1(n10172), .A2(n14996), .B1(n9834), .B2(n14994), .ZN(
        n10015) );
  INV_X1 U12561 ( .A(n10015), .ZN(n10016) );
  OAI211_X1 U12562 ( .C1(n10175), .C2(n14937), .A(n10170), .B(n10016), .ZN(
        n10019) );
  NAND2_X1 U12563 ( .A1(n10019), .A2(n15019), .ZN(n10017) );
  OAI21_X1 U12564 ( .B1(n15019), .B2(n10018), .A(n10017), .ZN(P2_U3500) );
  INV_X1 U12565 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n10021) );
  NAND2_X1 U12566 ( .A1(n10019), .A2(n15004), .ZN(n10020) );
  OAI21_X1 U12567 ( .B1(n14953), .B2(n10021), .A(n10020), .ZN(P2_U3433) );
  MUX2_X1 U12568 ( .A(n10024), .B(n10023), .S(n10022), .Z(n10025) );
  NAND2_X1 U12569 ( .A1(n10026), .A2(n10025), .ZN(n10030) );
  NAND2_X1 U12570 ( .A1(n10029), .A2(n13106), .ZN(n10034) );
  INV_X1 U12571 ( .A(n10030), .ZN(n10031) );
  NOR2_X1 U12572 ( .A1(n15170), .A2(n12695), .ZN(n15105) );
  INV_X1 U12573 ( .A(n13094), .ZN(n13108) );
  AOI22_X1 U12574 ( .A1(n13108), .A2(n10032), .B1(n13092), .B2(
        P3_REG3_REG_0__SCAN_IN), .ZN(n10033) );
  OAI211_X1 U12575 ( .C1(n10035), .C2(n13106), .A(n10034), .B(n10033), .ZN(
        P3_U3233) );
  NAND2_X1 U12576 ( .A1(n8833), .A2(n12159), .ZN(n10347) );
  XNOR2_X1 U12577 ( .A(n13270), .B(n12098), .ZN(n10045) );
  NAND2_X1 U12578 ( .A1(n13395), .A2(n12163), .ZN(n10040) );
  NOR2_X1 U12579 ( .A1(n10045), .A2(n10040), .ZN(n10041) );
  AOI21_X1 U12580 ( .B1(n10045), .B2(n10040), .A(n10041), .ZN(n13268) );
  INV_X1 U12581 ( .A(n10041), .ZN(n10042) );
  OAI21_X1 U12582 ( .B1(n10044), .B2(n13267), .A(n11716), .ZN(n10054) );
  NOR4_X1 U12583 ( .A1(n13327), .A2(n10191), .A3(n10045), .A4(n10044), .ZN(
        n10053) );
  INV_X1 U12584 ( .A(n10046), .ZN(n10047) );
  INV_X1 U12585 ( .A(n13366), .ZN(n13308) );
  OAI22_X1 U12586 ( .A1(n10377), .A2(n13657), .B1(n10191), .B2(n13655), .ZN(
        n10251) );
  AOI22_X1 U12587 ( .A1(n13308), .A2(n10251), .B1(P2_REG3_REG_4__SCAN_IN), 
        .B2(P2_U3088), .ZN(n10051) );
  NAND2_X1 U12588 ( .A1(n9820), .A2(n10299), .ZN(n10050) );
  OAI211_X1 U12589 ( .C1(n13352), .C2(n10296), .A(n10051), .B(n10050), .ZN(
        n10052) );
  AOI211_X1 U12590 ( .C1(n10054), .C2(n13359), .A(n10053), .B(n10052), .ZN(
        n10055) );
  INV_X1 U12591 ( .A(n10055), .ZN(P2_U3202) );
  MUX2_X1 U12592 ( .A(P3_REG2_REG_6__SCAN_IN), .B(P3_REG1_REG_6__SCAN_IN), .S(
        n12836), .Z(n10156) );
  XNOR2_X1 U12593 ( .A(n10156), .B(n10155), .ZN(n10157) );
  NAND2_X1 U12594 ( .A1(n10124), .A2(n10122), .ZN(n10060) );
  INV_X1 U12595 ( .A(P3_REG2_REG_2__SCAN_IN), .ZN(n10056) );
  INV_X1 U12596 ( .A(P3_REG1_REG_2__SCAN_IN), .ZN(n10075) );
  MUX2_X1 U12597 ( .A(n10056), .B(n10075), .S(n12836), .Z(n10057) );
  NAND2_X1 U12598 ( .A1(n10057), .A2(n10111), .ZN(n15029) );
  INV_X1 U12599 ( .A(n10057), .ZN(n10058) );
  NAND2_X1 U12600 ( .A1(n10058), .A2(n10088), .ZN(n10059) );
  AND2_X1 U12601 ( .A1(n15029), .A2(n10059), .ZN(n10121) );
  NAND2_X1 U12602 ( .A1(n10060), .A2(n10121), .ZN(n15030) );
  NAND2_X1 U12603 ( .A1(n15030), .A2(n15029), .ZN(n10066) );
  INV_X1 U12604 ( .A(P3_REG2_REG_3__SCAN_IN), .ZN(n10062) );
  INV_X1 U12605 ( .A(P3_REG1_REG_3__SCAN_IN), .ZN(n10061) );
  MUX2_X1 U12606 ( .A(n10062), .B(n10061), .S(n12836), .Z(n10063) );
  NAND2_X1 U12607 ( .A1(n10063), .A2(n15035), .ZN(n10067) );
  INV_X1 U12608 ( .A(n10063), .ZN(n10064) );
  INV_X1 U12609 ( .A(n15035), .ZN(n14312) );
  NAND2_X1 U12610 ( .A1(n10064), .A2(n14312), .ZN(n10065) );
  AND2_X1 U12611 ( .A1(n10067), .A2(n10065), .ZN(n15027) );
  NAND2_X1 U12612 ( .A1(n10066), .A2(n15027), .ZN(n15032) );
  NAND2_X1 U12613 ( .A1(n15032), .A2(n10067), .ZN(n15040) );
  MUX2_X1 U12614 ( .A(P3_REG2_REG_4__SCAN_IN), .B(P3_REG1_REG_4__SCAN_IN), .S(
        n12836), .Z(n10068) );
  XNOR2_X1 U12615 ( .A(n10068), .B(n10091), .ZN(n15039) );
  NAND2_X1 U12616 ( .A1(n15040), .A2(n15039), .ZN(n15038) );
  INV_X1 U12617 ( .A(n10068), .ZN(n10069) );
  NAND2_X1 U12618 ( .A1(n10069), .A2(n10091), .ZN(n10070) );
  NAND2_X1 U12619 ( .A1(n15038), .A2(n10070), .ZN(n15063) );
  INV_X1 U12620 ( .A(P3_REG2_REG_5__SCAN_IN), .ZN(n10072) );
  INV_X1 U12621 ( .A(P3_REG1_REG_5__SCAN_IN), .ZN(n10071) );
  MUX2_X1 U12622 ( .A(n10072), .B(n10071), .S(n12836), .Z(n10074) );
  INV_X1 U12623 ( .A(n10074), .ZN(n10073) );
  NAND2_X1 U12624 ( .A1(n10073), .A2(n10093), .ZN(n15059) );
  AND2_X1 U12625 ( .A1(n10074), .A2(n15069), .ZN(n15060) );
  AOI21_X1 U12626 ( .B1(n15063), .B2(n15059), .A(n15060), .ZN(n10158) );
  XOR2_X1 U12627 ( .A(n10157), .B(n10158), .Z(n10103) );
  INV_X1 U12628 ( .A(P3_REG1_REG_6__SCAN_IN), .ZN(n15184) );
  AOI22_X1 U12629 ( .A1(n10160), .A2(n15184), .B1(P3_REG1_REG_6__SCAN_IN), 
        .B2(n10155), .ZN(n10083) );
  INV_X1 U12630 ( .A(P3_REG1_REG_4__SCAN_IN), .ZN(n15181) );
  AOI22_X1 U12631 ( .A1(P3_REG1_REG_4__SCAN_IN), .A2(n15051), .B1(n10091), 
        .B2(n15181), .ZN(n15043) );
  MUX2_X1 U12632 ( .A(n10075), .B(P3_REG1_REG_2__SCAN_IN), .S(n10111), .Z(
        n10114) );
  OAI21_X1 U12633 ( .B1(P3_IR_REG_1__SCAN_IN), .B2(n10077), .A(n10076), .ZN(
        n10113) );
  NAND2_X1 U12634 ( .A1(n10114), .A2(n10113), .ZN(n10112) );
  OAI21_X1 U12635 ( .B1(n10111), .B2(n10075), .A(n10112), .ZN(n10078) );
  NAND2_X1 U12636 ( .A1(n14312), .A2(n10078), .ZN(n10079) );
  XNOR2_X1 U12637 ( .A(n15035), .B(n10078), .ZN(n15023) );
  NAND2_X1 U12638 ( .A1(P3_REG1_REG_3__SCAN_IN), .A2(n15023), .ZN(n15022) );
  NAND2_X1 U12639 ( .A1(n10093), .A2(n10080), .ZN(n10081) );
  NAND2_X1 U12640 ( .A1(P3_REG1_REG_5__SCAN_IN), .A2(n15067), .ZN(n15066) );
  OAI21_X1 U12641 ( .B1(n10083), .B2(n10082), .A(n10159), .ZN(n10101) );
  NOR2_X1 U12642 ( .A1(n10084), .A2(P3_STATE_REG_SCAN_IN), .ZN(n10814) );
  AOI21_X1 U12643 ( .B1(n15094), .B2(P3_ADDR_REG_6__SCAN_IN), .A(n10814), .ZN(
        n10085) );
  OAI21_X1 U12644 ( .B1(n15088), .B2(n10155), .A(n10085), .ZN(n10100) );
  AOI21_X1 U12645 ( .B1(P3_REG2_REG_0__SCAN_IN), .B2(n10087), .A(n10086), .ZN(
        n10110) );
  AOI22_X1 U12646 ( .A1(n10111), .A2(P3_REG2_REG_2__SCAN_IN), .B1(n10056), 
        .B2(n10088), .ZN(n10109) );
  NOR2_X1 U12647 ( .A1(n10110), .A2(n10109), .ZN(n10108) );
  NOR2_X1 U12648 ( .A1(n15035), .A2(n10089), .ZN(n10090) );
  XNOR2_X1 U12649 ( .A(n10089), .B(n15035), .ZN(n15021) );
  INV_X1 U12650 ( .A(P3_REG2_REG_4__SCAN_IN), .ZN(n10524) );
  AOI22_X1 U12651 ( .A1(P3_REG2_REG_4__SCAN_IN), .A2(n10091), .B1(n15051), 
        .B2(n10524), .ZN(n15045) );
  NOR2_X1 U12652 ( .A1(n15069), .A2(n10092), .ZN(n10094) );
  INV_X1 U12653 ( .A(P3_REG2_REG_6__SCAN_IN), .ZN(n10095) );
  AOI22_X1 U12654 ( .A1(n10160), .A2(P3_REG2_REG_6__SCAN_IN), .B1(n10095), 
        .B2(n10155), .ZN(n10096) );
  AOI21_X1 U12655 ( .B1(n10097), .B2(n10096), .A(n10152), .ZN(n10098) );
  NOR2_X1 U12656 ( .A1(n10098), .A2(n15101), .ZN(n10099) );
  AOI211_X1 U12657 ( .C1(n15097), .C2(n10101), .A(n10100), .B(n10099), .ZN(
        n10102) );
  OAI21_X1 U12658 ( .B1(n10103), .B2(n15090), .A(n10102), .ZN(P3_U3188) );
  INV_X1 U12659 ( .A(n12497), .ZN(n12452) );
  NAND2_X1 U12660 ( .A1(n12452), .A2(P3_STATE_REG_SCAN_IN), .ZN(n10293) );
  INV_X1 U12661 ( .A(n10293), .ZN(n10208) );
  INV_X1 U12662 ( .A(n12471), .ZN(n12443) );
  OAI22_X1 U12663 ( .A1(n12443), .A2(n15110), .B1(n10104), .B2(n12500), .ZN(
        n10105) );
  AOI21_X1 U12664 ( .B1(n12502), .B2(n12699), .A(n10105), .ZN(n10106) );
  OAI21_X1 U12665 ( .B1(n10208), .B2(n10107), .A(n10106), .ZN(P3_U3172) );
  AOI21_X1 U12666 ( .B1(n10110), .B2(n10109), .A(n10108), .ZN(n10120) );
  INV_X1 U12667 ( .A(n15088), .ZN(n15070) );
  NAND2_X1 U12668 ( .A1(n15070), .A2(n10111), .ZN(n10119) );
  OAI21_X1 U12669 ( .B1(n10114), .B2(n10113), .A(n10112), .ZN(n10115) );
  NAND2_X1 U12670 ( .A1(n15097), .A2(n10115), .ZN(n10117) );
  AOI22_X1 U12671 ( .A1(n15094), .A2(P3_ADDR_REG_2__SCAN_IN), .B1(
        P3_REG3_REG_2__SCAN_IN), .B2(P3_U3151), .ZN(n10116) );
  AND2_X1 U12672 ( .A1(n10117), .A2(n10116), .ZN(n10118) );
  OAI211_X1 U12673 ( .C1(n10120), .C2(n15101), .A(n10119), .B(n10118), .ZN(
        n10127) );
  INV_X1 U12674 ( .A(n10121), .ZN(n10123) );
  NAND3_X1 U12675 ( .A1(n10124), .A2(n10123), .A3(n10122), .ZN(n10125) );
  AOI21_X1 U12676 ( .B1(n15030), .B2(n10125), .A(n15090), .ZN(n10126) );
  OR2_X1 U12677 ( .A1(n10127), .A2(n10126), .ZN(P3_U3184) );
  INV_X1 U12678 ( .A(n11163), .ZN(n10133) );
  NOR2_X1 U12679 ( .A1(n6668), .A2(n10128), .ZN(n10129) );
  MUX2_X1 U12680 ( .A(n10128), .B(n10129), .S(P1_IR_REG_15__SCAN_IN), .Z(
        n10131) );
  INV_X1 U12681 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n10130) );
  AND2_X1 U12682 ( .A1(n6668), .A2(n10130), .ZN(n10308) );
  OAI222_X1 U12683 ( .A1(n14292), .A2(n10132), .B1(n12152), .B2(n10133), .C1(
        n14036), .C2(P1_U3086), .ZN(P1_U3340) );
  OAI222_X1 U12684 ( .A1(n13822), .A2(n10134), .B1(n13820), .B2(n10133), .C1(
        n14904), .C2(P2_U3088), .ZN(P2_U3312) );
  INV_X1 U12685 ( .A(n10135), .ZN(n10137) );
  NAND4_X1 U12686 ( .A1(n10137), .A2(n10136), .A3(n14932), .A4(n14931), .ZN(
        n10138) );
  INV_X1 U12687 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n10139) );
  OAI22_X1 U12688 ( .A1(n13606), .A2(n10140), .B1(n10139), .B2(n13607), .ZN(
        n10145) );
  INV_X1 U12689 ( .A(n10141), .ZN(n10142) );
  NOR2_X1 U12690 ( .A1(n13688), .A2(n10143), .ZN(n10144) );
  AOI211_X1 U12691 ( .C1(n10146), .C2(n13669), .A(n10145), .B(n10144), .ZN(
        n10150) );
  NAND2_X1 U12692 ( .A1(n9832), .A2(n13490), .ZN(n10173) );
  NAND2_X1 U12693 ( .A1(n13654), .A2(n10173), .ZN(n10147) );
  INV_X1 U12694 ( .A(n13649), .ZN(n13690) );
  NAND2_X1 U12695 ( .A1(n13690), .A2(n10148), .ZN(n10149) );
  OAI211_X1 U12696 ( .C1(n13671), .C2(n10151), .A(n10150), .B(n10149), .ZN(
        P2_U3263) );
  INV_X1 U12697 ( .A(n10269), .ZN(n10273) );
  INV_X1 U12698 ( .A(P3_REG2_REG_7__SCAN_IN), .ZN(n10153) );
  NOR2_X1 U12699 ( .A1(n10153), .A2(n10154), .ZN(n10262) );
  AOI21_X1 U12700 ( .B1(n10154), .B2(n10153), .A(n10262), .ZN(n10168) );
  MUX2_X1 U12701 ( .A(P3_REG2_REG_7__SCAN_IN), .B(P3_REG1_REG_7__SCAN_IN), .S(
        n12836), .Z(n10267) );
  XNOR2_X1 U12702 ( .A(n10267), .B(n10269), .ZN(n10270) );
  XNOR2_X1 U12703 ( .A(n10271), .B(n10270), .ZN(n10166) );
  NAND2_X1 U12704 ( .A1(P3_REG1_REG_7__SCAN_IN), .A2(n10161), .ZN(n10274) );
  OAI21_X1 U12705 ( .B1(P3_REG1_REG_7__SCAN_IN), .B2(n10161), .A(n10274), .ZN(
        n10162) );
  NAND2_X1 U12706 ( .A1(n10162), .A2(n15097), .ZN(n10164) );
  AOI22_X1 U12707 ( .A1(n15094), .A2(P3_ADDR_REG_7__SCAN_IN), .B1(
        P3_REG3_REG_7__SCAN_IN), .B2(P3_U3151), .ZN(n10163) );
  OAI211_X1 U12708 ( .C1(n15088), .C2(n10273), .A(n10164), .B(n10163), .ZN(
        n10165) );
  AOI21_X1 U12709 ( .B1(n10166), .B2(n15064), .A(n10165), .ZN(n10167) );
  OAI21_X1 U12710 ( .B1(n10168), .B2(n15101), .A(n10167), .ZN(P3_U3189) );
  OAI22_X1 U12711 ( .A1(n10170), .A2(n13671), .B1(n10169), .B2(n13607), .ZN(
        n10178) );
  INV_X1 U12712 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n10171) );
  OAI22_X1 U12713 ( .A1(n11660), .A2(n10172), .B1(n13606), .B2(n10171), .ZN(
        n10177) );
  INV_X1 U12714 ( .A(n10173), .ZN(n10174) );
  NAND2_X1 U12715 ( .A1(n13606), .A2(n10174), .ZN(n13666) );
  OAI22_X1 U12716 ( .A1(n10175), .A2(n13666), .B1(n13688), .B2(n9834), .ZN(
        n10176) );
  OR3_X1 U12717 ( .A1(n10178), .A2(n10177), .A3(n10176), .ZN(P2_U3264) );
  INV_X1 U12718 ( .A(n10196), .ZN(n10184) );
  NAND2_X1 U12719 ( .A1(n10180), .A2(n10179), .ZN(n10182) );
  NAND2_X1 U12720 ( .A1(n10191), .A2(n13270), .ZN(n10181) );
  NAND2_X1 U12721 ( .A1(n10182), .A2(n10181), .ZN(n10248) );
  NAND2_X1 U12722 ( .A1(n10248), .A2(n10249), .ZN(n10247) );
  OAI21_X1 U12723 ( .B1(n10184), .B2(n10183), .A(n10374), .ZN(n10185) );
  NAND2_X1 U12724 ( .A1(n10185), .A2(n13677), .ZN(n10187) );
  AOI22_X1 U12725 ( .A1(n13642), .A2(n13393), .B1(n8833), .B2(n13640), .ZN(
        n10186) );
  AND2_X1 U12726 ( .A1(n10187), .A2(n10186), .ZN(n14950) );
  XNOR2_X1 U12727 ( .A(n10323), .B(n10317), .ZN(n14948) );
  OAI22_X1 U12728 ( .A1(n13606), .A2(n10188), .B1(n11712), .B2(n13607), .ZN(
        n10190) );
  NOR2_X1 U12729 ( .A1(n13688), .A2(n10317), .ZN(n10189) );
  AOI211_X1 U12730 ( .C1(n14948), .C2(n13669), .A(n10190), .B(n10189), .ZN(
        n10198) );
  NAND2_X1 U12731 ( .A1(n10191), .A2(n10238), .ZN(n10192) );
  NAND2_X1 U12732 ( .A1(n10193), .A2(n10192), .ZN(n10244) );
  INV_X1 U12733 ( .A(n10249), .ZN(n10243) );
  NAND2_X1 U12734 ( .A1(n10244), .A2(n10243), .ZN(n10246) );
  NAND2_X1 U12735 ( .A1(n11710), .A2(n10194), .ZN(n10195) );
  NAND2_X1 U12736 ( .A1(n10246), .A2(n10195), .ZN(n10316) );
  XNOR2_X1 U12737 ( .A(n10316), .B(n10196), .ZN(n14945) );
  NAND2_X1 U12738 ( .A1(n14945), .A2(n13690), .ZN(n10197) );
  OAI211_X1 U12739 ( .C1(n14950), .C2(n13671), .A(n10198), .B(n10197), .ZN(
        P2_U3260) );
  INV_X1 U12740 ( .A(n12553), .ZN(n10200) );
  NAND3_X1 U12741 ( .A1(n10200), .A2(n12703), .A3(n11671), .ZN(n10201) );
  OAI211_X1 U12742 ( .C1(n10202), .C2(n10412), .A(n10199), .B(n10201), .ZN(
        n10203) );
  NAND2_X1 U12743 ( .A1(n10203), .A2(n12502), .ZN(n10207) );
  OAI22_X1 U12744 ( .A1(n12443), .A2(n10204), .B1(n15125), .B2(n12500), .ZN(
        n10205) );
  AOI21_X1 U12745 ( .B1(n12441), .B2(n12766), .A(n10205), .ZN(n10206) );
  OAI211_X1 U12746 ( .C1(n10208), .C2(n10417), .A(n10207), .B(n10206), .ZN(
        P3_U3162) );
  INV_X1 U12747 ( .A(n11180), .ZN(n10211) );
  OR2_X1 U12748 ( .A1(n10308), .A2(n10128), .ZN(n10209) );
  XNOR2_X1 U12749 ( .A(n10209), .B(P1_IR_REG_16__SCAN_IN), .ZN(n14625) );
  INV_X1 U12750 ( .A(n14625), .ZN(n14025) );
  OAI222_X1 U12751 ( .A1(n14292), .A2(n10210), .B1(n12152), .B2(n10211), .C1(
        n14025), .C2(P1_U3086), .ZN(P1_U3339) );
  INV_X1 U12752 ( .A(n13467), .ZN(n10932) );
  OAI222_X1 U12753 ( .A1(n13822), .A2(n10212), .B1(n13820), .B2(n10211), .C1(
        n10932), .C2(P2_U3088), .ZN(P2_U3311) );
  INV_X1 U12754 ( .A(n13607), .ZN(n13685) );
  INV_X1 U12755 ( .A(n13654), .ZN(n13570) );
  NOR2_X1 U12756 ( .A1(n13570), .A2(n13677), .ZN(n10213) );
  OAI22_X1 U12757 ( .A1(n14936), .A2(n10213), .B1(n7122), .B2(n13657), .ZN(
        n14941) );
  AOI21_X1 U12758 ( .B1(P2_REG3_REG_0__SCAN_IN), .B2(n13685), .A(n14941), .ZN(
        n10214) );
  NOR2_X1 U12759 ( .A1(n13671), .A2(n10214), .ZN(n10215) );
  AOI21_X1 U12760 ( .B1(n13671), .B2(P2_REG2_REG_0__SCAN_IN), .A(n10215), .ZN(
        n10218) );
  OAI21_X1 U12761 ( .B1(n13553), .B2(n13669), .A(n10216), .ZN(n10217) );
  OAI211_X1 U12762 ( .C1(n13666), .C2(n14936), .A(n10218), .B(n10217), .ZN(
        P2_U3265) );
  MUX2_X1 U12763 ( .A(P1_REG1_REG_9__SCAN_IN), .B(n14795), .S(n10563), .Z(
        n10221) );
  OAI21_X1 U12764 ( .B1(P1_REG1_REG_8__SCAN_IN), .B2(n10462), .A(n10219), .ZN(
        n10220) );
  NAND2_X1 U12765 ( .A1(n10220), .A2(n10221), .ZN(n10534) );
  OAI21_X1 U12766 ( .B1(n10221), .B2(n10220), .A(n10534), .ZN(n10232) );
  NAND2_X1 U12767 ( .A1(n14658), .A2(n10563), .ZN(n10223) );
  NAND2_X1 U12768 ( .A1(P1_REG3_REG_9__SCAN_IN), .A2(P1_U3086), .ZN(n10222) );
  OAI211_X1 U12769 ( .C1(n10224), .C2(n14661), .A(n10223), .B(n10222), .ZN(
        n10231) );
  INV_X1 U12770 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n10226) );
  MUX2_X1 U12771 ( .A(P1_REG2_REG_9__SCAN_IN), .B(n10226), .S(n10563), .Z(
        n10227) );
  INV_X1 U12772 ( .A(n10227), .ZN(n10228) );
  AOI211_X1 U12773 ( .C1(n10229), .C2(n10228), .A(n14651), .B(n10528), .ZN(
        n10230) );
  AOI211_X1 U12774 ( .C1(n14633), .C2(n10232), .A(n10231), .B(n10230), .ZN(
        n10233) );
  INV_X1 U12775 ( .A(n10233), .ZN(P1_U3252) );
  INV_X1 U12776 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n10234) );
  AOI22_X1 U12777 ( .A1(n13671), .A2(P2_REG2_REG_3__SCAN_IN), .B1(n13685), 
        .B2(n10234), .ZN(n10237) );
  NAND2_X1 U12778 ( .A1(n13669), .A2(n10235), .ZN(n10236) );
  OAI211_X1 U12779 ( .C1(n10238), .C2(n13688), .A(n10237), .B(n10236), .ZN(
        n10239) );
  AOI21_X1 U12780 ( .B1(n13690), .B2(n10240), .A(n10239), .ZN(n10241) );
  OAI21_X1 U12781 ( .B1(n13671), .B2(n10242), .A(n10241), .ZN(P2_U3262) );
  INV_X1 U12782 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n10257) );
  OR2_X1 U12783 ( .A1(n10244), .A2(n10243), .ZN(n10245) );
  AND2_X1 U12784 ( .A1(n10246), .A2(n10245), .ZN(n10303) );
  OAI21_X1 U12785 ( .B1(n10249), .B2(n10248), .A(n10247), .ZN(n10252) );
  NOR2_X1 U12786 ( .A1(n10303), .A2(n13654), .ZN(n10250) );
  AOI211_X1 U12787 ( .C1(n13645), .C2(n10252), .A(n10251), .B(n10250), .ZN(
        n10306) );
  NAND2_X1 U12788 ( .A1(n10253), .A2(n10299), .ZN(n10254) );
  AND2_X1 U12789 ( .A1(n10323), .A2(n10254), .ZN(n10300) );
  AOI22_X1 U12790 ( .A1(n10300), .A2(n14988), .B1(n10299), .B2(n14986), .ZN(
        n10255) );
  OAI211_X1 U12791 ( .C1(n10303), .C2(n14937), .A(n10306), .B(n10255), .ZN(
        n10258) );
  NAND2_X1 U12792 ( .A1(n10258), .A2(n14953), .ZN(n10256) );
  OAI21_X1 U12793 ( .B1(n15004), .B2(n10257), .A(n10256), .ZN(P2_U3442) );
  NAND2_X1 U12794 ( .A1(n10258), .A2(n15019), .ZN(n10259) );
  OAI21_X1 U12795 ( .B1(n15019), .B2(n10260), .A(n10259), .ZN(P2_U3503) );
  NOR2_X1 U12796 ( .A1(n10269), .A2(n10261), .ZN(n10263) );
  INV_X1 U12797 ( .A(P3_REG2_REG_8__SCAN_IN), .ZN(n10264) );
  AOI22_X1 U12798 ( .A1(P3_REG2_REG_8__SCAN_IN), .A2(n10699), .B1(n10709), 
        .B2(n10264), .ZN(n10265) );
  AOI21_X1 U12799 ( .B1(n10266), .B2(n10265), .A(n10693), .ZN(n10285) );
  INV_X1 U12800 ( .A(n10267), .ZN(n10268) );
  AOI22_X1 U12801 ( .A1(n10271), .A2(n10270), .B1(n10269), .B2(n10268), .ZN(
        n10712) );
  MUX2_X1 U12802 ( .A(P3_REG2_REG_8__SCAN_IN), .B(P3_REG1_REG_8__SCAN_IN), .S(
        n12836), .Z(n10710) );
  XNOR2_X1 U12803 ( .A(n10710), .B(n10709), .ZN(n10711) );
  XNOR2_X1 U12804 ( .A(n10712), .B(n10711), .ZN(n10283) );
  INV_X1 U12805 ( .A(P3_REG1_REG_8__SCAN_IN), .ZN(n15188) );
  AOI22_X1 U12806 ( .A1(P3_REG1_REG_8__SCAN_IN), .A2(n10709), .B1(n10699), 
        .B2(n15188), .ZN(n10277) );
  NAND2_X1 U12807 ( .A1(n10273), .A2(n10272), .ZN(n10275) );
  OAI21_X1 U12808 ( .B1(n10277), .B2(n10276), .A(n10698), .ZN(n10278) );
  NAND2_X1 U12809 ( .A1(n10278), .A2(n15097), .ZN(n10281) );
  NOR2_X1 U12810 ( .A1(n10279), .A2(P3_STATE_REG_SCAN_IN), .ZN(n11044) );
  AOI21_X1 U12811 ( .B1(n15094), .B2(P3_ADDR_REG_8__SCAN_IN), .A(n11044), .ZN(
        n10280) );
  OAI211_X1 U12812 ( .C1(n15088), .C2(n10709), .A(n10281), .B(n10280), .ZN(
        n10282) );
  AOI21_X1 U12813 ( .B1(n10283), .B2(n15064), .A(n10282), .ZN(n10284) );
  OAI21_X1 U12814 ( .B1(n10285), .B2(n15101), .A(n10284), .ZN(P3_U3190) );
  OAI222_X1 U12815 ( .A1(P3_U3151), .A2(n10288), .B1(n13247), .B2(n10287), 
        .C1(n13250), .C2(n10286), .ZN(P3_U3275) );
  XOR2_X1 U12816 ( .A(n10290), .B(n10289), .Z(n10295) );
  AOI22_X1 U12817 ( .A1(n12471), .A2(n12763), .B1(n12476), .B2(n15130), .ZN(
        n10291) );
  OAI21_X1 U12818 ( .B1(n15110), .B2(n12474), .A(n10291), .ZN(n10292) );
  AOI21_X1 U12819 ( .B1(P3_REG3_REG_2__SCAN_IN), .B2(n10293), .A(n10292), .ZN(
        n10294) );
  OAI21_X1 U12820 ( .B1(n10295), .B2(n12478), .A(n10294), .ZN(P3_U3177) );
  OAI22_X1 U12821 ( .A1(n13606), .A2(n10297), .B1(n10296), .B2(n13607), .ZN(
        n10298) );
  AOI21_X1 U12822 ( .B1(n13553), .B2(n10299), .A(n10298), .ZN(n10302) );
  NAND2_X1 U12823 ( .A1(n13669), .A2(n10300), .ZN(n10301) );
  OAI211_X1 U12824 ( .C1(n10303), .C2(n13666), .A(n10302), .B(n10301), .ZN(
        n10304) );
  INV_X1 U12825 ( .A(n10304), .ZN(n10305) );
  OAI21_X1 U12826 ( .B1(n10306), .B2(n13671), .A(n10305), .ZN(P2_U3261) );
  INV_X1 U12827 ( .A(n11240), .ZN(n10313) );
  INV_X1 U12828 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n10307) );
  NAND2_X1 U12829 ( .A1(n10308), .A2(n10307), .ZN(n10310) );
  NAND2_X1 U12830 ( .A1(n10310), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10309) );
  MUX2_X1 U12831 ( .A(P1_IR_REG_31__SCAN_IN), .B(n10309), .S(
        P1_IR_REG_17__SCAN_IN), .Z(n10311) );
  AND2_X1 U12832 ( .A1(n10311), .A2(n10679), .ZN(n14042) );
  INV_X1 U12833 ( .A(n14042), .ZN(n14641) );
  OAI222_X1 U12834 ( .A1(n14292), .A2(n10312), .B1(n12152), .B2(n10313), .C1(
        n14641), .C2(P1_U3086), .ZN(P1_U3338) );
  INV_X1 U12835 ( .A(n13468), .ZN(n14921) );
  OAI222_X1 U12836 ( .A1(n13822), .A2(n10314), .B1(n13820), .B2(n10313), .C1(
        n14921), .C2(P2_U3088), .ZN(P2_U3310) );
  NAND2_X1 U12837 ( .A1(n13394), .A2(n14947), .ZN(n10315) );
  NAND2_X1 U12838 ( .A1(n10316), .A2(n10315), .ZN(n10319) );
  NAND2_X1 U12839 ( .A1(n10377), .A2(n10317), .ZN(n10318) );
  NAND2_X1 U12840 ( .A1(n10319), .A2(n10318), .ZN(n10370) );
  NAND2_X1 U12841 ( .A1(n10380), .A2(n13393), .ZN(n10320) );
  OAI21_X1 U12842 ( .B1(n10321), .B2(n10328), .A(n10619), .ZN(n14961) );
  OAI22_X1 U12843 ( .A1(n13606), .A2(n10322), .B1(n10600), .B2(n13607), .ZN(
        n10326) );
  INV_X1 U12844 ( .A(n10624), .ZN(n14962) );
  INV_X1 U12845 ( .A(n11505), .ZN(n10324) );
  OAI21_X1 U12846 ( .B1(n14962), .B2(n10382), .A(n10324), .ZN(n14963) );
  NOR2_X1 U12847 ( .A1(n14963), .A2(n11660), .ZN(n10325) );
  AOI211_X1 U12848 ( .C1(n13553), .C2(n10624), .A(n10326), .B(n10325), .ZN(
        n10334) );
  INV_X1 U12849 ( .A(n13393), .ZN(n11709) );
  NAND2_X1 U12850 ( .A1(n10380), .A2(n11709), .ZN(n10327) );
  NAND2_X1 U12851 ( .A1(n10376), .A2(n10327), .ZN(n10623) );
  INV_X1 U12852 ( .A(n10328), .ZN(n10329) );
  XNOR2_X1 U12853 ( .A(n10623), .B(n10329), .ZN(n10330) );
  NAND2_X1 U12854 ( .A1(n10330), .A2(n13677), .ZN(n10332) );
  AOI22_X1 U12855 ( .A1(n13640), .A2(n13393), .B1(n13391), .B2(n13642), .ZN(
        n10331) );
  NAND2_X1 U12856 ( .A1(n10332), .A2(n10331), .ZN(n14964) );
  NAND2_X1 U12857 ( .A1(n14964), .A2(n13606), .ZN(n10333) );
  OAI211_X1 U12858 ( .C1(n14961), .C2(n13649), .A(n10334), .B(n10333), .ZN(
        P2_U3258) );
  AOI22_X1 U12859 ( .A1(n12303), .A2(n11798), .B1(n10746), .B2(n13993), .ZN(
        n10335) );
  XOR2_X1 U12860 ( .A(n11452), .B(n10335), .Z(n10647) );
  INV_X1 U12861 ( .A(n13993), .ZN(n10424) );
  OAI22_X1 U12862 ( .A1(n12276), .A2(n10424), .B1(n10484), .B2(n12223), .ZN(
        n10645) );
  XOR2_X1 U12863 ( .A(n10647), .B(n10648), .Z(n10344) );
  INV_X1 U12864 ( .A(n10612), .ZN(n10342) );
  AOI21_X1 U12865 ( .B1(n14466), .B2(n10610), .A(n10339), .ZN(n10341) );
  NAND2_X1 U12866 ( .A1(n14463), .A2(n11798), .ZN(n10340) );
  OAI211_X1 U12867 ( .C1(n14469), .C2(n10342), .A(n10341), .B(n10340), .ZN(
        n10343) );
  AOI21_X1 U12868 ( .B1(n10344), .B2(n14465), .A(n10343), .ZN(n10345) );
  INV_X1 U12869 ( .A(n10345), .ZN(P1_U3230) );
  XNOR2_X1 U12870 ( .A(n10380), .B(n6485), .ZN(n10594) );
  AND2_X1 U12871 ( .A1(n13393), .A2(n12163), .ZN(n10346) );
  NAND2_X1 U12872 ( .A1(n10594), .A2(n10346), .ZN(n10542) );
  OAI21_X1 U12873 ( .B1(n10594), .B2(n10346), .A(n10542), .ZN(n10355) );
  NAND2_X1 U12874 ( .A1(n13394), .A2(n12159), .ZN(n10350) );
  INV_X1 U12875 ( .A(n10350), .ZN(n10353) );
  XNOR2_X1 U12876 ( .A(n14947), .B(n6485), .ZN(n10352) );
  INV_X1 U12877 ( .A(n10347), .ZN(n10348) );
  OR2_X1 U12878 ( .A1(n10348), .A2(n11706), .ZN(n10349) );
  NAND2_X1 U12879 ( .A1(n11716), .A2(n10349), .ZN(n10351) );
  XNOR2_X1 U12880 ( .A(n10352), .B(n10350), .ZN(n11707) );
  AOI211_X1 U12881 ( .C1(n10355), .C2(n10354), .A(n13334), .B(n10596), .ZN(
        n10359) );
  OAI22_X1 U12882 ( .A1(n10377), .A2(n13353), .B1(n13351), .B2(n11766), .ZN(
        n10358) );
  NAND2_X1 U12883 ( .A1(n9820), .A2(n10380), .ZN(n10356) );
  NAND2_X1 U12884 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_U3088), .ZN(n13432) );
  OAI211_X1 U12885 ( .C1(n13352), .C2(n10385), .A(n10356), .B(n13432), .ZN(
        n10357) );
  OR3_X1 U12886 ( .A1(n10359), .A2(n10358), .A3(n10357), .ZN(P2_U3211) );
  OAI211_X1 U12887 ( .C1(n10362), .C2(n10361), .A(n10360), .B(n12502), .ZN(
        n10367) );
  MUX2_X1 U12888 ( .A(n12497), .B(P3_U3151), .S(P3_REG3_REG_3__SCAN_IN), .Z(
        n10365) );
  OAI22_X1 U12889 ( .A1(n12443), .A2(n10363), .B1(n12500), .B2(n15135), .ZN(
        n10364) );
  AOI211_X1 U12890 ( .C1(n12441), .C2(n6469), .A(n10365), .B(n10364), .ZN(
        n10366) );
  NAND2_X1 U12891 ( .A1(n10367), .A2(n10366), .ZN(P3_U3158) );
  INV_X1 U12892 ( .A(n10368), .ZN(n10369) );
  AOI21_X1 U12893 ( .B1(n10371), .B2(n10370), .A(n10369), .ZN(n14959) );
  INV_X1 U12894 ( .A(n14959), .ZN(n10390) );
  INV_X1 U12895 ( .A(n10371), .ZN(n10373) );
  NAND3_X1 U12896 ( .A1(n10374), .A2(n10373), .A3(n10372), .ZN(n10375) );
  AOI21_X1 U12897 ( .B1(n10376), .B2(n10375), .A(n13594), .ZN(n10379) );
  OAI22_X1 U12898 ( .A1(n10377), .A2(n13655), .B1(n11766), .B2(n13657), .ZN(
        n10378) );
  AOI211_X1 U12899 ( .C1(n14959), .C2(n13570), .A(n10379), .B(n10378), .ZN(
        n14956) );
  MUX2_X1 U12900 ( .A(n9714), .B(n14956), .S(n13606), .Z(n10389) );
  INV_X1 U12901 ( .A(n10380), .ZN(n14954) );
  INV_X1 U12902 ( .A(n10381), .ZN(n10384) );
  INV_X1 U12903 ( .A(n10382), .ZN(n10383) );
  OAI21_X1 U12904 ( .B1(n14954), .B2(n10384), .A(n10383), .ZN(n14955) );
  INV_X1 U12905 ( .A(n14955), .ZN(n10387) );
  OAI22_X1 U12906 ( .A1(n13688), .A2(n14954), .B1(n10385), .B2(n13607), .ZN(
        n10386) );
  AOI21_X1 U12907 ( .B1(n13669), .B2(n10387), .A(n10386), .ZN(n10388) );
  OAI211_X1 U12908 ( .C1(n10390), .C2(n13666), .A(n10389), .B(n10388), .ZN(
        P2_U3259) );
  OR2_X1 U12909 ( .A1(n10391), .A2(n10404), .ZN(n10392) );
  NAND2_X1 U12910 ( .A1(n10393), .A2(n10392), .ZN(n10405) );
  INV_X1 U12911 ( .A(n10405), .ZN(n14731) );
  NAND2_X1 U12912 ( .A1(n10395), .A2(n10394), .ZN(n11622) );
  OR2_X1 U12913 ( .A1(n11781), .A2(n14149), .ZN(n11976) );
  OR2_X1 U12914 ( .A1(n14706), .A2(n11976), .ZN(n14175) );
  NAND2_X1 U12915 ( .A1(n14728), .A2(n10396), .ZN(n10397) );
  NAND2_X1 U12916 ( .A1(n10397), .A2(n7114), .ZN(n10398) );
  NOR2_X1 U12917 ( .A1(n10399), .A2(n10398), .ZN(n14727) );
  INV_X1 U12918 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n14010) );
  OAI22_X1 U12919 ( .A1(n14708), .A2(n10401), .B1(n14010), .B2(n14188), .ZN(
        n10402) );
  AOI21_X1 U12920 ( .B1(n14713), .B2(n14727), .A(n10402), .ZN(n10411) );
  XNOR2_X1 U12921 ( .A(n10404), .B(n10403), .ZN(n10408) );
  NAND2_X1 U12922 ( .A1(n10405), .A2(n14743), .ZN(n10407) );
  AOI22_X1 U12923 ( .A1(n13994), .A2(n14455), .B1(n14457), .B2(n14187), .ZN(
        n10406) );
  OAI211_X1 U12924 ( .C1(n14780), .C2(n10408), .A(n10407), .B(n10406), .ZN(
        n14733) );
  INV_X1 U12925 ( .A(n14733), .ZN(n10409) );
  MUX2_X1 U12926 ( .A(n10409), .B(n9576), .S(n14706), .Z(n10410) );
  OAI211_X1 U12927 ( .C1(n14731), .C2(n14175), .A(n10411), .B(n10410), .ZN(
        P1_U3291) );
  XNOR2_X1 U12928 ( .A(n12703), .B(n12553), .ZN(n15126) );
  INV_X1 U12929 ( .A(n15120), .ZN(n12920) );
  AOI22_X1 U12930 ( .A1(n13098), .A2(n12766), .B1(n6469), .B2(n13100), .ZN(
        n10415) );
  OAI21_X1 U12931 ( .B1(n12703), .B2(n10412), .A(n15114), .ZN(n10413) );
  NAND2_X1 U12932 ( .A1(n10413), .A2(n13103), .ZN(n10414) );
  OAI211_X1 U12933 ( .C1(n15126), .C2(n12920), .A(n10415), .B(n10414), .ZN(
        n15128) );
  AOI21_X1 U12934 ( .B1(n15105), .B2(n10416), .A(n15128), .ZN(n10421) );
  INV_X1 U12935 ( .A(n15126), .ZN(n10419) );
  AND2_X1 U12936 ( .A1(n12695), .A2(n12547), .ZN(n15123) );
  OAI22_X1 U12937 ( .A1(n13106), .A2(n9772), .B1(n10417), .B2(n15108), .ZN(
        n10418) );
  AOI21_X1 U12938 ( .B1(n10419), .B2(n12926), .A(n10418), .ZN(n10420) );
  OAI21_X1 U12939 ( .B1(n10421), .B2(n13116), .A(n10420), .ZN(P3_U3232) );
  OAI222_X1 U12940 ( .A1(P3_U3151), .A2(n12552), .B1(n13247), .B2(n10423), 
        .C1(n13250), .C2(n10422), .ZN(P3_U3274) );
  OAI21_X1 U12941 ( .B1(n10425), .B2(n10424), .A(n10484), .ZN(n10427) );
  NAND2_X1 U12942 ( .A1(n10425), .A2(n10424), .ZN(n10426) );
  NAND2_X1 U12943 ( .A1(n10428), .A2(n11960), .ZN(n10431) );
  AOI22_X1 U12944 ( .A1(n11430), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n6479), 
        .B2(n10429), .ZN(n10430) );
  NAND2_X1 U12945 ( .A1(n10431), .A2(n10430), .ZN(n11807) );
  XNOR2_X1 U12946 ( .A(n11807), .B(n10650), .ZN(n14700) );
  OR2_X1 U12947 ( .A1(n13992), .A2(n11807), .ZN(n10432) );
  NAND2_X1 U12948 ( .A1(n10433), .A2(n11960), .ZN(n10436) );
  AOI22_X1 U12949 ( .A1(n11430), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n6479), 
        .B2(n10434), .ZN(n10435) );
  NAND2_X1 U12950 ( .A1(n10436), .A2(n10435), .ZN(n13945) );
  NAND2_X1 U12951 ( .A1(n11587), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n10445) );
  NAND2_X1 U12952 ( .A1(n10452), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n10444) );
  INV_X1 U12953 ( .A(n10439), .ZN(n10437) );
  AOI21_X1 U12954 ( .B1(n10437), .B2(P1_REG3_REG_5__SCAN_IN), .A(
        P1_REG3_REG_6__SCAN_IN), .ZN(n10440) );
  NAND2_X1 U12955 ( .A1(P1_REG3_REG_6__SCAN_IN), .A2(P1_REG3_REG_5__SCAN_IN), 
        .ZN(n10438) );
  NOR2_X1 U12956 ( .A1(n10439), .A2(n10438), .ZN(n10453) );
  OR2_X1 U12957 ( .A1(n10440), .A2(n10453), .ZN(n13944) );
  INV_X1 U12958 ( .A(n13944), .ZN(n10441) );
  NAND2_X1 U12959 ( .A1(n6475), .A2(n10441), .ZN(n10443) );
  NAND2_X1 U12960 ( .A1(n11526), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n10442) );
  NAND4_X1 U12961 ( .A1(n10445), .A2(n10444), .A3(n10443), .A4(n10442), .ZN(
        n13991) );
  XNOR2_X1 U12962 ( .A(n13945), .B(n13991), .ZN(n12001) );
  OR2_X1 U12963 ( .A1(n13945), .A2(n13991), .ZN(n10446) );
  NAND2_X1 U12964 ( .A1(n10448), .A2(n11960), .ZN(n10451) );
  AOI22_X1 U12965 ( .A1(n11430), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n6478), 
        .B2(n10449), .ZN(n10450) );
  NAND2_X1 U12966 ( .A1(n10451), .A2(n10450), .ZN(n11817) );
  NAND2_X1 U12967 ( .A1(n11587), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n10458) );
  INV_X2 U12968 ( .A(n10999), .ZN(n11616) );
  NAND2_X1 U12969 ( .A1(n11616), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n10457) );
  NAND2_X1 U12970 ( .A1(n10453), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n10465) );
  OR2_X1 U12971 ( .A1(n10453), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n10454) );
  AND2_X1 U12972 ( .A1(n10465), .A2(n10454), .ZN(n14690) );
  NAND2_X1 U12973 ( .A1(n9893), .A2(n14690), .ZN(n10456) );
  NAND2_X1 U12974 ( .A1(n11526), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n10455) );
  NAND4_X1 U12975 ( .A1(n10458), .A2(n10457), .A3(n10456), .A4(n10455), .ZN(
        n13990) );
  XNOR2_X1 U12976 ( .A(n11817), .B(n13990), .ZN(n12002) );
  INV_X1 U12977 ( .A(n12002), .ZN(n14687) );
  OR2_X1 U12978 ( .A1(n11817), .A2(n13990), .ZN(n10459) );
  NAND2_X1 U12979 ( .A1(n10461), .A2(n11960), .ZN(n10464) );
  AOI22_X1 U12980 ( .A1(n11430), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n6479), 
        .B2(n10462), .ZN(n10463) );
  NAND2_X1 U12981 ( .A1(n10464), .A2(n10463), .ZN(n11826) );
  NAND2_X1 U12982 ( .A1(n11587), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n10470) );
  NAND2_X1 U12983 ( .A1(n11616), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n10469) );
  NAND2_X1 U12984 ( .A1(n10465), .A2(n10827), .ZN(n10466) );
  AND2_X1 U12985 ( .A1(n10476), .A2(n10466), .ZN(n10831) );
  NAND2_X1 U12986 ( .A1(n9893), .A2(n10831), .ZN(n10468) );
  NAND2_X1 U12987 ( .A1(n11954), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n10467) );
  NAND4_X1 U12988 ( .A1(n10470), .A2(n10469), .A3(n10468), .A4(n10467), .ZN(
        n13989) );
  XNOR2_X1 U12989 ( .A(n11826), .B(n13989), .ZN(n12004) );
  INV_X1 U12990 ( .A(n12004), .ZN(n10578) );
  XNOR2_X1 U12991 ( .A(n10579), .B(n10578), .ZN(n14765) );
  INV_X1 U12992 ( .A(n14765), .ZN(n10502) );
  INV_X1 U12993 ( .A(n10831), .ZN(n10472) );
  OAI22_X1 U12994 ( .A1(n14179), .A2(n9977), .B1(n10472), .B2(n14188), .ZN(
        n10473) );
  AOI21_X1 U12995 ( .B1(n14476), .B2(n11826), .A(n10473), .ZN(n10501) );
  INV_X1 U12996 ( .A(n11817), .ZN(n14754) );
  AOI21_X1 U12997 ( .B1(n14693), .B2(n11826), .A(n14493), .ZN(n10483) );
  OR2_X1 U12998 ( .A1(n14693), .A2(n11826), .ZN(n14673) );
  NAND2_X1 U12999 ( .A1(n11587), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n10481) );
  NAND2_X1 U13000 ( .A1(n11616), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n10480) );
  NAND2_X1 U13001 ( .A1(n10476), .A2(n10475), .ZN(n10477) );
  NAND2_X1 U13002 ( .A1(n10572), .A2(n10477), .ZN(n11117) );
  INV_X1 U13003 ( .A(n11117), .ZN(n14668) );
  NAND2_X1 U13004 ( .A1(n9893), .A2(n14668), .ZN(n10479) );
  NAND2_X1 U13005 ( .A1(n11526), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n10478) );
  NAND4_X1 U13006 ( .A1(n10481), .A2(n10480), .A3(n10479), .A4(n10478), .ZN(
        n13988) );
  AOI22_X1 U13007 ( .A1(n14457), .A2(n13990), .B1(n13988), .B2(n14455), .ZN(
        n10828) );
  INV_X1 U13008 ( .A(n10828), .ZN(n10482) );
  AOI21_X1 U13009 ( .B1(n10483), .B2(n14673), .A(n10482), .ZN(n14762) );
  INV_X1 U13010 ( .A(n11798), .ZN(n10484) );
  NAND2_X1 U13011 ( .A1(n10486), .A2(n10485), .ZN(n10488) );
  NAND2_X1 U13012 ( .A1(n10484), .A2(n13993), .ZN(n10487) );
  NAND2_X1 U13013 ( .A1(n10488), .A2(n10487), .ZN(n14699) );
  NAND2_X1 U13014 ( .A1(n11807), .A2(n10650), .ZN(n10489) );
  NAND2_X1 U13015 ( .A1(n14699), .A2(n10489), .ZN(n10491) );
  OR2_X1 U13016 ( .A1(n10650), .A2(n11807), .ZN(n10490) );
  NAND2_X1 U13017 ( .A1(n10491), .A2(n10490), .ZN(n10510) );
  INV_X1 U13018 ( .A(n13991), .ZN(n10493) );
  NOR2_X1 U13019 ( .A1(n13945), .A2(n10493), .ZN(n10492) );
  OR2_X1 U13020 ( .A1(n10510), .A2(n10492), .ZN(n10495) );
  NAND2_X1 U13021 ( .A1(n13945), .A2(n10493), .ZN(n10494) );
  NAND2_X1 U13022 ( .A1(n10495), .A2(n10494), .ZN(n14686) );
  INV_X1 U13023 ( .A(n13990), .ZN(n10496) );
  OR2_X1 U13024 ( .A1(n11817), .A2(n10496), .ZN(n10497) );
  OAI211_X1 U13025 ( .C1(n10498), .C2(n12004), .A(n14701), .B(n10561), .ZN(
        n14763) );
  OAI21_X1 U13026 ( .B1(n12035), .B2(n14762), .A(n14763), .ZN(n10499) );
  NAND2_X1 U13027 ( .A1(n10499), .A2(n14179), .ZN(n10500) );
  OAI211_X1 U13028 ( .C1(n10502), .C2(n14174), .A(n10501), .B(n10500), .ZN(
        P1_U3285) );
  XNOR2_X1 U13029 ( .A(n10503), .B(n10509), .ZN(n14750) );
  INV_X1 U13030 ( .A(n14750), .ZN(n10516) );
  NAND2_X1 U13031 ( .A1(n14711), .A2(n13945), .ZN(n10504) );
  NAND2_X1 U13032 ( .A1(n10504), .A2(n7114), .ZN(n10505) );
  OR2_X1 U13033 ( .A1(n10505), .A2(n14694), .ZN(n14745) );
  INV_X1 U13034 ( .A(n14745), .ZN(n10508) );
  INV_X1 U13035 ( .A(n13945), .ZN(n10506) );
  OAI22_X1 U13036 ( .A1(n14708), .A2(n10506), .B1(n13944), .B2(n14188), .ZN(
        n10507) );
  AOI21_X1 U13037 ( .B1(n14713), .B2(n10508), .A(n10507), .ZN(n10515) );
  XNOR2_X1 U13038 ( .A(n10510), .B(n10509), .ZN(n10513) );
  NAND2_X1 U13039 ( .A1(n13990), .A2(n14455), .ZN(n10512) );
  NAND2_X1 U13040 ( .A1(n13992), .A2(n14457), .ZN(n10511) );
  NAND2_X1 U13041 ( .A1(n10512), .A2(n10511), .ZN(n13943) );
  AOI21_X1 U13042 ( .B1(n10513), .B2(n14701), .A(n13943), .ZN(n14747) );
  MUX2_X1 U13043 ( .A(n9596), .B(n14747), .S(n14179), .Z(n10514) );
  OAI211_X1 U13044 ( .C1(n10516), .C2(n14174), .A(n10515), .B(n10514), .ZN(
        P1_U3287) );
  XNOR2_X1 U13045 ( .A(n12698), .B(n10517), .ZN(n10522) );
  AOI22_X1 U13046 ( .A1(n13098), .A2(n12763), .B1(n12761), .B2(n13100), .ZN(
        n10521) );
  NAND3_X1 U13047 ( .A1(n10726), .A2(n12698), .A3(n12563), .ZN(n10518) );
  NAND2_X1 U13048 ( .A1(n10519), .A2(n10518), .ZN(n15143) );
  NAND2_X1 U13049 ( .A1(n15143), .A2(n15120), .ZN(n10520) );
  OAI211_X1 U13050 ( .C1(n10522), .C2(n15115), .A(n10521), .B(n10520), .ZN(
        n15141) );
  INV_X1 U13051 ( .A(n15141), .ZN(n10527) );
  AOI22_X1 U13052 ( .A1(n13108), .A2(n10661), .B1(n13092), .B2(n10665), .ZN(
        n10523) );
  OAI21_X1 U13053 ( .B1(n10524), .B2(n13106), .A(n10523), .ZN(n10525) );
  AOI21_X1 U13054 ( .B1(n15143), .B2(n12926), .A(n10525), .ZN(n10526) );
  OAI21_X1 U13055 ( .B1(n10527), .B2(n13116), .A(n10526), .ZN(P3_U3229) );
  INV_X1 U13056 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n10529) );
  MUX2_X1 U13057 ( .A(P1_REG2_REG_10__SCAN_IN), .B(n10529), .S(n11411), .Z(
        n10530) );
  INV_X1 U13058 ( .A(n10530), .ZN(n10531) );
  NOR2_X1 U13059 ( .A1(n10532), .A2(n10531), .ZN(n11403) );
  AOI211_X1 U13060 ( .C1(n10532), .C2(n10531), .A(n14651), .B(n11403), .ZN(
        n10541) );
  INV_X1 U13061 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n10533) );
  MUX2_X1 U13062 ( .A(n10533), .B(P1_REG1_REG_10__SCAN_IN), .S(n11411), .Z(
        n10536) );
  OAI21_X1 U13063 ( .B1(n10563), .B2(P1_REG1_REG_9__SCAN_IN), .A(n10534), .ZN(
        n10535) );
  NOR2_X1 U13064 ( .A1(n10535), .A2(n10536), .ZN(n11410) );
  AOI211_X1 U13065 ( .C1(n10536), .C2(n10535), .A(n14647), .B(n11410), .ZN(
        n10540) );
  NAND2_X1 U13066 ( .A1(n14658), .A2(n11411), .ZN(n10537) );
  NAND2_X1 U13067 ( .A1(P1_REG3_REG_10__SCAN_IN), .A2(P1_U3086), .ZN(n11232)
         );
  OAI211_X1 U13068 ( .C1(n10538), .C2(n14661), .A(n10537), .B(n11232), .ZN(
        n10539) );
  OR3_X1 U13069 ( .A1(n10541), .A2(n10540), .A3(n10539), .ZN(P1_U3253) );
  INV_X1 U13070 ( .A(n10542), .ZN(n10547) );
  XNOR2_X1 U13071 ( .A(n10624), .B(n6485), .ZN(n11760) );
  AND2_X1 U13072 ( .A1(n13392), .A2(n12163), .ZN(n10543) );
  NAND2_X1 U13073 ( .A1(n11760), .A2(n10543), .ZN(n10548) );
  INV_X1 U13074 ( .A(n11760), .ZN(n10545) );
  INV_X1 U13075 ( .A(n10543), .ZN(n10544) );
  NAND2_X1 U13076 ( .A1(n10545), .A2(n10544), .ZN(n10546) );
  AND2_X1 U13077 ( .A1(n10548), .A2(n10546), .ZN(n10595) );
  XNOR2_X1 U13078 ( .A(n11771), .B(n6485), .ZN(n10549) );
  NAND2_X1 U13079 ( .A1(n13391), .A2(n12159), .ZN(n10550) );
  XNOR2_X1 U13080 ( .A(n10549), .B(n10550), .ZN(n11763) );
  INV_X1 U13081 ( .A(n10549), .ZN(n10554) );
  NAND2_X1 U13082 ( .A1(n10554), .A2(n10550), .ZN(n10551) );
  XNOR2_X1 U13083 ( .A(n10779), .B(n12098), .ZN(n10766) );
  NAND2_X1 U13084 ( .A1(n13390), .A2(n12159), .ZN(n10765) );
  XNOR2_X1 U13085 ( .A(n10766), .B(n10765), .ZN(n10556) );
  INV_X1 U13086 ( .A(n13391), .ZN(n10632) );
  NAND2_X1 U13087 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(P2_U3088), .ZN(n14850) );
  OAI21_X1 U13088 ( .B1(n13353), .B2(n10632), .A(n14850), .ZN(n10553) );
  INV_X1 U13089 ( .A(n13389), .ZN(n10842) );
  OAI22_X1 U13090 ( .A1(n13351), .A2(n10842), .B1(n13352), .B2(n10633), .ZN(
        n10552) );
  AOI211_X1 U13091 ( .C1(n10779), .C2(n9820), .A(n10553), .B(n10552), .ZN(
        n10558) );
  OAI22_X1 U13092 ( .A1(n13327), .A2(n10632), .B1(n10554), .B2(n13334), .ZN(
        n10555) );
  NAND3_X1 U13093 ( .A1(n11774), .A2(n10556), .A3(n10555), .ZN(n10557) );
  OAI211_X1 U13094 ( .C1(n6638), .C2(n13334), .A(n10558), .B(n10557), .ZN(
        P2_U3203) );
  INV_X1 U13095 ( .A(n13989), .ZN(n10559) );
  OR2_X1 U13096 ( .A1(n11826), .A2(n10559), .ZN(n10560) );
  NAND2_X1 U13097 ( .A1(n10561), .A2(n10560), .ZN(n14665) );
  INV_X1 U13098 ( .A(n14665), .ZN(n10566) );
  AOI22_X1 U13099 ( .A1(n11430), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n10563), 
        .B2(n6478), .ZN(n10564) );
  INV_X1 U13100 ( .A(n14664), .ZN(n10565) );
  NAND2_X1 U13101 ( .A1(n14672), .A2(n11109), .ZN(n10567) );
  NAND2_X1 U13102 ( .A1(n10568), .A2(n11960), .ZN(n10570) );
  AOI22_X1 U13103 ( .A1(n11411), .A2(n6478), .B1(n11430), .B2(
        P2_DATAO_REG_10__SCAN_IN), .ZN(n10569) );
  NAND2_X1 U13104 ( .A1(n11587), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n10577) );
  NAND2_X1 U13105 ( .A1(n11616), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n10576) );
  AND2_X1 U13106 ( .A1(n10572), .A2(n10571), .ZN(n10573) );
  NOR2_X1 U13107 ( .A1(n10582), .A2(n10573), .ZN(n11231) );
  NAND2_X1 U13108 ( .A1(n9893), .A2(n11231), .ZN(n10575) );
  NAND2_X1 U13109 ( .A1(n11526), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n10574) );
  NAND4_X1 U13110 ( .A1(n10577), .A2(n10576), .A3(n10575), .A4(n10574), .ZN(
        n14458) );
  INV_X1 U13111 ( .A(n14458), .ZN(n10956) );
  XNOR2_X1 U13112 ( .A(n14778), .B(n10956), .ZN(n12006) );
  XNOR2_X1 U13113 ( .A(n10957), .B(n12006), .ZN(n14781) );
  OR2_X1 U13114 ( .A1(n14706), .A2(n14780), .ZN(n14135) );
  OR2_X1 U13115 ( .A1(n14672), .A2(n13988), .ZN(n10580) );
  NAND2_X1 U13116 ( .A1(n10581), .A2(n10580), .ZN(n10936) );
  XNOR2_X1 U13117 ( .A(n10936), .B(n12006), .ZN(n14784) );
  NAND2_X1 U13118 ( .A1(n14784), .A2(n14483), .ZN(n10593) );
  INV_X1 U13119 ( .A(n14778), .ZN(n10953) );
  XNOR2_X1 U13120 ( .A(n14676), .B(n10953), .ZN(n10588) );
  NAND2_X1 U13121 ( .A1(n10582), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n10947) );
  OR2_X1 U13122 ( .A1(n10582), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n10583) );
  NAND2_X1 U13123 ( .A1(n10947), .A2(n10583), .ZN(n14468) );
  INV_X1 U13124 ( .A(n14468), .ZN(n14475) );
  NAND2_X1 U13125 ( .A1(n6475), .A2(n14475), .ZN(n10587) );
  NAND2_X1 U13126 ( .A1(n11616), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n10586) );
  NAND2_X1 U13127 ( .A1(n11526), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n10585) );
  NAND2_X1 U13128 ( .A1(n11587), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n10584) );
  NAND4_X1 U13129 ( .A1(n10587), .A2(n10586), .A3(n10585), .A4(n10584), .ZN(
        n13987) );
  OAI22_X1 U13130 ( .A1(n10588), .A2(n14493), .B1(n11234), .B2(n14167), .ZN(
        n14775) );
  NOR2_X1 U13131 ( .A1(n11109), .A2(n14169), .ZN(n14776) );
  AOI22_X1 U13132 ( .A1(n14179), .A2(n14776), .B1(n11231), .B2(n14704), .ZN(
        n10590) );
  NAND2_X1 U13133 ( .A1(n14681), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n10589) );
  OAI211_X1 U13134 ( .C1(n10953), .C2(n14708), .A(n10590), .B(n10589), .ZN(
        n10591) );
  AOI21_X1 U13135 ( .B1(n14775), .B2(n14713), .A(n10591), .ZN(n10592) );
  OAI211_X1 U13136 ( .C1(n14781), .C2(n14135), .A(n10593), .B(n10592), .ZN(
        P1_U3283) );
  NAND3_X1 U13137 ( .A1(n13347), .A2(n13393), .A3(n10594), .ZN(n10599) );
  OAI21_X1 U13138 ( .B1(n10596), .B2(n10595), .A(n13359), .ZN(n10598) );
  INV_X1 U13139 ( .A(n11762), .ZN(n10597) );
  AOI21_X1 U13140 ( .B1(n10599), .B2(n10598), .A(n10597), .ZN(n10604) );
  OAI22_X1 U13141 ( .A1(n13353), .A2(n11709), .B1(n13352), .B2(n10600), .ZN(
        n10603) );
  AOI22_X1 U13142 ( .A1(n11753), .A2(n13391), .B1(P2_REG3_REG_7__SCAN_IN), 
        .B2(P2_U3088), .ZN(n10601) );
  OAI21_X1 U13143 ( .B1(n14962), .B2(n13371), .A(n10601), .ZN(n10602) );
  OR3_X1 U13144 ( .A1(n10604), .A2(n10603), .A3(n10602), .ZN(P2_U3185) );
  INV_X1 U13145 ( .A(n10605), .ZN(n10607) );
  OAI22_X1 U13146 ( .A1(n12739), .A2(P3_U3151), .B1(SI_22_), .B2(n13247), .ZN(
        n10606) );
  AOI21_X1 U13147 ( .B1(n10607), .B2(n14317), .A(n10606), .ZN(P3_U3273) );
  INV_X1 U13148 ( .A(n10608), .ZN(n10611) );
  AOI211_X1 U13149 ( .C1(n10611), .C2(n14149), .A(n10610), .B(n10609), .ZN(
        n10617) );
  AOI22_X1 U13150 ( .A1(n14706), .A2(P1_REG2_REG_4__SCAN_IN), .B1(n10612), 
        .B2(n14704), .ZN(n10613) );
  OAI21_X1 U13151 ( .B1(n14708), .B2(n10484), .A(n10613), .ZN(n10614) );
  AOI21_X1 U13152 ( .B1(n10615), .B2(n14483), .A(n10614), .ZN(n10616) );
  OAI21_X1 U13153 ( .B1(n10617), .B2(n14706), .A(n10616), .ZN(P1_U3289) );
  NAND2_X1 U13154 ( .A1(n10624), .A2(n13392), .ZN(n10618) );
  NAND2_X1 U13155 ( .A1(n11771), .A2(n13391), .ZN(n10620) );
  INV_X1 U13156 ( .A(n10777), .ZN(n10630) );
  NAND2_X1 U13157 ( .A1(n10621), .A2(n10630), .ZN(n10775) );
  OAI21_X1 U13158 ( .B1(n10621), .B2(n10630), .A(n10775), .ZN(n14977) );
  OR2_X1 U13159 ( .A1(n10624), .A2(n11766), .ZN(n10622) );
  NAND2_X1 U13160 ( .A1(n10623), .A2(n10622), .ZN(n10626) );
  NAND2_X1 U13161 ( .A1(n10624), .A2(n11766), .ZN(n10625) );
  NAND2_X1 U13162 ( .A1(n10626), .A2(n10625), .ZN(n11497) );
  NAND2_X1 U13163 ( .A1(n11497), .A2(n10627), .ZN(n10629) );
  NAND2_X1 U13164 ( .A1(n11771), .A2(n10632), .ZN(n10628) );
  NAND2_X1 U13165 ( .A1(n10629), .A2(n10628), .ZN(n10778) );
  XNOR2_X1 U13166 ( .A(n10778), .B(n10630), .ZN(n10631) );
  OAI222_X1 U13167 ( .A1(n13657), .A2(n10842), .B1(n13655), .B2(n10632), .C1(
        n13594), .C2(n10631), .ZN(n14980) );
  NAND2_X1 U13168 ( .A1(n14980), .A2(n13606), .ZN(n10638) );
  OAI22_X1 U13169 ( .A1(n13606), .A2(n10634), .B1(n10633), .B2(n13607), .ZN(
        n10636) );
  INV_X1 U13170 ( .A(n11771), .ZN(n14970) );
  INV_X1 U13171 ( .A(n10779), .ZN(n14978) );
  NAND2_X1 U13172 ( .A1(n11507), .A2(n14978), .ZN(n10799) );
  OAI21_X1 U13173 ( .B1(n11507), .B2(n14978), .A(n10799), .ZN(n14979) );
  NOR2_X1 U13174 ( .A1(n14979), .A2(n11660), .ZN(n10635) );
  AOI211_X1 U13175 ( .C1(n13553), .C2(n10779), .A(n10636), .B(n10635), .ZN(
        n10637) );
  OAI211_X1 U13176 ( .C1(n13649), .C2(n14977), .A(n10638), .B(n10637), .ZN(
        P2_U3256) );
  NAND2_X1 U13177 ( .A1(n12765), .A2(P3_DATAO_REG_30__SCAN_IN), .ZN(n10639) );
  OAI21_X1 U13178 ( .B1(n12529), .B2(n12765), .A(n10639), .ZN(P3_U3521) );
  INV_X1 U13179 ( .A(n13946), .ZN(n10826) );
  NAND2_X1 U13180 ( .A1(n14777), .A2(n11807), .ZN(n14737) );
  NAND2_X1 U13181 ( .A1(n13991), .A2(n14455), .ZN(n10641) );
  NAND2_X1 U13182 ( .A1(n13993), .A2(n14457), .ZN(n10640) );
  NAND2_X1 U13183 ( .A1(n10641), .A2(n10640), .ZN(n14735) );
  NAND2_X1 U13184 ( .A1(n14466), .A2(n14735), .ZN(n10643) );
  OAI211_X1 U13185 ( .C1(n10826), .C2(n14737), .A(n10643), .B(n10642), .ZN(
        n10655) );
  INV_X1 U13186 ( .A(n10644), .ZN(n10646) );
  OAI22_X1 U13187 ( .A1(n6904), .A2(n9342), .B1(n12223), .B2(n10650), .ZN(
        n10649) );
  XNOR2_X1 U13188 ( .A(n10649), .B(n11452), .ZN(n10652) );
  OAI22_X1 U13189 ( .A1(n12276), .A2(n10650), .B1(n6904), .B2(n12223), .ZN(
        n10651) );
  NAND2_X1 U13190 ( .A1(n10652), .A2(n10651), .ZN(n10740) );
  NOR2_X1 U13191 ( .A1(n10653), .A2(n13938), .ZN(n10654) );
  AOI211_X1 U13192 ( .C1(n14705), .C2(n13955), .A(n10655), .B(n10654), .ZN(
        n10656) );
  INV_X1 U13193 ( .A(n10656), .ZN(P1_U3227) );
  INV_X1 U13194 ( .A(n10657), .ZN(n10658) );
  AOI21_X1 U13195 ( .B1(n10660), .B2(n10659), .A(n10658), .ZN(n10667) );
  AOI22_X1 U13196 ( .A1(n12441), .A2(n12763), .B1(n12471), .B2(n12761), .ZN(
        n10663) );
  AOI22_X1 U13197 ( .A1(n12476), .A2(n10661), .B1(P3_REG3_REG_4__SCAN_IN), 
        .B2(P3_U3151), .ZN(n10662) );
  NAND2_X1 U13198 ( .A1(n10663), .A2(n10662), .ZN(n10664) );
  AOI21_X1 U13199 ( .B1(n10665), .B2(n12497), .A(n10664), .ZN(n10666) );
  OAI21_X1 U13200 ( .B1(n10667), .B2(n12478), .A(n10666), .ZN(P3_U3170) );
  OAI22_X1 U13201 ( .A1(n14681), .A2(n10668), .B1(P1_REG3_REG_3__SCAN_IN), 
        .B2(n14188), .ZN(n10671) );
  NOR2_X1 U13202 ( .A1(n14708), .A2(n10669), .ZN(n10670) );
  AOI211_X1 U13203 ( .C1(n14706), .C2(P1_REG2_REG_3__SCAN_IN), .A(n10671), .B(
        n10670), .ZN(n10672) );
  OAI21_X1 U13204 ( .B1(n11701), .B2(n10673), .A(n10672), .ZN(n10674) );
  AOI21_X1 U13205 ( .B1(n14483), .B2(n10675), .A(n10674), .ZN(n10676) );
  OAI21_X1 U13206 ( .B1(n14135), .B2(n10677), .A(n10676), .ZN(P1_U3290) );
  INV_X1 U13207 ( .A(n11373), .ZN(n10681) );
  OAI222_X1 U13208 ( .A1(n13822), .A2(n10678), .B1(n13820), .B2(n10681), .C1(
        P2_U3088), .C2(n13479), .ZN(P2_U3309) );
  NAND2_X1 U13209 ( .A1(n10679), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10680) );
  XNOR2_X1 U13210 ( .A(n10680), .B(P1_IR_REG_18__SCAN_IN), .ZN(n14657) );
  INV_X1 U13211 ( .A(n14657), .ZN(n14043) );
  OAI222_X1 U13212 ( .A1(n14292), .A2(n10682), .B1(n12152), .B2(n10681), .C1(
        P1_U3086), .C2(n14043), .ZN(P1_U3337) );
  NAND2_X1 U13213 ( .A1(n10683), .A2(n12701), .ZN(n10684) );
  AND2_X1 U13214 ( .A1(n10879), .A2(n10684), .ZN(n10688) );
  XNOR2_X1 U13215 ( .A(n10685), .B(n12701), .ZN(n15145) );
  NAND2_X1 U13216 ( .A1(n15145), .A2(n15120), .ZN(n10687) );
  AOI22_X1 U13217 ( .A1(n13098), .A2(n12762), .B1(n12760), .B2(n13100), .ZN(
        n10686) );
  OAI211_X1 U13218 ( .C1(n10688), .C2(n15115), .A(n10687), .B(n10686), .ZN(
        n15149) );
  INV_X1 U13219 ( .A(n15149), .ZN(n10692) );
  AOI22_X1 U13220 ( .A1(n13108), .A2(n10755), .B1(n13092), .B2(n10759), .ZN(
        n10689) );
  OAI21_X1 U13221 ( .B1(n10072), .B2(n13106), .A(n10689), .ZN(n10690) );
  AOI21_X1 U13222 ( .B1(n15145), .B2(n12926), .A(n10690), .ZN(n10691) );
  OAI21_X1 U13223 ( .B1(n10692), .B2(n13116), .A(n10691), .ZN(P3_U3228) );
  INV_X1 U13224 ( .A(P3_REG2_REG_9__SCAN_IN), .ZN(n15081) );
  NOR2_X1 U13225 ( .A1(n10714), .A2(n10694), .ZN(n10695) );
  INV_X1 U13226 ( .A(P3_REG2_REG_10__SCAN_IN), .ZN(n10696) );
  AOI22_X1 U13227 ( .A1(n11025), .A2(P3_REG2_REG_10__SCAN_IN), .B1(n10696), 
        .B2(n11021), .ZN(n10697) );
  AOI21_X1 U13228 ( .B1(n6636), .B2(n10697), .A(n11020), .ZN(n10723) );
  INV_X1 U13229 ( .A(P3_REG1_REG_10__SCAN_IN), .ZN(n13178) );
  AOI22_X1 U13230 ( .A1(n11025), .A2(n13178), .B1(P3_REG1_REG_10__SCAN_IN), 
        .B2(n11021), .ZN(n10703) );
  NAND2_X1 U13231 ( .A1(n15089), .A2(n10700), .ZN(n10701) );
  NAND2_X1 U13232 ( .A1(P3_REG1_REG_9__SCAN_IN), .A2(n15096), .ZN(n15095) );
  OAI21_X1 U13233 ( .B1(n10703), .B2(n10702), .A(n11024), .ZN(n10708) );
  NOR2_X1 U13234 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n10704), .ZN(n10705) );
  AOI21_X1 U13235 ( .B1(n15094), .B2(P3_ADDR_REG_10__SCAN_IN), .A(n10705), 
        .ZN(n10706) );
  OAI21_X1 U13236 ( .B1(n15088), .B2(n11021), .A(n10706), .ZN(n10707) );
  AOI21_X1 U13237 ( .B1(n10708), .B2(n15097), .A(n10707), .ZN(n10722) );
  OAI22_X1 U13238 ( .A1(n10712), .A2(n10711), .B1(n10710), .B2(n10709), .ZN(
        n15083) );
  MUX2_X1 U13239 ( .A(P3_REG2_REG_9__SCAN_IN), .B(P3_REG1_REG_9__SCAN_IN), .S(
        n12836), .Z(n10713) );
  NAND2_X1 U13240 ( .A1(n10713), .A2(n15089), .ZN(n15084) );
  NAND2_X1 U13241 ( .A1(n15083), .A2(n15084), .ZN(n15082) );
  INV_X1 U13242 ( .A(n10713), .ZN(n10715) );
  NAND2_X1 U13243 ( .A1(n10715), .A2(n10714), .ZN(n15086) );
  MUX2_X1 U13244 ( .A(n10696), .B(n13178), .S(n12836), .Z(n10716) );
  NAND2_X1 U13245 ( .A1(n10716), .A2(n11025), .ZN(n11028) );
  INV_X1 U13246 ( .A(n10716), .ZN(n10717) );
  NAND2_X1 U13247 ( .A1(n10717), .A2(n11021), .ZN(n10718) );
  NAND2_X1 U13248 ( .A1(n11028), .A2(n10718), .ZN(n10719) );
  AOI21_X1 U13249 ( .B1(n15082), .B2(n15086), .A(n10719), .ZN(n11030) );
  AND3_X1 U13250 ( .A1(n15082), .A2(n15086), .A3(n10719), .ZN(n10720) );
  OAI21_X1 U13251 ( .B1(n11030), .B2(n10720), .A(n15064), .ZN(n10721) );
  OAI211_X1 U13252 ( .C1(n10723), .C2(n15101), .A(n10722), .B(n10721), .ZN(
        P3_U3192) );
  OR2_X1 U13253 ( .A1(n10724), .A2(n12705), .ZN(n10725) );
  NAND2_X1 U13254 ( .A1(n10726), .A2(n10725), .ZN(n15138) );
  OAI22_X1 U13255 ( .A1(n13094), .A2(n15135), .B1(P3_REG3_REG_3__SCAN_IN), 
        .B2(n15108), .ZN(n10735) );
  AOI21_X1 U13256 ( .B1(n15117), .B2(n10728), .A(n10727), .ZN(n10733) );
  NAND2_X1 U13257 ( .A1(n10729), .A2(n13103), .ZN(n10732) );
  NAND2_X1 U13258 ( .A1(n15138), .A2(n15120), .ZN(n10731) );
  AOI22_X1 U13259 ( .A1(n13098), .A2(n6469), .B1(n12762), .B2(n13100), .ZN(
        n10730) );
  OAI211_X1 U13260 ( .C1(n10733), .C2(n10732), .A(n10731), .B(n10730), .ZN(
        n15136) );
  MUX2_X1 U13261 ( .A(n15136), .B(P3_REG2_REG_3__SCAN_IN), .S(n13043), .Z(
        n10734) );
  AOI211_X1 U13262 ( .C1(n12926), .C2(n15138), .A(n10735), .B(n10734), .ZN(
        n10736) );
  INV_X1 U13263 ( .A(n10736), .ZN(P3_U3230) );
  AOI22_X1 U13264 ( .A1(n12301), .A2(n13991), .B1(n10746), .B2(n13945), .ZN(
        n10742) );
  NAND2_X1 U13265 ( .A1(n13945), .A2(n12303), .ZN(n10738) );
  NAND2_X1 U13266 ( .A1(n10746), .A2(n13991), .ZN(n10737) );
  NAND2_X1 U13267 ( .A1(n10738), .A2(n10737), .ZN(n10739) );
  XNOR2_X1 U13268 ( .A(n10739), .B(n11452), .ZN(n10741) );
  XNOR2_X1 U13269 ( .A(n10742), .B(n10741), .ZN(n13941) );
  NAND2_X1 U13270 ( .A1(n13942), .A2(n13941), .ZN(n13940) );
  NAND2_X1 U13271 ( .A1(n11817), .A2(n12303), .ZN(n10744) );
  NAND2_X1 U13272 ( .A1(n10746), .A2(n13990), .ZN(n10743) );
  NAND2_X1 U13273 ( .A1(n10744), .A2(n10743), .ZN(n10745) );
  XNOR2_X1 U13274 ( .A(n10745), .B(n11452), .ZN(n10819) );
  AOI22_X1 U13275 ( .A1(n11817), .A2(n10746), .B1(n12301), .B2(n13990), .ZN(
        n10820) );
  XNOR2_X1 U13276 ( .A(n10819), .B(n10820), .ZN(n10747) );
  OAI211_X1 U13277 ( .C1(n10748), .C2(n10747), .A(n10823), .B(n14465), .ZN(
        n10752) );
  AOI22_X1 U13278 ( .A1(n14457), .A2(n13991), .B1(n13989), .B2(n14455), .ZN(
        n14683) );
  INV_X1 U13279 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n10749) );
  OAI22_X1 U13280 ( .A1(n13934), .A2(n14683), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n10749), .ZN(n10750) );
  AOI21_X1 U13281 ( .B1(n14690), .B2(n13955), .A(n10750), .ZN(n10751) );
  OAI211_X1 U13282 ( .C1(n14754), .C2(n13972), .A(n10752), .B(n10751), .ZN(
        P1_U3213) );
  XOR2_X1 U13283 ( .A(n10754), .B(n10753), .Z(n10761) );
  AOI22_X1 U13284 ( .A1(n12441), .A2(n12762), .B1(n12471), .B2(n12760), .ZN(
        n10757) );
  AOI22_X1 U13285 ( .A1(n12476), .A2(n10755), .B1(P3_REG3_REG_5__SCAN_IN), 
        .B2(P3_U3151), .ZN(n10756) );
  NAND2_X1 U13286 ( .A1(n10757), .A2(n10756), .ZN(n10758) );
  AOI21_X1 U13287 ( .B1(n10759), .B2(n12497), .A(n10758), .ZN(n10760) );
  OAI21_X1 U13288 ( .B1(n10761), .B2(n12478), .A(n10760), .ZN(P3_U3167) );
  NAND2_X1 U13289 ( .A1(n10762), .A2(n14317), .ZN(n10763) );
  OAI211_X1 U13290 ( .C1(n9113), .C2(n13247), .A(n10763), .B(n12741), .ZN(
        P3_U3272) );
  INV_X1 U13291 ( .A(n11428), .ZN(n11653) );
  OAI222_X1 U13292 ( .A1(n13822), .A2(n10764), .B1(n13820), .B2(n11653), .C1(
        P2_U3088), .C2(n13680), .ZN(P2_U3308) );
  INV_X1 U13293 ( .A(n14987), .ZN(n10803) );
  XNOR2_X1 U13294 ( .A(n14987), .B(n12098), .ZN(n10834) );
  NAND2_X1 U13295 ( .A1(n13389), .A2(n12159), .ZN(n10767) );
  NOR2_X1 U13296 ( .A1(n10834), .A2(n10767), .ZN(n10837) );
  AOI21_X1 U13297 ( .B1(n10834), .B2(n10767), .A(n10837), .ZN(n10768) );
  OAI211_X1 U13298 ( .C1(n10769), .C2(n10768), .A(n10840), .B(n13359), .ZN(
        n10773) );
  NAND2_X1 U13299 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(P2_U3088), .ZN(n14864)
         );
  INV_X1 U13300 ( .A(n14864), .ZN(n10771) );
  OAI22_X1 U13301 ( .A1(n13353), .A2(n11768), .B1(n13352), .B2(n10800), .ZN(
        n10770) );
  AOI211_X1 U13302 ( .C1(n11753), .C2(n13388), .A(n10771), .B(n10770), .ZN(
        n10772) );
  OAI211_X1 U13303 ( .C1(n10803), .C2(n13371), .A(n10773), .B(n10772), .ZN(
        P2_U3189) );
  NAND2_X1 U13304 ( .A1(n10779), .A2(n13390), .ZN(n10774) );
  NAND2_X1 U13305 ( .A1(n10775), .A2(n10774), .ZN(n10852) );
  INV_X1 U13306 ( .A(n10794), .ZN(n10850) );
  NAND2_X1 U13307 ( .A1(n10852), .A2(n10850), .ZN(n10805) );
  NAND2_X1 U13308 ( .A1(n14987), .A2(n13389), .ZN(n10856) );
  NAND2_X1 U13309 ( .A1(n10805), .A2(n10856), .ZN(n10776) );
  XOR2_X1 U13310 ( .A(n10860), .B(n10776), .Z(n15001) );
  INV_X1 U13311 ( .A(n15001), .ZN(n10793) );
  NAND2_X1 U13312 ( .A1(n10778), .A2(n10777), .ZN(n10781) );
  NAND2_X1 U13313 ( .A1(n10779), .A2(n11768), .ZN(n10780) );
  NAND2_X1 U13314 ( .A1(n10781), .A2(n10780), .ZN(n10795) );
  AND2_X1 U13315 ( .A1(n14987), .A2(n10842), .ZN(n10782) );
  AOI21_X1 U13316 ( .B1(n10795), .B2(n10794), .A(n10782), .ZN(n10861) );
  XNOR2_X1 U13317 ( .A(n10861), .B(n10860), .ZN(n10783) );
  NAND2_X1 U13318 ( .A1(n10783), .A2(n13677), .ZN(n10785) );
  AOI22_X1 U13319 ( .A1(n13640), .A2(n13389), .B1(n13387), .B2(n13642), .ZN(
        n10784) );
  NAND2_X1 U13320 ( .A1(n10785), .A2(n10784), .ZN(n14999) );
  INV_X1 U13321 ( .A(n10854), .ZN(n14995) );
  INV_X1 U13322 ( .A(n10864), .ZN(n10787) );
  OAI21_X1 U13323 ( .B1(n14995), .B2(n6677), .A(n10787), .ZN(n14997) );
  OAI22_X1 U13324 ( .A1(n13606), .A2(n10788), .B1(n10843), .B2(n13607), .ZN(
        n10789) );
  AOI21_X1 U13325 ( .B1(n10854), .B2(n13553), .A(n10789), .ZN(n10790) );
  OAI21_X1 U13326 ( .B1(n14997), .B2(n11660), .A(n10790), .ZN(n10791) );
  AOI21_X1 U13327 ( .B1(n14999), .B2(n13606), .A(n10791), .ZN(n10792) );
  OAI21_X1 U13328 ( .B1(n10793), .B2(n13649), .A(n10792), .ZN(P2_U3254) );
  XNOR2_X1 U13329 ( .A(n10795), .B(n10794), .ZN(n10796) );
  NAND2_X1 U13330 ( .A1(n10796), .A2(n13677), .ZN(n10798) );
  AOI22_X1 U13331 ( .A1(n13642), .A2(n13388), .B1(n13390), .B2(n13640), .ZN(
        n10797) );
  XNOR2_X1 U13332 ( .A(n10799), .B(n10803), .ZN(n14989) );
  INV_X1 U13333 ( .A(n10800), .ZN(n10801) );
  AOI22_X1 U13334 ( .A1(n13671), .A2(P2_REG2_REG_10__SCAN_IN), .B1(n10801), 
        .B2(n13685), .ZN(n10802) );
  OAI21_X1 U13335 ( .B1(n10803), .B2(n13688), .A(n10802), .ZN(n10807) );
  OR2_X1 U13336 ( .A1(n10852), .A2(n10850), .ZN(n10804) );
  NAND2_X1 U13337 ( .A1(n10805), .A2(n10804), .ZN(n14985) );
  NOR2_X1 U13338 ( .A1(n14985), .A2(n13649), .ZN(n10806) );
  AOI211_X1 U13339 ( .C1(n13669), .C2(n14989), .A(n10807), .B(n10806), .ZN(
        n10808) );
  OAI21_X1 U13340 ( .B1(n13671), .B2(n14991), .A(n10808), .ZN(P2_U3255) );
  INV_X1 U13341 ( .A(n10884), .ZN(n10817) );
  AOI21_X1 U13342 ( .B1(n10810), .B2(n10809), .A(n12478), .ZN(n10812) );
  NAND2_X1 U13343 ( .A1(n10812), .A2(n10811), .ZN(n10816) );
  OAI22_X1 U13344 ( .A1(n12443), .A2(n12587), .B1(n10876), .B2(n12474), .ZN(
        n10813) );
  AOI211_X1 U13345 ( .C1(n12476), .C2(n15151), .A(n10814), .B(n10813), .ZN(
        n10815) );
  OAI211_X1 U13346 ( .C1(n10817), .C2(n12452), .A(n10816), .B(n10815), .ZN(
        P3_U3179) );
  AOI22_X1 U13347 ( .A1(n11826), .A2(n12303), .B1(n10746), .B2(n13989), .ZN(
        n10818) );
  XNOR2_X1 U13348 ( .A(n10818), .B(n11452), .ZN(n11107) );
  AOI22_X1 U13349 ( .A1(n11826), .A2(n10746), .B1(n12301), .B2(n13989), .ZN(
        n11106) );
  XNOR2_X1 U13350 ( .A(n11107), .B(n11106), .ZN(n10825) );
  INV_X1 U13351 ( .A(n10820), .ZN(n10821) );
  AOI21_X1 U13352 ( .B1(n10825), .B2(n10824), .A(n11108), .ZN(n10833) );
  NAND2_X1 U13353 ( .A1(n11826), .A2(n14777), .ZN(n14761) );
  NOR2_X1 U13354 ( .A1(n10826), .A2(n14761), .ZN(n10830) );
  OAI22_X1 U13355 ( .A1(n13934), .A2(n10828), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n10827), .ZN(n10829) );
  AOI211_X1 U13356 ( .C1(n10831), .C2(n13955), .A(n10830), .B(n10829), .ZN(
        n10832) );
  OAI21_X1 U13357 ( .B1(n10833), .B2(n13938), .A(n10832), .ZN(P1_U3221) );
  INV_X1 U13358 ( .A(n10840), .ZN(n10836) );
  NOR3_X1 U13359 ( .A1(n10834), .A2(n13327), .A3(n10842), .ZN(n10835) );
  AOI21_X1 U13360 ( .B1(n10836), .B2(n13359), .A(n10835), .ZN(n10849) );
  XNOR2_X1 U13361 ( .A(n10854), .B(n6485), .ZN(n11724) );
  NAND2_X1 U13362 ( .A1(n13388), .A2(n12159), .ZN(n11087) );
  XNOR2_X1 U13363 ( .A(n11724), .B(n11087), .ZN(n10848) );
  INV_X1 U13364 ( .A(n10837), .ZN(n10838) );
  INV_X1 U13365 ( .A(n11090), .ZN(n11727) );
  NAND2_X1 U13366 ( .A1(n11727), .A2(n13359), .ZN(n10847) );
  OAI21_X1 U13367 ( .B1(n13353), .B2(n10842), .A(n10841), .ZN(n10845) );
  OAI22_X1 U13368 ( .A1(n13351), .A2(n11123), .B1(n13352), .B2(n10843), .ZN(
        n10844) );
  AOI211_X1 U13369 ( .C1(n10854), .C2(n9820), .A(n10845), .B(n10844), .ZN(
        n10846) );
  OAI211_X1 U13370 ( .C1(n10849), .C2(n10848), .A(n10847), .B(n10846), .ZN(
        P2_U3208) );
  OR2_X1 U13371 ( .A1(n10854), .A2(n13388), .ZN(n10853) );
  AND2_X1 U13372 ( .A1(n10850), .A2(n10853), .ZN(n10851) );
  INV_X1 U13373 ( .A(n10853), .ZN(n10858) );
  NAND2_X1 U13374 ( .A1(n10854), .A2(n13388), .ZN(n10855) );
  AND2_X1 U13375 ( .A1(n10856), .A2(n10855), .ZN(n10857) );
  OR2_X1 U13376 ( .A1(n10858), .A2(n10857), .ZN(n10859) );
  XNOR2_X1 U13377 ( .A(n11121), .B(n10862), .ZN(n10904) );
  XOR2_X1 U13378 ( .A(n10862), .B(n11127), .Z(n10863) );
  AOI222_X1 U13379 ( .A1(n13645), .A2(n10863), .B1(n13386), .B2(n13642), .C1(
        n13388), .C2(n13640), .ZN(n10903) );
  OR2_X1 U13380 ( .A1(n10903), .A2(n13671), .ZN(n10870) );
  NOR2_X1 U13381 ( .A1(n10864), .A2(n11124), .ZN(n10865) );
  NOR2_X1 U13382 ( .A1(n11124), .A2(n13688), .ZN(n10868) );
  INV_X1 U13383 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n10866) );
  OAI22_X1 U13384 ( .A1(n13606), .A2(n10866), .B1(n11719), .B2(n13607), .ZN(
        n10867) );
  AOI211_X1 U13385 ( .C1(n6634), .C2(n13669), .A(n10868), .B(n10867), .ZN(
        n10869) );
  OAI211_X1 U13386 ( .C1(n10904), .C2(n13649), .A(n10870), .B(n10869), .ZN(
        P2_U3253) );
  INV_X1 U13387 ( .A(n11469), .ZN(n10901) );
  OAI222_X1 U13388 ( .A1(n13822), .A2(n10872), .B1(n13820), .B2(n10901), .C1(
        n10871), .C2(P2_U3088), .ZN(P2_U3307) );
  OAI21_X1 U13389 ( .B1(n10875), .B2(n10874), .A(n10873), .ZN(n15153) );
  INV_X1 U13390 ( .A(n15153), .ZN(n10887) );
  OAI22_X1 U13391 ( .A1(n10876), .A2(n15109), .B1(n12587), .B2(n15111), .ZN(
        n10883) );
  INV_X1 U13392 ( .A(n10877), .ZN(n10881) );
  AOI21_X1 U13393 ( .B1(n10879), .B2(n10878), .A(n12704), .ZN(n10880) );
  NOR3_X1 U13394 ( .A1(n10881), .A2(n10880), .A3(n15115), .ZN(n10882) );
  AOI211_X1 U13395 ( .C1(n15120), .C2(n15153), .A(n10883), .B(n10882), .ZN(
        n15155) );
  MUX2_X1 U13396 ( .A(n10095), .B(n15155), .S(n13106), .Z(n10886) );
  AOI22_X1 U13397 ( .A1(n13108), .A2(n15151), .B1(n13092), .B2(n10884), .ZN(
        n10885) );
  OAI211_X1 U13398 ( .C1(n10887), .C2(n11074), .A(n10886), .B(n10885), .ZN(
        P3_U3227) );
  OR2_X1 U13399 ( .A1(n10888), .A2(n12706), .ZN(n10889) );
  NAND2_X1 U13400 ( .A1(n10890), .A2(n10889), .ZN(n15160) );
  INV_X1 U13401 ( .A(n15160), .ZN(n10900) );
  XNOR2_X1 U13402 ( .A(n10892), .B(n10891), .ZN(n10895) );
  NAND2_X1 U13403 ( .A1(n15160), .A2(n15120), .ZN(n10894) );
  AOI22_X1 U13404 ( .A1(n13098), .A2(n12760), .B1(n12758), .B2(n13100), .ZN(
        n10893) );
  OAI211_X1 U13405 ( .C1(n15115), .C2(n10895), .A(n10894), .B(n10893), .ZN(
        n15158) );
  NAND2_X1 U13406 ( .A1(n15158), .A2(n13106), .ZN(n10899) );
  INV_X1 U13407 ( .A(n12322), .ZN(n10896) );
  OAI22_X1 U13408 ( .A1(n13094), .A2(n15157), .B1(n10896), .B2(n15108), .ZN(
        n10897) );
  AOI21_X1 U13409 ( .B1(P3_REG2_REG_7__SCAN_IN), .B2(n13116), .A(n10897), .ZN(
        n10898) );
  OAI211_X1 U13410 ( .C1(n10900), .C2(n11074), .A(n10899), .B(n10898), .ZN(
        P3_U3226) );
  INV_X1 U13411 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n11470) );
  OAI222_X1 U13412 ( .A1(n14292), .A2(n11470), .B1(P1_U3086), .B2(n11972), 
        .C1(n12152), .C2(n10901), .ZN(P1_U3335) );
  INV_X1 U13413 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n10906) );
  AOI22_X1 U13414 ( .A1(n6634), .A2(n14988), .B1(n11730), .B2(n14986), .ZN(
        n10902) );
  OAI211_X1 U13415 ( .C1(n14984), .C2(n10904), .A(n10903), .B(n10902), .ZN(
        n10907) );
  NAND2_X1 U13416 ( .A1(n10907), .A2(n14953), .ZN(n10905) );
  OAI21_X1 U13417 ( .B1(n15004), .B2(n10906), .A(n10905), .ZN(P2_U3466) );
  NAND2_X1 U13418 ( .A1(n10907), .A2(n15019), .ZN(n10908) );
  OAI21_X1 U13419 ( .B1(n15019), .B2(n9867), .A(n10908), .ZN(P2_U3511) );
  INV_X1 U13420 ( .A(n10909), .ZN(n10911) );
  OAI222_X1 U13421 ( .A1(P3_U3151), .A2(n10912), .B1(n13250), .B2(n10911), 
        .C1(n10910), .C2(n13247), .ZN(P3_U3271) );
  OAI21_X1 U13422 ( .B1(P2_REG2_REG_12__SCAN_IN), .B2(n10925), .A(n10913), 
        .ZN(n14868) );
  XNOR2_X1 U13423 ( .A(n14875), .B(P2_REG2_REG_13__SCAN_IN), .ZN(n14869) );
  NOR2_X1 U13424 ( .A1(n14868), .A2(n14869), .ZN(n14867) );
  AOI21_X1 U13425 ( .B1(n14875), .B2(P2_REG2_REG_13__SCAN_IN), .A(n14867), 
        .ZN(n10915) );
  NOR2_X1 U13426 ( .A1(n10915), .A2(n10914), .ZN(n10917) );
  AOI21_X1 U13427 ( .B1(n10915), .B2(n10914), .A(n10917), .ZN(n10916) );
  INV_X1 U13428 ( .A(n10916), .ZN(n14881) );
  INV_X1 U13429 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n14882) );
  NOR2_X1 U13430 ( .A1(n14881), .A2(n14882), .ZN(n14879) );
  NOR2_X1 U13431 ( .A1(n10917), .A2(n14879), .ZN(n10918) );
  NOR2_X1 U13432 ( .A1(n10918), .A2(n14904), .ZN(n10919) );
  XNOR2_X1 U13433 ( .A(n14904), .B(n10918), .ZN(n14900) );
  NOR2_X1 U13434 ( .A1(n14899), .A2(n14900), .ZN(n14898) );
  NOR2_X1 U13435 ( .A1(n10919), .A2(n14898), .ZN(n10923) );
  INV_X1 U13436 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n10920) );
  MUX2_X1 U13437 ( .A(P2_REG2_REG_16__SCAN_IN), .B(n10920), .S(n13467), .Z(
        n10921) );
  INV_X1 U13438 ( .A(n10921), .ZN(n10922) );
  NOR2_X1 U13439 ( .A1(n10923), .A2(n10922), .ZN(n13458) );
  AOI211_X1 U13440 ( .C1(n10923), .C2(n10922), .A(n13458), .B(n14880), .ZN(
        n10935) );
  OAI21_X1 U13441 ( .B1(P2_REG1_REG_12__SCAN_IN), .B2(n10925), .A(n10924), 
        .ZN(n14871) );
  INV_X1 U13442 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n10926) );
  MUX2_X1 U13443 ( .A(n10926), .B(P2_REG1_REG_13__SCAN_IN), .S(n14875), .Z(
        n14872) );
  NOR2_X1 U13444 ( .A1(n14871), .A2(n14872), .ZN(n14870) );
  XNOR2_X1 U13445 ( .A(n14889), .B(P2_REG1_REG_14__SCAN_IN), .ZN(n14885) );
  NOR2_X1 U13446 ( .A1(n14886), .A2(n14885), .ZN(n14883) );
  NOR2_X1 U13447 ( .A1(n10927), .A2(n14904), .ZN(n10928) );
  XNOR2_X1 U13448 ( .A(n14904), .B(n10927), .ZN(n14896) );
  NOR2_X1 U13449 ( .A1(n14895), .A2(n14896), .ZN(n14894) );
  XNOR2_X1 U13450 ( .A(n13467), .B(P2_REG1_REG_16__SCAN_IN), .ZN(n10929) );
  NOR2_X1 U13451 ( .A1(n10930), .A2(n10929), .ZN(n13466) );
  AOI211_X1 U13452 ( .C1(n10930), .C2(n10929), .A(n13466), .B(n14884), .ZN(
        n10934) );
  NAND2_X1 U13453 ( .A1(P2_REG3_REG_16__SCAN_IN), .A2(P2_U3088), .ZN(n13315)
         );
  NAND2_X1 U13454 ( .A1(n14800), .A2(P2_ADDR_REG_16__SCAN_IN), .ZN(n10931) );
  OAI211_X1 U13455 ( .C1(n14922), .C2(n10932), .A(n13315), .B(n10931), .ZN(
        n10933) );
  OR3_X1 U13456 ( .A1(n10935), .A2(n10934), .A3(n10933), .ZN(P2_U3230) );
  NAND2_X1 U13457 ( .A1(n10936), .A2(n12006), .ZN(n10938) );
  OR2_X1 U13458 ( .A1(n14778), .A2(n14458), .ZN(n10937) );
  NAND2_X1 U13459 ( .A1(n10939), .A2(n11960), .ZN(n10941) );
  AOI22_X1 U13460 ( .A1(n11413), .A2(n6479), .B1(n11430), .B2(
        P2_DATAO_REG_11__SCAN_IN), .ZN(n10940) );
  XNOR2_X1 U13461 ( .A(n14477), .B(n11234), .ZN(n14479) );
  OR2_X1 U13462 ( .A1(n14477), .A2(n13987), .ZN(n10942) );
  NAND2_X1 U13463 ( .A1(n10943), .A2(n11960), .ZN(n10945) );
  AOI22_X1 U13464 ( .A1(n14582), .A2(n6478), .B1(n11430), .B2(
        P2_DATAO_REG_12__SCAN_IN), .ZN(n10944) );
  NAND2_X1 U13465 ( .A1(n11587), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n10952) );
  NAND2_X1 U13466 ( .A1(n11616), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n10951) );
  NAND2_X1 U13467 ( .A1(n10947), .A2(n10946), .ZN(n10948) );
  AND2_X1 U13468 ( .A1(n10963), .A2(n10948), .ZN(n11355) );
  NAND2_X1 U13469 ( .A1(n6475), .A2(n11355), .ZN(n10950) );
  NAND2_X1 U13470 ( .A1(n11526), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n10949) );
  NAND4_X1 U13471 ( .A1(n10952), .A2(n10951), .A3(n10950), .A4(n10949), .ZN(
        n14456) );
  INV_X1 U13472 ( .A(n14456), .ZN(n11346) );
  XNOR2_X1 U13473 ( .A(n11849), .B(n11346), .ZN(n12008) );
  XNOR2_X1 U13474 ( .A(n11013), .B(n12008), .ZN(n14337) );
  INV_X1 U13475 ( .A(n14337), .ZN(n10975) );
  AND2_X1 U13476 ( .A1(n14676), .A2(n10953), .ZN(n14481) );
  INV_X1 U13477 ( .A(n14477), .ZN(n14526) );
  NAND2_X1 U13478 ( .A1(n14481), .A2(n14526), .ZN(n14480) );
  INV_X1 U13479 ( .A(n14480), .ZN(n10954) );
  INV_X1 U13480 ( .A(n11849), .ZN(n14333) );
  OAI211_X1 U13481 ( .C1(n10954), .C2(n14333), .A(n7114), .B(n11049), .ZN(
        n14332) );
  INV_X1 U13482 ( .A(n14332), .ZN(n10973) );
  AOI22_X1 U13483 ( .A1(n14681), .A2(P1_REG2_REG_12__SCAN_IN), .B1(n11355), 
        .B2(n14704), .ZN(n10955) );
  OAI21_X1 U13484 ( .B1(n14333), .B2(n14708), .A(n10955), .ZN(n10972) );
  INV_X1 U13485 ( .A(n14479), .ZN(n10958) );
  OR2_X1 U13486 ( .A1(n14477), .A2(n11234), .ZN(n10959) );
  INV_X1 U13487 ( .A(n12008), .ZN(n10960) );
  NAND2_X1 U13488 ( .A1(n10961), .A2(n10960), .ZN(n10980) );
  OAI211_X1 U13489 ( .C1(n10961), .C2(n10960), .A(n14701), .B(n10980), .ZN(
        n14334) );
  NAND2_X1 U13490 ( .A1(n11616), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n10968) );
  NAND2_X1 U13491 ( .A1(n11526), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n10967) );
  AND2_X1 U13492 ( .A1(n10963), .A2(n10962), .ZN(n10964) );
  NOR2_X1 U13493 ( .A1(n10989), .A2(n10964), .ZN(n11463) );
  NAND2_X1 U13494 ( .A1(n9893), .A2(n11463), .ZN(n10966) );
  NAND2_X1 U13495 ( .A1(n11587), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n10965) );
  NAND4_X1 U13496 ( .A1(n10968), .A2(n10967), .A3(n10966), .A4(n10965), .ZN(
        n13986) );
  NAND2_X1 U13497 ( .A1(n13986), .A2(n14455), .ZN(n10970) );
  NAND2_X1 U13498 ( .A1(n13987), .A2(n14457), .ZN(n10969) );
  AND2_X1 U13499 ( .A1(n10970), .A2(n10969), .ZN(n14331) );
  AOI21_X1 U13500 ( .B1(n14334), .B2(n14331), .A(n14681), .ZN(n10971) );
  AOI211_X1 U13501 ( .C1(n10973), .C2(n14713), .A(n10972), .B(n10971), .ZN(
        n10974) );
  OAI21_X1 U13502 ( .B1(n14174), .B2(n10975), .A(n10974), .ZN(P1_U3281) );
  INV_X1 U13503 ( .A(n11514), .ZN(n10978) );
  OAI222_X1 U13504 ( .A1(n13822), .A2(n10977), .B1(n13820), .B2(n10978), .C1(
        n10976), .C2(P2_U3088), .ZN(P2_U3306) );
  OAI222_X1 U13505 ( .A1(n14292), .A2(n11515), .B1(P1_U3086), .B2(n11979), 
        .C1(n12152), .C2(n10978), .ZN(P1_U3334) );
  OR2_X1 U13506 ( .A1(n11849), .A2(n11346), .ZN(n10979) );
  NAND2_X1 U13507 ( .A1(n10981), .A2(n11960), .ZN(n10985) );
  NOR2_X1 U13508 ( .A1(n9371), .A2(n10982), .ZN(n10983) );
  AOI21_X1 U13509 ( .B1(n11416), .B2(n6479), .A(n10983), .ZN(n10984) );
  NAND2_X1 U13510 ( .A1(n10985), .A2(n10984), .ZN(n11858) );
  INV_X1 U13511 ( .A(n13986), .ZN(n11859) );
  XNOR2_X1 U13512 ( .A(n11858), .B(n11859), .ZN(n12009) );
  OR2_X1 U13513 ( .A1(n11858), .A2(n11859), .ZN(n10995) );
  NAND2_X1 U13514 ( .A1(n10986), .A2(n11960), .ZN(n10988) );
  AOI22_X1 U13515 ( .A1(n14610), .A2(n6478), .B1(n11430), .B2(
        P2_DATAO_REG_14__SCAN_IN), .ZN(n10987) );
  NAND2_X1 U13516 ( .A1(n10989), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n10997) );
  OR2_X1 U13517 ( .A1(n10989), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n10990) );
  NAND2_X1 U13518 ( .A1(n10997), .A2(n10990), .ZN(n14446) );
  INV_X1 U13519 ( .A(n14446), .ZN(n11010) );
  NAND2_X1 U13520 ( .A1(n11010), .A2(n6475), .ZN(n10994) );
  NAND2_X1 U13521 ( .A1(n11616), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n10993) );
  NAND2_X1 U13522 ( .A1(n11526), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n10992) );
  NAND2_X1 U13523 ( .A1(n11587), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n10991) );
  OR2_X1 U13524 ( .A1(n14442), .A2(n13965), .ZN(n11862) );
  NAND2_X1 U13525 ( .A1(n14442), .A2(n13965), .ZN(n11863) );
  NAND2_X1 U13526 ( .A1(n11862), .A2(n11863), .ZN(n12011) );
  NAND3_X1 U13527 ( .A1(n11054), .A2(n12011), .A3(n10995), .ZN(n10996) );
  NAND3_X1 U13528 ( .A1(n11170), .A2(n14701), .A3(n10996), .ZN(n11005) );
  NAND2_X1 U13529 ( .A1(n10997), .A2(n11419), .ZN(n10998) );
  AND2_X1 U13530 ( .A1(n11173), .A2(n10998), .ZN(n13963) );
  AOI22_X1 U13531 ( .A1(n13963), .A2(n6475), .B1(n11587), .B2(
        P1_REG2_REG_15__SCAN_IN), .ZN(n11001) );
  AOI22_X1 U13532 ( .A1(n11616), .A2(P1_REG1_REG_15__SCAN_IN), .B1(n11526), 
        .B2(P1_REG0_REG_15__SCAN_IN), .ZN(n11000) );
  OR2_X1 U13533 ( .A1(n12188), .A2(n14167), .ZN(n11003) );
  NAND2_X1 U13534 ( .A1(n13986), .A2(n14457), .ZN(n11002) );
  NAND2_X1 U13535 ( .A1(n11003), .A2(n11002), .ZN(n14444) );
  INV_X1 U13536 ( .A(n14444), .ZN(n11004) );
  NAND2_X1 U13537 ( .A1(n11005), .A2(n11004), .ZN(n14518) );
  NAND2_X1 U13538 ( .A1(n14442), .A2(n11050), .ZN(n11008) );
  NAND2_X1 U13539 ( .A1(n11008), .A2(n7114), .ZN(n11009) );
  OR2_X1 U13540 ( .A1(n6624), .A2(n11009), .ZN(n14514) );
  AOI22_X1 U13541 ( .A1(n14681), .A2(P1_REG2_REG_14__SCAN_IN), .B1(n11010), 
        .B2(n14704), .ZN(n11012) );
  NAND2_X1 U13542 ( .A1(n14442), .A2(n14476), .ZN(n11011) );
  OAI211_X1 U13543 ( .C1(n14514), .C2(n11701), .A(n11012), .B(n11011), .ZN(
        n11018) );
  OR2_X1 U13544 ( .A1(n11858), .A2(n13986), .ZN(n11014) );
  NAND2_X1 U13545 ( .A1(n11016), .A2(n11015), .ZN(n14512) );
  AND3_X1 U13546 ( .A1(n14513), .A2(n14483), .A3(n14512), .ZN(n11017) );
  AOI211_X1 U13547 ( .C1(n14179), .C2(n14518), .A(n11018), .B(n11017), .ZN(
        n11019) );
  INV_X1 U13548 ( .A(n11019), .ZN(P1_U3279) );
  INV_X1 U13549 ( .A(P3_REG2_REG_11__SCAN_IN), .ZN(n11023) );
  AOI21_X1 U13550 ( .B1(n11023), .B2(n11022), .A(n11140), .ZN(n11038) );
  NAND2_X1 U13551 ( .A1(P3_REG1_REG_11__SCAN_IN), .A2(n11026), .ZN(n11146) );
  OAI21_X1 U13552 ( .B1(n11026), .B2(P3_REG1_REG_11__SCAN_IN), .A(n11146), 
        .ZN(n11036) );
  NAND2_X1 U13553 ( .A1(P3_REG3_REG_11__SCAN_IN), .A2(P3_U3151), .ZN(n12457)
         );
  NAND2_X1 U13554 ( .A1(n15094), .A2(P3_ADDR_REG_11__SCAN_IN), .ZN(n11027) );
  OAI211_X1 U13555 ( .C1(n15088), .C2(n14320), .A(n12457), .B(n11027), .ZN(
        n11035) );
  INV_X1 U13556 ( .A(n11028), .ZN(n11029) );
  NOR2_X1 U13557 ( .A1(n11030), .A2(n11029), .ZN(n11032) );
  MUX2_X1 U13558 ( .A(P3_REG2_REG_11__SCAN_IN), .B(P3_REG1_REG_11__SCAN_IN), 
        .S(n12836), .Z(n11152) );
  XNOR2_X1 U13559 ( .A(n11152), .B(n14320), .ZN(n11031) );
  AOI21_X1 U13560 ( .B1(n11032), .B2(n11031), .A(n11154), .ZN(n11033) );
  NOR2_X1 U13561 ( .A1(n11033), .A2(n15090), .ZN(n11034) );
  AOI211_X1 U13562 ( .C1(n15097), .C2(n11036), .A(n11035), .B(n11034), .ZN(
        n11037) );
  OAI21_X1 U13563 ( .B1(n11038), .B2(n15101), .A(n11037), .ZN(P3_U3193) );
  INV_X1 U13564 ( .A(n11039), .ZN(n11081) );
  OAI211_X1 U13565 ( .C1(n11042), .C2(n11041), .A(n11040), .B(n12502), .ZN(
        n11047) );
  OAI22_X1 U13566 ( .A1(n12443), .A2(n12352), .B1(n12587), .B2(n12474), .ZN(
        n11043) );
  AOI211_X1 U13567 ( .C1(n12476), .C2(n11045), .A(n11044), .B(n11043), .ZN(
        n11046) );
  OAI211_X1 U13568 ( .C1(n11081), .C2(n12452), .A(n11047), .B(n11046), .ZN(
        P3_U3161) );
  XNOR2_X1 U13569 ( .A(n11048), .B(n12009), .ZN(n14523) );
  OAI211_X1 U13570 ( .C1(n11007), .C2(n11006), .A(n7114), .B(n11050), .ZN(
        n14520) );
  AOI22_X1 U13571 ( .A1(n14681), .A2(P1_REG2_REG_13__SCAN_IN), .B1(n11463), 
        .B2(n14704), .ZN(n11052) );
  NAND2_X1 U13572 ( .A1(n11858), .A2(n14476), .ZN(n11051) );
  OAI211_X1 U13573 ( .C1(n14520), .C2(n11701), .A(n11052), .B(n11051), .ZN(
        n11061) );
  INV_X1 U13574 ( .A(n11053), .ZN(n11056) );
  INV_X1 U13575 ( .A(n11054), .ZN(n11055) );
  AOI211_X1 U13576 ( .C1(n12009), .C2(n11056), .A(n14780), .B(n11055), .ZN(
        n14521) );
  INV_X1 U13577 ( .A(n14521), .ZN(n11059) );
  OR2_X1 U13578 ( .A1(n13965), .A2(n14167), .ZN(n11058) );
  NAND2_X1 U13579 ( .A1(n14456), .A2(n14457), .ZN(n11057) );
  AND2_X1 U13580 ( .A1(n11058), .A2(n11057), .ZN(n14519) );
  AOI21_X1 U13581 ( .B1(n11059), .B2(n14519), .A(n14706), .ZN(n11060) );
  AOI211_X1 U13582 ( .C1(n14523), .C2(n14483), .A(n11061), .B(n11060), .ZN(
        n11062) );
  INV_X1 U13583 ( .A(n11062), .ZN(P1_U3280) );
  XNOR2_X1 U13584 ( .A(n11063), .B(n12593), .ZN(n15172) );
  AOI22_X1 U13585 ( .A1(n13098), .A2(n12758), .B1(n13086), .B2(n13100), .ZN(
        n11068) );
  AND2_X1 U13586 ( .A1(n11077), .A2(n11064), .ZN(n11066) );
  OAI211_X1 U13587 ( .C1(n11066), .C2(n12593), .A(n13103), .B(n11065), .ZN(
        n11067) );
  OAI211_X1 U13588 ( .C1(n15172), .C2(n12920), .A(n11068), .B(n11067), .ZN(
        n15174) );
  NAND2_X1 U13589 ( .A1(n15174), .A2(n13106), .ZN(n11072) );
  INV_X1 U13590 ( .A(n12427), .ZN(n11069) );
  OAI22_X1 U13591 ( .A1(n13094), .A2(n15169), .B1(n11069), .B2(n15108), .ZN(
        n11070) );
  AOI21_X1 U13592 ( .B1(P3_REG2_REG_9__SCAN_IN), .B2(n13116), .A(n11070), .ZN(
        n11071) );
  OAI211_X1 U13593 ( .C1(n15172), .C2(n11074), .A(n11072), .B(n11071), .ZN(
        P3_U3224) );
  NAND2_X1 U13594 ( .A1(n13106), .A2(n15120), .ZN(n11073) );
  INV_X1 U13595 ( .A(n13113), .ZN(n13084) );
  OAI21_X1 U13596 ( .B1(n11076), .B2(n12707), .A(n11075), .ZN(n15166) );
  INV_X1 U13597 ( .A(n15166), .ZN(n11085) );
  INV_X1 U13598 ( .A(n11077), .ZN(n11078) );
  AOI21_X1 U13599 ( .B1(n12707), .B2(n11079), .A(n11078), .ZN(n11080) );
  OAI222_X1 U13600 ( .A1(n15111), .A2(n12352), .B1(n15109), .B2(n12587), .C1(
        n15115), .C2(n11080), .ZN(n15164) );
  NAND2_X1 U13601 ( .A1(n15164), .A2(n13106), .ZN(n11084) );
  OAI22_X1 U13602 ( .A1(n13094), .A2(n15163), .B1(n11081), .B2(n15108), .ZN(
        n11082) );
  AOI21_X1 U13603 ( .B1(P3_REG2_REG_8__SCAN_IN), .B2(n13116), .A(n11082), .ZN(
        n11083) );
  OAI211_X1 U13604 ( .C1(n13084), .C2(n11085), .A(n11084), .B(n11083), .ZN(
        P3_U3225) );
  XNOR2_X1 U13605 ( .A(n11281), .B(n6485), .ZN(n11212) );
  AND2_X1 U13606 ( .A1(n13386), .A2(n12163), .ZN(n11086) );
  NAND2_X1 U13607 ( .A1(n11212), .A2(n11086), .ZN(n11214) );
  OAI21_X1 U13608 ( .B1(n11212), .B2(n11086), .A(n11214), .ZN(n11096) );
  NAND2_X1 U13609 ( .A1(n13387), .A2(n12159), .ZN(n11091) );
  INV_X1 U13610 ( .A(n11091), .ZN(n11094) );
  XNOR2_X1 U13611 ( .A(n11730), .B(n6485), .ZN(n11093) );
  INV_X1 U13612 ( .A(n11087), .ZN(n11088) );
  NAND2_X1 U13613 ( .A1(n11090), .A2(n11089), .ZN(n11092) );
  XNOR2_X1 U13614 ( .A(n11093), .B(n11091), .ZN(n11725) );
  AOI211_X1 U13615 ( .C1(n11096), .C2(n11095), .A(n13334), .B(n6625), .ZN(
        n11101) );
  AOI22_X1 U13616 ( .A1(n11753), .A2(n13385), .B1(P2_REG3_REG_13__SCAN_IN), 
        .B2(P2_U3088), .ZN(n11099) );
  INV_X1 U13617 ( .A(n13353), .ZN(n11754) );
  INV_X1 U13618 ( .A(n13352), .ZN(n13368) );
  INV_X1 U13619 ( .A(n11097), .ZN(n11204) );
  AOI22_X1 U13620 ( .A1(n11754), .A2(n13387), .B1(n13368), .B2(n11204), .ZN(
        n11098) );
  OAI211_X1 U13621 ( .C1(n7176), .C2(n13371), .A(n11099), .B(n11098), .ZN(
        n11100) );
  OR2_X1 U13622 ( .A1(n11101), .A2(n11100), .ZN(P2_U3206) );
  INV_X1 U13623 ( .A(n11102), .ZN(n11103) );
  OAI222_X1 U13624 ( .A1(n11105), .A2(P3_U3151), .B1(n13247), .B2(n11104), 
        .C1(n13250), .C2(n11103), .ZN(P3_U3270) );
  NOR2_X1 U13625 ( .A1(n12276), .A2(n11109), .ZN(n11110) );
  AOI21_X1 U13626 ( .B1(n14672), .B2(n10746), .A(n11110), .ZN(n11224) );
  AOI22_X1 U13627 ( .A1(n14672), .A2(n12303), .B1(n10746), .B2(n13988), .ZN(
        n11112) );
  XOR2_X1 U13628 ( .A(n11452), .B(n11112), .Z(n11226) );
  XNOR2_X1 U13629 ( .A(n11227), .B(n11226), .ZN(n11119) );
  NAND2_X1 U13630 ( .A1(n14458), .A2(n14455), .ZN(n11114) );
  NAND2_X1 U13631 ( .A1(n13989), .A2(n14457), .ZN(n11113) );
  NAND2_X1 U13632 ( .A1(n11114), .A2(n11113), .ZN(n14767) );
  AOI22_X1 U13633 ( .A1(n14466), .A2(n14767), .B1(P1_REG3_REG_9__SCAN_IN), 
        .B2(P1_U3086), .ZN(n11116) );
  AND2_X1 U13634 ( .A1(n14672), .A2(n14777), .ZN(n14768) );
  NAND2_X1 U13635 ( .A1(n14768), .A2(n13946), .ZN(n11115) );
  OAI211_X1 U13636 ( .C1(n14469), .C2(n11117), .A(n11116), .B(n11115), .ZN(
        n11118) );
  AOI21_X1 U13637 ( .B1(n11119), .B2(n14465), .A(n11118), .ZN(n11120) );
  INV_X1 U13638 ( .A(n11120), .ZN(P1_U3231) );
  INV_X1 U13639 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n11135) );
  OR2_X1 U13640 ( .A1(n11730), .A2(n13387), .ZN(n11122) );
  XOR2_X1 U13641 ( .A(n11128), .B(n11275), .Z(n11211) );
  NAND2_X1 U13642 ( .A1(n11124), .A2(n13387), .ZN(n11125) );
  XOR2_X1 U13643 ( .A(n11280), .B(n11128), .Z(n11129) );
  AOI222_X1 U13644 ( .A1(n13677), .A2(n11129), .B1(n13385), .B2(n13642), .C1(
        n13387), .C2(n13640), .ZN(n11206) );
  INV_X1 U13645 ( .A(n11130), .ZN(n11132) );
  INV_X1 U13646 ( .A(n11277), .ZN(n11131) );
  AOI21_X1 U13647 ( .B1(n11281), .B2(n11132), .A(n11131), .ZN(n11209) );
  AOI22_X1 U13648 ( .A1(n11209), .A2(n14988), .B1(n11281), .B2(n14986), .ZN(
        n11133) );
  OAI211_X1 U13649 ( .C1(n14984), .C2(n11211), .A(n11206), .B(n11133), .ZN(
        n11136) );
  NAND2_X1 U13650 ( .A1(n11136), .A2(n14953), .ZN(n11134) );
  OAI21_X1 U13651 ( .B1(n15004), .B2(n11135), .A(n11134), .ZN(P2_U3469) );
  NAND2_X1 U13652 ( .A1(n11136), .A2(n15019), .ZN(n11137) );
  OAI21_X1 U13653 ( .B1(n15019), .B2(n10926), .A(n11137), .ZN(P2_U3512) );
  NOR2_X1 U13654 ( .A1(n11139), .A2(n11138), .ZN(n11141) );
  INV_X1 U13655 ( .A(P3_REG2_REG_12__SCAN_IN), .ZN(n11142) );
  AOI22_X1 U13656 ( .A1(P3_REG2_REG_12__SCAN_IN), .A2(n12770), .B1(n12773), 
        .B2(n11142), .ZN(n11143) );
  NOR2_X1 U13657 ( .A1(n11144), .A2(n11143), .ZN(n12767) );
  AOI21_X1 U13658 ( .B1(n11144), .B2(n11143), .A(n12767), .ZN(n11161) );
  INV_X1 U13659 ( .A(P3_REG1_REG_12__SCAN_IN), .ZN(n14426) );
  AOI22_X1 U13660 ( .A1(P3_REG1_REG_12__SCAN_IN), .A2(n12773), .B1(n12770), 
        .B2(n14426), .ZN(n11149) );
  NAND2_X1 U13661 ( .A1(n14320), .A2(n11145), .ZN(n11147) );
  OAI21_X1 U13662 ( .B1(n11149), .B2(n11148), .A(n12769), .ZN(n11159) );
  INV_X1 U13663 ( .A(P3_REG3_REG_12__SCAN_IN), .ZN(n12377) );
  NOR2_X1 U13664 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n12377), .ZN(n11150) );
  AOI21_X1 U13665 ( .B1(n15094), .B2(P3_ADDR_REG_12__SCAN_IN), .A(n11150), 
        .ZN(n11151) );
  OAI21_X1 U13666 ( .B1(n15088), .B2(n12773), .A(n11151), .ZN(n11158) );
  MUX2_X1 U13667 ( .A(P3_REG2_REG_12__SCAN_IN), .B(P3_REG1_REG_12__SCAN_IN), 
        .S(n12836), .Z(n12774) );
  XNOR2_X1 U13668 ( .A(n12774), .B(n12773), .ZN(n11156) );
  NOR2_X1 U13669 ( .A1(n11152), .A2(n14320), .ZN(n11153) );
  OR2_X1 U13670 ( .A1(n11154), .A2(n11153), .ZN(n11155) );
  NOR3_X1 U13671 ( .A1(n11154), .A2(n11153), .A3(n11156), .ZN(n12772) );
  AOI211_X1 U13672 ( .C1(n11156), .C2(n11155), .A(n15090), .B(n12772), .ZN(
        n11157) );
  AOI211_X1 U13673 ( .C1(n11159), .C2(n15097), .A(n11158), .B(n11157), .ZN(
        n11160) );
  OAI21_X1 U13674 ( .B1(n11161), .B2(n15101), .A(n11160), .ZN(P3_U3194) );
  INV_X1 U13675 ( .A(n13965), .ZN(n13985) );
  NAND2_X1 U13676 ( .A1(n14442), .A2(n13985), .ZN(n11162) );
  NAND2_X1 U13677 ( .A1(n11163), .A2(n11960), .ZN(n11166) );
  INV_X1 U13678 ( .A(n14036), .ZN(n11164) );
  AOI22_X1 U13679 ( .A1(n11430), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n6479), 
        .B2(n11164), .ZN(n11165) );
  NAND2_X1 U13680 ( .A1(n12184), .A2(n12188), .ZN(n11866) );
  INV_X1 U13681 ( .A(n12014), .ZN(n11167) );
  OAI21_X1 U13682 ( .B1(n6626), .B2(n11167), .A(n11197), .ZN(n14510) );
  OAI211_X1 U13683 ( .C1(n14506), .C2(n6624), .A(n7114), .B(n11187), .ZN(
        n14505) );
  AOI22_X1 U13684 ( .A1(n14681), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n13963), 
        .B2(n14704), .ZN(n11169) );
  NAND2_X1 U13685 ( .A1(n12184), .A2(n14476), .ZN(n11168) );
  OAI211_X1 U13686 ( .C1(n14505), .C2(n11701), .A(n11169), .B(n11168), .ZN(
        n11178) );
  OAI211_X1 U13687 ( .C1(n11171), .C2(n12014), .A(n14701), .B(n11183), .ZN(
        n14507) );
  AND2_X1 U13688 ( .A1(n11173), .A2(n11172), .ZN(n11174) );
  OR2_X1 U13689 ( .A1(n11174), .A2(n11188), .ZN(n14454) );
  AOI22_X1 U13690 ( .A1(n11587), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n11526), 
        .B2(P1_REG0_REG_16__SCAN_IN), .ZN(n11176) );
  NAND2_X1 U13691 ( .A1(n11616), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n11175) );
  OAI211_X1 U13692 ( .C1(n14454), .C2(n11384), .A(n11176), .B(n11175), .ZN(
        n13983) );
  AOI22_X1 U13693 ( .A1(n13983), .A2(n14455), .B1(n13985), .B2(n14457), .ZN(
        n14504) );
  AOI21_X1 U13694 ( .B1(n14507), .B2(n14504), .A(n14706), .ZN(n11177) );
  AOI211_X1 U13695 ( .C1(n14483), .C2(n14510), .A(n11178), .B(n11177), .ZN(
        n11179) );
  INV_X1 U13696 ( .A(n11179), .ZN(P1_U3278) );
  NAND2_X1 U13697 ( .A1(n11180), .A2(n11960), .ZN(n11182) );
  AOI22_X1 U13698 ( .A1(n11430), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n6478), 
        .B2(n14625), .ZN(n11181) );
  XNOR2_X1 U13699 ( .A(n14498), .B(n13983), .ZN(n12012) );
  NAND2_X1 U13700 ( .A1(n11183), .A2(n11867), .ZN(n11186) );
  INV_X1 U13701 ( .A(n11186), .ZN(n11184) );
  NAND2_X1 U13702 ( .A1(n11184), .A2(n12012), .ZN(n11260) );
  INV_X1 U13703 ( .A(n11260), .ZN(n11185) );
  AOI21_X1 U13704 ( .B1(n11238), .B2(n11186), .A(n11185), .ZN(n14500) );
  AOI211_X1 U13705 ( .C1(n14498), .C2(n11187), .A(n14493), .B(n11243), .ZN(
        n14496) );
  NAND2_X1 U13706 ( .A1(n14681), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n11194) );
  NOR2_X1 U13707 ( .A1(n14188), .A2(n14454), .ZN(n11192) );
  NOR2_X1 U13708 ( .A1(n11188), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n11189) );
  OR2_X1 U13709 ( .A1(n11245), .A2(n11189), .ZN(n13885) );
  AOI22_X1 U13710 ( .A1(n11616), .A2(P1_REG1_REG_17__SCAN_IN), .B1(n11954), 
        .B2(P1_REG0_REG_17__SCAN_IN), .ZN(n11191) );
  NAND2_X1 U13711 ( .A1(n9377), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n11190) );
  OAI211_X1 U13712 ( .C1(n13885), .C2(n11384), .A(n11191), .B(n11190), .ZN(
        n13982) );
  INV_X1 U13713 ( .A(n13982), .ZN(n12201) );
  OAI22_X1 U13714 ( .A1(n12201), .A2(n14167), .B1(n12188), .B2(n14169), .ZN(
        n14497) );
  OAI21_X1 U13715 ( .B1(n11192), .B2(n14497), .A(n14179), .ZN(n11193) );
  OAI211_X1 U13716 ( .C1(n6911), .C2(n14708), .A(n11194), .B(n11193), .ZN(
        n11195) );
  AOI21_X1 U13717 ( .B1(n14496), .B2(n14713), .A(n11195), .ZN(n11199) );
  INV_X1 U13718 ( .A(n12188), .ZN(n13984) );
  OR2_X1 U13719 ( .A1(n12184), .A2(n13984), .ZN(n11196) );
  XNOR2_X1 U13720 ( .A(n11239), .B(n11238), .ZN(n14502) );
  NAND2_X1 U13721 ( .A1(n14502), .A2(n14483), .ZN(n11198) );
  OAI211_X1 U13722 ( .C1(n14500), .C2(n14135), .A(n11199), .B(n11198), .ZN(
        P1_U3277) );
  INV_X1 U13723 ( .A(n11200), .ZN(n11201) );
  OAI222_X1 U13724 ( .A1(n11203), .A2(P3_U3151), .B1(n13247), .B2(n11202), 
        .C1(n13250), .C2(n11201), .ZN(P3_U3269) );
  AOI22_X1 U13725 ( .A1(n13671), .A2(P2_REG2_REG_13__SCAN_IN), .B1(n11204), 
        .B2(n13685), .ZN(n11205) );
  OAI21_X1 U13726 ( .B1(n7176), .B2(n13688), .A(n11205), .ZN(n11208) );
  NOR2_X1 U13727 ( .A1(n11206), .A2(n13671), .ZN(n11207) );
  AOI211_X1 U13728 ( .C1(n11209), .C2(n13669), .A(n11208), .B(n11207), .ZN(
        n11210) );
  OAI21_X1 U13729 ( .B1(n13649), .B2(n11211), .A(n11210), .ZN(P2_U3252) );
  NOR2_X1 U13730 ( .A1(n13327), .A2(n11282), .ZN(n11213) );
  AOI22_X1 U13731 ( .A1(n6625), .A2(n13359), .B1(n11213), .B2(n11212), .ZN(
        n11223) );
  XNOR2_X1 U13732 ( .A(n13784), .B(n12098), .ZN(n11323) );
  NAND2_X1 U13733 ( .A1(n13385), .A2(n12159), .ZN(n11322) );
  XNOR2_X1 U13734 ( .A(n11323), .B(n11322), .ZN(n11215) );
  INV_X1 U13735 ( .A(n11215), .ZN(n11222) );
  INV_X1 U13736 ( .A(n11214), .ZN(n11216) );
  INV_X1 U13737 ( .A(n13784), .ZN(n11289) );
  NOR2_X1 U13738 ( .A1(n11289), .A2(n13371), .ZN(n11220) );
  INV_X1 U13739 ( .A(n11217), .ZN(n11278) );
  AOI22_X1 U13740 ( .A1(n11753), .A2(n13384), .B1(n13368), .B2(n11278), .ZN(
        n11218) );
  NAND2_X1 U13741 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(P2_U3088), .ZN(n14891)
         );
  OAI211_X1 U13742 ( .C1(n11282), .C2(n13353), .A(n11218), .B(n14891), .ZN(
        n11219) );
  AOI211_X1 U13743 ( .C1(n11324), .C2(n13359), .A(n11220), .B(n11219), .ZN(
        n11221) );
  OAI21_X1 U13744 ( .B1(n11223), .B2(n11222), .A(n11221), .ZN(P2_U3187) );
  NAND2_X1 U13745 ( .A1(n14778), .A2(n12303), .ZN(n11229) );
  NAND2_X1 U13746 ( .A1(n10746), .A2(n14458), .ZN(n11228) );
  NAND2_X1 U13747 ( .A1(n11229), .A2(n11228), .ZN(n11230) );
  XNOR2_X1 U13748 ( .A(n11230), .B(n9355), .ZN(n11335) );
  AOI22_X1 U13749 ( .A1(n14778), .A2(n10746), .B1(n12301), .B2(n14458), .ZN(
        n11336) );
  XNOR2_X1 U13750 ( .A(n11335), .B(n11336), .ZN(n11338) );
  XOR2_X1 U13751 ( .A(n11339), .B(n11338), .Z(n11237) );
  NAND2_X1 U13752 ( .A1(n14466), .A2(n14457), .ZN(n13966) );
  INV_X1 U13753 ( .A(n13966), .ZN(n13956) );
  AOI22_X1 U13754 ( .A1(n13956), .A2(n13988), .B1(n13955), .B2(n11231), .ZN(
        n11233) );
  OAI211_X1 U13755 ( .C1(n11234), .C2(n12312), .A(n11233), .B(n11232), .ZN(
        n11235) );
  AOI21_X1 U13756 ( .B1(n14463), .B2(n14778), .A(n11235), .ZN(n11236) );
  OAI21_X1 U13757 ( .B1(n11237), .B2(n13938), .A(n11236), .ZN(P1_U3217) );
  NAND2_X1 U13758 ( .A1(n11240), .A2(n11960), .ZN(n11242) );
  AOI22_X1 U13759 ( .A1(n11430), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n6479), 
        .B2(n14042), .ZN(n11241) );
  XNOR2_X1 U13760 ( .A(n14489), .B(n13982), .ZN(n12015) );
  XNOR2_X1 U13761 ( .A(n11372), .B(n11261), .ZN(n14495) );
  INV_X1 U13762 ( .A(n14495), .ZN(n11265) );
  NOR2_X1 U13763 ( .A1(n11243), .A2(n12203), .ZN(n11244) );
  OR2_X1 U13764 ( .A1(n11387), .A2(n11244), .ZN(n14492) );
  INV_X1 U13765 ( .A(n14492), .ZN(n11258) );
  NOR2_X1 U13766 ( .A1(n11701), .A2(n14493), .ZN(n14191) );
  NOR2_X1 U13767 ( .A1(n11245), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n11246) );
  NOR2_X1 U13768 ( .A1(n11378), .A2(n11246), .ZN(n13932) );
  NAND2_X1 U13769 ( .A1(n13932), .A2(n6475), .ZN(n11251) );
  INV_X1 U13770 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n14649) );
  NAND2_X1 U13771 ( .A1(n11587), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n11248) );
  NAND2_X1 U13772 ( .A1(n11526), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n11247) );
  OAI211_X1 U13773 ( .C1(n10999), .C2(n14649), .A(n11248), .B(n11247), .ZN(
        n11249) );
  INV_X1 U13774 ( .A(n11249), .ZN(n11250) );
  OR2_X1 U13775 ( .A1(n13851), .A2(n14167), .ZN(n11253) );
  NAND2_X1 U13776 ( .A1(n13983), .A2(n14457), .ZN(n11252) );
  NAND2_X1 U13777 ( .A1(n11253), .A2(n11252), .ZN(n14488) );
  INV_X1 U13778 ( .A(n14488), .ZN(n11254) );
  OAI22_X1 U13779 ( .A1(n14681), .A2(n11254), .B1(n13885), .B2(n14188), .ZN(
        n11255) );
  AOI21_X1 U13780 ( .B1(P1_REG2_REG_17__SCAN_IN), .B2(n14706), .A(n11255), 
        .ZN(n11256) );
  OAI21_X1 U13781 ( .B1(n12203), .B2(n14708), .A(n11256), .ZN(n11257) );
  AOI21_X1 U13782 ( .B1(n11258), .B2(n14191), .A(n11257), .ZN(n11264) );
  INV_X1 U13783 ( .A(n13983), .ZN(n12195) );
  NAND2_X1 U13784 ( .A1(n14498), .A2(n12195), .ZN(n11259) );
  NAND2_X1 U13785 ( .A1(n11260), .A2(n11259), .ZN(n11262) );
  NAND2_X1 U13786 ( .A1(n11262), .A2(n11261), .ZN(n14486) );
  INV_X1 U13787 ( .A(n14135), .ZN(n14186) );
  NAND3_X1 U13788 ( .A1(n14487), .A2(n14486), .A3(n14186), .ZN(n11263) );
  OAI211_X1 U13789 ( .C1(n11265), .C2(n14174), .A(n11264), .B(n11263), .ZN(
        P1_U3276) );
  NAND2_X1 U13790 ( .A1(n11532), .A2(n11266), .ZN(n11268) );
  OAI211_X1 U13791 ( .C1(n11269), .C2(n13822), .A(n11268), .B(n11267), .ZN(
        P2_U3304) );
  INV_X1 U13792 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n11533) );
  NAND2_X1 U13793 ( .A1(n11532), .A2(n11270), .ZN(n11271) );
  OAI211_X1 U13794 ( .C1(n11533), .C2(n11652), .A(n11271), .B(n12060), .ZN(
        P1_U3332) );
  INV_X1 U13795 ( .A(n11272), .ZN(n11274) );
  OAI222_X1 U13796 ( .A1(P3_U3151), .A2(n12836), .B1(n13250), .B2(n11274), 
        .C1(n11273), .C2(n13247), .ZN(P3_U3268) );
  XNOR2_X1 U13797 ( .A(n11297), .B(n11283), .ZN(n13788) );
  INV_X1 U13798 ( .A(n11363), .ZN(n11276) );
  AOI21_X1 U13799 ( .B1(n13784), .B2(n11277), .A(n11276), .ZN(n13785) );
  AOI22_X1 U13800 ( .A1(n13671), .A2(P2_REG2_REG_14__SCAN_IN), .B1(n11278), 
        .B2(n13685), .ZN(n11279) );
  OAI21_X1 U13801 ( .B1(n11289), .B2(n13688), .A(n11279), .ZN(n11286) );
  XOR2_X1 U13802 ( .A(n11283), .B(n11288), .Z(n11284) );
  AOI222_X1 U13803 ( .A1(n13677), .A2(n11284), .B1(n13384), .B2(n13642), .C1(
        n13386), .C2(n13640), .ZN(n13787) );
  NOR2_X1 U13804 ( .A1(n13787), .A2(n13671), .ZN(n11285) );
  AOI211_X1 U13805 ( .C1(n13785), .C2(n13669), .A(n11286), .B(n11285), .ZN(
        n11287) );
  OAI21_X1 U13806 ( .B1(n13788), .B2(n13649), .A(n11287), .ZN(P2_U3251) );
  INV_X1 U13807 ( .A(n11299), .ZN(n11361) );
  XNOR2_X1 U13808 ( .A(n11307), .B(n11301), .ZN(n11291) );
  AOI222_X1 U13809 ( .A1(n13645), .A2(n11291), .B1(n13382), .B2(n13642), .C1(
        n13384), .C2(n13640), .ZN(n13778) );
  INV_X1 U13810 ( .A(n11366), .ZN(n11293) );
  INV_X1 U13811 ( .A(n13772), .ZN(n11305) );
  NAND2_X1 U13812 ( .A1(n11305), .A2(n11366), .ZN(n11316) );
  INV_X1 U13813 ( .A(n11316), .ZN(n11292) );
  AOI21_X1 U13814 ( .B1(n13772), .B2(n11293), .A(n11292), .ZN(n13773) );
  NOR2_X1 U13815 ( .A1(n11305), .A2(n13688), .ZN(n11295) );
  OAI22_X1 U13816 ( .A1(n13606), .A2(n10920), .B1(n13317), .B2(n13607), .ZN(
        n11294) );
  AOI211_X1 U13817 ( .C1(n13773), .C2(n13669), .A(n11295), .B(n11294), .ZN(
        n11304) );
  AND2_X1 U13818 ( .A1(n13784), .A2(n13385), .ZN(n11296) );
  OR2_X1 U13819 ( .A1(n13784), .A2(n13385), .ZN(n11298) );
  OR2_X1 U13820 ( .A1(n13780), .A2(n13384), .ZN(n11300) );
  NAND2_X1 U13821 ( .A1(n11302), .A2(n11301), .ZN(n13774) );
  NAND3_X1 U13822 ( .A1(n13775), .A2(n13774), .A3(n13690), .ZN(n11303) );
  OAI211_X1 U13823 ( .C1(n13778), .C2(n13671), .A(n11304), .B(n11303), .ZN(
        P2_U3249) );
  NAND2_X1 U13824 ( .A1(n11305), .A2(n13383), .ZN(n11306) );
  INV_X1 U13825 ( .A(n13383), .ZN(n13328) );
  NAND2_X1 U13826 ( .A1(n11308), .A2(n11311), .ZN(n12113) );
  OAI211_X1 U13827 ( .C1(n11308), .C2(n11311), .A(n12113), .B(n13645), .ZN(
        n11310) );
  AOI22_X1 U13828 ( .A1(n13381), .A2(n13642), .B1(n13640), .B2(n13383), .ZN(
        n11309) );
  AND2_X1 U13829 ( .A1(n11310), .A2(n11309), .ZN(n13770) );
  INV_X1 U13830 ( .A(n11311), .ZN(n11312) );
  NAND2_X1 U13831 ( .A1(n11313), .A2(n11312), .ZN(n12131) );
  OAI21_X1 U13832 ( .B1(n11313), .B2(n11312), .A(n12131), .ZN(n13771) );
  INV_X1 U13833 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n11314) );
  OAI22_X1 U13834 ( .A1(n13606), .A2(n11314), .B1(n13324), .B2(n13607), .ZN(
        n11315) );
  AOI21_X1 U13835 ( .B1(n13767), .B2(n13553), .A(n11315), .ZN(n11319) );
  NAND2_X1 U13836 ( .A1(n11316), .A2(n13767), .ZN(n11317) );
  AND2_X1 U13837 ( .A1(n13674), .A2(n11317), .ZN(n13768) );
  NAND2_X1 U13838 ( .A1(n13768), .A2(n13669), .ZN(n11318) );
  OAI211_X1 U13839 ( .C1(n13771), .C2(n13649), .A(n11319), .B(n11318), .ZN(
        n11320) );
  INV_X1 U13840 ( .A(n11320), .ZN(n11321) );
  OAI21_X1 U13841 ( .B1(n13770), .B2(n13671), .A(n11321), .ZN(P2_U3248) );
  XNOR2_X1 U13842 ( .A(n13780), .B(n12098), .ZN(n11733) );
  INV_X1 U13843 ( .A(n11733), .ZN(n11325) );
  AND2_X1 U13844 ( .A1(n13384), .A2(n12159), .ZN(n11326) );
  INV_X1 U13845 ( .A(n11736), .ZN(n11334) );
  AOI22_X1 U13846 ( .A1(n11327), .A2(n13359), .B1(n13347), .B2(n13384), .ZN(
        n11333) );
  OAI22_X1 U13847 ( .A1(n13351), .A2(n13328), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n11328), .ZN(n11331) );
  OAI22_X1 U13848 ( .A1(n13353), .A2(n11329), .B1(n13352), .B2(n11368), .ZN(
        n11330) );
  AOI211_X1 U13849 ( .C1(n13780), .C2(n9820), .A(n11331), .B(n11330), .ZN(
        n11332) );
  OAI21_X1 U13850 ( .B1(n11334), .B2(n11333), .A(n11332), .ZN(P2_U3213) );
  INV_X1 U13851 ( .A(n11335), .ZN(n11337) );
  AOI22_X1 U13852 ( .A1(n14477), .A2(n10746), .B1(n12301), .B2(n13987), .ZN(
        n11343) );
  NAND2_X1 U13853 ( .A1(n14477), .A2(n12303), .ZN(n11341) );
  NAND2_X1 U13854 ( .A1(n10746), .A2(n13987), .ZN(n11340) );
  NAND2_X1 U13855 ( .A1(n11341), .A2(n11340), .ZN(n11342) );
  XNOR2_X1 U13856 ( .A(n11342), .B(n11452), .ZN(n11345) );
  XOR2_X1 U13857 ( .A(n11343), .B(n11345), .Z(n14461) );
  INV_X1 U13858 ( .A(n11343), .ZN(n11344) );
  NOR2_X1 U13859 ( .A1(n12276), .A2(n11346), .ZN(n11347) );
  AOI21_X1 U13860 ( .B1(n11849), .B2(n10746), .A(n11347), .ZN(n11455) );
  NAND2_X1 U13861 ( .A1(n11849), .A2(n12303), .ZN(n11349) );
  NAND2_X1 U13862 ( .A1(n10746), .A2(n14456), .ZN(n11348) );
  NAND2_X1 U13863 ( .A1(n11349), .A2(n11348), .ZN(n11350) );
  XNOR2_X1 U13864 ( .A(n11350), .B(n11452), .ZN(n11454) );
  XOR2_X1 U13865 ( .A(n11455), .B(n11454), .Z(n11352) );
  AOI21_X1 U13866 ( .B1(n11351), .B2(n11352), .A(n13938), .ZN(n11353) );
  NAND2_X1 U13867 ( .A1(n11353), .A2(n11458), .ZN(n11357) );
  NAND2_X1 U13868 ( .A1(P1_REG3_REG_12__SCAN_IN), .A2(P1_U3086), .ZN(n14584)
         );
  OAI21_X1 U13869 ( .B1(n13934), .B2(n14331), .A(n14584), .ZN(n11354) );
  AOI21_X1 U13870 ( .B1(n11355), .B2(n13955), .A(n11354), .ZN(n11356) );
  OAI211_X1 U13871 ( .C1(n14333), .C2(n13972), .A(n11357), .B(n11356), .ZN(
        P1_U3224) );
  XNOR2_X1 U13872 ( .A(n11358), .B(n11361), .ZN(n13783) );
  OAI21_X1 U13873 ( .B1(n11361), .B2(n11360), .A(n11359), .ZN(n11362) );
  AOI222_X1 U13874 ( .A1(n13677), .A2(n11362), .B1(n13383), .B2(n13642), .C1(
        n13385), .C2(n13640), .ZN(n13782) );
  NAND2_X1 U13875 ( .A1(n13780), .A2(n11363), .ZN(n11364) );
  NAND2_X1 U13876 ( .A1(n11364), .A2(n14988), .ZN(n11365) );
  NOR2_X1 U13877 ( .A1(n11366), .A2(n11365), .ZN(n13779) );
  NAND2_X1 U13878 ( .A1(n13779), .A2(n13680), .ZN(n11367) );
  OAI211_X1 U13879 ( .C1(n13607), .C2(n11368), .A(n13782), .B(n11367), .ZN(
        n11369) );
  NAND2_X1 U13880 ( .A1(n11369), .A2(n13606), .ZN(n11371) );
  AOI22_X1 U13881 ( .A1(n13780), .A2(n13553), .B1(P2_REG2_REG_15__SCAN_IN), 
        .B2(n13671), .ZN(n11370) );
  OAI211_X1 U13882 ( .C1(n13783), .C2(n13649), .A(n11371), .B(n11370), .ZN(
        P2_U3250) );
  NAND2_X1 U13883 ( .A1(n11373), .A2(n11960), .ZN(n11375) );
  AOI22_X1 U13884 ( .A1(n11430), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n6479), 
        .B2(n14657), .ZN(n11374) );
  INV_X1 U13885 ( .A(n13851), .ZN(n13981) );
  XNOR2_X1 U13886 ( .A(n14270), .B(n13981), .ZN(n12018) );
  XOR2_X1 U13887 ( .A(n11427), .B(n12018), .Z(n14272) );
  NAND2_X1 U13888 ( .A1(n12203), .A2(n13982), .ZN(n11376) );
  NAND2_X1 U13889 ( .A1(n14487), .A2(n11376), .ZN(n11377) );
  NAND2_X1 U13890 ( .A1(n11377), .A2(n12018), .ZN(n11434) );
  OAI211_X1 U13891 ( .C1(n11377), .C2(n12018), .A(n11434), .B(n14701), .ZN(
        n11386) );
  NOR2_X1 U13892 ( .A1(n11378), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n11379) );
  OR2_X1 U13893 ( .A1(n11437), .A2(n11379), .ZN(n13850) );
  INV_X1 U13894 ( .A(n6475), .ZN(n11384) );
  INV_X1 U13895 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n14045) );
  NAND2_X1 U13896 ( .A1(n11526), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n11381) );
  NAND2_X1 U13897 ( .A1(n9377), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n11380) );
  OAI211_X1 U13898 ( .C1(n10999), .C2(n14045), .A(n11381), .B(n11380), .ZN(
        n11382) );
  INV_X1 U13899 ( .A(n11382), .ZN(n11383) );
  OAI21_X1 U13900 ( .B1(n13850), .B2(n11384), .A(n11383), .ZN(n13980) );
  AND2_X1 U13901 ( .A1(n13982), .A2(n14457), .ZN(n11385) );
  AOI21_X1 U13902 ( .B1(n13980), .B2(n14455), .A(n11385), .ZN(n13935) );
  NAND2_X1 U13903 ( .A1(n11386), .A2(n13935), .ZN(n14268) );
  INV_X1 U13904 ( .A(n11387), .ZN(n11389) );
  INV_X1 U13905 ( .A(n11435), .ZN(n11388) );
  AOI211_X1 U13906 ( .C1(n14270), .C2(n11389), .A(n14493), .B(n11388), .ZN(
        n14269) );
  NAND2_X1 U13907 ( .A1(n14269), .A2(n14713), .ZN(n11391) );
  AOI22_X1 U13908 ( .A1(n14681), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n13932), 
        .B2(n14704), .ZN(n11390) );
  OAI211_X1 U13909 ( .C1(n12209), .C2(n14708), .A(n11391), .B(n11390), .ZN(
        n11392) );
  AOI21_X1 U13910 ( .B1(n14179), .B2(n14268), .A(n11392), .ZN(n11393) );
  OAI21_X1 U13911 ( .B1(n14174), .B2(n14272), .A(n11393), .ZN(P1_U3275) );
  INV_X1 U13912 ( .A(n11543), .ZN(n12151) );
  INV_X1 U13913 ( .A(n11394), .ZN(n11395) );
  OAI222_X1 U13914 ( .A1(n13822), .A2(n11396), .B1(n13820), .B2(n12151), .C1(
        P2_U3088), .C2(n11395), .ZN(P2_U3303) );
  INV_X1 U13915 ( .A(n11563), .ZN(n11425) );
  OAI222_X1 U13916 ( .A1(P2_U3088), .A2(n11398), .B1(n13820), .B2(n11425), 
        .C1(n11397), .C2(n13822), .ZN(P2_U3301) );
  INV_X1 U13917 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n11399) );
  MUX2_X1 U13918 ( .A(P1_REG2_REG_14__SCAN_IN), .B(n11399), .S(n14610), .Z(
        n14605) );
  NAND2_X1 U13919 ( .A1(P1_REG2_REG_13__SCAN_IN), .A2(n11416), .ZN(n11400) );
  OAI21_X1 U13920 ( .B1(P1_REG2_REG_13__SCAN_IN), .B2(n11416), .A(n11400), 
        .ZN(n14588) );
  INV_X1 U13921 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n11402) );
  AOI22_X1 U13922 ( .A1(n14582), .A2(P1_REG2_REG_12__SCAN_IN), .B1(n11402), 
        .B2(n11401), .ZN(n14580) );
  NAND2_X1 U13923 ( .A1(P1_REG2_REG_11__SCAN_IN), .A2(n11413), .ZN(n11404) );
  OAI21_X1 U13924 ( .B1(n11413), .B2(P1_REG2_REG_11__SCAN_IN), .A(n11404), 
        .ZN(n14567) );
  OAI21_X1 U13925 ( .B1(n14582), .B2(P1_REG2_REG_12__SCAN_IN), .A(n14578), 
        .ZN(n14587) );
  NOR2_X1 U13926 ( .A1(n14588), .A2(n14587), .ZN(n14589) );
  AOI21_X1 U13927 ( .B1(n11416), .B2(P1_REG2_REG_13__SCAN_IN), .A(n14589), 
        .ZN(n11405) );
  INV_X1 U13928 ( .A(n11405), .ZN(n14604) );
  NAND2_X1 U13929 ( .A1(n14605), .A2(n14604), .ZN(n14603) );
  INV_X1 U13930 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n11406) );
  OAI21_X1 U13931 ( .B1(n11407), .B2(n11406), .A(n14028), .ZN(n11423) );
  INV_X1 U13932 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n11408) );
  MUX2_X1 U13933 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n11408), .S(n14610), .Z(
        n14607) );
  OR2_X1 U13934 ( .A1(n14582), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n11414) );
  INV_X1 U13935 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n11409) );
  MUX2_X1 U13936 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n11409), .S(n14582), .Z(
        n14576) );
  INV_X1 U13937 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n11412) );
  MUX2_X1 U13938 ( .A(P1_REG1_REG_11__SCAN_IN), .B(n11412), .S(n11413), .Z(
        n14564) );
  NAND2_X1 U13939 ( .A1(n11414), .A2(n14575), .ZN(n14593) );
  INV_X1 U13940 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n11415) );
  MUX2_X1 U13941 ( .A(n11415), .B(P1_REG1_REG_13__SCAN_IN), .S(n11416), .Z(
        n14594) );
  NOR2_X1 U13942 ( .A1(n14593), .A2(n14594), .ZN(n14592) );
  INV_X1 U13943 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n14511) );
  NAND2_X1 U13944 ( .A1(n11417), .A2(n14511), .ZN(n14037) );
  OAI21_X1 U13945 ( .B1(n11417), .B2(n14511), .A(n14037), .ZN(n11418) );
  NAND2_X1 U13946 ( .A1(n11418), .A2(n14633), .ZN(n11421) );
  NOR2_X1 U13947 ( .A1(n11419), .A2(P1_STATE_REG_SCAN_IN), .ZN(n13968) );
  AOI21_X1 U13948 ( .B1(n14003), .B2(P1_ADDR_REG_15__SCAN_IN), .A(n13968), 
        .ZN(n11420) );
  OAI211_X1 U13949 ( .C1(n14642), .C2(n14036), .A(n11421), .B(n11420), .ZN(
        n11422) );
  AOI21_X1 U13950 ( .B1(n14638), .B2(n11423), .A(n11422), .ZN(n11424) );
  INV_X1 U13951 ( .A(n11424), .ZN(P1_U3258) );
  OAI222_X1 U13952 ( .A1(n14292), .A2(n11564), .B1(P1_U3086), .B2(n9389), .C1(
        n12152), .C2(n11425), .ZN(P1_U3329) );
  NAND2_X1 U13953 ( .A1(n14270), .A2(n13981), .ZN(n11896) );
  INV_X1 U13954 ( .A(n11896), .ZN(n11426) );
  OR2_X1 U13955 ( .A1(n14270), .A2(n13981), .ZN(n11893) );
  OAI21_X2 U13956 ( .B1(n11427), .B2(n11426), .A(n11893), .ZN(n11491) );
  NAND2_X1 U13957 ( .A1(n11428), .A2(n11960), .ZN(n11432) );
  AOI22_X1 U13958 ( .A1(n11430), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n12035), 
        .B2(n6478), .ZN(n11431) );
  XNOR2_X1 U13959 ( .A(n11899), .B(n13980), .ZN(n12020) );
  XNOR2_X1 U13960 ( .A(n11491), .B(n12020), .ZN(n14267) );
  NAND2_X1 U13961 ( .A1(n12209), .A2(n13981), .ZN(n11433) );
  INV_X1 U13962 ( .A(n12020), .ZN(n11490) );
  OAI21_X1 U13963 ( .B1(n6632), .B2(n12020), .A(n11468), .ZN(n14262) );
  AOI21_X1 U13964 ( .B1(n11435), .B2(n11899), .A(n14493), .ZN(n11436) );
  AND2_X1 U13965 ( .A1(n11436), .A2(n11485), .ZN(n14263) );
  NAND2_X1 U13966 ( .A1(n14263), .A2(n14713), .ZN(n11449) );
  OR2_X1 U13967 ( .A1(n11437), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n11438) );
  AND2_X1 U13968 ( .A1(n11438), .A2(n11475), .ZN(n13908) );
  NAND2_X1 U13969 ( .A1(n13908), .A2(n9893), .ZN(n11444) );
  INV_X1 U13970 ( .A(P1_REG2_REG_20__SCAN_IN), .ZN(n11441) );
  NAND2_X1 U13971 ( .A1(n11526), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n11440) );
  NAND2_X1 U13972 ( .A1(n11616), .A2(P1_REG1_REG_20__SCAN_IN), .ZN(n11439) );
  OAI211_X1 U13973 ( .C1(n9420), .C2(n11441), .A(n11440), .B(n11439), .ZN(
        n11442) );
  INV_X1 U13974 ( .A(n11442), .ZN(n11443) );
  OAI22_X1 U13975 ( .A1(n14170), .A2(n14167), .B1(n13851), .B2(n14169), .ZN(
        n14264) );
  NAND2_X1 U13976 ( .A1(n14179), .A2(n14264), .ZN(n11446) );
  NAND2_X1 U13977 ( .A1(n14681), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n11445) );
  OAI211_X1 U13978 ( .C1(n14188), .C2(n13850), .A(n11446), .B(n11445), .ZN(
        n11447) );
  AOI21_X1 U13979 ( .B1(n11899), .B2(n14476), .A(n11447), .ZN(n11448) );
  NAND2_X1 U13980 ( .A1(n11449), .A2(n11448), .ZN(n11450) );
  AOI21_X1 U13981 ( .B1(n14262), .B2(n14186), .A(n11450), .ZN(n11451) );
  OAI21_X1 U13982 ( .B1(n14174), .B2(n14267), .A(n11451), .ZN(P1_U3274) );
  OAI22_X1 U13983 ( .A1(n11006), .A2(n9342), .B1(n11859), .B2(n12223), .ZN(
        n11453) );
  XNOR2_X1 U13984 ( .A(n11453), .B(n11452), .ZN(n12174) );
  OAI22_X1 U13985 ( .A1(n11006), .A2(n12223), .B1(n11859), .B2(n12276), .ZN(
        n12173) );
  XNOR2_X1 U13986 ( .A(n12174), .B(n12173), .ZN(n11462) );
  INV_X1 U13987 ( .A(n11455), .ZN(n11456) );
  NAND2_X1 U13988 ( .A1(n11454), .A2(n11456), .ZN(n11457) );
  INV_X1 U13989 ( .A(n11462), .ZN(n11459) );
  INV_X1 U13990 ( .A(n12176), .ZN(n11460) );
  AOI21_X1 U13991 ( .B1(n11462), .B2(n11461), .A(n11460), .ZN(n11467) );
  AOI22_X1 U13992 ( .A1(n13956), .A2(n14456), .B1(n13955), .B2(n11463), .ZN(
        n11464) );
  NAND2_X1 U13993 ( .A1(P1_REG3_REG_13__SCAN_IN), .A2(P1_U3086), .ZN(n14600)
         );
  OAI211_X1 U13994 ( .C1(n13965), .C2(n12312), .A(n11464), .B(n14600), .ZN(
        n11465) );
  AOI21_X1 U13995 ( .B1(n14463), .B2(n11858), .A(n11465), .ZN(n11466) );
  OAI21_X1 U13996 ( .B1(n11467), .B2(n13938), .A(n11466), .ZN(P1_U3234) );
  INV_X1 U13997 ( .A(n13980), .ZN(n11898) );
  NAND2_X1 U13998 ( .A1(n11899), .A2(n11898), .ZN(n11900) );
  NAND2_X1 U13999 ( .A1(n11469), .A2(n11960), .ZN(n11472) );
  OR2_X1 U14000 ( .A1(n9371), .A2(n11470), .ZN(n11471) );
  XNOR2_X1 U14001 ( .A(n14256), .B(n13978), .ZN(n12019) );
  AOI21_X1 U14002 ( .B1(n11473), .B2(n11493), .A(n14780), .ZN(n11484) );
  NAND2_X1 U14003 ( .A1(n11616), .A2(P1_REG1_REG_21__SCAN_IN), .ZN(n11481) );
  NAND2_X1 U14004 ( .A1(n9377), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n11480) );
  INV_X1 U14005 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n11474) );
  NAND2_X1 U14006 ( .A1(n11474), .A2(n11475), .ZN(n11477) );
  INV_X1 U14007 ( .A(n11522), .ZN(n11523) );
  NAND2_X1 U14008 ( .A1(n9893), .A2(n14160), .ZN(n11479) );
  NAND2_X1 U14009 ( .A1(n11526), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n11478) );
  NAND4_X1 U14010 ( .A1(n11481), .A2(n11480), .A3(n11479), .A4(n11478), .ZN(
        n13977) );
  AND2_X1 U14011 ( .A1(n13977), .A2(n14455), .ZN(n11482) );
  AOI21_X1 U14012 ( .B1(n13980), .B2(n14457), .A(n11482), .ZN(n13904) );
  INV_X1 U14013 ( .A(n13904), .ZN(n11483) );
  AOI21_X1 U14014 ( .B1(n11484), .B2(n11603), .A(n11483), .ZN(n14261) );
  AOI21_X1 U14015 ( .B1(n14256), .B2(n11485), .A(n14493), .ZN(n11486) );
  NAND2_X1 U14016 ( .A1(n11486), .A2(n6622), .ZN(n14258) );
  INV_X1 U14017 ( .A(n14258), .ZN(n11489) );
  AOI22_X1 U14018 ( .A1(n14681), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n13908), 
        .B2(n14704), .ZN(n11487) );
  OAI21_X1 U14019 ( .B1(n13905), .B2(n14708), .A(n11487), .ZN(n11488) );
  AOI21_X1 U14020 ( .B1(n11489), .B2(n14713), .A(n11488), .ZN(n11496) );
  OR2_X1 U14021 ( .A1(n11899), .A2(n13980), .ZN(n11492) );
  NAND2_X1 U14022 ( .A1(n11494), .A2(n12019), .ZN(n14257) );
  NAND3_X1 U14023 ( .A1(n11513), .A2(n14257), .A3(n14483), .ZN(n11495) );
  OAI211_X1 U14024 ( .C1(n14261), .C2(n14706), .A(n11496), .B(n11495), .ZN(
        P1_U3273) );
  XNOR2_X1 U14025 ( .A(n11497), .B(n11498), .ZN(n11504) );
  OR2_X1 U14026 ( .A1(n11499), .A2(n11498), .ZN(n11500) );
  NAND2_X1 U14027 ( .A1(n11501), .A2(n11500), .ZN(n14968) );
  OR2_X1 U14028 ( .A1(n14968), .A2(n13654), .ZN(n11503) );
  AOI22_X1 U14029 ( .A1(n13640), .A2(n13392), .B1(n13390), .B2(n13642), .ZN(
        n11502) );
  OAI211_X1 U14030 ( .C1(n13594), .C2(n11504), .A(n11503), .B(n11502), .ZN(
        n14972) );
  MUX2_X1 U14031 ( .A(n14972), .B(P2_REG2_REG_8__SCAN_IN), .S(n13671), .Z(
        n11511) );
  NOR2_X1 U14032 ( .A1(n11505), .A2(n14970), .ZN(n11506) );
  NOR2_X1 U14033 ( .A1(n11507), .A2(n11506), .ZN(n14969) );
  OAI22_X1 U14034 ( .A1(n13688), .A2(n14970), .B1(n11767), .B2(n13607), .ZN(
        n11508) );
  AOI21_X1 U14035 ( .B1(n14969), .B2(n13669), .A(n11508), .ZN(n11509) );
  OAI21_X1 U14036 ( .B1(n14968), .B2(n13666), .A(n11509), .ZN(n11510) );
  OR2_X1 U14037 ( .A1(n11511), .A2(n11510), .ZN(P2_U3257) );
  OR2_X1 U14038 ( .A1(n13905), .A2(n14170), .ZN(n11512) );
  NAND2_X1 U14039 ( .A1(n11514), .A2(n11960), .ZN(n11517) );
  OR2_X1 U14040 ( .A1(n9371), .A2(n11515), .ZN(n11516) );
  INV_X1 U14041 ( .A(n13977), .ZN(n11604) );
  XNOR2_X1 U14042 ( .A(n14252), .B(n11604), .ZN(n12017) );
  OR2_X1 U14043 ( .A1(n14252), .A2(n13977), .ZN(n11518) );
  NAND2_X1 U14044 ( .A1(n14155), .A2(n11518), .ZN(n14137) );
  NAND2_X1 U14045 ( .A1(n8591), .A2(n11519), .ZN(n11520) );
  XNOR2_X1 U14046 ( .A(n11520), .B(P2_DATAO_REG_22__SCAN_IN), .ZN(n14298) );
  NAND2_X1 U14047 ( .A1(n11587), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n11530) );
  NAND2_X1 U14048 ( .A1(n11616), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n11529) );
  INV_X1 U14049 ( .A(n11536), .ZN(n11525) );
  INV_X1 U14050 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n13916) );
  NAND2_X1 U14051 ( .A1(n11523), .A2(n13916), .ZN(n11524) );
  NAND2_X1 U14052 ( .A1(n6475), .A2(n14148), .ZN(n11528) );
  NAND2_X1 U14053 ( .A1(n11526), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n11527) );
  NAND4_X1 U14054 ( .A1(n11530), .A2(n11529), .A3(n11528), .A4(n11527), .ZN(
        n14120) );
  INV_X1 U14055 ( .A(n14138), .ZN(n14142) );
  OR2_X1 U14056 ( .A1(n14247), .A2(n14120), .ZN(n11531) );
  NAND2_X1 U14057 ( .A1(n11532), .A2(n11960), .ZN(n11535) );
  OR2_X1 U14058 ( .A1(n9371), .A2(n11533), .ZN(n11534) );
  NAND2_X1 U14059 ( .A1(n11616), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n11541) );
  NAND2_X1 U14060 ( .A1(n11954), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n11540) );
  NOR2_X1 U14061 ( .A1(n11536), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n11537) );
  NOR2_X1 U14062 ( .A1(n11546), .A2(n11537), .ZN(n14124) );
  NAND2_X1 U14063 ( .A1(n9893), .A2(n14124), .ZN(n11539) );
  NAND2_X1 U14064 ( .A1(n9377), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n11538) );
  NAND4_X1 U14065 ( .A1(n11541), .A2(n11540), .A3(n11539), .A4(n11538), .ZN(
        n13976) );
  INV_X1 U14066 ( .A(n13976), .ZN(n12251) );
  XNOR2_X1 U14067 ( .A(n14239), .B(n12251), .ZN(n12024) );
  NAND2_X1 U14068 ( .A1(n14239), .A2(n13976), .ZN(n11542) );
  NAND2_X1 U14069 ( .A1(n11543), .A2(n11960), .ZN(n11545) );
  OR2_X1 U14070 ( .A1(n9371), .A2(n12153), .ZN(n11544) );
  NAND2_X2 U14071 ( .A1(n11545), .A2(n11544), .ZN(n14233) );
  NAND2_X1 U14072 ( .A1(n11587), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n11551) );
  NAND2_X1 U14073 ( .A1(n11616), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n11550) );
  INV_X1 U14074 ( .A(n11546), .ZN(n11547) );
  INV_X1 U14075 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n13898) );
  NAND2_X1 U14076 ( .A1(n11546), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n11556) );
  AOI21_X1 U14077 ( .B1(n11547), .B2(n13898), .A(n11555), .ZN(n14109) );
  NAND2_X1 U14078 ( .A1(n6475), .A2(n14109), .ZN(n11549) );
  NAND2_X1 U14079 ( .A1(n11526), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n11548) );
  NAND4_X1 U14080 ( .A1(n11551), .A2(n11550), .A3(n11549), .A4(n11548), .ZN(
        n14121) );
  OR2_X1 U14081 ( .A1(n14233), .A2(n14121), .ZN(n11552) );
  NAND2_X1 U14082 ( .A1(n12317), .A2(n11960), .ZN(n11554) );
  OR2_X1 U14083 ( .A1(n9371), .A2(n12318), .ZN(n11553) );
  NAND2_X1 U14084 ( .A1(n11616), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n11561) );
  NAND2_X1 U14085 ( .A1(n9377), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n11560) );
  INV_X1 U14086 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n11557) );
  NAND2_X1 U14087 ( .A1(n11555), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n11568) );
  INV_X1 U14088 ( .A(n11568), .ZN(n11567) );
  AOI21_X1 U14089 ( .B1(n11557), .B2(n11556), .A(n11567), .ZN(n14091) );
  NAND2_X1 U14090 ( .A1(n6475), .A2(n14091), .ZN(n11559) );
  NAND2_X1 U14091 ( .A1(n11526), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n11558) );
  NAND4_X1 U14092 ( .A1(n11561), .A2(n11560), .A3(n11559), .A4(n11558), .ZN(
        n14068) );
  INV_X1 U14093 ( .A(n14068), .ZN(n12275) );
  INV_X1 U14094 ( .A(n14082), .ZN(n14097) );
  NAND2_X1 U14095 ( .A1(n14226), .A2(n14068), .ZN(n11562) );
  NAND2_X1 U14096 ( .A1(n11563), .A2(n11960), .ZN(n11566) );
  OR2_X1 U14097 ( .A1(n9371), .A2(n11564), .ZN(n11565) );
  NAND2_X1 U14098 ( .A1(n11587), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n11573) );
  NAND2_X1 U14099 ( .A1(n11616), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n11572) );
  INV_X1 U14100 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n11569) );
  NAND2_X1 U14101 ( .A1(n11567), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n11577) );
  INV_X1 U14102 ( .A(n11577), .ZN(n11579) );
  AOI21_X1 U14103 ( .B1(n11569), .B2(n11568), .A(n11579), .ZN(n14073) );
  NAND2_X1 U14104 ( .A1(n6475), .A2(n14073), .ZN(n11571) );
  NAND2_X1 U14105 ( .A1(n11526), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n11570) );
  NAND4_X1 U14106 ( .A1(n11573), .A2(n11572), .A3(n11571), .A4(n11570), .ZN(
        n14085) );
  XNOR2_X1 U14107 ( .A(n14221), .B(n14085), .ZN(n12026) );
  NAND2_X1 U14108 ( .A1(n14221), .A2(n14085), .ZN(n11574) );
  NAND2_X1 U14109 ( .A1(n11664), .A2(n11960), .ZN(n11576) );
  OR2_X1 U14110 ( .A1(n9371), .A2(n11665), .ZN(n11575) );
  NAND2_X1 U14111 ( .A1(n9377), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n11584) );
  NAND2_X1 U14112 ( .A1(n11616), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n11583) );
  INV_X1 U14113 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n11578) );
  NAND2_X1 U14114 ( .A1(n11578), .A2(n11577), .ZN(n11580) );
  NAND2_X1 U14115 ( .A1(P1_REG3_REG_27__SCAN_IN), .A2(n11579), .ZN(n11596) );
  NAND2_X1 U14116 ( .A1(n9893), .A2(n13828), .ZN(n11582) );
  NAND2_X1 U14117 ( .A1(n11526), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n11581) );
  NAND2_X1 U14118 ( .A1(n11655), .A2(n11960), .ZN(n11586) );
  INV_X1 U14119 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n11656) );
  OR2_X1 U14120 ( .A1(n9371), .A2(n11656), .ZN(n11585) );
  NAND2_X1 U14121 ( .A1(n11587), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n11591) );
  NAND2_X1 U14122 ( .A1(n11616), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n11590) );
  XNOR2_X1 U14123 ( .A(n11596), .B(P1_REG3_REG_28__SCAN_IN), .ZN(n11696) );
  NAND2_X1 U14124 ( .A1(n6475), .A2(n11696), .ZN(n11589) );
  NAND2_X1 U14125 ( .A1(n11526), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n11588) );
  NAND4_X1 U14126 ( .A1(n11591), .A2(n11590), .A3(n11589), .A4(n11588), .ZN(
        n13975) );
  NAND2_X1 U14127 ( .A1(n14209), .A2(n13975), .ZN(n11594) );
  OR2_X1 U14128 ( .A1(n14209), .A2(n13975), .ZN(n11592) );
  NAND2_X1 U14129 ( .A1(n11594), .A2(n11592), .ZN(n12029) );
  NAND2_X1 U14130 ( .A1(n11694), .A2(n11594), .ZN(n11601) );
  INV_X1 U14131 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n14293) );
  NOR2_X1 U14132 ( .A1(n9371), .A2(n14293), .ZN(n11595) );
  NAND2_X1 U14133 ( .A1(n9377), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n11600) );
  NAND2_X1 U14134 ( .A1(n11616), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n11599) );
  INV_X1 U14135 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n12308) );
  NOR2_X1 U14136 ( .A1(n11596), .A2(n12308), .ZN(n11620) );
  NAND2_X1 U14137 ( .A1(n6475), .A2(n11620), .ZN(n11598) );
  NAND2_X1 U14138 ( .A1(n11526), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n11597) );
  INV_X1 U14139 ( .A(n12311), .ZN(n13974) );
  XNOR2_X1 U14140 ( .A(n11613), .B(n13974), .ZN(n12031) );
  NAND2_X1 U14141 ( .A1(n13905), .A2(n13978), .ZN(n11602) );
  OR2_X1 U14142 ( .A1(n14252), .A2(n11604), .ZN(n11605) );
  NAND2_X1 U14143 ( .A1(n14247), .A2(n14168), .ZN(n11606) );
  NAND2_X1 U14144 ( .A1(n14239), .A2(n12251), .ZN(n11607) );
  INV_X1 U14145 ( .A(n14103), .ZN(n11608) );
  INV_X1 U14146 ( .A(n14121), .ZN(n12261) );
  OR2_X1 U14147 ( .A1(n14233), .A2(n12261), .ZN(n11609) );
  INV_X1 U14148 ( .A(n14221), .ZN(n14075) );
  INV_X1 U14149 ( .A(n14069), .ZN(n12309) );
  INV_X1 U14150 ( .A(n13975), .ZN(n11611) );
  INV_X1 U14151 ( .A(n14209), .ZN(n11692) );
  INV_X1 U14152 ( .A(n14239), .ZN(n14127) );
  NOR2_X1 U14153 ( .A1(n14247), .A2(n14158), .ZN(n14147) );
  NAND2_X1 U14154 ( .A1(n14127), .A2(n14147), .ZN(n14119) );
  NAND2_X1 U14155 ( .A1(n14206), .A2(n14713), .ZN(n11626) );
  INV_X1 U14156 ( .A(P1_B_REG_SCAN_IN), .ZN(n11614) );
  OR2_X1 U14157 ( .A1(n6484), .A2(n11614), .ZN(n11615) );
  AND2_X1 U14158 ( .A1(n14455), .A2(n11615), .ZN(n14058) );
  INV_X1 U14159 ( .A(P1_REG2_REG_30__SCAN_IN), .ZN(n11619) );
  NAND2_X1 U14160 ( .A1(n11616), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n11618) );
  NAND2_X1 U14161 ( .A1(n11954), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n11617) );
  OAI211_X1 U14162 ( .C1(n9420), .C2(n11619), .A(n11618), .B(n11617), .ZN(
        n13973) );
  NAND2_X1 U14163 ( .A1(n14058), .A2(n13973), .ZN(n14202) );
  INV_X1 U14164 ( .A(n11620), .ZN(n11621) );
  OAI22_X1 U14165 ( .A1(n11622), .A2(n14202), .B1(n14188), .B2(n11621), .ZN(
        n11624) );
  NAND2_X1 U14166 ( .A1(n13975), .A2(n14457), .ZN(n14203) );
  NOR2_X1 U14167 ( .A1(n14681), .A2(n14203), .ZN(n11623) );
  AOI211_X1 U14168 ( .C1(n14706), .C2(P1_REG2_REG_29__SCAN_IN), .A(n11624), 
        .B(n11623), .ZN(n11625) );
  OAI211_X1 U14169 ( .C1(n14204), .C2(n14708), .A(n11626), .B(n11625), .ZN(
        n11627) );
  AOI21_X1 U14170 ( .B1(n14207), .B2(n14186), .A(n11627), .ZN(n11628) );
  OAI21_X1 U14171 ( .B1(n14208), .B2(n14174), .A(n11628), .ZN(P1_U3356) );
  XNOR2_X1 U14172 ( .A(n11631), .B(n12027), .ZN(n11634) );
  AOI22_X1 U14173 ( .A1(n14455), .A2(n13975), .B1(n14085), .B2(n14457), .ZN(
        n11632) );
  AOI211_X1 U14174 ( .C1(n14216), .C2(n14071), .A(n14493), .B(n11693), .ZN(
        n14215) );
  INV_X1 U14175 ( .A(n14216), .ZN(n11638) );
  AOI22_X1 U14176 ( .A1(n14681), .A2(P1_REG2_REG_27__SCAN_IN), .B1(n13828), 
        .B2(n14704), .ZN(n11637) );
  OAI21_X1 U14177 ( .B1(n11638), .B2(n14708), .A(n11637), .ZN(n11640) );
  NOR2_X1 U14178 ( .A1(n14219), .A2(n14175), .ZN(n11639) );
  AOI211_X1 U14179 ( .C1(n14215), .C2(n14713), .A(n11640), .B(n11639), .ZN(
        n11641) );
  OAI21_X1 U14180 ( .B1(n14706), .B2(n14218), .A(n11641), .ZN(P1_U3266) );
  INV_X1 U14181 ( .A(n11642), .ZN(n11643) );
  XNOR2_X1 U14182 ( .A(n12506), .B(P2_DATAO_REG_30__SCAN_IN), .ZN(n11645) );
  XNOR2_X1 U14183 ( .A(n12509), .B(n11645), .ZN(n12521) );
  INV_X1 U14184 ( .A(n12521), .ZN(n11646) );
  OAI222_X1 U14185 ( .A1(P3_U3151), .A2(n11647), .B1(n13247), .B2(n12522), 
        .C1(n13250), .C2(n11646), .ZN(P3_U3265) );
  INV_X1 U14186 ( .A(n11648), .ZN(n11650) );
  OAI222_X1 U14187 ( .A1(n13822), .A2(n11651), .B1(n13820), .B2(n11650), .C1(
        n11649), .C2(P2_U3088), .ZN(P2_U3305) );
  INV_X1 U14188 ( .A(n11961), .ZN(n11704) );
  INV_X1 U14189 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n12507) );
  OAI222_X1 U14190 ( .A1(n14296), .A2(n11704), .B1(P1_U3086), .B2(n9328), .C1(
        n12507), .C2(n11652), .ZN(P1_U3325) );
  OAI222_X1 U14191 ( .A1(n14292), .A2(n11654), .B1(n14296), .B2(n11653), .C1(
        n14149), .C2(P1_U3086), .ZN(P1_U3336) );
  INV_X1 U14192 ( .A(n11655), .ZN(n13815) );
  OAI222_X1 U14193 ( .A1(n14292), .A2(n11656), .B1(n14296), .B2(n13815), .C1(
        n9428), .C2(P1_U3086), .ZN(P1_U3327) );
  INV_X1 U14194 ( .A(n13700), .ZN(n12129) );
  AOI21_X1 U14195 ( .B1(n11657), .B2(P2_B_REG_SCAN_IN), .A(n13657), .ZN(n12122) );
  NAND2_X1 U14196 ( .A1(n12122), .A2(n13372), .ZN(n13697) );
  NOR2_X1 U14197 ( .A1(n13671), .A2(n13697), .ZN(n13499) );
  AOI21_X1 U14198 ( .B1(P2_REG2_REG_31__SCAN_IN), .B2(n13671), .A(n13499), 
        .ZN(n11659) );
  NAND2_X1 U14199 ( .A1(n13694), .A2(n13553), .ZN(n11658) );
  OAI211_X1 U14200 ( .C1(n13695), .C2(n11660), .A(n11659), .B(n11658), .ZN(
        P2_U3234) );
  INV_X1 U14201 ( .A(n11661), .ZN(n14295) );
  OAI222_X1 U14202 ( .A1(n13822), .A2(n11663), .B1(n13820), .B2(n14295), .C1(
        n11662), .C2(P2_U3088), .ZN(P2_U3298) );
  INV_X1 U14203 ( .A(n11664), .ZN(n13816) );
  OAI222_X1 U14204 ( .A1(n14292), .A2(n11665), .B1(n14296), .B2(n13816), .C1(
        n6484), .C2(P1_U3086), .ZN(P1_U3328) );
  INV_X1 U14205 ( .A(n11666), .ZN(n11669) );
  OAI222_X1 U14206 ( .A1(n13247), .A2(n11670), .B1(n13250), .B2(n11669), .C1(
        P3_U3151), .C2(n11667), .ZN(P3_U3266) );
  XNOR2_X1 U14207 ( .A(n12542), .B(n11671), .ZN(n11679) );
  INV_X1 U14208 ( .A(n11679), .ZN(n11672) );
  NAND2_X1 U14209 ( .A1(n11672), .A2(n12502), .ZN(n11685) );
  INV_X1 U14210 ( .A(n11673), .ZN(n11674) );
  NAND4_X1 U14211 ( .A1(n11684), .A2(n12502), .A3(n11674), .A4(n11679), .ZN(
        n11683) );
  AOI22_X1 U14212 ( .A1(n12441), .A2(n12746), .B1(P3_REG3_REG_28__SCAN_IN), 
        .B2(P3_U3151), .ZN(n11676) );
  NAND2_X1 U14213 ( .A1(n12497), .A2(n12875), .ZN(n11675) );
  OAI211_X1 U14214 ( .C1(n11677), .C2(n12443), .A(n11676), .B(n11675), .ZN(
        n11681) );
  NOR4_X1 U14215 ( .A1(n11679), .A2(n11678), .A3(n12478), .A4(n12746), .ZN(
        n11680) );
  AOI211_X1 U14216 ( .C1(n12476), .C2(n7954), .A(n11681), .B(n11680), .ZN(
        n11682) );
  OAI211_X1 U14217 ( .C1(n11685), .C2(n11684), .A(n11683), .B(n11682), .ZN(
        P3_U3160) );
  XNOR2_X1 U14218 ( .A(n11686), .B(n11593), .ZN(n11690) );
  NAND2_X1 U14219 ( .A1(n13974), .A2(n14455), .ZN(n11688) );
  NAND2_X1 U14220 ( .A1(n14069), .A2(n14457), .ZN(n11687) );
  OAI211_X1 U14221 ( .C1(n11693), .C2(n11692), .A(n7114), .B(n11691), .ZN(
        n14211) );
  NAND2_X1 U14222 ( .A1(n11695), .A2(n12029), .ZN(n14210) );
  NAND3_X1 U14223 ( .A1(n11694), .A2(n14483), .A3(n14210), .ZN(n11700) );
  INV_X1 U14224 ( .A(n11696), .ZN(n12310) );
  NAND2_X1 U14225 ( .A1(n14681), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n11697) );
  OAI21_X1 U14226 ( .B1(n14188), .B2(n12310), .A(n11697), .ZN(n11698) );
  AOI21_X1 U14227 ( .B1(n14209), .B2(n14476), .A(n11698), .ZN(n11699) );
  OAI211_X1 U14228 ( .C1(n11701), .C2(n14211), .A(n11700), .B(n11699), .ZN(
        n11702) );
  INV_X1 U14229 ( .A(n11702), .ZN(n11703) );
  OAI21_X1 U14230 ( .B1(n14214), .B2(n14706), .A(n11703), .ZN(P1_U3265) );
  OAI222_X1 U14231 ( .A1(n11705), .A2(P2_U3088), .B1(n13820), .B2(n11704), 
        .C1(n12506), .C2(n13822), .ZN(P2_U3297) );
  AOI22_X1 U14232 ( .A1(n13347), .A2(n8833), .B1(n13359), .B2(n11706), .ZN(
        n11708) );
  NOR2_X1 U14233 ( .A1(n11708), .A2(n11707), .ZN(n11715) );
  OAI22_X1 U14234 ( .A1(n11710), .A2(n13353), .B1(n13351), .B2(n11709), .ZN(
        n11714) );
  NAND2_X1 U14235 ( .A1(n9820), .A2(n14947), .ZN(n11711) );
  NAND2_X1 U14236 ( .A1(P2_REG3_REG_5__SCAN_IN), .A2(P2_U3088), .ZN(n14823) );
  OAI211_X1 U14237 ( .C1(n13352), .C2(n11712), .A(n11711), .B(n14823), .ZN(
        n11713) );
  AOI211_X1 U14238 ( .C1(n11716), .C2(n11715), .A(n11714), .B(n11713), .ZN(
        n11717) );
  OAI21_X1 U14239 ( .B1(n11718), .B2(n13334), .A(n11717), .ZN(P2_U3199) );
  INV_X1 U14240 ( .A(n11719), .ZN(n11720) );
  AOI22_X1 U14241 ( .A1(n11753), .A2(n13386), .B1(n13368), .B2(n11720), .ZN(
        n11722) );
  OAI211_X1 U14242 ( .C1(n11723), .C2(n13353), .A(n11722), .B(n11721), .ZN(
        n11729) );
  AOI22_X1 U14243 ( .A1(n11724), .A2(n13359), .B1(n13347), .B2(n13388), .ZN(
        n11726) );
  NOR3_X1 U14244 ( .A1(n11727), .A2(n11726), .A3(n11725), .ZN(n11728) );
  AOI211_X1 U14245 ( .C1(n11730), .C2(n9820), .A(n11729), .B(n11728), .ZN(
        n11731) );
  OAI21_X1 U14246 ( .B1(n11732), .B2(n13334), .A(n11731), .ZN(P2_U3196) );
  INV_X1 U14247 ( .A(n13313), .ZN(n11738) );
  NAND2_X1 U14248 ( .A1(n13383), .A2(n12163), .ZN(n11740) );
  XNOR2_X1 U14249 ( .A(n13772), .B(n6485), .ZN(n11739) );
  XOR2_X1 U14250 ( .A(n11740), .B(n11739), .Z(n13314) );
  INV_X1 U14251 ( .A(n13314), .ZN(n11737) );
  INV_X1 U14252 ( .A(n11739), .ZN(n13329) );
  NAND2_X1 U14253 ( .A1(n13382), .A2(n12159), .ZN(n11741) );
  XNOR2_X1 U14254 ( .A(n13767), .B(n6485), .ZN(n11743) );
  XOR2_X1 U14255 ( .A(n11741), .B(n11743), .Z(n13331) );
  INV_X1 U14256 ( .A(n11741), .ZN(n11742) );
  XNOR2_X1 U14257 ( .A(n13763), .B(n12098), .ZN(n13281) );
  NAND2_X1 U14258 ( .A1(n13381), .A2(n12159), .ZN(n11744) );
  NOR2_X1 U14259 ( .A1(n13281), .A2(n11744), .ZN(n11745) );
  AOI21_X1 U14260 ( .B1(n13281), .B2(n11744), .A(n11745), .ZN(n13360) );
  NAND2_X1 U14261 ( .A1(n13641), .A2(n12159), .ZN(n11746) );
  XNOR2_X1 U14262 ( .A(n13757), .B(n6485), .ZN(n11750) );
  XOR2_X1 U14263 ( .A(n11746), .B(n11750), .Z(n13283) );
  INV_X1 U14264 ( .A(n11746), .ZN(n11747) );
  XNOR2_X1 U14265 ( .A(n13752), .B(n6485), .ZN(n12062) );
  NAND2_X1 U14266 ( .A1(n13624), .A2(n12159), .ZN(n12063) );
  XNOR2_X1 U14267 ( .A(n12062), .B(n12063), .ZN(n11752) );
  AOI22_X1 U14268 ( .A1(n11750), .A2(n13359), .B1(n13347), .B2(n13641), .ZN(
        n11751) );
  NOR2_X1 U14269 ( .A1(n11752), .A2(n11751), .ZN(n11758) );
  INV_X1 U14270 ( .A(n13752), .ZN(n13634) );
  AOI22_X1 U14271 ( .A1(n11753), .A2(n13643), .B1(P2_REG3_REG_20__SCAN_IN), 
        .B2(P2_U3088), .ZN(n11756) );
  AOI22_X1 U14272 ( .A1(n11754), .A2(n13641), .B1(n13368), .B2(n13632), .ZN(
        n11755) );
  OAI211_X1 U14273 ( .C1(n13634), .C2(n13371), .A(n11756), .B(n11755), .ZN(
        n11757) );
  AOI21_X1 U14274 ( .B1(n13277), .B2(n11758), .A(n11757), .ZN(n11759) );
  OAI21_X1 U14275 ( .B1(n12066), .B2(n13334), .A(n11759), .ZN(P2_U3205) );
  NAND3_X1 U14276 ( .A1(n13347), .A2(n13392), .A3(n11760), .ZN(n11761) );
  OAI21_X1 U14277 ( .B1(n11762), .B2(n13334), .A(n11761), .ZN(n11765) );
  INV_X1 U14278 ( .A(n11763), .ZN(n11764) );
  NAND2_X1 U14279 ( .A1(n11765), .A2(n11764), .ZN(n11773) );
  NAND2_X1 U14280 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(P2_U3088), .ZN(n14835) );
  OAI21_X1 U14281 ( .B1(n13353), .B2(n11766), .A(n14835), .ZN(n11770) );
  OAI22_X1 U14282 ( .A1(n13351), .A2(n11768), .B1(n13352), .B2(n11767), .ZN(
        n11769) );
  AOI211_X1 U14283 ( .C1(n11771), .C2(n9820), .A(n11770), .B(n11769), .ZN(
        n11772) );
  OAI211_X1 U14284 ( .C1(n11774), .C2(n13334), .A(n11773), .B(n11772), .ZN(
        P2_U3193) );
  NAND2_X1 U14285 ( .A1(n11779), .A2(n11776), .ZN(n14185) );
  NAND2_X1 U14286 ( .A1(n11778), .A2(n11777), .ZN(n11963) );
  XNOR2_X1 U14287 ( .A(n11779), .B(n11797), .ZN(n11780) );
  OAI211_X1 U14288 ( .C1(n14185), .C2(n11781), .A(n11780), .B(n11998), .ZN(
        n11785) );
  NAND2_X1 U14289 ( .A1(n11792), .A2(n6473), .ZN(n11783) );
  NAND2_X1 U14290 ( .A1(n11797), .A2(n6906), .ZN(n11782) );
  MUX2_X1 U14291 ( .A(n11783), .B(n11782), .S(n14187), .Z(n11784) );
  NAND2_X1 U14292 ( .A1(n11789), .A2(n11788), .ZN(n11796) );
  INV_X1 U14293 ( .A(n11791), .ZN(n11793) );
  MUX2_X1 U14294 ( .A(n7233), .B(n11793), .S(n11792), .Z(n11794) );
  INV_X1 U14295 ( .A(n11794), .ZN(n11795) );
  NAND2_X1 U14296 ( .A1(n11796), .A2(n11795), .ZN(n11801) );
  MUX2_X1 U14297 ( .A(n11798), .B(n13993), .S(n11792), .Z(n11802) );
  NAND2_X1 U14298 ( .A1(n11801), .A2(n11802), .ZN(n11800) );
  MUX2_X1 U14299 ( .A(n13993), .B(n11798), .S(n11792), .Z(n11799) );
  NAND2_X1 U14300 ( .A1(n11800), .A2(n11799), .ZN(n11806) );
  INV_X1 U14301 ( .A(n11801), .ZN(n11804) );
  INV_X1 U14302 ( .A(n11802), .ZN(n11803) );
  NAND2_X1 U14303 ( .A1(n11804), .A2(n11803), .ZN(n11805) );
  NAND2_X1 U14304 ( .A1(n11806), .A2(n11805), .ZN(n11811) );
  MUX2_X1 U14305 ( .A(n13992), .B(n11807), .S(n6476), .Z(n11810) );
  NAND2_X1 U14306 ( .A1(n11811), .A2(n11810), .ZN(n11809) );
  MUX2_X1 U14307 ( .A(n11807), .B(n13992), .S(n11792), .Z(n11808) );
  NAND2_X1 U14308 ( .A1(n11809), .A2(n11808), .ZN(n11813) );
  OR2_X2 U14309 ( .A1(n11811), .A2(n11810), .ZN(n11812) );
  MUX2_X1 U14310 ( .A(n13991), .B(n13945), .S(n6483), .Z(n11815) );
  MUX2_X1 U14311 ( .A(n13991), .B(n13945), .S(n6476), .Z(n11814) );
  INV_X1 U14312 ( .A(n11815), .ZN(n11816) );
  MUX2_X1 U14313 ( .A(n13990), .B(n11817), .S(n11980), .Z(n11821) );
  NAND2_X1 U14314 ( .A1(n11820), .A2(n11821), .ZN(n11819) );
  MUX2_X1 U14315 ( .A(n13990), .B(n11817), .S(n6483), .Z(n11818) );
  NAND2_X1 U14316 ( .A1(n11819), .A2(n11818), .ZN(n11825) );
  INV_X1 U14317 ( .A(n11820), .ZN(n11823) );
  INV_X1 U14318 ( .A(n11821), .ZN(n11822) );
  NAND2_X1 U14319 ( .A1(n11823), .A2(n11822), .ZN(n11824) );
  MUX2_X1 U14320 ( .A(n13989), .B(n11826), .S(n6483), .Z(n11830) );
  NAND2_X1 U14321 ( .A1(n11829), .A2(n11830), .ZN(n11828) );
  MUX2_X1 U14322 ( .A(n13989), .B(n11826), .S(n11980), .Z(n11827) );
  NAND2_X1 U14323 ( .A1(n11828), .A2(n11827), .ZN(n11834) );
  INV_X1 U14324 ( .A(n11829), .ZN(n11832) );
  INV_X1 U14325 ( .A(n11830), .ZN(n11831) );
  NAND2_X1 U14326 ( .A1(n11832), .A2(n11831), .ZN(n11833) );
  MUX2_X1 U14327 ( .A(n13988), .B(n14672), .S(n11980), .Z(n11836) );
  MUX2_X1 U14328 ( .A(n13988), .B(n14672), .S(n6483), .Z(n11835) );
  INV_X1 U14329 ( .A(n11836), .ZN(n11837) );
  MUX2_X1 U14330 ( .A(n14458), .B(n14778), .S(n6483), .Z(n11841) );
  NAND2_X1 U14331 ( .A1(n11840), .A2(n11841), .ZN(n11839) );
  MUX2_X1 U14332 ( .A(n14458), .B(n14778), .S(n11980), .Z(n11838) );
  NAND2_X1 U14333 ( .A1(n11839), .A2(n11838), .ZN(n11845) );
  INV_X1 U14334 ( .A(n11840), .ZN(n11843) );
  INV_X1 U14335 ( .A(n11841), .ZN(n11842) );
  NAND2_X1 U14336 ( .A1(n11843), .A2(n11842), .ZN(n11844) );
  MUX2_X1 U14337 ( .A(n13987), .B(n14477), .S(n11980), .Z(n11847) );
  MUX2_X1 U14338 ( .A(n13987), .B(n14477), .S(n6483), .Z(n11846) );
  INV_X1 U14339 ( .A(n11847), .ZN(n11848) );
  MUX2_X1 U14340 ( .A(n14456), .B(n11849), .S(n6483), .Z(n11853) );
  NAND2_X1 U14341 ( .A1(n11852), .A2(n11853), .ZN(n11851) );
  MUX2_X1 U14342 ( .A(n14456), .B(n11849), .S(n11980), .Z(n11850) );
  NAND2_X1 U14343 ( .A1(n11851), .A2(n11850), .ZN(n11857) );
  INV_X1 U14344 ( .A(n11852), .ZN(n11855) );
  INV_X1 U14345 ( .A(n11853), .ZN(n11854) );
  NAND2_X1 U14346 ( .A1(n11855), .A2(n11854), .ZN(n11856) );
  MUX2_X1 U14347 ( .A(n13986), .B(n11858), .S(n11980), .Z(n11861) );
  MUX2_X1 U14348 ( .A(n11859), .B(n11006), .S(n6483), .Z(n11860) );
  NAND2_X1 U14349 ( .A1(n11867), .A2(n11862), .ZN(n11865) );
  NAND2_X1 U14350 ( .A1(n11866), .A2(n11863), .ZN(n11864) );
  MUX2_X1 U14351 ( .A(n11865), .B(n11864), .S(n11980), .Z(n11869) );
  MUX2_X1 U14352 ( .A(n11867), .B(n11866), .S(n6483), .Z(n11868) );
  MUX2_X1 U14353 ( .A(n13983), .B(n14498), .S(n6483), .Z(n11885) );
  OR2_X1 U14354 ( .A1(n13983), .A2(n11980), .ZN(n11871) );
  INV_X1 U14355 ( .A(n11871), .ZN(n11881) );
  AOI21_X1 U14356 ( .B1(n11885), .B2(n13982), .A(n11881), .ZN(n11874) );
  NAND2_X1 U14357 ( .A1(n11885), .A2(n12201), .ZN(n11870) );
  OR2_X1 U14358 ( .A1(n14498), .A2(n6483), .ZN(n11877) );
  NAND2_X1 U14359 ( .A1(n11870), .A2(n11877), .ZN(n11872) );
  NAND2_X1 U14360 ( .A1(n13982), .A2(n11980), .ZN(n11878) );
  OAI22_X1 U14361 ( .A1(n14498), .A2(n11878), .B1(n13982), .B2(n11871), .ZN(
        n11884) );
  AOI21_X1 U14362 ( .B1(n11872), .B2(n12203), .A(n11884), .ZN(n11873) );
  OAI21_X1 U14363 ( .B1(n12203), .B2(n11874), .A(n11873), .ZN(n11875) );
  NAND2_X1 U14364 ( .A1(n11876), .A2(n11875), .ZN(n11891) );
  INV_X1 U14365 ( .A(n11877), .ZN(n11880) );
  INV_X1 U14366 ( .A(n11878), .ZN(n11879) );
  AOI21_X1 U14367 ( .B1(n11885), .B2(n11880), .A(n11879), .ZN(n11888) );
  NAND2_X1 U14368 ( .A1(n11885), .A2(n11881), .ZN(n11882) );
  OAI21_X1 U14369 ( .B1(n11980), .B2(n13982), .A(n11882), .ZN(n11883) );
  NAND2_X1 U14370 ( .A1(n11883), .A2(n14489), .ZN(n11887) );
  NAND2_X1 U14371 ( .A1(n11885), .A2(n11884), .ZN(n11886) );
  OAI211_X1 U14372 ( .C1(n11888), .C2(n14489), .A(n11887), .B(n11886), .ZN(
        n11889) );
  INV_X1 U14373 ( .A(n11889), .ZN(n11890) );
  NAND2_X1 U14374 ( .A1(n11891), .A2(n11890), .ZN(n11894) );
  INV_X1 U14375 ( .A(n11894), .ZN(n11897) );
  MUX2_X1 U14376 ( .A(n13851), .B(n12209), .S(n11980), .Z(n11892) );
  OAI211_X1 U14377 ( .C1(n11897), .C2(n11896), .A(n11895), .B(n12020), .ZN(
        n11903) );
  OR2_X1 U14378 ( .A1(n11899), .A2(n11898), .ZN(n11901) );
  MUX2_X1 U14379 ( .A(n11901), .B(n11900), .S(n11980), .Z(n11902) );
  NAND2_X1 U14380 ( .A1(n11903), .A2(n11902), .ZN(n11906) );
  MUX2_X1 U14381 ( .A(n14170), .B(n13905), .S(n6483), .Z(n11905) );
  MUX2_X1 U14382 ( .A(n13978), .B(n14256), .S(n11980), .Z(n11904) );
  NAND2_X1 U14383 ( .A1(n11906), .A2(n11905), .ZN(n11907) );
  MUX2_X1 U14384 ( .A(n13977), .B(n14252), .S(n11980), .Z(n11910) );
  MUX2_X1 U14385 ( .A(n14252), .B(n13977), .S(n11980), .Z(n11909) );
  MUX2_X1 U14386 ( .A(n14120), .B(n14247), .S(n6483), .Z(n11914) );
  NAND2_X1 U14387 ( .A1(n11913), .A2(n11914), .ZN(n11912) );
  MUX2_X1 U14388 ( .A(n14120), .B(n14247), .S(n11980), .Z(n11911) );
  NAND2_X1 U14389 ( .A1(n11912), .A2(n11911), .ZN(n11918) );
  INV_X1 U14390 ( .A(n11913), .ZN(n11916) );
  INV_X1 U14391 ( .A(n11914), .ZN(n11915) );
  NAND2_X1 U14392 ( .A1(n11916), .A2(n11915), .ZN(n11917) );
  NAND2_X1 U14393 ( .A1(n11918), .A2(n11917), .ZN(n11921) );
  MUX2_X1 U14394 ( .A(n13976), .B(n14239), .S(n11980), .Z(n11922) );
  NAND2_X1 U14395 ( .A1(n11921), .A2(n11922), .ZN(n11920) );
  MUX2_X1 U14396 ( .A(n13976), .B(n14239), .S(n6483), .Z(n11919) );
  NAND2_X1 U14397 ( .A1(n11920), .A2(n11919), .ZN(n11926) );
  INV_X1 U14398 ( .A(n11921), .ZN(n11924) );
  INV_X1 U14399 ( .A(n11922), .ZN(n11923) );
  NAND2_X1 U14400 ( .A1(n11924), .A2(n11923), .ZN(n11925) );
  MUX2_X1 U14401 ( .A(n14121), .B(n14233), .S(n6483), .Z(n11928) );
  INV_X1 U14402 ( .A(n11928), .ZN(n11929) );
  MUX2_X1 U14403 ( .A(n14068), .B(n14226), .S(n11980), .Z(n11933) );
  NAND2_X1 U14404 ( .A1(n11932), .A2(n11933), .ZN(n11931) );
  MUX2_X1 U14405 ( .A(n14068), .B(n14226), .S(n6483), .Z(n11930) );
  NAND2_X1 U14406 ( .A1(n11931), .A2(n11930), .ZN(n11937) );
  INV_X1 U14407 ( .A(n11932), .ZN(n11935) );
  INV_X1 U14408 ( .A(n11933), .ZN(n11934) );
  NAND2_X1 U14409 ( .A1(n11935), .A2(n11934), .ZN(n11936) );
  MUX2_X1 U14410 ( .A(n14085), .B(n14221), .S(n6483), .Z(n11939) );
  MUX2_X1 U14411 ( .A(n14085), .B(n14221), .S(n11980), .Z(n11938) );
  MUX2_X1 U14412 ( .A(n14069), .B(n14216), .S(n11980), .Z(n11943) );
  NAND2_X1 U14413 ( .A1(n11942), .A2(n11943), .ZN(n11941) );
  MUX2_X1 U14414 ( .A(n14069), .B(n14216), .S(n6483), .Z(n11940) );
  NAND2_X1 U14415 ( .A1(n11941), .A2(n11940), .ZN(n11947) );
  INV_X1 U14416 ( .A(n11942), .ZN(n11945) );
  INV_X1 U14417 ( .A(n11943), .ZN(n11944) );
  NAND2_X1 U14418 ( .A1(n11945), .A2(n11944), .ZN(n11946) );
  MUX2_X1 U14419 ( .A(n13975), .B(n14209), .S(n6483), .Z(n11949) );
  MUX2_X1 U14420 ( .A(n13975), .B(n14209), .S(n11980), .Z(n11948) );
  MUX2_X1 U14421 ( .A(n12311), .B(n14204), .S(n11980), .Z(n11950) );
  MUX2_X1 U14422 ( .A(n12311), .B(n14204), .S(n6483), .Z(n11952) );
  OAI22_X1 U14423 ( .A1(n11953), .A2(n11952), .B1(n11951), .B2(n6676), .ZN(
        n11987) );
  NAND2_X1 U14424 ( .A1(n11616), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n11957) );
  NAND2_X1 U14425 ( .A1(n9377), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n11956) );
  NAND2_X1 U14426 ( .A1(n11954), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n11955) );
  AND3_X1 U14427 ( .A1(n11957), .A2(n11956), .A3(n11955), .ZN(n11989) );
  INV_X1 U14428 ( .A(n11989), .ZN(n14059) );
  OAI21_X1 U14429 ( .B1(n14059), .B2(n11958), .A(n13973), .ZN(n11962) );
  NOR2_X1 U14430 ( .A1(n9371), .A2(n12507), .ZN(n11959) );
  MUX2_X1 U14431 ( .A(n11962), .B(n14201), .S(n11980), .Z(n11984) );
  INV_X1 U14432 ( .A(n14201), .ZN(n14062) );
  NAND2_X1 U14433 ( .A1(n14062), .A2(n6483), .ZN(n11968) );
  INV_X1 U14434 ( .A(n11963), .ZN(n11964) );
  OAI22_X1 U14435 ( .A1(n6483), .A2(n11989), .B1(n11965), .B2(n11964), .ZN(
        n11966) );
  NAND2_X1 U14436 ( .A1(n11966), .A2(n13973), .ZN(n11967) );
  NAND2_X1 U14437 ( .A1(n11968), .A2(n11967), .ZN(n11983) );
  AND2_X1 U14438 ( .A1(n11984), .A2(n11983), .ZN(n12040) );
  NAND2_X1 U14439 ( .A1(n13807), .A2(n11960), .ZN(n11971) );
  INV_X1 U14440 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n11969) );
  OR2_X1 U14441 ( .A1(n9371), .A2(n11969), .ZN(n11970) );
  NAND2_X1 U14442 ( .A1(n12045), .A2(n11980), .ZN(n11990) );
  NAND2_X1 U14443 ( .A1(n11973), .A2(n11972), .ZN(n11974) );
  NAND2_X1 U14444 ( .A1(n11975), .A2(n11974), .ZN(n11977) );
  NAND2_X1 U14445 ( .A1(n11977), .A2(n11976), .ZN(n12043) );
  NAND2_X1 U14446 ( .A1(n11979), .A2(n11978), .ZN(n12046) );
  AND2_X1 U14447 ( .A1(n12043), .A2(n12046), .ZN(n11988) );
  OR2_X1 U14448 ( .A1(n12045), .A2(n11980), .ZN(n12044) );
  OR2_X1 U14449 ( .A1(n12044), .A2(n11989), .ZN(n11981) );
  OAI211_X1 U14450 ( .C1(n11990), .C2(n14059), .A(n11988), .B(n11981), .ZN(
        n11994) );
  NOR3_X1 U14451 ( .A1(n11987), .A2(n12040), .A3(n11994), .ZN(n12054) );
  XNOR2_X1 U14452 ( .A(n12045), .B(n14059), .ZN(n12034) );
  INV_X1 U14453 ( .A(n12043), .ZN(n11982) );
  AND2_X1 U14454 ( .A1(n12034), .A2(n11982), .ZN(n12039) );
  INV_X1 U14455 ( .A(n11983), .ZN(n11986) );
  INV_X1 U14456 ( .A(n11984), .ZN(n11985) );
  NAND2_X1 U14457 ( .A1(n11986), .A2(n11985), .ZN(n11993) );
  OR3_X1 U14458 ( .A1(n11990), .A2(n14059), .A3(n12043), .ZN(n11992) );
  NAND4_X1 U14459 ( .A1(n11990), .A2(n11989), .A3(n11988), .A4(n12045), .ZN(
        n11991) );
  OAI211_X1 U14460 ( .C1(n11994), .C2(n11993), .A(n11992), .B(n11991), .ZN(
        n11995) );
  INV_X1 U14461 ( .A(n11995), .ZN(n12051) );
  INV_X1 U14462 ( .A(n14185), .ZN(n14720) );
  NAND4_X1 U14463 ( .A1(n14720), .A2(n11998), .A3(n11997), .A4(n11996), .ZN(
        n12000) );
  NOR3_X1 U14464 ( .A1(n12000), .A2(n14700), .A3(n11999), .ZN(n12003) );
  NAND4_X1 U14465 ( .A1(n12004), .A2(n12003), .A3(n12002), .A4(n12001), .ZN(
        n12005) );
  OR4_X1 U14466 ( .A1(n14479), .A2(n12006), .A3(n14664), .A4(n12005), .ZN(
        n12007) );
  OR3_X1 U14467 ( .A1(n12009), .A2(n12008), .A3(n12007), .ZN(n12010) );
  NOR2_X1 U14468 ( .A1(n12011), .A2(n12010), .ZN(n12013) );
  NAND4_X1 U14469 ( .A1(n12015), .A2(n12014), .A3(n12013), .A4(n12012), .ZN(
        n12016) );
  NOR2_X1 U14470 ( .A1(n12017), .A2(n12016), .ZN(n12022) );
  AND2_X1 U14471 ( .A1(n12019), .A2(n12018), .ZN(n12021) );
  NAND4_X1 U14472 ( .A1(n14138), .A2(n12022), .A3(n12021), .A4(n12020), .ZN(
        n12023) );
  NOR2_X1 U14473 ( .A1(n12024), .A2(n12023), .ZN(n12025) );
  AND2_X1 U14474 ( .A1(n12026), .A2(n12025), .ZN(n12028) );
  NAND4_X1 U14475 ( .A1(n12029), .A2(n12028), .A3(n14102), .A4(n12027), .ZN(
        n12030) );
  NOR2_X1 U14476 ( .A1(n12030), .A2(n14082), .ZN(n12033) );
  XNOR2_X1 U14477 ( .A(n14062), .B(n13973), .ZN(n12032) );
  NAND4_X1 U14478 ( .A1(n12034), .A2(n12033), .A3(n12032), .A4(n12031), .ZN(
        n12036) );
  XNOR2_X1 U14479 ( .A(n12036), .B(n12035), .ZN(n12038) );
  INV_X1 U14480 ( .A(n12046), .ZN(n12037) );
  NAND2_X1 U14481 ( .A1(n12038), .A2(n12037), .ZN(n12050) );
  INV_X1 U14482 ( .A(n12039), .ZN(n12042) );
  INV_X1 U14483 ( .A(n12040), .ZN(n12041) );
  OR2_X1 U14484 ( .A1(n12042), .A2(n12041), .ZN(n12049) );
  XNOR2_X1 U14485 ( .A(n12044), .B(n12043), .ZN(n12047) );
  NAND4_X1 U14486 ( .A1(n12047), .A2(n14197), .A3(n14059), .A4(n12046), .ZN(
        n12048) );
  NAND4_X1 U14487 ( .A1(n12051), .A2(n12050), .A3(n12049), .A4(n12048), .ZN(
        n12052) );
  NOR3_X1 U14488 ( .A1(n12054), .A2(n12053), .A3(n12052), .ZN(n12061) );
  NAND4_X1 U14489 ( .A1(n12057), .A2(n12056), .A3(n14457), .A4(n12055), .ZN(
        n12058) );
  OAI211_X1 U14490 ( .C1(n14297), .C2(n12060), .A(n12058), .B(P1_B_REG_SCAN_IN), .ZN(n12059) );
  OAI21_X1 U14491 ( .B1(n12061), .B2(n12060), .A(n12059), .ZN(P1_U3242) );
  INV_X1 U14492 ( .A(n12062), .ZN(n12064) );
  NAND2_X1 U14493 ( .A1(n12064), .A2(n12063), .ZN(n12065) );
  XNOR2_X1 U14494 ( .A(n13747), .B(n6485), .ZN(n12068) );
  NAND2_X1 U14495 ( .A1(n13643), .A2(n12159), .ZN(n12069) );
  XNOR2_X1 U14496 ( .A(n12068), .B(n12069), .ZN(n13290) );
  INV_X1 U14497 ( .A(n12069), .ZN(n12067) );
  NAND2_X1 U14498 ( .A1(n12068), .A2(n12067), .ZN(n12077) );
  XNOR2_X1 U14499 ( .A(n13740), .B(n6485), .ZN(n12074) );
  NAND2_X1 U14500 ( .A1(n13346), .A2(n12074), .ZN(n12082) );
  INV_X1 U14501 ( .A(n12068), .ZN(n12070) );
  AND2_X1 U14502 ( .A1(n12070), .A2(n12069), .ZN(n12072) );
  INV_X1 U14503 ( .A(n12072), .ZN(n12071) );
  NAND2_X1 U14504 ( .A1(n12074), .A2(n12071), .ZN(n12080) );
  INV_X1 U14505 ( .A(n12074), .ZN(n13345) );
  NAND2_X1 U14506 ( .A1(n13345), .A2(n12072), .ZN(n12076) );
  INV_X1 U14507 ( .A(n12077), .ZN(n12073) );
  NAND2_X1 U14508 ( .A1(n12074), .A2(n12073), .ZN(n12075) );
  AND4_X1 U14509 ( .A1(n12076), .A2(n12075), .A3(n13625), .A4(n12159), .ZN(
        n12079) );
  NAND3_X1 U14510 ( .A1(n12081), .A2(n13345), .A3(n12077), .ZN(n12078) );
  OAI211_X1 U14511 ( .C1(n12081), .C2(n12080), .A(n12079), .B(n12078), .ZN(
        n13349) );
  XNOR2_X1 U14512 ( .A(n13735), .B(n12098), .ZN(n12086) );
  NOR2_X1 U14513 ( .A1(n13598), .A2(n12083), .ZN(n13260) );
  XNOR2_X1 U14514 ( .A(n13729), .B(n12098), .ZN(n13301) );
  NAND2_X1 U14515 ( .A1(n13379), .A2(n12159), .ZN(n12084) );
  NOR2_X1 U14516 ( .A1(n13301), .A2(n12084), .ZN(n12090) );
  AOI21_X1 U14517 ( .B1(n13301), .B2(n12084), .A(n12090), .ZN(n13339) );
  AND2_X1 U14518 ( .A1(n13260), .A2(n13339), .ZN(n12085) );
  INV_X1 U14519 ( .A(n12086), .ZN(n12087) );
  NAND2_X1 U14520 ( .A1(n12088), .A2(n12087), .ZN(n13335) );
  INV_X1 U14521 ( .A(n13339), .ZN(n12089) );
  INV_X1 U14522 ( .A(n12090), .ZN(n12091) );
  NAND3_X1 U14523 ( .A1(n13298), .A2(n13297), .A3(n12091), .ZN(n12096) );
  XNOR2_X1 U14524 ( .A(n13724), .B(n6485), .ZN(n12092) );
  AND2_X1 U14525 ( .A1(n13378), .A2(n12159), .ZN(n12093) );
  NAND2_X1 U14526 ( .A1(n12092), .A2(n12093), .ZN(n12097) );
  INV_X1 U14527 ( .A(n12092), .ZN(n12102) );
  INV_X1 U14528 ( .A(n12093), .ZN(n12094) );
  NAND2_X1 U14529 ( .A1(n12102), .A2(n12094), .ZN(n12095) );
  INV_X1 U14530 ( .A(n12097), .ZN(n12099) );
  XNOR2_X1 U14531 ( .A(n13719), .B(n12098), .ZN(n12154) );
  NAND2_X1 U14532 ( .A1(n13377), .A2(n12163), .ZN(n12155) );
  XNOR2_X1 U14533 ( .A(n12154), .B(n12155), .ZN(n12103) );
  NOR2_X1 U14534 ( .A1(n12099), .A2(n12103), .ZN(n12100) );
  NOR2_X1 U14535 ( .A1(n12101), .A2(n13334), .ZN(n12105) );
  NOR3_X1 U14536 ( .A1(n12102), .A2(n7152), .A3(n13327), .ZN(n12104) );
  OAI21_X1 U14537 ( .B1(n12105), .B2(n12104), .A(n12103), .ZN(n12111) );
  OAI22_X1 U14538 ( .A1(n12143), .A2(n13657), .B1(n7152), .B2(n13655), .ZN(
        n13532) );
  INV_X1 U14539 ( .A(n13532), .ZN(n12108) );
  INV_X1 U14540 ( .A(n12106), .ZN(n13535) );
  AOI22_X1 U14541 ( .A1(n13535), .A2(n13368), .B1(P2_REG3_REG_26__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12107) );
  OAI21_X1 U14542 ( .B1(n12108), .B2(n13366), .A(n12107), .ZN(n12109) );
  AOI21_X1 U14543 ( .B1(n13719), .B2(n9820), .A(n12109), .ZN(n12110) );
  OAI211_X1 U14544 ( .C1(n13334), .C2(n12158), .A(n12111), .B(n12110), .ZN(
        P2_U3212) );
  INV_X1 U14545 ( .A(n13719), .ZN(n13537) );
  INV_X1 U14546 ( .A(n13740), .ZN(n13604) );
  INV_X1 U14547 ( .A(n13624), .ZN(n13658) );
  NAND2_X1 U14548 ( .A1(n12113), .A2(n12112), .ZN(n13675) );
  NAND2_X1 U14549 ( .A1(n13763), .A2(n13656), .ZN(n12114) );
  INV_X1 U14550 ( .A(n13612), .ZN(n13596) );
  AOI21_X1 U14551 ( .B1(n13604), .B2(n13625), .A(n13593), .ZN(n13579) );
  INV_X1 U14552 ( .A(n13583), .ZN(n13578) );
  NAND2_X1 U14553 ( .A1(n13579), .A2(n13578), .ZN(n13577) );
  INV_X1 U14554 ( .A(n13735), .ZN(n13590) );
  NAND2_X1 U14555 ( .A1(n13577), .A2(n7358), .ZN(n13566) );
  INV_X1 U14556 ( .A(n13565), .ZN(n13561) );
  INV_X1 U14557 ( .A(n12118), .ZN(n13538) );
  INV_X1 U14558 ( .A(n13502), .ZN(n13505) );
  NAND2_X1 U14559 ( .A1(n13504), .A2(n12119), .ZN(n12121) );
  INV_X1 U14560 ( .A(n12144), .ZN(n12120) );
  XNOR2_X1 U14561 ( .A(n12121), .B(n12120), .ZN(n12125) );
  AOI22_X1 U14562 ( .A1(n13375), .A2(n13640), .B1(n12122), .B2(n13373), .ZN(
        n12123) );
  AOI21_X2 U14563 ( .B1(n12125), .B2(n13645), .A(n12124), .ZN(n13704) );
  XNOR2_X1 U14564 ( .A(n13509), .B(n13700), .ZN(n13701) );
  INV_X1 U14565 ( .A(n12126), .ZN(n12127) );
  AOI22_X1 U14566 ( .A1(n12127), .A2(n13685), .B1(P2_REG2_REG_29__SCAN_IN), 
        .B2(n13671), .ZN(n12128) );
  OAI21_X1 U14567 ( .B1(n12129), .B2(n13688), .A(n12128), .ZN(n12147) );
  NAND2_X1 U14568 ( .A1(n13767), .A2(n13382), .ZN(n12130) );
  NAND2_X1 U14569 ( .A1(n12131), .A2(n12130), .ZN(n13683) );
  OR2_X1 U14570 ( .A1(n13763), .A2(n13381), .ZN(n12134) );
  NOR2_X1 U14571 ( .A1(n13757), .A2(n13641), .ZN(n12136) );
  NAND2_X1 U14572 ( .A1(n13757), .A2(n13641), .ZN(n12135) );
  OR2_X1 U14573 ( .A1(n13752), .A2(n13624), .ZN(n12137) );
  INV_X1 U14574 ( .A(n13616), .ZN(n13622) );
  OR2_X1 U14575 ( .A1(n13747), .A2(n13643), .ZN(n12138) );
  NAND2_X1 U14576 ( .A1(n12139), .A2(n12138), .ZN(n13613) );
  NOR2_X1 U14577 ( .A1(n13613), .A2(n13612), .ZN(n13611) );
  NAND2_X1 U14578 ( .A1(n13584), .A2(n13583), .ZN(n13582) );
  OR2_X1 U14579 ( .A1(n13735), .A2(n13380), .ZN(n12140) );
  NAND2_X1 U14580 ( .A1(n13582), .A2(n12140), .ZN(n13562) );
  NOR2_X1 U14581 ( .A1(n13562), .A2(n13561), .ZN(n13564) );
  AOI22_X1 U14582 ( .A1(n13503), .A2(n13502), .B1(n13706), .B2(n13375), .ZN(
        n12145) );
  XNOR2_X1 U14583 ( .A(n12145), .B(n12144), .ZN(n13703) );
  NOR2_X1 U14584 ( .A1(n13703), .A2(n13649), .ZN(n12146) );
  OAI21_X1 U14585 ( .B1(n13704), .B2(n13671), .A(n12148), .ZN(P2_U3236) );
  OAI222_X1 U14586 ( .A1(n14292), .A2(n12153), .B1(n12152), .B2(n12151), .C1(
        n12150), .C2(P1_U3086), .ZN(P1_U3331) );
  INV_X1 U14587 ( .A(n12154), .ZN(n12157) );
  INV_X1 U14588 ( .A(n12155), .ZN(n12156) );
  XNOR2_X1 U14589 ( .A(n13711), .B(n6485), .ZN(n12161) );
  AND2_X1 U14590 ( .A1(n13376), .A2(n12159), .ZN(n12160) );
  NAND2_X1 U14591 ( .A1(n12161), .A2(n12160), .ZN(n12162) );
  OAI21_X1 U14592 ( .B1(n12161), .B2(n12160), .A(n12162), .ZN(n13252) );
  NAND2_X1 U14593 ( .A1(n13257), .A2(n12162), .ZN(n12167) );
  NAND2_X1 U14594 ( .A1(n13375), .A2(n12163), .ZN(n12164) );
  XNOR2_X1 U14595 ( .A(n12164), .B(n6485), .ZN(n12165) );
  XNOR2_X1 U14596 ( .A(n13706), .B(n12165), .ZN(n12166) );
  XNOR2_X1 U14597 ( .A(n12167), .B(n12166), .ZN(n12172) );
  AOI22_X1 U14598 ( .A1(n13374), .A2(n13642), .B1(n13376), .B2(n13640), .ZN(
        n13507) );
  NOR2_X1 U14599 ( .A1(n13507), .A2(n13366), .ZN(n12170) );
  OAI22_X1 U14600 ( .A1(n13511), .A2(n13352), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n12168), .ZN(n12169) );
  AOI211_X1 U14601 ( .C1(n13706), .C2(n9820), .A(n12170), .B(n12169), .ZN(
        n12171) );
  OAI21_X1 U14602 ( .B1(n12172), .B2(n13334), .A(n12171), .ZN(P2_U3192) );
  OR2_X1 U14603 ( .A1(n12174), .A2(n12173), .ZN(n12175) );
  INV_X1 U14604 ( .A(n14442), .ZN(n14515) );
  OAI22_X1 U14605 ( .A1(n14515), .A2(n12223), .B1(n13965), .B2(n12276), .ZN(
        n12180) );
  NAND2_X1 U14606 ( .A1(n14442), .A2(n12303), .ZN(n12178) );
  NAND2_X1 U14607 ( .A1(n10746), .A2(n13985), .ZN(n12177) );
  NAND2_X1 U14608 ( .A1(n12178), .A2(n12177), .ZN(n12179) );
  XNOR2_X1 U14609 ( .A(n12179), .B(n9355), .ZN(n12181) );
  XOR2_X1 U14610 ( .A(n12180), .B(n12181), .Z(n14440) );
  NAND2_X1 U14611 ( .A1(n14441), .A2(n14440), .ZN(n12183) );
  NAND2_X1 U14612 ( .A1(n12184), .A2(n12303), .ZN(n12186) );
  NAND2_X1 U14613 ( .A1(n10746), .A2(n13984), .ZN(n12185) );
  NAND2_X1 U14614 ( .A1(n12186), .A2(n12185), .ZN(n12187) );
  XNOR2_X1 U14615 ( .A(n12187), .B(n9355), .ZN(n12190) );
  OAI22_X1 U14616 ( .A1(n14506), .A2(n12223), .B1(n12188), .B2(n12276), .ZN(
        n13961) );
  INV_X1 U14617 ( .A(n12189), .ZN(n12191) );
  NAND2_X1 U14618 ( .A1(n12191), .A2(n12190), .ZN(n14447) );
  NAND2_X1 U14619 ( .A1(n14498), .A2(n12303), .ZN(n12193) );
  NAND2_X1 U14620 ( .A1(n10746), .A2(n13983), .ZN(n12192) );
  NAND2_X1 U14621 ( .A1(n12193), .A2(n12192), .ZN(n12194) );
  XNOR2_X1 U14622 ( .A(n12194), .B(n9355), .ZN(n12197) );
  NOR2_X1 U14623 ( .A1(n12276), .A2(n12195), .ZN(n12196) );
  AOI21_X1 U14624 ( .B1(n14498), .B2(n10746), .A(n12196), .ZN(n12198) );
  XNOR2_X1 U14625 ( .A(n12197), .B(n12198), .ZN(n14450) );
  INV_X1 U14626 ( .A(n12197), .ZN(n12199) );
  NAND2_X1 U14627 ( .A1(n12199), .A2(n12198), .ZN(n12200) );
  OAI22_X1 U14628 ( .A1(n12203), .A2(n9342), .B1(n12201), .B2(n12223), .ZN(
        n12202) );
  XNOR2_X1 U14629 ( .A(n12202), .B(n9355), .ZN(n13880) );
  OR2_X1 U14630 ( .A1(n12203), .A2(n12223), .ZN(n12205) );
  NAND2_X1 U14631 ( .A1(n12301), .A2(n13982), .ZN(n12204) );
  NAND2_X1 U14632 ( .A1(n12205), .A2(n12204), .ZN(n13881) );
  NAND2_X1 U14633 ( .A1(n13880), .A2(n13881), .ZN(n12207) );
  OAI22_X1 U14634 ( .A1(n12209), .A2(n9342), .B1(n13851), .B2(n12223), .ZN(
        n12208) );
  XNOR2_X1 U14635 ( .A(n12208), .B(n9355), .ZN(n12219) );
  OAI22_X1 U14636 ( .A1(n12209), .A2(n12223), .B1(n13851), .B2(n12276), .ZN(
        n12218) );
  XNOR2_X1 U14637 ( .A(n12219), .B(n12218), .ZN(n13931) );
  NAND2_X1 U14638 ( .A1(n11899), .A2(n12303), .ZN(n12211) );
  NAND2_X1 U14639 ( .A1(n13980), .A2(n10746), .ZN(n12210) );
  NAND2_X1 U14640 ( .A1(n12211), .A2(n12210), .ZN(n12212) );
  XNOR2_X1 U14641 ( .A(n12212), .B(n12273), .ZN(n12217) );
  INV_X1 U14642 ( .A(n12217), .ZN(n12215) );
  AND2_X1 U14643 ( .A1(n13980), .A2(n12301), .ZN(n12213) );
  AOI21_X1 U14644 ( .B1(n11899), .B2(n10746), .A(n12213), .ZN(n12216) );
  INV_X1 U14645 ( .A(n12216), .ZN(n12214) );
  OR2_X1 U14646 ( .A1(n13931), .A2(n7350), .ZN(n12220) );
  XNOR2_X1 U14647 ( .A(n12217), .B(n12216), .ZN(n13844) );
  NOR2_X1 U14648 ( .A1(n12219), .A2(n12218), .ZN(n13845) );
  NOR2_X1 U14649 ( .A1(n13844), .A2(n13845), .ZN(n13846) );
  OR2_X1 U14650 ( .A1(n13905), .A2(n12223), .ZN(n12222) );
  NAND2_X1 U14651 ( .A1(n13978), .A2(n12301), .ZN(n12221) );
  NAND2_X1 U14652 ( .A1(n12222), .A2(n12221), .ZN(n12225) );
  OAI22_X1 U14653 ( .A1(n13905), .A2(n9342), .B1(n14170), .B2(n12223), .ZN(
        n12224) );
  XNOR2_X1 U14654 ( .A(n12224), .B(n9355), .ZN(n12226) );
  XOR2_X1 U14655 ( .A(n12225), .B(n12226), .Z(n13902) );
  NAND2_X1 U14656 ( .A1(n12226), .A2(n12225), .ZN(n12227) );
  NAND2_X1 U14657 ( .A1(n14252), .A2(n12303), .ZN(n12229) );
  NAND2_X1 U14658 ( .A1(n10746), .A2(n13977), .ZN(n12228) );
  NAND2_X1 U14659 ( .A1(n12229), .A2(n12228), .ZN(n12230) );
  XNOR2_X1 U14660 ( .A(n12230), .B(n9355), .ZN(n12234) );
  NAND2_X1 U14661 ( .A1(n14252), .A2(n10746), .ZN(n12232) );
  NAND2_X1 U14662 ( .A1(n12301), .A2(n13977), .ZN(n12231) );
  NAND2_X1 U14663 ( .A1(n12232), .A2(n12231), .ZN(n12233) );
  NOR2_X1 U14664 ( .A1(n12234), .A2(n12233), .ZN(n13913) );
  AOI21_X1 U14665 ( .B1(n12234), .B2(n12233), .A(n13913), .ZN(n13863) );
  NAND2_X1 U14666 ( .A1(n14247), .A2(n12303), .ZN(n12236) );
  NAND2_X1 U14667 ( .A1(n10746), .A2(n14120), .ZN(n12235) );
  NAND2_X1 U14668 ( .A1(n12236), .A2(n12235), .ZN(n12237) );
  XNOR2_X1 U14669 ( .A(n12237), .B(n12273), .ZN(n12239) );
  NOR2_X1 U14670 ( .A1(n12276), .A2(n14168), .ZN(n12238) );
  AOI21_X1 U14671 ( .B1(n14247), .B2(n10746), .A(n12238), .ZN(n12240) );
  NAND2_X1 U14672 ( .A1(n12239), .A2(n12240), .ZN(n13835) );
  INV_X1 U14673 ( .A(n12239), .ZN(n12242) );
  INV_X1 U14674 ( .A(n12240), .ZN(n12241) );
  NAND2_X1 U14675 ( .A1(n12242), .A2(n12241), .ZN(n12243) );
  AND2_X1 U14676 ( .A1(n13863), .A2(n13912), .ZN(n12244) );
  INV_X1 U14677 ( .A(n13912), .ZN(n12246) );
  INV_X1 U14678 ( .A(n13913), .ZN(n12245) );
  AND2_X1 U14679 ( .A1(n13833), .A2(n13835), .ZN(n12247) );
  NAND2_X1 U14680 ( .A1(n14239), .A2(n12303), .ZN(n12249) );
  NAND2_X1 U14681 ( .A1(n10746), .A2(n13976), .ZN(n12248) );
  NAND2_X1 U14682 ( .A1(n12249), .A2(n12248), .ZN(n12250) );
  XNOR2_X1 U14683 ( .A(n12250), .B(n12273), .ZN(n12253) );
  NOR2_X1 U14684 ( .A1(n12276), .A2(n12251), .ZN(n12252) );
  AOI21_X1 U14685 ( .B1(n14239), .B2(n10746), .A(n12252), .ZN(n12254) );
  NAND2_X1 U14686 ( .A1(n12253), .A2(n12254), .ZN(n13889) );
  INV_X1 U14687 ( .A(n12253), .ZN(n12256) );
  INV_X1 U14688 ( .A(n12254), .ZN(n12255) );
  NAND2_X1 U14689 ( .A1(n12256), .A2(n12255), .ZN(n12257) );
  NAND2_X1 U14690 ( .A1(n14233), .A2(n12303), .ZN(n12259) );
  NAND2_X1 U14691 ( .A1(n10746), .A2(n14121), .ZN(n12258) );
  NAND2_X1 U14692 ( .A1(n12259), .A2(n12258), .ZN(n12260) );
  XNOR2_X1 U14693 ( .A(n12260), .B(n12273), .ZN(n12263) );
  NOR2_X1 U14694 ( .A1(n12276), .A2(n12261), .ZN(n12262) );
  AOI21_X1 U14695 ( .B1(n14233), .B2(n10746), .A(n12262), .ZN(n12264) );
  NAND2_X1 U14696 ( .A1(n12263), .A2(n12264), .ZN(n13873) );
  INV_X1 U14697 ( .A(n12263), .ZN(n12266) );
  INV_X1 U14698 ( .A(n12264), .ZN(n12265) );
  NAND2_X1 U14699 ( .A1(n12266), .A2(n12265), .ZN(n12267) );
  AND2_X1 U14700 ( .A1(n13837), .A2(n13890), .ZN(n12268) );
  INV_X1 U14701 ( .A(n13890), .ZN(n12269) );
  OR2_X1 U14702 ( .A1(n12269), .A2(n13889), .ZN(n13869) );
  AND2_X1 U14703 ( .A1(n13869), .A2(n13873), .ZN(n12270) );
  NAND2_X1 U14704 ( .A1(n13870), .A2(n12270), .ZN(n12283) );
  NAND2_X1 U14705 ( .A1(n14226), .A2(n12303), .ZN(n12272) );
  NAND2_X1 U14706 ( .A1(n10746), .A2(n14068), .ZN(n12271) );
  NAND2_X1 U14707 ( .A1(n12272), .A2(n12271), .ZN(n12274) );
  XNOR2_X1 U14708 ( .A(n12274), .B(n12273), .ZN(n12278) );
  NOR2_X1 U14709 ( .A1(n12276), .A2(n12275), .ZN(n12277) );
  AOI21_X1 U14710 ( .B1(n14226), .B2(n10746), .A(n12277), .ZN(n12279) );
  NAND2_X1 U14711 ( .A1(n12278), .A2(n12279), .ZN(n12284) );
  INV_X1 U14712 ( .A(n12278), .ZN(n12281) );
  INV_X1 U14713 ( .A(n12279), .ZN(n12280) );
  NAND2_X1 U14714 ( .A1(n12281), .A2(n12280), .ZN(n12282) );
  NAND2_X1 U14715 ( .A1(n12283), .A2(n13871), .ZN(n13875) );
  NAND2_X1 U14716 ( .A1(n14221), .A2(n12303), .ZN(n12286) );
  NAND2_X1 U14717 ( .A1(n10746), .A2(n14085), .ZN(n12285) );
  NAND2_X1 U14718 ( .A1(n12286), .A2(n12285), .ZN(n12287) );
  XNOR2_X1 U14719 ( .A(n12287), .B(n9355), .ZN(n12291) );
  NAND2_X1 U14720 ( .A1(n14221), .A2(n10746), .ZN(n12289) );
  NAND2_X1 U14721 ( .A1(n12301), .A2(n14085), .ZN(n12288) );
  NAND2_X1 U14722 ( .A1(n12289), .A2(n12288), .ZN(n12290) );
  NOR2_X1 U14723 ( .A1(n12291), .A2(n12290), .ZN(n12292) );
  AOI21_X1 U14724 ( .B1(n12291), .B2(n12290), .A(n12292), .ZN(n13953) );
  NAND2_X1 U14725 ( .A1(n14216), .A2(n12303), .ZN(n12294) );
  NAND2_X1 U14726 ( .A1(n10746), .A2(n14069), .ZN(n12293) );
  NAND2_X1 U14727 ( .A1(n12294), .A2(n12293), .ZN(n12295) );
  XNOR2_X1 U14728 ( .A(n12295), .B(n9355), .ZN(n12299) );
  NAND2_X1 U14729 ( .A1(n14216), .A2(n10746), .ZN(n12297) );
  NAND2_X1 U14730 ( .A1(n12301), .A2(n14069), .ZN(n12296) );
  NAND2_X1 U14731 ( .A1(n12297), .A2(n12296), .ZN(n12298) );
  NOR2_X1 U14732 ( .A1(n12299), .A2(n12298), .ZN(n12300) );
  AOI21_X1 U14733 ( .B1(n12299), .B2(n12298), .A(n12300), .ZN(n13826) );
  AOI22_X1 U14734 ( .A1(n14209), .A2(n10746), .B1(n12301), .B2(n13975), .ZN(
        n12302) );
  XNOR2_X1 U14735 ( .A(n12302), .B(n9355), .ZN(n12305) );
  AOI22_X1 U14736 ( .A1(n14209), .A2(n12303), .B1(n10746), .B2(n13975), .ZN(
        n12304) );
  XNOR2_X1 U14737 ( .A(n12305), .B(n12304), .ZN(n12306) );
  XNOR2_X1 U14738 ( .A(n12307), .B(n12306), .ZN(n12316) );
  OAI22_X1 U14739 ( .A1(n13966), .A2(n12309), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n12308), .ZN(n12314) );
  OAI22_X1 U14740 ( .A1(n12312), .A2(n12311), .B1(n14469), .B2(n12310), .ZN(
        n12313) );
  AOI211_X1 U14741 ( .C1(n14209), .C2(n14463), .A(n12314), .B(n12313), .ZN(
        n12315) );
  OAI21_X1 U14742 ( .B1(n12316), .B2(n13938), .A(n12315), .ZN(P1_U3220) );
  INV_X1 U14743 ( .A(n12317), .ZN(n13819) );
  OAI222_X1 U14744 ( .A1(n14292), .A2(n12318), .B1(n14296), .B2(n13819), .C1(
        n9387), .C2(P1_U3086), .ZN(P1_U3330) );
  OAI211_X1 U14745 ( .C1(n12321), .C2(n12320), .A(n12319), .B(n12502), .ZN(
        n12326) );
  AOI22_X1 U14746 ( .A1(n12476), .A2(n12588), .B1(P3_U3151), .B2(
        P3_REG3_REG_7__SCAN_IN), .ZN(n12325) );
  AOI22_X1 U14747 ( .A1(n12441), .A2(n12760), .B1(n12471), .B2(n12758), .ZN(
        n12324) );
  NAND2_X1 U14748 ( .A1(n12497), .A2(n12322), .ZN(n12323) );
  NAND4_X1 U14749 ( .A1(n12326), .A2(n12325), .A3(n12324), .A4(n12323), .ZN(
        P3_U3153) );
  OAI21_X1 U14750 ( .B1(n12329), .B2(n12328), .A(n12327), .ZN(n12330) );
  NAND2_X1 U14751 ( .A1(n12330), .A2(n12502), .ZN(n12335) );
  NAND2_X1 U14752 ( .A1(n13050), .A2(n12441), .ZN(n12331) );
  NAND2_X1 U14753 ( .A1(P3_REG3_REG_14__SCAN_IN), .A2(P3_U3151), .ZN(n12798)
         );
  OAI211_X1 U14754 ( .C1(n12332), .C2(n12443), .A(n12331), .B(n12798), .ZN(
        n12333) );
  AOI21_X1 U14755 ( .B1(n13053), .B2(n12497), .A(n12333), .ZN(n12334) );
  OAI211_X1 U14756 ( .C1(n12500), .C2(n14413), .A(n12335), .B(n12334), .ZN(
        P3_U3155) );
  INV_X1 U14757 ( .A(n13134), .ZN(n12942) );
  OAI21_X1 U14758 ( .B1(n12450), .B2(n12337), .A(n12336), .ZN(n12338) );
  NAND2_X1 U14759 ( .A1(n12338), .A2(n12502), .ZN(n12343) );
  NOR2_X1 U14760 ( .A1(n12389), .A2(n15111), .ZN(n12339) );
  AOI21_X1 U14761 ( .B1(n12751), .B2(n13098), .A(n12339), .ZN(n12938) );
  OAI22_X1 U14762 ( .A1(n12938), .A2(n12486), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n12340), .ZN(n12341) );
  AOI21_X1 U14763 ( .B1(n12940), .B2(n12497), .A(n12341), .ZN(n12342) );
  OAI211_X1 U14764 ( .C1(n12942), .C2(n12500), .A(n12343), .B(n12342), .ZN(
        P3_U3156) );
  NAND2_X1 U14765 ( .A1(n12344), .A2(n12345), .ZN(n12347) );
  AOI21_X1 U14766 ( .B1(n12347), .B2(n12346), .A(n12478), .ZN(n12350) );
  CLKBUF_X1 U14767 ( .A(n12348), .Z(n12349) );
  NAND2_X1 U14768 ( .A1(n12350), .A2(n12349), .ZN(n12355) );
  INV_X1 U14769 ( .A(n12464), .ZN(n13101) );
  AOI22_X1 U14770 ( .A1(n13101), .A2(n12471), .B1(P3_REG3_REG_10__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12351) );
  OAI21_X1 U14771 ( .B1(n12352), .B2(n12474), .A(n12351), .ZN(n12353) );
  AOI21_X1 U14772 ( .B1(n13104), .B2(n12497), .A(n12353), .ZN(n12354) );
  OAI211_X1 U14773 ( .C1(n12500), .C2(n13233), .A(n12355), .B(n12354), .ZN(
        P3_U3157) );
  XNOR2_X1 U14774 ( .A(n12357), .B(n12356), .ZN(n12362) );
  NAND2_X1 U14775 ( .A1(n12753), .A2(n12471), .ZN(n12358) );
  NAND2_X1 U14776 ( .A1(P3_U3151), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n12856)
         );
  OAI211_X1 U14777 ( .C1(n13018), .C2(n12474), .A(n12358), .B(n12856), .ZN(
        n12359) );
  AOI21_X1 U14778 ( .B1(n12992), .B2(n12497), .A(n12359), .ZN(n12361) );
  NAND2_X1 U14779 ( .A1(n12991), .A2(n12476), .ZN(n12360) );
  OAI211_X1 U14780 ( .C1(n12362), .C2(n12478), .A(n12361), .B(n12360), .ZN(
        P3_U3159) );
  OAI21_X1 U14781 ( .B1(n12365), .B2(n12364), .A(n12363), .ZN(n12366) );
  NAND2_X1 U14782 ( .A1(n12366), .A2(n12502), .ZN(n12370) );
  AOI22_X1 U14783 ( .A1(n12751), .A2(n13100), .B1(n13098), .B2(n12753), .ZN(
        n12964) );
  OAI22_X1 U14784 ( .A1(n12964), .A2(n12486), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n12367), .ZN(n12368) );
  AOI21_X1 U14785 ( .B1(n12966), .B2(n12497), .A(n12368), .ZN(n12369) );
  OAI211_X1 U14786 ( .C1(n13210), .C2(n12500), .A(n12370), .B(n12369), .ZN(
        P3_U3163) );
  INV_X1 U14787 ( .A(n12371), .ZN(n12372) );
  XOR2_X1 U14788 ( .A(n12371), .B(n12373), .Z(n12463) );
  NOR2_X1 U14789 ( .A1(n12463), .A2(n12464), .ZN(n12462) );
  AOI21_X1 U14790 ( .B1(n12373), .B2(n12372), .A(n12462), .ZN(n12376) );
  XNOR2_X1 U14791 ( .A(n12374), .B(n13087), .ZN(n12375) );
  XNOR2_X1 U14792 ( .A(n12376), .B(n12375), .ZN(n12381) );
  AOI22_X1 U14793 ( .A1(n13098), .A2(n13101), .B1(n13050), .B2(n13100), .ZN(
        n13077) );
  OAI22_X1 U14794 ( .A1(n13077), .A2(n12486), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n12377), .ZN(n12378) );
  AOI21_X1 U14795 ( .B1(n13079), .B2(n12497), .A(n12378), .ZN(n12380) );
  NAND2_X1 U14796 ( .A1(n14425), .A2(n12476), .ZN(n12379) );
  OAI211_X1 U14797 ( .C1(n12381), .C2(n12478), .A(n12380), .B(n12379), .ZN(
        P3_U3164) );
  INV_X1 U14798 ( .A(n12383), .ZN(n12388) );
  NOR3_X1 U14799 ( .A1(n12384), .A2(n12386), .A3(n12385), .ZN(n12387) );
  OAI21_X1 U14800 ( .B1(n12388), .B2(n12387), .A(n12502), .ZN(n12395) );
  OR2_X1 U14801 ( .A1(n12389), .A2(n15109), .ZN(n12391) );
  NAND2_X1 U14802 ( .A1(n12747), .A2(n13100), .ZN(n12390) );
  AND2_X1 U14803 ( .A1(n12391), .A2(n12390), .ZN(n12904) );
  OAI22_X1 U14804 ( .A1(n12904), .A2(n12486), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n12392), .ZN(n12393) );
  AOI21_X1 U14805 ( .B1(n12906), .B2(n12497), .A(n12393), .ZN(n12394) );
  OAI211_X1 U14806 ( .C1(n13197), .C2(n12500), .A(n12395), .B(n12394), .ZN(
        P3_U3165) );
  OR2_X1 U14807 ( .A1(n12398), .A2(n12397), .ZN(n12400) );
  AOI22_X1 U14808 ( .A1(n12396), .A2(n12400), .B1(n12399), .B2(n12398), .ZN(
        n12405) );
  AOI22_X1 U14809 ( .A1(n13051), .A2(n13098), .B1(n13100), .B2(n12756), .ZN(
        n13029) );
  OAI22_X1 U14810 ( .A1(n13029), .A2(n12486), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n12401), .ZN(n12402) );
  AOI21_X1 U14811 ( .B1(n13031), .B2(n12497), .A(n12402), .ZN(n12404) );
  NAND2_X1 U14812 ( .A1(n13167), .A2(n12476), .ZN(n12403) );
  OAI211_X1 U14813 ( .C1(n12405), .C2(n12478), .A(n12404), .B(n12403), .ZN(
        P3_U3166) );
  XNOR2_X1 U14814 ( .A(n12396), .B(n12406), .ZN(n12411) );
  AOI22_X1 U14815 ( .A1(n12471), .A2(n12755), .B1(P3_REG3_REG_17__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12407) );
  OAI21_X1 U14816 ( .B1(n13017), .B2(n12474), .A(n12407), .ZN(n12409) );
  NOR2_X1 U14817 ( .A1(n13226), .A2(n12500), .ZN(n12408) );
  AOI211_X1 U14818 ( .C1(n13019), .C2(n12497), .A(n12409), .B(n12408), .ZN(
        n12410) );
  OAI21_X1 U14819 ( .B1(n12411), .B2(n12478), .A(n12410), .ZN(P3_U3168) );
  AND3_X1 U14820 ( .A1(n12336), .A2(n6490), .A3(n12412), .ZN(n12413) );
  OAI21_X1 U14821 ( .B1(n12384), .B2(n12413), .A(n12502), .ZN(n12419) );
  OR2_X1 U14822 ( .A1(n12450), .A2(n15109), .ZN(n12414) );
  OAI21_X1 U14823 ( .B1(n12415), .B2(n15111), .A(n12414), .ZN(n12914) );
  AOI22_X1 U14824 ( .A1(n12914), .A2(n12496), .B1(P3_REG3_REG_24__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12418) );
  NAND2_X1 U14825 ( .A1(n12922), .A2(n12476), .ZN(n12417) );
  NAND2_X1 U14826 ( .A1(n12497), .A2(n12923), .ZN(n12416) );
  NAND4_X1 U14827 ( .A1(n12419), .A2(n12418), .A3(n12417), .A4(n12416), .ZN(
        P3_U3169) );
  INV_X1 U14828 ( .A(n12344), .ZN(n12420) );
  AOI21_X1 U14829 ( .B1(n12422), .B2(n12421), .A(n12420), .ZN(n12429) );
  AOI22_X1 U14830 ( .A1(n12441), .A2(n12758), .B1(n12471), .B2(n13086), .ZN(
        n12425) );
  AOI22_X1 U14831 ( .A1(n12476), .A2(n12423), .B1(P3_REG3_REG_9__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12424) );
  NAND2_X1 U14832 ( .A1(n12425), .A2(n12424), .ZN(n12426) );
  AOI21_X1 U14833 ( .B1(n12427), .B2(n12497), .A(n12426), .ZN(n12428) );
  OAI21_X1 U14834 ( .B1(n12429), .B2(n12478), .A(n12428), .ZN(P3_U3171) );
  XNOR2_X1 U14835 ( .A(n12431), .B(n12430), .ZN(n12436) );
  AOI22_X1 U14836 ( .A1(n12752), .A2(n12471), .B1(P3_REG3_REG_20__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12433) );
  NAND2_X1 U14837 ( .A1(n12977), .A2(n12497), .ZN(n12432) );
  OAI211_X1 U14838 ( .C1(n13003), .C2(n12474), .A(n12433), .B(n12432), .ZN(
        n12434) );
  AOI21_X1 U14839 ( .B1(n13145), .B2(n12476), .A(n12434), .ZN(n12435) );
  OAI21_X1 U14840 ( .B1(n12436), .B2(n12478), .A(n12435), .ZN(P3_U3173) );
  XNOR2_X1 U14841 ( .A(n12438), .B(n12437), .ZN(n12439) );
  XNOR2_X1 U14842 ( .A(n12440), .B(n12439), .ZN(n12447) );
  AOI22_X1 U14843 ( .A1(n12441), .A2(n13087), .B1(P3_REG3_REG_13__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12442) );
  OAI21_X1 U14844 ( .B1(n12493), .B2(n12443), .A(n12442), .ZN(n12445) );
  NOR2_X1 U14845 ( .A1(n14417), .A2(n12500), .ZN(n12444) );
  AOI211_X1 U14846 ( .C1(n13065), .C2(n12497), .A(n12445), .B(n12444), .ZN(
        n12446) );
  OAI21_X1 U14847 ( .B1(n12447), .B2(n12478), .A(n12446), .ZN(P3_U3174) );
  AOI21_X1 U14848 ( .B1(n12751), .B2(n12449), .A(n12448), .ZN(n12456) );
  INV_X1 U14849 ( .A(n12955), .ZN(n12453) );
  OAI22_X1 U14850 ( .A1(n12973), .A2(n15109), .B1(n12450), .B2(n15111), .ZN(
        n12951) );
  AOI22_X1 U14851 ( .A1(n12951), .A2(n12496), .B1(P3_REG3_REG_22__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12451) );
  OAI21_X1 U14852 ( .B1(n12453), .B2(n12452), .A(n12451), .ZN(n12454) );
  AOI21_X1 U14853 ( .B1(n12954), .B2(n12476), .A(n12454), .ZN(n12455) );
  OAI21_X1 U14854 ( .B1(n12456), .B2(n12478), .A(n12455), .ZN(P3_U3175) );
  INV_X1 U14855 ( .A(n12457), .ZN(n12458) );
  AOI21_X1 U14856 ( .B1(n12471), .B2(n13087), .A(n12458), .ZN(n12460) );
  NAND2_X1 U14857 ( .A1(n12497), .A2(n13091), .ZN(n12459) );
  OAI211_X1 U14858 ( .C1(n12461), .C2(n12474), .A(n12460), .B(n12459), .ZN(
        n12466) );
  AOI211_X1 U14859 ( .C1(n12464), .C2(n12463), .A(n12478), .B(n12462), .ZN(
        n12465) );
  AOI211_X1 U14860 ( .C1(n12476), .C2(n12467), .A(n12466), .B(n12465), .ZN(
        n12468) );
  INV_X1 U14861 ( .A(n12468), .ZN(P3_U3176) );
  XNOR2_X1 U14862 ( .A(n12469), .B(n12470), .ZN(n12479) );
  AOI22_X1 U14863 ( .A1(n12754), .A2(n12471), .B1(P3_REG3_REG_18__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12473) );
  NAND2_X1 U14864 ( .A1(n12497), .A2(n13005), .ZN(n12472) );
  OAI211_X1 U14865 ( .C1(n13002), .C2(n12474), .A(n12473), .B(n12472), .ZN(
        n12475) );
  AOI21_X1 U14866 ( .B1(n13004), .B2(n12476), .A(n12475), .ZN(n12477) );
  OAI21_X1 U14867 ( .B1(n12479), .B2(n12478), .A(n12477), .ZN(P3_U3178) );
  OAI21_X1 U14868 ( .B1(n12483), .B2(n12482), .A(n12481), .ZN(n12484) );
  NAND2_X1 U14869 ( .A1(n12484), .A2(n12502), .ZN(n12489) );
  AOI22_X1 U14870 ( .A1(n12748), .A2(n13098), .B1(n13100), .B2(n12746), .ZN(
        n12890) );
  OAI22_X1 U14871 ( .A1(n12890), .A2(n12486), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n12485), .ZN(n12487) );
  AOI21_X1 U14872 ( .B1(n12894), .B2(n12497), .A(n12487), .ZN(n12488) );
  OAI211_X1 U14873 ( .C1(n13193), .C2(n12500), .A(n12489), .B(n12488), .ZN(
        P3_U3180) );
  XNOR2_X1 U14874 ( .A(n12490), .B(n13051), .ZN(n12491) );
  XNOR2_X1 U14875 ( .A(n12492), .B(n12491), .ZN(n12503) );
  OR2_X1 U14876 ( .A1(n13017), .A2(n15111), .ZN(n12495) );
  OR2_X1 U14877 ( .A1(n12493), .A2(n15109), .ZN(n12494) );
  NAND2_X1 U14878 ( .A1(n12495), .A2(n12494), .ZN(n13039) );
  AOI22_X1 U14879 ( .A1(n13039), .A2(n12496), .B1(P3_REG3_REG_15__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12499) );
  NAND2_X1 U14880 ( .A1(n12497), .A2(n13042), .ZN(n12498) );
  OAI211_X1 U14881 ( .C1(n13231), .C2(n12500), .A(n12499), .B(n12498), .ZN(
        n12501) );
  AOI21_X1 U14882 ( .B1(n12503), .B2(n12502), .A(n12501), .ZN(n12504) );
  INV_X1 U14883 ( .A(n12504), .ZN(P3_U3181) );
  INV_X1 U14884 ( .A(n12505), .ZN(n12528) );
  NOR2_X1 U14885 ( .A1(n12506), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n12508) );
  OAI22_X1 U14886 ( .A1(n12509), .A2(n12508), .B1(P1_DATAO_REG_30__SCAN_IN), 
        .B2(n12507), .ZN(n12511) );
  XNOR2_X1 U14887 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(P2_DATAO_REG_31__SCAN_IN), 
        .ZN(n12510) );
  XNOR2_X1 U14888 ( .A(n12511), .B(n12510), .ZN(n13240) );
  NAND2_X1 U14889 ( .A1(n13240), .A2(n12520), .ZN(n12513) );
  OR2_X1 U14890 ( .A1(n6480), .A2(n13245), .ZN(n12512) );
  NAND2_X1 U14891 ( .A1(n12513), .A2(n12512), .ZN(n12530) );
  NAND2_X1 U14892 ( .A1(n12514), .A2(P3_REG2_REG_31__SCAN_IN), .ZN(n12518) );
  NAND2_X1 U14893 ( .A1(n7522), .A2(P3_REG1_REG_31__SCAN_IN), .ZN(n12517) );
  NAND2_X1 U14894 ( .A1(n7454), .A2(P3_REG0_REG_31__SCAN_IN), .ZN(n12516) );
  OR2_X1 U14895 ( .A1(n12530), .A2(n12861), .ZN(n12526) );
  NAND2_X1 U14896 ( .A1(n12521), .A2(n12520), .ZN(n12524) );
  OR2_X1 U14897 ( .A1(n6481), .A2(n12522), .ZN(n12523) );
  NAND2_X1 U14898 ( .A1(n13186), .A2(n12529), .ZN(n12525) );
  NAND2_X1 U14899 ( .A1(n12526), .A2(n12525), .ZN(n12722) );
  INV_X1 U14900 ( .A(n13186), .ZN(n12866) );
  INV_X1 U14901 ( .A(n12861), .ZN(n12743) );
  OAI21_X1 U14902 ( .B1(n12866), .B2(n12743), .A(n12686), .ZN(n12527) );
  NOR2_X1 U14903 ( .A1(n13184), .A2(n12743), .ZN(n12696) );
  NOR2_X1 U14904 ( .A1(n13186), .A2(n12529), .ZN(n12721) );
  XNOR2_X1 U14905 ( .A(n12533), .B(n12857), .ZN(n12734) );
  INV_X1 U14906 ( .A(n12534), .ZN(n12541) );
  NOR2_X1 U14907 ( .A1(n12541), .A2(n12539), .ZN(n12538) );
  OAI22_X1 U14908 ( .A1(n12541), .A2(n12540), .B1(n12536), .B2(n12535), .ZN(
        n12537) );
  MUX2_X1 U14909 ( .A(n12538), .B(n12537), .S(n12671), .Z(n12684) );
  NAND2_X1 U14910 ( .A1(n12540), .A2(n12539), .ZN(n12893) );
  NAND2_X1 U14911 ( .A1(n12660), .A2(n12658), .ZN(n12949) );
  INV_X1 U14912 ( .A(n12949), .ZN(n12657) );
  NAND2_X1 U14913 ( .A1(n12752), .A2(n12671), .ZN(n12544) );
  NAND2_X1 U14914 ( .A1(n12973), .A2(n12689), .ZN(n12543) );
  MUX2_X1 U14915 ( .A(n12544), .B(n12543), .S(n12545), .Z(n12656) );
  XNOR2_X1 U14916 ( .A(n12545), .B(n12973), .ZN(n12962) );
  INV_X1 U14917 ( .A(n12962), .ZN(n12654) );
  INV_X1 U14918 ( .A(n12546), .ZN(n12549) );
  NAND2_X1 U14919 ( .A1(n12549), .A2(n12547), .ZN(n12548) );
  NAND2_X1 U14920 ( .A1(n12548), .A2(n12671), .ZN(n12551) );
  NAND3_X1 U14921 ( .A1(n12557), .A2(n12549), .A3(n12739), .ZN(n12550) );
  NAND2_X1 U14922 ( .A1(n12551), .A2(n12550), .ZN(n12555) );
  NAND2_X1 U14923 ( .A1(n12553), .A2(n12552), .ZN(n12554) );
  NAND3_X1 U14924 ( .A1(n12555), .A2(n12554), .A3(n12559), .ZN(n12560) );
  NAND3_X1 U14925 ( .A1(n12560), .A2(n12556), .A3(n12557), .ZN(n12558) );
  NAND3_X1 U14926 ( .A1(n12558), .A2(n12563), .A3(n7436), .ZN(n12568) );
  NAND3_X1 U14927 ( .A1(n12560), .A2(n12556), .A3(n12559), .ZN(n12566) );
  AND2_X1 U14928 ( .A1(n12562), .A2(n12561), .ZN(n12565) );
  INV_X1 U14929 ( .A(n12563), .ZN(n12564) );
  AOI21_X1 U14930 ( .B1(n12566), .B2(n12565), .A(n12564), .ZN(n12567) );
  MUX2_X1 U14931 ( .A(n12568), .B(n12567), .S(n12689), .Z(n12571) );
  NAND3_X1 U14932 ( .A1(n12763), .A2(n12671), .A3(n15135), .ZN(n12569) );
  NAND3_X1 U14933 ( .A1(n12571), .A2(n12570), .A3(n12569), .ZN(n12575) );
  MUX2_X1 U14934 ( .A(n12573), .B(n12572), .S(n12689), .Z(n12574) );
  NAND3_X1 U14935 ( .A1(n12575), .A2(n12701), .A3(n12574), .ZN(n12582) );
  NAND2_X1 U14936 ( .A1(n12584), .A2(n12576), .ZN(n12579) );
  NAND2_X1 U14937 ( .A1(n12583), .A2(n12577), .ZN(n12578) );
  MUX2_X1 U14938 ( .A(n12579), .B(n12578), .S(n12671), .Z(n12580) );
  INV_X1 U14939 ( .A(n12580), .ZN(n12581) );
  NAND2_X1 U14940 ( .A1(n12582), .A2(n12581), .ZN(n12586) );
  MUX2_X1 U14941 ( .A(n12584), .B(n12583), .S(n12689), .Z(n12585) );
  NAND3_X1 U14942 ( .A1(n12586), .A2(n12706), .A3(n12585), .ZN(n12592) );
  NAND2_X1 U14943 ( .A1(n12759), .A2(n12671), .ZN(n12590) );
  NAND2_X1 U14944 ( .A1(n12587), .A2(n12689), .ZN(n12589) );
  MUX2_X1 U14945 ( .A(n12590), .B(n12589), .S(n12588), .Z(n12591) );
  NAND3_X1 U14946 ( .A1(n12592), .A2(n12707), .A3(n12591), .ZN(n12597) );
  INV_X1 U14947 ( .A(n12593), .ZN(n12700) );
  MUX2_X1 U14948 ( .A(n12595), .B(n12594), .S(n12689), .Z(n12596) );
  NAND3_X1 U14949 ( .A1(n12597), .A2(n12700), .A3(n12596), .ZN(n12601) );
  MUX2_X1 U14950 ( .A(n12599), .B(n12598), .S(n12689), .Z(n12600) );
  NAND4_X1 U14951 ( .A1(n12601), .A2(n7573), .A3(n7587), .A4(n12600), .ZN(
        n12616) );
  OAI211_X1 U14952 ( .C1(n12606), .C2(n12603), .A(n12610), .B(n12602), .ZN(
        n12608) );
  OAI211_X1 U14953 ( .C1(n12606), .C2(n12605), .A(n12611), .B(n12604), .ZN(
        n12607) );
  MUX2_X1 U14954 ( .A(n12608), .B(n12607), .S(n12671), .Z(n12609) );
  INV_X1 U14955 ( .A(n12609), .ZN(n12615) );
  INV_X1 U14956 ( .A(n12610), .ZN(n12613) );
  INV_X1 U14957 ( .A(n12611), .ZN(n12612) );
  MUX2_X1 U14958 ( .A(n12613), .B(n12612), .S(n12689), .Z(n12614) );
  AOI21_X1 U14959 ( .B1(n12616), .B2(n12615), .A(n12614), .ZN(n12620) );
  INV_X1 U14960 ( .A(n13058), .ZN(n13049) );
  MUX2_X1 U14961 ( .A(n12618), .B(n12617), .S(n12689), .Z(n12619) );
  OAI211_X1 U14962 ( .C1(n12620), .C2(n13070), .A(n13049), .B(n12619), .ZN(
        n12624) );
  MUX2_X1 U14963 ( .A(n12622), .B(n12621), .S(n12671), .Z(n12623) );
  NAND3_X1 U14964 ( .A1(n12624), .A2(n13038), .A3(n12623), .ZN(n12629) );
  OAI21_X1 U14965 ( .B1(n13167), .B2(n13017), .A(n12625), .ZN(n12626) );
  NAND2_X1 U14966 ( .A1(n12626), .A2(n12671), .ZN(n12628) );
  AOI21_X1 U14967 ( .B1(n12629), .B2(n12628), .A(n12627), .ZN(n12633) );
  AOI21_X1 U14968 ( .B1(n12630), .B2(n13024), .A(n12671), .ZN(n12632) );
  OR3_X1 U14969 ( .A1(n13167), .A2(n13017), .A3(n12671), .ZN(n12631) );
  OAI21_X1 U14970 ( .B1(n12633), .B2(n12632), .A(n12631), .ZN(n12640) );
  INV_X1 U14971 ( .A(n12634), .ZN(n12635) );
  AOI21_X1 U14972 ( .B1(n12641), .B2(n12635), .A(n12671), .ZN(n12636) );
  NAND2_X1 U14973 ( .A1(n12637), .A2(n12636), .ZN(n12643) );
  INV_X1 U14974 ( .A(n12638), .ZN(n12639) );
  AOI22_X1 U14975 ( .A1(n12640), .A2(n13013), .B1(n12643), .B2(n12639), .ZN(
        n12645) );
  NAND3_X1 U14976 ( .A1(n12647), .A2(n12671), .A3(n12641), .ZN(n12642) );
  NAND2_X1 U14977 ( .A1(n12643), .A2(n12642), .ZN(n12644) );
  OAI21_X1 U14978 ( .B1(n12645), .B2(n7893), .A(n12644), .ZN(n12649) );
  MUX2_X1 U14979 ( .A(n12647), .B(n12646), .S(n12671), .Z(n12648) );
  NAND3_X1 U14980 ( .A1(n12649), .A2(n12971), .A3(n12648), .ZN(n12653) );
  MUX2_X1 U14981 ( .A(n12651), .B(n12650), .S(n12689), .Z(n12652) );
  NAND3_X1 U14982 ( .A1(n12654), .A2(n12653), .A3(n12652), .ZN(n12655) );
  NAND3_X1 U14983 ( .A1(n12657), .A2(n12656), .A3(n12655), .ZN(n12659) );
  NAND3_X1 U14984 ( .A1(n12930), .A2(n12658), .A3(n12659), .ZN(n12664) );
  NAND3_X1 U14985 ( .A1(n12930), .A2(n12660), .A3(n12659), .ZN(n12662) );
  AND2_X1 U14986 ( .A1(n12662), .A2(n12661), .ZN(n12663) );
  MUX2_X1 U14987 ( .A(n12664), .B(n12663), .S(n12689), .Z(n12666) );
  OAI21_X1 U14988 ( .B1(n12916), .B2(n12666), .A(n12665), .ZN(n12676) );
  INV_X1 U14989 ( .A(n12916), .ZN(n12670) );
  XNOR2_X1 U14990 ( .A(n12667), .B(n12689), .ZN(n12668) );
  AOI21_X1 U14991 ( .B1(n12670), .B2(n12669), .A(n12668), .ZN(n12675) );
  MUX2_X1 U14992 ( .A(n12673), .B(n12672), .S(n12671), .Z(n12674) );
  OAI21_X1 U14993 ( .B1(n12676), .B2(n12675), .A(n12674), .ZN(n12682) );
  INV_X1 U14994 ( .A(n12719), .ZN(n12681) );
  NAND2_X1 U14995 ( .A1(n12677), .A2(n12679), .ZN(n12678) );
  MUX2_X1 U14996 ( .A(n12679), .B(n12678), .S(n12689), .Z(n12680) );
  OAI211_X1 U14997 ( .C1(n12720), .C2(n12682), .A(n12681), .B(n12680), .ZN(
        n12683) );
  AOI21_X1 U14998 ( .B1(n12685), .B2(n12684), .A(n12683), .ZN(n12693) );
  NAND2_X1 U14999 ( .A1(n12687), .A2(n12689), .ZN(n12688) );
  NAND2_X1 U15000 ( .A1(n12686), .A2(n12688), .ZN(n12692) );
  NAND2_X1 U15001 ( .A1(n12693), .A2(n12689), .ZN(n12690) );
  INV_X1 U15002 ( .A(n12696), .ZN(n12723) );
  NAND3_X1 U15003 ( .A1(n12694), .A2(n12735), .A3(n12723), .ZN(n12731) );
  OAI21_X1 U15004 ( .B1(n12697), .B2(n12696), .A(n12695), .ZN(n12730) );
  INV_X1 U15005 ( .A(n12930), .ZN(n12936) );
  XNOR2_X1 U15006 ( .A(n12991), .B(n13003), .ZN(n12988) );
  NOR2_X1 U15007 ( .A1(n12699), .A2(n12698), .ZN(n12702) );
  NAND4_X1 U15008 ( .A1(n12702), .A2(n12701), .A3(n12556), .A4(n12700), .ZN(
        n12710) );
  NOR2_X1 U15009 ( .A1(n12704), .A2(n12703), .ZN(n12708) );
  NAND4_X1 U15010 ( .A1(n12708), .A2(n12707), .A3(n12706), .A4(n12705), .ZN(
        n12709) );
  NOR2_X1 U15011 ( .A1(n12710), .A2(n12709), .ZN(n12712) );
  NAND4_X1 U15012 ( .A1(n12712), .A2(n12711), .A3(n7587), .A4(n7573), .ZN(
        n12713) );
  NOR2_X1 U15013 ( .A1(n12713), .A2(n13070), .ZN(n12714) );
  NAND4_X1 U15014 ( .A1(n13027), .A2(n13038), .A3(n13049), .A4(n12714), .ZN(
        n12715) );
  OR4_X1 U15015 ( .A1(n7893), .A2(n12988), .A3(n13015), .A4(n12715), .ZN(
        n12716) );
  OR4_X1 U15016 ( .A1(n12949), .A2(n12962), .A3(n12982), .A4(n12716), .ZN(
        n12717) );
  OR4_X1 U15017 ( .A1(n12901), .A2(n12916), .A3(n12936), .A4(n12717), .ZN(
        n12718) );
  NOR4_X1 U15018 ( .A1(n12721), .A2(n12720), .A3(n12719), .A4(n12718), .ZN(
        n12725) );
  INV_X1 U15019 ( .A(n12722), .ZN(n12724) );
  NAND3_X1 U15020 ( .A1(n12725), .A2(n12724), .A3(n12723), .ZN(n12726) );
  XNOR2_X1 U15021 ( .A(n12726), .B(n12825), .ZN(n12728) );
  NAND3_X1 U15022 ( .A1(n12731), .A2(n12730), .A3(n12729), .ZN(n12732) );
  AOI21_X1 U15023 ( .B1(n12734), .B2(n12733), .A(n12732), .ZN(n12742) );
  NAND4_X1 U15024 ( .A1(n13098), .A2(n12737), .A3(n12736), .A4(n12735), .ZN(
        n12738) );
  OAI211_X1 U15025 ( .C1(n12739), .C2(n12741), .A(n12738), .B(P3_B_REG_SCAN_IN), .ZN(n12740) );
  OAI21_X1 U15026 ( .B1(n12742), .B2(n12741), .A(n12740), .ZN(P3_U3296) );
  MUX2_X1 U15027 ( .A(P3_DATAO_REG_31__SCAN_IN), .B(n12743), .S(P3_U3897), .Z(
        P3_U3522) );
  MUX2_X1 U15028 ( .A(P3_DATAO_REG_29__SCAN_IN), .B(n12744), .S(P3_U3897), .Z(
        P3_U3520) );
  MUX2_X1 U15029 ( .A(n12745), .B(P3_DATAO_REG_28__SCAN_IN), .S(n12765), .Z(
        P3_U3519) );
  MUX2_X1 U15030 ( .A(n12746), .B(P3_DATAO_REG_27__SCAN_IN), .S(n12765), .Z(
        P3_U3518) );
  MUX2_X1 U15031 ( .A(n12747), .B(P3_DATAO_REG_26__SCAN_IN), .S(n12765), .Z(
        P3_U3517) );
  MUX2_X1 U15032 ( .A(P3_DATAO_REG_25__SCAN_IN), .B(n12748), .S(P3_U3897), .Z(
        P3_U3516) );
  MUX2_X1 U15033 ( .A(P3_DATAO_REG_24__SCAN_IN), .B(n12749), .S(P3_U3897), .Z(
        P3_U3515) );
  MUX2_X1 U15034 ( .A(P3_DATAO_REG_23__SCAN_IN), .B(n12750), .S(P3_U3897), .Z(
        P3_U3514) );
  MUX2_X1 U15035 ( .A(P3_DATAO_REG_22__SCAN_IN), .B(n12751), .S(P3_U3897), .Z(
        P3_U3513) );
  MUX2_X1 U15036 ( .A(n12752), .B(P3_DATAO_REG_21__SCAN_IN), .S(n12765), .Z(
        P3_U3512) );
  MUX2_X1 U15037 ( .A(n12753), .B(P3_DATAO_REG_20__SCAN_IN), .S(n12765), .Z(
        P3_U3511) );
  MUX2_X1 U15038 ( .A(n12754), .B(P3_DATAO_REG_19__SCAN_IN), .S(n12765), .Z(
        P3_U3510) );
  MUX2_X1 U15039 ( .A(n12755), .B(P3_DATAO_REG_18__SCAN_IN), .S(n12765), .Z(
        P3_U3509) );
  MUX2_X1 U15040 ( .A(n12756), .B(P3_DATAO_REG_17__SCAN_IN), .S(n12765), .Z(
        P3_U3508) );
  MUX2_X1 U15041 ( .A(n12757), .B(P3_DATAO_REG_16__SCAN_IN), .S(n12765), .Z(
        P3_U3507) );
  MUX2_X1 U15042 ( .A(P3_DATAO_REG_15__SCAN_IN), .B(n13051), .S(P3_U3897), .Z(
        P3_U3506) );
  MUX2_X1 U15043 ( .A(n13063), .B(P3_DATAO_REG_14__SCAN_IN), .S(n12765), .Z(
        P3_U3505) );
  MUX2_X1 U15044 ( .A(n13050), .B(P3_DATAO_REG_13__SCAN_IN), .S(n12765), .Z(
        P3_U3504) );
  MUX2_X1 U15045 ( .A(n13087), .B(P3_DATAO_REG_12__SCAN_IN), .S(n12765), .Z(
        P3_U3503) );
  MUX2_X1 U15046 ( .A(P3_DATAO_REG_11__SCAN_IN), .B(n13101), .S(P3_U3897), .Z(
        P3_U3502) );
  MUX2_X1 U15047 ( .A(n13086), .B(P3_DATAO_REG_10__SCAN_IN), .S(n12765), .Z(
        P3_U3501) );
  MUX2_X1 U15048 ( .A(n13099), .B(P3_DATAO_REG_9__SCAN_IN), .S(n12765), .Z(
        P3_U3500) );
  MUX2_X1 U15049 ( .A(n12758), .B(P3_DATAO_REG_8__SCAN_IN), .S(n12765), .Z(
        P3_U3499) );
  MUX2_X1 U15050 ( .A(n12759), .B(P3_DATAO_REG_7__SCAN_IN), .S(n12765), .Z(
        P3_U3498) );
  MUX2_X1 U15051 ( .A(n12760), .B(P3_DATAO_REG_6__SCAN_IN), .S(n12765), .Z(
        P3_U3497) );
  MUX2_X1 U15052 ( .A(n12761), .B(P3_DATAO_REG_5__SCAN_IN), .S(n12765), .Z(
        P3_U3496) );
  MUX2_X1 U15053 ( .A(n12762), .B(P3_DATAO_REG_4__SCAN_IN), .S(n12765), .Z(
        P3_U3495) );
  MUX2_X1 U15054 ( .A(n12763), .B(P3_DATAO_REG_3__SCAN_IN), .S(n12765), .Z(
        P3_U3494) );
  MUX2_X1 U15055 ( .A(n6469), .B(P3_DATAO_REG_2__SCAN_IN), .S(n12765), .Z(
        P3_U3493) );
  MUX2_X1 U15056 ( .A(P3_DATAO_REG_1__SCAN_IN), .B(n12764), .S(P3_U3897), .Z(
        P3_U3492) );
  MUX2_X1 U15057 ( .A(n12766), .B(P3_DATAO_REG_0__SCAN_IN), .S(n12765), .Z(
        P3_U3491) );
  INV_X1 U15058 ( .A(P3_REG2_REG_13__SCAN_IN), .ZN(n13067) );
  AOI21_X1 U15059 ( .B1(n13067), .B2(n12768), .A(n12787), .ZN(n12784) );
  NAND2_X1 U15060 ( .A1(P3_REG1_REG_13__SCAN_IN), .A2(n12771), .ZN(n12794) );
  OAI21_X1 U15061 ( .B1(P3_REG1_REG_13__SCAN_IN), .B2(n12771), .A(n12794), 
        .ZN(n12782) );
  AOI21_X1 U15062 ( .B1(n12774), .B2(n12773), .A(n12772), .ZN(n12776) );
  MUX2_X1 U15063 ( .A(P3_REG2_REG_13__SCAN_IN), .B(P3_REG1_REG_13__SCAN_IN), 
        .S(n12836), .Z(n12801) );
  XNOR2_X1 U15064 ( .A(n12801), .B(n12802), .ZN(n12775) );
  NAND2_X1 U15065 ( .A1(n12776), .A2(n12775), .ZN(n12809) );
  OAI21_X1 U15066 ( .B1(n12776), .B2(n12775), .A(n12809), .ZN(n12777) );
  NAND2_X1 U15067 ( .A1(n12777), .A2(n15064), .ZN(n12780) );
  NOR2_X1 U15068 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n7620), .ZN(n12778) );
  AOI21_X1 U15069 ( .B1(n15094), .B2(P3_ADDR_REG_13__SCAN_IN), .A(n12778), 
        .ZN(n12779) );
  OAI211_X1 U15070 ( .C1(n15088), .C2(n12793), .A(n12780), .B(n12779), .ZN(
        n12781) );
  AOI21_X1 U15071 ( .B1(n15097), .B2(n12782), .A(n12781), .ZN(n12783) );
  OAI21_X1 U15072 ( .B1(n12784), .B2(n15101), .A(n12783), .ZN(P3_U3195) );
  NOR2_X1 U15073 ( .A1(n12802), .A2(n12785), .ZN(n12786) );
  NAND2_X1 U15074 ( .A1(n12790), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n12827) );
  OAI21_X1 U15075 ( .B1(n12790), .B2(P3_REG2_REG_14__SCAN_IN), .A(n12827), 
        .ZN(n12804) );
  NOR2_X2 U15076 ( .A1(n12788), .A2(n12804), .ZN(n12817) );
  AOI21_X1 U15077 ( .B1(n12788), .B2(n12804), .A(n12817), .ZN(n12816) );
  INV_X1 U15078 ( .A(n12790), .ZN(n12797) );
  INV_X1 U15079 ( .A(P3_REG1_REG_14__SCAN_IN), .ZN(n12789) );
  NAND2_X1 U15080 ( .A1(n12797), .A2(n12789), .ZN(n12791) );
  NAND2_X1 U15081 ( .A1(n12790), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n12844) );
  AND2_X1 U15082 ( .A1(n12791), .A2(n12844), .ZN(n12806) );
  NAND2_X1 U15083 ( .A1(n12793), .A2(n12792), .ZN(n12795) );
  NAND2_X1 U15084 ( .A1(n12795), .A2(n12794), .ZN(n12796) );
  NAND2_X1 U15085 ( .A1(n12796), .A2(n12806), .ZN(n12843) );
  OAI21_X1 U15086 ( .B1(n12806), .B2(n12796), .A(n12843), .ZN(n12814) );
  NAND2_X1 U15087 ( .A1(n15070), .A2(n12797), .ZN(n12799) );
  OAI211_X1 U15088 ( .C1(n12800), .C2(n15077), .A(n12799), .B(n12798), .ZN(
        n12813) );
  INV_X1 U15089 ( .A(n12801), .ZN(n12803) );
  NAND2_X1 U15090 ( .A1(n12803), .A2(n12802), .ZN(n12808) );
  INV_X1 U15091 ( .A(n12804), .ZN(n12805) );
  MUX2_X1 U15092 ( .A(n12806), .B(n12805), .S(n12826), .Z(n12807) );
  NAND3_X1 U15093 ( .A1(n12809), .A2(n12808), .A3(n12807), .ZN(n12829) );
  INV_X1 U15094 ( .A(n12829), .ZN(n12811) );
  AOI21_X1 U15095 ( .B1(n12809), .B2(n12808), .A(n12807), .ZN(n12810) );
  NOR3_X1 U15096 ( .A1(n12811), .A2(n12810), .A3(n15090), .ZN(n12812) );
  AOI211_X1 U15097 ( .C1(n15097), .C2(n12814), .A(n12813), .B(n12812), .ZN(
        n12815) );
  OAI21_X1 U15098 ( .B1(n12816), .B2(n15101), .A(n12815), .ZN(P3_U3196) );
  INV_X1 U15099 ( .A(P3_REG2_REG_15__SCAN_IN), .ZN(n14353) );
  AND2_X1 U15100 ( .A1(n12818), .A2(n12819), .ZN(n12820) );
  NOR2_X2 U15101 ( .A1(n14352), .A2(n12820), .ZN(n14373) );
  NAND2_X1 U15102 ( .A1(P3_REG2_REG_16__SCAN_IN), .A2(n12842), .ZN(n12821) );
  OAI21_X1 U15103 ( .B1(P3_REG2_REG_16__SCAN_IN), .B2(n12842), .A(n12821), 
        .ZN(n14372) );
  NOR2_X1 U15104 ( .A1(n14379), .A2(n12822), .ZN(n12823) );
  INV_X1 U15105 ( .A(P3_REG2_REG_17__SCAN_IN), .ZN(n14388) );
  INV_X1 U15106 ( .A(P3_REG2_REG_18__SCAN_IN), .ZN(n12824) );
  AOI22_X1 U15107 ( .A1(P3_REG2_REG_18__SCAN_IN), .A2(n14394), .B1(n12840), 
        .B2(n12824), .ZN(n14405) );
  XNOR2_X1 U15108 ( .A(n12825), .B(P3_REG2_REG_19__SCAN_IN), .ZN(n12835) );
  MUX2_X1 U15109 ( .A(P3_REG2_REG_17__SCAN_IN), .B(P3_REG1_REG_17__SCAN_IN), 
        .S(n12836), .Z(n12833) );
  MUX2_X1 U15110 ( .A(n12844), .B(n12827), .S(n12826), .Z(n12828) );
  NAND2_X1 U15111 ( .A1(n12829), .A2(n12828), .ZN(n12830) );
  INV_X1 U15112 ( .A(n12830), .ZN(n12831) );
  XNOR2_X1 U15113 ( .A(n12830), .B(n12818), .ZN(n14348) );
  MUX2_X1 U15114 ( .A(P3_REG2_REG_15__SCAN_IN), .B(P3_REG1_REG_15__SCAN_IN), 
        .S(n12836), .Z(n14349) );
  AOI21_X1 U15115 ( .B1(n12831), .B2(n14344), .A(n14347), .ZN(n14366) );
  INV_X1 U15116 ( .A(P3_REG1_REG_16__SCAN_IN), .ZN(n12841) );
  MUX2_X1 U15117 ( .A(n7204), .B(n12841), .S(n12836), .Z(n12832) );
  NOR2_X1 U15118 ( .A1(n12832), .A2(n14361), .ZN(n14362) );
  NAND2_X1 U15119 ( .A1(n12832), .A2(n14361), .ZN(n14363) );
  OAI21_X1 U15120 ( .B1(n14366), .B2(n14362), .A(n14363), .ZN(n14383) );
  XNOR2_X1 U15121 ( .A(n12833), .B(n12848), .ZN(n14384) );
  NOR2_X1 U15122 ( .A1(n14383), .A2(n14384), .ZN(n14382) );
  XNOR2_X1 U15123 ( .A(n12834), .B(n14394), .ZN(n14399) );
  MUX2_X1 U15124 ( .A(P3_REG2_REG_18__SCAN_IN), .B(P3_REG1_REG_18__SCAN_IN), 
        .S(n12836), .Z(n14400) );
  NOR2_X1 U15125 ( .A1(n14399), .A2(n14400), .ZN(n14398) );
  AOI21_X1 U15126 ( .B1(n12834), .B2(n14394), .A(n14398), .ZN(n12839) );
  INV_X1 U15127 ( .A(n12835), .ZN(n12837) );
  XNOR2_X1 U15128 ( .A(n12857), .B(P3_REG1_REG_19__SCAN_IN), .ZN(n12851) );
  MUX2_X1 U15129 ( .A(n12837), .B(n12851), .S(n12836), .Z(n12838) );
  XNOR2_X1 U15130 ( .A(n12839), .B(n12838), .ZN(n12859) );
  INV_X1 U15131 ( .A(P3_REG1_REG_18__SCAN_IN), .ZN(n13160) );
  AOI22_X1 U15132 ( .A1(P3_REG1_REG_18__SCAN_IN), .A2(n12840), .B1(n14394), 
        .B2(n13160), .ZN(n14397) );
  NAND2_X1 U15133 ( .A1(P3_REG1_REG_16__SCAN_IN), .A2(n12842), .ZN(n12847) );
  AOI22_X1 U15134 ( .A1(P3_REG1_REG_16__SCAN_IN), .A2(n12842), .B1(n14361), 
        .B2(n12841), .ZN(n14369) );
  NAND2_X1 U15135 ( .A1(n12844), .A2(n12843), .ZN(n12845) );
  NAND2_X1 U15136 ( .A1(n12818), .A2(n12845), .ZN(n12846) );
  XNOR2_X1 U15137 ( .A(n14344), .B(n12845), .ZN(n14346) );
  NAND2_X1 U15138 ( .A1(P3_REG1_REG_15__SCAN_IN), .A2(n14346), .ZN(n14345) );
  NAND2_X1 U15139 ( .A1(n12848), .A2(n12849), .ZN(n12850) );
  NAND2_X1 U15140 ( .A1(P3_REG1_REG_17__SCAN_IN), .A2(n14381), .ZN(n14380) );
  NAND2_X1 U15141 ( .A1(n12850), .A2(n14380), .ZN(n14396) );
  NAND2_X1 U15142 ( .A1(n14397), .A2(n14396), .ZN(n14395) );
  OAI21_X1 U15143 ( .B1(n14394), .B2(n13160), .A(n14395), .ZN(n12852) );
  XNOR2_X1 U15144 ( .A(n12852), .B(n12851), .ZN(n12854) );
  NAND2_X1 U15145 ( .A1(n15094), .A2(P3_ADDR_REG_19__SCAN_IN), .ZN(n12855) );
  OAI211_X1 U15146 ( .C1(n15088), .C2(n12857), .A(n12856), .B(n12855), .ZN(
        n12858) );
  NOR2_X1 U15147 ( .A1(n12861), .A2(n12860), .ZN(n13182) );
  NOR2_X1 U15148 ( .A1(n15108), .A2(n12862), .ZN(n12868) );
  AOI21_X1 U15149 ( .B1(n13182), .B2(n13106), .A(n12868), .ZN(n12865) );
  NAND2_X1 U15150 ( .A1(n13116), .A2(P3_REG2_REG_31__SCAN_IN), .ZN(n12863) );
  OAI211_X1 U15151 ( .C1(n13184), .C2(n13094), .A(n12865), .B(n12863), .ZN(
        P3_U3202) );
  NAND2_X1 U15152 ( .A1(n13116), .A2(P3_REG2_REG_30__SCAN_IN), .ZN(n12864) );
  OAI211_X1 U15153 ( .C1(n12866), .C2(n13094), .A(n12865), .B(n12864), .ZN(
        P3_U3203) );
  INV_X1 U15154 ( .A(n12867), .ZN(n12874) );
  AOI21_X1 U15155 ( .B1(n13116), .B2(P3_REG2_REG_29__SCAN_IN), .A(n12868), 
        .ZN(n12869) );
  OAI21_X1 U15156 ( .B1(n12870), .B2(n13094), .A(n12869), .ZN(n12871) );
  AOI21_X1 U15157 ( .B1(n12872), .B2(n13113), .A(n12871), .ZN(n12873) );
  OAI21_X1 U15158 ( .B1(n12874), .B2(n13116), .A(n12873), .ZN(P3_U3204) );
  INV_X1 U15159 ( .A(P3_REG2_REG_28__SCAN_IN), .ZN(n12877) );
  INV_X1 U15160 ( .A(n12875), .ZN(n12876) );
  OAI22_X1 U15161 ( .A1(n13106), .A2(n12877), .B1(n12876), .B2(n15108), .ZN(
        n12878) );
  AOI21_X1 U15162 ( .B1(n7954), .B2(n13108), .A(n12878), .ZN(n12881) );
  NAND2_X1 U15163 ( .A1(n12879), .A2(n13113), .ZN(n12880) );
  OAI211_X1 U15164 ( .C1(n12882), .C2(n13116), .A(n12881), .B(n12880), .ZN(
        P3_U3205) );
  INV_X1 U15165 ( .A(n13106), .ZN(n13043) );
  AOI22_X1 U15166 ( .A1(n13043), .A2(P3_REG2_REG_27__SCAN_IN), .B1(n13092), 
        .B2(n12883), .ZN(n12884) );
  OAI21_X1 U15167 ( .B1(n12885), .B2(n13094), .A(n12884), .ZN(n12886) );
  AOI21_X1 U15168 ( .B1(n12887), .B2(n12926), .A(n12886), .ZN(n12888) );
  OAI21_X1 U15169 ( .B1(n6558), .B2(n13116), .A(n12888), .ZN(P3_U3206) );
  XNOR2_X1 U15170 ( .A(n12889), .B(n12893), .ZN(n12891) );
  OAI21_X1 U15171 ( .B1(n12891), .B2(n15115), .A(n12890), .ZN(n13121) );
  INV_X1 U15172 ( .A(n13121), .ZN(n12898) );
  XOR2_X1 U15173 ( .A(n12892), .B(n12893), .Z(n13122) );
  AOI22_X1 U15174 ( .A1(n13043), .A2(P3_REG2_REG_26__SCAN_IN), .B1(n13092), 
        .B2(n12894), .ZN(n12895) );
  OAI21_X1 U15175 ( .B1(n13193), .B2(n13094), .A(n12895), .ZN(n12896) );
  AOI21_X1 U15176 ( .B1(n13122), .B2(n13113), .A(n12896), .ZN(n12897) );
  OAI21_X1 U15177 ( .B1(n13116), .B2(n12898), .A(n12897), .ZN(P3_U3207) );
  XNOR2_X1 U15178 ( .A(n12899), .B(n12901), .ZN(n12905) );
  OAI211_X1 U15179 ( .C1(n12902), .C2(n12901), .A(n12900), .B(n13103), .ZN(
        n12903) );
  OAI211_X1 U15180 ( .C1(n12905), .C2(n12920), .A(n12904), .B(n12903), .ZN(
        n13125) );
  INV_X1 U15181 ( .A(n13125), .ZN(n12910) );
  INV_X1 U15182 ( .A(n12905), .ZN(n13126) );
  AOI22_X1 U15183 ( .A1(n13043), .A2(P3_REG2_REG_25__SCAN_IN), .B1(n13092), 
        .B2(n12906), .ZN(n12907) );
  OAI21_X1 U15184 ( .B1(n13197), .B2(n13094), .A(n12907), .ZN(n12908) );
  AOI21_X1 U15185 ( .B1(n13126), .B2(n12926), .A(n12908), .ZN(n12909) );
  OAI21_X1 U15186 ( .B1(n12910), .B2(n13116), .A(n12909), .ZN(P3_U3208) );
  INV_X1 U15187 ( .A(n12911), .ZN(n12912) );
  AOI21_X1 U15188 ( .B1(n12916), .B2(n12913), .A(n12912), .ZN(n12921) );
  INV_X1 U15189 ( .A(n12914), .ZN(n12919) );
  OAI211_X1 U15190 ( .C1(n12917), .C2(n12916), .A(n12915), .B(n13103), .ZN(
        n12918) );
  OAI211_X1 U15191 ( .C1(n12921), .C2(n12920), .A(n12919), .B(n12918), .ZN(
        n13129) );
  INV_X1 U15192 ( .A(n13129), .ZN(n12928) );
  INV_X1 U15193 ( .A(n12921), .ZN(n13130) );
  INV_X1 U15194 ( .A(n12922), .ZN(n13201) );
  AOI22_X1 U15195 ( .A1(n13043), .A2(P3_REG2_REG_24__SCAN_IN), .B1(n13092), 
        .B2(n12923), .ZN(n12924) );
  OAI21_X1 U15196 ( .B1(n13201), .B2(n13094), .A(n12924), .ZN(n12925) );
  AOI21_X1 U15197 ( .B1(n13130), .B2(n12926), .A(n12925), .ZN(n12927) );
  OAI21_X1 U15198 ( .B1(n12928), .B2(n13116), .A(n12927), .ZN(P3_U3209) );
  OAI21_X1 U15199 ( .B1(n12931), .B2(n12930), .A(n12929), .ZN(n13136) );
  OR2_X1 U15200 ( .A1(n12972), .A2(n12932), .ZN(n12934) );
  NAND2_X1 U15201 ( .A1(n12934), .A2(n12933), .ZN(n12937) );
  OAI211_X1 U15202 ( .C1(n12937), .C2(n12936), .A(n13103), .B(n12935), .ZN(
        n12939) );
  NAND2_X1 U15203 ( .A1(n12939), .A2(n12938), .ZN(n13133) );
  AOI22_X1 U15204 ( .A1(n13043), .A2(P3_REG2_REG_23__SCAN_IN), .B1(n13092), 
        .B2(n12940), .ZN(n12941) );
  OAI21_X1 U15205 ( .B1(n12942), .B2(n13094), .A(n12941), .ZN(n12943) );
  AOI21_X1 U15206 ( .B1(n13133), .B2(n13106), .A(n12943), .ZN(n12944) );
  OAI21_X1 U15207 ( .B1(n13084), .B2(n13136), .A(n12944), .ZN(P3_U3210) );
  XNOR2_X1 U15208 ( .A(n12945), .B(n12949), .ZN(n13138) );
  INV_X1 U15209 ( .A(n13138), .ZN(n12959) );
  OR2_X1 U15210 ( .A1(n12972), .A2(n12946), .ZN(n12948) );
  NAND2_X1 U15211 ( .A1(n12948), .A2(n12947), .ZN(n12950) );
  XNOR2_X1 U15212 ( .A(n12950), .B(n12949), .ZN(n12953) );
  INV_X1 U15213 ( .A(n12951), .ZN(n12952) );
  OAI21_X1 U15214 ( .B1(n12953), .B2(n15115), .A(n12952), .ZN(n13137) );
  INV_X1 U15215 ( .A(n12954), .ZN(n13206) );
  AOI22_X1 U15216 ( .A1(n12955), .A2(n13092), .B1(n13043), .B2(
        P3_REG2_REG_22__SCAN_IN), .ZN(n12956) );
  OAI21_X1 U15217 ( .B1(n13206), .B2(n13094), .A(n12956), .ZN(n12957) );
  AOI21_X1 U15218 ( .B1(n13137), .B2(n13106), .A(n12957), .ZN(n12958) );
  OAI21_X1 U15219 ( .B1(n12959), .B2(n13084), .A(n12958), .ZN(P3_U3211) );
  XNOR2_X1 U15220 ( .A(n12960), .B(n12962), .ZN(n13142) );
  INV_X1 U15221 ( .A(n13142), .ZN(n12970) );
  NAND2_X1 U15222 ( .A1(n12975), .A2(n12961), .ZN(n12963) );
  XNOR2_X1 U15223 ( .A(n12963), .B(n12962), .ZN(n12965) );
  OAI21_X1 U15224 ( .B1(n12965), .B2(n15115), .A(n12964), .ZN(n13141) );
  AOI22_X1 U15225 ( .A1(n12966), .A2(n13092), .B1(n13043), .B2(
        P3_REG2_REG_21__SCAN_IN), .ZN(n12967) );
  OAI21_X1 U15226 ( .B1(n13210), .B2(n13094), .A(n12967), .ZN(n12968) );
  AOI21_X1 U15227 ( .B1(n13141), .B2(n13106), .A(n12968), .ZN(n12969) );
  OAI21_X1 U15228 ( .B1(n12970), .B2(n13084), .A(n12969), .ZN(P3_U3212) );
  AOI21_X1 U15229 ( .B1(n12972), .B2(n12971), .A(n15115), .ZN(n12976) );
  OAI22_X1 U15230 ( .A1(n12973), .A2(n15111), .B1(n13003), .B2(n15109), .ZN(
        n12974) );
  AOI21_X1 U15231 ( .B1(n12976), .B2(n12975), .A(n12974), .ZN(n13148) );
  INV_X1 U15232 ( .A(n12977), .ZN(n12979) );
  INV_X1 U15233 ( .A(P3_REG2_REG_20__SCAN_IN), .ZN(n12978) );
  OAI22_X1 U15234 ( .A1(n12979), .A2(n15108), .B1(n12978), .B2(n13106), .ZN(
        n12980) );
  AOI21_X1 U15235 ( .B1(n13145), .B2(n13108), .A(n12980), .ZN(n12984) );
  NAND2_X1 U15236 ( .A1(n12981), .A2(n12982), .ZN(n13146) );
  NAND3_X1 U15237 ( .A1(n13147), .A2(n13146), .A3(n13113), .ZN(n12983) );
  OAI211_X1 U15238 ( .C1(n13148), .C2(n13116), .A(n12984), .B(n12983), .ZN(
        P3_U3213) );
  NAND2_X1 U15239 ( .A1(n13158), .A2(n12985), .ZN(n12986) );
  XNOR2_X1 U15240 ( .A(n12986), .B(n12988), .ZN(n13153) );
  INV_X1 U15241 ( .A(n13153), .ZN(n12996) );
  XOR2_X1 U15242 ( .A(n12988), .B(n12987), .Z(n12989) );
  OAI222_X1 U15243 ( .A1(n15111), .A2(n12990), .B1(n15109), .B2(n13018), .C1(
        n12989), .C2(n15115), .ZN(n13152) );
  INV_X1 U15244 ( .A(n12991), .ZN(n13218) );
  AOI22_X1 U15245 ( .A1(n13043), .A2(P3_REG2_REG_19__SCAN_IN), .B1(n13092), 
        .B2(n12992), .ZN(n12993) );
  OAI21_X1 U15246 ( .B1(n13218), .B2(n13094), .A(n12993), .ZN(n12994) );
  AOI21_X1 U15247 ( .B1(n13152), .B2(n13106), .A(n12994), .ZN(n12995) );
  OAI21_X1 U15248 ( .B1(n13084), .B2(n12996), .A(n12995), .ZN(P3_U3214) );
  INV_X1 U15249 ( .A(n12997), .ZN(n12998) );
  AOI21_X1 U15250 ( .B1(n13000), .B2(n12999), .A(n12998), .ZN(n13001) );
  OAI222_X1 U15251 ( .A1(n15111), .A2(n13003), .B1(n15109), .B2(n13002), .C1(
        n15115), .C2(n13001), .ZN(n13157) );
  INV_X1 U15252 ( .A(n13004), .ZN(n13222) );
  AOI22_X1 U15253 ( .A1(n13043), .A2(P3_REG2_REG_18__SCAN_IN), .B1(n13092), 
        .B2(n13005), .ZN(n13006) );
  OAI21_X1 U15254 ( .B1(n13222), .B2(n13094), .A(n13006), .ZN(n13010) );
  INV_X1 U15255 ( .A(n13158), .ZN(n13008) );
  AND2_X1 U15256 ( .A1(n13007), .A2(n7893), .ZN(n13156) );
  NOR3_X1 U15257 ( .A1(n13008), .A2(n13156), .A3(n13084), .ZN(n13009) );
  AOI211_X1 U15258 ( .C1(n13157), .C2(n13106), .A(n13010), .B(n13009), .ZN(
        n13011) );
  INV_X1 U15259 ( .A(n13011), .ZN(P3_U3215) );
  XNOR2_X1 U15260 ( .A(n13012), .B(n13013), .ZN(n13163) );
  INV_X1 U15261 ( .A(n13163), .ZN(n13023) );
  XNOR2_X1 U15262 ( .A(n13014), .B(n13015), .ZN(n13016) );
  OAI222_X1 U15263 ( .A1(n15111), .A2(n13018), .B1(n15109), .B2(n13017), .C1(
        n13016), .C2(n15115), .ZN(n13162) );
  AOI22_X1 U15264 ( .A1(n13043), .A2(P3_REG2_REG_17__SCAN_IN), .B1(n13092), 
        .B2(n13019), .ZN(n13020) );
  OAI21_X1 U15265 ( .B1(n13226), .B2(n13094), .A(n13020), .ZN(n13021) );
  AOI21_X1 U15266 ( .B1(n13162), .B2(n13106), .A(n13021), .ZN(n13022) );
  OAI21_X1 U15267 ( .B1(n13084), .B2(n13023), .A(n13022), .ZN(P3_U3216) );
  NAND2_X1 U15268 ( .A1(n13036), .A2(n13038), .ZN(n13025) );
  NAND2_X1 U15269 ( .A1(n13025), .A2(n13024), .ZN(n13026) );
  XOR2_X1 U15270 ( .A(n13027), .B(n13026), .Z(n13169) );
  XNOR2_X1 U15271 ( .A(n13028), .B(n13027), .ZN(n13030) );
  OAI21_X1 U15272 ( .B1(n13030), .B2(n15115), .A(n13029), .ZN(n13166) );
  INV_X1 U15273 ( .A(n13167), .ZN(n13033) );
  AOI22_X1 U15274 ( .A1(n13043), .A2(P3_REG2_REG_16__SCAN_IN), .B1(n13092), 
        .B2(n13031), .ZN(n13032) );
  OAI21_X1 U15275 ( .B1(n13033), .B2(n13094), .A(n13032), .ZN(n13034) );
  AOI21_X1 U15276 ( .B1(n13166), .B2(n13106), .A(n13034), .ZN(n13035) );
  OAI21_X1 U15277 ( .B1(n13169), .B2(n13084), .A(n13035), .ZN(P3_U3217) );
  XNOR2_X1 U15278 ( .A(n13036), .B(n13038), .ZN(n13171) );
  INV_X1 U15279 ( .A(n13171), .ZN(n13047) );
  XOR2_X1 U15280 ( .A(n13038), .B(n13037), .Z(n13041) );
  INV_X1 U15281 ( .A(n13039), .ZN(n13040) );
  OAI21_X1 U15282 ( .B1(n13041), .B2(n15115), .A(n13040), .ZN(n13170) );
  AOI22_X1 U15283 ( .A1(n13043), .A2(P3_REG2_REG_15__SCAN_IN), .B1(n13092), 
        .B2(n13042), .ZN(n13044) );
  OAI21_X1 U15284 ( .B1(n13231), .B2(n13094), .A(n13044), .ZN(n13045) );
  AOI21_X1 U15285 ( .B1(n13170), .B2(n13106), .A(n13045), .ZN(n13046) );
  OAI21_X1 U15286 ( .B1(n13047), .B2(n13084), .A(n13046), .ZN(P3_U3218) );
  XNOR2_X1 U15287 ( .A(n13048), .B(n13049), .ZN(n13052) );
  AOI222_X1 U15288 ( .A1(n13103), .A2(n13052), .B1(n13051), .B2(n13100), .C1(
        n13050), .C2(n13098), .ZN(n14412) );
  INV_X1 U15289 ( .A(n14413), .ZN(n13057) );
  INV_X1 U15290 ( .A(P3_REG2_REG_14__SCAN_IN), .ZN(n13055) );
  INV_X1 U15291 ( .A(n13053), .ZN(n13054) );
  OAI22_X1 U15292 ( .A1(n13106), .A2(n13055), .B1(n13054), .B2(n15108), .ZN(
        n13056) );
  AOI21_X1 U15293 ( .B1(n13057), .B2(n13108), .A(n13056), .ZN(n13061) );
  XNOR2_X1 U15294 ( .A(n13059), .B(n13058), .ZN(n14415) );
  NAND2_X1 U15295 ( .A1(n14415), .A2(n13113), .ZN(n13060) );
  OAI211_X1 U15296 ( .C1(n14412), .C2(n13116), .A(n13061), .B(n13060), .ZN(
        P3_U3219) );
  XOR2_X1 U15297 ( .A(n13062), .B(n13070), .Z(n13064) );
  AOI222_X1 U15298 ( .A1(n13103), .A2(n13064), .B1(n13063), .B2(n13100), .C1(
        n13087), .C2(n13098), .ZN(n14416) );
  INV_X1 U15299 ( .A(n14417), .ZN(n13069) );
  INV_X1 U15300 ( .A(n13065), .ZN(n13066) );
  OAI22_X1 U15301 ( .A1(n13106), .A2(n13067), .B1(n13066), .B2(n15108), .ZN(
        n13068) );
  AOI21_X1 U15302 ( .B1(n13069), .B2(n13108), .A(n13068), .ZN(n13073) );
  XOR2_X1 U15303 ( .A(n13071), .B(n13070), .Z(n14419) );
  NAND2_X1 U15304 ( .A1(n14419), .A2(n13113), .ZN(n13072) );
  OAI211_X1 U15305 ( .C1(n14416), .C2(n13116), .A(n13073), .B(n13072), .ZN(
        P3_U3220) );
  XNOR2_X1 U15306 ( .A(n13074), .B(n13076), .ZN(n14422) );
  XNOR2_X1 U15307 ( .A(n13075), .B(n13076), .ZN(n13078) );
  OAI21_X1 U15308 ( .B1(n13078), .B2(n15115), .A(n13077), .ZN(n14424) );
  INV_X1 U15309 ( .A(n14425), .ZN(n13081) );
  AOI22_X1 U15310 ( .A1(n13116), .A2(P3_REG2_REG_12__SCAN_IN), .B1(n13092), 
        .B2(n13079), .ZN(n13080) );
  OAI21_X1 U15311 ( .B1(n13081), .B2(n13094), .A(n13080), .ZN(n13082) );
  AOI21_X1 U15312 ( .B1(n14424), .B2(n13106), .A(n13082), .ZN(n13083) );
  OAI21_X1 U15313 ( .B1(n14422), .B2(n13084), .A(n13083), .ZN(P3_U3221) );
  XNOR2_X1 U15314 ( .A(n13085), .B(n7587), .ZN(n13088) );
  AOI222_X1 U15315 ( .A1(n13103), .A2(n13088), .B1(n13087), .B2(n13100), .C1(
        n13086), .C2(n13098), .ZN(n14427) );
  OAI21_X1 U15316 ( .B1(n13090), .B2(n7587), .A(n13089), .ZN(n14430) );
  AOI22_X1 U15317 ( .A1(n13116), .A2(P3_REG2_REG_11__SCAN_IN), .B1(n13092), 
        .B2(n13091), .ZN(n13093) );
  OAI21_X1 U15318 ( .B1(n14428), .B2(n13094), .A(n13093), .ZN(n13095) );
  AOI21_X1 U15319 ( .B1(n14430), .B2(n13113), .A(n13095), .ZN(n13096) );
  OAI21_X1 U15320 ( .B1(n14427), .B2(n13116), .A(n13096), .ZN(P3_U3222) );
  XNOR2_X1 U15321 ( .A(n13097), .B(n7573), .ZN(n13102) );
  AOI222_X1 U15322 ( .A1(n13103), .A2(n13102), .B1(n13101), .B2(n13100), .C1(
        n13099), .C2(n13098), .ZN(n13177) );
  INV_X1 U15323 ( .A(n13104), .ZN(n13105) );
  OAI22_X1 U15324 ( .A1(n13106), .A2(n10696), .B1(n13105), .B2(n15108), .ZN(
        n13107) );
  AOI21_X1 U15325 ( .B1(n13109), .B2(n13108), .A(n13107), .ZN(n13115) );
  NAND2_X1 U15326 ( .A1(n13111), .A2(n13112), .ZN(n13174) );
  NAND3_X1 U15327 ( .A1(n13175), .A2(n13174), .A3(n13113), .ZN(n13114) );
  OAI211_X1 U15328 ( .C1(n13177), .C2(n13116), .A(n13115), .B(n13114), .ZN(
        P3_U3223) );
  NAND2_X1 U15329 ( .A1(n15190), .A2(P3_REG1_REG_31__SCAN_IN), .ZN(n13117) );
  NAND2_X1 U15330 ( .A1(n13182), .A2(n15193), .ZN(n13118) );
  OAI211_X1 U15331 ( .C1(n13184), .C2(n13179), .A(n13117), .B(n13118), .ZN(
        P3_U3490) );
  INV_X1 U15332 ( .A(P3_REG1_REG_30__SCAN_IN), .ZN(n13120) );
  NAND2_X1 U15333 ( .A1(n13186), .A2(n8900), .ZN(n13119) );
  OAI211_X1 U15334 ( .C1(n15193), .C2(n13120), .A(n13119), .B(n13118), .ZN(
        P3_U3489) );
  INV_X1 U15335 ( .A(P3_REG1_REG_26__SCAN_IN), .ZN(n13123) );
  AOI21_X1 U15336 ( .B1(n13122), .B2(n15167), .A(n13121), .ZN(n13190) );
  MUX2_X1 U15337 ( .A(n13123), .B(n13190), .S(n15193), .Z(n13124) );
  OAI21_X1 U15338 ( .B1(n13193), .B2(n13179), .A(n13124), .ZN(P3_U3485) );
  INV_X1 U15339 ( .A(P3_REG1_REG_25__SCAN_IN), .ZN(n13127) );
  AOI21_X1 U15340 ( .B1(n15161), .B2(n13126), .A(n13125), .ZN(n13194) );
  MUX2_X1 U15341 ( .A(n13127), .B(n13194), .S(n15193), .Z(n13128) );
  OAI21_X1 U15342 ( .B1(n13197), .B2(n13179), .A(n13128), .ZN(P3_U3484) );
  INV_X1 U15343 ( .A(P3_REG1_REG_24__SCAN_IN), .ZN(n13131) );
  AOI21_X1 U15344 ( .B1(n15161), .B2(n13130), .A(n13129), .ZN(n13198) );
  MUX2_X1 U15345 ( .A(n13131), .B(n13198), .S(n15193), .Z(n13132) );
  OAI21_X1 U15346 ( .B1(n13201), .B2(n13179), .A(n13132), .ZN(P3_U3483) );
  INV_X1 U15347 ( .A(n15167), .ZN(n14421) );
  AOI21_X1 U15348 ( .B1(n15152), .B2(n13134), .A(n13133), .ZN(n13135) );
  OAI21_X1 U15349 ( .B1(n14421), .B2(n13136), .A(n13135), .ZN(n13202) );
  MUX2_X1 U15350 ( .A(P3_REG1_REG_23__SCAN_IN), .B(n13202), .S(n15193), .Z(
        P3_U3482) );
  INV_X1 U15351 ( .A(P3_REG1_REG_22__SCAN_IN), .ZN(n13139) );
  AOI21_X1 U15352 ( .B1(n15167), .B2(n13138), .A(n13137), .ZN(n13203) );
  MUX2_X1 U15353 ( .A(n13139), .B(n13203), .S(n15193), .Z(n13140) );
  OAI21_X1 U15354 ( .B1(n13206), .B2(n13179), .A(n13140), .ZN(P3_U3481) );
  INV_X1 U15355 ( .A(P3_REG1_REG_21__SCAN_IN), .ZN(n13143) );
  AOI21_X1 U15356 ( .B1(n13142), .B2(n15167), .A(n13141), .ZN(n13207) );
  MUX2_X1 U15357 ( .A(n13143), .B(n13207), .S(n15193), .Z(n13144) );
  OAI21_X1 U15358 ( .B1(n13210), .B2(n13179), .A(n13144), .ZN(P3_U3480) );
  INV_X1 U15359 ( .A(n13145), .ZN(n13214) );
  NAND3_X1 U15360 ( .A1(n13147), .A2(n13146), .A3(n15167), .ZN(n13149) );
  AND2_X1 U15361 ( .A1(n13149), .A2(n13148), .ZN(n13212) );
  INV_X1 U15362 ( .A(P3_REG1_REG_20__SCAN_IN), .ZN(n13150) );
  MUX2_X1 U15363 ( .A(n13212), .B(n13150), .S(n15190), .Z(n13151) );
  OAI21_X1 U15364 ( .B1(n13214), .B2(n13179), .A(n13151), .ZN(P3_U3479) );
  INV_X1 U15365 ( .A(P3_REG1_REG_19__SCAN_IN), .ZN(n13154) );
  AOI21_X1 U15366 ( .B1(n13153), .B2(n15167), .A(n13152), .ZN(n13215) );
  MUX2_X1 U15367 ( .A(n13154), .B(n13215), .S(n15193), .Z(n13155) );
  OAI21_X1 U15368 ( .B1(n13218), .B2(n13179), .A(n13155), .ZN(P3_U3478) );
  NOR2_X1 U15369 ( .A1(n13156), .A2(n14421), .ZN(n13159) );
  AOI21_X1 U15370 ( .B1(n13159), .B2(n13158), .A(n13157), .ZN(n13219) );
  MUX2_X1 U15371 ( .A(n13160), .B(n13219), .S(n15193), .Z(n13161) );
  OAI21_X1 U15372 ( .B1(n13222), .B2(n13179), .A(n13161), .ZN(P3_U3477) );
  INV_X1 U15373 ( .A(P3_REG1_REG_17__SCAN_IN), .ZN(n13164) );
  AOI21_X1 U15374 ( .B1(n13163), .B2(n15167), .A(n13162), .ZN(n13223) );
  MUX2_X1 U15375 ( .A(n13164), .B(n13223), .S(n15193), .Z(n13165) );
  OAI21_X1 U15376 ( .B1(n13179), .B2(n13226), .A(n13165), .ZN(P3_U3476) );
  AOI21_X1 U15377 ( .B1(n15152), .B2(n13167), .A(n13166), .ZN(n13168) );
  OAI21_X1 U15378 ( .B1(n13169), .B2(n14421), .A(n13168), .ZN(n13227) );
  MUX2_X1 U15379 ( .A(P3_REG1_REG_16__SCAN_IN), .B(n13227), .S(n15193), .Z(
        P3_U3475) );
  INV_X1 U15380 ( .A(P3_REG1_REG_15__SCAN_IN), .ZN(n13172) );
  AOI21_X1 U15381 ( .B1(n13171), .B2(n15167), .A(n13170), .ZN(n13228) );
  MUX2_X1 U15382 ( .A(n13172), .B(n13228), .S(n15193), .Z(n13173) );
  OAI21_X1 U15383 ( .B1(n13179), .B2(n13231), .A(n13173), .ZN(P3_U3474) );
  NAND3_X1 U15384 ( .A1(n13175), .A2(n13174), .A3(n15167), .ZN(n13176) );
  NAND2_X1 U15385 ( .A1(n13177), .A2(n13176), .ZN(n13236) );
  OAI22_X1 U15386 ( .A1(n13179), .A2(n13233), .B1(n15193), .B2(n13178), .ZN(
        n13180) );
  AOI21_X1 U15387 ( .B1(n13236), .B2(n15193), .A(n13180), .ZN(n13181) );
  INV_X1 U15388 ( .A(n13181), .ZN(P3_U3469) );
  NAND2_X1 U15389 ( .A1(n15175), .A2(P3_REG0_REG_31__SCAN_IN), .ZN(n13183) );
  NAND2_X1 U15390 ( .A1(n13182), .A2(n15177), .ZN(n13187) );
  OAI211_X1 U15391 ( .C1(n13184), .C2(n13234), .A(n13183), .B(n13187), .ZN(
        P3_U3458) );
  INV_X1 U15392 ( .A(P3_REG0_REG_30__SCAN_IN), .ZN(n13189) );
  NAND2_X1 U15393 ( .A1(n13186), .A2(n13185), .ZN(n13188) );
  OAI211_X1 U15394 ( .C1(n15177), .C2(n13189), .A(n13188), .B(n13187), .ZN(
        P3_U3457) );
  INV_X1 U15395 ( .A(P3_REG0_REG_26__SCAN_IN), .ZN(n13191) );
  MUX2_X1 U15396 ( .A(n13191), .B(n13190), .S(n15177), .Z(n13192) );
  OAI21_X1 U15397 ( .B1(n13193), .B2(n13234), .A(n13192), .ZN(P3_U3453) );
  INV_X1 U15398 ( .A(P3_REG0_REG_25__SCAN_IN), .ZN(n13195) );
  MUX2_X1 U15399 ( .A(n13195), .B(n13194), .S(n15177), .Z(n13196) );
  OAI21_X1 U15400 ( .B1(n13197), .B2(n13234), .A(n13196), .ZN(P3_U3452) );
  INV_X1 U15401 ( .A(P3_REG0_REG_24__SCAN_IN), .ZN(n13199) );
  MUX2_X1 U15402 ( .A(n13199), .B(n13198), .S(n15177), .Z(n13200) );
  OAI21_X1 U15403 ( .B1(n13201), .B2(n13234), .A(n13200), .ZN(P3_U3451) );
  MUX2_X1 U15404 ( .A(P3_REG0_REG_23__SCAN_IN), .B(n13202), .S(n15177), .Z(
        P3_U3450) );
  INV_X1 U15405 ( .A(P3_REG0_REG_22__SCAN_IN), .ZN(n13204) );
  MUX2_X1 U15406 ( .A(n13204), .B(n13203), .S(n15177), .Z(n13205) );
  OAI21_X1 U15407 ( .B1(n13206), .B2(n13234), .A(n13205), .ZN(P3_U3449) );
  MUX2_X1 U15408 ( .A(n13208), .B(n13207), .S(n15177), .Z(n13209) );
  OAI21_X1 U15409 ( .B1(n13210), .B2(n13234), .A(n13209), .ZN(P3_U3448) );
  MUX2_X1 U15410 ( .A(n13212), .B(n13211), .S(n15175), .Z(n13213) );
  OAI21_X1 U15411 ( .B1(n13214), .B2(n13234), .A(n13213), .ZN(P3_U3447) );
  MUX2_X1 U15412 ( .A(n13216), .B(n13215), .S(n15177), .Z(n13217) );
  OAI21_X1 U15413 ( .B1(n13218), .B2(n13234), .A(n13217), .ZN(P3_U3446) );
  INV_X1 U15414 ( .A(P3_REG0_REG_18__SCAN_IN), .ZN(n13220) );
  MUX2_X1 U15415 ( .A(n13220), .B(n13219), .S(n15177), .Z(n13221) );
  OAI21_X1 U15416 ( .B1(n13222), .B2(n13234), .A(n13221), .ZN(P3_U3444) );
  INV_X1 U15417 ( .A(P3_REG0_REG_17__SCAN_IN), .ZN(n13224) );
  MUX2_X1 U15418 ( .A(n13224), .B(n13223), .S(n15177), .Z(n13225) );
  OAI21_X1 U15419 ( .B1(n13234), .B2(n13226), .A(n13225), .ZN(P3_U3441) );
  MUX2_X1 U15420 ( .A(P3_REG0_REG_16__SCAN_IN), .B(n13227), .S(n15177), .Z(
        P3_U3438) );
  INV_X1 U15421 ( .A(P3_REG0_REG_15__SCAN_IN), .ZN(n13229) );
  MUX2_X1 U15422 ( .A(n13229), .B(n13228), .S(n15177), .Z(n13230) );
  OAI21_X1 U15423 ( .B1(n13234), .B2(n13231), .A(n13230), .ZN(P3_U3435) );
  INV_X1 U15424 ( .A(P3_REG0_REG_10__SCAN_IN), .ZN(n13232) );
  OAI22_X1 U15425 ( .A1(n13234), .A2(n13233), .B1(n15177), .B2(n13232), .ZN(
        n13235) );
  AOI21_X1 U15426 ( .B1(n13236), .B2(n15177), .A(n13235), .ZN(n13237) );
  INV_X1 U15427 ( .A(n13237), .ZN(P3_U3420) );
  MUX2_X1 U15428 ( .A(n13239), .B(P3_D_REG_0__SCAN_IN), .S(n13238), .Z(
        P3_U3376) );
  NAND2_X1 U15429 ( .A1(n13240), .A2(n14317), .ZN(n13244) );
  OR4_X1 U15430 ( .A1(n13242), .A2(P3_IR_REG_30__SCAN_IN), .A3(P3_U3151), .A4(
        n13241), .ZN(n13243) );
  OAI211_X1 U15431 ( .C1(n13245), .C2(n13247), .A(n13244), .B(n13243), .ZN(
        P3_U3264) );
  INV_X1 U15432 ( .A(n13246), .ZN(n13249) );
  OAI222_X1 U15433 ( .A1(n13250), .A2(n13249), .B1(P3_U3151), .B2(n7915), .C1(
        n13248), .C2(n13247), .ZN(P3_U3267) );
  MUX2_X1 U15434 ( .A(n13251), .B(P3_IR_REG_0__SCAN_IN), .S(
        P3_STATE_REG_SCAN_IN), .Z(P3_U3295) );
  AOI21_X1 U15435 ( .B1(n13253), .B2(n13252), .A(n13334), .ZN(n13258) );
  AOI22_X1 U15436 ( .A1(n13375), .A2(n13642), .B1(n13640), .B2(n13377), .ZN(
        n13520) );
  NAND2_X1 U15437 ( .A1(n13711), .A2(n9820), .ZN(n13255) );
  AOI22_X1 U15438 ( .A1(n13524), .A2(n13368), .B1(P2_REG3_REG_27__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13254) );
  OAI211_X1 U15439 ( .C1(n13520), .C2(n13366), .A(n13255), .B(n13254), .ZN(
        n13256) );
  AOI21_X1 U15440 ( .B1(n13258), .B2(n13257), .A(n13256), .ZN(n13259) );
  INV_X1 U15441 ( .A(n13259), .ZN(P2_U3186) );
  AOI22_X1 U15442 ( .A1(n13261), .A2(n13359), .B1(n13347), .B2(n13380), .ZN(
        n13266) );
  NAND2_X1 U15443 ( .A1(n13261), .A2(n13260), .ZN(n13336) );
  INV_X1 U15444 ( .A(n13336), .ZN(n13265) );
  OAI22_X1 U15445 ( .A1(n13304), .A2(n13657), .B1(n13292), .B2(n13655), .ZN(
        n13580) );
  AOI22_X1 U15446 ( .A1(n13580), .A2(n13308), .B1(P2_REG3_REG_23__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13262) );
  OAI21_X1 U15447 ( .B1(n13586), .B2(n13352), .A(n13262), .ZN(n13263) );
  AOI21_X1 U15448 ( .B1(n13735), .B2(n9820), .A(n13263), .ZN(n13264) );
  OAI21_X1 U15449 ( .B1(n13266), .B2(n13265), .A(n13264), .ZN(P2_U3188) );
  OAI211_X1 U15450 ( .C1(n13269), .C2(n13268), .A(n13267), .B(n13359), .ZN(
        n13274) );
  AOI22_X1 U15451 ( .A1(n13308), .A2(n13271), .B1(n9820), .B2(n13270), .ZN(
        n13273) );
  MUX2_X1 U15452 ( .A(n13352), .B(P2_STATE_REG_SCAN_IN), .S(
        P2_REG3_REG_3__SCAN_IN), .Z(n13272) );
  NAND3_X1 U15453 ( .A1(n13274), .A2(n13273), .A3(n13272), .ZN(P2_U3190) );
  INV_X1 U15454 ( .A(n13277), .ZN(n13278) );
  AOI21_X1 U15455 ( .B1(n13283), .B2(n13276), .A(n13278), .ZN(n13288) );
  INV_X1 U15456 ( .A(n13279), .ZN(n13664) );
  NAND2_X1 U15457 ( .A1(n13368), .A2(n13664), .ZN(n13280) );
  NAND2_X1 U15458 ( .A1(P2_U3088), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n13493)
         );
  OAI211_X1 U15459 ( .C1(n13351), .C2(n13658), .A(n13280), .B(n13493), .ZN(
        n13286) );
  INV_X1 U15460 ( .A(n13281), .ZN(n13282) );
  NAND3_X1 U15461 ( .A1(n13283), .A2(n13347), .A3(n13282), .ZN(n13284) );
  AOI21_X1 U15462 ( .B1(n13284), .B2(n13353), .A(n13656), .ZN(n13285) );
  AOI211_X1 U15463 ( .C1(n13757), .C2(n9820), .A(n13286), .B(n13285), .ZN(
        n13287) );
  OAI21_X1 U15464 ( .B1(n13288), .B2(n13334), .A(n13287), .ZN(P2_U3191) );
  OAI211_X1 U15465 ( .C1(n13291), .C2(n13290), .A(n13289), .B(n13359), .ZN(
        n13296) );
  OAI22_X1 U15466 ( .A1(n13353), .A2(n13658), .B1(n13352), .B2(n13618), .ZN(
        n13294) );
  NOR2_X1 U15467 ( .A1(n13292), .A2(n13351), .ZN(n13293) );
  AOI211_X1 U15468 ( .C1(P2_REG3_REG_21__SCAN_IN), .C2(P2_U3088), .A(n13294), 
        .B(n13293), .ZN(n13295) );
  OAI211_X1 U15469 ( .C1(n13621), .C2(n13371), .A(n13296), .B(n13295), .ZN(
        P2_U3195) );
  AND2_X1 U15470 ( .A1(n13298), .A2(n13297), .ZN(n13337) );
  INV_X1 U15471 ( .A(n13299), .ZN(n13300) );
  AOI21_X1 U15472 ( .B1(n13337), .B2(n13300), .A(n13334), .ZN(n13303) );
  NOR3_X1 U15473 ( .A1(n13301), .A2(n13304), .A3(n13327), .ZN(n13302) );
  OAI21_X1 U15474 ( .B1(n13303), .B2(n13302), .A(n12101), .ZN(n13310) );
  OAI22_X1 U15475 ( .A1(n13305), .A2(n13657), .B1(n13304), .B2(n13655), .ZN(
        n13544) );
  OAI22_X1 U15476 ( .A1(n13551), .A2(n13352), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13306), .ZN(n13307) );
  AOI21_X1 U15477 ( .B1(n13544), .B2(n13308), .A(n13307), .ZN(n13309) );
  OAI211_X1 U15478 ( .C1(n6955), .C2(n13371), .A(n13310), .B(n13309), .ZN(
        P2_U3197) );
  INV_X1 U15479 ( .A(n13311), .ZN(n13312) );
  AOI21_X1 U15480 ( .B1(n13314), .B2(n13313), .A(n13312), .ZN(n13322) );
  OAI21_X1 U15481 ( .B1(n13351), .B2(n13316), .A(n13315), .ZN(n13320) );
  OAI22_X1 U15482 ( .A1(n13353), .A2(n13318), .B1(n13352), .B2(n13317), .ZN(
        n13319) );
  AOI211_X1 U15483 ( .C1(n13772), .C2(n9820), .A(n13320), .B(n13319), .ZN(
        n13321) );
  OAI21_X1 U15484 ( .B1(n13322), .B2(n13334), .A(n13321), .ZN(P2_U3198) );
  OAI22_X1 U15485 ( .A1(n13351), .A2(n13656), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13323), .ZN(n13326) );
  OAI22_X1 U15486 ( .A1(n13353), .A2(n13328), .B1(n13352), .B2(n13324), .ZN(
        n13325) );
  AOI211_X1 U15487 ( .C1(n13767), .C2(n9820), .A(n13326), .B(n13325), .ZN(
        n13333) );
  OAI22_X1 U15488 ( .A1(n13329), .A2(n13334), .B1(n13328), .B2(n13327), .ZN(
        n13330) );
  NAND3_X1 U15489 ( .A1(n13311), .A2(n13331), .A3(n13330), .ZN(n13332) );
  OAI211_X1 U15490 ( .C1(n6630), .C2(n13334), .A(n13333), .B(n13332), .ZN(
        P2_U3200) );
  NAND2_X1 U15491 ( .A1(n13336), .A2(n13335), .ZN(n13338) );
  OAI211_X1 U15492 ( .C1(n13339), .C2(n13338), .A(n13337), .B(n13359), .ZN(
        n13344) );
  NOR2_X1 U15493 ( .A1(n13598), .A2(n13353), .ZN(n13342) );
  OAI22_X1 U15494 ( .A1(n7152), .A2(n13351), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13340), .ZN(n13341) );
  AOI211_X1 U15495 ( .C1(n13368), .C2(n13571), .A(n13342), .B(n13341), .ZN(
        n13343) );
  OAI211_X1 U15496 ( .C1(n6957), .C2(n13371), .A(n13344), .B(n13343), .ZN(
        P2_U3201) );
  XNOR2_X1 U15497 ( .A(n13346), .B(n13345), .ZN(n13348) );
  AOI22_X1 U15498 ( .A1(n13348), .A2(n13359), .B1(n13347), .B2(n13625), .ZN(
        n13358) );
  INV_X1 U15499 ( .A(n13349), .ZN(n13357) );
  OAI22_X1 U15500 ( .A1(n13598), .A2(n13351), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13350), .ZN(n13355) );
  OAI22_X1 U15501 ( .A1(n13353), .A2(n13597), .B1(n13352), .B2(n13608), .ZN(
        n13354) );
  AOI211_X1 U15502 ( .C1(n13740), .C2(n9820), .A(n13355), .B(n13354), .ZN(
        n13356) );
  OAI21_X1 U15503 ( .B1(n13358), .B2(n13357), .A(n13356), .ZN(P2_U3207) );
  OAI211_X1 U15504 ( .C1(n13361), .C2(n13360), .A(n13275), .B(n13359), .ZN(
        n13370) );
  NAND2_X1 U15505 ( .A1(n13641), .A2(n13642), .ZN(n13363) );
  NAND2_X1 U15506 ( .A1(n13382), .A2(n13640), .ZN(n13362) );
  NAND2_X1 U15507 ( .A1(n13363), .A2(n13362), .ZN(n13676) );
  INV_X1 U15508 ( .A(n13676), .ZN(n13365) );
  OAI22_X1 U15509 ( .A1(n13366), .A2(n13365), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13364), .ZN(n13367) );
  AOI21_X1 U15510 ( .B1(n13686), .B2(n13368), .A(n13367), .ZN(n13369) );
  OAI211_X1 U15511 ( .C1(n6953), .C2(n13371), .A(n13370), .B(n13369), .ZN(
        P2_U3210) );
  MUX2_X1 U15512 ( .A(n13372), .B(P2_DATAO_REG_31__SCAN_IN), .S(n13397), .Z(
        P2_U3562) );
  MUX2_X1 U15513 ( .A(n13373), .B(P2_DATAO_REG_30__SCAN_IN), .S(n13397), .Z(
        P2_U3561) );
  MUX2_X1 U15514 ( .A(n13374), .B(P2_DATAO_REG_29__SCAN_IN), .S(n13397), .Z(
        P2_U3560) );
  MUX2_X1 U15515 ( .A(n13375), .B(P2_DATAO_REG_28__SCAN_IN), .S(n13397), .Z(
        P2_U3559) );
  MUX2_X1 U15516 ( .A(n13376), .B(P2_DATAO_REG_27__SCAN_IN), .S(n13397), .Z(
        P2_U3558) );
  MUX2_X1 U15517 ( .A(n13377), .B(P2_DATAO_REG_26__SCAN_IN), .S(n13397), .Z(
        P2_U3557) );
  MUX2_X1 U15518 ( .A(n13378), .B(P2_DATAO_REG_25__SCAN_IN), .S(n13397), .Z(
        P2_U3556) );
  MUX2_X1 U15519 ( .A(n13379), .B(P2_DATAO_REG_24__SCAN_IN), .S(n13397), .Z(
        P2_U3555) );
  MUX2_X1 U15520 ( .A(n13380), .B(P2_DATAO_REG_23__SCAN_IN), .S(n13397), .Z(
        P2_U3554) );
  MUX2_X1 U15521 ( .A(n13625), .B(P2_DATAO_REG_22__SCAN_IN), .S(n13397), .Z(
        P2_U3553) );
  MUX2_X1 U15522 ( .A(n13643), .B(P2_DATAO_REG_21__SCAN_IN), .S(n13397), .Z(
        P2_U3552) );
  MUX2_X1 U15523 ( .A(n13624), .B(P2_DATAO_REG_20__SCAN_IN), .S(n13397), .Z(
        P2_U3551) );
  INV_X2 U15524 ( .A(P2_U3947), .ZN(n13397) );
  MUX2_X1 U15525 ( .A(n13641), .B(P2_DATAO_REG_19__SCAN_IN), .S(n13397), .Z(
        P2_U3550) );
  MUX2_X1 U15526 ( .A(n13381), .B(P2_DATAO_REG_18__SCAN_IN), .S(n13397), .Z(
        P2_U3549) );
  MUX2_X1 U15527 ( .A(n13382), .B(P2_DATAO_REG_17__SCAN_IN), .S(n13397), .Z(
        P2_U3548) );
  MUX2_X1 U15528 ( .A(n13383), .B(P2_DATAO_REG_16__SCAN_IN), .S(n13397), .Z(
        P2_U3547) );
  MUX2_X1 U15529 ( .A(n13384), .B(P2_DATAO_REG_15__SCAN_IN), .S(n13397), .Z(
        P2_U3546) );
  MUX2_X1 U15530 ( .A(n13385), .B(P2_DATAO_REG_14__SCAN_IN), .S(n13397), .Z(
        P2_U3545) );
  MUX2_X1 U15531 ( .A(n13386), .B(P2_DATAO_REG_13__SCAN_IN), .S(n13397), .Z(
        P2_U3544) );
  MUX2_X1 U15532 ( .A(n13387), .B(P2_DATAO_REG_12__SCAN_IN), .S(n13397), .Z(
        P2_U3543) );
  MUX2_X1 U15533 ( .A(n13388), .B(P2_DATAO_REG_11__SCAN_IN), .S(n13397), .Z(
        P2_U3542) );
  MUX2_X1 U15534 ( .A(n13389), .B(P2_DATAO_REG_10__SCAN_IN), .S(n13397), .Z(
        P2_U3541) );
  MUX2_X1 U15535 ( .A(n13390), .B(P2_DATAO_REG_9__SCAN_IN), .S(n13397), .Z(
        P2_U3540) );
  MUX2_X1 U15536 ( .A(n13391), .B(P2_DATAO_REG_8__SCAN_IN), .S(n13397), .Z(
        P2_U3539) );
  MUX2_X1 U15537 ( .A(n13392), .B(P2_DATAO_REG_7__SCAN_IN), .S(n13397), .Z(
        P2_U3538) );
  MUX2_X1 U15538 ( .A(n13393), .B(P2_DATAO_REG_6__SCAN_IN), .S(n13397), .Z(
        P2_U3537) );
  MUX2_X1 U15539 ( .A(n13394), .B(P2_DATAO_REG_5__SCAN_IN), .S(n13397), .Z(
        P2_U3536) );
  MUX2_X1 U15540 ( .A(n8833), .B(P2_DATAO_REG_4__SCAN_IN), .S(n13397), .Z(
        P2_U3535) );
  MUX2_X1 U15541 ( .A(n13395), .B(P2_DATAO_REG_3__SCAN_IN), .S(n13397), .Z(
        P2_U3534) );
  MUX2_X1 U15542 ( .A(n8841), .B(P2_DATAO_REG_2__SCAN_IN), .S(n13397), .Z(
        P2_U3533) );
  MUX2_X1 U15543 ( .A(n13396), .B(P2_DATAO_REG_1__SCAN_IN), .S(n13397), .Z(
        P2_U3532) );
  MUX2_X1 U15544 ( .A(n8838), .B(P2_DATAO_REG_0__SCAN_IN), .S(n13397), .Z(
        P2_U3531) );
  OAI211_X1 U15545 ( .C1(n13400), .C2(n13399), .A(n14913), .B(n13398), .ZN(
        n13407) );
  OAI211_X1 U15546 ( .C1(n13403), .C2(n13402), .A(n14918), .B(n13401), .ZN(
        n13406) );
  AOI22_X1 U15547 ( .A1(n14800), .A2(P2_ADDR_REG_1__SCAN_IN), .B1(
        P2_REG3_REG_1__SCAN_IN), .B2(P2_U3088), .ZN(n13405) );
  NAND2_X1 U15548 ( .A1(n14890), .A2(n8037), .ZN(n13404) );
  NAND4_X1 U15549 ( .A1(n13407), .A2(n13406), .A3(n13405), .A4(n13404), .ZN(
        P2_U3215) );
  NAND2_X1 U15550 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_U3088), .ZN(n13408) );
  OAI21_X1 U15551 ( .B1(n14922), .B2(n13409), .A(n13408), .ZN(n13410) );
  AOI21_X1 U15552 ( .B1(n14800), .B2(P2_ADDR_REG_3__SCAN_IN), .A(n13410), .ZN(
        n13419) );
  OAI211_X1 U15553 ( .C1(n13413), .C2(n13412), .A(n14918), .B(n13411), .ZN(
        n13418) );
  OAI211_X1 U15554 ( .C1(n13416), .C2(n13415), .A(n14913), .B(n13414), .ZN(
        n13417) );
  NAND3_X1 U15555 ( .A1(n13419), .A2(n13418), .A3(n13417), .ZN(P2_U3217) );
  NAND2_X1 U15556 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_U3088), .ZN(n13420) );
  OAI21_X1 U15557 ( .B1(n14922), .B2(n13421), .A(n13420), .ZN(n13422) );
  AOI21_X1 U15558 ( .B1(n14800), .B2(P2_ADDR_REG_4__SCAN_IN), .A(n13422), .ZN(
        n13431) );
  OAI211_X1 U15559 ( .C1(n13425), .C2(n13424), .A(n14918), .B(n13423), .ZN(
        n13430) );
  OAI211_X1 U15560 ( .C1(n13428), .C2(n13427), .A(n14913), .B(n13426), .ZN(
        n13429) );
  NAND3_X1 U15561 ( .A1(n13431), .A2(n13430), .A3(n13429), .ZN(P2_U3218) );
  OAI21_X1 U15562 ( .B1(n14922), .B2(n13433), .A(n13432), .ZN(n13434) );
  AOI21_X1 U15563 ( .B1(n14800), .B2(P2_ADDR_REG_6__SCAN_IN), .A(n13434), .ZN(
        n13443) );
  OAI211_X1 U15564 ( .C1(n13437), .C2(n13436), .A(n14918), .B(n13435), .ZN(
        n13442) );
  OAI211_X1 U15565 ( .C1(n13440), .C2(n13439), .A(n14913), .B(n13438), .ZN(
        n13441) );
  NAND3_X1 U15566 ( .A1(n13443), .A2(n13442), .A3(n13441), .ZN(P2_U3220) );
  NAND2_X1 U15567 ( .A1(n14890), .A2(n13444), .ZN(n13446) );
  NAND2_X1 U15568 ( .A1(P2_REG3_REG_7__SCAN_IN), .A2(P2_U3088), .ZN(n13445) );
  OAI211_X1 U15569 ( .C1(n13447), .C2(n14926), .A(n13446), .B(n13445), .ZN(
        n13448) );
  INV_X1 U15570 ( .A(n13448), .ZN(n13457) );
  OAI211_X1 U15571 ( .C1(n13451), .C2(n13450), .A(n14913), .B(n13449), .ZN(
        n13456) );
  OAI211_X1 U15572 ( .C1(n13454), .C2(n13453), .A(n14918), .B(n13452), .ZN(
        n13455) );
  NAND3_X1 U15573 ( .A1(n13457), .A2(n13456), .A3(n13455), .ZN(P2_U3221) );
  AOI21_X1 U15574 ( .B1(n13467), .B2(P2_REG2_REG_16__SCAN_IN), .A(n13458), 
        .ZN(n14915) );
  OR2_X1 U15575 ( .A1(n13468), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n13460) );
  NAND2_X1 U15576 ( .A1(n13468), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n13459) );
  NAND2_X1 U15577 ( .A1(n13460), .A2(n13459), .ZN(n14916) );
  NOR2_X1 U15578 ( .A1(n14915), .A2(n14916), .ZN(n14914) );
  AOI21_X1 U15579 ( .B1(P2_REG2_REG_17__SCAN_IN), .B2(n13468), .A(n14914), 
        .ZN(n13480) );
  INV_X1 U15580 ( .A(n13480), .ZN(n13461) );
  XNOR2_X1 U15581 ( .A(n13479), .B(n13461), .ZN(n13463) );
  INV_X1 U15582 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n13462) );
  NAND2_X1 U15583 ( .A1(n13463), .A2(n13462), .ZN(n13482) );
  OAI21_X1 U15584 ( .B1(n13463), .B2(n13462), .A(n13482), .ZN(n13473) );
  NAND2_X1 U15585 ( .A1(P2_REG3_REG_18__SCAN_IN), .A2(P2_U3088), .ZN(n13465)
         );
  NAND2_X1 U15586 ( .A1(n14800), .A2(P2_ADDR_REG_18__SCAN_IN), .ZN(n13464) );
  OAI211_X1 U15587 ( .C1(n14922), .C2(n13479), .A(n13465), .B(n13464), .ZN(
        n13472) );
  AOI21_X1 U15588 ( .B1(n13467), .B2(P2_REG1_REG_16__SCAN_IN), .A(n13466), 
        .ZN(n14910) );
  XNOR2_X1 U15589 ( .A(n13468), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n14911) );
  NOR2_X1 U15590 ( .A1(n14910), .A2(n14911), .ZN(n14909) );
  XNOR2_X1 U15591 ( .A(n13479), .B(n13475), .ZN(n13470) );
  NOR2_X1 U15592 ( .A1(n13469), .A2(n13470), .ZN(n13477) );
  AOI211_X1 U15593 ( .C1(n13470), .C2(n13469), .A(n13477), .B(n14884), .ZN(
        n13471) );
  AOI211_X1 U15594 ( .C1(n14918), .C2(n13473), .A(n13472), .B(n13471), .ZN(
        n13474) );
  INV_X1 U15595 ( .A(n13474), .ZN(P2_U3232) );
  NOR2_X1 U15596 ( .A1(n13475), .A2(n13479), .ZN(n13476) );
  NOR2_X1 U15597 ( .A1(n13477), .A2(n13476), .ZN(n13478) );
  XOR2_X1 U15598 ( .A(n13478), .B(P2_REG1_REG_19__SCAN_IN), .Z(n13485) );
  NAND2_X1 U15599 ( .A1(n13480), .A2(n13479), .ZN(n13481) );
  NAND2_X1 U15600 ( .A1(n13482), .A2(n13481), .ZN(n13483) );
  XNOR2_X1 U15601 ( .A(P2_REG2_REG_19__SCAN_IN), .B(n13483), .ZN(n13489) );
  INV_X1 U15602 ( .A(n13489), .ZN(n13484) );
  OAI22_X1 U15603 ( .A1(n13485), .A2(n14884), .B1(n13484), .B2(n14880), .ZN(
        n13492) );
  INV_X1 U15604 ( .A(n13485), .ZN(n13486) );
  OAI21_X1 U15605 ( .B1(n14884), .B2(n13486), .A(n14922), .ZN(n13487) );
  INV_X1 U15606 ( .A(n13487), .ZN(n13488) );
  OAI21_X1 U15607 ( .B1(n13489), .B2(n14880), .A(n13488), .ZN(n13491) );
  OAI21_X1 U15608 ( .B1(n14926), .B2(n7399), .A(n13493), .ZN(n13494) );
  INV_X1 U15609 ( .A(n13498), .ZN(n13699) );
  AOI21_X1 U15610 ( .B1(n13498), .B2(n13497), .A(n13496), .ZN(n13696) );
  NAND2_X1 U15611 ( .A1(n13696), .A2(n13669), .ZN(n13501) );
  AOI21_X1 U15612 ( .B1(n13671), .B2(P2_REG2_REG_30__SCAN_IN), .A(n13499), 
        .ZN(n13500) );
  OAI211_X1 U15613 ( .C1(n13699), .C2(n13688), .A(n13501), .B(n13500), .ZN(
        P2_U3235) );
  XNOR2_X1 U15614 ( .A(n13503), .B(n13502), .ZN(n13709) );
  OAI211_X1 U15615 ( .C1(n13506), .C2(n13505), .A(n13504), .B(n13645), .ZN(
        n13508) );
  AOI211_X1 U15616 ( .C1(n13706), .C2(n13515), .A(n14996), .B(n13509), .ZN(
        n13705) );
  NAND2_X1 U15617 ( .A1(n13705), .A2(n13680), .ZN(n13510) );
  OAI211_X1 U15618 ( .C1(n13511), .C2(n13607), .A(n13708), .B(n13510), .ZN(
        n13512) );
  NAND2_X1 U15619 ( .A1(n13512), .A2(n13606), .ZN(n13514) );
  AOI22_X1 U15620 ( .A1(n13706), .A2(n13553), .B1(n13671), .B2(
        P2_REG2_REG_28__SCAN_IN), .ZN(n13513) );
  OAI211_X1 U15621 ( .C1(n13649), .C2(n13709), .A(n13514), .B(n13513), .ZN(
        P2_U3237) );
  INV_X1 U15622 ( .A(n13534), .ZN(n13517) );
  INV_X1 U15623 ( .A(n13515), .ZN(n13516) );
  AOI211_X1 U15624 ( .C1(n13711), .C2(n13517), .A(n14996), .B(n13516), .ZN(
        n13713) );
  XNOR2_X1 U15625 ( .A(n13519), .B(n13518), .ZN(n13521) );
  OAI21_X1 U15626 ( .B1(n13521), .B2(n13594), .A(n13520), .ZN(n13710) );
  AOI21_X1 U15627 ( .B1(n13713), .B2(n13680), .A(n13710), .ZN(n13530) );
  XNOR2_X1 U15628 ( .A(n13523), .B(n13522), .ZN(n13715) );
  INV_X1 U15629 ( .A(n13715), .ZN(n13528) );
  AOI22_X1 U15630 ( .A1(n13524), .A2(n13685), .B1(P2_REG2_REG_27__SCAN_IN), 
        .B2(n13671), .ZN(n13525) );
  OAI21_X1 U15631 ( .B1(n13526), .B2(n13688), .A(n13525), .ZN(n13527) );
  AOI21_X1 U15632 ( .B1(n13528), .B2(n13690), .A(n13527), .ZN(n13529) );
  OAI21_X1 U15633 ( .B1(n13530), .B2(n13671), .A(n13529), .ZN(P2_U3238) );
  XNOR2_X1 U15634 ( .A(n13531), .B(n13538), .ZN(n13533) );
  AOI21_X1 U15635 ( .B1(n13533), .B2(n13677), .A(n13532), .ZN(n13722) );
  AOI21_X1 U15636 ( .B1(n13719), .B2(n13556), .A(n13534), .ZN(n13720) );
  AOI22_X1 U15637 ( .A1(n13535), .A2(n13685), .B1(P2_REG2_REG_26__SCAN_IN), 
        .B2(n13671), .ZN(n13536) );
  OAI21_X1 U15638 ( .B1(n13537), .B2(n13688), .A(n13536), .ZN(n13541) );
  XNOR2_X1 U15639 ( .A(n13539), .B(n13538), .ZN(n13723) );
  NOR2_X1 U15640 ( .A1(n13723), .A2(n13649), .ZN(n13540) );
  AOI211_X1 U15641 ( .C1(n13720), .C2(n13669), .A(n13541), .B(n13540), .ZN(
        n13542) );
  OAI21_X1 U15642 ( .B1(n13722), .B2(n13671), .A(n13542), .ZN(P2_U3239) );
  XNOR2_X1 U15643 ( .A(n13543), .B(n13547), .ZN(n13545) );
  AOI21_X1 U15644 ( .B1(n13545), .B2(n13677), .A(n13544), .ZN(n13727) );
  OAI21_X1 U15645 ( .B1(n13548), .B2(n13547), .A(n13546), .ZN(n13549) );
  INV_X1 U15646 ( .A(n13549), .ZN(n13728) );
  INV_X1 U15647 ( .A(P2_REG2_REG_25__SCAN_IN), .ZN(n13550) );
  OAI22_X1 U15648 ( .A1(n13551), .A2(n13607), .B1(n13550), .B2(n13606), .ZN(
        n13552) );
  AOI21_X1 U15649 ( .B1(n13724), .B2(n13553), .A(n13552), .ZN(n13558) );
  NAND2_X1 U15650 ( .A1(n13724), .A2(n13554), .ZN(n13555) );
  AND2_X1 U15651 ( .A1(n13556), .A2(n13555), .ZN(n13725) );
  NAND2_X1 U15652 ( .A1(n13725), .A2(n13669), .ZN(n13557) );
  OAI211_X1 U15653 ( .C1(n13728), .C2(n13649), .A(n13558), .B(n13557), .ZN(
        n13559) );
  INV_X1 U15654 ( .A(n13559), .ZN(n13560) );
  OAI21_X1 U15655 ( .B1(n13727), .B2(n13671), .A(n13560), .ZN(P2_U3240) );
  AND2_X1 U15656 ( .A1(n13562), .A2(n13561), .ZN(n13563) );
  NOR2_X1 U15657 ( .A1(n13564), .A2(n13563), .ZN(n13573) );
  OAI22_X1 U15658 ( .A1(n7152), .A2(n13657), .B1(n13598), .B2(n13655), .ZN(
        n13569) );
  XNOR2_X1 U15659 ( .A(n13566), .B(n13565), .ZN(n13567) );
  NOR2_X1 U15660 ( .A1(n13567), .A2(n13594), .ZN(n13568) );
  AOI211_X1 U15661 ( .C1(n13570), .C2(n13573), .A(n13569), .B(n13568), .ZN(
        n13732) );
  XOR2_X1 U15662 ( .A(n13585), .B(n13729), .Z(n13730) );
  AOI22_X1 U15663 ( .A1(n13571), .A2(n13685), .B1(P2_REG2_REG_24__SCAN_IN), 
        .B2(n13671), .ZN(n13572) );
  OAI21_X1 U15664 ( .B1(n6957), .B2(n13688), .A(n13572), .ZN(n13575) );
  INV_X1 U15665 ( .A(n13573), .ZN(n13733) );
  NOR2_X1 U15666 ( .A1(n13733), .A2(n13666), .ZN(n13574) );
  AOI211_X1 U15667 ( .C1(n13730), .C2(n13669), .A(n13575), .B(n13574), .ZN(
        n13576) );
  OAI21_X1 U15668 ( .B1(n13732), .B2(n13671), .A(n13576), .ZN(P2_U3241) );
  OAI21_X1 U15669 ( .B1(n13579), .B2(n13578), .A(n13577), .ZN(n13581) );
  AOI21_X1 U15670 ( .B1(n13581), .B2(n13677), .A(n13580), .ZN(n13738) );
  OAI21_X1 U15671 ( .B1(n13584), .B2(n13583), .A(n13582), .ZN(n13734) );
  AOI21_X1 U15672 ( .B1(n13735), .B2(n13601), .A(n6958), .ZN(n13736) );
  NAND2_X1 U15673 ( .A1(n13736), .A2(n13669), .ZN(n13589) );
  INV_X1 U15674 ( .A(n13586), .ZN(n13587) );
  AOI22_X1 U15675 ( .A1(n13587), .A2(n13685), .B1(P2_REG2_REG_23__SCAN_IN), 
        .B2(n13671), .ZN(n13588) );
  OAI211_X1 U15676 ( .C1(n13590), .C2(n13688), .A(n13589), .B(n13588), .ZN(
        n13591) );
  AOI21_X1 U15677 ( .B1(n13734), .B2(n13690), .A(n13591), .ZN(n13592) );
  OAI21_X1 U15678 ( .B1(n13738), .B2(n13671), .A(n13592), .ZN(P2_U3242) );
  AOI211_X1 U15679 ( .C1(n13596), .C2(n13595), .A(n13594), .B(n13593), .ZN(
        n13600) );
  OAI22_X1 U15680 ( .A1(n13598), .A2(n13657), .B1(n13597), .B2(n13655), .ZN(
        n13599) );
  NOR2_X1 U15681 ( .A1(n13600), .A2(n13599), .ZN(n13746) );
  INV_X1 U15682 ( .A(n13601), .ZN(n13602) );
  AOI21_X1 U15683 ( .B1(n13740), .B2(n13603), .A(n13602), .ZN(n13741) );
  NOR2_X1 U15684 ( .A1(n13604), .A2(n13688), .ZN(n13610) );
  INV_X1 U15685 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n13605) );
  OAI22_X1 U15686 ( .A1(n13608), .A2(n13607), .B1(n13606), .B2(n13605), .ZN(
        n13609) );
  AOI211_X1 U15687 ( .C1(n13741), .C2(n13669), .A(n13610), .B(n13609), .ZN(
        n13615) );
  NAND2_X1 U15688 ( .A1(n13613), .A2(n13612), .ZN(n13742) );
  NAND3_X1 U15689 ( .A1(n13743), .A2(n13742), .A3(n13690), .ZN(n13614) );
  OAI211_X1 U15690 ( .C1(n13746), .C2(n13671), .A(n13615), .B(n13614), .ZN(
        P2_U3243) );
  XNOR2_X1 U15691 ( .A(n13617), .B(n13616), .ZN(n13751) );
  XNOR2_X1 U15692 ( .A(n13631), .B(n13747), .ZN(n13748) );
  INV_X1 U15693 ( .A(n13618), .ZN(n13619) );
  AOI22_X1 U15694 ( .A1(n13671), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n13619), 
        .B2(n13685), .ZN(n13620) );
  OAI21_X1 U15695 ( .B1(n13621), .B2(n13688), .A(n13620), .ZN(n13628) );
  XNOR2_X1 U15696 ( .A(n13623), .B(n13622), .ZN(n13626) );
  AOI222_X1 U15697 ( .A1(n13645), .A2(n13626), .B1(n13625), .B2(n13642), .C1(
        n13624), .C2(n13640), .ZN(n13750) );
  NOR2_X1 U15698 ( .A1(n13750), .A2(n13671), .ZN(n13627) );
  AOI211_X1 U15699 ( .C1(n13748), .C2(n13669), .A(n13628), .B(n13627), .ZN(
        n13629) );
  OAI21_X1 U15700 ( .B1(n13649), .B2(n13751), .A(n13629), .ZN(P2_U3244) );
  XNOR2_X1 U15701 ( .A(n13630), .B(n13637), .ZN(n13756) );
  AOI21_X1 U15702 ( .B1(n13752), .B2(n13662), .A(n13631), .ZN(n13753) );
  AOI22_X1 U15703 ( .A1(n13671), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n13632), 
        .B2(n13685), .ZN(n13633) );
  OAI21_X1 U15704 ( .B1(n13634), .B2(n13688), .A(n13633), .ZN(n13647) );
  INV_X1 U15705 ( .A(n13635), .ZN(n13639) );
  NAND3_X1 U15706 ( .A1(n13650), .A2(n13637), .A3(n13636), .ZN(n13638) );
  NAND2_X1 U15707 ( .A1(n13639), .A2(n13638), .ZN(n13644) );
  AOI222_X1 U15708 ( .A1(n13645), .A2(n13644), .B1(n13643), .B2(n13642), .C1(
        n13641), .C2(n13640), .ZN(n13755) );
  NOR2_X1 U15709 ( .A1(n13755), .A2(n13671), .ZN(n13646) );
  AOI211_X1 U15710 ( .C1(n13753), .C2(n13669), .A(n13647), .B(n13646), .ZN(
        n13648) );
  OAI21_X1 U15711 ( .B1(n13756), .B2(n13649), .A(n13648), .ZN(P2_U3245) );
  OAI21_X1 U15712 ( .B1(n13652), .B2(n13651), .A(n13650), .ZN(n13661) );
  XNOR2_X1 U15713 ( .A(n13653), .B(n13652), .ZN(n13761) );
  NOR2_X1 U15714 ( .A1(n13761), .A2(n13654), .ZN(n13660) );
  OAI22_X1 U15715 ( .A1(n13658), .A2(n13657), .B1(n13656), .B2(n13655), .ZN(
        n13659) );
  AOI211_X1 U15716 ( .C1(n13661), .C2(n13677), .A(n13660), .B(n13659), .ZN(
        n13760) );
  INV_X1 U15717 ( .A(n13662), .ZN(n13663) );
  AOI21_X1 U15718 ( .B1(n13757), .B2(n13672), .A(n13663), .ZN(n13758) );
  AOI22_X1 U15719 ( .A1(n13671), .A2(P2_REG2_REG_19__SCAN_IN), .B1(n13664), 
        .B2(n13685), .ZN(n13665) );
  OAI21_X1 U15720 ( .B1(n6951), .B2(n13688), .A(n13665), .ZN(n13668) );
  NOR2_X1 U15721 ( .A1(n13761), .A2(n13666), .ZN(n13667) );
  AOI211_X1 U15722 ( .C1(n13758), .C2(n13669), .A(n13668), .B(n13667), .ZN(
        n13670) );
  OAI21_X1 U15723 ( .B1(n13760), .B2(n13671), .A(n13670), .ZN(P2_U3246) );
  INV_X1 U15724 ( .A(n13672), .ZN(n13673) );
  AOI211_X1 U15725 ( .C1(n13763), .C2(n13674), .A(n14996), .B(n13673), .ZN(
        n13762) );
  XOR2_X1 U15726 ( .A(n13675), .B(n13684), .Z(n13678) );
  AOI21_X1 U15727 ( .B1(n13678), .B2(n13677), .A(n13676), .ZN(n13765) );
  INV_X1 U15728 ( .A(n13765), .ZN(n13679) );
  AOI21_X1 U15729 ( .B1(n13762), .B2(n13680), .A(n13679), .ZN(n13693) );
  INV_X1 U15730 ( .A(n13681), .ZN(n13682) );
  AOI21_X1 U15731 ( .B1(n13684), .B2(n13683), .A(n13682), .ZN(n13766) );
  INV_X1 U15732 ( .A(n13766), .ZN(n13691) );
  AOI22_X1 U15733 ( .A1(n13671), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n13686), 
        .B2(n13685), .ZN(n13687) );
  OAI21_X1 U15734 ( .B1(n6953), .B2(n13688), .A(n13687), .ZN(n13689) );
  AOI21_X1 U15735 ( .B1(n13691), .B2(n13690), .A(n13689), .ZN(n13692) );
  OAI21_X1 U15736 ( .B1(n13693), .B2(n13671), .A(n13692), .ZN(P2_U3247) );
  MUX2_X1 U15737 ( .A(P2_REG1_REG_31__SCAN_IN), .B(n13789), .S(n15019), .Z(
        P2_U3530) );
  NAND2_X1 U15738 ( .A1(n13696), .A2(n14988), .ZN(n13698) );
  OAI211_X1 U15739 ( .C1(n14994), .C2(n13699), .A(n13698), .B(n13697), .ZN(
        n13790) );
  MUX2_X1 U15740 ( .A(P2_REG1_REG_30__SCAN_IN), .B(n13790), .S(n15019), .Z(
        P2_U3529) );
  AOI22_X1 U15741 ( .A1(n13701), .A2(n14988), .B1(n13700), .B2(n14986), .ZN(
        n13702) );
  MUX2_X1 U15742 ( .A(P2_REG1_REG_29__SCAN_IN), .B(n13791), .S(n15019), .Z(
        P2_U3528) );
  OAI211_X1 U15743 ( .C1(n14984), .C2(n13709), .A(n13708), .B(n13707), .ZN(
        n13792) );
  MUX2_X1 U15744 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n13792), .S(n15019), .Z(
        P2_U3527) );
  INV_X1 U15745 ( .A(n13716), .ZN(n13717) );
  MUX2_X1 U15746 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n13793), .S(n15019), .Z(
        P2_U3526) );
  AOI22_X1 U15747 ( .A1(n13720), .A2(n14988), .B1(n13719), .B2(n14986), .ZN(
        n13721) );
  OAI211_X1 U15748 ( .C1(n14984), .C2(n13723), .A(n13722), .B(n13721), .ZN(
        n13794) );
  MUX2_X1 U15749 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n13794), .S(n15019), .Z(
        P2_U3525) );
  AOI22_X1 U15750 ( .A1(n13725), .A2(n14988), .B1(n13724), .B2(n14986), .ZN(
        n13726) );
  OAI211_X1 U15751 ( .C1(n14984), .C2(n13728), .A(n13727), .B(n13726), .ZN(
        n13795) );
  MUX2_X1 U15752 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n13795), .S(n15019), .Z(
        P2_U3524) );
  AOI22_X1 U15753 ( .A1(n13730), .A2(n14988), .B1(n13729), .B2(n14986), .ZN(
        n13731) );
  OAI211_X1 U15754 ( .C1(n14937), .C2(n13733), .A(n13732), .B(n13731), .ZN(
        n13796) );
  MUX2_X1 U15755 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n13796), .S(n15019), .Z(
        P2_U3523) );
  INV_X1 U15756 ( .A(n13734), .ZN(n13739) );
  AOI22_X1 U15757 ( .A1(n13736), .A2(n14988), .B1(n13735), .B2(n14986), .ZN(
        n13737) );
  OAI211_X1 U15758 ( .C1(n14984), .C2(n13739), .A(n13738), .B(n13737), .ZN(
        n13797) );
  MUX2_X1 U15759 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n13797), .S(n15019), .Z(
        P2_U3522) );
  AOI22_X1 U15760 ( .A1(n13741), .A2(n14988), .B1(n13740), .B2(n14986), .ZN(
        n13745) );
  NAND3_X1 U15761 ( .A1(n13743), .A2(n15000), .A3(n13742), .ZN(n13744) );
  NAND3_X1 U15762 ( .A1(n13746), .A2(n13745), .A3(n13744), .ZN(n13798) );
  MUX2_X1 U15763 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n13798), .S(n15019), .Z(
        P2_U3521) );
  AOI22_X1 U15764 ( .A1(n13748), .A2(n14988), .B1(n13747), .B2(n14986), .ZN(
        n13749) );
  OAI211_X1 U15765 ( .C1(n14984), .C2(n13751), .A(n13750), .B(n13749), .ZN(
        n13799) );
  MUX2_X1 U15766 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n13799), .S(n15019), .Z(
        P2_U3520) );
  AOI22_X1 U15767 ( .A1(n13753), .A2(n14988), .B1(n13752), .B2(n14986), .ZN(
        n13754) );
  OAI211_X1 U15768 ( .C1(n14984), .C2(n13756), .A(n13755), .B(n13754), .ZN(
        n13800) );
  MUX2_X1 U15769 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n13800), .S(n15019), .Z(
        P2_U3519) );
  AOI22_X1 U15770 ( .A1(n13758), .A2(n14988), .B1(n13757), .B2(n14986), .ZN(
        n13759) );
  OAI211_X1 U15771 ( .C1(n13761), .C2(n14937), .A(n13760), .B(n13759), .ZN(
        n13801) );
  MUX2_X1 U15772 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n13801), .S(n15019), .Z(
        P2_U3518) );
  AOI21_X1 U15773 ( .B1(n13763), .B2(n14986), .A(n13762), .ZN(n13764) );
  OAI211_X1 U15774 ( .C1(n14984), .C2(n13766), .A(n13765), .B(n13764), .ZN(
        n13802) );
  MUX2_X1 U15775 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n13802), .S(n15019), .Z(
        P2_U3517) );
  AOI22_X1 U15776 ( .A1(n13768), .A2(n14988), .B1(n13767), .B2(n14986), .ZN(
        n13769) );
  OAI211_X1 U15777 ( .C1(n14984), .C2(n13771), .A(n13770), .B(n13769), .ZN(
        n13803) );
  MUX2_X1 U15778 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n13803), .S(n15019), .Z(
        P2_U3516) );
  AOI22_X1 U15779 ( .A1(n13773), .A2(n14988), .B1(n13772), .B2(n14986), .ZN(
        n13777) );
  NAND3_X1 U15780 ( .A1(n13775), .A2(n13774), .A3(n15000), .ZN(n13776) );
  NAND3_X1 U15781 ( .A1(n13778), .A2(n13777), .A3(n13776), .ZN(n13804) );
  MUX2_X1 U15782 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n13804), .S(n15019), .Z(
        P2_U3515) );
  AOI21_X1 U15783 ( .B1(n13780), .B2(n14986), .A(n13779), .ZN(n13781) );
  OAI211_X1 U15784 ( .C1(n14984), .C2(n13783), .A(n13782), .B(n13781), .ZN(
        n13805) );
  MUX2_X1 U15785 ( .A(P2_REG1_REG_15__SCAN_IN), .B(n13805), .S(n15019), .Z(
        P2_U3514) );
  AOI22_X1 U15786 ( .A1(n13785), .A2(n14988), .B1(n13784), .B2(n14986), .ZN(
        n13786) );
  OAI211_X1 U15787 ( .C1(n14984), .C2(n13788), .A(n13787), .B(n13786), .ZN(
        n13806) );
  MUX2_X1 U15788 ( .A(P2_REG1_REG_14__SCAN_IN), .B(n13806), .S(n15019), .Z(
        P2_U3513) );
  MUX2_X1 U15789 ( .A(P2_REG0_REG_31__SCAN_IN), .B(n13789), .S(n14953), .Z(
        P2_U3498) );
  MUX2_X1 U15790 ( .A(P2_REG0_REG_30__SCAN_IN), .B(n13790), .S(n15004), .Z(
        P2_U3497) );
  MUX2_X1 U15791 ( .A(P2_REG0_REG_29__SCAN_IN), .B(n13791), .S(n15004), .Z(
        P2_U3496) );
  MUX2_X1 U15792 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n13792), .S(n15004), .Z(
        P2_U3495) );
  MUX2_X1 U15793 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n13793), .S(n15004), .Z(
        P2_U3494) );
  MUX2_X1 U15794 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n13794), .S(n15004), .Z(
        P2_U3493) );
  MUX2_X1 U15795 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n13795), .S(n15004), .Z(
        P2_U3492) );
  MUX2_X1 U15796 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n13796), .S(n15004), .Z(
        P2_U3491) );
  MUX2_X1 U15797 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n13797), .S(n15004), .Z(
        P2_U3490) );
  MUX2_X1 U15798 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n13798), .S(n14953), .Z(
        P2_U3489) );
  MUX2_X1 U15799 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n13799), .S(n14953), .Z(
        P2_U3488) );
  MUX2_X1 U15800 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n13800), .S(n14953), .Z(
        P2_U3487) );
  MUX2_X1 U15801 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n13801), .S(n14953), .Z(
        P2_U3486) );
  MUX2_X1 U15802 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n13802), .S(n14953), .Z(
        P2_U3484) );
  MUX2_X1 U15803 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n13803), .S(n14953), .Z(
        P2_U3481) );
  MUX2_X1 U15804 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n13804), .S(n14953), .Z(
        P2_U3478) );
  MUX2_X1 U15805 ( .A(P2_REG0_REG_15__SCAN_IN), .B(n13805), .S(n14953), .Z(
        P2_U3475) );
  MUX2_X1 U15806 ( .A(P2_REG0_REG_14__SCAN_IN), .B(n13806), .S(n14953), .Z(
        P2_U3472) );
  INV_X1 U15807 ( .A(n13807), .ZN(n14291) );
  NOR4_X1 U15808 ( .A1(n13809), .A2(P2_IR_REG_30__SCAN_IN), .A3(n13808), .A4(
        P2_U3088), .ZN(n13810) );
  AOI21_X1 U15809 ( .B1(n13813), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n13810), 
        .ZN(n13811) );
  OAI21_X1 U15810 ( .B1(n14291), .B2(n13820), .A(n13811), .ZN(P2_U3296) );
  AOI21_X1 U15811 ( .B1(n13813), .B2(P1_DATAO_REG_28__SCAN_IN), .A(n13812), 
        .ZN(n13814) );
  OAI21_X1 U15812 ( .B1(n13815), .B2(n13820), .A(n13814), .ZN(P2_U3299) );
  OAI222_X1 U15813 ( .A1(n13822), .A2(n13817), .B1(n13820), .B2(n13816), .C1(
        n8820), .C2(P2_U3088), .ZN(P2_U3300) );
  INV_X1 U15814 ( .A(n13818), .ZN(n13821) );
  OAI222_X1 U15815 ( .A1(n13823), .A2(n13822), .B1(P2_U3088), .B2(n13821), 
        .C1(n13820), .C2(n13819), .ZN(P2_U3302) );
  MUX2_X1 U15816 ( .A(n13824), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3327) );
  NAND2_X1 U15817 ( .A1(n13827), .A2(n14465), .ZN(n13832) );
  AOI22_X1 U15818 ( .A1(n13969), .A2(n13975), .B1(P1_REG3_REG_27__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13831) );
  AOI22_X1 U15819 ( .A1(n13956), .A2(n14085), .B1(n13955), .B2(n13828), .ZN(
        n13830) );
  NAND2_X1 U15820 ( .A1(n14216), .A2(n14463), .ZN(n13829) );
  NAND4_X1 U15821 ( .A1(n13832), .A2(n13831), .A3(n13830), .A4(n13829), .ZN(
        P1_U3214) );
  INV_X1 U15822 ( .A(n13835), .ZN(n13836) );
  NOR3_X1 U15823 ( .A1(n6540), .A2(n13836), .A3(n13837), .ZN(n13839) );
  OAI21_X1 U15824 ( .B1(n13839), .B2(n13892), .A(n14465), .ZN(n13843) );
  AOI22_X1 U15825 ( .A1(n13969), .A2(n14121), .B1(P1_REG3_REG_23__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13842) );
  AOI22_X1 U15826 ( .A1(n13956), .A2(n14120), .B1(n13955), .B2(n14124), .ZN(
        n13841) );
  NAND2_X1 U15827 ( .A1(n14239), .A2(n14463), .ZN(n13840) );
  NAND4_X1 U15828 ( .A1(n13843), .A2(n13842), .A3(n13841), .A4(n13840), .ZN(
        P1_U3216) );
  INV_X1 U15829 ( .A(n11899), .ZN(n13855) );
  INV_X1 U15830 ( .A(n13847), .ZN(n13929) );
  OAI21_X1 U15831 ( .B1(n13929), .B2(n13845), .A(n13844), .ZN(n13849) );
  NAND2_X1 U15832 ( .A1(n13847), .A2(n13846), .ZN(n13848) );
  NAND3_X1 U15833 ( .A1(n13849), .A2(n14465), .A3(n13848), .ZN(n13854) );
  AND2_X1 U15834 ( .A1(P1_U3086), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n14053) );
  OAI22_X1 U15835 ( .A1(n13966), .A2(n13851), .B1(n14469), .B2(n13850), .ZN(
        n13852) );
  AOI211_X1 U15836 ( .C1(n13969), .C2(n13978), .A(n14053), .B(n13852), .ZN(
        n13853) );
  OAI211_X1 U15837 ( .C1(n13855), .C2(n13972), .A(n13854), .B(n13853), .ZN(
        P1_U3219) );
  OAI21_X1 U15838 ( .B1(n13858), .B2(n13857), .A(n13856), .ZN(n13859) );
  NAND2_X1 U15839 ( .A1(n13859), .A2(n14465), .ZN(n13862) );
  AOI22_X1 U15840 ( .A1(n13969), .A2(n13995), .B1(P1_REG3_REG_1__SCAN_IN), 
        .B2(n13925), .ZN(n13861) );
  AOI22_X1 U15841 ( .A1(n13956), .A2(n13996), .B1(n14463), .B2(n6473), .ZN(
        n13860) );
  NAND3_X1 U15842 ( .A1(n13862), .A2(n13861), .A3(n13860), .ZN(P1_U3222) );
  NAND2_X1 U15843 ( .A1(n6524), .A2(n13863), .ZN(n13911) );
  OAI21_X1 U15844 ( .B1(n6524), .B2(n13863), .A(n13911), .ZN(n13864) );
  NAND2_X1 U15845 ( .A1(n13864), .A2(n14465), .ZN(n13868) );
  AOI22_X1 U15846 ( .A1(n13969), .A2(n14120), .B1(P1_REG3_REG_21__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13867) );
  AOI22_X1 U15847 ( .A1(n13956), .A2(n13978), .B1(n13955), .B2(n14160), .ZN(
        n13866) );
  NAND2_X1 U15848 ( .A1(n14252), .A2(n14463), .ZN(n13865) );
  NAND4_X1 U15849 ( .A1(n13868), .A2(n13867), .A3(n13866), .A4(n13865), .ZN(
        P1_U3223) );
  AND2_X1 U15850 ( .A1(n13870), .A2(n13869), .ZN(n13893) );
  INV_X1 U15851 ( .A(n13871), .ZN(n13872) );
  NAND3_X1 U15852 ( .A1(n13893), .A2(n13873), .A3(n13872), .ZN(n13874) );
  AOI21_X1 U15853 ( .B1(n13875), .B2(n13874), .A(n13938), .ZN(n13879) );
  INV_X1 U15854 ( .A(n14226), .ZN(n14093) );
  AOI22_X1 U15855 ( .A1(n13969), .A2(n14085), .B1(P1_REG3_REG_25__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13877) );
  AOI22_X1 U15856 ( .A1(n13956), .A2(n14121), .B1(n13955), .B2(n14091), .ZN(
        n13876) );
  OAI211_X1 U15857 ( .C1(n14093), .C2(n13972), .A(n13877), .B(n13876), .ZN(
        n13878) );
  OR2_X1 U15858 ( .A1(n13879), .A2(n13878), .ZN(P1_U3225) );
  XOR2_X1 U15859 ( .A(n13881), .B(n13880), .Z(n13882) );
  XNOR2_X1 U15860 ( .A(n13883), .B(n13882), .ZN(n13888) );
  NAND2_X1 U15861 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n14644)
         );
  NAND2_X1 U15862 ( .A1(n14466), .A2(n14488), .ZN(n13884) );
  OAI211_X1 U15863 ( .C1(n14469), .C2(n13885), .A(n14644), .B(n13884), .ZN(
        n13886) );
  AOI21_X1 U15864 ( .B1(n14489), .B2(n14463), .A(n13886), .ZN(n13887) );
  OAI21_X1 U15865 ( .B1(n13888), .B2(n13938), .A(n13887), .ZN(P1_U3228) );
  INV_X1 U15866 ( .A(n14233), .ZN(n14111) );
  INV_X1 U15867 ( .A(n13889), .ZN(n13891) );
  NOR3_X1 U15868 ( .A1(n13892), .A2(n13891), .A3(n13890), .ZN(n13895) );
  INV_X1 U15869 ( .A(n13893), .ZN(n13894) );
  OAI21_X1 U15870 ( .B1(n13895), .B2(n13894), .A(n14465), .ZN(n13901) );
  NAND2_X1 U15871 ( .A1(n13976), .A2(n14457), .ZN(n13897) );
  NAND2_X1 U15872 ( .A1(n14068), .A2(n14455), .ZN(n13896) );
  AND2_X1 U15873 ( .A1(n13897), .A2(n13896), .ZN(n14104) );
  OAI22_X1 U15874 ( .A1(n13934), .A2(n14104), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13898), .ZN(n13899) );
  AOI21_X1 U15875 ( .B1(n14109), .B2(n13955), .A(n13899), .ZN(n13900) );
  OAI211_X1 U15876 ( .C1(n14111), .C2(n13972), .A(n13901), .B(n13900), .ZN(
        P1_U3229) );
  XNOR2_X1 U15877 ( .A(n6531), .B(n13902), .ZN(n13910) );
  INV_X1 U15878 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n13903) );
  OAI22_X1 U15879 ( .A1(n13934), .A2(n13904), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13903), .ZN(n13907) );
  NOR2_X1 U15880 ( .A1(n13905), .A2(n13972), .ZN(n13906) );
  AOI211_X1 U15881 ( .C1(n13908), .C2(n13955), .A(n13907), .B(n13906), .ZN(
        n13909) );
  OAI21_X1 U15882 ( .B1(n13910), .B2(n13938), .A(n13909), .ZN(P1_U3233) );
  INV_X1 U15883 ( .A(n13911), .ZN(n13914) );
  NOR3_X1 U15884 ( .A1(n13914), .A2(n13913), .A3(n13912), .ZN(n13915) );
  OAI21_X1 U15885 ( .B1(n13915), .B2(n6540), .A(n14465), .ZN(n13919) );
  AOI22_X1 U15886 ( .A1(n14457), .A2(n13977), .B1(n13976), .B2(n14455), .ZN(
        n14143) );
  OAI22_X1 U15887 ( .A1(n13934), .A2(n14143), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13916), .ZN(n13917) );
  AOI21_X1 U15888 ( .B1(n14148), .B2(n13955), .A(n13917), .ZN(n13918) );
  OAI211_X1 U15889 ( .C1(n13972), .C2(n13920), .A(n13919), .B(n13918), .ZN(
        P1_U3235) );
  OAI21_X1 U15890 ( .B1(n13923), .B2(n13922), .A(n13921), .ZN(n13924) );
  NAND2_X1 U15891 ( .A1(n13924), .A2(n14465), .ZN(n13928) );
  AOI22_X1 U15892 ( .A1(n13969), .A2(n13994), .B1(P1_REG3_REG_2__SCAN_IN), 
        .B2(n13925), .ZN(n13927) );
  AOI22_X1 U15893 ( .A1(n13956), .A2(n14187), .B1(n14463), .B2(n14728), .ZN(
        n13926) );
  NAND3_X1 U15894 ( .A1(n13928), .A2(n13927), .A3(n13926), .ZN(P1_U3237) );
  AOI21_X1 U15895 ( .B1(n13931), .B2(n13930), .A(n13929), .ZN(n13939) );
  NAND2_X1 U15896 ( .A1(n13955), .A2(n13932), .ZN(n13933) );
  NAND2_X1 U15897 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n14659)
         );
  OAI211_X1 U15898 ( .C1(n13935), .C2(n13934), .A(n13933), .B(n14659), .ZN(
        n13936) );
  AOI21_X1 U15899 ( .B1(n14270), .B2(n14463), .A(n13936), .ZN(n13937) );
  OAI21_X1 U15900 ( .B1(n13939), .B2(n13938), .A(n13937), .ZN(P1_U3238) );
  OAI211_X1 U15901 ( .C1(n13942), .C2(n13941), .A(n13940), .B(n14465), .ZN(
        n13950) );
  AOI22_X1 U15902 ( .A1(n14466), .A2(n13943), .B1(P1_REG3_REG_6__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13949) );
  OR2_X1 U15903 ( .A1(n14469), .A2(n13944), .ZN(n13948) );
  AND2_X1 U15904 ( .A1(n13945), .A2(n14777), .ZN(n14744) );
  NAND2_X1 U15905 ( .A1(n13946), .A2(n14744), .ZN(n13947) );
  NAND4_X1 U15906 ( .A1(n13950), .A2(n13949), .A3(n13948), .A4(n13947), .ZN(
        P1_U3239) );
  OAI21_X1 U15907 ( .B1(n13953), .B2(n13952), .A(n13951), .ZN(n13954) );
  NAND2_X1 U15908 ( .A1(n13954), .A2(n14465), .ZN(n13960) );
  AOI22_X1 U15909 ( .A1(n13969), .A2(n14069), .B1(P1_REG3_REG_26__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13959) );
  AOI22_X1 U15910 ( .A1(n13956), .A2(n14068), .B1(n13955), .B2(n14073), .ZN(
        n13958) );
  NAND2_X1 U15911 ( .A1(n14221), .A2(n14463), .ZN(n13957) );
  NAND4_X1 U15912 ( .A1(n13960), .A2(n13959), .A3(n13958), .A4(n13957), .ZN(
        P1_U3240) );
  OAI211_X1 U15913 ( .C1(n13962), .C2(n13961), .A(n14448), .B(n14465), .ZN(
        n13971) );
  INV_X1 U15914 ( .A(n13963), .ZN(n13964) );
  OAI22_X1 U15915 ( .A1(n13966), .A2(n13965), .B1(n14469), .B2(n13964), .ZN(
        n13967) );
  AOI211_X1 U15916 ( .C1(n13969), .C2(n13983), .A(n13968), .B(n13967), .ZN(
        n13970) );
  OAI211_X1 U15917 ( .C1(n14506), .C2(n13972), .A(n13971), .B(n13970), .ZN(
        P1_U3241) );
  MUX2_X1 U15918 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(n14059), .S(P1_U4016), .Z(
        P1_U3591) );
  MUX2_X1 U15919 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n13973), .S(P1_U4016), .Z(
        P1_U3590) );
  MUX2_X1 U15920 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n13974), .S(P1_U4016), .Z(
        P1_U3589) );
  MUX2_X1 U15921 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n13975), .S(P1_U4016), .Z(
        P1_U3588) );
  MUX2_X1 U15922 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n14069), .S(P1_U4016), .Z(
        P1_U3587) );
  MUX2_X1 U15923 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n14085), .S(P1_U4016), .Z(
        P1_U3586) );
  MUX2_X1 U15924 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n14068), .S(P1_U4016), .Z(
        P1_U3585) );
  MUX2_X1 U15925 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n14121), .S(P1_U4016), .Z(
        P1_U3584) );
  MUX2_X1 U15926 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n13976), .S(P1_U4016), .Z(
        P1_U3583) );
  MUX2_X1 U15927 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n14120), .S(P1_U4016), .Z(
        P1_U3582) );
  MUX2_X1 U15928 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n13977), .S(P1_U4016), .Z(
        P1_U3581) );
  MUX2_X1 U15929 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n13978), .S(P1_U4016), .Z(
        P1_U3580) );
  MUX2_X1 U15930 ( .A(n13980), .B(P1_DATAO_REG_19__SCAN_IN), .S(n13979), .Z(
        P1_U3579) );
  MUX2_X1 U15931 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n13981), .S(P1_U4016), .Z(
        P1_U3578) );
  MUX2_X1 U15932 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n13982), .S(P1_U4016), .Z(
        P1_U3577) );
  MUX2_X1 U15933 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n13983), .S(P1_U4016), .Z(
        P1_U3576) );
  MUX2_X1 U15934 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n13984), .S(P1_U4016), .Z(
        P1_U3575) );
  MUX2_X1 U15935 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n13985), .S(P1_U4016), .Z(
        P1_U3574) );
  MUX2_X1 U15936 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n13986), .S(P1_U4016), .Z(
        P1_U3573) );
  MUX2_X1 U15937 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n14456), .S(P1_U4016), .Z(
        P1_U3572) );
  MUX2_X1 U15938 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n13987), .S(P1_U4016), .Z(
        P1_U3571) );
  MUX2_X1 U15939 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n14458), .S(P1_U4016), .Z(
        P1_U3570) );
  MUX2_X1 U15940 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n13988), .S(P1_U4016), .Z(
        P1_U3569) );
  MUX2_X1 U15941 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n13989), .S(P1_U4016), .Z(
        P1_U3568) );
  MUX2_X1 U15942 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n13990), .S(P1_U4016), .Z(
        P1_U3567) );
  MUX2_X1 U15943 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n13991), .S(P1_U4016), .Z(
        P1_U3566) );
  MUX2_X1 U15944 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n13992), .S(P1_U4016), .Z(
        P1_U3565) );
  MUX2_X1 U15945 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n13993), .S(P1_U4016), .Z(
        P1_U3564) );
  MUX2_X1 U15946 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n13994), .S(P1_U4016), .Z(
        P1_U3563) );
  MUX2_X1 U15947 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n13995), .S(P1_U4016), .Z(
        P1_U3562) );
  MUX2_X1 U15948 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n14187), .S(P1_U4016), .Z(
        P1_U3561) );
  MUX2_X1 U15949 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(n13996), .S(P1_U4016), .Z(
        P1_U3560) );
  OAI211_X1 U15950 ( .C1(n13999), .C2(n13998), .A(n14633), .B(n13997), .ZN(
        n14008) );
  OAI211_X1 U15951 ( .C1(n14002), .C2(n14001), .A(n14638), .B(n14000), .ZN(
        n14007) );
  AOI22_X1 U15952 ( .A1(n14003), .A2(P1_ADDR_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(P1_U3086), .ZN(n14006) );
  NAND2_X1 U15953 ( .A1(n14658), .A2(n14004), .ZN(n14005) );
  NAND4_X1 U15954 ( .A1(n14008), .A2(n14007), .A3(n14006), .A4(n14005), .ZN(
        P1_U3244) );
  INV_X1 U15955 ( .A(n14009), .ZN(n14024) );
  OAI22_X1 U15956 ( .A1(n14661), .A2(n8902), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14010), .ZN(n14011) );
  AOI21_X1 U15957 ( .B1(n6470), .B2(n14658), .A(n14011), .ZN(n14023) );
  INV_X1 U15958 ( .A(n14013), .ZN(n14014) );
  OAI211_X1 U15959 ( .C1(n14016), .C2(n14015), .A(n14638), .B(n14014), .ZN(
        n14022) );
  INV_X1 U15960 ( .A(n14017), .ZN(n14018) );
  OAI211_X1 U15961 ( .C1(n14020), .C2(n14019), .A(n14633), .B(n14018), .ZN(
        n14021) );
  NAND4_X1 U15962 ( .A1(n14024), .A2(n14023), .A3(n14022), .A4(n14021), .ZN(
        P1_U3245) );
  INV_X1 U15963 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n14026) );
  AOI22_X1 U15964 ( .A1(n14625), .A2(n14026), .B1(P1_REG2_REG_16__SCAN_IN), 
        .B2(n14025), .ZN(n14621) );
  NAND2_X1 U15965 ( .A1(n14027), .A2(n14036), .ZN(n14029) );
  NAND2_X1 U15966 ( .A1(n14029), .A2(n14028), .ZN(n14622) );
  NOR2_X1 U15967 ( .A1(n14621), .A2(n14622), .ZN(n14620) );
  NAND2_X1 U15968 ( .A1(n14042), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n14030) );
  OAI21_X1 U15969 ( .B1(n14042), .B2(P1_REG2_REG_17__SCAN_IN), .A(n14030), 
        .ZN(n14636) );
  NOR2_X1 U15970 ( .A1(n14635), .A2(n14636), .ZN(n14634) );
  NOR2_X1 U15971 ( .A1(n14031), .A2(n14043), .ZN(n14032) );
  INV_X1 U15972 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n14653) );
  XNOR2_X1 U15973 ( .A(P1_REG2_REG_19__SCAN_IN), .B(n14033), .ZN(n14050) );
  INV_X1 U15974 ( .A(n14050), .ZN(n14048) );
  INV_X1 U15975 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n14503) );
  NOR2_X1 U15976 ( .A1(n14625), .A2(n14503), .ZN(n14034) );
  AOI21_X1 U15977 ( .B1(n14625), .B2(n14503), .A(n14034), .ZN(n14618) );
  NAND2_X1 U15978 ( .A1(n14036), .A2(n14035), .ZN(n14038) );
  NAND2_X1 U15979 ( .A1(n14038), .A2(n14037), .ZN(n14619) );
  INV_X1 U15980 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n14039) );
  OR2_X1 U15981 ( .A1(n14042), .A2(n14039), .ZN(n14041) );
  NAND2_X1 U15982 ( .A1(n14042), .A2(n14039), .ZN(n14040) );
  AND2_X1 U15983 ( .A1(n14041), .A2(n14040), .ZN(n14631) );
  XNOR2_X1 U15984 ( .A(n14043), .B(n6532), .ZN(n14650) );
  NOR2_X1 U15985 ( .A1(n14649), .A2(n14650), .ZN(n14648) );
  NOR2_X1 U15986 ( .A1(n6532), .A2(n14043), .ZN(n14044) );
  NOR2_X1 U15987 ( .A1(n14648), .A2(n14044), .ZN(n14046) );
  XOR2_X1 U15988 ( .A(n14046), .B(n14045), .Z(n14049) );
  OAI21_X1 U15989 ( .B1(n14049), .B2(n14647), .A(n14642), .ZN(n14047) );
  AOI21_X1 U15990 ( .B1(n14048), .B2(n14638), .A(n14047), .ZN(n14052) );
  AOI22_X1 U15991 ( .A1(n14050), .A2(n14638), .B1(n14633), .B2(n14049), .ZN(
        n14051) );
  MUX2_X1 U15992 ( .A(n14052), .B(n14051), .S(n14149), .Z(n14055) );
  INV_X1 U15993 ( .A(n14053), .ZN(n14054) );
  OAI211_X1 U15994 ( .C1(n14056), .C2(n14661), .A(n14055), .B(n14054), .ZN(
        P1_U3262) );
  NAND2_X1 U15995 ( .A1(n14063), .A2(n14201), .ZN(n14057) );
  XNOR2_X1 U15996 ( .A(n14057), .B(n14197), .ZN(n14195) );
  NAND2_X1 U15997 ( .A1(n14195), .A2(n14191), .ZN(n14061) );
  NAND2_X1 U15998 ( .A1(n14059), .A2(n14058), .ZN(n14199) );
  NOR2_X1 U15999 ( .A1(n14706), .A2(n14199), .ZN(n14064) );
  AOI21_X1 U16000 ( .B1(n14706), .B2(P1_REG2_REG_31__SCAN_IN), .A(n14064), 
        .ZN(n14060) );
  OAI211_X1 U16001 ( .C1(n14197), .C2(n14708), .A(n14061), .B(n14060), .ZN(
        P1_U3263) );
  XNOR2_X1 U16002 ( .A(n14063), .B(n14062), .ZN(n14198) );
  NAND2_X1 U16003 ( .A1(n14198), .A2(n14191), .ZN(n14066) );
  AOI21_X1 U16004 ( .B1(n14706), .B2(P1_REG2_REG_30__SCAN_IN), .A(n14064), 
        .ZN(n14065) );
  OAI211_X1 U16005 ( .C1(n14201), .C2(n14708), .A(n14066), .B(n14065), .ZN(
        P1_U3264) );
  XNOR2_X1 U16006 ( .A(n14067), .B(n14077), .ZN(n14070) );
  AOI222_X1 U16007 ( .A1(n14701), .A2(n14070), .B1(n14069), .B2(n14455), .C1(
        n14068), .C2(n14457), .ZN(n14223) );
  INV_X1 U16008 ( .A(n14071), .ZN(n14072) );
  AOI211_X1 U16009 ( .C1(n14221), .C2(n14089), .A(n14493), .B(n14072), .ZN(
        n14220) );
  AOI22_X1 U16010 ( .A1(n14681), .A2(P1_REG2_REG_26__SCAN_IN), .B1(n14073), 
        .B2(n14704), .ZN(n14074) );
  OAI21_X1 U16011 ( .B1(n14075), .B2(n14708), .A(n14074), .ZN(n14080) );
  OAI21_X1 U16012 ( .B1(n14078), .B2(n14077), .A(n14076), .ZN(n14224) );
  NOR2_X1 U16013 ( .A1(n14224), .A2(n14174), .ZN(n14079) );
  AOI211_X1 U16014 ( .C1(n14220), .C2(n14713), .A(n14080), .B(n14079), .ZN(
        n14081) );
  OAI21_X1 U16015 ( .B1(n14223), .B2(n14706), .A(n14081), .ZN(P1_U3267) );
  AND2_X1 U16016 ( .A1(n14083), .A2(n14082), .ZN(n14084) );
  OAI21_X1 U16017 ( .B1(n6549), .B2(n14084), .A(n14701), .ZN(n14087) );
  AOI22_X1 U16018 ( .A1(n14457), .A2(n14121), .B1(n14085), .B2(n14455), .ZN(
        n14086) );
  NAND2_X1 U16019 ( .A1(n14087), .A2(n14086), .ZN(n14231) );
  INV_X1 U16020 ( .A(n14231), .ZN(n14101) );
  AOI21_X1 U16021 ( .B1(n14226), .B2(n14108), .A(n14493), .ZN(n14090) );
  NAND2_X1 U16022 ( .A1(n14090), .A2(n14089), .ZN(n14227) );
  INV_X1 U16023 ( .A(n14227), .ZN(n14095) );
  AOI22_X1 U16024 ( .A1(n14681), .A2(P1_REG2_REG_25__SCAN_IN), .B1(n14091), 
        .B2(n14704), .ZN(n14092) );
  OAI21_X1 U16025 ( .B1(n14093), .B2(n14708), .A(n14092), .ZN(n14094) );
  AOI21_X1 U16026 ( .B1(n14095), .B2(n14713), .A(n14094), .ZN(n14100) );
  NAND2_X1 U16027 ( .A1(n14098), .A2(n14097), .ZN(n14225) );
  NAND3_X1 U16028 ( .A1(n14096), .A2(n14225), .A3(n14483), .ZN(n14099) );
  OAI211_X1 U16029 ( .C1(n14101), .C2(n14706), .A(n14100), .B(n14099), .ZN(
        P1_U3268) );
  AOI21_X1 U16030 ( .B1(n14103), .B2(n7265), .A(n14780), .ZN(n14107) );
  INV_X1 U16031 ( .A(n14104), .ZN(n14105) );
  AOI21_X1 U16032 ( .B1(n14107), .B2(n14106), .A(n14105), .ZN(n14235) );
  AOI211_X1 U16033 ( .C1(n14233), .C2(n14119), .A(n14493), .B(n14088), .ZN(
        n14232) );
  AOI22_X1 U16034 ( .A1(n14681), .A2(P1_REG2_REG_24__SCAN_IN), .B1(n14109), 
        .B2(n14704), .ZN(n14110) );
  OAI21_X1 U16035 ( .B1(n14111), .B2(n14708), .A(n14110), .ZN(n14116) );
  INV_X1 U16036 ( .A(n14112), .ZN(n14113) );
  AOI21_X1 U16037 ( .B1(n14102), .B2(n14114), .A(n14113), .ZN(n14236) );
  NOR2_X1 U16038 ( .A1(n14236), .A2(n14174), .ZN(n14115) );
  AOI211_X1 U16039 ( .C1(n14232), .C2(n14713), .A(n14116), .B(n14115), .ZN(
        n14117) );
  OAI21_X1 U16040 ( .B1(n14706), .B2(n14235), .A(n14117), .ZN(P1_U3269) );
  XNOR2_X1 U16041 ( .A(n14118), .B(n14131), .ZN(n14237) );
  INV_X1 U16042 ( .A(n14237), .ZN(n14136) );
  OAI211_X1 U16043 ( .C1(n14127), .C2(n14147), .A(n7114), .B(n14119), .ZN(
        n14241) );
  INV_X1 U16044 ( .A(n14241), .ZN(n14129) );
  NAND2_X1 U16045 ( .A1(n14120), .A2(n14457), .ZN(n14123) );
  NAND2_X1 U16046 ( .A1(n14121), .A2(n14455), .ZN(n14122) );
  NAND2_X1 U16047 ( .A1(n14123), .A2(n14122), .ZN(n14238) );
  AOI22_X1 U16048 ( .A1(n14179), .A2(n14238), .B1(n14124), .B2(n14704), .ZN(
        n14126) );
  NAND2_X1 U16049 ( .A1(n14681), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n14125) );
  OAI211_X1 U16050 ( .C1(n14127), .C2(n14708), .A(n14126), .B(n14125), .ZN(
        n14128) );
  AOI21_X1 U16051 ( .B1(n14129), .B2(n14713), .A(n14128), .ZN(n14134) );
  NAND2_X1 U16052 ( .A1(n14132), .A2(n14131), .ZN(n14240) );
  NAND3_X1 U16053 ( .A1(n14130), .A2(n14240), .A3(n14483), .ZN(n14133) );
  OAI211_X1 U16054 ( .C1(n14136), .C2(n14135), .A(n14134), .B(n14133), .ZN(
        P1_U3270) );
  XNOR2_X1 U16055 ( .A(n14137), .B(n14138), .ZN(n14249) );
  INV_X1 U16056 ( .A(n14139), .ZN(n14140) );
  AOI21_X1 U16057 ( .B1(n14142), .B2(n14141), .A(n14140), .ZN(n14144) );
  OAI21_X1 U16058 ( .B1(n14144), .B2(n14780), .A(n14143), .ZN(n14245) );
  INV_X1 U16059 ( .A(n14245), .ZN(n14151) );
  NAND2_X1 U16060 ( .A1(n14247), .A2(n14158), .ZN(n14145) );
  NAND2_X1 U16061 ( .A1(n14145), .A2(n7114), .ZN(n14146) );
  NOR2_X1 U16062 ( .A1(n14147), .A2(n14146), .ZN(n14246) );
  AOI22_X1 U16063 ( .A1(n14246), .A2(n14149), .B1(n14704), .B2(n14148), .ZN(
        n14150) );
  AOI21_X1 U16064 ( .B1(n14151), .B2(n14150), .A(n14706), .ZN(n14152) );
  INV_X1 U16065 ( .A(n14152), .ZN(n14154) );
  AOI22_X1 U16066 ( .A1(n14247), .A2(n14476), .B1(P1_REG2_REG_22__SCAN_IN), 
        .B2(n14706), .ZN(n14153) );
  OAI211_X1 U16067 ( .C1(n14249), .C2(n14174), .A(n14154), .B(n14153), .ZN(
        P1_U3271) );
  INV_X1 U16068 ( .A(n14155), .ZN(n14156) );
  AOI21_X1 U16069 ( .B1(n14165), .B2(n14157), .A(n14156), .ZN(n14255) );
  INV_X1 U16070 ( .A(n14158), .ZN(n14159) );
  AOI211_X1 U16071 ( .C1(n14252), .C2(n6622), .A(n14493), .B(n14159), .ZN(
        n14250) );
  INV_X1 U16072 ( .A(n14252), .ZN(n14162) );
  AOI22_X1 U16073 ( .A1(n14681), .A2(P1_REG2_REG_21__SCAN_IN), .B1(n14160), 
        .B2(n14704), .ZN(n14161) );
  OAI21_X1 U16074 ( .B1(n14162), .B2(n14708), .A(n14161), .ZN(n14163) );
  AOI21_X1 U16075 ( .B1(n14250), .B2(n14713), .A(n14163), .ZN(n14173) );
  OAI211_X1 U16076 ( .C1(n14166), .C2(n14165), .A(n14701), .B(n14164), .ZN(
        n14253) );
  INV_X1 U16077 ( .A(n14253), .ZN(n14171) );
  OAI22_X1 U16078 ( .A1(n14170), .A2(n14169), .B1(n14168), .B2(n14167), .ZN(
        n14251) );
  OAI21_X1 U16079 ( .B1(n14171), .B2(n14251), .A(n14179), .ZN(n14172) );
  OAI211_X1 U16080 ( .C1(n14255), .C2(n14174), .A(n14173), .B(n14172), .ZN(
        P1_U3272) );
  INV_X1 U16081 ( .A(n14175), .ZN(n14714) );
  AOI22_X1 U16082 ( .A1(n14714), .A2(n14177), .B1(n14476), .B2(n6473), .ZN(
        n14184) );
  AOI22_X1 U16083 ( .A1(n14706), .A2(P1_REG2_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(n14704), .ZN(n14183) );
  NAND2_X1 U16084 ( .A1(n14179), .A2(n14178), .ZN(n14182) );
  NAND2_X1 U16085 ( .A1(n14191), .A2(n14180), .ZN(n14181) );
  NAND4_X1 U16086 ( .A1(n14184), .A2(n14183), .A3(n14182), .A4(n14181), .ZN(
        P1_U3292) );
  OAI21_X1 U16087 ( .B1(n14483), .B2(n14186), .A(n14185), .ZN(n14194) );
  NAND2_X1 U16088 ( .A1(n14187), .A2(n14455), .ZN(n14719) );
  INV_X1 U16089 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n14189) );
  OAI22_X1 U16090 ( .A1(n14681), .A2(n14719), .B1(n14189), .B2(n14188), .ZN(
        n14190) );
  AOI21_X1 U16091 ( .B1(P1_REG2_REG_0__SCAN_IN), .B2(n14706), .A(n14190), .ZN(
        n14193) );
  OAI21_X1 U16092 ( .B1(n14476), .B2(n14191), .A(n14725), .ZN(n14192) );
  NAND3_X1 U16093 ( .A1(n14194), .A2(n14193), .A3(n14192), .ZN(P1_U3293) );
  NAND2_X1 U16094 ( .A1(n14195), .A2(n7114), .ZN(n14196) );
  OAI211_X1 U16095 ( .C1(n14753), .C2(n14197), .A(n14196), .B(n14199), .ZN(
        n14273) );
  MUX2_X1 U16096 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n14273), .S(n14799), .Z(
        P1_U3559) );
  NAND2_X1 U16097 ( .A1(n14198), .A2(n7114), .ZN(n14200) );
  OAI211_X1 U16098 ( .C1(n14753), .C2(n14201), .A(n14200), .B(n14199), .ZN(
        n14274) );
  MUX2_X1 U16099 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n14274), .S(n14799), .Z(
        P1_U3558) );
  OAI211_X1 U16100 ( .C1(n14204), .C2(n14753), .A(n14203), .B(n14202), .ZN(
        n14205) );
  MUX2_X1 U16101 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n14275), .S(n14799), .Z(
        P1_U3557) );
  NAND2_X1 U16102 ( .A1(n14209), .A2(n14777), .ZN(n14213) );
  NAND3_X1 U16103 ( .A1(n11694), .A2(n14783), .A3(n14210), .ZN(n14212) );
  NAND4_X1 U16104 ( .A1(n14214), .A2(n14213), .A3(n14212), .A4(n14211), .ZN(
        n14276) );
  MUX2_X1 U16105 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n14276), .S(n14799), .Z(
        P1_U3556) );
  AOI21_X1 U16106 ( .B1(n14216), .B2(n14777), .A(n14215), .ZN(n14217) );
  OAI211_X1 U16107 ( .C1(n14219), .C2(n14730), .A(n14218), .B(n14217), .ZN(
        n14277) );
  MUX2_X1 U16108 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n14277), .S(n14799), .Z(
        P1_U3555) );
  AOI21_X1 U16109 ( .B1(n14221), .B2(n14777), .A(n14220), .ZN(n14222) );
  OAI211_X1 U16110 ( .C1(n14721), .C2(n14224), .A(n14223), .B(n14222), .ZN(
        n14278) );
  MUX2_X1 U16111 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n14278), .S(n14799), .Z(
        P1_U3554) );
  NAND3_X1 U16112 ( .A1(n14096), .A2(n14783), .A3(n14225), .ZN(n14229) );
  NAND2_X1 U16113 ( .A1(n14226), .A2(n14777), .ZN(n14228) );
  NAND3_X1 U16114 ( .A1(n14229), .A2(n14228), .A3(n14227), .ZN(n14230) );
  MUX2_X1 U16115 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n14279), .S(n14799), .Z(
        P1_U3553) );
  AOI21_X1 U16116 ( .B1(n14233), .B2(n14777), .A(n14232), .ZN(n14234) );
  OAI211_X1 U16117 ( .C1(n14236), .C2(n14721), .A(n14235), .B(n14234), .ZN(
        n14280) );
  MUX2_X1 U16118 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n14280), .S(n14799), .Z(
        P1_U3552) );
  NAND2_X1 U16119 ( .A1(n14237), .A2(n14701), .ZN(n14244) );
  AOI21_X1 U16120 ( .B1(n14239), .B2(n14777), .A(n14238), .ZN(n14243) );
  NAND3_X1 U16121 ( .A1(n14130), .A2(n14240), .A3(n14783), .ZN(n14242) );
  NAND4_X1 U16122 ( .A1(n14244), .A2(n14243), .A3(n14242), .A4(n14241), .ZN(
        n14281) );
  MUX2_X1 U16123 ( .A(n14281), .B(P1_REG1_REG_23__SCAN_IN), .S(n14797), .Z(
        P1_U3551) );
  AOI211_X1 U16124 ( .C1(n14247), .C2(n14777), .A(n14246), .B(n14245), .ZN(
        n14248) );
  OAI21_X1 U16125 ( .B1(n14721), .B2(n14249), .A(n14248), .ZN(n14282) );
  MUX2_X1 U16126 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n14282), .S(n14799), .Z(
        P1_U3550) );
  AOI211_X1 U16127 ( .C1(n14252), .C2(n14777), .A(n14251), .B(n14250), .ZN(
        n14254) );
  OAI211_X1 U16128 ( .C1(n14255), .C2(n14721), .A(n14254), .B(n14253), .ZN(
        n14283) );
  MUX2_X1 U16129 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n14283), .S(n14799), .Z(
        P1_U3549) );
  NAND2_X1 U16130 ( .A1(n14256), .A2(n14777), .ZN(n14260) );
  NAND3_X1 U16131 ( .A1(n11513), .A2(n14257), .A3(n14783), .ZN(n14259) );
  NAND4_X1 U16132 ( .A1(n14261), .A2(n14260), .A3(n14259), .A4(n14258), .ZN(
        n14284) );
  MUX2_X1 U16133 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n14284), .S(n14799), .Z(
        P1_U3548) );
  NAND2_X1 U16134 ( .A1(n14262), .A2(n14701), .ZN(n14266) );
  AOI211_X1 U16135 ( .C1(n11899), .C2(n14777), .A(n14264), .B(n14263), .ZN(
        n14265) );
  OAI211_X1 U16136 ( .C1(n14721), .C2(n14267), .A(n14266), .B(n14265), .ZN(
        n14285) );
  MUX2_X1 U16137 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n14285), .S(n14799), .Z(
        P1_U3547) );
  AOI211_X1 U16138 ( .C1(n14270), .C2(n14777), .A(n14269), .B(n14268), .ZN(
        n14271) );
  OAI21_X1 U16139 ( .B1(n14721), .B2(n14272), .A(n14271), .ZN(n14286) );
  MUX2_X1 U16140 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n14286), .S(n14799), .Z(
        P1_U3546) );
  MUX2_X1 U16141 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n14273), .S(n14787), .Z(
        P1_U3527) );
  MUX2_X1 U16142 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n14274), .S(n14787), .Z(
        P1_U3526) );
  MUX2_X1 U16143 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n14276), .S(n14787), .Z(
        P1_U3524) );
  MUX2_X1 U16144 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n14277), .S(n14787), .Z(
        P1_U3523) );
  MUX2_X1 U16145 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n14278), .S(n14787), .Z(
        P1_U3522) );
  MUX2_X1 U16146 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n14279), .S(n14787), .Z(
        P1_U3521) );
  MUX2_X1 U16147 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n14280), .S(n14787), .Z(
        P1_U3520) );
  MUX2_X1 U16148 ( .A(n14281), .B(P1_REG0_REG_23__SCAN_IN), .S(n14785), .Z(
        P1_U3519) );
  MUX2_X1 U16149 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n14282), .S(n14787), .Z(
        P1_U3518) );
  MUX2_X1 U16150 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n14283), .S(n14787), .Z(
        P1_U3517) );
  MUX2_X1 U16151 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n14284), .S(n14787), .Z(
        P1_U3516) );
  MUX2_X1 U16152 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n14285), .S(n14787), .Z(
        P1_U3515) );
  MUX2_X1 U16153 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n14286), .S(n14787), .Z(
        P1_U3513) );
  NOR4_X1 U16154 ( .A1(n14287), .A2(P1_IR_REG_30__SCAN_IN), .A3(n10128), .A4(
        P1_U3086), .ZN(n14288) );
  AOI21_X1 U16155 ( .B1(n14289), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n14288), 
        .ZN(n14290) );
  OAI21_X1 U16156 ( .B1(n14291), .B2(n14296), .A(n14290), .ZN(P1_U3324) );
  OAI222_X1 U16157 ( .A1(n14296), .A2(n14295), .B1(P1_U3086), .B2(n14294), 
        .C1(n14293), .C2(n14292), .ZN(P1_U3326) );
  MUX2_X1 U16158 ( .A(n14298), .B(n14297), .S(P1_STATE_REG_SCAN_IN), .Z(
        P1_U3333) );
  MUX2_X1 U16159 ( .A(n14300), .B(n14299), .S(P1_STATE_REG_SCAN_IN), .Z(
        P1_U3355) );
  AOI21_X1 U16160 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(
        P3_WR_REG_SCAN_IN), .ZN(n14303) );
  OAI21_X1 U16161 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(n14303), 
        .ZN(U28) );
  OAI221_X1 U16162 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .C1(
        n14305), .C2(n7398), .A(n14304), .ZN(U29) );
  AOI21_X1 U16163 ( .B1(n14308), .B2(n14307), .A(n14306), .ZN(n14309) );
  XOR2_X1 U16164 ( .A(n14309), .B(P2_ADDR_REG_2__SCAN_IN), .Z(SUB_1596_U61) );
  AOI22_X1 U16165 ( .A1(n14310), .A2(n14317), .B1(SI_3_), .B2(n14316), .ZN(
        n14311) );
  OAI21_X1 U16166 ( .B1(P3_U3151), .B2(n14312), .A(n14311), .ZN(P3_U3292) );
  AOI22_X1 U16167 ( .A1(n14317), .A2(n14313), .B1(n14316), .B2(SI_2_), .ZN(
        n14314) );
  OAI21_X1 U16168 ( .B1(P3_U3151), .B2(n10088), .A(n14314), .ZN(P3_U3293) );
  INV_X1 U16169 ( .A(n14315), .ZN(n14318) );
  AOI22_X1 U16170 ( .A1(n14318), .A2(n14317), .B1(SI_11_), .B2(n14316), .ZN(
        n14319) );
  OAI21_X1 U16171 ( .B1(P3_U3151), .B2(n14320), .A(n14319), .ZN(P3_U3284) );
  XOR2_X1 U16172 ( .A(n14322), .B(n14321), .Z(SUB_1596_U57) );
  XOR2_X1 U16173 ( .A(n14323), .B(P2_ADDR_REG_8__SCAN_IN), .Z(SUB_1596_U55) );
  OAI21_X1 U16174 ( .B1(n14326), .B2(n14325), .A(n14324), .ZN(n14327) );
  XOR2_X1 U16175 ( .A(n14327), .B(n14852), .Z(SUB_1596_U54) );
  INV_X1 U16176 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n14866) );
  NOR2_X1 U16177 ( .A1(n14329), .A2(n14328), .ZN(n14330) );
  XNOR2_X1 U16178 ( .A(n14866), .B(n14330), .ZN(SUB_1596_U70) );
  OAI211_X1 U16179 ( .C1(n14333), .C2(n14753), .A(n14332), .B(n14331), .ZN(
        n14336) );
  INV_X1 U16180 ( .A(n14334), .ZN(n14335) );
  AOI211_X1 U16181 ( .C1(n14337), .C2(n14783), .A(n14336), .B(n14335), .ZN(
        n14339) );
  INV_X1 U16182 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n14338) );
  AOI22_X1 U16183 ( .A1(n14787), .A2(n14339), .B1(n14338), .B2(n14785), .ZN(
        P1_U3495) );
  AOI22_X1 U16184 ( .A1(n14799), .A2(n14339), .B1(n11409), .B2(n14797), .ZN(
        P1_U3540) );
  OAI21_X1 U16185 ( .B1(n14342), .B2(n14341), .A(n14340), .ZN(n14343) );
  INV_X1 U16186 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n14927) );
  XOR2_X1 U16187 ( .A(n14343), .B(n14927), .Z(SUB_1596_U63) );
  INV_X1 U16188 ( .A(P3_REG3_REG_15__SCAN_IN), .ZN(n14360) );
  AOI22_X1 U16189 ( .A1(n15070), .A2(n14344), .B1(n15094), .B2(
        P3_ADDR_REG_15__SCAN_IN), .ZN(n14359) );
  OAI21_X1 U16190 ( .B1(P3_REG1_REG_15__SCAN_IN), .B2(n14346), .A(n14345), 
        .ZN(n14357) );
  AOI21_X1 U16191 ( .B1(n14349), .B2(n14348), .A(n14347), .ZN(n14350) );
  NOR2_X1 U16192 ( .A1(n14350), .A2(n15090), .ZN(n14356) );
  AOI21_X1 U16193 ( .B1(n14353), .B2(n14351), .A(n14352), .ZN(n14354) );
  NOR2_X1 U16194 ( .A1(n14354), .A2(n15101), .ZN(n14355) );
  AOI211_X1 U16195 ( .C1(n15097), .C2(n14357), .A(n14356), .B(n14355), .ZN(
        n14358) );
  OAI211_X1 U16196 ( .C1(P3_STATE_REG_SCAN_IN), .C2(n14360), .A(n14359), .B(
        n14358), .ZN(P3_U3197) );
  AOI22_X1 U16197 ( .A1(n15070), .A2(n14361), .B1(n15094), .B2(
        P3_ADDR_REG_16__SCAN_IN), .ZN(n14378) );
  INV_X1 U16198 ( .A(n14362), .ZN(n14364) );
  NAND2_X1 U16199 ( .A1(n14364), .A2(n14363), .ZN(n14365) );
  XNOR2_X1 U16200 ( .A(n14366), .B(n14365), .ZN(n14371) );
  OAI21_X1 U16201 ( .B1(n14369), .B2(n14368), .A(n14367), .ZN(n14370) );
  AOI22_X1 U16202 ( .A1(n14371), .A2(n15064), .B1(n15097), .B2(n14370), .ZN(
        n14377) );
  NAND2_X1 U16203 ( .A1(P3_REG3_REG_16__SCAN_IN), .A2(P3_U3151), .ZN(n14376)
         );
  OAI221_X1 U16204 ( .B1(n14374), .B2(n14373), .C1(n14374), .C2(n14372), .A(
        n14404), .ZN(n14375) );
  NAND4_X1 U16205 ( .A1(n14378), .A2(n14377), .A3(n14376), .A4(n14375), .ZN(
        P3_U3198) );
  AOI22_X1 U16206 ( .A1(n15070), .A2(n14379), .B1(n15094), .B2(
        P3_ADDR_REG_17__SCAN_IN), .ZN(n14393) );
  OAI21_X1 U16207 ( .B1(P3_REG1_REG_17__SCAN_IN), .B2(n14381), .A(n14380), 
        .ZN(n14386) );
  AOI211_X1 U16208 ( .C1(n14384), .C2(n14383), .A(n15090), .B(n14382), .ZN(
        n14385) );
  AOI21_X1 U16209 ( .B1(n15097), .B2(n14386), .A(n14385), .ZN(n14392) );
  NAND2_X1 U16210 ( .A1(P3_REG3_REG_17__SCAN_IN), .A2(P3_U3151), .ZN(n14391)
         );
  OAI221_X1 U16211 ( .B1(n14389), .B2(n14388), .C1(n14389), .C2(n14387), .A(
        n14404), .ZN(n14390) );
  NAND4_X1 U16212 ( .A1(n14393), .A2(n14392), .A3(n14391), .A4(n14390), .ZN(
        P3_U3199) );
  AOI22_X1 U16213 ( .A1(n15070), .A2(n14394), .B1(n15094), .B2(
        P3_ADDR_REG_18__SCAN_IN), .ZN(n14411) );
  OAI21_X1 U16214 ( .B1(n14397), .B2(n14396), .A(n14395), .ZN(n14403) );
  AOI21_X1 U16215 ( .B1(n14400), .B2(n14399), .A(n14398), .ZN(n14401) );
  NOR2_X1 U16216 ( .A1(n14401), .A2(n15090), .ZN(n14402) );
  AOI21_X1 U16217 ( .B1(n15097), .B2(n14403), .A(n14402), .ZN(n14410) );
  NAND2_X1 U16218 ( .A1(P3_REG3_REG_18__SCAN_IN), .A2(P3_U3151), .ZN(n14409)
         );
  OAI221_X1 U16219 ( .B1(n14407), .B2(n14406), .C1(n14407), .C2(n14405), .A(
        n14404), .ZN(n14408) );
  OAI21_X1 U16220 ( .B1(n15170), .B2(n14413), .A(n14412), .ZN(n14414) );
  AOI21_X1 U16221 ( .B1(n15167), .B2(n14415), .A(n14414), .ZN(n14433) );
  AOI22_X1 U16222 ( .A1(n15193), .A2(n14433), .B1(n12789), .B2(n15190), .ZN(
        P3_U3473) );
  OAI21_X1 U16223 ( .B1(n15170), .B2(n14417), .A(n14416), .ZN(n14418) );
  AOI21_X1 U16224 ( .B1(n14419), .B2(n15167), .A(n14418), .ZN(n14435) );
  INV_X1 U16225 ( .A(P3_REG1_REG_13__SCAN_IN), .ZN(n14420) );
  AOI22_X1 U16226 ( .A1(n15193), .A2(n14435), .B1(n14420), .B2(n15190), .ZN(
        P3_U3472) );
  NOR2_X1 U16227 ( .A1(n14422), .A2(n14421), .ZN(n14423) );
  AOI211_X1 U16228 ( .C1(n15152), .C2(n14425), .A(n14424), .B(n14423), .ZN(
        n14437) );
  AOI22_X1 U16229 ( .A1(n15193), .A2(n14437), .B1(n14426), .B2(n15190), .ZN(
        P3_U3471) );
  OAI21_X1 U16230 ( .B1(n15170), .B2(n14428), .A(n14427), .ZN(n14429) );
  AOI21_X1 U16231 ( .B1(n15167), .B2(n14430), .A(n14429), .ZN(n14439) );
  INV_X1 U16232 ( .A(P3_REG1_REG_11__SCAN_IN), .ZN(n14431) );
  AOI22_X1 U16233 ( .A1(n15193), .A2(n14439), .B1(n14431), .B2(n15190), .ZN(
        P3_U3470) );
  INV_X1 U16234 ( .A(P3_REG0_REG_14__SCAN_IN), .ZN(n14432) );
  AOI22_X1 U16235 ( .A1(n15177), .A2(n14433), .B1(n14432), .B2(n15175), .ZN(
        P3_U3432) );
  INV_X1 U16236 ( .A(P3_REG0_REG_13__SCAN_IN), .ZN(n14434) );
  AOI22_X1 U16237 ( .A1(n15177), .A2(n14435), .B1(n14434), .B2(n15175), .ZN(
        P3_U3429) );
  INV_X1 U16238 ( .A(P3_REG0_REG_12__SCAN_IN), .ZN(n14436) );
  AOI22_X1 U16239 ( .A1(n15177), .A2(n14437), .B1(n14436), .B2(n15175), .ZN(
        P3_U3426) );
  INV_X1 U16240 ( .A(P3_REG0_REG_11__SCAN_IN), .ZN(n14438) );
  AOI22_X1 U16241 ( .A1(n15177), .A2(n14439), .B1(n14438), .B2(n15175), .ZN(
        P3_U3423) );
  XNOR2_X1 U16242 ( .A(n14441), .B(n14440), .ZN(n14443) );
  AOI222_X1 U16243 ( .A1(n14444), .A2(n14466), .B1(n14465), .B2(n14443), .C1(
        n14442), .C2(n14463), .ZN(n14445) );
  NAND2_X1 U16244 ( .A1(P1_REG3_REG_14__SCAN_IN), .A2(P1_U3086), .ZN(n14614)
         );
  OAI211_X1 U16245 ( .C1(n14469), .C2(n14446), .A(n14445), .B(n14614), .ZN(
        P1_U3215) );
  AND2_X1 U16246 ( .A1(n14448), .A2(n14447), .ZN(n14451) );
  OAI21_X1 U16247 ( .B1(n14451), .B2(n14450), .A(n14449), .ZN(n14452) );
  AOI222_X1 U16248 ( .A1(n14497), .A2(n14466), .B1(n14452), .B2(n14465), .C1(
        n14498), .C2(n14463), .ZN(n14453) );
  NAND2_X1 U16249 ( .A1(P1_REG3_REG_16__SCAN_IN), .A2(P1_U3086), .ZN(n14626)
         );
  OAI211_X1 U16250 ( .C1(n14469), .C2(n14454), .A(n14453), .B(n14626), .ZN(
        P1_U3226) );
  NAND2_X1 U16251 ( .A1(n14456), .A2(n14455), .ZN(n14460) );
  NAND2_X1 U16252 ( .A1(n14458), .A2(n14457), .ZN(n14459) );
  NAND2_X1 U16253 ( .A1(n14460), .A2(n14459), .ZN(n14472) );
  XNOR2_X1 U16254 ( .A(n14462), .B(n14461), .ZN(n14464) );
  AOI222_X1 U16255 ( .A1(n14472), .A2(n14466), .B1(n14465), .B2(n14464), .C1(
        n14477), .C2(n14463), .ZN(n14467) );
  NAND2_X1 U16256 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_U3086), .ZN(n14572)
         );
  OAI211_X1 U16257 ( .C1(n14469), .C2(n14468), .A(n14467), .B(n14572), .ZN(
        P1_U3236) );
  INV_X1 U16258 ( .A(n14470), .ZN(n14471) );
  AOI21_X1 U16259 ( .B1(n14471), .B2(n14479), .A(n14780), .ZN(n14474) );
  AOI21_X1 U16260 ( .B1(n14474), .B2(n14473), .A(n14472), .ZN(n14525) );
  AOI222_X1 U16261 ( .A1(n14477), .A2(n14476), .B1(P1_REG2_REG_11__SCAN_IN), 
        .B2(n14706), .C1(n14475), .C2(n14704), .ZN(n14485) );
  XNOR2_X1 U16262 ( .A(n14478), .B(n14479), .ZN(n14528) );
  OAI211_X1 U16263 ( .C1(n14481), .C2(n14526), .A(n7114), .B(n14480), .ZN(
        n14524) );
  INV_X1 U16264 ( .A(n14524), .ZN(n14482) );
  AOI22_X1 U16265 ( .A1(n14528), .A2(n14483), .B1(n14713), .B2(n14482), .ZN(
        n14484) );
  OAI211_X1 U16266 ( .C1(n14706), .C2(n14525), .A(n14485), .B(n14484), .ZN(
        P1_U3282) );
  NAND3_X1 U16267 ( .A1(n14487), .A2(n14486), .A3(n14701), .ZN(n14491) );
  AOI21_X1 U16268 ( .B1(n14489), .B2(n14777), .A(n14488), .ZN(n14490) );
  OAI211_X1 U16269 ( .C1(n14493), .C2(n14492), .A(n14491), .B(n14490), .ZN(
        n14494) );
  AOI21_X1 U16270 ( .B1(n14495), .B2(n14783), .A(n14494), .ZN(n14530) );
  AOI22_X1 U16271 ( .A1(n14799), .A2(n14530), .B1(n14039), .B2(n14797), .ZN(
        P1_U3545) );
  AOI211_X1 U16272 ( .C1(n14498), .C2(n14777), .A(n14497), .B(n14496), .ZN(
        n14499) );
  OAI21_X1 U16273 ( .B1(n14500), .B2(n14780), .A(n14499), .ZN(n14501) );
  AOI21_X1 U16274 ( .B1(n14502), .B2(n14783), .A(n14501), .ZN(n14532) );
  AOI22_X1 U16275 ( .A1(n14799), .A2(n14532), .B1(n14503), .B2(n14797), .ZN(
        P1_U3544) );
  OAI211_X1 U16276 ( .C1(n14506), .C2(n14753), .A(n14505), .B(n14504), .ZN(
        n14509) );
  INV_X1 U16277 ( .A(n14507), .ZN(n14508) );
  AOI211_X1 U16278 ( .C1(n14783), .C2(n14510), .A(n14509), .B(n14508), .ZN(
        n14534) );
  AOI22_X1 U16279 ( .A1(n14799), .A2(n14534), .B1(n14511), .B2(n14797), .ZN(
        P1_U3543) );
  AND3_X1 U16280 ( .A1(n14513), .A2(n14512), .A3(n14783), .ZN(n14517) );
  OAI21_X1 U16281 ( .B1(n14515), .B2(n14753), .A(n14514), .ZN(n14516) );
  NOR3_X1 U16282 ( .A1(n14518), .A2(n14517), .A3(n14516), .ZN(n14536) );
  AOI22_X1 U16283 ( .A1(n14799), .A2(n14536), .B1(n11408), .B2(n14797), .ZN(
        P1_U3542) );
  OAI211_X1 U16284 ( .C1(n11006), .C2(n14753), .A(n14520), .B(n14519), .ZN(
        n14522) );
  AOI211_X1 U16285 ( .C1(n14523), .C2(n14783), .A(n14522), .B(n14521), .ZN(
        n14538) );
  AOI22_X1 U16286 ( .A1(n14799), .A2(n14538), .B1(n11415), .B2(n14797), .ZN(
        P1_U3541) );
  OAI211_X1 U16287 ( .C1(n14526), .C2(n14753), .A(n14525), .B(n14524), .ZN(
        n14527) );
  AOI21_X1 U16288 ( .B1(n14528), .B2(n14783), .A(n14527), .ZN(n14540) );
  AOI22_X1 U16289 ( .A1(n14799), .A2(n14540), .B1(n11412), .B2(n14797), .ZN(
        P1_U3539) );
  INV_X1 U16290 ( .A(P1_REG0_REG_17__SCAN_IN), .ZN(n14529) );
  AOI22_X1 U16291 ( .A1(n14787), .A2(n14530), .B1(n14529), .B2(n14785), .ZN(
        P1_U3510) );
  INV_X1 U16292 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n14531) );
  AOI22_X1 U16293 ( .A1(n14787), .A2(n14532), .B1(n14531), .B2(n14785), .ZN(
        P1_U3507) );
  INV_X1 U16294 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n14533) );
  AOI22_X1 U16295 ( .A1(n14787), .A2(n14534), .B1(n14533), .B2(n14785), .ZN(
        P1_U3504) );
  INV_X1 U16296 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n14535) );
  AOI22_X1 U16297 ( .A1(n14787), .A2(n14536), .B1(n14535), .B2(n14785), .ZN(
        P1_U3501) );
  INV_X1 U16298 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n14537) );
  AOI22_X1 U16299 ( .A1(n14787), .A2(n14538), .B1(n14537), .B2(n14785), .ZN(
        P1_U3498) );
  INV_X1 U16300 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n14539) );
  AOI22_X1 U16301 ( .A1(n14787), .A2(n14540), .B1(n14539), .B2(n14785), .ZN(
        P1_U3492) );
  AOI21_X1 U16302 ( .B1(n14543), .B2(n14542), .A(n14541), .ZN(n14544) );
  XOR2_X1 U16303 ( .A(n14544), .B(P2_ADDR_REG_11__SCAN_IN), .Z(SUB_1596_U69)
         );
  XNOR2_X1 U16304 ( .A(P2_ADDR_REG_12__SCAN_IN), .B(n14545), .ZN(SUB_1596_U68)
         );
  AOI21_X1 U16305 ( .B1(n14548), .B2(n14547), .A(n14546), .ZN(n14549) );
  XOR2_X1 U16306 ( .A(n14549), .B(P2_ADDR_REG_13__SCAN_IN), .Z(SUB_1596_U67)
         );
  AOI21_X1 U16307 ( .B1(n14552), .B2(n14551), .A(n14550), .ZN(n14553) );
  XOR2_X1 U16308 ( .A(n14553), .B(P2_ADDR_REG_14__SCAN_IN), .Z(SUB_1596_U66)
         );
  AOI21_X1 U16309 ( .B1(n14556), .B2(n14555), .A(n14554), .ZN(n14557) );
  XOR2_X1 U16310 ( .A(n14557), .B(P2_ADDR_REG_15__SCAN_IN), .Z(SUB_1596_U65)
         );
  OAI222_X1 U16311 ( .A1(n14562), .A2(n14561), .B1(n14562), .B2(n14560), .C1(
        n14559), .C2(n14558), .ZN(SUB_1596_U64) );
  OAI21_X1 U16312 ( .B1(n14565), .B2(n14564), .A(n14563), .ZN(n14571) );
  NOR2_X1 U16313 ( .A1(n14642), .A2(n6856), .ZN(n14570) );
  AOI211_X1 U16314 ( .C1(n14568), .C2(n14567), .A(n14651), .B(n14566), .ZN(
        n14569) );
  AOI211_X1 U16315 ( .C1(n14633), .C2(n14571), .A(n14570), .B(n14569), .ZN(
        n14573) );
  OAI211_X1 U16316 ( .C1(n14574), .C2(n14661), .A(n14573), .B(n14572), .ZN(
        P1_U3254) );
  OAI21_X1 U16317 ( .B1(n14577), .B2(n14576), .A(n14575), .ZN(n14583) );
  OAI21_X1 U16318 ( .B1(n14580), .B2(n14579), .A(n14578), .ZN(n14581) );
  AOI222_X1 U16319 ( .A1(n14583), .A2(n14633), .B1(n14582), .B2(n14658), .C1(
        n14581), .C2(n14638), .ZN(n14585) );
  OAI211_X1 U16320 ( .C1(n14586), .C2(n14661), .A(n14585), .B(n14584), .ZN(
        P1_U3255) );
  NAND2_X1 U16321 ( .A1(n14588), .A2(n14587), .ZN(n14591) );
  INV_X1 U16322 ( .A(n14589), .ZN(n14590) );
  NAND3_X1 U16323 ( .A1(n14638), .A2(n14591), .A3(n14590), .ZN(n14597) );
  AOI21_X1 U16324 ( .B1(n14594), .B2(n14593), .A(n14592), .ZN(n14595) );
  NAND2_X1 U16325 ( .A1(n14633), .A2(n14595), .ZN(n14596) );
  OAI211_X1 U16326 ( .C1(n14642), .C2(n14598), .A(n14597), .B(n14596), .ZN(
        n14599) );
  INV_X1 U16327 ( .A(n14599), .ZN(n14601) );
  OAI211_X1 U16328 ( .C1(n14602), .C2(n14661), .A(n14601), .B(n14600), .ZN(
        P1_U3256) );
  OAI211_X1 U16329 ( .C1(n14605), .C2(n14604), .A(n14638), .B(n14603), .ZN(
        n14613) );
  OAI21_X1 U16330 ( .B1(n14608), .B2(n14607), .A(n14606), .ZN(n14609) );
  NAND2_X1 U16331 ( .A1(n14633), .A2(n14609), .ZN(n14612) );
  NAND2_X1 U16332 ( .A1(n14658), .A2(n14610), .ZN(n14611) );
  AND3_X1 U16333 ( .A1(n14613), .A2(n14612), .A3(n14611), .ZN(n14615) );
  OAI211_X1 U16334 ( .C1(n14616), .C2(n14661), .A(n14615), .B(n14614), .ZN(
        P1_U3257) );
  AOI211_X1 U16335 ( .C1(n14619), .C2(n14618), .A(n14617), .B(n14647), .ZN(
        n14624) );
  AOI211_X1 U16336 ( .C1(n14622), .C2(n14621), .A(n14620), .B(n14651), .ZN(
        n14623) );
  AOI211_X1 U16337 ( .C1(n14658), .C2(n14625), .A(n14624), .B(n14623), .ZN(
        n14627) );
  OAI211_X1 U16338 ( .C1(n14628), .C2(n14661), .A(n14627), .B(n14626), .ZN(
        P1_U3259) );
  AOI21_X1 U16339 ( .B1(n14631), .B2(n14630), .A(n14629), .ZN(n14632) );
  NAND2_X1 U16340 ( .A1(n14633), .A2(n14632), .ZN(n14640) );
  AOI21_X1 U16341 ( .B1(n14636), .B2(n14635), .A(n14634), .ZN(n14637) );
  NAND2_X1 U16342 ( .A1(n14638), .A2(n14637), .ZN(n14639) );
  OAI211_X1 U16343 ( .C1(n14642), .C2(n14641), .A(n14640), .B(n14639), .ZN(
        n14643) );
  INV_X1 U16344 ( .A(n14643), .ZN(n14645) );
  OAI211_X1 U16345 ( .C1(n14646), .C2(n14661), .A(n14645), .B(n14644), .ZN(
        P1_U3260) );
  INV_X1 U16346 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n14662) );
  AOI211_X1 U16347 ( .C1(n14650), .C2(n14649), .A(n14648), .B(n14647), .ZN(
        n14656) );
  AOI211_X1 U16348 ( .C1(n14654), .C2(n14653), .A(n14652), .B(n14651), .ZN(
        n14655) );
  AOI211_X1 U16349 ( .C1(n14658), .C2(n14657), .A(n14656), .B(n14655), .ZN(
        n14660) );
  OAI211_X1 U16350 ( .C1(n14662), .C2(n14661), .A(n14660), .B(n14659), .ZN(
        P1_U3261) );
  XNOR2_X1 U16351 ( .A(n14663), .B(n14664), .ZN(n14773) );
  NAND2_X1 U16352 ( .A1(n14665), .A2(n14664), .ZN(n14666) );
  AOI21_X1 U16353 ( .B1(n14667), .B2(n14666), .A(n14780), .ZN(n14771) );
  AOI211_X1 U16354 ( .C1(n14743), .C2(n14773), .A(n14767), .B(n14771), .ZN(
        n14680) );
  INV_X1 U16355 ( .A(n14672), .ZN(n14670) );
  AOI22_X1 U16356 ( .A1(n14681), .A2(P1_REG2_REG_9__SCAN_IN), .B1(n14668), 
        .B2(n14704), .ZN(n14669) );
  OAI21_X1 U16357 ( .B1(n14708), .B2(n14670), .A(n14669), .ZN(n14671) );
  INV_X1 U16358 ( .A(n14671), .ZN(n14679) );
  NAND2_X1 U16359 ( .A1(n14673), .A2(n14672), .ZN(n14674) );
  NAND2_X1 U16360 ( .A1(n14674), .A2(n7114), .ZN(n14675) );
  OR2_X1 U16361 ( .A1(n14676), .A2(n14675), .ZN(n14770) );
  INV_X1 U16362 ( .A(n14770), .ZN(n14677) );
  AOI22_X1 U16363 ( .A1(n14773), .A2(n14714), .B1(n14713), .B2(n14677), .ZN(
        n14678) );
  OAI211_X1 U16364 ( .C1(n14681), .C2(n14680), .A(n14679), .B(n14678), .ZN(
        P1_U3284) );
  XNOR2_X1 U16365 ( .A(n14682), .B(n14687), .ZN(n14758) );
  INV_X1 U16366 ( .A(n14683), .ZN(n14689) );
  INV_X1 U16367 ( .A(n14684), .ZN(n14685) );
  AOI211_X1 U16368 ( .C1(n14687), .C2(n14686), .A(n14780), .B(n14685), .ZN(
        n14688) );
  AOI211_X1 U16369 ( .C1(n14743), .C2(n14758), .A(n14689), .B(n14688), .ZN(
        n14755) );
  AOI22_X1 U16370 ( .A1(n14706), .A2(P1_REG2_REG_7__SCAN_IN), .B1(n14690), 
        .B2(n14704), .ZN(n14691) );
  OAI21_X1 U16371 ( .B1(n14708), .B2(n14754), .A(n14691), .ZN(n14692) );
  INV_X1 U16372 ( .A(n14692), .ZN(n14697) );
  OAI211_X1 U16373 ( .C1(n14694), .C2(n14754), .A(n14693), .B(n7114), .ZN(
        n14752) );
  INV_X1 U16374 ( .A(n14752), .ZN(n14695) );
  AOI22_X1 U16375 ( .A1(n14758), .A2(n14714), .B1(n14713), .B2(n14695), .ZN(
        n14696) );
  OAI211_X1 U16376 ( .C1(n14706), .C2(n14755), .A(n14697), .B(n14696), .ZN(
        P1_U3286) );
  XNOR2_X1 U16377 ( .A(n14698), .B(n14700), .ZN(n14741) );
  XNOR2_X1 U16378 ( .A(n14699), .B(n14700), .ZN(n14702) );
  NAND2_X1 U16379 ( .A1(n14702), .A2(n14701), .ZN(n14739) );
  INV_X1 U16380 ( .A(n14739), .ZN(n14703) );
  AOI211_X1 U16381 ( .C1(n14741), .C2(n14743), .A(n14735), .B(n14703), .ZN(
        n14717) );
  AOI22_X1 U16382 ( .A1(n14706), .A2(P1_REG2_REG_5__SCAN_IN), .B1(n14705), 
        .B2(n14704), .ZN(n14707) );
  OAI21_X1 U16383 ( .B1(n14708), .B2(n6904), .A(n14707), .ZN(n14709) );
  INV_X1 U16384 ( .A(n14709), .ZN(n14716) );
  OAI211_X1 U16385 ( .C1(n6905), .C2(n6904), .A(n7114), .B(n14711), .ZN(n14736) );
  INV_X1 U16386 ( .A(n14736), .ZN(n14712) );
  AOI22_X1 U16387 ( .A1(n14741), .A2(n14714), .B1(n14713), .B2(n14712), .ZN(
        n14715) );
  OAI211_X1 U16388 ( .C1(n14706), .C2(n14717), .A(n14716), .B(n14715), .ZN(
        P1_U3288) );
  AND2_X1 U16389 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n14718), .ZN(P1_U3294) );
  AND2_X1 U16390 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n14718), .ZN(P1_U3295) );
  AND2_X1 U16391 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n14718), .ZN(P1_U3296) );
  AND2_X1 U16392 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n14718), .ZN(P1_U3297) );
  AND2_X1 U16393 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n14718), .ZN(P1_U3298) );
  AND2_X1 U16394 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n14718), .ZN(P1_U3299) );
  AND2_X1 U16395 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n14718), .ZN(P1_U3300) );
  AND2_X1 U16396 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n14718), .ZN(P1_U3301) );
  AND2_X1 U16397 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n14718), .ZN(P1_U3302) );
  AND2_X1 U16398 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n14718), .ZN(P1_U3303) );
  AND2_X1 U16399 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n14718), .ZN(P1_U3304) );
  AND2_X1 U16400 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n14718), .ZN(P1_U3305) );
  AND2_X1 U16401 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n14718), .ZN(P1_U3306) );
  AND2_X1 U16402 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n14718), .ZN(P1_U3307) );
  AND2_X1 U16403 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n14718), .ZN(P1_U3308) );
  AND2_X1 U16404 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n14718), .ZN(P1_U3309) );
  AND2_X1 U16405 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n14718), .ZN(P1_U3310) );
  AND2_X1 U16406 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n14718), .ZN(P1_U3311) );
  AND2_X1 U16407 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n14718), .ZN(P1_U3312) );
  AND2_X1 U16408 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n14718), .ZN(P1_U3313) );
  AND2_X1 U16409 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n14718), .ZN(P1_U3314) );
  AND2_X1 U16410 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n14718), .ZN(P1_U3315) );
  AND2_X1 U16411 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n14718), .ZN(P1_U3316) );
  AND2_X1 U16412 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n14718), .ZN(P1_U3317) );
  AND2_X1 U16413 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n14718), .ZN(P1_U3318) );
  AND2_X1 U16414 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n14718), .ZN(P1_U3319) );
  AND2_X1 U16415 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n14718), .ZN(P1_U3320) );
  AND2_X1 U16416 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n14718), .ZN(P1_U3321) );
  AND2_X1 U16417 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n14718), .ZN(P1_U3322) );
  AND2_X1 U16418 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n14718), .ZN(P1_U3323) );
  INV_X1 U16419 ( .A(n14719), .ZN(n14723) );
  AOI21_X1 U16420 ( .B1(n14780), .B2(n14721), .A(n14720), .ZN(n14722) );
  AOI211_X1 U16421 ( .C1(n14725), .C2(n14724), .A(n14723), .B(n14722), .ZN(
        n14788) );
  INV_X1 U16422 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n14726) );
  AOI22_X1 U16423 ( .A1(n14787), .A2(n14788), .B1(n14726), .B2(n14785), .ZN(
        P1_U3459) );
  AOI21_X1 U16424 ( .B1(n14728), .B2(n14777), .A(n14727), .ZN(n14729) );
  OAI21_X1 U16425 ( .B1(n14731), .B2(n14730), .A(n14729), .ZN(n14732) );
  NOR2_X1 U16426 ( .A1(n14733), .A2(n14732), .ZN(n14790) );
  INV_X1 U16427 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n14734) );
  AOI22_X1 U16428 ( .A1(n14787), .A2(n14790), .B1(n14734), .B2(n14785), .ZN(
        P1_U3465) );
  INV_X1 U16429 ( .A(n14735), .ZN(n14738) );
  NAND4_X1 U16430 ( .A1(n14739), .A2(n14738), .A3(n14737), .A4(n14736), .ZN(
        n14740) );
  AOI21_X1 U16431 ( .B1(n14741), .B2(n14783), .A(n14740), .ZN(n14791) );
  INV_X1 U16432 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n14742) );
  AOI22_X1 U16433 ( .A1(n14787), .A2(n14791), .B1(n14742), .B2(n14785), .ZN(
        P1_U3474) );
  NAND2_X1 U16434 ( .A1(n14750), .A2(n14743), .ZN(n14748) );
  INV_X1 U16435 ( .A(n14744), .ZN(n14746) );
  NAND4_X1 U16436 ( .A1(n14748), .A2(n14747), .A3(n14746), .A4(n14745), .ZN(
        n14749) );
  AOI21_X1 U16437 ( .B1(n14759), .B2(n14750), .A(n14749), .ZN(n14792) );
  INV_X1 U16438 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n14751) );
  AOI22_X1 U16439 ( .A1(n14787), .A2(n14792), .B1(n14751), .B2(n14785), .ZN(
        P1_U3477) );
  OAI21_X1 U16440 ( .B1(n14754), .B2(n14753), .A(n14752), .ZN(n14757) );
  INV_X1 U16441 ( .A(n14755), .ZN(n14756) );
  AOI211_X1 U16442 ( .C1(n14759), .C2(n14758), .A(n14757), .B(n14756), .ZN(
        n14793) );
  INV_X1 U16443 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n14760) );
  AOI22_X1 U16444 ( .A1(n14787), .A2(n14793), .B1(n14760), .B2(n14785), .ZN(
        P1_U3480) );
  NAND3_X1 U16445 ( .A1(n14763), .A2(n14762), .A3(n14761), .ZN(n14764) );
  AOI21_X1 U16446 ( .B1(n14765), .B2(n14783), .A(n14764), .ZN(n14794) );
  INV_X1 U16447 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n14766) );
  AOI22_X1 U16448 ( .A1(n14787), .A2(n14794), .B1(n14766), .B2(n14785), .ZN(
        P1_U3483) );
  NOR2_X1 U16449 ( .A1(n14768), .A2(n14767), .ZN(n14769) );
  NAND2_X1 U16450 ( .A1(n14770), .A2(n14769), .ZN(n14772) );
  AOI211_X1 U16451 ( .C1(n14773), .C2(n14783), .A(n14772), .B(n14771), .ZN(
        n14796) );
  INV_X1 U16452 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n14774) );
  AOI22_X1 U16453 ( .A1(n14787), .A2(n14796), .B1(n14774), .B2(n14785), .ZN(
        P1_U3486) );
  AOI211_X1 U16454 ( .C1(n14778), .C2(n14777), .A(n14776), .B(n14775), .ZN(
        n14779) );
  OAI21_X1 U16455 ( .B1(n14781), .B2(n14780), .A(n14779), .ZN(n14782) );
  AOI21_X1 U16456 ( .B1(n14784), .B2(n14783), .A(n14782), .ZN(n14798) );
  INV_X1 U16457 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n14786) );
  AOI22_X1 U16458 ( .A1(n14787), .A2(n14798), .B1(n14786), .B2(n14785), .ZN(
        P1_U3489) );
  AOI22_X1 U16459 ( .A1(n14799), .A2(n14788), .B1(n9507), .B2(n14797), .ZN(
        P1_U3528) );
  AOI22_X1 U16460 ( .A1(n14799), .A2(n14790), .B1(n14789), .B2(n14797), .ZN(
        P1_U3530) );
  AOI22_X1 U16461 ( .A1(n14799), .A2(n14791), .B1(n9602), .B2(n14797), .ZN(
        P1_U3533) );
  AOI22_X1 U16462 ( .A1(n14799), .A2(n14792), .B1(n6868), .B2(n14797), .ZN(
        P1_U3534) );
  AOI22_X1 U16463 ( .A1(n14799), .A2(n14793), .B1(n9687), .B2(n14797), .ZN(
        P1_U3535) );
  AOI22_X1 U16464 ( .A1(n14799), .A2(n14794), .B1(n9970), .B2(n14797), .ZN(
        P1_U3536) );
  INV_X1 U16465 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n14795) );
  AOI22_X1 U16466 ( .A1(n14799), .A2(n14796), .B1(n14795), .B2(n14797), .ZN(
        P1_U3537) );
  AOI22_X1 U16467 ( .A1(n14799), .A2(n14798), .B1(n10533), .B2(n14797), .ZN(
        P1_U3538) );
  NOR2_X1 U16468 ( .A1(n14800), .A2(P2_U3947), .ZN(P2_U3087) );
  AOI22_X1 U16469 ( .A1(n14800), .A2(P2_ADDR_REG_2__SCAN_IN), .B1(
        P2_REG3_REG_2__SCAN_IN), .B2(P2_U3088), .ZN(n14812) );
  OAI211_X1 U16470 ( .C1(n14803), .C2(n14802), .A(n14913), .B(n14801), .ZN(
        n14810) );
  OAI211_X1 U16471 ( .C1(n14806), .C2(n14805), .A(n14918), .B(n14804), .ZN(
        n14809) );
  NAND2_X1 U16472 ( .A1(n14890), .A2(n14807), .ZN(n14808) );
  AND3_X1 U16473 ( .A1(n14810), .A2(n14809), .A3(n14808), .ZN(n14811) );
  NAND2_X1 U16474 ( .A1(n14812), .A2(n14811), .ZN(P2_U3216) );
  INV_X1 U16475 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n15197) );
  OAI211_X1 U16476 ( .C1(n14815), .C2(n14814), .A(n14918), .B(n14813), .ZN(
        n14822) );
  OAI211_X1 U16477 ( .C1(n14818), .C2(n14817), .A(n14913), .B(n14816), .ZN(
        n14821) );
  NAND2_X1 U16478 ( .A1(n14890), .A2(n14819), .ZN(n14820) );
  AND3_X1 U16479 ( .A1(n14822), .A2(n14821), .A3(n14820), .ZN(n14824) );
  OAI211_X1 U16480 ( .C1(n14926), .C2(n15197), .A(n14824), .B(n14823), .ZN(
        P2_U3219) );
  INV_X1 U16481 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n14837) );
  OAI211_X1 U16482 ( .C1(n14827), .C2(n14826), .A(n14918), .B(n14825), .ZN(
        n14832) );
  OAI211_X1 U16483 ( .C1(n14830), .C2(n14829), .A(n14913), .B(n14828), .ZN(
        n14831) );
  OAI211_X1 U16484 ( .C1(n14922), .C2(n14833), .A(n14832), .B(n14831), .ZN(
        n14834) );
  INV_X1 U16485 ( .A(n14834), .ZN(n14836) );
  OAI211_X1 U16486 ( .C1(n14837), .C2(n14926), .A(n14836), .B(n14835), .ZN(
        P2_U3222) );
  AND2_X1 U16487 ( .A1(n14839), .A2(n14838), .ZN(n14840) );
  OAI21_X1 U16488 ( .B1(n14841), .B2(n14840), .A(n14913), .ZN(n14849) );
  AND2_X1 U16489 ( .A1(n14843), .A2(n14842), .ZN(n14844) );
  OAI21_X1 U16490 ( .B1(n14845), .B2(n14844), .A(n14918), .ZN(n14848) );
  NAND2_X1 U16491 ( .A1(n14890), .A2(n14846), .ZN(n14847) );
  AND3_X1 U16492 ( .A1(n14849), .A2(n14848), .A3(n14847), .ZN(n14851) );
  OAI211_X1 U16493 ( .C1(n14852), .C2(n14926), .A(n14851), .B(n14850), .ZN(
        P2_U3223) );
  OAI21_X1 U16494 ( .B1(n14854), .B2(n14853), .A(n14918), .ZN(n14856) );
  NOR2_X1 U16495 ( .A1(n14856), .A2(n14855), .ZN(n14862) );
  OAI21_X1 U16496 ( .B1(n14858), .B2(n14857), .A(n14913), .ZN(n14860) );
  NOR2_X1 U16497 ( .A1(n14860), .A2(n14859), .ZN(n14861) );
  AOI211_X1 U16498 ( .C1(n14890), .C2(n14863), .A(n14862), .B(n14861), .ZN(
        n14865) );
  OAI211_X1 U16499 ( .C1(n14866), .C2(n14926), .A(n14865), .B(n14864), .ZN(
        P2_U3224) );
  AOI211_X1 U16500 ( .C1(n14869), .C2(n14868), .A(n14880), .B(n14867), .ZN(
        n14874) );
  AOI211_X1 U16501 ( .C1(n14872), .C2(n14871), .A(n14884), .B(n14870), .ZN(
        n14873) );
  AOI211_X1 U16502 ( .C1(n14890), .C2(n14875), .A(n14874), .B(n14873), .ZN(
        n14877) );
  NAND2_X1 U16503 ( .A1(P2_REG3_REG_13__SCAN_IN), .A2(P2_U3088), .ZN(n14876)
         );
  OAI211_X1 U16504 ( .C1(n14878), .C2(n14926), .A(n14877), .B(n14876), .ZN(
        P2_U3227) );
  AOI211_X1 U16505 ( .C1(n14882), .C2(n14881), .A(n14880), .B(n14879), .ZN(
        n14888) );
  AOI211_X1 U16506 ( .C1(n14886), .C2(n14885), .A(n14884), .B(n14883), .ZN(
        n14887) );
  AOI211_X1 U16507 ( .C1(n14890), .C2(n14889), .A(n14888), .B(n14887), .ZN(
        n14892) );
  OAI211_X1 U16508 ( .C1(n14893), .C2(n14926), .A(n14892), .B(n14891), .ZN(
        P2_U3228) );
  AOI21_X1 U16509 ( .B1(n14896), .B2(n14895), .A(n14894), .ZN(n14897) );
  NAND2_X1 U16510 ( .A1(n14913), .A2(n14897), .ZN(n14903) );
  AOI21_X1 U16511 ( .B1(n14900), .B2(n14899), .A(n14898), .ZN(n14901) );
  NAND2_X1 U16512 ( .A1(n14918), .A2(n14901), .ZN(n14902) );
  OAI211_X1 U16513 ( .C1(n14922), .C2(n14904), .A(n14903), .B(n14902), .ZN(
        n14905) );
  INV_X1 U16514 ( .A(n14905), .ZN(n14907) );
  NAND2_X1 U16515 ( .A1(P2_REG3_REG_15__SCAN_IN), .A2(P2_U3088), .ZN(n14906)
         );
  OAI211_X1 U16516 ( .C1(n14908), .C2(n14926), .A(n14907), .B(n14906), .ZN(
        P2_U3229) );
  AOI21_X1 U16517 ( .B1(n14911), .B2(n14910), .A(n14909), .ZN(n14912) );
  NAND2_X1 U16518 ( .A1(n14913), .A2(n14912), .ZN(n14920) );
  AOI21_X1 U16519 ( .B1(n14916), .B2(n14915), .A(n14914), .ZN(n14917) );
  NAND2_X1 U16520 ( .A1(n14918), .A2(n14917), .ZN(n14919) );
  OAI211_X1 U16521 ( .C1(n14922), .C2(n14921), .A(n14920), .B(n14919), .ZN(
        n14923) );
  INV_X1 U16522 ( .A(n14923), .ZN(n14925) );
  NAND2_X1 U16523 ( .A1(P2_REG3_REG_17__SCAN_IN), .A2(P2_U3088), .ZN(n14924)
         );
  OAI211_X1 U16524 ( .C1(n14927), .C2(n14926), .A(n14925), .B(n14924), .ZN(
        P2_U3231) );
  AND2_X1 U16525 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n14929), .ZN(P2_U3266) );
  AND2_X1 U16526 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n14929), .ZN(P2_U3267) );
  AND2_X1 U16527 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n14929), .ZN(P2_U3268) );
  AND2_X1 U16528 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n14929), .ZN(P2_U3269) );
  AND2_X1 U16529 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n14929), .ZN(P2_U3270) );
  AND2_X1 U16530 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n14929), .ZN(P2_U3271) );
  AND2_X1 U16531 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n14929), .ZN(P2_U3272) );
  AND2_X1 U16532 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n14929), .ZN(P2_U3273) );
  AND2_X1 U16533 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n14929), .ZN(P2_U3274) );
  AND2_X1 U16534 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n14929), .ZN(P2_U3275) );
  AND2_X1 U16535 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n14929), .ZN(P2_U3276) );
  AND2_X1 U16536 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n14929), .ZN(P2_U3277) );
  AND2_X1 U16537 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n14929), .ZN(P2_U3278) );
  AND2_X1 U16538 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n14929), .ZN(P2_U3279) );
  AND2_X1 U16539 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n14929), .ZN(P2_U3280) );
  AND2_X1 U16540 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n14929), .ZN(P2_U3281) );
  AND2_X1 U16541 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n14929), .ZN(P2_U3282) );
  AND2_X1 U16542 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n14929), .ZN(P2_U3283) );
  AND2_X1 U16543 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n14929), .ZN(P2_U3284) );
  AND2_X1 U16544 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n14929), .ZN(P2_U3285) );
  AND2_X1 U16545 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n14929), .ZN(P2_U3286) );
  AND2_X1 U16546 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n14929), .ZN(P2_U3287) );
  AND2_X1 U16547 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n14929), .ZN(P2_U3288) );
  AND2_X1 U16548 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n14929), .ZN(P2_U3289) );
  AND2_X1 U16549 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n14929), .ZN(P2_U3290) );
  AND2_X1 U16550 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n14929), .ZN(P2_U3291) );
  AND2_X1 U16551 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n14929), .ZN(P2_U3292) );
  AND2_X1 U16552 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n14929), .ZN(P2_U3293) );
  AND2_X1 U16553 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n14929), .ZN(P2_U3294) );
  AND2_X1 U16554 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n14929), .ZN(P2_U3295) );
  AOI22_X1 U16555 ( .A1(n14932), .A2(n14931), .B1(n14930), .B2(n14934), .ZN(
        P2_U3416) );
  AOI21_X1 U16556 ( .B1(n14935), .B2(n14934), .A(n14933), .ZN(P2_U3417) );
  INV_X1 U16557 ( .A(n14936), .ZN(n14943) );
  INV_X1 U16558 ( .A(n14937), .ZN(n14975) );
  NOR3_X1 U16559 ( .A1(n14940), .A2(n14939), .A3(n14938), .ZN(n14942) );
  AOI211_X1 U16560 ( .C1(n14943), .C2(n14975), .A(n14942), .B(n14941), .ZN(
        n15005) );
  INV_X1 U16561 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n14944) );
  AOI22_X1 U16562 ( .A1(n14953), .A2(n15005), .B1(n14944), .B2(n15002), .ZN(
        P2_U3430) );
  NAND2_X1 U16563 ( .A1(n14945), .A2(n15000), .ZN(n14951) );
  AOI22_X1 U16564 ( .A1(n14948), .A2(n14988), .B1(n14947), .B2(n14986), .ZN(
        n14949) );
  AND3_X1 U16565 ( .A1(n14951), .A2(n14950), .A3(n14949), .ZN(n15006) );
  INV_X1 U16566 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n14952) );
  AOI22_X1 U16567 ( .A1(n14953), .A2(n15006), .B1(n14952), .B2(n15002), .ZN(
        P2_U3445) );
  OAI22_X1 U16568 ( .A1(n14955), .A2(n14996), .B1(n14954), .B2(n14994), .ZN(
        n14958) );
  INV_X1 U16569 ( .A(n14956), .ZN(n14957) );
  AOI211_X1 U16570 ( .C1(n14975), .C2(n14959), .A(n14958), .B(n14957), .ZN(
        n15008) );
  INV_X1 U16571 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n14960) );
  AOI22_X1 U16572 ( .A1(n15004), .A2(n15008), .B1(n14960), .B2(n15002), .ZN(
        P2_U3448) );
  INV_X1 U16573 ( .A(n14961), .ZN(n14966) );
  OAI22_X1 U16574 ( .A1(n14963), .A2(n14996), .B1(n14962), .B2(n14994), .ZN(
        n14965) );
  AOI211_X1 U16575 ( .C1(n14966), .C2(n15000), .A(n14965), .B(n14964), .ZN(
        n15010) );
  INV_X1 U16576 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n14967) );
  AOI22_X1 U16577 ( .A1(n15004), .A2(n15010), .B1(n14967), .B2(n15002), .ZN(
        P2_U3451) );
  INV_X1 U16578 ( .A(n14968), .ZN(n14974) );
  INV_X1 U16579 ( .A(n14969), .ZN(n14971) );
  OAI22_X1 U16580 ( .A1(n14971), .A2(n14996), .B1(n14970), .B2(n14994), .ZN(
        n14973) );
  AOI211_X1 U16581 ( .C1(n14975), .C2(n14974), .A(n14973), .B(n14972), .ZN(
        n15012) );
  INV_X1 U16582 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n14976) );
  AOI22_X1 U16583 ( .A1(n15004), .A2(n15012), .B1(n14976), .B2(n15002), .ZN(
        P2_U3454) );
  INV_X1 U16584 ( .A(n14977), .ZN(n14982) );
  OAI22_X1 U16585 ( .A1(n14979), .A2(n14996), .B1(n14978), .B2(n14994), .ZN(
        n14981) );
  AOI211_X1 U16586 ( .C1(n14982), .C2(n15000), .A(n14981), .B(n14980), .ZN(
        n15014) );
  INV_X1 U16587 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n14983) );
  AOI22_X1 U16588 ( .A1(n15004), .A2(n15014), .B1(n14983), .B2(n15002), .ZN(
        P2_U3457) );
  OR2_X1 U16589 ( .A1(n14985), .A2(n14984), .ZN(n14992) );
  AOI22_X1 U16590 ( .A1(n14989), .A2(n14988), .B1(n14987), .B2(n14986), .ZN(
        n14990) );
  INV_X1 U16591 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n14993) );
  AOI22_X1 U16592 ( .A1(n15004), .A2(n15016), .B1(n14993), .B2(n15002), .ZN(
        P2_U3460) );
  OAI22_X1 U16593 ( .A1(n14997), .A2(n14996), .B1(n14995), .B2(n14994), .ZN(
        n14998) );
  AOI211_X1 U16594 ( .C1(n15001), .C2(n15000), .A(n14999), .B(n14998), .ZN(
        n15018) );
  INV_X1 U16595 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n15003) );
  AOI22_X1 U16596 ( .A1(n15004), .A2(n15018), .B1(n15003), .B2(n15002), .ZN(
        P2_U3463) );
  AOI22_X1 U16597 ( .A1(n15019), .A2(n15005), .B1(n9646), .B2(n15017), .ZN(
        P2_U3499) );
  AOI22_X1 U16598 ( .A1(n15019), .A2(n15006), .B1(n9731), .B2(n15017), .ZN(
        P2_U3504) );
  AOI22_X1 U16599 ( .A1(n15019), .A2(n15008), .B1(n15007), .B2(n15017), .ZN(
        P2_U3505) );
  AOI22_X1 U16600 ( .A1(n15019), .A2(n15010), .B1(n15009), .B2(n15017), .ZN(
        P2_U3506) );
  AOI22_X1 U16601 ( .A1(n15019), .A2(n15012), .B1(n15011), .B2(n15017), .ZN(
        P2_U3507) );
  AOI22_X1 U16602 ( .A1(n15019), .A2(n15014), .B1(n15013), .B2(n15017), .ZN(
        P2_U3508) );
  AOI22_X1 U16603 ( .A1(n15019), .A2(n15016), .B1(n15015), .B2(n15017), .ZN(
        P2_U3509) );
  AOI22_X1 U16604 ( .A1(n15019), .A2(n15018), .B1(n9739), .B2(n15017), .ZN(
        P2_U3510) );
  NOR2_X1 U16605 ( .A1(P3_U3897), .A2(n15094), .ZN(P3_U3150) );
  AOI21_X1 U16606 ( .B1(n15021), .B2(n10062), .A(n15020), .ZN(n15026) );
  OAI21_X1 U16607 ( .B1(P3_REG1_REG_3__SCAN_IN), .B2(n15023), .A(n15022), .ZN(
        n15024) );
  NAND2_X1 U16608 ( .A1(n15097), .A2(n15024), .ZN(n15025) );
  OAI21_X1 U16609 ( .B1(n15101), .B2(n15026), .A(n15025), .ZN(n15034) );
  INV_X1 U16610 ( .A(n15027), .ZN(n15028) );
  NAND3_X1 U16611 ( .A1(n15030), .A2(n15029), .A3(n15028), .ZN(n15031) );
  AOI21_X1 U16612 ( .B1(n15032), .B2(n15031), .A(n15090), .ZN(n15033) );
  AOI211_X1 U16613 ( .C1(n15070), .C2(n15035), .A(n15034), .B(n15033), .ZN(
        n15037) );
  NAND2_X1 U16614 ( .A1(P3_REG3_REG_3__SCAN_IN), .A2(P3_U3151), .ZN(n15036) );
  OAI211_X1 U16615 ( .C1(n7090), .C2(n15077), .A(n15037), .B(n15036), .ZN(
        P3_U3185) );
  OAI21_X1 U16616 ( .B1(n15040), .B2(n15039), .A(n15038), .ZN(n15053) );
  OAI21_X1 U16617 ( .B1(n15043), .B2(n15042), .A(n15041), .ZN(n15049) );
  AOI21_X1 U16618 ( .B1(n15046), .B2(n15045), .A(n15044), .ZN(n15047) );
  NOR2_X1 U16619 ( .A1(n15101), .A2(n15047), .ZN(n15048) );
  AOI21_X1 U16620 ( .B1(n15097), .B2(n15049), .A(n15048), .ZN(n15050) );
  OAI21_X1 U16621 ( .B1(n15051), .B2(n15088), .A(n15050), .ZN(n15052) );
  AOI21_X1 U16622 ( .B1(n15064), .B2(n15053), .A(n15052), .ZN(n15055) );
  NAND2_X1 U16623 ( .A1(P3_REG3_REG_4__SCAN_IN), .A2(P3_U3151), .ZN(n15054) );
  OAI211_X1 U16624 ( .C1(n15056), .C2(n15077), .A(n15055), .B(n15054), .ZN(
        P3_U3186) );
  AOI21_X1 U16625 ( .B1(n15058), .B2(n10072), .A(n15057), .ZN(n15073) );
  INV_X1 U16626 ( .A(n15059), .ZN(n15061) );
  NOR2_X1 U16627 ( .A1(n15061), .A2(n15060), .ZN(n15062) );
  XNOR2_X1 U16628 ( .A(n15063), .B(n15062), .ZN(n15065) );
  NAND2_X1 U16629 ( .A1(n15065), .A2(n15064), .ZN(n15072) );
  OAI21_X1 U16630 ( .B1(P3_REG1_REG_5__SCAN_IN), .B2(n15067), .A(n15066), .ZN(
        n15068) );
  AOI22_X1 U16631 ( .A1(n15070), .A2(n15069), .B1(n15097), .B2(n15068), .ZN(
        n15071) );
  OAI211_X1 U16632 ( .C1(n15073), .C2(n15101), .A(n15072), .B(n15071), .ZN(
        n15074) );
  INV_X1 U16633 ( .A(n15074), .ZN(n15076) );
  NAND2_X1 U16634 ( .A1(P3_REG3_REG_5__SCAN_IN), .A2(P3_U3151), .ZN(n15075) );
  OAI211_X1 U16635 ( .C1(n15078), .C2(n15077), .A(n15076), .B(n15075), .ZN(
        P3_U3187) );
  AOI21_X1 U16636 ( .B1(n15081), .B2(n15080), .A(n15079), .ZN(n15102) );
  NOR2_X1 U16637 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n7540), .ZN(n15093) );
  INV_X1 U16638 ( .A(n15082), .ZN(n15087) );
  AOI21_X1 U16639 ( .B1(n15084), .B2(n15086), .A(n15083), .ZN(n15085) );
  AOI21_X1 U16640 ( .B1(n15087), .B2(n15086), .A(n15085), .ZN(n15091) );
  OAI22_X1 U16641 ( .A1(n15091), .A2(n15090), .B1(n15089), .B2(n15088), .ZN(
        n15092) );
  AOI211_X1 U16642 ( .C1(P3_ADDR_REG_9__SCAN_IN), .C2(n15094), .A(n15093), .B(
        n15092), .ZN(n15100) );
  OAI21_X1 U16643 ( .B1(P3_REG1_REG_9__SCAN_IN), .B2(n15096), .A(n15095), .ZN(
        n15098) );
  NAND2_X1 U16644 ( .A1(n15098), .A2(n15097), .ZN(n15099) );
  OAI211_X1 U16645 ( .C1(n15102), .C2(n15101), .A(n15100), .B(n15099), .ZN(
        P3_U3191) );
  OAI21_X1 U16646 ( .B1(n15104), .B2(n12556), .A(n15103), .ZN(n15131) );
  INV_X1 U16647 ( .A(n15105), .ZN(n15106) );
  OAI22_X1 U16648 ( .A1(n7389), .A2(n15108), .B1(n15107), .B2(n15106), .ZN(
        n15122) );
  OAI22_X1 U16649 ( .A1(n15112), .A2(n15111), .B1(n15110), .B2(n15109), .ZN(
        n15119) );
  NAND3_X1 U16650 ( .A1(n15114), .A2(n12556), .A3(n15113), .ZN(n15116) );
  AOI21_X1 U16651 ( .B1(n15117), .B2(n15116), .A(n15115), .ZN(n15118) );
  AOI211_X1 U16652 ( .C1(n15120), .C2(n15131), .A(n15119), .B(n15118), .ZN(
        n15133) );
  INV_X1 U16653 ( .A(n15133), .ZN(n15121) );
  AOI211_X1 U16654 ( .C1(n15123), .C2(n15131), .A(n15122), .B(n15121), .ZN(
        n15124) );
  AOI22_X1 U16655 ( .A1(n13116), .A2(n10056), .B1(n15124), .B2(n13106), .ZN(
        P3_U3231) );
  OAI22_X1 U16656 ( .A1(n15126), .A2(n15171), .B1(n15125), .B2(n15170), .ZN(
        n15127) );
  NOR2_X1 U16657 ( .A1(n15128), .A2(n15127), .ZN(n15178) );
  INV_X1 U16658 ( .A(P3_REG0_REG_1__SCAN_IN), .ZN(n15129) );
  AOI22_X1 U16659 ( .A1(n15177), .A2(n15178), .B1(n15129), .B2(n15175), .ZN(
        P3_U3393) );
  AOI22_X1 U16660 ( .A1(n15131), .A2(n15161), .B1(n15152), .B2(n15130), .ZN(
        n15132) );
  AND2_X1 U16661 ( .A1(n15133), .A2(n15132), .ZN(n15179) );
  INV_X1 U16662 ( .A(P3_REG0_REG_2__SCAN_IN), .ZN(n15134) );
  AOI22_X1 U16663 ( .A1(n15177), .A2(n15179), .B1(n15134), .B2(n15175), .ZN(
        P3_U3396) );
  NOR2_X1 U16664 ( .A1(n15135), .A2(n15170), .ZN(n15137) );
  AOI211_X1 U16665 ( .C1(n15161), .C2(n15138), .A(n15137), .B(n15136), .ZN(
        n15180) );
  INV_X1 U16666 ( .A(P3_REG0_REG_3__SCAN_IN), .ZN(n15139) );
  AOI22_X1 U16667 ( .A1(n15177), .A2(n15180), .B1(n15139), .B2(n15175), .ZN(
        P3_U3399) );
  NOR2_X1 U16668 ( .A1(n15140), .A2(n15170), .ZN(n15142) );
  AOI211_X1 U16669 ( .C1(n15161), .C2(n15143), .A(n15142), .B(n15141), .ZN(
        n15182) );
  INV_X1 U16670 ( .A(P3_REG0_REG_4__SCAN_IN), .ZN(n15144) );
  AOI22_X1 U16671 ( .A1(n15177), .A2(n15182), .B1(n15144), .B2(n15175), .ZN(
        P3_U3402) );
  INV_X1 U16672 ( .A(n15145), .ZN(n15147) );
  OAI22_X1 U16673 ( .A1(n15147), .A2(n15171), .B1(n15170), .B2(n15146), .ZN(
        n15148) );
  NOR2_X1 U16674 ( .A1(n15149), .A2(n15148), .ZN(n15183) );
  INV_X1 U16675 ( .A(P3_REG0_REG_5__SCAN_IN), .ZN(n15150) );
  AOI22_X1 U16676 ( .A1(n15177), .A2(n15183), .B1(n15150), .B2(n15175), .ZN(
        P3_U3405) );
  AOI22_X1 U16677 ( .A1(n15153), .A2(n15161), .B1(n15152), .B2(n15151), .ZN(
        n15154) );
  AND2_X1 U16678 ( .A1(n15155), .A2(n15154), .ZN(n15185) );
  INV_X1 U16679 ( .A(P3_REG0_REG_6__SCAN_IN), .ZN(n15156) );
  AOI22_X1 U16680 ( .A1(n15177), .A2(n15185), .B1(n15156), .B2(n15175), .ZN(
        P3_U3408) );
  NOR2_X1 U16681 ( .A1(n15157), .A2(n15170), .ZN(n15159) );
  AOI211_X1 U16682 ( .C1(n15161), .C2(n15160), .A(n15159), .B(n15158), .ZN(
        n15187) );
  INV_X1 U16683 ( .A(P3_REG0_REG_7__SCAN_IN), .ZN(n15162) );
  AOI22_X1 U16684 ( .A1(n15177), .A2(n15187), .B1(n15162), .B2(n15175), .ZN(
        P3_U3411) );
  NOR2_X1 U16685 ( .A1(n15163), .A2(n15170), .ZN(n15165) );
  AOI211_X1 U16686 ( .C1(n15167), .C2(n15166), .A(n15165), .B(n15164), .ZN(
        n15189) );
  INV_X1 U16687 ( .A(P3_REG0_REG_8__SCAN_IN), .ZN(n15168) );
  AOI22_X1 U16688 ( .A1(n15177), .A2(n15189), .B1(n15168), .B2(n15175), .ZN(
        P3_U3414) );
  OAI22_X1 U16689 ( .A1(n15172), .A2(n15171), .B1(n15170), .B2(n15169), .ZN(
        n15173) );
  NOR2_X1 U16690 ( .A1(n15174), .A2(n15173), .ZN(n15192) );
  INV_X1 U16691 ( .A(P3_REG0_REG_9__SCAN_IN), .ZN(n15176) );
  AOI22_X1 U16692 ( .A1(n15177), .A2(n15192), .B1(n15176), .B2(n15175), .ZN(
        P3_U3417) );
  AOI22_X1 U16693 ( .A1(n15193), .A2(n15178), .B1(n9771), .B2(n15190), .ZN(
        P3_U3460) );
  AOI22_X1 U16694 ( .A1(n15193), .A2(n15179), .B1(n10075), .B2(n15190), .ZN(
        P3_U3461) );
  AOI22_X1 U16695 ( .A1(n15193), .A2(n15180), .B1(n10061), .B2(n15190), .ZN(
        P3_U3462) );
  AOI22_X1 U16696 ( .A1(n15193), .A2(n15182), .B1(n15181), .B2(n15190), .ZN(
        P3_U3463) );
  AOI22_X1 U16697 ( .A1(n15193), .A2(n15183), .B1(n10071), .B2(n15190), .ZN(
        P3_U3464) );
  AOI22_X1 U16698 ( .A1(n15193), .A2(n15185), .B1(n15184), .B2(n15190), .ZN(
        P3_U3465) );
  INV_X1 U16699 ( .A(P3_REG1_REG_7__SCAN_IN), .ZN(n15186) );
  AOI22_X1 U16700 ( .A1(n15193), .A2(n15187), .B1(n15186), .B2(n15190), .ZN(
        P3_U3466) );
  AOI22_X1 U16701 ( .A1(n15193), .A2(n15189), .B1(n15188), .B2(n15190), .ZN(
        P3_U3467) );
  INV_X1 U16702 ( .A(P3_REG1_REG_9__SCAN_IN), .ZN(n15191) );
  AOI22_X1 U16703 ( .A1(n15193), .A2(n15192), .B1(n15191), .B2(n15190), .ZN(
        P3_U3468) );
  XOR2_X1 U16704 ( .A(n15195), .B(n15194), .Z(SUB_1596_U59) );
  XOR2_X1 U16705 ( .A(n15197), .B(n15196), .Z(SUB_1596_U58) );
  AOI21_X1 U16706 ( .B1(n15199), .B2(n15198), .A(n15208), .ZN(SUB_1596_U53) );
  XNOR2_X1 U16707 ( .A(n15201), .B(n15200), .ZN(SUB_1596_U56) );
  OAI21_X1 U16708 ( .B1(n15204), .B2(n15203), .A(n15202), .ZN(n15206) );
  XOR2_X1 U16709 ( .A(n15206), .B(n15205), .Z(SUB_1596_U60) );
  XOR2_X1 U16710 ( .A(n15208), .B(n15207), .Z(SUB_1596_U5) );
  CLKBUF_X1 U7232 ( .A(n7462), .Z(n6481) );
  CLKBUF_X1 U7325 ( .A(n8835), .Z(n10012) );
  CLKBUF_X1 U8294 ( .A(n8821), .Z(n8822) );
  CLKBUF_X1 U9110 ( .A(n7462), .Z(n6480) );
  NAND2_X1 U9545 ( .A1(n9334), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9335) );
endmodule

