

module b22_C_2inp_gates_syn ( P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN, 
        P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN, 
        P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN, 
        P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN, 
        P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN, 
        P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN, 
        P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN, 
        P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN, 
        P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN, 
        P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN, P3_REG3_REG_0__SCAN_IN, 
        P3_REG3_REG_20__SCAN_IN, P3_REG3_REG_13__SCAN_IN, 
        P3_REG3_REG_22__SCAN_IN, P3_REG3_REG_11__SCAN_IN, 
        P3_REG3_REG_2__SCAN_IN, P3_REG3_REG_18__SCAN_IN, 
        P3_REG3_REG_6__SCAN_IN, P3_REG3_REG_26__SCAN_IN, 
        P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_ADDR_REG_0__SCAN_IN, 
        P3_ADDR_REG_1__SCAN_IN, P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN, 
        P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN, P3_ADDR_REG_6__SCAN_IN, 
        P3_ADDR_REG_7__SCAN_IN, P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, 
        P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, 
        P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, 
        P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, 
        P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, 
        P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, 
        P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, 
        P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, 
        P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, 
        P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, 
        P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, 
        P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, 
        P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, 
        P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, 
        P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, 
        P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, 
        P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, 
        P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, 
        P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, 
        P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, 
        P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, 
        P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, 
        P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, 
        P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, 
        P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, 
        P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, 
        P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN, 
        P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN, 
        P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN, 
        P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN, 
        P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN, 
        P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN, 
        P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN, 
        P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN, 
        P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN, 
        P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN, 
        P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN, 
        P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN, 
        P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN, 
        P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN, 
        P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN, 
        P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN, 
        P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN, 
        P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_4__SCAN_IN, 
        P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_17__SCAN_IN, 
        P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_16__SCAN_IN, 
        P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_12__SCAN_IN, 
        P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_1__SCAN_IN, 
        P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_28__SCAN_IN, 
        P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_3__SCAN_IN, 
        P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_23__SCAN_IN, 
        P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_27__SCAN_IN, 
        P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN, P2_RD_REG_SCAN_IN, 
        P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN, P3_IR_REG_1__SCAN_IN, 
        P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN, P3_IR_REG_4__SCAN_IN, 
        P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN, P3_IR_REG_7__SCAN_IN, 
        P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN, P3_IR_REG_10__SCAN_IN, 
        P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN, P3_IR_REG_13__SCAN_IN, 
        P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN, P3_IR_REG_16__SCAN_IN, 
        P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN, P3_IR_REG_19__SCAN_IN, 
        P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN, P3_IR_REG_22__SCAN_IN, 
        P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN, P3_IR_REG_25__SCAN_IN, 
        P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN, P3_IR_REG_28__SCAN_IN, 
        P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN, P3_IR_REG_31__SCAN_IN, 
        P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN, P3_D_REG_2__SCAN_IN, 
        P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN, P3_D_REG_5__SCAN_IN, 
        P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN, P3_D_REG_8__SCAN_IN, 
        P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN, P3_D_REG_11__SCAN_IN, 
        P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN, P3_D_REG_14__SCAN_IN, 
        P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN, P3_D_REG_17__SCAN_IN, 
        P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN, P3_D_REG_20__SCAN_IN, 
        P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN, P3_D_REG_23__SCAN_IN, 
        P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN, P3_D_REG_26__SCAN_IN, 
        P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN, P3_D_REG_29__SCAN_IN, 
        P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN, P3_REG0_REG_0__SCAN_IN, 
        P3_REG0_REG_1__SCAN_IN, P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN, 
        P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN, P3_REG0_REG_6__SCAN_IN, 
        P3_REG0_REG_7__SCAN_IN, P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN, 
        P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN, 
        P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN, 
        P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN, 
        P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN, 
        P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN, 
        P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN, 
        P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN, 
        P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN, 
        P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN, 
        P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN, 
        P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN, 
        P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN, P3_REG1_REG_2__SCAN_IN, 
        P3_REG1_REG_3__SCAN_IN, P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN, 
        P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN, P3_REG1_REG_8__SCAN_IN, 
        P3_REG1_REG_9__SCAN_IN, P3_REG1_REG_10__SCAN_IN, 
        P3_REG1_REG_11__SCAN_IN, P3_REG1_REG_12__SCAN_IN, 
        P3_REG1_REG_13__SCAN_IN, P3_REG1_REG_14__SCAN_IN, 
        P3_REG1_REG_15__SCAN_IN, P3_REG1_REG_16__SCAN_IN, 
        P3_REG1_REG_17__SCAN_IN, P3_REG1_REG_18__SCAN_IN, 
        P3_REG1_REG_19__SCAN_IN, P3_REG1_REG_20__SCAN_IN, 
        P3_REG1_REG_21__SCAN_IN, P3_REG1_REG_22__SCAN_IN, 
        P3_REG1_REG_23__SCAN_IN, P3_REG1_REG_24__SCAN_IN, 
        P3_REG1_REG_25__SCAN_IN, P3_REG1_REG_26__SCAN_IN, 
        P3_REG1_REG_27__SCAN_IN, P3_REG1_REG_28__SCAN_IN, 
        P3_REG1_REG_29__SCAN_IN, P3_REG1_REG_30__SCAN_IN, 
        P3_REG1_REG_31__SCAN_IN, P3_REG2_REG_0__SCAN_IN, 
        P3_REG2_REG_1__SCAN_IN, P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN, 
        P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN, P3_REG2_REG_6__SCAN_IN, 
        P3_REG2_REG_7__SCAN_IN, P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN, 
        P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN, 
        P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN, 
        P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN, 
        P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN, 
        P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN, 
        P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN, 
        P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN, 
        P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN, 
        P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN, 
        P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN, 
        P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN, 
        P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN, 
        P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN, 
        P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN, 
        P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN, 
        P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, SUB_1596_U4, 
        SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65, SUB_1596_U66, 
        SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70, SUB_1596_U54, 
        SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58, SUB_1596_U59, 
        SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53, U29, U28, 
        P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349, 
        P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342, 
        P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335, 
        P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328, 
        P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446, P1_U3323, 
        P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316, 
        P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309, 
        P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302, 
        P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295, 
        P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471, P1_U3474, 
        P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492, P1_U3495, 
        P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513, P1_U3515, 
        P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, 
        P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, 
        P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, 
        P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, 
        P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, 
        P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556, P1_U3557, 
        P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290, P1_U3289, 
        P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282, 
        P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275, 
        P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268, 
        P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, P1_U3262, 
        P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255, 
        P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248, 
        P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560, P1_U3561, 
        P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, 
        P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, 
        P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, 
        P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588, P1_U3589, 
        P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239, P1_U3238, 
        P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231, 
        P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224, 
        P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, 
        P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, P1_U4016, 
        P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321, 
        P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314, 
        P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307, 
        P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300, 
        P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417, P2_U3295, 
        P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, 
        P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, 
        P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, 
        P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, 
        P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442, P2_U3445, 
        P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463, P2_U3466, 
        P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484, P2_U3486, 
        P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492, P2_U3493, 
        P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499, P2_U3500, 
        P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506, P2_U3507, 
        P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, P2_U3514, 
        P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, P2_U3521, 
        P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527, P2_U3528, 
        P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, 
        P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, 
        P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, 
        P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241, P2_U3240, 
        P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, 
        P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, 
        P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, 
        P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531, P2_U3532, 
        P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, 
        P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, 
        P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552, P2_U3553, 
        P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559, P2_U3560, 
        P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211, P2_U3210, 
        P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, 
        P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, 
        P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, 
        P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087, P2_U3947, 
        P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290, P3_U3289, 
        P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283, P3_U3282, 
        P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276, P3_U3275, 
        P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269, P3_U3268, 
        P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377, P3_U3263, 
        P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257, P3_U3256, 
        P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250, P3_U3249, 
        P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243, P3_U3242, 
        P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236, P3_U3235, 
        P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402, P3_U3405, 
        P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423, P3_U3426, 
        P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444, P3_U3446, 
        P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452, P3_U3453, 
        P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459, P3_U3460, 
        P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466, P3_U3467, 
        P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473, P3_U3474, 
        P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480, P3_U3481, 
        P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487, P3_U3488, 
        P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230, P3_U3229, 
        P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223, P3_U3222, 
        P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216, P3_U3215, 
        P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209, P3_U3208, 
        P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202, P3_U3201, 
        P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195, P3_U3194, 
        P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188, P3_U3187, 
        P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491, P3_U3492, 
        P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498, P3_U3499, 
        P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505, P3_U3506, 
        P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512, P3_U3513, 
        P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519, P3_U3520, 
        P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179, P3_U3178, 
        P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172, P3_U3171, 
        P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165, P3_U3164, 
        P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158, P3_U3157, 
        P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150, P3_U3897, 
        keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, 
        keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, 
        keyinput12, keyinput13, keyinput14, keyinput15, keyinput16, keyinput17, 
        keyinput18, keyinput19, keyinput20, keyinput21, keyinput22, keyinput23, 
        keyinput24, keyinput25, keyinput26, keyinput27, keyinput28, keyinput29, 
        keyinput30, keyinput31, keyinput32, keyinput33, keyinput34, keyinput35, 
        keyinput36, keyinput37, keyinput38, keyinput39, keyinput40, keyinput41, 
        keyinput42, keyinput43, keyinput44, keyinput45, keyinput46, keyinput47, 
        keyinput48, keyinput49, keyinput50, keyinput51, keyinput52, keyinput53, 
        keyinput54, keyinput55, keyinput56, keyinput57, keyinput58, keyinput59, 
        keyinput60, keyinput61, keyinput62, keyinput63, keyinput64, keyinput65, 
        keyinput66, keyinput67, keyinput68, keyinput69, keyinput70, keyinput71, 
        keyinput72, keyinput73, keyinput74, keyinput75, keyinput76, keyinput77, 
        keyinput78, keyinput79, keyinput80, keyinput81, keyinput82, keyinput83, 
        keyinput84, keyinput85, keyinput86, keyinput87, keyinput88, keyinput89, 
        keyinput90, keyinput91, keyinput92, keyinput93, keyinput94, keyinput95, 
        keyinput96, keyinput97, keyinput98, keyinput99, keyinput100, 
        keyinput101, keyinput102, keyinput103, keyinput104, keyinput105, 
        keyinput106, keyinput107, keyinput108, keyinput109, keyinput110, 
        keyinput111, keyinput112, keyinput113, keyinput114, keyinput115, 
        keyinput116, keyinput117, keyinput118, keyinput119, keyinput120, 
        keyinput121, keyinput122, keyinput123, keyinput124, keyinput125, 
        keyinput126, keyinput127 );
  input P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN,
         P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN,
         P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN,
         P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN,
         P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN,
         P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN,
         P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN,
         P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN,
         P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN,
         P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN,
         P3_REG3_REG_0__SCAN_IN, P3_REG3_REG_20__SCAN_IN,
         P3_REG3_REG_13__SCAN_IN, P3_REG3_REG_22__SCAN_IN,
         P3_REG3_REG_11__SCAN_IN, P3_REG3_REG_2__SCAN_IN,
         P3_REG3_REG_18__SCAN_IN, P3_REG3_REG_6__SCAN_IN,
         P3_REG3_REG_26__SCAN_IN, P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN,
         P3_DATAO_REG_31__SCAN_IN, P3_DATAO_REG_30__SCAN_IN,
         P3_DATAO_REG_29__SCAN_IN, P3_DATAO_REG_28__SCAN_IN,
         P3_DATAO_REG_27__SCAN_IN, P3_DATAO_REG_26__SCAN_IN,
         P3_DATAO_REG_25__SCAN_IN, P3_DATAO_REG_24__SCAN_IN,
         P3_DATAO_REG_23__SCAN_IN, P3_DATAO_REG_22__SCAN_IN,
         P3_DATAO_REG_21__SCAN_IN, P3_DATAO_REG_20__SCAN_IN,
         P3_DATAO_REG_19__SCAN_IN, P3_DATAO_REG_18__SCAN_IN,
         P3_DATAO_REG_17__SCAN_IN, P3_DATAO_REG_16__SCAN_IN,
         P3_DATAO_REG_15__SCAN_IN, P3_DATAO_REG_14__SCAN_IN,
         P3_DATAO_REG_13__SCAN_IN, P3_DATAO_REG_12__SCAN_IN,
         P3_DATAO_REG_11__SCAN_IN, P3_DATAO_REG_10__SCAN_IN,
         P3_DATAO_REG_9__SCAN_IN, P3_DATAO_REG_8__SCAN_IN,
         P3_DATAO_REG_7__SCAN_IN, P3_DATAO_REG_6__SCAN_IN,
         P3_DATAO_REG_5__SCAN_IN, P3_DATAO_REG_4__SCAN_IN,
         P3_DATAO_REG_3__SCAN_IN, P3_DATAO_REG_2__SCAN_IN,
         P3_DATAO_REG_1__SCAN_IN, P3_DATAO_REG_0__SCAN_IN,
         P3_ADDR_REG_0__SCAN_IN, P3_ADDR_REG_1__SCAN_IN,
         P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN,
         P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN,
         P3_ADDR_REG_6__SCAN_IN, P3_ADDR_REG_7__SCAN_IN,
         P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, P1_IR_REG_0__SCAN_IN,
         P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN,
         P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN,
         P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN,
         P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN,
         P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN,
         P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN,
         P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN,
         P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN,
         P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN,
         P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN,
         P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN,
         P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN,
         P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN,
         P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN,
         P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN,
         P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN,
         P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN,
         P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN,
         P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN,
         P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN,
         P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN,
         P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN,
         P2_RD_REG_SCAN_IN, P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN,
         P3_IR_REG_1__SCAN_IN, P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN,
         P3_IR_REG_4__SCAN_IN, P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN,
         P3_IR_REG_7__SCAN_IN, P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN,
         P3_IR_REG_10__SCAN_IN, P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN,
         P3_IR_REG_13__SCAN_IN, P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN,
         P3_IR_REG_16__SCAN_IN, P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN,
         P3_IR_REG_19__SCAN_IN, P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN,
         P3_IR_REG_22__SCAN_IN, P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN,
         P3_IR_REG_25__SCAN_IN, P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN,
         P3_IR_REG_28__SCAN_IN, P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN,
         P3_IR_REG_31__SCAN_IN, P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN,
         P3_D_REG_2__SCAN_IN, P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN,
         P3_D_REG_5__SCAN_IN, P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN,
         P3_D_REG_8__SCAN_IN, P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN,
         P3_D_REG_11__SCAN_IN, P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN,
         P3_D_REG_14__SCAN_IN, P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN,
         P3_D_REG_17__SCAN_IN, P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN,
         P3_D_REG_20__SCAN_IN, P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN,
         P3_D_REG_23__SCAN_IN, P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN,
         P3_D_REG_26__SCAN_IN, P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN,
         P3_D_REG_29__SCAN_IN, P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN,
         P3_REG0_REG_0__SCAN_IN, P3_REG0_REG_1__SCAN_IN,
         P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN,
         P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN,
         P3_REG0_REG_6__SCAN_IN, P3_REG0_REG_7__SCAN_IN,
         P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN,
         P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN,
         P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN,
         P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN,
         P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN,
         P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN,
         P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN,
         P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN,
         P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN,
         P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN,
         P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN,
         P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN,
         P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN,
         P3_REG1_REG_2__SCAN_IN, P3_REG1_REG_3__SCAN_IN,
         P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN,
         P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN,
         P3_REG1_REG_8__SCAN_IN, P3_REG1_REG_9__SCAN_IN,
         P3_REG1_REG_10__SCAN_IN, P3_REG1_REG_11__SCAN_IN,
         P3_REG1_REG_12__SCAN_IN, P3_REG1_REG_13__SCAN_IN,
         P3_REG1_REG_14__SCAN_IN, P3_REG1_REG_15__SCAN_IN,
         P3_REG1_REG_16__SCAN_IN, P3_REG1_REG_17__SCAN_IN,
         P3_REG1_REG_18__SCAN_IN, P3_REG1_REG_19__SCAN_IN,
         P3_REG1_REG_20__SCAN_IN, P3_REG1_REG_21__SCAN_IN,
         P3_REG1_REG_22__SCAN_IN, P3_REG1_REG_23__SCAN_IN,
         P3_REG1_REG_24__SCAN_IN, P3_REG1_REG_25__SCAN_IN,
         P3_REG1_REG_26__SCAN_IN, P3_REG1_REG_27__SCAN_IN,
         P3_REG1_REG_28__SCAN_IN, P3_REG1_REG_29__SCAN_IN,
         P3_REG1_REG_30__SCAN_IN, P3_REG1_REG_31__SCAN_IN,
         P3_REG2_REG_0__SCAN_IN, P3_REG2_REG_1__SCAN_IN,
         P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN,
         P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN,
         P3_REG2_REG_6__SCAN_IN, P3_REG2_REG_7__SCAN_IN,
         P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN,
         P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN,
         P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN,
         P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN,
         P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN,
         P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN,
         P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN,
         P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN,
         P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN,
         P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN,
         P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN,
         P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN,
         P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN,
         P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN,
         P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN,
         P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN,
         P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, keyinput0,
         keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, keyinput6,
         keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, keyinput12,
         keyinput13, keyinput14, keyinput15, keyinput16, keyinput17,
         keyinput18, keyinput19, keyinput20, keyinput21, keyinput22,
         keyinput23, keyinput24, keyinput25, keyinput26, keyinput27,
         keyinput28, keyinput29, keyinput30, keyinput31, keyinput32,
         keyinput33, keyinput34, keyinput35, keyinput36, keyinput37,
         keyinput38, keyinput39, keyinput40, keyinput41, keyinput42,
         keyinput43, keyinput44, keyinput45, keyinput46, keyinput47,
         keyinput48, keyinput49, keyinput50, keyinput51, keyinput52,
         keyinput53, keyinput54, keyinput55, keyinput56, keyinput57,
         keyinput58, keyinput59, keyinput60, keyinput61, keyinput62,
         keyinput63, keyinput64, keyinput65, keyinput66, keyinput67,
         keyinput68, keyinput69, keyinput70, keyinput71, keyinput72,
         keyinput73, keyinput74, keyinput75, keyinput76, keyinput77,
         keyinput78, keyinput79, keyinput80, keyinput81, keyinput82,
         keyinput83, keyinput84, keyinput85, keyinput86, keyinput87,
         keyinput88, keyinput89, keyinput90, keyinput91, keyinput92,
         keyinput93, keyinput94, keyinput95, keyinput96, keyinput97,
         keyinput98, keyinput99, keyinput100, keyinput101, keyinput102,
         keyinput103, keyinput104, keyinput105, keyinput106, keyinput107,
         keyinput108, keyinput109, keyinput110, keyinput111, keyinput112,
         keyinput113, keyinput114, keyinput115, keyinput116, keyinput117,
         keyinput118, keyinput119, keyinput120, keyinput121, keyinput122,
         keyinput123, keyinput124, keyinput125, keyinput126, keyinput127;
  output SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65,
         SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70,
         SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58,
         SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53,
         U29, U28, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350,
         P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343,
         P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336,
         P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329,
         P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446,
         P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317,
         P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310,
         P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303,
         P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296,
         P1_U3295, P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471,
         P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492,
         P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556,
         P1_U3557, P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290,
         P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283,
         P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276,
         P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269,
         P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263,
         P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256,
         P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249,
         P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588,
         P1_U3589, P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239,
         P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232,
         P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085,
         P1_U4016, P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322,
         P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315,
         P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308,
         P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301,
         P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417,
         P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289,
         P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282,
         P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275,
         P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268,
         P2_U3267, P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442,
         P2_U3445, P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463,
         P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484,
         P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492,
         P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499,
         P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506,
         P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513,
         P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520,
         P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527,
         P2_U3528, P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262,
         P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255,
         P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248,
         P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241,
         P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234,
         P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227,
         P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220,
         P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531,
         P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538,
         P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545,
         P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552,
         P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559,
         P2_U3560, P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204,
         P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197,
         P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190,
         P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087,
         P2_U3947, P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290,
         P3_U3289, P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283,
         P3_U3282, P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276,
         P3_U3275, P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269,
         P3_U3268, P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377,
         P3_U3263, P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257,
         P3_U3256, P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250,
         P3_U3249, P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243,
         P3_U3242, P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236,
         P3_U3235, P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402,
         P3_U3405, P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423,
         P3_U3426, P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444,
         P3_U3446, P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452,
         P3_U3453, P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459,
         P3_U3460, P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466,
         P3_U3467, P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473,
         P3_U3474, P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480,
         P3_U3481, P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487,
         P3_U3488, P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230,
         P3_U3229, P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223,
         P3_U3222, P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216,
         P3_U3215, P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209,
         P3_U3208, P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202,
         P3_U3201, P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195,
         P3_U3194, P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188,
         P3_U3187, P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491,
         P3_U3492, P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498,
         P3_U3499, P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505,
         P3_U3506, P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512,
         P3_U3513, P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519,
         P3_U3520, P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179,
         P3_U3178, P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172,
         P3_U3171, P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165,
         P3_U3164, P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158,
         P3_U3157, P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150,
         P3_U3897;
  wire   n6547, n6548, n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557,
         n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567,
         n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577,
         n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587,
         n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597,
         n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607,
         n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617,
         n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627,
         n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637,
         n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647,
         n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657,
         n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667,
         n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677,
         n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687,
         n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697,
         n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707,
         n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6716, n6717, n6718,
         n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728,
         n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738,
         n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748,
         n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758,
         n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768,
         n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778,
         n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788,
         n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798,
         n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808,
         n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818,
         n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828,
         n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838,
         n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848,
         n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858,
         n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868,
         n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878,
         n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888,
         n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898,
         n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908,
         n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918,
         n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928,
         n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938,
         n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948,
         n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958,
         n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968,
         n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978,
         n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988,
         n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998,
         n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008,
         n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018,
         n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028,
         n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038,
         n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048,
         n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058,
         n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068,
         n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078,
         n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088,
         n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098,
         n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108,
         n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118,
         n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128,
         n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138,
         n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148,
         n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158,
         n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168,
         n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178,
         n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188,
         n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198,
         n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208,
         n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218,
         n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228,
         n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238,
         n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248,
         n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258,
         n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268,
         n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7279,
         n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289,
         n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299,
         n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309,
         n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319,
         n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329,
         n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339,
         n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349,
         n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359,
         n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369,
         n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379,
         n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389,
         n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399,
         n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409,
         n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419,
         n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429,
         n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439,
         n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449,
         n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459,
         n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469,
         n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479,
         n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489,
         n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499,
         n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509,
         n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519,
         n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529,
         n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539,
         n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549,
         n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559,
         n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569,
         n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579,
         n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589,
         n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599,
         n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609,
         n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619,
         n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629,
         n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639,
         n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649,
         n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659,
         n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669,
         n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679,
         n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689,
         n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699,
         n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709,
         n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719,
         n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729,
         n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739,
         n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749,
         n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759,
         n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769,
         n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779,
         n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789,
         n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799,
         n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809,
         n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819,
         n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829,
         n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839,
         n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849,
         n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859,
         n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869,
         n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879,
         n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889,
         n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899,
         n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909,
         n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919,
         n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929,
         n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939,
         n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949,
         n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959,
         n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969,
         n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979,
         n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989,
         n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999,
         n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009,
         n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019,
         n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029,
         n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039,
         n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049,
         n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059,
         n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069,
         n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079,
         n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089,
         n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099,
         n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109,
         n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119,
         n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129,
         n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139,
         n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149,
         n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159,
         n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169,
         n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179,
         n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189,
         n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199,
         n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209,
         n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219,
         n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229,
         n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239,
         n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249,
         n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259,
         n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269,
         n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279,
         n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289,
         n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299,
         n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309,
         n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319,
         n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329,
         n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339,
         n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349,
         n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359,
         n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369,
         n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379,
         n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389,
         n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399,
         n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409,
         n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419,
         n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429,
         n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439,
         n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449,
         n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459,
         n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469,
         n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479,
         n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489,
         n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499,
         n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509,
         n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519,
         n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529,
         n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539,
         n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549,
         n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559,
         n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569,
         n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579,
         n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589,
         n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599,
         n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609,
         n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619,
         n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629,
         n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639,
         n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649,
         n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659,
         n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669,
         n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679,
         n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689,
         n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699,
         n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709,
         n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719,
         n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729,
         n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739,
         n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749,
         n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759,
         n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769,
         n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779,
         n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789,
         n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799,
         n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809,
         n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819,
         n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829,
         n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839,
         n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849,
         n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859,
         n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869,
         n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879,
         n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889,
         n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899,
         n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909,
         n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919,
         n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929,
         n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939,
         n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949,
         n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959,
         n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969,
         n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979,
         n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989,
         n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999,
         n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009,
         n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019,
         n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029,
         n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039,
         n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049,
         n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059,
         n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069,
         n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079,
         n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089,
         n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099,
         n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109,
         n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119,
         n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129,
         n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139,
         n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149,
         n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159,
         n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169,
         n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179,
         n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189,
         n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199,
         n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209,
         n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219,
         n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229,
         n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239,
         n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249,
         n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259,
         n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269,
         n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279,
         n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289,
         n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299,
         n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309,
         n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319,
         n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329,
         n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339,
         n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349,
         n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359,
         n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369,
         n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379,
         n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389,
         n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399,
         n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409,
         n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419,
         n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429,
         n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439,
         n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449,
         n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459,
         n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469,
         n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479,
         n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489,
         n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499,
         n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509,
         n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519,
         n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529,
         n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539,
         n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549,
         n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559,
         n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569,
         n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579,
         n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589,
         n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9599, n9600,
         n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610,
         n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620,
         n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630,
         n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640,
         n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650,
         n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660,
         n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670,
         n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680,
         n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690,
         n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700,
         n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710,
         n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720,
         n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730,
         n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740,
         n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750,
         n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760,
         n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770,
         n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780,
         n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790,
         n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800,
         n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810,
         n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820,
         n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830,
         n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840,
         n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850,
         n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860,
         n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870,
         n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880,
         n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890,
         n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900,
         n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910,
         n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920,
         n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930,
         n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940,
         n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950,
         n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960,
         n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970,
         n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980,
         n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990,
         n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000,
         n10001, n10002, n10003, n10004, n10005, n10006, n10007, n10008,
         n10009, n10010, n10011, n10012, n10013, n10014, n10015, n10016,
         n10017, n10018, n10019, n10020, n10021, n10022, n10023, n10024,
         n10025, n10026, n10027, n10028, n10029, n10030, n10031, n10032,
         n10033, n10034, n10035, n10036, n10037, n10038, n10039, n10040,
         n10041, n10042, n10043, n10044, n10045, n10046, n10047, n10048,
         n10049, n10050, n10051, n10052, n10053, n10054, n10055, n10056,
         n10057, n10058, n10059, n10060, n10061, n10062, n10063, n10064,
         n10065, n10066, n10067, n10068, n10069, n10070, n10071, n10072,
         n10073, n10074, n10075, n10076, n10077, n10078, n10079, n10080,
         n10081, n10082, n10083, n10084, n10085, n10086, n10087, n10088,
         n10089, n10090, n10091, n10092, n10093, n10094, n10095, n10096,
         n10097, n10098, n10099, n10100, n10101, n10102, n10103, n10104,
         n10105, n10106, n10107, n10108, n10109, n10110, n10111, n10112,
         n10113, n10114, n10115, n10116, n10117, n10118, n10119, n10120,
         n10121, n10122, n10123, n10124, n10125, n10126, n10127, n10128,
         n10129, n10130, n10131, n10132, n10133, n10134, n10135, n10136,
         n10137, n10138, n10139, n10140, n10141, n10142, n10143, n10144,
         n10145, n10146, n10147, n10148, n10149, n10150, n10151, n10152,
         n10153, n10154, n10155, n10156, n10157, n10158, n10159, n10160,
         n10161, n10162, n10163, n10164, n10165, n10166, n10167, n10168,
         n10169, n10170, n10171, n10172, n10173, n10174, n10175, n10176,
         n10177, n10178, n10179, n10180, n10181, n10182, n10183, n10184,
         n10185, n10186, n10187, n10188, n10189, n10190, n10191, n10192,
         n10193, n10194, n10195, n10196, n10197, n10198, n10199, n10200,
         n10201, n10202, n10203, n10204, n10205, n10206, n10207, n10208,
         n10209, n10210, n10211, n10212, n10213, n10214, n10215, n10216,
         n10217, n10218, n10219, n10220, n10221, n10222, n10223, n10224,
         n10225, n10226, n10227, n10228, n10229, n10230, n10231, n10232,
         n10233, n10234, n10235, n10236, n10237, n10238, n10239, n10240,
         n10241, n10242, n10243, n10244, n10245, n10246, n10247, n10248,
         n10249, n10250, n10251, n10252, n10253, n10254, n10255, n10256,
         n10257, n10258, n10259, n10260, n10261, n10262, n10263, n10264,
         n10265, n10266, n10267, n10268, n10269, n10270, n10271, n10272,
         n10273, n10274, n10275, n10276, n10277, n10278, n10279, n10280,
         n10281, n10282, n10283, n10284, n10285, n10286, n10287, n10288,
         n10289, n10290, n10291, n10292, n10293, n10294, n10295, n10296,
         n10297, n10298, n10299, n10300, n10301, n10302, n10303, n10304,
         n10305, n10306, n10307, n10308, n10309, n10310, n10311, n10312,
         n10313, n10314, n10315, n10316, n10317, n10318, n10319, n10320,
         n10321, n10322, n10323, n10324, n10325, n10326, n10327, n10328,
         n10329, n10330, n10331, n10332, n10333, n10334, n10335, n10336,
         n10337, n10338, n10339, n10340, n10341, n10342, n10343, n10344,
         n10345, n10346, n10347, n10348, n10349, n10350, n10351, n10352,
         n10353, n10354, n10355, n10356, n10357, n10358, n10359, n10360,
         n10361, n10362, n10363, n10364, n10365, n10366, n10367, n10368,
         n10369, n10370, n10371, n10372, n10373, n10374, n10375, n10376,
         n10377, n10378, n10379, n10380, n10381, n10382, n10383, n10384,
         n10385, n10386, n10387, n10388, n10389, n10390, n10391, n10392,
         n10393, n10394, n10395, n10396, n10397, n10398, n10399, n10400,
         n10401, n10402, n10403, n10404, n10405, n10406, n10407, n10408,
         n10409, n10410, n10411, n10412, n10413, n10414, n10415, n10416,
         n10417, n10418, n10419, n10420, n10421, n10422, n10423, n10424,
         n10425, n10426, n10427, n10428, n10429, n10430, n10431, n10432,
         n10433, n10434, n10435, n10436, n10437, n10438, n10439, n10440,
         n10441, n10442, n10443, n10444, n10445, n10446, n10447, n10448,
         n10449, n10450, n10451, n10452, n10453, n10454, n10455, n10456,
         n10457, n10458, n10459, n10460, n10461, n10462, n10463, n10464,
         n10465, n10466, n10467, n10468, n10469, n10470, n10471, n10472,
         n10473, n10474, n10475, n10476, n10477, n10478, n10479, n10480,
         n10481, n10482, n10483, n10484, n10485, n10486, n10487, n10488,
         n10489, n10490, n10491, n10492, n10493, n10494, n10495, n10496,
         n10497, n10498, n10499, n10500, n10501, n10502, n10503, n10504,
         n10505, n10506, n10507, n10508, n10509, n10510, n10511, n10512,
         n10513, n10514, n10515, n10516, n10517, n10518, n10519, n10520,
         n10521, n10522, n10523, n10524, n10525, n10526, n10527, n10528,
         n10529, n10530, n10531, n10532, n10533, n10534, n10535, n10536,
         n10537, n10538, n10539, n10540, n10541, n10542, n10543, n10544,
         n10545, n10546, n10547, n10548, n10549, n10550, n10551, n10552,
         n10553, n10554, n10555, n10556, n10557, n10558, n10559, n10560,
         n10561, n10562, n10563, n10564, n10565, n10566, n10567, n10568,
         n10569, n10570, n10571, n10572, n10573, n10574, n10575, n10576,
         n10577, n10578, n10579, n10580, n10581, n10582, n10583, n10584,
         n10585, n10586, n10587, n10588, n10589, n10590, n10591, n10592,
         n10593, n10594, n10595, n10596, n10597, n10598, n10599, n10600,
         n10601, n10602, n10603, n10604, n10605, n10606, n10607, n10608,
         n10609, n10610, n10611, n10612, n10613, n10614, n10615, n10616,
         n10617, n10618, n10619, n10620, n10621, n10622, n10623, n10624,
         n10625, n10626, n10627, n10628, n10629, n10630, n10631, n10632,
         n10633, n10634, n10635, n10636, n10637, n10638, n10639, n10640,
         n10641, n10642, n10643, n10644, n10645, n10646, n10647, n10648,
         n10649, n10650, n10651, n10652, n10653, n10654, n10655, n10656,
         n10657, n10658, n10659, n10660, n10661, n10662, n10663, n10664,
         n10665, n10666, n10667, n10668, n10669, n10670, n10671, n10672,
         n10673, n10674, n10675, n10676, n10677, n10678, n10679, n10680,
         n10681, n10682, n10683, n10684, n10685, n10686, n10687, n10688,
         n10689, n10690, n10691, n10692, n10693, n10694, n10695, n10696,
         n10697, n10698, n10699, n10700, n10701, n10702, n10703, n10704,
         n10705, n10706, n10707, n10708, n10709, n10710, n10711, n10712,
         n10713, n10714, n10715, n10716, n10717, n10718, n10719, n10720,
         n10721, n10722, n10723, n10724, n10725, n10726, n10727, n10728,
         n10729, n10730, n10731, n10732, n10733, n10734, n10735, n10736,
         n10737, n10738, n10739, n10740, n10741, n10742, n10743, n10744,
         n10745, n10746, n10747, n10748, n10749, n10750, n10751, n10752,
         n10753, n10754, n10755, n10756, n10757, n10758, n10759, n10760,
         n10761, n10762, n10763, n10764, n10765, n10766, n10767, n10768,
         n10769, n10770, n10771, n10772, n10773, n10774, n10775, n10776,
         n10777, n10778, n10779, n10780, n10781, n10782, n10783, n10784,
         n10785, n10786, n10787, n10788, n10789, n10790, n10791, n10792,
         n10793, n10794, n10795, n10796, n10797, n10798, n10799, n10800,
         n10801, n10802, n10803, n10804, n10805, n10806, n10807, n10808,
         n10809, n10810, n10811, n10812, n10813, n10814, n10815, n10816,
         n10817, n10818, n10819, n10820, n10821, n10822, n10823, n10824,
         n10825, n10826, n10827, n10828, n10829, n10830, n10831, n10832,
         n10833, n10834, n10835, n10836, n10837, n10838, n10839, n10840,
         n10841, n10842, n10843, n10844, n10845, n10846, n10847, n10848,
         n10849, n10850, n10851, n10852, n10853, n10854, n10855, n10856,
         n10857, n10858, n10859, n10860, n10861, n10862, n10863, n10864,
         n10865, n10866, n10867, n10868, n10869, n10870, n10871, n10872,
         n10873, n10874, n10875, n10876, n10877, n10878, n10879, n10880,
         n10881, n10882, n10883, n10884, n10885, n10886, n10887, n10888,
         n10889, n10890, n10891, n10892, n10893, n10894, n10895, n10896,
         n10897, n10898, n10899, n10900, n10901, n10902, n10903, n10904,
         n10905, n10906, n10907, n10908, n10909, n10910, n10911, n10912,
         n10913, n10914, n10915, n10916, n10917, n10918, n10919, n10920,
         n10921, n10922, n10923, n10924, n10925, n10926, n10927, n10928,
         n10929, n10930, n10931, n10932, n10933, n10934, n10935, n10936,
         n10937, n10938, n10939, n10940, n10941, n10942, n10943, n10944,
         n10945, n10946, n10947, n10948, n10949, n10950, n10951, n10952,
         n10953, n10954, n10955, n10956, n10957, n10958, n10959, n10960,
         n10961, n10962, n10963, n10964, n10965, n10966, n10967, n10968,
         n10969, n10970, n10971, n10972, n10973, n10974, n10975, n10976,
         n10977, n10978, n10979, n10980, n10981, n10982, n10983, n10984,
         n10985, n10986, n10987, n10988, n10989, n10990, n10991, n10992,
         n10993, n10994, n10995, n10996, n10997, n10998, n10999, n11000,
         n11001, n11002, n11003, n11004, n11005, n11006, n11007, n11008,
         n11009, n11010, n11011, n11012, n11013, n11014, n11015, n11016,
         n11017, n11018, n11019, n11020, n11021, n11022, n11023, n11024,
         n11025, n11026, n11027, n11028, n11029, n11030, n11031, n11032,
         n11033, n11034, n11035, n11036, n11037, n11038, n11039, n11040,
         n11041, n11042, n11043, n11044, n11045, n11046, n11047, n11048,
         n11049, n11050, n11051, n11052, n11053, n11054, n11055, n11056,
         n11057, n11058, n11059, n11060, n11061, n11062, n11063, n11064,
         n11065, n11066, n11067, n11068, n11069, n11070, n11071, n11072,
         n11073, n11074, n11075, n11076, n11077, n11078, n11079, n11080,
         n11081, n11082, n11083, n11084, n11085, n11086, n11087, n11088,
         n11089, n11090, n11091, n11092, n11093, n11094, n11095, n11096,
         n11097, n11098, n11099, n11100, n11101, n11102, n11103, n11104,
         n11105, n11106, n11107, n11108, n11109, n11110, n11111, n11112,
         n11113, n11114, n11115, n11116, n11117, n11118, n11119, n11120,
         n11121, n11122, n11123, n11124, n11125, n11126, n11127, n11128,
         n11129, n11130, n11131, n11132, n11133, n11134, n11135, n11136,
         n11137, n11138, n11139, n11140, n11141, n11142, n11143, n11144,
         n11145, n11146, n11147, n11148, n11149, n11150, n11151, n11152,
         n11153, n11154, n11155, n11156, n11157, n11158, n11159, n11160,
         n11161, n11162, n11163, n11164, n11165, n11166, n11167, n11168,
         n11169, n11170, n11171, n11172, n11173, n11174, n11175, n11176,
         n11177, n11178, n11179, n11180, n11181, n11182, n11183, n11184,
         n11185, n11186, n11187, n11188, n11189, n11190, n11191, n11192,
         n11193, n11194, n11195, n11196, n11197, n11198, n11199, n11200,
         n11201, n11202, n11203, n11204, n11205, n11206, n11207, n11208,
         n11209, n11210, n11211, n11212, n11213, n11214, n11215, n11216,
         n11217, n11218, n11219, n11220, n11221, n11222, n11223, n11224,
         n11225, n11226, n11227, n11228, n11229, n11230, n11231, n11232,
         n11233, n11234, n11235, n11236, n11237, n11238, n11239, n11240,
         n11241, n11242, n11243, n11244, n11245, n11246, n11247, n11248,
         n11249, n11250, n11251, n11252, n11253, n11254, n11255, n11256,
         n11257, n11258, n11259, n11260, n11261, n11262, n11263, n11264,
         n11265, n11266, n11267, n11268, n11269, n11270, n11271, n11272,
         n11273, n11274, n11275, n11276, n11277, n11278, n11279, n11280,
         n11281, n11282, n11283, n11284, n11285, n11286, n11287, n11288,
         n11289, n11290, n11291, n11292, n11293, n11294, n11295, n11296,
         n11297, n11298, n11299, n11300, n11301, n11302, n11303, n11304,
         n11305, n11306, n11307, n11308, n11309, n11310, n11311, n11312,
         n11313, n11314, n11315, n11316, n11317, n11318, n11319, n11320,
         n11321, n11322, n11323, n11324, n11325, n11326, n11327, n11328,
         n11329, n11330, n11331, n11332, n11333, n11334, n11335, n11336,
         n11337, n11338, n11339, n11340, n11341, n11342, n11343, n11344,
         n11345, n11346, n11347, n11348, n11349, n11350, n11351, n11352,
         n11353, n11354, n11355, n11356, n11357, n11358, n11359, n11360,
         n11361, n11362, n11363, n11364, n11365, n11366, n11367, n11368,
         n11369, n11370, n11371, n11372, n11373, n11374, n11375, n11376,
         n11377, n11378, n11379, n11380, n11381, n11382, n11383, n11384,
         n11385, n11386, n11387, n11388, n11389, n11390, n11391, n11392,
         n11393, n11394, n11395, n11396, n11397, n11398, n11399, n11400,
         n11401, n11402, n11403, n11404, n11405, n11406, n11407, n11408,
         n11409, n11410, n11411, n11412, n11413, n11414, n11415, n11416,
         n11417, n11418, n11419, n11420, n11421, n11422, n11423, n11424,
         n11425, n11426, n11427, n11428, n11429, n11430, n11431, n11432,
         n11433, n11434, n11435, n11436, n11437, n11438, n11439, n11440,
         n11441, n11442, n11443, n11444, n11445, n11446, n11447, n11448,
         n11449, n11450, n11451, n11452, n11453, n11454, n11455, n11456,
         n11457, n11458, n11459, n11460, n11461, n11462, n11463, n11464,
         n11465, n11466, n11467, n11468, n11469, n11470, n11471, n11472,
         n11473, n11474, n11475, n11476, n11477, n11478, n11479, n11480,
         n11481, n11482, n11483, n11484, n11485, n11486, n11487, n11488,
         n11489, n11490, n11491, n11492, n11493, n11494, n11495, n11496,
         n11497, n11498, n11499, n11500, n11501, n11502, n11503, n11504,
         n11505, n11506, n11507, n11508, n11509, n11510, n11511, n11512,
         n11513, n11514, n11515, n11516, n11517, n11518, n11519, n11520,
         n11521, n11522, n11523, n11524, n11525, n11526, n11527, n11528,
         n11529, n11530, n11531, n11532, n11533, n11534, n11535, n11536,
         n11537, n11538, n11539, n11540, n11541, n11542, n11543, n11544,
         n11545, n11546, n11547, n11548, n11549, n11550, n11551, n11552,
         n11553, n11554, n11555, n11556, n11557, n11558, n11559, n11560,
         n11561, n11562, n11563, n11564, n11565, n11566, n11567, n11568,
         n11569, n11570, n11571, n11572, n11573, n11574, n11575, n11576,
         n11577, n11578, n11579, n11580, n11581, n11582, n11583, n11584,
         n11585, n11586, n11587, n11588, n11589, n11590, n11591, n11592,
         n11593, n11594, n11595, n11596, n11597, n11598, n11599, n11600,
         n11601, n11602, n11603, n11604, n11605, n11606, n11607, n11608,
         n11609, n11610, n11611, n11612, n11613, n11614, n11615, n11616,
         n11617, n11618, n11619, n11620, n11621, n11622, n11623, n11624,
         n11625, n11626, n11627, n11628, n11629, n11630, n11631, n11632,
         n11633, n11634, n11635, n11636, n11637, n11638, n11639, n11640,
         n11641, n11642, n11643, n11644, n11645, n11646, n11647, n11648,
         n11649, n11650, n11651, n11652, n11653, n11654, n11655, n11656,
         n11657, n11658, n11659, n11660, n11661, n11662, n11663, n11664,
         n11665, n11666, n11667, n11668, n11669, n11670, n11671, n11672,
         n11673, n11674, n11675, n11676, n11677, n11678, n11679, n11680,
         n11681, n11682, n11683, n11684, n11685, n11686, n11687, n11688,
         n11689, n11690, n11691, n11692, n11693, n11694, n11695, n11696,
         n11697, n11698, n11699, n11700, n11701, n11702, n11703, n11704,
         n11705, n11706, n11707, n11708, n11709, n11710, n11711, n11712,
         n11713, n11714, n11715, n11716, n11717, n11718, n11719, n11720,
         n11721, n11722, n11723, n11724, n11725, n11726, n11727, n11728,
         n11729, n11730, n11731, n11732, n11733, n11734, n11735, n11736,
         n11737, n11738, n11739, n11740, n11741, n11742, n11743, n11744,
         n11745, n11746, n11747, n11748, n11749, n11750, n11751, n11752,
         n11753, n11754, n11755, n11756, n11757, n11758, n11759, n11760,
         n11761, n11762, n11763, n11764, n11765, n11766, n11767, n11768,
         n11769, n11770, n11771, n11772, n11773, n11774, n11775, n11776,
         n11777, n11778, n11779, n11780, n11781, n11782, n11783, n11784,
         n11785, n11786, n11787, n11788, n11789, n11790, n11791, n11792,
         n11793, n11794, n11795, n11796, n11797, n11798, n11799, n11800,
         n11801, n11802, n11803, n11804, n11805, n11806, n11807, n11808,
         n11809, n11810, n11811, n11812, n11813, n11814, n11815, n11816,
         n11817, n11818, n11819, n11820, n11821, n11822, n11823, n11824,
         n11825, n11826, n11827, n11828, n11829, n11830, n11831, n11832,
         n11833, n11834, n11835, n11836, n11837, n11838, n11839, n11840,
         n11841, n11842, n11843, n11844, n11845, n11846, n11847, n11848,
         n11849, n11850, n11851, n11852, n11853, n11854, n11855, n11856,
         n11857, n11858, n11859, n11860, n11861, n11862, n11863, n11864,
         n11865, n11866, n11867, n11868, n11869, n11870, n11871, n11872,
         n11873, n11874, n11875, n11876, n11877, n11878, n11879, n11880,
         n11881, n11882, n11883, n11884, n11885, n11886, n11887, n11888,
         n11889, n11890, n11891, n11892, n11893, n11894, n11895, n11896,
         n11897, n11898, n11899, n11900, n11901, n11902, n11903, n11904,
         n11905, n11906, n11907, n11908, n11909, n11910, n11911, n11912,
         n11913, n11914, n11915, n11916, n11917, n11918, n11919, n11920,
         n11921, n11922, n11923, n11924, n11925, n11926, n11927, n11928,
         n11929, n11930, n11931, n11932, n11933, n11934, n11935, n11936,
         n11937, n11938, n11939, n11940, n11941, n11942, n11943, n11944,
         n11945, n11946, n11947, n11948, n11949, n11950, n11951, n11952,
         n11953, n11954, n11955, n11956, n11957, n11958, n11959, n11960,
         n11961, n11962, n11963, n11964, n11965, n11966, n11967, n11968,
         n11969, n11970, n11971, n11972, n11973, n11974, n11975, n11976,
         n11977, n11978, n11979, n11980, n11981, n11982, n11983, n11984,
         n11985, n11986, n11987, n11988, n11989, n11990, n11991, n11992,
         n11993, n11994, n11995, n11996, n11997, n11998, n11999, n12000,
         n12001, n12002, n12003, n12004, n12005, n12006, n12007, n12008,
         n12009, n12010, n12011, n12012, n12013, n12014, n12015, n12016,
         n12017, n12018, n12019, n12020, n12021, n12022, n12023, n12024,
         n12025, n12026, n12027, n12028, n12029, n12030, n12031, n12032,
         n12033, n12034, n12035, n12036, n12037, n12038, n12039, n12040,
         n12041, n12042, n12043, n12044, n12045, n12046, n12047, n12048,
         n12049, n12050, n12051, n12052, n12053, n12054, n12055, n12056,
         n12057, n12058, n12059, n12060, n12061, n12062, n12063, n12064,
         n12065, n12066, n12067, n12068, n12069, n12070, n12071, n12072,
         n12073, n12074, n12075, n12076, n12077, n12078, n12079, n12080,
         n12081, n12082, n12083, n12084, n12085, n12086, n12087, n12088,
         n12089, n12090, n12091, n12092, n12093, n12094, n12095, n12096,
         n12097, n12098, n12099, n12100, n12101, n12102, n12103, n12104,
         n12105, n12106, n12107, n12108, n12109, n12110, n12111, n12112,
         n12113, n12114, n12115, n12116, n12117, n12118, n12119, n12120,
         n12121, n12122, n12123, n12124, n12125, n12126, n12127, n12128,
         n12129, n12130, n12131, n12132, n12133, n12134, n12135, n12136,
         n12137, n12138, n12139, n12140, n12141, n12142, n12143, n12144,
         n12145, n12146, n12147, n12148, n12149, n12150, n12151, n12152,
         n12153, n12154, n12155, n12156, n12157, n12158, n12159, n12160,
         n12161, n12162, n12163, n12164, n12165, n12166, n12167, n12168,
         n12169, n12170, n12171, n12172, n12173, n12174, n12175, n12176,
         n12177, n12178, n12179, n12180, n12181, n12182, n12183, n12184,
         n12185, n12186, n12187, n12188, n12189, n12190, n12191, n12192,
         n12193, n12194, n12195, n12196, n12197, n12198, n12199, n12200,
         n12201, n12202, n12203, n12204, n12205, n12206, n12207, n12208,
         n12209, n12210, n12211, n12212, n12213, n12214, n12215, n12216,
         n12217, n12218, n12219, n12220, n12221, n12222, n12223, n12224,
         n12225, n12226, n12227, n12228, n12229, n12230, n12231, n12232,
         n12233, n12234, n12235, n12236, n12237, n12238, n12239, n12240,
         n12241, n12242, n12243, n12244, n12245, n12246, n12247, n12248,
         n12249, n12250, n12251, n12252, n12253, n12254, n12255, n12256,
         n12257, n12258, n12259, n12260, n12261, n12262, n12263, n12264,
         n12265, n12266, n12267, n12268, n12269, n12270, n12271, n12272,
         n12273, n12274, n12275, n12276, n12277, n12278, n12279, n12280,
         n12281, n12282, n12283, n12284, n12285, n12286, n12287, n12288,
         n12289, n12290, n12291, n12292, n12293, n12294, n12295, n12296,
         n12297, n12298, n12299, n12300, n12301, n12302, n12303, n12304,
         n12305, n12306, n12307, n12308, n12309, n12310, n12311, n12312,
         n12313, n12314, n12315, n12316, n12317, n12318, n12319, n12320,
         n12321, n12322, n12323, n12324, n12325, n12326, n12327, n12328,
         n12329, n12330, n12331, n12332, n12333, n12334, n12335, n12336,
         n12337, n12338, n12339, n12340, n12341, n12342, n12343, n12344,
         n12345, n12346, n12347, n12348, n12349, n12350, n12351, n12352,
         n12353, n12354, n12355, n12356, n12357, n12358, n12359, n12360,
         n12361, n12362, n12363, n12364, n12365, n12366, n12367, n12368,
         n12369, n12370, n12371, n12372, n12373, n12374, n12375, n12376,
         n12377, n12378, n12379, n12380, n12381, n12382, n12383, n12384,
         n12385, n12386, n12387, n12388, n12389, n12390, n12391, n12392,
         n12393, n12394, n12395, n12396, n12397, n12398, n12399, n12400,
         n12401, n12402, n12403, n12404, n12405, n12406, n12407, n12408,
         n12409, n12410, n12411, n12412, n12413, n12414, n12415, n12416,
         n12417, n12418, n12419, n12420, n12421, n12422, n12423, n12424,
         n12425, n12426, n12427, n12428, n12429, n12430, n12431, n12432,
         n12433, n12434, n12435, n12436, n12437, n12438, n12439, n12440,
         n12441, n12442, n12443, n12444, n12445, n12446, n12447, n12448,
         n12449, n12450, n12451, n12452, n12453, n12454, n12455, n12456,
         n12457, n12458, n12459, n12460, n12461, n12462, n12463, n12464,
         n12465, n12466, n12467, n12468, n12469, n12470, n12471, n12472,
         n12473, n12474, n12475, n12476, n12477, n12478, n12479, n12480,
         n12481, n12482, n12483, n12484, n12485, n12486, n12487, n12488,
         n12489, n12490, n12491, n12492, n12493, n12494, n12495, n12496,
         n12497, n12498, n12499, n12500, n12501, n12502, n12503, n12504,
         n12505, n12506, n12507, n12508, n12509, n12510, n12511, n12512,
         n12513, n12514, n12515, n12516, n12517, n12518, n12519, n12520,
         n12521, n12522, n12523, n12524, n12525, n12526, n12527, n12528,
         n12529, n12530, n12531, n12532, n12533, n12534, n12535, n12536,
         n12537, n12538, n12539, n12540, n12541, n12542, n12543, n12544,
         n12545, n12546, n12547, n12548, n12549, n12550, n12551, n12552,
         n12553, n12554, n12555, n12556, n12557, n12558, n12559, n12560,
         n12561, n12562, n12563, n12564, n12565, n12566, n12567, n12568,
         n12569, n12570, n12571, n12572, n12573, n12574, n12575, n12576,
         n12577, n12578, n12579, n12580, n12581, n12582, n12583, n12584,
         n12585, n12586, n12587, n12588, n12589, n12590, n12591, n12592,
         n12593, n12594, n12595, n12596, n12597, n12598, n12599, n12600,
         n12601, n12602, n12603, n12604, n12605, n12606, n12607, n12608,
         n12609, n12610, n12611, n12612, n12613, n12614, n12615, n12616,
         n12617, n12618, n12619, n12620, n12621, n12622, n12623, n12624,
         n12625, n12626, n12627, n12628, n12629, n12630, n12631, n12632,
         n12633, n12634, n12635, n12636, n12637, n12638, n12639, n12640,
         n12641, n12642, n12643, n12644, n12645, n12646, n12647, n12648,
         n12649, n12650, n12651, n12652, n12653, n12654, n12655, n12656,
         n12657, n12658, n12659, n12660, n12661, n12662, n12663, n12664,
         n12665, n12666, n12667, n12668, n12669, n12670, n12671, n12672,
         n12673, n12674, n12675, n12676, n12677, n12678, n12679, n12680,
         n12681, n12682, n12683, n12684, n12685, n12686, n12687, n12688,
         n12689, n12690, n12691, n12692, n12693, n12694, n12695, n12696,
         n12697, n12698, n12699, n12700, n12701, n12702, n12703, n12704,
         n12705, n12706, n12707, n12708, n12709, n12710, n12711, n12712,
         n12713, n12714, n12715, n12716, n12717, n12718, n12719, n12720,
         n12721, n12722, n12723, n12724, n12725, n12726, n12727, n12728,
         n12729, n12730, n12731, n12732, n12733, n12734, n12735, n12736,
         n12737, n12738, n12739, n12740, n12741, n12742, n12743, n12744,
         n12745, n12746, n12747, n12748, n12749, n12750, n12751, n12752,
         n12753, n12754, n12755, n12756, n12757, n12758, n12759, n12760,
         n12761, n12762, n12763, n12764, n12765, n12766, n12767, n12768,
         n12769, n12770, n12771, n12772, n12773, n12774, n12775, n12776,
         n12777, n12778, n12779, n12780, n12781, n12782, n12783, n12784,
         n12785, n12786, n12787, n12788, n12789, n12790, n12791, n12792,
         n12793, n12794, n12795, n12796, n12797, n12798, n12799, n12800,
         n12801, n12802, n12803, n12804, n12805, n12806, n12807, n12808,
         n12809, n12810, n12811, n12812, n12813, n12814, n12815, n12816,
         n12817, n12818, n12819, n12820, n12821, n12822, n12823, n12824,
         n12825, n12826, n12827, n12828, n12829, n12830, n12831, n12832,
         n12833, n12834, n12835, n12836, n12837, n12838, n12839, n12840,
         n12841, n12842, n12843, n12844, n12845, n12846, n12847, n12848,
         n12849, n12850, n12851, n12852, n12853, n12854, n12855, n12856,
         n12857, n12858, n12859, n12860, n12861, n12862, n12863, n12864,
         n12865, n12866, n12867, n12868, n12869, n12870, n12871, n12872,
         n12873, n12874, n12875, n12876, n12877, n12878, n12879, n12880,
         n12881, n12882, n12883, n12884, n12885, n12886, n12887, n12888,
         n12889, n12890, n12891, n12892, n12893, n12894, n12895, n12896,
         n12897, n12898, n12899, n12900, n12901, n12902, n12903, n12904,
         n12905, n12906, n12907, n12908, n12909, n12910, n12911, n12912,
         n12913, n12914, n12915, n12916, n12917, n12918, n12919, n12920,
         n12921, n12922, n12923, n12924, n12925, n12926, n12927, n12928,
         n12929, n12930, n12931, n12932, n12933, n12934, n12935, n12936,
         n12937, n12938, n12939, n12940, n12941, n12942, n12943, n12944,
         n12945, n12946, n12947, n12948, n12949, n12950, n12951, n12952,
         n12953, n12954, n12955, n12956, n12957, n12958, n12959, n12960,
         n12961, n12962, n12963, n12964, n12965, n12966, n12967, n12968,
         n12969, n12970, n12971, n12972, n12973, n12974, n12975, n12976,
         n12977, n12978, n12979, n12980, n12981, n12982, n12983, n12984,
         n12985, n12986, n12987, n12988, n12989, n12990, n12991, n12992,
         n12993, n12994, n12995, n12996, n12997, n12998, n12999, n13000,
         n13001, n13002, n13003, n13004, n13005, n13006, n13007, n13008,
         n13009, n13010, n13011, n13012, n13013, n13014, n13015, n13016,
         n13017, n13018, n13019, n13020, n13021, n13022, n13023, n13024,
         n13025, n13026, n13027, n13028, n13029, n13030, n13031, n13032,
         n13033, n13034, n13035, n13036, n13037, n13038, n13039, n13040,
         n13041, n13042, n13043, n13044, n13045, n13046, n13047, n13048,
         n13049, n13050, n13051, n13052, n13053, n13054, n13055, n13056,
         n13057, n13058, n13059, n13060, n13061, n13062, n13063, n13064,
         n13065, n13066, n13067, n13068, n13069, n13070, n13071, n13072,
         n13073, n13074, n13075, n13076, n13077, n13078, n13079, n13080,
         n13081, n13082, n13083, n13084, n13085, n13086, n13087, n13088,
         n13089, n13090, n13091, n13092, n13093, n13094, n13095, n13096,
         n13097, n13098, n13099, n13100, n13101, n13102, n13103, n13104,
         n13105, n13106, n13107, n13108, n13109, n13110, n13111, n13112,
         n13113, n13114, n13115, n13116, n13117, n13118, n13119, n13120,
         n13121, n13122, n13123, n13124, n13125, n13126, n13127, n13128,
         n13129, n13130, n13131, n13132, n13133, n13134, n13135, n13136,
         n13137, n13138, n13139, n13140, n13141, n13142, n13143, n13144,
         n13145, n13146, n13147, n13148, n13149, n13150, n13151, n13152,
         n13153, n13154, n13155, n13156, n13157, n13158, n13159, n13160,
         n13161, n13162, n13163, n13164, n13165, n13166, n13167, n13168,
         n13169, n13170, n13171, n13172, n13173, n13174, n13175, n13176,
         n13177, n13178, n13179, n13180, n13181, n13182, n13183, n13184,
         n13185, n13186, n13187, n13188, n13189, n13190, n13191, n13192,
         n13193, n13194, n13195, n13196, n13197, n13198, n13199, n13200,
         n13201, n13202, n13203, n13204, n13205, n13206, n13207, n13208,
         n13209, n13210, n13211, n13212, n13213, n13214, n13215, n13216,
         n13217, n13218, n13219, n13220, n13221, n13222, n13223, n13224,
         n13225, n13226, n13227, n13228, n13229, n13230, n13231, n13232,
         n13233, n13234, n13235, n13236, n13237, n13238, n13239, n13240,
         n13241, n13242, n13243, n13244, n13245, n13246, n13247, n13248,
         n13249, n13250, n13251, n13252, n13253, n13254, n13255, n13256,
         n13257, n13258, n13259, n13260, n13261, n13262, n13263, n13264,
         n13265, n13266, n13267, n13268, n13269, n13270, n13271, n13272,
         n13273, n13274, n13275, n13276, n13277, n13278, n13279, n13280,
         n13281, n13282, n13283, n13284, n13285, n13286, n13287, n13288,
         n13289, n13290, n13291, n13292, n13293, n13294, n13295, n13296,
         n13297, n13298, n13299, n13300, n13301, n13302, n13303, n13304,
         n13305, n13306, n13307, n13308, n13309, n13310, n13311, n13312,
         n13313, n13314, n13315, n13316, n13317, n13318, n13319, n13320,
         n13321, n13322, n13323, n13324, n13325, n13326, n13327, n13328,
         n13329, n13330, n13331, n13332, n13333, n13334, n13335, n13336,
         n13337, n13338, n13339, n13340, n13341, n13342, n13343, n13344,
         n13345, n13346, n13347, n13348, n13349, n13350, n13351, n13352,
         n13353, n13354, n13355, n13356, n13357, n13358, n13359, n13360,
         n13361, n13362, n13363, n13364, n13365, n13366, n13367, n13368,
         n13369, n13370, n13371, n13372, n13373, n13374, n13375, n13376,
         n13377, n13378, n13379, n13380, n13381, n13382, n13383, n13384,
         n13385, n13386, n13387, n13388, n13389, n13390, n13391, n13392,
         n13393, n13394, n13395, n13396, n13397, n13398, n13399, n13400,
         n13401, n13402, n13403, n13404, n13405, n13406, n13407, n13408,
         n13409, n13410, n13411, n13412, n13413, n13414, n13415, n13416,
         n13417, n13418, n13419, n13420, n13421, n13422, n13423, n13424,
         n13425, n13426, n13427, n13428, n13429, n13430, n13431, n13432,
         n13433, n13434, n13435, n13436, n13437, n13438, n13439, n13440,
         n13441, n13442, n13443, n13444, n13445, n13446, n13447, n13448,
         n13449, n13450, n13451, n13452, n13453, n13454, n13455, n13456,
         n13457, n13458, n13459, n13460, n13461, n13462, n13463, n13464,
         n13465, n13466, n13467, n13468, n13469, n13470, n13471, n13472,
         n13473, n13474, n13475, n13476, n13477, n13478, n13479, n13480,
         n13481, n13482, n13483, n13484, n13485, n13486, n13487, n13488,
         n13489, n13490, n13491, n13492, n13493, n13494, n13495, n13496,
         n13497, n13498, n13499, n13500, n13501, n13502, n13503, n13504,
         n13505, n13506, n13507, n13508, n13509, n13510, n13511, n13512,
         n13513, n13514, n13515, n13516, n13517, n13518, n13519, n13520,
         n13521, n13522, n13523, n13524, n13525, n13526, n13527, n13528,
         n13529, n13530, n13531, n13532, n13533, n13534, n13535, n13536,
         n13537, n13538, n13539, n13540, n13541, n13542, n13543, n13544,
         n13545, n13546, n13547, n13548, n13549, n13550, n13551, n13552,
         n13553, n13554, n13555, n13556, n13557, n13558, n13559, n13560,
         n13561, n13562, n13563, n13564, n13565, n13566, n13567, n13568,
         n13569, n13570, n13571, n13572, n13573, n13574, n13575, n13576,
         n13577, n13578, n13579, n13580, n13581, n13582, n13583, n13584,
         n13585, n13586, n13587, n13588, n13589, n13590, n13591, n13592,
         n13593, n13594, n13595, n13596, n13597, n13598, n13599, n13600,
         n13601, n13602, n13603, n13604, n13605, n13606, n13607, n13608,
         n13609, n13610, n13611, n13612, n13613, n13614, n13615, n13616,
         n13617, n13618, n13619, n13620, n13621, n13622, n13623, n13624,
         n13625, n13626, n13627, n13628, n13629, n13630, n13631, n13632,
         n13633, n13634, n13635, n13636, n13637, n13638, n13639, n13640,
         n13641, n13642, n13643, n13644, n13645, n13646, n13647, n13648,
         n13649, n13650, n13651, n13652, n13653, n13654, n13655, n13656,
         n13657, n13658, n13659, n13660, n13661, n13662, n13663, n13664,
         n13665, n13666, n13667, n13668, n13669, n13670, n13671, n13672,
         n13673, n13674, n13675, n13676, n13677, n13678, n13679, n13680,
         n13681, n13682, n13683, n13684, n13685, n13686, n13687, n13688,
         n13689, n13690, n13691, n13692, n13693, n13694, n13695, n13696,
         n13697, n13698, n13699, n13700, n13701, n13702, n13703, n13704,
         n13705, n13706, n13707, n13708, n13709, n13710, n13711, n13712,
         n13713, n13714, n13715, n13716, n13717, n13718, n13719, n13720,
         n13721, n13722, n13723, n13724, n13725, n13726, n13727, n13728,
         n13729, n13730, n13731, n13732, n13733, n13734, n13735, n13736,
         n13737, n13738, n13739, n13740, n13741, n13742, n13743, n13744,
         n13745, n13746, n13747, n13748, n13749, n13750, n13751, n13752,
         n13753, n13754, n13755, n13756, n13757, n13758, n13759, n13760,
         n13761, n13762, n13763, n13764, n13765, n13766, n13767, n13768,
         n13769, n13770, n13771, n13772, n13773, n13774, n13775, n13776,
         n13777, n13778, n13779, n13780, n13781, n13782, n13783, n13784,
         n13785, n13786, n13787, n13788, n13789, n13790, n13791, n13792,
         n13793, n13794, n13795, n13796, n13797, n13798, n13799, n13800,
         n13801, n13802, n13803, n13804, n13805, n13806, n13807, n13808,
         n13809, n13810, n13811, n13812, n13813, n13814, n13815, n13816,
         n13817, n13818, n13819, n13820, n13821, n13822, n13823, n13824,
         n13825, n13826, n13827, n13828, n13829, n13830, n13831, n13832,
         n13833, n13834, n13835, n13836, n13837, n13838, n13839, n13840,
         n13841, n13842, n13843, n13844, n13845, n13846, n13847, n13848,
         n13849, n13850, n13851, n13852, n13853, n13854, n13855, n13856,
         n13857, n13858, n13859, n13860, n13861, n13862, n13863, n13864,
         n13865, n13866, n13867, n13868, n13869, n13870, n13871, n13872,
         n13873, n13874, n13875, n13876, n13877, n13878, n13879, n13880,
         n13881, n13882, n13883, n13884, n13885, n13886, n13887, n13888,
         n13889, n13890, n13891, n13892, n13893, n13894, n13895, n13896,
         n13897, n13898, n13899, n13900, n13901, n13902, n13903, n13904,
         n13905, n13906, n13907, n13908, n13909, n13910, n13911, n13912,
         n13913, n13914, n13915, n13916, n13917, n13918, n13919, n13920,
         n13921, n13922, n13923, n13924, n13925, n13926, n13927, n13928,
         n13929, n13930, n13931, n13932, n13933, n13934, n13935, n13936,
         n13937, n13938, n13939, n13940, n13941, n13942, n13943, n13944,
         n13945, n13946, n13947, n13948, n13949, n13950, n13951, n13952,
         n13953, n13954, n13955, n13956, n13957, n13958, n13959, n13960,
         n13961, n13962, n13963, n13964, n13965, n13966, n13967, n13968,
         n13969, n13970, n13971, n13972, n13973, n13974, n13975, n13976,
         n13977, n13978, n13979, n13980, n13981, n13982, n13983, n13984,
         n13985, n13986, n13987, n13988, n13989, n13990, n13991, n13992,
         n13993, n13994, n13995, n13996, n13997, n13998, n13999, n14000,
         n14001, n14002, n14003, n14004, n14005, n14006, n14007, n14008,
         n14009, n14010, n14011, n14012, n14013, n14014, n14015, n14016,
         n14017, n14018, n14019, n14020, n14021, n14022, n14023, n14024,
         n14025, n14026, n14027, n14028, n14029, n14030, n14031, n14032,
         n14033, n14034, n14035, n14036, n14037, n14038, n14039, n14040,
         n14041, n14042, n14043, n14044, n14045, n14046, n14047, n14048,
         n14049, n14050, n14051, n14052, n14053, n14054, n14055, n14056,
         n14057, n14058, n14059, n14060, n14061, n14062, n14063, n14064,
         n14065, n14066, n14067, n14068, n14069, n14070, n14071, n14072,
         n14073, n14074, n14075, n14076, n14077, n14078, n14079, n14080,
         n14081, n14082, n14083, n14084, n14085, n14086, n14087, n14088,
         n14089, n14090, n14091, n14092, n14093, n14094, n14095, n14096,
         n14097, n14098, n14099, n14100, n14101, n14102, n14103, n14104,
         n14105, n14106, n14107, n14108, n14109, n14110, n14111, n14112,
         n14113, n14114, n14115, n14116, n14117, n14118, n14119, n14120,
         n14121, n14122, n14123, n14124, n14125, n14126, n14127, n14128,
         n14129, n14130, n14131, n14132, n14133, n14134, n14135, n14136,
         n14137, n14138, n14139, n14140, n14141, n14142, n14143, n14144,
         n14145, n14146, n14147, n14148, n14149, n14150, n14151, n14152,
         n14153, n14154, n14155, n14156, n14157, n14158, n14159, n14160,
         n14161, n14162, n14163, n14164, n14165, n14166, n14167, n14168,
         n14169, n14170, n14171, n14172, n14173, n14174, n14175, n14176,
         n14177, n14178, n14179, n14180, n14181, n14182, n14183, n14184,
         n14185, n14186, n14187, n14188, n14189, n14190, n14191, n14192,
         n14193, n14194, n14195, n14196, n14197, n14198, n14199, n14200,
         n14201, n14202, n14203, n14204, n14205, n14206, n14207, n14208,
         n14209, n14210, n14211, n14212, n14213, n14214, n14215, n14216,
         n14217, n14218, n14219, n14220, n14221, n14222, n14223, n14224,
         n14225, n14226, n14227, n14228, n14229, n14230, n14231, n14232,
         n14233, n14234, n14235, n14236, n14237, n14238, n14239, n14240,
         n14241, n14242, n14243, n14244, n14245, n14246, n14247, n14248,
         n14249, n14250, n14251, n14252, n14253, n14254, n14255, n14256,
         n14257, n14258, n14259, n14260, n14261, n14262, n14263, n14264,
         n14265, n14266, n14267, n14268, n14269, n14270, n14271, n14272,
         n14273, n14274, n14275, n14276, n14277, n14278, n14279, n14280,
         n14281, n14282, n14283, n14284, n14285, n14286, n14287, n14288,
         n14289, n14290, n14291, n14292, n14293, n14294, n14295, n14296,
         n14297, n14298, n14299, n14300, n14301, n14302, n14303, n14304,
         n14305, n14306, n14307, n14308, n14309, n14310, n14311, n14312,
         n14313, n14314, n14315, n14316, n14317, n14318, n14319, n14320,
         n14321, n14322, n14323, n14324, n14325, n14326, n14327, n14328,
         n14329, n14330, n14331, n14332, n14333, n14334, n14335, n14336,
         n14337, n14338, n14339, n14340, n14341, n14342, n14343, n14344,
         n14345, n14346, n14347, n14348, n14349, n14350, n14351, n14352,
         n14353, n14354, n14355, n14356, n14357, n14358, n14359, n14360,
         n14361, n14362, n14363, n14364, n14365, n14366, n14367, n14368,
         n14369, n14370, n14371, n14372, n14373, n14374, n14375, n14376,
         n14377, n14378, n14379, n14380, n14381, n14382, n14383, n14384,
         n14385, n14386, n14387, n14388, n14389, n14390, n14391, n14392,
         n14393, n14394, n14395, n14396, n14397, n14398, n14399, n14400,
         n14401, n14402, n14403, n14404, n14405, n14406, n14407, n14408,
         n14409, n14410, n14411, n14412, n14413, n14414, n14415, n14416,
         n14417, n14418, n14419, n14420, n14421, n14422, n14423, n14424,
         n14425, n14426, n14427, n14428, n14429, n14430, n14431, n14432,
         n14433, n14434, n14435, n14436, n14437, n14438, n14439, n14440,
         n14441, n14442, n14443, n14444, n14445, n14446, n14447, n14448,
         n14449, n14450, n14451, n14452, n14453, n14454, n14455, n14456,
         n14457, n14458, n14459, n14460, n14461, n14462, n14463, n14464,
         n14465, n14466, n14467, n14468, n14469, n14470, n14471, n14472,
         n14473, n14474, n14475, n14476, n14477, n14478, n14479, n14480,
         n14481, n14482, n14483, n14484, n14485, n14486, n14487, n14488,
         n14489, n14490, n14491, n14492, n14493, n14494, n14495, n14496,
         n14497, n14498, n14499, n14500, n14501, n14502, n14503, n14504,
         n14505, n14506, n14507, n14508, n14509, n14510, n14511, n14512,
         n14513, n14514, n14515, n14516, n14517, n14518, n14519, n14520,
         n14521, n14522, n14523, n14524, n14525, n14526, n14527, n14528,
         n14529, n14530, n14531, n14532, n14533, n14534, n14535, n14536,
         n14537, n14538, n14539, n14540, n14541, n14542, n14543, n14544,
         n14545, n14546, n14547, n14548, n14549, n14550, n14551, n14552,
         n14553, n14554, n14555, n14556, n14557, n14558, n14559, n14560,
         n14561, n14562, n14563, n14564, n14565, n14566, n14567, n14568,
         n14569, n14570, n14571, n14572, n14573, n14574, n14575, n14576,
         n14577, n14578, n14579, n14580, n14581, n14582, n14583, n14584,
         n14585, n14586, n14587, n14588, n14589, n14590, n14591, n14592,
         n14593, n14594, n14595, n14596, n14597, n14598, n14599, n14600,
         n14601, n14602, n14603, n14604, n14605, n14606, n14607, n14608,
         n14609, n14610, n14611, n14612, n14613, n14614, n14615, n14616,
         n14617, n14618, n14619, n14620, n14621, n14622, n14623, n14624,
         n14625, n14626, n14627, n14628, n14629, n14630, n14631, n14632,
         n14633, n14634, n14635, n14636, n14637, n14638, n14639, n14640,
         n14641, n14642, n14643, n14644, n14645, n14646, n14647, n14648,
         n14649, n14650, n14651, n14652, n14653, n14654, n14655, n14656,
         n14657, n14658, n14659, n14660, n14661, n14662, n14663, n14664,
         n14665, n14666, n14667, n14668, n14669, n14670, n14671, n14672,
         n14673, n14674, n14675, n14676, n14677, n14678, n14679, n14680,
         n14681, n14682, n14683, n14684, n14685, n14686, n14687, n14688,
         n14689, n14690, n14691, n14692, n14693, n14694, n14695, n14696,
         n14697, n14698, n14699, n14700, n14701, n14702, n14703, n14704,
         n14705, n14706, n14707, n14708, n14709, n14710, n14711, n14712,
         n14713, n14714, n14715, n14716, n14717, n14718, n14719, n14720,
         n14721, n14722, n14723, n14724, n14725, n14726, n14727, n14728,
         n14729, n14730, n14731, n14732, n14733, n14734, n14735, n14736,
         n14737, n14738, n14739, n14740, n14741, n14742, n14743, n14744,
         n14745, n14746, n14747, n14748, n14749, n14750, n14751, n14752,
         n14753, n14754, n14755, n14756, n14757, n14758, n14759, n14760,
         n14761, n14762, n14763, n14764, n14765, n14766, n14767, n14768,
         n14769, n14770, n14771, n14772, n14773, n14774, n14775, n14776,
         n14777, n14778, n14779, n14780, n14781, n14782, n14783, n14784,
         n14785, n14786, n14787, n14788, n14789, n14790, n14791, n14792,
         n14793, n14794, n14795, n14796, n14797, n14798, n14799, n14800,
         n14801, n14802, n14803, n14804, n14805, n14806, n14807, n14808,
         n14809, n14810, n14811, n14812, n14813, n14814, n14815, n14816,
         n14817, n14818, n14819, n14820, n14821, n14822, n14823, n14824,
         n14825, n14826, n14827, n14828, n14829, n14830, n14831, n14832,
         n14833, n14834, n14835, n14836, n14837, n14838, n14839, n14840,
         n14841, n14842, n14843, n14844, n14845, n14846, n14847, n14848,
         n14849, n14850, n14851, n14852, n14853, n14854, n14855, n14856,
         n14857, n14858, n14859, n14860, n14861, n14862, n14863, n14864,
         n14865, n14866, n14867, n14868, n14869, n14870, n14871, n14872,
         n14873, n14874, n14875, n14876, n14877, n14878, n14879, n14880,
         n14881, n14882, n14883, n14884, n14885, n14886, n14887, n14888,
         n14889, n14890, n14891, n14892, n14893, n14894, n14895, n14896,
         n14897, n14898, n14899, n14900, n14901, n14902, n14903, n14904,
         n14905, n14906, n14907, n14908, n14909, n14910, n14911, n14912,
         n14913, n14914, n14915, n14916, n14917, n14918, n14920, n14921,
         n14922, n14923, n14924, n14925, n14926, n14927, n14928, n14929,
         n14930, n14931, n14932, n14933, n14934, n14935, n14936, n14937,
         n14938, n14939, n14940, n14941, n14942, n14943, n14944, n14945,
         n14946, n14947, n14948, n14949, n14950, n14951, n14952, n14953,
         n14954, n14955, n14956, n14957, n14958, n14959, n14960, n14961,
         n14962, n14963, n14964, n14965, n14966, n14967, n14968, n14969,
         n14970, n14971, n14972, n14973, n14974, n14975, n14976, n14977,
         n14978, n14979, n14980, n14981, n14982, n14983, n14984, n14985,
         n14986, n14987, n14988, n14989, n14990, n14991, n14992, n14993,
         n14994, n14995, n14996, n14997, n14998, n14999, n15000, n15001,
         n15002, n15003, n15004, n15005, n15006, n15007, n15008, n15009,
         n15010, n15011, n15012, n15013, n15014, n15015, n15016, n15017,
         n15018, n15019, n15020, n15021, n15022, n15023, n15024, n15025,
         n15026, n15027, n15028, n15029, n15030, n15031, n15032, n15033,
         n15034, n15035, n15036, n15037, n15038, n15039, n15040, n15041,
         n15042, n15043, n15044, n15045, n15046, n15047, n15048, n15049,
         n15050, n15051, n15052, n15053, n15054, n15055, n15056, n15057,
         n15058, n15059, n15060, n15061, n15062, n15063, n15064, n15065,
         n15066, n15067, n15068, n15069, n15070, n15071, n15072, n15073,
         n15074, n15075, n15076, n15077, n15078, n15079, n15080, n15081,
         n15082, n15083, n15084, n15085, n15086, n15087, n15088, n15089,
         n15090, n15091, n15092, n15093, n15094, n15095, n15096, n15097,
         n15098, n15099, n15100, n15101, n15102, n15103, n15104, n15105,
         n15106, n15107, n15108, n15109, n15110, n15111, n15112, n15113,
         n15114, n15115, n15116, n15117, n15118, n15119, n15120, n15121,
         n15122, n15123, n15124, n15125, n15126, n15127, n15128, n15129,
         n15130, n15131, n15132, n15133, n15134, n15135, n15136, n15137,
         n15138, n15139, n15140, n15141, n15142, n15143, n15144, n15145,
         n15146, n15147, n15148, n15149, n15150, n15151, n15152, n15153,
         n15154, n15155, n15156, n15157, n15158, n15159, n15160, n15161,
         n15162, n15163, n15164, n15165, n15166, n15167, n15168, n15169,
         n15170, n15171, n15172, n15173, n15174, n15175, n15176, n15177,
         n15178, n15179, n15180, n15181, n15182, n15183, n15184, n15185,
         n15186, n15187, n15188, n15189, n15190, n15191, n15192, n15193,
         n15194, n15195, n15196, n15197, n15198, n15199, n15200, n15201,
         n15202, n15203, n15204, n15205, n15206, n15207, n15208, n15209,
         n15210, n15211, n15212, n15213, n15214, n15215, n15216, n15217,
         n15218, n15219, n15220, n15221, n15222, n15223, n15224, n15225,
         n15226, n15227, n15228, n15229, n15230, n15231, n15232, n15233,
         n15234, n15235, n15236, n15237, n15238, n15239, n15240, n15241,
         n15242, n15243, n15244, n15245, n15246, n15247, n15248, n15249,
         n15250, n15251, n15252, n15253, n15254, n15255, n15256, n15257,
         n15258, n15259, n15260, n15261, n15262, n15263, n15264, n15265,
         n15266, n15267, n15268, n15269, n15270, n15271, n15272, n15273,
         n15274, n15275, n15276, n15277, n15278, n15279, n15280, n15281,
         n15282, n15283, n15284, n15285, n15286, n15287, n15288, n15289,
         n15290, n15291, n15292, n15293, n15294, n15295, n15296, n15297,
         n15298, n15299, n15300, n15301, n15302, n15303, n15304, n15305,
         n15306, n15307, n15308, n15309, n15310, n15311, n15312, n15313,
         n15314, n15315, n15316, n15317, n15318, n15319, n15320, n15321,
         n15322, n15323, n15324, n15325, n15326, n15327, n15328, n15329,
         n15330, n15331, n15332, n15333, n15334, n15335, n15336, n15337,
         n15338, n15339, n15340, n15341, n15342, n15343, n15344, n15345,
         n15346, n15347, n15348, n15349, n15350, n15351, n15352, n15353,
         n15354, n15355, n15356, n15357, n15358, n15359, n15360, n15361,
         n15362, n15363, n15364, n15365, n15366, n15367, n15368, n15369,
         n15370, n15371, n15372, n15373, n15374, n15375, n15376, n15377,
         n15378, n15379, n15380, n15381, n15382, n15383, n15384, n15385,
         n15386, n15387, n15388, n15389, n15390, n15391, n15392, n15393,
         n15394, n15395, n15396, n15397, n15398, n15399, n15400, n15401,
         n15402, n15403, n15404, n15405, n15406, n15407, n15408, n15409,
         n15410, n15411, n15412, n15413, n15414, n15415, n15416, n15417,
         n15418, n15419, n15420, n15421, n15422, n15423, n15424, n15425,
         n15426, n15427, n15428, n15429, n15430, n15431, n15432, n15433,
         n15434, n15435, n15436, n15437, n15438, n15439, n15440, n15441,
         n15442, n15443, n15444, n15445, n15446, n15447, n15448, n15449,
         n15450, n15451, n15452, n15453, n15454, n15455, n15456, n15457,
         n15458, n15459, n15460, n15461, n15462, n15463, n15464, n15465,
         n15466, n15467, n15468, n15469, n15470, n15471, n15472, n15473,
         n15474, n15475, n15476, n15477, n15478, n15479, n15480, n15481,
         n15482, n15483, n15484, n15485, n15486, n15487, n15488, n15489,
         n15490, n15491, n15492, n15493, n15494, n15495, n15496, n15497,
         n15498, n15499, n15500, n15501, n15502, n15503, n15504, n15505,
         n15506, n15507, n15508, n15509, n15510, n15511, n15512, n15513,
         n15514, n15515, n15516, n15517, n15518, n15519, n15520, n15521,
         n15522, n15523, n15524, n15525, n15526, n15527, n15528, n15529,
         n15530, n15531, n15532, n15533, n15534, n15535, n15536, n15537,
         n15538, n15539, n15540, n15541, n15542, n15543, n15544, n15545,
         n15546, n15547, n15548, n15549, n15550, n15551, n15552, n15553,
         n15554, n15555, n15556, n15557, n15558, n15559, n15560, n15561,
         n15562, n15563, n15564, n15565, n15566, n15567, n15568, n15569,
         n15570, n15571, n15572, n15573, n15574, n15575, n15576, n15577,
         n15578, n15579, n15580, n15581, n15582, n15583, n15584, n15585,
         n15586, n15587, n15588, n15589, n15590, n15591, n15592, n15593,
         n15594, n15595, n15596, n15597, n15598, n15599, n15600, n15601,
         n15602, n15603, n15604, n15605, n15606, n15607, n15608, n15609,
         n15610, n15611, n15612, n15613, n15614, n15615, n15616, n15617,
         n15618, n15619, n15620, n15621, n15622, n15623, n15624, n15625,
         n15626, n15627, n15628, n15629, n15630, n15631, n15632, n15633,
         n15634, n15635, n15636, n15637, n15638, n15639, n15640, n15641,
         n15642, n15643, n15644, n15645, n15646, n15647, n15648, n15649,
         n15650, n15651, n15652, n15653, n15654, n15655, n15656, n15657,
         n15658, n15659, n15660, n15661, n15662, n15663, n15664, n15665,
         n15666, n15667, n15668, n15669, n15670, n15671, n15672, n15673,
         n15674, n15675, n15676, n15677, n15678, n15679, n15680, n15681,
         n15682, n15683, n15684, n15685, n15686, n15687, n15689, n15690,
         n15691, n15692, n15693, n15694, n15695, n15696, n15697, n15698,
         n15699, n15700, n15701, n15702, n15703, n15704, n15705, n15706,
         n15707, n15708, n15709, n15710, n15711, n15712, n15713, n15714,
         n15715, n15716, n15717, n15718, n15719, n15720, n15721, n15722,
         n15723, n15724, n15725, n15726, n15727, n15728, n15729, n15730,
         n15731, n15732, n15733, n15734, n15735, n15736, n15737, n15738,
         n15739, n15740, n15741, n15742, n15743, n15744, n15745, n15746,
         n15747, n15748, n15749, n15750, n15751, n15752, n15753, n15754,
         n15755, n15756, n15757, n15758, n15759, n15760, n15761, n15762,
         n15763, n15764, n15765, n15766, n15767, n15768, n15769, n15770,
         n15771, n15772, n15773, n15774, n15775, n15776, n15777, n15778,
         n15779, n15780, n15781, n15782, n15783, n15784, n15785, n15786,
         n15787, n15788, n15789, n15790, n15791, n15792, n15793, n15794,
         n15795, n15796, n15797, n15798, n15799, n15800, n15801, n15802,
         n15803, n15804, n15805, n15806, n15807, n15808, n15809, n15810,
         n15811, n15812, n15813, n15814, n15815, n15816, n15817, n15818,
         n15819, n15820, n15821, n15822, n15823, n15824, n15825, n15826,
         n15827, n15828, n15829, n15830, n15831, n15832, n15833, n15834,
         n15835, n15836, n15837, n15838, n15839, n15840, n15841, n15842,
         n15843, n15844, n15845, n15846, n15847, n15848, n15849, n15850,
         n15851, n15852, n15853, n15854, n15855, n15856, n15857, n15858,
         n15859, n15860, n15861, n15862, n15863, n15864, n15865, n15866,
         n15867, n15868, n15869, n15870, n15871, n15872, n15873, n15874,
         n15875, n15876, n15877, n15878, n15879, n15880, n15881, n15882,
         n15883, n15884, n15885, n15886, n15887, n15888, n15889, n15890,
         n15891, n15892, n15893, n15894, n15895, n15896, n15897, n15898,
         n15899, n15900, n15901, n15902, n15903, n15904, n15905, n15906,
         n15907, n15908, n15909, n15910, n15911, n15912, n15913, n15914,
         n15915, n15916, n15917, n15918, n15919, n15920, n15921, n15922,
         n15923, n15924, n15925, n15926, n15927, n15928, n15929, n15930,
         n15931, n15932, n15933, n15934, n15935, n15936, n15937, n15938,
         n15939, n15940, n15941, n15942, n15943, n15944, n15945, n15946,
         n15947, n15948, n15949, n15950, n15951, n15952, n15953, n15954,
         n15955, n15956, n15957, n15958, n15959, n15960, n15961, n15962,
         n15963, n15964, n15965, n15966, n15967, n15968, n15969, n15970,
         n15971, n15972, n15973, n15974, n15975, n15976, n15977, n15978,
         n15979, n15980, n15981, n15982, n15983, n15984, n15985, n15986,
         n15987, n15988, n15989, n15990, n15991, n15992, n15993, n15994,
         n15995, n15996, n15997, n15998, n15999, n16000, n16001, n16002,
         n16003, n16004, n16005, n16006, n16007, n16008, n16009, n16010,
         n16011, n16012, n16013, n16014, n16015, n16016, n16017, n16018,
         n16019, n16021, n16022, n16023, n16024, n16025, n16026, n16027,
         n16028, n16029, n16030, n16031, n16032, n16033, n16034, n16035,
         n16036, n16037, n16038, n16039, n16040, n16041, n16042, n16043,
         n16044, n16045, n16046, n16047, n16048, n16049, n16050, n16051,
         n16052, n16053, n16054, n16055, n16056, n16057, n16058, n16059,
         n16060, n16061, n16062, n16063, n16064, n16065, n16066, n16067,
         n16068, n16069, n16070, n16071, n16072, n16073, n16074, n16075,
         n16076, n16077, n16078, n16079, n16080, n16081, n16082, n16083,
         n16084, n16085, n16086, n16087, n16088, n16089, n16090, n16091,
         n16092, n16093, n16094, n16095, n16096, n16097, n16098, n16099,
         n16100, n16101, n16102, n16103, n16104, n16105, n16106;

  OR2_X1 U7295 ( .A1(n11830), .A2(n11829), .ZN(n15804) );
  NAND2_X1 U7296 ( .A1(n8538), .A2(n8537), .ZN(n14395) );
  AND3_X1 U7297 ( .A1(n12368), .A2(n12340), .A3(n7453), .ZN(n12567) );
  OR2_X1 U7298 ( .A1(n8423), .A2(n14013), .ZN(n8458) );
  INV_X1 U7299 ( .A(n15983), .ZN(n8585) );
  INV_X1 U7300 ( .A(n12028), .ZN(n15792) );
  INV_X1 U7301 ( .A(n14136), .ZN(n7190) );
  INV_X1 U7302 ( .A(n14316), .ZN(n14267) );
  NAND4_X2 U7304 ( .A1(n8933), .A2(n8932), .A3(n8931), .A4(n8930), .ZN(n16047)
         );
  BUF_X1 U7305 ( .A(n9526), .Z(n6552) );
  INV_X1 U7306 ( .A(n10123), .ZN(n10118) );
  NAND2_X1 U7307 ( .A1(n10064), .A2(n10067), .ZN(n12794) );
  NAND2_X1 U7308 ( .A1(n12097), .A2(n10011), .ZN(n11472) );
  INV_X1 U7309 ( .A(n8376), .ZN(n8554) );
  AND2_X1 U7310 ( .A1(n14899), .A2(n14904), .ZN(n8108) );
  XNOR2_X1 U7311 ( .A(n9471), .B(P1_IR_REG_22__SCAN_IN), .ZN(n15705) );
  NAND2_X2 U7312 ( .A1(n7791), .A2(n7792), .ZN(n15699) );
  AND2_X1 U7313 ( .A1(n9457), .A2(n6711), .ZN(n7791) );
  CLKBUF_X1 U7314 ( .A(n15118), .Z(n6547) );
  NOR2_X1 U7315 ( .A1(n10607), .A2(n10606), .ZN(n15118) );
  CLKBUF_X1 U7316 ( .A(n14614), .Z(n6548) );
  OAI21_X1 U7317 ( .B1(n10398), .B2(n10397), .A(n14736), .ZN(n14614) );
  INV_X1 U7318 ( .A(n14263), .ZN(n14238) );
  NAND2_X1 U7319 ( .A1(n11431), .A2(n10104), .ZN(n13482) );
  OR2_X1 U7320 ( .A1(n8784), .A2(n8697), .ZN(n9363) );
  INV_X1 U7321 ( .A(n8056), .ZN(n8141) );
  NAND2_X1 U7322 ( .A1(n8533), .A2(n8532), .ZN(n14749) );
  INV_X2 U7323 ( .A(n10348), .ZN(n10340) );
  INV_X1 U7324 ( .A(n15696), .ZN(n9450) );
  INV_X1 U7325 ( .A(n12140), .ZN(n10011) );
  INV_X1 U7326 ( .A(n11708), .ZN(n13487) );
  AND2_X1 U7327 ( .A1(n13533), .A2(P3_REG1_REG_13__SCAN_IN), .ZN(n13566) );
  INV_X1 U7329 ( .A(n14120), .ZN(n7166) );
  NAND2_X1 U7330 ( .A1(n6633), .A2(n13010), .ZN(n15434) );
  NAND3_X1 U7331 ( .A1(n6765), .A2(n12254), .A3(n12255), .ZN(n12256) );
  OAI21_X1 U7332 ( .B1(n6775), .B2(n6774), .A(n6772), .ZN(n13244) );
  AND3_X1 U7333 ( .A1(n13625), .A2(n13624), .A3(n13623), .ZN(n13626) );
  OR2_X1 U7334 ( .A1(n8796), .A2(n6998), .ZN(n8798) );
  AND2_X1 U7335 ( .A1(n10401), .A2(n10400), .ZN(n14743) );
  XNOR2_X1 U7336 ( .A(n8069), .B(P2_IR_REG_3__SCAN_IN), .ZN(n14428) );
  AOI21_X1 U7337 ( .B1(n15050), .B2(n15051), .A(n7971), .ZN(n14951) );
  OAI211_X1 U7338 ( .C1(n9812), .C2(n10702), .A(n9520), .B(n9519), .ZN(n11798)
         );
  NAND2_X1 U7339 ( .A1(n13032), .A2(n10036), .ZN(n15485) );
  NAND2_X1 U7340 ( .A1(n10060), .A2(n10059), .ZN(n15611) );
  OAI211_X1 U7341 ( .C1(n15551), .C2(n15874), .A(n15550), .B(n7060), .ZN(
        n15668) );
  INV_X1 U7342 ( .A(n13683), .ZN(n7128) );
  NOR2_X1 U7343 ( .A1(n13626), .A2(n13627), .ZN(n13644) );
  XNOR2_X1 U7344 ( .A(n8798), .B(n8797), .ZN(n11431) );
  NAND2_X1 U7345 ( .A1(n8560), .A2(n8559), .ZN(n14394) );
  INV_X1 U7346 ( .A(n14231), .ZN(n14877) );
  INV_X1 U7347 ( .A(n11798), .ZN(n15834) );
  OR2_X4 U7348 ( .A1(n16030), .A2(n16056), .ZN(n9402) );
  NAND2_X2 U7349 ( .A1(n7984), .A2(n15348), .ZN(n15347) );
  AND2_X2 U7350 ( .A1(n15378), .A2(n13017), .ZN(n7984) );
  OR2_X2 U7351 ( .A1(n9353), .A2(n10730), .ZN(n8915) );
  INV_X1 U7352 ( .A(n12091), .ZN(n15843) );
  NAND2_X2 U7353 ( .A1(n13338), .A2(n7538), .ZN(n13347) );
  NAND4_X4 U7354 ( .A1(n8029), .A2(n8028), .A3(n8026), .A4(n8027), .ZN(n8040)
         );
  BUF_X8 U7356 ( .A(n9957), .Z(n6550) );
  NAND2_X2 U7357 ( .A1(n6880), .A2(n9450), .ZN(n9957) );
  NAND2_X2 U7358 ( .A1(n6996), .A2(n8739), .ZN(n8836) );
  NOR2_X2 U7359 ( .A1(n15490), .A2(n15628), .ZN(n15471) );
  NAND2_X2 U7360 ( .A1(n8804), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n6784) );
  NAND2_X2 U7361 ( .A1(n15003), .A2(n10278), .ZN(n15050) );
  OAI222_X1 U7362 ( .A1(P3_U3151), .A2(n8808), .B1(n13102), .B2(n13972), .C1(
        n13971), .C2(n13970), .ZN(P3_U3267) );
  NAND2_X1 U7363 ( .A1(n8808), .A2(n8809), .ZN(n8912) );
  AOI21_X2 U7364 ( .B1(n14335), .B2(n8129), .A(n8128), .ZN(n12230) );
  CLKBUF_X1 U7365 ( .A(n9526), .Z(n6551) );
  OAI222_X1 U7368 ( .A1(P1_U3086), .A2(n15696), .B1(n15703), .B2(n15695), .C1(
        n15694), .C2(n15700), .ZN(P1_U3326) );
  XNOR2_X2 U7369 ( .A(n8904), .B(n8903), .ZN(n8905) );
  NAND2_X1 U7370 ( .A1(n7476), .A2(n7474), .ZN(n6554) );
  AND2_X4 U7371 ( .A1(n6805), .A2(n6803), .ZN(n8096) );
  XNOR2_X2 U7372 ( .A(n10144), .B(n7348), .ZN(n11859) );
  XNOR2_X1 U7373 ( .A(n15307), .B(n13021), .ZN(n15576) );
  AND2_X1 U7374 ( .A1(n7576), .A2(n10082), .ZN(n7575) );
  NAND2_X1 U7375 ( .A1(n7823), .A2(n6626), .ZN(n15352) );
  NAND2_X1 U7376 ( .A1(n13769), .A2(n7031), .ZN(n13760) );
  INV_X1 U7377 ( .A(n15301), .ZN(n15565) );
  NAND2_X1 U7378 ( .A1(n6985), .A2(n6986), .ZN(n12594) );
  AND2_X1 U7379 ( .A1(n6987), .A2(P3_REG2_REG_11__SCAN_IN), .ZN(n6985) );
  NAND2_X1 U7380 ( .A1(n9755), .A2(n9754), .ZN(n15616) );
  INV_X1 U7381 ( .A(n14697), .ZN(n14882) );
  NAND2_X2 U7382 ( .A1(n13358), .A2(n13361), .ZN(n13355) );
  NAND2_X1 U7383 ( .A1(n16048), .A2(n11600), .ZN(n16043) );
  OR2_X1 U7384 ( .A1(n11264), .A2(n7644), .ZN(n7643) );
  INV_X2 U7385 ( .A(n15099), .ZN(n7219) );
  INV_X1 U7386 ( .A(n15096), .ZN(n12199) );
  INV_X4 U7387 ( .A(n13468), .ZN(n13450) );
  NAND2_X1 U7388 ( .A1(n10607), .A2(n10117), .ZN(n10348) );
  NAND2_X1 U7389 ( .A1(n10607), .A2(n11472), .ZN(n10151) );
  NAND4_X1 U7390 ( .A1(n9016), .A2(n9015), .A3(n9014), .A4(n9013), .ZN(n13507)
         );
  INV_X1 U7391 ( .A(n14265), .ZN(n14316) );
  CLKBUF_X2 U7393 ( .A(n8108), .Z(n12989) );
  NOR2_X1 U7394 ( .A1(n8746), .A2(n7229), .ZN(n11315) );
  CLKBUF_X2 U7395 ( .A(n9506), .Z(n9947) );
  XNOR2_X1 U7396 ( .A(n9446), .B(n9445), .ZN(n9451) );
  CLKBUF_X1 U7397 ( .A(n10695), .Z(n7218) );
  AND2_X1 U7398 ( .A1(n6796), .A2(n6795), .ZN(n14374) );
  NAND2_X1 U7399 ( .A1(n7153), .A2(n15561), .ZN(n15670) );
  NAND2_X1 U7400 ( .A1(n9985), .A2(n7240), .ZN(n10010) );
  AND3_X1 U7401 ( .A1(n7063), .A2(n13075), .A3(n7062), .ZN(n15551) );
  NOR2_X1 U7402 ( .A1(n8651), .A2(n14516), .ZN(n14851) );
  NAND2_X1 U7403 ( .A1(n10083), .A2(n7575), .ZN(n13657) );
  OR2_X1 U7404 ( .A1(n13611), .A2(n7652), .ZN(n13625) );
  OR2_X1 U7405 ( .A1(n10084), .A2(n16034), .ZN(n7576) );
  NAND2_X1 U7406 ( .A1(n7807), .A2(n7806), .ZN(n7227) );
  XNOR2_X1 U7407 ( .A(n7061), .B(n13067), .ZN(n15545) );
  AOI21_X1 U7408 ( .B1(n9428), .B2(n9427), .A(n9426), .ZN(n9429) );
  NAND2_X1 U7409 ( .A1(n13052), .A2(n7991), .ZN(n15295) );
  NAND2_X1 U7410 ( .A1(n7023), .A2(n7027), .ZN(n15011) );
  XNOR2_X1 U7411 ( .A(n9414), .B(n6607), .ZN(n10113) );
  NAND2_X1 U7412 ( .A1(n14017), .A2(n6575), .ZN(n14083) );
  INV_X1 U7413 ( .A(n13590), .ZN(n6555) );
  OAI21_X1 U7414 ( .B1(n14017), .B2(n6634), .A(n7289), .ZN(n10556) );
  AOI21_X1 U7415 ( .B1(n6916), .B2(n13631), .A(n6915), .ZN(n7164) );
  XNOR2_X1 U7416 ( .A(n8830), .B(n8897), .ZN(n6916) );
  NAND2_X1 U7417 ( .A1(n8506), .A2(n7621), .ZN(n7620) );
  NAND2_X1 U7418 ( .A1(n15540), .A2(n7104), .ZN(n15666) );
  NAND2_X1 U7419 ( .A1(n13042), .A2(n7824), .ZN(n7823) );
  OR2_X1 U7420 ( .A1(n13633), .A2(n8829), .ZN(n8830) );
  AOI21_X1 U7421 ( .B1(n13990), .B2(n10531), .A(n10530), .ZN(n10532) );
  INV_X1 U7422 ( .A(n7105), .ZN(n7104) );
  NAND2_X1 U7423 ( .A1(n14556), .A2(n14560), .ZN(n14555) );
  NAND2_X1 U7424 ( .A1(n13703), .A2(n13710), .ZN(n9275) );
  NAND2_X1 U7425 ( .A1(n13173), .A2(n12960), .ZN(n12963) );
  NAND2_X1 U7426 ( .A1(n13212), .A2(n6782), .ZN(n13173) );
  INV_X1 U7427 ( .A(n7290), .ZN(n7289) );
  OAI21_X1 U7428 ( .B1(n15541), .B2(n15844), .A(n15542), .ZN(n7105) );
  OAI21_X1 U7429 ( .B1(n6575), .B2(n6634), .A(n10553), .ZN(n7290) );
  NAND2_X1 U7430 ( .A1(n13214), .A2(n13213), .ZN(n13212) );
  NOR2_X1 U7431 ( .A1(n15277), .A2(n15553), .ZN(n15280) );
  AOI21_X1 U7432 ( .B1(n7806), .B2(n13051), .A(n7808), .ZN(n7804) );
  NAND2_X1 U7433 ( .A1(n15430), .A2(n15434), .ZN(n13038) );
  NAND2_X1 U7434 ( .A1(n14546), .A2(n14531), .ZN(n14530) );
  NAND2_X1 U7435 ( .A1(n7825), .A2(n6658), .ZN(n15454) );
  NAND2_X1 U7436 ( .A1(n13760), .A2(n9210), .ZN(n13744) );
  OAI21_X1 U7437 ( .B1(n13572), .B2(n13604), .A(n13603), .ZN(n13602) );
  NAND3_X1 U7438 ( .A1(n7667), .A2(n7078), .A3(n14646), .ZN(n14649) );
  AND3_X1 U7439 ( .A1(n7707), .A2(P3_REG1_REG_15__SCAN_IN), .A3(n7717), .ZN(
        n13572) );
  NAND2_X1 U7440 ( .A1(n7623), .A2(n7624), .ZN(n14668) );
  INV_X1 U7441 ( .A(n13195), .ZN(n6775) );
  NAND2_X1 U7442 ( .A1(n14692), .A2(n8341), .ZN(n7623) );
  OAI22_X1 U7443 ( .A1(n13784), .A2(n7254), .B1(n7255), .B2(n13425), .ZN(
        n13742) );
  XNOR2_X1 U7444 ( .A(n6794), .B(n8531), .ZN(n14911) );
  NAND2_X1 U7445 ( .A1(n8283), .A2(n8282), .ZN(n14726) );
  AND2_X1 U7446 ( .A1(n8629), .A2(n14647), .ZN(n14657) );
  NAND2_X1 U7447 ( .A1(n9461), .A2(n9460), .ZN(n15597) );
  NAND2_X1 U7448 ( .A1(n8422), .A2(n8421), .ZN(n14628) );
  NAND2_X1 U7449 ( .A1(n9783), .A2(n9782), .ZN(n15605) );
  OAI21_X2 U7450 ( .B1(n14616), .B2(n8648), .A(n8465), .ZN(n14400) );
  AOI21_X1 U7451 ( .B1(n7814), .B2(n12555), .A(n7175), .ZN(n7811) );
  INV_X1 U7452 ( .A(n7333), .ZN(n12360) );
  NOR2_X1 U7453 ( .A1(n12855), .A2(n12854), .ZN(n12880) );
  AND2_X1 U7454 ( .A1(n13030), .A2(n9770), .ZN(n13029) );
  NAND2_X1 U7455 ( .A1(n8365), .A2(n8349), .ZN(n11973) );
  NAND2_X1 U7456 ( .A1(n9700), .A2(n9699), .ZN(n15639) );
  NAND2_X1 U7457 ( .A1(n8273), .A2(n8272), .ZN(n14824) );
  OAI21_X1 U7458 ( .B1(n12615), .B2(n7676), .A(n7674), .ZN(n12189) );
  NAND2_X1 U7459 ( .A1(n8334), .A2(n8333), .ZN(n14697) );
  NAND2_X1 U7460 ( .A1(n9144), .A2(n9143), .ZN(n13952) );
  NAND2_X1 U7461 ( .A1(n8200), .A2(n8199), .ZN(n14842) );
  NAND2_X1 U7462 ( .A1(n8183), .A2(n8182), .ZN(n14159) );
  OAI21_X1 U7463 ( .B1(n8344), .B2(n7883), .A(n7880), .ZN(n8474) );
  XNOR2_X1 U7464 ( .A(n8310), .B(SI_14_), .ZN(n7058) );
  NAND2_X2 U7465 ( .A1(n9634), .A2(n9633), .ZN(n15662) );
  NAND2_X1 U7466 ( .A1(n6935), .A2(n9107), .ZN(n9139) );
  AOI21_X1 U7467 ( .B1(n11643), .B2(n9405), .A(n9404), .ZN(n12098) );
  INV_X1 U7468 ( .A(n12246), .ZN(n13370) );
  NAND2_X1 U7469 ( .A1(n9672), .A2(n9671), .ZN(n12902) );
  NAND2_X1 U7470 ( .A1(n6988), .A2(n6990), .ZN(n7663) );
  OR2_X1 U7471 ( .A1(n13505), .A2(n12274), .ZN(n13379) );
  INV_X1 U7472 ( .A(n11958), .ZN(n11804) );
  AND3_X1 U7473 ( .A1(n9037), .A2(n9036), .A3(n9035), .ZN(n12274) );
  NAND2_X1 U7474 ( .A1(n8597), .A2(n8598), .ZN(n14335) );
  INV_X2 U7475 ( .A(n15528), .ZN(n6556) );
  NAND2_X1 U7476 ( .A1(n9603), .A2(n9602), .ZN(n15780) );
  INV_X2 U7477 ( .A(n11965), .ZN(n7220) );
  NAND2_X2 U7478 ( .A1(n9402), .A2(n13342), .ZN(n16052) );
  NAND4_X2 U7479 ( .A1(n8113), .A2(n8112), .A3(n8111), .A4(n8110), .ZN(n14416)
         );
  NAND4_X1 U7480 ( .A1(n8122), .A2(n8121), .A3(n8120), .A4(n8119), .ZN(n14417)
         );
  NAND2_X1 U7481 ( .A1(n9559), .A2(n9558), .ZN(n12091) );
  NAND2_X1 U7482 ( .A1(n7803), .A2(n9536), .ZN(n11965) );
  NAND3_X1 U7483 ( .A1(n7645), .A2(n7643), .A3(n7642), .ZN(n11244) );
  NAND2_X1 U7484 ( .A1(n8243), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n8260) );
  NAND2_X1 U7485 ( .A1(n8521), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n8112) );
  NAND2_X1 U7486 ( .A1(n8136), .A2(n8135), .ZN(n8153) );
  NAND2_X2 U7487 ( .A1(n11835), .A2(n10140), .ZN(n10342) );
  OR2_X1 U7488 ( .A1(n13509), .A2(n11974), .ZN(n13361) );
  AND3_X1 U7489 ( .A1(n9021), .A2(n9020), .A3(n9019), .ZN(n12245) );
  NAND4_X1 U7490 ( .A1(n8993), .A2(n8992), .A3(n8991), .A4(n8990), .ZN(n13506)
         );
  INV_X2 U7491 ( .A(n8141), .ZN(n12988) );
  OAI211_X1 U7492 ( .C1(n8981), .C2(n9367), .A(n8983), .B(n8982), .ZN(n11647)
         );
  NAND4_X1 U7493 ( .A1(n9054), .A2(n9053), .A3(n9052), .A4(n9051), .ZN(n13504)
         );
  NAND4_X2 U7494 ( .A1(n9028), .A2(n9027), .A3(n9026), .A4(n9025), .ZN(n13505)
         );
  NAND3_X1 U7495 ( .A1(n7969), .A2(n8973), .A3(n8970), .ZN(n11974) );
  INV_X2 U7496 ( .A(n10151), .ZN(n10346) );
  BUF_X2 U7497 ( .A(n10154), .Z(n10329) );
  NAND2_X2 U7498 ( .A1(n7737), .A2(n14379), .ZN(n13111) );
  AND2_X2 U7499 ( .A1(n13487), .A2(n13333), .ZN(n13468) );
  NAND4_X2 U7500 ( .A1(n8969), .A2(n8968), .A3(n8967), .A4(n8966), .ZN(n13509)
         );
  NAND2_X2 U7501 ( .A1(n10420), .A2(n14323), .ZN(n10436) );
  NAND4_X1 U7502 ( .A1(n9547), .A2(n9546), .A3(n9545), .A4(n9544), .ZN(n15795)
         );
  OAI21_X2 U7503 ( .B1(n7827), .B2(n7444), .A(n7443), .ZN(n7137) );
  AND2_X1 U7504 ( .A1(n14899), .A2(n8009), .ZN(n8056) );
  AND2_X1 U7505 ( .A1(n8008), .A2(n8009), .ZN(n8071) );
  INV_X2 U7506 ( .A(n8108), .ZN(n8557) );
  INV_X1 U7507 ( .A(n8062), .ZN(n8099) );
  INV_X4 U7508 ( .A(n11146), .ZN(n8368) );
  INV_X1 U7509 ( .A(n9367), .ZN(n9197) );
  CLKBUF_X1 U7510 ( .A(n9372), .Z(n7094) );
  NAND2_X1 U7511 ( .A1(n7475), .A2(n11750), .ZN(n7474) );
  NAND2_X1 U7512 ( .A1(n10356), .A2(n10071), .ZN(n10607) );
  BUF_X2 U7513 ( .A(n13292), .Z(n6568) );
  INV_X2 U7514 ( .A(n9812), .ZN(n10006) );
  CLKBUF_X1 U7515 ( .A(n8420), .Z(n7140) );
  INV_X2 U7516 ( .A(n9486), .ZN(n9524) );
  CLKBUF_X3 U7517 ( .A(n8974), .Z(n9372) );
  CLKBUF_X3 U7518 ( .A(n8036), .Z(n11146) );
  BUF_X2 U7519 ( .A(n8912), .Z(n9367) );
  INV_X1 U7520 ( .A(n6552), .ZN(n9838) );
  NAND2_X1 U7521 ( .A1(n7615), .A2(n7310), .ZN(n14904) );
  AND2_X1 U7522 ( .A1(n14329), .A2(n14105), .ZN(n14107) );
  AND2_X1 U7523 ( .A1(n10353), .A2(n12097), .ZN(n7133) );
  XNOR2_X1 U7525 ( .A(n9364), .B(P3_IR_REG_20__SCAN_IN), .ZN(n10104) );
  NAND2_X1 U7526 ( .A1(n9480), .A2(n9479), .ZN(n12097) );
  OR2_X1 U7527 ( .A1(n8185), .A2(n8184), .ZN(n8202) );
  NAND2_X1 U7528 ( .A1(n8020), .A2(n8021), .ZN(n11179) );
  NOR2_X1 U7529 ( .A1(n11299), .A2(n11298), .ZN(n11297) );
  MUX2_X1 U7530 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8022), .S(
        P2_IR_REG_27__SCAN_IN), .Z(n8025) );
  OAI211_X2 U7531 ( .C1(n8583), .C2(n8582), .A(n8658), .B(n8581), .ZN(n14379)
         );
  XNOR2_X1 U7532 ( .A(n8367), .B(P2_IR_REG_19__SCAN_IN), .ZN(n14322) );
  OAI211_X2 U7533 ( .C1(n8573), .C2(n8572), .A(n7537), .B(n7536), .ZN(n14329)
         );
  NAND2_X1 U7534 ( .A1(n13960), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8902) );
  XNOR2_X1 U7535 ( .A(n9473), .B(n9472), .ZN(n12140) );
  NAND2_X1 U7536 ( .A1(n8019), .A2(n8018), .ZN(n8020) );
  NAND2_X1 U7537 ( .A1(n9474), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7208) );
  NAND2_X2 U7538 ( .A1(n7218), .A2(P1_U3086), .ZN(n15703) );
  OR2_X1 U7539 ( .A1(n8571), .A2(n8569), .ZN(n7537) );
  OR2_X1 U7540 ( .A1(n9739), .A2(n9470), .ZN(n9476) );
  AND2_X1 U7541 ( .A1(n7970), .A2(n6887), .ZN(n6886) );
  AND2_X1 U7542 ( .A1(n7778), .A2(n7970), .ZN(n7777) );
  OR2_X1 U7543 ( .A1(n8743), .A2(P3_IR_REG_3__SCAN_IN), .ZN(n8732) );
  AND2_X1 U7544 ( .A1(n7862), .A2(n8903), .ZN(n7861) );
  AND3_X1 U7545 ( .A1(n6888), .A2(n9467), .A3(n9437), .ZN(n7778) );
  NOR2_X1 U7546 ( .A1(n8290), .A2(n7998), .ZN(n6969) );
  AND4_X1 U7547 ( .A1(n9442), .A2(n7053), .A3(n10061), .A4(n9443), .ZN(n7970)
         );
  AND3_X1 U7548 ( .A1(n7340), .A2(n7339), .A3(n7338), .ZN(n7780) );
  AND2_X1 U7549 ( .A1(n9438), .A2(n6802), .ZN(n6888) );
  NAND2_X1 U7550 ( .A1(n8005), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8018) );
  AND2_X1 U7551 ( .A1(n8707), .A2(n7569), .ZN(n7568) );
  AND2_X1 U7552 ( .A1(n9515), .A2(n9438), .ZN(n9531) );
  NOR2_X1 U7553 ( .A1(P1_IR_REG_5__SCAN_IN), .A2(P1_IR_REG_4__SCAN_IN), .ZN(
        n9462) );
  INV_X4 U7554 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  NOR2_X1 U7555 ( .A1(P3_IR_REG_21__SCAN_IN), .A2(P3_IR_REG_23__SCAN_IN), .ZN(
        n8703) );
  NOR3_X1 U7556 ( .A1(P3_IR_REG_17__SCAN_IN), .A2(P3_IR_REG_16__SCAN_IN), .A3(
        P3_IR_REG_24__SCAN_IN), .ZN(n8707) );
  NOR2_X1 U7557 ( .A1(P3_IR_REG_18__SCAN_IN), .A2(P3_IR_REG_22__SCAN_IN), .ZN(
        n8702) );
  INV_X1 U7558 ( .A(P3_IR_REG_7__SCAN_IN), .ZN(n8723) );
  INV_X1 U7559 ( .A(P3_IR_REG_8__SCAN_IN), .ZN(n8726) );
  NOR2_X1 U7560 ( .A1(P1_IR_REG_17__SCAN_IN), .A2(P1_IR_REG_20__SCAN_IN), .ZN(
        n9467) );
  NOR2_X1 U7561 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P1_IR_REG_16__SCAN_IN), .ZN(
        n9469) );
  NOR2_X1 U7562 ( .A1(P3_IR_REG_5__SCAN_IN), .A2(P3_IR_REG_4__SCAN_IN), .ZN(
        n8695) );
  NOR2_X1 U7563 ( .A1(P3_IR_REG_3__SCAN_IN), .A2(P3_IR_REG_2__SCAN_IN), .ZN(
        n8694) );
  NOR2_X2 U7564 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(P1_IR_REG_7__SCAN_IN), .ZN(
        n10816) );
  INV_X4 U7565 ( .A(P3_STATE_REG_SCAN_IN), .ZN(P3_U3151) );
  NOR2_X1 U7566 ( .A1(P1_IR_REG_15__SCAN_IN), .A2(P1_IR_REG_3__SCAN_IN), .ZN(
        n9437) );
  INV_X1 U7567 ( .A(P3_IR_REG_1__SCAN_IN), .ZN(n6770) );
  INV_X2 U7568 ( .A(P3_IR_REG_0__SCAN_IN), .ZN(n6771) );
  NOR2_X1 U7569 ( .A1(P3_IR_REG_17__SCAN_IN), .A2(P3_IR_REG_16__SCAN_IN), .ZN(
        n7485) );
  NOR2_X1 U7570 ( .A1(P3_IR_REG_14__SCAN_IN), .A2(P3_IR_REG_10__SCAN_IN), .ZN(
        n8691) );
  NOR2_X1 U7571 ( .A1(P1_IR_REG_12__SCAN_IN), .A2(P1_IR_REG_11__SCAN_IN), .ZN(
        n9441) );
  INV_X1 U7572 ( .A(P3_IR_REG_11__SCAN_IN), .ZN(n8762) );
  INV_X1 U7573 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n7339) );
  INV_X1 U7574 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n8575) );
  INV_X1 U7575 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n10965) );
  NOR2_X1 U7576 ( .A1(P2_IR_REG_2__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n7665) );
  NOR2_X1 U7577 ( .A1(P2_IR_REG_5__SCAN_IN), .A2(P2_IR_REG_8__SCAN_IN), .ZN(
        n7993) );
  NOR2_X1 U7578 ( .A1(P2_IR_REG_3__SCAN_IN), .A2(P2_IR_REG_4__SCAN_IN), .ZN(
        n7664) );
  INV_X1 U7579 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n8568) );
  INV_X1 U7580 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n8653) );
  INV_X1 U7581 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n8659) );
  NOR2_X1 U7582 ( .A1(P1_IR_REG_14__SCAN_IN), .A2(P1_IR_REG_13__SCAN_IN), .ZN(
        n9440) );
  INV_X4 U7583 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3088) );
  INV_X1 U7584 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n8158) );
  INV_X2 U7585 ( .A(P3_ADDR_REG_19__SCAN_IN), .ZN(n15768) );
  NAND2_X1 U7586 ( .A1(n12368), .A2(n15093), .ZN(n12553) );
  XNOR2_X1 U7587 ( .A(n8212), .B(n8211), .ZN(n11036) );
  AND3_X1 U7588 ( .A1(n7263), .A2(n7568), .A3(n8696), .ZN(n6557) );
  AND3_X1 U7589 ( .A1(n7263), .A2(n7568), .A3(n8696), .ZN(n6558) );
  NAND2_X1 U7590 ( .A1(n13744), .A2(n13329), .ZN(n6559) );
  AND3_X2 U7591 ( .A1(n8811), .A2(n8695), .A3(n8694), .ZN(n6560) );
  AND3_X1 U7592 ( .A1(n7263), .A2(n7568), .A3(n8696), .ZN(n8801) );
  NOR2_X4 U7593 ( .A1(n7174), .A2(n8693), .ZN(n8696) );
  NAND2_X1 U7594 ( .A1(n13744), .A2(n13329), .ZN(n13747) );
  AND3_X1 U7595 ( .A1(n8811), .A2(n8695), .A3(n8694), .ZN(n8722) );
  AND2_X2 U7596 ( .A1(n6771), .A2(n6770), .ZN(n8811) );
  OR2_X2 U7597 ( .A1(n8906), .A2(n8905), .ZN(n8974) );
  INV_X1 U7598 ( .A(n8906), .ZN(n13103) );
  INV_X1 U7599 ( .A(n8905), .ZN(n8907) );
  AND2_X2 U7600 ( .A1(n14696), .A2(n14681), .ZN(n14676) );
  INV_X2 U7601 ( .A(n9555), .ZN(n6561) );
  AND2_X1 U7602 ( .A1(n9514), .A2(n10696), .ZN(n9513) );
  NAND2_X2 U7603 ( .A1(n9042), .A2(n9041), .ZN(n12113) );
  NAND2_X2 U7604 ( .A1(n13790), .A2(n6596), .ZN(n13769) );
  AND2_X1 U7605 ( .A1(n6560), .A2(n7485), .ZN(n7110) );
  OR2_X2 U7606 ( .A1(n6563), .A2(n8836), .ZN(n8914) );
  OAI222_X1 U7607 ( .A1(P3_U3151), .A2(n6771), .B1(n13102), .B2(n10736), .C1(
        n10735), .C2(n13962), .ZN(P3_U3295) );
  OAI222_X1 U7608 ( .A1(n13970), .A2(n13291), .B1(P3_U3151), .B2(n13103), .C1(
        n13102), .C2(n13101), .ZN(P3_U3265) );
  NAND2_X2 U7609 ( .A1(n13103), .A2(n8905), .ZN(n9007) );
  NAND2_X1 U7610 ( .A1(n8808), .A2(n8809), .ZN(n6562) );
  NAND2_X1 U7611 ( .A1(n8808), .A2(n8809), .ZN(n6563) );
  NAND2_X1 U7612 ( .A1(n8928), .A2(n8927), .ZN(n16025) );
  NAND2_X1 U7613 ( .A1(n13103), .A2(n8905), .ZN(n6565) );
  NOR2_X2 U7614 ( .A1(n12917), .A2(n14824), .ZN(n14730) );
  INV_X2 U7615 ( .A(n16047), .ZN(n7260) );
  INV_X1 U7616 ( .A(n9007), .ZN(n6566) );
  INV_X1 U7617 ( .A(n9007), .ZN(n6567) );
  NAND2_X1 U7618 ( .A1(n7845), .A2(n7843), .ZN(n12498) );
  NAND2_X2 U7619 ( .A1(n12701), .A2(n12700), .ZN(n12699) );
  NAND2_X4 U7620 ( .A1(n7476), .A2(n7474), .ZN(n11436) );
  NAND2_X2 U7621 ( .A1(n8941), .A2(n8940), .ZN(n11638) );
  NAND2_X2 U7622 ( .A1(n7839), .A2(n7838), .ZN(n13800) );
  NAND3_X2 U7623 ( .A1(n7120), .A2(n8986), .A3(n8985), .ZN(n11868) );
  NAND2_X1 U7624 ( .A1(n6562), .A2(n10696), .ZN(n13292) );
  OR2_X1 U7625 ( .A1(n13911), .A2(n13733), .ZN(n13441) );
  INV_X1 U7626 ( .A(n9157), .ZN(n7593) );
  AOI21_X1 U7627 ( .B1(n7527), .B2(n7526), .A(n7524), .ZN(n7523) );
  NAND2_X1 U7628 ( .A1(n7866), .A2(n7865), .ZN(n9976) );
  OR2_X1 U7629 ( .A1(n9953), .A2(n9954), .ZN(n7865) );
  NAND2_X1 U7630 ( .A1(n9942), .A2(n7867), .ZN(n7866) );
  NOR2_X1 U7631 ( .A1(n9953), .A2(n7868), .ZN(n7867) );
  OAI21_X1 U7632 ( .B1(n8096), .B2(n10655), .A(n7167), .ZN(n8094) );
  NAND2_X1 U7633 ( .A1(n8096), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n7167) );
  NAND2_X1 U7634 ( .A1(n10628), .A2(n10629), .ZN(n7500) );
  INV_X2 U7635 ( .A(n9007), .ZN(n13285) );
  NAND2_X1 U7636 ( .A1(n7250), .A2(n7252), .ZN(n7249) );
  AND2_X1 U7637 ( .A1(n7557), .A2(n7251), .ZN(n7250) );
  INV_X1 U7638 ( .A(n7592), .ZN(n7591) );
  OAI21_X1 U7639 ( .B1(n9155), .B2(n7593), .A(n9168), .ZN(n7592) );
  NAND2_X1 U7640 ( .A1(n14657), .A2(n6573), .ZN(n7669) );
  INV_X1 U7641 ( .A(n9451), .ZN(n6880) );
  NAND2_X1 U7642 ( .A1(n9968), .A2(n9967), .ZN(n10005) );
  INV_X1 U7643 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n10061) );
  NAND2_X1 U7644 ( .A1(n8529), .A2(n6646), .ZN(n8530) );
  OAI21_X1 U7645 ( .B1(n8231), .B2(n8230), .A(n8229), .ZN(n8252) );
  INV_X1 U7646 ( .A(n9311), .ZN(n9368) );
  INV_X1 U7647 ( .A(n9126), .ZN(n9355) );
  NAND2_X1 U7648 ( .A1(n6925), .A2(n7246), .ZN(n6924) );
  NAND2_X1 U7649 ( .A1(n7244), .A2(n7242), .ZN(n6926) );
  XNOR2_X1 U7650 ( .A(n13460), .B(n13666), .ZN(n13458) );
  XNOR2_X1 U7651 ( .A(n14628), .B(n10436), .ZN(n10522) );
  INV_X1 U7652 ( .A(n14398), .ZN(n14261) );
  OR2_X1 U7653 ( .A1(n14562), .A2(n14397), .ZN(n8504) );
  AND2_X1 U7654 ( .A1(n9451), .A2(n15696), .ZN(n9506) );
  NAND2_X2 U7655 ( .A1(n9514), .A2(n7218), .ZN(n9812) );
  INV_X2 U7656 ( .A(n9555), .ZN(n9940) );
  NAND2_X1 U7657 ( .A1(n7227), .A2(n7965), .ZN(n15557) );
  OAI21_X1 U7658 ( .B1(n9743), .B2(n15843), .A(n7108), .ZN(n9570) );
  NAND2_X1 U7659 ( .A1(n9743), .A2(n15098), .ZN(n7108) );
  NAND2_X1 U7660 ( .A1(n9569), .A2(n7921), .ZN(n7920) );
  INV_X1 U7661 ( .A(n9570), .ZN(n7921) );
  NAND2_X1 U7662 ( .A1(n14131), .A2(n14130), .ZN(n7295) );
  INV_X1 U7663 ( .A(n14149), .ZN(n7529) );
  AOI21_X1 U7664 ( .B1(n7400), .B2(n13412), .A(n6582), .ZN(n7399) );
  MUX2_X1 U7665 ( .A(n14406), .B(n14809), .S(n14263), .Z(n14216) );
  AOI22_X1 U7666 ( .A1(n7930), .A2(n7926), .B1(n9825), .B2(n7925), .ZN(n7924)
         );
  INV_X1 U7667 ( .A(n7928), .ZN(n7926) );
  NOR2_X1 U7668 ( .A1(n9287), .A2(n7851), .ZN(n7850) );
  INV_X1 U7669 ( .A(n9274), .ZN(n7851) );
  NAND2_X1 U7670 ( .A1(n16036), .A2(n16047), .ZN(n7538) );
  OAI21_X1 U7671 ( .B1(n14240), .B2(n7527), .A(n7307), .ZN(n14246) );
  NOR2_X1 U7672 ( .A1(n14245), .A2(n7308), .ZN(n7307) );
  AOI21_X1 U7673 ( .B1(n7681), .B2(n7680), .A(n14577), .ZN(n7679) );
  INV_X1 U7674 ( .A(n7683), .ZN(n7680) );
  NAND2_X1 U7675 ( .A1(n9971), .A2(n9972), .ZN(n7871) );
  INV_X1 U7676 ( .A(n7878), .ZN(n7877) );
  OAI21_X1 U7677 ( .B1(n7978), .B2(n7879), .A(n8309), .ZN(n7878) );
  NAND2_X1 U7678 ( .A1(n8254), .A2(n11056), .ZN(n8269) );
  NAND2_X1 U7679 ( .A1(n8214), .A2(n10683), .ZN(n8229) );
  OR2_X1 U7680 ( .A1(n12970), .A2(n13257), .ZN(n12972) );
  NOR2_X1 U7681 ( .A1(n12938), .A2(n7834), .ZN(n7833) );
  INV_X1 U7682 ( .A(n7837), .ZN(n7834) );
  AND2_X1 U7683 ( .A1(n7080), .A2(n7079), .ZN(n13479) );
  NAND2_X1 U7684 ( .A1(n13296), .A2(n13297), .ZN(n7079) );
  NAND2_X1 U7685 ( .A1(n13299), .A2(n6636), .ZN(n7148) );
  XNOR2_X1 U7686 ( .A(n10662), .B(P3_REG1_REG_4__SCAN_IN), .ZN(n11271) );
  NAND3_X1 U7687 ( .A1(n6910), .A2(n6908), .A3(n6659), .ZN(n8819) );
  NAND2_X1 U7688 ( .A1(n6909), .A2(n7718), .ZN(n6908) );
  INV_X1 U7689 ( .A(n11697), .ZN(n7732) );
  NAND2_X1 U7690 ( .A1(n7656), .A2(n7655), .ZN(n8764) );
  AOI21_X1 U7691 ( .B1(n8756), .B2(n7658), .A(n8758), .ZN(n7655) );
  NOR2_X1 U7692 ( .A1(n6905), .A2(n6902), .ZN(n8823) );
  NOR2_X1 U7693 ( .A1(n6904), .A2(n6903), .ZN(n6902) );
  INV_X1 U7694 ( .A(P3_REG1_REG_12__SCAN_IN), .ZN(n6903) );
  NAND2_X1 U7695 ( .A1(n13664), .A2(n9317), .ZN(n9319) );
  NAND2_X1 U7696 ( .A1(n13453), .A2(n13676), .ZN(n6946) );
  NAND2_X1 U7697 ( .A1(n7260), .A2(n7259), .ZN(n13338) );
  INV_X1 U7698 ( .A(n16036), .ZN(n7259) );
  NAND2_X1 U7699 ( .A1(n7129), .A2(n7128), .ZN(n13311) );
  OR2_X1 U7700 ( .A1(n13922), .A2(n13761), .ZN(n13431) );
  INV_X1 U7701 ( .A(n7602), .ZN(n7601) );
  OAI21_X1 U7702 ( .B1(n9032), .B2(n7603), .A(n9056), .ZN(n7602) );
  NAND2_X1 U7703 ( .A1(n10699), .A2(P2_DATAO_REG_5__SCAN_IN), .ZN(n8996) );
  NAND2_X1 U7704 ( .A1(n10705), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n8955) );
  INV_X1 U7705 ( .A(n7266), .ZN(n6973) );
  OAI21_X1 U7706 ( .B1(n7750), .B2(n7751), .A(n10494), .ZN(n7266) );
  NOR2_X1 U7707 ( .A1(n14744), .A2(n14519), .ZN(n7904) );
  NOR2_X1 U7708 ( .A1(n6643), .A2(n7360), .ZN(n7359) );
  NOR2_X1 U7709 ( .A1(n14560), .A2(n7361), .ZN(n7360) );
  INV_X1 U7710 ( .A(n7980), .ZN(n7629) );
  NOR2_X1 U7711 ( .A1(n14626), .A2(n7631), .ZN(n7630) );
  INV_X1 U7712 ( .A(n8402), .ZN(n7631) );
  NAND2_X1 U7713 ( .A1(n11744), .A2(n14148), .ZN(n8598) );
  INV_X1 U7714 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n7992) );
  OR2_X1 U7715 ( .A1(n10123), .A2(n10342), .ZN(n10125) );
  OAI21_X1 U7716 ( .B1(n10248), .B2(n7962), .A(n10264), .ZN(n7961) );
  OAI21_X1 U7717 ( .B1(n14990), .B2(n14988), .A(n10265), .ZN(n10263) );
  AND2_X1 U7718 ( .A1(n10172), .A2(n10171), .ZN(n12066) );
  NAND2_X1 U7719 ( .A1(n6737), .A2(n7209), .ZN(n7084) );
  INV_X1 U7720 ( .A(n12097), .ZN(n7209) );
  OR2_X1 U7721 ( .A1(n15553), .A2(n14927), .ZN(n10024) );
  OR2_X1 U7722 ( .A1(n9883), .A2(n10935), .ZN(n9870) );
  OAI21_X1 U7723 ( .B1(n15467), .B2(n7071), .A(n13007), .ZN(n7070) );
  AND2_X1 U7724 ( .A1(n13004), .A2(n13003), .ZN(n7096) );
  OR2_X1 U7725 ( .A1(n15633), .A2(n15501), .ZN(n13003) );
  INV_X1 U7726 ( .A(n7795), .ZN(n7794) );
  OAI21_X1 U7727 ( .B1(n7175), .B2(n7796), .A(n15532), .ZN(n7795) );
  INV_X1 U7728 ( .A(n7884), .ZN(n7883) );
  AND2_X1 U7729 ( .A1(n7881), .A2(n8438), .ZN(n7880) );
  NAND2_X1 U7730 ( .A1(n7884), .A2(n7882), .ZN(n7881) );
  NOR2_X1 U7731 ( .A1(n8382), .A2(SI_18_), .ZN(n8407) );
  NAND2_X1 U7732 ( .A1(n8387), .A2(n11461), .ZN(n8411) );
  OAI21_X1 U7733 ( .B1(SI_21_), .B2(n8403), .A(n8434), .ZN(n8416) );
  AND2_X1 U7734 ( .A1(n7877), .A2(n7366), .ZN(n7365) );
  NAND2_X1 U7735 ( .A1(n7367), .A2(n8253), .ZN(n7366) );
  NAND2_X1 U7736 ( .A1(n8211), .A2(n7065), .ZN(n6809) );
  AOI21_X1 U7737 ( .B1(n8097), .B2(n7265), .A(n6672), .ZN(n7264) );
  INV_X1 U7738 ( .A(n8095), .ZN(n7265) );
  INV_X1 U7739 ( .A(n8096), .ZN(n7057) );
  NAND2_X1 U7740 ( .A1(n10625), .A2(n10624), .ZN(n6844) );
  INV_X1 U7741 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n6845) );
  NAND2_X1 U7742 ( .A1(n7499), .A2(P3_ADDR_REG_4__SCAN_IN), .ZN(n10675) );
  NAND2_X1 U7743 ( .A1(n7500), .A2(n10646), .ZN(n7499) );
  NOR2_X1 U7744 ( .A1(n13152), .A2(n7836), .ZN(n7831) );
  XNOR2_X1 U7745 ( .A(n16056), .B(n6554), .ZN(n6776) );
  OAI21_X1 U7746 ( .B1(n6598), .B2(n7471), .A(n7468), .ZN(n7467) );
  NAND2_X1 U7747 ( .A1(n6598), .A2(n7469), .ZN(n7468) );
  OR2_X1 U7748 ( .A1(n7473), .A2(n7471), .ZN(n7469) );
  AND2_X1 U7749 ( .A1(n12282), .A2(n6767), .ZN(n6766) );
  NAND2_X1 U7750 ( .A1(n12249), .A2(n12310), .ZN(n6767) );
  AND2_X1 U7751 ( .A1(n8816), .A2(n11270), .ZN(n7704) );
  OR2_X1 U7752 ( .A1(n8815), .A2(n7696), .ZN(n8816) );
  NOR2_X1 U7753 ( .A1(n8820), .A2(n12601), .ZN(n8821) );
  NAND2_X1 U7754 ( .A1(n13511), .A2(n8773), .ZN(n6976) );
  AOI21_X1 U7755 ( .B1(n8889), .B2(n13582), .A(n13576), .ZN(n13597) );
  AND2_X1 U7756 ( .A1(n16021), .A2(n13332), .ZN(n7439) );
  NOR2_X1 U7757 ( .A1(n13300), .A2(n13817), .ZN(n10580) );
  OAI21_X1 U7758 ( .B1(n13719), .B2(n9256), .A(n9255), .ZN(n13703) );
  INV_X1 U7759 ( .A(n13440), .ZN(n13312) );
  NAND2_X1 U7760 ( .A1(n7860), .A2(n13747), .ZN(n13728) );
  AND2_X1 U7761 ( .A1(n9236), .A2(n9223), .ZN(n7860) );
  NOR2_X1 U7762 ( .A1(n7563), .A2(n7561), .ZN(n7560) );
  INV_X1 U7763 ( .A(n13359), .ZN(n7561) );
  OR2_X1 U7764 ( .A1(n13145), .A2(n12979), .ZN(n13462) );
  INV_X1 U7765 ( .A(n13775), .ZN(n13748) );
  NOR2_X1 U7766 ( .A1(n13758), .A2(n7032), .ZN(n7031) );
  INV_X1 U7767 ( .A(n9192), .ZN(n7032) );
  OR2_X1 U7768 ( .A1(n13868), .A2(n13791), .ZN(n13755) );
  NAND2_X1 U7769 ( .A1(n13796), .A2(n13415), .ZN(n13784) );
  INV_X1 U7770 ( .A(n7546), .ZN(n7545) );
  OAI21_X1 U7771 ( .B1(n13325), .B2(n13405), .A(n7547), .ZN(n7546) );
  AOI21_X1 U7772 ( .B1(n7545), .B2(n13405), .A(n7544), .ZN(n7543) );
  INV_X1 U7773 ( .A(n13414), .ZN(n7544) );
  AND2_X1 U7774 ( .A1(n7194), .A2(n13408), .ZN(n7838) );
  INV_X1 U7775 ( .A(n6569), .ZN(n9198) );
  INV_X1 U7776 ( .A(n13323), .ZN(n9409) );
  INV_X1 U7777 ( .A(n9353), .ZN(n13294) );
  AND2_X1 U7778 ( .A1(n13468), .A2(n11440), .ZN(n16049) );
  NAND2_X1 U7779 ( .A1(n10085), .A2(n13308), .ZN(n16044) );
  NOR2_X1 U7780 ( .A1(n9407), .A2(n7556), .ZN(n7555) );
  AOI21_X1 U7781 ( .B1(n13384), .B2(n13387), .A(n7554), .ZN(n7553) );
  INV_X1 U7782 ( .A(n13388), .ZN(n7554) );
  NAND2_X1 U7783 ( .A1(n7249), .A2(n13379), .ZN(n12110) );
  NAND2_X2 U7784 ( .A1(n8912), .A2(n7218), .ZN(n9353) );
  OR2_X1 U7785 ( .A1(n13450), .A2(n11440), .ZN(n13817) );
  NAND2_X1 U7786 ( .A1(n11708), .A2(n11431), .ZN(n16055) );
  INV_X1 U7787 ( .A(P3_IR_REG_9__SCAN_IN), .ZN(n8690) );
  AOI21_X1 U7788 ( .B1(n9320), .B2(n7613), .A(n6606), .ZN(n7612) );
  XNOR2_X1 U7789 ( .A(n9289), .B(P1_DATAO_REG_24__SCAN_IN), .ZN(n9288) );
  NAND2_X1 U7790 ( .A1(n6945), .A2(n9213), .ZN(n9239) );
  NAND2_X1 U7791 ( .A1(n9212), .A2(n9211), .ZN(n6945) );
  AND2_X1 U7792 ( .A1(n6923), .A2(n9184), .ZN(n6922) );
  OR2_X1 U7793 ( .A1(n7589), .A2(n9181), .ZN(n6923) );
  NAND2_X1 U7794 ( .A1(n10716), .A2(P1_DATAO_REG_8__SCAN_IN), .ZN(n9043) );
  NAND2_X1 U7795 ( .A1(n10710), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n8958) );
  AOI21_X1 U7796 ( .B1(n7756), .B2(n7758), .A(n6686), .ZN(n7755) );
  AOI21_X1 U7797 ( .B1(n12428), .B2(n7774), .A(n7773), .ZN(n7772) );
  INV_X1 U7798 ( .A(n10470), .ZN(n7773) );
  INV_X1 U7799 ( .A(n10464), .ZN(n7774) );
  INV_X1 U7800 ( .A(n12428), .ZN(n7775) );
  NAND2_X1 U7801 ( .A1(n10436), .A2(n14110), .ZN(n10429) );
  XNOR2_X1 U7802 ( .A(n14562), .B(n10436), .ZN(n10540) );
  NAND2_X1 U7803 ( .A1(n14009), .A2(n10523), .ZN(n10527) );
  OAI21_X1 U7804 ( .B1(n6800), .B2(n14258), .A(n14268), .ZN(n6797) );
  AOI21_X1 U7805 ( .B1(n14277), .B2(n14278), .A(n14279), .ZN(n14268) );
  AND2_X1 U7806 ( .A1(n14259), .A2(n14260), .ZN(n6800) );
  INV_X1 U7807 ( .A(n8553), .ZN(n8648) );
  INV_X1 U7808 ( .A(n14472), .ZN(n6889) );
  OR2_X1 U7809 ( .A1(n11176), .A2(n11175), .ZN(n11213) );
  OR2_X1 U7810 ( .A1(n11237), .A2(n11236), .ZN(n11234) );
  NAND2_X1 U7811 ( .A1(n8517), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n8551) );
  INV_X1 U7812 ( .A(n8519), .ZN(n8517) );
  XNOR2_X1 U7813 ( .A(n14549), .B(n14396), .ZN(n14545) );
  NAND2_X1 U7814 ( .A1(n14580), .A2(n8492), .ZN(n14559) );
  NAND2_X1 U7815 ( .A1(n7362), .A2(n8633), .ZN(n14605) );
  OR2_X1 U7816 ( .A1(n14231), .A2(n14076), .ZN(n8629) );
  NAND2_X1 U7817 ( .A1(n8628), .A2(n8627), .ZN(n7672) );
  NAND2_X1 U7818 ( .A1(n7020), .A2(n6657), .ZN(n12754) );
  NAND2_X1 U7819 ( .A1(n8609), .A2(n6644), .ZN(n7020) );
  OR2_X1 U7820 ( .A1(n14829), .A2(n14410), .ZN(n7638) );
  INV_X1 U7821 ( .A(n8227), .ZN(n7637) );
  NAND2_X1 U7822 ( .A1(n7014), .A2(n7012), .ZN(n6826) );
  AND2_X1 U7823 ( .A1(n7013), .A2(n12232), .ZN(n7012) );
  NOR2_X1 U7824 ( .A1(n14421), .A2(n14110), .ZN(n11771) );
  INV_X1 U7825 ( .A(n14110), .ZN(n14108) );
  OR2_X1 U7826 ( .A1(n10554), .A2(n8681), .ZN(n10398) );
  NAND2_X1 U7827 ( .A1(n13128), .A2(n13127), .ZN(n14318) );
  INV_X2 U7828 ( .A(n8099), .ZN(n13126) );
  INV_X4 U7829 ( .A(n8420), .ZN(n13125) );
  NAND2_X1 U7830 ( .A1(n8688), .A2(n15978), .ZN(n11633) );
  XNOR2_X1 U7831 ( .A(n7160), .B(P2_IR_REG_30__SCAN_IN), .ZN(n8008) );
  NAND2_X1 U7832 ( .A1(n7310), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7160) );
  OR2_X1 U7833 ( .A1(n9826), .A2(n8471), .ZN(n8455) );
  OR2_X1 U7834 ( .A1(n8291), .A2(P2_IR_REG_10__SCAN_IN), .ZN(n8235) );
  NAND2_X1 U7835 ( .A1(n6880), .A2(n15696), .ZN(n9486) );
  NAND2_X1 U7836 ( .A1(n9859), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n9883) );
  INV_X1 U7837 ( .A(n9881), .ZN(n9859) );
  OR2_X1 U7838 ( .A1(n14959), .A2(n14960), .ZN(n14957) );
  NAND2_X1 U7839 ( .A1(n7028), .A2(n6608), .ZN(n7027) );
  INV_X1 U7840 ( .A(n14942), .ZN(n7028) );
  AOI21_X1 U7841 ( .B1(n14960), .B2(n10303), .A(n7957), .ZN(n7956) );
  INV_X1 U7842 ( .A(n15042), .ZN(n7957) );
  AND2_X1 U7843 ( .A1(n15705), .A2(n10011), .ZN(n10719) );
  BUF_X1 U7844 ( .A(n9486), .Z(n9960) );
  NAND2_X1 U7845 ( .A1(n6866), .A2(n6865), .ZN(n11110) );
  INV_X1 U7846 ( .A(n11113), .ZN(n6865) );
  INV_X1 U7847 ( .A(n11112), .ZN(n6866) );
  AOI21_X1 U7848 ( .B1(n7346), .B2(n13054), .A(n13065), .ZN(n7345) );
  NAND2_X1 U7849 ( .A1(n9868), .A2(n9867), .ZN(n15559) );
  NAND2_X1 U7850 ( .A1(n14911), .A2(n10006), .ZN(n9868) );
  OR2_X1 U7851 ( .A1(n15290), .A2(n13049), .ZN(n13050) );
  NAND2_X1 U7852 ( .A1(n15329), .A2(n7072), .ZN(n15308) );
  NOR2_X1 U7853 ( .A1(n15311), .A2(n7073), .ZN(n7072) );
  INV_X1 U7854 ( .A(n13020), .ZN(n7073) );
  NAND2_X1 U7855 ( .A1(n15347), .A2(n7797), .ZN(n15329) );
  NOR2_X1 U7856 ( .A1(n15326), .A2(n7798), .ZN(n7797) );
  INV_X1 U7857 ( .A(n13018), .ZN(n7798) );
  OR2_X1 U7858 ( .A1(n15597), .A2(n15045), .ZN(n13041) );
  NAND2_X1 U7859 ( .A1(n7226), .A2(n6633), .ZN(n13011) );
  NAND2_X1 U7860 ( .A1(n15454), .A2(n13036), .ZN(n15430) );
  OAI21_X1 U7861 ( .B1(n12196), .B2(n7335), .A(n7334), .ZN(n7333) );
  NAND2_X1 U7862 ( .A1(n6571), .A2(n7206), .ZN(n7335) );
  AOI21_X1 U7863 ( .B1(n7336), .B2(n7206), .A(n12202), .ZN(n7334) );
  INV_X1 U7864 ( .A(n15516), .ZN(n15500) );
  NAND2_X1 U7865 ( .A1(n7132), .A2(n15250), .ZN(n11829) );
  INV_X1 U7866 ( .A(n15258), .ZN(n15541) );
  OR2_X1 U7867 ( .A1(n12183), .A2(n9812), .ZN(n9814) );
  INV_X1 U7868 ( .A(n15870), .ZN(n15844) );
  AND2_X1 U7869 ( .A1(n15436), .A2(n15620), .ZN(n15874) );
  NOR2_X1 U7870 ( .A1(P1_IR_REG_18__SCAN_IN), .A2(P1_IR_REG_21__SCAN_IN), .ZN(
        n9439) );
  INV_X1 U7871 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n9442) );
  AND2_X1 U7872 ( .A1(n8530), .A2(n8514), .ZN(n14915) );
  INV_X2 U7873 ( .A(n10695), .ZN(n9991) );
  NAND2_X1 U7874 ( .A1(n7095), .A2(n8414), .ZN(n8406) );
  INV_X1 U7875 ( .A(n8390), .ZN(n7095) );
  NAND2_X1 U7876 ( .A1(n9334), .A2(n9333), .ZN(n13666) );
  NAND2_X1 U7877 ( .A1(n15981), .A2(n10396), .ZN(n14736) );
  INV_X1 U7878 ( .A(n11483), .ZN(n11795) );
  NAND2_X1 U7879 ( .A1(n9847), .A2(n9846), .ZN(n15341) );
  INV_X1 U7880 ( .A(n15363), .ZN(n15045) );
  NAND2_X1 U7881 ( .A1(n9858), .A2(n9857), .ZN(n15306) );
  NAND2_X1 U7882 ( .A1(n9843), .A2(n9842), .ZN(n15362) );
  NAND2_X1 U7883 ( .A1(n7227), .A2(n6635), .ZN(n7062) );
  NAND2_X1 U7884 ( .A1(n7064), .A2(n13070), .ZN(n7063) );
  AND2_X1 U7885 ( .A1(n7173), .A2(n6695), .ZN(n15561) );
  OAI21_X1 U7886 ( .B1(n12333), .B2(n6609), .A(n7513), .ZN(n12843) );
  NAND2_X1 U7887 ( .A1(n11802), .A2(n9743), .ZN(n9504) );
  NAND2_X1 U7888 ( .A1(n14421), .A2(n7297), .ZN(n7296) );
  INV_X1 U7889 ( .A(n9542), .ZN(n6742) );
  NOR2_X1 U7890 ( .A1(n9635), .A2(n7219), .ZN(n9541) );
  AND2_X1 U7891 ( .A1(n7923), .A2(n9570), .ZN(n7922) );
  OR2_X1 U7892 ( .A1(n7917), .A2(n7207), .ZN(n9589) );
  OAI21_X1 U7893 ( .B1(n9605), .B2(n6577), .A(n7089), .ZN(n9622) );
  AND2_X1 U7894 ( .A1(n7912), .A2(n7090), .ZN(n7089) );
  INV_X1 U7895 ( .A(n9621), .ZN(n7090) );
  NAND2_X1 U7896 ( .A1(n7293), .A2(n7292), .ZN(n14142) );
  OR2_X1 U7897 ( .A1(n7531), .A2(n14138), .ZN(n7292) );
  INV_X1 U7898 ( .A(n14137), .ZN(n7531) );
  NAND2_X1 U7899 ( .A1(n14142), .A2(n14143), .ZN(n14141) );
  AOI21_X1 U7900 ( .B1(n7318), .B2(n7317), .A(n7315), .ZN(n7314) );
  INV_X1 U7901 ( .A(n14152), .ZN(n7315) );
  NOR2_X1 U7902 ( .A1(n7317), .A2(n14153), .ZN(n7313) );
  AOI22_X1 U7903 ( .A1(n7314), .A2(n7316), .B1(n7313), .B2(n7530), .ZN(n7311)
         );
  INV_X1 U7904 ( .A(n7318), .ZN(n7316) );
  NOR2_X1 U7905 ( .A1(n7314), .A2(n7313), .ZN(n7312) );
  AND2_X1 U7906 ( .A1(n9675), .A2(n7916), .ZN(n7915) );
  NAND2_X1 U7907 ( .A1(n9673), .A2(n9676), .ZN(n7914) );
  AOI21_X1 U7908 ( .B1(n6590), .B2(n13415), .A(n13416), .ZN(n7400) );
  INV_X1 U7909 ( .A(n13402), .ZN(n7385) );
  INV_X1 U7910 ( .A(n13399), .ZN(n7389) );
  MUX2_X1 U7911 ( .A(n14177), .B(n14176), .S(n14263), .Z(n14207) );
  AOI21_X1 U7912 ( .B1(n7399), .B2(n7397), .A(n13783), .ZN(n7396) );
  INV_X1 U7913 ( .A(n7400), .ZN(n7397) );
  NAND2_X1 U7914 ( .A1(n7306), .A2(n14170), .ZN(n7305) );
  NAND2_X1 U7915 ( .A1(n14168), .A2(n7533), .ZN(n7532) );
  AND2_X1 U7916 ( .A1(n14175), .A2(n7302), .ZN(n7301) );
  NAND2_X1 U7917 ( .A1(n7303), .A2(n14172), .ZN(n7302) );
  INV_X1 U7918 ( .A(n14170), .ZN(n7303) );
  INV_X1 U7919 ( .A(n14219), .ZN(n7142) );
  AOI21_X1 U7920 ( .B1(n7392), .B2(n7394), .A(n6592), .ZN(n7391) );
  NOR2_X1 U7921 ( .A1(n7930), .A2(n9825), .ZN(n7927) );
  NOR2_X1 U7922 ( .A1(n7931), .A2(n9823), .ZN(n7929) );
  MUX2_X1 U7923 ( .A(n13450), .B(n13449), .S(n13676), .Z(n13451) );
  INV_X1 U7924 ( .A(n9836), .ZN(n7107) );
  NAND2_X1 U7925 ( .A1(n7873), .A2(n7872), .ZN(n9972) );
  NAND2_X1 U7926 ( .A1(n10046), .A2(n9956), .ZN(n7872) );
  OR2_X1 U7927 ( .A1(n13076), .A2(n9956), .ZN(n7873) );
  INV_X1 U7928 ( .A(n12257), .ZN(n7481) );
  OR2_X1 U7929 ( .A1(n13460), .A2(n13461), .ZN(n7232) );
  AND2_X1 U7930 ( .A1(n6560), .A2(n8800), .ZN(n7411) );
  INV_X1 U7931 ( .A(n8887), .ZN(n7423) );
  NAND2_X1 U7932 ( .A1(n13677), .A2(n9286), .ZN(n7010) );
  INV_X1 U7933 ( .A(n13028), .ZN(n6885) );
  INV_X1 U7934 ( .A(n8508), .ZN(n7893) );
  INV_X1 U7935 ( .A(n7365), .ZN(n6788) );
  NAND2_X1 U7936 ( .A1(n8317), .A2(n11211), .ZN(n8330) );
  AND2_X1 U7937 ( .A1(n8086), .A2(n8085), .ZN(n8087) );
  INV_X1 U7938 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n10810) );
  INV_X1 U7939 ( .A(P3_REG3_REG_8__SCAN_IN), .ZN(n7326) );
  INV_X1 U7940 ( .A(P3_REG3_REG_7__SCAN_IN), .ZN(n8987) );
  INV_X1 U7941 ( .A(n9011), .ZN(n8988) );
  INV_X1 U7942 ( .A(n13482), .ZN(n7477) );
  INV_X1 U7943 ( .A(n13477), .ZN(n7597) );
  AND2_X1 U7944 ( .A1(n13469), .A2(n7596), .ZN(n7595) );
  NOR2_X1 U7945 ( .A1(n13330), .A2(n7330), .ZN(n7596) );
  OR2_X1 U7946 ( .A1(n6565), .A2(n7172), .ZN(n8911) );
  OR2_X1 U7947 ( .A1(n8962), .A2(n6619), .ZN(n7644) );
  INV_X1 U7948 ( .A(n11396), .ZN(n7721) );
  AOI21_X1 U7949 ( .B1(n11692), .B2(n7419), .A(n7418), .ZN(n7417) );
  INV_X1 U7950 ( .A(n12055), .ZN(n7418) );
  INV_X1 U7951 ( .A(n11693), .ZN(n7419) );
  INV_X1 U7952 ( .A(n8886), .ZN(n7714) );
  NOR2_X1 U7953 ( .A1(n7706), .A2(n12711), .ZN(n7705) );
  INV_X1 U7954 ( .A(n13564), .ZN(n7706) );
  NAND2_X1 U7955 ( .A1(n7716), .A2(n8886), .ZN(n7715) );
  NAND2_X1 U7956 ( .A1(n7640), .A2(P3_REG2_REG_16__SCAN_IN), .ZN(n7639) );
  NOR2_X1 U7957 ( .A1(n13836), .A2(n13684), .ZN(n13456) );
  NOR2_X1 U7958 ( .A1(n7010), .A2(n7005), .ZN(n7004) );
  OR2_X1 U7959 ( .A1(n13704), .A2(n7006), .ZN(n7005) );
  NOR2_X1 U7960 ( .A1(n7008), .A2(n7007), .ZN(n7006) );
  INV_X1 U7961 ( .A(n9256), .ZN(n7008) );
  INV_X1 U7962 ( .A(n7850), .ZN(n7847) );
  INV_X1 U7963 ( .A(n13677), .ZN(n13679) );
  NAND2_X1 U7964 ( .A1(n9275), .A2(n7850), .ZN(n7849) );
  NOR2_X1 U7965 ( .A1(n9279), .A2(P3_REG3_REG_24__SCAN_IN), .ZN(n9295) );
  NOR2_X1 U7966 ( .A1(n9162), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n7324) );
  OR2_X1 U7967 ( .A1(n9065), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n9092) );
  NAND2_X1 U7968 ( .A1(n7564), .A2(n13375), .ZN(n7563) );
  NAND2_X1 U7969 ( .A1(n13370), .A2(n7565), .ZN(n7564) );
  AND2_X1 U7970 ( .A1(n13313), .A2(n13359), .ZN(n7562) );
  NAND2_X1 U7971 ( .A1(n10100), .A2(n13300), .ZN(n13472) );
  OR2_X1 U7972 ( .A1(n10100), .A2(n13300), .ZN(n13475) );
  OR2_X1 U7973 ( .A1(n12859), .A2(n13502), .ZN(n13391) );
  NAND2_X1 U7974 ( .A1(n16027), .A2(n16026), .ZN(n16029) );
  AND2_X1 U7975 ( .A1(n8720), .A2(n8719), .ZN(n8792) );
  NAND2_X1 U7976 ( .A1(n9277), .A2(n9276), .ZN(n9289) );
  INV_X1 U7977 ( .A(n9107), .ZN(n6938) );
  INV_X1 U7978 ( .A(n6928), .ZN(n6927) );
  OAI21_X1 U7979 ( .B1(n6930), .B2(n6929), .A(n7601), .ZN(n6928) );
  INV_X1 U7980 ( .A(n9029), .ZN(n6929) );
  INV_X1 U7981 ( .A(n9043), .ZN(n7603) );
  AND2_X1 U7982 ( .A1(n6931), .A2(n8998), .ZN(n6930) );
  INV_X1 U7983 ( .A(n9001), .ZN(n6931) );
  NOR2_X1 U7984 ( .A1(n14074), .A2(n7766), .ZN(n7765) );
  INV_X1 U7985 ( .A(n10509), .ZN(n7766) );
  NOR2_X1 U7986 ( .A1(n8372), .A2(n8371), .ZN(n7171) );
  AND2_X1 U7987 ( .A1(n7763), .A2(n6624), .ZN(n6966) );
  NOR2_X1 U7988 ( .A1(n10492), .A2(n7752), .ZN(n7751) );
  INV_X1 U7989 ( .A(n10484), .ZN(n7752) );
  AND2_X1 U7990 ( .A1(n7267), .A2(n10486), .ZN(n7750) );
  INV_X1 U7991 ( .A(n13976), .ZN(n7267) );
  INV_X1 U7992 ( .A(n14904), .ZN(n8009) );
  INV_X1 U7993 ( .A(n7359), .ZN(n7357) );
  NAND2_X1 U7994 ( .A1(n7041), .A2(n6585), .ZN(n7358) );
  NAND2_X1 U7995 ( .A1(n14605), .A2(n7679), .ZN(n7041) );
  INV_X1 U7996 ( .A(n7685), .ZN(n7684) );
  OAI21_X1 U7997 ( .B1(n14609), .B2(n7686), .A(n8636), .ZN(n7685) );
  NAND2_X1 U7998 ( .A1(n14657), .A2(n7077), .ZN(n7670) );
  AND2_X1 U7999 ( .A1(n8625), .A2(n6573), .ZN(n7077) );
  NAND2_X1 U8000 ( .A1(n8324), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n8336) );
  NOR2_X1 U8001 ( .A1(n8260), .A2(n12925), .ZN(n7170) );
  NAND2_X1 U8002 ( .A1(n6655), .A2(n7638), .ZN(n7636) );
  INV_X1 U8003 ( .A(n8602), .ZN(n7677) );
  NOR2_X1 U8004 ( .A1(n8596), .A2(n8602), .ZN(n7675) );
  INV_X1 U8005 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n9243) );
  NAND2_X1 U8006 ( .A1(n8051), .A2(n8050), .ZN(n8067) );
  INV_X1 U8007 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n8050) );
  NAND2_X1 U8008 ( .A1(n10118), .A2(n10340), .ZN(n10135) );
  INV_X1 U8009 ( .A(n9678), .ZN(n6828) );
  NOR2_X1 U8010 ( .A1(n9828), .A2(n15044), .ZN(n6829) );
  NOR2_X1 U8011 ( .A1(n9975), .A2(n9976), .ZN(n9983) );
  INV_X1 U8012 ( .A(n9989), .ZN(n9986) );
  NAND2_X1 U8013 ( .A1(n15565), .A2(n7460), .ZN(n7459) );
  INV_X1 U8014 ( .A(n7461), .ZN(n7460) );
  INV_X1 U8015 ( .A(n15086), .ZN(n13055) );
  NAND2_X1 U8016 ( .A1(n13040), .A2(n10026), .ZN(n13039) );
  AND2_X1 U8017 ( .A1(n15485), .A2(n15482), .ZN(n13002) );
  NOR2_X1 U8018 ( .A1(n7454), .A2(n12902), .ZN(n7453) );
  INV_X1 U8019 ( .A(n7455), .ZN(n7454) );
  INV_X1 U8020 ( .A(n9591), .ZN(n9432) );
  INV_X1 U8021 ( .A(n15095), .ZN(n12201) );
  NAND2_X1 U8022 ( .A1(n12029), .A2(n15098), .ZN(n12032) );
  OR2_X1 U8023 ( .A1(n12028), .A2(n15795), .ZN(n12029) );
  NAND2_X1 U8024 ( .A1(n13058), .A2(n6814), .ZN(n15277) );
  NOR2_X1 U8025 ( .A1(n7459), .A2(n15559), .ZN(n6814) );
  XNOR2_X1 U8026 ( .A(n15586), .B(n15362), .ZN(n15351) );
  NAND2_X1 U8027 ( .A1(n15352), .A2(n15351), .ZN(n15350) );
  OR2_X1 U8028 ( .A1(n8510), .A2(n12507), .ZN(n8529) );
  AND2_X1 U8029 ( .A1(n9443), .A2(n10061), .ZN(n7054) );
  OR2_X1 U8030 ( .A1(n8476), .A2(n12984), .ZN(n8493) );
  INV_X1 U8031 ( .A(n7895), .ZN(n7894) );
  INV_X1 U8032 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n9468) );
  OR2_X1 U8033 ( .A1(n8432), .A2(n11459), .ZN(n8364) );
  AND2_X1 U8034 ( .A1(n7364), .A2(n7874), .ZN(n7363) );
  AOI21_X1 U8035 ( .B1(n7877), .B2(n7879), .A(n7875), .ZN(n7874) );
  INV_X1 U8036 ( .A(n8316), .ZN(n7875) );
  NAND2_X1 U8037 ( .A1(n8286), .A2(SI_15_), .ZN(n8314) );
  NAND2_X1 U8038 ( .A1(n7058), .A2(n8311), .ZN(n8285) );
  NAND2_X1 U8039 ( .A1(n8229), .A2(n8216), .ZN(n8230) );
  NAND2_X1 U8040 ( .A1(n7067), .A2(n8177), .ZN(n8194) );
  AND2_X1 U8042 ( .A1(n10626), .A2(n10618), .ZN(n10624) );
  OR2_X1 U8043 ( .A1(n11337), .A2(P3_ADDR_REG_7__SCAN_IN), .ZN(n11578) );
  OAI21_X1 U8044 ( .B1(n11579), .B2(n15161), .A(n11578), .ZN(n11583) );
  NAND2_X1 U8045 ( .A1(n11947), .A2(n11946), .ZN(n12007) );
  AND2_X1 U8046 ( .A1(n12971), .A2(n7856), .ZN(n7855) );
  OR2_X1 U8047 ( .A1(n7858), .A2(n7857), .ZN(n7856) );
  NAND2_X1 U8048 ( .A1(n12935), .A2(n7833), .ZN(n7832) );
  NAND2_X1 U8049 ( .A1(n8988), .A2(n6627), .ZN(n9049) );
  NOR2_X1 U8050 ( .A1(n13175), .A2(n6783), .ZN(n6782) );
  INV_X1 U8051 ( .A(n12956), .ZN(n6783) );
  INV_X1 U8052 ( .A(n7831), .ZN(n7830) );
  AND2_X1 U8053 ( .A1(n11607), .A2(n11608), .ZN(n11605) );
  INV_X1 U8054 ( .A(n11652), .ZN(n7488) );
  NOR2_X1 U8055 ( .A1(n16048), .A2(n11845), .ZN(n13339) );
  AOI21_X1 U8056 ( .B1(n7831), .B2(n7829), .A(n6678), .ZN(n7828) );
  INV_X1 U8057 ( .A(n7833), .ZN(n7829) );
  AND2_X1 U8058 ( .A1(n7828), .A2(n7492), .ZN(n7491) );
  INV_X1 U8059 ( .A(n13265), .ZN(n7492) );
  OR2_X1 U8060 ( .A1(n12935), .A2(n7830), .ZN(n7493) );
  NAND2_X1 U8061 ( .A1(n9356), .A2(n9355), .ZN(n13290) );
  INV_X1 U8062 ( .A(n9423), .ZN(n9356) );
  AOI21_X1 U8063 ( .B1(n8834), .B2(n8812), .A(n8813), .ZN(n11287) );
  NAND2_X1 U8064 ( .A1(n8838), .A2(n11300), .ZN(n11282) );
  NAND2_X1 U8065 ( .A1(n7704), .A2(P3_REG1_REG_3__SCAN_IN), .ZN(n11320) );
  NOR2_X1 U8066 ( .A1(n11271), .A2(n11317), .ZN(n7698) );
  NAND2_X1 U8067 ( .A1(n7703), .A2(n7701), .ZN(n7700) );
  INV_X1 U8068 ( .A(n11270), .ZN(n7701) );
  AND2_X1 U8069 ( .A1(n7702), .A2(n7646), .ZN(n8817) );
  NAND2_X1 U8070 ( .A1(n7647), .A2(n7646), .ZN(n11391) );
  INV_X1 U8071 ( .A(n7406), .ZN(n7408) );
  OAI21_X1 U8072 ( .B1(n11325), .B2(n7407), .A(n11261), .ZN(n7406) );
  NAND2_X1 U8073 ( .A1(n8862), .A2(n11540), .ZN(n11694) );
  AND2_X1 U8074 ( .A1(n7196), .A2(n7195), .ZN(n12052) );
  NAND2_X1 U8075 ( .A1(n6690), .A2(n7728), .ZN(n6912) );
  NAND2_X1 U8076 ( .A1(n12061), .A2(n7732), .ZN(n7722) );
  NAND2_X1 U8077 ( .A1(n12052), .A2(P3_REG2_REG_9__SCAN_IN), .ZN(n12051) );
  NAND2_X1 U8078 ( .A1(n7429), .A2(n7428), .ZN(n13536) );
  INV_X1 U8079 ( .A(n13520), .ZN(n7428) );
  INV_X1 U8080 ( .A(n13519), .ZN(n7429) );
  NOR2_X1 U8081 ( .A1(n8824), .A2(n13565), .ZN(n13533) );
  NAND2_X1 U8082 ( .A1(n13536), .A2(n8882), .ZN(n13558) );
  NOR2_X1 U8083 ( .A1(n7427), .A2(n6683), .ZN(n7426) );
  AND2_X1 U8084 ( .A1(n8882), .A2(n13520), .ZN(n7427) );
  INV_X1 U8085 ( .A(n13557), .ZN(n7430) );
  NAND2_X1 U8086 ( .A1(n7641), .A2(n13589), .ZN(n13590) );
  INV_X1 U8087 ( .A(n13597), .ZN(n7437) );
  NOR2_X1 U8088 ( .A1(n13613), .A2(n7434), .ZN(n7433) );
  XNOR2_X1 U8089 ( .A(n8899), .B(n7441), .ZN(n7440) );
  INV_X1 U8090 ( .A(n8898), .ZN(n7441) );
  OR2_X1 U8091 ( .A1(n9342), .A2(P3_REG3_REG_28__SCAN_IN), .ZN(n9423) );
  NAND2_X1 U8092 ( .A1(n9319), .A2(n9318), .ZN(n10080) );
  OR2_X1 U8093 ( .A1(n9308), .A2(P3_REG3_REG_26__SCAN_IN), .ZN(n9328) );
  NAND2_X1 U8094 ( .A1(n6570), .A2(n6647), .ZN(n7244) );
  NAND2_X1 U8095 ( .A1(n6570), .A2(n13704), .ZN(n7246) );
  NAND2_X1 U8096 ( .A1(n13435), .A2(n13436), .ZN(n9236) );
  INV_X1 U8097 ( .A(n9236), .ZN(n13731) );
  NAND2_X1 U8098 ( .A1(n9202), .A2(n9201), .ZN(n9216) );
  INV_X1 U8099 ( .A(n7324), .ZN(n9175) );
  OR2_X1 U8100 ( .A1(n9127), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n9147) );
  AOI21_X1 U8101 ( .B1(n13381), .B2(n9055), .A(n7844), .ZN(n7843) );
  NAND2_X1 U8102 ( .A1(n7567), .A2(n7566), .ZN(n11866) );
  NOR2_X1 U8103 ( .A1(n7562), .A2(n9406), .ZN(n7566) );
  NAND2_X1 U8104 ( .A1(n13359), .A2(n12098), .ZN(n7567) );
  NOR2_X1 U8105 ( .A1(n9396), .A2(n10088), .ZN(n10109) );
  OR3_X1 U8106 ( .A1(n11422), .A2(n10091), .A3(n10087), .ZN(n9396) );
  AND2_X1 U8107 ( .A1(n13311), .A2(n13676), .ZN(n13696) );
  NAND2_X1 U8108 ( .A1(n13784), .A2(n13788), .ZN(n7258) );
  NAND2_X1 U8109 ( .A1(n7258), .A2(n7257), .ZN(n13767) );
  AND3_X1 U8110 ( .A1(n9191), .A2(n9190), .A3(n9189), .ZN(n13791) );
  INV_X1 U8111 ( .A(n7035), .ZN(n7034) );
  OAI21_X1 U8112 ( .B1(n13802), .B2(n7039), .A(n13783), .ZN(n7035) );
  AND3_X1 U8113 ( .A1(n9179), .A2(n9178), .A3(n9177), .ZN(n13805) );
  AOI21_X1 U8114 ( .B1(n7543), .B2(n7541), .A(n13802), .ZN(n7540) );
  INV_X1 U8115 ( .A(n7543), .ZN(n7542) );
  INV_X1 U8116 ( .A(n7545), .ZN(n7541) );
  INV_X1 U8117 ( .A(n16044), .ZN(n16034) );
  NAND2_X1 U8118 ( .A1(n9136), .A2(n9135), .ZN(n13325) );
  INV_X1 U8119 ( .A(n16049), .ZN(n13815) );
  AOI21_X1 U8120 ( .B1(n7551), .B2(n7553), .A(n7550), .ZN(n7549) );
  NAND2_X1 U8121 ( .A1(n7249), .A2(n7247), .ZN(n7253) );
  INV_X1 U8122 ( .A(n7555), .ZN(n7551) );
  OR2_X1 U8123 ( .A1(n11422), .A2(n11595), .ZN(n13486) );
  NAND2_X1 U8124 ( .A1(n13100), .A2(n13099), .ZN(n13280) );
  NAND2_X1 U8125 ( .A1(n9352), .A2(n9351), .ZN(n13100) );
  INV_X1 U8126 ( .A(P3_IR_REG_25__SCAN_IN), .ZN(n7569) );
  AND2_X1 U8127 ( .A1(n8803), .A2(n8805), .ZN(n7862) );
  OR2_X1 U8128 ( .A1(n9289), .A2(n12580), .ZN(n9290) );
  NAND2_X1 U8129 ( .A1(n9288), .A2(n12578), .ZN(n7580) );
  INV_X1 U8130 ( .A(P3_IR_REG_24__SCAN_IN), .ZN(n8704) );
  NOR2_X1 U8131 ( .A1(P3_IR_REG_24__SCAN_IN), .A2(P3_IR_REG_31__SCAN_IN), .ZN(
        n8710) );
  INV_X1 U8132 ( .A(P3_IR_REG_19__SCAN_IN), .ZN(n8700) );
  AOI21_X1 U8133 ( .B1(n6922), .B2(n9181), .A(n9193), .ZN(n6921) );
  OR2_X1 U8134 ( .A1(n8784), .A2(P3_IR_REG_18__SCAN_IN), .ZN(n8789) );
  AOI21_X1 U8135 ( .B1(n7591), .B2(n7593), .A(n6724), .ZN(n7589) );
  NAND2_X1 U8136 ( .A1(n6934), .A2(n6932), .ZN(n9156) );
  AOI21_X1 U8137 ( .B1(n6936), .B2(n6938), .A(n6933), .ZN(n6932) );
  NAND2_X1 U8138 ( .A1(n9105), .A2(n6936), .ZN(n6934) );
  INV_X1 U8139 ( .A(n9142), .ZN(n6933) );
  XNOR2_X1 U8140 ( .A(n9139), .B(P2_DATAO_REG_13__SCAN_IN), .ZN(n9119) );
  NOR2_X1 U8141 ( .A1(n8766), .A2(P3_IR_REG_11__SCAN_IN), .ZN(n8770) );
  AND2_X1 U8142 ( .A1(n9058), .A2(n9045), .ZN(n9056) );
  NAND2_X1 U8143 ( .A1(n9030), .A2(n9029), .ZN(n9033) );
  AND2_X1 U8144 ( .A1(n9043), .A2(n9031), .ZN(n9032) );
  NAND2_X1 U8145 ( .A1(n9033), .A2(n9032), .ZN(n9044) );
  NAND2_X1 U8146 ( .A1(n8999), .A2(n6930), .ZN(n9030) );
  AOI21_X1 U8147 ( .B1(n7585), .B2(n7587), .A(n7582), .ZN(n7581) );
  INV_X1 U8148 ( .A(n8996), .ZN(n7582) );
  AND2_X1 U8149 ( .A1(n8996), .A2(n8959), .ZN(n8994) );
  AND2_X1 U8150 ( .A1(n8958), .A2(n8957), .ZN(n8971) );
  NAND2_X1 U8151 ( .A1(n6995), .A2(n6994), .ZN(n8939) );
  AND2_X1 U8152 ( .A1(n8952), .A2(n8936), .ZN(n8950) );
  NAND2_X1 U8153 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(P3_IR_REG_0__SCAN_IN), .ZN(
        n8736) );
  NAND2_X1 U8154 ( .A1(n8913), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n8934) );
  INV_X1 U8155 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n8666) );
  NAND2_X1 U8156 ( .A1(n7753), .A2(n7121), .ZN(n6959) );
  NAND2_X1 U8157 ( .A1(n11740), .A2(n7755), .ZN(n7121) );
  INV_X1 U8158 ( .A(n11979), .ZN(n7754) );
  NAND2_X1 U8159 ( .A1(n7168), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n8245) );
  INV_X1 U8160 ( .A(n8221), .ZN(n7168) );
  NAND2_X1 U8161 ( .A1(n11616), .A2(n10443), .ZN(n11740) );
  NAND2_X1 U8162 ( .A1(n8445), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n8484) );
  AND2_X1 U8163 ( .A1(n10527), .A2(n10526), .ZN(n13990) );
  INV_X1 U8164 ( .A(n11771), .ZN(n11906) );
  AND2_X1 U8165 ( .A1(n10516), .A2(n14001), .ZN(n7279) );
  NAND2_X1 U8166 ( .A1(n12890), .A2(n12891), .ZN(n12889) );
  NOR2_X1 U8167 ( .A1(n7771), .A2(n12819), .ZN(n7770) );
  INV_X1 U8168 ( .A(n7772), .ZN(n7771) );
  INV_X1 U8169 ( .A(n12819), .ZN(n7769) );
  OR2_X1 U8170 ( .A1(n12870), .A2(n12869), .ZN(n12867) );
  OR2_X1 U8171 ( .A1(n8336), .A2(n8335), .ZN(n8355) );
  INV_X1 U8172 ( .A(n6964), .ZN(n6963) );
  OAI21_X1 U8173 ( .B1(n14047), .B2(n6965), .A(n14018), .ZN(n6964) );
  INV_X1 U8174 ( .A(n10539), .ZN(n6965) );
  INV_X1 U8175 ( .A(n10545), .ZN(n6962) );
  NOR2_X1 U8176 ( .A1(n14322), .A2(n7738), .ZN(n7737) );
  NAND2_X1 U8177 ( .A1(n14329), .A2(n7517), .ZN(n7738) );
  AND2_X1 U8178 ( .A1(n14367), .A2(n7517), .ZN(n14387) );
  OR2_X1 U8179 ( .A1(n8376), .A2(n11157), .ZN(n8042) );
  OR2_X1 U8180 ( .A1(n8376), .A2(n11154), .ZN(n8026) );
  NAND2_X1 U8181 ( .A1(n6891), .A2(n6890), .ZN(n11925) );
  INV_X1 U8182 ( .A(n11731), .ZN(n6890) );
  INV_X1 U8183 ( .A(n11732), .ZN(n6891) );
  INV_X1 U8184 ( .A(n6878), .ZN(n6877) );
  OAI21_X1 U8185 ( .B1(n15939), .B2(n6879), .A(n12688), .ZN(n6878) );
  INV_X1 U8186 ( .A(n12686), .ZN(n6879) );
  AOI21_X1 U8187 ( .B1(n14536), .B2(n7695), .A(n6645), .ZN(n7694) );
  INV_X1 U8188 ( .A(n8638), .ZN(n7695) );
  OR2_X1 U8189 ( .A1(n8551), .A2(n8550), .ZN(n10402) );
  INV_X1 U8190 ( .A(n14749), .ZN(n14531) );
  NAND2_X1 U8191 ( .A1(n7620), .A2(n8527), .ZN(n14537) );
  NAND2_X1 U8192 ( .A1(n7627), .A2(n8469), .ZN(n6817) );
  NAND2_X1 U8193 ( .A1(n14637), .A2(n7630), .ZN(n6819) );
  INV_X1 U8194 ( .A(n7627), .ZN(n6818) );
  AND2_X1 U8195 ( .A1(n7687), .A2(n8634), .ZN(n7683) );
  AND2_X1 U8196 ( .A1(n14358), .A2(n14357), .ZN(n14592) );
  OR2_X1 U8197 ( .A1(n14618), .A2(n14248), .ZN(n8634) );
  NAND2_X1 U8198 ( .A1(n7688), .A2(n14609), .ZN(n14607) );
  INV_X1 U8199 ( .A(n14605), .ZN(n7688) );
  NAND2_X1 U8200 ( .A1(n8401), .A2(n7980), .ZN(n7632) );
  NAND2_X1 U8201 ( .A1(n7672), .A2(n7671), .ZN(n14645) );
  NAND2_X1 U8202 ( .A1(n7048), .A2(n7046), .ZN(n8628) );
  OR2_X1 U8203 ( .A1(n8622), .A2(n7047), .ZN(n7046) );
  NAND2_X1 U8204 ( .A1(n8619), .A2(n7049), .ZN(n7048) );
  INV_X1 U8205 ( .A(n8624), .ZN(n7047) );
  NOR2_X1 U8206 ( .A1(n8306), .A2(n7692), .ZN(n7690) );
  XNOR2_X1 U8207 ( .A(n14824), .B(n14188), .ZN(n14328) );
  NAND2_X1 U8208 ( .A1(n6824), .A2(n7015), .ZN(n8228) );
  AOI21_X1 U8209 ( .B1(n7016), .B2(n8610), .A(n6674), .ZN(n7015) );
  NAND2_X1 U8210 ( .A1(n12376), .A2(n7016), .ZN(n6824) );
  NAND2_X1 U8211 ( .A1(n8597), .A2(n12614), .ZN(n8599) );
  NAND2_X1 U8212 ( .A1(n12615), .A2(n8596), .ZN(n7673) );
  AND2_X1 U8213 ( .A1(n7055), .A2(n15983), .ZN(n12614) );
  INV_X1 U8214 ( .A(n14417), .ZN(n7055) );
  XNOR2_X1 U8215 ( .A(n14419), .B(n11713), .ZN(n11671) );
  NAND2_X1 U8216 ( .A1(n8590), .A2(n8589), .ZN(n11673) );
  NAND2_X1 U8217 ( .A1(n11676), .A2(n11713), .ZN(n11816) );
  OAI21_X2 U8218 ( .B1(n14379), .B2(n8584), .A(n14372), .ZN(n14675) );
  XNOR2_X1 U8219 ( .A(n7166), .B(n14420), .ZN(n11625) );
  XNOR2_X1 U8220 ( .A(n14107), .B(n14379), .ZN(n6958) );
  NAND2_X1 U8221 ( .A1(n10394), .A2(n10393), .ZN(n14744) );
  NAND2_X1 U8222 ( .A1(n8496), .A2(n8495), .ZN(n14562) );
  OR2_X1 U8223 ( .A1(n12143), .A2(n7140), .ZN(n8422) );
  NAND2_X1 U8224 ( .A1(n8370), .A2(n8369), .ZN(n14231) );
  INV_X1 U8225 ( .A(n11909), .ZN(n7739) );
  NAND2_X1 U8226 ( .A1(n8242), .A2(n8241), .ZN(n14829) );
  AND2_X1 U8227 ( .A1(n10420), .A2(n14846), .ZN(n16000) );
  NAND2_X1 U8228 ( .A1(n14383), .A2(n14379), .ZN(n14846) );
  NAND2_X1 U8229 ( .A1(n8023), .A2(n8005), .ZN(n8021) );
  AND2_X2 U8230 ( .A1(n7908), .A2(n6949), .ZN(n8023) );
  AND2_X1 U8231 ( .A1(n8657), .A2(n8656), .ZN(n8683) );
  OR2_X1 U8232 ( .A1(n8576), .A2(P2_IR_REG_22__SCAN_IN), .ZN(n8658) );
  AND2_X1 U8233 ( .A1(n8181), .A2(n8291), .ZN(n11221) );
  AND2_X1 U8234 ( .A1(n10179), .A2(n7942), .ZN(n7935) );
  NAND2_X1 U8235 ( .A1(n10249), .A2(n10248), .ZN(n14931) );
  INV_X1 U8236 ( .A(n11756), .ZN(n10158) );
  OR2_X1 U8237 ( .A1(n6553), .A2(n10725), .ZN(n9493) );
  AND2_X1 U8238 ( .A1(n6608), .A2(n10307), .ZN(n7029) );
  NAND2_X1 U8239 ( .A1(n9433), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n9640) );
  INV_X1 U8240 ( .A(n9624), .ZN(n9433) );
  OAI21_X1 U8241 ( .B1(n7961), .B2(n14933), .A(n7959), .ZN(n10274) );
  AOI21_X1 U8242 ( .B1(n7960), .B2(n7962), .A(n10269), .ZN(n7959) );
  AND2_X1 U8243 ( .A1(n10178), .A2(n10177), .ZN(n7941) );
  CLKBUF_X1 U8244 ( .A(n12079), .Z(n7155) );
  NAND3_X1 U8245 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .A3(P1_REG3_REG_5__SCAN_IN), .ZN(n9573) );
  NAND2_X1 U8246 ( .A1(n9431), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n9591) );
  INV_X1 U8247 ( .A(n9573), .ZN(n9431) );
  NAND2_X1 U8248 ( .A1(n10022), .A2(n7210), .ZN(n10053) );
  NOR2_X1 U8249 ( .A1(n7212), .A2(n7211), .ZN(n7210) );
  NOR2_X1 U8250 ( .A1(n10023), .A2(n15256), .ZN(n7211) );
  INV_X1 U8251 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n15122) );
  NAND2_X1 U8252 ( .A1(n11090), .A2(n6870), .ZN(n11195) );
  NOR2_X1 U8253 ( .A1(n11198), .A2(n6871), .ZN(n6870) );
  INV_X1 U8254 ( .A(n11089), .ZN(n6871) );
  NAND2_X1 U8255 ( .A1(n11559), .A2(n11558), .ZN(n11560) );
  NAND2_X1 U8256 ( .A1(n11560), .A2(n11561), .ZN(n11891) );
  OR2_X1 U8257 ( .A1(n11893), .A2(n11894), .ZN(n12166) );
  NAND2_X1 U8258 ( .A1(n9860), .A2(P1_REG3_REG_27__SCAN_IN), .ZN(n13079) );
  INV_X1 U8259 ( .A(n13088), .ZN(n7343) );
  AND2_X1 U8260 ( .A1(n9870), .A2(n9869), .ZN(n15298) );
  INV_X1 U8261 ( .A(n13058), .ZN(n15336) );
  NAND2_X1 U8262 ( .A1(n15388), .A2(n15387), .ZN(n13042) );
  NAND2_X1 U8263 ( .A1(n9435), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n9817) );
  INV_X1 U8264 ( .A(n9815), .ZN(n9435) );
  INV_X1 U8265 ( .A(n15421), .ZN(n15390) );
  NAND2_X1 U8266 ( .A1(n15403), .A2(n13040), .ZN(n15388) );
  AND2_X1 U8267 ( .A1(n13012), .A2(n13037), .ZN(n7820) );
  NAND2_X1 U8268 ( .A1(n7819), .A2(n7818), .ZN(n15403) );
  AND2_X1 U8269 ( .A1(n15404), .A2(n6638), .ZN(n7818) );
  INV_X1 U8270 ( .A(n13039), .ZN(n15404) );
  NAND2_X1 U8271 ( .A1(n13005), .A2(n7096), .ZN(n15468) );
  NAND2_X1 U8272 ( .A1(n15468), .A2(n15467), .ZN(n15466) );
  INV_X1 U8273 ( .A(n13029), .ZN(n15505) );
  AOI21_X1 U8274 ( .B1(n7811), .B2(n7812), .A(n6670), .ZN(n7809) );
  INV_X1 U8275 ( .A(n13023), .ZN(n7175) );
  NAND2_X1 U8276 ( .A1(n12566), .A2(n7175), .ZN(n13000) );
  XNOR2_X1 U8277 ( .A(n15651), .B(n15520), .ZN(n13023) );
  OR2_X1 U8278 ( .A1(n12556), .A2(n7815), .ZN(n7814) );
  INV_X1 U8279 ( .A(n12361), .ZN(n7815) );
  NAND2_X1 U8280 ( .A1(n12360), .A2(n12359), .ZN(n12362) );
  XNOR2_X1 U8281 ( .A(n15869), .B(n12201), .ZN(n12337) );
  OAI21_X1 U8282 ( .B1(n12195), .B2(n7337), .A(n12200), .ZN(n7336) );
  XNOR2_X1 U8283 ( .A(n15780), .B(n12199), .ZN(n15776) );
  NAND2_X1 U8284 ( .A1(n11960), .A2(n11806), .ZN(n12019) );
  AND2_X1 U8285 ( .A1(n10719), .A2(n11071), .ZN(n15521) );
  NAND2_X1 U8286 ( .A1(n9759), .A2(n9758), .ZN(n15622) );
  NAND2_X1 U8287 ( .A1(n9718), .A2(n9717), .ZN(n15645) );
  OAI211_X1 U8288 ( .C1(n10005), .C2(n10004), .A(n10003), .B(n10002), .ZN(
        n14895) );
  XNOR2_X1 U8289 ( .A(n9939), .B(n9938), .ZN(n13133) );
  NAND2_X1 U8290 ( .A1(n10005), .A2(n9993), .ZN(n9939) );
  AND2_X1 U8291 ( .A1(n7778), .A2(n7779), .ZN(n7349) );
  AND3_X2 U8292 ( .A1(n7779), .A2(n9465), .A3(n7777), .ZN(n9459) );
  NAND2_X1 U8293 ( .A1(n10056), .A2(n7052), .ZN(n10067) );
  AND2_X1 U8294 ( .A1(n7054), .A2(n7053), .ZN(n7052) );
  NAND2_X1 U8295 ( .A1(n10056), .A2(n7054), .ZN(n10063) );
  XNOR2_X1 U8296 ( .A(n8442), .B(n8441), .ZN(n12317) );
  NAND2_X1 U8297 ( .A1(n7886), .A2(n8346), .ZN(n8432) );
  AOI21_X1 U8298 ( .B1(n8412), .B2(n8411), .A(n8410), .ZN(n8433) );
  NAND2_X1 U8299 ( .A1(n8408), .A2(n8411), .ZN(n8430) );
  NOR2_X1 U8300 ( .A1(n8416), .A2(n8415), .ZN(n8436) );
  INV_X1 U8301 ( .A(n9476), .ZN(n9478) );
  NOR2_X1 U8302 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), .ZN(
        n9477) );
  OR2_X1 U8303 ( .A1(n9647), .A2(P1_IR_REG_9__SCAN_IN), .ZN(n9668) );
  NAND4_X1 U8304 ( .A1(n8014), .A2(n6807), .A3(P3_ADDR_REG_19__SCAN_IN), .A4(
        n6806), .ZN(n6805) );
  NAND4_X1 U8305 ( .A1(n15768), .A2(P1_ADDR_REG_19__SCAN_IN), .A3(n6804), .A4(
        P2_ADDR_REG_19__SCAN_IN), .ZN(n6803) );
  INV_X1 U8306 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n6807) );
  NAND2_X1 U8307 ( .A1(n9499), .A2(n8031), .ZN(n8048) );
  NAND2_X1 U8308 ( .A1(n10676), .A2(n10649), .ZN(n10679) );
  NAND2_X1 U8309 ( .A1(n10675), .A2(n6846), .ZN(n10648) );
  NAND2_X1 U8310 ( .A1(n11048), .A2(n11047), .ZN(n11339) );
  INV_X1 U8311 ( .A(n11576), .ZN(n6841) );
  NAND2_X1 U8312 ( .A1(n11945), .A2(n6842), .ZN(n12001) );
  NAND2_X1 U8313 ( .A1(n12329), .A2(n12328), .ZN(n12527) );
  NAND2_X1 U8314 ( .A1(n12848), .A2(n12847), .ZN(n15714) );
  OR2_X1 U8315 ( .A1(n12845), .A2(n12844), .ZN(n12848) );
  OAI21_X1 U8316 ( .B1(n15743), .B2(P2_ADDR_REG_16__SCAN_IN), .A(n15742), .ZN(
        n15751) );
  INV_X1 U8317 ( .A(n15764), .ZN(n7123) );
  AND2_X1 U8318 ( .A1(n9222), .A2(n9221), .ZN(n13761) );
  NAND2_X1 U8319 ( .A1(n9341), .A2(n9340), .ZN(n13145) );
  AND2_X1 U8320 ( .A1(n9254), .A2(n9253), .ZN(n13733) );
  NOR2_X1 U8321 ( .A1(n6602), .A2(n13264), .ZN(n7463) );
  INV_X1 U8322 ( .A(n7473), .ZN(n7466) );
  NAND2_X1 U8323 ( .A1(n7467), .A2(n7470), .ZN(n7465) );
  NAND2_X1 U8324 ( .A1(n6598), .A2(n7472), .ZN(n7470) );
  AND2_X1 U8325 ( .A1(n11653), .A2(n7487), .ZN(n11913) );
  NAND2_X1 U8326 ( .A1(n6768), .A2(n6632), .ZN(n6765) );
  NAND2_X1 U8327 ( .A1(n9186), .A2(n9185), .ZN(n13868) );
  OAI21_X1 U8328 ( .B1(n7854), .B2(n6780), .A(n6778), .ZN(n6781) );
  AOI21_X1 U8329 ( .B1(n13254), .B2(n7857), .A(n6779), .ZN(n6778) );
  INV_X1 U8330 ( .A(n13254), .ZN(n6780) );
  INV_X1 U8331 ( .A(n13256), .ZN(n6779) );
  INV_X1 U8332 ( .A(n13257), .ZN(n7109) );
  INV_X1 U8333 ( .A(n13261), .ZN(n13276) );
  OR2_X1 U8334 ( .A1(n11610), .A2(n11609), .ZN(n13273) );
  NAND2_X1 U8335 ( .A1(n13480), .A2(n10086), .ZN(n7373) );
  INV_X1 U8336 ( .A(n13761), .ZN(n13495) );
  INV_X1 U8337 ( .A(n13791), .ZN(n13496) );
  OR2_X1 U8338 ( .A1(n9126), .A2(n11658), .ZN(n8967) );
  OAI21_X1 U8339 ( .B1(n8821), .B2(n7734), .A(n7733), .ZN(n6905) );
  OR2_X1 U8340 ( .A1(n13524), .A2(n12593), .ZN(n7734) );
  NAND2_X1 U8341 ( .A1(n6975), .A2(n8822), .ZN(n7659) );
  NAND3_X1 U8342 ( .A1(n7659), .A2(P3_REG2_REG_13__SCAN_IN), .A3(n13548), .ZN(
        n13552) );
  NOR2_X1 U8343 ( .A1(n10580), .A2(n7981), .ZN(n10581) );
  NAND2_X1 U8344 ( .A1(n9266), .A2(n9265), .ZN(n13850) );
  AOI21_X1 U8345 ( .B1(n12110), .B2(n13383), .A(n13384), .ZN(n12497) );
  OR3_X1 U8346 ( .A1(n11422), .A2(n16055), .A3(n16057), .ZN(n12707) );
  NAND2_X1 U8347 ( .A1(n13284), .A2(n13283), .ZN(n13825) );
  NAND2_X1 U8348 ( .A1(n16106), .A2(n13869), .ZN(n13860) );
  NAND2_X1 U8349 ( .A1(n6919), .A2(n6663), .ZN(n6918) );
  NAND2_X1 U8350 ( .A1(n13655), .A2(n16070), .ZN(n6919) );
  NAND2_X1 U8351 ( .A1(n7074), .A2(n9278), .ZN(n13899) );
  NAND2_X1 U8352 ( .A1(n9247), .A2(n9246), .ZN(n13911) );
  NAND2_X1 U8353 ( .A1(n9173), .A2(n9172), .ZN(n13939) );
  NAND2_X1 U8354 ( .A1(n9159), .A2(n9158), .ZN(n13942) );
  NAND2_X1 U8355 ( .A1(n9078), .A2(n9079), .ZN(n12886) );
  XNOR2_X1 U8356 ( .A(n8795), .B(n8794), .ZN(n11708) );
  NOR2_X1 U8357 ( .A1(n10553), .A2(n6634), .ZN(n7747) );
  NAND2_X1 U8358 ( .A1(n7746), .A2(n6576), .ZN(n7745) );
  INV_X1 U8359 ( .A(n7747), .ZN(n7746) );
  NAND2_X1 U8360 ( .A1(n11146), .A2(n14920), .ZN(n7180) );
  NAND2_X1 U8361 ( .A1(n14421), .A2(n14110), .ZN(n14106) );
  OAI21_X2 U8362 ( .B1(n12183), .B2(n7140), .A(n8392), .ZN(n14790) );
  NAND2_X1 U8363 ( .A1(n8516), .A2(n8515), .ZN(n14549) );
  NAND2_X1 U8364 ( .A1(n14915), .A2(n13125), .ZN(n8516) );
  NAND2_X1 U8365 ( .A1(n10560), .A2(n14736), .ZN(n14101) );
  AND2_X1 U8366 ( .A1(n14324), .A2(n14382), .ZN(n7093) );
  NAND2_X1 U8367 ( .A1(n8526), .A2(n8525), .ZN(n14396) );
  OR2_X1 U8368 ( .A1(n14087), .A2(n8648), .ZN(n8526) );
  NAND2_X1 U8369 ( .A1(n8491), .A2(n8490), .ZN(n14398) );
  CLKBUF_X2 U8370 ( .A(P2_U3947), .Z(n15887) );
  NAND2_X1 U8371 ( .A1(n11161), .A2(n11160), .ZN(n14443) );
  OAI21_X1 U8372 ( .B1(n15922), .B2(n6889), .A(n6677), .ZN(n14487) );
  NAND2_X1 U8373 ( .A1(n11234), .A2(n11214), .ZN(n11218) );
  NAND2_X1 U8374 ( .A1(n7126), .A2(n14501), .ZN(n6900) );
  INV_X1 U8375 ( .A(n7127), .ZN(n7126) );
  OAI21_X1 U8376 ( .B1(n14502), .B2(n15904), .A(n15919), .ZN(n7127) );
  XNOR2_X1 U8377 ( .A(n7183), .B(n10416), .ZN(n14747) );
  NAND2_X1 U8378 ( .A1(n10392), .A2(n10391), .ZN(n7183) );
  NOR2_X1 U8379 ( .A1(n10415), .A2(n6620), .ZN(n14746) );
  NAND2_X1 U8380 ( .A1(n7623), .A2(n7626), .ZN(n14670) );
  INV_X1 U8381 ( .A(n7625), .ZN(n7626) );
  CLKBUF_X1 U8382 ( .A(n14719), .Z(n14738) );
  INV_X1 U8383 ( .A(n11713), .ZN(n14129) );
  INV_X1 U8384 ( .A(n14703), .ZN(n14721) );
  INV_X1 U8385 ( .A(n14742), .ZN(n14723) );
  OR2_X1 U8386 ( .A1(n10395), .A2(n15980), .ZN(n10397) );
  INV_X1 U8387 ( .A(n14736), .ZN(n14713) );
  INV_X1 U8388 ( .A(n8039), .ZN(n14114) );
  INV_X1 U8389 ( .A(n14318), .ZN(n14849) );
  INV_X1 U8390 ( .A(n14519), .ZN(n14853) );
  AND2_X1 U8391 ( .A1(n7908), .A2(n6699), .ZN(n7165) );
  INV_X1 U8392 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n7309) );
  INV_X1 U8393 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n12356) );
  INV_X1 U8394 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n12184) );
  INV_X1 U8395 ( .A(n7947), .ZN(n7946) );
  AND2_X1 U8396 ( .A1(n7952), .A2(n7944), .ZN(n7943) );
  INV_X1 U8397 ( .A(n7953), .ZN(n7952) );
  AND2_X1 U8398 ( .A1(n15080), .A2(n15521), .ZN(n15062) );
  NAND2_X2 U8399 ( .A1(n9921), .A2(n9920), .ZN(n15553) );
  NAND2_X1 U8400 ( .A1(n15019), .A2(n10299), .ZN(n14959) );
  OR2_X1 U8401 ( .A1(n12143), .A2(n9812), .ZN(n9461) );
  OR2_X1 U8402 ( .A1(n15011), .A2(n15012), .ZN(n7949) );
  INV_X1 U8403 ( .A(n14980), .ZN(n7157) );
  NAND2_X1 U8404 ( .A1(n9742), .A2(n9741), .ZN(n15628) );
  INV_X1 U8405 ( .A(n15362), .ZN(n15332) );
  INV_X1 U8406 ( .A(n15080), .ZN(n15025) );
  OR2_X1 U8407 ( .A1(n10381), .A2(n12318), .ZN(n15061) );
  INV_X1 U8408 ( .A(n15062), .ZN(n15056) );
  OR2_X1 U8409 ( .A1(n11973), .A2(n9812), .ZN(n9755) );
  OR2_X1 U8410 ( .A1(n15025), .A2(n15516), .ZN(n15065) );
  AND2_X1 U8411 ( .A1(n12910), .A2(n15870), .ZN(n15068) );
  NAND2_X1 U8412 ( .A1(n9889), .A2(n9888), .ZN(n15330) );
  NAND2_X1 U8413 ( .A1(n9456), .A2(n9455), .ZN(n15363) );
  OR3_X1 U8414 ( .A1(n9729), .A2(n9728), .A3(n9727), .ZN(n15501) );
  NAND4_X2 U8415 ( .A1(n9509), .A2(n9510), .A3(n9512), .A4(n9511), .ZN(n10144)
         );
  OR2_X1 U8416 ( .A1(n6550), .A2(n15121), .ZN(n9512) );
  NAND2_X1 U8417 ( .A1(n9524), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n9511) );
  NAND2_X1 U8418 ( .A1(n11110), .A2(n11094), .ZN(n11361) );
  NAND2_X1 U8419 ( .A1(n6792), .A2(n7132), .ZN(n15540) );
  XNOR2_X1 U8420 ( .A(n15253), .B(n15541), .ZN(n6792) );
  AOI21_X1 U8421 ( .B1(n15276), .B2(n15611), .A(n15275), .ZN(n15555) );
  NAND2_X1 U8422 ( .A1(n15274), .A2(n15273), .ZN(n15275) );
  NAND2_X1 U8423 ( .A1(n9891), .A2(n9890), .ZN(n15318) );
  NAND2_X1 U8424 ( .A1(n15347), .A2(n13018), .ZN(n15327) );
  NAND2_X2 U8425 ( .A1(n7442), .A2(n9484), .ZN(n11483) );
  AND2_X1 U8426 ( .A1(n7445), .A2(n9483), .ZN(n7442) );
  OR2_X1 U8427 ( .A1(n9514), .A2(n9482), .ZN(n9483) );
  AOI21_X1 U8428 ( .B1(n15549), .B2(n7132), .A(n15548), .ZN(n15550) );
  NAND2_X1 U8429 ( .A1(n15545), .A2(n15611), .ZN(n7060) );
  OAI21_X1 U8430 ( .B1(n15562), .B2(n15620), .A(n15560), .ZN(n7154) );
  INV_X1 U8431 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n12096) );
  XNOR2_X1 U8432 ( .A(n11575), .B(n14464), .ZN(n11343) );
  NOR2_X1 U8433 ( .A1(n6841), .A2(n11942), .ZN(n6840) );
  XNOR2_X1 U8434 ( .A(n12001), .B(n12002), .ZN(n11949) );
  OAI21_X1 U8435 ( .B1(n12843), .B2(P2_ADDR_REG_12__SCAN_IN), .A(n7085), .ZN(
        n7509) );
  INV_X1 U8436 ( .A(n7510), .ZN(n7086) );
  XNOR2_X1 U8437 ( .A(n15751), .B(n15749), .ZN(n15753) );
  AND2_X1 U8438 ( .A1(n14107), .A2(n14110), .ZN(n7297) );
  OR2_X1 U8439 ( .A1(n9635), .A2(n10118), .ZN(n7241) );
  NAND2_X1 U8440 ( .A1(n7922), .A2(n7920), .ZN(n7919) );
  INV_X1 U8441 ( .A(n9584), .ZN(n7207) );
  INV_X1 U8442 ( .A(n7922), .ZN(n7238) );
  INV_X1 U8443 ( .A(n7920), .ZN(n7237) );
  INV_X1 U8444 ( .A(n9604), .ZN(n7913) );
  NAND2_X1 U8445 ( .A1(n6577), .A2(n7912), .ZN(n7911) );
  OR2_X1 U8446 ( .A1(n7913), .A2(n9606), .ZN(n7912) );
  NAND2_X1 U8447 ( .A1(n14135), .A2(n14134), .ZN(n7294) );
  NAND2_X1 U8448 ( .A1(n9636), .A2(n9638), .ZN(n7213) );
  AOI21_X1 U8449 ( .B1(n7530), .B2(n7320), .A(n7319), .ZN(n7318) );
  NOR2_X1 U8450 ( .A1(n6580), .A2(n13385), .ZN(n7387) );
  NOR2_X1 U8451 ( .A1(n14158), .A2(n14155), .ZN(n7535) );
  INV_X1 U8452 ( .A(n14155), .ZN(n7534) );
  NAND2_X1 U8453 ( .A1(n6755), .A2(n6754), .ZN(n6753) );
  AOI21_X1 U8454 ( .B1(n7396), .B2(n7398), .A(n6684), .ZN(n7395) );
  INV_X1 U8455 ( .A(n7399), .ZN(n7398) );
  OAI21_X1 U8456 ( .B1(n7386), .B2(n7384), .A(n7385), .ZN(n7383) );
  INV_X1 U8457 ( .A(n13403), .ZN(n7384) );
  AND2_X1 U8458 ( .A1(n6591), .A2(n7388), .ZN(n7386) );
  AOI21_X1 U8459 ( .B1(n7395), .B2(n7393), .A(n13426), .ZN(n7392) );
  INV_X1 U8460 ( .A(n7396), .ZN(n7393) );
  INV_X1 U8461 ( .A(n7395), .ZN(n7394) );
  NAND2_X1 U8462 ( .A1(n7301), .A2(n7304), .ZN(n7300) );
  NAND2_X1 U8463 ( .A1(n7532), .A2(n7305), .ZN(n7304) );
  NAND2_X1 U8464 ( .A1(n7143), .A2(n6640), .ZN(n14220) );
  NAND2_X1 U8465 ( .A1(n7142), .A2(n14697), .ZN(n7141) );
  NOR2_X1 U8466 ( .A1(n14203), .A2(n14189), .ZN(n14226) );
  INV_X1 U8467 ( .A(n13720), .ZN(n13438) );
  NAND2_X1 U8468 ( .A1(n14242), .A2(n14239), .ZN(n7526) );
  NAND2_X1 U8469 ( .A1(n9823), .A2(n7931), .ZN(n7928) );
  NAND2_X1 U8470 ( .A1(n6685), .A2(n7236), .ZN(n7235) );
  INV_X1 U8471 ( .A(n9810), .ZN(n7236) );
  INV_X1 U8472 ( .A(n6688), .ZN(n7930) );
  NAND2_X1 U8473 ( .A1(n6688), .A2(n7928), .ZN(n7925) );
  INV_X1 U8474 ( .A(n13454), .ZN(n7375) );
  OR2_X1 U8475 ( .A1(n7381), .A2(n13696), .ZN(n7380) );
  INV_X1 U8476 ( .A(n7526), .ZN(n7308) );
  OR2_X1 U8477 ( .A1(n14235), .A2(n14234), .ZN(n14236) );
  AND2_X1 U8478 ( .A1(n14241), .A2(n7528), .ZN(n7527) );
  INV_X1 U8479 ( .A(n14239), .ZN(n7528) );
  MUX2_X1 U8480 ( .A(n14759), .B(n14266), .S(n14265), .Z(n14285) );
  INV_X1 U8481 ( .A(n9941), .ZN(n7868) );
  NOR2_X1 U8482 ( .A1(n13331), .A2(n13677), .ZN(n7331) );
  INV_X1 U8483 ( .A(n7720), .ZN(n6909) );
  NOR2_X1 U8484 ( .A1(n10589), .A2(n12117), .ZN(n7657) );
  INV_X1 U8485 ( .A(n9255), .ZN(n7007) );
  NAND2_X1 U8486 ( .A1(n13506), .A2(n12134), .ZN(n13374) );
  AND2_X1 U8487 ( .A1(n9242), .A2(n7609), .ZN(n7608) );
  INV_X1 U8488 ( .A(n9257), .ZN(n7609) );
  MUX2_X1 U8489 ( .A(n14264), .B(n14531), .S(n14263), .Z(n14290) );
  INV_X1 U8490 ( .A(n8608), .ZN(n7022) );
  NOR2_X1 U8491 ( .A1(n6720), .A2(n7870), .ZN(n7869) );
  NOR2_X1 U8492 ( .A1(n9941), .A2(n9954), .ZN(n7870) );
  OR2_X1 U8493 ( .A1(n6749), .A2(n7107), .ZN(n6746) );
  NAND2_X1 U8494 ( .A1(n6750), .A2(n6748), .ZN(n6747) );
  NAND2_X1 U8495 ( .A1(n6749), .A2(n7107), .ZN(n6748) );
  NAND2_X1 U8496 ( .A1(n11471), .A2(n6738), .ZN(n9481) );
  OR2_X1 U8497 ( .A1(n9780), .A2(n15705), .ZN(n6738) );
  NOR2_X1 U8498 ( .A1(n9763), .A2(n15052), .ZN(n6831) );
  NOR2_X1 U8499 ( .A1(n7975), .A2(n7885), .ZN(n7884) );
  OR2_X1 U8500 ( .A1(n8431), .A2(n8430), .ZN(n7975) );
  INV_X1 U8501 ( .A(n8343), .ZN(n7882) );
  NAND2_X1 U8502 ( .A1(n8403), .A2(SI_21_), .ZN(n8434) );
  AOI21_X1 U8503 ( .B1(n8315), .B2(n8314), .A(n8313), .ZN(n8316) );
  INV_X1 U8504 ( .A(n8269), .ZN(n7879) );
  INV_X1 U8505 ( .A(n7978), .ZN(n7282) );
  AOI21_X1 U8506 ( .B1(n8230), .B2(n8229), .A(n7367), .ZN(n7288) );
  OAI21_X1 U8507 ( .B1(n9991), .B2(P2_DATAO_REG_12__SCAN_IN), .A(n7161), .ZN(
        n8232) );
  NAND2_X1 U8508 ( .A1(n9991), .A2(n11259), .ZN(n7161) );
  INV_X1 U8509 ( .A(n8177), .ZN(n7066) );
  AND2_X1 U8510 ( .A1(n8196), .A2(n8155), .ZN(n6811) );
  INV_X1 U8511 ( .A(n6618), .ZN(n7065) );
  OAI21_X1 U8512 ( .B1(n10696), .B2(n10674), .A(n7217), .ZN(n8154) );
  NAND2_X1 U8513 ( .A1(n10696), .A2(P1_DATAO_REG_7__SCAN_IN), .ZN(n7217) );
  OAI21_X1 U8514 ( .B1(n9991), .B2(n10779), .A(n7186), .ZN(n8134) );
  NAND2_X1 U8515 ( .A1(n9991), .A2(P1_DATAO_REG_6__SCAN_IN), .ZN(n7186) );
  OAI21_X1 U8516 ( .B1(n8096), .B2(n10692), .A(n7188), .ZN(n8098) );
  NAND2_X1 U8517 ( .A1(n8096), .A2(P1_DATAO_REG_5__SCAN_IN), .ZN(n7188) );
  NAND2_X1 U8518 ( .A1(n7481), .A2(n6613), .ZN(n7480) );
  NAND2_X1 U8519 ( .A1(n7482), .A2(n6613), .ZN(n7479) );
  NOR2_X1 U8520 ( .A1(n12968), .A2(n7859), .ZN(n7858) );
  INV_X1 U8521 ( .A(n12962), .ZN(n7859) );
  INV_X1 U8522 ( .A(n7147), .ZN(n7146) );
  XNOR2_X1 U8523 ( .A(n7412), .B(n8802), .ZN(n8809) );
  NAND2_X1 U8524 ( .A1(n7413), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7412) );
  NAND2_X1 U8525 ( .A1(n7403), .A2(n7402), .ZN(n8835) );
  OR2_X1 U8526 ( .A1(n8895), .A2(P3_REG2_REG_1__SCAN_IN), .ZN(n7403) );
  NAND2_X1 U8527 ( .A1(n8895), .A2(n16095), .ZN(n7402) );
  OR2_X1 U8528 ( .A1(n8939), .A2(n8929), .ZN(n7697) );
  NOR2_X1 U8529 ( .A1(n6617), .A2(n11297), .ZN(n8745) );
  NAND2_X1 U8530 ( .A1(n8835), .A2(n8834), .ZN(n11300) );
  AOI21_X1 U8531 ( .B1(n11325), .B2(n7405), .A(n7407), .ZN(n7410) );
  NOR2_X1 U8532 ( .A1(n6579), .A2(n7730), .ZN(n7726) );
  INV_X1 U8533 ( .A(n13556), .ZN(n7431) );
  NAND2_X1 U8534 ( .A1(n8779), .A2(n7979), .ZN(n8782) );
  AOI21_X1 U8535 ( .B1(n7426), .B2(n7424), .A(n7423), .ZN(n7422) );
  INV_X1 U8536 ( .A(n7426), .ZN(n7425) );
  INV_X1 U8537 ( .A(n8882), .ZN(n7424) );
  NAND2_X1 U8538 ( .A1(n13602), .A2(n7987), .ZN(n8826) );
  OAI21_X1 U8539 ( .B1(n13597), .B2(n6725), .A(n7432), .ZN(n8893) );
  OR2_X1 U8540 ( .A1(n7433), .A2(n6603), .ZN(n7432) );
  INV_X1 U8541 ( .A(n13456), .ZN(n7242) );
  AND2_X1 U8542 ( .A1(n9201), .A2(n7323), .ZN(n7322) );
  INV_X1 U8543 ( .A(P3_REG3_REG_20__SCAN_IN), .ZN(n7323) );
  INV_X1 U8544 ( .A(n6614), .ZN(n9202) );
  NOR2_X1 U8545 ( .A1(n9092), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n7321) );
  AND2_X1 U8546 ( .A1(n6627), .A2(n9048), .ZN(n7325) );
  INV_X1 U8547 ( .A(P3_REG3_REG_9__SCAN_IN), .ZN(n9048) );
  INV_X1 U8548 ( .A(P3_REG3_REG_5__SCAN_IN), .ZN(n8943) );
  INV_X1 U8549 ( .A(P3_REG3_REG_4__SCAN_IN), .ZN(n8942) );
  OR2_X1 U8550 ( .A1(n13450), .A2(n10086), .ZN(n11404) );
  OR2_X1 U8551 ( .A1(n13841), .A2(n13209), .ZN(n13452) );
  NAND2_X1 U8552 ( .A1(n13841), .A2(n13209), .ZN(n13453) );
  NAND2_X1 U8553 ( .A1(n13733), .A2(n13911), .ZN(n13440) );
  NOR2_X1 U8554 ( .A1(n7039), .A2(n7040), .ZN(n7037) );
  NOR2_X1 U8555 ( .A1(n7842), .A2(n7841), .ZN(n7840) );
  INV_X1 U8556 ( .A(n9118), .ZN(n7841) );
  NOR2_X1 U8557 ( .A1(n7552), .A2(n7248), .ZN(n7247) );
  INV_X1 U8558 ( .A(n13379), .ZN(n7248) );
  INV_X1 U8559 ( .A(n7553), .ZN(n7552) );
  AND2_X1 U8560 ( .A1(n7478), .A2(n13958), .ZN(n10088) );
  INV_X1 U8561 ( .A(n9322), .ZN(n7614) );
  NOR2_X1 U8562 ( .A1(n7607), .A2(n6944), .ZN(n6943) );
  INV_X1 U8563 ( .A(n9213), .ZN(n6944) );
  INV_X1 U8564 ( .A(n7608), .ZN(n7607) );
  INV_X1 U8565 ( .A(n7604), .ZN(n6940) );
  AOI21_X1 U8566 ( .B1(n7608), .B2(n7606), .A(n7605), .ZN(n7604) );
  INV_X1 U8567 ( .A(n9259), .ZN(n7605) );
  INV_X1 U8568 ( .A(n9238), .ZN(n7606) );
  OR2_X1 U8569 ( .A1(P3_IR_REG_18__SCAN_IN), .A2(P3_IR_REG_19__SCAN_IN), .ZN(
        n8697) );
  INV_X1 U8570 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n9183) );
  INV_X1 U8571 ( .A(n6937), .ZN(n6936) );
  OAI21_X1 U8572 ( .B1(n9104), .B2(n6938), .A(n9138), .ZN(n6937) );
  AND2_X1 U8573 ( .A1(n9140), .A2(n9137), .ZN(n9138) );
  NOR2_X1 U8574 ( .A1(n8752), .A2(P3_IR_REG_9__SCAN_IN), .ZN(n8761) );
  INV_X1 U8575 ( .A(n7586), .ZN(n7585) );
  OAI21_X1 U8576 ( .B1(n8971), .B2(n7587), .A(n8994), .ZN(n7586) );
  INV_X1 U8577 ( .A(n8958), .ZN(n7587) );
  NOR2_X1 U8578 ( .A1(n11761), .A2(n7759), .ZN(n7758) );
  INV_X1 U8579 ( .A(n10449), .ZN(n7759) );
  NOR2_X1 U8580 ( .A1(n13112), .A2(n7276), .ZN(n7275) );
  INV_X1 U8581 ( .A(n8272), .ZN(n7276) );
  NAND2_X1 U8582 ( .A1(n7268), .A2(n13112), .ZN(n7277) );
  NAND2_X1 U8583 ( .A1(n8273), .A2(n8272), .ZN(n7268) );
  XNOR2_X1 U8584 ( .A(n14749), .B(n10436), .ZN(n10548) );
  XNOR2_X1 U8585 ( .A(n7907), .B(n13112), .ZN(n10512) );
  OAI21_X1 U8586 ( .B1(n14251), .B2(n14250), .A(n14249), .ZN(n14253) );
  INV_X1 U8587 ( .A(n8527), .ZN(n7619) );
  NOR2_X1 U8588 ( .A1(n8528), .A2(n7622), .ZN(n7621) );
  INV_X1 U8589 ( .A(n8505), .ZN(n7622) );
  AOI21_X1 U8590 ( .B1(n7679), .B2(n7682), .A(n6652), .ZN(n7042) );
  NOR2_X1 U8591 ( .A1(n6673), .A2(n7179), .ZN(n7178) );
  NOR2_X1 U8592 ( .A1(n7907), .A2(n14790), .ZN(n7906) );
  AND2_X1 U8593 ( .A1(n7689), .A2(n8624), .ZN(n7049) );
  AND2_X1 U8594 ( .A1(n14353), .A2(n7691), .ZN(n7689) );
  NOR2_X1 U8595 ( .A1(n7692), .A2(n8623), .ZN(n7691) );
  NAND2_X1 U8596 ( .A1(n6825), .A2(n8306), .ZN(n14692) );
  INV_X1 U8597 ( .A(n14726), .ZN(n6825) );
  AND2_X1 U8598 ( .A1(n8299), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n8324) );
  INV_X1 U8599 ( .A(n8300), .ZN(n8299) );
  INV_X1 U8600 ( .A(n8618), .ZN(n7692) );
  NAND2_X1 U8601 ( .A1(n7169), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n8221) );
  INV_X1 U8602 ( .A(n8202), .ZN(n7169) );
  OR2_X1 U8603 ( .A1(n14154), .A2(n14159), .ZN(n6955) );
  INV_X1 U8604 ( .A(n7899), .ZN(n7897) );
  NAND2_X1 U8605 ( .A1(n8585), .A2(n7900), .ZN(n7899) );
  NAND2_X1 U8606 ( .A1(n7224), .A2(n6950), .ZN(n12917) );
  NOR2_X1 U8607 ( .A1(n14191), .A2(n14829), .ZN(n6950) );
  NOR2_X1 U8608 ( .A1(n8003), .A2(n8002), .ZN(n8004) );
  NAND4_X1 U8609 ( .A1(n8568), .A2(n8001), .A3(n8659), .A4(n8653), .ZN(n8002)
         );
  AND2_X1 U8610 ( .A1(n8001), .A2(n8568), .ZN(n7776) );
  INV_X1 U8611 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n8001) );
  INV_X1 U8612 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n8294) );
  NOR2_X1 U8613 ( .A1(n9735), .A2(n12651), .ZN(n7163) );
  INV_X1 U8614 ( .A(n10252), .ZN(n7962) );
  INV_X1 U8615 ( .A(n11467), .ZN(n10367) );
  INV_X1 U8616 ( .A(n10021), .ZN(n7212) );
  AND2_X1 U8617 ( .A1(n7990), .A2(n6626), .ZN(n7822) );
  AND2_X1 U8618 ( .A1(n15374), .A2(n13041), .ZN(n7824) );
  NAND2_X1 U8619 ( .A1(n15572), .A2(n15578), .ZN(n7461) );
  OR2_X1 U8620 ( .A1(n15602), .A2(n15390), .ZN(n13040) );
  NAND2_X1 U8621 ( .A1(n6831), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n9815) );
  AND2_X1 U8622 ( .A1(n7456), .A2(n15471), .ZN(n7458) );
  INV_X1 U8623 ( .A(n6831), .ZN(n9785) );
  NAND2_X1 U8624 ( .A1(n15633), .A2(n14993), .ZN(n10036) );
  OR2_X1 U8625 ( .A1(n15633), .A2(n14993), .ZN(n13032) );
  INV_X1 U8626 ( .A(n12555), .ZN(n7812) );
  NAND2_X1 U8627 ( .A1(n6828), .A2(n6722), .ZN(n9710) );
  AND2_X1 U8628 ( .A1(n7205), .A2(n12357), .ZN(n7788) );
  NOR2_X1 U8629 ( .A1(n15662), .A2(n15869), .ZN(n7455) );
  NOR2_X1 U8630 ( .A1(n12206), .A2(n15780), .ZN(n12340) );
  AND2_X1 U8631 ( .A1(n15792), .A2(n15843), .ZN(n7448) );
  AND2_X1 U8632 ( .A1(n7450), .A2(n7220), .ZN(n7449) );
  NAND2_X1 U8633 ( .A1(n9780), .A2(n15705), .ZN(n11471) );
  AOI21_X1 U8634 ( .B1(n13029), .B2(n6885), .A(n6883), .ZN(n6882) );
  INV_X1 U8635 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n7338) );
  INV_X1 U8636 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n7340) );
  NOR2_X1 U8637 ( .A1(n6599), .A2(n7891), .ZN(n7890) );
  XNOR2_X1 U8638 ( .A(n8507), .B(SI_25_), .ZN(n8508) );
  AOI21_X1 U8639 ( .B1(n6682), .B2(n8409), .A(n7354), .ZN(n7353) );
  INV_X1 U8640 ( .A(n8411), .ZN(n7354) );
  NAND2_X1 U8641 ( .A1(n8252), .A2(n6786), .ZN(n6785) );
  NOR2_X1 U8642 ( .A1(n6788), .A2(n6787), .ZN(n6786) );
  INV_X1 U8643 ( .A(n7988), .ZN(n6787) );
  AOI21_X1 U8644 ( .B1(n7288), .B2(n7286), .A(n7285), .ZN(n7284) );
  INV_X1 U8645 ( .A(n8229), .ZN(n7286) );
  INV_X1 U8646 ( .A(n7288), .ZN(n7287) );
  NAND2_X1 U8647 ( .A1(n8156), .A2(n8155), .ZN(n8175) );
  XNOR2_X1 U8648 ( .A(n8134), .B(SI_6_), .ZN(n8131) );
  NOR2_X1 U8649 ( .A1(n8091), .A2(n8090), .ZN(n8092) );
  NAND2_X1 U8650 ( .A1(n8089), .A2(SI_3_), .ZN(n8086) );
  INV_X1 U8651 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n9438) );
  OAI21_X1 U8652 ( .B1(n8096), .B2(P2_DATAO_REG_2__SCAN_IN), .A(n7189), .ZN(
        n8065) );
  AND2_X1 U8653 ( .A1(n10729), .A2(P3_ADDR_REG_0__SCAN_IN), .ZN(n10614) );
  XNOR2_X1 U8654 ( .A(P1_ADDR_REG_1__SCAN_IN), .B(P3_ADDR_REG_1__SCAN_IN), 
        .ZN(n10615) );
  NAND2_X1 U8655 ( .A1(n7494), .A2(n11049), .ZN(n11050) );
  NAND2_X1 U8656 ( .A1(n6835), .A2(n11943), .ZN(n6834) );
  INV_X1 U8657 ( .A(n11577), .ZN(n6835) );
  INV_X1 U8658 ( .A(n6840), .ZN(n6833) );
  NAND2_X1 U8659 ( .A1(n7484), .A2(n7483), .ZN(n7482) );
  INV_X1 U8660 ( .A(n12485), .ZN(n7483) );
  INV_X1 U8661 ( .A(n12488), .ZN(n7484) );
  NAND2_X1 U8662 ( .A1(n8988), .A2(n8987), .ZN(n9023) );
  NAND2_X1 U8663 ( .A1(n7478), .A2(n7477), .ZN(n7476) );
  NAND2_X1 U8664 ( .A1(n11431), .A2(n13332), .ZN(n7475) );
  NAND2_X1 U8665 ( .A1(n13444), .A2(n12964), .ZN(n7473) );
  XNOR2_X1 U8666 ( .A(n11436), .B(n12123), .ZN(n11650) );
  INV_X1 U8667 ( .A(n11914), .ZN(n6763) );
  NAND2_X1 U8668 ( .A1(n12933), .A2(n12934), .ZN(n7837) );
  XNOR2_X1 U8669 ( .A(n7594), .B(n13306), .ZN(n7159) );
  AND2_X1 U8670 ( .A1(n13479), .A2(n7329), .ZN(n7328) );
  AOI21_X1 U8671 ( .B1(n13478), .B2(n13479), .A(n13477), .ZN(n13480) );
  AND2_X1 U8672 ( .A1(n13290), .A2(n13289), .ZN(n13309) );
  OR2_X1 U8673 ( .A1(n9126), .A2(n11445), .ZN(n8910) );
  AND2_X1 U8674 ( .A1(n8811), .A2(P3_REG1_REG_0__SCAN_IN), .ZN(n8813) );
  XNOR2_X1 U8675 ( .A(n8939), .B(n7654), .ZN(n11299) );
  NAND2_X1 U8676 ( .A1(n8962), .A2(n6619), .ZN(n7642) );
  NAND2_X1 U8677 ( .A1(n11245), .A2(P3_REG1_REG_5__SCAN_IN), .ZN(n11397) );
  AND3_X1 U8678 ( .A1(n7720), .A2(n6628), .A3(n7719), .ZN(n8818) );
  AND2_X1 U8679 ( .A1(n9006), .A2(n6629), .ZN(n6990) );
  NAND2_X1 U8680 ( .A1(n11535), .A2(P3_REG1_REG_7__SCAN_IN), .ZN(n11698) );
  INV_X1 U8681 ( .A(n6629), .ZN(n6989) );
  NAND2_X1 U8682 ( .A1(n7415), .A2(n6660), .ZN(n12058) );
  NAND2_X1 U8683 ( .A1(n11694), .A2(n7417), .ZN(n7415) );
  NAND2_X1 U8684 ( .A1(n7417), .A2(n7420), .ZN(n7414) );
  NAND2_X1 U8685 ( .A1(n8765), .A2(n8878), .ZN(n6986) );
  NAND2_X1 U8686 ( .A1(n7736), .A2(n7735), .ZN(n13525) );
  AND2_X1 U8687 ( .A1(n13523), .A2(P3_REG1_REG_11__SCAN_IN), .ZN(n7735) );
  NOR2_X1 U8688 ( .A1(n7713), .A2(n12711), .ZN(n7708) );
  NAND2_X1 U8689 ( .A1(n13533), .A2(n7705), .ZN(n7710) );
  NAND2_X1 U8690 ( .A1(n6993), .A2(P3_REG2_REG_15__SCAN_IN), .ZN(n6992) );
  AOI21_X1 U8691 ( .B1(n6906), .B2(n6907), .A(n7713), .ZN(n13604) );
  INV_X1 U8692 ( .A(n7715), .ZN(n6907) );
  NAND2_X1 U8693 ( .A1(n8696), .A2(n6560), .ZN(n8709) );
  OR2_X1 U8694 ( .A1(n9171), .A2(n7639), .ZN(n6983) );
  AND2_X1 U8695 ( .A1(n7639), .A2(n9171), .ZN(n6984) );
  XNOR2_X1 U8696 ( .A(n8893), .B(n13641), .ZN(n13636) );
  NAND3_X1 U8697 ( .A1(n6981), .A2(n6979), .A3(n6978), .ZN(n7648) );
  NOR2_X1 U8698 ( .A1(n7651), .A2(n6980), .ZN(n6979) );
  INV_X1 U8699 ( .A(n6983), .ZN(n6980) );
  NAND2_X1 U8700 ( .A1(n7653), .A2(P3_REG2_REG_17__SCAN_IN), .ZN(n7651) );
  INV_X1 U8701 ( .A(n13623), .ZN(n7653) );
  NAND2_X1 U8702 ( .A1(n6982), .A2(n13616), .ZN(n13624) );
  NAND2_X1 U8703 ( .A1(n13590), .A2(n7639), .ZN(n6982) );
  NAND2_X1 U8704 ( .A1(n9327), .A2(n9326), .ZN(n9342) );
  NAND2_X1 U8705 ( .A1(n7846), .A2(n7003), .ZN(n13664) );
  AOI21_X1 U8706 ( .B1(n7848), .B2(n7847), .A(n6679), .ZN(n7846) );
  NAND2_X1 U8707 ( .A1(n7009), .A2(n7004), .ZN(n7003) );
  NAND2_X1 U8708 ( .A1(n9295), .A2(n9294), .ZN(n9308) );
  NAND2_X1 U8709 ( .A1(n7849), .A2(n9286), .ZN(n13680) );
  NAND2_X1 U8710 ( .A1(n7849), .A2(n7848), .ZN(n13682) );
  OR2_X1 U8711 ( .A1(n9267), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n9279) );
  NAND2_X1 U8712 ( .A1(n13707), .A2(n13704), .ZN(n13708) );
  OR2_X1 U8713 ( .A1(n9248), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n9267) );
  NAND2_X1 U8714 ( .A1(n9202), .A2(n7322), .ZN(n9231) );
  NAND2_X1 U8715 ( .A1(n13790), .A2(n9180), .ZN(n13771) );
  NAND2_X1 U8716 ( .A1(n7324), .A2(n9174), .ZN(n9187) );
  NAND2_X1 U8717 ( .A1(n9146), .A2(n9145), .ZN(n9162) );
  INV_X1 U8718 ( .A(n9147), .ZN(n9146) );
  NAND2_X1 U8719 ( .A1(n9111), .A2(n9110), .ZN(n9127) );
  INV_X1 U8720 ( .A(P3_REG3_REG_13__SCAN_IN), .ZN(n9110) );
  INV_X1 U8721 ( .A(n9112), .ZN(n9111) );
  NAND2_X1 U8722 ( .A1(n7321), .A2(n9081), .ZN(n9112) );
  INV_X1 U8723 ( .A(P3_REG3_REG_12__SCAN_IN), .ZN(n9081) );
  INV_X1 U8724 ( .A(n7321), .ZN(n9094) );
  NAND2_X1 U8725 ( .A1(n13315), .A2(n13370), .ZN(n7559) );
  INV_X1 U8726 ( .A(n7563), .ZN(n7558) );
  NAND4_X1 U8727 ( .A1(n8942), .A2(n11684), .A3(n7327), .A4(n8943), .ZN(n9011)
         );
  INV_X1 U8728 ( .A(P3_REG3_REG_6__SCAN_IN), .ZN(n7327) );
  INV_X1 U8729 ( .A(n13358), .ZN(n9403) );
  NAND2_X1 U8730 ( .A1(n11684), .A2(n8942), .ZN(n8965) );
  INV_X1 U8731 ( .A(n13347), .ZN(n16027) );
  AND2_X1 U8732 ( .A1(n11404), .A2(n9397), .ZN(n10108) );
  AND2_X1 U8733 ( .A1(n13646), .A2(n13645), .ZN(n13888) );
  OAI21_X1 U8734 ( .B1(n13132), .B2(n9353), .A(n9354), .ZN(n10100) );
  NAND2_X1 U8735 ( .A1(n13452), .A2(n13453), .ZN(n13677) );
  NAND2_X1 U8736 ( .A1(n13441), .A2(n13440), .ZN(n13720) );
  AOI21_X1 U8737 ( .B1(n13735), .B2(n9355), .A(n9235), .ZN(n13749) );
  NAND2_X1 U8738 ( .A1(n7257), .A2(n13427), .ZN(n7254) );
  AOI21_X1 U8739 ( .B1(n7257), .B2(n13783), .A(n7256), .ZN(n7255) );
  INV_X1 U8740 ( .A(n13420), .ZN(n7256) );
  AND2_X1 U8741 ( .A1(n13431), .A2(n13432), .ZN(n13745) );
  NAND2_X1 U8742 ( .A1(n13800), .A2(n13801), .ZN(n7038) );
  AND3_X1 U8743 ( .A1(n9166), .A2(n9165), .A3(n9164), .ZN(n13818) );
  NAND2_X1 U8744 ( .A1(n12699), .A2(n9118), .ZN(n12767) );
  NAND2_X1 U8745 ( .A1(n12767), .A2(n13402), .ZN(n12766) );
  INV_X1 U8746 ( .A(n13325), .ZN(n13402) );
  AND4_X1 U8747 ( .A1(n9134), .A2(n9133), .A3(n9132), .A4(n9131), .ZN(n13816)
         );
  NAND2_X1 U8748 ( .A1(n12403), .A2(n13391), .ZN(n12447) );
  NAND2_X1 U8749 ( .A1(n13395), .A2(n13396), .ZN(n13323) );
  OR2_X1 U8750 ( .A1(n13959), .A2(n8792), .ZN(n11422) );
  AND2_X1 U8751 ( .A1(n10088), .A2(n10090), .ZN(n11424) );
  OAI21_X1 U8752 ( .B1(n9350), .B2(n9349), .A(n9348), .ZN(n9352) );
  XNOR2_X1 U8753 ( .A(n8714), .B(P3_IR_REG_26__SCAN_IN), .ZN(n9381) );
  AND2_X1 U8754 ( .A1(n9290), .A2(n6736), .ZN(n7579) );
  INV_X1 U8755 ( .A(n6558), .ZN(n8716) );
  OAI21_X1 U8756 ( .B1(n9212), .B2(n6942), .A(n6939), .ZN(n9263) );
  AOI21_X1 U8757 ( .B1(n6943), .B2(n6941), .A(n6940), .ZN(n6939) );
  INV_X1 U8758 ( .A(n6943), .ZN(n6942) );
  INV_X1 U8759 ( .A(n9211), .ZN(n6941) );
  NAND2_X1 U8760 ( .A1(n9263), .A2(n9262), .ZN(n9277) );
  INV_X1 U8761 ( .A(P3_IR_REG_21__SCAN_IN), .ZN(n8797) );
  OR2_X1 U8762 ( .A1(n8776), .A2(P3_IR_REG_13__SCAN_IN), .ZN(n8780) );
  NAND2_X1 U8763 ( .A1(n9105), .A2(n9104), .ZN(n6935) );
  AOI21_X1 U8764 ( .B1(n7601), .B2(n7603), .A(n7600), .ZN(n7599) );
  OAI21_X1 U8765 ( .B1(n8999), .B2(n6929), .A(n6927), .ZN(n7598) );
  INV_X1 U8766 ( .A(n9058), .ZN(n7600) );
  INV_X1 U8767 ( .A(n8761), .ZN(n8759) );
  XNOR2_X1 U8768 ( .A(n15995), .B(n10436), .ZN(n10456) );
  INV_X1 U8769 ( .A(n7758), .ZN(n7757) );
  NAND2_X1 U8770 ( .A1(n8142), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n8165) );
  INV_X1 U8771 ( .A(n8144), .ZN(n8142) );
  NOR2_X1 U8772 ( .A1(n7273), .A2(n7269), .ZN(n13980) );
  AOI21_X1 U8773 ( .B1(n7274), .B2(n7277), .A(n7272), .ZN(n7273) );
  AND2_X1 U8774 ( .A1(n7277), .A2(n7271), .ZN(n7269) );
  AND2_X1 U8775 ( .A1(n7274), .A2(n7272), .ZN(n7271) );
  AOI21_X1 U8776 ( .B1(n7765), .B2(n14040), .A(n6681), .ZN(n7763) );
  INV_X1 U8777 ( .A(n7765), .ZN(n7764) );
  NAND2_X1 U8778 ( .A1(n10512), .A2(n10513), .ZN(n14002) );
  NAND2_X1 U8779 ( .A1(n6973), .A2(n7750), .ZN(n6968) );
  NAND2_X1 U8780 ( .A1(n12889), .A2(n6973), .ZN(n6967) );
  XNOR2_X1 U8781 ( .A(n14769), .B(n10436), .ZN(n10534) );
  XNOR2_X1 U8782 ( .A(n10436), .B(n14129), .ZN(n10433) );
  NAND2_X1 U8783 ( .A1(n8163), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n8185) );
  INV_X1 U8784 ( .A(n8165), .ZN(n8163) );
  INV_X1 U8785 ( .A(n7171), .ZN(n8394) );
  NAND2_X1 U8786 ( .A1(n7171), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n8423) );
  INV_X1 U8787 ( .A(n8245), .ZN(n8243) );
  INV_X1 U8788 ( .A(n7170), .ZN(n8275) );
  INV_X1 U8789 ( .A(n14376), .ZN(n14095) );
  AND2_X1 U8790 ( .A1(n11513), .A2(n11512), .ZN(n10430) );
  NAND2_X1 U8791 ( .A1(n8353), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n8372) );
  XNOR2_X1 U8792 ( .A(n14800), .B(n13112), .ZN(n10511) );
  NAND2_X1 U8793 ( .A1(n11740), .A2(n11741), .ZN(n11739) );
  AOI21_X1 U8794 ( .B1(n12889), .B2(n7751), .A(n7750), .ZN(n7749) );
  NOR2_X1 U8795 ( .A1(n10564), .A2(n10554), .ZN(n10559) );
  INV_X1 U8796 ( .A(n14107), .ZN(n14323) );
  AND2_X1 U8797 ( .A1(n6799), .A2(n6584), .ZN(n6798) );
  INV_X1 U8798 ( .A(n14314), .ZN(n6799) );
  AND2_X1 U8799 ( .A1(n8453), .A2(n8452), .ZN(n14254) );
  OR2_X1 U8800 ( .A1(n11232), .A2(n11233), .ZN(n11230) );
  OR2_X1 U8801 ( .A1(n11218), .A2(n11217), .ZN(n11528) );
  OR2_X1 U8802 ( .A1(n11723), .A2(n11724), .ZN(n11929) );
  INV_X1 U8803 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n12925) );
  NAND2_X1 U8804 ( .A1(n11925), .A2(n11924), .ZN(n11987) );
  NAND2_X1 U8805 ( .A1(n6876), .A2(n6874), .ZN(n12797) );
  AOI21_X1 U8806 ( .B1(n6877), .B2(n6879), .A(n6875), .ZN(n6874) );
  INV_X1 U8807 ( .A(n12795), .ZN(n6875) );
  OR2_X1 U8808 ( .A1(n12797), .A2(n12806), .ZN(n14497) );
  OR2_X1 U8809 ( .A1(n12800), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n14498) );
  AND2_X1 U8810 ( .A1(n7904), .A2(n14511), .ZN(n7901) );
  INV_X1 U8811 ( .A(n14530), .ZN(n7903) );
  NOR2_X1 U8812 ( .A1(n14530), .A2(n7902), .ZN(n12987) );
  INV_X1 U8813 ( .A(n7904), .ZN(n7902) );
  INV_X1 U8814 ( .A(n10412), .ZN(n10413) );
  OR2_X1 U8815 ( .A1(n14363), .A2(n8640), .ZN(n10414) );
  OAI211_X1 U8816 ( .C1(n7620), .C2(n7051), .A(n14362), .B(n7050), .ZN(n10392)
         );
  INV_X1 U8817 ( .A(n8540), .ZN(n7051) );
  NAND2_X1 U8818 ( .A1(n7618), .A2(n8540), .ZN(n7050) );
  NAND2_X1 U8819 ( .A1(n7355), .A2(n6649), .ZN(n10418) );
  NOR2_X1 U8820 ( .A1(n8539), .A2(n7357), .ZN(n7356) );
  AND2_X1 U8821 ( .A1(n8649), .A2(n11151), .ZN(n14376) );
  AND2_X1 U8822 ( .A1(n8649), .A2(n11179), .ZN(n14086) );
  NAND2_X1 U8823 ( .A1(n7358), .A2(n7359), .ZN(n8639) );
  INV_X1 U8824 ( .A(n14549), .ZN(n14759) );
  NOR2_X2 U8825 ( .A1(n14572), .A2(n14562), .ZN(n14561) );
  OR2_X1 U8826 ( .A1(n8497), .A2(n14020), .ZN(n8519) );
  NAND2_X1 U8827 ( .A1(n8483), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n8497) );
  INV_X1 U8828 ( .A(n8484), .ZN(n8483) );
  NAND2_X1 U8829 ( .A1(n7041), .A2(n7042), .ZN(n14556) );
  NAND2_X1 U8830 ( .A1(n6581), .A2(n14676), .ZN(n14596) );
  NAND2_X1 U8831 ( .A1(n7632), .A2(n7630), .ZN(n14589) );
  OR2_X1 U8832 ( .A1(n14610), .A2(n14609), .ZN(n14612) );
  NAND2_X1 U8833 ( .A1(n7668), .A2(n8628), .ZN(n7667) );
  AND2_X1 U8834 ( .A1(n7670), .A2(n14647), .ZN(n7668) );
  NAND2_X1 U8835 ( .A1(n7906), .A2(n14676), .ZN(n14639) );
  NAND2_X1 U8836 ( .A1(n7099), .A2(n6666), .ZN(n7625) );
  NAND2_X1 U8837 ( .A1(n8341), .A2(n14693), .ZN(n7099) );
  NOR2_X1 U8838 ( .A1(n14671), .A2(n7625), .ZN(n7624) );
  NOR2_X1 U8839 ( .A1(n7989), .A2(n14697), .ZN(n14696) );
  NAND2_X1 U8840 ( .A1(n7115), .A2(n7114), .ZN(n7989) );
  NAND2_X1 U8841 ( .A1(n7170), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n8300) );
  INV_X1 U8842 ( .A(n7635), .ZN(n7634) );
  OAI21_X1 U8843 ( .B1(n7636), .B2(n6616), .A(n8267), .ZN(n7635) );
  NAND2_X1 U8844 ( .A1(n7224), .A2(n14173), .ZN(n12834) );
  AOI21_X1 U8845 ( .B1(n14344), .B2(n7018), .A(n7017), .ZN(n7016) );
  INV_X1 U8846 ( .A(n8191), .ZN(n7018) );
  INV_X1 U8847 ( .A(n8210), .ZN(n7017) );
  NAND2_X1 U8848 ( .A1(n12456), .A2(n8610), .ZN(n12659) );
  NAND2_X1 U8849 ( .A1(n8609), .A2(n8608), .ZN(n12456) );
  AOI21_X1 U8850 ( .B1(n7675), .B2(n8600), .A(n6669), .ZN(n7674) );
  NAND2_X1 U8851 ( .A1(n8600), .A2(n7677), .ZN(n7676) );
  NAND2_X1 U8852 ( .A1(n6954), .A2(n7233), .ZN(n12384) );
  NOR2_X1 U8853 ( .A1(n7616), .A2(n14341), .ZN(n7011) );
  INV_X1 U8854 ( .A(n8150), .ZN(n7616) );
  INV_X1 U8855 ( .A(n11816), .ZN(n7191) );
  NOR2_X1 U8856 ( .A1(n14846), .A2(n7516), .ZN(n10396) );
  NAND2_X1 U8857 ( .A1(n14331), .A2(n11771), .ZN(n8588) );
  INV_X1 U8858 ( .A(n11625), .ZN(n14332) );
  NOR2_X2 U8859 ( .A1(n11769), .A2(n14120), .ZN(n11676) );
  NOR2_X1 U8860 ( .A1(n7741), .A2(n7516), .ZN(n11909) );
  INV_X1 U8861 ( .A(n11633), .ZN(n10395) );
  AOI22_X1 U8862 ( .A1(n13126), .A2(P1_DATAO_REG_4__SCAN_IN), .B1(n8368), .B2(
        n14440), .ZN(n8084) );
  AND2_X1 U8863 ( .A1(n8004), .A2(n7909), .ZN(n7908) );
  INV_X1 U8864 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n7909) );
  INV_X1 U8865 ( .A(n8661), .ZN(n8654) );
  INV_X1 U8866 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n8567) );
  OR2_X1 U8867 ( .A1(n8239), .A2(P2_IR_REG_12__SCAN_IN), .ZN(n8270) );
  OR2_X1 U8868 ( .A1(n8137), .A2(P2_IR_REG_6__SCAN_IN), .ZN(n8157) );
  NAND3_X1 U8869 ( .A1(n7665), .A2(n7664), .A3(n8051), .ZN(n8100) );
  NAND2_X1 U8870 ( .A1(n6893), .A2(n8068), .ZN(n8077) );
  INV_X1 U8871 ( .A(n8067), .ZN(n6893) );
  XNOR2_X1 U8872 ( .A(n8034), .B(P2_IR_REG_1__SCAN_IN), .ZN(n11155) );
  NOR2_X1 U8873 ( .A1(n15060), .A2(n7948), .ZN(n7947) );
  INV_X1 U8874 ( .A(n7950), .ZN(n7948) );
  OAI21_X1 U8875 ( .B1(n15060), .B2(n7954), .A(n10334), .ZN(n7953) );
  NAND2_X1 U8876 ( .A1(n7947), .A2(n7945), .ZN(n7944) );
  INV_X1 U8877 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n9639) );
  OR2_X1 U8878 ( .A1(n9640), .A2(n9639), .ZN(n9661) );
  NAND2_X1 U8879 ( .A1(n10340), .A2(n11798), .ZN(n10145) );
  NAND2_X1 U8880 ( .A1(n7162), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n9678) );
  INV_X1 U8881 ( .A(n9661), .ZN(n7162) );
  NAND2_X1 U8882 ( .A1(n6828), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n9708) );
  NAND2_X1 U8883 ( .A1(n6829), .A2(n9848), .ZN(n9881) );
  NAND2_X1 U8884 ( .A1(n7163), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n9763) );
  INV_X1 U8885 ( .A(n7163), .ZN(n9761) );
  INV_X1 U8886 ( .A(n7200), .ZN(n10202) );
  INV_X1 U8887 ( .A(n6829), .ZN(n9851) );
  AND2_X1 U8888 ( .A1(n7951), .A2(n14980), .ZN(n7950) );
  NAND2_X1 U8889 ( .A1(n15012), .A2(n7955), .ZN(n7951) );
  AOI21_X1 U8890 ( .B1(n7025), .B2(n7027), .A(n7945), .ZN(n7024) );
  INV_X1 U8891 ( .A(n7029), .ZN(n7025) );
  AOI21_X1 U8892 ( .B1(n10367), .B2(n10686), .A(n10685), .ZN(n11827) );
  NAND2_X1 U8893 ( .A1(n14931), .A2(n10252), .ZN(n14989) );
  AND2_X1 U8894 ( .A1(n10257), .A2(n10256), .ZN(n14988) );
  AND2_X1 U8895 ( .A1(n6631), .A2(n9984), .ZN(n7240) );
  NAND2_X1 U8896 ( .A1(n7083), .A2(n6661), .ZN(n9985) );
  NOR2_X1 U8897 ( .A1(n9983), .A2(n9982), .ZN(n9984) );
  AND4_X1 U8898 ( .A1(n9568), .A2(n9567), .A3(n9566), .A4(n9565), .ZN(n12030)
         );
  INV_X1 U8899 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n15101) );
  NOR2_X2 U8900 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n9515) );
  NAND2_X1 U8901 ( .A1(n6861), .A2(n6860), .ZN(n11559) );
  INV_X1 U8902 ( .A(n11366), .ZN(n6860) );
  INV_X1 U8903 ( .A(n11365), .ZN(n6861) );
  OR2_X1 U8904 ( .A1(n11553), .A2(n11554), .ZN(n11897) );
  AND2_X1 U8905 ( .A1(n12166), .A2(n12165), .ZN(n15186) );
  OR2_X1 U8906 ( .A1(n11899), .A2(n11900), .ZN(n12161) );
  INV_X1 U8907 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n14935) );
  XNOR2_X1 U8908 ( .A(n12634), .B(n12644), .ZN(n12632) );
  NAND2_X1 U8909 ( .A1(n12632), .A2(n12631), .ZN(n6864) );
  AND2_X1 U8910 ( .A1(n10720), .A2(n7827), .ZN(n10722) );
  NAND2_X1 U8911 ( .A1(n6864), .A2(n6862), .ZN(n15199) );
  NOR2_X1 U8912 ( .A1(n6863), .A2(n12638), .ZN(n6862) );
  INV_X1 U8913 ( .A(n12635), .ZN(n6863) );
  OR2_X1 U8914 ( .A1(n12649), .A2(n12650), .ZN(n15207) );
  NAND2_X1 U8915 ( .A1(n15216), .A2(n15215), .ZN(n15217) );
  INV_X1 U8916 ( .A(n7227), .ZN(n7064) );
  NOR2_X1 U8917 ( .A1(n13067), .A2(n13069), .ZN(n13070) );
  NAND2_X1 U8918 ( .A1(n9970), .A2(n9969), .ZN(n13076) );
  AND2_X1 U8919 ( .A1(n15280), .A2(n15547), .ZN(n15260) );
  AND2_X1 U8920 ( .A1(n13054), .A2(n6637), .ZN(n7806) );
  INV_X1 U8921 ( .A(n15267), .ZN(n7808) );
  NAND2_X1 U8922 ( .A1(n7341), .A2(n7345), .ZN(n15271) );
  AOI21_X1 U8923 ( .B1(n15295), .B2(n13053), .A(n13054), .ZN(n15270) );
  NAND2_X1 U8924 ( .A1(n13065), .A2(n6578), .ZN(n7139) );
  NAND2_X1 U8925 ( .A1(n15297), .A2(n15521), .ZN(n15273) );
  NAND2_X1 U8926 ( .A1(n15288), .A2(n15293), .ZN(n7807) );
  OAI21_X1 U8927 ( .B1(n15270), .B2(n7817), .A(n15611), .ZN(n7816) );
  AND3_X1 U8928 ( .A1(n15295), .A2(n13054), .A3(n13053), .ZN(n7817) );
  NOR2_X1 U8929 ( .A1(n15336), .A2(n7461), .ZN(n15312) );
  NOR2_X1 U8930 ( .A1(n15336), .A2(n15341), .ZN(n15338) );
  NOR2_X1 U8931 ( .A1(n13012), .A2(n7800), .ZN(n7799) );
  INV_X1 U8932 ( .A(n13010), .ZN(n7800) );
  OR2_X1 U8933 ( .A1(n9817), .A2(n14961), .ZN(n9828) );
  NOR2_X1 U8934 ( .A1(n15408), .A2(n15597), .ZN(n15392) );
  XNOR2_X1 U8935 ( .A(n15597), .B(n15045), .ZN(n15385) );
  NAND3_X1 U8936 ( .A1(n7458), .A2(n6572), .A3(n7457), .ZN(n15408) );
  OR2_X1 U8937 ( .A1(n15400), .A2(n15404), .ZN(n15402) );
  NAND2_X1 U8938 ( .A1(n7458), .A2(n6572), .ZN(n15418) );
  NAND2_X1 U8939 ( .A1(n7068), .A2(n7069), .ZN(n13009) );
  INV_X1 U8940 ( .A(n7070), .ZN(n7069) );
  OR2_X1 U8941 ( .A1(n9710), .A2(n14935), .ZN(n9724) );
  NAND2_X1 U8942 ( .A1(n9434), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n9735) );
  INV_X1 U8943 ( .A(n9724), .ZN(n9434) );
  NAND2_X1 U8944 ( .A1(n12367), .A2(n12368), .ZN(n12723) );
  NAND2_X1 U8945 ( .A1(n12340), .A2(n12207), .ZN(n12342) );
  NAND2_X1 U8946 ( .A1(n9432), .A2(n6668), .ZN(n9624) );
  NAND2_X1 U8947 ( .A1(n9432), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n9609) );
  AOI22_X1 U8948 ( .A1(n9513), .A2(P2_DATAO_REG_4__SCAN_IN), .B1(n9781), .B2(
        n11079), .ZN(n9551) );
  NAND2_X1 U8949 ( .A1(n11849), .A2(n11799), .ZN(n11955) );
  NAND2_X1 U8950 ( .A1(n11956), .A2(n15834), .ZN(n11799) );
  AOI21_X1 U8951 ( .B1(n9513), .B2(P2_DATAO_REG_3__SCAN_IN), .A(n7801), .ZN(
        n7803) );
  NOR2_X1 U8952 ( .A1(n9812), .A2(n7802), .ZN(n7801) );
  INV_X1 U8953 ( .A(n7449), .ZN(n11964) );
  AND2_X1 U8954 ( .A1(n7133), .A2(n12140), .ZN(n15810) );
  NOR2_X1 U8955 ( .A1(n11483), .A2(n7137), .ZN(n11853) );
  NAND2_X1 U8956 ( .A1(n7136), .A2(n12043), .ZN(n10028) );
  OR2_X1 U8957 ( .A1(n10378), .A2(n11071), .ZN(n15516) );
  AOI211_X1 U8958 ( .C1(n7122), .C2(n6625), .A(n15608), .B(n13059), .ZN(n15558) );
  NAND2_X1 U8959 ( .A1(n13000), .A2(n12999), .ZN(n15533) );
  AND2_X1 U8960 ( .A1(n11469), .A2(n11468), .ZN(n11828) );
  AND2_X1 U8961 ( .A1(n10607), .A2(n10687), .ZN(n10684) );
  NAND2_X1 U8962 ( .A1(n15689), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9446) );
  XNOR2_X1 U8963 ( .A(n9968), .B(n9967), .ZN(n14902) );
  NAND2_X1 U8964 ( .A1(n7889), .A2(n7887), .ZN(n9934) );
  INV_X1 U8965 ( .A(n7888), .ZN(n7887) );
  NAND2_X1 U8966 ( .A1(n8512), .A2(n7890), .ZN(n7889) );
  OAI21_X1 U8967 ( .B1(n8529), .B2(n6599), .A(n8542), .ZN(n7888) );
  XNOR2_X1 U8968 ( .A(n7790), .B(n9458), .ZN(n10073) );
  NAND2_X1 U8969 ( .A1(n9457), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7790) );
  NAND2_X1 U8970 ( .A1(n9459), .A2(n9444), .ZN(n9457) );
  NAND2_X1 U8971 ( .A1(n8530), .A2(n8529), .ZN(n6794) );
  AND2_X1 U8972 ( .A1(n10070), .A2(n10069), .ZN(n10356) );
  MUX2_X1 U8973 ( .A(P1_IR_REG_31__SCAN_IN), .B(n10068), .S(
        P1_IR_REG_26__SCAN_IN), .Z(n10070) );
  NAND2_X1 U8974 ( .A1(n10067), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10068) );
  XNOR2_X1 U8975 ( .A(n8509), .B(n8508), .ZN(n12789) );
  NAND2_X1 U8976 ( .A1(n8493), .A2(n7895), .ZN(n8509) );
  AND2_X1 U8977 ( .A1(n8494), .A2(n8480), .ZN(n12577) );
  NAND2_X1 U8978 ( .A1(n8493), .A2(n7894), .ZN(n8494) );
  NAND2_X1 U8979 ( .A1(n8493), .A2(n8477), .ZN(n8479) );
  XNOR2_X1 U8980 ( .A(n8366), .B(n8385), .ZN(n12141) );
  NAND2_X1 U8981 ( .A1(n8364), .A2(n8347), .ZN(n8348) );
  OR2_X2 U8982 ( .A1(n8348), .A2(n8383), .ZN(n8365) );
  INV_X1 U8983 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n6759) );
  NAND2_X1 U8984 ( .A1(n6789), .A2(n7363), .ZN(n8329) );
  NAND2_X1 U8985 ( .A1(n8252), .A2(n7365), .ZN(n6789) );
  XNOR2_X1 U8986 ( .A(n8289), .B(n8288), .ZN(n11666) );
  NAND2_X1 U8987 ( .A1(n7863), .A2(n8196), .ZN(n8212) );
  NAND2_X1 U8988 ( .A1(n8194), .A2(n8193), .ZN(n7863) );
  OR2_X1 U8989 ( .A1(n9631), .A2(n9630), .ZN(n9647) );
  XNOR2_X1 U8990 ( .A(n8175), .B(n8173), .ZN(n10711) );
  OR2_X1 U8991 ( .A1(n9580), .A2(P1_IR_REG_5__SCAN_IN), .ZN(n9720) );
  NAND2_X1 U8992 ( .A1(n7352), .A2(n7350), .ZN(n8063) );
  XNOR2_X1 U8993 ( .A(n8065), .B(SI_2_), .ZN(n8064) );
  NAND2_X1 U8994 ( .A1(n7057), .A2(n8030), .ZN(n9499) );
  NAND2_X1 U8995 ( .A1(n6844), .A2(n10626), .ZN(n10627) );
  NAND2_X1 U8996 ( .A1(n6844), .A2(n6588), .ZN(n10628) );
  INV_X1 U8997 ( .A(P3_ADDR_REG_3__SCAN_IN), .ZN(n6843) );
  XNOR2_X1 U8998 ( .A(n11050), .B(n10678), .ZN(n11045) );
  NAND2_X1 U8999 ( .A1(n11342), .A2(n11341), .ZN(n11575) );
  NAND2_X1 U9000 ( .A1(n11578), .A2(n11338), .ZN(n11579) );
  NAND2_X1 U9001 ( .A1(n12010), .A2(n12009), .ZN(n12015) );
  OR2_X1 U9002 ( .A1(n12007), .A2(n12006), .ZN(n12010) );
  OR2_X1 U9003 ( .A1(n12015), .A2(n12014), .ZN(n12329) );
  NAND2_X1 U9004 ( .A1(n7514), .A2(P2_ADDR_REG_11__SCAN_IN), .ZN(n7513) );
  INV_X1 U9005 ( .A(n12332), .ZN(n7514) );
  OAI21_X1 U9006 ( .B1(n7513), .B2(n7512), .A(n7511), .ZN(n7510) );
  INV_X1 U9007 ( .A(n12842), .ZN(n7511) );
  INV_X1 U9008 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n7515) );
  AOI21_X1 U9009 ( .B1(n13652), .B2(n9355), .A(n9346), .ZN(n12979) );
  AOI21_X1 U9010 ( .B1(n7855), .B2(n7857), .A(n6676), .ZN(n7853) );
  NAND2_X1 U9011 ( .A1(n9325), .A2(n9324), .ZN(n13460) );
  NAND2_X1 U9012 ( .A1(n7832), .A2(n7835), .ZN(n13151) );
  NAND2_X1 U9013 ( .A1(n9200), .A2(n9199), .ZN(n13172) );
  AND2_X1 U9014 ( .A1(n13290), .A2(n9361), .ZN(n13300) );
  NAND2_X1 U9015 ( .A1(n13212), .A2(n12956), .ZN(n13174) );
  AND2_X1 U9016 ( .A1(n9316), .A2(n9315), .ZN(n13684) );
  NAND2_X1 U9017 ( .A1(n7854), .A2(n12967), .ZN(n13255) );
  AOI21_X1 U9018 ( .B1(n7491), .B2(n7830), .A(n6664), .ZN(n7489) );
  NAND2_X1 U9019 ( .A1(n7486), .A2(n6764), .ZN(n11915) );
  NAND2_X1 U9020 ( .A1(n6775), .A2(n12945), .ZN(n13196) );
  NOR2_X1 U9021 ( .A1(n12256), .A2(n12257), .ZN(n12486) );
  NAND2_X1 U9022 ( .A1(n12935), .A2(n7837), .ZN(n13222) );
  OAI211_X2 U9023 ( .C1(n8939), .C2(n9367), .A(n8938), .B(n8937), .ZN(n16036)
         );
  OR2_X1 U9024 ( .A1(n6568), .A2(SI_2_), .ZN(n8937) );
  INV_X1 U9025 ( .A(n6773), .ZN(n6772) );
  OAI21_X1 U9026 ( .B1(n12945), .B2(n6774), .A(n13245), .ZN(n6773) );
  INV_X1 U9027 ( .A(n12948), .ZN(n6774) );
  NAND2_X1 U9028 ( .A1(n13196), .A2(n12948), .ZN(n13246) );
  NAND2_X1 U9029 ( .A1(n7493), .A2(n7828), .ZN(n13266) );
  INV_X1 U9030 ( .A(n13684), .ZN(n13494) );
  INV_X1 U9031 ( .A(n13733), .ZN(n13705) );
  NAND2_X1 U9032 ( .A1(n9208), .A2(n9207), .ZN(n13775) );
  OR2_X1 U9033 ( .A1(n9372), .A2(n16104), .ZN(n9027) );
  OR2_X1 U9034 ( .A1(n9311), .A2(n7654), .ZN(n8931) );
  CLKBUF_X1 U9035 ( .A(n16030), .Z(n7149) );
  INV_X1 U9036 ( .A(P3_ADDR_REG_2__SCAN_IN), .ZN(n11307) );
  INV_X1 U9037 ( .A(n7704), .ZN(n11318) );
  NAND2_X1 U9038 ( .A1(n7699), .A2(n7700), .ZN(n11273) );
  NAND2_X1 U9039 ( .A1(n7409), .A2(n11325), .ZN(n11327) );
  NAND2_X1 U9040 ( .A1(n11303), .A2(n11324), .ZN(n7409) );
  NAND2_X1 U9041 ( .A1(n8853), .A2(n11252), .ZN(n11388) );
  NAND2_X1 U9042 ( .A1(n7416), .A2(n11692), .ZN(n12056) );
  NAND2_X1 U9043 ( .A1(n11694), .A2(n11693), .ZN(n7416) );
  NAND2_X1 U9044 ( .A1(n7723), .A2(n6912), .ZN(n12049) );
  NAND2_X1 U9045 ( .A1(n6914), .A2(n7723), .ZN(n6913) );
  AOI21_X1 U9046 ( .B1(n12051), .B2(n7196), .A(n10589), .ZN(n10588) );
  NAND2_X1 U9047 ( .A1(n7736), .A2(n13523), .ZN(n12592) );
  AOI21_X1 U9048 ( .B1(n13552), .B2(n13548), .A(n8885), .ZN(n13551) );
  NAND2_X1 U9049 ( .A1(n13519), .A2(n8882), .ZN(n7421) );
  OR2_X1 U9050 ( .A1(n6992), .A2(n6991), .ZN(n13591) );
  NAND2_X1 U9051 ( .A1(n7435), .A2(n13594), .ZN(n13612) );
  NAND2_X1 U9052 ( .A1(n7437), .A2(n7436), .ZN(n7435) );
  NAND2_X1 U9053 ( .A1(n7648), .A2(n7649), .ZN(n13627) );
  NAND2_X1 U9054 ( .A1(n7650), .A2(n7653), .ZN(n7649) );
  INV_X1 U9055 ( .A(n13624), .ZN(n7650) );
  NAND2_X1 U9056 ( .A1(n6593), .A2(n7438), .ZN(n6915) );
  NOR2_X1 U9057 ( .A1(n7439), .A2(n8900), .ZN(n7438) );
  INV_X1 U9058 ( .A(n10113), .ZN(n9428) );
  NAND2_X1 U9059 ( .A1(n7243), .A2(n7244), .ZN(n13669) );
  NAND2_X1 U9060 ( .A1(n13707), .A2(n7245), .ZN(n7243) );
  NAND2_X1 U9061 ( .A1(n6559), .A2(n9223), .ZN(n13730) );
  NAND2_X1 U9062 ( .A1(n12114), .A2(n9055), .ZN(n12500) );
  NAND2_X1 U9063 ( .A1(n11866), .A2(n13365), .ZN(n12125) );
  INV_X1 U9064 ( .A(n13814), .ZN(n13737) );
  INV_X1 U9065 ( .A(P3_REG3_REG_3__SCAN_IN), .ZN(n11684) );
  OR2_X1 U9066 ( .A1(n10104), .A2(n13306), .ZN(n16057) );
  AND2_X1 U9067 ( .A1(n9422), .A2(n12707), .ZN(n16066) );
  INV_X1 U9068 ( .A(n11647), .ZN(n12123) );
  INV_X1 U9069 ( .A(n13860), .ZN(n13880) );
  NOR2_X1 U9070 ( .A1(n13657), .A2(n7574), .ZN(n13833) );
  AND2_X1 U9071 ( .A1(n13661), .A2(n16090), .ZN(n7574) );
  NAND2_X1 U9072 ( .A1(n9275), .A2(n9274), .ZN(n13697) );
  NAND2_X1 U9073 ( .A1(n9215), .A2(n9214), .ZN(n13922) );
  INV_X1 U9074 ( .A(n13172), .ZN(n13929) );
  NAND2_X1 U9075 ( .A1(n13769), .A2(n9192), .ZN(n13759) );
  AND2_X1 U9076 ( .A1(n7258), .A2(n9411), .ZN(n13768) );
  NAND2_X1 U9077 ( .A1(n7539), .A2(n7543), .ZN(n13798) );
  NAND2_X1 U9078 ( .A1(n12765), .A2(n7545), .ZN(n7539) );
  AOI21_X1 U9079 ( .B1(n12765), .B2(n13325), .A(n13405), .ZN(n13812) );
  NAND2_X1 U9080 ( .A1(n9109), .A2(n9108), .ZN(n13223) );
  NAND2_X1 U9081 ( .A1(n7548), .A2(n7553), .ZN(n12404) );
  NAND2_X1 U9082 ( .A1(n12110), .A2(n7555), .ZN(n7548) );
  INV_X1 U9083 ( .A(n13918), .ZN(n13953) );
  OR2_X1 U9084 ( .A1(n8912), .A2(n6771), .ZN(n8924) );
  INV_X1 U9085 ( .A(n10106), .ZN(n13958) );
  NAND2_X1 U9086 ( .A1(n8799), .A2(P3_STATE_REG_SCAN_IN), .ZN(n13959) );
  XNOR2_X1 U9087 ( .A(n13282), .B(n13281), .ZN(n13967) );
  OAI22_X1 U9088 ( .A1(n13280), .A2(n13279), .B1(P1_DATAO_REG_30__SCAN_IN), 
        .B2(n13278), .ZN(n13282) );
  OAI21_X1 U9089 ( .B1(n9352), .B2(n9351), .A(n13100), .ZN(n13132) );
  NAND2_X1 U9090 ( .A1(n7176), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8904) );
  XNOR2_X1 U9091 ( .A(n9303), .B(n9291), .ZN(n12293) );
  NAND2_X1 U9092 ( .A1(n7580), .A2(n9290), .ZN(n9303) );
  NOR2_X1 U9093 ( .A1(n8704), .A2(n6998), .ZN(n8705) );
  NAND2_X1 U9094 ( .A1(n7610), .A2(n9242), .ZN(n9258) );
  INV_X1 U9095 ( .A(n10104), .ZN(n11750) );
  INV_X1 U9096 ( .A(SI_19_), .ZN(n11461) );
  OAI21_X1 U9097 ( .B1(n7588), .B2(n9181), .A(n6922), .ZN(n9194) );
  NAND2_X1 U9098 ( .A1(n7588), .A2(n7589), .ZN(n9182) );
  NAND2_X1 U9099 ( .A1(n7590), .A2(n9157), .ZN(n9169) );
  NAND2_X1 U9100 ( .A1(n9156), .A2(n9155), .ZN(n7590) );
  INV_X1 U9101 ( .A(SI_14_), .ZN(n11128) );
  INV_X1 U9102 ( .A(n8770), .ZN(n8768) );
  INV_X1 U9103 ( .A(SI_12_), .ZN(n10744) );
  INV_X1 U9104 ( .A(SI_11_), .ZN(n10683) );
  NAND2_X1 U9105 ( .A1(n9044), .A2(n9043), .ZN(n9057) );
  NAND2_X1 U9106 ( .A1(n8999), .A2(n8998), .ZN(n9002) );
  NAND2_X1 U9107 ( .A1(n7584), .A2(n8958), .ZN(n8995) );
  NAND2_X1 U9108 ( .A1(n8972), .A2(n8971), .ZN(n7584) );
  NAND2_X1 U9109 ( .A1(n8738), .A2(n8737), .ZN(n8739) );
  NAND2_X1 U9110 ( .A1(n6770), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8737) );
  OAI21_X1 U9111 ( .B1(n12298), .B2(n7775), .A(n7772), .ZN(n12820) );
  INV_X1 U9112 ( .A(n14877), .ZN(n7907) );
  AND2_X1 U9113 ( .A1(n14010), .A2(n10519), .ZN(n6974) );
  AND2_X1 U9114 ( .A1(n14055), .A2(n10519), .ZN(n14011) );
  NAND2_X1 U9115 ( .A1(n14046), .A2(n10539), .ZN(n14019) );
  AND2_X1 U9116 ( .A1(n10545), .A2(n10544), .ZN(n14018) );
  NAND2_X1 U9117 ( .A1(n8127), .A2(n8126), .ZN(n15983) );
  NAND2_X1 U9118 ( .A1(n14048), .A2(n14047), .ZN(n14046) );
  NAND2_X1 U9119 ( .A1(n6970), .A2(n10442), .ZN(n11616) );
  NAND2_X1 U9120 ( .A1(n12427), .A2(n12428), .ZN(n12426) );
  NAND2_X1 U9121 ( .A1(n12298), .A2(n10464), .ZN(n12427) );
  AND2_X1 U9122 ( .A1(n11906), .A2(n10428), .ZN(n7985) );
  INV_X1 U9123 ( .A(n13111), .ZN(n14733) );
  NAND2_X1 U9124 ( .A1(n7280), .A2(n14001), .ZN(n14057) );
  NAND2_X1 U9125 ( .A1(n12889), .A2(n10484), .ZN(n13974) );
  NAND2_X1 U9126 ( .A1(n6971), .A2(n6656), .ZN(n12870) );
  NAND2_X1 U9127 ( .A1(n12298), .A2(n7770), .ZN(n6971) );
  OR2_X1 U9128 ( .A1(n10472), .A2(n10471), .ZN(n7767) );
  NAND2_X1 U9129 ( .A1(n8219), .A2(n8218), .ZN(n14171) );
  INV_X1 U9130 ( .A(n14090), .ZN(n14097) );
  XNOR2_X1 U9131 ( .A(n10511), .B(n10510), .ZN(n14074) );
  NAND2_X1 U9132 ( .A1(n14038), .A2(n10509), .ZN(n14075) );
  NAND2_X1 U9133 ( .A1(n11739), .A2(n10449), .ZN(n11762) );
  AND2_X1 U9134 ( .A1(n11356), .A2(P2_STATE_REG_SCAN_IN), .ZN(n14088) );
  AOI21_X1 U9135 ( .B1(n6963), .B2(n6965), .A(n6962), .ZN(n6961) );
  INV_X1 U9136 ( .A(n14254), .ZN(n14399) );
  OR2_X1 U9137 ( .A1(n8557), .A2(n8109), .ZN(n8110) );
  NAND4_X1 U9138 ( .A1(n8061), .A2(n8060), .A3(n8059), .A4(n8058), .ZN(n14419)
         );
  NAND4_X1 U9139 ( .A1(n8045), .A2(n8044), .A3(n8043), .A4(n8042), .ZN(n14420)
         );
  NAND2_X1 U9140 ( .A1(n8056), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n8044) );
  NAND2_X1 U9141 ( .A1(n8056), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n8028) );
  NAND2_X1 U9142 ( .A1(n8071), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n8027) );
  NAND2_X1 U9143 ( .A1(n8554), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n8013) );
  AND3_X1 U9144 ( .A1(n8012), .A2(n8010), .A3(n8011), .ZN(n7075) );
  NAND2_X1 U9145 ( .A1(n11164), .A2(n11163), .ZN(n14454) );
  NAND2_X1 U9146 ( .A1(n15922), .A2(n15923), .ZN(n15921) );
  NAND2_X1 U9147 ( .A1(n14487), .A2(n14486), .ZN(n11172) );
  OR2_X1 U9148 ( .A1(n11144), .A2(n11145), .ZN(n11223) );
  NAND2_X1 U9149 ( .A1(n11213), .A2(n11212), .ZN(n11237) );
  OR2_X1 U9150 ( .A1(n11520), .A2(n11521), .ZN(n11721) );
  NAND2_X1 U9151 ( .A1(n11728), .A2(n11727), .ZN(n11732) );
  XNOR2_X1 U9152 ( .A(n11987), .B(n11926), .ZN(n11986) );
  NAND2_X1 U9153 ( .A1(n15940), .A2(n15939), .ZN(n15938) );
  NAND2_X1 U9154 ( .A1(n6873), .A2(n6877), .ZN(n12796) );
  OR2_X1 U9155 ( .A1(n15940), .A2(n6879), .ZN(n6873) );
  INV_X1 U9156 ( .A(n14504), .ZN(n15937) );
  AND2_X1 U9157 ( .A1(n8552), .A2(n10402), .ZN(n14517) );
  XNOR2_X1 U9158 ( .A(n6823), .B(n14545), .ZN(n14757) );
  NAND2_X1 U9159 ( .A1(n6816), .A2(n8469), .ZN(n14578) );
  NAND2_X1 U9160 ( .A1(n14605), .A2(n7683), .ZN(n7678) );
  NAND2_X1 U9161 ( .A1(n14607), .A2(n8634), .ZN(n14584) );
  NAND2_X1 U9162 ( .A1(n8444), .A2(n8443), .ZN(n14600) );
  NAND2_X1 U9163 ( .A1(n7632), .A2(n8402), .ZN(n14627) );
  AND2_X1 U9164 ( .A1(n7672), .A2(n6573), .ZN(n14656) );
  INV_X1 U9165 ( .A(n8628), .ZN(n14667) );
  NAND2_X1 U9166 ( .A1(n8619), .A2(n8618), .ZN(n14727) );
  NAND2_X1 U9167 ( .A1(n7633), .A2(n7638), .ZN(n12752) );
  NAND2_X1 U9168 ( .A1(n8228), .A2(n6616), .ZN(n7633) );
  NAND2_X1 U9169 ( .A1(n12457), .A2(n14344), .ZN(n12459) );
  NAND2_X1 U9170 ( .A1(n12376), .A2(n8191), .ZN(n12457) );
  NAND2_X1 U9171 ( .A1(n7673), .A2(n8600), .ZN(n12234) );
  INV_X1 U9172 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n7118) );
  AND2_X2 U9173 ( .A1(n11634), .A2(n10395), .ZN(n16011) );
  AND2_X1 U9174 ( .A1(n14744), .A2(n15996), .ZN(n7177) );
  AND2_X1 U9175 ( .A1(n14529), .A2(n6999), .ZN(n14854) );
  NOR2_X1 U9176 ( .A1(n14753), .A2(n7000), .ZN(n6999) );
  INV_X1 U9177 ( .A(n14528), .ZN(n7000) );
  OR2_X1 U9178 ( .A1(n14761), .A2(n6820), .ZN(n14856) );
  NAND2_X1 U9179 ( .A1(n6822), .A2(n6821), .ZN(n6820) );
  INV_X1 U9180 ( .A(n14760), .ZN(n6821) );
  NAND2_X1 U9181 ( .A1(n14757), .A2(n15993), .ZN(n6822) );
  INV_X1 U9182 ( .A(n14600), .ZN(n14865) );
  INV_X1 U9183 ( .A(n14171), .ZN(n14893) );
  NAND2_X1 U9184 ( .A1(n7193), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n7192) );
  NAND2_X1 U9185 ( .A1(n13125), .A2(n10637), .ZN(n6827) );
  AND2_X2 U9186 ( .A1(n8038), .A2(n7184), .ZN(n8039) );
  NAND2_X1 U9187 ( .A1(n8062), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n8038) );
  OAI21_X1 U9188 ( .B1(n8420), .B2(n10751), .A(n8037), .ZN(n7185) );
  MUX2_X1 U9190 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8007), .S(
        P2_IR_REG_29__SCAN_IN), .Z(n7615) );
  INV_X1 U9191 ( .A(n8683), .ZN(n14918) );
  XNOR2_X1 U9192 ( .A(n8660), .B(n8659), .ZN(n12582) );
  AND2_X1 U9193 ( .A1(n8574), .A2(P2_IR_REG_22__SCAN_IN), .ZN(n8583) );
  NAND2_X1 U9194 ( .A1(n8580), .A2(n8579), .ZN(n8581) );
  AND2_X1 U9195 ( .A1(n8455), .A2(n8454), .ZN(n12354) );
  INV_X1 U9196 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n11972) );
  INV_X1 U9197 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n11664) );
  INV_X1 U9198 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n11587) );
  INV_X1 U9199 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n11381) );
  INV_X1 U9200 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n11259) );
  INV_X1 U9201 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n11058) );
  INV_X1 U9202 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n11041) );
  AND2_X1 U9203 ( .A1(n8198), .A2(n8235), .ZN(n11238) );
  INV_X1 U9204 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n10749) );
  INV_X1 U9205 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n10713) );
  INV_X1 U9206 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n10964) );
  INV_X1 U9207 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n10707) );
  INV_X1 U9208 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n10699) );
  INV_X1 U9209 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n10710) );
  XNOR2_X1 U9210 ( .A(n6892), .B(P2_IR_REG_4__SCAN_IN), .ZN(n14440) );
  OAI21_X1 U9211 ( .B1(n8077), .B2(P2_IR_REG_3__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n6892) );
  INV_X1 U9212 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n10703) );
  INV_X1 U9213 ( .A(n7056), .ZN(n7936) );
  OAI21_X1 U9214 ( .B1(n7941), .B2(n12179), .A(n10187), .ZN(n7056) );
  AND2_X1 U9215 ( .A1(n9919), .A2(n9918), .ZN(n14927) );
  CLKBUF_X1 U9216 ( .A(n15559), .Z(n7122) );
  INV_X1 U9217 ( .A(n15501), .ZN(n14993) );
  NAND2_X1 U9218 ( .A1(n15031), .A2(n10243), .ZN(n14933) );
  NAND2_X1 U9219 ( .A1(n9845), .A2(n9844), .ZN(n15586) );
  AOI21_X1 U9220 ( .B1(n7964), .B2(n12410), .A(n6671), .ZN(n7963) );
  NAND2_X1 U9221 ( .A1(n14951), .A2(n14950), .ZN(n14949) );
  INV_X1 U9222 ( .A(n15094), .ZN(n12413) );
  CLKBUF_X1 U9223 ( .A(n12409), .Z(n7200) );
  AOI22_X1 U9224 ( .A1(n9513), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n9781), .B2(
        n11097), .ZN(n9559) );
  NAND2_X1 U9225 ( .A1(n15040), .A2(n7029), .ZN(n7023) );
  AND2_X1 U9226 ( .A1(n12407), .A2(n10205), .ZN(n12512) );
  AND2_X1 U9227 ( .A1(n7044), .A2(n15020), .ZN(n7043) );
  OR2_X1 U9228 ( .A1(n14950), .A2(n7045), .ZN(n7044) );
  INV_X1 U9229 ( .A(n10292), .ZN(n7045) );
  NAND2_X1 U9230 ( .A1(n14949), .A2(n10292), .ZN(n15021) );
  INV_X1 U9231 ( .A(n15091), .ZN(n15517) );
  NAND2_X1 U9232 ( .A1(n14957), .A2(n10303), .ZN(n15041) );
  NAND2_X1 U9233 ( .A1(n12740), .A2(n10220), .ZN(n12900) );
  NAND2_X1 U9234 ( .A1(n9524), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n9489) );
  INV_X1 U9235 ( .A(n7941), .ZN(n7938) );
  NAND2_X1 U9236 ( .A1(n7155), .A2(n10179), .ZN(n7939) );
  AND2_X1 U9237 ( .A1(n6830), .A2(n9866), .ZN(n15066) );
  OR2_X1 U9238 ( .A1(n13060), .A2(n6550), .ZN(n6830) );
  AOI21_X1 U9239 ( .B1(n7030), .B2(n7950), .A(n7158), .ZN(n7135) );
  INV_X1 U9240 ( .A(n7954), .ZN(n7158) );
  OAI21_X1 U9241 ( .B1(n15040), .B2(n7026), .A(n7024), .ZN(n7030) );
  INV_X1 U9242 ( .A(n7027), .ZN(n7026) );
  INV_X1 U9243 ( .A(n15060), .ZN(n7134) );
  INV_X1 U9244 ( .A(n15705), .ZN(n10353) );
  INV_X1 U9245 ( .A(n15066), .ZN(n15297) );
  NAND2_X1 U9246 ( .A1(n9876), .A2(n9875), .ZN(n15086) );
  INV_X1 U9247 ( .A(n15391), .ZN(n15087) );
  NAND2_X1 U9248 ( .A1(n9822), .A2(n9821), .ZN(n15421) );
  INV_X1 U9249 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n10729) );
  XNOR2_X1 U9250 ( .A(n6872), .B(P1_IR_REG_1__SCAN_IN), .ZN(n15103) );
  NAND2_X1 U9251 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), .ZN(
        n6872) );
  NAND2_X1 U9252 ( .A1(n11090), .A2(n11089), .ZN(n11197) );
  NAND2_X1 U9253 ( .A1(n11195), .A2(n11092), .ZN(n15168) );
  NAND2_X1 U9254 ( .A1(n15168), .A2(n15169), .ZN(n15167) );
  AOI21_X1 U9255 ( .B1(n11361), .B2(n11360), .A(n11359), .ZN(n15175) );
  NAND2_X1 U9256 ( .A1(n15175), .A2(n15174), .ZN(n15173) );
  NAND2_X1 U9257 ( .A1(n11891), .A2(n11890), .ZN(n11893) );
  NAND2_X1 U9258 ( .A1(n6864), .A2(n12635), .ZN(n12637) );
  AND2_X1 U9259 ( .A1(n6867), .A2(n15235), .ZN(n15219) );
  NAND2_X1 U9260 ( .A1(n6869), .A2(n6868), .ZN(n6867) );
  INV_X1 U9261 ( .A(n15217), .ZN(n6869) );
  NAND2_X1 U9262 ( .A1(n15219), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n15236) );
  OAI21_X1 U9263 ( .B1(n15249), .B2(n15248), .A(n6675), .ZN(n6857) );
  OAI21_X1 U9264 ( .B1(n15252), .B2(n8014), .A(n15251), .ZN(n6856) );
  NAND2_X1 U9265 ( .A1(n10008), .A2(n10007), .ZN(n15258) );
  INV_X1 U9266 ( .A(n13076), .ZN(n15547) );
  OAI21_X1 U9267 ( .B1(n7344), .B2(n15295), .A(n7342), .ZN(n7061) );
  AOI21_X1 U9268 ( .B1(n7345), .B2(n7347), .A(n7343), .ZN(n7342) );
  NAND2_X1 U9269 ( .A1(n9878), .A2(n9877), .ZN(n15301) );
  NAND2_X1 U9270 ( .A1(n15329), .A2(n13020), .ZN(n15310) );
  NOR2_X1 U9271 ( .A1(n15325), .A2(n6665), .ZN(n15307) );
  AND2_X1 U9272 ( .A1(n15335), .A2(n15334), .ZN(n15582) );
  NAND2_X1 U9273 ( .A1(n13042), .A2(n13041), .ZN(n15360) );
  AND2_X1 U9274 ( .A1(n7819), .A2(n6638), .ZN(n15405) );
  NAND2_X1 U9275 ( .A1(n13038), .A2(n13037), .ZN(n15417) );
  NAND2_X1 U9276 ( .A1(n13011), .A2(n13010), .ZN(n15415) );
  NAND2_X1 U9277 ( .A1(n7825), .A2(n13034), .ZN(n15451) );
  NAND2_X1 U9278 ( .A1(n15466), .A2(n13006), .ZN(n15449) );
  NAND2_X1 U9279 ( .A1(n15518), .A2(n13026), .ZN(n6884) );
  CLKBUF_X1 U9280 ( .A(n15518), .Z(n15519) );
  INV_X1 U9281 ( .A(n15526), .ZN(n12568) );
  NAND2_X1 U9282 ( .A1(n7810), .A2(n12555), .ZN(n13024) );
  NAND2_X1 U9283 ( .A1(n12362), .A2(n7813), .ZN(n7810) );
  INV_X1 U9284 ( .A(n7814), .ZN(n7813) );
  NAND2_X1 U9285 ( .A1(n12216), .A2(n7787), .ZN(n12358) );
  NAND2_X1 U9286 ( .A1(n12336), .A2(n12337), .ZN(n7787) );
  OAI21_X1 U9287 ( .B1(n12196), .B2(n7337), .A(n6901), .ZN(n12338) );
  INV_X1 U9288 ( .A(n7336), .ZN(n6901) );
  NAND2_X1 U9289 ( .A1(n7821), .A2(n12198), .ZN(n15777) );
  NAND2_X1 U9290 ( .A1(n12196), .A2(n12195), .ZN(n7821) );
  NAND2_X1 U9291 ( .A1(n12212), .A2(n12211), .ZN(n7783) );
  INV_X1 U9292 ( .A(n15344), .ZN(n15812) );
  INV_X1 U9293 ( .A(n15807), .ZN(n15496) );
  INV_X1 U9294 ( .A(n15535), .ZN(n15513) );
  OR2_X1 U9295 ( .A1(n15556), .A2(n15874), .ZN(n7138) );
  AND2_X2 U9296 ( .A1(n11828), .A2(n11495), .ZN(n15877) );
  AND2_X1 U9297 ( .A1(n10718), .A2(P1_STATE_REG_SCAN_IN), .ZN(n10687) );
  NAND2_X1 U9298 ( .A1(n10684), .A2(n11467), .ZN(n15821) );
  NAND2_X1 U9299 ( .A1(n7933), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9449) );
  AND2_X1 U9300 ( .A1(n7970), .A2(n6583), .ZN(n7932) );
  BUF_X1 U9301 ( .A(n10073), .Z(n15119) );
  INV_X1 U9302 ( .A(n10356), .ZN(n15704) );
  MUX2_X1 U9303 ( .A(P1_IR_REG_31__SCAN_IN), .B(n10062), .S(
        P1_IR_REG_25__SCAN_IN), .Z(n10064) );
  XNOR2_X1 U9304 ( .A(n9827), .B(P2_DATAO_REG_22__SCAN_IN), .ZN(n15706) );
  NAND2_X1 U9305 ( .A1(n8419), .A2(n8418), .ZN(n12143) );
  NAND2_X1 U9306 ( .A1(n8406), .A2(n8405), .ZN(n8419) );
  NOR2_X1 U9307 ( .A1(n9478), .A2(n9477), .ZN(n9479) );
  NOR2_X1 U9308 ( .A1(n9475), .A2(n9447), .ZN(n7201) );
  NAND2_X1 U9309 ( .A1(n8406), .A2(n8391), .ZN(n12183) );
  INV_X1 U9310 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n11971) );
  INV_X1 U9311 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n11669) );
  XNOR2_X1 U9312 ( .A(n9698), .B(P1_IR_REG_14__SCAN_IN), .ZN(n15191) );
  INV_X1 U9313 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n11383) );
  INV_X1 U9314 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n11061) );
  INV_X1 U9315 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n11038) );
  INV_X1 U9316 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n10747) );
  INV_X1 U9317 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n10716) );
  XNOR2_X1 U9318 ( .A(n10679), .B(n10650), .ZN(n10651) );
  XNOR2_X1 U9319 ( .A(n11045), .B(n11044), .ZN(n11043) );
  XNOR2_X1 U9320 ( .A(n11339), .B(P2_ADDR_REG_6__SCAN_IN), .ZN(n11053) );
  NAND2_X1 U9321 ( .A1(n12005), .A2(n12004), .ZN(n12324) );
  NOR2_X1 U9322 ( .A1(n12333), .A2(n12332), .ZN(n12334) );
  AOI21_X1 U9323 ( .B1(n7509), .B2(n7508), .A(n6623), .ZN(n15720) );
  NAND2_X1 U9324 ( .A1(n15710), .A2(P2_ADDR_REG_13__SCAN_IN), .ZN(n7508) );
  INV_X1 U9325 ( .A(n15738), .ZN(n6851) );
  OR2_X1 U9326 ( .A1(n7506), .A2(n7504), .ZN(n7503) );
  AOI21_X1 U9327 ( .B1(n7124), .B2(n15750), .A(n7123), .ZN(n6848) );
  NAND2_X1 U9328 ( .A1(n7465), .A2(n13243), .ZN(n7464) );
  NAND2_X1 U9329 ( .A1(n11653), .A2(n11652), .ZN(n11657) );
  XNOR2_X1 U9330 ( .A(n6781), .B(n7109), .ZN(n13263) );
  OR2_X1 U9331 ( .A1(n13489), .A2(n13488), .ZN(n7372) );
  NAND2_X1 U9332 ( .A1(n7659), .A2(n13548), .ZN(n13531) );
  OAI21_X1 U9333 ( .B1(n6918), .B2(n16103), .A(n6600), .ZN(n13831) );
  OAI21_X1 U9334 ( .B1(n13833), .B2(n16103), .A(n7571), .ZN(P3_U3486) );
  NOR2_X1 U9335 ( .A1(n7573), .A2(n7572), .ZN(n7571) );
  NOR2_X1 U9336 ( .A1(n16106), .A2(n13834), .ZN(n7572) );
  NOR2_X1 U9337 ( .A1(n13835), .A2(n13860), .ZN(n7573) );
  NAND2_X1 U9338 ( .A1(n6918), .A2(n16094), .ZN(n10586) );
  OAI22_X1 U9339 ( .A1(n13832), .A2(n13918), .B1(n16094), .B2(n10583), .ZN(
        n10584) );
  NOR2_X1 U9340 ( .A1(n11150), .A2(n10587), .ZN(P2_U3947) );
  AND2_X1 U9341 ( .A1(n14083), .A2(n7747), .ZN(n13124) );
  AND2_X1 U9342 ( .A1(n13123), .A2(n7745), .ZN(n7744) );
  NAND2_X1 U9343 ( .A1(n14083), .A2(n6642), .ZN(n7748) );
  AND2_X1 U9344 ( .A1(n14388), .A2(n14389), .ZN(n7091) );
  NAND2_X1 U9345 ( .A1(n14325), .A2(n7093), .ZN(n7092) );
  AOI21_X1 U9346 ( .B1(n15899), .B2(P2_ADDR_REG_19__SCAN_IN), .A(n14506), .ZN(
        n6898) );
  NAND2_X1 U9347 ( .A1(n6897), .A2(n8584), .ZN(n6896) );
  NAND2_X1 U9348 ( .A1(n6900), .A2(n14322), .ZN(n6899) );
  NAND2_X1 U9349 ( .A1(n14529), .A2(n14528), .ZN(n14754) );
  NAND2_X1 U9350 ( .A1(n7119), .A2(n7116), .ZN(P2_U3530) );
  INV_X1 U9351 ( .A(n7117), .ZN(n7116) );
  OAI22_X1 U9352 ( .A1(n14849), .A2(n14840), .B1(n16011), .B2(n7118), .ZN(
        n7117) );
  MUX2_X1 U9353 ( .A(P2_REG1_REG_30__SCAN_IN), .B(n12996), .S(n16011), .Z(
        n12997) );
  OAI21_X1 U9354 ( .B1(n14847), .B2(n16002), .A(n7111), .ZN(n14848) );
  NAND2_X1 U9355 ( .A1(n16002), .A2(n7112), .ZN(n7111) );
  INV_X1 U9356 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n7112) );
  MUX2_X1 U9357 ( .A(n12996), .B(P2_REG0_REG_30__SCAN_IN), .S(n16002), .Z(
        n12994) );
  OAI21_X1 U9358 ( .B1(n14851), .B2(n16002), .A(n7181), .ZN(P2_U3495) );
  NOR2_X1 U9359 ( .A1(n6662), .A2(n7182), .ZN(n7181) );
  NOR2_X1 U9360 ( .A1(n16004), .A2(n14852), .ZN(n7182) );
  NAND2_X1 U9361 ( .A1(n7002), .A2(n7001), .ZN(P2_U3494) );
  OR2_X1 U9362 ( .A1(n16004), .A2(n14855), .ZN(n7001) );
  OR2_X1 U9363 ( .A1(n14854), .A2(n16002), .ZN(n7002) );
  CLKBUF_X1 U9364 ( .A(n6547), .Z(P1_U4016) );
  OAI22_X1 U9365 ( .A1(n15065), .A2(n11956), .B1(n11476), .B2(n15056), .ZN(
        n11487) );
  XNOR2_X1 U9366 ( .A(n14979), .B(n7157), .ZN(n7156) );
  NAND2_X1 U9367 ( .A1(n6858), .A2(n6855), .ZN(P1_U3262) );
  NAND2_X1 U9368 ( .A1(n6859), .A2(n9780), .ZN(n6858) );
  AOI21_X1 U9369 ( .B1(n6857), .B2(n15250), .A(n6856), .ZN(n6855) );
  OAI22_X1 U9370 ( .A1(n15243), .A2(n15248), .B1(n15245), .B2(n15242), .ZN(
        n6859) );
  NAND2_X1 U9371 ( .A1(n7103), .A2(n7102), .ZN(P1_U3559) );
  NAND2_X1 U9372 ( .A1(n15884), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n7102) );
  NAND2_X1 U9373 ( .A1(n15666), .A2(n15886), .ZN(n7103) );
  NAND2_X1 U9374 ( .A1(n15884), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n7202) );
  NAND2_X1 U9375 ( .A1(n6895), .A2(n6894), .ZN(P1_U3556) );
  NAND2_X1 U9376 ( .A1(n15884), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n6894) );
  NAND2_X1 U9377 ( .A1(n15669), .A2(n15886), .ZN(n6895) );
  NAND2_X1 U9378 ( .A1(n15884), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n7151) );
  NAND2_X1 U9379 ( .A1(n6791), .A2(n6731), .ZN(P1_U3527) );
  NAND2_X1 U9380 ( .A1(n15666), .A2(n15877), .ZN(n6791) );
  INV_X1 U9381 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n6790) );
  INV_X1 U9382 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n7451) );
  INV_X1 U9383 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n7097) );
  NAND2_X1 U9384 ( .A1(n6837), .A2(n6836), .ZN(n11941) );
  INV_X1 U9385 ( .A(n6838), .ZN(n6837) );
  INV_X2 U9386 ( .A(n9651), .ZN(n9635) );
  INV_X1 U9387 ( .A(n14148), .ZN(n7900) );
  NAND3_X2 U9388 ( .A1(n7516), .A2(n14383), .A3(n14379), .ZN(n14265) );
  NAND2_X1 U9389 ( .A1(n13452), .A2(n6946), .ZN(n6570) );
  NAND2_X2 U9390 ( .A1(n8906), .A2(n8907), .ZN(n9126) );
  AND2_X1 U9391 ( .A1(n7967), .A2(n12198), .ZN(n6571) );
  AND2_X1 U9392 ( .A1(n15444), .A2(n15459), .ZN(n6572) );
  OR2_X1 U9393 ( .A1(n14800), .A2(n8626), .ZN(n6573) );
  AND2_X1 U9394 ( .A1(n8619), .A2(n7690), .ZN(n6574) );
  AND2_X1 U9395 ( .A1(n7291), .A2(n10545), .ZN(n6575) );
  AND3_X1 U9396 ( .A1(n13120), .A2(n14065), .A3(n13119), .ZN(n6576) );
  INV_X1 U9397 ( .A(n10589), .ZN(n7658) );
  AND2_X1 U9398 ( .A1(n9606), .A2(n7913), .ZN(n6577) );
  OR2_X1 U9399 ( .A1(n13087), .A2(n15297), .ZN(n6578) );
  AND2_X1 U9400 ( .A1(n7732), .A2(P3_REG1_REG_7__SCAN_IN), .ZN(n6579) );
  NAND2_X1 U9401 ( .A1(n13390), .A2(n13389), .ZN(n6580) );
  AND2_X1 U9402 ( .A1(n7178), .A2(n14865), .ZN(n6581) );
  INV_X1 U9403 ( .A(n7320), .ZN(n7317) );
  NOR3_X1 U9404 ( .A1(n13942), .A2(n13818), .A3(n13450), .ZN(n6582) );
  INV_X1 U9405 ( .A(n7570), .ZN(n8713) );
  INV_X1 U9406 ( .A(n13383), .ZN(n7556) );
  AND2_X1 U9407 ( .A1(n9444), .A2(n9458), .ZN(n6583) );
  INV_X1 U9408 ( .A(n14037), .ZN(n10508) );
  AND2_X1 U9409 ( .A1(n14320), .A2(n14319), .ZN(n6584) );
  AND2_X1 U9410 ( .A1(n7042), .A2(n8637), .ZN(n6585) );
  NOR2_X1 U9411 ( .A1(n7684), .A2(n8635), .ZN(n7682) );
  AND2_X1 U9412 ( .A1(n6813), .A2(n8196), .ZN(n6586) );
  NAND2_X1 U9413 ( .A1(n8273), .A2(n7275), .ZN(n7274) );
  AND2_X1 U9414 ( .A1(n12766), .A2(n9136), .ZN(n6587) );
  AND2_X1 U9415 ( .A1(n6843), .A2(n10626), .ZN(n6588) );
  NAND2_X1 U9416 ( .A1(n11703), .A2(P3_REG1_REG_8__SCAN_IN), .ZN(n7731) );
  OR2_X1 U9417 ( .A1(n7159), .A2(n13482), .ZN(n6589) );
  AND2_X1 U9418 ( .A1(n13411), .A2(n13450), .ZN(n6590) );
  XNOR2_X1 U9419 ( .A(n10527), .B(n10525), .ZN(n13988) );
  AND2_X1 U9420 ( .A1(n13398), .A2(n13397), .ZN(n6591) );
  AND2_X1 U9421 ( .A1(n6691), .A2(n13422), .ZN(n6592) );
  NAND2_X1 U9422 ( .A1(n7440), .A2(n13537), .ZN(n6593) );
  INV_X1 U9423 ( .A(n9673), .ZN(n7916) );
  INV_X1 U9424 ( .A(n9636), .ZN(n7910) );
  INV_X1 U9425 ( .A(n14169), .ZN(n7533) );
  NOR2_X1 U9426 ( .A1(n15764), .A2(P2_ADDR_REG_17__SCAN_IN), .ZN(n6594) );
  NOR2_X1 U9427 ( .A1(n13524), .A2(n8878), .ZN(n6595) );
  AND2_X1 U9428 ( .A1(n10391), .A2(n8561), .ZN(n14362) );
  INV_X1 U9429 ( .A(n14362), .ZN(n7693) );
  INV_X1 U9430 ( .A(n8192), .ZN(n8193) );
  XNOR2_X1 U9431 ( .A(n8195), .B(SI_9_), .ZN(n8192) );
  AND2_X1 U9432 ( .A1(n13426), .A2(n9180), .ZN(n6596) );
  AND2_X1 U9433 ( .A1(n10463), .A2(n10457), .ZN(n6597) );
  XOR2_X1 U9434 ( .A(n13206), .B(n13683), .Z(n6598) );
  NOR2_X1 U9435 ( .A1(n8541), .A2(SI_27_), .ZN(n6599) );
  OR2_X1 U9436 ( .A1(n16106), .A2(P3_REG1_REG_28__SCAN_IN), .ZN(n6600) );
  NAND2_X1 U9437 ( .A1(n9273), .A2(n9272), .ZN(n13722) );
  INV_X1 U9438 ( .A(n13722), .ZN(n13444) );
  AND2_X1 U9439 ( .A1(n12333), .A2(n12332), .ZN(n6601) );
  NAND2_X1 U9440 ( .A1(n14730), .A2(n14176), .ZN(n14731) );
  INV_X1 U9441 ( .A(n14731), .ZN(n7115) );
  AND2_X1 U9442 ( .A1(n7467), .A2(n6718), .ZN(n6602) );
  AND2_X1 U9443 ( .A1(n8891), .A2(n13616), .ZN(n6603) );
  OAI21_X1 U9444 ( .B1(n9383), .B2(P3_D_REG_0__SCAN_IN), .A(n9382), .ZN(n11430) );
  OR2_X1 U9445 ( .A1(n12225), .A2(n7899), .ZN(n6604) );
  AND2_X1 U9446 ( .A1(n7449), .A2(n15792), .ZN(n6605) );
  AND2_X1 U9447 ( .A1(n14913), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n6606) );
  INV_X1 U9448 ( .A(n13601), .ZN(n7640) );
  XNOR2_X1 U9449 ( .A(n8790), .B(P3_IR_REG_19__SCAN_IN), .ZN(n13332) );
  INV_X1 U9450 ( .A(n13332), .ZN(n13306) );
  INV_X1 U9451 ( .A(n11324), .ZN(n7405) );
  INV_X1 U9452 ( .A(n9513), .ZN(n9555) );
  INV_X1 U9453 ( .A(n10739), .ZN(n7234) );
  AND2_X1 U9454 ( .A1(n8566), .A2(n8576), .ZN(n14105) );
  NAND2_X1 U9455 ( .A1(n9307), .A2(n9306), .ZN(n13836) );
  NAND2_X1 U9456 ( .A1(n9125), .A2(n9124), .ZN(n13404) );
  INV_X1 U9457 ( .A(n8962), .ZN(n7646) );
  AND2_X1 U9458 ( .A1(n13475), .A2(n13472), .ZN(n6607) );
  NAND2_X1 U9459 ( .A1(n10313), .A2(n10312), .ZN(n6608) );
  NAND2_X1 U9460 ( .A1(n8735), .A2(n8747), .ZN(n10662) );
  NAND2_X1 U9461 ( .A1(n8259), .A2(n8258), .ZN(n14191) );
  INV_X1 U9462 ( .A(n14191), .ZN(n6951) );
  NAND2_X1 U9463 ( .A1(n9293), .A2(n9292), .ZN(n13841) );
  INV_X1 U9464 ( .A(n7749), .ZN(n14027) );
  XNOR2_X1 U9465 ( .A(n14744), .B(n14393), .ZN(n14363) );
  NAND2_X1 U9466 ( .A1(n9230), .A2(n9229), .ZN(n13734) );
  AND2_X1 U9467 ( .A1(n12332), .A2(n7515), .ZN(n6609) );
  NAND2_X1 U9468 ( .A1(n12362), .A2(n12361), .ZN(n12557) );
  NAND2_X1 U9469 ( .A1(n14676), .A2(n14877), .ZN(n14638) );
  AND3_X1 U9470 ( .A1(n7906), .A2(n14676), .A3(n7905), .ZN(n6610) );
  OR2_X1 U9471 ( .A1(n14530), .A2(n14519), .ZN(n6611) );
  INV_X1 U9472 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n8051) );
  AND2_X1 U9473 ( .A1(n6572), .A2(n15471), .ZN(n6612) );
  XNOR2_X1 U9474 ( .A(n15559), .B(n15066), .ZN(n13054) );
  INV_X1 U9475 ( .A(n7347), .ZN(n7346) );
  NAND2_X1 U9476 ( .A1(n12853), .A2(n13503), .ZN(n6613) );
  OR2_X1 U9477 ( .A1(n9187), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n6614) );
  AND2_X1 U9478 ( .A1(n9402), .A2(n13340), .ZN(n6615) );
  NOR2_X1 U9479 ( .A1(n8251), .A2(n7637), .ZN(n6616) );
  AND2_X1 U9480 ( .A1(n13427), .A2(n13428), .ZN(n13758) );
  AND2_X1 U9481 ( .A1(n11312), .A2(P3_REG2_REG_2__SCAN_IN), .ZN(n6617) );
  AND2_X1 U9482 ( .A1(n8213), .A2(SI_10_), .ZN(n6618) );
  AND2_X1 U9483 ( .A1(n10662), .A2(P3_REG2_REG_4__SCAN_IN), .ZN(n6619) );
  AND2_X1 U9484 ( .A1(n10418), .A2(n10417), .ZN(n6620) );
  OR2_X1 U9485 ( .A1(n12913), .A2(n14328), .ZN(n8619) );
  INV_X1 U9486 ( .A(n14379), .ZN(n7741) );
  OR2_X1 U9487 ( .A1(n11146), .A2(n8053), .ZN(n6621) );
  NAND4_X1 U9488 ( .A1(n9530), .A2(n9529), .A3(n9528), .A4(n9527), .ZN(n15099)
         );
  NOR2_X1 U9489 ( .A1(n12901), .A2(n10234), .ZN(n6622) );
  AND2_X1 U9490 ( .A1(n15712), .A2(n15711), .ZN(n6623) );
  XNOR2_X1 U9491 ( .A(n8744), .B(P3_IR_REG_3__SCAN_IN), .ZN(n8981) );
  INV_X1 U9492 ( .A(n8981), .ZN(n7696) );
  NAND2_X1 U9493 ( .A1(n15040), .A2(n10307), .ZN(n14941) );
  AND2_X1 U9494 ( .A1(n6968), .A2(n10501), .ZN(n6624) );
  OR2_X1 U9495 ( .A1(n15336), .A2(n7459), .ZN(n6625) );
  OR2_X1 U9496 ( .A1(n15370), .A2(n15087), .ZN(n6626) );
  AND2_X1 U9497 ( .A1(n8987), .A2(n7326), .ZN(n6627) );
  NAND2_X1 U9498 ( .A1(n7678), .A2(n7681), .ZN(n14568) );
  NAND2_X1 U9499 ( .A1(n10739), .A2(P3_REG1_REG_6__SCAN_IN), .ZN(n6628) );
  OR2_X1 U9500 ( .A1(n7234), .A2(n9012), .ZN(n6629) );
  XOR2_X1 U9501 ( .A(n12253), .B(n13505), .Z(n6630) );
  OR3_X1 U9502 ( .A1(n9989), .A2(n9988), .A3(n9987), .ZN(n6631) );
  AND3_X1 U9503 ( .A1(n6630), .A2(n12472), .A3(n6766), .ZN(n6632) );
  OR2_X1 U9504 ( .A1(n15616), .A2(n15419), .ZN(n6633) );
  INV_X1 U9505 ( .A(n11859), .ZN(n7826) );
  AND2_X1 U9506 ( .A1(n10547), .A2(n10546), .ZN(n6634) );
  AND2_X1 U9507 ( .A1(n13067), .A2(n13066), .ZN(n6635) );
  AND3_X1 U9508 ( .A1(n13298), .A2(n13462), .A3(n13475), .ZN(n6636) );
  XNOR2_X1 U9509 ( .A(n14749), .B(n14395), .ZN(n14536) );
  INV_X1 U9510 ( .A(n14646), .ZN(n7666) );
  INV_X1 U9511 ( .A(n8346), .ZN(n7885) );
  NAND2_X1 U9512 ( .A1(n10508), .A2(n10507), .ZN(n14038) );
  NAND2_X1 U9513 ( .A1(n8457), .A2(n8456), .ZN(n14618) );
  INV_X1 U9514 ( .A(n15093), .ZN(n12904) );
  NAND2_X1 U9515 ( .A1(n15301), .A2(n15086), .ZN(n6637) );
  NAND2_X1 U9516 ( .A1(n15605), .A2(n15433), .ZN(n6638) );
  INV_X1 U9517 ( .A(n7669), .ZN(n7671) );
  INV_X1 U9518 ( .A(n13566), .ZN(n6906) );
  INV_X1 U9519 ( .A(n15341), .ZN(n15578) );
  AND2_X1 U9520 ( .A1(n12230), .A2(n12220), .ZN(n6639) );
  INV_X1 U9521 ( .A(n13365), .ZN(n7565) );
  AND2_X1 U9522 ( .A1(n14218), .A2(n7141), .ZN(n6640) );
  AND2_X1 U9523 ( .A1(n7721), .A2(P3_REG1_REG_5__SCAN_IN), .ZN(n6641) );
  AND2_X1 U9524 ( .A1(n7747), .A2(n13116), .ZN(n6642) );
  AND4_X1 U9525 ( .A1(n9086), .A2(n9085), .A3(n9084), .A4(n9083), .ZN(n12934)
         );
  NOR2_X1 U9526 ( .A1(n14549), .A2(n14266), .ZN(n6643) );
  AND2_X1 U9527 ( .A1(n12735), .A2(n13503), .ZN(n9407) );
  INV_X1 U9528 ( .A(n8253), .ZN(n7285) );
  AND2_X1 U9529 ( .A1(n7021), .A2(n8612), .ZN(n6644) );
  AND2_X1 U9530 ( .A1(n9285), .A2(n9284), .ZN(n13683) );
  AND2_X1 U9531 ( .A1(n14749), .A2(n14264), .ZN(n6645) );
  AND2_X1 U9532 ( .A1(n8511), .A2(n8513), .ZN(n6646) );
  NAND2_X1 U9533 ( .A1(n13053), .A2(n10025), .ZN(n15293) );
  OR2_X1 U9534 ( .A1(n13677), .A2(n13448), .ZN(n6647) );
  AND2_X1 U9535 ( .A1(n6852), .A2(n6851), .ZN(n6648) );
  AND2_X1 U9536 ( .A1(n7693), .A2(n7694), .ZN(n6649) );
  OR2_X1 U9537 ( .A1(n15923), .A2(n6889), .ZN(n6650) );
  AND2_X1 U9538 ( .A1(n14147), .A2(n14146), .ZN(n6651) );
  AND2_X1 U9539 ( .A1(n14769), .A2(n14261), .ZN(n6652) );
  AND2_X1 U9540 ( .A1(n7435), .A2(n7433), .ZN(n6653) );
  AND2_X1 U9541 ( .A1(n9335), .A2(n9318), .ZN(n6654) );
  INV_X1 U9542 ( .A(n9837), .ZN(n6749) );
  OR2_X1 U9543 ( .A1(n14191), .A2(n14409), .ZN(n6655) );
  AND2_X1 U9544 ( .A1(n7768), .A2(n7767), .ZN(n6656) );
  AND2_X1 U9545 ( .A1(n7019), .A2(n8616), .ZN(n6657) );
  AND2_X1 U9546 ( .A1(n13035), .A2(n13034), .ZN(n6658) );
  NOR2_X1 U9547 ( .A1(n7149), .A2(n6776), .ZN(n11499) );
  OR2_X1 U9548 ( .A1(n6628), .A2(n9006), .ZN(n6659) );
  NOR2_X1 U9549 ( .A1(n14151), .A2(n14149), .ZN(n7530) );
  AND2_X1 U9550 ( .A1(n7414), .A2(n12053), .ZN(n6660) );
  OAI21_X1 U9551 ( .B1(n6580), .B2(n7844), .A(n7389), .ZN(n7388) );
  NOR2_X1 U9552 ( .A1(n8385), .A2(n8384), .ZN(n8409) );
  AND2_X1 U9553 ( .A1(n7986), .A2(n9986), .ZN(n6661) );
  OR2_X1 U9554 ( .A1(n15639), .A2(n15517), .ZN(n13030) );
  INV_X1 U9555 ( .A(n13030), .ZN(n6883) );
  INV_X1 U9556 ( .A(n14245), .ZN(n7524) );
  NOR2_X1 U9557 ( .A1(n14853), .A2(n14892), .ZN(n6662) );
  INV_X1 U9558 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n9458) );
  AND2_X1 U9559 ( .A1(n10582), .A2(n10581), .ZN(n6663) );
  INV_X1 U9560 ( .A(n14172), .ZN(n7306) );
  AND2_X1 U9561 ( .A1(n12942), .A2(n13498), .ZN(n6664) );
  AND2_X1 U9562 ( .A1(n15578), .A2(n15306), .ZN(n6665) );
  NAND2_X1 U9563 ( .A1(n14697), .A2(n14405), .ZN(n6666) );
  INV_X1 U9564 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n8578) );
  OR2_X1 U9565 ( .A1(n13506), .A2(n12134), .ZN(n13375) );
  AND2_X1 U9566 ( .A1(n14535), .A2(n8540), .ZN(n6667) );
  AND2_X1 U9567 ( .A1(P1_REG3_REG_7__SCAN_IN), .A2(P1_REG3_REG_8__SCAN_IN), 
        .ZN(n6668) );
  NAND2_X1 U9568 ( .A1(n8482), .A2(n8481), .ZN(n14769) );
  INV_X1 U9569 ( .A(n14769), .ZN(n6952) );
  NOR2_X1 U9570 ( .A1(n8601), .A2(n15995), .ZN(n6669) );
  NOR2_X1 U9571 ( .A1(n15651), .A2(n13025), .ZN(n6670) );
  NOR2_X1 U9572 ( .A1(n10212), .A2(n10211), .ZN(n6671) );
  INV_X1 U9573 ( .A(n8637), .ZN(n7361) );
  AND2_X1 U9574 ( .A1(n8098), .A2(SI_5_), .ZN(n6672) );
  AND4_X2 U9575 ( .A1(n9488), .A2(n9490), .A3(n9489), .A4(n9491), .ZN(n10123)
         );
  INV_X1 U9576 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n8201) );
  INV_X1 U9577 ( .A(n7836), .ZN(n7835) );
  NOR2_X1 U9578 ( .A1(n12936), .A2(n12937), .ZN(n7836) );
  AND2_X1 U9579 ( .A1(n13417), .A2(n9411), .ZN(n13788) );
  INV_X1 U9580 ( .A(n13788), .ZN(n13783) );
  AND2_X1 U9581 ( .A1(n13755), .A2(n13423), .ZN(n13770) );
  INV_X1 U9582 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n12903) );
  OR2_X1 U9583 ( .A1(n10319), .A2(n10318), .ZN(n7955) );
  INV_X1 U9584 ( .A(n7955), .ZN(n7945) );
  INV_X1 U9585 ( .A(n14153), .ZN(n7319) );
  OR2_X1 U9586 ( .A1(n14618), .A2(n14628), .ZN(n6673) );
  NOR2_X1 U9587 ( .A1(n14171), .A2(n14411), .ZN(n6674) );
  AND2_X1 U9588 ( .A1(n14676), .A2(n7178), .ZN(n14595) );
  AND2_X1 U9589 ( .A1(n15247), .A2(n15246), .ZN(n6675) );
  AND2_X1 U9590 ( .A1(n13801), .A2(n9153), .ZN(n13408) );
  INV_X1 U9591 ( .A(n13408), .ZN(n7547) );
  NOR2_X1 U9592 ( .A1(n12976), .A2(n12975), .ZN(n6676) );
  AND2_X1 U9593 ( .A1(n9465), .A2(n7349), .ZN(n10056) );
  AND2_X1 U9594 ( .A1(n11169), .A2(n6650), .ZN(n6677) );
  AND2_X1 U9595 ( .A1(n13929), .A2(n13748), .ZN(n13425) );
  AND2_X1 U9596 ( .A1(n12940), .A2(n13816), .ZN(n6678) );
  AND2_X1 U9597 ( .A1(n13391), .A2(n13392), .ZN(n13390) );
  INV_X1 U9598 ( .A(n13390), .ZN(n7550) );
  AND2_X1 U9599 ( .A1(n13841), .A2(n6947), .ZN(n6679) );
  NAND2_X1 U9600 ( .A1(n8529), .A2(n8511), .ZN(n6793) );
  NAND2_X1 U9601 ( .A1(n10056), .A2(n9443), .ZN(n6680) );
  NOR2_X1 U9602 ( .A1(n10511), .A2(n10510), .ZN(n6681) );
  OR2_X1 U9603 ( .A1(n7885), .A2(n8407), .ZN(n6682) );
  INV_X1 U9604 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n10655) );
  INV_X1 U9605 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n10779) );
  INV_X1 U9606 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n10692) );
  INV_X1 U9607 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n10674) );
  OR2_X1 U9608 ( .A1(n7431), .A2(n7430), .ZN(n6683) );
  INV_X1 U9609 ( .A(n7731), .ZN(n7730) );
  AND2_X1 U9610 ( .A1(n13422), .A2(n13421), .ZN(n6684) );
  NOR2_X1 U9611 ( .A1(n7927), .A2(n7929), .ZN(n6685) );
  AND2_X1 U9612 ( .A1(n13410), .A2(n13415), .ZN(n13797) );
  XNOR2_X1 U9613 ( .A(n8213), .B(SI_10_), .ZN(n8211) );
  AND2_X1 U9614 ( .A1(n10453), .A2(n10452), .ZN(n6686) );
  OR2_X1 U9615 ( .A1(n13480), .A2(n16057), .ZN(n6687) );
  INV_X1 U9616 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n9106) );
  INV_X1 U9617 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n10820) );
  INV_X1 U9618 ( .A(n13065), .ZN(n15269) );
  AND2_X1 U9619 ( .A1(n6745), .A2(n6744), .ZN(n6688) );
  AND2_X1 U9620 ( .A1(n6591), .A2(n7387), .ZN(n6689) );
  AND2_X1 U9621 ( .A1(n7725), .A2(n8867), .ZN(n6690) );
  OR2_X1 U9622 ( .A1(n13425), .A2(n13424), .ZN(n6691) );
  NAND2_X1 U9623 ( .A1(n8084), .A2(n8083), .ZN(n14136) );
  AND2_X1 U9624 ( .A1(n9411), .A2(n13770), .ZN(n7257) );
  INV_X1 U9625 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n8005) );
  INV_X1 U9626 ( .A(n6571), .ZN(n7337) );
  INV_X1 U9627 ( .A(n9569), .ZN(n7923) );
  OR2_X1 U9628 ( .A1(n14536), .A2(n7619), .ZN(n7618) );
  NAND2_X1 U9629 ( .A1(n13379), .A2(n13378), .ZN(n13373) );
  INV_X1 U9630 ( .A(n13373), .ZN(n7251) );
  AND3_X1 U9631 ( .A1(n8564), .A2(n8568), .A3(n8567), .ZN(n6692) );
  NOR2_X1 U9632 ( .A1(n15662), .A2(n15094), .ZN(n6693) );
  OR2_X1 U9633 ( .A1(n13456), .A2(n13455), .ZN(n13668) );
  INV_X1 U9634 ( .A(n13668), .ZN(n13665) );
  NAND2_X1 U9635 ( .A1(n8782), .A2(n11126), .ZN(n13588) );
  INV_X1 U9636 ( .A(n13588), .ZN(n6991) );
  INV_X1 U9637 ( .A(n12213), .ZN(n7784) );
  AND2_X1 U9638 ( .A1(n13462), .A2(n9413), .ZN(n13469) );
  INV_X1 U9639 ( .A(n13469), .ZN(n7215) );
  AND2_X1 U9640 ( .A1(n6993), .A2(n13588), .ZN(n6694) );
  AND2_X1 U9641 ( .A1(n7816), .A2(n13057), .ZN(n6695) );
  AND2_X1 U9642 ( .A1(n13343), .A2(n13450), .ZN(n6696) );
  AND2_X1 U9643 ( .A1(n13893), .A2(n13491), .ZN(n13474) );
  INV_X1 U9644 ( .A(n13474), .ZN(n7329) );
  NOR2_X1 U9645 ( .A1(n14298), .A2(n14297), .ZN(n6697) );
  AND4_X2 U9646 ( .A1(n9494), .A2(n9495), .A3(n9496), .A4(n9493), .ZN(n11476)
         );
  INV_X1 U9647 ( .A(n12999), .ZN(n7796) );
  AND2_X1 U9648 ( .A1(n13665), .A2(n13454), .ZN(n6698) );
  INV_X1 U9649 ( .A(n13006), .ZN(n7071) );
  AND2_X1 U9650 ( .A1(n8005), .A2(n7309), .ZN(n6699) );
  INV_X1 U9651 ( .A(n8634), .ZN(n7686) );
  AND2_X1 U9652 ( .A1(n9302), .A2(n9301), .ZN(n13209) );
  INV_X1 U9653 ( .A(n13209), .ZN(n6947) );
  AND2_X1 U9654 ( .A1(n7911), .A2(n9621), .ZN(n6700) );
  OR2_X1 U9655 ( .A1(n14139), .A2(n14137), .ZN(n6701) );
  AND2_X1 U9656 ( .A1(n6622), .A2(n10220), .ZN(n6702) );
  AND2_X1 U9657 ( .A1(n7100), .A2(n13629), .ZN(n6703) );
  AND2_X1 U9658 ( .A1(n13341), .A2(n6615), .ZN(n6704) );
  OR2_X1 U9659 ( .A1(n14168), .A2(n7533), .ZN(n6705) );
  OR2_X1 U9660 ( .A1(n13026), .A2(n6885), .ZN(n6706) );
  INV_X1 U9661 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n9448) );
  AND2_X1 U9662 ( .A1(n7776), .A2(n8578), .ZN(n6707) );
  INV_X1 U9663 ( .A(n8625), .ZN(n8627) );
  INV_X1 U9664 ( .A(P3_IR_REG_29__SCAN_IN), .ZN(n8903) );
  AND2_X1 U9665 ( .A1(n7597), .A2(n6607), .ZN(n6708) );
  AND2_X1 U9666 ( .A1(n12511), .A2(n10205), .ZN(n7964) );
  AND2_X1 U9667 ( .A1(n6689), .A2(n7385), .ZN(n6709) );
  INV_X1 U9668 ( .A(n10485), .ZN(n7272) );
  INV_X1 U9669 ( .A(P3_IR_REG_28__SCAN_IN), .ZN(n8805) );
  NAND2_X1 U9670 ( .A1(n9637), .A2(n7910), .ZN(n6710) );
  OR2_X1 U9671 ( .A1(P1_IR_REG_27__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), .ZN(
        n6711) );
  INV_X1 U9672 ( .A(P3_IR_REG_2__SCAN_IN), .ZN(n6997) );
  INV_X1 U9673 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n9444) );
  OR2_X1 U9674 ( .A1(n8539), .A2(n7693), .ZN(n6712) );
  INV_X1 U9675 ( .A(P3_IR_REG_6__SCAN_IN), .ZN(n7082) );
  INV_X1 U9676 ( .A(P3_IR_REG_31__SCAN_IN), .ZN(n6998) );
  OR2_X1 U9677 ( .A1(n6609), .A2(n7512), .ZN(n6713) );
  NAND2_X1 U9678 ( .A1(n10662), .A2(P3_REG1_REG_4__SCAN_IN), .ZN(n6714) );
  INV_X1 U9679 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n7053) );
  NAND3_X1 U9680 ( .A1(n6899), .A2(n6898), .A3(n6896), .ZN(P2_U3233) );
  INV_X1 U9681 ( .A(n11436), .ZN(n12957) );
  INV_X1 U9682 ( .A(n14628), .ZN(n7905) );
  INV_X1 U9683 ( .A(n9006), .ZN(n7718) );
  INV_X1 U9684 ( .A(n15605), .ZN(n7456) );
  INV_X1 U9685 ( .A(n7196), .ZN(n8756) );
  NAND2_X1 U9686 ( .A1(n8754), .A2(n12061), .ZN(n7196) );
  INV_X1 U9687 ( .A(P3_REG2_REG_2__SCAN_IN), .ZN(n7654) );
  INV_X1 U9688 ( .A(n12967), .ZN(n7857) );
  NAND2_X1 U9689 ( .A1(n8595), .A2(n8594), .ZN(n12615) );
  NOR2_X1 U9690 ( .A1(n6953), .A2(n6955), .ZN(n12465) );
  AND2_X1 U9691 ( .A1(n15471), .A2(n15459), .ZN(n15440) );
  NAND2_X1 U9692 ( .A1(n9814), .A2(n9813), .ZN(n15602) );
  INV_X1 U9693 ( .A(n15602), .ZN(n7457) );
  AND2_X1 U9694 ( .A1(n12340), .A2(n7455), .ZN(n12367) );
  INV_X2 U9695 ( .A(n16092), .ZN(n16094) );
  NAND2_X1 U9696 ( .A1(n15527), .A2(n15511), .ZN(n15489) );
  AOI21_X1 U9697 ( .B1(n13295), .B2(n6564), .A(n13293), .ZN(n13893) );
  INV_X1 U9698 ( .A(n11430), .ZN(n7478) );
  NAND2_X1 U9699 ( .A1(n6976), .A2(n13543), .ZN(n13548) );
  OAI21_X1 U9700 ( .B1(n12376), .B2(n8610), .A(n7016), .ZN(n12657) );
  NAND2_X1 U9701 ( .A1(n8228), .A2(n8227), .ZN(n12825) );
  NAND2_X1 U9702 ( .A1(n6884), .A2(n13028), .ZN(n15499) );
  INV_X1 U9703 ( .A(n13801), .ZN(n7040) );
  NAND2_X1 U9704 ( .A1(n6826), .A2(n7011), .ZN(n12185) );
  OR2_X1 U9705 ( .A1(n12113), .A2(n13381), .ZN(n12114) );
  AND2_X1 U9706 ( .A1(n7421), .A2(n7426), .ZN(n6716) );
  NAND2_X1 U9707 ( .A1(n12407), .A2(n7964), .ZN(n12510) );
  NAND2_X1 U9708 ( .A1(n6967), .A2(n6624), .ZN(n14037) );
  NAND2_X1 U9709 ( .A1(n7493), .A2(n7491), .ZN(n13267) );
  NAND2_X1 U9710 ( .A1(n6959), .A2(n10457), .ZN(n12297) );
  INV_X1 U9711 ( .A(n12836), .ZN(n7224) );
  INV_X1 U9712 ( .A(n13595), .ZN(n7436) );
  NOR2_X1 U9713 ( .A1(n12486), .A2(n7482), .ZN(n6717) );
  OR2_X1 U9714 ( .A1(n6598), .A2(n7466), .ZN(n6718) );
  AND2_X1 U9715 ( .A1(n7832), .A2(n7831), .ZN(n6719) );
  NOR2_X1 U9716 ( .A1(n9956), .A2(n9955), .ZN(n6720) );
  OR2_X1 U9717 ( .A1(n13404), .A2(n13816), .ZN(n9136) );
  OR2_X1 U9718 ( .A1(n12334), .A2(P2_ADDR_REG_11__SCAN_IN), .ZN(n6721) );
  INV_X1 U9719 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n10639) );
  INV_X1 U9720 ( .A(n7472), .ZN(n7471) );
  NAND2_X1 U9721 ( .A1(n13204), .A2(n13722), .ZN(n7472) );
  AND2_X1 U9722 ( .A1(P1_REG3_REG_12__SCAN_IN), .A2(P1_REG3_REG_13__SCAN_IN), 
        .ZN(n6722) );
  NAND2_X1 U9723 ( .A1(n10202), .A2(n10201), .ZN(n12407) );
  INV_X1 U9724 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n10705) );
  INV_X1 U9725 ( .A(n7713), .ZN(n7712) );
  OR2_X1 U9726 ( .A1(n8709), .A2(P3_IR_REG_16__SCAN_IN), .ZN(n6723) );
  AND2_X1 U9727 ( .A1(n9170), .A2(P1_DATAO_REG_16__SCAN_IN), .ZN(n6724) );
  OR2_X1 U9728 ( .A1(n13595), .A2(n6603), .ZN(n6725) );
  OR2_X1 U9729 ( .A1(n8475), .A2(SI_23_), .ZN(n6726) );
  OR2_X1 U9730 ( .A1(n8507), .A2(SI_25_), .ZN(n6727) );
  AND2_X1 U9731 ( .A1(n7939), .A2(n7941), .ZN(n6728) );
  AND2_X1 U9732 ( .A1(n7322), .A2(n10861), .ZN(n6729) );
  INV_X1 U9733 ( .A(n12179), .ZN(n7942) );
  INV_X1 U9735 ( .A(n14103), .ZN(n14065) );
  NAND2_X1 U9736 ( .A1(n6958), .A2(n8584), .ZN(n10420) );
  INV_X1 U9737 ( .A(n13264), .ZN(n13243) );
  INV_X1 U9738 ( .A(n14809), .ZN(n7114) );
  AND2_X2 U9739 ( .A1(n11495), .A2(n11494), .ZN(n15886) );
  NAND2_X1 U9740 ( .A1(n8162), .A2(n8161), .ZN(n14154) );
  INV_X1 U9741 ( .A(n14154), .ZN(n7233) );
  INV_X1 U9742 ( .A(n7401), .ZN(n11281) );
  NOR2_X1 U9743 ( .A1(n16016), .A2(n11282), .ZN(n7401) );
  INV_X1 U9744 ( .A(n14329), .ZN(n7740) );
  INV_X1 U9745 ( .A(n13594), .ZN(n7434) );
  AND2_X1 U9746 ( .A1(n7898), .A2(n8585), .ZN(n6730) );
  AOI21_X1 U9747 ( .B1(n8818), .B2(n9006), .A(n8819), .ZN(n11535) );
  NAND2_X1 U9748 ( .A1(n7783), .A2(n12213), .ZN(n15775) );
  OR2_X1 U9749 ( .A1(n13510), .A2(n9375), .ZN(n16013) );
  INV_X1 U9750 ( .A(n8513), .ZN(n7891) );
  INV_X1 U9751 ( .A(n11692), .ZN(n7420) );
  NAND2_X1 U9752 ( .A1(n11417), .A2(n11416), .ZN(n13264) );
  AOI21_X1 U9753 ( .B1(n11243), .B2(n11391), .A(n11392), .ZN(n11390) );
  NAND2_X1 U9754 ( .A1(n6841), .A2(n11942), .ZN(n6839) );
  OR2_X1 U9755 ( .A1(n15877), .A2(n6790), .ZN(n6731) );
  NAND2_X1 U9756 ( .A1(n8819), .A2(n7732), .ZN(n7729) );
  NAND2_X1 U9757 ( .A1(n11606), .A2(n11605), .ZN(n11653) );
  INV_X1 U9758 ( .A(n11963), .ZN(n7450) );
  AND2_X1 U9759 ( .A1(n7720), .A2(n7719), .ZN(n6732) );
  INV_X1 U9760 ( .A(n7517), .ZN(n7516) );
  INV_X1 U9761 ( .A(n7661), .ZN(n11689) );
  OAI21_X1 U9762 ( .B1(n11390), .B2(n6989), .A(n7718), .ZN(n7661) );
  INV_X1 U9763 ( .A(n15633), .ZN(n6801) );
  INV_X1 U9764 ( .A(n7447), .ZN(n15809) );
  NAND2_X1 U9765 ( .A1(n7191), .A2(n7190), .ZN(n12225) );
  NOR2_X1 U9766 ( .A1(n7662), .A2(n11689), .ZN(n6733) );
  OR2_X1 U9767 ( .A1(n15877), .A2(n7097), .ZN(n6734) );
  OR2_X1 U9768 ( .A1(n15877), .A2(n7451), .ZN(n6735) );
  NAND2_X1 U9769 ( .A1(n12792), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n6736) );
  NOR2_X1 U9770 ( .A1(n9337), .A2(n7614), .ZN(n7613) );
  INV_X1 U9771 ( .A(n15227), .ZN(n6868) );
  NAND2_X1 U9772 ( .A1(n15810), .A2(n9780), .ZN(n11835) );
  NAND2_X1 U9773 ( .A1(n11315), .A2(P3_REG2_REG_3__SCAN_IN), .ZN(n11265) );
  INV_X1 U9774 ( .A(n14322), .ZN(n8584) );
  NAND2_X1 U9775 ( .A1(n8771), .A2(n8776), .ZN(n13515) );
  INV_X1 U9776 ( .A(n13515), .ZN(n6904) );
  INV_X1 U9777 ( .A(n11260), .ZN(n7407) );
  INV_X1 U9778 ( .A(n9780), .ZN(n15250) );
  INV_X1 U9779 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n7512) );
  INV_X1 U9780 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n7444) );
  INV_X1 U9781 ( .A(P3_REG2_REG_17__SCAN_IN), .ZN(n7652) );
  INV_X1 U9782 ( .A(P3_REG0_REG_1__SCAN_IN), .ZN(n7172) );
  INV_X1 U9783 ( .A(P3_ADDR_REG_5__SCAN_IN), .ZN(n7495) );
  INV_X1 U9784 ( .A(n9481), .ZN(n6737) );
  AND2_X1 U9785 ( .A1(n6741), .A2(n6739), .ZN(n9571) );
  NAND3_X1 U9786 ( .A1(n6740), .A2(n6743), .A3(n6742), .ZN(n6739) );
  NAND2_X1 U9787 ( .A1(n9554), .A2(n9553), .ZN(n6740) );
  OR2_X1 U9788 ( .A1(n9553), .A2(n9554), .ZN(n6741) );
  NAND3_X1 U9789 ( .A1(n9538), .A2(n11804), .A3(n9539), .ZN(n6743) );
  NAND2_X1 U9790 ( .A1(n15045), .A2(n9635), .ZN(n6744) );
  NAND2_X1 U9791 ( .A1(n15393), .A2(n9956), .ZN(n6745) );
  NAND2_X1 U9792 ( .A1(n6747), .A2(n6746), .ZN(n9895) );
  NAND2_X1 U9793 ( .A1(n6751), .A2(n7924), .ZN(n6750) );
  OR2_X1 U9794 ( .A1(n9811), .A2(n7235), .ZN(n6751) );
  NAND2_X1 U9795 ( .A1(n6756), .A2(n6752), .ZN(n9769) );
  NAND2_X1 U9796 ( .A1(n6753), .A2(n9692), .ZN(n6752) );
  INV_X1 U9797 ( .A(n7915), .ZN(n6754) );
  NAND2_X1 U9798 ( .A1(n9674), .A2(n7914), .ZN(n6755) );
  NAND2_X1 U9799 ( .A1(n6757), .A2(n9690), .ZN(n6756) );
  NAND2_X1 U9800 ( .A1(n6758), .A2(n9691), .ZN(n6757) );
  OAI21_X1 U9801 ( .B1(n9674), .B2(n7915), .A(n7914), .ZN(n6758) );
  NAND3_X1 U9802 ( .A1(n9534), .A2(n9465), .A3(n9464), .ZN(n9739) );
  NAND4_X1 U9803 ( .A1(n9534), .A2(n9465), .A3(n9464), .A4(n6759), .ZN(n9756)
         );
  NOR2_X2 U9804 ( .A1(n9756), .A2(P1_IR_REG_17__SCAN_IN), .ZN(n9751) );
  NAND3_X1 U9805 ( .A1(n9622), .A2(n6710), .A3(n6760), .ZN(n7214) );
  NAND2_X1 U9806 ( .A1(n6761), .A2(n9620), .ZN(n6760) );
  NAND2_X1 U9807 ( .A1(n6762), .A2(n6700), .ZN(n6761) );
  NAND2_X1 U9808 ( .A1(n9605), .A2(n7912), .ZN(n6762) );
  NAND3_X1 U9809 ( .A1(n7486), .A2(n6764), .A3(n6763), .ZN(n6768) );
  NAND2_X1 U9810 ( .A1(n6769), .A2(n11912), .ZN(n6764) );
  INV_X1 U9811 ( .A(n6768), .ZN(n12281) );
  OAI21_X2 U9812 ( .B1(n12256), .B2(n7480), .A(n7479), .ZN(n12855) );
  INV_X1 U9813 ( .A(n7487), .ZN(n6769) );
  INV_X1 U9814 ( .A(n8811), .ZN(n6996) );
  OAI21_X1 U9815 ( .B1(n8811), .B2(n6998), .A(P3_IR_REG_2__SCAN_IN), .ZN(n6994) );
  NOR2_X1 U9816 ( .A1(n11433), .A2(n11499), .ZN(n11438) );
  AND2_X4 U9817 ( .A1(n6777), .A2(n8915), .ZN(n16056) );
  AND2_X2 U9818 ( .A1(n8916), .A2(n8914), .ZN(n6777) );
  XNOR2_X2 U9819 ( .A(n6784), .B(n8805), .ZN(n8808) );
  OAI211_X2 U9820 ( .C1(n6787), .C2(n7363), .A(n6785), .B(n8330), .ZN(n8344)
         );
  INV_X1 U9821 ( .A(n6793), .ZN(n8512) );
  NAND2_X1 U9822 ( .A1(n9513), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n9520) );
  NAND2_X2 U9823 ( .A1(n10073), .A2(n15699), .ZN(n9514) );
  NAND2_X1 U9824 ( .A1(n14315), .A2(n6584), .ZN(n6795) );
  NAND3_X1 U9825 ( .A1(n6697), .A2(n6798), .A3(n6797), .ZN(n6796) );
  NAND2_X1 U9826 ( .A1(n10140), .A2(n11798), .ZN(n10141) );
  NAND3_X1 U9827 ( .A1(n15527), .A2(n15511), .A3(n6801), .ZN(n15490) );
  INV_X1 U9828 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n6802) );
  INV_X1 U9829 ( .A(P2_RD_REG_SCAN_IN), .ZN(n6804) );
  INV_X1 U9830 ( .A(P1_RD_REG_SCAN_IN), .ZN(n6806) );
  INV_X1 U9831 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n8014) );
  AND4_X2 U9832 ( .A1(n6812), .A2(n6810), .A3(n6809), .A4(n6808), .ZN(n8231)
         );
  NAND3_X1 U9833 ( .A1(n8196), .A2(n7065), .A3(n8192), .ZN(n6808) );
  NAND3_X1 U9834 ( .A1(n6811), .A2(n8156), .A3(n6813), .ZN(n6810) );
  NAND2_X1 U9835 ( .A1(n8173), .A2(n6586), .ZN(n6812) );
  NOR2_X2 U9836 ( .A1(n7066), .A2(n6618), .ZN(n6813) );
  NAND3_X1 U9837 ( .A1(n7448), .A2(n7449), .A3(n12035), .ZN(n12206) );
  NAND3_X1 U9838 ( .A1(n6817), .A2(n14577), .A3(n6815), .ZN(n14580) );
  NAND3_X1 U9839 ( .A1(n14637), .A2(n7630), .A3(n8469), .ZN(n6815) );
  NAND2_X1 U9840 ( .A1(n6819), .A2(n6818), .ZN(n6816) );
  NAND2_X1 U9841 ( .A1(n8506), .A2(n8505), .ZN(n6823) );
  OAI21_X2 U9842 ( .B1(n8228), .B2(n7636), .A(n7634), .ZN(n12916) );
  NAND2_X2 U9843 ( .A1(n12374), .A2(n12379), .ZN(n12376) );
  NAND2_X1 U9844 ( .A1(n6826), .A2(n8150), .ZN(n12187) );
  AND3_X2 U9845 ( .A1(n6948), .A2(n7192), .A3(n6827), .ZN(n11713) );
  NAND2_X1 U9846 ( .A1(n11577), .A2(n11576), .ZN(n11944) );
  NAND3_X1 U9847 ( .A1(n6834), .A2(n6832), .A3(n14478), .ZN(n6842) );
  NAND3_X1 U9848 ( .A1(n11577), .A2(n6833), .A3(n6839), .ZN(n6832) );
  NAND2_X1 U9849 ( .A1(n6840), .A2(n11577), .ZN(n6836) );
  OAI21_X1 U9850 ( .B1(n11577), .B2(n11943), .A(n6839), .ZN(n6838) );
  NAND3_X1 U9851 ( .A1(n10675), .A2(n6846), .A3(n6845), .ZN(n10676) );
  NAND2_X1 U9852 ( .A1(n7497), .A2(n7500), .ZN(n6846) );
  XNOR2_X1 U9853 ( .A(n6847), .B(P2_ADDR_REG_18__SCAN_IN), .ZN(SUB_1596_U62)
         );
  NAND3_X1 U9854 ( .A1(n15765), .A2(n7503), .A3(n7502), .ZN(n6847) );
  NAND2_X1 U9855 ( .A1(n15753), .A2(n6594), .ZN(n7502) );
  NAND2_X1 U9856 ( .A1(n6849), .A2(n6848), .ZN(n15765) );
  NAND2_X1 U9857 ( .A1(n15753), .A2(n15752), .ZN(n6849) );
  INV_X1 U9858 ( .A(n6852), .ZN(n15740) );
  INV_X1 U9859 ( .A(n6850), .ZN(n15743) );
  NAND2_X1 U9860 ( .A1(n6854), .A2(n6648), .ZN(n6850) );
  NAND2_X1 U9861 ( .A1(n7507), .A2(n6853), .ZN(n6852) );
  INV_X1 U9862 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n6853) );
  NAND2_X1 U9863 ( .A1(n15737), .A2(n15739), .ZN(n6854) );
  NAND2_X1 U9864 ( .A1(n15736), .A2(P2_ADDR_REG_15__SCAN_IN), .ZN(n15737) );
  INV_X1 U9865 ( .A(n7507), .ZN(n15736) );
  OAI21_X2 U9866 ( .B1(n12324), .B2(n12323), .A(n12327), .ZN(n12333) );
  NAND2_X1 U9867 ( .A1(n15940), .A2(n6877), .ZN(n6876) );
  NAND2_X1 U9868 ( .A1(n6881), .A2(n6882), .ZN(n15484) );
  NAND3_X1 U9869 ( .A1(n15518), .A2(n13029), .A3(n6706), .ZN(n6881) );
  NAND4_X1 U9870 ( .A1(n9465), .A2(n6886), .A3(n7779), .A4(n7778), .ZN(n15689)
         );
  AND2_X1 U9871 ( .A1(n6583), .A2(n9448), .ZN(n6887) );
  AND4_X2 U9872 ( .A1(n7780), .A2(n10816), .A3(n9441), .A4(n9440), .ZN(n9465)
         );
  INV_X1 U9873 ( .A(n9465), .ZN(n9719) );
  OR2_X2 U9874 ( .A1(n15465), .A2(n15467), .ZN(n7825) );
  NAND3_X1 U9875 ( .A1(n15555), .A2(n7138), .A3(n15554), .ZN(n15669) );
  OAI22_X1 U9876 ( .A1(n14505), .A2(n14504), .B1(n14503), .B2(n15904), .ZN(
        n6897) );
  OAI21_X1 U9877 ( .B1(n13526), .B2(n6905), .A(n13631), .ZN(n13527) );
  NAND2_X1 U9878 ( .A1(n7707), .A2(n7717), .ZN(n13573) );
  INV_X1 U9879 ( .A(n8817), .ZN(n11395) );
  NAND2_X1 U9880 ( .A1(n8817), .A2(n7721), .ZN(n7720) );
  NAND3_X1 U9881 ( .A1(n11245), .A2(n7718), .A3(n6641), .ZN(n6910) );
  NOR2_X2 U9882 ( .A1(n8817), .A2(n6911), .ZN(n11245) );
  NOR2_X1 U9883 ( .A1(n7702), .A2(n7646), .ZN(n6911) );
  NAND3_X1 U9884 ( .A1(n7723), .A2(n6912), .A3(P3_REG1_REG_9__SCAN_IN), .ZN(
        n6914) );
  INV_X1 U9885 ( .A(n6914), .ZN(n12048) );
  NAND2_X1 U9886 ( .A1(n6913), .A2(n10592), .ZN(n10595) );
  NAND3_X1 U9887 ( .A1(n7100), .A2(P3_REG1_REG_17__SCAN_IN), .A3(n13629), .ZN(
        n13630) );
  OAI21_X1 U9888 ( .B1(P3_REG1_REG_17__SCAN_IN), .B2(n6703), .A(n13630), .ZN(
        n13620) );
  NAND2_X1 U9889 ( .A1(n7578), .A2(n6917), .ZN(n7577) );
  XNOR2_X1 U9890 ( .A(n6917), .B(n8934), .ZN(n10730) );
  XNOR2_X1 U9891 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(P1_DATAO_REG_1__SCAN_IN), 
        .ZN(n6917) );
  NAND2_X1 U9892 ( .A1(n6920), .A2(n6921), .ZN(n9196) );
  NAND2_X1 U9893 ( .A1(n7588), .A2(n6922), .ZN(n6920) );
  INV_X1 U9894 ( .A(n6926), .ZN(n6925) );
  OAI211_X1 U9895 ( .C1(n13707), .C2(n6926), .A(n6924), .B(n13310), .ZN(n10077) );
  INV_X1 U9896 ( .A(n7246), .ZN(n7245) );
  NAND2_X1 U9897 ( .A1(n8368), .A2(n14428), .ZN(n6948) );
  NAND2_X1 U9898 ( .A1(n6949), .A2(n8004), .ZN(n8656) );
  NAND2_X1 U9899 ( .A1(n6949), .A2(n6692), .ZN(n6972) );
  NAND2_X1 U9900 ( .A1(n6949), .A2(n8001), .ZN(n8571) );
  NAND2_X1 U9901 ( .A1(n6949), .A2(n7776), .ZN(n8577) );
  NAND2_X1 U9902 ( .A1(n6949), .A2(n8565), .ZN(n8576) );
  NAND2_X1 U9903 ( .A1(n6949), .A2(n6707), .ZN(n8580) );
  OR2_X1 U9904 ( .A1(n6949), .A2(n8006), .ZN(n8332) );
  NAND2_X1 U9905 ( .A1(n7165), .A2(n6949), .ZN(n7310) );
  AND2_X4 U9906 ( .A1(n6969), .A2(n8180), .ZN(n6949) );
  NAND3_X1 U9907 ( .A1(n6581), .A2(n14676), .A3(n6952), .ZN(n14572) );
  INV_X1 U9908 ( .A(n12188), .ZN(n6954) );
  NOR2_X1 U9909 ( .A1(n6955), .A2(n12188), .ZN(n12464) );
  NAND2_X1 U9910 ( .A1(n6954), .A2(n12468), .ZN(n6953) );
  NAND2_X1 U9911 ( .A1(n6956), .A2(n10435), .ZN(n11619) );
  NAND3_X1 U9912 ( .A1(n6957), .A2(n10431), .A3(n11568), .ZN(n6956) );
  NAND2_X1 U9913 ( .A1(n10430), .A2(n11448), .ZN(n6957) );
  NAND2_X1 U9914 ( .A1(n6959), .A2(n6597), .ZN(n12298) );
  NAND2_X1 U9915 ( .A1(n6960), .A2(n6961), .ZN(n14082) );
  NAND2_X1 U9916 ( .A1(n14048), .A2(n6963), .ZN(n6960) );
  OAI21_X2 U9917 ( .B1(n14048), .B2(n6965), .A(n6963), .ZN(n14017) );
  NAND2_X1 U9918 ( .A1(n6967), .A2(n6966), .ZN(n7762) );
  NOR2_X2 U9919 ( .A1(n8100), .A2(n7994), .ZN(n8180) );
  INV_X1 U9920 ( .A(n11619), .ZN(n6970) );
  XNOR2_X1 U9921 ( .A(n7166), .B(n10436), .ZN(n10425) );
  NAND2_X1 U9922 ( .A1(n6972), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8563) );
  NAND2_X1 U9923 ( .A1(n14055), .A2(n6974), .ZN(n14009) );
  INV_X1 U9924 ( .A(n6976), .ZN(n6975) );
  NAND2_X1 U9925 ( .A1(n13590), .A2(n6984), .ZN(n6978) );
  NAND2_X1 U9926 ( .A1(n6555), .A2(n13616), .ZN(n6981) );
  NAND2_X1 U9927 ( .A1(n6977), .A2(n7649), .ZN(n8791) );
  AND2_X1 U9928 ( .A1(n7648), .A2(n8788), .ZN(n6977) );
  NAND3_X1 U9929 ( .A1(n6981), .A2(n6983), .A3(n6978), .ZN(n13611) );
  NAND2_X1 U9930 ( .A1(n12594), .A2(n6987), .ZN(n13512) );
  NAND2_X1 U9931 ( .A1(n8764), .A2(n12601), .ZN(n6987) );
  AND2_X1 U9932 ( .A1(n6986), .A2(n6987), .ZN(n12595) );
  INV_X1 U9933 ( .A(n11390), .ZN(n6988) );
  NAND2_X1 U9934 ( .A1(n7663), .A2(P3_REG2_REG_7__SCAN_IN), .ZN(n7662) );
  NAND2_X1 U9935 ( .A1(n7662), .A2(n7661), .ZN(n7660) );
  NAND2_X1 U9936 ( .A1(n6992), .A2(n13588), .ZN(n7641) );
  NAND2_X1 U9937 ( .A1(n7113), .A2(n13582), .ZN(n6993) );
  NAND3_X1 U9938 ( .A1(n6996), .A2(n6997), .A3(P3_IR_REG_31__SCAN_IN), .ZN(
        n6995) );
  INV_X1 U9939 ( .A(n7010), .ZN(n7848) );
  NAND2_X1 U9940 ( .A1(n13719), .A2(n9255), .ZN(n7009) );
  NAND2_X1 U9941 ( .A1(n12230), .A2(n12231), .ZN(n7013) );
  NAND2_X1 U9942 ( .A1(n12221), .A2(n6639), .ZN(n7014) );
  NAND2_X1 U9943 ( .A1(n11815), .A2(n14338), .ZN(n12221) );
  NAND3_X1 U9944 ( .A1(n7021), .A2(n8612), .A3(n14344), .ZN(n7019) );
  NAND2_X1 U9945 ( .A1(n8610), .A2(n7022), .ZN(n7021) );
  NAND2_X2 U9946 ( .A1(n7033), .A2(n8381), .ZN(n14637) );
  NAND2_X1 U9947 ( .A1(n14655), .A2(n8380), .ZN(n7033) );
  NAND2_X1 U9948 ( .A1(n13800), .A2(n7037), .ZN(n7036) );
  NAND2_X2 U9949 ( .A1(n7036), .A2(n7034), .ZN(n13790) );
  NAND2_X1 U9950 ( .A1(n7038), .A2(n13802), .ZN(n13786) );
  INV_X1 U9951 ( .A(n13787), .ZN(n7039) );
  OAI21_X2 U9952 ( .B1(n14951), .B2(n7045), .A(n7043), .ZN(n15019) );
  NAND2_X1 U9953 ( .A1(n7620), .A2(n7617), .ZN(n14535) );
  INV_X2 U9954 ( .A(n10151), .ZN(n10140) );
  NAND2_X1 U9955 ( .A1(n7057), .A2(n10656), .ZN(n7351) );
  XNOR2_X1 U9956 ( .A(n7058), .B(n8307), .ZN(n11588) );
  NAND2_X1 U9957 ( .A1(n7059), .A2(n8095), .ZN(n8124) );
  OAI21_X2 U9958 ( .B1(n7059), .B2(n8125), .A(n7264), .ZN(n8133) );
  NAND2_X1 U9959 ( .A1(n8093), .A2(n8092), .ZN(n7059) );
  NAND2_X1 U9960 ( .A1(n8175), .A2(n8174), .ZN(n7067) );
  NAND3_X1 U9961 ( .A1(n13005), .A2(n7096), .A3(n13006), .ZN(n7068) );
  NAND2_X1 U9962 ( .A1(n12983), .A2(n6564), .ZN(n7074) );
  NAND2_X1 U9964 ( .A1(n11626), .A2(n11625), .ZN(n11624) );
  NAND2_X2 U9965 ( .A1(n7075), .A2(n8013), .ZN(n14421) );
  OAI21_X1 U9967 ( .B1(n14518), .B2(n16000), .A(n14521), .ZN(n8651) );
  NAND2_X1 U9968 ( .A1(n6667), .A2(n7693), .ZN(n8562) );
  NAND2_X1 U9969 ( .A1(n7076), .A2(n11609), .ZN(n7261) );
  NAND4_X1 U9970 ( .A1(n6687), .A2(n7262), .A3(n7373), .A4(n6589), .ZN(n7076)
         );
  NAND2_X1 U9971 ( .A1(n7146), .A2(n7148), .ZN(n13307) );
  OAI21_X1 U9972 ( .B1(n13479), .B2(n13305), .A(n13304), .ZN(n7147) );
  INV_X1 U9973 ( .A(n8472), .ZN(n7198) );
  NAND2_X1 U9974 ( .A1(n7280), .A2(n7279), .ZN(n14055) );
  NAND2_X1 U9975 ( .A1(n7760), .A2(n7762), .ZN(n7280) );
  NAND2_X1 U9976 ( .A1(n10711), .A2(n10006), .ZN(n9619) );
  INV_X1 U9977 ( .A(n13899), .ZN(n7129) );
  INV_X1 U9978 ( .A(n12216), .ZN(n7789) );
  OAI21_X1 U9979 ( .B1(n13053), .B2(n13054), .A(n6578), .ZN(n7347) );
  NAND3_X1 U9980 ( .A1(n7328), .A2(n6708), .A3(n7595), .ZN(n7594) );
  AND4_X2 U9981 ( .A1(n9515), .A2(n9462), .A3(n9469), .A4(n9439), .ZN(n7779)
         );
  NAND2_X1 U9982 ( .A1(n7668), .A2(n7669), .ZN(n7078) );
  NAND3_X1 U9983 ( .A1(n15485), .A2(n13029), .A3(n15482), .ZN(n13004) );
  NAND2_X1 U9984 ( .A1(n13890), .A2(n13646), .ZN(n7080) );
  NOR2_X1 U9985 ( .A1(n14743), .A2(n7177), .ZN(n14745) );
  INV_X1 U9986 ( .A(n7906), .ZN(n7179) );
  AOI22_X1 U9987 ( .A1(n13533), .A2(n7708), .B1(n7712), .B2(n7715), .ZN(n7707)
         );
  INV_X1 U9988 ( .A(n8826), .ZN(n7101) );
  NOR2_X1 U9989 ( .A1(n8823), .A2(n8822), .ZN(n13565) );
  AOI21_X1 U9990 ( .B1(n7378), .B2(n7380), .A(n13457), .ZN(n7377) );
  NAND2_X1 U9991 ( .A1(n13311), .A2(n13675), .ZN(n13448) );
  NAND2_X2 U9992 ( .A1(n13728), .A2(n9237), .ZN(n13719) );
  NAND2_X1 U9993 ( .A1(n13451), .A2(n13679), .ZN(n7381) );
  NAND2_X1 U9994 ( .A1(n11868), .A2(n7966), .ZN(n9042) );
  NAND2_X1 U9995 ( .A1(n14555), .A2(n8637), .ZN(n14541) );
  NAND2_X1 U9996 ( .A1(n7081), .A2(n8723), .ZN(n8725) );
  INV_X1 U9997 ( .A(n8749), .ZN(n7081) );
  NAND2_X1 U9998 ( .A1(n6560), .A2(n7082), .ZN(n8749) );
  AND3_X2 U9999 ( .A1(n8926), .A2(n8924), .A3(n8925), .ZN(n11845) );
  OR2_X1 U10000 ( .A1(n9224), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n9226) );
  INV_X1 U10001 ( .A(n7506), .ZN(n7124) );
  NAND3_X1 U10002 ( .A1(n9896), .A2(n9897), .A3(n9929), .ZN(n7083) );
  NAND2_X2 U10003 ( .A1(n7084), .A2(n9945), .ZN(n9651) );
  AND2_X1 U10004 ( .A1(n13509), .A2(n11886), .ZN(n8984) );
  OAI21_X1 U10005 ( .B1(n12333), .B2(n6713), .A(n7086), .ZN(n7085) );
  AOI21_X1 U10006 ( .B1(n7239), .B2(n7238), .A(n7237), .ZN(n9587) );
  NAND2_X1 U10007 ( .A1(n7087), .A2(n10076), .ZN(P1_U3242) );
  NAND2_X1 U10008 ( .A1(n7088), .A2(n12318), .ZN(n7087) );
  NAND4_X1 U10009 ( .A1(n10053), .A2(n10055), .A3(n10052), .A4(n10054), .ZN(
        n7088) );
  NAND2_X1 U10010 ( .A1(n8755), .A2(n8867), .ZN(n7195) );
  INV_X1 U10011 ( .A(n10010), .ZN(n10022) );
  NAND3_X1 U10012 ( .A1(n7092), .A2(n14390), .A3(n7091), .ZN(P2_U3328) );
  INV_X1 U10013 ( .A(n10430), .ZN(n11446) );
  AOI21_X2 U10014 ( .B1(n12246), .B2(n12126), .A(n9022), .ZN(n12267) );
  INV_X1 U10015 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n10750) );
  OAI21_X1 U10016 ( .B1(n9321), .B2(n9320), .A(n9322), .ZN(n9338) );
  NAND2_X1 U10017 ( .A1(n7137), .A2(n7136), .ZN(n11794) );
  NAND2_X1 U10018 ( .A1(n15531), .A2(n13001), .ZN(n15481) );
  OAI21_X2 U10019 ( .B1(n12722), .B2(n12564), .A(n12563), .ZN(n12565) );
  NAND3_X1 U10020 ( .A1(n7349), .A2(n7932), .A3(n9465), .ZN(n7933) );
  NAND2_X1 U10021 ( .A1(n7793), .A2(n7794), .ZN(n15531) );
  NAND2_X1 U10022 ( .A1(n7098), .A2(n6734), .ZN(P1_U3523) );
  NAND2_X1 U10023 ( .A1(n15670), .A2(n15877), .ZN(n7098) );
  NAND2_X1 U10024 ( .A1(n11666), .A2(n10006), .ZN(n7106) );
  INV_X1 U10025 ( .A(n14637), .ZN(n8401) );
  AND2_X1 U10026 ( .A1(n12033), .A2(n12213), .ZN(n7223) );
  NAND2_X1 U10027 ( .A1(n7704), .A2(n7698), .ZN(n7699) );
  NAND2_X1 U10028 ( .A1(n7101), .A2(n9171), .ZN(n7100) );
  AND2_X2 U10029 ( .A1(n15526), .A2(n15530), .ZN(n15527) );
  AND2_X2 U10030 ( .A1(n12567), .A2(n14978), .ZN(n15526) );
  NAND2_X1 U10031 ( .A1(n8365), .A2(n8364), .ZN(n8366) );
  NAND2_X2 U10032 ( .A1(n7106), .A2(n9722), .ZN(n15633) );
  INV_X1 U10033 ( .A(n7961), .ZN(n7960) );
  NAND2_X1 U10034 ( .A1(n7919), .A2(n9585), .ZN(n7918) );
  OAI21_X2 U10035 ( .B1(n12880), .B2(n13502), .A(n12879), .ZN(n12932) );
  NAND2_X1 U10036 ( .A1(n7110), .A2(n8696), .ZN(n8784) );
  NAND2_X1 U10037 ( .A1(n13164), .A2(n12953), .ZN(n13214) );
  NAND2_X1 U10038 ( .A1(n7490), .A2(n7489), .ZN(n13186) );
  AOI211_X2 U10039 ( .C1(n15993), .C2(n14765), .A(n14764), .B(n14763), .ZN(
        n14857) );
  OAI21_X4 U10040 ( .B1(n11973), .B2(n7140), .A(n8352), .ZN(n14800) );
  OAI21_X1 U10041 ( .B1(n15270), .B2(n7139), .A(n15271), .ZN(n15276) );
  NAND2_X1 U10042 ( .A1(n12052), .A2(n7657), .ZN(n7656) );
  NAND2_X1 U10043 ( .A1(n7346), .A2(n15295), .ZN(n7341) );
  INV_X1 U10044 ( .A(n8782), .ZN(n7113) );
  NAND2_X1 U10045 ( .A1(n8826), .A2(n13616), .ZN(n13629) );
  INV_X1 U10046 ( .A(n14083), .ZN(n7743) );
  NAND2_X1 U10047 ( .A1(n12215), .A2(n12214), .ZN(n12336) );
  NAND2_X1 U10048 ( .A1(n14237), .A2(n14236), .ZN(n14240) );
  NAND2_X1 U10049 ( .A1(n12562), .A2(n12561), .ZN(n12722) );
  NAND3_X1 U10050 ( .A1(n14226), .A2(n14196), .A3(n14197), .ZN(n7522) );
  NAND2_X2 U10051 ( .A1(n11179), .A2(n14912), .ZN(n8036) );
  NAND2_X1 U10052 ( .A1(n14847), .A2(n16011), .ZN(n7119) );
  NAND3_X1 U10053 ( .A1(n11638), .A2(n13313), .A3(n12101), .ZN(n7120) );
  NAND2_X1 U10054 ( .A1(n14082), .A2(n14084), .ZN(n7187) );
  MUX2_X1 U10055 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8563), .S(
        P2_IR_REG_21__SCAN_IN), .Z(n8566) );
  NAND2_X1 U10056 ( .A1(n11793), .A2(n11794), .ZN(n11797) );
  NAND2_X1 U10057 ( .A1(n7628), .A2(n8467), .ZN(n7627) );
  INV_X1 U10058 ( .A(n9136), .ZN(n7842) );
  NAND2_X1 U10059 ( .A1(n7199), .A2(n7198), .ZN(n7197) );
  NAND2_X1 U10060 ( .A1(n9136), .A2(n13325), .ZN(n7194) );
  NAND2_X1 U10061 ( .A1(n11803), .A2(n7826), .ZN(n11856) );
  NAND2_X1 U10062 ( .A1(n13033), .A2(n13032), .ZN(n15465) );
  NAND2_X1 U10063 ( .A1(n7809), .A2(n7125), .ZN(n15518) );
  NAND2_X1 U10064 ( .A1(n7811), .A2(n12362), .ZN(n7125) );
  NAND2_X1 U10065 ( .A1(n11528), .A2(n11526), .ZN(n11524) );
  OAI21_X1 U10066 ( .B1(n15720), .B2(n15719), .A(n15724), .ZN(n7507) );
  OAI21_X4 U10067 ( .B1(n11146), .B2(P2_IR_REG_0__SCAN_IN), .A(n7180), .ZN(
        n14110) );
  NAND2_X2 U10068 ( .A1(n8298), .A2(n8297), .ZN(n14817) );
  NAND2_X1 U10069 ( .A1(n7377), .A2(n7379), .ZN(n13459) );
  AND2_X1 U10070 ( .A1(n7374), .A2(n13665), .ZN(n7378) );
  NAND2_X2 U10071 ( .A1(n13375), .A2(n13374), .ZN(n12246) );
  NAND2_X1 U10072 ( .A1(n7131), .A2(n7130), .ZN(n8689) );
  OR2_X1 U10073 ( .A1(n16011), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n7130) );
  NAND2_X1 U10074 ( .A1(n14851), .A2(n16011), .ZN(n7131) );
  NAND2_X2 U10075 ( .A1(n8036), .A2(n10696), .ZN(n8420) );
  NOR2_X1 U10076 ( .A1(n15322), .A2(n13019), .ZN(n15325) );
  AND2_X2 U10077 ( .A1(n7222), .A2(n7221), .ZN(n12555) );
  NAND2_X1 U10078 ( .A1(n8474), .A2(n8473), .ZN(n7199) );
  NAND2_X1 U10079 ( .A1(n12716), .A2(n15092), .ZN(n7221) );
  NAND2_X2 U10080 ( .A1(n9650), .A2(n9649), .ZN(n12560) );
  NAND2_X1 U10081 ( .A1(n12742), .A2(n12741), .ZN(n12740) );
  NAND2_X1 U10082 ( .A1(n10125), .A2(n10124), .ZN(n10133) );
  NAND2_X1 U10083 ( .A1(n12147), .A2(n12146), .ZN(n12145) );
  XNOR2_X1 U10084 ( .A(n7135), .B(n7134), .ZN(n15071) );
  BUF_X1 U10085 ( .A(n15810), .Z(n7132) );
  NAND2_X1 U10086 ( .A1(n7934), .A2(n7936), .ZN(n12147) );
  NAND2_X1 U10087 ( .A1(n7228), .A2(n7963), .ZN(n12742) );
  NAND2_X1 U10088 ( .A1(n13094), .A2(n13095), .ZN(n13093) );
  NAND2_X1 U10089 ( .A1(n11351), .A2(n11350), .ZN(n11349) );
  NAND2_X1 U10090 ( .A1(n11753), .A2(n10162), .ZN(n12079) );
  NAND2_X1 U10091 ( .A1(n12409), .A2(n7964), .ZN(n7228) );
  AOI22_X1 U10092 ( .A1(n12032), .A2(n15843), .B1(n12031), .B2(n12030), .ZN(
        n12033) );
  NAND2_X2 U10093 ( .A1(n9551), .A2(n9550), .ZN(n12028) );
  NAND2_X2 U10094 ( .A1(n13011), .A2(n7799), .ZN(n15383) );
  NAND2_X1 U10095 ( .A1(n11848), .A2(n11859), .ZN(n11849) );
  INV_X2 U10096 ( .A(n11476), .ZN(n7136) );
  NAND2_X1 U10097 ( .A1(n7220), .A2(n7219), .ZN(n11800) );
  NOR2_X1 U10098 ( .A1(n7498), .A2(P3_ADDR_REG_4__SCAN_IN), .ZN(n7497) );
  NAND2_X2 U10099 ( .A1(n12022), .A2(n12021), .ZN(n12196) );
  NAND2_X1 U10100 ( .A1(n8096), .A2(n10703), .ZN(n7189) );
  NAND2_X1 U10101 ( .A1(n14559), .A2(n8504), .ZN(n8506) );
  NAND2_X1 U10102 ( .A1(n11624), .A2(n8055), .ZN(n11672) );
  INV_X1 U10103 ( .A(n7185), .ZN(n7184) );
  NAND2_X1 U10104 ( .A1(n7525), .A2(n7523), .ZN(n14244) );
  NAND3_X1 U10105 ( .A1(n7522), .A2(n14227), .A3(n14228), .ZN(n7521) );
  NAND3_X1 U10106 ( .A1(n14210), .A2(n14208), .A3(n14209), .ZN(n7143) );
  NAND2_X1 U10107 ( .A1(n7144), .A2(n14092), .ZN(P2_U3212) );
  NAND2_X1 U10108 ( .A1(n7145), .A2(n14065), .ZN(n7144) );
  NAND2_X1 U10109 ( .A1(n7187), .A2(n14083), .ZN(n7145) );
  NAND2_X1 U10110 ( .A1(n8956), .A2(n8955), .ZN(n8972) );
  NAND2_X1 U10111 ( .A1(n9061), .A2(n9060), .ZN(n9073) );
  NAND2_X1 U10112 ( .A1(n13484), .A2(n13483), .ZN(n7262) );
  NAND2_X1 U10113 ( .A1(n9076), .A2(n9075), .ZN(n9105) );
  NAND2_X1 U10114 ( .A1(n10077), .A2(n13458), .ZN(n10575) );
  NAND2_X1 U10115 ( .A1(n7216), .A2(n7215), .ZN(n10579) );
  NAND3_X2 U10116 ( .A1(n8909), .A2(n8910), .A3(n7150), .ZN(n16030) );
  AND2_X1 U10117 ( .A1(n8908), .A2(n8911), .ZN(n7150) );
  NAND3_X1 U10118 ( .A1(n12101), .A2(n12102), .A3(n13313), .ZN(n8986) );
  NAND2_X1 U10119 ( .A1(n11974), .A2(n13509), .ZN(n13358) );
  NAND2_X1 U10120 ( .A1(n13009), .A2(n13008), .ZN(n15435) );
  INV_X1 U10121 ( .A(n10637), .ZN(n7802) );
  NAND2_X1 U10122 ( .A1(n15670), .A2(n15886), .ZN(n7152) );
  INV_X1 U10123 ( .A(n7154), .ZN(n7153) );
  AOI21_X1 U10124 ( .B1(n7788), .B2(n7789), .A(n6693), .ZN(n7785) );
  INV_X1 U10125 ( .A(n12337), .ZN(n7206) );
  NAND2_X1 U10126 ( .A1(n7152), .A2(n7151), .ZN(P1_U3555) );
  NAND2_X1 U10127 ( .A1(n12145), .A2(n10196), .ZN(n12409) );
  OAI21_X1 U10128 ( .B1(n7156), .B2(n15070), .A(n14984), .ZN(P1_U3225) );
  NAND2_X1 U10129 ( .A1(n7958), .A2(n7956), .ZN(n15040) );
  NAND2_X1 U10130 ( .A1(n7660), .A2(n11688), .ZN(n11691) );
  NAND2_X1 U10131 ( .A1(n14668), .A2(n8363), .ZN(n14655) );
  NAND2_X1 U10132 ( .A1(n15668), .A2(n15886), .ZN(n7203) );
  INV_X1 U10133 ( .A(n7983), .ZN(n7367) );
  INV_X1 U10134 ( .A(n7509), .ZN(n15709) );
  INV_X1 U10135 ( .A(n10646), .ZN(n7498) );
  NAND2_X1 U10136 ( .A1(n7496), .A2(n7495), .ZN(n7494) );
  OAI21_X1 U10137 ( .B1(n8901), .B2(n16014), .A(n7164), .ZN(P3_U3201) );
  NAND3_X1 U10138 ( .A1(n7699), .A2(n7700), .A3(n6714), .ZN(n7702) );
  AND2_X1 U10139 ( .A1(n7711), .A2(n13582), .ZN(n7709) );
  NAND2_X1 U10140 ( .A1(n14649), .A2(n8631), .ZN(n14623) );
  NAND2_X1 U10141 ( .A1(n11768), .A2(n11772), .ZN(n11767) );
  NAND2_X1 U10142 ( .A1(n11672), .A2(n11671), .ZN(n11670) );
  NAND2_X1 U10143 ( .A1(n8106), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n8144) );
  INV_X1 U10144 ( .A(n7682), .ZN(n7681) );
  NAND2_X1 U10145 ( .A1(n7225), .A2(n10043), .ZN(n7965) );
  NAND2_X1 U10146 ( .A1(n12027), .A2(n12026), .ZN(n12034) );
  NAND2_X1 U10147 ( .A1(n15557), .A2(n15850), .ZN(n7173) );
  NAND2_X1 U10148 ( .A1(n9514), .A2(n15707), .ZN(n7443) );
  NAND2_X1 U10149 ( .A1(n15484), .A2(n13031), .ZN(n13033) );
  NAND4_X1 U10150 ( .A1(n8692), .A2(n8691), .A3(n8723), .A4(n8690), .ZN(n7174)
         );
  NAND2_X1 U10151 ( .A1(n12554), .A2(n12726), .ZN(n7222) );
  NAND2_X1 U10152 ( .A1(n7807), .A2(n6637), .ZN(n7225) );
  NAND4_X1 U10153 ( .A1(n8696), .A2(n7263), .A3(n7862), .A4(n7568), .ZN(n7176)
         );
  NAND2_X1 U10154 ( .A1(n10392), .A2(n8562), .ZN(n14518) );
  XNOR2_X2 U10155 ( .A(n8040), .B(n8039), .ZN(n11772) );
  NAND2_X1 U10156 ( .A1(n12185), .A2(n8172), .ZN(n12374) );
  NAND2_X1 U10157 ( .A1(n7197), .A2(n6726), .ZN(n8476) );
  INV_X1 U10158 ( .A(n7618), .ZN(n7617) );
  AND2_X2 U10159 ( .A1(n11800), .A2(n9537), .ZN(n11958) );
  NAND2_X1 U10160 ( .A1(n7332), .A2(n12020), .ZN(n15798) );
  INV_X1 U10161 ( .A(n14002), .ZN(n7761) );
  INV_X2 U10162 ( .A(n8099), .ZN(n7193) );
  NAND2_X1 U10163 ( .A1(n8656), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8022) );
  NOR2_X1 U10164 ( .A1(n8745), .A2(n8981), .ZN(n8746) );
  INV_X1 U10165 ( .A(n7345), .ZN(n7344) );
  NAND2_X1 U10166 ( .A1(n7203), .A2(n7202), .ZN(P1_U3557) );
  NAND2_X1 U10167 ( .A1(n10159), .A2(n10158), .ZN(n11753) );
  NAND2_X1 U10168 ( .A1(n7214), .A2(n7213), .ZN(n9654) );
  INV_X1 U10169 ( .A(n14933), .ZN(n10249) );
  OAI21_X1 U10170 ( .B1(n9474), .B2(P1_IR_REG_19__SCAN_IN), .A(n7201), .ZN(
        n9480) );
  NAND2_X1 U10171 ( .A1(n7949), .A2(n7955), .ZN(n14979) );
  OAI211_X1 U10172 ( .C1(n9743), .C2(n11483), .A(n7241), .B(n11793), .ZN(n9522) );
  NAND2_X1 U10173 ( .A1(n7204), .A2(n7781), .ZN(n12215) );
  NAND2_X1 U10174 ( .A1(n12034), .A2(n7223), .ZN(n7204) );
  NAND2_X1 U10175 ( .A1(n12216), .A2(n7206), .ZN(n7205) );
  XNOR2_X2 U10176 ( .A(n7208), .B(n9466), .ZN(n9780) );
  NAND2_X1 U10177 ( .A1(n7630), .A2(n7629), .ZN(n7628) );
  OR2_X1 U10178 ( .A1(n8388), .A2(n11751), .ZN(n8404) );
  NAND2_X1 U10179 ( .A1(n8404), .A2(n8389), .ZN(n8390) );
  NAND2_X1 U10180 ( .A1(n10579), .A2(n9347), .ZN(n9362) );
  INV_X1 U10181 ( .A(n10577), .ZN(n7216) );
  NAND2_X1 U10182 ( .A1(n15668), .A2(n15877), .ZN(n7452) );
  NAND2_X1 U10184 ( .A1(n7611), .A2(n7612), .ZN(n9350) );
  NAND2_X1 U10185 ( .A1(n11955), .A2(n11958), .ZN(n11954) );
  INV_X1 U10186 ( .A(n10677), .ZN(n7496) );
  NAND2_X1 U10187 ( .A1(n7452), .A2(n6735), .ZN(P1_U3525) );
  NAND2_X1 U10188 ( .A1(n14623), .A2(n8632), .ZN(n7362) );
  NAND2_X1 U10189 ( .A1(n10078), .A2(n9336), .ZN(n10577) );
  OR2_X2 U10190 ( .A1(n13508), .A2(n12099), .ZN(n13359) );
  NOR2_X2 U10191 ( .A1(n10341), .A2(n14922), .ZN(n10374) );
  OAI21_X2 U10192 ( .B1(n15011), .B2(n7946), .A(n7943), .ZN(n14923) );
  INV_X8 U10193 ( .A(n10695), .ZN(n10696) );
  NAND2_X1 U10194 ( .A1(n7710), .A2(n7709), .ZN(n7717) );
  NAND2_X1 U10195 ( .A1(n7283), .A2(n7281), .ZN(n7876) );
  NAND2_X1 U10196 ( .A1(n7876), .A2(n8269), .ZN(n8310) );
  INV_X1 U10197 ( .A(n7782), .ZN(n7781) );
  INV_X1 U10198 ( .A(n15435), .ZN(n7226) );
  NAND2_X1 U10199 ( .A1(n12079), .A2(n7935), .ZN(n7934) );
  NAND2_X1 U10200 ( .A1(n15030), .A2(n10239), .ZN(n15031) );
  NAND2_X1 U10201 ( .A1(n12336), .A2(n7788), .ZN(n7786) );
  OAI21_X1 U10202 ( .B1(n7784), .B2(n12211), .A(n15776), .ZN(n7782) );
  AND2_X1 U10203 ( .A1(n8745), .A2(n8981), .ZN(n7229) );
  NAND2_X1 U10204 ( .A1(n8801), .A2(n8803), .ZN(n8804) );
  NAND2_X1 U10205 ( .A1(n7583), .A2(n7581), .ZN(n9018) );
  NAND2_X1 U10206 ( .A1(n7230), .A2(n9304), .ZN(n9321) );
  NAND2_X1 U10207 ( .A1(n7579), .A2(n7580), .ZN(n7230) );
  NAND2_X1 U10208 ( .A1(n7261), .A2(n7372), .ZN(P3_U3296) );
  NOR2_X1 U10209 ( .A1(n7376), .A2(n7375), .ZN(n7374) );
  NAND2_X1 U10210 ( .A1(n7231), .A2(n13469), .ZN(n13466) );
  NAND2_X1 U10211 ( .A1(n13467), .A2(n7232), .ZN(n7231) );
  NAND2_X1 U10212 ( .A1(n8588), .A2(n8587), .ZN(n11629) );
  INV_X1 U10213 ( .A(n11741), .ZN(n7756) );
  INV_X4 U10214 ( .A(n10436), .ZN(n13112) );
  NAND2_X1 U10215 ( .A1(n8039), .A2(n14110), .ZN(n11769) );
  OAI211_X1 U10216 ( .C1(n14747), .C2(n16000), .A(n14746), .B(n14745), .ZN(
        n14850) );
  INV_X1 U10217 ( .A(n8764), .ZN(n8765) );
  AOI21_X2 U10218 ( .B1(n11265), .B2(n11266), .A(n11267), .ZN(n11264) );
  INV_X1 U10219 ( .A(n9571), .ZN(n7239) );
  NAND2_X1 U10220 ( .A1(n7786), .A2(n7785), .ZN(n12559) );
  NAND2_X1 U10221 ( .A1(n7557), .A2(n7252), .ZN(n12266) );
  NAND2_X1 U10222 ( .A1(n7560), .A2(n12098), .ZN(n7252) );
  NAND2_X1 U10223 ( .A1(n7253), .A2(n7549), .ZN(n12403) );
  NAND2_X1 U10224 ( .A1(n13742), .A2(n13745), .ZN(n13741) );
  AND2_X2 U10225 ( .A1(n8708), .A2(n8722), .ZN(n7263) );
  NAND2_X1 U10226 ( .A1(n7270), .A2(n10485), .ZN(n10486) );
  NAND2_X1 U10227 ( .A1(n7277), .A2(n7274), .ZN(n7270) );
  NAND2_X1 U10228 ( .A1(n8231), .A2(n7284), .ZN(n7283) );
  OAI21_X1 U10229 ( .B1(n8231), .B2(n7287), .A(n7284), .ZN(n8268) );
  AOI21_X1 U10230 ( .B1(n7284), .B2(n7287), .A(n7282), .ZN(n7281) );
  INV_X1 U10231 ( .A(n14084), .ZN(n7291) );
  NAND3_X1 U10232 ( .A1(n7295), .A2(n7294), .A3(n6701), .ZN(n7293) );
  NAND2_X1 U10233 ( .A1(n14265), .A2(n14107), .ZN(n7298) );
  NAND3_X1 U10234 ( .A1(n7298), .A2(n14109), .A3(n7296), .ZN(n14112) );
  AND2_X1 U10235 ( .A1(n7299), .A2(n7300), .ZN(n14197) );
  NAND4_X1 U10236 ( .A1(n14167), .A2(n14166), .A3(n7301), .A4(n6705), .ZN(
        n7299) );
  OAI21_X1 U10237 ( .B1(n6651), .B2(n7312), .A(n7311), .ZN(n14156) );
  OR2_X1 U10238 ( .A1(n7529), .A2(n14150), .ZN(n7320) );
  NAND2_X1 U10239 ( .A1(n9202), .A2(n6729), .ZN(n9248) );
  NAND2_X1 U10240 ( .A1(n8988), .A2(n7325), .ZN(n9065) );
  NAND3_X1 U10241 ( .A1(n8943), .A2(n11684), .A3(n8942), .ZN(n9009) );
  NAND3_X1 U10242 ( .A1(n13665), .A2(n13458), .A3(n7331), .ZN(n7330) );
  NAND2_X1 U10243 ( .A1(n15798), .A2(n15799), .ZN(n12022) );
  NAND2_X1 U10244 ( .A1(n12019), .A2(n12018), .ZN(n7332) );
  INV_X1 U10245 ( .A(n11798), .ZN(n7348) );
  NAND2_X1 U10246 ( .A1(n8063), .A2(n8064), .ZN(n8088) );
  NAND3_X1 U10247 ( .A1(n7351), .A2(n8049), .A3(SI_1_), .ZN(n7350) );
  NAND2_X1 U10248 ( .A1(n8048), .A2(n8047), .ZN(n7352) );
  OAI21_X1 U10249 ( .B1(n7886), .B2(n8412), .A(n7353), .ZN(n8388) );
  NAND2_X1 U10250 ( .A1(n7358), .A2(n7356), .ZN(n7355) );
  NAND2_X1 U10251 ( .A1(n7365), .A2(n7285), .ZN(n7364) );
  NAND2_X1 U10252 ( .A1(n7368), .A2(n13357), .ZN(n13363) );
  NAND2_X1 U10253 ( .A1(n7369), .A2(n13353), .ZN(n7368) );
  NAND4_X1 U10254 ( .A1(n13349), .A2(n13350), .A3(n7371), .A4(n7370), .ZN(
        n7369) );
  NAND2_X1 U10255 ( .A1(n13344), .A2(n6696), .ZN(n7370) );
  NAND2_X1 U10256 ( .A1(n13344), .A2(n6704), .ZN(n7371) );
  INV_X1 U10257 ( .A(n7381), .ZN(n7376) );
  NAND3_X1 U10258 ( .A1(n13447), .A2(n6698), .A3(n7380), .ZN(n7379) );
  NAND2_X1 U10259 ( .A1(n13386), .A2(n6709), .ZN(n7382) );
  NAND2_X1 U10260 ( .A1(n7382), .A2(n7383), .ZN(n13409) );
  NAND2_X1 U10261 ( .A1(n13413), .A2(n7392), .ZN(n7390) );
  NAND2_X1 U10262 ( .A1(n7390), .A2(n7391), .ZN(n13430) );
  NAND2_X1 U10263 ( .A1(n11303), .A2(n7410), .ZN(n7404) );
  NAND2_X1 U10264 ( .A1(n7408), .A2(n7404), .ZN(n11250) );
  NAND4_X1 U10265 ( .A1(n7568), .A2(n7411), .A3(n8708), .A4(n8696), .ZN(n7413)
         );
  OAI21_X1 U10266 ( .B1(n13519), .B2(n7425), .A(n7422), .ZN(n8888) );
  NAND2_X1 U10267 ( .A1(n7446), .A2(n9514), .ZN(n7445) );
  NOR2_X1 U10268 ( .A1(n10751), .A2(n9991), .ZN(n7446) );
  NAND2_X1 U10269 ( .A1(n7449), .A2(n7448), .ZN(n7447) );
  NAND2_X1 U10270 ( .A1(n13203), .A2(n7463), .ZN(n7462) );
  OAI211_X1 U10271 ( .C1(n13203), .C2(n7464), .A(n7462), .B(n13211), .ZN(
        P3_U3169) );
  XNOR2_X1 U10272 ( .A(n13203), .B(n13204), .ZN(n13205) );
  NAND3_X1 U10273 ( .A1(n11606), .A2(n11605), .A3(n11912), .ZN(n7486) );
  NOR2_X1 U10274 ( .A1(n11656), .A2(n7488), .ZN(n7487) );
  NAND2_X1 U10275 ( .A1(n12935), .A2(n7491), .ZN(n7490) );
  NAND2_X1 U10276 ( .A1(n10628), .A2(n10646), .ZN(n10647) );
  NAND2_X1 U10277 ( .A1(n15765), .A2(n7501), .ZN(n7505) );
  NAND3_X1 U10278 ( .A1(n7502), .A2(n7503), .A3(P2_ADDR_REG_18__SCAN_IN), .ZN(
        n7501) );
  OR2_X1 U10279 ( .A1(n15764), .A2(n15749), .ZN(n7504) );
  XNOR2_X1 U10280 ( .A(n7505), .B(n15772), .ZN(SUB_1596_U4) );
  INV_X1 U10281 ( .A(n15751), .ZN(n7506) );
  INV_X1 U10282 ( .A(n14105), .ZN(n7517) );
  NAND2_X1 U10283 ( .A1(n7519), .A2(n7518), .ZN(n14235) );
  OR2_X1 U10284 ( .A1(n7521), .A2(n14229), .ZN(n7518) );
  NAND2_X1 U10285 ( .A1(n7520), .A2(n14230), .ZN(n7519) );
  NAND2_X1 U10286 ( .A1(n7521), .A2(n14229), .ZN(n7520) );
  NAND2_X1 U10287 ( .A1(n14240), .A2(n7526), .ZN(n7525) );
  OAI22_X2 U10288 ( .A1(n14156), .A2(n7535), .B1(n14157), .B2(n7534), .ZN(
        n14162) );
  NAND2_X1 U10289 ( .A1(n14162), .A2(n14163), .ZN(n14161) );
  NAND2_X1 U10290 ( .A1(n8571), .A2(n8570), .ZN(n7536) );
  NAND2_X1 U10291 ( .A1(n13351), .A2(n7538), .ZN(n13352) );
  OAI21_X2 U10292 ( .B1(n12765), .B2(n7542), .A(n7540), .ZN(n13796) );
  OAI21_X1 U10293 ( .B1(n7562), .B2(n7559), .A(n7558), .ZN(n7557) );
  OAI21_X1 U10294 ( .B1(n12098), .B2(n13313), .A(n13359), .ZN(n11867) );
  NAND4_X1 U10295 ( .A1(n8696), .A2(n8708), .A3(n6560), .A4(n8707), .ZN(n7570)
         );
  NAND2_X1 U10296 ( .A1(n7577), .A2(n8935), .ZN(n8951) );
  INV_X1 U10297 ( .A(n8934), .ZN(n7578) );
  NAND2_X1 U10298 ( .A1(n8972), .A2(n7585), .ZN(n7583) );
  NAND2_X1 U10299 ( .A1(n9156), .A2(n7591), .ZN(n7588) );
  NAND2_X1 U10300 ( .A1(n7598), .A2(n7599), .ZN(n9061) );
  NAND2_X1 U10301 ( .A1(n9239), .A2(n9238), .ZN(n7610) );
  NAND2_X1 U10302 ( .A1(n9321), .A2(n7613), .ZN(n7611) );
  INV_X1 U10303 ( .A(n11772), .ZN(n14331) );
  NAND2_X1 U10304 ( .A1(n8953), .A2(n8952), .ZN(n8980) );
  AOI21_X1 U10305 ( .B1(n13727), .B2(n13436), .A(n9412), .ZN(n13717) );
  OAI21_X2 U10306 ( .B1(n13717), .B2(n13312), .A(n13441), .ZN(n13707) );
  NAND2_X1 U10307 ( .A1(n16029), .A2(n13338), .ZN(n11643) );
  NAND2_X1 U10308 ( .A1(n11670), .A2(n8070), .ZN(n11815) );
  NAND2_X1 U10309 ( .A1(n9073), .A2(n9072), .ZN(n9088) );
  OR2_X1 U10310 ( .A1(n11264), .A2(n6619), .ZN(n7647) );
  NAND2_X1 U10311 ( .A1(n11264), .A2(n8962), .ZN(n7645) );
  NAND2_X1 U10312 ( .A1(n11244), .A2(P3_REG2_REG_5__SCAN_IN), .ZN(n11243) );
  NAND2_X1 U10313 ( .A1(n7661), .A2(n7663), .ZN(n11534) );
  NAND2_X2 U10314 ( .A1(n8025), .A2(n8024), .ZN(n14912) );
  NAND2_X1 U10315 ( .A1(n12189), .A2(n8603), .ZN(n8606) );
  INV_X1 U10316 ( .A(n8635), .ZN(n7687) );
  OAI22_X1 U10317 ( .A1(n8639), .A2(n6712), .B1(n7694), .B2(n7693), .ZN(n8641)
         );
  NAND2_X1 U10318 ( .A1(n8639), .A2(n8638), .ZN(n14526) );
  NAND2_X1 U10319 ( .A1(n11294), .A2(n7697), .ZN(n8815) );
  NAND2_X1 U10320 ( .A1(n11295), .A2(n11296), .ZN(n11294) );
  INV_X1 U10321 ( .A(n11271), .ZN(n7703) );
  OAI21_X1 U10322 ( .B1(n13566), .B2(n13565), .A(n13564), .ZN(n13563) );
  AOI21_X1 U10323 ( .B1(n13565), .B2(n13564), .A(n7714), .ZN(n7711) );
  OAI21_X1 U10324 ( .B1(n13564), .B2(n7714), .A(n11126), .ZN(n7713) );
  INV_X1 U10325 ( .A(n13565), .ZN(n7716) );
  NAND2_X1 U10326 ( .A1(n11245), .A2(n6641), .ZN(n7719) );
  INV_X1 U10327 ( .A(n7727), .ZN(n7725) );
  NAND2_X1 U10328 ( .A1(n7729), .A2(n7731), .ZN(n7727) );
  OAI22_X1 U10329 ( .A1(n11696), .A2(n7722), .B1(n8867), .B2(n7726), .ZN(n7724) );
  NAND2_X1 U10330 ( .A1(n11535), .A2(n6579), .ZN(n7728) );
  INV_X1 U10331 ( .A(n7723), .ZN(n10593) );
  OAI21_X1 U10332 ( .B1(n7727), .B2(n11535), .A(n7724), .ZN(n7723) );
  NAND2_X1 U10333 ( .A1(n7728), .A2(n7729), .ZN(n11700) );
  NAND2_X1 U10334 ( .A1(n8820), .A2(n6595), .ZN(n7733) );
  NAND2_X1 U10335 ( .A1(n8820), .A2(n12601), .ZN(n13523) );
  INV_X1 U10336 ( .A(n8821), .ZN(n7736) );
  NOR2_X2 U10337 ( .A1(n7739), .A2(n7740), .ZN(n14818) );
  NAND3_X1 U10338 ( .A1(n7748), .A2(n7744), .A3(n7742), .ZN(P2_U3192) );
  NAND2_X1 U10339 ( .A1(n7743), .A2(n6576), .ZN(n7742) );
  OAI21_X1 U10340 ( .B1(n11740), .B2(n7757), .A(n7755), .ZN(n11978) );
  AOI21_X1 U10341 ( .B1(n7755), .B2(n7757), .A(n7754), .ZN(n7753) );
  OAI21_X1 U10342 ( .B1(n10508), .B2(n7764), .A(n7763), .ZN(n14003) );
  AOI21_X1 U10343 ( .B1(n7763), .B2(n7764), .A(n7761), .ZN(n7760) );
  NAND3_X1 U10344 ( .A1(n7769), .A2(n7772), .A3(n7775), .ZN(n7768) );
  NAND2_X1 U10345 ( .A1(n12034), .A2(n12033), .ZN(n12212) );
  INV_X1 U10346 ( .A(n12565), .ZN(n12566) );
  NAND2_X1 U10347 ( .A1(n12565), .A2(n12999), .ZN(n7793) );
  NAND2_X1 U10348 ( .A1(n15383), .A2(n13013), .ZN(n13016) );
  OAI21_X2 U10349 ( .B1(n15288), .B2(n7805), .A(n7804), .ZN(n15268) );
  INV_X1 U10350 ( .A(n7806), .ZN(n7805) );
  NAND2_X1 U10351 ( .A1(n13038), .A2(n7820), .ZN(n7819) );
  NAND2_X1 U10352 ( .A1(n7823), .A2(n7822), .ZN(n13052) );
  CLKBUF_X1 U10353 ( .A(n9514), .Z(n7827) );
  OR2_X1 U10354 ( .A1(n9514), .A2(n9518), .ZN(n9519) );
  INV_X2 U10355 ( .A(n9514), .ZN(n9781) );
  NAND2_X1 U10356 ( .A1(n15706), .A2(n7827), .ZN(n15370) );
  NAND2_X1 U10357 ( .A1(n12699), .A2(n7840), .ZN(n7839) );
  NAND2_X1 U10358 ( .A1(n9319), .A2(n6654), .ZN(n10078) );
  INV_X1 U10359 ( .A(n12499), .ZN(n7844) );
  NAND2_X1 U10360 ( .A1(n12113), .A2(n9055), .ZN(n7845) );
  NAND2_X1 U10361 ( .A1(n12963), .A2(n7855), .ZN(n7852) );
  NAND2_X1 U10362 ( .A1(n7852), .A2(n7853), .ZN(n13139) );
  NAND2_X1 U10363 ( .A1(n12963), .A2(n7858), .ZN(n7854) );
  NAND2_X1 U10364 ( .A1(n12963), .A2(n12962), .ZN(n13203) );
  OAI21_X2 U10365 ( .B1(n13186), .B2(n12943), .A(n12944), .ZN(n13195) );
  NAND2_X1 U10366 ( .A1(n6557), .A2(n7861), .ZN(n13960) );
  OAI21_X1 U10367 ( .B1(n9942), .B2(n9954), .A(n7869), .ZN(n9977) );
  NAND2_X1 U10368 ( .A1(n9942), .A2(n9941), .ZN(n15265) );
  NAND2_X1 U10369 ( .A1(n9976), .A2(n9977), .ZN(n7864) );
  NAND2_X1 U10370 ( .A1(n7864), .A2(n7871), .ZN(n9989) );
  NAND2_X1 U10371 ( .A1(n8344), .A2(n8343), .ZN(n7886) );
  NAND2_X1 U10372 ( .A1(n8477), .A2(n7896), .ZN(n7895) );
  NAND2_X1 U10373 ( .A1(n7892), .A2(n6727), .ZN(n8510) );
  NAND3_X1 U10374 ( .A1(n8493), .A2(n7893), .A3(n7895), .ZN(n7892) );
  INV_X1 U10375 ( .A(n8478), .ZN(n7896) );
  INV_X1 U10376 ( .A(n12225), .ZN(n7898) );
  NAND3_X1 U10377 ( .A1(n7898), .A2(n12241), .A3(n7897), .ZN(n12188) );
  NAND2_X1 U10378 ( .A1(n7903), .A2(n7901), .ZN(n13129) );
  NAND2_X1 U10379 ( .A1(n9654), .A2(n9655), .ZN(n9653) );
  AOI21_X1 U10380 ( .B1(n9571), .B2(n7920), .A(n7918), .ZN(n7917) );
  INV_X1 U10381 ( .A(n9824), .ZN(n7931) );
  INV_X1 U10382 ( .A(n10179), .ZN(n7940) );
  OAI211_X1 U10383 ( .C1(n7938), .C2(n7155), .A(n7937), .B(n7942), .ZN(n12177)
         );
  NAND2_X1 U10384 ( .A1(n7940), .A2(n7941), .ZN(n7937) );
  INV_X1 U10385 ( .A(n14923), .ZN(n10341) );
  NAND2_X1 U10386 ( .A1(n10325), .A2(n10324), .ZN(n7954) );
  NAND2_X1 U10387 ( .A1(n14959), .A2(n10303), .ZN(n7958) );
  NAND2_X1 U10388 ( .A1(n12740), .A2(n6702), .ZN(n15030) );
  OR2_X1 U10389 ( .A1(n9372), .A2(n8929), .ZN(n8930) );
  NAND2_X1 U10390 ( .A1(n10556), .A2(n14065), .ZN(n10573) );
  CLKBUF_X1 U10391 ( .A(n15484), .Z(n15486) );
  NAND2_X1 U10392 ( .A1(n8736), .A2(P3_IR_REG_1__SCAN_IN), .ZN(n8738) );
  INV_X1 U10393 ( .A(n8974), .ZN(n9357) );
  OR2_X1 U10394 ( .A1(n8658), .A2(n8652), .ZN(n8661) );
  OAI21_X1 U10395 ( .B1(n13124), .B2(n10573), .A(n10572), .ZN(P2_U3186) );
  NAND2_X1 U10396 ( .A1(n10027), .A2(n9503), .ZN(n11802) );
  OR2_X1 U10397 ( .A1(n14547), .A2(n14546), .ZN(n14758) );
  NAND2_X1 U10398 ( .A1(n10577), .A2(n13469), .ZN(n10578) );
  OR2_X1 U10399 ( .A1(n9311), .A2(n16064), .ZN(n8909) );
  OR2_X1 U10400 ( .A1(n11350), .A2(n11474), .ZN(n10132) );
  NAND2_X1 U10401 ( .A1(n9502), .A2(n9635), .ZN(n9505) );
  OAI21_X1 U10402 ( .B1(n8023), .B2(n8006), .A(P2_IR_REG_28__SCAN_IN), .ZN(
        n8019) );
  NAND2_X1 U10403 ( .A1(n9501), .A2(n11801), .ZN(n9502) );
  NAND2_X1 U10404 ( .A1(n9774), .A2(n7968), .ZN(n9775) );
  OR2_X1 U10405 ( .A1(n15314), .A2(n6550), .ZN(n9889) );
  OR2_X1 U10406 ( .A1(n15013), .A2(n6550), .ZN(n9858) );
  INV_X1 U10407 ( .A(n6550), .ZN(n9913) );
  OR2_X1 U10408 ( .A1(n6550), .A2(n12041), .ZN(n9494) );
  OR2_X1 U10409 ( .A1(n9957), .A2(n15100), .ZN(n9491) );
  OR2_X1 U10410 ( .A1(n15394), .A2(n6550), .ZN(n9456) );
  INV_X1 U10411 ( .A(n12987), .ZN(n10400) );
  OR2_X1 U10412 ( .A1(n10123), .A2(n11483), .ZN(n11801) );
  NAND2_X1 U10413 ( .A1(n10559), .A2(n10555), .ZN(n14103) );
  AND2_X1 U10414 ( .A1(n12267), .A2(n13373), .ZN(n7966) );
  NAND2_X1 U10415 ( .A1(n15780), .A2(n12199), .ZN(n7967) );
  AND4_X1 U10416 ( .A1(n13029), .A2(n9954), .A3(n15502), .A4(n10036), .ZN(
        n7968) );
  INV_X1 U10417 ( .A(n13824), .ZN(n9427) );
  INV_X2 U10418 ( .A(n16103), .ZN(n16106) );
  INV_X1 U10419 ( .A(n8008), .ZN(n14899) );
  OR2_X1 U10420 ( .A1(n9367), .A2(n11278), .ZN(n7969) );
  AND2_X1 U10421 ( .A1(n10284), .A2(n10283), .ZN(n7971) );
  OR2_X1 U10422 ( .A1(n14746), .A2(n14738), .ZN(n7972) );
  OR2_X1 U10423 ( .A1(n14747), .A2(n14742), .ZN(n7973) );
  OR2_X1 U10424 ( .A1(n14853), .A2(n14840), .ZN(n7974) );
  AND2_X1 U10425 ( .A1(n13323), .A2(n12448), .ZN(n7976) );
  OR2_X1 U10426 ( .A1(n16106), .A2(P3_REG1_REG_29__SCAN_IN), .ZN(n7977) );
  INV_X1 U10427 ( .A(n13758), .ZN(n9209) );
  AND2_X1 U10428 ( .A1(n8269), .A2(n8256), .ZN(n7978) );
  OR2_X1 U10429 ( .A1(n13562), .A2(n9130), .ZN(n7979) );
  OR2_X1 U10430 ( .A1(n14790), .A2(n14402), .ZN(n7980) );
  AND2_X1 U10431 ( .A1(n13666), .A2(n16049), .ZN(n7981) );
  AND2_X1 U10432 ( .A1(n13126), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n7982) );
  INV_X1 U10433 ( .A(P3_IR_REG_30__SCAN_IN), .ZN(n13961) );
  AND2_X1 U10434 ( .A1(n8253), .A2(n8234), .ZN(n7983) );
  XNOR2_X1 U10435 ( .A(n13076), .B(n10046), .ZN(n13068) );
  INV_X1 U10436 ( .A(n13068), .ZN(n13067) );
  AND2_X1 U10437 ( .A1(n9931), .A2(n9930), .ZN(n7986) );
  INV_X1 U10438 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n9443) );
  OR2_X1 U10439 ( .A1(n13601), .A2(n13876), .ZN(n7987) );
  AND2_X1 U10440 ( .A1(n8330), .A2(n8319), .ZN(n7988) );
  INV_X1 U10441 ( .A(n15869), .ZN(n12207) );
  XNOR2_X1 U10442 ( .A(n15341), .B(n15306), .ZN(n15326) );
  INV_X1 U10443 ( .A(n15326), .ZN(n13019) );
  AND2_X1 U10444 ( .A1(n15292), .A2(n15289), .ZN(n7990) );
  AND2_X1 U10445 ( .A1(n13051), .A2(n13050), .ZN(n7991) );
  XNOR2_X1 U10446 ( .A(n15318), .B(n15330), .ZN(n15311) );
  INV_X1 U10447 ( .A(n15311), .ZN(n13021) );
  NAND2_X1 U10448 ( .A1(n11852), .A2(n15804), .ZN(n15528) );
  NAND2_X1 U10449 ( .A1(n14126), .A2(n14125), .ZN(n14127) );
  NAND2_X1 U10450 ( .A1(n9505), .A2(n9504), .ZN(n9521) );
  OR2_X1 U10451 ( .A1(n15416), .A2(n9804), .ZN(n9805) );
  NAND2_X1 U10452 ( .A1(n14251), .A2(n14250), .ZN(n14252) );
  INV_X1 U10453 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n7997) );
  INV_X1 U10454 ( .A(n13458), .ZN(n9335) );
  AOI21_X1 U10455 ( .B1(n8437), .B2(n8436), .A(n8435), .ZN(n8438) );
  OR2_X1 U10456 ( .A1(n13899), .A2(n7128), .ZN(n9286) );
  NOR2_X1 U10457 ( .A1(P3_IR_REG_27__SCAN_IN), .A2(P3_IR_REG_26__SCAN_IN), 
        .ZN(n8803) );
  INV_X1 U10458 ( .A(n14040), .ZN(n10507) );
  NAND2_X1 U10459 ( .A1(n14311), .A2(n14310), .ZN(n14312) );
  AND2_X1 U10460 ( .A1(n12613), .A2(n8597), .ZN(n8596) );
  INV_X1 U10461 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n7995) );
  NAND2_X1 U10462 ( .A1(n10118), .A2(n11483), .ZN(n11793) );
  INV_X1 U10463 ( .A(P3_IR_REG_27__SCAN_IN), .ZN(n8802) );
  INV_X1 U10464 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n9170) );
  NAND2_X1 U10465 ( .A1(n9018), .A2(n8997), .ZN(n8999) );
  OAI21_X1 U10466 ( .B1(n14314), .B2(n14313), .A(n14312), .ZN(n14315) );
  INV_X1 U10467 ( .A(n14675), .ZN(n8640) );
  INV_X1 U10468 ( .A(n14536), .ZN(n8539) );
  INV_X1 U10469 ( .A(n14353), .ZN(n8306) );
  INV_X1 U10470 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n8236) );
  INV_X1 U10471 ( .A(n15502), .ZN(n13027) );
  OAI21_X1 U10472 ( .B1(n11336), .B2(P1_ADDR_REG_6__SCAN_IN), .A(n11335), .ZN(
        n11337) );
  OR2_X1 U10473 ( .A1(n12252), .A2(n12251), .ZN(n12255) );
  INV_X1 U10474 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n10785) );
  AND2_X1 U10475 ( .A1(n8823), .A2(n8822), .ZN(n8824) );
  INV_X1 U10476 ( .A(P3_IR_REG_20__SCAN_IN), .ZN(n8701) );
  NAND2_X1 U10477 ( .A1(n10674), .A2(P1_DATAO_REG_7__SCAN_IN), .ZN(n9029) );
  NAND2_X1 U10478 ( .A1(n10703), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n8952) );
  INV_X1 U10479 ( .A(n12300), .ZN(n10463) );
  INV_X1 U10480 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n8184) );
  INV_X1 U10481 ( .A(n12410), .ZN(n10201) );
  INV_X1 U10482 ( .A(n10342), .ZN(n10338) );
  INV_X1 U10483 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n12651) );
  INV_X1 U10484 ( .A(n13071), .ZN(n13066) );
  INV_X1 U10485 ( .A(n12340), .ZN(n15785) );
  NOR2_X1 U10486 ( .A1(n8414), .A2(SI_20_), .ZN(n8415) );
  NAND2_X1 U10487 ( .A1(n11651), .A2(n16031), .ZN(n11652) );
  AND2_X1 U10488 ( .A1(n11420), .A2(n11419), .ZN(n11441) );
  OR2_X1 U10489 ( .A1(n11421), .A2(n11440), .ZN(n13271) );
  AND2_X1 U10490 ( .A1(n8833), .A2(n8807), .ZN(n8831) );
  INV_X1 U10491 ( .A(n11431), .ZN(n13333) );
  INV_X1 U10492 ( .A(n9406), .ZN(n13315) );
  AND2_X1 U10493 ( .A1(n10091), .A2(n10090), .ZN(n11419) );
  AND2_X1 U10494 ( .A1(n9072), .A2(n9059), .ZN(n9060) );
  AND2_X1 U10495 ( .A1(n8955), .A2(n8954), .ZN(n8979) );
  NAND2_X1 U10496 ( .A1(n10559), .A2(n14375), .ZN(n14090) );
  AND2_X1 U10497 ( .A1(n8519), .A2(n8498), .ZN(n14563) );
  OAI21_X1 U10498 ( .B1(n12754), .B2(n14350), .A(n8617), .ZN(n12913) );
  XNOR2_X1 U10499 ( .A(n8601), .B(n15995), .ZN(n12232) );
  NAND2_X1 U10500 ( .A1(n6548), .A2(n10558), .ZN(n14698) );
  INV_X1 U10501 ( .A(n14086), .ZN(n14096) );
  OR2_X1 U10502 ( .A1(n8036), .A2(n8035), .ZN(n8037) );
  INV_X1 U10503 ( .A(n14818), .ZN(n14717) );
  OR2_X1 U10504 ( .A1(n10333), .A2(n10332), .ZN(n10334) );
  OR2_X1 U10505 ( .A1(n12097), .A2(n15824), .ZN(n11832) );
  NAND2_X1 U10506 ( .A1(n10384), .A2(n15072), .ZN(n10370) );
  OAI21_X1 U10507 ( .B1(n11476), .B2(n10348), .A(n10131), .ZN(n11350) );
  OR2_X1 U10508 ( .A1(n12900), .A2(n12901), .ZN(n14969) );
  INV_X1 U10509 ( .A(n10684), .ZN(n11830) );
  NAND2_X1 U10510 ( .A1(n13133), .A2(n10006), .ZN(n9942) );
  OR2_X1 U10511 ( .A1(n12551), .A2(n12550), .ZN(n12556) );
  INV_X1 U10512 ( .A(n15521), .ZN(n15431) );
  OR2_X1 U10513 ( .A1(n6556), .A2(n11832), .ZN(n15807) );
  INV_X1 U10514 ( .A(n12357), .ZN(n12359) );
  AND2_X1 U10515 ( .A1(n15721), .A2(P2_ADDR_REG_14__SCAN_IN), .ZN(n15719) );
  AND2_X1 U10516 ( .A1(n11441), .A2(n11440), .ZN(n13269) );
  NAND2_X1 U10517 ( .A1(n11425), .A2(n12707), .ZN(n13261) );
  AND2_X1 U10518 ( .A1(n8831), .A2(n8892), .ZN(n13631) );
  NAND2_X1 U10519 ( .A1(n9425), .A2(n9424), .ZN(n9426) );
  OR2_X1 U10520 ( .A1(n16066), .A2(n12503), .ZN(n9421) );
  INV_X1 U10521 ( .A(n13817), .ZN(n16046) );
  AND2_X1 U10522 ( .A1(n11708), .A2(n16038), .ZN(n16090) );
  OR2_X1 U10523 ( .A1(n16054), .A2(n16090), .ZN(n16070) );
  NOR2_X1 U10524 ( .A1(n8713), .A2(n8710), .ZN(n8711) );
  NAND2_X1 U10525 ( .A1(n9196), .A2(n9195), .ZN(n9212) );
  INV_X1 U10526 ( .A(P3_IR_REG_13__SCAN_IN), .ZN(n8774) );
  AND2_X1 U10527 ( .A1(n13115), .A2(n14065), .ZN(n13116) );
  AND3_X1 U10528 ( .A1(n12992), .A2(n12991), .A3(n12990), .ZN(n14317) );
  OR2_X1 U10529 ( .A1(n14574), .A2(n8648), .ZN(n8491) );
  INV_X1 U10530 ( .A(n15919), .ZN(n15936) );
  INV_X1 U10531 ( .A(n14698), .ZN(n14739) );
  AND2_X1 U10532 ( .A1(n6548), .A2(n8584), .ZN(n14703) );
  INV_X1 U10533 ( .A(n15989), .ZN(n15996) );
  INV_X1 U10534 ( .A(n16000), .ZN(n15993) );
  NOR2_X1 U10535 ( .A1(n10398), .A2(n8686), .ZN(n11634) );
  AND2_X1 U10536 ( .A1(n8678), .A2(n8683), .ZN(n15945) );
  AND2_X1 U10537 ( .A1(n11150), .A2(n12320), .ZN(n10566) );
  AND2_X1 U10538 ( .A1(n8240), .A2(n8270), .ZN(n11523) );
  NAND2_X1 U10539 ( .A1(n11829), .A2(n11832), .ZN(n15870) );
  INV_X1 U10540 ( .A(n15070), .ZN(n15072) );
  AND2_X1 U10541 ( .A1(n9835), .A2(n9834), .ZN(n15391) );
  NAND2_X1 U10542 ( .A1(n9524), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n9530) );
  AND2_X1 U10543 ( .A1(n11082), .A2(n11081), .ZN(n15244) );
  INV_X1 U10544 ( .A(n13074), .ZN(n13075) );
  INV_X1 U10545 ( .A(n13012), .ZN(n15416) );
  OR2_X1 U10546 ( .A1(n11474), .A2(n11473), .ZN(n11831) );
  INV_X1 U10547 ( .A(n15611), .ZN(n15826) );
  AND2_X1 U10548 ( .A1(n11470), .A2(n11829), .ZN(n11495) );
  NAND2_X1 U10549 ( .A1(n10355), .A2(n10356), .ZN(n11467) );
  AND2_X1 U10550 ( .A1(n9616), .A2(n9601), .ZN(n15163) );
  NAND2_X1 U10551 ( .A1(n15723), .A2(n15722), .ZN(n15724) );
  AND2_X1 U10552 ( .A1(n8833), .A2(n8832), .ZN(n16012) );
  INV_X1 U10553 ( .A(n13273), .ZN(n13226) );
  INV_X1 U10554 ( .A(n13309), .ZN(n13646) );
  INV_X1 U10555 ( .A(n13816), .ZN(n13499) );
  INV_X1 U10556 ( .A(n16021), .ZN(n13617) );
  INV_X1 U10557 ( .A(n13631), .ZN(n16015) );
  OR2_X1 U10558 ( .A1(n8810), .A2(n9366), .ZN(n16014) );
  OR2_X1 U10559 ( .A1(n16066), .A2(n16039), .ZN(n12629) );
  AND2_X1 U10560 ( .A1(n12629), .A2(n9421), .ZN(n13824) );
  NAND2_X1 U10561 ( .A1(n16106), .A2(n16070), .ZN(n13883) );
  NAND2_X1 U10562 ( .A1(n10110), .A2(n10109), .ZN(n16103) );
  INV_X1 U10563 ( .A(n10584), .ZN(n10585) );
  OR2_X1 U10564 ( .A1(n16092), .A2(n11790), .ZN(n13955) );
  AND2_X1 U10565 ( .A1(n10093), .A2(n10092), .ZN(n16092) );
  OR2_X1 U10566 ( .A1(n16092), .A2(n16055), .ZN(n13918) );
  INV_X1 U10567 ( .A(SI_16_), .ZN(n11211) );
  INV_X1 U10568 ( .A(SI_13_), .ZN(n11056) );
  INV_X1 U10569 ( .A(n14088), .ZN(n14099) );
  INV_X1 U10570 ( .A(n14101), .ZN(n14073) );
  OAI21_X1 U10571 ( .B1(n10402), .B2(n8648), .A(n8647), .ZN(n14393) );
  NAND2_X1 U10572 ( .A1(n8503), .A2(n8502), .ZN(n14397) );
  NAND2_X1 U10573 ( .A1(n13130), .A2(n14818), .ZN(n14510) );
  INV_X1 U10574 ( .A(n6548), .ZN(n14719) );
  OR2_X1 U10575 ( .A1(n14738), .A2(n12153), .ZN(n14682) );
  NAND2_X1 U10576 ( .A1(n16011), .A2(n15996), .ZN(n14840) );
  INV_X1 U10577 ( .A(n16011), .ZN(n16008) );
  INV_X1 U10578 ( .A(n14618), .ZN(n14869) );
  NAND2_X1 U10579 ( .A1(n16004), .A2(n15996), .ZN(n14892) );
  INV_X1 U10580 ( .A(n16004), .ZN(n16002) );
  AND2_X2 U10581 ( .A1(n11634), .A2(n11633), .ZN(n16004) );
  NOR2_X1 U10582 ( .A1(n15945), .A2(n15979), .ZN(n15960) );
  AND2_X1 U10583 ( .A1(n10566), .A2(P2_STATE_REG_SCAN_IN), .ZN(n15981) );
  INV_X1 U10584 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n11592) );
  INV_X1 U10585 ( .A(n15061), .ZN(n15077) );
  NAND3_X1 U10586 ( .A1(n15844), .A2(n10369), .A3(n10368), .ZN(n15070) );
  INV_X1 U10587 ( .A(n14927), .ZN(n15085) );
  OR2_X1 U10588 ( .A1(n11072), .A2(n15113), .ZN(n15248) );
  OR2_X1 U10589 ( .A1(n11852), .A2(n15250), .ZN(n15344) );
  OR2_X1 U10590 ( .A1(n6556), .A2(n11831), .ZN(n15535) );
  INV_X1 U10591 ( .A(n15886), .ZN(n15884) );
  INV_X1 U10592 ( .A(n15877), .ZN(n15876) );
  INV_X1 U10593 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n11590) );
  INV_X1 U10594 ( .A(n13510), .ZN(P3_U3897) );
  NAND4_X1 U10595 ( .A1(n7993), .A2(n8158), .A3(n7992), .A4(n10965), .ZN(n7994) );
  NOR2_X1 U10596 ( .A1(P2_IR_REG_12__SCAN_IN), .A2(P2_IR_REG_14__SCAN_IN), 
        .ZN(n7996) );
  NAND4_X1 U10597 ( .A1(n7996), .A2(n10785), .A3(n8236), .A4(n7995), .ZN(n8290) );
  NAND2_X1 U10598 ( .A1(n8294), .A2(n7997), .ZN(n7998) );
  NOR2_X1 U10599 ( .A1(P2_IR_REG_23__SCAN_IN), .A2(P2_IR_REG_26__SCAN_IN), 
        .ZN(n8000) );
  NOR2_X1 U10600 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_21__SCAN_IN), 
        .ZN(n7999) );
  NAND4_X1 U10601 ( .A1(n8000), .A2(n7999), .A3(n8575), .A4(n8567), .ZN(n8003)
         );
  INV_X1 U10602 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n8006) );
  NAND2_X1 U10603 ( .A1(n8021), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8007) );
  NAND2_X1 U10604 ( .A1(n8056), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n8012) );
  NAND2_X1 U10605 ( .A1(n8071), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n8011) );
  NAND2_X1 U10606 ( .A1(n8108), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n8010) );
  INV_X2 U10607 ( .A(n8096), .ZN(n10695) );
  NAND2_X1 U10608 ( .A1(n10696), .A2(SI_0_), .ZN(n8015) );
  INV_X1 U10609 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n8913) );
  NAND2_X1 U10610 ( .A1(n8015), .A2(n8913), .ZN(n8017) );
  AND2_X1 U10611 ( .A1(SI_0_), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n8016) );
  NAND2_X1 U10612 ( .A1(n8096), .A2(n8016), .ZN(n8031) );
  NAND2_X1 U10613 ( .A1(n8017), .A2(n8031), .ZN(n14920) );
  INV_X1 U10614 ( .A(n8023), .ZN(n8024) );
  NAND2_X1 U10615 ( .A1(n14421), .A2(n14108), .ZN(n11768) );
  NAND2_X1 U10616 ( .A1(n8108), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n8029) );
  INV_X1 U10617 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n11154) );
  AND2_X1 U10618 ( .A1(P2_DATAO_REG_0__SCAN_IN), .A2(SI_0_), .ZN(n8030) );
  INV_X1 U10619 ( .A(SI_1_), .ZN(n10731) );
  XNOR2_X1 U10620 ( .A(n8048), .B(n10731), .ZN(n8033) );
  MUX2_X1 U10621 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(P1_DATAO_REG_1__SCAN_IN), 
        .S(n8096), .Z(n8032) );
  XNOR2_X1 U10622 ( .A(n8033), .B(n8032), .ZN(n10751) );
  AND2_X2 U10623 ( .A1(n8036), .A2(n7218), .ZN(n8062) );
  NAND2_X1 U10624 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), 
        .ZN(n8034) );
  INV_X1 U10625 ( .A(n11155), .ZN(n8035) );
  INV_X1 U10626 ( .A(n8040), .ZN(n11453) );
  NAND2_X1 U10627 ( .A1(n11453), .A2(n8039), .ZN(n8041) );
  NAND2_X1 U10628 ( .A1(n11767), .A2(n8041), .ZN(n11626) );
  NAND2_X1 U10629 ( .A1(n8108), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n8045) );
  NAND2_X1 U10630 ( .A1(n8071), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n8043) );
  INV_X1 U10631 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n11157) );
  INV_X1 U10632 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n10656) );
  NAND2_X1 U10633 ( .A1(n8096), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n8046) );
  OAI211_X1 U10634 ( .C1(n8096), .C2(n10656), .A(n8046), .B(n10731), .ZN(n8047) );
  NAND2_X1 U10635 ( .A1(n8096), .A2(n10750), .ZN(n8049) );
  XNOR2_X1 U10636 ( .A(n8063), .B(n8064), .ZN(n10702) );
  NAND2_X1 U10637 ( .A1(n8062), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n8054) );
  NAND2_X1 U10638 ( .A1(n8067), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8052) );
  XNOR2_X1 U10639 ( .A(n8052), .B(P2_IR_REG_2__SCAN_IN), .ZN(n11158) );
  INV_X1 U10640 ( .A(n11158), .ZN(n8053) );
  OAI211_X2 U10641 ( .C1(n8420), .C2(n10702), .A(n8054), .B(n6621), .ZN(n14120) );
  INV_X1 U10642 ( .A(n14420), .ZN(n11570) );
  NAND2_X1 U10643 ( .A1(n11570), .A2(n7166), .ZN(n8055) );
  NAND2_X1 U10644 ( .A1(n12989), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n8061) );
  NAND2_X1 U10646 ( .A1(n8521), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n8060) );
  INV_X1 U10647 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n8057) );
  NAND2_X1 U10648 ( .A1(n8553), .A2(n8057), .ZN(n8059) );
  INV_X1 U10649 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n11159) );
  OR2_X1 U10650 ( .A1(n8376), .A2(n11159), .ZN(n8058) );
  INV_X1 U10651 ( .A(n8065), .ZN(n8066) );
  NAND2_X1 U10652 ( .A1(n8066), .A2(SI_2_), .ZN(n8085) );
  NAND2_X1 U10653 ( .A1(n8088), .A2(n8085), .ZN(n8080) );
  MUX2_X1 U10654 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(P1_DATAO_REG_3__SCAN_IN), 
        .S(n8096), .Z(n8089) );
  XNOR2_X1 U10655 ( .A(n8089), .B(SI_3_), .ZN(n8078) );
  XNOR2_X1 U10656 ( .A(n8080), .B(n8078), .ZN(n10637) );
  INV_X1 U10657 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n8068) );
  NAND2_X1 U10658 ( .A1(n8077), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8069) );
  INV_X1 U10659 ( .A(n14419), .ZN(n11452) );
  NAND2_X1 U10660 ( .A1(n11452), .A2(n11713), .ZN(n8070) );
  NAND2_X1 U10661 ( .A1(n12989), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n8076) );
  NAND2_X1 U10662 ( .A1(n8521), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n8075) );
  INV_X1 U10663 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n8072) );
  XNOR2_X1 U10664 ( .A(n8072), .B(P2_REG3_REG_3__SCAN_IN), .ZN(n12534) );
  NAND2_X1 U10665 ( .A1(n8553), .A2(n12534), .ZN(n8074) );
  INV_X1 U10666 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n11162) );
  OR2_X1 U10667 ( .A1(n8376), .A2(n11162), .ZN(n8073) );
  NAND4_X1 U10668 ( .A1(n8076), .A2(n8075), .A3(n8074), .A4(n8073), .ZN(n14418) );
  INV_X1 U10669 ( .A(n8078), .ZN(n8079) );
  NAND2_X1 U10670 ( .A1(n8080), .A2(n8079), .ZN(n8081) );
  NAND2_X1 U10671 ( .A1(n8081), .A2(n8086), .ZN(n8082) );
  XNOR2_X1 U10672 ( .A(n8094), .B(SI_4_), .ZN(n8091) );
  XNOR2_X1 U10673 ( .A(n8082), .B(n8091), .ZN(n10654) );
  NAND2_X1 U10674 ( .A1(n10654), .A2(n13125), .ZN(n8083) );
  XNOR2_X1 U10675 ( .A(n14418), .B(n7190), .ZN(n14338) );
  NAND2_X1 U10676 ( .A1(n8088), .A2(n8087), .ZN(n8093) );
  NOR2_X1 U10677 ( .A1(n8089), .A2(SI_3_), .ZN(n8090) );
  NAND2_X1 U10678 ( .A1(n8094), .A2(SI_4_), .ZN(n8095) );
  XNOR2_X1 U10679 ( .A(n8098), .B(SI_5_), .ZN(n8125) );
  INV_X1 U10680 ( .A(n8125), .ZN(n8097) );
  XNOR2_X1 U10681 ( .A(n8133), .B(n8131), .ZN(n10693) );
  NAND2_X1 U10682 ( .A1(n10693), .A2(n13125), .ZN(n8105) );
  INV_X1 U10683 ( .A(n8100), .ZN(n8102) );
  INV_X1 U10684 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n8101) );
  NAND2_X1 U10685 ( .A1(n8102), .A2(n8101), .ZN(n8137) );
  NAND2_X1 U10686 ( .A1(n8137), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8103) );
  XNOR2_X1 U10687 ( .A(n8103), .B(P2_IR_REG_6__SCAN_IN), .ZN(n11168) );
  AOI22_X1 U10688 ( .A1(n13126), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n8368), 
        .B2(n11168), .ZN(n8104) );
  NAND2_X2 U10689 ( .A1(n8105), .A2(n8104), .ZN(n14148) );
  NAND2_X1 U10690 ( .A1(n8554), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n8113) );
  NAND3_X1 U10691 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .A3(P2_REG3_REG_5__SCAN_IN), .ZN(n8117) );
  INV_X1 U10692 ( .A(n8117), .ZN(n8106) );
  INV_X1 U10693 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n10791) );
  NAND2_X1 U10694 ( .A1(n8117), .A2(n10791), .ZN(n8107) );
  AND2_X1 U10695 ( .A1(n8144), .A2(n8107), .ZN(n12611) );
  NAND2_X1 U10696 ( .A1(n8553), .A2(n12611), .ZN(n8111) );
  INV_X1 U10697 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n8109) );
  NAND2_X1 U10698 ( .A1(n7900), .A2(n14416), .ZN(n8597) );
  INV_X1 U10699 ( .A(n14416), .ZN(n11744) );
  NAND2_X1 U10700 ( .A1(n8554), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n8122) );
  NAND2_X1 U10701 ( .A1(n8521), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n8121) );
  INV_X1 U10702 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n8115) );
  NAND2_X1 U10703 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n8114) );
  NAND2_X1 U10704 ( .A1(n8115), .A2(n8114), .ZN(n8116) );
  AND2_X1 U10705 ( .A1(n8117), .A2(n8116), .ZN(n11738) );
  NAND2_X1 U10706 ( .A1(n8553), .A2(n11738), .ZN(n8120) );
  INV_X1 U10707 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n8118) );
  OR2_X1 U10708 ( .A1(n8557), .A2(n8118), .ZN(n8119) );
  NAND2_X1 U10709 ( .A1(n8100), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8123) );
  XNOR2_X1 U10710 ( .A(n8123), .B(P2_IR_REG_5__SCAN_IN), .ZN(n14451) );
  AOI22_X1 U10711 ( .A1(n13126), .A2(P1_DATAO_REG_5__SCAN_IN), .B1(n8368), 
        .B2(n14451), .ZN(n8127) );
  XNOR2_X1 U10712 ( .A(n8125), .B(n8124), .ZN(n10690) );
  NAND2_X1 U10713 ( .A1(n10690), .A2(n13125), .ZN(n8126) );
  NOR2_X1 U10714 ( .A1(n14417), .A2(n15983), .ZN(n8129) );
  NOR2_X1 U10715 ( .A1(n14148), .A2(n14416), .ZN(n8128) );
  INV_X1 U10716 ( .A(n14418), .ZN(n11743) );
  NAND2_X1 U10717 ( .A1(n11743), .A2(n7190), .ZN(n12220) );
  NAND2_X1 U10718 ( .A1(n14417), .A2(n15983), .ZN(n8130) );
  NAND2_X1 U10719 ( .A1(n14335), .A2(n8130), .ZN(n12231) );
  INV_X1 U10720 ( .A(n8131), .ZN(n8132) );
  NAND2_X1 U10721 ( .A1(n8133), .A2(n8132), .ZN(n8136) );
  NAND2_X1 U10722 ( .A1(n8134), .A2(SI_6_), .ZN(n8135) );
  XNOR2_X1 U10723 ( .A(n8154), .B(SI_7_), .ZN(n8151) );
  XNOR2_X1 U10724 ( .A(n8153), .B(n8151), .ZN(n10672) );
  NAND2_X1 U10725 ( .A1(n10672), .A2(n13125), .ZN(n8140) );
  NAND2_X1 U10726 ( .A1(n8157), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8138) );
  XNOR2_X1 U10727 ( .A(n8138), .B(P2_IR_REG_7__SCAN_IN), .ZN(n14470) );
  AOI22_X1 U10728 ( .A1(n13126), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n8368), 
        .B2(n14470), .ZN(n8139) );
  NAND2_X1 U10729 ( .A1(n8140), .A2(n8139), .ZN(n15995) );
  NAND2_X1 U10730 ( .A1(n12989), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n8149) );
  NAND2_X1 U10731 ( .A1(n12988), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n8148) );
  INV_X1 U10732 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n8143) );
  NAND2_X1 U10733 ( .A1(n8144), .A2(n8143), .ZN(n8145) );
  AND2_X1 U10734 ( .A1(n8165), .A2(n8145), .ZN(n12239) );
  NAND2_X1 U10735 ( .A1(n8553), .A2(n12239), .ZN(n8147) );
  INV_X1 U10736 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n12238) );
  OR2_X1 U10737 ( .A1(n8376), .A2(n12238), .ZN(n8146) );
  NAND4_X1 U10738 ( .A1(n8149), .A2(n8148), .A3(n8147), .A4(n8146), .ZN(n14415) );
  INV_X1 U10739 ( .A(n14415), .ZN(n8601) );
  OR2_X1 U10740 ( .A1(n15995), .A2(n14415), .ZN(n8150) );
  INV_X1 U10741 ( .A(n8151), .ZN(n8152) );
  NAND2_X1 U10742 ( .A1(n8153), .A2(n8152), .ZN(n8156) );
  NAND2_X1 U10743 ( .A1(n8154), .A2(SI_7_), .ZN(n8155) );
  MUX2_X1 U10744 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(P1_DATAO_REG_8__SCAN_IN), 
        .S(n10696), .Z(n8176) );
  XNOR2_X1 U10745 ( .A(n8176), .B(SI_8_), .ZN(n8173) );
  NAND2_X1 U10746 ( .A1(n10711), .A2(n13125), .ZN(n8162) );
  INV_X1 U10747 ( .A(n8157), .ZN(n8159) );
  NAND2_X1 U10748 ( .A1(n8159), .A2(n8158), .ZN(n8178) );
  NAND2_X1 U10749 ( .A1(n8178), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8160) );
  XNOR2_X1 U10750 ( .A(n8160), .B(P2_IR_REG_8__SCAN_IN), .ZN(n14484) );
  AOI22_X1 U10751 ( .A1(n13126), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n8368), 
        .B2(n14484), .ZN(n8161) );
  NAND2_X1 U10752 ( .A1(n8554), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n8171) );
  NAND2_X1 U10753 ( .A1(n8521), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n8170) );
  INV_X1 U10754 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n8164) );
  NAND2_X1 U10755 ( .A1(n8165), .A2(n8164), .ZN(n8166) );
  AND2_X1 U10756 ( .A1(n8185), .A2(n8166), .ZN(n12583) );
  NAND2_X1 U10757 ( .A1(n8553), .A2(n12583), .ZN(n8169) );
  INV_X1 U10758 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n8167) );
  OR2_X1 U10759 ( .A1(n8557), .A2(n8167), .ZN(n8168) );
  NAND4_X1 U10760 ( .A1(n8171), .A2(n8170), .A3(n8169), .A4(n8168), .ZN(n14414) );
  XNOR2_X1 U10761 ( .A(n14154), .B(n14414), .ZN(n14341) );
  NAND2_X1 U10762 ( .A1(n14154), .A2(n14414), .ZN(n8172) );
  INV_X1 U10763 ( .A(n8173), .ZN(n8174) );
  NAND2_X1 U10764 ( .A1(n8176), .A2(SI_8_), .ZN(n8177) );
  MUX2_X1 U10765 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(P1_DATAO_REG_9__SCAN_IN), 
        .S(n10696), .Z(n8195) );
  XNOR2_X1 U10766 ( .A(n8194), .B(n8192), .ZN(n10745) );
  NAND2_X1 U10767 ( .A1(n10745), .A2(n13125), .ZN(n8183) );
  OAI21_X1 U10768 ( .B1(n8178), .B2(P2_IR_REG_8__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n8179) );
  MUX2_X1 U10769 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8179), .S(
        P2_IR_REG_9__SCAN_IN), .Z(n8181) );
  INV_X1 U10770 ( .A(n8180), .ZN(n8291) );
  AOI22_X1 U10771 ( .A1(n7193), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n8368), .B2(
        n11221), .ZN(n8182) );
  NAND2_X1 U10772 ( .A1(n8643), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n8190) );
  NAND2_X1 U10773 ( .A1(n8521), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n8189) );
  NAND2_X1 U10774 ( .A1(n8185), .A2(n8184), .ZN(n8186) );
  AND2_X1 U10775 ( .A1(n8202), .A2(n8186), .ZN(n12433) );
  NAND2_X1 U10776 ( .A1(n8553), .A2(n12433), .ZN(n8188) );
  INV_X1 U10777 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n12396) );
  OR2_X1 U10778 ( .A1(n8557), .A2(n12396), .ZN(n8187) );
  NAND4_X1 U10779 ( .A1(n8190), .A2(n8189), .A3(n8188), .A4(n8187), .ZN(n14413) );
  INV_X1 U10780 ( .A(n14413), .ZN(n8607) );
  XNOR2_X1 U10781 ( .A(n14159), .B(n8607), .ZN(n12379) );
  NAND2_X1 U10782 ( .A1(n14159), .A2(n14413), .ZN(n8191) );
  NAND2_X1 U10783 ( .A1(n8195), .A2(SI_9_), .ZN(n8196) );
  MUX2_X1 U10784 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(P1_DATAO_REG_10__SCAN_IN), 
        .S(n10696), .Z(n8213) );
  NAND2_X1 U10785 ( .A1(n11036), .A2(n13125), .ZN(n8200) );
  NAND2_X1 U10786 ( .A1(n8291), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8197) );
  MUX2_X1 U10787 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8197), .S(
        P2_IR_REG_10__SCAN_IN), .Z(n8198) );
  AOI22_X1 U10788 ( .A1(n7193), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n8368), 
        .B2(n11238), .ZN(n8199) );
  NAND2_X1 U10789 ( .A1(n12989), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n8208) );
  NAND2_X1 U10790 ( .A1(n12988), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n8207) );
  NAND2_X1 U10791 ( .A1(n8202), .A2(n8201), .ZN(n8203) );
  AND2_X1 U10792 ( .A1(n8221), .A2(n8203), .ZN(n12815) );
  NAND2_X1 U10793 ( .A1(n8553), .A2(n12815), .ZN(n8206) );
  INV_X1 U10794 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n8204) );
  OR2_X1 U10795 ( .A1(n8376), .A2(n8204), .ZN(n8205) );
  NAND4_X1 U10796 ( .A1(n8208), .A2(n8207), .A3(n8206), .A4(n8205), .ZN(n14412) );
  NAND2_X1 U10797 ( .A1(n14842), .A2(n14412), .ZN(n8210) );
  OR2_X1 U10798 ( .A1(n14842), .A2(n14412), .ZN(n8209) );
  AND2_X2 U10799 ( .A1(n8210), .A2(n8209), .ZN(n14344) );
  MUX2_X1 U10800 ( .A(n11061), .B(n11058), .S(n10696), .Z(n8214) );
  INV_X1 U10801 ( .A(n8214), .ZN(n8215) );
  NAND2_X1 U10802 ( .A1(n8215), .A2(SI_11_), .ZN(n8216) );
  XNOR2_X1 U10803 ( .A(n8231), .B(n8230), .ZN(n11057) );
  NAND2_X1 U10804 ( .A1(n11057), .A2(n13125), .ZN(n8219) );
  NAND2_X1 U10805 ( .A1(n8235), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8217) );
  XNOR2_X1 U10806 ( .A(n8217), .B(P2_IR_REG_11__SCAN_IN), .ZN(n11522) );
  AOI22_X1 U10807 ( .A1(n13126), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n8368), 
        .B2(n11522), .ZN(n8218) );
  NAND2_X1 U10808 ( .A1(n8554), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n8226) );
  NAND2_X1 U10809 ( .A1(n12988), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n8225) );
  INV_X1 U10810 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n8220) );
  NAND2_X1 U10811 ( .A1(n8221), .A2(n8220), .ZN(n8222) );
  AND2_X1 U10812 ( .A1(n8245), .A2(n8222), .ZN(n12871) );
  NAND2_X1 U10813 ( .A1(n8553), .A2(n12871), .ZN(n8224) );
  INV_X1 U10814 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n14890) );
  OR2_X1 U10815 ( .A1(n8557), .A2(n14890), .ZN(n8223) );
  NAND4_X1 U10816 ( .A1(n8226), .A2(n8225), .A3(n8224), .A4(n8223), .ZN(n14411) );
  NAND2_X1 U10817 ( .A1(n14171), .A2(n14411), .ZN(n8227) );
  NAND2_X1 U10818 ( .A1(n8232), .A2(n10744), .ZN(n8253) );
  INV_X1 U10819 ( .A(n8232), .ZN(n8233) );
  NAND2_X1 U10820 ( .A1(n8233), .A2(SI_12_), .ZN(n8234) );
  XNOR2_X1 U10821 ( .A(n8252), .B(n7983), .ZN(n11207) );
  NAND2_X1 U10822 ( .A1(n11207), .A2(n13125), .ZN(n8242) );
  INV_X1 U10823 ( .A(n8235), .ZN(n8237) );
  NAND2_X1 U10824 ( .A1(n8237), .A2(n8236), .ZN(n8239) );
  NAND2_X1 U10825 ( .A1(n8239), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8238) );
  MUX2_X1 U10826 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8238), .S(
        P2_IR_REG_12__SCAN_IN), .Z(n8240) );
  AOI22_X1 U10827 ( .A1(n7193), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n8368), 
        .B2(n11523), .ZN(n8241) );
  NAND2_X1 U10828 ( .A1(n12988), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n8250) );
  INV_X1 U10829 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n8244) );
  NAND2_X1 U10830 ( .A1(n8245), .A2(n8244), .ZN(n8246) );
  AND2_X1 U10831 ( .A1(n8260), .A2(n8246), .ZN(n12896) );
  NAND2_X1 U10832 ( .A1(n8553), .A2(n12896), .ZN(n8249) );
  NAND2_X1 U10833 ( .A1(n12989), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n8248) );
  INV_X1 U10834 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n11725) );
  OR2_X1 U10835 ( .A1(n8376), .A2(n11725), .ZN(n8247) );
  NAND4_X1 U10836 ( .A1(n8250), .A2(n8249), .A3(n8248), .A4(n8247), .ZN(n14410) );
  AND2_X1 U10837 ( .A1(n14829), .A2(n14410), .ZN(n8251) );
  MUX2_X1 U10838 ( .A(n11383), .B(n11381), .S(n10696), .Z(n8254) );
  INV_X1 U10839 ( .A(n8254), .ZN(n8255) );
  NAND2_X1 U10840 ( .A1(n8255), .A2(SI_13_), .ZN(n8256) );
  XNOR2_X1 U10841 ( .A(n8268), .B(n7978), .ZN(n11379) );
  NAND2_X1 U10842 ( .A1(n11379), .A2(n13125), .ZN(n8259) );
  NAND2_X1 U10843 ( .A1(n8270), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8257) );
  XNOR2_X1 U10844 ( .A(n8257), .B(P2_IR_REG_13__SCAN_IN), .ZN(n11927) );
  AOI22_X1 U10845 ( .A1(n13126), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n8368), 
        .B2(n11927), .ZN(n8258) );
  NAND2_X1 U10846 ( .A1(n8643), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n8266) );
  NAND2_X1 U10847 ( .A1(n12988), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n8265) );
  NAND2_X1 U10848 ( .A1(n8260), .A2(n12925), .ZN(n8261) );
  AND2_X1 U10849 ( .A1(n8275), .A2(n8261), .ZN(n12929) );
  NAND2_X1 U10850 ( .A1(n8553), .A2(n12929), .ZN(n8264) );
  INV_X1 U10851 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n8262) );
  OR2_X1 U10852 ( .A1(n8557), .A2(n8262), .ZN(n8263) );
  NAND4_X1 U10853 ( .A1(n8266), .A2(n8265), .A3(n8264), .A4(n8263), .ZN(n14409) );
  NAND2_X1 U10854 ( .A1(n14191), .A2(n14409), .ZN(n8267) );
  MUX2_X1 U10855 ( .A(n11590), .B(n11592), .S(n9991), .Z(n8307) );
  NAND2_X1 U10856 ( .A1(n11588), .A2(n13125), .ZN(n8273) );
  OAI21_X1 U10857 ( .B1(n8270), .B2(P2_IR_REG_13__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n8271) );
  XNOR2_X1 U10858 ( .A(n8271), .B(P2_IR_REG_14__SCAN_IN), .ZN(n11993) );
  AOI22_X1 U10859 ( .A1(n7193), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n8368), 
        .B2(n11993), .ZN(n8272) );
  NAND2_X1 U10860 ( .A1(n12988), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n8281) );
  INV_X1 U10861 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n8274) );
  NAND2_X1 U10862 ( .A1(n8275), .A2(n8274), .ZN(n8276) );
  AND2_X1 U10863 ( .A1(n8300), .A2(n8276), .ZN(n13985) );
  NAND2_X1 U10864 ( .A1(n13985), .A2(n8553), .ZN(n8280) );
  NAND2_X1 U10865 ( .A1(n8643), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n8279) );
  INV_X1 U10866 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n8277) );
  OR2_X1 U10867 ( .A1(n8557), .A2(n8277), .ZN(n8278) );
  NAND4_X1 U10868 ( .A1(n8281), .A2(n8280), .A3(n8279), .A4(n8278), .ZN(n14408) );
  INV_X1 U10869 ( .A(n14408), .ZN(n14188) );
  NAND2_X1 U10870 ( .A1(n12916), .A2(n14328), .ZN(n8283) );
  NAND2_X1 U10871 ( .A1(n14824), .A2(n14408), .ZN(n8282) );
  INV_X1 U10872 ( .A(n8307), .ZN(n8311) );
  OR2_X1 U10873 ( .A1(n8310), .A2(n11128), .ZN(n8284) );
  NAND2_X1 U10874 ( .A1(n8285), .A2(n8284), .ZN(n8289) );
  MUX2_X1 U10875 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(P1_DATAO_REG_15__SCAN_IN), 
        .S(n10696), .Z(n8286) );
  INV_X1 U10876 ( .A(n8286), .ZN(n8287) );
  INV_X1 U10877 ( .A(SI_15_), .ZN(n11125) );
  NAND2_X1 U10878 ( .A1(n8287), .A2(n11125), .ZN(n8312) );
  NAND2_X1 U10879 ( .A1(n8314), .A2(n8312), .ZN(n8288) );
  NAND2_X1 U10880 ( .A1(n11666), .A2(n13125), .ZN(n8298) );
  OR2_X1 U10881 ( .A1(n8291), .A2(n8290), .ZN(n8293) );
  NAND2_X1 U10882 ( .A1(n8293), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8292) );
  MUX2_X1 U10883 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8292), .S(
        P2_IR_REG_15__SCAN_IN), .Z(n8296) );
  INV_X1 U10884 ( .A(n8293), .ZN(n8295) );
  NAND2_X1 U10885 ( .A1(n8295), .A2(n8294), .ZN(n8320) );
  NAND2_X1 U10886 ( .A1(n8296), .A2(n8320), .ZN(n11996) );
  INV_X1 U10887 ( .A(n11996), .ZN(n12679) );
  AOI22_X1 U10888 ( .A1(n13126), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n8368), 
        .B2(n12679), .ZN(n8297) );
  INV_X1 U10889 ( .A(n8324), .ZN(n8325) );
  INV_X1 U10890 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n11990) );
  NAND2_X1 U10891 ( .A1(n8300), .A2(n11990), .ZN(n8301) );
  NAND2_X1 U10892 ( .A1(n8325), .A2(n8301), .ZN(n14735) );
  NAND2_X1 U10893 ( .A1(n12988), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n8303) );
  NAND2_X1 U10894 ( .A1(n12989), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n8302) );
  AND2_X1 U10895 ( .A1(n8303), .A2(n8302), .ZN(n8305) );
  NAND2_X1 U10896 ( .A1(n8554), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n8304) );
  OAI211_X1 U10897 ( .C1(n14735), .C2(n8648), .A(n8305), .B(n8304), .ZN(n14407) );
  XNOR2_X1 U10898 ( .A(n14817), .B(n14407), .ZN(n14353) );
  OAI21_X1 U10899 ( .B1(n11128), .B2(n8307), .A(n8314), .ZN(n8308) );
  INV_X1 U10900 ( .A(n8308), .ZN(n8309) );
  NOR2_X1 U10901 ( .A1(n8311), .A2(SI_14_), .ZN(n8315) );
  INV_X1 U10902 ( .A(n8312), .ZN(n8313) );
  MUX2_X1 U10903 ( .A(n9170), .B(n11587), .S(n9991), .Z(n8317) );
  INV_X1 U10904 ( .A(n8317), .ZN(n8318) );
  NAND2_X1 U10905 ( .A1(n8318), .A2(SI_16_), .ZN(n8319) );
  XNOR2_X1 U10906 ( .A(n8329), .B(n7988), .ZN(n11548) );
  NAND2_X1 U10907 ( .A1(n11548), .A2(n13125), .ZN(n8323) );
  NAND2_X1 U10908 ( .A1(n8320), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8321) );
  XNOR2_X1 U10909 ( .A(n8321), .B(P2_IR_REG_16__SCAN_IN), .ZN(n15935) );
  AOI22_X1 U10910 ( .A1(n7193), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n8368), 
        .B2(n15935), .ZN(n8322) );
  NAND2_X2 U10911 ( .A1(n8323), .A2(n8322), .ZN(n14809) );
  INV_X1 U10912 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n14884) );
  INV_X1 U10913 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n15927) );
  NAND2_X1 U10914 ( .A1(n8325), .A2(n15927), .ZN(n8326) );
  NAND2_X1 U10915 ( .A1(n8336), .A2(n8326), .ZN(n14707) );
  OR2_X1 U10916 ( .A1(n14707), .A2(n8648), .ZN(n8328) );
  AOI22_X1 U10917 ( .A1(n8643), .A2(P2_REG2_REG_16__SCAN_IN), .B1(n12988), 
        .B2(P2_REG1_REG_16__SCAN_IN), .ZN(n8327) );
  OAI211_X1 U10918 ( .C1(n8557), .C2(n14884), .A(n8328), .B(n8327), .ZN(n14406) );
  AND2_X1 U10919 ( .A1(n14809), .A2(n14406), .ZN(n14693) );
  OR2_X1 U10920 ( .A1(n14817), .A2(n14407), .ZN(n14691) );
  OAI22_X1 U10921 ( .A1(n14691), .A2(n14693), .B1(n14809), .B2(n14406), .ZN(
        n8340) );
  MUX2_X1 U10922 ( .A(n9183), .B(n11664), .S(n10696), .Z(n8345) );
  XNOR2_X1 U10923 ( .A(n8345), .B(SI_17_), .ZN(n8331) );
  XNOR2_X1 U10924 ( .A(n8344), .B(n8331), .ZN(n11593) );
  NAND2_X1 U10925 ( .A1(n11593), .A2(n13125), .ZN(n8334) );
  XNOR2_X1 U10926 ( .A(n8332), .B(P2_IR_REG_17__SCAN_IN), .ZN(n12803) );
  AOI22_X1 U10927 ( .A1(n7193), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n8368), 
        .B2(n12803), .ZN(n8333) );
  INV_X1 U10928 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n8335) );
  NAND2_X1 U10929 ( .A1(n8336), .A2(n8335), .ZN(n8337) );
  NAND2_X1 U10930 ( .A1(n8355), .A2(n8337), .ZN(n14699) );
  AOI22_X1 U10931 ( .A1(n8643), .A2(P2_REG2_REG_17__SCAN_IN), .B1(n12988), 
        .B2(P2_REG1_REG_17__SCAN_IN), .ZN(n8339) );
  NAND2_X1 U10932 ( .A1(n12989), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n8338) );
  OAI211_X1 U10933 ( .C1(n14699), .C2(n8648), .A(n8339), .B(n8338), .ZN(n14405) );
  XNOR2_X1 U10934 ( .A(n14697), .B(n14405), .ZN(n14695) );
  NOR2_X1 U10935 ( .A1(n8340), .A2(n14695), .ZN(n8341) );
  INV_X1 U10936 ( .A(n8345), .ZN(n8342) );
  NAND2_X1 U10937 ( .A1(n8342), .A2(SI_17_), .ZN(n8343) );
  INV_X1 U10938 ( .A(SI_17_), .ZN(n11348) );
  NAND2_X1 U10939 ( .A1(n8345), .A2(n11348), .ZN(n8346) );
  INV_X1 U10940 ( .A(SI_18_), .ZN(n11459) );
  NAND2_X1 U10941 ( .A1(n8432), .A2(n11459), .ZN(n8347) );
  MUX2_X1 U10942 ( .A(n11971), .B(n11972), .S(n10696), .Z(n8383) );
  NAND2_X1 U10943 ( .A1(n8348), .A2(n8383), .ZN(n8349) );
  NAND2_X1 U10944 ( .A1(n8571), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8350) );
  MUX2_X1 U10945 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8350), .S(
        P2_IR_REG_18__SCAN_IN), .Z(n8351) );
  AND2_X1 U10946 ( .A1(n8351), .A2(n8577), .ZN(n12806) );
  AOI22_X1 U10947 ( .A1(n7193), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n8368), 
        .B2(n12806), .ZN(n8352) );
  INV_X1 U10948 ( .A(n8355), .ZN(n8353) );
  INV_X1 U10949 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n8354) );
  NAND2_X1 U10950 ( .A1(n8355), .A2(n8354), .ZN(n8356) );
  NAND2_X1 U10951 ( .A1(n8372), .A2(n8356), .ZN(n14678) );
  OR2_X1 U10952 ( .A1(n14678), .A2(n8648), .ZN(n8362) );
  INV_X1 U10953 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n8359) );
  NAND2_X1 U10954 ( .A1(n8643), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n8358) );
  NAND2_X1 U10955 ( .A1(n12988), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n8357) );
  OAI211_X1 U10956 ( .C1(n8359), .C2(n8557), .A(n8358), .B(n8357), .ZN(n8360)
         );
  INV_X1 U10957 ( .A(n8360), .ZN(n8361) );
  NAND2_X1 U10958 ( .A1(n8362), .A2(n8361), .ZN(n14404) );
  XNOR2_X1 U10959 ( .A(n14800), .B(n14404), .ZN(n14671) );
  OR2_X1 U10960 ( .A1(n14800), .A2(n14404), .ZN(n8363) );
  MUX2_X1 U10961 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(P1_DATAO_REG_19__SCAN_IN), 
        .S(n10696), .Z(n8386) );
  XNOR2_X1 U10962 ( .A(n8386), .B(SI_19_), .ZN(n8385) );
  NAND2_X1 U10963 ( .A1(n12141), .A2(n13125), .ZN(n8370) );
  NAND2_X1 U10964 ( .A1(n8577), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8367) );
  AOI22_X1 U10965 ( .A1(n7193), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n14322), 
        .B2(n8368), .ZN(n8369) );
  INV_X1 U10966 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n8371) );
  NAND2_X1 U10967 ( .A1(n8372), .A2(n8371), .ZN(n8373) );
  AND2_X1 U10968 ( .A1(n8394), .A2(n8373), .ZN(n14661) );
  NAND2_X1 U10969 ( .A1(n14661), .A2(n8553), .ZN(n8379) );
  INV_X1 U10970 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n14499) );
  NAND2_X1 U10971 ( .A1(n12988), .A2(P2_REG1_REG_19__SCAN_IN), .ZN(n8375) );
  NAND2_X1 U10972 ( .A1(n12989), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n8374) );
  OAI211_X1 U10973 ( .C1(n8376), .C2(n14499), .A(n8375), .B(n8374), .ZN(n8377)
         );
  INV_X1 U10974 ( .A(n8377), .ZN(n8378) );
  NAND2_X1 U10975 ( .A1(n8379), .A2(n8378), .ZN(n14403) );
  NAND2_X1 U10976 ( .A1(n7907), .A2(n14403), .ZN(n8380) );
  OR2_X1 U10977 ( .A1(n7907), .A2(n14403), .ZN(n8381) );
  INV_X1 U10978 ( .A(n8383), .ZN(n8382) );
  NOR2_X1 U10979 ( .A1(n8383), .A2(n11459), .ZN(n8384) );
  INV_X1 U10980 ( .A(n8386), .ZN(n8387) );
  INV_X1 U10981 ( .A(SI_20_), .ZN(n11751) );
  NAND2_X1 U10982 ( .A1(n8388), .A2(n11751), .ZN(n8389) );
  MUX2_X1 U10983 ( .A(n12096), .B(n12184), .S(n10696), .Z(n8413) );
  NAND2_X1 U10984 ( .A1(n8390), .A2(n8413), .ZN(n8391) );
  NAND2_X1 U10985 ( .A1(n13126), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n8392) );
  INV_X1 U10986 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n8393) );
  NAND2_X1 U10987 ( .A1(n8394), .A2(n8393), .ZN(n8395) );
  NAND2_X1 U10988 ( .A1(n8423), .A2(n8395), .ZN(n14641) );
  OR2_X1 U10989 ( .A1(n14641), .A2(n8648), .ZN(n8400) );
  INV_X1 U10990 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n10811) );
  NAND2_X1 U10991 ( .A1(n8643), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n8397) );
  NAND2_X1 U10992 ( .A1(n12989), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n8396) );
  OAI211_X1 U10993 ( .C1(n8141), .C2(n10811), .A(n8397), .B(n8396), .ZN(n8398)
         );
  INV_X1 U10994 ( .A(n8398), .ZN(n8399) );
  NAND2_X1 U10995 ( .A1(n8400), .A2(n8399), .ZN(n14402) );
  NAND2_X1 U10996 ( .A1(n14790), .A2(n14402), .ZN(n8402) );
  MUX2_X1 U10997 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(P1_DATAO_REG_21__SCAN_IN), 
        .S(n10696), .Z(n8403) );
  AND2_X1 U10998 ( .A1(n8404), .A2(n8416), .ZN(n8405) );
  INV_X1 U10999 ( .A(n8407), .ZN(n8408) );
  INV_X1 U11000 ( .A(n8409), .ZN(n8412) );
  NOR2_X1 U11001 ( .A1(n8413), .A2(n11751), .ZN(n8410) );
  OAI21_X1 U11002 ( .B1(n8432), .B2(n8430), .A(n8433), .ZN(n8417) );
  INV_X1 U11003 ( .A(n8413), .ZN(n8414) );
  NAND2_X1 U11004 ( .A1(n8417), .A2(n8436), .ZN(n8418) );
  NAND2_X1 U11005 ( .A1(n7193), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n8421) );
  INV_X1 U11006 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n14013) );
  NAND2_X1 U11007 ( .A1(n8423), .A2(n14013), .ZN(n8424) );
  NAND2_X1 U11008 ( .A1(n8458), .A2(n8424), .ZN(n14012) );
  OR2_X1 U11009 ( .A1(n14012), .A2(n8648), .ZN(n8429) );
  INV_X1 U11010 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n14787) );
  NAND2_X1 U11011 ( .A1(n12989), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n8426) );
  NAND2_X1 U11012 ( .A1(n8554), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n8425) );
  OAI211_X1 U11013 ( .C1(n8141), .C2(n14787), .A(n8426), .B(n8425), .ZN(n8427)
         );
  INV_X1 U11014 ( .A(n8427), .ZN(n8428) );
  NAND2_X1 U11015 ( .A1(n8429), .A2(n8428), .ZN(n14401) );
  XNOR2_X1 U11016 ( .A(n14628), .B(n14401), .ZN(n14626) );
  INV_X1 U11017 ( .A(n8436), .ZN(n8431) );
  INV_X1 U11018 ( .A(n8433), .ZN(n8437) );
  INV_X1 U11019 ( .A(n8434), .ZN(n8435) );
  NAND2_X1 U11020 ( .A1(n8474), .A2(SI_22_), .ZN(n8440) );
  OR2_X1 U11021 ( .A1(n8474), .A2(SI_22_), .ZN(n8439) );
  NAND2_X1 U11022 ( .A1(n8440), .A2(n8439), .ZN(n9826) );
  MUX2_X1 U11023 ( .A(n9243), .B(n12356), .S(n9991), .Z(n8471) );
  NAND2_X1 U11024 ( .A1(n8455), .A2(n8440), .ZN(n8442) );
  MUX2_X1 U11025 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(P1_DATAO_REG_23__SCAN_IN), 
        .S(n10696), .Z(n8475) );
  XNOR2_X1 U11026 ( .A(n8475), .B(SI_23_), .ZN(n8441) );
  NAND2_X1 U11027 ( .A1(n12317), .A2(n13125), .ZN(n8444) );
  NAND2_X1 U11028 ( .A1(n7193), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n8443) );
  INV_X1 U11029 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n14069) );
  NOR2_X2 U11030 ( .A1(n8458), .A2(n14069), .ZN(n8445) );
  INV_X1 U11031 ( .A(n8445), .ZN(n8460) );
  INV_X1 U11032 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n8446) );
  NAND2_X1 U11033 ( .A1(n8460), .A2(n8446), .ZN(n8447) );
  NAND2_X1 U11034 ( .A1(n8484), .A2(n8447), .ZN(n14598) );
  OR2_X1 U11035 ( .A1(n14598), .A2(n8648), .ZN(n8453) );
  INV_X1 U11036 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n8450) );
  NAND2_X1 U11037 ( .A1(n12988), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n8449) );
  NAND2_X1 U11038 ( .A1(n8643), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n8448) );
  OAI211_X1 U11039 ( .C1(n8557), .C2(n8450), .A(n8449), .B(n8448), .ZN(n8451)
         );
  INV_X1 U11040 ( .A(n8451), .ZN(n8452) );
  OR2_X1 U11041 ( .A1(n14600), .A2(n14399), .ZN(n14358) );
  NAND2_X1 U11042 ( .A1(n9826), .A2(n8471), .ZN(n8454) );
  NAND2_X1 U11043 ( .A1(n12354), .A2(n13125), .ZN(n8457) );
  NAND2_X1 U11044 ( .A1(n7193), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n8456) );
  NAND2_X1 U11045 ( .A1(n8458), .A2(n14069), .ZN(n8459) );
  NAND2_X1 U11046 ( .A1(n8460), .A2(n8459), .ZN(n14616) );
  INV_X1 U11047 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n8463) );
  NAND2_X1 U11048 ( .A1(n12988), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n8462) );
  NAND2_X1 U11049 ( .A1(n8643), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n8461) );
  OAI211_X1 U11050 ( .C1(n8463), .C2(n8557), .A(n8462), .B(n8461), .ZN(n8464)
         );
  INV_X1 U11051 ( .A(n8464), .ZN(n8465) );
  INV_X1 U11052 ( .A(n14400), .ZN(n14248) );
  NAND2_X1 U11053 ( .A1(n14618), .A2(n14248), .ZN(n8466) );
  NAND2_X1 U11054 ( .A1(n8634), .A2(n8466), .ZN(n14604) );
  OR2_X1 U11055 ( .A1(n14628), .A2(n14401), .ZN(n14588) );
  AND3_X1 U11056 ( .A1(n14358), .A2(n14604), .A3(n14588), .ZN(n8467) );
  AND2_X1 U11057 ( .A1(n14618), .A2(n14400), .ZN(n14590) );
  NAND2_X1 U11058 ( .A1(n14358), .A2(n14590), .ZN(n8468) );
  NAND2_X1 U11059 ( .A1(n14600), .A2(n14399), .ZN(n14357) );
  AND2_X1 U11060 ( .A1(n8468), .A2(n14357), .ZN(n8469) );
  INV_X1 U11061 ( .A(SI_22_), .ZN(n9245) );
  NAND2_X1 U11062 ( .A1(n8471), .A2(n9245), .ZN(n8473) );
  INV_X1 U11063 ( .A(n8475), .ZN(n8470) );
  INV_X1 U11064 ( .A(SI_23_), .ZN(n11940) );
  OAI22_X1 U11065 ( .A1(n8471), .A2(n9245), .B1(n8470), .B2(n11940), .ZN(n8472) );
  INV_X1 U11066 ( .A(SI_24_), .ZN(n12984) );
  NAND2_X1 U11067 ( .A1(n8476), .A2(n12984), .ZN(n8477) );
  INV_X1 U11068 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n12578) );
  INV_X1 U11069 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n12580) );
  MUX2_X1 U11070 ( .A(n12578), .B(n12580), .S(n10696), .Z(n8478) );
  NAND2_X1 U11071 ( .A1(n8479), .A2(n8478), .ZN(n8480) );
  NAND2_X1 U11072 ( .A1(n12577), .A2(n13125), .ZN(n8482) );
  NAND2_X1 U11073 ( .A1(n7193), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n8481) );
  INV_X1 U11074 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n14051) );
  NAND2_X1 U11075 ( .A1(n8484), .A2(n14051), .ZN(n8485) );
  NAND2_X1 U11076 ( .A1(n8497), .A2(n8485), .ZN(n14574) );
  INV_X1 U11077 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n8488) );
  NAND2_X1 U11078 ( .A1(n8554), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n8487) );
  NAND2_X1 U11079 ( .A1(n12988), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n8486) );
  OAI211_X1 U11080 ( .C1(n8488), .C2(n8557), .A(n8487), .B(n8486), .ZN(n8489)
         );
  INV_X1 U11081 ( .A(n8489), .ZN(n8490) );
  XNOR2_X1 U11082 ( .A(n14769), .B(n14261), .ZN(n14577) );
  NAND2_X1 U11083 ( .A1(n14769), .A2(n14398), .ZN(n8492) );
  MUX2_X1 U11084 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(P1_DATAO_REG_25__SCAN_IN), 
        .S(n10696), .Z(n8507) );
  NAND2_X1 U11085 ( .A1(n12789), .A2(n13125), .ZN(n8496) );
  NAND2_X1 U11086 ( .A1(n13126), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n8495) );
  INV_X1 U11087 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n14020) );
  NAND2_X1 U11088 ( .A1(n8497), .A2(n14020), .ZN(n8498) );
  NAND2_X1 U11089 ( .A1(n14563), .A2(n8553), .ZN(n8503) );
  INV_X1 U11090 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n14858) );
  NAND2_X1 U11091 ( .A1(n8643), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n8500) );
  NAND2_X1 U11092 ( .A1(n12988), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n8499) );
  OAI211_X1 U11093 ( .C1(n14858), .C2(n8557), .A(n8500), .B(n8499), .ZN(n8501)
         );
  INV_X1 U11094 ( .A(n8501), .ZN(n8502) );
  NAND2_X1 U11095 ( .A1(n14562), .A2(n14397), .ZN(n8505) );
  INV_X1 U11096 ( .A(SI_26_), .ZN(n12507) );
  NAND2_X1 U11097 ( .A1(n8510), .A2(n12507), .ZN(n8511) );
  MUX2_X1 U11098 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(P1_DATAO_REG_26__SCAN_IN), 
        .S(n10696), .Z(n8513) );
  NAND2_X1 U11099 ( .A1(n6793), .A2(n7891), .ZN(n8514) );
  NAND2_X1 U11100 ( .A1(n13126), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n8515) );
  INV_X1 U11101 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n8518) );
  NAND2_X1 U11102 ( .A1(n8519), .A2(n8518), .ZN(n8520) );
  NAND2_X1 U11103 ( .A1(n8551), .A2(n8520), .ZN(n14087) );
  INV_X1 U11104 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n10995) );
  NAND2_X1 U11105 ( .A1(n8643), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n8523) );
  NAND2_X1 U11106 ( .A1(n12989), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n8522) );
  OAI211_X1 U11107 ( .C1(n8141), .C2(n10995), .A(n8523), .B(n8522), .ZN(n8524)
         );
  INV_X1 U11108 ( .A(n8524), .ZN(n8525) );
  AND2_X1 U11109 ( .A1(n14549), .A2(n14396), .ZN(n8528) );
  OR2_X1 U11110 ( .A1(n14549), .A2(n14396), .ZN(n8527) );
  MUX2_X1 U11111 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(P1_DATAO_REG_27__SCAN_IN), 
        .S(n10696), .Z(n8541) );
  XNOR2_X1 U11112 ( .A(n8541), .B(SI_27_), .ZN(n8531) );
  NAND2_X1 U11113 ( .A1(n14911), .A2(n13125), .ZN(n8533) );
  NAND2_X1 U11114 ( .A1(n7193), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n8532) );
  XNOR2_X1 U11115 ( .A(n8551), .B(P2_REG3_REG_27__SCAN_IN), .ZN(n14532) );
  NAND2_X1 U11116 ( .A1(n14532), .A2(n8553), .ZN(n8538) );
  INV_X1 U11117 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n14855) );
  NAND2_X1 U11118 ( .A1(n8643), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n8535) );
  NAND2_X1 U11119 ( .A1(n12988), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n8534) );
  OAI211_X1 U11120 ( .C1(n14855), .C2(n8557), .A(n8535), .B(n8534), .ZN(n8536)
         );
  INV_X1 U11121 ( .A(n8536), .ZN(n8537) );
  NAND2_X1 U11122 ( .A1(n14749), .A2(n14395), .ZN(n8540) );
  NAND2_X1 U11123 ( .A1(n8541), .A2(SI_27_), .ZN(n8542) );
  INV_X1 U11124 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n13106) );
  INV_X1 U11125 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n14910) );
  MUX2_X1 U11126 ( .A(n13106), .B(n14910), .S(n9991), .Z(n8543) );
  INV_X1 U11127 ( .A(SI_28_), .ZN(n13971) );
  NAND2_X1 U11128 ( .A1(n8543), .A2(n13971), .ZN(n9932) );
  INV_X1 U11129 ( .A(n8543), .ZN(n8544) );
  NAND2_X1 U11130 ( .A1(n8544), .A2(SI_28_), .ZN(n8545) );
  NAND2_X1 U11131 ( .A1(n9932), .A2(n8545), .ZN(n9933) );
  XNOR2_X2 U11132 ( .A(n9934), .B(n9933), .ZN(n14907) );
  NAND2_X1 U11133 ( .A1(n14907), .A2(n13125), .ZN(n8547) );
  NAND2_X1 U11134 ( .A1(n7193), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n8546) );
  NAND2_X2 U11135 ( .A1(n8547), .A2(n8546), .ZN(n14519) );
  INV_X1 U11136 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n8549) );
  INV_X1 U11137 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n8548) );
  OAI21_X1 U11138 ( .B1(n8551), .B2(n8549), .A(n8548), .ZN(n8552) );
  NAND2_X1 U11139 ( .A1(P2_REG3_REG_27__SCAN_IN), .A2(P2_REG3_REG_28__SCAN_IN), 
        .ZN(n8550) );
  NAND2_X1 U11140 ( .A1(n14517), .A2(n8553), .ZN(n8560) );
  INV_X1 U11141 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n14852) );
  NAND2_X1 U11142 ( .A1(n8643), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n8556) );
  NAND2_X1 U11143 ( .A1(n12988), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n8555) );
  OAI211_X1 U11144 ( .C1(n14852), .C2(n8557), .A(n8556), .B(n8555), .ZN(n8558)
         );
  INV_X1 U11145 ( .A(n8558), .ZN(n8559) );
  NAND2_X1 U11146 ( .A1(n14519), .A2(n14394), .ZN(n10391) );
  OR2_X1 U11147 ( .A1(n14519), .A2(n14394), .ZN(n8561) );
  NOR2_X1 U11148 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_17__SCAN_IN), 
        .ZN(n8564) );
  NOR2_X1 U11149 ( .A1(P2_IR_REG_20__SCAN_IN), .A2(P2_IR_REG_21__SCAN_IN), 
        .ZN(n8574) );
  AND3_X1 U11150 ( .A1(n8574), .A2(n8564), .A3(n8568), .ZN(n8565) );
  AND3_X1 U11151 ( .A1(n8578), .A2(n8568), .A3(P2_IR_REG_20__SCAN_IN), .ZN(
        n8573) );
  XNOR2_X1 U11152 ( .A(n8567), .B(P2_IR_REG_31__SCAN_IN), .ZN(n8572) );
  NAND3_X1 U11153 ( .A1(n8578), .A2(n8568), .A3(n8567), .ZN(n8569) );
  AND2_X1 U11154 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_20__SCAN_IN), 
        .ZN(n8570) );
  XNOR2_X1 U11155 ( .A(n8575), .B(P2_IR_REG_31__SCAN_IN), .ZN(n8582) );
  AND2_X1 U11156 ( .A1(P2_IR_REG_22__SCAN_IN), .A2(P2_IR_REG_31__SCAN_IN), 
        .ZN(n8579) );
  AND2_X2 U11157 ( .A1(n14322), .A2(n14329), .ZN(n14383) );
  INV_X1 U11158 ( .A(n15995), .ZN(n12241) );
  INV_X1 U11159 ( .A(n14842), .ZN(n12468) );
  NAND2_X1 U11160 ( .A1(n12465), .A2(n14893), .ZN(n12836) );
  INV_X1 U11161 ( .A(n14817), .ZN(n14176) );
  INV_X1 U11162 ( .A(n14800), .ZN(n14681) );
  AND2_X2 U11163 ( .A1(n14561), .A2(n14759), .ZN(n14546) );
  AOI21_X1 U11164 ( .B1(n14530), .B2(n14519), .A(n14717), .ZN(n8586) );
  NAND2_X1 U11165 ( .A1(n8586), .A2(n6611), .ZN(n14521) );
  NAND2_X1 U11166 ( .A1(n11453), .A2(n14114), .ZN(n8587) );
  NAND2_X1 U11167 ( .A1(n11629), .A2(n14332), .ZN(n8590) );
  NAND2_X1 U11168 ( .A1(n11570), .A2(n14120), .ZN(n8589) );
  INV_X1 U11169 ( .A(n11671), .ZN(n14333) );
  NAND2_X1 U11170 ( .A1(n11673), .A2(n14333), .ZN(n8592) );
  NAND2_X1 U11171 ( .A1(n11452), .A2(n14129), .ZN(n8591) );
  NAND2_X1 U11172 ( .A1(n8592), .A2(n8591), .ZN(n11817) );
  INV_X1 U11173 ( .A(n14338), .ZN(n8593) );
  NAND2_X1 U11174 ( .A1(n11817), .A2(n8593), .ZN(n8595) );
  NAND2_X1 U11175 ( .A1(n11743), .A2(n14136), .ZN(n8594) );
  NAND2_X1 U11176 ( .A1(n14417), .A2(n8585), .ZN(n12613) );
  AND2_X1 U11177 ( .A1(n8599), .A2(n8598), .ZN(n8600) );
  AND2_X1 U11178 ( .A1(n15995), .A2(n8601), .ZN(n8602) );
  INV_X1 U11179 ( .A(n14414), .ZN(n8604) );
  NAND2_X1 U11180 ( .A1(n14154), .A2(n8604), .ZN(n8603) );
  OR2_X1 U11181 ( .A1(n14154), .A2(n8604), .ZN(n8605) );
  NAND2_X1 U11182 ( .A1(n8606), .A2(n8605), .ZN(n12380) );
  INV_X1 U11183 ( .A(n12379), .ZN(n14346) );
  NAND2_X1 U11184 ( .A1(n12380), .A2(n14346), .ZN(n8609) );
  OR2_X1 U11185 ( .A1(n14159), .A2(n8607), .ZN(n8608) );
  INV_X1 U11186 ( .A(n14344), .ZN(n8610) );
  INV_X1 U11187 ( .A(n14829), .ZN(n14173) );
  INV_X1 U11188 ( .A(n14411), .ZN(n8613) );
  INV_X1 U11189 ( .A(n14412), .ZN(n12661) );
  OR2_X1 U11190 ( .A1(n14842), .A2(n12661), .ZN(n12658) );
  OAI21_X1 U11191 ( .B1(n14171), .B2(n8613), .A(n12658), .ZN(n8611) );
  AOI21_X1 U11192 ( .B1(n14173), .B2(n14410), .A(n8611), .ZN(n8612) );
  NAND2_X1 U11193 ( .A1(n14171), .A2(n8613), .ZN(n12826) );
  NAND2_X1 U11194 ( .A1(n12826), .A2(n14410), .ZN(n8615) );
  NOR2_X1 U11195 ( .A1(n14410), .A2(n14411), .ZN(n8614) );
  AOI22_X1 U11196 ( .A1(n14829), .A2(n8615), .B1(n8614), .B2(n14171), .ZN(
        n8616) );
  INV_X1 U11197 ( .A(n14409), .ZN(n14190) );
  XNOR2_X1 U11198 ( .A(n14191), .B(n14190), .ZN(n14350) );
  OR2_X1 U11199 ( .A1(n14191), .A2(n14190), .ZN(n8617) );
  NAND2_X1 U11200 ( .A1(n14824), .A2(n14188), .ZN(n8618) );
  INV_X1 U11201 ( .A(n14406), .ZN(n14178) );
  NAND2_X1 U11202 ( .A1(n14809), .A2(n14178), .ZN(n8621) );
  INV_X1 U11203 ( .A(n8621), .ZN(n8623) );
  INV_X1 U11204 ( .A(n14407), .ZN(n14177) );
  NOR2_X1 U11205 ( .A1(n14817), .A2(n14177), .ZN(n14686) );
  INV_X1 U11206 ( .A(n14405), .ZN(n14204) );
  OR2_X1 U11207 ( .A1(n14809), .A2(n14178), .ZN(n14687) );
  OAI21_X1 U11208 ( .B1(n14697), .B2(n14204), .A(n14687), .ZN(n8620) );
  AOI21_X1 U11209 ( .B1(n14686), .B2(n8621), .A(n8620), .ZN(n8622) );
  NAND2_X1 U11210 ( .A1(n14697), .A2(n14204), .ZN(n8624) );
  INV_X1 U11211 ( .A(n14404), .ZN(n8626) );
  AND2_X1 U11212 ( .A1(n14800), .A2(n8626), .ZN(n8625) );
  INV_X1 U11213 ( .A(n14403), .ZN(n14076) );
  NAND2_X1 U11214 ( .A1(n14231), .A2(n14076), .ZN(n14647) );
  XNOR2_X1 U11215 ( .A(n14790), .B(n14402), .ZN(n14646) );
  INV_X1 U11216 ( .A(n14402), .ZN(n8630) );
  NAND2_X1 U11217 ( .A1(n14790), .A2(n8630), .ZN(n8631) );
  INV_X1 U11218 ( .A(n14401), .ZN(n14068) );
  OR2_X1 U11219 ( .A1(n14628), .A2(n14068), .ZN(n8632) );
  NAND2_X1 U11220 ( .A1(n14628), .A2(n14068), .ZN(n8633) );
  NAND2_X1 U11221 ( .A1(n14600), .A2(n14254), .ZN(n8636) );
  NOR2_X1 U11222 ( .A1(n14600), .A2(n14254), .ZN(n8635) );
  INV_X1 U11223 ( .A(n14577), .ZN(n14569) );
  XNOR2_X1 U11224 ( .A(n14562), .B(n14397), .ZN(n14560) );
  INV_X1 U11225 ( .A(n14397), .ZN(n14262) );
  NAND2_X1 U11226 ( .A1(n14562), .A2(n14262), .ZN(n8637) );
  INV_X1 U11227 ( .A(n14396), .ZN(n14266) );
  NAND2_X1 U11228 ( .A1(n14549), .A2(n14266), .ZN(n8638) );
  INV_X1 U11229 ( .A(n14395), .ZN(n14264) );
  NAND2_X1 U11230 ( .A1(n14105), .A2(n7740), .ZN(n14372) );
  NOR2_X1 U11231 ( .A1(n8641), .A2(n8640), .ZN(n8642) );
  NAND2_X1 U11232 ( .A1(n10418), .A2(n8642), .ZN(n8650) );
  NAND2_X1 U11233 ( .A1(n7741), .A2(n14105), .ZN(n11147) );
  INV_X1 U11234 ( .A(n11147), .ZN(n8649) );
  INV_X1 U11235 ( .A(n11179), .ZN(n11151) );
  NAND2_X1 U11236 ( .A1(n12989), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n8646) );
  NAND2_X1 U11237 ( .A1(n8643), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n8645) );
  NAND2_X1 U11238 ( .A1(n12988), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n8644) );
  AND3_X1 U11239 ( .A1(n8646), .A2(n8645), .A3(n8644), .ZN(n8647) );
  AOI22_X1 U11240 ( .A1(n14395), .A2(n14376), .B1(n14393), .B2(n14086), .ZN(
        n13118) );
  NAND2_X1 U11241 ( .A1(n8650), .A2(n13118), .ZN(n14516) );
  NAND2_X1 U11242 ( .A1(n8659), .A2(n8666), .ZN(n8652) );
  NAND2_X1 U11243 ( .A1(n8654), .A2(n8653), .ZN(n8663) );
  NAND2_X1 U11244 ( .A1(n8663), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8655) );
  MUX2_X1 U11245 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8655), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n8657) );
  NAND2_X1 U11246 ( .A1(n8658), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8667) );
  NAND2_X1 U11247 ( .A1(n8667), .A2(n8666), .ZN(n8669) );
  NAND2_X1 U11248 ( .A1(n8669), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8660) );
  NAND2_X1 U11249 ( .A1(n8661), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8662) );
  MUX2_X1 U11250 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8662), .S(
        P2_IR_REG_25__SCAN_IN), .Z(n8664) );
  NAND2_X1 U11251 ( .A1(n8664), .A2(n8663), .ZN(n12790) );
  NOR2_X1 U11252 ( .A1(n12582), .A2(n12790), .ZN(n8665) );
  NAND2_X1 U11253 ( .A1(n8683), .A2(n8665), .ZN(n11150) );
  OR2_X1 U11254 ( .A1(n8667), .A2(n8666), .ZN(n8668) );
  NAND2_X1 U11255 ( .A1(n8669), .A2(n8668), .ZN(n12320) );
  NOR4_X1 U11256 ( .A1(P2_D_REG_14__SCAN_IN), .A2(P2_D_REG_15__SCAN_IN), .A3(
        P2_D_REG_17__SCAN_IN), .A4(P2_D_REG_18__SCAN_IN), .ZN(n8673) );
  NOR4_X1 U11257 ( .A1(P2_D_REG_10__SCAN_IN), .A2(P2_D_REG_12__SCAN_IN), .A3(
        P2_D_REG_13__SCAN_IN), .A4(P2_D_REG_16__SCAN_IN), .ZN(n8672) );
  NOR4_X1 U11258 ( .A1(P2_D_REG_22__SCAN_IN), .A2(P2_D_REG_27__SCAN_IN), .A3(
        P2_D_REG_24__SCAN_IN), .A4(P2_D_REG_25__SCAN_IN), .ZN(n8671) );
  NOR4_X1 U11259 ( .A1(P2_D_REG_19__SCAN_IN), .A2(P2_D_REG_20__SCAN_IN), .A3(
        P2_D_REG_23__SCAN_IN), .A4(P2_D_REG_21__SCAN_IN), .ZN(n8670) );
  NAND4_X1 U11260 ( .A1(n8673), .A2(n8672), .A3(n8671), .A4(n8670), .ZN(n8680)
         );
  NOR4_X1 U11261 ( .A1(P2_D_REG_30__SCAN_IN), .A2(P2_D_REG_11__SCAN_IN), .A3(
        P2_D_REG_4__SCAN_IN), .A4(P2_D_REG_29__SCAN_IN), .ZN(n10828) );
  NOR2_X1 U11262 ( .A1(P2_D_REG_28__SCAN_IN), .A2(P2_D_REG_31__SCAN_IN), .ZN(
        n8676) );
  NOR4_X1 U11263 ( .A1(P2_D_REG_8__SCAN_IN), .A2(P2_D_REG_6__SCAN_IN), .A3(
        P2_D_REG_7__SCAN_IN), .A4(P2_D_REG_9__SCAN_IN), .ZN(n8675) );
  NOR4_X1 U11264 ( .A1(P2_D_REG_26__SCAN_IN), .A2(P2_D_REG_2__SCAN_IN), .A3(
        P2_D_REG_3__SCAN_IN), .A4(P2_D_REG_5__SCAN_IN), .ZN(n8674) );
  NAND4_X1 U11265 ( .A1(n10828), .A2(n8676), .A3(n8675), .A4(n8674), .ZN(n8679) );
  XNOR2_X1 U11266 ( .A(n12582), .B(P2_B_REG_SCAN_IN), .ZN(n8677) );
  NAND2_X1 U11267 ( .A1(n8677), .A2(n12790), .ZN(n8678) );
  OAI21_X1 U11268 ( .B1(n8680), .B2(n8679), .A(n15945), .ZN(n10561) );
  NAND2_X1 U11269 ( .A1(n15981), .A2(n10561), .ZN(n10554) );
  NAND2_X1 U11270 ( .A1(n8584), .A2(n14329), .ZN(n10557) );
  NAND2_X1 U11271 ( .A1(n10557), .A2(n7516), .ZN(n14270) );
  OR2_X1 U11272 ( .A1(n14270), .A2(n14379), .ZN(n10565) );
  INV_X1 U11273 ( .A(n10565), .ZN(n8681) );
  INV_X1 U11274 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n8682) );
  NAND2_X1 U11275 ( .A1(n15945), .A2(n8682), .ZN(n8685) );
  NAND2_X1 U11276 ( .A1(n14918), .A2(n12790), .ZN(n8684) );
  NAND2_X1 U11277 ( .A1(n8685), .A2(n8684), .ZN(n15980) );
  INV_X1 U11278 ( .A(n10396), .ZN(n10562) );
  NAND2_X1 U11279 ( .A1(n15980), .A2(n10562), .ZN(n8686) );
  INV_X1 U11280 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n8687) );
  NAND2_X1 U11281 ( .A1(n15945), .A2(n8687), .ZN(n8688) );
  NAND2_X1 U11282 ( .A1(n14918), .A2(n12582), .ZN(n15978) );
  NAND2_X1 U11283 ( .A1(n11909), .A2(n10557), .ZN(n15989) );
  NAND2_X1 U11284 ( .A1(n8689), .A2(n7974), .ZN(P2_U3527) );
  NOR2_X1 U11285 ( .A1(P3_IR_REG_12__SCAN_IN), .A2(P3_IR_REG_15__SCAN_IN), 
        .ZN(n8692) );
  NAND4_X1 U11286 ( .A1(n8774), .A2(n8726), .A3(n8762), .A4(n7082), .ZN(n8693)
         );
  NOR2_X2 U11287 ( .A1(n9363), .A2(P3_IR_REG_20__SCAN_IN), .ZN(n8796) );
  NAND2_X1 U11288 ( .A1(n8796), .A2(n8797), .ZN(n8793) );
  OAI21_X1 U11289 ( .B1(n8793), .B2(P3_IR_REG_22__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n8699) );
  INV_X1 U11290 ( .A(P3_IR_REG_23__SCAN_IN), .ZN(n8698) );
  XNOR2_X1 U11291 ( .A(n8699), .B(n8698), .ZN(n8799) );
  NAND4_X1 U11292 ( .A1(n8703), .A2(n8702), .A3(n8701), .A4(n8700), .ZN(n8706)
         );
  OAI21_X1 U11293 ( .B1(n8784), .B2(n8706), .A(n8705), .ZN(n8712) );
  INV_X1 U11294 ( .A(n8706), .ZN(n8708) );
  NAND2_X1 U11295 ( .A1(n8712), .A2(n8711), .ZN(n12986) );
  INV_X1 U11296 ( .A(n12986), .ZN(n8720) );
  NAND2_X1 U11297 ( .A1(n8716), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8714) );
  NAND2_X1 U11298 ( .A1(n7570), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8715) );
  MUX2_X1 U11299 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8715), .S(
        P3_IR_REG_25__SCAN_IN), .Z(n8717) );
  NAND2_X1 U11300 ( .A1(n8717), .A2(n8716), .ZN(n12296) );
  INV_X1 U11301 ( .A(n12296), .ZN(n8718) );
  AND2_X1 U11302 ( .A1(n9381), .A2(n8718), .ZN(n8719) );
  INV_X1 U11303 ( .A(n8792), .ZN(n11403) );
  OR2_X2 U11304 ( .A1(n13959), .A2(n11403), .ZN(n13510) );
  NAND2_X1 U11305 ( .A1(n8709), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8721) );
  XNOR2_X1 U11306 ( .A(n8721), .B(P3_IR_REG_16__SCAN_IN), .ZN(n13601) );
  INV_X1 U11307 ( .A(P3_REG2_REG_16__SCAN_IN), .ZN(n13808) );
  INV_X1 U11308 ( .A(n6560), .ZN(n8729) );
  NAND2_X1 U11309 ( .A1(n8725), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8724) );
  MUX2_X1 U11310 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8724), .S(
        P3_IR_REG_8__SCAN_IN), .Z(n8728) );
  INV_X1 U11311 ( .A(n8725), .ZN(n8727) );
  NAND2_X1 U11312 ( .A1(n8727), .A2(n8726), .ZN(n8752) );
  NAND2_X1 U11313 ( .A1(n8728), .A2(n8752), .ZN(n11703) );
  INV_X1 U11314 ( .A(n11703), .ZN(n8863) );
  INV_X1 U11315 ( .A(P3_REG2_REG_8__SCAN_IN), .ZN(n12273) );
  NAND2_X1 U11316 ( .A1(n8729), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8730) );
  XNOR2_X1 U11317 ( .A(n7082), .B(n8730), .ZN(n10739) );
  NAND2_X1 U11318 ( .A1(n8811), .A2(n6997), .ZN(n8743) );
  NAND2_X1 U11319 ( .A1(n8732), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8731) );
  MUX2_X1 U11320 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8731), .S(
        P3_IR_REG_4__SCAN_IN), .Z(n8735) );
  INV_X1 U11321 ( .A(n8732), .ZN(n8734) );
  INV_X1 U11322 ( .A(P3_IR_REG_4__SCAN_IN), .ZN(n8733) );
  NAND2_X1 U11323 ( .A1(n8734), .A2(n8733), .ZN(n8747) );
  INV_X1 U11324 ( .A(n8939), .ZN(n11312) );
  INV_X1 U11325 ( .A(P3_REG2_REG_0__SCAN_IN), .ZN(n8917) );
  NOR2_X1 U11326 ( .A1(n8917), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n8740) );
  NAND2_X1 U11327 ( .A1(n8811), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n8741) );
  OAI21_X1 U11328 ( .B1(n8836), .B2(n8740), .A(n8741), .ZN(n11285) );
  INV_X1 U11329 ( .A(P3_REG2_REG_1__SCAN_IN), .ZN(n16064) );
  NOR2_X1 U11330 ( .A1(n11285), .A2(n16064), .ZN(n11284) );
  INV_X1 U11331 ( .A(n8741), .ZN(n8742) );
  NOR2_X1 U11332 ( .A1(n11284), .A2(n8742), .ZN(n11298) );
  NAND2_X1 U11333 ( .A1(n8743), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8744) );
  INV_X1 U11334 ( .A(n8746), .ZN(n11266) );
  XNOR2_X1 U11335 ( .A(n10662), .B(P3_REG2_REG_4__SCAN_IN), .ZN(n11267) );
  NAND2_X1 U11336 ( .A1(n8747), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8748) );
  XNOR2_X1 U11337 ( .A(n8748), .B(P3_IR_REG_5__SCAN_IN), .ZN(n8962) );
  XNOR2_X1 U11338 ( .A(n10739), .B(P3_REG2_REG_6__SCAN_IN), .ZN(n11392) );
  NAND2_X1 U11339 ( .A1(n8749), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8750) );
  XNOR2_X1 U11340 ( .A(n8750), .B(P3_IR_REG_7__SCAN_IN), .ZN(n9006) );
  INV_X1 U11341 ( .A(P3_REG2_REG_7__SCAN_IN), .ZN(n12132) );
  XNOR2_X1 U11342 ( .A(n11703), .B(n12273), .ZN(n11688) );
  OAI21_X1 U11343 ( .B1(n8863), .B2(n12273), .A(n11691), .ZN(n8754) );
  INV_X1 U11344 ( .A(n8754), .ZN(n8755) );
  NAND2_X1 U11345 ( .A1(n8752), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8751) );
  MUX2_X1 U11346 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8751), .S(
        P3_IR_REG_9__SCAN_IN), .Z(n8753) );
  NAND2_X1 U11347 ( .A1(n8753), .A2(n8759), .ZN(n12061) );
  INV_X1 U11348 ( .A(n12061), .ZN(n8867) );
  NAND2_X1 U11349 ( .A1(n8759), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8757) );
  INV_X1 U11350 ( .A(P3_IR_REG_10__SCAN_IN), .ZN(n8760) );
  XNOR2_X1 U11351 ( .A(n8757), .B(n8760), .ZN(n10671) );
  XNOR2_X1 U11352 ( .A(n10671), .B(P3_REG2_REG_10__SCAN_IN), .ZN(n10589) );
  INV_X1 U11353 ( .A(n10671), .ZN(n8871) );
  INV_X1 U11354 ( .A(P3_REG2_REG_10__SCAN_IN), .ZN(n12624) );
  NOR2_X1 U11355 ( .A1(n8871), .A2(n12624), .ZN(n8758) );
  NAND2_X1 U11356 ( .A1(n8761), .A2(n8760), .ZN(n8766) );
  NAND2_X1 U11357 ( .A1(n8766), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8763) );
  XNOR2_X1 U11358 ( .A(n8763), .B(n8762), .ZN(n12601) );
  INV_X1 U11359 ( .A(n12601), .ZN(n8878) );
  NAND2_X1 U11360 ( .A1(n8768), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8767) );
  MUX2_X1 U11361 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8767), .S(
        P3_IR_REG_12__SCAN_IN), .Z(n8771) );
  INV_X1 U11362 ( .A(P3_IR_REG_12__SCAN_IN), .ZN(n8769) );
  NAND2_X1 U11363 ( .A1(n8770), .A2(n8769), .ZN(n8776) );
  NAND2_X1 U11364 ( .A1(n13515), .A2(P3_REG2_REG_12__SCAN_IN), .ZN(n8773) );
  OAI21_X1 U11365 ( .B1(n13515), .B2(P3_REG2_REG_12__SCAN_IN), .A(n8773), .ZN(
        n8772) );
  INV_X1 U11366 ( .A(n8772), .ZN(n13513) );
  NAND2_X1 U11367 ( .A1(n13512), .A2(n13513), .ZN(n13511) );
  NAND2_X1 U11368 ( .A1(n8776), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8775) );
  XNOR2_X1 U11369 ( .A(n8775), .B(n8774), .ZN(n13543) );
  INV_X1 U11370 ( .A(P3_REG2_REG_13__SCAN_IN), .ZN(n13532) );
  NAND2_X1 U11371 ( .A1(n8780), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8778) );
  INV_X1 U11372 ( .A(P3_IR_REG_14__SCAN_IN), .ZN(n8777) );
  XNOR2_X1 U11373 ( .A(n8778), .B(n8777), .ZN(n11129) );
  XNOR2_X1 U11374 ( .A(n11129), .B(P3_REG2_REG_14__SCAN_IN), .ZN(n8885) );
  INV_X1 U11375 ( .A(n13551), .ZN(n8779) );
  INV_X1 U11376 ( .A(n11129), .ZN(n13562) );
  INV_X1 U11377 ( .A(P3_REG2_REG_14__SCAN_IN), .ZN(n9130) );
  OAI21_X1 U11378 ( .B1(n8780), .B2(P3_IR_REG_14__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n8781) );
  XNOR2_X1 U11379 ( .A(n8781), .B(P3_IR_REG_15__SCAN_IN), .ZN(n13582) );
  INV_X1 U11380 ( .A(n13582), .ZN(n11126) );
  INV_X1 U11381 ( .A(P3_REG2_REG_15__SCAN_IN), .ZN(n13821) );
  XNOR2_X1 U11382 ( .A(n13601), .B(P3_REG2_REG_16__SCAN_IN), .ZN(n13589) );
  NAND2_X1 U11383 ( .A1(n6723), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8783) );
  XNOR2_X1 U11384 ( .A(n8783), .B(P3_IR_REG_17__SCAN_IN), .ZN(n9171) );
  INV_X1 U11385 ( .A(n9171), .ZN(n13616) );
  NAND2_X1 U11386 ( .A1(n8784), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8785) );
  XNOR2_X1 U11387 ( .A(n8785), .B(P3_IR_REG_18__SCAN_IN), .ZN(n13641) );
  INV_X1 U11388 ( .A(P3_REG2_REG_18__SCAN_IN), .ZN(n8786) );
  OR2_X1 U11389 ( .A1(n13641), .A2(n8786), .ZN(n8788) );
  NAND2_X1 U11390 ( .A1(n13641), .A2(n8786), .ZN(n8787) );
  NAND2_X1 U11391 ( .A1(n8788), .A2(n8787), .ZN(n13623) );
  NAND2_X1 U11392 ( .A1(n8789), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8790) );
  XNOR2_X1 U11393 ( .A(n13306), .B(P3_REG2_REG_19__SCAN_IN), .ZN(n8894) );
  XNOR2_X1 U11394 ( .A(n8791), .B(n8894), .ZN(n8901) );
  OR2_X1 U11395 ( .A1(n8799), .A2(P3_U3151), .ZN(n13490) );
  NAND2_X1 U11396 ( .A1(n11422), .A2(n13490), .ZN(n8833) );
  NAND2_X1 U11397 ( .A1(n8793), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8795) );
  INV_X1 U11398 ( .A(P3_IR_REG_22__SCAN_IN), .ZN(n8794) );
  NAND2_X1 U11399 ( .A1(n13468), .A2(n8799), .ZN(n8806) );
  INV_X1 U11400 ( .A(P3_IR_REG_26__SCAN_IN), .ZN(n8800) );
  NAND2_X1 U11401 ( .A1(n8806), .A2(n9367), .ZN(n8832) );
  INV_X1 U11402 ( .A(n8832), .ZN(n8807) );
  INV_X1 U11403 ( .A(n8831), .ZN(n8810) );
  INV_X1 U11404 ( .A(n8808), .ZN(n9375) );
  NAND2_X1 U11405 ( .A1(n9375), .A2(n13485), .ZN(n9366) );
  INV_X1 U11406 ( .A(P3_REG1_REG_10__SCAN_IN), .ZN(n12733) );
  INV_X1 U11407 ( .A(n8836), .ZN(n8834) );
  NAND2_X1 U11408 ( .A1(n6771), .A2(P3_REG1_REG_0__SCAN_IN), .ZN(n8812) );
  NAND2_X1 U11409 ( .A1(n11287), .A2(P3_REG1_REG_1__SCAN_IN), .ZN(n11286) );
  INV_X1 U11410 ( .A(n8813), .ZN(n8814) );
  NAND2_X1 U11411 ( .A1(n11286), .A2(n8814), .ZN(n11295) );
  XNOR2_X1 U11412 ( .A(n8939), .B(P3_REG1_REG_2__SCAN_IN), .ZN(n11296) );
  INV_X1 U11413 ( .A(P3_REG1_REG_2__SCAN_IN), .ZN(n8929) );
  NAND2_X1 U11414 ( .A1(n8815), .A2(n7696), .ZN(n11270) );
  INV_X1 U11415 ( .A(P3_REG1_REG_3__SCAN_IN), .ZN(n11317) );
  XNOR2_X1 U11416 ( .A(n10739), .B(P3_REG1_REG_6__SCAN_IN), .ZN(n11396) );
  INV_X1 U11417 ( .A(n8819), .ZN(n11696) );
  XNOR2_X1 U11418 ( .A(n11703), .B(P3_REG1_REG_8__SCAN_IN), .ZN(n11697) );
  INV_X1 U11419 ( .A(P3_REG1_REG_9__SCAN_IN), .ZN(n12050) );
  XNOR2_X1 U11420 ( .A(n10671), .B(n12733), .ZN(n10592) );
  OAI21_X1 U11421 ( .B1(n8871), .B2(n12733), .A(n10595), .ZN(n8820) );
  INV_X1 U11422 ( .A(P3_REG1_REG_11__SCAN_IN), .ZN(n12593) );
  XNOR2_X1 U11423 ( .A(n13515), .B(P3_REG1_REG_12__SCAN_IN), .ZN(n13524) );
  INV_X1 U11424 ( .A(n13543), .ZN(n8822) );
  NAND2_X1 U11425 ( .A1(n11129), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n8886) );
  OR2_X1 U11426 ( .A1(n11129), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n8825) );
  AND2_X1 U11427 ( .A1(n8886), .A2(n8825), .ZN(n13564) );
  INV_X1 U11428 ( .A(P3_REG1_REG_15__SCAN_IN), .ZN(n13879) );
  XNOR2_X1 U11429 ( .A(n13601), .B(P3_REG1_REG_16__SCAN_IN), .ZN(n13603) );
  INV_X1 U11430 ( .A(P3_REG1_REG_16__SCAN_IN), .ZN(n13876) );
  INV_X1 U11431 ( .A(P3_REG1_REG_17__SCAN_IN), .ZN(n13872) );
  INV_X1 U11432 ( .A(P3_REG1_REG_18__SCAN_IN), .ZN(n13870) );
  OR2_X1 U11433 ( .A1(n13641), .A2(n13870), .ZN(n8828) );
  NAND2_X1 U11434 ( .A1(n13641), .A2(n13870), .ZN(n8827) );
  NAND2_X1 U11435 ( .A1(n8828), .A2(n8827), .ZN(n13628) );
  AOI21_X1 U11436 ( .B1(n13630), .B2(n13629), .A(n13628), .ZN(n13633) );
  INV_X1 U11437 ( .A(n8828), .ZN(n8829) );
  XNOR2_X1 U11438 ( .A(n13332), .B(P3_REG1_REG_19__SCAN_IN), .ZN(n8897) );
  INV_X2 U11439 ( .A(n13485), .ZN(n8892) );
  MUX2_X1 U11440 ( .A(P3_U3897), .B(n8831), .S(n8808), .Z(n16021) );
  INV_X1 U11441 ( .A(n16012), .ZN(n16024) );
  NAND2_X1 U11442 ( .A1(P3_U3151), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n13167)
         );
  OAI21_X1 U11443 ( .B1(n16024), .B2(n15768), .A(n13167), .ZN(n8900) );
  MUX2_X1 U11444 ( .A(P3_REG2_REG_17__SCAN_IN), .B(P3_REG1_REG_17__SCAN_IN), 
        .S(n8892), .Z(n8891) );
  INV_X1 U11445 ( .A(P3_REG1_REG_1__SCAN_IN), .ZN(n16095) );
  INV_X1 U11446 ( .A(n8835), .ZN(n8837) );
  NAND2_X1 U11447 ( .A1(n8837), .A2(n8836), .ZN(n8838) );
  INV_X1 U11448 ( .A(P3_REG1_REG_0__SCAN_IN), .ZN(n8918) );
  MUX2_X1 U11449 ( .A(n8917), .B(n8918), .S(n8895), .Z(n16017) );
  NAND2_X1 U11450 ( .A1(n16017), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n16016) );
  NAND2_X1 U11451 ( .A1(n11281), .A2(n11300), .ZN(n8842) );
  MUX2_X1 U11452 ( .A(n7654), .B(n8929), .S(n8895), .Z(n8839) );
  NAND2_X1 U11453 ( .A1(n8839), .A2(n8939), .ZN(n11324) );
  INV_X1 U11454 ( .A(n8839), .ZN(n8840) );
  NAND2_X1 U11455 ( .A1(n8840), .A2(n11312), .ZN(n8841) );
  AND2_X1 U11456 ( .A1(n11324), .A2(n8841), .ZN(n11301) );
  NAND2_X1 U11457 ( .A1(n8842), .A2(n11301), .ZN(n11303) );
  INV_X1 U11458 ( .A(P3_REG2_REG_3__SCAN_IN), .ZN(n11682) );
  MUX2_X1 U11459 ( .A(n11682), .B(n11317), .S(n8895), .Z(n8843) );
  NAND2_X1 U11460 ( .A1(n8843), .A2(n8981), .ZN(n11260) );
  INV_X1 U11461 ( .A(n8843), .ZN(n8844) );
  NAND2_X1 U11462 ( .A1(n8844), .A2(n7696), .ZN(n8845) );
  AND2_X1 U11463 ( .A1(n11260), .A2(n8845), .ZN(n11325) );
  INV_X1 U11464 ( .A(P3_REG2_REG_4__SCAN_IN), .ZN(n11883) );
  INV_X1 U11465 ( .A(P3_REG1_REG_4__SCAN_IN), .ZN(n8846) );
  MUX2_X1 U11466 ( .A(n11883), .B(n8846), .S(n8895), .Z(n8847) );
  INV_X1 U11467 ( .A(n10662), .ZN(n11278) );
  NAND2_X1 U11468 ( .A1(n8847), .A2(n11278), .ZN(n11251) );
  INV_X1 U11469 ( .A(n8847), .ZN(n8848) );
  NAND2_X1 U11470 ( .A1(n8848), .A2(n10662), .ZN(n8849) );
  AND2_X1 U11471 ( .A1(n11251), .A2(n8849), .ZN(n11261) );
  NAND2_X1 U11472 ( .A1(n11250), .A2(n11251), .ZN(n8853) );
  INV_X1 U11473 ( .A(P3_REG2_REG_5__SCAN_IN), .ZN(n8945) );
  INV_X1 U11474 ( .A(P3_REG1_REG_5__SCAN_IN), .ZN(n16099) );
  MUX2_X1 U11475 ( .A(n8945), .B(n16099), .S(n8892), .Z(n8850) );
  NAND2_X1 U11476 ( .A1(n8850), .A2(n8962), .ZN(n11384) );
  INV_X1 U11477 ( .A(n8850), .ZN(n8851) );
  NAND2_X1 U11478 ( .A1(n8851), .A2(n7646), .ZN(n8852) );
  AND2_X1 U11479 ( .A1(n11384), .A2(n8852), .ZN(n11252) );
  NAND2_X1 U11480 ( .A1(n11388), .A2(n11384), .ZN(n8858) );
  INV_X1 U11481 ( .A(P3_REG2_REG_6__SCAN_IN), .ZN(n9012) );
  INV_X1 U11482 ( .A(P3_REG1_REG_6__SCAN_IN), .ZN(n8854) );
  MUX2_X1 U11483 ( .A(n9012), .B(n8854), .S(n8892), .Z(n8855) );
  NAND2_X1 U11484 ( .A1(n8855), .A2(n7234), .ZN(n11539) );
  INV_X1 U11485 ( .A(n8855), .ZN(n8856) );
  NAND2_X1 U11486 ( .A1(n8856), .A2(n10739), .ZN(n8857) );
  AND2_X1 U11487 ( .A1(n11539), .A2(n8857), .ZN(n11386) );
  NAND2_X1 U11488 ( .A1(n8858), .A2(n11386), .ZN(n11387) );
  NAND2_X1 U11489 ( .A1(n11387), .A2(n11539), .ZN(n8862) );
  INV_X1 U11490 ( .A(P3_REG1_REG_7__SCAN_IN), .ZN(n16101) );
  MUX2_X1 U11491 ( .A(n12132), .B(n16101), .S(n8892), .Z(n8859) );
  NAND2_X1 U11492 ( .A1(n8859), .A2(n9006), .ZN(n11693) );
  INV_X1 U11493 ( .A(n8859), .ZN(n8860) );
  NAND2_X1 U11494 ( .A1(n8860), .A2(n7718), .ZN(n8861) );
  AND2_X1 U11495 ( .A1(n11693), .A2(n8861), .ZN(n11540) );
  INV_X1 U11496 ( .A(P3_REG1_REG_8__SCAN_IN), .ZN(n16104) );
  MUX2_X1 U11497 ( .A(n12273), .B(n16104), .S(n8892), .Z(n8864) );
  NAND2_X1 U11498 ( .A1(n8864), .A2(n8863), .ZN(n12055) );
  INV_X1 U11499 ( .A(n8864), .ZN(n8865) );
  NAND2_X1 U11500 ( .A1(n8865), .A2(n11703), .ZN(n8866) );
  AND2_X1 U11501 ( .A1(n12055), .A2(n8866), .ZN(n11692) );
  INV_X1 U11502 ( .A(P3_REG2_REG_9__SCAN_IN), .ZN(n12117) );
  MUX2_X1 U11503 ( .A(n12117), .B(n12050), .S(n8892), .Z(n8868) );
  NAND2_X1 U11504 ( .A1(n8868), .A2(n8867), .ZN(n10598) );
  INV_X1 U11505 ( .A(n8868), .ZN(n8869) );
  NAND2_X1 U11506 ( .A1(n8869), .A2(n12061), .ZN(n8870) );
  AND2_X1 U11507 ( .A1(n10598), .A2(n8870), .ZN(n12053) );
  NAND2_X1 U11508 ( .A1(n12058), .A2(n10598), .ZN(n8875) );
  MUX2_X1 U11509 ( .A(n12624), .B(n12733), .S(n8892), .Z(n8872) );
  NAND2_X1 U11510 ( .A1(n8872), .A2(n8871), .ZN(n8876) );
  INV_X1 U11511 ( .A(n8872), .ZN(n8873) );
  NAND2_X1 U11512 ( .A1(n8873), .A2(n10671), .ZN(n8874) );
  AND2_X1 U11513 ( .A1(n8876), .A2(n8874), .ZN(n10596) );
  NAND2_X1 U11514 ( .A1(n8875), .A2(n10596), .ZN(n10600) );
  NAND2_X1 U11515 ( .A1(n10600), .A2(n8876), .ZN(n12599) );
  MUX2_X1 U11516 ( .A(P3_REG2_REG_11__SCAN_IN), .B(P3_REG1_REG_11__SCAN_IN), 
        .S(n8892), .Z(n8877) );
  XNOR2_X1 U11517 ( .A(n8877), .B(n8878), .ZN(n12598) );
  NAND2_X1 U11518 ( .A1(n12599), .A2(n12598), .ZN(n12597) );
  INV_X1 U11519 ( .A(n8877), .ZN(n8879) );
  NAND2_X1 U11520 ( .A1(n8879), .A2(n8878), .ZN(n8880) );
  NAND2_X1 U11521 ( .A1(n12597), .A2(n8880), .ZN(n13519) );
  MUX2_X1 U11522 ( .A(P3_REG2_REG_12__SCAN_IN), .B(P3_REG1_REG_12__SCAN_IN), 
        .S(n8892), .Z(n8881) );
  XNOR2_X1 U11523 ( .A(n8881), .B(n13515), .ZN(n13520) );
  INV_X1 U11524 ( .A(P3_REG1_REG_13__SCAN_IN), .ZN(n12711) );
  MUX2_X1 U11525 ( .A(n13532), .B(n12711), .S(n8892), .Z(n8883) );
  XNOR2_X1 U11526 ( .A(n13543), .B(n8883), .ZN(n13534) );
  NAND2_X1 U11527 ( .A1(n8881), .A2(n13515), .ZN(n13535) );
  AND2_X1 U11528 ( .A1(n13534), .A2(n13535), .ZN(n8882) );
  INV_X1 U11529 ( .A(n8883), .ZN(n8884) );
  OR2_X1 U11530 ( .A1(n13543), .A2(n8884), .ZN(n13557) );
  INV_X1 U11531 ( .A(n8885), .ZN(n13549) );
  MUX2_X1 U11532 ( .A(n13549), .B(n13564), .S(n8892), .Z(n13556) );
  MUX2_X1 U11533 ( .A(n7979), .B(n8886), .S(n8892), .Z(n8887) );
  INV_X1 U11534 ( .A(n8888), .ZN(n8889) );
  XOR2_X1 U11535 ( .A(n13582), .B(n8888), .Z(n13578) );
  MUX2_X1 U11536 ( .A(P3_REG2_REG_15__SCAN_IN), .B(P3_REG1_REG_15__SCAN_IN), 
        .S(n8892), .Z(n13577) );
  NOR2_X1 U11537 ( .A1(n13578), .A2(n13577), .ZN(n13576) );
  MUX2_X1 U11538 ( .A(n13808), .B(n13876), .S(n8892), .Z(n8890) );
  NOR2_X1 U11539 ( .A1(n8890), .A2(n13601), .ZN(n13595) );
  NAND2_X1 U11540 ( .A1(n8890), .A2(n13601), .ZN(n13594) );
  XOR2_X1 U11541 ( .A(n9171), .B(n8891), .Z(n13613) );
  MUX2_X1 U11542 ( .A(P3_REG2_REG_18__SCAN_IN), .B(P3_REG1_REG_18__SCAN_IN), 
        .S(n8892), .Z(n13637) );
  NOR2_X1 U11543 ( .A1(n13636), .A2(n13637), .ZN(n13635) );
  AOI21_X1 U11544 ( .B1(n8893), .B2(n13641), .A(n13635), .ZN(n8899) );
  INV_X1 U11545 ( .A(n8894), .ZN(n8896) );
  INV_X1 U11546 ( .A(n8895), .ZN(n13485) );
  MUX2_X1 U11547 ( .A(n8897), .B(n8896), .S(n13485), .Z(n8898) );
  XNOR2_X2 U11548 ( .A(n8902), .B(P3_IR_REG_30__SCAN_IN), .ZN(n8906) );
  INV_X1 U11549 ( .A(P3_REG3_REG_1__SCAN_IN), .ZN(n11445) );
  NAND2_X2 U11550 ( .A1(n8906), .A2(n8905), .ZN(n9311) );
  OR2_X1 U11551 ( .A1(n8974), .A2(n16095), .ZN(n8908) );
  OR2_X1 U11552 ( .A1(n13292), .A2(n10731), .ZN(n8916) );
  NAND2_X2 U11553 ( .A1(n16030), .A2(n16056), .ZN(n13342) );
  NAND2_X1 U11554 ( .A1(n13285), .A2(P3_REG0_REG_0__SCAN_IN), .ZN(n8922) );
  INV_X1 U11555 ( .A(P3_REG3_REG_0__SCAN_IN), .ZN(n11429) );
  OR2_X1 U11556 ( .A1(n9126), .A2(n11429), .ZN(n8921) );
  OR2_X1 U11557 ( .A1(n9311), .A2(n8917), .ZN(n8920) );
  OR2_X1 U11558 ( .A1(n8974), .A2(n8918), .ZN(n8919) );
  NAND4_X2 U11559 ( .A1(n8922), .A2(n8921), .A3(n8920), .A4(n8919), .ZN(n16048) );
  INV_X1 U11560 ( .A(SI_0_), .ZN(n10735) );
  OR2_X1 U11561 ( .A1(n13292), .A2(n10735), .ZN(n8926) );
  INV_X1 U11562 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n9497) );
  NAND2_X1 U11563 ( .A1(n9497), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n8923) );
  AND2_X1 U11564 ( .A1(n8934), .A2(n8923), .ZN(n10736) );
  OR2_X1 U11565 ( .A1(n9353), .A2(n10736), .ZN(n8925) );
  INV_X1 U11566 ( .A(n11845), .ZN(n11600) );
  NAND2_X1 U11567 ( .A1(n16052), .A2(n16043), .ZN(n8928) );
  INV_X1 U11568 ( .A(n16030), .ZN(n11432) );
  NAND2_X1 U11569 ( .A1(n16056), .A2(n11432), .ZN(n8927) );
  NAND2_X1 U11570 ( .A1(n6567), .A2(P3_REG0_REG_2__SCAN_IN), .ZN(n8933) );
  INV_X1 U11571 ( .A(P3_REG3_REG_2__SCAN_IN), .ZN(n11508) );
  OR2_X1 U11572 ( .A1(n9126), .A2(n11508), .ZN(n8932) );
  NAND2_X1 U11573 ( .A1(n10750), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n8935) );
  NAND2_X1 U11574 ( .A1(n10820), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n8936) );
  XNOR2_X1 U11575 ( .A(n8951), .B(n8950), .ZN(n10666) );
  OR2_X1 U11576 ( .A1(n9353), .A2(n10666), .ZN(n8938) );
  NAND2_X1 U11577 ( .A1(n16025), .A2(n13347), .ZN(n8941) );
  NAND2_X1 U11578 ( .A1(n7260), .A2(n16036), .ZN(n8940) );
  NAND2_X1 U11579 ( .A1(n13285), .A2(P3_REG0_REG_5__SCAN_IN), .ZN(n8949) );
  OR2_X1 U11580 ( .A1(n9372), .A2(n16099), .ZN(n8948) );
  NAND2_X1 U11581 ( .A1(n8965), .A2(P3_REG3_REG_5__SCAN_IN), .ZN(n8944) );
  AND2_X1 U11582 ( .A1(n9009), .A2(n8944), .ZN(n12100) );
  OR2_X1 U11583 ( .A1(n9126), .A2(n12100), .ZN(n8947) );
  OR2_X1 U11584 ( .A1(n9311), .A2(n8945), .ZN(n8946) );
  NAND4_X2 U11585 ( .A1(n8949), .A2(n8948), .A3(n8947), .A4(n8946), .ZN(n13508) );
  NAND2_X1 U11586 ( .A1(n8951), .A2(n8950), .ZN(n8953) );
  NAND2_X1 U11587 ( .A1(n10639), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n8954) );
  NAND2_X1 U11588 ( .A1(n8980), .A2(n8979), .ZN(n8956) );
  NAND2_X1 U11589 ( .A1(n10655), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n8957) );
  NAND2_X1 U11590 ( .A1(n10692), .A2(P1_DATAO_REG_5__SCAN_IN), .ZN(n8959) );
  XNOR2_X1 U11591 ( .A(n8995), .B(n8994), .ZN(n10657) );
  OR2_X1 U11592 ( .A1(n9353), .A2(n10657), .ZN(n8961) );
  OR2_X1 U11593 ( .A1(n6568), .A2(SI_5_), .ZN(n8960) );
  OAI211_X1 U11594 ( .C1(n8962), .C2(n9367), .A(n8961), .B(n8960), .ZN(n12099)
         );
  NAND2_X1 U11595 ( .A1(n13508), .A2(n12099), .ZN(n13364) );
  NAND2_X2 U11596 ( .A1(n13359), .A2(n13364), .ZN(n13313) );
  NAND2_X1 U11597 ( .A1(n9357), .A2(P3_REG1_REG_4__SCAN_IN), .ZN(n8969) );
  INV_X1 U11598 ( .A(P3_REG0_REG_4__SCAN_IN), .ZN(n8963) );
  OR2_X1 U11599 ( .A1(n9007), .A2(n8963), .ZN(n8968) );
  NAND2_X1 U11600 ( .A1(P3_REG3_REG_3__SCAN_IN), .A2(P3_REG3_REG_4__SCAN_IN), 
        .ZN(n8964) );
  AND2_X1 U11601 ( .A1(n8965), .A2(n8964), .ZN(n11658) );
  OR2_X1 U11602 ( .A1(n9311), .A2(n11883), .ZN(n8966) );
  OR2_X1 U11603 ( .A1(n6569), .A2(SI_4_), .ZN(n8970) );
  XNOR2_X1 U11604 ( .A(n8972), .B(n8971), .ZN(n10660) );
  OR2_X1 U11605 ( .A1(n9353), .A2(n10660), .ZN(n8973) );
  NAND2_X1 U11606 ( .A1(n6566), .A2(P3_REG0_REG_3__SCAN_IN), .ZN(n8978) );
  OR2_X1 U11607 ( .A1(n9126), .A2(P3_REG3_REG_3__SCAN_IN), .ZN(n8977) );
  OR2_X1 U11608 ( .A1(n9311), .A2(n11682), .ZN(n8976) );
  OR2_X1 U11609 ( .A1(n8974), .A2(n11317), .ZN(n8975) );
  NAND4_X1 U11610 ( .A1(n8978), .A2(n8977), .A3(n8976), .A4(n8975), .ZN(n16031) );
  OR2_X1 U11611 ( .A1(n6568), .A2(SI_3_), .ZN(n8983) );
  XNOR2_X1 U11612 ( .A(n8980), .B(n8979), .ZN(n10732) );
  OR2_X1 U11613 ( .A1(n9353), .A2(n10732), .ZN(n8982) );
  AND2_X1 U11614 ( .A1(n16031), .A2(n12123), .ZN(n11783) );
  INV_X1 U11615 ( .A(n11974), .ZN(n11886) );
  AOI21_X2 U11616 ( .B1(n13355), .B2(n11783), .A(n8984), .ZN(n12101) );
  OR2_X1 U11617 ( .A1(n16031), .A2(n11647), .ZN(n13354) );
  NAND2_X1 U11618 ( .A1(n16031), .A2(n11647), .ZN(n13351) );
  NAND2_X1 U11619 ( .A1(n13354), .A2(n13351), .ZN(n11639) );
  NAND2_X1 U11620 ( .A1(n11639), .A2(n13355), .ZN(n12102) );
  INV_X1 U11621 ( .A(n13508), .ZN(n12286) );
  NAND2_X1 U11622 ( .A1(n12286), .A2(n12099), .ZN(n8985) );
  NAND2_X1 U11623 ( .A1(n13285), .A2(P3_REG0_REG_7__SCAN_IN), .ZN(n8993) );
  OR2_X1 U11624 ( .A1(n9372), .A2(n16101), .ZN(n8992) );
  NAND2_X1 U11625 ( .A1(n9011), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n8989) );
  AND2_X1 U11626 ( .A1(n9023), .A2(n8989), .ZN(n12316) );
  OR2_X1 U11627 ( .A1(n9126), .A2(n12316), .ZN(n8991) );
  OR2_X1 U11628 ( .A1(n9311), .A2(n12132), .ZN(n8990) );
  OR2_X1 U11629 ( .A1(n6568), .A2(SI_7_), .ZN(n9005) );
  NAND2_X1 U11630 ( .A1(n10779), .A2(P1_DATAO_REG_6__SCAN_IN), .ZN(n8997) );
  NAND2_X1 U11631 ( .A1(n10707), .A2(P2_DATAO_REG_6__SCAN_IN), .ZN(n8998) );
  NAND2_X1 U11632 ( .A1(n10964), .A2(P2_DATAO_REG_7__SCAN_IN), .ZN(n9000) );
  NAND2_X1 U11633 ( .A1(n9029), .A2(n9000), .ZN(n9001) );
  NAND2_X1 U11634 ( .A1(n9002), .A2(n9001), .ZN(n9003) );
  AND2_X1 U11635 ( .A1(n9030), .A2(n9003), .ZN(n10663) );
  OR2_X1 U11636 ( .A1(n9353), .A2(n10663), .ZN(n9004) );
  OAI211_X1 U11637 ( .C1(n9006), .C2(n9367), .A(n9005), .B(n9004), .ZN(n12134)
         );
  NAND2_X1 U11638 ( .A1(n9357), .A2(P3_REG1_REG_6__SCAN_IN), .ZN(n9016) );
  INV_X1 U11639 ( .A(P3_REG0_REG_6__SCAN_IN), .ZN(n9008) );
  OR2_X1 U11640 ( .A1(n9007), .A2(n9008), .ZN(n9015) );
  NAND2_X1 U11641 ( .A1(n9009), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n9010) );
  AND2_X1 U11642 ( .A1(n9011), .A2(n9010), .ZN(n12292) );
  OR2_X1 U11643 ( .A1(n9126), .A2(n12292), .ZN(n9014) );
  OR2_X1 U11644 ( .A1(n9311), .A2(n9012), .ZN(n9013) );
  XNOR2_X1 U11645 ( .A(n10779), .B(P1_DATAO_REG_6__SCAN_IN), .ZN(n9017) );
  XNOR2_X1 U11646 ( .A(n9018), .B(n9017), .ZN(n10738) );
  OR2_X1 U11647 ( .A1(n9353), .A2(n10738), .ZN(n9021) );
  INV_X1 U11648 ( .A(SI_6_), .ZN(n10737) );
  OR2_X1 U11649 ( .A1(n6568), .A2(n10737), .ZN(n9020) );
  OR2_X1 U11650 ( .A1(n9367), .A2(n10739), .ZN(n9019) );
  INV_X1 U11651 ( .A(n12245), .ZN(n12289) );
  AND2_X1 U11652 ( .A1(n13507), .A2(n12289), .ZN(n12126) );
  INV_X1 U11653 ( .A(n12134), .ZN(n12313) );
  AND2_X1 U11654 ( .A1(n13506), .A2(n12313), .ZN(n9022) );
  NAND2_X1 U11655 ( .A1(n6567), .A2(P3_REG0_REG_8__SCAN_IN), .ZN(n9028) );
  NAND2_X1 U11656 ( .A1(n9023), .A2(P3_REG3_REG_8__SCAN_IN), .ZN(n9024) );
  AND2_X1 U11657 ( .A1(n9049), .A2(n9024), .ZN(n12483) );
  OR2_X1 U11658 ( .A1(n9126), .A2(n12483), .ZN(n9026) );
  OR2_X1 U11659 ( .A1(n9311), .A2(n12273), .ZN(n9025) );
  NAND2_X1 U11660 ( .A1(n10713), .A2(P2_DATAO_REG_8__SCAN_IN), .ZN(n9031) );
  OR2_X1 U11661 ( .A1(n9033), .A2(n9032), .ZN(n9034) );
  NAND2_X1 U11662 ( .A1(n9044), .A2(n9034), .ZN(n10640) );
  OR2_X1 U11663 ( .A1(n10640), .A2(n9353), .ZN(n9037) );
  INV_X1 U11664 ( .A(SI_8_), .ZN(n10641) );
  OR2_X1 U11665 ( .A1(n6568), .A2(n10641), .ZN(n9036) );
  OR2_X1 U11666 ( .A1(n9367), .A2(n11703), .ZN(n9035) );
  NAND2_X1 U11667 ( .A1(n13505), .A2(n12274), .ZN(n13378) );
  OR2_X1 U11668 ( .A1(n13507), .A2(n12245), .ZN(n13365) );
  NAND2_X1 U11669 ( .A1(n13507), .A2(n12245), .ZN(n13372) );
  NAND2_X1 U11670 ( .A1(n13365), .A2(n13372), .ZN(n9406) );
  NAND2_X1 U11671 ( .A1(n9406), .A2(n12246), .ZN(n12268) );
  NAND2_X1 U11672 ( .A1(n12268), .A2(n13373), .ZN(n9039) );
  INV_X1 U11673 ( .A(n12267), .ZN(n9038) );
  INV_X1 U11674 ( .A(n12274), .ZN(n12480) );
  OAI22_X1 U11675 ( .A1(n9039), .A2(n9038), .B1(n12480), .B2(n13505), .ZN(
        n9040) );
  INV_X1 U11676 ( .A(n9040), .ZN(n9041) );
  NAND2_X1 U11677 ( .A1(n10747), .A2(P1_DATAO_REG_9__SCAN_IN), .ZN(n9058) );
  NAND2_X1 U11678 ( .A1(n10749), .A2(P2_DATAO_REG_9__SCAN_IN), .ZN(n9045) );
  XNOR2_X1 U11679 ( .A(n9057), .B(n9056), .ZN(n10741) );
  NAND2_X1 U11680 ( .A1(n10741), .A2(n6564), .ZN(n9047) );
  INV_X1 U11681 ( .A(SI_9_), .ZN(n10740) );
  AOI22_X1 U11682 ( .A1(n9198), .A2(n10740), .B1(n9197), .B2(n12061), .ZN(
        n9046) );
  NAND2_X1 U11683 ( .A1(n9047), .A2(n9046), .ZN(n13887) );
  INV_X1 U11684 ( .A(n13887), .ZN(n12112) );
  NAND2_X1 U11685 ( .A1(n13285), .A2(P3_REG0_REG_9__SCAN_IN), .ZN(n9054) );
  OR2_X1 U11686 ( .A1(n9372), .A2(n12050), .ZN(n9053) );
  NAND2_X1 U11687 ( .A1(n9049), .A2(P3_REG3_REG_9__SCAN_IN), .ZN(n9050) );
  AND2_X1 U11688 ( .A1(n9065), .A2(n9050), .ZN(n12111) );
  OR2_X1 U11689 ( .A1(n9126), .A2(n12111), .ZN(n9052) );
  OR2_X1 U11690 ( .A1(n9311), .A2(n12117), .ZN(n9051) );
  XNOR2_X1 U11691 ( .A(n12112), .B(n13504), .ZN(n13381) );
  NAND2_X1 U11692 ( .A1(n12112), .A2(n13504), .ZN(n9055) );
  NAND2_X1 U11693 ( .A1(n11038), .A2(P1_DATAO_REG_10__SCAN_IN), .ZN(n9072) );
  NAND2_X1 U11694 ( .A1(n11041), .A2(P2_DATAO_REG_10__SCAN_IN), .ZN(n9059) );
  OR2_X1 U11695 ( .A1(n9061), .A2(n9060), .ZN(n9062) );
  NAND2_X1 U11696 ( .A1(n9073), .A2(n9062), .ZN(n10669) );
  NAND2_X1 U11697 ( .A1(n10669), .A2(n6564), .ZN(n9064) );
  INV_X1 U11698 ( .A(SI_10_), .ZN(n10670) );
  AOI22_X1 U11699 ( .A1(n9198), .A2(n10670), .B1(n9197), .B2(n10671), .ZN(
        n9063) );
  NAND2_X1 U11700 ( .A1(n9064), .A2(n9063), .ZN(n12735) );
  NAND2_X1 U11701 ( .A1(n6567), .A2(P3_REG0_REG_10__SCAN_IN), .ZN(n9070) );
  OR2_X1 U11702 ( .A1(n9372), .A2(n12733), .ZN(n9069) );
  NAND2_X1 U11703 ( .A1(n9065), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n9066) );
  AND2_X1 U11704 ( .A1(n9092), .A2(n9066), .ZN(n12489) );
  OR2_X1 U11705 ( .A1(n9126), .A2(n12489), .ZN(n9068) );
  OR2_X1 U11706 ( .A1(n9311), .A2(n12624), .ZN(n9067) );
  NAND4_X1 U11707 ( .A1(n9070), .A2(n9069), .A3(n9068), .A4(n9067), .ZN(n13503) );
  OR2_X1 U11708 ( .A1(n12735), .A2(n13503), .ZN(n13388) );
  INV_X1 U11709 ( .A(n9407), .ZN(n13387) );
  NAND2_X1 U11710 ( .A1(n13388), .A2(n13387), .ZN(n12499) );
  INV_X1 U11711 ( .A(n13503), .ZN(n12258) );
  OR2_X1 U11712 ( .A1(n12735), .A2(n12258), .ZN(n9071) );
  NAND2_X1 U11713 ( .A1(n12498), .A2(n9071), .ZN(n12400) );
  NAND2_X1 U11714 ( .A1(n11058), .A2(P2_DATAO_REG_11__SCAN_IN), .ZN(n9074) );
  NAND2_X1 U11715 ( .A1(n9088), .A2(n9074), .ZN(n9076) );
  NAND2_X1 U11716 ( .A1(n11061), .A2(P1_DATAO_REG_11__SCAN_IN), .ZN(n9075) );
  XNOR2_X1 U11717 ( .A(n11259), .B(P2_DATAO_REG_12__SCAN_IN), .ZN(n9103) );
  XNOR2_X1 U11718 ( .A(n9105), .B(n9103), .ZN(n10742) );
  NAND2_X1 U11719 ( .A1(n10742), .A2(n6564), .ZN(n9079) );
  OAI22_X1 U11720 ( .A1(n6569), .A2(n10744), .B1(n13515), .B2(n9367), .ZN(
        n9077) );
  INV_X1 U11721 ( .A(n9077), .ZN(n9078) );
  NAND2_X1 U11722 ( .A1(n9357), .A2(P3_REG1_REG_12__SCAN_IN), .ZN(n9086) );
  INV_X1 U11723 ( .A(P3_REG0_REG_12__SCAN_IN), .ZN(n9080) );
  OR2_X1 U11724 ( .A1(n9007), .A2(n9080), .ZN(n9085) );
  NAND2_X1 U11725 ( .A1(n9094), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n9082) );
  AND2_X1 U11726 ( .A1(n9112), .A2(n9082), .ZN(n12883) );
  OR2_X1 U11727 ( .A1(n9126), .A2(n12883), .ZN(n9084) );
  INV_X1 U11728 ( .A(P3_REG2_REG_12__SCAN_IN), .ZN(n12694) );
  OR2_X1 U11729 ( .A1(n9311), .A2(n12694), .ZN(n9083) );
  OR2_X1 U11730 ( .A1(n12886), .A2(n12934), .ZN(n13395) );
  NAND2_X1 U11731 ( .A1(n12886), .A2(n12934), .ZN(n13396) );
  XNOR2_X1 U11732 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(P2_DATAO_REG_11__SCAN_IN), 
        .ZN(n9087) );
  XNOR2_X1 U11733 ( .A(n9088), .B(n9087), .ZN(n10682) );
  NAND2_X1 U11734 ( .A1(n10682), .A2(n6564), .ZN(n9090) );
  AOI22_X1 U11735 ( .A1(n9198), .A2(n10683), .B1(n9197), .B2(n12601), .ZN(
        n9089) );
  NAND2_X1 U11736 ( .A1(n9090), .A2(n9089), .ZN(n12859) );
  NAND2_X1 U11737 ( .A1(n9357), .A2(P3_REG1_REG_11__SCAN_IN), .ZN(n9098) );
  INV_X1 U11738 ( .A(P3_REG0_REG_11__SCAN_IN), .ZN(n9091) );
  OR2_X1 U11739 ( .A1(n9007), .A2(n9091), .ZN(n9097) );
  NAND2_X1 U11740 ( .A1(n9092), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n9093) );
  AND2_X1 U11741 ( .A1(n9094), .A2(n9093), .ZN(n12437) );
  OR2_X1 U11742 ( .A1(n9126), .A2(n12437), .ZN(n9096) );
  INV_X1 U11743 ( .A(P3_REG2_REG_11__SCAN_IN), .ZN(n12439) );
  OR2_X1 U11744 ( .A1(n9311), .A2(n12439), .ZN(n9095) );
  NAND4_X1 U11745 ( .A1(n9098), .A2(n9097), .A3(n9096), .A4(n9095), .ZN(n13502) );
  INV_X1 U11746 ( .A(n13502), .ZN(n12857) );
  NAND2_X1 U11747 ( .A1(n12859), .A2(n12857), .ZN(n12448) );
  NAND2_X1 U11748 ( .A1(n12400), .A2(n7976), .ZN(n9102) );
  NAND2_X1 U11749 ( .A1(n12859), .A2(n13502), .ZN(n13392) );
  INV_X1 U11750 ( .A(n12448), .ZN(n9099) );
  NOR2_X1 U11751 ( .A1(n7550), .A2(n9099), .ZN(n9100) );
  INV_X1 U11752 ( .A(n12934), .ZN(n13501) );
  AOI22_X1 U11753 ( .A1(n13323), .A2(n9100), .B1(n13501), .B2(n12886), .ZN(
        n9101) );
  NAND2_X1 U11754 ( .A1(n9102), .A2(n9101), .ZN(n12701) );
  INV_X1 U11755 ( .A(n9103), .ZN(n9104) );
  NAND2_X1 U11756 ( .A1(n9106), .A2(P1_DATAO_REG_12__SCAN_IN), .ZN(n9107) );
  XNOR2_X1 U11757 ( .A(n9119), .B(P1_DATAO_REG_13__SCAN_IN), .ZN(n11055) );
  NAND2_X1 U11758 ( .A1(n11055), .A2(n6564), .ZN(n9109) );
  AOI22_X1 U11759 ( .A1(n9197), .A2(n13543), .B1(n9198), .B2(n11056), .ZN(
        n9108) );
  NAND2_X1 U11760 ( .A1(n9357), .A2(P3_REG1_REG_13__SCAN_IN), .ZN(n9117) );
  INV_X1 U11761 ( .A(P3_REG0_REG_13__SCAN_IN), .ZN(n12704) );
  OR2_X1 U11762 ( .A1(n9007), .A2(n12704), .ZN(n9116) );
  NAND2_X1 U11763 ( .A1(n9112), .A2(P3_REG3_REG_13__SCAN_IN), .ZN(n9113) );
  AND2_X1 U11764 ( .A1(n9127), .A2(n9113), .ZN(n13227) );
  OR2_X1 U11765 ( .A1(n9126), .A2(n13227), .ZN(n9115) );
  OR2_X1 U11766 ( .A1(n9311), .A2(n13532), .ZN(n9114) );
  NAND4_X1 U11767 ( .A1(n9117), .A2(n9116), .A3(n9115), .A4(n9114), .ZN(n13500) );
  OR2_X1 U11768 ( .A1(n13223), .A2(n13500), .ZN(n13401) );
  AND2_X1 U11769 ( .A1(n13223), .A2(n13500), .ZN(n9410) );
  INV_X1 U11770 ( .A(n9410), .ZN(n13400) );
  NAND2_X1 U11771 ( .A1(n13401), .A2(n13400), .ZN(n12700) );
  INV_X1 U11772 ( .A(n13500), .ZN(n12937) );
  OR2_X1 U11773 ( .A1(n13223), .A2(n12937), .ZN(n9118) );
  NAND2_X1 U11774 ( .A1(n9119), .A2(P1_DATAO_REG_13__SCAN_IN), .ZN(n9121) );
  NAND2_X1 U11775 ( .A1(n9139), .A2(n11383), .ZN(n9120) );
  NAND2_X1 U11776 ( .A1(n9121), .A2(n9120), .ZN(n9123) );
  XNOR2_X1 U11777 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(P2_DATAO_REG_14__SCAN_IN), 
        .ZN(n9122) );
  XNOR2_X1 U11778 ( .A(n9123), .B(n9122), .ZN(n11127) );
  NAND2_X1 U11779 ( .A1(n11127), .A2(n6564), .ZN(n9125) );
  AOI22_X1 U11780 ( .A1(n11129), .A2(n9197), .B1(n9198), .B2(n11128), .ZN(
        n9124) );
  NAND2_X1 U11781 ( .A1(n9127), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n9128) );
  NAND2_X1 U11782 ( .A1(n9147), .A2(n9128), .ZN(n13156) );
  NAND2_X1 U11783 ( .A1(n9355), .A2(n13156), .ZN(n9134) );
  INV_X1 U11784 ( .A(P3_REG1_REG_14__SCAN_IN), .ZN(n9129) );
  OR2_X1 U11785 ( .A1(n7094), .A2(n9129), .ZN(n9133) );
  INV_X1 U11786 ( .A(P3_REG0_REG_14__SCAN_IN), .ZN(n12770) );
  OR2_X1 U11787 ( .A1(n9007), .A2(n12770), .ZN(n9132) );
  OR2_X1 U11788 ( .A1(n9311), .A2(n9130), .ZN(n9131) );
  NAND2_X1 U11789 ( .A1(n13404), .A2(n13816), .ZN(n9135) );
  NAND2_X1 U11790 ( .A1(n11592), .A2(P2_DATAO_REG_14__SCAN_IN), .ZN(n9140) );
  NAND2_X1 U11791 ( .A1(n11381), .A2(P2_DATAO_REG_13__SCAN_IN), .ZN(n9137) );
  AND2_X1 U11792 ( .A1(n11383), .A2(P1_DATAO_REG_13__SCAN_IN), .ZN(n9141) );
  AOI22_X1 U11793 ( .A1(n9141), .A2(n9140), .B1(P1_DATAO_REG_14__SCAN_IN), 
        .B2(n11590), .ZN(n9142) );
  XNOR2_X1 U11794 ( .A(n11669), .B(P1_DATAO_REG_15__SCAN_IN), .ZN(n9154) );
  XNOR2_X1 U11795 ( .A(n9156), .B(n9154), .ZN(n11123) );
  NAND2_X1 U11796 ( .A1(n11123), .A2(n6564), .ZN(n9144) );
  AOI22_X1 U11797 ( .A1(n13582), .A2(n9197), .B1(SI_15_), .B2(n9198), .ZN(
        n9143) );
  INV_X1 U11798 ( .A(P3_REG3_REG_15__SCAN_IN), .ZN(n9145) );
  NAND2_X1 U11799 ( .A1(n9147), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n9148) );
  NAND2_X1 U11800 ( .A1(n9162), .A2(n9148), .ZN(n13813) );
  NAND2_X1 U11801 ( .A1(n13813), .A2(n9355), .ZN(n9152) );
  NAND2_X1 U11802 ( .A1(n9357), .A2(P3_REG1_REG_15__SCAN_IN), .ZN(n9151) );
  INV_X1 U11803 ( .A(P3_REG0_REG_15__SCAN_IN), .ZN(n10983) );
  OR2_X1 U11804 ( .A1(n9007), .A2(n10983), .ZN(n9150) );
  OR2_X1 U11805 ( .A1(n9311), .A2(n13821), .ZN(n9149) );
  NAND4_X1 U11806 ( .A1(n9152), .A2(n9151), .A3(n9150), .A4(n9149), .ZN(n13498) );
  NAND2_X1 U11807 ( .A1(n13952), .A2(n13498), .ZN(n13801) );
  OR2_X1 U11808 ( .A1(n13952), .A2(n13498), .ZN(n9153) );
  INV_X1 U11809 ( .A(n9154), .ZN(n9155) );
  NAND2_X1 U11810 ( .A1(n11669), .A2(P1_DATAO_REG_15__SCAN_IN), .ZN(n9157) );
  XNOR2_X1 U11811 ( .A(n11587), .B(P2_DATAO_REG_16__SCAN_IN), .ZN(n9167) );
  XNOR2_X1 U11812 ( .A(n9169), .B(n9167), .ZN(n11209) );
  NAND2_X1 U11813 ( .A1(n11209), .A2(n6564), .ZN(n9159) );
  AOI22_X1 U11814 ( .A1(n9198), .A2(SI_16_), .B1(n9197), .B2(n13601), .ZN(
        n9158) );
  NAND2_X1 U11815 ( .A1(n9357), .A2(P3_REG1_REG_16__SCAN_IN), .ZN(n9161) );
  NAND2_X1 U11816 ( .A1(n13285), .A2(P3_REG0_REG_16__SCAN_IN), .ZN(n9160) );
  AND2_X1 U11817 ( .A1(n9161), .A2(n9160), .ZN(n9166) );
  NAND2_X1 U11818 ( .A1(n9162), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n9163) );
  NAND2_X1 U11819 ( .A1(n9175), .A2(n9163), .ZN(n13799) );
  NAND2_X1 U11820 ( .A1(n13799), .A2(n9355), .ZN(n9165) );
  OR2_X1 U11821 ( .A1(n9311), .A2(n13808), .ZN(n9164) );
  OR2_X1 U11822 ( .A1(n13942), .A2(n13818), .ZN(n13410) );
  NAND2_X1 U11823 ( .A1(n13942), .A2(n13818), .ZN(n13415) );
  INV_X1 U11824 ( .A(n13797), .ZN(n13802) );
  INV_X1 U11825 ( .A(n13818), .ZN(n13497) );
  NAND2_X1 U11826 ( .A1(n13942), .A2(n13497), .ZN(n13787) );
  INV_X1 U11827 ( .A(n9167), .ZN(n9168) );
  XNOR2_X1 U11828 ( .A(n11664), .B(P2_DATAO_REG_17__SCAN_IN), .ZN(n9181) );
  XNOR2_X1 U11829 ( .A(n9182), .B(n9181), .ZN(n11346) );
  NAND2_X1 U11830 ( .A1(n11346), .A2(n6564), .ZN(n9173) );
  AOI22_X1 U11831 ( .A1(n9198), .A2(SI_17_), .B1(n9197), .B2(n9171), .ZN(n9172) );
  INV_X1 U11832 ( .A(P3_REG3_REG_17__SCAN_IN), .ZN(n9174) );
  NAND2_X1 U11833 ( .A1(n9175), .A2(P3_REG3_REG_17__SCAN_IN), .ZN(n9176) );
  NAND2_X1 U11834 ( .A1(n9187), .A2(n9176), .ZN(n13785) );
  NAND2_X1 U11835 ( .A1(n13785), .A2(n9355), .ZN(n9179) );
  AOI22_X1 U11836 ( .A1(n9357), .A2(P3_REG1_REG_17__SCAN_IN), .B1(n6567), .B2(
        P3_REG0_REG_17__SCAN_IN), .ZN(n9178) );
  NAND2_X1 U11837 ( .A1(n9368), .A2(P3_REG2_REG_17__SCAN_IN), .ZN(n9177) );
  OR2_X1 U11838 ( .A1(n13939), .A2(n13805), .ZN(n13417) );
  NAND2_X1 U11839 ( .A1(n13939), .A2(n13805), .ZN(n9411) );
  INV_X1 U11840 ( .A(n13805), .ZN(n13774) );
  NAND2_X1 U11841 ( .A1(n13939), .A2(n13774), .ZN(n9180) );
  NAND2_X1 U11842 ( .A1(n9183), .A2(P1_DATAO_REG_17__SCAN_IN), .ZN(n9184) );
  XNOR2_X1 U11843 ( .A(n11972), .B(P2_DATAO_REG_18__SCAN_IN), .ZN(n9193) );
  XNOR2_X1 U11844 ( .A(n9194), .B(n9193), .ZN(n11457) );
  NAND2_X1 U11845 ( .A1(n11457), .A2(n6564), .ZN(n9186) );
  AOI22_X1 U11846 ( .A1(n9198), .A2(SI_18_), .B1(n9197), .B2(n13641), .ZN(
        n9185) );
  NAND2_X1 U11847 ( .A1(n9187), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n9188) );
  NAND2_X1 U11848 ( .A1(n6614), .A2(n9188), .ZN(n13778) );
  NAND2_X1 U11849 ( .A1(n13778), .A2(n9355), .ZN(n9191) );
  AOI22_X1 U11850 ( .A1(n9357), .A2(P3_REG1_REG_18__SCAN_IN), .B1(n13285), 
        .B2(P3_REG0_REG_18__SCAN_IN), .ZN(n9190) );
  NAND2_X1 U11851 ( .A1(n9368), .A2(P3_REG2_REG_18__SCAN_IN), .ZN(n9189) );
  NAND2_X1 U11852 ( .A1(n13868), .A2(n13791), .ZN(n13423) );
  OR2_X1 U11853 ( .A1(n13868), .A2(n13496), .ZN(n9192) );
  NAND2_X1 U11854 ( .A1(n11971), .A2(P1_DATAO_REG_18__SCAN_IN), .ZN(n9195) );
  XNOR2_X1 U11855 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(P2_DATAO_REG_19__SCAN_IN), 
        .ZN(n9211) );
  XNOR2_X1 U11856 ( .A(n9212), .B(n9211), .ZN(n11462) );
  NAND2_X1 U11857 ( .A1(n11462), .A2(n6564), .ZN(n9200) );
  AOI22_X1 U11858 ( .A1(n9198), .A2(n11461), .B1(n9197), .B2(n13306), .ZN(
        n9199) );
  INV_X1 U11859 ( .A(P3_REG3_REG_19__SCAN_IN), .ZN(n9201) );
  NAND2_X1 U11860 ( .A1(n6614), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n9203) );
  NAND2_X1 U11861 ( .A1(n9216), .A2(n9203), .ZN(n13757) );
  NAND2_X1 U11862 ( .A1(n13757), .A2(n9355), .ZN(n9208) );
  INV_X1 U11863 ( .A(P3_REG1_REG_19__SCAN_IN), .ZN(n13864) );
  NAND2_X1 U11864 ( .A1(n9368), .A2(P3_REG2_REG_19__SCAN_IN), .ZN(n9205) );
  NAND2_X1 U11865 ( .A1(n6567), .A2(P3_REG0_REG_19__SCAN_IN), .ZN(n9204) );
  OAI211_X1 U11866 ( .C1(n9372), .C2(n13864), .A(n9205), .B(n9204), .ZN(n9206)
         );
  INV_X1 U11867 ( .A(n9206), .ZN(n9207) );
  INV_X1 U11868 ( .A(n13425), .ZN(n13427) );
  NAND2_X1 U11869 ( .A1(n13172), .A2(n13775), .ZN(n13428) );
  OR2_X1 U11870 ( .A1(n13172), .A2(n13748), .ZN(n9210) );
  INV_X1 U11871 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n12142) );
  NAND2_X1 U11872 ( .A1(n12142), .A2(P1_DATAO_REG_19__SCAN_IN), .ZN(n9213) );
  XNOR2_X1 U11873 ( .A(n9239), .B(P1_DATAO_REG_20__SCAN_IN), .ZN(n9224) );
  XNOR2_X1 U11874 ( .A(n9224), .B(n12096), .ZN(n11749) );
  NAND2_X1 U11875 ( .A1(n11749), .A2(n6564), .ZN(n9215) );
  OR2_X1 U11876 ( .A1(n6568), .A2(n11751), .ZN(n9214) );
  NAND2_X1 U11877 ( .A1(n9216), .A2(P3_REG3_REG_20__SCAN_IN), .ZN(n9217) );
  NAND2_X1 U11878 ( .A1(n9231), .A2(n9217), .ZN(n13743) );
  NAND2_X1 U11879 ( .A1(n13743), .A2(n9355), .ZN(n9222) );
  INV_X1 U11880 ( .A(P3_REG1_REG_20__SCAN_IN), .ZN(n13861) );
  NAND2_X1 U11881 ( .A1(n9368), .A2(P3_REG2_REG_20__SCAN_IN), .ZN(n9219) );
  NAND2_X1 U11882 ( .A1(n13285), .A2(P3_REG0_REG_20__SCAN_IN), .ZN(n9218) );
  OAI211_X1 U11883 ( .C1(n7094), .C2(n13861), .A(n9219), .B(n9218), .ZN(n9220)
         );
  INV_X1 U11884 ( .A(n9220), .ZN(n9221) );
  NAND2_X1 U11885 ( .A1(n13922), .A2(n13761), .ZN(n13432) );
  INV_X1 U11886 ( .A(n13745), .ZN(n13329) );
  NAND2_X1 U11887 ( .A1(n13922), .A2(n13495), .ZN(n9223) );
  NAND2_X1 U11888 ( .A1(n9239), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n9225) );
  NAND2_X1 U11889 ( .A1(n9226), .A2(n9225), .ZN(n9228) );
  INV_X1 U11890 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n12144) );
  XNOR2_X1 U11891 ( .A(n12144), .B(P2_DATAO_REG_21__SCAN_IN), .ZN(n9227) );
  XNOR2_X1 U11892 ( .A(n9228), .B(n9227), .ZN(n13148) );
  NAND2_X1 U11893 ( .A1(n13148), .A2(n6564), .ZN(n9230) );
  INV_X1 U11894 ( .A(SI_21_), .ZN(n13149) );
  OR2_X1 U11895 ( .A1(n6569), .A2(n13149), .ZN(n9229) );
  INV_X1 U11896 ( .A(P3_REG3_REG_21__SCAN_IN), .ZN(n10861) );
  NAND2_X1 U11897 ( .A1(n9231), .A2(P3_REG3_REG_21__SCAN_IN), .ZN(n9232) );
  NAND2_X1 U11898 ( .A1(n9248), .A2(n9232), .ZN(n13735) );
  INV_X1 U11899 ( .A(P3_REG1_REG_21__SCAN_IN), .ZN(n13858) );
  NAND2_X1 U11900 ( .A1(n9368), .A2(P3_REG2_REG_21__SCAN_IN), .ZN(n9234) );
  NAND2_X1 U11901 ( .A1(n13285), .A2(P3_REG0_REG_21__SCAN_IN), .ZN(n9233) );
  OAI211_X1 U11902 ( .C1(n7094), .C2(n13858), .A(n9234), .B(n9233), .ZN(n9235)
         );
  NOR2_X1 U11903 ( .A1(n13734), .A2(n13749), .ZN(n9412) );
  INV_X1 U11904 ( .A(n9412), .ZN(n13435) );
  NAND2_X1 U11905 ( .A1(n13734), .A2(n13749), .ZN(n13436) );
  INV_X1 U11906 ( .A(n13749), .ZN(n13721) );
  OR2_X1 U11907 ( .A1(n13734), .A2(n13721), .ZN(n9237) );
  AOI22_X1 U11908 ( .A1(P2_DATAO_REG_21__SCAN_IN), .A2(n12144), .B1(n12184), 
        .B2(P2_DATAO_REG_20__SCAN_IN), .ZN(n9238) );
  OAI21_X1 U11909 ( .B1(n12184), .B2(P2_DATAO_REG_20__SCAN_IN), .A(
        P2_DATAO_REG_21__SCAN_IN), .ZN(n9241) );
  NOR2_X1 U11910 ( .A1(P2_DATAO_REG_20__SCAN_IN), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n9240) );
  AOI22_X1 U11911 ( .A1(n9241), .A2(P1_DATAO_REG_21__SCAN_IN), .B1(n9240), 
        .B2(P1_DATAO_REG_20__SCAN_IN), .ZN(n9242) );
  NAND2_X1 U11912 ( .A1(n12356), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n9259) );
  NAND2_X1 U11913 ( .A1(n9243), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n9244) );
  NAND2_X1 U11914 ( .A1(n9259), .A2(n9244), .ZN(n9257) );
  XNOR2_X1 U11915 ( .A(n9258), .B(n9257), .ZN(n11710) );
  NAND2_X1 U11916 ( .A1(n11710), .A2(n6564), .ZN(n9247) );
  OR2_X1 U11917 ( .A1(n6568), .A2(n9245), .ZN(n9246) );
  NAND2_X1 U11918 ( .A1(n9248), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n9249) );
  NAND2_X1 U11919 ( .A1(n9267), .A2(n9249), .ZN(n13718) );
  NAND2_X1 U11920 ( .A1(n13718), .A2(n9355), .ZN(n9254) );
  INV_X1 U11921 ( .A(P3_REG1_REG_22__SCAN_IN), .ZN(n13853) );
  NAND2_X1 U11922 ( .A1(n13285), .A2(P3_REG0_REG_22__SCAN_IN), .ZN(n9251) );
  NAND2_X1 U11923 ( .A1(n9368), .A2(P3_REG2_REG_22__SCAN_IN), .ZN(n9250) );
  OAI211_X1 U11924 ( .C1(n13853), .C2(n9372), .A(n9251), .B(n9250), .ZN(n9252)
         );
  INV_X1 U11925 ( .A(n9252), .ZN(n9253) );
  NOR2_X1 U11926 ( .A1(n13911), .A2(n13705), .ZN(n9256) );
  NAND2_X1 U11927 ( .A1(n13911), .A2(n13705), .ZN(n9255) );
  INV_X1 U11928 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n9260) );
  NAND2_X1 U11929 ( .A1(n9260), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n9276) );
  INV_X1 U11930 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n10934) );
  NAND2_X1 U11931 ( .A1(n10934), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n9261) );
  AND2_X1 U11932 ( .A1(n9276), .A2(n9261), .ZN(n9262) );
  OR2_X1 U11933 ( .A1(n9263), .A2(n9262), .ZN(n9264) );
  NAND2_X1 U11934 ( .A1(n9277), .A2(n9264), .ZN(n11938) );
  NAND2_X1 U11935 ( .A1(n11938), .A2(n6564), .ZN(n9266) );
  OR2_X1 U11936 ( .A1(n6569), .A2(n11940), .ZN(n9265) );
  NAND2_X1 U11937 ( .A1(n9267), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n9268) );
  NAND2_X1 U11938 ( .A1(n9279), .A2(n9268), .ZN(n13712) );
  NAND2_X1 U11939 ( .A1(n13712), .A2(n9355), .ZN(n9273) );
  INV_X1 U11940 ( .A(P3_REG1_REG_23__SCAN_IN), .ZN(n13851) );
  NAND2_X1 U11941 ( .A1(n9368), .A2(P3_REG2_REG_23__SCAN_IN), .ZN(n9270) );
  INV_X1 U11942 ( .A(P3_REG0_REG_23__SCAN_IN), .ZN(n13906) );
  OR2_X1 U11943 ( .A1(n9007), .A2(n13906), .ZN(n9269) );
  OAI211_X1 U11944 ( .C1(n9372), .C2(n13851), .A(n9270), .B(n9269), .ZN(n9271)
         );
  INV_X1 U11945 ( .A(n9271), .ZN(n9272) );
  XNOR2_X1 U11946 ( .A(n13850), .B(n13722), .ZN(n13704) );
  INV_X1 U11947 ( .A(n13704), .ZN(n13710) );
  NAND2_X1 U11948 ( .A1(n13850), .A2(n13722), .ZN(n9274) );
  XNOR2_X1 U11949 ( .A(n9288), .B(P2_DATAO_REG_24__SCAN_IN), .ZN(n12983) );
  OR2_X1 U11950 ( .A1(n6568), .A2(n12984), .ZN(n9278) );
  INV_X1 U11951 ( .A(n9295), .ZN(n9296) );
  NAND2_X1 U11952 ( .A1(n9279), .A2(P3_REG3_REG_24__SCAN_IN), .ZN(n9280) );
  NAND2_X1 U11953 ( .A1(n9296), .A2(n9280), .ZN(n13695) );
  NAND2_X1 U11954 ( .A1(n13695), .A2(n9355), .ZN(n9285) );
  INV_X1 U11955 ( .A(P3_REG1_REG_24__SCAN_IN), .ZN(n13844) );
  NAND2_X1 U11956 ( .A1(n6567), .A2(P3_REG0_REG_24__SCAN_IN), .ZN(n9282) );
  INV_X1 U11957 ( .A(P3_REG2_REG_24__SCAN_IN), .ZN(n13699) );
  OR2_X1 U11958 ( .A1(n9311), .A2(n13699), .ZN(n9281) );
  OAI211_X1 U11959 ( .C1(n9372), .C2(n13844), .A(n9282), .B(n9281), .ZN(n9283)
         );
  INV_X1 U11960 ( .A(n9283), .ZN(n9284) );
  AND2_X1 U11961 ( .A1(n13899), .A2(n7128), .ZN(n9287) );
  INV_X1 U11962 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n12791) );
  XNOR2_X1 U11963 ( .A(n12791), .B(P2_DATAO_REG_25__SCAN_IN), .ZN(n9291) );
  NAND2_X1 U11964 ( .A1(n12293), .A2(n6564), .ZN(n9293) );
  INV_X1 U11965 ( .A(SI_25_), .ZN(n12294) );
  OR2_X1 U11966 ( .A1(n6568), .A2(n12294), .ZN(n9292) );
  INV_X1 U11967 ( .A(P3_REG3_REG_25__SCAN_IN), .ZN(n9294) );
  NAND2_X1 U11968 ( .A1(n9296), .A2(P3_REG3_REG_25__SCAN_IN), .ZN(n9297) );
  NAND2_X1 U11969 ( .A1(n9308), .A2(n9297), .ZN(n13688) );
  NAND2_X1 U11970 ( .A1(n13688), .A2(n9355), .ZN(n9302) );
  INV_X1 U11971 ( .A(P3_REG1_REG_25__SCAN_IN), .ZN(n13842) );
  NAND2_X1 U11972 ( .A1(n9368), .A2(P3_REG2_REG_25__SCAN_IN), .ZN(n9299) );
  NAND2_X1 U11973 ( .A1(n13285), .A2(P3_REG0_REG_25__SCAN_IN), .ZN(n9298) );
  OAI211_X1 U11974 ( .C1(n9372), .C2(n13842), .A(n9299), .B(n9298), .ZN(n9300)
         );
  INV_X1 U11975 ( .A(n9300), .ZN(n9301) );
  INV_X1 U11976 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n12792) );
  NAND2_X1 U11977 ( .A1(n12791), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n9304) );
  XNOR2_X1 U11978 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(P2_DATAO_REG_26__SCAN_IN), 
        .ZN(n9305) );
  XNOR2_X1 U11979 ( .A(n9321), .B(n9305), .ZN(n12506) );
  NAND2_X1 U11980 ( .A1(n12506), .A2(n6564), .ZN(n9307) );
  OR2_X1 U11981 ( .A1(n6568), .A2(n12507), .ZN(n9306) );
  NAND2_X1 U11982 ( .A1(n9308), .A2(P3_REG3_REG_26__SCAN_IN), .ZN(n9309) );
  NAND2_X1 U11983 ( .A1(n9328), .A2(n9309), .ZN(n13670) );
  NAND2_X1 U11984 ( .A1(n13670), .A2(n9355), .ZN(n9316) );
  INV_X1 U11985 ( .A(P3_REG1_REG_26__SCAN_IN), .ZN(n10914) );
  NAND2_X1 U11986 ( .A1(n13285), .A2(P3_REG0_REG_26__SCAN_IN), .ZN(n9313) );
  INV_X1 U11987 ( .A(P3_REG2_REG_26__SCAN_IN), .ZN(n9310) );
  OR2_X1 U11988 ( .A1(n9311), .A2(n9310), .ZN(n9312) );
  OAI211_X1 U11989 ( .C1(n10914), .C2(n7094), .A(n9313), .B(n9312), .ZN(n9314)
         );
  INV_X1 U11990 ( .A(n9314), .ZN(n9315) );
  OR2_X1 U11991 ( .A1(n13836), .A2(n13494), .ZN(n9317) );
  NAND2_X1 U11992 ( .A1(n13836), .A2(n13494), .ZN(n9318) );
  INV_X1 U11993 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n15701) );
  NOR2_X1 U11994 ( .A1(n15701), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n9320) );
  NAND2_X1 U11995 ( .A1(n15701), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n9322) );
  INV_X1 U11996 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n14913) );
  XNOR2_X1 U11997 ( .A(n14913), .B(P2_DATAO_REG_27__SCAN_IN), .ZN(n9323) );
  XNOR2_X1 U11998 ( .A(n9338), .B(n9323), .ZN(n13108) );
  NAND2_X1 U11999 ( .A1(n13108), .A2(n6564), .ZN(n9325) );
  INV_X1 U12000 ( .A(SI_27_), .ZN(n13109) );
  OR2_X1 U12001 ( .A1(n6569), .A2(n13109), .ZN(n9324) );
  INV_X1 U12002 ( .A(n9328), .ZN(n9327) );
  INV_X1 U12003 ( .A(P3_REG3_REG_27__SCAN_IN), .ZN(n9326) );
  NAND2_X1 U12004 ( .A1(n9328), .A2(P3_REG3_REG_27__SCAN_IN), .ZN(n9329) );
  NAND2_X1 U12005 ( .A1(n9342), .A2(n9329), .ZN(n13658) );
  NAND2_X1 U12006 ( .A1(n13658), .A2(n9355), .ZN(n9334) );
  INV_X1 U12007 ( .A(P3_REG1_REG_27__SCAN_IN), .ZN(n13834) );
  NAND2_X1 U12008 ( .A1(n13285), .A2(P3_REG0_REG_27__SCAN_IN), .ZN(n9331) );
  NAND2_X1 U12009 ( .A1(n9368), .A2(P3_REG2_REG_27__SCAN_IN), .ZN(n9330) );
  OAI211_X1 U12010 ( .C1(n9372), .C2(n13834), .A(n9331), .B(n9330), .ZN(n9332)
         );
  INV_X1 U12011 ( .A(n9332), .ZN(n9333) );
  OR2_X1 U12012 ( .A1(n13460), .A2(n13666), .ZN(n9336) );
  INV_X1 U12013 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n15697) );
  AND2_X1 U12014 ( .A1(n15697), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n9337) );
  XNOR2_X1 U12015 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(P2_DATAO_REG_28__SCAN_IN), 
        .ZN(n9339) );
  XNOR2_X1 U12016 ( .A(n9350), .B(n9339), .ZN(n13969) );
  NAND2_X1 U12017 ( .A1(n13969), .A2(n6564), .ZN(n9341) );
  OR2_X1 U12018 ( .A1(n6568), .A2(n13971), .ZN(n9340) );
  NAND2_X1 U12019 ( .A1(n9342), .A2(P3_REG3_REG_28__SCAN_IN), .ZN(n9343) );
  NAND2_X1 U12020 ( .A1(n9423), .A2(n9343), .ZN(n13652) );
  INV_X1 U12021 ( .A(P3_REG1_REG_28__SCAN_IN), .ZN(n13830) );
  NAND2_X1 U12022 ( .A1(n6567), .A2(P3_REG0_REG_28__SCAN_IN), .ZN(n9345) );
  NAND2_X1 U12023 ( .A1(n9368), .A2(P3_REG2_REG_28__SCAN_IN), .ZN(n9344) );
  OAI211_X1 U12024 ( .C1(n13830), .C2(n7094), .A(n9345), .B(n9344), .ZN(n9346)
         );
  NAND2_X1 U12025 ( .A1(n13145), .A2(n12979), .ZN(n9413) );
  INV_X1 U12026 ( .A(n12979), .ZN(n13493) );
  NAND2_X1 U12027 ( .A1(n13145), .A2(n13493), .ZN(n9347) );
  AND2_X1 U12028 ( .A1(n14910), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n9349) );
  NAND2_X1 U12029 ( .A1(n13106), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n9348) );
  XNOR2_X1 U12030 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(P2_DATAO_REG_29__SCAN_IN), 
        .ZN(n9351) );
  INV_X1 U12031 ( .A(SI_29_), .ZN(n13131) );
  OR2_X1 U12032 ( .A1(n6569), .A2(n13131), .ZN(n9354) );
  INV_X1 U12033 ( .A(P3_REG0_REG_29__SCAN_IN), .ZN(n10905) );
  NAND2_X1 U12034 ( .A1(n9357), .A2(P3_REG1_REG_29__SCAN_IN), .ZN(n9359) );
  NAND2_X1 U12035 ( .A1(n9368), .A2(P3_REG2_REG_29__SCAN_IN), .ZN(n9358) );
  OAI211_X1 U12036 ( .C1(n9007), .C2(n10905), .A(n9359), .B(n9358), .ZN(n9360)
         );
  INV_X1 U12037 ( .A(n9360), .ZN(n9361) );
  XNOR2_X1 U12038 ( .A(n9362), .B(n6607), .ZN(n9365) );
  NAND2_X1 U12039 ( .A1(n13487), .A2(n13332), .ZN(n10085) );
  NAND2_X1 U12040 ( .A1(n9363), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9364) );
  NAND2_X1 U12041 ( .A1(n13333), .A2(n10104), .ZN(n13308) );
  NAND2_X1 U12042 ( .A1(n9365), .A2(n16044), .ZN(n9378) );
  AND2_X1 U12043 ( .A1(n9367), .A2(n9366), .ZN(n11440) );
  INV_X1 U12044 ( .A(P3_REG1_REG_30__SCAN_IN), .ZN(n9371) );
  NAND2_X1 U12045 ( .A1(n9368), .A2(P3_REG2_REG_30__SCAN_IN), .ZN(n9370) );
  NAND2_X1 U12046 ( .A1(n13285), .A2(P3_REG0_REG_30__SCAN_IN), .ZN(n9369) );
  OAI211_X1 U12047 ( .C1(n9372), .C2(n9371), .A(n9370), .B(n9369), .ZN(n9373)
         );
  INV_X1 U12048 ( .A(n9373), .ZN(n9374) );
  NAND2_X1 U12049 ( .A1(n13290), .A2(n9374), .ZN(n13491) );
  AND2_X1 U12050 ( .A1(n9375), .A2(P3_B_REG_SCAN_IN), .ZN(n9376) );
  NOR2_X1 U12051 ( .A1(n13817), .A2(n9376), .ZN(n13645) );
  AOI22_X1 U12052 ( .A1(n16049), .A2(n13493), .B1(n13491), .B2(n13645), .ZN(
        n9377) );
  NAND2_X1 U12053 ( .A1(n9378), .A2(n9377), .ZN(n10111) );
  XNOR2_X1 U12054 ( .A(n12986), .B(P3_B_REG_SCAN_IN), .ZN(n9379) );
  NAND2_X1 U12055 ( .A1(n9379), .A2(n12296), .ZN(n9380) );
  NAND2_X1 U12056 ( .A1(n9380), .A2(n9381), .ZN(n9383) );
  INV_X1 U12057 ( .A(n9381), .ZN(n12509) );
  NAND2_X1 U12058 ( .A1(n12986), .A2(n12509), .ZN(n9382) );
  OR2_X1 U12059 ( .A1(n9383), .A2(P3_D_REG_1__SCAN_IN), .ZN(n9385) );
  NAND2_X1 U12060 ( .A1(n12509), .A2(n12296), .ZN(n9384) );
  NAND2_X1 U12061 ( .A1(n9385), .A2(n9384), .ZN(n10106) );
  AND2_X1 U12062 ( .A1(n11430), .A2(n10106), .ZN(n10091) );
  NOR2_X1 U12063 ( .A1(P3_D_REG_7__SCAN_IN), .A2(P3_D_REG_3__SCAN_IN), .ZN(
        n10801) );
  NOR4_X1 U12064 ( .A1(P3_D_REG_4__SCAN_IN), .A2(P3_D_REG_2__SCAN_IN), .A3(
        P3_D_REG_13__SCAN_IN), .A4(P3_D_REG_9__SCAN_IN), .ZN(n9388) );
  NOR4_X1 U12065 ( .A1(P3_D_REG_17__SCAN_IN), .A2(P3_D_REG_22__SCAN_IN), .A3(
        P3_D_REG_25__SCAN_IN), .A4(P3_D_REG_20__SCAN_IN), .ZN(n9387) );
  NOR4_X1 U12066 ( .A1(P3_D_REG_14__SCAN_IN), .A2(P3_D_REG_27__SCAN_IN), .A3(
        P3_D_REG_8__SCAN_IN), .A4(P3_D_REG_10__SCAN_IN), .ZN(n9386) );
  NAND4_X1 U12067 ( .A1(n10801), .A2(n9388), .A3(n9387), .A4(n9386), .ZN(n9394) );
  NOR4_X1 U12068 ( .A1(P3_D_REG_29__SCAN_IN), .A2(P3_D_REG_21__SCAN_IN), .A3(
        P3_D_REG_12__SCAN_IN), .A4(P3_D_REG_11__SCAN_IN), .ZN(n9392) );
  NOR4_X1 U12069 ( .A1(P3_D_REG_19__SCAN_IN), .A2(P3_D_REG_18__SCAN_IN), .A3(
        P3_D_REG_31__SCAN_IN), .A4(P3_D_REG_24__SCAN_IN), .ZN(n9391) );
  NOR4_X1 U12070 ( .A1(P3_D_REG_28__SCAN_IN), .A2(P3_D_REG_23__SCAN_IN), .A3(
        P3_D_REG_6__SCAN_IN), .A4(P3_D_REG_5__SCAN_IN), .ZN(n9390) );
  NOR4_X1 U12071 ( .A1(P3_D_REG_26__SCAN_IN), .A2(P3_D_REG_30__SCAN_IN), .A3(
        P3_D_REG_16__SCAN_IN), .A4(P3_D_REG_15__SCAN_IN), .ZN(n9389) );
  NAND4_X1 U12072 ( .A1(n9392), .A2(n9391), .A3(n9390), .A4(n9389), .ZN(n9393)
         );
  NOR2_X1 U12073 ( .A1(n9394), .A2(n9393), .ZN(n9395) );
  NOR2_X1 U12074 ( .A1(n9383), .A2(n9395), .ZN(n10087) );
  NAND2_X1 U12075 ( .A1(n11750), .A2(n13306), .ZN(n13481) );
  INV_X1 U12076 ( .A(n13481), .ZN(n10086) );
  OR3_X1 U12077 ( .A1(n11708), .A2(n13332), .A3(n11750), .ZN(n9419) );
  NAND2_X1 U12078 ( .A1(n13450), .A2(n9419), .ZN(n9397) );
  NAND2_X1 U12079 ( .A1(n9397), .A2(n13958), .ZN(n9398) );
  OAI21_X1 U12080 ( .B1(n10108), .B2(n13958), .A(n9398), .ZN(n9399) );
  INV_X1 U12081 ( .A(n9399), .ZN(n9400) );
  NAND2_X1 U12082 ( .A1(n10109), .A2(n9400), .ZN(n9422) );
  INV_X2 U12083 ( .A(n16066), .ZN(n9401) );
  NAND2_X1 U12084 ( .A1(n10111), .A2(n9401), .ZN(n9430) );
  NAND2_X1 U12085 ( .A1(n13339), .A2(n13342), .ZN(n11434) );
  NAND2_X1 U12086 ( .A1(n11434), .A2(n9402), .ZN(n16026) );
  AND2_X1 U12087 ( .A1(n13358), .A2(n13351), .ZN(n9405) );
  OAI21_X1 U12088 ( .B1(n9403), .B2(n13354), .A(n13361), .ZN(n9404) );
  NAND2_X1 U12089 ( .A1(n13504), .A2(n13887), .ZN(n13383) );
  NOR2_X1 U12090 ( .A1(n13504), .A2(n13887), .ZN(n13384) );
  INV_X1 U12091 ( .A(n13396), .ZN(n9408) );
  AOI21_X2 U12092 ( .B1(n12447), .B2(n9409), .A(n9408), .ZN(n12698) );
  AOI21_X2 U12093 ( .B1(n12698), .B2(n13401), .A(n9410), .ZN(n12765) );
  NOR2_X1 U12094 ( .A1(n13404), .A2(n13499), .ZN(n13405) );
  INV_X1 U12095 ( .A(n13498), .ZN(n13804) );
  NAND2_X1 U12096 ( .A1(n13952), .A2(n13804), .ZN(n13414) );
  INV_X1 U12097 ( .A(n9411), .ZN(n13421) );
  AND2_X1 U12098 ( .A1(n13428), .A2(n13755), .ZN(n13420) );
  NAND2_X1 U12099 ( .A1(n13741), .A2(n13431), .ZN(n13727) );
  OR2_X1 U12100 ( .A1(n13850), .A2(n13444), .ZN(n13675) );
  NAND2_X1 U12101 ( .A1(n13899), .A2(n13683), .ZN(n13676) );
  NAND2_X1 U12102 ( .A1(n13836), .A2(n13684), .ZN(n13310) );
  INV_X1 U12103 ( .A(n13666), .ZN(n13461) );
  NAND2_X1 U12104 ( .A1(n13460), .A2(n13461), .ZN(n10574) );
  AND2_X1 U12105 ( .A1(n9413), .A2(n10574), .ZN(n13464) );
  NAND2_X1 U12106 ( .A1(n10575), .A2(n13464), .ZN(n13299) );
  NAND2_X1 U12107 ( .A1(n13299), .A2(n13462), .ZN(n9414) );
  INV_X1 U12108 ( .A(n16057), .ZN(n16038) );
  NAND2_X1 U12109 ( .A1(n13333), .A2(n16038), .ZN(n16039) );
  OAI21_X1 U12110 ( .B1(n11708), .B2(n10104), .A(n13332), .ZN(n9415) );
  NAND2_X1 U12111 ( .A1(n9415), .A2(n11431), .ZN(n9417) );
  OAI21_X1 U12112 ( .B1(n13333), .B2(n10104), .A(n11708), .ZN(n9416) );
  NAND2_X1 U12113 ( .A1(n9417), .A2(n9416), .ZN(n11411) );
  AND2_X1 U12114 ( .A1(n16055), .A2(n10086), .ZN(n9418) );
  NAND2_X1 U12115 ( .A1(n11411), .A2(n9418), .ZN(n9420) );
  NAND2_X1 U12116 ( .A1(n9420), .A2(n9419), .ZN(n16054) );
  INV_X1 U12117 ( .A(n16054), .ZN(n12503) );
  OR2_X1 U12118 ( .A1(n9422), .A2(n16038), .ZN(n12133) );
  NOR2_X2 U12119 ( .A1(n12133), .A2(n16055), .ZN(n13814) );
  NOR2_X1 U12120 ( .A1(n9423), .A2(n12707), .ZN(n13647) );
  AOI21_X1 U12121 ( .B1(n10100), .B2(n13814), .A(n13647), .ZN(n9425) );
  NAND2_X1 U12122 ( .A1(n16066), .A2(P3_REG2_REG_29__SCAN_IN), .ZN(n9424) );
  NAND2_X1 U12123 ( .A1(n9430), .A2(n9429), .ZN(P3_U3204) );
  INV_X1 U12124 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n15052) );
  INV_X1 U12125 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n14961) );
  NAND2_X1 U12126 ( .A1(n9817), .A2(n14961), .ZN(n9436) );
  NAND2_X1 U12127 ( .A1(n9828), .A2(n9436), .ZN(n15394) );
  INV_X1 U12128 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n9445) );
  INV_X1 U12129 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n9447) );
  XNOR2_X2 U12130 ( .A(n9449), .B(n9448), .ZN(n15696) );
  INV_X1 U12131 ( .A(P1_REG2_REG_21__SCAN_IN), .ZN(n15395) );
  NAND2_X1 U12133 ( .A1(n9838), .A2(P1_REG1_REG_21__SCAN_IN), .ZN(n9453) );
  NAND2_X1 U12134 ( .A1(n9947), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n9452) );
  OAI211_X1 U12135 ( .C1(n9960), .C2(n15395), .A(n9453), .B(n9452), .ZN(n9454)
         );
  INV_X1 U12136 ( .A(n9454), .ZN(n9455) );
  NAND2_X1 U12137 ( .A1(n9940), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n9460) );
  INV_X1 U12138 ( .A(n15597), .ZN(n15393) );
  AND2_X2 U12139 ( .A1(n9531), .A2(n10810), .ZN(n9534) );
  INV_X1 U12140 ( .A(n9462), .ZN(n9463) );
  NOR2_X1 U12141 ( .A1(n9463), .A2(P1_IR_REG_15__SCAN_IN), .ZN(n9464) );
  NAND2_X1 U12142 ( .A1(n9751), .A2(n9468), .ZN(n9474) );
  INV_X1 U12143 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n9466) );
  NAND3_X1 U12144 ( .A1(n9469), .A2(n9467), .A3(n9468), .ZN(n9470) );
  OAI21_X2 U12145 ( .B1(n9476), .B2(P1_IR_REG_21__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n9471) );
  NAND2_X1 U12146 ( .A1(n9476), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9473) );
  INV_X1 U12147 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n9472) );
  NAND2_X1 U12148 ( .A1(n9481), .A2(n12140), .ZN(n9945) );
  INV_X1 U12149 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n9475) );
  NAND2_X1 U12150 ( .A1(n9513), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n9484) );
  INV_X1 U12151 ( .A(n15103), .ZN(n9482) );
  INV_X1 U12152 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n15100) );
  INV_X1 U12153 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n9485) );
  OR2_X1 U12154 ( .A1(n9832), .A2(n9485), .ZN(n9490) );
  INV_X1 U12155 ( .A(n6551), .ZN(n9487) );
  NAND2_X1 U12156 ( .A1(n9487), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n9488) );
  INV_X4 U12157 ( .A(n9635), .ZN(n9743) );
  NAND2_X1 U12158 ( .A1(n9506), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n9496) );
  INV_X1 U12159 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n9492) );
  OR2_X1 U12160 ( .A1(n9486), .A2(n9492), .ZN(n9495) );
  INV_X1 U12161 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n12041) );
  INV_X1 U12162 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n10725) );
  OAI21_X1 U12163 ( .B1(n10696), .B2(n10735), .A(n9497), .ZN(n9498) );
  AND2_X1 U12164 ( .A1(n9499), .A2(n9498), .ZN(n15707) );
  INV_X1 U12165 ( .A(n11472), .ZN(n10117) );
  NAND2_X1 U12166 ( .A1(n10028), .A2(n10117), .ZN(n9500) );
  NAND2_X1 U12167 ( .A1(n11476), .A2(n7137), .ZN(n10027) );
  NAND2_X1 U12168 ( .A1(n9500), .A2(n10027), .ZN(n9501) );
  NAND2_X1 U12169 ( .A1(n10123), .A2(n11483), .ZN(n9503) );
  INV_X1 U12170 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n15121) );
  INV_X2 U12171 ( .A(n9506), .ZN(n9832) );
  INV_X1 U12172 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n9507) );
  OR2_X1 U12173 ( .A1(n9832), .A2(n9507), .ZN(n9510) );
  INV_X1 U12174 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n9508) );
  OR2_X1 U12175 ( .A1(n6553), .A2(n9508), .ZN(n9509) );
  INV_X1 U12176 ( .A(n9515), .ZN(n9516) );
  NAND2_X1 U12177 ( .A1(n9516), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9517) );
  XNOR2_X1 U12178 ( .A(n9517), .B(P1_IR_REG_2__SCAN_IN), .ZN(n15124) );
  INV_X1 U12179 ( .A(n15124), .ZN(n9518) );
  NAND3_X1 U12180 ( .A1(n9522), .A2(n9521), .A3(n7826), .ZN(n9539) );
  NAND2_X1 U12181 ( .A1(n10144), .A2(n15834), .ZN(n9523) );
  OR2_X1 U12182 ( .A1(n10144), .A2(n15834), .ZN(n11957) );
  MUX2_X1 U12183 ( .A(n9523), .B(n11957), .S(n9743), .Z(n9538) );
  OR2_X1 U12184 ( .A1(n6550), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n9529) );
  INV_X1 U12185 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n9525) );
  OR2_X1 U12186 ( .A1(n9832), .A2(n9525), .ZN(n9528) );
  INV_X1 U12187 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n11064) );
  OR2_X1 U12188 ( .A1(n6553), .A2(n11064), .ZN(n9527) );
  INV_X1 U12189 ( .A(n9531), .ZN(n9532) );
  NAND2_X1 U12190 ( .A1(n9532), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9533) );
  MUX2_X1 U12191 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9533), .S(
        P1_IR_REG_3__SCAN_IN), .Z(n9535) );
  INV_X1 U12192 ( .A(n9534), .ZN(n9548) );
  AND2_X1 U12193 ( .A1(n9535), .A2(n9548), .ZN(n15136) );
  NAND2_X1 U12194 ( .A1(n9781), .A2(n15136), .ZN(n9536) );
  NAND2_X1 U12195 ( .A1(n15099), .A2(n11965), .ZN(n9537) );
  NOR2_X1 U12196 ( .A1(n15099), .A2(n9743), .ZN(n9540) );
  MUX2_X1 U12197 ( .A(n9541), .B(n9540), .S(n11965), .Z(n9542) );
  NAND2_X1 U12198 ( .A1(n9524), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n9547) );
  INV_X1 U12199 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n11066) );
  OR2_X1 U12200 ( .A1(n6552), .A2(n11066), .ZN(n9546) );
  XNOR2_X1 U12201 ( .A(P1_REG3_REG_3__SCAN_IN), .B(P1_REG3_REG_4__SCAN_IN), 
        .ZN(n12073) );
  OR2_X1 U12202 ( .A1(n6550), .A2(n12073), .ZN(n9545) );
  INV_X1 U12203 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n9543) );
  OR2_X1 U12204 ( .A1(n9832), .A2(n9543), .ZN(n9544) );
  NAND2_X1 U12205 ( .A1(n9548), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9549) );
  XNOR2_X1 U12206 ( .A(n9549), .B(P1_IR_REG_4__SCAN_IN), .ZN(n11079) );
  NAND2_X1 U12207 ( .A1(n10654), .A2(n10006), .ZN(n9550) );
  MUX2_X1 U12208 ( .A(n15795), .B(n12028), .S(n9743), .Z(n9552) );
  INV_X1 U12209 ( .A(n9552), .ZN(n9554) );
  MUX2_X1 U12210 ( .A(n12028), .B(n15795), .S(n9743), .Z(n9553) );
  INV_X1 U12211 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n9556) );
  NAND2_X1 U12212 ( .A1(n9534), .A2(n9556), .ZN(n9580) );
  NAND2_X1 U12213 ( .A1(n9580), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9557) );
  XNOR2_X1 U12214 ( .A(n9557), .B(P1_IR_REG_5__SCAN_IN), .ZN(n11097) );
  NAND2_X1 U12215 ( .A1(n10690), .A2(n10006), .ZN(n9558) );
  NAND2_X1 U12216 ( .A1(n9947), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n9568) );
  INV_X1 U12217 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n9560) );
  OR2_X1 U12218 ( .A1(n6552), .A2(n9560), .ZN(n9567) );
  INV_X1 U12219 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n9561) );
  OR2_X1 U12220 ( .A1(n9960), .A2(n9561), .ZN(n9566) );
  INV_X1 U12221 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n9563) );
  NAND2_X1 U12222 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .ZN(n9562) );
  NAND2_X1 U12223 ( .A1(n9563), .A2(n9562), .ZN(n9564) );
  NAND2_X1 U12224 ( .A1(n9573), .A2(n9564), .ZN(n15803) );
  OR2_X1 U12225 ( .A1(n6550), .A2(n15803), .ZN(n9565) );
  INV_X1 U12226 ( .A(n12030), .ZN(n15098) );
  MUX2_X1 U12227 ( .A(n12091), .B(n15098), .S(n9635), .Z(n9569) );
  NAND2_X1 U12228 ( .A1(n9838), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n9579) );
  INV_X1 U12229 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n12036) );
  OR2_X1 U12230 ( .A1(n9960), .A2(n12036), .ZN(n9578) );
  INV_X1 U12231 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n9572) );
  NAND2_X1 U12232 ( .A1(n9573), .A2(n9572), .ZN(n9574) );
  NAND2_X1 U12233 ( .A1(n9591), .A2(n9574), .ZN(n12176) );
  OR2_X1 U12234 ( .A1(n6550), .A2(n12176), .ZN(n9577) );
  INV_X1 U12235 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n9575) );
  OR2_X1 U12236 ( .A1(n9832), .A2(n9575), .ZN(n9576) );
  NAND4_X1 U12237 ( .A1(n9579), .A2(n9578), .A3(n9577), .A4(n9576), .ZN(n15097) );
  NAND2_X1 U12238 ( .A1(n10693), .A2(n10006), .ZN(n9583) );
  NAND2_X1 U12239 ( .A1(n9720), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9581) );
  XNOR2_X1 U12240 ( .A(n9581), .B(P1_IR_REG_6__SCAN_IN), .ZN(n11201) );
  AOI22_X1 U12241 ( .A1(n9940), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n9781), .B2(
        n11201), .ZN(n9582) );
  NAND2_X1 U12242 ( .A1(n9583), .A2(n9582), .ZN(n15853) );
  MUX2_X1 U12243 ( .A(n15097), .B(n15853), .S(n9743), .Z(n9585) );
  MUX2_X1 U12244 ( .A(n15853), .B(n15097), .S(n9743), .Z(n9584) );
  INV_X1 U12245 ( .A(n9585), .ZN(n9586) );
  NAND2_X1 U12246 ( .A1(n9587), .A2(n9586), .ZN(n9588) );
  NAND2_X1 U12247 ( .A1(n9589), .A2(n9588), .ZN(n9605) );
  NAND2_X1 U12248 ( .A1(n9947), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n9597) );
  INV_X1 U12249 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n9590) );
  OR2_X1 U12250 ( .A1(n9960), .A2(n9590), .ZN(n9596) );
  INV_X1 U12251 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n12148) );
  NAND2_X1 U12252 ( .A1(n9591), .A2(n12148), .ZN(n9592) );
  NAND2_X1 U12253 ( .A1(n9609), .A2(n9592), .ZN(n15781) );
  OR2_X1 U12254 ( .A1(n6550), .A2(n15781), .ZN(n9595) );
  INV_X1 U12255 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n9593) );
  OR2_X1 U12256 ( .A1(n6552), .A2(n9593), .ZN(n9594) );
  NAND4_X1 U12257 ( .A1(n9597), .A2(n9596), .A3(n9595), .A4(n9594), .ZN(n15096) );
  NAND2_X1 U12258 ( .A1(n10672), .A2(n10006), .ZN(n9603) );
  INV_X1 U12259 ( .A(n9720), .ZN(n9599) );
  NAND2_X1 U12260 ( .A1(n9599), .A2(n7338), .ZN(n9631) );
  NAND2_X1 U12261 ( .A1(n9631), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9600) );
  INV_X1 U12262 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n10868) );
  NAND2_X1 U12263 ( .A1(n9600), .A2(n10868), .ZN(n9616) );
  OR2_X1 U12264 ( .A1(n9600), .A2(n10868), .ZN(n9601) );
  AOI22_X1 U12265 ( .A1(n6561), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n9781), .B2(
        n15163), .ZN(n9602) );
  MUX2_X1 U12266 ( .A(n15096), .B(n15780), .S(n9635), .Z(n9606) );
  MUX2_X1 U12267 ( .A(n15096), .B(n15780), .S(n9743), .Z(n9604) );
  NAND2_X1 U12268 ( .A1(n9524), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n9615) );
  INV_X1 U12269 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n9607) );
  OR2_X1 U12270 ( .A1(n6553), .A2(n9607), .ZN(n9614) );
  INV_X1 U12271 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n9608) );
  NAND2_X1 U12272 ( .A1(n9609), .A2(n9608), .ZN(n9610) );
  NAND2_X1 U12273 ( .A1(n9624), .A2(n9610), .ZN(n12414) );
  OR2_X1 U12274 ( .A1(n6550), .A2(n12414), .ZN(n9613) );
  INV_X1 U12275 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n9611) );
  OR2_X1 U12276 ( .A1(n9832), .A2(n9611), .ZN(n9612) );
  NAND4_X1 U12277 ( .A1(n9615), .A2(n9614), .A3(n9613), .A4(n9612), .ZN(n15095) );
  NAND2_X1 U12278 ( .A1(n9616), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9617) );
  XNOR2_X1 U12279 ( .A(n9617), .B(P1_IR_REG_8__SCAN_IN), .ZN(n11116) );
  AOI22_X1 U12280 ( .A1(n9940), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n11116), 
        .B2(n9781), .ZN(n9618) );
  NAND2_X2 U12281 ( .A1(n9619), .A2(n9618), .ZN(n15869) );
  MUX2_X1 U12282 ( .A(n15095), .B(n15869), .S(n9743), .Z(n9621) );
  MUX2_X1 U12283 ( .A(n15095), .B(n15869), .S(n9635), .Z(n9620) );
  NAND2_X1 U12284 ( .A1(n9524), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n9629) );
  INV_X1 U12285 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n11088) );
  OR2_X1 U12286 ( .A1(n6552), .A2(n11088), .ZN(n9628) );
  INV_X1 U12287 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n9623) );
  NAND2_X1 U12288 ( .A1(n9624), .A2(n9623), .ZN(n9625) );
  NAND2_X1 U12289 ( .A1(n9640), .A2(n9625), .ZN(n12515) );
  OR2_X1 U12290 ( .A1(n6550), .A2(n12515), .ZN(n9627) );
  INV_X1 U12291 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n10993) );
  OR2_X1 U12292 ( .A1(n9832), .A2(n10993), .ZN(n9626) );
  NAND4_X1 U12293 ( .A1(n9629), .A2(n9628), .A3(n9627), .A4(n9626), .ZN(n15094) );
  NAND2_X1 U12294 ( .A1(n10745), .A2(n10006), .ZN(n9634) );
  INV_X1 U12295 ( .A(n10816), .ZN(n9630) );
  NAND2_X1 U12296 ( .A1(n9647), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9632) );
  XNOR2_X1 U12297 ( .A(n9632), .B(P1_IR_REG_9__SCAN_IN), .ZN(n11370) );
  AOI22_X1 U12298 ( .A1(n6561), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n9781), .B2(
        n11370), .ZN(n9633) );
  MUX2_X1 U12299 ( .A(n15094), .B(n15662), .S(n9635), .Z(n9637) );
  MUX2_X1 U12300 ( .A(n15094), .B(n15662), .S(n9743), .Z(n9636) );
  INV_X1 U12301 ( .A(n9637), .ZN(n9638) );
  NAND2_X1 U12302 ( .A1(n9838), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n9646) );
  INV_X1 U12303 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n12366) );
  OR2_X1 U12304 ( .A1(n9960), .A2(n12366), .ZN(n9645) );
  NAND2_X1 U12305 ( .A1(n9640), .A2(n9639), .ZN(n9641) );
  NAND2_X1 U12306 ( .A1(n9661), .A2(n9641), .ZN(n12743) );
  OR2_X1 U12307 ( .A1(n6550), .A2(n12743), .ZN(n9644) );
  INV_X1 U12308 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n9642) );
  OR2_X1 U12309 ( .A1(n9832), .A2(n9642), .ZN(n9643) );
  NAND4_X1 U12310 ( .A1(n9646), .A2(n9645), .A3(n9644), .A4(n9643), .ZN(n15093) );
  NAND2_X1 U12311 ( .A1(n11036), .A2(n10006), .ZN(n9650) );
  NAND2_X1 U12312 ( .A1(n9668), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9648) );
  XNOR2_X1 U12313 ( .A(n9648), .B(P1_IR_REG_10__SCAN_IN), .ZN(n15178) );
  AOI22_X1 U12314 ( .A1(n6561), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n15178), 
        .B2(n9781), .ZN(n9649) );
  MUX2_X1 U12315 ( .A(n15093), .B(n12560), .S(n9743), .Z(n9655) );
  INV_X1 U12316 ( .A(n9651), .ZN(n9954) );
  MUX2_X1 U12317 ( .A(n15093), .B(n12560), .S(n9954), .Z(n9652) );
  NAND2_X1 U12318 ( .A1(n9653), .A2(n9652), .ZN(n9659) );
  INV_X1 U12319 ( .A(n9654), .ZN(n9657) );
  INV_X1 U12320 ( .A(n9655), .ZN(n9656) );
  NAND2_X1 U12321 ( .A1(n9657), .A2(n9656), .ZN(n9658) );
  NAND2_X1 U12322 ( .A1(n9659), .A2(n9658), .ZN(n9674) );
  NAND2_X1 U12323 ( .A1(n9524), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n9667) );
  INV_X1 U12324 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n9660) );
  OR2_X1 U12325 ( .A1(n6553), .A2(n9660), .ZN(n9666) );
  NAND2_X1 U12326 ( .A1(n9661), .A2(n12903), .ZN(n9662) );
  NAND2_X1 U12327 ( .A1(n9678), .A2(n9662), .ZN(n12907) );
  OR2_X1 U12328 ( .A1(n6550), .A2(n12907), .ZN(n9665) );
  INV_X1 U12329 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n9663) );
  OR2_X1 U12330 ( .A1(n9832), .A2(n9663), .ZN(n9664) );
  NAND4_X1 U12331 ( .A1(n9667), .A2(n9666), .A3(n9665), .A4(n9664), .ZN(n15092) );
  NAND2_X1 U12332 ( .A1(n11057), .A2(n10006), .ZN(n9672) );
  INV_X1 U12333 ( .A(n9668), .ZN(n9669) );
  NAND2_X1 U12334 ( .A1(n9669), .A2(n7339), .ZN(n9684) );
  NAND2_X1 U12335 ( .A1(n9684), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9670) );
  XNOR2_X1 U12336 ( .A(n9670), .B(P1_IR_REG_11__SCAN_IN), .ZN(n11557) );
  AOI22_X1 U12337 ( .A1(n11557), .A2(n9781), .B1(n9940), .B2(
        P2_DATAO_REG_11__SCAN_IN), .ZN(n9671) );
  MUX2_X1 U12338 ( .A(n15092), .B(n12902), .S(n9954), .Z(n9675) );
  MUX2_X1 U12339 ( .A(n15092), .B(n12902), .S(n9743), .Z(n9673) );
  INV_X1 U12340 ( .A(n9675), .ZN(n9676) );
  NAND2_X1 U12341 ( .A1(n9947), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n9683) );
  INV_X1 U12342 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n11556) );
  OR2_X1 U12343 ( .A1(n6552), .A2(n11556), .ZN(n9682) );
  INV_X1 U12344 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n9677) );
  OR2_X1 U12345 ( .A1(n9960), .A2(n9677), .ZN(n9681) );
  INV_X1 U12346 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n10812) );
  NAND2_X1 U12347 ( .A1(n9678), .A2(n10812), .ZN(n9679) );
  NAND2_X1 U12348 ( .A1(n9708), .A2(n9679), .ZN(n14973) );
  OR2_X1 U12349 ( .A1(n6550), .A2(n14973), .ZN(n9680) );
  NAND4_X1 U12350 ( .A1(n9683), .A2(n9682), .A3(n9681), .A4(n9680), .ZN(n15520) );
  NAND2_X1 U12351 ( .A1(n11207), .A2(n10006), .ZN(n9689) );
  INV_X1 U12352 ( .A(n9684), .ZN(n9686) );
  INV_X1 U12353 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n9685) );
  NAND2_X1 U12354 ( .A1(n9686), .A2(n9685), .ZN(n9687) );
  NAND2_X1 U12355 ( .A1(n9687), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9694) );
  XNOR2_X1 U12356 ( .A(n9694), .B(P1_IR_REG_12__SCAN_IN), .ZN(n11895) );
  AOI22_X1 U12357 ( .A1(n11895), .A2(n9781), .B1(n9940), .B2(
        P2_DATAO_REG_12__SCAN_IN), .ZN(n9688) );
  NAND2_X2 U12358 ( .A1(n9689), .A2(n9688), .ZN(n15651) );
  MUX2_X1 U12359 ( .A(n15520), .B(n15651), .S(n9743), .Z(n9691) );
  MUX2_X1 U12360 ( .A(n15520), .B(n15651), .S(n9954), .Z(n9690) );
  INV_X1 U12361 ( .A(n9691), .ZN(n9692) );
  INV_X1 U12362 ( .A(n9769), .ZN(n9731) );
  NAND2_X1 U12363 ( .A1(n11588), .A2(n10006), .ZN(n9700) );
  INV_X1 U12364 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n9693) );
  NAND2_X1 U12365 ( .A1(n9694), .A2(n9693), .ZN(n9695) );
  NAND2_X1 U12366 ( .A1(n9695), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9716) );
  INV_X1 U12367 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n9696) );
  NAND2_X1 U12368 ( .A1(n9716), .A2(n9696), .ZN(n9697) );
  NAND2_X1 U12369 ( .A1(n9697), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9698) );
  AOI22_X1 U12370 ( .A1(n15191), .A2(n9781), .B1(n6561), .B2(
        P2_DATAO_REG_14__SCAN_IN), .ZN(n9699) );
  NAND2_X1 U12371 ( .A1(n9710), .A2(n14935), .ZN(n9701) );
  AND2_X1 U12372 ( .A1(n9724), .A2(n9701), .ZN(n15508) );
  NAND2_X1 U12373 ( .A1(n9913), .A2(n15508), .ZN(n9706) );
  INV_X1 U12374 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n12162) );
  OR2_X1 U12375 ( .A1(n9960), .A2(n12162), .ZN(n9705) );
  INV_X1 U12376 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n12167) );
  OR2_X1 U12377 ( .A1(n6552), .A2(n12167), .ZN(n9704) );
  INV_X1 U12378 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n9702) );
  OR2_X1 U12379 ( .A1(n9832), .A2(n9702), .ZN(n9703) );
  NAND4_X1 U12380 ( .A1(n9706), .A2(n9705), .A3(n9704), .A4(n9703), .ZN(n15091) );
  NAND2_X1 U12381 ( .A1(n15639), .A2(n15517), .ZN(n9770) );
  NAND2_X1 U12382 ( .A1(n9838), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n9715) );
  INV_X1 U12383 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n15529) );
  OR2_X1 U12384 ( .A1(n9960), .A2(n15529), .ZN(n9714) );
  INV_X1 U12385 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n9707) );
  NAND2_X1 U12386 ( .A1(n9708), .A2(n9707), .ZN(n9709) );
  NAND2_X1 U12387 ( .A1(n9710), .A2(n9709), .ZN(n15034) );
  OR2_X1 U12388 ( .A1(n6550), .A2(n15034), .ZN(n9713) );
  INV_X1 U12389 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n9711) );
  OR2_X1 U12390 ( .A1(n9832), .A2(n9711), .ZN(n9712) );
  NAND4_X1 U12391 ( .A1(n9715), .A2(n9714), .A3(n9713), .A4(n9712), .ZN(n15502) );
  NAND2_X1 U12392 ( .A1(n11379), .A2(n10006), .ZN(n9718) );
  XNOR2_X1 U12393 ( .A(n9716), .B(P1_IR_REG_13__SCAN_IN), .ZN(n12164) );
  AOI22_X1 U12394 ( .A1(n12164), .A2(n9781), .B1(n9940), .B2(
        P2_DATAO_REG_13__SCAN_IN), .ZN(n9717) );
  MUX2_X1 U12395 ( .A(n15502), .B(n15645), .S(n9954), .Z(n9768) );
  INV_X1 U12396 ( .A(n9768), .ZN(n9730) );
  OAI21_X1 U12397 ( .B1(n9720), .B2(n9719), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n9721) );
  XNOR2_X1 U12398 ( .A(n9721), .B(P1_IR_REG_15__SCAN_IN), .ZN(n12644) );
  AOI22_X1 U12399 ( .A1(n9940), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n9781), 
        .B2(n12644), .ZN(n9722) );
  INV_X1 U12400 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n9723) );
  NAND2_X1 U12401 ( .A1(n9724), .A2(n9723), .ZN(n9725) );
  NAND2_X1 U12402 ( .A1(n9735), .A2(n9725), .ZN(n15492) );
  NOR2_X1 U12403 ( .A1(n15492), .A2(n6550), .ZN(n9729) );
  INV_X1 U12404 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n9726) );
  NOR2_X1 U12405 ( .A1(n9832), .A2(n9726), .ZN(n9728) );
  INV_X1 U12406 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n12631) );
  INV_X1 U12407 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n12642) );
  OAI22_X1 U12408 ( .A1(n6553), .A2(n12631), .B1(n9960), .B2(n12642), .ZN(
        n9727) );
  NAND4_X1 U12409 ( .A1(n9731), .A2(n13029), .A3(n9730), .A4(n10036), .ZN(
        n9734) );
  OAI21_X1 U12410 ( .B1(n13030), .B2(n14993), .A(n15633), .ZN(n9732) );
  OAI211_X1 U12411 ( .C1(n6883), .C2(n15501), .A(n9732), .B(n9954), .ZN(n9733)
         );
  NOR2_X1 U12412 ( .A1(n13032), .A2(n9954), .ZN(n9777) );
  AOI21_X1 U12413 ( .B1(n9734), .B2(n9733), .A(n9777), .ZN(n9767) );
  NAND2_X1 U12414 ( .A1(n9735), .A2(n12651), .ZN(n9736) );
  NAND2_X1 U12415 ( .A1(n9761), .A2(n9736), .ZN(n15472) );
  AOI22_X1 U12416 ( .A1(n9838), .A2(P1_REG1_REG_16__SCAN_IN), .B1(n9524), .B2(
        P1_REG2_REG_16__SCAN_IN), .ZN(n9738) );
  NAND2_X1 U12417 ( .A1(n9947), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n9737) );
  OAI211_X1 U12418 ( .C1(n15472), .C2(n6550), .A(n9738), .B(n9737), .ZN(n15090) );
  INV_X1 U12419 ( .A(n15090), .ZN(n15076) );
  NAND2_X1 U12420 ( .A1(n11548), .A2(n10006), .ZN(n9742) );
  NAND2_X1 U12421 ( .A1(n9739), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9740) );
  XNOR2_X1 U12422 ( .A(n9740), .B(P1_IR_REG_16__SCAN_IN), .ZN(n15205) );
  AOI22_X1 U12423 ( .A1(n6561), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n9781), 
        .B2(n15205), .ZN(n9741) );
  INV_X1 U12424 ( .A(n15628), .ZN(n15477) );
  MUX2_X1 U12425 ( .A(n15076), .B(n15477), .S(n9743), .Z(n9796) );
  INV_X1 U12426 ( .A(n9954), .ZN(n9956) );
  MUX2_X1 U12427 ( .A(n15628), .B(n15090), .S(n9956), .Z(n9795) );
  NAND2_X1 U12428 ( .A1(n9763), .A2(n15052), .ZN(n9744) );
  AND2_X1 U12429 ( .A1(n9785), .A2(n9744), .ZN(n15442) );
  NAND2_X1 U12430 ( .A1(n15442), .A2(n9913), .ZN(n9750) );
  INV_X1 U12431 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n9747) );
  NAND2_X1 U12432 ( .A1(n9838), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n9746) );
  NAND2_X1 U12433 ( .A1(n9947), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n9745) );
  OAI211_X1 U12434 ( .C1(n9960), .C2(n9747), .A(n9746), .B(n9745), .ZN(n9748)
         );
  INV_X1 U12435 ( .A(n9748), .ZN(n9749) );
  NAND2_X1 U12436 ( .A1(n9750), .A2(n9749), .ZN(n15419) );
  INV_X1 U12437 ( .A(n9751), .ZN(n9752) );
  NAND2_X1 U12438 ( .A1(n9752), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9753) );
  XNOR2_X1 U12439 ( .A(n9753), .B(P1_IR_REG_18__SCAN_IN), .ZN(n15227) );
  AOI22_X1 U12440 ( .A1(n9940), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n9781), 
        .B2(n15227), .ZN(n9754) );
  MUX2_X1 U12441 ( .A(n15419), .B(n15616), .S(n9956), .Z(n9798) );
  NAND2_X1 U12442 ( .A1(n15616), .A2(n15419), .ZN(n13010) );
  NAND2_X1 U12443 ( .A1(n11593), .A2(n10006), .ZN(n9759) );
  NAND2_X1 U12444 ( .A1(n9756), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9757) );
  XNOR2_X1 U12445 ( .A(n9757), .B(P1_IR_REG_17__SCAN_IN), .ZN(n15224) );
  AOI22_X1 U12446 ( .A1(n6561), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n9781), 
        .B2(n15224), .ZN(n9758) );
  INV_X1 U12447 ( .A(P1_REG0_REG_17__SCAN_IN), .ZN(n10848) );
  INV_X1 U12448 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n9760) );
  NAND2_X1 U12449 ( .A1(n9761), .A2(n9760), .ZN(n9762) );
  NAND2_X1 U12450 ( .A1(n9763), .A2(n9762), .ZN(n15457) );
  OR2_X1 U12451 ( .A1(n15457), .A2(n6550), .ZN(n9765) );
  AOI22_X1 U12452 ( .A1(n9838), .A2(P1_REG1_REG_17__SCAN_IN), .B1(n9524), .B2(
        P1_REG2_REG_17__SCAN_IN), .ZN(n9764) );
  OAI211_X1 U12453 ( .C1(n9832), .C2(n10848), .A(n9765), .B(n9764), .ZN(n15089) );
  INV_X1 U12454 ( .A(n15089), .ZN(n15432) );
  XNOR2_X1 U12455 ( .A(n15622), .B(n15432), .ZN(n15450) );
  AOI21_X1 U12456 ( .B1(n9798), .B2(n13010), .A(n15450), .ZN(n9797) );
  OAI21_X1 U12457 ( .B1(n9796), .B2(n9795), .A(n9797), .ZN(n9766) );
  NOR2_X1 U12458 ( .A1(n9767), .A2(n9766), .ZN(n9807) );
  NAND2_X1 U12459 ( .A1(n9769), .A2(n9768), .ZN(n9774) );
  AND2_X1 U12460 ( .A1(n10036), .A2(n9770), .ZN(n9771) );
  INV_X1 U12461 ( .A(n9771), .ZN(n9773) );
  INV_X1 U12462 ( .A(n15645), .ZN(n15530) );
  OAI21_X1 U12463 ( .B1(n15505), .B2(n15530), .A(n9771), .ZN(n9772) );
  OAI211_X1 U12464 ( .C1(n9774), .C2(n9773), .A(n9651), .B(n9772), .ZN(n9776)
         );
  NAND2_X1 U12465 ( .A1(n9776), .A2(n9775), .ZN(n9779) );
  INV_X1 U12466 ( .A(n9777), .ZN(n9778) );
  NAND2_X1 U12467 ( .A1(n9779), .A2(n9778), .ZN(n9806) );
  NAND2_X1 U12468 ( .A1(n12141), .A2(n10006), .ZN(n9783) );
  AOI22_X1 U12469 ( .A1(n6561), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n15250), 
        .B2(n9781), .ZN(n9782) );
  INV_X1 U12470 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n9784) );
  NAND2_X1 U12471 ( .A1(n9785), .A2(n9784), .ZN(n9786) );
  NAND2_X1 U12472 ( .A1(n9815), .A2(n9786), .ZN(n15422) );
  OR2_X1 U12473 ( .A1(n15422), .A2(n6550), .ZN(n9791) );
  INV_X1 U12474 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n15237) );
  NAND2_X1 U12475 ( .A1(n9947), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n9788) );
  NAND2_X1 U12476 ( .A1(n9524), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n9787) );
  OAI211_X1 U12477 ( .C1(n6552), .C2(n15237), .A(n9788), .B(n9787), .ZN(n9789)
         );
  INV_X1 U12478 ( .A(n9789), .ZN(n9790) );
  NAND2_X1 U12479 ( .A1(n9791), .A2(n9790), .ZN(n15088) );
  XNOR2_X1 U12480 ( .A(n15605), .B(n15088), .ZN(n13012) );
  NOR2_X1 U12481 ( .A1(n15089), .A2(n9956), .ZN(n9794) );
  NAND2_X1 U12482 ( .A1(n15089), .A2(n9956), .ZN(n9792) );
  NOR2_X1 U12483 ( .A1(n15622), .A2(n9792), .ZN(n9793) );
  AOI21_X1 U12484 ( .B1(n9794), .B2(n15622), .A(n9793), .ZN(n9803) );
  NAND3_X1 U12485 ( .A1(n9797), .A2(n9796), .A3(n9795), .ZN(n9802) );
  INV_X1 U12486 ( .A(n9803), .ZN(n9800) );
  INV_X1 U12487 ( .A(n9798), .ZN(n9799) );
  OAI21_X1 U12488 ( .B1(n6633), .B2(n9800), .A(n9799), .ZN(n9801) );
  OAI211_X1 U12489 ( .C1(n9803), .C2(n13010), .A(n9802), .B(n9801), .ZN(n9804)
         );
  AOI21_X1 U12490 ( .B1(n9807), .B2(n9806), .A(n9805), .ZN(n9811) );
  INV_X1 U12491 ( .A(n15088), .ZN(n15433) );
  NOR2_X1 U12492 ( .A1(n15433), .A2(n9956), .ZN(n9809) );
  NOR2_X1 U12493 ( .A1(n15088), .A2(n9954), .ZN(n9808) );
  MUX2_X1 U12494 ( .A(n9809), .B(n9808), .S(n15605), .Z(n9810) );
  NAND2_X1 U12495 ( .A1(n9940), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n9813) );
  INV_X1 U12496 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n15024) );
  NAND2_X1 U12497 ( .A1(n9815), .A2(n15024), .ZN(n9816) );
  NAND2_X1 U12498 ( .A1(n9817), .A2(n9816), .ZN(n15022) );
  OR2_X1 U12499 ( .A1(n15022), .A2(n6550), .ZN(n9822) );
  INV_X1 U12500 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n10802) );
  NAND2_X1 U12501 ( .A1(n9947), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n9819) );
  NAND2_X1 U12502 ( .A1(n9524), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n9818) );
  OAI211_X1 U12503 ( .C1(n6553), .C2(n10802), .A(n9819), .B(n9818), .ZN(n9820)
         );
  INV_X1 U12504 ( .A(n9820), .ZN(n9821) );
  MUX2_X1 U12505 ( .A(n15602), .B(n15421), .S(n9956), .Z(n9823) );
  MUX2_X1 U12506 ( .A(n15421), .B(n15602), .S(n9956), .Z(n9824) );
  MUX2_X1 U12507 ( .A(n15597), .B(n15363), .S(n9956), .Z(n9825) );
  OR2_X1 U12508 ( .A1(n9826), .A2(n9991), .ZN(n9827) );
  INV_X1 U12509 ( .A(n15370), .ZN(n15591) );
  INV_X1 U12510 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n15044) );
  NAND2_X1 U12511 ( .A1(n9828), .A2(n15044), .ZN(n9829) );
  AND2_X1 U12512 ( .A1(n9851), .A2(n9829), .ZN(n15368) );
  NAND2_X1 U12513 ( .A1(n15368), .A2(n9913), .ZN(n9835) );
  INV_X1 U12514 ( .A(P1_REG0_REG_22__SCAN_IN), .ZN(n11016) );
  NAND2_X1 U12515 ( .A1(n9838), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n9831) );
  NAND2_X1 U12516 ( .A1(n9524), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n9830) );
  OAI211_X1 U12517 ( .C1(n9832), .C2(n11016), .A(n9831), .B(n9830), .ZN(n9833)
         );
  INV_X1 U12518 ( .A(n9833), .ZN(n9834) );
  MUX2_X1 U12519 ( .A(n15591), .B(n15087), .S(n9956), .Z(n9837) );
  MUX2_X1 U12520 ( .A(n15391), .B(n15370), .S(n9956), .Z(n9836) );
  XNOR2_X1 U12521 ( .A(n9851), .B(P1_REG3_REG_23__SCAN_IN), .ZN(n15349) );
  NAND2_X1 U12522 ( .A1(n15349), .A2(n9913), .ZN(n9843) );
  INV_X1 U12523 ( .A(P1_REG0_REG_23__SCAN_IN), .ZN(n10947) );
  NAND2_X1 U12524 ( .A1(n9524), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n9840) );
  NAND2_X1 U12525 ( .A1(n9838), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n9839) );
  OAI211_X1 U12526 ( .C1(n9832), .C2(n10947), .A(n9840), .B(n9839), .ZN(n9841)
         );
  INV_X1 U12527 ( .A(n9841), .ZN(n9842) );
  NAND2_X1 U12528 ( .A1(n12317), .A2(n10006), .ZN(n9845) );
  NAND2_X1 U12529 ( .A1(n9940), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n9844) );
  INV_X1 U12530 ( .A(n15586), .ZN(n15356) );
  MUX2_X1 U12531 ( .A(n15332), .B(n15356), .S(n9956), .Z(n9894) );
  NAND2_X1 U12532 ( .A1(n12577), .A2(n10006), .ZN(n9847) );
  NAND2_X1 U12533 ( .A1(n9940), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n9846) );
  AND2_X1 U12534 ( .A1(P1_REG3_REG_24__SCAN_IN), .A2(P1_REG3_REG_23__SCAN_IN), 
        .ZN(n9848) );
  INV_X1 U12535 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n9850) );
  INV_X1 U12536 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n9849) );
  OAI21_X1 U12537 ( .B1(n9851), .B2(n9850), .A(n9849), .ZN(n9852) );
  NAND2_X1 U12538 ( .A1(n9881), .A2(n9852), .ZN(n15013) );
  INV_X1 U12539 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n9855) );
  NAND2_X1 U12540 ( .A1(n9524), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n9854) );
  NAND2_X1 U12541 ( .A1(n9947), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n9853) );
  OAI211_X1 U12542 ( .C1(n6553), .C2(n9855), .A(n9854), .B(n9853), .ZN(n9856)
         );
  INV_X1 U12543 ( .A(n9856), .ZN(n9857) );
  INV_X1 U12544 ( .A(n15306), .ZN(n13045) );
  MUX2_X1 U12545 ( .A(n15578), .B(n13045), .S(n9954), .Z(n9926) );
  MUX2_X1 U12546 ( .A(n15341), .B(n15306), .S(n9956), .Z(n9925) );
  AOI22_X1 U12547 ( .A1(n9895), .A2(n9894), .B1(n9926), .B2(n9925), .ZN(n9897)
         );
  INV_X1 U12548 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n10935) );
  INV_X1 U12549 ( .A(n9870), .ZN(n9860) );
  INV_X1 U12550 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n9861) );
  NAND2_X1 U12551 ( .A1(n9870), .A2(n9861), .ZN(n9862) );
  NAND2_X1 U12552 ( .A1(n13079), .A2(n9862), .ZN(n13060) );
  INV_X1 U12553 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n10985) );
  NAND2_X1 U12554 ( .A1(n9524), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n9864) );
  NAND2_X1 U12555 ( .A1(n9947), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n9863) );
  OAI211_X1 U12556 ( .C1(n6553), .C2(n10985), .A(n9864), .B(n9863), .ZN(n9865)
         );
  INV_X1 U12557 ( .A(n9865), .ZN(n9866) );
  NAND2_X1 U12558 ( .A1(n6561), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n9867) );
  INV_X1 U12559 ( .A(n15559), .ZN(n13087) );
  MUX2_X1 U12560 ( .A(n15066), .B(n13087), .S(n9956), .Z(n9908) );
  MUX2_X1 U12561 ( .A(n15297), .B(n15559), .S(n9954), .Z(n9906) );
  NAND2_X1 U12562 ( .A1(n9908), .A2(n9906), .ZN(n9880) );
  NAND2_X1 U12563 ( .A1(n9883), .A2(n10935), .ZN(n9869) );
  NAND2_X1 U12564 ( .A1(n15298), .A2(n9913), .ZN(n9876) );
  INV_X1 U12565 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n9873) );
  NAND2_X1 U12566 ( .A1(n9947), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n9872) );
  NAND2_X1 U12567 ( .A1(n9524), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n9871) );
  OAI211_X1 U12568 ( .C1(n6552), .C2(n9873), .A(n9872), .B(n9871), .ZN(n9874)
         );
  INV_X1 U12569 ( .A(n9874), .ZN(n9875) );
  NAND2_X1 U12570 ( .A1(n14915), .A2(n10006), .ZN(n9878) );
  NAND2_X1 U12571 ( .A1(n6561), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n9877) );
  MUX2_X1 U12572 ( .A(n13055), .B(n15565), .S(n9956), .Z(n9903) );
  MUX2_X1 U12573 ( .A(n15301), .B(n15086), .S(n9956), .Z(n9902) );
  NAND2_X1 U12574 ( .A1(n9903), .A2(n9902), .ZN(n9879) );
  NAND2_X1 U12575 ( .A1(n9880), .A2(n9879), .ZN(n9898) );
  INV_X1 U12576 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n14981) );
  NAND2_X1 U12577 ( .A1(n9881), .A2(n14981), .ZN(n9882) );
  NAND2_X1 U12578 ( .A1(n9883), .A2(n9882), .ZN(n15314) );
  INV_X1 U12579 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n9886) );
  NAND2_X1 U12580 ( .A1(n9947), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n9885) );
  NAND2_X1 U12581 ( .A1(n9524), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n9884) );
  OAI211_X1 U12582 ( .C1(n6552), .C2(n9886), .A(n9885), .B(n9884), .ZN(n9887)
         );
  INV_X1 U12583 ( .A(n9887), .ZN(n9888) );
  INV_X1 U12584 ( .A(n15330), .ZN(n13043) );
  NAND2_X1 U12585 ( .A1(n12789), .A2(n10006), .ZN(n9891) );
  NAND2_X1 U12586 ( .A1(n6561), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n9890) );
  INV_X1 U12587 ( .A(n15318), .ZN(n15572) );
  MUX2_X1 U12588 ( .A(n13043), .B(n15572), .S(n9954), .Z(n9900) );
  MUX2_X1 U12589 ( .A(n15318), .B(n15330), .S(n9954), .Z(n9899) );
  NOR2_X1 U12590 ( .A1(n9900), .A2(n9899), .ZN(n9892) );
  NOR2_X1 U12591 ( .A1(n9898), .A2(n9892), .ZN(n9929) );
  MUX2_X1 U12592 ( .A(n15586), .B(n15362), .S(n9956), .Z(n9893) );
  OAI21_X1 U12593 ( .B1(n9895), .B2(n9894), .A(n9893), .ZN(n9896) );
  INV_X1 U12594 ( .A(n9898), .ZN(n9901) );
  NAND3_X1 U12595 ( .A1(n9901), .A2(n9900), .A3(n9899), .ZN(n9924) );
  INV_X1 U12596 ( .A(n9902), .ZN(n9905) );
  INV_X1 U12597 ( .A(n9903), .ZN(n9904) );
  NAND2_X1 U12598 ( .A1(n9905), .A2(n9904), .ZN(n9907) );
  NAND2_X1 U12599 ( .A1(n9908), .A2(n9907), .ZN(n9912) );
  INV_X1 U12600 ( .A(n9906), .ZN(n9911) );
  INV_X1 U12601 ( .A(n9907), .ZN(n9910) );
  INV_X1 U12602 ( .A(n9908), .ZN(n9909) );
  AOI22_X1 U12603 ( .A1(n9912), .A2(n9911), .B1(n9910), .B2(n9909), .ZN(n9923)
         );
  XNOR2_X1 U12604 ( .A(n13079), .B(P1_REG3_REG_28__SCAN_IN), .ZN(n15281) );
  NAND2_X1 U12605 ( .A1(n15281), .A2(n9913), .ZN(n9919) );
  INV_X1 U12606 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n9916) );
  NAND2_X1 U12607 ( .A1(n9524), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n9915) );
  NAND2_X1 U12608 ( .A1(n9947), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n9914) );
  OAI211_X1 U12609 ( .C1(n6553), .C2(n9916), .A(n9915), .B(n9914), .ZN(n9917)
         );
  INV_X1 U12610 ( .A(n9917), .ZN(n9918) );
  NAND2_X1 U12611 ( .A1(n14907), .A2(n10006), .ZN(n9921) );
  NAND2_X1 U12612 ( .A1(n6561), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n9920) );
  INV_X1 U12613 ( .A(n15553), .ZN(n15284) );
  MUX2_X1 U12614 ( .A(n14927), .B(n15284), .S(n9954), .Z(n9988) );
  MUX2_X1 U12615 ( .A(n15085), .B(n15553), .S(n9651), .Z(n9987) );
  NAND2_X1 U12616 ( .A1(n9988), .A2(n9987), .ZN(n9922) );
  AND3_X1 U12617 ( .A1(n9924), .A2(n9923), .A3(n9922), .ZN(n9931) );
  INV_X1 U12618 ( .A(n9925), .ZN(n9928) );
  INV_X1 U12619 ( .A(n9926), .ZN(n9927) );
  NAND3_X1 U12620 ( .A1(n9929), .A2(n9928), .A3(n9927), .ZN(n9930) );
  OAI21_X2 U12621 ( .B1(n9934), .B2(n9933), .A(n9932), .ZN(n9968) );
  INV_X1 U12622 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n15694) );
  INV_X1 U12623 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n14905) );
  MUX2_X1 U12624 ( .A(n15694), .B(n14905), .S(n10696), .Z(n9935) );
  XNOR2_X1 U12625 ( .A(n9935), .B(SI_29_), .ZN(n9967) );
  NAND2_X1 U12626 ( .A1(n9935), .A2(n13131), .ZN(n9993) );
  MUX2_X1 U12627 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(P1_DATAO_REG_30__SCAN_IN), 
        .S(n10696), .Z(n9936) );
  NAND2_X1 U12628 ( .A1(n9936), .A2(SI_30_), .ZN(n9997) );
  INV_X1 U12629 ( .A(n9936), .ZN(n9937) );
  INV_X1 U12630 ( .A(SI_30_), .ZN(n13291) );
  NAND2_X1 U12631 ( .A1(n9937), .A2(n13291), .ZN(n9994) );
  AND2_X1 U12632 ( .A1(n9997), .A2(n9994), .ZN(n9938) );
  NAND2_X1 U12633 ( .A1(n6561), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n9941) );
  INV_X1 U12634 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n10894) );
  NAND2_X1 U12635 ( .A1(n9947), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n9944) );
  INV_X1 U12636 ( .A(P1_REG2_REG_31__SCAN_IN), .ZN(n15254) );
  OR2_X1 U12637 ( .A1(n9960), .A2(n15254), .ZN(n9943) );
  OAI211_X1 U12638 ( .C1(n6553), .C2(n10894), .A(n9944), .B(n9943), .ZN(n15256) );
  INV_X1 U12639 ( .A(n9945), .ZN(n9946) );
  AOI21_X1 U12640 ( .B1(n15256), .B2(n9956), .A(n9946), .ZN(n9952) );
  INV_X1 U12641 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n9950) );
  NAND2_X1 U12642 ( .A1(n9947), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n9949) );
  INV_X1 U12643 ( .A(P1_REG2_REG_30__SCAN_IN), .ZN(n15262) );
  OR2_X1 U12644 ( .A1(n9960), .A2(n15262), .ZN(n9948) );
  OAI211_X1 U12645 ( .C1(n6552), .C2(n9950), .A(n9949), .B(n9948), .ZN(n15084)
         );
  INV_X1 U12646 ( .A(n15084), .ZN(n9951) );
  NOR2_X1 U12647 ( .A1(n9952), .A2(n9951), .ZN(n9953) );
  OR2_X1 U12648 ( .A1(n12097), .A2(n12140), .ZN(n10060) );
  OAI21_X1 U12649 ( .B1(n15256), .B2(n10060), .A(n15084), .ZN(n9955) );
  INV_X1 U12650 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n13078) );
  OR2_X1 U12651 ( .A1(n6550), .A2(n13078), .ZN(n9958) );
  OR2_X1 U12652 ( .A1(n13079), .A2(n9958), .ZN(n9966) );
  INV_X1 U12653 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n9963) );
  NAND2_X1 U12654 ( .A1(n9947), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n9962) );
  INV_X1 U12655 ( .A(P1_REG2_REG_29__SCAN_IN), .ZN(n9959) );
  OR2_X1 U12656 ( .A1(n9960), .A2(n9959), .ZN(n9961) );
  OAI211_X1 U12657 ( .C1(n9963), .C2(n6552), .A(n9962), .B(n9961), .ZN(n9964)
         );
  INV_X1 U12658 ( .A(n9964), .ZN(n9965) );
  NAND2_X1 U12659 ( .A1(n9966), .A2(n9965), .ZN(n15272) );
  INV_X1 U12660 ( .A(n15272), .ZN(n10046) );
  NAND2_X1 U12661 ( .A1(n14902), .A2(n10006), .ZN(n9970) );
  NAND2_X1 U12662 ( .A1(n9940), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n9969) );
  MUX2_X1 U12663 ( .A(n15272), .B(n13076), .S(n9651), .Z(n9971) );
  INV_X1 U12664 ( .A(n9971), .ZN(n9974) );
  INV_X1 U12665 ( .A(n9972), .ZN(n9973) );
  AND2_X1 U12666 ( .A1(n9974), .A2(n9973), .ZN(n9980) );
  INV_X1 U12667 ( .A(n9980), .ZN(n9975) );
  INV_X1 U12668 ( .A(n9976), .ZN(n9979) );
  INV_X1 U12669 ( .A(n9977), .ZN(n9978) );
  OAI21_X1 U12670 ( .B1(n9980), .B2(n9979), .A(n9978), .ZN(n9981) );
  INV_X1 U12671 ( .A(n9981), .ZN(n9982) );
  OR2_X1 U12672 ( .A1(n7133), .A2(n10719), .ZN(n9990) );
  OR2_X1 U12673 ( .A1(n11472), .A2(n9780), .ZN(n11850) );
  NAND2_X1 U12674 ( .A1(n9990), .A2(n11850), .ZN(n10012) );
  INV_X1 U12675 ( .A(n10012), .ZN(n10009) );
  MUX2_X1 U12676 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n9991), .Z(n9992) );
  INV_X1 U12677 ( .A(SI_31_), .ZN(n13963) );
  XNOR2_X1 U12678 ( .A(n9992), .B(n13963), .ZN(n9996) );
  NAND2_X1 U12679 ( .A1(n9996), .A2(n9997), .ZN(n10004) );
  NAND2_X1 U12680 ( .A1(n9994), .A2(n9993), .ZN(n10000) );
  NOR2_X1 U12681 ( .A1(n10000), .A2(n9996), .ZN(n9995) );
  NAND2_X1 U12682 ( .A1(n10005), .A2(n9995), .ZN(n10003) );
  INV_X1 U12683 ( .A(n9996), .ZN(n10001) );
  INV_X1 U12684 ( .A(n9997), .ZN(n9998) );
  XNOR2_X1 U12685 ( .A(n10001), .B(n9998), .ZN(n9999) );
  OAI21_X1 U12686 ( .B1(n10001), .B2(n10000), .A(n9999), .ZN(n10002) );
  NAND2_X1 U12687 ( .A1(n14895), .A2(n10006), .ZN(n10008) );
  NAND2_X1 U12688 ( .A1(n9940), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(n10007) );
  XNOR2_X1 U12689 ( .A(n15258), .B(n15256), .ZN(n10045) );
  NAND3_X1 U12690 ( .A1(n10010), .A2(n10009), .A3(n10045), .ZN(n10055) );
  OR2_X1 U12691 ( .A1(n12097), .A2(n10011), .ZN(n10013) );
  NAND2_X1 U12692 ( .A1(n10012), .A2(n10013), .ZN(n10019) );
  NOR3_X1 U12693 ( .A1(n15541), .A2(n15256), .A3(n10019), .ZN(n10018) );
  NAND2_X1 U12694 ( .A1(n15258), .A2(n9651), .ZN(n10023) );
  NOR3_X1 U12695 ( .A1(n10023), .A2(n15256), .A3(n10012), .ZN(n10017) );
  NOR2_X1 U12696 ( .A1(n15258), .A2(n9743), .ZN(n10020) );
  XNOR2_X1 U12697 ( .A(n10020), .B(n10012), .ZN(n10015) );
  INV_X1 U12698 ( .A(n15256), .ZN(n10014) );
  INV_X1 U12699 ( .A(n10013), .ZN(n10050) );
  NOR4_X1 U12700 ( .A1(n10015), .A2(n10014), .A3(n10050), .A4(n15258), .ZN(
        n10016) );
  AOI211_X1 U12701 ( .C1(n10018), .C2(n10023), .A(n10017), .B(n10016), .ZN(
        n10054) );
  AOI21_X1 U12702 ( .B1(n10020), .B2(n15256), .A(n10019), .ZN(n10021) );
  XOR2_X1 U12703 ( .A(n15084), .B(n15265), .Z(n10048) );
  NAND2_X1 U12704 ( .A1(n15553), .A2(n14927), .ZN(n13088) );
  NAND2_X1 U12705 ( .A1(n13088), .A2(n10024), .ZN(n13065) );
  NAND2_X1 U12706 ( .A1(n15301), .A2(n13055), .ZN(n13053) );
  OR2_X1 U12707 ( .A1(n15301), .A2(n13055), .ZN(n10025) );
  INV_X1 U12708 ( .A(n15351), .ZN(n15348) );
  XNOR2_X1 U12709 ( .A(n15370), .B(n15391), .ZN(n15374) );
  AND2_X1 U12710 ( .A1(n13012), .A2(n15374), .ZN(n10041) );
  NAND2_X1 U12711 ( .A1(n15602), .A2(n15390), .ZN(n10026) );
  XNOR2_X1 U12712 ( .A(n15628), .B(n15076), .ZN(n15467) );
  XNOR2_X1 U12713 ( .A(n15645), .B(n13027), .ZN(n15532) );
  XNOR2_X1 U12714 ( .A(n12902), .B(n15092), .ZN(n12720) );
  NAND2_X1 U12715 ( .A1(n12560), .A2(n12904), .ZN(n12549) );
  NAND2_X1 U12716 ( .A1(n12553), .A2(n12549), .ZN(n12558) );
  INV_X1 U12717 ( .A(n12558), .ZN(n12363) );
  AND2_X1 U12718 ( .A1(n10028), .A2(n10027), .ZN(n15825) );
  XNOR2_X1 U12719 ( .A(n10123), .B(n11795), .ZN(n11478) );
  NAND4_X1 U12720 ( .A1(n15825), .A2(n11804), .A3(n7826), .A4(n11478), .ZN(
        n10029) );
  XNOR2_X1 U12721 ( .A(n15795), .B(n15792), .ZN(n11807) );
  NOR2_X1 U12722 ( .A1(n10029), .A2(n11807), .ZN(n10031) );
  INV_X1 U12723 ( .A(n15776), .ZN(n10030) );
  INV_X1 U12724 ( .A(n15097), .ZN(n12197) );
  XNOR2_X1 U12725 ( .A(n12197), .B(n15853), .ZN(n12211) );
  INV_X1 U12726 ( .A(n12211), .ZN(n12195) );
  XNOR2_X1 U12727 ( .A(n12030), .B(n15843), .ZN(n15799) );
  NAND4_X1 U12728 ( .A1(n10031), .A2(n10030), .A3(n12195), .A4(n15799), .ZN(
        n10032) );
  NOR2_X1 U12729 ( .A1(n10032), .A2(n12337), .ZN(n10033) );
  XNOR2_X1 U12730 ( .A(n15662), .B(n12413), .ZN(n12357) );
  NAND4_X1 U12731 ( .A1(n12720), .A2(n12363), .A3(n10033), .A4(n12359), .ZN(
        n10034) );
  OR3_X1 U12732 ( .A1(n15532), .A2(n7175), .A3(n10034), .ZN(n10035) );
  NOR2_X1 U12733 ( .A1(n15467), .A2(n10035), .ZN(n10038) );
  NOR2_X1 U12734 ( .A1(n15485), .A2(n15450), .ZN(n10037) );
  NAND4_X1 U12735 ( .A1(n15434), .A2(n13029), .A3(n10038), .A4(n10037), .ZN(
        n10039) );
  NOR2_X1 U12736 ( .A1(n13039), .A2(n10039), .ZN(n10040) );
  INV_X1 U12737 ( .A(n15385), .ZN(n15387) );
  NAND4_X1 U12738 ( .A1(n15326), .A2(n10041), .A3(n10040), .A4(n15387), .ZN(
        n10042) );
  NOR4_X1 U12739 ( .A1(n15293), .A2(n15348), .A3(n13021), .A4(n10042), .ZN(
        n10044) );
  INV_X1 U12740 ( .A(n13054), .ZN(n10043) );
  NAND4_X1 U12741 ( .A1(n10045), .A2(n15269), .A3(n10044), .A4(n10043), .ZN(
        n10047) );
  NOR3_X1 U12742 ( .A1(n10048), .A2(n10047), .A3(n13068), .ZN(n10049) );
  XNOR2_X1 U12743 ( .A(n10049), .B(n9780), .ZN(n10051) );
  NAND2_X1 U12744 ( .A1(n10051), .A2(n10050), .ZN(n10052) );
  INV_X1 U12745 ( .A(n10056), .ZN(n10057) );
  NAND2_X1 U12746 ( .A1(n10057), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10058) );
  XNOR2_X1 U12747 ( .A(n10058), .B(P1_IR_REG_23__SCAN_IN), .ZN(n10072) );
  AND2_X1 U12748 ( .A1(n10072), .A2(P1_STATE_REG_SCAN_IN), .ZN(n12318) );
  INV_X1 U12749 ( .A(P1_B_REG_SCAN_IN), .ZN(n13080) );
  NAND2_X1 U12750 ( .A1(n15250), .A2(n15705), .ZN(n10059) );
  NAND2_X1 U12751 ( .A1(n15611), .A2(n10719), .ZN(n11352) );
  NAND2_X1 U12752 ( .A1(n10063), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10062) );
  NAND2_X1 U12753 ( .A1(n6680), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10065) );
  MUX2_X1 U12754 ( .A(P1_IR_REG_31__SCAN_IN), .B(n10065), .S(
        P1_IR_REG_24__SCAN_IN), .Z(n10066) );
  NAND2_X1 U12755 ( .A1(n10066), .A2(n10063), .ZN(n12579) );
  NOR2_X1 U12756 ( .A1(n12794), .A2(n12579), .ZN(n10071) );
  INV_X1 U12757 ( .A(n9459), .ZN(n10069) );
  INV_X1 U12758 ( .A(n10072), .ZN(n10718) );
  NAND2_X1 U12759 ( .A1(n11352), .A2(n10684), .ZN(n11465) );
  INV_X1 U12760 ( .A(n15119), .ZN(n11071) );
  NOR3_X1 U12761 ( .A1(n11465), .A2(n15699), .A3(n15431), .ZN(n10074) );
  AOI211_X1 U12762 ( .C1(n12318), .C2(n10353), .A(n13080), .B(n10074), .ZN(
        n10075) );
  INV_X1 U12763 ( .A(n10075), .ZN(n10076) );
  OAI21_X1 U12764 ( .B1(n10077), .B2(n13458), .A(n10575), .ZN(n13661) );
  INV_X1 U12765 ( .A(n10078), .ZN(n10079) );
  AOI21_X1 U12766 ( .B1(n13458), .B2(n10080), .A(n10079), .ZN(n10084) );
  NAND2_X1 U12767 ( .A1(n13661), .A2(n16054), .ZN(n10083) );
  OAI22_X1 U12768 ( .A1(n12979), .A2(n13817), .B1(n13684), .B2(n13815), .ZN(
        n10081) );
  INV_X1 U12769 ( .A(n10081), .ZN(n10082) );
  OR2_X1 U12770 ( .A1(n10085), .A2(n13482), .ZN(n11412) );
  NAND2_X1 U12771 ( .A1(n13468), .A2(n10086), .ZN(n11595) );
  OAI21_X1 U12772 ( .B1(n11422), .B2(n11412), .A(n13486), .ZN(n10089) );
  INV_X1 U12773 ( .A(n10087), .ZN(n10090) );
  NAND2_X1 U12774 ( .A1(n10089), .A2(n11424), .ZN(n10093) );
  INV_X1 U12775 ( .A(n11422), .ZN(n11416) );
  NAND3_X1 U12776 ( .A1(n11419), .A2(n11416), .A3(n11411), .ZN(n10092) );
  OR2_X1 U12777 ( .A1(n13833), .A2(n16092), .ZN(n10097) );
  INV_X1 U12778 ( .A(n13460), .ZN(n13835) );
  INV_X1 U12779 ( .A(P3_REG0_REG_27__SCAN_IN), .ZN(n10094) );
  OAI22_X1 U12780 ( .A1(n13835), .A2(n13918), .B1(n16094), .B2(n10094), .ZN(
        n10095) );
  INV_X1 U12781 ( .A(n10095), .ZN(n10096) );
  NAND2_X1 U12782 ( .A1(n10097), .A2(n10096), .ZN(P3_U3454) );
  OR2_X1 U12783 ( .A1(n10111), .A2(n16092), .ZN(n10099) );
  NAND2_X1 U12784 ( .A1(n16092), .A2(n10905), .ZN(n10098) );
  NAND2_X1 U12785 ( .A1(n10099), .A2(n10098), .ZN(n10103) );
  INV_X1 U12786 ( .A(n16070), .ZN(n11790) );
  INV_X1 U12787 ( .A(n10100), .ZN(n13301) );
  OAI22_X1 U12788 ( .A1(n10113), .A2(n13955), .B1(n13301), .B2(n13918), .ZN(
        n10101) );
  INV_X1 U12789 ( .A(n10101), .ZN(n10102) );
  NAND2_X1 U12790 ( .A1(n10103), .A2(n10102), .ZN(P3_U3456) );
  OAI22_X1 U12791 ( .A1(n16055), .A2(n10104), .B1(n13332), .B2(n11708), .ZN(
        n10105) );
  AOI21_X1 U12792 ( .B1(n10105), .B2(n13481), .A(n13468), .ZN(n10107) );
  MUX2_X1 U12793 ( .A(n10108), .B(n10107), .S(n10106), .Z(n10110) );
  OR2_X1 U12794 ( .A1(n10111), .A2(n16103), .ZN(n10112) );
  NAND2_X1 U12795 ( .A1(n10112), .A2(n7977), .ZN(n10116) );
  INV_X1 U12796 ( .A(n16055), .ZN(n13869) );
  OAI22_X1 U12797 ( .A1(n10113), .A2(n13883), .B1(n13301), .B2(n13860), .ZN(
        n10114) );
  INV_X1 U12798 ( .A(n10114), .ZN(n10115) );
  NAND2_X1 U12799 ( .A1(n10116), .A2(n10115), .ZN(P3_U3488) );
  NAND2_X1 U12800 ( .A1(n10140), .A2(n11483), .ZN(n10134) );
  AND2_X2 U12801 ( .A1(n11472), .A2(n11471), .ZN(n11474) );
  INV_X1 U12802 ( .A(n11474), .ZN(n10154) );
  AND2_X1 U12803 ( .A1(n10134), .A2(n10154), .ZN(n10119) );
  NAND2_X1 U12804 ( .A1(n10135), .A2(n10119), .ZN(n10122) );
  INV_X1 U12805 ( .A(n10134), .ZN(n10120) );
  NAND2_X1 U12806 ( .A1(n10120), .A2(n11474), .ZN(n10121) );
  NAND2_X1 U12807 ( .A1(n10122), .A2(n10121), .ZN(n10126) );
  NAND2_X1 U12808 ( .A1(n10340), .A2(n11483), .ZN(n10124) );
  XNOR2_X1 U12809 ( .A(n10133), .B(n10126), .ZN(n11488) );
  INV_X1 U12810 ( .A(n10342), .ZN(n10127) );
  NAND2_X1 U12811 ( .A1(n7136), .A2(n10127), .ZN(n10129) );
  INV_X1 U12812 ( .A(n10607), .ZN(n10130) );
  AOI22_X1 U12813 ( .A1(n10340), .A2(n7137), .B1(n10130), .B2(
        P1_IR_REG_0__SCAN_IN), .ZN(n10128) );
  AND2_X1 U12814 ( .A1(n10129), .A2(n10128), .ZN(n11351) );
  AOI22_X1 U12815 ( .A1(n10140), .A2(n7137), .B1(n10130), .B2(
        P1_REG1_REG_0__SCAN_IN), .ZN(n10131) );
  NAND2_X1 U12816 ( .A1(n11349), .A2(n10132), .ZN(n11490) );
  NAND2_X1 U12817 ( .A1(n11488), .A2(n11490), .ZN(n11489) );
  INV_X1 U12818 ( .A(n10133), .ZN(n10138) );
  NAND2_X1 U12819 ( .A1(n10135), .A2(n10134), .ZN(n10136) );
  XNOR2_X1 U12820 ( .A(n10136), .B(n11474), .ZN(n10137) );
  NAND2_X1 U12821 ( .A1(n10138), .A2(n10137), .ZN(n10139) );
  NAND2_X1 U12822 ( .A1(n11489), .A2(n10139), .ZN(n13094) );
  INV_X2 U12823 ( .A(n10348), .ZN(n10326) );
  NAND2_X1 U12824 ( .A1(n10144), .A2(n10326), .ZN(n10142) );
  NAND2_X1 U12825 ( .A1(n10142), .A2(n10141), .ZN(n10143) );
  XNOR2_X1 U12826 ( .A(n10143), .B(n11474), .ZN(n10149) );
  INV_X1 U12827 ( .A(n10144), .ZN(n11956) );
  OR2_X1 U12828 ( .A1(n11956), .A2(n10342), .ZN(n10146) );
  NAND2_X1 U12829 ( .A1(n10146), .A2(n10145), .ZN(n10147) );
  XNOR2_X1 U12830 ( .A(n10149), .B(n10147), .ZN(n13095) );
  INV_X1 U12831 ( .A(n10147), .ZN(n10148) );
  NAND2_X1 U12832 ( .A1(n10149), .A2(n10148), .ZN(n10150) );
  NAND2_X1 U12833 ( .A1(n13093), .A2(n10150), .ZN(n11755) );
  INV_X1 U12834 ( .A(n11755), .ZN(n10159) );
  NAND2_X1 U12835 ( .A1(n15099), .A2(n10326), .ZN(n10153) );
  NAND2_X1 U12836 ( .A1(n10346), .A2(n11965), .ZN(n10152) );
  NAND2_X1 U12837 ( .A1(n10153), .A2(n10152), .ZN(n10155) );
  XNOR2_X1 U12838 ( .A(n10155), .B(n10329), .ZN(n10161) );
  OR2_X1 U12839 ( .A1(n7219), .A2(n10342), .ZN(n10157) );
  NAND2_X1 U12840 ( .A1(n10340), .A2(n11965), .ZN(n10156) );
  NAND2_X1 U12841 ( .A1(n10157), .A2(n10156), .ZN(n10160) );
  XNOR2_X1 U12842 ( .A(n10161), .B(n10160), .ZN(n11756) );
  NAND2_X1 U12843 ( .A1(n10161), .A2(n10160), .ZN(n10162) );
  NAND2_X1 U12844 ( .A1(n15098), .A2(n10326), .ZN(n10164) );
  NAND2_X1 U12845 ( .A1(n12091), .A2(n10346), .ZN(n10163) );
  NAND2_X1 U12846 ( .A1(n10164), .A2(n10163), .ZN(n10165) );
  XNOR2_X1 U12847 ( .A(n10165), .B(n10329), .ZN(n10174) );
  INV_X1 U12848 ( .A(n10174), .ZN(n12085) );
  OR2_X1 U12849 ( .A1(n12030), .A2(n10342), .ZN(n10167) );
  NAND2_X1 U12850 ( .A1(n10340), .A2(n12091), .ZN(n10166) );
  AND2_X1 U12851 ( .A1(n10167), .A2(n10166), .ZN(n12084) );
  NAND2_X1 U12852 ( .A1(n12085), .A2(n12084), .ZN(n12083) );
  NAND2_X1 U12853 ( .A1(n15795), .A2(n10326), .ZN(n10169) );
  NAND2_X1 U12854 ( .A1(n12028), .A2(n10346), .ZN(n10168) );
  NAND2_X1 U12855 ( .A1(n10169), .A2(n10168), .ZN(n10170) );
  XNOR2_X1 U12856 ( .A(n10170), .B(n11474), .ZN(n12067) );
  INV_X1 U12857 ( .A(n15795), .ZN(n15793) );
  OR2_X1 U12858 ( .A1(n15793), .A2(n10342), .ZN(n10172) );
  NAND2_X1 U12859 ( .A1(n10340), .A2(n12028), .ZN(n10171) );
  NAND2_X1 U12860 ( .A1(n12067), .A2(n12066), .ZN(n10173) );
  AND2_X1 U12861 ( .A1(n12083), .A2(n10173), .ZN(n10179) );
  OAI21_X1 U12862 ( .B1(n12067), .B2(n12066), .A(n12084), .ZN(n10175) );
  NAND2_X1 U12863 ( .A1(n10175), .A2(n10174), .ZN(n10178) );
  INV_X1 U12864 ( .A(n12067), .ZN(n12081) );
  INV_X1 U12865 ( .A(n12066), .ZN(n12080) );
  INV_X1 U12866 ( .A(n12084), .ZN(n10176) );
  NAND3_X1 U12867 ( .A1(n12081), .A2(n12080), .A3(n10176), .ZN(n10177) );
  NAND2_X1 U12868 ( .A1(n15853), .A2(n10346), .ZN(n10181) );
  NAND2_X1 U12869 ( .A1(n15097), .A2(n10326), .ZN(n10180) );
  NAND2_X1 U12870 ( .A1(n10181), .A2(n10180), .ZN(n10182) );
  XNOR2_X1 U12871 ( .A(n10182), .B(n10329), .ZN(n10186) );
  OR2_X1 U12872 ( .A1(n12197), .A2(n10342), .ZN(n10184) );
  NAND2_X1 U12873 ( .A1(n15853), .A2(n10326), .ZN(n10183) );
  NAND2_X1 U12874 ( .A1(n10184), .A2(n10183), .ZN(n10185) );
  XNOR2_X1 U12875 ( .A(n10186), .B(n10185), .ZN(n12179) );
  NAND2_X1 U12876 ( .A1(n10186), .A2(n10185), .ZN(n10187) );
  NAND2_X1 U12877 ( .A1(n15780), .A2(n10346), .ZN(n10189) );
  NAND2_X1 U12878 ( .A1(n15096), .A2(n10326), .ZN(n10188) );
  NAND2_X1 U12879 ( .A1(n10189), .A2(n10188), .ZN(n10190) );
  XNOR2_X1 U12880 ( .A(n10190), .B(n11474), .ZN(n10193) );
  NAND2_X1 U12881 ( .A1(n15780), .A2(n10340), .ZN(n10192) );
  OR2_X1 U12882 ( .A1(n12199), .A2(n10342), .ZN(n10191) );
  NAND2_X1 U12883 ( .A1(n10192), .A2(n10191), .ZN(n10194) );
  XNOR2_X1 U12884 ( .A(n10193), .B(n10194), .ZN(n12146) );
  INV_X1 U12885 ( .A(n10193), .ZN(n10195) );
  NAND2_X1 U12886 ( .A1(n10195), .A2(n10194), .ZN(n10196) );
  NAND2_X1 U12887 ( .A1(n15869), .A2(n10346), .ZN(n10198) );
  NAND2_X1 U12888 ( .A1(n15095), .A2(n10340), .ZN(n10197) );
  NAND2_X1 U12889 ( .A1(n10198), .A2(n10197), .ZN(n10199) );
  XNOR2_X1 U12890 ( .A(n10199), .B(n11474), .ZN(n10204) );
  NOR2_X1 U12891 ( .A1(n12201), .A2(n10342), .ZN(n10200) );
  AOI21_X1 U12892 ( .B1(n15869), .B2(n10326), .A(n10200), .ZN(n10203) );
  XNOR2_X1 U12893 ( .A(n10204), .B(n10203), .ZN(n12410) );
  NAND2_X1 U12894 ( .A1(n10204), .A2(n10203), .ZN(n10205) );
  NAND2_X1 U12895 ( .A1(n15662), .A2(n10346), .ZN(n10207) );
  NAND2_X1 U12896 ( .A1(n15094), .A2(n10326), .ZN(n10206) );
  NAND2_X1 U12897 ( .A1(n10207), .A2(n10206), .ZN(n10208) );
  XNOR2_X1 U12898 ( .A(n10208), .B(n10329), .ZN(n10210) );
  NOR2_X1 U12899 ( .A1(n12413), .A2(n10342), .ZN(n10209) );
  AOI21_X1 U12900 ( .B1(n15662), .B2(n10326), .A(n10209), .ZN(n10211) );
  XNOR2_X1 U12901 ( .A(n10210), .B(n10211), .ZN(n12511) );
  INV_X1 U12902 ( .A(n10210), .ZN(n10212) );
  NAND2_X1 U12903 ( .A1(n12560), .A2(n10346), .ZN(n10214) );
  NAND2_X1 U12904 ( .A1(n15093), .A2(n10326), .ZN(n10213) );
  NAND2_X1 U12905 ( .A1(n10214), .A2(n10213), .ZN(n10215) );
  XNOR2_X1 U12906 ( .A(n10215), .B(n10329), .ZN(n10217) );
  NOR2_X1 U12907 ( .A1(n12904), .A2(n10342), .ZN(n10216) );
  AOI21_X1 U12908 ( .B1(n12560), .B2(n10340), .A(n10216), .ZN(n10218) );
  XNOR2_X1 U12909 ( .A(n10217), .B(n10218), .ZN(n12741) );
  INV_X1 U12910 ( .A(n10217), .ZN(n10219) );
  OR2_X1 U12911 ( .A1(n10219), .A2(n10218), .ZN(n10220) );
  NAND2_X1 U12912 ( .A1(n12902), .A2(n10346), .ZN(n10222) );
  NAND2_X1 U12913 ( .A1(n15092), .A2(n10326), .ZN(n10221) );
  NAND2_X1 U12914 ( .A1(n10222), .A2(n10221), .ZN(n10223) );
  XNOR2_X1 U12915 ( .A(n10223), .B(n11474), .ZN(n10231) );
  INV_X1 U12916 ( .A(n15092), .ZN(n12552) );
  NOR2_X1 U12917 ( .A1(n12552), .A2(n10342), .ZN(n10224) );
  AOI21_X1 U12918 ( .B1(n12902), .B2(n10326), .A(n10224), .ZN(n10230) );
  XNOR2_X1 U12919 ( .A(n10231), .B(n10230), .ZN(n12901) );
  NAND2_X1 U12920 ( .A1(n15651), .A2(n10346), .ZN(n10226) );
  NAND2_X1 U12921 ( .A1(n15520), .A2(n10340), .ZN(n10225) );
  NAND2_X1 U12922 ( .A1(n10226), .A2(n10225), .ZN(n10227) );
  XNOR2_X1 U12923 ( .A(n10227), .B(n10329), .ZN(n10233) );
  INV_X1 U12924 ( .A(n10233), .ZN(n10229) );
  INV_X1 U12925 ( .A(n15520), .ZN(n13025) );
  NOR2_X1 U12926 ( .A1(n13025), .A2(n10342), .ZN(n10228) );
  AOI21_X1 U12927 ( .B1(n15651), .B2(n10340), .A(n10228), .ZN(n10232) );
  NOR2_X1 U12928 ( .A1(n10229), .A2(n10232), .ZN(n10234) );
  NAND2_X1 U12929 ( .A1(n10231), .A2(n10230), .ZN(n14967) );
  XNOR2_X1 U12930 ( .A(n10233), .B(n10232), .ZN(n14971) );
  AND2_X1 U12931 ( .A1(n14967), .A2(n14971), .ZN(n14968) );
  OR2_X1 U12932 ( .A1(n10234), .A2(n14968), .ZN(n15029) );
  NAND2_X1 U12933 ( .A1(n15645), .A2(n10346), .ZN(n10236) );
  NAND2_X1 U12934 ( .A1(n15502), .A2(n10326), .ZN(n10235) );
  NAND2_X1 U12935 ( .A1(n10236), .A2(n10235), .ZN(n10237) );
  XNOR2_X1 U12936 ( .A(n10237), .B(n10329), .ZN(n10240) );
  NOR2_X1 U12937 ( .A1(n13027), .A2(n10342), .ZN(n10238) );
  AOI21_X1 U12938 ( .B1(n15645), .B2(n10340), .A(n10238), .ZN(n10241) );
  XNOR2_X1 U12939 ( .A(n10240), .B(n10241), .ZN(n15032) );
  AND2_X1 U12940 ( .A1(n15029), .A2(n15032), .ZN(n10239) );
  INV_X1 U12941 ( .A(n10240), .ZN(n10242) );
  OR2_X1 U12942 ( .A1(n10242), .A2(n10241), .ZN(n10243) );
  NAND2_X1 U12943 ( .A1(n15639), .A2(n10346), .ZN(n10245) );
  NAND2_X1 U12944 ( .A1(n15091), .A2(n10326), .ZN(n10244) );
  NAND2_X1 U12945 ( .A1(n10245), .A2(n10244), .ZN(n10246) );
  XNOR2_X1 U12946 ( .A(n10246), .B(n11474), .ZN(n10251) );
  NOR2_X1 U12947 ( .A1(n15517), .A2(n10342), .ZN(n10247) );
  AOI21_X1 U12948 ( .B1(n15639), .B2(n10340), .A(n10247), .ZN(n10250) );
  XNOR2_X1 U12949 ( .A(n10251), .B(n10250), .ZN(n14934) );
  INV_X1 U12950 ( .A(n14934), .ZN(n10248) );
  NAND2_X1 U12951 ( .A1(n10251), .A2(n10250), .ZN(n10252) );
  NAND2_X1 U12952 ( .A1(n15633), .A2(n10346), .ZN(n10254) );
  NAND2_X1 U12953 ( .A1(n15501), .A2(n10326), .ZN(n10253) );
  NAND2_X1 U12954 ( .A1(n10254), .A2(n10253), .ZN(n10255) );
  XNOR2_X1 U12955 ( .A(n10255), .B(n11474), .ZN(n14990) );
  NAND2_X1 U12956 ( .A1(n15633), .A2(n10326), .ZN(n10257) );
  NAND2_X1 U12957 ( .A1(n10338), .A2(n15501), .ZN(n10256) );
  NAND2_X1 U12958 ( .A1(n15628), .A2(n10346), .ZN(n10259) );
  NAND2_X1 U12959 ( .A1(n15090), .A2(n10340), .ZN(n10258) );
  NAND2_X1 U12960 ( .A1(n10259), .A2(n10258), .ZN(n10260) );
  XNOR2_X1 U12961 ( .A(n10260), .B(n10329), .ZN(n14986) );
  NAND2_X1 U12962 ( .A1(n15628), .A2(n10326), .ZN(n10262) );
  NAND2_X1 U12963 ( .A1(n15090), .A2(n10338), .ZN(n10261) );
  NAND2_X1 U12964 ( .A1(n10262), .A2(n10261), .ZN(n14985) );
  NAND2_X1 U12965 ( .A1(n14986), .A2(n14985), .ZN(n10265) );
  INV_X1 U12966 ( .A(n10263), .ZN(n10264) );
  NAND2_X1 U12967 ( .A1(n10265), .A2(n14988), .ZN(n10268) );
  INV_X1 U12968 ( .A(n14990), .ZN(n14987) );
  INV_X1 U12969 ( .A(n14986), .ZN(n10267) );
  INV_X1 U12970 ( .A(n14985), .ZN(n10266) );
  NAND2_X1 U12971 ( .A1(n10267), .A2(n10266), .ZN(n14999) );
  OAI21_X1 U12972 ( .B1(n10268), .B2(n14987), .A(n14999), .ZN(n10269) );
  NAND2_X1 U12973 ( .A1(n15622), .A2(n10346), .ZN(n10271) );
  NAND2_X1 U12974 ( .A1(n15089), .A2(n10340), .ZN(n10270) );
  NAND2_X1 U12975 ( .A1(n10271), .A2(n10270), .ZN(n10272) );
  XNOR2_X1 U12976 ( .A(n10272), .B(n10329), .ZN(n10277) );
  AND2_X1 U12977 ( .A1(n15089), .A2(n10338), .ZN(n10273) );
  AOI21_X1 U12978 ( .B1(n15622), .B2(n10326), .A(n10273), .ZN(n10275) );
  XNOR2_X1 U12979 ( .A(n10277), .B(n10275), .ZN(n15000) );
  NAND2_X1 U12980 ( .A1(n10274), .A2(n15000), .ZN(n15003) );
  INV_X1 U12981 ( .A(n10275), .ZN(n10276) );
  OR2_X1 U12982 ( .A1(n10277), .A2(n10276), .ZN(n10278) );
  NAND2_X1 U12983 ( .A1(n15616), .A2(n10346), .ZN(n10280) );
  NAND2_X1 U12984 ( .A1(n15419), .A2(n10326), .ZN(n10279) );
  NAND2_X1 U12985 ( .A1(n10280), .A2(n10279), .ZN(n10281) );
  XNOR2_X1 U12986 ( .A(n10281), .B(n10329), .ZN(n10282) );
  AOI22_X1 U12987 ( .A1(n15616), .A2(n10326), .B1(n10338), .B2(n15419), .ZN(
        n10283) );
  XNOR2_X1 U12988 ( .A(n10282), .B(n10283), .ZN(n15051) );
  INV_X1 U12989 ( .A(n10282), .ZN(n10284) );
  NAND2_X1 U12990 ( .A1(n15605), .A2(n10346), .ZN(n10286) );
  NAND2_X1 U12991 ( .A1(n15088), .A2(n10326), .ZN(n10285) );
  NAND2_X1 U12992 ( .A1(n10286), .A2(n10285), .ZN(n10287) );
  XNOR2_X1 U12993 ( .A(n10287), .B(n10329), .ZN(n10289) );
  AND2_X1 U12994 ( .A1(n15088), .A2(n10338), .ZN(n10288) );
  AOI21_X1 U12995 ( .B1(n15605), .B2(n10340), .A(n10288), .ZN(n10290) );
  XNOR2_X1 U12996 ( .A(n10289), .B(n10290), .ZN(n14950) );
  INV_X1 U12997 ( .A(n10290), .ZN(n10291) );
  NAND2_X1 U12998 ( .A1(n10289), .A2(n10291), .ZN(n10292) );
  AND2_X1 U12999 ( .A1(n15421), .A2(n10338), .ZN(n10293) );
  AOI21_X1 U13000 ( .B1(n15602), .B2(n10340), .A(n10293), .ZN(n10296) );
  AOI22_X1 U13001 ( .A1(n15602), .A2(n10346), .B1(n10340), .B2(n15421), .ZN(
        n10294) );
  XNOR2_X1 U13002 ( .A(n10294), .B(n10329), .ZN(n10295) );
  XOR2_X1 U13003 ( .A(n10296), .B(n10295), .Z(n15020) );
  INV_X1 U13004 ( .A(n10295), .ZN(n10298) );
  INV_X1 U13005 ( .A(n10296), .ZN(n10297) );
  NAND2_X1 U13006 ( .A1(n10298), .A2(n10297), .ZN(n10299) );
  AOI22_X1 U13007 ( .A1(n15597), .A2(n10346), .B1(n10340), .B2(n15363), .ZN(
        n10300) );
  XNOR2_X1 U13008 ( .A(n10300), .B(n10329), .ZN(n10301) );
  AOI22_X1 U13009 ( .A1(n15597), .A2(n10326), .B1(n10338), .B2(n15363), .ZN(
        n10302) );
  XNOR2_X1 U13010 ( .A(n10301), .B(n10302), .ZN(n14960) );
  NAND2_X1 U13011 ( .A1(n10301), .A2(n10302), .ZN(n10303) );
  OAI22_X1 U13012 ( .A1(n15370), .A2(n10348), .B1(n15391), .B2(n10342), .ZN(
        n10305) );
  OAI22_X1 U13013 ( .A1(n15370), .A2(n10151), .B1(n15391), .B2(n10348), .ZN(
        n10304) );
  XNOR2_X1 U13014 ( .A(n10304), .B(n10329), .ZN(n10306) );
  XOR2_X1 U13015 ( .A(n10305), .B(n10306), .Z(n15042) );
  OR2_X1 U13016 ( .A1(n10306), .A2(n10305), .ZN(n10307) );
  NAND2_X1 U13017 ( .A1(n15586), .A2(n10346), .ZN(n10309) );
  NAND2_X1 U13018 ( .A1(n15362), .A2(n10326), .ZN(n10308) );
  NAND2_X1 U13019 ( .A1(n10309), .A2(n10308), .ZN(n10310) );
  XNOR2_X1 U13020 ( .A(n10310), .B(n10329), .ZN(n10311) );
  AOI22_X1 U13021 ( .A1(n15586), .A2(n10326), .B1(n10338), .B2(n15362), .ZN(
        n10312) );
  XNOR2_X1 U13022 ( .A(n10311), .B(n10312), .ZN(n14942) );
  INV_X1 U13023 ( .A(n10311), .ZN(n10313) );
  AOI22_X1 U13024 ( .A1(n15341), .A2(n10326), .B1(n10338), .B2(n15306), .ZN(
        n10317) );
  NAND2_X1 U13025 ( .A1(n15341), .A2(n10346), .ZN(n10315) );
  NAND2_X1 U13026 ( .A1(n15306), .A2(n10326), .ZN(n10314) );
  NAND2_X1 U13027 ( .A1(n10315), .A2(n10314), .ZN(n10316) );
  XNOR2_X1 U13028 ( .A(n10316), .B(n10329), .ZN(n10319) );
  XOR2_X1 U13029 ( .A(n10317), .B(n10319), .Z(n15012) );
  INV_X1 U13030 ( .A(n10317), .ZN(n10318) );
  NAND2_X1 U13031 ( .A1(n15318), .A2(n10346), .ZN(n10321) );
  NAND2_X1 U13032 ( .A1(n15330), .A2(n10326), .ZN(n10320) );
  NAND2_X1 U13033 ( .A1(n10321), .A2(n10320), .ZN(n10322) );
  XNOR2_X1 U13034 ( .A(n10322), .B(n10329), .ZN(n10323) );
  AOI22_X1 U13035 ( .A1(n15318), .A2(n10326), .B1(n10338), .B2(n15330), .ZN(
        n10324) );
  XNOR2_X1 U13036 ( .A(n10323), .B(n10324), .ZN(n14980) );
  INV_X1 U13037 ( .A(n10323), .ZN(n10325) );
  AOI22_X1 U13038 ( .A1(n15301), .A2(n10326), .B1(n10338), .B2(n15086), .ZN(
        n10331) );
  NAND2_X1 U13039 ( .A1(n15301), .A2(n10346), .ZN(n10328) );
  NAND2_X1 U13040 ( .A1(n15086), .A2(n10340), .ZN(n10327) );
  NAND2_X1 U13041 ( .A1(n10328), .A2(n10327), .ZN(n10330) );
  XNOR2_X1 U13042 ( .A(n10330), .B(n10329), .ZN(n10333) );
  XOR2_X1 U13043 ( .A(n10331), .B(n10333), .Z(n15060) );
  INV_X1 U13044 ( .A(n10331), .ZN(n10332) );
  NAND2_X1 U13045 ( .A1(n7122), .A2(n10346), .ZN(n10336) );
  NAND2_X1 U13046 ( .A1(n15297), .A2(n10340), .ZN(n10335) );
  NAND2_X1 U13047 ( .A1(n10336), .A2(n10335), .ZN(n10337) );
  XNOR2_X1 U13048 ( .A(n10337), .B(n11474), .ZN(n10352) );
  AND2_X1 U13049 ( .A1(n15297), .A2(n10338), .ZN(n10339) );
  AOI21_X1 U13050 ( .B1(n7122), .B2(n10340), .A(n10339), .ZN(n10351) );
  XNOR2_X1 U13051 ( .A(n10352), .B(n10351), .ZN(n14922) );
  INV_X1 U13052 ( .A(n10374), .ZN(n10372) );
  NAND2_X1 U13053 ( .A1(n15553), .A2(n10340), .ZN(n10344) );
  OR2_X1 U13054 ( .A1(n14927), .A2(n10342), .ZN(n10343) );
  NAND2_X1 U13055 ( .A1(n10344), .A2(n10343), .ZN(n10345) );
  XNOR2_X1 U13056 ( .A(n10345), .B(n11474), .ZN(n10350) );
  NAND2_X1 U13057 ( .A1(n15553), .A2(n10346), .ZN(n10347) );
  OAI21_X1 U13058 ( .B1(n14927), .B2(n10348), .A(n10347), .ZN(n10349) );
  XNOR2_X1 U13059 ( .A(n10350), .B(n10349), .ZN(n10373) );
  INV_X1 U13060 ( .A(n10373), .ZN(n10385) );
  NAND2_X1 U13061 ( .A1(n10352), .A2(n10351), .ZN(n10384) );
  NAND2_X1 U13062 ( .A1(n10353), .A2(n12140), .ZN(n15824) );
  NAND2_X1 U13063 ( .A1(n12794), .A2(P1_B_REG_SCAN_IN), .ZN(n10354) );
  MUX2_X1 U13064 ( .A(P1_B_REG_SCAN_IN), .B(n10354), .S(n12579), .Z(n10355) );
  INV_X1 U13065 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n10686) );
  AND2_X1 U13066 ( .A1(n15704), .A2(n12794), .ZN(n10685) );
  NOR4_X1 U13067 ( .A1(P1_D_REG_13__SCAN_IN), .A2(P1_D_REG_15__SCAN_IN), .A3(
        P1_D_REG_17__SCAN_IN), .A4(P1_D_REG_18__SCAN_IN), .ZN(n10360) );
  NOR4_X1 U13068 ( .A1(P1_D_REG_9__SCAN_IN), .A2(P1_D_REG_11__SCAN_IN), .A3(
        P1_D_REG_14__SCAN_IN), .A4(P1_D_REG_12__SCAN_IN), .ZN(n10359) );
  NOR4_X1 U13069 ( .A1(P1_D_REG_24__SCAN_IN), .A2(P1_D_REG_25__SCAN_IN), .A3(
        P1_D_REG_26__SCAN_IN), .A4(P1_D_REG_28__SCAN_IN), .ZN(n10358) );
  NOR4_X1 U13070 ( .A1(P1_D_REG_19__SCAN_IN), .A2(P1_D_REG_23__SCAN_IN), .A3(
        P1_D_REG_20__SCAN_IN), .A4(P1_D_REG_22__SCAN_IN), .ZN(n10357) );
  NAND4_X1 U13071 ( .A1(n10360), .A2(n10359), .A3(n10358), .A4(n10357), .ZN(
        n10365) );
  NOR2_X1 U13072 ( .A1(P1_D_REG_27__SCAN_IN), .A2(P1_D_REG_21__SCAN_IN), .ZN(
        n10800) );
  NOR4_X1 U13073 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_31__SCAN_IN), .A3(
        P1_D_REG_16__SCAN_IN), .A4(P1_D_REG_30__SCAN_IN), .ZN(n10363) );
  NOR4_X1 U13074 ( .A1(P1_D_REG_5__SCAN_IN), .A2(P1_D_REG_6__SCAN_IN), .A3(
        P1_D_REG_7__SCAN_IN), .A4(P1_D_REG_8__SCAN_IN), .ZN(n10362) );
  NOR4_X1 U13075 ( .A1(P1_D_REG_10__SCAN_IN), .A2(P1_D_REG_2__SCAN_IN), .A3(
        P1_D_REG_3__SCAN_IN), .A4(P1_D_REG_4__SCAN_IN), .ZN(n10361) );
  NAND4_X1 U13076 ( .A1(n10800), .A2(n10363), .A3(n10362), .A4(n10361), .ZN(
        n10364) );
  NOR2_X1 U13077 ( .A1(n10365), .A2(n10364), .ZN(n11463) );
  NAND2_X1 U13078 ( .A1(n11463), .A2(P1_D_REG_0__SCAN_IN), .ZN(n10366) );
  NAND2_X1 U13079 ( .A1(n15704), .A2(n12579), .ZN(n11466) );
  INV_X1 U13080 ( .A(n11466), .ZN(n10688) );
  AOI21_X1 U13081 ( .B1(n10367), .B2(n10366), .A(n10688), .ZN(n10376) );
  NAND2_X1 U13082 ( .A1(n11827), .A2(n10376), .ZN(n10375) );
  INV_X1 U13083 ( .A(n10375), .ZN(n10369) );
  NOR2_X1 U13084 ( .A1(n11830), .A2(n10719), .ZN(n10368) );
  NOR2_X1 U13085 ( .A1(n10373), .A2(n10370), .ZN(n10371) );
  NAND2_X1 U13086 ( .A1(n10372), .A2(n10371), .ZN(n10390) );
  NAND3_X1 U13087 ( .A1(n10374), .A2(n15072), .A3(n10373), .ZN(n10389) );
  NAND2_X1 U13088 ( .A1(n10375), .A2(n11829), .ZN(n10380) );
  AND2_X1 U13089 ( .A1(n10380), .A2(n10684), .ZN(n12910) );
  INV_X1 U13090 ( .A(n10376), .ZN(n10377) );
  NOR2_X1 U13091 ( .A1(n11465), .A2(n10377), .ZN(n11494) );
  AND2_X1 U13092 ( .A1(n11494), .A2(n11827), .ZN(n15080) );
  INV_X1 U13093 ( .A(n10719), .ZN(n10378) );
  INV_X1 U13094 ( .A(n15065), .ZN(n15053) );
  AOI22_X1 U13095 ( .A1(n15272), .A2(n15053), .B1(P1_REG3_REG_28__SCAN_IN), 
        .B2(P1_U3086), .ZN(n10383) );
  AND2_X1 U13096 ( .A1(n11352), .A2(n10607), .ZN(n10379) );
  AOI21_X1 U13097 ( .B1(n10380), .B2(n10379), .A(P1_U3086), .ZN(n10381) );
  NAND2_X1 U13098 ( .A1(n15281), .A2(n15061), .ZN(n10382) );
  OAI211_X1 U13099 ( .C1(n15066), .C2(n15056), .A(n10383), .B(n10382), .ZN(
        n10387) );
  NOR3_X1 U13100 ( .A1(n10385), .A2(n15070), .A3(n10384), .ZN(n10386) );
  AOI211_X1 U13101 ( .C1(n15068), .C2(n15553), .A(n10387), .B(n10386), .ZN(
        n10388) );
  NAND3_X1 U13102 ( .A1(n10390), .A2(n10389), .A3(n10388), .ZN(P1_U3220) );
  NAND2_X1 U13103 ( .A1(n14902), .A2(n13125), .ZN(n10394) );
  NAND2_X1 U13104 ( .A1(n13126), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n10393) );
  NAND2_X1 U13105 ( .A1(n14383), .A2(n14105), .ZN(n12153) );
  NAND2_X1 U13106 ( .A1(n10420), .A2(n12153), .ZN(n10399) );
  NAND2_X1 U13107 ( .A1(n6548), .A2(n10399), .ZN(n14742) );
  AOI21_X1 U13108 ( .B1(n14744), .B2(n6611), .A(n14717), .ZN(n10401) );
  INV_X1 U13109 ( .A(n14744), .ZN(n14272) );
  AND2_X1 U13110 ( .A1(n7517), .A2(n7740), .ZN(n14321) );
  AND2_X1 U13111 ( .A1(n14379), .A2(n14321), .ZN(n10558) );
  INV_X1 U13112 ( .A(n10402), .ZN(n10403) );
  AOI22_X1 U13113 ( .A1(n10403), .A2(n14713), .B1(P2_REG2_REG_29__SCAN_IN), 
        .B2(n14738), .ZN(n10404) );
  OAI21_X1 U13114 ( .B1(n14272), .B2(n14698), .A(n10404), .ZN(n10405) );
  AOI21_X1 U13115 ( .B1(n14743), .B2(n14703), .A(n10405), .ZN(n10419) );
  NAND2_X1 U13116 ( .A1(n12988), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n10408) );
  NAND2_X1 U13117 ( .A1(n8643), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n10407) );
  NAND2_X1 U13118 ( .A1(n12989), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n10406) );
  AND3_X1 U13119 ( .A1(n10408), .A2(n10407), .A3(n10406), .ZN(n14326) );
  INV_X1 U13120 ( .A(P2_B_REG_SCAN_IN), .ZN(n14378) );
  OR2_X1 U13121 ( .A1(n14912), .A2(n14378), .ZN(n10409) );
  NAND2_X1 U13122 ( .A1(n14086), .A2(n10409), .ZN(n12993) );
  INV_X1 U13123 ( .A(n14363), .ZN(n10416) );
  NAND4_X1 U13124 ( .A1(n10416), .A2(n14853), .A3(n14394), .A4(n14675), .ZN(
        n10411) );
  NAND2_X1 U13125 ( .A1(n14394), .A2(n14376), .ZN(n10410) );
  OAI211_X1 U13126 ( .C1(n14326), .C2(n12993), .A(n10411), .B(n10410), .ZN(
        n10412) );
  OAI21_X1 U13127 ( .B1(n10418), .B2(n10414), .A(n10413), .ZN(n10415) );
  AOI211_X1 U13128 ( .C1(n14853), .C2(n14394), .A(n8640), .B(n10416), .ZN(
        n10417) );
  NAND3_X1 U13129 ( .A1(n7973), .A2(n10419), .A3(n7972), .ZN(P2_U3236) );
  NAND2_X1 U13130 ( .A1(n8040), .A2(n13111), .ZN(n10427) );
  XNOR2_X1 U13131 ( .A(n10436), .B(n14114), .ZN(n10426) );
  INV_X1 U13132 ( .A(n10426), .ZN(n10421) );
  AND2_X1 U13133 ( .A1(n10427), .A2(n10421), .ZN(n11447) );
  NAND2_X1 U13134 ( .A1(n14420), .A2(n13111), .ZN(n10424) );
  INV_X1 U13135 ( .A(n10424), .ZN(n10423) );
  INV_X1 U13136 ( .A(n10425), .ZN(n10422) );
  NAND2_X1 U13137 ( .A1(n10423), .A2(n10422), .ZN(n11448) );
  AND2_X1 U13138 ( .A1(n10425), .A2(n10424), .ZN(n11566) );
  AOI21_X1 U13139 ( .B1(n11447), .B2(n11448), .A(n11566), .ZN(n10431) );
  XNOR2_X1 U13140 ( .A(n10427), .B(n10426), .ZN(n11513) );
  NAND2_X1 U13141 ( .A1(n14733), .A2(n14108), .ZN(n10428) );
  NAND2_X1 U13142 ( .A1(n7985), .A2(n10429), .ZN(n11512) );
  NAND2_X1 U13143 ( .A1(n14419), .A2(n13111), .ZN(n10432) );
  XNOR2_X1 U13144 ( .A(n10432), .B(n10433), .ZN(n11568) );
  INV_X1 U13145 ( .A(n10432), .ZN(n10434) );
  NAND2_X1 U13146 ( .A1(n10434), .A2(n10433), .ZN(n10435) );
  XNOR2_X1 U13147 ( .A(n14136), .B(n13112), .ZN(n10438) );
  NAND2_X1 U13148 ( .A1(n14418), .A2(n13111), .ZN(n10437) );
  NAND2_X1 U13149 ( .A1(n10438), .A2(n10437), .ZN(n10443) );
  INV_X1 U13150 ( .A(n10437), .ZN(n10440) );
  INV_X1 U13151 ( .A(n10438), .ZN(n10439) );
  NAND2_X1 U13152 ( .A1(n10440), .A2(n10439), .ZN(n10441) );
  NAND2_X1 U13153 ( .A1(n10443), .A2(n10441), .ZN(n11618) );
  INV_X1 U13154 ( .A(n11618), .ZN(n10442) );
  XNOR2_X1 U13155 ( .A(n15983), .B(n13112), .ZN(n10445) );
  NAND2_X1 U13156 ( .A1(n14417), .A2(n13111), .ZN(n10444) );
  NAND2_X1 U13157 ( .A1(n10445), .A2(n10444), .ZN(n10449) );
  INV_X1 U13158 ( .A(n10444), .ZN(n10447) );
  INV_X1 U13159 ( .A(n10445), .ZN(n10446) );
  NAND2_X1 U13160 ( .A1(n10447), .A2(n10446), .ZN(n10448) );
  AND2_X1 U13161 ( .A1(n10449), .A2(n10448), .ZN(n11741) );
  XNOR2_X1 U13162 ( .A(n14148), .B(n13112), .ZN(n10450) );
  NAND2_X1 U13163 ( .A1(n14416), .A2(n13111), .ZN(n10451) );
  XNOR2_X1 U13164 ( .A(n10450), .B(n10451), .ZN(n11761) );
  INV_X1 U13165 ( .A(n10450), .ZN(n10453) );
  INV_X1 U13166 ( .A(n10451), .ZN(n10452) );
  NAND2_X1 U13167 ( .A1(n14415), .A2(n13111), .ZN(n10454) );
  XNOR2_X1 U13168 ( .A(n10456), .B(n10454), .ZN(n11979) );
  INV_X1 U13169 ( .A(n10454), .ZN(n10455) );
  NAND2_X1 U13170 ( .A1(n10456), .A2(n10455), .ZN(n10457) );
  XNOR2_X1 U13171 ( .A(n14154), .B(n13112), .ZN(n10458) );
  NAND2_X1 U13172 ( .A1(n14414), .A2(n13111), .ZN(n10459) );
  NAND2_X1 U13173 ( .A1(n10458), .A2(n10459), .ZN(n10464) );
  INV_X1 U13174 ( .A(n10458), .ZN(n10461) );
  INV_X1 U13175 ( .A(n10459), .ZN(n10460) );
  NAND2_X1 U13176 ( .A1(n10461), .A2(n10460), .ZN(n10462) );
  NAND2_X1 U13177 ( .A1(n10464), .A2(n10462), .ZN(n12300) );
  XNOR2_X1 U13178 ( .A(n14159), .B(n13112), .ZN(n10465) );
  NAND2_X1 U13179 ( .A1(n14413), .A2(n13111), .ZN(n10466) );
  NAND2_X1 U13180 ( .A1(n10465), .A2(n10466), .ZN(n10470) );
  INV_X1 U13181 ( .A(n10465), .ZN(n10468) );
  INV_X1 U13182 ( .A(n10466), .ZN(n10467) );
  NAND2_X1 U13183 ( .A1(n10468), .A2(n10467), .ZN(n10469) );
  AND2_X1 U13184 ( .A1(n10470), .A2(n10469), .ZN(n12428) );
  XNOR2_X1 U13185 ( .A(n14842), .B(n13112), .ZN(n10472) );
  NAND2_X1 U13186 ( .A1(n14412), .A2(n13111), .ZN(n10471) );
  XNOR2_X1 U13187 ( .A(n10472), .B(n10471), .ZN(n12819) );
  XNOR2_X1 U13188 ( .A(n14171), .B(n13112), .ZN(n10473) );
  NAND2_X1 U13189 ( .A1(n14411), .A2(n13111), .ZN(n10474) );
  NAND2_X1 U13190 ( .A1(n10473), .A2(n10474), .ZN(n10478) );
  INV_X1 U13191 ( .A(n10473), .ZN(n10476) );
  INV_X1 U13192 ( .A(n10474), .ZN(n10475) );
  NAND2_X1 U13193 ( .A1(n10476), .A2(n10475), .ZN(n10477) );
  NAND2_X1 U13194 ( .A1(n10478), .A2(n10477), .ZN(n12869) );
  NAND2_X1 U13195 ( .A1(n12867), .A2(n10478), .ZN(n12890) );
  XNOR2_X1 U13196 ( .A(n14829), .B(n13112), .ZN(n10479) );
  NAND2_X1 U13197 ( .A1(n14410), .A2(n13111), .ZN(n10480) );
  NAND2_X1 U13198 ( .A1(n10479), .A2(n10480), .ZN(n10484) );
  INV_X1 U13199 ( .A(n10479), .ZN(n10482) );
  INV_X1 U13200 ( .A(n10480), .ZN(n10481) );
  NAND2_X1 U13201 ( .A1(n10482), .A2(n10481), .ZN(n10483) );
  AND2_X1 U13202 ( .A1(n10484), .A2(n10483), .ZN(n12891) );
  XNOR2_X1 U13203 ( .A(n14191), .B(n13112), .ZN(n10487) );
  NAND2_X1 U13204 ( .A1(n14409), .A2(n13111), .ZN(n10488) );
  XNOR2_X1 U13205 ( .A(n10487), .B(n10488), .ZN(n13973) );
  NAND2_X1 U13206 ( .A1(n14408), .A2(n13111), .ZN(n10485) );
  INV_X1 U13207 ( .A(n10486), .ZN(n10491) );
  OR2_X1 U13208 ( .A1(n13973), .A2(n10491), .ZN(n10492) );
  INV_X1 U13209 ( .A(n10487), .ZN(n10490) );
  INV_X1 U13210 ( .A(n10488), .ZN(n10489) );
  NAND2_X1 U13211 ( .A1(n10490), .A2(n10489), .ZN(n13975) );
  AND2_X1 U13212 ( .A1(n13980), .A2(n13975), .ZN(n13976) );
  XNOR2_X1 U13213 ( .A(n14817), .B(n13112), .ZN(n14028) );
  XNOR2_X1 U13214 ( .A(n14809), .B(n13112), .ZN(n10496) );
  NAND2_X1 U13215 ( .A1(n14406), .A2(n13111), .ZN(n10497) );
  NAND2_X1 U13216 ( .A1(n10496), .A2(n10497), .ZN(n10493) );
  INV_X1 U13217 ( .A(n10493), .ZN(n14026) );
  AND2_X1 U13218 ( .A1(n14407), .A2(n13111), .ZN(n14093) );
  NAND2_X1 U13219 ( .A1(n10493), .A2(n14093), .ZN(n10495) );
  OAI21_X1 U13220 ( .B1(n14028), .B2(n14026), .A(n10495), .ZN(n10494) );
  INV_X1 U13221 ( .A(n10495), .ZN(n10500) );
  INV_X1 U13222 ( .A(n14028), .ZN(n14029) );
  INV_X1 U13223 ( .A(n10496), .ZN(n10499) );
  INV_X1 U13224 ( .A(n10497), .ZN(n10498) );
  AND2_X1 U13225 ( .A1(n10499), .A2(n10498), .ZN(n14025) );
  AOI21_X1 U13226 ( .B1(n10500), .B2(n14029), .A(n14025), .ZN(n10501) );
  XNOR2_X1 U13227 ( .A(n14697), .B(n13112), .ZN(n10502) );
  NAND2_X1 U13228 ( .A1(n14405), .A2(n13111), .ZN(n10503) );
  NAND2_X1 U13229 ( .A1(n10502), .A2(n10503), .ZN(n10509) );
  INV_X1 U13230 ( .A(n10502), .ZN(n10505) );
  INV_X1 U13231 ( .A(n10503), .ZN(n10504) );
  NAND2_X1 U13232 ( .A1(n10505), .A2(n10504), .ZN(n10506) );
  NAND2_X1 U13233 ( .A1(n10509), .A2(n10506), .ZN(n14040) );
  NAND2_X1 U13234 ( .A1(n14404), .A2(n13111), .ZN(n10510) );
  NAND2_X1 U13235 ( .A1(n14403), .A2(n13111), .ZN(n10513) );
  INV_X1 U13236 ( .A(n10512), .ZN(n10515) );
  INV_X1 U13237 ( .A(n10513), .ZN(n10514) );
  NAND2_X1 U13238 ( .A1(n10515), .A2(n10514), .ZN(n14001) );
  XNOR2_X1 U13239 ( .A(n14790), .B(n13112), .ZN(n10518) );
  NAND2_X1 U13240 ( .A1(n14402), .A2(n13111), .ZN(n10517) );
  XNOR2_X1 U13241 ( .A(n10518), .B(n10517), .ZN(n14058) );
  INV_X1 U13242 ( .A(n14058), .ZN(n10516) );
  NAND2_X1 U13243 ( .A1(n10518), .A2(n10517), .ZN(n10519) );
  NAND2_X1 U13244 ( .A1(n14401), .A2(n13111), .ZN(n10520) );
  XNOR2_X1 U13245 ( .A(n10522), .B(n10520), .ZN(n14010) );
  INV_X1 U13246 ( .A(n10520), .ZN(n10521) );
  NAND2_X1 U13247 ( .A1(n10522), .A2(n10521), .ZN(n10523) );
  XNOR2_X1 U13248 ( .A(n14618), .B(n13112), .ZN(n10525) );
  XNOR2_X1 U13249 ( .A(n14600), .B(n13112), .ZN(n13992) );
  NAND2_X1 U13250 ( .A1(n14400), .A2(n13111), .ZN(n14063) );
  AOI21_X1 U13251 ( .B1(n13992), .B2(n14254), .A(n14063), .ZN(n10524) );
  NAND2_X1 U13252 ( .A1(n13988), .A2(n10524), .ZN(n10533) );
  INV_X1 U13253 ( .A(n10525), .ZN(n10526) );
  AND2_X1 U13254 ( .A1(n14399), .A2(n13111), .ZN(n10528) );
  INV_X1 U13255 ( .A(n10528), .ZN(n13991) );
  NAND2_X1 U13256 ( .A1(n13992), .A2(n13991), .ZN(n10531) );
  INV_X1 U13257 ( .A(n13992), .ZN(n10529) );
  AND2_X1 U13258 ( .A1(n10529), .A2(n10528), .ZN(n10530) );
  NAND2_X1 U13259 ( .A1(n10533), .A2(n10532), .ZN(n14048) );
  AND2_X1 U13260 ( .A1(n14398), .A2(n13111), .ZN(n10535) );
  NAND2_X1 U13261 ( .A1(n10534), .A2(n10535), .ZN(n10539) );
  INV_X1 U13262 ( .A(n10534), .ZN(n10537) );
  INV_X1 U13263 ( .A(n10535), .ZN(n10536) );
  NAND2_X1 U13264 ( .A1(n10537), .A2(n10536), .ZN(n10538) );
  AND2_X1 U13265 ( .A1(n10539), .A2(n10538), .ZN(n14047) );
  AND2_X1 U13266 ( .A1(n14397), .A2(n13111), .ZN(n10541) );
  NAND2_X1 U13267 ( .A1(n10540), .A2(n10541), .ZN(n10545) );
  INV_X1 U13268 ( .A(n10540), .ZN(n10543) );
  INV_X1 U13269 ( .A(n10541), .ZN(n10542) );
  NAND2_X1 U13270 ( .A1(n10543), .A2(n10542), .ZN(n10544) );
  XNOR2_X1 U13271 ( .A(n14549), .B(n13112), .ZN(n10547) );
  NAND2_X1 U13272 ( .A1(n14396), .A2(n13111), .ZN(n10546) );
  XNOR2_X1 U13273 ( .A(n10547), .B(n10546), .ZN(n14084) );
  AND2_X1 U13274 ( .A1(n14395), .A2(n13111), .ZN(n10549) );
  NAND2_X1 U13275 ( .A1(n10548), .A2(n10549), .ZN(n13119) );
  INV_X1 U13276 ( .A(n10548), .ZN(n10551) );
  INV_X1 U13277 ( .A(n10549), .ZN(n10550) );
  NAND2_X1 U13278 ( .A1(n10551), .A2(n10550), .ZN(n10552) );
  NAND2_X1 U13279 ( .A1(n13119), .A2(n10552), .ZN(n10553) );
  OR2_X1 U13280 ( .A1(n15980), .A2(n11633), .ZN(n10564) );
  AND2_X1 U13281 ( .A1(n15989), .A2(n11147), .ZN(n10555) );
  AOI22_X1 U13282 ( .A1(n14394), .A2(n14086), .B1(n14376), .B2(n14396), .ZN(
        n14528) );
  INV_X1 U13283 ( .A(n10557), .ZN(n14375) );
  NAND2_X1 U13284 ( .A1(n10559), .A2(n10558), .ZN(n10560) );
  NAND2_X1 U13285 ( .A1(n14749), .A2(n14101), .ZN(n10570) );
  INV_X1 U13286 ( .A(n10561), .ZN(n10563) );
  OAI21_X1 U13287 ( .B1(n10564), .B2(n10563), .A(n10562), .ZN(n10568) );
  AND2_X1 U13288 ( .A1(n10566), .A2(n10565), .ZN(n10567) );
  NAND2_X1 U13289 ( .A1(n10568), .A2(n10567), .ZN(n11356) );
  AOI22_X1 U13290 ( .A1(n14532), .A2(n14088), .B1(P2_REG3_REG_27__SCAN_IN), 
        .B2(P2_U3088), .ZN(n10569) );
  OAI211_X1 U13291 ( .C1(n14528), .C2(n14090), .A(n10570), .B(n10569), .ZN(
        n10571) );
  INV_X1 U13292 ( .A(n10571), .ZN(n10572) );
  NAND2_X1 U13293 ( .A1(n10575), .A2(n10574), .ZN(n10576) );
  XNOR2_X1 U13294 ( .A(n10576), .B(n13469), .ZN(n13655) );
  NAND3_X1 U13295 ( .A1(n10579), .A2(n16044), .A3(n10578), .ZN(n10582) );
  INV_X1 U13296 ( .A(n13145), .ZN(n13832) );
  INV_X1 U13297 ( .A(P3_REG0_REG_28__SCAN_IN), .ZN(n10583) );
  NAND2_X1 U13298 ( .A1(n10586), .A2(n10585), .ZN(P3_U3455) );
  NAND2_X1 U13299 ( .A1(n12320), .A2(P2_STATE_REG_SCAN_IN), .ZN(n10587) );
  INV_X1 U13300 ( .A(n10588), .ZN(n10591) );
  NAND3_X1 U13301 ( .A1(n12051), .A2(n10589), .A3(n7196), .ZN(n10590) );
  AOI21_X1 U13302 ( .B1(n10591), .B2(n10590), .A(n16014), .ZN(n10605) );
  OR3_X1 U13303 ( .A1(n10593), .A2(n12048), .A3(n10592), .ZN(n10594) );
  AOI21_X1 U13304 ( .B1(n10595), .B2(n10594), .A(n16015), .ZN(n10604) );
  INV_X1 U13305 ( .A(n10596), .ZN(n10597) );
  NAND3_X1 U13306 ( .A1(n12058), .A2(n10598), .A3(n10597), .ZN(n10599) );
  AOI21_X1 U13307 ( .B1(n10600), .B2(n10599), .A(n16013), .ZN(n10603) );
  AND2_X1 U13308 ( .A1(P3_U3151), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n12490) );
  AOI21_X1 U13309 ( .B1(n16012), .B2(P3_ADDR_REG_10__SCAN_IN), .A(n12490), 
        .ZN(n10601) );
  OAI21_X1 U13310 ( .B1(n13617), .B2(n10671), .A(n10601), .ZN(n10602) );
  OR4_X1 U13311 ( .A1(n10605), .A2(n10604), .A3(n10603), .A4(n10602), .ZN(
        P3_U3192) );
  INV_X1 U13312 ( .A(n10687), .ZN(n10606) );
  INV_X1 U13313 ( .A(n10614), .ZN(n10610) );
  XNOR2_X1 U13314 ( .A(n10615), .B(n10610), .ZN(n10619) );
  XNOR2_X1 U13315 ( .A(n10619), .B(P2_ADDR_REG_1__SCAN_IN), .ZN(n10612) );
  INV_X1 U13316 ( .A(P3_ADDR_REG_0__SCAN_IN), .ZN(n10608) );
  NAND2_X1 U13317 ( .A1(n10608), .A2(P1_ADDR_REG_0__SCAN_IN), .ZN(n10609) );
  NAND2_X1 U13318 ( .A1(n10610), .A2(n10609), .ZN(n15708) );
  AND2_X1 U13319 ( .A1(n15708), .A2(P2_ADDR_REG_0__SCAN_IN), .ZN(n10611) );
  NAND2_X1 U13320 ( .A1(n10612), .A2(n10611), .ZN(n10622) );
  OAI21_X1 U13321 ( .B1(n10612), .B2(n10611), .A(n10622), .ZN(n10613) );
  INV_X1 U13322 ( .A(n10613), .ZN(SUB_1596_U5) );
  NAND2_X1 U13323 ( .A1(n10615), .A2(n10614), .ZN(n10617) );
  NAND2_X1 U13324 ( .A1(n15101), .A2(P3_ADDR_REG_1__SCAN_IN), .ZN(n10616) );
  NAND2_X1 U13325 ( .A1(n10617), .A2(n10616), .ZN(n10625) );
  NAND2_X1 U13326 ( .A1(n15122), .A2(P3_ADDR_REG_2__SCAN_IN), .ZN(n10626) );
  NAND2_X1 U13327 ( .A1(n11307), .A2(P1_ADDR_REG_2__SCAN_IN), .ZN(n10618) );
  XNOR2_X1 U13328 ( .A(n10625), .B(n10624), .ZN(n10630) );
  INV_X1 U13329 ( .A(n10630), .ZN(n10633) );
  INV_X1 U13330 ( .A(P2_ADDR_REG_2__SCAN_IN), .ZN(n10970) );
  XNOR2_X1 U13331 ( .A(n10633), .B(n10970), .ZN(n10623) );
  INV_X1 U13332 ( .A(n10619), .ZN(n10620) );
  NAND2_X1 U13333 ( .A1(n10620), .A2(P2_ADDR_REG_1__SCAN_IN), .ZN(n10621) );
  NAND2_X1 U13334 ( .A1(n10622), .A2(n10621), .ZN(n10632) );
  XNOR2_X1 U13335 ( .A(n10623), .B(n10632), .ZN(SUB_1596_U61) );
  NAND2_X1 U13336 ( .A1(n10627), .A2(P3_ADDR_REG_3__SCAN_IN), .ZN(n10646) );
  INV_X1 U13337 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n10629) );
  XNOR2_X1 U13338 ( .A(n10647), .B(n10629), .ZN(n10642) );
  XNOR2_X1 U13339 ( .A(n10642), .B(P2_ADDR_REG_3__SCAN_IN), .ZN(n10636) );
  AND2_X1 U13340 ( .A1(n10630), .A2(P2_ADDR_REG_2__SCAN_IN), .ZN(n10631) );
  OR2_X1 U13341 ( .A1(n10632), .A2(n10631), .ZN(n10635) );
  NAND2_X1 U13342 ( .A1(n10633), .A2(n10970), .ZN(n10634) );
  NAND2_X1 U13343 ( .A1(n10635), .A2(n10634), .ZN(n10643) );
  XNOR2_X1 U13344 ( .A(n10636), .B(n10643), .ZN(SUB_1596_U60) );
  NAND2_X1 U13345 ( .A1(n10696), .A2(P1_U3086), .ZN(n15700) );
  INV_X1 U13346 ( .A(n15136), .ZN(n10638) );
  OAI222_X1 U13347 ( .A1(n15700), .A2(n10639), .B1(n15703), .B2(n7802), .C1(
        n10638), .C2(P1_U3086), .ZN(P1_U3352) );
  NAND2_X1 U13348 ( .A1(n10696), .A2(P3_U3151), .ZN(n13970) );
  NOR2_X1 U13349 ( .A1(n10696), .A2(P3_STATE_REG_SCAN_IN), .ZN(n13966) );
  INV_X2 U13350 ( .A(n13966), .ZN(n13102) );
  OAI222_X1 U13351 ( .A1(P3_U3151), .A2(n11703), .B1(n13970), .B2(n10641), 
        .C1(n13102), .C2(n10640), .ZN(P3_U3287) );
  INV_X1 U13352 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n14422) );
  OAI21_X1 U13353 ( .B1(n10643), .B2(n14422), .A(n10642), .ZN(n10645) );
  NAND2_X1 U13354 ( .A1(n10643), .A2(n14422), .ZN(n10644) );
  AND2_X1 U13355 ( .A1(n10645), .A2(n10644), .ZN(n10652) );
  NAND2_X1 U13356 ( .A1(n10648), .A2(P1_ADDR_REG_4__SCAN_IN), .ZN(n10649) );
  INV_X1 U13357 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n10650) );
  NAND2_X1 U13358 ( .A1(n10651), .A2(n10652), .ZN(n10681) );
  OAI21_X1 U13359 ( .B1(n10652), .B2(n10651), .A(n10681), .ZN(n10653) );
  INV_X1 U13360 ( .A(n10653), .ZN(SUB_1596_U59) );
  INV_X1 U13361 ( .A(n10654), .ZN(n10709) );
  INV_X1 U13362 ( .A(n11079), .ZN(n15146) );
  OAI222_X1 U13363 ( .A1(n15700), .A2(n10655), .B1(n15703), .B2(n10709), .C1(
        n15146), .C2(P1_U3086), .ZN(P1_U3351) );
  OAI222_X1 U13364 ( .A1(P1_U3086), .A2(n9482), .B1(n15703), .B2(n10751), .C1(
        n10656), .C2(n15700), .ZN(P1_U3354) );
  CLKBUF_X1 U13365 ( .A(n13970), .Z(n13962) );
  INV_X1 U13366 ( .A(SI_5_), .ZN(n10659) );
  INV_X1 U13367 ( .A(n10657), .ZN(n10658) );
  OAI222_X1 U13368 ( .A1(P3_U3151), .A2(n7646), .B1(n13962), .B2(n10659), .C1(
        n13102), .C2(n10658), .ZN(P3_U3290) );
  INV_X1 U13369 ( .A(SI_4_), .ZN(n10821) );
  INV_X1 U13370 ( .A(n10660), .ZN(n10661) );
  OAI222_X1 U13371 ( .A1(P3_U3151), .A2(n10662), .B1(n13962), .B2(n10821), 
        .C1(n13102), .C2(n10661), .ZN(P3_U3291) );
  INV_X1 U13372 ( .A(SI_7_), .ZN(n10665) );
  INV_X1 U13373 ( .A(n10663), .ZN(n10664) );
  OAI222_X1 U13374 ( .A1(P3_U3151), .A2(n7718), .B1(n13962), .B2(n10665), .C1(
        n13102), .C2(n10664), .ZN(P3_U3288) );
  INV_X1 U13375 ( .A(SI_2_), .ZN(n10668) );
  INV_X1 U13376 ( .A(n10666), .ZN(n10667) );
  OAI222_X1 U13377 ( .A1(P3_U3151), .A2(n11312), .B1(n13962), .B2(n10668), 
        .C1(n13102), .C2(n10667), .ZN(P3_U3293) );
  OAI222_X1 U13378 ( .A1(P3_U3151), .A2(n10671), .B1(n13962), .B2(n10670), 
        .C1(n13102), .C2(n10669), .ZN(P3_U3285) );
  INV_X1 U13379 ( .A(n10672), .ZN(n10701) );
  INV_X1 U13380 ( .A(n15163), .ZN(n10673) );
  OAI222_X1 U13381 ( .A1(n15700), .A2(n10674), .B1(n15703), .B2(n10701), .C1(
        n10673), .C2(P1_U3086), .ZN(P1_U3348) );
  NAND2_X1 U13382 ( .A1(n10676), .A2(n10675), .ZN(n10677) );
  NAND2_X1 U13383 ( .A1(n10677), .A2(P3_ADDR_REG_5__SCAN_IN), .ZN(n11049) );
  INV_X1 U13384 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n10678) );
  NAND2_X1 U13385 ( .A1(n10679), .A2(P2_ADDR_REG_4__SCAN_IN), .ZN(n10680) );
  NAND2_X1 U13386 ( .A1(n10681), .A2(n10680), .ZN(n11044) );
  INV_X1 U13387 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n11042) );
  XNOR2_X1 U13388 ( .A(n11043), .B(n11042), .ZN(SUB_1596_U58) );
  OAI222_X1 U13389 ( .A1(P3_U3151), .A2(n12601), .B1(n13962), .B2(n10683), 
        .C1(n13102), .C2(n10682), .ZN(P3_U3284) );
  AOI22_X1 U13390 ( .A1(n15821), .A2(n10686), .B1(n10685), .B2(n10687), .ZN(
        P1_U3446) );
  INV_X1 U13391 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n10689) );
  AOI22_X1 U13392 ( .A1(n15821), .A2(n10689), .B1(n10688), .B2(n10687), .ZN(
        P1_U3445) );
  CLKBUF_X1 U13393 ( .A(n15700), .Z(n13134) );
  INV_X1 U13394 ( .A(n10690), .ZN(n10698) );
  INV_X1 U13395 ( .A(n11097), .ZN(n10691) );
  OAI222_X1 U13396 ( .A1(n13134), .A2(n10692), .B1(n15703), .B2(n10698), .C1(
        n10691), .C2(P1_U3086), .ZN(P1_U3350) );
  INV_X1 U13397 ( .A(n10693), .ZN(n10706) );
  INV_X1 U13398 ( .A(n11201), .ZN(n10694) );
  OAI222_X1 U13399 ( .A1(n13134), .A2(n10779), .B1(n15703), .B2(n10706), .C1(
        n10694), .C2(P1_U3086), .ZN(P1_U3349) );
  OAI222_X1 U13400 ( .A1(n13134), .A2(n10820), .B1(n15703), .B2(n10702), .C1(
        n9518), .C2(P1_U3086), .ZN(P1_U3353) );
  AND2_X1 U13401 ( .A1(n7218), .A2(P2_U3088), .ZN(n14897) );
  INV_X2 U13402 ( .A(n14897), .ZN(n14914) );
  NAND2_X1 U13403 ( .A1(n10696), .A2(P2_U3088), .ZN(n14917) );
  INV_X1 U13404 ( .A(n14451), .ZN(n10697) );
  OAI222_X1 U13405 ( .A1(n14914), .A2(n10699), .B1(n14917), .B2(n10698), .C1(
        P2_U3088), .C2(n10697), .ZN(P2_U3322) );
  INV_X1 U13406 ( .A(n14470), .ZN(n10700) );
  OAI222_X1 U13407 ( .A1(n14914), .A2(n10964), .B1(n14917), .B2(n10701), .C1(
        P2_U3088), .C2(n10700), .ZN(P2_U3320) );
  OAI222_X1 U13408 ( .A1(n14914), .A2(n10703), .B1(n14917), .B2(n10702), .C1(
        P2_U3088), .C2(n8053), .ZN(P2_U3325) );
  INV_X1 U13409 ( .A(n14428), .ZN(n10704) );
  OAI222_X1 U13410 ( .A1(n14914), .A2(n10705), .B1(n14917), .B2(n7802), .C1(
        P2_U3088), .C2(n10704), .ZN(P2_U3324) );
  INV_X1 U13411 ( .A(n11168), .ZN(n15918) );
  OAI222_X1 U13412 ( .A1(n14914), .A2(n10707), .B1(n14917), .B2(n10706), .C1(
        P2_U3088), .C2(n15918), .ZN(P2_U3321) );
  INV_X1 U13413 ( .A(n14440), .ZN(n10708) );
  OAI222_X1 U13414 ( .A1(n14914), .A2(n10710), .B1(n14917), .B2(n10709), .C1(
        P2_U3088), .C2(n10708), .ZN(P2_U3323) );
  INV_X1 U13415 ( .A(n10711), .ZN(n10715) );
  INV_X1 U13416 ( .A(n14484), .ZN(n10712) );
  OAI222_X1 U13417 ( .A1(n14914), .A2(n10713), .B1(n14917), .B2(n10715), .C1(
        P2_U3088), .C2(n10712), .ZN(P2_U3319) );
  INV_X1 U13418 ( .A(n11116), .ZN(n10714) );
  OAI222_X1 U13419 ( .A1(n15700), .A2(n10716), .B1(n15703), .B2(n10715), .C1(
        n10714), .C2(P1_U3086), .ZN(P1_U3347) );
  INV_X1 U13420 ( .A(n12318), .ZN(n10717) );
  NAND2_X1 U13421 ( .A1(n11830), .A2(n10717), .ZN(n10723) );
  NAND2_X1 U13422 ( .A1(n10719), .A2(n10718), .ZN(n10720) );
  INV_X1 U13423 ( .A(n10722), .ZN(n10721) );
  NAND2_X1 U13424 ( .A1(n10723), .A2(n10721), .ZN(n15252) );
  AND2_X1 U13425 ( .A1(n10723), .A2(n10722), .ZN(n11082) );
  INV_X1 U13426 ( .A(n15699), .ZN(n15113) );
  NAND2_X1 U13427 ( .A1(n15113), .A2(n9492), .ZN(n10724) );
  NAND2_X1 U13428 ( .A1(n11071), .A2(n10724), .ZN(n15116) );
  AOI21_X1 U13429 ( .B1(n15699), .B2(n10725), .A(n15116), .ZN(n10726) );
  XNOR2_X1 U13430 ( .A(n10726), .B(n7444), .ZN(n10727) );
  AOI22_X1 U13431 ( .A1(n11082), .A2(n10727), .B1(P1_REG3_REG_0__SCAN_IN), 
        .B2(P1_U3086), .ZN(n10728) );
  OAI21_X1 U13432 ( .B1(n10729), .B2(n15252), .A(n10728), .ZN(P1_U3243) );
  OAI222_X1 U13433 ( .A1(P3_U3151), .A2(n8836), .B1(n13962), .B2(n10731), .C1(
        n13102), .C2(n10730), .ZN(P3_U3294) );
  INV_X1 U13434 ( .A(SI_3_), .ZN(n10734) );
  INV_X1 U13435 ( .A(n10732), .ZN(n10733) );
  OAI222_X1 U13436 ( .A1(P3_U3151), .A2(n7696), .B1(n13962), .B2(n10734), .C1(
        n13102), .C2(n10733), .ZN(P3_U3292) );
  OAI222_X1 U13437 ( .A1(n10739), .A2(P3_U3151), .B1(n13102), .B2(n10738), 
        .C1(n10737), .C2(n13962), .ZN(P3_U3289) );
  OAI222_X1 U13438 ( .A1(n12061), .A2(P3_U3151), .B1(n13102), .B2(n10741), 
        .C1(n10740), .C2(n13962), .ZN(P3_U3286) );
  INV_X1 U13439 ( .A(n10742), .ZN(n10743) );
  OAI222_X1 U13440 ( .A1(P3_U3151), .A2(n13515), .B1(n13962), .B2(n10744), 
        .C1(n13102), .C2(n10743), .ZN(P3_U3283) );
  INV_X1 U13441 ( .A(n10745), .ZN(n10748) );
  INV_X1 U13442 ( .A(n11370), .ZN(n10746) );
  OAI222_X1 U13443 ( .A1(n13134), .A2(n10747), .B1(n15703), .B2(n10748), .C1(
        n10746), .C2(P1_U3086), .ZN(P1_U3346) );
  INV_X1 U13444 ( .A(n11221), .ZN(n11183) );
  OAI222_X1 U13445 ( .A1(n14914), .A2(n10749), .B1(n14917), .B2(n10748), .C1(
        P2_U3088), .C2(n11183), .ZN(P2_U3318) );
  INV_X1 U13446 ( .A(n14917), .ZN(n14906) );
  INV_X1 U13447 ( .A(n14906), .ZN(n14903) );
  OAI222_X1 U13448 ( .A1(n8035), .A2(P2_U3088), .B1(n14903), .B2(n10751), .C1(
        n10750), .C2(n14914), .ZN(P2_U3326) );
  INV_X1 U13449 ( .A(n9383), .ZN(n10752) );
  NOR2_X1 U13450 ( .A1(n13959), .A2(n10752), .ZN(n10755) );
  CLKBUF_X1 U13451 ( .A(n10755), .Z(n10775) );
  INV_X1 U13452 ( .A(P3_D_REG_2__SCAN_IN), .ZN(n10753) );
  NOR2_X1 U13453 ( .A1(n10775), .A2(n10753), .ZN(P3_U3263) );
  INV_X1 U13454 ( .A(P3_D_REG_16__SCAN_IN), .ZN(n10754) );
  NOR2_X1 U13455 ( .A1(n10775), .A2(n10754), .ZN(P3_U3249) );
  INV_X1 U13456 ( .A(P3_D_REG_23__SCAN_IN), .ZN(n10756) );
  NOR2_X1 U13457 ( .A1(n10775), .A2(n10756), .ZN(P3_U3242) );
  INV_X1 U13458 ( .A(P3_D_REG_28__SCAN_IN), .ZN(n10757) );
  NOR2_X1 U13459 ( .A1(n10755), .A2(n10757), .ZN(P3_U3237) );
  INV_X1 U13460 ( .A(P3_D_REG_24__SCAN_IN), .ZN(n10758) );
  NOR2_X1 U13461 ( .A1(n10755), .A2(n10758), .ZN(P3_U3241) );
  INV_X1 U13462 ( .A(P3_D_REG_3__SCAN_IN), .ZN(n10923) );
  NOR2_X1 U13463 ( .A1(n10755), .A2(n10923), .ZN(P3_U3262) );
  INV_X1 U13464 ( .A(P3_D_REG_26__SCAN_IN), .ZN(n10759) );
  NOR2_X1 U13465 ( .A1(n10755), .A2(n10759), .ZN(P3_U3239) );
  INV_X1 U13466 ( .A(P3_D_REG_4__SCAN_IN), .ZN(n10760) );
  NOR2_X1 U13467 ( .A1(n10775), .A2(n10760), .ZN(P3_U3261) );
  INV_X1 U13468 ( .A(P3_D_REG_21__SCAN_IN), .ZN(n10761) );
  NOR2_X1 U13469 ( .A1(n10755), .A2(n10761), .ZN(P3_U3244) );
  INV_X1 U13470 ( .A(P3_D_REG_8__SCAN_IN), .ZN(n10892) );
  NOR2_X1 U13471 ( .A1(n10775), .A2(n10892), .ZN(P3_U3257) );
  INV_X1 U13472 ( .A(P3_D_REG_9__SCAN_IN), .ZN(n10857) );
  NOR2_X1 U13473 ( .A1(n10775), .A2(n10857), .ZN(P3_U3256) );
  INV_X1 U13474 ( .A(P3_D_REG_10__SCAN_IN), .ZN(n10921) );
  NOR2_X1 U13475 ( .A1(n10775), .A2(n10921), .ZN(P3_U3255) );
  INV_X1 U13476 ( .A(P3_D_REG_7__SCAN_IN), .ZN(n10916) );
  NOR2_X1 U13477 ( .A1(n10755), .A2(n10916), .ZN(P3_U3258) );
  INV_X1 U13478 ( .A(P3_D_REG_6__SCAN_IN), .ZN(n10762) );
  NOR2_X1 U13479 ( .A1(n10775), .A2(n10762), .ZN(P3_U3259) );
  INV_X1 U13480 ( .A(P3_D_REG_5__SCAN_IN), .ZN(n10763) );
  NOR2_X1 U13481 ( .A1(n10755), .A2(n10763), .ZN(P3_U3260) );
  INV_X1 U13482 ( .A(P3_D_REG_12__SCAN_IN), .ZN(n10764) );
  NOR2_X1 U13483 ( .A1(n10775), .A2(n10764), .ZN(P3_U3253) );
  INV_X1 U13484 ( .A(P3_D_REG_13__SCAN_IN), .ZN(n10837) );
  NOR2_X1 U13485 ( .A1(n10775), .A2(n10837), .ZN(P3_U3252) );
  INV_X1 U13486 ( .A(P3_D_REG_14__SCAN_IN), .ZN(n10867) );
  NOR2_X1 U13487 ( .A1(n10775), .A2(n10867), .ZN(P3_U3251) );
  INV_X1 U13488 ( .A(P3_D_REG_15__SCAN_IN), .ZN(n10765) );
  NOR2_X1 U13489 ( .A1(n10775), .A2(n10765), .ZN(P3_U3250) );
  INV_X1 U13490 ( .A(P3_D_REG_31__SCAN_IN), .ZN(n10766) );
  NOR2_X1 U13491 ( .A1(n10755), .A2(n10766), .ZN(P3_U3234) );
  INV_X1 U13492 ( .A(P3_D_REG_17__SCAN_IN), .ZN(n10767) );
  NOR2_X1 U13493 ( .A1(n10775), .A2(n10767), .ZN(P3_U3248) );
  INV_X1 U13494 ( .A(P3_D_REG_18__SCAN_IN), .ZN(n10768) );
  NOR2_X1 U13495 ( .A1(n10775), .A2(n10768), .ZN(P3_U3247) );
  INV_X1 U13496 ( .A(P3_D_REG_19__SCAN_IN), .ZN(n10769) );
  NOR2_X1 U13497 ( .A1(n10775), .A2(n10769), .ZN(P3_U3246) );
  INV_X1 U13498 ( .A(P3_D_REG_20__SCAN_IN), .ZN(n10770) );
  NOR2_X1 U13499 ( .A1(n10755), .A2(n10770), .ZN(P3_U3245) );
  INV_X1 U13500 ( .A(P3_D_REG_25__SCAN_IN), .ZN(n10771) );
  NOR2_X1 U13501 ( .A1(n10755), .A2(n10771), .ZN(P3_U3240) );
  INV_X1 U13502 ( .A(P3_D_REG_22__SCAN_IN), .ZN(n10772) );
  NOR2_X1 U13503 ( .A1(n10755), .A2(n10772), .ZN(P3_U3243) );
  INV_X1 U13504 ( .A(P3_D_REG_27__SCAN_IN), .ZN(n10883) );
  NOR2_X1 U13505 ( .A1(n10775), .A2(n10883), .ZN(P3_U3238) );
  INV_X1 U13506 ( .A(P3_D_REG_29__SCAN_IN), .ZN(n10773) );
  NOR2_X1 U13507 ( .A1(n10775), .A2(n10773), .ZN(P3_U3236) );
  INV_X1 U13508 ( .A(P3_D_REG_11__SCAN_IN), .ZN(n10774) );
  NOR2_X1 U13509 ( .A1(n10775), .A2(n10774), .ZN(P3_U3254) );
  INV_X1 U13510 ( .A(P3_D_REG_30__SCAN_IN), .ZN(n10776) );
  NOR2_X1 U13511 ( .A1(n10775), .A2(n10776), .ZN(P3_U3235) );
  MUX2_X1 U13512 ( .A(n7149), .B(P3_DATAO_REG_1__SCAN_IN), .S(n13510), .Z(
        n11035) );
  INV_X1 U13513 ( .A(P3_ADDR_REG_13__SCAN_IN), .ZN(n12850) );
  INV_X1 U13514 ( .A(P3_REG3_REG_16__SCAN_IN), .ZN(n10945) );
  NAND4_X1 U13515 ( .A1(P2_DATAO_REG_9__SCAN_IN), .A2(P3_REG1_REG_24__SCAN_IN), 
        .A3(n12925), .A4(n10945), .ZN(n10778) );
  NAND4_X1 U13516 ( .A1(P1_DATAO_REG_28__SCAN_IN), .A2(P3_REG3_REG_23__SCAN_IN), .A3(P3_REG2_REG_10__SCAN_IN), .A4(n14890), .ZN(n10777) );
  OR4_X1 U13517 ( .A1(n12850), .A2(n10934), .A3(n10778), .A4(n10777), .ZN(
        n10781) );
  NAND4_X1 U13518 ( .A1(n10779), .A2(n10965), .A3(P2_IR_REG_2__SCAN_IN), .A4(
        SI_27_), .ZN(n10780) );
  NOR4_X1 U13519 ( .A1(n10781), .A2(n10780), .A3(n14884), .A4(n10935), .ZN(
        n10834) );
  INV_X1 U13520 ( .A(P3_DATAO_REG_23__SCAN_IN), .ZN(n12095) );
  INV_X1 U13521 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n12846) );
  INV_X1 U13522 ( .A(P3_ADDR_REG_12__SCAN_IN), .ZN(n13517) );
  NAND4_X1 U13523 ( .A1(P1_REG0_REG_23__SCAN_IN), .A2(P2_DATAO_REG_18__SCAN_IN), .A3(n12846), .A4(n13517), .ZN(n10784) );
  NAND4_X1 U13524 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P3_REG2_REG_26__SCAN_IN), 
        .A3(P2_REG2_REG_31__SCAN_IN), .A4(n11556), .ZN(n10783) );
  NAND4_X1 U13525 ( .A1(P3_IR_REG_8__SCAN_IN), .A2(P1_REG1_REG_25__SCAN_IN), 
        .A3(P1_REG0_REG_22__SCAN_IN), .A4(n12507), .ZN(n10782) );
  NOR4_X1 U13526 ( .A1(P1_REG2_REG_23__SCAN_IN), .A2(n10784), .A3(n10783), 
        .A4(n10782), .ZN(n10786) );
  AND4_X1 U13527 ( .A1(n12095), .A2(P3_REG0_REG_6__SCAN_IN), .A3(n10786), .A4(
        n10785), .ZN(n10833) );
  NOR4_X1 U13528 ( .A1(P2_REG1_REG_16__SCAN_IN), .A2(P3_D_REG_14__SCAN_IN), 
        .A3(P1_D_REG_10__SCAN_IN), .A4(n13080), .ZN(n10787) );
  NAND3_X1 U13529 ( .A1(P3_REG3_REG_21__SCAN_IN), .A2(P1_REG2_REG_7__SCAN_IN), 
        .A3(n10787), .ZN(n10799) );
  NAND4_X1 U13530 ( .A1(n11041), .A2(P2_REG1_REG_21__SCAN_IN), .A3(
        P3_IR_REG_12__SCAN_IN), .A4(P3_REG2_REG_16__SCAN_IN), .ZN(n10789) );
  INV_X1 U13531 ( .A(P3_DATAO_REG_3__SCAN_IN), .ZN(n10788) );
  NOR3_X1 U13532 ( .A1(n10789), .A2(n10788), .A3(P3_D_REG_27__SCAN_IN), .ZN(
        n10797) );
  INV_X1 U13533 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n10922) );
  NAND4_X1 U13534 ( .A1(P3_D_REG_10__SCAN_IN), .A2(P1_D_REG_2__SCAN_IN), .A3(
        n10922), .A4(n9747), .ZN(n10795) );
  NAND4_X1 U13535 ( .A1(P3_D_REG_8__SCAN_IN), .A2(P3_IR_REG_4__SCAN_IN), .A3(
        n13699), .A4(n8917), .ZN(n10794) );
  INV_X1 U13536 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n11141) );
  INV_X1 U13537 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n11911) );
  NAND4_X1 U13538 ( .A1(P1_IR_REG_6__SCAN_IN), .A2(n14913), .A3(n11141), .A4(
        n11911), .ZN(n10790) );
  NOR2_X1 U13539 ( .A1(P3_REG1_REG_26__SCAN_IN), .A2(n10790), .ZN(n10792) );
  NAND4_X1 U13540 ( .A1(n10792), .A2(P2_REG2_REG_20__SCAN_IN), .A3(n10791), 
        .A4(P3_REG0_REG_29__SCAN_IN), .ZN(n10793) );
  NOR3_X1 U13541 ( .A1(n10795), .A2(n10794), .A3(n10793), .ZN(n10796) );
  NAND4_X1 U13542 ( .A1(P1_REG1_REG_31__SCAN_IN), .A2(n10797), .A3(n10796), 
        .A4(n11669), .ZN(n10798) );
  NOR4_X1 U13543 ( .A1(P1_DATAO_REG_19__SCAN_IN), .A2(n14378), .A3(n10799), 
        .A4(n10798), .ZN(n10832) );
  NAND4_X1 U13544 ( .A1(n10801), .A2(n10800), .A3(P1_ADDR_REG_3__SCAN_IN), 
        .A4(P2_ADDR_REG_2__SCAN_IN), .ZN(n10808) );
  NOR4_X1 U13545 ( .A1(P2_REG1_REG_26__SCAN_IN), .A2(P2_REG2_REG_10__SCAN_IN), 
        .A3(P1_REG3_REG_1__SCAN_IN), .A4(n10993), .ZN(n10806) );
  INV_X1 U13546 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n15161) );
  INV_X1 U13547 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n14464) );
  NOR4_X1 U13548 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(n10802), .A3(n15161), .A4(
        n14464), .ZN(n10805) );
  NOR4_X1 U13549 ( .A1(P2_DATAO_REG_24__SCAN_IN), .A2(P3_REG0_REG_15__SCAN_IN), 
        .A3(P1_REG3_REG_22__SCAN_IN), .A4(P1_REG1_REG_8__SCAN_IN), .ZN(n10804)
         );
  NOR4_X1 U13550 ( .A1(P1_REG1_REG_27__SCAN_IN), .A2(P3_REG1_REG_7__SCAN_IN), 
        .A3(P1_REG0_REG_8__SCAN_IN), .A4(n12144), .ZN(n10803) );
  NAND4_X1 U13551 ( .A1(n10806), .A2(n10805), .A3(n10804), .A4(n10803), .ZN(
        n10807) );
  OR4_X1 U13552 ( .A1(P1_ADDR_REG_2__SCAN_IN), .A2(P3_ADDR_REG_2__SCAN_IN), 
        .A3(n10808), .A4(n10807), .ZN(n10830) );
  NAND4_X1 U13553 ( .A1(P3_D_REG_9__SCAN_IN), .A2(P2_D_REG_26__SCAN_IN), .A3(
        P1_REG1_REG_3__SCAN_IN), .A4(n10848), .ZN(n10809) );
  NOR3_X1 U13554 ( .A1(P3_DATAO_REG_17__SCAN_IN), .A2(n11128), .A3(n10809), 
        .ZN(n10827) );
  NAND4_X1 U13555 ( .A1(n8006), .A2(n10811), .A3(n10810), .A4(
        P2_IR_REG_24__SCAN_IN), .ZN(n10814) );
  INV_X1 U13556 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n15943) );
  NAND4_X1 U13557 ( .A1(n10812), .A2(n15943), .A3(P3_D_REG_13__SCAN_IN), .A4(
        P1_D_REG_30__SCAN_IN), .ZN(n10813) );
  NOR2_X1 U13558 ( .A1(n10814), .A2(n10813), .ZN(n10826) );
  NAND4_X1 U13559 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P1_DATAO_REG_7__SCAN_IN), 
        .A3(P1_DATAO_REG_26__SCAN_IN), .A4(P1_D_REG_16__SCAN_IN), .ZN(n10824)
         );
  INV_X1 U13560 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n10956) );
  AND4_X1 U13561 ( .A1(P1_REG3_REG_25__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .A3(n10956), .A4(n13851), .ZN(n10815) );
  INV_X1 U13562 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n10846) );
  NAND4_X1 U13563 ( .A1(n10815), .A2(n11157), .A3(n10846), .A4(n9485), .ZN(
        n10818) );
  NAND2_X1 U13564 ( .A1(n10816), .A2(n15395), .ZN(n10817) );
  NOR2_X1 U13565 ( .A1(n10818), .A2(n10817), .ZN(n10819) );
  NAND4_X1 U13566 ( .A1(n11259), .A2(n10820), .A3(n13906), .A4(n10819), .ZN(
        n10823) );
  NAND4_X1 U13567 ( .A1(n10821), .A2(P2_IR_REG_18__SCAN_IN), .A3(
        P3_REG1_REG_10__SCAN_IN), .A4(P3_REG3_REG_0__SCAN_IN), .ZN(n10822) );
  NOR3_X1 U13568 ( .A1(n10824), .A2(n10823), .A3(n10822), .ZN(n10825) );
  NAND4_X1 U13569 ( .A1(n10828), .A2(n10827), .A3(n10826), .A4(n10825), .ZN(
        n10829) );
  NOR2_X1 U13570 ( .A1(n10830), .A2(n10829), .ZN(n10831) );
  NAND4_X1 U13571 ( .A1(n10834), .A2(n10833), .A3(n10832), .A4(n10831), .ZN(
        n11033) );
  AOI22_X1 U13572 ( .A1(n15395), .A2(keyinput21), .B1(n11157), .B2(keyinput115), .ZN(n10835) );
  OAI221_X1 U13573 ( .B1(n15395), .B2(keyinput21), .C1(n11157), .C2(
        keyinput115), .A(n10835), .ZN(n10844) );
  INV_X1 U13574 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n15732) );
  AOI22_X1 U13575 ( .A1(n15732), .A2(keyinput24), .B1(n10837), .B2(keyinput82), 
        .ZN(n10836) );
  OAI221_X1 U13576 ( .B1(n15732), .B2(keyinput24), .C1(n10837), .C2(keyinput82), .A(n10836), .ZN(n10843) );
  XNOR2_X1 U13577 ( .A(P1_REG3_REG_12__SCAN_IN), .B(keyinput121), .ZN(n10841)
         );
  XNOR2_X1 U13578 ( .A(P2_IR_REG_31__SCAN_IN), .B(keyinput45), .ZN(n10840) );
  XNOR2_X1 U13579 ( .A(P2_REG1_REG_20__SCAN_IN), .B(keyinput92), .ZN(n10839)
         );
  XNOR2_X1 U13580 ( .A(P1_IR_REG_3__SCAN_IN), .B(keyinput71), .ZN(n10838) );
  NAND4_X1 U13581 ( .A1(n10841), .A2(n10840), .A3(n10839), .A4(n10838), .ZN(
        n10842) );
  NOR3_X1 U13582 ( .A1(n10844), .A2(n10843), .A3(n10842), .ZN(n10880) );
  INV_X1 U13583 ( .A(P1_D_REG_30__SCAN_IN), .ZN(n15816) );
  AOI22_X1 U13584 ( .A1(n15816), .A2(keyinput107), .B1(n10846), .B2(keyinput58), .ZN(n10845) );
  OAI221_X1 U13585 ( .B1(n15816), .B2(keyinput107), .C1(n10846), .C2(
        keyinput58), .A(n10845), .ZN(n10855) );
  AOI22_X1 U13586 ( .A1(n9485), .A2(keyinput83), .B1(n10848), .B2(keyinput79), 
        .ZN(n10847) );
  OAI221_X1 U13587 ( .B1(n9485), .B2(keyinput83), .C1(n10848), .C2(keyinput79), 
        .A(n10847), .ZN(n10854) );
  AOI22_X1 U13588 ( .A1(n15943), .A2(keyinput81), .B1(n12733), .B2(keyinput51), 
        .ZN(n10849) );
  OAI221_X1 U13589 ( .B1(n15943), .B2(keyinput81), .C1(n12733), .C2(keyinput51), .A(n10849), .ZN(n10853) );
  XNOR2_X1 U13590 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(keyinput102), .ZN(n10851)
         );
  XNOR2_X1 U13591 ( .A(P2_IR_REG_18__SCAN_IN), .B(keyinput29), .ZN(n10850) );
  NAND2_X1 U13592 ( .A1(n10851), .A2(n10850), .ZN(n10852) );
  NOR4_X1 U13593 ( .A1(n10855), .A2(n10854), .A3(n10853), .A4(n10852), .ZN(
        n10879) );
  INV_X1 U13594 ( .A(P2_D_REG_11__SCAN_IN), .ZN(n15967) );
  AOI22_X1 U13595 ( .A1(n15967), .A2(keyinput16), .B1(keyinput86), .B2(n10857), 
        .ZN(n10856) );
  OAI221_X1 U13596 ( .B1(n15967), .B2(keyinput16), .C1(n10857), .C2(keyinput86), .A(n10856), .ZN(n10865) );
  INV_X1 U13597 ( .A(P3_DATAO_REG_17__SCAN_IN), .ZN(n11314) );
  AOI22_X1 U13598 ( .A1(n11314), .A2(keyinput68), .B1(n11128), .B2(keyinput39), 
        .ZN(n10858) );
  OAI221_X1 U13599 ( .B1(n11314), .B2(keyinput68), .C1(n11128), .C2(keyinput39), .A(n10858), .ZN(n10864) );
  AOI22_X1 U13600 ( .A1(n11064), .A2(keyinput7), .B1(keyinput47), .B2(n15161), 
        .ZN(n10859) );
  OAI221_X1 U13601 ( .B1(n11064), .B2(keyinput7), .C1(n15161), .C2(keyinput47), 
        .A(n10859), .ZN(n10863) );
  INV_X1 U13602 ( .A(P2_D_REG_26__SCAN_IN), .ZN(n15951) );
  AOI22_X1 U13603 ( .A1(n15951), .A2(keyinput41), .B1(keyinput54), .B2(n10861), 
        .ZN(n10860) );
  OAI221_X1 U13604 ( .B1(n15951), .B2(keyinput41), .C1(n10861), .C2(keyinput54), .A(n10860), .ZN(n10862) );
  NOR4_X1 U13605 ( .A1(n10865), .A2(n10864), .A3(n10863), .A4(n10862), .ZN(
        n10878) );
  AOI22_X1 U13606 ( .A1(n9590), .A2(keyinput55), .B1(n10867), .B2(keyinput57), 
        .ZN(n10866) );
  OAI221_X1 U13607 ( .B1(n9590), .B2(keyinput55), .C1(n10867), .C2(keyinput57), 
        .A(n10866), .ZN(n10872) );
  INV_X1 U13608 ( .A(P2_D_REG_4__SCAN_IN), .ZN(n15974) );
  XNOR2_X1 U13609 ( .A(n15974), .B(keyinput22), .ZN(n10871) );
  XOR2_X1 U13610 ( .A(P1_IR_REG_8__SCAN_IN), .B(keyinput93), .Z(n10870) );
  XNOR2_X1 U13611 ( .A(n10868), .B(keyinput32), .ZN(n10869) );
  OR4_X1 U13612 ( .A1(n10872), .A2(n10871), .A3(n10870), .A4(n10869), .ZN(
        n10876) );
  INV_X1 U13613 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n14815) );
  INV_X1 U13614 ( .A(P1_D_REG_10__SCAN_IN), .ZN(n15820) );
  AOI22_X1 U13615 ( .A1(n14815), .A2(keyinput35), .B1(keyinput89), .B2(n15820), 
        .ZN(n10873) );
  OAI221_X1 U13616 ( .B1(n14815), .B2(keyinput35), .C1(n15820), .C2(keyinput89), .A(n10873), .ZN(n10875) );
  INV_X1 U13617 ( .A(P1_D_REG_21__SCAN_IN), .ZN(n15818) );
  XNOR2_X1 U13618 ( .A(n15818), .B(keyinput49), .ZN(n10874) );
  NOR3_X1 U13619 ( .A1(n10876), .A2(n10875), .A3(n10874), .ZN(n10877) );
  NAND4_X1 U13620 ( .A1(n10880), .A2(n10879), .A3(n10878), .A4(n10877), .ZN(
        n11031) );
  AOI22_X1 U13621 ( .A1(n13080), .A2(keyinput53), .B1(keyinput36), .B2(n10629), 
        .ZN(n10881) );
  OAI221_X1 U13622 ( .B1(n13080), .B2(keyinput53), .C1(n10629), .C2(keyinput36), .A(n10881), .ZN(n10890) );
  AOI22_X1 U13623 ( .A1(n10883), .A2(keyinput43), .B1(n14787), .B2(keyinput127), .ZN(n10882) );
  OAI221_X1 U13624 ( .B1(n10883), .B2(keyinput43), .C1(n14787), .C2(
        keyinput127), .A(n10882), .ZN(n10889) );
  INV_X1 U13625 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n13105) );
  AOI22_X1 U13626 ( .A1(n14378), .A2(keyinput100), .B1(keyinput14), .B2(n13105), .ZN(n10884) );
  OAI221_X1 U13627 ( .B1(n14378), .B2(keyinput100), .C1(n13105), .C2(
        keyinput14), .A(n10884), .ZN(n10888) );
  XOR2_X1 U13628 ( .A(n10788), .B(keyinput8), .Z(n10886) );
  XNOR2_X1 U13629 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(keyinput66), .ZN(n10885)
         );
  NAND2_X1 U13630 ( .A1(n10886), .A2(n10885), .ZN(n10887) );
  NOR4_X1 U13631 ( .A1(n10890), .A2(n10889), .A3(n10888), .A4(n10887), .ZN(
        n10930) );
  AOI22_X1 U13632 ( .A1(n10892), .A2(keyinput46), .B1(keyinput117), .B2(n8917), 
        .ZN(n10891) );
  OAI221_X1 U13633 ( .B1(n10892), .B2(keyinput46), .C1(n8917), .C2(keyinput117), .A(n10891), .ZN(n10901) );
  INV_X1 U13634 ( .A(P2_D_REG_29__SCAN_IN), .ZN(n15948) );
  AOI22_X1 U13635 ( .A1(n10894), .A2(keyinput80), .B1(n15948), .B2(keyinput99), 
        .ZN(n10893) );
  OAI221_X1 U13636 ( .B1(n10894), .B2(keyinput80), .C1(n15948), .C2(keyinput99), .A(n10893), .ZN(n10900) );
  AOI22_X1 U13637 ( .A1(n11669), .A2(keyinput125), .B1(keyinput73), .B2(n13808), .ZN(n10895) );
  OAI221_X1 U13638 ( .B1(n11669), .B2(keyinput125), .C1(n13808), .C2(
        keyinput73), .A(n10895), .ZN(n10899) );
  XNOR2_X1 U13639 ( .A(P3_IR_REG_12__SCAN_IN), .B(keyinput63), .ZN(n10897) );
  XNOR2_X1 U13640 ( .A(P3_IR_REG_4__SCAN_IN), .B(keyinput70), .ZN(n10896) );
  NAND2_X1 U13641 ( .A1(n10897), .A2(n10896), .ZN(n10898) );
  NOR4_X1 U13642 ( .A1(n10901), .A2(n10900), .A3(n10899), .A4(n10898), .ZN(
        n10929) );
  AOI22_X1 U13643 ( .A1(n11141), .A2(keyinput19), .B1(keyinput10), .B2(n11911), 
        .ZN(n10902) );
  OAI221_X1 U13644 ( .B1(n11141), .B2(keyinput19), .C1(n11911), .C2(keyinput10), .A(n10902), .ZN(n10912) );
  INV_X1 U13645 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n10904) );
  AOI22_X1 U13646 ( .A1(n10905), .A2(keyinput95), .B1(n10904), .B2(keyinput120), .ZN(n10903) );
  OAI221_X1 U13647 ( .B1(n10905), .B2(keyinput95), .C1(n10904), .C2(
        keyinput120), .A(n10903), .ZN(n10911) );
  XNOR2_X1 U13648 ( .A(P1_IR_REG_6__SCAN_IN), .B(keyinput123), .ZN(n10909) );
  XNOR2_X1 U13649 ( .A(P3_REG2_REG_24__SCAN_IN), .B(keyinput113), .ZN(n10908)
         );
  XNOR2_X1 U13650 ( .A(P2_REG3_REG_6__SCAN_IN), .B(keyinput72), .ZN(n10907) );
  XNOR2_X1 U13651 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(keyinput103), .ZN(n10906)
         );
  NAND4_X1 U13652 ( .A1(n10909), .A2(n10908), .A3(n10907), .A4(n10906), .ZN(
        n10910) );
  NOR3_X1 U13653 ( .A1(n10912), .A2(n10911), .A3(n10910), .ZN(n10928) );
  AOI22_X1 U13654 ( .A1(n10914), .A2(keyinput84), .B1(keyinput27), .B2(n9747), 
        .ZN(n10913) );
  OAI221_X1 U13655 ( .B1(n10914), .B2(keyinput84), .C1(n9747), .C2(keyinput27), 
        .A(n10913), .ZN(n10919) );
  INV_X1 U13656 ( .A(P1_D_REG_2__SCAN_IN), .ZN(n15822) );
  AOI22_X1 U13657 ( .A1(n10916), .A2(keyinput37), .B1(keyinput116), .B2(n15822), .ZN(n10915) );
  OAI221_X1 U13658 ( .B1(n10916), .B2(keyinput37), .C1(n15822), .C2(
        keyinput116), .A(n10915), .ZN(n10918) );
  XNOR2_X1 U13659 ( .A(n11259), .B(keyinput109), .ZN(n10917) );
  OR3_X1 U13660 ( .A1(n10919), .A2(n10918), .A3(n10917), .ZN(n10926) );
  AOI22_X1 U13661 ( .A1(n10922), .A2(keyinput6), .B1(keyinput5), .B2(n10921), 
        .ZN(n10920) );
  OAI221_X1 U13662 ( .B1(n10922), .B2(keyinput6), .C1(n10921), .C2(keyinput5), 
        .A(n10920), .ZN(n10925) );
  XNOR2_X1 U13663 ( .A(n10923), .B(keyinput67), .ZN(n10924) );
  NOR3_X1 U13664 ( .A1(n10926), .A2(n10925), .A3(n10924), .ZN(n10927) );
  NAND4_X1 U13665 ( .A1(n10930), .A2(n10929), .A3(n10928), .A4(n10927), .ZN(
        n11030) );
  AOI22_X1 U13666 ( .A1(n14884), .A2(keyinput18), .B1(n13109), .B2(keyinput96), 
        .ZN(n10931) );
  OAI221_X1 U13667 ( .B1(n14884), .B2(keyinput18), .C1(n13109), .C2(keyinput96), .A(n10931), .ZN(n10941) );
  AOI22_X1 U13668 ( .A1(n14910), .A2(keyinput105), .B1(keyinput94), .B2(n12624), .ZN(n10932) );
  OAI221_X1 U13669 ( .B1(n14910), .B2(keyinput105), .C1(n12624), .C2(
        keyinput94), .A(n10932), .ZN(n10940) );
  AOI22_X1 U13670 ( .A1(n10935), .A2(keyinput91), .B1(n10934), .B2(keyinput2), 
        .ZN(n10933) );
  OAI221_X1 U13671 ( .B1(n10935), .B2(keyinput91), .C1(n10934), .C2(keyinput2), 
        .A(n10933), .ZN(n10939) );
  XNOR2_X1 U13672 ( .A(P3_ADDR_REG_13__SCAN_IN), .B(keyinput25), .ZN(n10937)
         );
  XNOR2_X1 U13673 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(keyinput15), .ZN(n10936)
         );
  NAND2_X1 U13674 ( .A1(n10937), .A2(n10936), .ZN(n10938) );
  NOR4_X1 U13675 ( .A1(n10941), .A2(n10940), .A3(n10939), .A4(n10938), .ZN(
        n10980) );
  INV_X1 U13676 ( .A(P3_REG3_REG_23__SCAN_IN), .ZN(n10943) );
  AOI22_X1 U13677 ( .A1(n10943), .A2(keyinput40), .B1(n14890), .B2(keyinput1), 
        .ZN(n10942) );
  OAI221_X1 U13678 ( .B1(n10943), .B2(keyinput40), .C1(n14890), .C2(keyinput1), 
        .A(n10942), .ZN(n10953) );
  AOI22_X1 U13679 ( .A1(n10945), .A2(keyinput65), .B1(keyinput61), .B2(n13844), 
        .ZN(n10944) );
  OAI221_X1 U13680 ( .B1(n10945), .B2(keyinput65), .C1(n13844), .C2(keyinput61), .A(n10944), .ZN(n10952) );
  AOI22_X1 U13681 ( .A1(n13517), .A2(keyinput38), .B1(n10947), .B2(keyinput75), 
        .ZN(n10946) );
  OAI221_X1 U13682 ( .B1(n13517), .B2(keyinput38), .C1(n10947), .C2(keyinput75), .A(n10946), .ZN(n10951) );
  XNOR2_X1 U13683 ( .A(P2_REG3_REG_13__SCAN_IN), .B(keyinput78), .ZN(n10949)
         );
  XNOR2_X1 U13684 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(keyinput64), .ZN(n10948)
         );
  NAND2_X1 U13685 ( .A1(n10949), .A2(n10948), .ZN(n10950) );
  NOR4_X1 U13686 ( .A1(n10953), .A2(n10952), .A3(n10951), .A4(n10950), .ZN(
        n10979) );
  INV_X1 U13687 ( .A(P1_D_REG_27__SCAN_IN), .ZN(n15817) );
  AOI22_X1 U13688 ( .A1(n15817), .A2(keyinput111), .B1(n11429), .B2(keyinput62), .ZN(n10954) );
  OAI221_X1 U13689 ( .B1(n15817), .B2(keyinput111), .C1(n11429), .C2(
        keyinput62), .A(n10954), .ZN(n10963) );
  AOI22_X1 U13690 ( .A1(n10956), .A2(keyinput124), .B1(keyinput97), .B2(n14981), .ZN(n10955) );
  OAI221_X1 U13691 ( .B1(n10956), .B2(keyinput124), .C1(n14981), .C2(
        keyinput97), .A(n10955), .ZN(n10962) );
  XNOR2_X1 U13692 ( .A(SI_4_), .B(keyinput26), .ZN(n10960) );
  XNOR2_X1 U13693 ( .A(P3_REG0_REG_23__SCAN_IN), .B(keyinput85), .ZN(n10959)
         );
  XNOR2_X1 U13694 ( .A(P3_REG1_REG_23__SCAN_IN), .B(keyinput69), .ZN(n10958)
         );
  XNOR2_X1 U13695 ( .A(P2_IR_REG_24__SCAN_IN), .B(keyinput126), .ZN(n10957) );
  NAND4_X1 U13696 ( .A1(n10960), .A2(n10959), .A3(n10958), .A4(n10957), .ZN(
        n10961) );
  NOR3_X1 U13697 ( .A1(n10963), .A2(n10962), .A3(n10961), .ZN(n10978) );
  XNOR2_X1 U13698 ( .A(n10964), .B(keyinput88), .ZN(n10969) );
  XOR2_X1 U13699 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(keyinput33), .Z(n10968) );
  XNOR2_X1 U13700 ( .A(n11307), .B(keyinput114), .ZN(n10967) );
  XNOR2_X1 U13701 ( .A(n10965), .B(keyinput108), .ZN(n10966) );
  NOR4_X1 U13702 ( .A1(n10969), .A2(n10968), .A3(n10967), .A4(n10966), .ZN(
        n10974) );
  XOR2_X1 U13703 ( .A(n10970), .B(keyinput17), .Z(n10973) );
  XNOR2_X1 U13704 ( .A(P2_IR_REG_0__SCAN_IN), .B(keyinput11), .ZN(n10972) );
  XNOR2_X1 U13705 ( .A(P2_IR_REG_2__SCAN_IN), .B(keyinput104), .ZN(n10971) );
  NAND4_X1 U13706 ( .A1(n10974), .A2(n10973), .A3(n10972), .A4(n10971), .ZN(
        n10976) );
  INV_X1 U13707 ( .A(P1_D_REG_16__SCAN_IN), .ZN(n15819) );
  XNOR2_X1 U13708 ( .A(n15819), .B(keyinput98), .ZN(n10975) );
  NOR2_X1 U13709 ( .A1(n10976), .A2(n10975), .ZN(n10977) );
  NAND4_X1 U13710 ( .A1(n10980), .A2(n10979), .A3(n10978), .A4(n10977), .ZN(
        n11029) );
  AOI22_X1 U13711 ( .A1(n16101), .A2(keyinput28), .B1(keyinput101), .B2(n9611), 
        .ZN(n10981) );
  OAI221_X1 U13712 ( .B1(n16101), .B2(keyinput28), .C1(n9611), .C2(keyinput101), .A(n10981), .ZN(n10991) );
  AOI22_X1 U13713 ( .A1(n9607), .A2(keyinput0), .B1(n10983), .B2(keyinput60), 
        .ZN(n10982) );
  OAI221_X1 U13714 ( .B1(n9607), .B2(keyinput0), .C1(n10983), .C2(keyinput60), 
        .A(n10982), .ZN(n10990) );
  AOI22_X1 U13715 ( .A1(n10985), .A2(keyinput12), .B1(n12578), .B2(keyinput9), 
        .ZN(n10984) );
  OAI221_X1 U13716 ( .B1(n10985), .B2(keyinput12), .C1(n12578), .C2(keyinput9), 
        .A(n10984), .ZN(n10989) );
  XNOR2_X1 U13717 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(keyinput112), .ZN(n10987)
         );
  XNOR2_X1 U13718 ( .A(P1_ADDR_REG_2__SCAN_IN), .B(keyinput50), .ZN(n10986) );
  NAND2_X1 U13719 ( .A1(n10987), .A2(n10986), .ZN(n10988) );
  NOR4_X1 U13720 ( .A1(n10991), .A2(n10990), .A3(n10989), .A4(n10988), .ZN(
        n11027) );
  AOI22_X1 U13721 ( .A1(n10993), .A2(keyinput118), .B1(keyinput110), .B2(
        n15100), .ZN(n10992) );
  OAI221_X1 U13722 ( .B1(n10993), .B2(keyinput118), .C1(n15100), .C2(
        keyinput110), .A(n10992), .ZN(n11002) );
  AOI22_X1 U13723 ( .A1(keyinput74), .A2(n10995), .B1(keyinput90), .B2(n10608), 
        .ZN(n10994) );
  OAI21_X1 U13724 ( .B1(n10995), .B2(keyinput74), .A(n10994), .ZN(n11001) );
  AOI22_X1 U13725 ( .A1(n8204), .A2(keyinput3), .B1(keyinput34), .B2(n14464), 
        .ZN(n10996) );
  OAI221_X1 U13726 ( .B1(n8204), .B2(keyinput3), .C1(n14464), .C2(keyinput34), 
        .A(n10996), .ZN(n11000) );
  XNOR2_X1 U13727 ( .A(P1_REG1_REG_20__SCAN_IN), .B(keyinput44), .ZN(n10998)
         );
  XNOR2_X1 U13728 ( .A(P1_IR_REG_0__SCAN_IN), .B(keyinput31), .ZN(n10997) );
  NAND2_X1 U13729 ( .A1(n10998), .A2(n10997), .ZN(n10999) );
  NOR4_X1 U13730 ( .A1(n11002), .A2(n11001), .A3(n11000), .A4(n10999), .ZN(
        n11026) );
  INV_X1 U13731 ( .A(P2_D_REG_30__SCAN_IN), .ZN(n15947) );
  AOI22_X1 U13732 ( .A1(n15947), .A2(keyinput56), .B1(keyinput77), .B2(n12846), 
        .ZN(n11003) );
  OAI221_X1 U13733 ( .B1(n15947), .B2(keyinput56), .C1(n12846), .C2(keyinput77), .A(n11003), .ZN(n11012) );
  AOI22_X1 U13734 ( .A1(n9008), .A2(keyinput48), .B1(keyinput20), .B2(n11556), 
        .ZN(n11004) );
  OAI221_X1 U13735 ( .B1(n9008), .B2(keyinput48), .C1(n11556), .C2(keyinput20), 
        .A(n11004), .ZN(n11011) );
  INV_X1 U13736 ( .A(P2_REG2_REG_31__SCAN_IN), .ZN(n11006) );
  AOI22_X1 U13737 ( .A1(n11006), .A2(keyinput30), .B1(n11971), .B2(keyinput87), 
        .ZN(n11005) );
  OAI221_X1 U13738 ( .B1(n11006), .B2(keyinput30), .C1(n11971), .C2(keyinput87), .A(n11005), .ZN(n11010) );
  XNOR2_X1 U13739 ( .A(P3_REG2_REG_26__SCAN_IN), .B(keyinput119), .ZN(n11008)
         );
  XNOR2_X1 U13740 ( .A(P1_IR_REG_1__SCAN_IN), .B(keyinput59), .ZN(n11007) );
  NAND2_X1 U13741 ( .A1(n11008), .A2(n11007), .ZN(n11009) );
  NOR4_X1 U13742 ( .A1(n11012), .A2(n11011), .A3(n11010), .A4(n11009), .ZN(
        n11025) );
  AOI22_X1 U13743 ( .A1(n12507), .A2(keyinput4), .B1(keyinput76), .B2(n12095), 
        .ZN(n11013) );
  OAI221_X1 U13744 ( .B1(n12507), .B2(keyinput4), .C1(n12095), .C2(keyinput76), 
        .A(n11013), .ZN(n11023) );
  INV_X1 U13745 ( .A(P1_REG2_REG_23__SCAN_IN), .ZN(n11015) );
  AOI22_X1 U13746 ( .A1(n11016), .A2(keyinput106), .B1(n11015), .B2(keyinput23), .ZN(n11014) );
  OAI221_X1 U13747 ( .B1(n11016), .B2(keyinput106), .C1(n11015), .C2(
        keyinput23), .A(n11014), .ZN(n11022) );
  XNOR2_X1 U13748 ( .A(P1_REG3_REG_22__SCAN_IN), .B(keyinput52), .ZN(n11020)
         );
  XNOR2_X1 U13749 ( .A(P3_IR_REG_8__SCAN_IN), .B(keyinput13), .ZN(n11019) );
  XNOR2_X1 U13750 ( .A(P2_IR_REG_13__SCAN_IN), .B(keyinput42), .ZN(n11018) );
  XNOR2_X1 U13751 ( .A(P1_REG1_REG_25__SCAN_IN), .B(keyinput122), .ZN(n11017)
         );
  NAND4_X1 U13752 ( .A1(n11020), .A2(n11019), .A3(n11018), .A4(n11017), .ZN(
        n11021) );
  NOR3_X1 U13753 ( .A1(n11023), .A2(n11022), .A3(n11021), .ZN(n11024) );
  NAND4_X1 U13754 ( .A1(n11027), .A2(n11026), .A3(n11025), .A4(n11024), .ZN(
        n11028) );
  NOR4_X1 U13755 ( .A1(n11031), .A2(n11030), .A3(n11029), .A4(n11028), .ZN(
        n11032) );
  OAI221_X1 U13756 ( .B1(n10608), .B2(keyinput90), .C1(n10608), .C2(n11033), 
        .A(n11032), .ZN(n11034) );
  XNOR2_X1 U13757 ( .A(n11035), .B(n11034), .ZN(P3_U3492) );
  INV_X1 U13758 ( .A(n11036), .ZN(n11040) );
  INV_X1 U13759 ( .A(n15178), .ZN(n11037) );
  OAI222_X1 U13760 ( .A1(n15700), .A2(n11038), .B1(n15703), .B2(n11040), .C1(
        n11037), .C2(P1_U3086), .ZN(P1_U3345) );
  INV_X1 U13761 ( .A(n11238), .ZN(n11039) );
  OAI222_X1 U13762 ( .A1(n14914), .A2(n11041), .B1(n14917), .B2(n11040), .C1(
        P2_U3088), .C2(n11039), .ZN(P2_U3317) );
  NAND2_X1 U13763 ( .A1(n11043), .A2(n11042), .ZN(n11048) );
  INV_X1 U13764 ( .A(n11044), .ZN(n11046) );
  NAND2_X1 U13765 ( .A1(n11046), .A2(n11045), .ZN(n11047) );
  OAI21_X1 U13766 ( .B1(n11050), .B2(P1_ADDR_REG_5__SCAN_IN), .A(n11049), .ZN(
        n11334) );
  XNOR2_X1 U13767 ( .A(P1_ADDR_REG_6__SCAN_IN), .B(P3_ADDR_REG_6__SCAN_IN), 
        .ZN(n11051) );
  XNOR2_X1 U13768 ( .A(n11334), .B(n11051), .ZN(n11052) );
  NAND2_X1 U13769 ( .A1(n11053), .A2(n11052), .ZN(n11342) );
  OAI21_X1 U13770 ( .B1(n11053), .B2(n11052), .A(n11342), .ZN(n11054) );
  INV_X1 U13771 ( .A(n11054), .ZN(SUB_1596_U57) );
  OAI222_X1 U13772 ( .A1(P3_U3151), .A2(n13543), .B1(n13962), .B2(n11056), 
        .C1(n13102), .C2(n11055), .ZN(P3_U3282) );
  INV_X1 U13773 ( .A(n11057), .ZN(n11060) );
  INV_X1 U13774 ( .A(n11522), .ZN(n11219) );
  OAI222_X1 U13775 ( .A1(n14914), .A2(n11058), .B1(n14917), .B2(n11060), .C1(
        P2_U3088), .C2(n11219), .ZN(P2_U3316) );
  INV_X1 U13776 ( .A(n11557), .ZN(n11059) );
  OAI222_X1 U13777 ( .A1(n15700), .A2(n11061), .B1(n15703), .B2(n11060), .C1(
        n11059), .C2(P1_U3086), .ZN(P1_U3344) );
  MUX2_X1 U13778 ( .A(n9560), .B(P1_REG1_REG_5__SCAN_IN), .S(n11097), .Z(
        n11070) );
  MUX2_X1 U13779 ( .A(P1_REG1_REG_2__SCAN_IN), .B(n9508), .S(n15124), .Z(
        n15127) );
  INV_X1 U13780 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n11498) );
  MUX2_X1 U13781 ( .A(P1_REG1_REG_1__SCAN_IN), .B(n11498), .S(n15103), .Z(
        n15108) );
  AND2_X1 U13782 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), 
        .ZN(n15107) );
  NAND2_X1 U13783 ( .A1(n15108), .A2(n15107), .ZN(n15106) );
  NAND2_X1 U13784 ( .A1(n15103), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n11062) );
  NAND2_X1 U13785 ( .A1(n15106), .A2(n11062), .ZN(n15126) );
  NAND2_X1 U13786 ( .A1(n15127), .A2(n15126), .ZN(n15125) );
  NAND2_X1 U13787 ( .A1(n15124), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n11063) );
  NAND2_X1 U13788 ( .A1(n15125), .A2(n11063), .ZN(n15138) );
  XNOR2_X1 U13789 ( .A(n15136), .B(n11064), .ZN(n15139) );
  NAND2_X1 U13790 ( .A1(n15138), .A2(n15139), .ZN(n15137) );
  NAND2_X1 U13791 ( .A1(n15136), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n11065) );
  NAND2_X1 U13792 ( .A1(n15137), .A2(n11065), .ZN(n15154) );
  XNOR2_X1 U13793 ( .A(n11079), .B(n11066), .ZN(n15155) );
  NAND2_X1 U13794 ( .A1(n15154), .A2(n15155), .ZN(n15153) );
  NAND2_X1 U13795 ( .A1(n11079), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n11067) );
  NAND2_X1 U13796 ( .A1(n15153), .A2(n11067), .ZN(n11069) );
  OR2_X1 U13797 ( .A1(n11069), .A2(n11070), .ZN(n11090) );
  INV_X1 U13798 ( .A(n11090), .ZN(n11068) );
  AOI21_X1 U13799 ( .B1(n11070), .B2(n11069), .A(n11068), .ZN(n11087) );
  INV_X1 U13800 ( .A(n11082), .ZN(n11072) );
  OR2_X1 U13801 ( .A1(n11072), .A2(n11071), .ZN(n15246) );
  INV_X1 U13802 ( .A(n15246), .ZN(n15223) );
  NAND2_X1 U13803 ( .A1(P1_REG3_REG_5__SCAN_IN), .A2(P1_U3086), .ZN(n12088) );
  OAI21_X1 U13804 ( .B1(n15252), .B2(n10678), .A(n12088), .ZN(n11073) );
  AOI21_X1 U13805 ( .B1(n15223), .B2(n11097), .A(n11073), .ZN(n11086) );
  MUX2_X1 U13806 ( .A(P1_REG2_REG_5__SCAN_IN), .B(n9561), .S(n11097), .Z(
        n11084) );
  INV_X1 U13807 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n11851) );
  MUX2_X1 U13808 ( .A(P1_REG2_REG_2__SCAN_IN), .B(n11851), .S(n15124), .Z(
        n15130) );
  INV_X1 U13809 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n11833) );
  MUX2_X1 U13810 ( .A(P1_REG2_REG_1__SCAN_IN), .B(n11833), .S(n15103), .Z(
        n15105) );
  AND2_X1 U13811 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n15112) );
  NAND2_X1 U13812 ( .A1(n15105), .A2(n15112), .ZN(n15104) );
  NAND2_X1 U13813 ( .A1(n15103), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n11074) );
  NAND2_X1 U13814 ( .A1(n15104), .A2(n11074), .ZN(n15129) );
  NAND2_X1 U13815 ( .A1(n15130), .A2(n15129), .ZN(n15128) );
  NAND2_X1 U13816 ( .A1(n15124), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n11075) );
  NAND2_X1 U13817 ( .A1(n15128), .A2(n11075), .ZN(n15141) );
  INV_X1 U13818 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n11076) );
  XNOR2_X1 U13819 ( .A(n15136), .B(n11076), .ZN(n15142) );
  NAND2_X1 U13820 ( .A1(n15141), .A2(n15142), .ZN(n15140) );
  NAND2_X1 U13821 ( .A1(n15136), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n11077) );
  NAND2_X1 U13822 ( .A1(n15140), .A2(n11077), .ZN(n15151) );
  INV_X1 U13823 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n11078) );
  XNOR2_X1 U13824 ( .A(n11079), .B(n11078), .ZN(n15152) );
  NAND2_X1 U13825 ( .A1(n15151), .A2(n15152), .ZN(n15150) );
  NAND2_X1 U13826 ( .A1(n11079), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n11080) );
  NAND2_X1 U13827 ( .A1(n15150), .A2(n11080), .ZN(n11083) );
  NOR2_X1 U13828 ( .A1(n15119), .A2(n15699), .ZN(n11081) );
  NAND2_X1 U13829 ( .A1(n11083), .A2(n11084), .ZN(n11099) );
  OAI211_X1 U13830 ( .C1(n11084), .C2(n11083), .A(n15244), .B(n11099), .ZN(
        n11085) );
  OAI211_X1 U13831 ( .C1(n11087), .C2(n15248), .A(n11086), .B(n11085), .ZN(
        P1_U3248) );
  XNOR2_X1 U13832 ( .A(n11370), .B(n11088), .ZN(n11360) );
  OR2_X1 U13833 ( .A1(n11097), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n11089) );
  INV_X1 U13834 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n11091) );
  MUX2_X1 U13835 ( .A(n11091), .B(P1_REG1_REG_6__SCAN_IN), .S(n11201), .Z(
        n11198) );
  NAND2_X1 U13836 ( .A1(n11201), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n11092) );
  MUX2_X1 U13837 ( .A(P1_REG1_REG_7__SCAN_IN), .B(n9593), .S(n15163), .Z(
        n15169) );
  NAND2_X1 U13838 ( .A1(n15163), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n11093) );
  NAND2_X1 U13839 ( .A1(n15167), .A2(n11093), .ZN(n11112) );
  MUX2_X1 U13840 ( .A(n9607), .B(P1_REG1_REG_8__SCAN_IN), .S(n11116), .Z(
        n11113) );
  OR2_X1 U13841 ( .A1(n11116), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n11094) );
  XOR2_X1 U13842 ( .A(n11360), .B(n11361), .Z(n11109) );
  INV_X1 U13843 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n12008) );
  NAND2_X1 U13844 ( .A1(P1_REG3_REG_9__SCAN_IN), .A2(P1_U3086), .ZN(n11095) );
  OAI21_X1 U13845 ( .B1(n15252), .B2(n12008), .A(n11095), .ZN(n11096) );
  AOI21_X1 U13846 ( .B1(n15223), .B2(n11370), .A(n11096), .ZN(n11108) );
  NAND2_X1 U13847 ( .A1(n11097), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n11098) );
  NAND2_X1 U13848 ( .A1(n11099), .A2(n11098), .ZN(n11203) );
  XNOR2_X1 U13849 ( .A(n11201), .B(n12036), .ZN(n11204) );
  NAND2_X1 U13850 ( .A1(n11203), .A2(n11204), .ZN(n11202) );
  NAND2_X1 U13851 ( .A1(n11201), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n11100) );
  NAND2_X1 U13852 ( .A1(n11202), .A2(n11100), .ZN(n15165) );
  MUX2_X1 U13853 ( .A(P1_REG2_REG_7__SCAN_IN), .B(n9590), .S(n15163), .Z(
        n15166) );
  NAND2_X1 U13854 ( .A1(n15165), .A2(n15166), .ZN(n15164) );
  NAND2_X1 U13855 ( .A1(n15163), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n11101) );
  NAND2_X1 U13856 ( .A1(n15164), .A2(n11101), .ZN(n11118) );
  INV_X1 U13857 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n11102) );
  MUX2_X1 U13858 ( .A(P1_REG2_REG_8__SCAN_IN), .B(n11102), .S(n11116), .Z(
        n11119) );
  NAND2_X1 U13859 ( .A1(n11118), .A2(n11119), .ZN(n11117) );
  NAND2_X1 U13860 ( .A1(n11116), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n11103) );
  NAND2_X1 U13861 ( .A1(n11117), .A2(n11103), .ZN(n11106) );
  INV_X1 U13862 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n11104) );
  MUX2_X1 U13863 ( .A(P1_REG2_REG_9__SCAN_IN), .B(n11104), .S(n11370), .Z(
        n11105) );
  NAND2_X1 U13864 ( .A1(n11106), .A2(n11105), .ZN(n11372) );
  OAI211_X1 U13865 ( .C1(n11106), .C2(n11105), .A(n11372), .B(n15244), .ZN(
        n11107) );
  OAI211_X1 U13866 ( .C1(n11109), .C2(n15248), .A(n11108), .B(n11107), .ZN(
        P1_U3252) );
  INV_X1 U13867 ( .A(n11110), .ZN(n11111) );
  AOI21_X1 U13868 ( .B1(n11113), .B2(n11112), .A(n11111), .ZN(n11122) );
  INV_X1 U13869 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n11114) );
  NAND2_X1 U13870 ( .A1(P1_REG3_REG_8__SCAN_IN), .A2(P1_U3086), .ZN(n12411) );
  OAI21_X1 U13871 ( .B1(n15252), .B2(n11114), .A(n12411), .ZN(n11115) );
  AOI21_X1 U13872 ( .B1(n15223), .B2(n11116), .A(n11115), .ZN(n11121) );
  OAI211_X1 U13873 ( .C1(n11119), .C2(n11118), .A(n15244), .B(n11117), .ZN(
        n11120) );
  OAI211_X1 U13874 ( .C1(n11122), .C2(n15248), .A(n11121), .B(n11120), .ZN(
        P1_U3251) );
  INV_X1 U13875 ( .A(n11123), .ZN(n11124) );
  OAI222_X1 U13876 ( .A1(P3_U3151), .A2(n11126), .B1(n13970), .B2(n11125), 
        .C1(n13102), .C2(n11124), .ZN(P3_U3280) );
  OAI222_X1 U13877 ( .A1(P3_U3151), .A2(n11129), .B1(n13962), .B2(n11128), 
        .C1(n13102), .C2(n11127), .ZN(P3_U3281) );
  XNOR2_X1 U13878 ( .A(n11221), .B(P2_REG1_REG_9__SCAN_IN), .ZN(n11145) );
  INV_X1 U13879 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n11130) );
  MUX2_X1 U13880 ( .A(P2_REG1_REG_2__SCAN_IN), .B(n11130), .S(n11158), .Z(
        n15902) );
  INV_X1 U13881 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n11131) );
  MUX2_X1 U13882 ( .A(P2_REG1_REG_1__SCAN_IN), .B(n11131), .S(n11155), .Z(
        n15889) );
  AND2_X1 U13883 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), 
        .ZN(n15888) );
  NAND2_X1 U13884 ( .A1(n15889), .A2(n15888), .ZN(n11133) );
  NAND2_X1 U13885 ( .A1(n11155), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n11132) );
  NAND2_X1 U13886 ( .A1(n11133), .A2(n11132), .ZN(n15901) );
  NAND2_X1 U13887 ( .A1(n15902), .A2(n15901), .ZN(n15900) );
  NAND2_X1 U13888 ( .A1(n11158), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n11134) );
  NAND2_X1 U13889 ( .A1(n15900), .A2(n11134), .ZN(n14426) );
  INV_X1 U13890 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n11712) );
  MUX2_X1 U13891 ( .A(P2_REG1_REG_3__SCAN_IN), .B(n11712), .S(n14428), .Z(
        n14427) );
  NAND2_X1 U13892 ( .A1(n14426), .A2(n14427), .ZN(n14425) );
  NAND2_X1 U13893 ( .A1(n14428), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n11135) );
  NAND2_X1 U13894 ( .A1(n14425), .A2(n11135), .ZN(n14438) );
  INV_X1 U13895 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n11823) );
  MUX2_X1 U13896 ( .A(P2_REG1_REG_4__SCAN_IN), .B(n11823), .S(n14440), .Z(
        n14439) );
  NAND2_X1 U13897 ( .A1(n14438), .A2(n14439), .ZN(n14437) );
  NAND2_X1 U13898 ( .A1(n14440), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n11136) );
  NAND2_X1 U13899 ( .A1(n14437), .A2(n11136), .ZN(n14458) );
  INV_X1 U13900 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n16005) );
  MUX2_X1 U13901 ( .A(P2_REG1_REG_5__SCAN_IN), .B(n16005), .S(n14451), .Z(
        n14459) );
  NAND2_X1 U13902 ( .A1(n14458), .A2(n14459), .ZN(n14457) );
  NAND2_X1 U13903 ( .A1(n14451), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n11137) );
  NAND2_X1 U13904 ( .A1(n14457), .A2(n11137), .ZN(n15914) );
  INV_X1 U13905 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n11138) );
  XNOR2_X1 U13906 ( .A(n11168), .B(n11138), .ZN(n15915) );
  NAND2_X1 U13907 ( .A1(n15914), .A2(n15915), .ZN(n15913) );
  NAND2_X1 U13908 ( .A1(n11168), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n11139) );
  NAND2_X1 U13909 ( .A1(n15913), .A2(n11139), .ZN(n14468) );
  INV_X1 U13910 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n16009) );
  MUX2_X1 U13911 ( .A(P2_REG1_REG_7__SCAN_IN), .B(n16009), .S(n14470), .Z(
        n14469) );
  NAND2_X1 U13912 ( .A1(n14468), .A2(n14469), .ZN(n14467) );
  NAND2_X1 U13913 ( .A1(n14470), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n11140) );
  NAND2_X1 U13914 ( .A1(n14467), .A2(n11140), .ZN(n14482) );
  XNOR2_X1 U13915 ( .A(n14484), .B(n11141), .ZN(n14483) );
  NAND2_X1 U13916 ( .A1(n14482), .A2(n14483), .ZN(n14481) );
  NAND2_X1 U13917 ( .A1(n14484), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n11142) );
  NAND2_X1 U13918 ( .A1(n14481), .A2(n11142), .ZN(n11144) );
  INV_X1 U13919 ( .A(n11223), .ZN(n11143) );
  AOI21_X1 U13920 ( .B1(n11145), .B2(n11144), .A(n11143), .ZN(n11187) );
  INV_X1 U13921 ( .A(n12320), .ZN(n11149) );
  OAI21_X1 U13922 ( .B1(n11147), .B2(n11149), .A(n11146), .ZN(n11148) );
  OAI21_X1 U13923 ( .B1(n11150), .B2(n11149), .A(n11148), .ZN(n11181) );
  NAND2_X1 U13924 ( .A1(n11151), .A2(P2_STATE_REG_SCAN_IN), .ZN(n14908) );
  INV_X1 U13925 ( .A(n14912), .ZN(n14377) );
  NOR2_X1 U13926 ( .A1(n14908), .A2(n14377), .ZN(n11152) );
  NAND2_X1 U13927 ( .A1(n11181), .A2(n11152), .ZN(n15904) );
  NOR2_X1 U13928 ( .A1(n14908), .A2(n14912), .ZN(n11153) );
  NAND2_X1 U13929 ( .A1(n11181), .A2(n11153), .ZN(n14504) );
  MUX2_X1 U13930 ( .A(P2_REG2_REG_1__SCAN_IN), .B(n11154), .S(n11155), .Z(
        n15894) );
  AND2_X1 U13931 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), 
        .ZN(n15895) );
  NAND2_X1 U13932 ( .A1(n15894), .A2(n15895), .ZN(n15893) );
  NAND2_X1 U13933 ( .A1(n11155), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n11156) );
  NAND2_X1 U13934 ( .A1(n15893), .A2(n11156), .ZN(n15908) );
  MUX2_X1 U13935 ( .A(P2_REG2_REG_2__SCAN_IN), .B(n11157), .S(n11158), .Z(
        n15909) );
  NAND2_X1 U13936 ( .A1(n15908), .A2(n15909), .ZN(n15907) );
  NAND2_X1 U13937 ( .A1(n11158), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n14430) );
  NAND2_X1 U13938 ( .A1(n15907), .A2(n14430), .ZN(n11161) );
  MUX2_X1 U13939 ( .A(P2_REG2_REG_3__SCAN_IN), .B(n11159), .S(n14428), .Z(
        n11160) );
  NAND2_X1 U13940 ( .A1(n14428), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n14442) );
  NAND2_X1 U13941 ( .A1(n14443), .A2(n14442), .ZN(n11164) );
  MUX2_X1 U13942 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n11162), .S(n14440), .Z(
        n11163) );
  NAND2_X1 U13943 ( .A1(n14440), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n14453) );
  NAND2_X1 U13944 ( .A1(n14454), .A2(n14453), .ZN(n11166) );
  INV_X1 U13945 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n12224) );
  MUX2_X1 U13946 ( .A(P2_REG2_REG_5__SCAN_IN), .B(n12224), .S(n14451), .Z(
        n11165) );
  NAND2_X1 U13947 ( .A1(n11166), .A2(n11165), .ZN(n14456) );
  NAND2_X1 U13948 ( .A1(n14451), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n11167) );
  NAND2_X1 U13949 ( .A1(n14456), .A2(n11167), .ZN(n15922) );
  MUX2_X1 U13950 ( .A(P2_REG2_REG_6__SCAN_IN), .B(n10956), .S(n11168), .Z(
        n15923) );
  NAND2_X1 U13951 ( .A1(n11168), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n14472) );
  MUX2_X1 U13952 ( .A(P2_REG2_REG_7__SCAN_IN), .B(n12238), .S(n14470), .Z(
        n11169) );
  NAND2_X1 U13953 ( .A1(n14470), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n14486) );
  INV_X1 U13954 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n11170) );
  MUX2_X1 U13955 ( .A(P2_REG2_REG_8__SCAN_IN), .B(n11170), .S(n14484), .Z(
        n11171) );
  NAND2_X1 U13956 ( .A1(n11172), .A2(n11171), .ZN(n14489) );
  NAND2_X1 U13957 ( .A1(n14484), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n11173) );
  NAND2_X1 U13958 ( .A1(n14489), .A2(n11173), .ZN(n11176) );
  INV_X1 U13959 ( .A(n11176), .ZN(n11178) );
  INV_X1 U13960 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n11174) );
  MUX2_X1 U13961 ( .A(P2_REG2_REG_9__SCAN_IN), .B(n11174), .S(n11221), .Z(
        n11177) );
  MUX2_X1 U13962 ( .A(n11174), .B(P2_REG2_REG_9__SCAN_IN), .S(n11221), .Z(
        n11175) );
  OAI21_X1 U13963 ( .B1(n11178), .B2(n11177), .A(n11213), .ZN(n11185) );
  AND2_X1 U13964 ( .A1(n11179), .A2(P2_STATE_REG_SCAN_IN), .ZN(n11180) );
  NAND2_X1 U13965 ( .A1(n11181), .A2(n11180), .ZN(n15919) );
  OR2_X1 U13966 ( .A1(n11181), .A2(P2_U3088), .ZN(n15944) );
  INV_X1 U13967 ( .A(n15944), .ZN(n15899) );
  NAND2_X1 U13968 ( .A1(n15899), .A2(P2_ADDR_REG_9__SCAN_IN), .ZN(n11182) );
  NAND2_X1 U13969 ( .A1(P2_U3088), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n12430) );
  OAI211_X1 U13970 ( .C1(n15919), .C2(n11183), .A(n11182), .B(n12430), .ZN(
        n11184) );
  AOI21_X1 U13971 ( .B1(n15937), .B2(n11185), .A(n11184), .ZN(n11186) );
  OAI21_X1 U13972 ( .B1(n11187), .B2(n15904), .A(n11186), .ZN(P2_U3223) );
  INV_X1 U13973 ( .A(n15904), .ZN(n15928) );
  AOI22_X1 U13974 ( .A1(P2_REG1_REG_0__SCAN_IN), .A2(n15928), .B1(n15937), 
        .B2(P2_REG2_REG_0__SCAN_IN), .ZN(n11191) );
  INV_X1 U13975 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n11189) );
  NOR2_X1 U13976 ( .A1(n14504), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n11188) );
  AOI211_X1 U13977 ( .C1(n15928), .C2(n11189), .A(n15936), .B(n11188), .ZN(
        n11190) );
  MUX2_X1 U13978 ( .A(n11191), .B(n11190), .S(P2_IR_REG_0__SCAN_IN), .Z(n11193) );
  AOI22_X1 U13979 ( .A1(n15899), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3088), .ZN(n11192) );
  NAND2_X1 U13980 ( .A1(n11193), .A2(n11192), .ZN(P2_U3214) );
  INV_X1 U13981 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n11332) );
  NAND2_X1 U13982 ( .A1(P1_REG3_REG_6__SCAN_IN), .A2(P1_U3086), .ZN(n11194) );
  OAI21_X1 U13983 ( .B1(n15252), .B2(n11332), .A(n11194), .ZN(n11200) );
  INV_X1 U13984 ( .A(n11195), .ZN(n11196) );
  AOI211_X1 U13985 ( .C1(n11198), .C2(n11197), .A(n11196), .B(n15248), .ZN(
        n11199) );
  AOI211_X1 U13986 ( .C1(n15223), .C2(n11201), .A(n11200), .B(n11199), .ZN(
        n11206) );
  OAI211_X1 U13987 ( .C1(n11204), .C2(n11203), .A(n15244), .B(n11202), .ZN(
        n11205) );
  NAND2_X1 U13988 ( .A1(n11206), .A2(n11205), .ZN(P1_U3249) );
  INV_X1 U13989 ( .A(n11207), .ZN(n11258) );
  INV_X1 U13990 ( .A(n15700), .ZN(n15691) );
  AOI22_X1 U13991 ( .A1(n11895), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(n15691), .ZN(n11208) );
  OAI21_X1 U13992 ( .B1(n11258), .B2(n15703), .A(n11208), .ZN(P1_U3343) );
  INV_X1 U13993 ( .A(n11209), .ZN(n11210) );
  OAI222_X1 U13994 ( .A1(P3_U3151), .A2(n7640), .B1(n13970), .B2(n11211), .C1(
        n13102), .C2(n11210), .ZN(P3_U3279) );
  OR2_X1 U13995 ( .A1(n11221), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n11212) );
  MUX2_X1 U13996 ( .A(n8204), .B(P2_REG2_REG_10__SCAN_IN), .S(n11238), .Z(
        n11236) );
  NAND2_X1 U13997 ( .A1(n11238), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n11214) );
  INV_X1 U13998 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n11215) );
  MUX2_X1 U13999 ( .A(n11215), .B(P2_REG2_REG_11__SCAN_IN), .S(n11522), .Z(
        n11217) );
  INV_X1 U14000 ( .A(n11528), .ZN(n11216) );
  AOI21_X1 U14001 ( .B1(n11218), .B2(n11217), .A(n11216), .ZN(n11229) );
  NAND2_X1 U14002 ( .A1(P2_U3088), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n12874)
         );
  OAI21_X1 U14003 ( .B1(n15919), .B2(n11219), .A(n12874), .ZN(n11220) );
  AOI21_X1 U14004 ( .B1(n15899), .B2(P2_ADDR_REG_11__SCAN_IN), .A(n11220), 
        .ZN(n11228) );
  OR2_X1 U14005 ( .A1(n11221), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n11222) );
  NAND2_X1 U14006 ( .A1(n11223), .A2(n11222), .ZN(n11232) );
  XNOR2_X1 U14007 ( .A(n11238), .B(P2_REG1_REG_10__SCAN_IN), .ZN(n11233) );
  NAND2_X1 U14008 ( .A1(n11238), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n11224) );
  NAND2_X1 U14009 ( .A1(n11230), .A2(n11224), .ZN(n11226) );
  INV_X1 U14010 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n14838) );
  XNOR2_X1 U14011 ( .A(n11522), .B(n14838), .ZN(n11225) );
  NAND2_X1 U14012 ( .A1(n11226), .A2(n11225), .ZN(n11518) );
  OAI211_X1 U14013 ( .C1(n11226), .C2(n11225), .A(n11518), .B(n15928), .ZN(
        n11227) );
  OAI211_X1 U14014 ( .C1(n11229), .C2(n14504), .A(n11228), .B(n11227), .ZN(
        P2_U3225) );
  INV_X1 U14015 ( .A(n11230), .ZN(n11231) );
  AOI211_X1 U14016 ( .C1(n11233), .C2(n11232), .A(n15904), .B(n11231), .ZN(
        n11242) );
  INV_X1 U14017 ( .A(n11234), .ZN(n11235) );
  AOI211_X1 U14018 ( .C1(n11237), .C2(n11236), .A(n14504), .B(n11235), .ZN(
        n11241) );
  INV_X1 U14019 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n12325) );
  NAND2_X1 U14020 ( .A1(n15936), .A2(n11238), .ZN(n11239) );
  NAND2_X1 U14021 ( .A1(P2_U3088), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n12816)
         );
  OAI211_X1 U14022 ( .C1(n15944), .C2(n12325), .A(n11239), .B(n12816), .ZN(
        n11240) );
  OR3_X1 U14023 ( .A1(n11242), .A2(n11241), .A3(n11240), .ZN(P2_U3224) );
  OAI21_X1 U14024 ( .B1(P3_REG2_REG_5__SCAN_IN), .B2(n11244), .A(n11243), .ZN(
        n11249) );
  INV_X1 U14025 ( .A(n16014), .ZN(n13583) );
  OAI21_X1 U14026 ( .B1(P3_REG1_REG_5__SCAN_IN), .B2(n11245), .A(n11397), .ZN(
        n11246) );
  NAND2_X1 U14027 ( .A1(n11246), .A2(n13631), .ZN(n11247) );
  NAND2_X1 U14028 ( .A1(P3_U3151), .A2(P3_REG3_REG_5__SCAN_IN), .ZN(n11916) );
  OAI211_X1 U14029 ( .C1(n16024), .C2(n7495), .A(n11247), .B(n11916), .ZN(
        n11248) );
  AOI21_X1 U14030 ( .B1(n11249), .B2(n13583), .A(n11248), .ZN(n11257) );
  INV_X1 U14031 ( .A(n11250), .ZN(n11262) );
  INV_X1 U14032 ( .A(n11251), .ZN(n11253) );
  NOR3_X1 U14033 ( .A1(n11262), .A2(n11253), .A3(n11252), .ZN(n11255) );
  INV_X1 U14034 ( .A(n11388), .ZN(n11254) );
  INV_X1 U14035 ( .A(n16013), .ZN(n13537) );
  OAI21_X1 U14036 ( .B1(n11255), .B2(n11254), .A(n13537), .ZN(n11256) );
  OAI211_X1 U14037 ( .C1(n13617), .C2(n7646), .A(n11257), .B(n11256), .ZN(
        P3_U3187) );
  INV_X1 U14038 ( .A(n11523), .ZN(n11726) );
  OAI222_X1 U14039 ( .A1(n14914), .A2(n11259), .B1(n14917), .B2(n11258), .C1(
        n11726), .C2(P2_U3088), .ZN(P2_U3315) );
  NOR2_X1 U14040 ( .A1(n11261), .A2(n7407), .ZN(n11263) );
  AOI21_X1 U14041 ( .B1(n11263), .B2(n11327), .A(n11262), .ZN(n11280) );
  INV_X1 U14042 ( .A(n11264), .ZN(n11269) );
  NAND3_X1 U14043 ( .A1(n11265), .A2(n11267), .A3(n11266), .ZN(n11268) );
  AOI21_X1 U14044 ( .B1(n11269), .B2(n11268), .A(n16014), .ZN(n11277) );
  INV_X1 U14045 ( .A(P3_ADDR_REG_4__SCAN_IN), .ZN(n11275) );
  AND3_X1 U14046 ( .A1(n11320), .A2(n11271), .A3(n11270), .ZN(n11272) );
  OAI21_X1 U14047 ( .B1(n11273), .B2(n11272), .A(n13631), .ZN(n11274) );
  NAND2_X1 U14048 ( .A1(P3_U3151), .A2(P3_REG3_REG_4__SCAN_IN), .ZN(n11659) );
  OAI211_X1 U14049 ( .C1(n16024), .C2(n11275), .A(n11274), .B(n11659), .ZN(
        n11276) );
  AOI211_X1 U14050 ( .C1(n16021), .C2(n11278), .A(n11277), .B(n11276), .ZN(
        n11279) );
  OAI21_X1 U14051 ( .B1(n11280), .B2(n16013), .A(n11279), .ZN(P3_U3186) );
  INV_X1 U14052 ( .A(n15252), .ZN(n15149) );
  NOR2_X1 U14053 ( .A1(n15149), .A2(P1_U4016), .ZN(P1_U3085) );
  AOI21_X1 U14054 ( .B1(n11282), .B2(n16016), .A(n7401), .ZN(n11283) );
  OAI22_X1 U14055 ( .A1(n11283), .A2(n16013), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n11445), .ZN(n11292) );
  AOI21_X1 U14056 ( .B1(n16064), .B2(n11285), .A(n11284), .ZN(n11290) );
  OAI21_X1 U14057 ( .B1(P3_REG1_REG_1__SCAN_IN), .B2(n11287), .A(n11286), .ZN(
        n11288) );
  NAND2_X1 U14058 ( .A1(n13631), .A2(n11288), .ZN(n11289) );
  OAI21_X1 U14059 ( .B1(n11290), .B2(n16014), .A(n11289), .ZN(n11291) );
  AOI211_X1 U14060 ( .C1(P3_ADDR_REG_1__SCAN_IN), .C2(n16012), .A(n11292), .B(
        n11291), .ZN(n11293) );
  OAI21_X1 U14061 ( .B1(n8836), .B2(n13617), .A(n11293), .ZN(P3_U3183) );
  OAI21_X1 U14062 ( .B1(n11296), .B2(n11295), .A(n11294), .ZN(n11310) );
  AOI21_X1 U14063 ( .B1(n11299), .B2(n11298), .A(n11297), .ZN(n11306) );
  INV_X1 U14064 ( .A(n11300), .ZN(n11302) );
  NOR3_X1 U14065 ( .A1(n7401), .A2(n11302), .A3(n11301), .ZN(n11304) );
  INV_X1 U14066 ( .A(n11303), .ZN(n11326) );
  OAI21_X1 U14067 ( .B1(n11304), .B2(n11326), .A(n13537), .ZN(n11305) );
  OAI21_X1 U14068 ( .B1(n16014), .B2(n11306), .A(n11305), .ZN(n11309) );
  OAI22_X1 U14069 ( .A1(n16024), .A2(n11307), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n11508), .ZN(n11308) );
  AOI211_X1 U14070 ( .C1(n13631), .C2(n11310), .A(n11309), .B(n11308), .ZN(
        n11311) );
  OAI21_X1 U14071 ( .B1(n11312), .B2(n13617), .A(n11311), .ZN(P3_U3184) );
  NAND2_X1 U14072 ( .A1(n13774), .A2(P3_U3897), .ZN(n11313) );
  OAI21_X1 U14073 ( .B1(P3_U3897), .B2(n11314), .A(n11313), .ZN(P3_U3508) );
  OAI21_X1 U14074 ( .B1(P3_REG2_REG_3__SCAN_IN), .B2(n11315), .A(n11265), .ZN(
        n11323) );
  AOI22_X1 U14075 ( .A1(n16012), .A2(P3_ADDR_REG_3__SCAN_IN), .B1(
        P3_REG3_REG_3__SCAN_IN), .B2(P3_U3151), .ZN(n11316) );
  INV_X1 U14076 ( .A(n11316), .ZN(n11322) );
  NAND2_X1 U14077 ( .A1(n11318), .A2(n11317), .ZN(n11319) );
  AOI21_X1 U14078 ( .B1(n11320), .B2(n11319), .A(n16015), .ZN(n11321) );
  AOI211_X1 U14079 ( .C1(n13583), .C2(n11323), .A(n11322), .B(n11321), .ZN(
        n11331) );
  NOR3_X1 U14080 ( .A1(n11326), .A2(n7405), .A3(n11325), .ZN(n11329) );
  INV_X1 U14081 ( .A(n11327), .ZN(n11328) );
  OAI21_X1 U14082 ( .B1(n11329), .B2(n11328), .A(n13537), .ZN(n11330) );
  OAI211_X1 U14083 ( .C1(n13617), .C2(n7696), .A(n11331), .B(n11330), .ZN(
        P3_U3185) );
  INV_X1 U14084 ( .A(P3_ADDR_REG_6__SCAN_IN), .ZN(n11336) );
  OR2_X1 U14085 ( .A1(P3_ADDR_REG_6__SCAN_IN), .A2(n11332), .ZN(n11333) );
  NAND2_X1 U14086 ( .A1(n11334), .A2(n11333), .ZN(n11335) );
  NAND2_X1 U14087 ( .A1(n11337), .A2(P3_ADDR_REG_7__SCAN_IN), .ZN(n11338) );
  XNOR2_X1 U14088 ( .A(n11579), .B(P1_ADDR_REG_7__SCAN_IN), .ZN(n11344) );
  INV_X1 U14089 ( .A(n11339), .ZN(n11340) );
  NAND2_X1 U14090 ( .A1(n11340), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n11341) );
  NAND2_X1 U14091 ( .A1(n11343), .A2(n11344), .ZN(n11577) );
  OAI21_X1 U14092 ( .B1(n11344), .B2(n11343), .A(n11577), .ZN(n11345) );
  INV_X1 U14093 ( .A(n11345), .ZN(SUB_1596_U56) );
  INV_X1 U14094 ( .A(n11346), .ZN(n11347) );
  OAI222_X1 U14095 ( .A1(P3_U3151), .A2(n13616), .B1(n13962), .B2(n11348), 
        .C1(n13102), .C2(n11347), .ZN(P3_U3278) );
  INV_X1 U14096 ( .A(n15068), .ZN(n15083) );
  INV_X1 U14097 ( .A(n7137), .ZN(n12043) );
  OAI21_X1 U14098 ( .B1(n11351), .B2(n11350), .A(n11349), .ZN(n15115) );
  OR2_X1 U14099 ( .A1(n10123), .A2(n15516), .ZN(n12042) );
  INV_X1 U14100 ( .A(n12042), .ZN(n15828) );
  AOI22_X1 U14101 ( .A1(n15115), .A2(n15072), .B1(n15080), .B2(n15828), .ZN(
        n11354) );
  NAND2_X1 U14102 ( .A1(n12910), .A2(n11352), .ZN(n13092) );
  NAND2_X1 U14103 ( .A1(n13092), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n11353) );
  OAI211_X1 U14104 ( .C1(n15083), .C2(n12043), .A(n11354), .B(n11353), .ZN(
        P1_U3232) );
  OAI21_X1 U14105 ( .B1(n14733), .B2(n14106), .A(n7985), .ZN(n11355) );
  AND2_X1 U14106 ( .A1(n8040), .A2(n14086), .ZN(n11907) );
  AOI22_X1 U14107 ( .A1(n14065), .A2(n11355), .B1(n14097), .B2(n11907), .ZN(
        n11358) );
  OR2_X1 U14108 ( .A1(n11356), .A2(P2_U3088), .ZN(n11511) );
  NAND2_X1 U14109 ( .A1(n11511), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n11357) );
  OAI211_X1 U14110 ( .C1(n14073), .C2(n14110), .A(n11358), .B(n11357), .ZN(
        P2_U3204) );
  XNOR2_X1 U14111 ( .A(n11557), .B(P1_REG1_REG_11__SCAN_IN), .ZN(n11366) );
  NOR2_X1 U14112 ( .A1(n11370), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n11359) );
  INV_X1 U14113 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n11362) );
  XNOR2_X1 U14114 ( .A(n15178), .B(n11362), .ZN(n15174) );
  NAND2_X1 U14115 ( .A1(n15178), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n11363) );
  NAND2_X1 U14116 ( .A1(n15173), .A2(n11363), .ZN(n11365) );
  INV_X1 U14117 ( .A(n11559), .ZN(n11364) );
  AOI21_X1 U14118 ( .B1(n11366), .B2(n11365), .A(n11364), .ZN(n11378) );
  INV_X1 U14119 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n11368) );
  NAND2_X1 U14120 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_U3086), .ZN(n11367)
         );
  OAI21_X1 U14121 ( .B1(n15252), .B2(n11368), .A(n11367), .ZN(n11369) );
  AOI21_X1 U14122 ( .B1(n15223), .B2(n11557), .A(n11369), .ZN(n11377) );
  NAND2_X1 U14123 ( .A1(n11370), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n11371) );
  NAND2_X1 U14124 ( .A1(n11372), .A2(n11371), .ZN(n15181) );
  MUX2_X1 U14125 ( .A(P1_REG2_REG_10__SCAN_IN), .B(n12366), .S(n15178), .Z(
        n15180) );
  NAND2_X1 U14126 ( .A1(n15181), .A2(n15180), .ZN(n15179) );
  NAND2_X1 U14127 ( .A1(n15178), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n11373) );
  NAND2_X1 U14128 ( .A1(n15179), .A2(n11373), .ZN(n11375) );
  INV_X1 U14129 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n12727) );
  XNOR2_X1 U14130 ( .A(n11557), .B(n12727), .ZN(n11374) );
  NAND2_X1 U14131 ( .A1(n11375), .A2(n11374), .ZN(n11551) );
  OAI211_X1 U14132 ( .C1(n11375), .C2(n11374), .A(n11551), .B(n15244), .ZN(
        n11376) );
  OAI211_X1 U14133 ( .C1(n11378), .C2(n15248), .A(n11377), .B(n11376), .ZN(
        P1_U3254) );
  INV_X1 U14134 ( .A(n11379), .ZN(n11382) );
  INV_X1 U14135 ( .A(n11927), .ZN(n11380) );
  OAI222_X1 U14136 ( .A1(n14914), .A2(n11381), .B1(n14903), .B2(n11382), .C1(
        n11380), .C2(P2_U3088), .ZN(P2_U3314) );
  INV_X1 U14137 ( .A(n12164), .ZN(n11902) );
  OAI222_X1 U14138 ( .A1(n15700), .A2(n11383), .B1(n15703), .B2(n11382), .C1(
        P1_U3086), .C2(n11902), .ZN(P1_U3342) );
  INV_X1 U14139 ( .A(n11384), .ZN(n11385) );
  NOR2_X1 U14140 ( .A1(n11386), .A2(n11385), .ZN(n11389) );
  INV_X1 U14141 ( .A(n11387), .ZN(n11542) );
  AOI21_X1 U14142 ( .B1(n11389), .B2(n11388), .A(n11542), .ZN(n11402) );
  NAND3_X1 U14143 ( .A1(n11243), .A2(n11392), .A3(n11391), .ZN(n11393) );
  AOI21_X1 U14144 ( .B1(n6988), .B2(n11393), .A(n16014), .ZN(n11394) );
  AOI21_X1 U14145 ( .B1(n16021), .B2(n7234), .A(n11394), .ZN(n11401) );
  AND2_X1 U14146 ( .A1(P3_U3151), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n12288) );
  NAND3_X1 U14147 ( .A1(n11397), .A2(n11396), .A3(n11395), .ZN(n11398) );
  AOI21_X1 U14148 ( .B1(n6732), .B2(n11398), .A(n16015), .ZN(n11399) );
  AOI211_X1 U14149 ( .C1(n16012), .C2(P3_ADDR_REG_6__SCAN_IN), .A(n12288), .B(
        n11399), .ZN(n11400) );
  OAI211_X1 U14150 ( .C1(n11402), .C2(n16013), .A(n11401), .B(n11400), .ZN(
        P3_U3188) );
  INV_X1 U14151 ( .A(n11411), .ZN(n11407) );
  AND2_X1 U14152 ( .A1(n11404), .A2(n11403), .ZN(n11406) );
  OR2_X1 U14153 ( .A1(n11419), .A2(n11412), .ZN(n11405) );
  OAI211_X1 U14154 ( .C1(n11424), .C2(n11407), .A(n11406), .B(n11405), .ZN(
        n11408) );
  NAND2_X1 U14155 ( .A1(n11408), .A2(P3_STATE_REG_SCAN_IN), .ZN(n11410) );
  OR2_X1 U14156 ( .A1(n13486), .A2(n11419), .ZN(n11409) );
  NAND2_X1 U14157 ( .A1(n11410), .A2(n11409), .ZN(n11610) );
  NOR2_X1 U14158 ( .A1(n11610), .A2(n13959), .ZN(n11509) );
  NAND3_X1 U14159 ( .A1(n11424), .A2(n16055), .A3(n11411), .ZN(n11415) );
  INV_X1 U14160 ( .A(n11412), .ZN(n11413) );
  NAND2_X1 U14161 ( .A1(n11419), .A2(n11413), .ZN(n11414) );
  NAND2_X1 U14162 ( .A1(n11415), .A2(n11414), .ZN(n11417) );
  NAND2_X1 U14163 ( .A1(n16048), .A2(n11845), .ZN(n13335) );
  INV_X1 U14164 ( .A(n13335), .ZN(n11418) );
  NOR2_X1 U14165 ( .A1(n13339), .A2(n11418), .ZN(n13314) );
  INV_X1 U14166 ( .A(n13314), .ZN(n11427) );
  INV_X1 U14167 ( .A(n13486), .ZN(n11420) );
  INV_X1 U14168 ( .A(n11441), .ZN(n11421) );
  NOR2_X1 U14169 ( .A1(n11422), .A2(n16055), .ZN(n11423) );
  NAND2_X1 U14170 ( .A1(n11424), .A2(n11423), .ZN(n11425) );
  OAI22_X1 U14171 ( .A1(n11432), .A2(n13271), .B1(n13276), .B2(n11845), .ZN(
        n11426) );
  AOI21_X1 U14172 ( .B1(n13243), .B2(n11427), .A(n11426), .ZN(n11428) );
  OAI21_X1 U14173 ( .B1(n11509), .B2(n11429), .A(n11428), .ZN(P3_U3172) );
  NOR3_X1 U14174 ( .A1(n11432), .A2(n16056), .A3(n11436), .ZN(n11433) );
  INV_X1 U14175 ( .A(n11434), .ZN(n11435) );
  OAI211_X1 U14176 ( .C1(n11435), .C2(n12957), .A(n11438), .B(n16043), .ZN(
        n11501) );
  INV_X1 U14177 ( .A(n13339), .ZN(n16053) );
  NAND3_X1 U14178 ( .A1(n16053), .A2(n16052), .A3(n11436), .ZN(n11437) );
  OAI211_X1 U14179 ( .C1(n11438), .C2(n16043), .A(n11501), .B(n11437), .ZN(
        n11439) );
  NAND2_X1 U14180 ( .A1(n11439), .A2(n13243), .ZN(n11444) );
  OAI22_X1 U14181 ( .A1(n7260), .A2(n13271), .B1(n13276), .B2(n16056), .ZN(
        n11442) );
  AOI21_X1 U14182 ( .B1(n13269), .B2(n16048), .A(n11442), .ZN(n11443) );
  OAI211_X1 U14183 ( .C1(n11509), .C2(n11445), .A(n11444), .B(n11443), .ZN(
        P3_U3162) );
  NOR2_X1 U14184 ( .A1(n10430), .A2(n11447), .ZN(n11451) );
  INV_X1 U14185 ( .A(n11566), .ZN(n11449) );
  NAND2_X1 U14186 ( .A1(n11449), .A2(n11448), .ZN(n11450) );
  NOR2_X1 U14187 ( .A1(n11451), .A2(n11450), .ZN(n11567) );
  AOI21_X1 U14188 ( .B1(n11451), .B2(n11450), .A(n11567), .ZN(n11456) );
  OAI22_X1 U14189 ( .A1(n11453), .A2(n14095), .B1(n11452), .B2(n14096), .ZN(
        n11630) );
  AOI22_X1 U14190 ( .A1(n14097), .A2(n11630), .B1(n14101), .B2(n14120), .ZN(
        n11455) );
  NAND2_X1 U14191 ( .A1(n11511), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n11454) );
  OAI211_X1 U14192 ( .C1(n11456), .C2(n14103), .A(n11455), .B(n11454), .ZN(
        P2_U3209) );
  INV_X1 U14193 ( .A(n13641), .ZN(n11460) );
  INV_X1 U14194 ( .A(n11457), .ZN(n11458) );
  OAI222_X1 U14195 ( .A1(P3_U3151), .A2(n11460), .B1(n13970), .B2(n11459), 
        .C1(n13102), .C2(n11458), .ZN(P3_U3277) );
  OAI222_X1 U14196 ( .A1(n13102), .A2(n11462), .B1(n13962), .B2(n11461), .C1(
        P3_U3151), .C2(n13306), .ZN(P3_U3276) );
  NOR2_X1 U14197 ( .A1(n11467), .A2(n11463), .ZN(n11464) );
  NOR2_X1 U14198 ( .A1(n11465), .A2(n11464), .ZN(n11469) );
  OAI21_X1 U14199 ( .B1(n11467), .B2(P1_D_REG_0__SCAN_IN), .A(n11466), .ZN(
        n11468) );
  INV_X1 U14200 ( .A(n11827), .ZN(n11470) );
  NOR2_X1 U14201 ( .A1(n11472), .A2(n11471), .ZN(n11473) );
  INV_X1 U14202 ( .A(n11831), .ZN(n11475) );
  NAND2_X1 U14203 ( .A1(n11475), .A2(n9780), .ZN(n15436) );
  NAND2_X1 U14204 ( .A1(n7133), .A2(n15250), .ZN(n15620) );
  XNOR2_X1 U14205 ( .A(n11478), .B(n11794), .ZN(n11841) );
  AND2_X1 U14206 ( .A1(n7137), .A2(n11483), .ZN(n11477) );
  OR2_X1 U14207 ( .A1(n11477), .A2(n11853), .ZN(n11837) );
  XNOR2_X1 U14208 ( .A(n11837), .B(n10123), .ZN(n11479) );
  MUX2_X1 U14209 ( .A(n11479), .B(n11478), .S(n7136), .Z(n11481) );
  AOI22_X1 U14210 ( .A1(n7136), .A2(n15521), .B1(n15500), .B2(n10144), .ZN(
        n11480) );
  OAI21_X1 U14211 ( .B1(n11481), .B2(n15826), .A(n11480), .ZN(n11482) );
  INV_X1 U14212 ( .A(n11482), .ZN(n11836) );
  INV_X1 U14213 ( .A(n11837), .ZN(n11484) );
  AOI22_X1 U14214 ( .A1(n11484), .A2(n7132), .B1(n15870), .B2(n11483), .ZN(
        n11485) );
  OAI211_X1 U14215 ( .C1(n15874), .C2(n11841), .A(n11836), .B(n11485), .ZN(
        n11496) );
  NAND2_X1 U14216 ( .A1(n11496), .A2(n15877), .ZN(n11486) );
  OAI21_X1 U14217 ( .B1(n15877), .B2(n9485), .A(n11486), .ZN(P1_U3462) );
  AOI21_X1 U14218 ( .B1(P1_REG3_REG_1__SCAN_IN), .B2(n13092), .A(n11487), .ZN(
        n11493) );
  OAI21_X1 U14219 ( .B1(n11488), .B2(n11490), .A(n11489), .ZN(n11491) );
  NAND2_X1 U14220 ( .A1(n11491), .A2(n15072), .ZN(n11492) );
  OAI211_X1 U14221 ( .C1(n11795), .C2(n15083), .A(n11493), .B(n11492), .ZN(
        P1_U3222) );
  NAND2_X1 U14222 ( .A1(n11496), .A2(n15886), .ZN(n11497) );
  OAI21_X1 U14223 ( .B1(n15886), .B2(n11498), .A(n11497), .ZN(P1_U3529) );
  XNOR2_X1 U14224 ( .A(n11436), .B(n16036), .ZN(n11603) );
  XNOR2_X1 U14225 ( .A(n11603), .B(n7260), .ZN(n11503) );
  INV_X1 U14226 ( .A(n11499), .ZN(n11500) );
  NAND2_X1 U14227 ( .A1(n11501), .A2(n11500), .ZN(n11502) );
  NAND2_X1 U14228 ( .A1(n11502), .A2(n11503), .ZN(n11606) );
  OAI21_X1 U14229 ( .B1(n11503), .B2(n11502), .A(n11606), .ZN(n11504) );
  NAND2_X1 U14230 ( .A1(n11504), .A2(n13243), .ZN(n11507) );
  INV_X1 U14231 ( .A(n16031), .ZN(n11787) );
  OAI22_X1 U14232 ( .A1(n11787), .A2(n13271), .B1(n13276), .B2(n16036), .ZN(
        n11505) );
  AOI21_X1 U14233 ( .B1(n13269), .B2(n7149), .A(n11505), .ZN(n11506) );
  OAI211_X1 U14234 ( .C1(n11509), .C2(n11508), .A(n11507), .B(n11506), .ZN(
        P3_U3177) );
  AOI22_X1 U14235 ( .A1(n14376), .A2(n14421), .B1(n14420), .B2(n14086), .ZN(
        n11773) );
  OAI22_X1 U14236 ( .A1(n14073), .A2(n8039), .B1(n11773), .B2(n14090), .ZN(
        n11510) );
  AOI21_X1 U14237 ( .B1(P2_REG3_REG_1__SCAN_IN), .B2(n11511), .A(n11510), .ZN(
        n11516) );
  OAI21_X1 U14238 ( .B1(n11513), .B2(n11512), .A(n11446), .ZN(n11514) );
  NAND2_X1 U14239 ( .A1(n14065), .A2(n11514), .ZN(n11515) );
  NAND2_X1 U14240 ( .A1(n11516), .A2(n11515), .ZN(P2_U3194) );
  XNOR2_X1 U14241 ( .A(n11523), .B(P2_REG1_REG_12__SCAN_IN), .ZN(n11521) );
  NAND2_X1 U14242 ( .A1(n11522), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n11517) );
  NAND2_X1 U14243 ( .A1(n11518), .A2(n11517), .ZN(n11520) );
  INV_X1 U14244 ( .A(n11721), .ZN(n11519) );
  AOI21_X1 U14245 ( .B1(n11521), .B2(n11520), .A(n11519), .ZN(n11533) );
  NAND2_X1 U14246 ( .A1(P2_U3088), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n12893)
         );
  OAI21_X1 U14247 ( .B1(n15919), .B2(n11726), .A(n12893), .ZN(n11531) );
  OR2_X1 U14248 ( .A1(n11522), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n11526) );
  MUX2_X1 U14249 ( .A(P2_REG2_REG_12__SCAN_IN), .B(n11725), .S(n11523), .Z(
        n11525) );
  NAND2_X1 U14250 ( .A1(n11524), .A2(n11525), .ZN(n11728) );
  INV_X1 U14251 ( .A(n11525), .ZN(n11527) );
  NAND3_X1 U14252 ( .A1(n11528), .A2(n11527), .A3(n11526), .ZN(n11529) );
  AOI21_X1 U14253 ( .B1(n11728), .B2(n11529), .A(n14504), .ZN(n11530) );
  AOI211_X1 U14254 ( .C1(n15899), .C2(P2_ADDR_REG_12__SCAN_IN), .A(n11531), 
        .B(n11530), .ZN(n11532) );
  OAI21_X1 U14255 ( .B1(n11533), .B2(n15904), .A(n11532), .ZN(P2_U3226) );
  AOI21_X1 U14256 ( .B1(n12132), .B2(n11534), .A(n6733), .ZN(n11547) );
  OAI21_X1 U14257 ( .B1(P3_REG1_REG_7__SCAN_IN), .B2(n11535), .A(n11698), .ZN(
        n11538) );
  AND2_X1 U14258 ( .A1(P3_U3151), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n12312) );
  AOI21_X1 U14259 ( .B1(n16012), .B2(P3_ADDR_REG_7__SCAN_IN), .A(n12312), .ZN(
        n11536) );
  OAI21_X1 U14260 ( .B1(n13617), .B2(n7718), .A(n11536), .ZN(n11537) );
  AOI21_X1 U14261 ( .B1(n11538), .B2(n13631), .A(n11537), .ZN(n11546) );
  INV_X1 U14262 ( .A(n11539), .ZN(n11541) );
  NOR3_X1 U14263 ( .A1(n11542), .A2(n11541), .A3(n11540), .ZN(n11544) );
  INV_X1 U14264 ( .A(n11694), .ZN(n11543) );
  OAI21_X1 U14265 ( .B1(n11544), .B2(n11543), .A(n13537), .ZN(n11545) );
  OAI211_X1 U14266 ( .C1(n11547), .C2(n16014), .A(n11546), .B(n11545), .ZN(
        P3_U3189) );
  INV_X1 U14267 ( .A(n11548), .ZN(n11586) );
  AOI22_X1 U14268 ( .A1(n15205), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(n15691), .ZN(n11549) );
  OAI21_X1 U14269 ( .B1(n11586), .B2(n15703), .A(n11549), .ZN(P1_U3339) );
  MUX2_X1 U14270 ( .A(n9677), .B(P1_REG2_REG_12__SCAN_IN), .S(n11895), .Z(
        n11554) );
  NAND2_X1 U14271 ( .A1(n11557), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n11550) );
  NAND2_X1 U14272 ( .A1(n11551), .A2(n11550), .ZN(n11553) );
  INV_X1 U14273 ( .A(n11897), .ZN(n11552) );
  AOI21_X1 U14274 ( .B1(n11554), .B2(n11553), .A(n11552), .ZN(n11565) );
  INV_X1 U14275 ( .A(n15244), .ZN(n15242) );
  AND2_X1 U14276 ( .A1(P1_U3086), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n14975) );
  NOR2_X1 U14277 ( .A1(n15252), .A2(n12846), .ZN(n11555) );
  AOI211_X1 U14278 ( .C1(n15223), .C2(n11895), .A(n14975), .B(n11555), .ZN(
        n11564) );
  XNOR2_X1 U14279 ( .A(n11895), .B(n11556), .ZN(n11561) );
  OR2_X1 U14280 ( .A1(n11557), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n11558) );
  OAI21_X1 U14281 ( .B1(n11561), .B2(n11560), .A(n11891), .ZN(n11562) );
  INV_X1 U14282 ( .A(n15248), .ZN(n15218) );
  NAND2_X1 U14283 ( .A1(n11562), .A2(n15218), .ZN(n11563) );
  OAI211_X1 U14284 ( .C1(n11565), .C2(n15242), .A(n11564), .B(n11563), .ZN(
        P1_U3255) );
  NOR2_X1 U14285 ( .A1(n11567), .A2(n11566), .ZN(n11569) );
  XNOR2_X1 U14286 ( .A(n11569), .B(n11568), .ZN(n11574) );
  OAI22_X1 U14287 ( .A1(n11570), .A2(n14095), .B1(n11743), .B2(n14096), .ZN(
        n11674) );
  AOI22_X1 U14288 ( .A1(n14097), .A2(n11674), .B1(P2_REG3_REG_3__SCAN_IN), 
        .B2(P2_U3088), .ZN(n11571) );
  OAI21_X1 U14289 ( .B1(n11713), .B2(n14073), .A(n11571), .ZN(n11572) );
  AOI21_X1 U14290 ( .B1(n14088), .B2(n8057), .A(n11572), .ZN(n11573) );
  OAI21_X1 U14291 ( .B1(n11574), .B2(n14103), .A(n11573), .ZN(P2_U3190) );
  NAND2_X1 U14292 ( .A1(n11575), .A2(P2_ADDR_REG_7__SCAN_IN), .ZN(n11576) );
  INV_X1 U14293 ( .A(P3_ADDR_REG_8__SCAN_IN), .ZN(n11580) );
  NAND2_X1 U14294 ( .A1(n11580), .A2(P1_ADDR_REG_8__SCAN_IN), .ZN(n11946) );
  NAND2_X1 U14295 ( .A1(n11114), .A2(P3_ADDR_REG_8__SCAN_IN), .ZN(n11581) );
  AND2_X1 U14296 ( .A1(n11946), .A2(n11581), .ZN(n11582) );
  NAND2_X1 U14297 ( .A1(n11583), .A2(n11582), .ZN(n11947) );
  OR2_X1 U14298 ( .A1(n11583), .A2(n11582), .ZN(n11584) );
  NAND2_X1 U14299 ( .A1(n11947), .A2(n11584), .ZN(n11942) );
  INV_X1 U14300 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n14478) );
  XNOR2_X1 U14301 ( .A(n11941), .B(n14478), .ZN(SUB_1596_U55) );
  INV_X1 U14302 ( .A(n15935), .ZN(n11585) );
  OAI222_X1 U14303 ( .A1(n14914), .A2(n11587), .B1(n14903), .B2(n11586), .C1(
        n11585), .C2(P2_U3088), .ZN(P2_U3311) );
  INV_X1 U14304 ( .A(n11588), .ZN(n11591) );
  INV_X1 U14305 ( .A(n15191), .ZN(n11589) );
  OAI222_X1 U14306 ( .A1(n15700), .A2(n11590), .B1(n15703), .B2(n11591), .C1(
        P1_U3086), .C2(n11589), .ZN(P1_U3341) );
  INV_X1 U14307 ( .A(n11993), .ZN(n11926) );
  OAI222_X1 U14308 ( .A1(n14914), .A2(n11592), .B1(n14903), .B2(n11591), .C1(
        n11926), .C2(P2_U3088), .ZN(P2_U3313) );
  INV_X1 U14309 ( .A(n11593), .ZN(n11665) );
  AOI22_X1 U14310 ( .A1(n15224), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n15691), .ZN(n11594) );
  OAI21_X1 U14311 ( .B1(n11665), .B2(n15703), .A(n11594), .ZN(P1_U3338) );
  NAND2_X1 U14312 ( .A1(n11595), .A2(n16055), .ZN(n11596) );
  OAI22_X1 U14313 ( .A1(n13314), .A2(n11596), .B1(n11432), .B2(n13817), .ZN(
        n11843) );
  INV_X1 U14314 ( .A(P3_REG0_REG_0__SCAN_IN), .ZN(n11597) );
  NOR2_X1 U14315 ( .A1(n16094), .A2(n11597), .ZN(n11598) );
  AOI21_X1 U14316 ( .B1(n16094), .B2(n11843), .A(n11598), .ZN(n11599) );
  OAI21_X1 U14317 ( .B1(n11845), .B2(n13918), .A(n11599), .ZN(P3_U3390) );
  INV_X2 U14318 ( .A(n12707), .ZN(n16061) );
  AOI22_X1 U14319 ( .A1(n11843), .A2(n9401), .B1(P3_REG3_REG_0__SCAN_IN), .B2(
        n16061), .ZN(n11602) );
  NAND2_X1 U14320 ( .A1(n13814), .A2(n11600), .ZN(n11601) );
  OAI211_X1 U14321 ( .C1(n8917), .C2(n9401), .A(n11602), .B(n11601), .ZN(
        P3_U3233) );
  XNOR2_X1 U14322 ( .A(n11650), .B(n16031), .ZN(n11607) );
  INV_X1 U14323 ( .A(n11603), .ZN(n11604) );
  NAND2_X1 U14324 ( .A1(n11604), .A2(n7260), .ZN(n11608) );
  NAND2_X1 U14325 ( .A1(n11653), .A2(n13243), .ZN(n11615) );
  AOI21_X1 U14326 ( .B1(n11606), .B2(n11608), .A(n11607), .ZN(n11614) );
  INV_X1 U14327 ( .A(n13509), .ZN(n11654) );
  OAI22_X1 U14328 ( .A1(n11654), .A2(n13271), .B1(n13276), .B2(n11647), .ZN(
        n11612) );
  INV_X1 U14329 ( .A(n13490), .ZN(n11609) );
  MUX2_X1 U14330 ( .A(n13273), .B(P3_U3151), .S(P3_REG3_REG_3__SCAN_IN), .Z(
        n11611) );
  AOI211_X1 U14331 ( .C1(n13269), .C2(n16047), .A(n11612), .B(n11611), .ZN(
        n11613) );
  OAI21_X1 U14332 ( .B1(n11615), .B2(n11614), .A(n11613), .ZN(P3_U3158) );
  INV_X1 U14333 ( .A(n11616), .ZN(n11617) );
  AOI21_X1 U14334 ( .B1(n11619), .B2(n11618), .A(n11617), .ZN(n11623) );
  AOI22_X1 U14335 ( .A1(n14086), .A2(n14417), .B1(n14419), .B2(n14376), .ZN(
        n11818) );
  NAND2_X1 U14336 ( .A1(n14101), .A2(n14136), .ZN(n11620) );
  NAND2_X1 U14337 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_U3088), .ZN(n14435) );
  OAI211_X1 U14338 ( .C1(n11818), .C2(n14090), .A(n11620), .B(n14435), .ZN(
        n11621) );
  AOI21_X1 U14339 ( .B1(n12534), .B2(n14088), .A(n11621), .ZN(n11622) );
  OAI21_X1 U14340 ( .B1(n11623), .B2(n14103), .A(n11622), .ZN(P2_U3202) );
  OAI21_X1 U14341 ( .B1(n11626), .B2(n11625), .A(n11624), .ZN(n12350) );
  NAND2_X1 U14342 ( .A1(n11769), .A2(n14120), .ZN(n11627) );
  NAND2_X1 U14343 ( .A1(n11627), .A2(n14818), .ZN(n11628) );
  NOR2_X1 U14344 ( .A1(n11676), .A2(n11628), .ZN(n12349) );
  XNOR2_X1 U14345 ( .A(n11629), .B(n14332), .ZN(n11631) );
  AOI21_X1 U14346 ( .B1(n11631), .B2(n14675), .A(n11630), .ZN(n12353) );
  INV_X1 U14347 ( .A(n12353), .ZN(n11632) );
  AOI211_X1 U14348 ( .C1(n15993), .C2(n12350), .A(n12349), .B(n11632), .ZN(
        n11718) );
  INV_X1 U14349 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n11635) );
  OAI22_X1 U14350 ( .A1(n14892), .A2(n7166), .B1(n16004), .B2(n11635), .ZN(
        n11636) );
  INV_X1 U14351 ( .A(n11636), .ZN(n11637) );
  OAI21_X1 U14352 ( .B1(n11718), .B2(n16002), .A(n11637), .ZN(P2_U3436) );
  INV_X1 U14353 ( .A(n11639), .ZN(n13316) );
  AOI21_X1 U14354 ( .B1(n11638), .B2(n13316), .A(n16034), .ZN(n11640) );
  OR2_X1 U14355 ( .A1(n11638), .A2(n13316), .ZN(n11785) );
  NAND2_X1 U14356 ( .A1(n11640), .A2(n11785), .ZN(n11642) );
  AOI22_X1 U14357 ( .A1(n16046), .A2(n13509), .B1(n16047), .B2(n16049), .ZN(
        n11641) );
  AND2_X1 U14358 ( .A1(n11642), .A2(n11641), .ZN(n11683) );
  NAND2_X1 U14359 ( .A1(n11643), .A2(n13316), .ZN(n11781) );
  OR2_X1 U14360 ( .A1(n11643), .A2(n13316), .ZN(n11644) );
  NAND2_X1 U14361 ( .A1(n11781), .A2(n11644), .ZN(n11681) );
  NAND2_X1 U14362 ( .A1(n11681), .A2(n16070), .ZN(n11645) );
  NAND2_X1 U14363 ( .A1(n11683), .A2(n11645), .ZN(n12121) );
  INV_X1 U14364 ( .A(P3_REG0_REG_3__SCAN_IN), .ZN(n11646) );
  OAI22_X1 U14365 ( .A1(n11647), .A2(n13918), .B1(n16094), .B2(n11646), .ZN(
        n11648) );
  AOI21_X1 U14366 ( .B1(n12121), .B2(n16094), .A(n11648), .ZN(n11649) );
  INV_X1 U14367 ( .A(n11649), .ZN(P3_U3399) );
  INV_X1 U14368 ( .A(n11650), .ZN(n11651) );
  XNOR2_X1 U14369 ( .A(n11436), .B(n11886), .ZN(n11655) );
  NAND2_X1 U14370 ( .A1(n11655), .A2(n11654), .ZN(n11912) );
  OAI21_X1 U14371 ( .B1(n11655), .B2(n11654), .A(n11912), .ZN(n11656) );
  AOI21_X1 U14372 ( .B1(n11657), .B2(n11656), .A(n11913), .ZN(n11663) );
  INV_X1 U14373 ( .A(n11658), .ZN(n11885) );
  INV_X1 U14374 ( .A(n13271), .ZN(n13247) );
  AOI22_X1 U14375 ( .A1(n13247), .A2(n13508), .B1(n13269), .B2(n16031), .ZN(
        n11660) );
  OAI211_X1 U14376 ( .C1(n13276), .C2(n11974), .A(n11660), .B(n11659), .ZN(
        n11661) );
  AOI21_X1 U14377 ( .B1(n11885), .B2(n13273), .A(n11661), .ZN(n11662) );
  OAI21_X1 U14378 ( .B1(n11663), .B2(n13264), .A(n11662), .ZN(P3_U3170) );
  INV_X1 U14379 ( .A(n12803), .ZN(n12685) );
  OAI222_X1 U14380 ( .A1(P2_U3088), .A2(n12685), .B1(n14903), .B2(n11665), 
        .C1(n11664), .C2(n14914), .ZN(P2_U3310) );
  INV_X1 U14381 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n11667) );
  INV_X1 U14382 ( .A(n11666), .ZN(n11668) );
  OAI222_X1 U14383 ( .A1(n14914), .A2(n11667), .B1(n14903), .B2(n11668), .C1(
        P2_U3088), .C2(n11996), .ZN(P2_U3312) );
  INV_X1 U14384 ( .A(n12644), .ZN(n12633) );
  OAI222_X1 U14385 ( .A1(n13134), .A2(n11669), .B1(n15703), .B2(n11668), .C1(
        n12633), .C2(P1_U3086), .ZN(P1_U3340) );
  OAI21_X1 U14386 ( .B1(n11672), .B2(n11671), .A(n11670), .ZN(n12546) );
  INV_X1 U14387 ( .A(n12546), .ZN(n11677) );
  XNOR2_X1 U14388 ( .A(n11673), .B(n14333), .ZN(n11675) );
  AOI21_X1 U14389 ( .B1(n11675), .B2(n14675), .A(n11674), .ZN(n12548) );
  OAI211_X1 U14390 ( .C1(n11676), .C2(n11713), .A(n14818), .B(n11816), .ZN(
        n12544) );
  OAI211_X1 U14391 ( .C1(n11677), .C2(n16000), .A(n12548), .B(n12544), .ZN(
        n11715) );
  INV_X1 U14392 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n11678) );
  OAI22_X1 U14393 ( .A1(n14892), .A2(n11713), .B1(n16004), .B2(n11678), .ZN(
        n11679) );
  AOI21_X1 U14394 ( .B1(n11715), .B2(n16004), .A(n11679), .ZN(n11680) );
  INV_X1 U14395 ( .A(n11680), .ZN(P2_U3439) );
  INV_X1 U14396 ( .A(n11681), .ZN(n11687) );
  MUX2_X1 U14397 ( .A(n11683), .B(n11682), .S(n16066), .Z(n11686) );
  AOI22_X1 U14398 ( .A1(n13814), .A2(n12123), .B1(n16061), .B2(n11684), .ZN(
        n11685) );
  OAI211_X1 U14399 ( .C1(n13824), .C2(n11687), .A(n11686), .B(n11685), .ZN(
        P3_U3230) );
  OR3_X1 U14400 ( .A1(n11689), .A2(n6733), .A3(n11688), .ZN(n11690) );
  AOI21_X1 U14401 ( .B1(n11691), .B2(n11690), .A(n16014), .ZN(n11706) );
  NAND3_X1 U14402 ( .A1(n11694), .A2(n11693), .A3(n7420), .ZN(n11695) );
  AOI21_X1 U14403 ( .B1(n12056), .B2(n11695), .A(n16013), .ZN(n11705) );
  AND3_X1 U14404 ( .A1(n11698), .A2(n11697), .A3(n11696), .ZN(n11699) );
  OAI21_X1 U14405 ( .B1(n11700), .B2(n11699), .A(n13631), .ZN(n11702) );
  AND2_X1 U14406 ( .A1(P3_U3151), .A2(P3_REG3_REG_8__SCAN_IN), .ZN(n12479) );
  AOI21_X1 U14407 ( .B1(n16012), .B2(P3_ADDR_REG_8__SCAN_IN), .A(n12479), .ZN(
        n11701) );
  OAI211_X1 U14408 ( .C1(n13617), .C2(n11703), .A(n11702), .B(n11701), .ZN(
        n11704) );
  OR3_X1 U14409 ( .A1(n11706), .A2(n11705), .A3(n11704), .ZN(P3_U3190) );
  NOR2_X1 U14410 ( .A1(n13970), .A2(SI_22_), .ZN(n11707) );
  AOI21_X1 U14411 ( .B1(n11708), .B2(P3_STATE_REG_SCAN_IN), .A(n11707), .ZN(
        n11709) );
  OAI21_X1 U14412 ( .B1(n11710), .B2(n13102), .A(n11709), .ZN(n11711) );
  INV_X1 U14413 ( .A(n11711), .ZN(P3_U3273) );
  OAI22_X1 U14414 ( .A1(n14840), .A2(n11713), .B1(n16011), .B2(n11712), .ZN(
        n11714) );
  AOI21_X1 U14415 ( .B1(n11715), .B2(n16011), .A(n11714), .ZN(n11716) );
  INV_X1 U14416 ( .A(n11716), .ZN(P2_U3502) );
  INV_X1 U14417 ( .A(n14840), .ZN(n12784) );
  AOI22_X1 U14418 ( .A1(n12784), .A2(n14120), .B1(n16008), .B2(
        P2_REG1_REG_2__SCAN_IN), .ZN(n11717) );
  OAI21_X1 U14419 ( .B1(n11718), .B2(n16008), .A(n11717), .ZN(P2_U3501) );
  XNOR2_X1 U14420 ( .A(n11927), .B(P2_REG1_REG_13__SCAN_IN), .ZN(n11724) );
  INV_X1 U14421 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n11719) );
  NAND2_X1 U14422 ( .A1(n11726), .A2(n11719), .ZN(n11720) );
  NAND2_X1 U14423 ( .A1(n11721), .A2(n11720), .ZN(n11723) );
  INV_X1 U14424 ( .A(n11929), .ZN(n11722) );
  AOI211_X1 U14425 ( .C1(n11724), .C2(n11723), .A(n15904), .B(n11722), .ZN(
        n11737) );
  NAND2_X1 U14426 ( .A1(n11726), .A2(n11725), .ZN(n11727) );
  INV_X1 U14427 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n11729) );
  MUX2_X1 U14428 ( .A(n11729), .B(P2_REG2_REG_13__SCAN_IN), .S(n11927), .Z(
        n11731) );
  INV_X1 U14429 ( .A(n11925), .ZN(n11730) );
  AOI211_X1 U14430 ( .C1(n11732), .C2(n11731), .A(n14504), .B(n11730), .ZN(
        n11736) );
  INV_X1 U14431 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n15711) );
  NOR2_X1 U14432 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n12925), .ZN(n11733) );
  AOI21_X1 U14433 ( .B1(n15936), .B2(n11927), .A(n11733), .ZN(n11734) );
  OAI21_X1 U14434 ( .B1(n15711), .B2(n15944), .A(n11734), .ZN(n11735) );
  OR3_X1 U14435 ( .A1(n11737), .A2(n11736), .A3(n11735), .ZN(P2_U3227) );
  INV_X1 U14436 ( .A(n11738), .ZN(n12226) );
  OAI21_X1 U14437 ( .B1(n11741), .B2(n11740), .A(n11739), .ZN(n11742) );
  NAND2_X1 U14438 ( .A1(n11742), .A2(n14065), .ZN(n11748) );
  OAI22_X1 U14439 ( .A1(n11744), .A2(n14096), .B1(n11743), .B2(n14095), .ZN(
        n12222) );
  INV_X1 U14440 ( .A(n12222), .ZN(n11745) );
  NAND2_X1 U14441 ( .A1(P2_REG3_REG_5__SCAN_IN), .A2(P2_U3088), .ZN(n14449) );
  OAI21_X1 U14442 ( .B1(n14090), .B2(n11745), .A(n14449), .ZN(n11746) );
  AOI21_X1 U14443 ( .B1(n15983), .B2(n14101), .A(n11746), .ZN(n11747) );
  OAI211_X1 U14444 ( .C1(n14099), .C2(n12226), .A(n11748), .B(n11747), .ZN(
        P2_U3199) );
  INV_X1 U14445 ( .A(n11749), .ZN(n11752) );
  OAI222_X1 U14446 ( .A1(n13102), .A2(n11752), .B1(n13962), .B2(n11751), .C1(
        P3_U3151), .C2(n11750), .ZN(P3_U3275) );
  INV_X1 U14447 ( .A(n11753), .ZN(n11754) );
  AOI211_X1 U14448 ( .C1(n11756), .C2(n11755), .A(n15070), .B(n11754), .ZN(
        n11760) );
  INV_X1 U14449 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n11966) );
  AOI22_X1 U14450 ( .A1(n15068), .A2(n11965), .B1(n15061), .B2(n11966), .ZN(
        n11758) );
  AOI22_X1 U14451 ( .A1(n15062), .A2(n10144), .B1(P1_REG3_REG_3__SCAN_IN), 
        .B2(P1_U3086), .ZN(n11757) );
  OAI211_X1 U14452 ( .C1(n15793), .C2(n15065), .A(n11758), .B(n11757), .ZN(
        n11759) );
  OR2_X1 U14453 ( .A1(n11760), .A2(n11759), .ZN(P1_U3218) );
  XNOR2_X1 U14454 ( .A(n11762), .B(n11761), .ZN(n11766) );
  AOI22_X1 U14455 ( .A1(n14376), .A2(n14417), .B1(n14415), .B2(n14086), .ZN(
        n12617) );
  NAND2_X1 U14456 ( .A1(n14101), .A2(n14148), .ZN(n11763) );
  NAND2_X1 U14457 ( .A1(P2_U3088), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n15916) );
  OAI211_X1 U14458 ( .C1(n12617), .C2(n14090), .A(n11763), .B(n15916), .ZN(
        n11764) );
  AOI21_X1 U14459 ( .B1(n12611), .B2(n14088), .A(n11764), .ZN(n11765) );
  OAI21_X1 U14460 ( .B1(n11766), .B2(n14103), .A(n11765), .ZN(P2_U3211) );
  OAI21_X1 U14461 ( .B1(n11772), .B2(n11768), .A(n11767), .ZN(n12524) );
  AOI21_X1 U14462 ( .B1(n14108), .B2(n14114), .A(n14717), .ZN(n11770) );
  NAND2_X1 U14463 ( .A1(n11770), .A2(n11769), .ZN(n12521) );
  INV_X1 U14464 ( .A(n12521), .ZN(n11775) );
  XNOR2_X1 U14465 ( .A(n11772), .B(n11771), .ZN(n11774) );
  OAI21_X1 U14466 ( .B1(n11774), .B2(n8640), .A(n11773), .ZN(n12519) );
  AOI211_X1 U14467 ( .C1(n15993), .C2(n12524), .A(n11775), .B(n12519), .ZN(
        n11780) );
  INV_X1 U14468 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n11776) );
  OAI22_X1 U14469 ( .A1(n14892), .A2(n8039), .B1(n16004), .B2(n11776), .ZN(
        n11777) );
  INV_X1 U14470 ( .A(n11777), .ZN(n11778) );
  OAI21_X1 U14471 ( .B1(n11780), .B2(n16002), .A(n11778), .ZN(P2_U3433) );
  AOI22_X1 U14472 ( .A1(n12784), .A2(n14114), .B1(n16008), .B2(
        P2_REG1_REG_1__SCAN_IN), .ZN(n11779) );
  OAI21_X1 U14473 ( .B1(n11780), .B2(n16008), .A(n11779), .ZN(P2_U3500) );
  NAND2_X1 U14474 ( .A1(n11781), .A2(n13354), .ZN(n11782) );
  XNOR2_X1 U14475 ( .A(n11782), .B(n13355), .ZN(n11889) );
  INV_X1 U14476 ( .A(n11783), .ZN(n11784) );
  NAND2_X1 U14477 ( .A1(n11785), .A2(n11784), .ZN(n11786) );
  INV_X1 U14478 ( .A(n13355), .ZN(n13317) );
  XNOR2_X1 U14479 ( .A(n11786), .B(n13317), .ZN(n11789) );
  OAI22_X1 U14480 ( .A1(n11787), .A2(n13815), .B1(n12286), .B2(n13817), .ZN(
        n11788) );
  AOI21_X1 U14481 ( .B1(n11789), .B2(n16044), .A(n11788), .ZN(n11884) );
  OAI21_X1 U14482 ( .B1(n11790), .B2(n11889), .A(n11884), .ZN(n11976) );
  OAI22_X1 U14483 ( .A1(n11974), .A2(n13918), .B1(n16094), .B2(n8963), .ZN(
        n11791) );
  AOI21_X1 U14484 ( .B1(n11976), .B2(n16094), .A(n11791), .ZN(n11792) );
  INV_X1 U14485 ( .A(n11792), .ZN(P3_U3402) );
  NAND2_X1 U14486 ( .A1(n10123), .A2(n11795), .ZN(n11796) );
  NAND2_X1 U14487 ( .A1(n11797), .A2(n11796), .ZN(n11848) );
  NAND2_X1 U14488 ( .A1(n11954), .A2(n11800), .ZN(n12027) );
  INV_X1 U14489 ( .A(n12027), .ZN(n15796) );
  XNOR2_X1 U14490 ( .A(n15796), .B(n11807), .ZN(n11882) );
  NAND2_X1 U14491 ( .A1(n11802), .A2(n11801), .ZN(n11858) );
  INV_X1 U14492 ( .A(n11858), .ZN(n11803) );
  NAND2_X1 U14493 ( .A1(n11856), .A2(n11957), .ZN(n11805) );
  NAND2_X1 U14494 ( .A1(n11805), .A2(n11804), .ZN(n11960) );
  OR2_X1 U14495 ( .A1(n15099), .A2(n7220), .ZN(n11806) );
  XOR2_X1 U14496 ( .A(n12019), .B(n11807), .Z(n11880) );
  NAND2_X1 U14497 ( .A1(n11853), .A2(n15834), .ZN(n11963) );
  NAND2_X1 U14498 ( .A1(n11964), .A2(n12028), .ZN(n11808) );
  NAND2_X1 U14499 ( .A1(n11808), .A2(n7132), .ZN(n11809) );
  NOR2_X1 U14500 ( .A1(n6605), .A2(n11809), .ZN(n11876) );
  OR2_X1 U14501 ( .A1(n12030), .A2(n15516), .ZN(n11811) );
  NAND2_X1 U14502 ( .A1(n15099), .A2(n15521), .ZN(n11810) );
  NAND2_X1 U14503 ( .A1(n11811), .A2(n11810), .ZN(n12070) );
  INV_X1 U14504 ( .A(n12070), .ZN(n11874) );
  OAI21_X1 U14505 ( .B1(n15844), .B2(n15792), .A(n11874), .ZN(n11812) );
  AOI211_X1 U14506 ( .C1(n11880), .C2(n15611), .A(n11876), .B(n11812), .ZN(
        n11813) );
  OAI21_X1 U14507 ( .B1(n15874), .B2(n11882), .A(n11813), .ZN(n11846) );
  NAND2_X1 U14508 ( .A1(n11846), .A2(n15877), .ZN(n11814) );
  OAI21_X1 U14509 ( .B1(n15877), .B2(n9543), .A(n11814), .ZN(P1_U3471) );
  OAI21_X1 U14510 ( .B1(n11815), .B2(n14338), .A(n12221), .ZN(n12540) );
  AOI211_X1 U14511 ( .C1(n14136), .C2(n11816), .A(n14717), .B(n7898), .ZN(
        n12533) );
  XNOR2_X1 U14512 ( .A(n11817), .B(n14338), .ZN(n11819) );
  OAI21_X1 U14513 ( .B1(n11819), .B2(n8640), .A(n11818), .ZN(n12537) );
  AOI211_X1 U14514 ( .C1(n15993), .C2(n12540), .A(n12533), .B(n12537), .ZN(
        n11826) );
  INV_X1 U14515 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n11820) );
  OAI22_X1 U14516 ( .A1(n14892), .A2(n7190), .B1(n16004), .B2(n11820), .ZN(
        n11821) );
  INV_X1 U14517 ( .A(n11821), .ZN(n11822) );
  OAI21_X1 U14518 ( .B1(n11826), .B2(n16002), .A(n11822), .ZN(P2_U3442) );
  OAI22_X1 U14519 ( .A1(n14840), .A2(n7190), .B1(n16011), .B2(n11823), .ZN(
        n11824) );
  INV_X1 U14520 ( .A(n11824), .ZN(n11825) );
  OAI21_X1 U14521 ( .B1(n11826), .B2(n16008), .A(n11825), .ZN(P2_U3503) );
  NAND2_X1 U14522 ( .A1(n11828), .A2(n11827), .ZN(n11852) );
  OAI22_X1 U14523 ( .A1(n15528), .A2(n11833), .B1(n15100), .B2(n15804), .ZN(
        n11834) );
  AOI21_X1 U14524 ( .B1(n15496), .B2(n11483), .A(n11834), .ZN(n11840) );
  OAI21_X1 U14525 ( .B1(n11835), .B2(n11837), .A(n11836), .ZN(n11838) );
  NAND2_X1 U14526 ( .A1(n11838), .A2(n15528), .ZN(n11839) );
  OAI211_X1 U14527 ( .C1(n15535), .C2(n11841), .A(n11840), .B(n11839), .ZN(
        P1_U3292) );
  NOR2_X1 U14528 ( .A1(n16106), .A2(n8918), .ZN(n11842) );
  AOI21_X1 U14529 ( .B1(n11843), .B2(n16106), .A(n11842), .ZN(n11844) );
  OAI21_X1 U14530 ( .B1(n11845), .B2(n13860), .A(n11844), .ZN(P3_U3459) );
  NAND2_X1 U14531 ( .A1(n11846), .A2(n15886), .ZN(n11847) );
  OAI21_X1 U14532 ( .B1(n15886), .B2(n11066), .A(n11847), .ZN(P1_U3532) );
  OAI21_X1 U14533 ( .B1(n11848), .B2(n11859), .A(n11849), .ZN(n15831) );
  INV_X1 U14534 ( .A(n15831), .ZN(n11865) );
  NOR2_X1 U14535 ( .A1(n6556), .A2(n11850), .ZN(n15813) );
  INV_X1 U14536 ( .A(n15813), .ZN(n15445) );
  OAI211_X1 U14537 ( .C1(n11853), .C2(n15834), .A(n7132), .B(n11963), .ZN(
        n15832) );
  OAI22_X1 U14538 ( .A1(n15344), .A2(n15832), .B1(n15121), .B2(n15804), .ZN(
        n11855) );
  NOR2_X1 U14539 ( .A1(n15807), .A2(n15834), .ZN(n11854) );
  AOI211_X1 U14540 ( .C1(n6556), .C2(P1_REG2_REG_2__SCAN_IN), .A(n11855), .B(
        n11854), .ZN(n11864) );
  INV_X1 U14541 ( .A(n11856), .ZN(n11857) );
  AOI21_X1 U14542 ( .B1(n11859), .B2(n11858), .A(n11857), .ZN(n11862) );
  AOI22_X1 U14543 ( .A1(n10118), .A2(n15521), .B1(n15500), .B2(n15099), .ZN(
        n11861) );
  INV_X1 U14544 ( .A(n15436), .ZN(n15850) );
  NAND2_X1 U14545 ( .A1(n15831), .A2(n15850), .ZN(n11860) );
  OAI211_X1 U14546 ( .C1(n11862), .C2(n15826), .A(n11861), .B(n11860), .ZN(
        n15836) );
  NAND2_X1 U14547 ( .A1(n15836), .A2(n15528), .ZN(n11863) );
  OAI211_X1 U14548 ( .C1(n11865), .C2(n15445), .A(n11864), .B(n11863), .ZN(
        P1_U3291) );
  OAI21_X1 U14549 ( .B1(n11867), .B2(n13315), .A(n11866), .ZN(n12077) );
  NOR2_X1 U14550 ( .A1(n11868), .A2(n13315), .ZN(n12127) );
  NAND2_X1 U14551 ( .A1(n11868), .A2(n13315), .ZN(n11869) );
  NAND2_X1 U14552 ( .A1(n11869), .A2(n16044), .ZN(n11870) );
  OR2_X1 U14553 ( .A1(n12127), .A2(n11870), .ZN(n11872) );
  AOI22_X1 U14554 ( .A1(n16046), .A2(n13506), .B1(n13508), .B2(n16049), .ZN(
        n11871) );
  NAND2_X1 U14555 ( .A1(n11872), .A2(n11871), .ZN(n12074) );
  AOI21_X1 U14556 ( .B1(n12077), .B2(n16070), .A(n12074), .ZN(n11953) );
  AOI22_X1 U14557 ( .A1(n13953), .A2(n12289), .B1(n16092), .B2(
        P3_REG0_REG_6__SCAN_IN), .ZN(n11873) );
  OAI21_X1 U14558 ( .B1(n11953), .B2(n16092), .A(n11873), .ZN(P3_U3408) );
  NOR2_X1 U14559 ( .A1(n6556), .A2(n15826), .ZN(n15428) );
  OAI22_X1 U14560 ( .A1(n6556), .A2(n11874), .B1(n12073), .B2(n15804), .ZN(
        n11875) );
  AOI21_X1 U14561 ( .B1(P1_REG2_REG_4__SCAN_IN), .B2(n6556), .A(n11875), .ZN(
        n11878) );
  NAND2_X1 U14562 ( .A1(n11876), .A2(n15812), .ZN(n11877) );
  OAI211_X1 U14563 ( .C1(n15792), .C2(n15807), .A(n11878), .B(n11877), .ZN(
        n11879) );
  AOI21_X1 U14564 ( .B1(n11880), .B2(n15428), .A(n11879), .ZN(n11881) );
  OAI21_X1 U14565 ( .B1(n15535), .B2(n11882), .A(n11881), .ZN(P1_U3289) );
  MUX2_X1 U14566 ( .A(n11884), .B(n11883), .S(n16066), .Z(n11888) );
  AOI22_X1 U14567 ( .A1(n13814), .A2(n11886), .B1(n16061), .B2(n11885), .ZN(
        n11887) );
  OAI211_X1 U14568 ( .C1(n13824), .C2(n11889), .A(n11888), .B(n11887), .ZN(
        P3_U3229) );
  XNOR2_X1 U14569 ( .A(n12164), .B(P1_REG1_REG_13__SCAN_IN), .ZN(n11894) );
  OR2_X1 U14570 ( .A1(n11895), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n11890) );
  INV_X1 U14571 ( .A(n12166), .ZN(n11892) );
  AOI211_X1 U14572 ( .C1(n11894), .C2(n11893), .A(n15248), .B(n11892), .ZN(
        n11905) );
  MUX2_X1 U14573 ( .A(n15529), .B(P1_REG2_REG_13__SCAN_IN), .S(n12164), .Z(
        n11900) );
  OR2_X1 U14574 ( .A1(n11895), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n11896) );
  NAND2_X1 U14575 ( .A1(n11897), .A2(n11896), .ZN(n11899) );
  INV_X1 U14576 ( .A(n12161), .ZN(n11898) );
  AOI211_X1 U14577 ( .C1(n11900), .C2(n11899), .A(n15242), .B(n11898), .ZN(
        n11904) );
  NAND2_X1 U14578 ( .A1(P1_U3086), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n15035)
         );
  NAND2_X1 U14579 ( .A1(n15149), .A2(P1_ADDR_REG_13__SCAN_IN), .ZN(n11901) );
  OAI211_X1 U14580 ( .C1(n15246), .C2(n11902), .A(n15035), .B(n11901), .ZN(
        n11903) );
  OR3_X1 U14581 ( .A1(n11905), .A2(n11904), .A3(n11903), .ZN(P1_U3256) );
  NAND2_X1 U14582 ( .A1(n11906), .A2(n14106), .ZN(n14330) );
  INV_X1 U14583 ( .A(n14330), .ZN(n12159) );
  NAND2_X1 U14584 ( .A1(n8640), .A2(n10420), .ZN(n11908) );
  AOI21_X1 U14585 ( .B1(n14330), .B2(n11908), .A(n11907), .ZN(n12154) );
  NAND2_X1 U14586 ( .A1(n14108), .A2(n11909), .ZN(n12155) );
  OAI211_X1 U14587 ( .C1(n12159), .C2(n14846), .A(n12154), .B(n12155), .ZN(
        n11922) );
  NAND2_X1 U14588 ( .A1(n16004), .A2(n11922), .ZN(n11910) );
  OAI21_X1 U14589 ( .B1(n16004), .B2(n11911), .A(n11910), .ZN(P2_U3430) );
  XNOR2_X1 U14590 ( .A(n11436), .B(n12099), .ZN(n12247) );
  XNOR2_X1 U14591 ( .A(n13508), .B(n12247), .ZN(n11914) );
  AOI21_X1 U14592 ( .B1(n11915), .B2(n11914), .A(n12281), .ZN(n11921) );
  INV_X1 U14593 ( .A(n12100), .ZN(n11919) );
  AOI22_X1 U14594 ( .A1(n13247), .A2(n13507), .B1(n13269), .B2(n13509), .ZN(
        n11917) );
  OAI211_X1 U14595 ( .C1(n13276), .C2(n12099), .A(n11917), .B(n11916), .ZN(
        n11918) );
  AOI21_X1 U14596 ( .B1(n11919), .B2(n13273), .A(n11918), .ZN(n11920) );
  OAI21_X1 U14597 ( .B1(n11921), .B2(n13264), .A(n11920), .ZN(P3_U3167) );
  NAND2_X1 U14598 ( .A1(n16011), .A2(n11922), .ZN(n11923) );
  OAI21_X1 U14599 ( .B1(n16011), .B2(n11189), .A(n11923), .ZN(P2_U3499) );
  NAND2_X1 U14600 ( .A1(n11927), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n11924) );
  XNOR2_X1 U14601 ( .A(n11986), .B(P2_REG2_REG_14__SCAN_IN), .ZN(n11937) );
  NAND2_X1 U14602 ( .A1(P2_U3088), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n13982)
         );
  OAI21_X1 U14603 ( .B1(n15919), .B2(n11926), .A(n13982), .ZN(n11935) );
  NAND2_X1 U14604 ( .A1(n11927), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n11928) );
  NAND2_X1 U14605 ( .A1(n11929), .A2(n11928), .ZN(n11932) );
  INV_X1 U14606 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n11930) );
  XNOR2_X1 U14607 ( .A(n11993), .B(n11930), .ZN(n11931) );
  NAND2_X1 U14608 ( .A1(n11932), .A2(n11931), .ZN(n11995) );
  OAI211_X1 U14609 ( .C1(n11932), .C2(n11931), .A(n11995), .B(n15928), .ZN(
        n11933) );
  INV_X1 U14610 ( .A(n11933), .ZN(n11934) );
  AOI211_X1 U14611 ( .C1(n15899), .C2(P2_ADDR_REG_14__SCAN_IN), .A(n11935), 
        .B(n11934), .ZN(n11936) );
  OAI21_X1 U14612 ( .B1(n11937), .B2(n14504), .A(n11936), .ZN(P2_U3228) );
  NAND2_X1 U14613 ( .A1(n11938), .A2(n13966), .ZN(n11939) );
  OAI211_X1 U14614 ( .C1(n11940), .C2(n13962), .A(n11939), .B(n13490), .ZN(
        P3_U3272) );
  INV_X1 U14615 ( .A(n11942), .ZN(n11943) );
  OR2_X1 U14616 ( .A1(n11944), .A2(n11943), .ZN(n11945) );
  INV_X1 U14617 ( .A(P3_ADDR_REG_9__SCAN_IN), .ZN(n11948) );
  XNOR2_X1 U14618 ( .A(n11948), .B(P1_ADDR_REG_9__SCAN_IN), .ZN(n12006) );
  XNOR2_X1 U14619 ( .A(n12007), .B(n12006), .ZN(n12002) );
  NAND2_X1 U14620 ( .A1(n11949), .A2(P2_ADDR_REG_9__SCAN_IN), .ZN(n12005) );
  OAI21_X1 U14621 ( .B1(n11949), .B2(P2_ADDR_REG_9__SCAN_IN), .A(n12005), .ZN(
        n11950) );
  INV_X1 U14622 ( .A(n11950), .ZN(SUB_1596_U54) );
  OAI22_X1 U14623 ( .A1(n13860), .A2(n12245), .B1(n16106), .B2(n8854), .ZN(
        n11951) );
  INV_X1 U14624 ( .A(n11951), .ZN(n11952) );
  OAI21_X1 U14625 ( .B1(n11953), .B2(n16103), .A(n11952), .ZN(P3_U3465) );
  OAI21_X1 U14626 ( .B1(n11955), .B2(n11958), .A(n11954), .ZN(n15841) );
  OAI22_X1 U14627 ( .A1(n11956), .A2(n15431), .B1(n15793), .B2(n15516), .ZN(
        n11962) );
  NAND3_X1 U14628 ( .A1(n11856), .A2(n11958), .A3(n11957), .ZN(n11959) );
  AOI21_X1 U14629 ( .B1(n11960), .B2(n11959), .A(n15826), .ZN(n11961) );
  AOI211_X1 U14630 ( .C1(n15850), .C2(n15841), .A(n11962), .B(n11961), .ZN(
        n15838) );
  OAI211_X1 U14631 ( .C1(n7450), .C2(n7220), .A(n7132), .B(n11964), .ZN(n15837) );
  NAND2_X1 U14632 ( .A1(n15496), .A2(n11965), .ZN(n11968) );
  INV_X1 U14633 ( .A(n15804), .ZN(n15525) );
  AOI22_X1 U14634 ( .A1(n6556), .A2(P1_REG2_REG_3__SCAN_IN), .B1(n15525), .B2(
        n11966), .ZN(n11967) );
  OAI211_X1 U14635 ( .C1(n15837), .C2(n15344), .A(n11968), .B(n11967), .ZN(
        n11969) );
  AOI21_X1 U14636 ( .B1(n15813), .B2(n15841), .A(n11969), .ZN(n11970) );
  OAI21_X1 U14637 ( .B1(n15838), .B2(n6556), .A(n11970), .ZN(P1_U3290) );
  OAI222_X1 U14638 ( .A1(n13134), .A2(n11971), .B1(n15703), .B2(n11973), .C1(
        P1_U3086), .C2(n6868), .ZN(P1_U3337) );
  INV_X1 U14639 ( .A(n12806), .ZN(n12801) );
  OAI222_X1 U14640 ( .A1(P2_U3088), .A2(n12801), .B1(n14903), .B2(n11973), 
        .C1(n11972), .C2(n14914), .ZN(P2_U3309) );
  OAI22_X1 U14641 ( .A1(n13860), .A2(n11974), .B1(n16106), .B2(n8846), .ZN(
        n11975) );
  AOI21_X1 U14642 ( .B1(n11976), .B2(n16106), .A(n11975), .ZN(n11977) );
  INV_X1 U14643 ( .A(n11977), .ZN(P3_U3463) );
  XNOR2_X1 U14644 ( .A(n11978), .B(n11979), .ZN(n11985) );
  NAND2_X1 U14645 ( .A1(n14414), .A2(n14086), .ZN(n11981) );
  NAND2_X1 U14646 ( .A1(n14416), .A2(n14376), .ZN(n11980) );
  AND2_X1 U14647 ( .A1(n11981), .A2(n11980), .ZN(n12235) );
  OAI22_X1 U14648 ( .A1(n14090), .A2(n12235), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8143), .ZN(n11983) );
  NOR2_X1 U14649 ( .A1(n14073), .A2(n12241), .ZN(n11982) );
  AOI211_X1 U14650 ( .C1(n14088), .C2(n12239), .A(n11983), .B(n11982), .ZN(
        n11984) );
  OAI21_X1 U14651 ( .B1(n11985), .B2(n14103), .A(n11984), .ZN(P2_U3185) );
  NAND2_X1 U14652 ( .A1(n11986), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n11989) );
  NAND2_X1 U14653 ( .A1(n11987), .A2(n11993), .ZN(n11988) );
  NAND2_X1 U14654 ( .A1(n11989), .A2(n11988), .ZN(n12680) );
  XNOR2_X1 U14655 ( .A(n12680), .B(n11996), .ZN(n12678) );
  XNOR2_X1 U14656 ( .A(n12678), .B(P2_REG2_REG_15__SCAN_IN), .ZN(n12000) );
  NOR2_X1 U14657 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n11990), .ZN(n11992) );
  NOR2_X1 U14658 ( .A1(n15919), .A2(n11996), .ZN(n11991) );
  AOI211_X1 U14659 ( .C1(n15899), .C2(P2_ADDR_REG_15__SCAN_IN), .A(n11992), 
        .B(n11991), .ZN(n11999) );
  NAND2_X1 U14660 ( .A1(n11993), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n11994) );
  NAND2_X1 U14661 ( .A1(n11995), .A2(n11994), .ZN(n12669) );
  XNOR2_X1 U14662 ( .A(n12669), .B(n11996), .ZN(n11997) );
  NAND2_X1 U14663 ( .A1(n11997), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n12671) );
  OAI211_X1 U14664 ( .C1(n11997), .C2(P2_REG1_REG_15__SCAN_IN), .A(n12671), 
        .B(n15928), .ZN(n11998) );
  OAI211_X1 U14665 ( .C1(n12000), .C2(n14504), .A(n11999), .B(n11998), .ZN(
        P2_U3229) );
  INV_X1 U14666 ( .A(n12001), .ZN(n12003) );
  NAND2_X1 U14667 ( .A1(n12003), .A2(n12002), .ZN(n12004) );
  NAND2_X1 U14668 ( .A1(n12008), .A2(P3_ADDR_REG_9__SCAN_IN), .ZN(n12009) );
  INV_X1 U14669 ( .A(P3_ADDR_REG_10__SCAN_IN), .ZN(n12011) );
  NAND2_X1 U14670 ( .A1(n12011), .A2(P1_ADDR_REG_10__SCAN_IN), .ZN(n12328) );
  INV_X1 U14671 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n12012) );
  NAND2_X1 U14672 ( .A1(n12012), .A2(P3_ADDR_REG_10__SCAN_IN), .ZN(n12013) );
  NAND2_X1 U14673 ( .A1(n12328), .A2(n12013), .ZN(n12014) );
  NAND2_X1 U14674 ( .A1(n12015), .A2(n12014), .ZN(n12016) );
  NAND2_X1 U14675 ( .A1(n12329), .A2(n12016), .ZN(n12326) );
  XNOR2_X1 U14676 ( .A(n12326), .B(n12325), .ZN(n12017) );
  XNOR2_X1 U14677 ( .A(n12324), .B(n12017), .ZN(SUB_1596_U70) );
  NAND2_X1 U14678 ( .A1(n15795), .A2(n15792), .ZN(n12018) );
  OR2_X1 U14679 ( .A1(n15795), .A2(n15792), .ZN(n12020) );
  NAND2_X1 U14680 ( .A1(n12030), .A2(n12091), .ZN(n12021) );
  XNOR2_X1 U14681 ( .A(n12196), .B(n12195), .ZN(n12025) );
  OR2_X1 U14682 ( .A1(n12030), .A2(n15431), .ZN(n12024) );
  NAND2_X1 U14683 ( .A1(n15096), .A2(n15500), .ZN(n12023) );
  NAND2_X1 U14684 ( .A1(n12024), .A2(n12023), .ZN(n12174) );
  AOI21_X1 U14685 ( .B1(n12025), .B2(n15611), .A(n12174), .ZN(n15859) );
  AOI22_X1 U14686 ( .A1(n15098), .A2(n12091), .B1(n12028), .B2(n15795), .ZN(
        n12026) );
  INV_X1 U14687 ( .A(n12029), .ZN(n12031) );
  XNOR2_X1 U14688 ( .A(n12212), .B(n12211), .ZN(n15852) );
  INV_X1 U14689 ( .A(n15853), .ZN(n12035) );
  OAI211_X1 U14690 ( .C1(n15809), .C2(n12035), .A(n7132), .B(n12206), .ZN(
        n15855) );
  OAI22_X1 U14691 ( .A1(n15528), .A2(n12036), .B1(n12176), .B2(n15804), .ZN(
        n12037) );
  AOI21_X1 U14692 ( .B1(n15496), .B2(n15853), .A(n12037), .ZN(n12038) );
  OAI21_X1 U14693 ( .B1(n15344), .B2(n15855), .A(n12038), .ZN(n12039) );
  AOI21_X1 U14694 ( .B1(n15852), .B2(n15513), .A(n12039), .ZN(n12040) );
  OAI21_X1 U14695 ( .B1(n15859), .B2(n6556), .A(n12040), .ZN(P1_U3287) );
  NOR2_X1 U14696 ( .A1(n15428), .A2(n15513), .ZN(n12047) );
  OAI22_X1 U14697 ( .A1(n6556), .A2(n12042), .B1(n12041), .B2(n15804), .ZN(
        n12045) );
  INV_X1 U14698 ( .A(n7132), .ZN(n15608) );
  NOR2_X1 U14699 ( .A1(n15344), .A2(n15608), .ZN(n13086) );
  INV_X1 U14700 ( .A(n13086), .ZN(n15426) );
  AOI21_X1 U14701 ( .B1(n15426), .B2(n15807), .A(n12043), .ZN(n12044) );
  AOI211_X1 U14702 ( .C1(n6556), .C2(P1_REG2_REG_0__SCAN_IN), .A(n12045), .B(
        n12044), .ZN(n12046) );
  OAI21_X1 U14703 ( .B1(n15825), .B2(n12047), .A(n12046), .ZN(P1_U3293) );
  AOI21_X1 U14704 ( .B1(n12050), .B2(n12049), .A(n12048), .ZN(n12065) );
  OAI21_X1 U14705 ( .B1(P3_REG2_REG_9__SCAN_IN), .B2(n12052), .A(n12051), .ZN(
        n12060) );
  INV_X1 U14706 ( .A(n12053), .ZN(n12054) );
  NAND3_X1 U14707 ( .A1(n12056), .A2(n12055), .A3(n12054), .ZN(n12057) );
  AOI21_X1 U14708 ( .B1(n12058), .B2(n12057), .A(n16013), .ZN(n12059) );
  AOI21_X1 U14709 ( .B1(n12060), .B2(n13583), .A(n12059), .ZN(n12064) );
  AND2_X1 U14710 ( .A1(P3_U3151), .A2(P3_REG3_REG_9__SCAN_IN), .ZN(n12260) );
  NOR2_X1 U14711 ( .A1(n13617), .A2(n12061), .ZN(n12062) );
  AOI211_X1 U14712 ( .C1(n16012), .C2(P3_ADDR_REG_9__SCAN_IN), .A(n12260), .B(
        n12062), .ZN(n12063) );
  OAI211_X1 U14713 ( .C1(n12065), .C2(n16015), .A(n12064), .B(n12063), .ZN(
        P3_U3191) );
  XNOR2_X1 U14714 ( .A(n7155), .B(n12066), .ZN(n12082) );
  XNOR2_X1 U14715 ( .A(n12082), .B(n12067), .ZN(n12068) );
  NAND2_X1 U14716 ( .A1(n12068), .A2(n15072), .ZN(n12072) );
  AND2_X1 U14717 ( .A1(P1_U3086), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n15148) );
  NOR2_X1 U14718 ( .A1(n15083), .A2(n15792), .ZN(n12069) );
  AOI211_X1 U14719 ( .C1(n15080), .C2(n12070), .A(n15148), .B(n12069), .ZN(
        n12071) );
  OAI211_X1 U14720 ( .C1(n15077), .C2(n12073), .A(n12072), .B(n12071), .ZN(
        P1_U3230) );
  OAI22_X1 U14721 ( .A1(n13737), .A2(n12245), .B1(n12292), .B2(n12707), .ZN(
        n12076) );
  MUX2_X1 U14722 ( .A(n12074), .B(P3_REG2_REG_6__SCAN_IN), .S(n16066), .Z(
        n12075) );
  AOI211_X1 U14723 ( .C1(n9427), .C2(n12077), .A(n12076), .B(n12075), .ZN(
        n12078) );
  INV_X1 U14724 ( .A(n12078), .ZN(P3_U3227) );
  AOI22_X1 U14725 ( .A1(n12082), .A2(n12081), .B1(n12080), .B2(n7155), .ZN(
        n12087) );
  OAI21_X1 U14726 ( .B1(n12085), .B2(n12084), .A(n12083), .ZN(n12086) );
  XNOR2_X1 U14727 ( .A(n12087), .B(n12086), .ZN(n12093) );
  AOI22_X1 U14728 ( .A1(n15521), .A2(n15795), .B1(n15097), .B2(n15500), .ZN(
        n15800) );
  OAI21_X1 U14729 ( .B1(n15025), .B2(n15800), .A(n12088), .ZN(n12090) );
  NOR2_X1 U14730 ( .A1(n15077), .A2(n15803), .ZN(n12089) );
  AOI211_X1 U14731 ( .C1(n15068), .C2(n12091), .A(n12090), .B(n12089), .ZN(
        n12092) );
  OAI21_X1 U14732 ( .B1(n12093), .B2(n15070), .A(n12092), .ZN(P1_U3227) );
  NAND2_X1 U14733 ( .A1(n13722), .A2(P3_U3897), .ZN(n12094) );
  OAI21_X1 U14734 ( .B1(P3_U3897), .B2(n12095), .A(n12094), .ZN(P3_U3514) );
  OAI222_X1 U14735 ( .A1(n12097), .A2(P1_U3086), .B1(n15703), .B2(n12183), 
        .C1(n12096), .C2(n15700), .ZN(P1_U3335) );
  XNOR2_X1 U14736 ( .A(n12098), .B(n13313), .ZN(n16077) );
  INV_X1 U14737 ( .A(n12629), .ZN(n16062) );
  OR2_X1 U14738 ( .A1(n12099), .A2(n16055), .ZN(n16076) );
  OAI22_X1 U14739 ( .A1(n12133), .A2(n16076), .B1(n12100), .B2(n12707), .ZN(
        n12108) );
  OAI21_X1 U14740 ( .B1(n11638), .B2(n12102), .A(n12101), .ZN(n12103) );
  XNOR2_X1 U14741 ( .A(n13313), .B(n12103), .ZN(n12106) );
  NAND2_X1 U14742 ( .A1(n16077), .A2(n16054), .ZN(n12105) );
  AOI22_X1 U14743 ( .A1(n16046), .A2(n13507), .B1(n13509), .B2(n16049), .ZN(
        n12104) );
  OAI211_X1 U14744 ( .C1(n16034), .C2(n12106), .A(n12105), .B(n12104), .ZN(
        n16080) );
  MUX2_X1 U14745 ( .A(P3_REG2_REG_5__SCAN_IN), .B(n16080), .S(n9401), .Z(
        n12107) );
  AOI211_X1 U14746 ( .C1(n16077), .C2(n16062), .A(n12108), .B(n12107), .ZN(
        n12109) );
  INV_X1 U14747 ( .A(n12109), .ZN(P3_U3228) );
  XNOR2_X1 U14748 ( .A(n12110), .B(n13381), .ZN(n13884) );
  INV_X1 U14749 ( .A(n13884), .ZN(n12120) );
  INV_X1 U14750 ( .A(n12111), .ZN(n12263) );
  AOI22_X1 U14751 ( .A1(n13814), .A2(n12112), .B1(n16061), .B2(n12263), .ZN(
        n12119) );
  AOI21_X1 U14752 ( .B1(n12113), .B2(n13381), .A(n16034), .ZN(n12116) );
  INV_X1 U14753 ( .A(n13505), .ZN(n12309) );
  OAI22_X1 U14754 ( .A1(n12309), .A2(n13815), .B1(n12258), .B2(n13817), .ZN(
        n12115) );
  AOI21_X1 U14755 ( .B1(n12116), .B2(n12114), .A(n12115), .ZN(n13885) );
  MUX2_X1 U14756 ( .A(n12117), .B(n13885), .S(n9401), .Z(n12118) );
  OAI211_X1 U14757 ( .C1(n12120), .C2(n13824), .A(n12119), .B(n12118), .ZN(
        P3_U3224) );
  MUX2_X1 U14758 ( .A(n12121), .B(P3_REG1_REG_3__SCAN_IN), .S(n16103), .Z(
        n12122) );
  AOI21_X1 U14759 ( .B1(n13880), .B2(n12123), .A(n12122), .ZN(n12124) );
  INV_X1 U14760 ( .A(n12124), .ZN(P3_U3462) );
  XNOR2_X1 U14761 ( .A(n12125), .B(n13370), .ZN(n16085) );
  INV_X1 U14762 ( .A(n16085), .ZN(n12138) );
  NOR2_X1 U14763 ( .A1(n12127), .A2(n12126), .ZN(n12128) );
  XNOR2_X1 U14764 ( .A(n12128), .B(n13370), .ZN(n12130) );
  AOI22_X1 U14765 ( .A1(n16049), .A2(n13507), .B1(n13505), .B2(n16046), .ZN(
        n12129) );
  OAI21_X1 U14766 ( .B1(n12130), .B2(n16034), .A(n12129), .ZN(n12131) );
  AOI21_X1 U14767 ( .B1(n16085), .B2(n16054), .A(n12131), .ZN(n16082) );
  MUX2_X1 U14768 ( .A(n12132), .B(n16082), .S(n9401), .Z(n12137) );
  INV_X1 U14769 ( .A(n12133), .ZN(n12276) );
  NOR2_X1 U14770 ( .A1(n12134), .A2(n16055), .ZN(n16084) );
  INV_X1 U14771 ( .A(n12316), .ZN(n12135) );
  AOI22_X1 U14772 ( .A1(n12276), .A2(n16084), .B1(n16061), .B2(n12135), .ZN(
        n12136) );
  OAI211_X1 U14773 ( .C1(n12138), .C2(n12629), .A(n12137), .B(n12136), .ZN(
        P3_U3226) );
  INV_X1 U14774 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n12139) );
  OAI222_X1 U14775 ( .A1(n12140), .A2(P1_U3086), .B1(n15703), .B2(n12143), 
        .C1(n12139), .C2(n13134), .ZN(P1_U3334) );
  INV_X1 U14776 ( .A(n12141), .ZN(n13104) );
  OAI222_X1 U14777 ( .A1(P1_U3086), .A2(n9780), .B1(n15703), .B2(n13104), .C1(
        n12142), .C2(n15700), .ZN(P1_U3336) );
  OAI222_X1 U14778 ( .A1(n14914), .A2(n12144), .B1(P2_U3088), .B2(n7517), .C1(
        n14903), .C2(n12143), .ZN(P2_U3306) );
  INV_X1 U14779 ( .A(n12910), .ZN(n12751) );
  NAND2_X1 U14780 ( .A1(n15780), .A2(n15870), .ZN(n15860) );
  OAI211_X1 U14781 ( .C1(n12147), .C2(n12146), .A(n12145), .B(n15072), .ZN(
        n12152) );
  INV_X1 U14782 ( .A(n15781), .ZN(n12150) );
  AOI22_X1 U14783 ( .A1(n15521), .A2(n15097), .B1(n15095), .B2(n15500), .ZN(
        n15861) );
  OAI22_X1 U14784 ( .A1(n15025), .A2(n15861), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n12148), .ZN(n12149) );
  AOI21_X1 U14785 ( .B1(n12150), .B2(n15061), .A(n12149), .ZN(n12151) );
  OAI211_X1 U14786 ( .C1(n12751), .C2(n15860), .A(n12152), .B(n12151), .ZN(
        P1_U3213) );
  OAI21_X1 U14787 ( .B1(n14383), .B2(n12155), .A(n12154), .ZN(n12156) );
  AOI22_X1 U14788 ( .A1(n6548), .A2(n12156), .B1(P2_REG3_REG_0__SCAN_IN), .B2(
        n14713), .ZN(n12158) );
  NAND2_X1 U14789 ( .A1(n14719), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n12157) );
  OAI211_X1 U14790 ( .C1(n14682), .C2(n12159), .A(n12158), .B(n12157), .ZN(
        P2_U3265) );
  NAND2_X1 U14791 ( .A1(n12164), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n12160) );
  NAND2_X1 U14792 ( .A1(n12161), .A2(n12160), .ZN(n15194) );
  XNOR2_X1 U14793 ( .A(n15191), .B(n12162), .ZN(n15193) );
  NAND2_X1 U14794 ( .A1(n15194), .A2(n15193), .ZN(n15192) );
  NAND2_X1 U14795 ( .A1(n15191), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n12163) );
  NAND2_X1 U14796 ( .A1(n15192), .A2(n12163), .ZN(n12645) );
  XNOR2_X1 U14797 ( .A(n12645), .B(n12633), .ZN(n12643) );
  XNOR2_X1 U14798 ( .A(n12643), .B(P1_REG2_REG_15__SCAN_IN), .ZN(n12173) );
  NAND2_X1 U14799 ( .A1(n12164), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n12165) );
  XNOR2_X1 U14800 ( .A(n15191), .B(n12167), .ZN(n15187) );
  NAND2_X1 U14801 ( .A1(n15186), .A2(n15187), .ZN(n15185) );
  OR2_X1 U14802 ( .A1(n15191), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n12168) );
  NAND2_X1 U14803 ( .A1(n15185), .A2(n12168), .ZN(n12634) );
  XNOR2_X1 U14804 ( .A(n12632), .B(n12631), .ZN(n12169) );
  NAND2_X1 U14805 ( .A1(n12169), .A2(n15218), .ZN(n12172) );
  AND2_X1 U14806 ( .A1(P1_U3086), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n15079) );
  NOR2_X1 U14807 ( .A1(n15252), .A2(n15732), .ZN(n12170) );
  AOI211_X1 U14808 ( .C1(n12644), .C2(n15223), .A(n15079), .B(n12170), .ZN(
        n12171) );
  OAI211_X1 U14809 ( .C1(n12173), .C2(n15242), .A(n12172), .B(n12171), .ZN(
        P1_U3258) );
  AOI22_X1 U14810 ( .A1(n15080), .A2(n12174), .B1(P1_REG3_REG_6__SCAN_IN), 
        .B2(P1_U3086), .ZN(n12175) );
  OAI21_X1 U14811 ( .B1(n15077), .B2(n12176), .A(n12175), .ZN(n12181) );
  INV_X1 U14812 ( .A(n12177), .ZN(n12178) );
  AOI211_X1 U14813 ( .C1(n6728), .C2(n12179), .A(n15070), .B(n12178), .ZN(
        n12180) );
  AOI211_X1 U14814 ( .C1(n15068), .C2(n15853), .A(n12181), .B(n12180), .ZN(
        n12182) );
  INV_X1 U14815 ( .A(n12182), .ZN(P1_U3239) );
  OAI222_X1 U14816 ( .A1(n14914), .A2(n12184), .B1(P2_U3088), .B2(n14329), 
        .C1(n14903), .C2(n12183), .ZN(P2_U3307) );
  INV_X1 U14817 ( .A(n12185), .ZN(n12186) );
  AOI21_X1 U14818 ( .B1(n14341), .B2(n12187), .A(n12186), .ZN(n12589) );
  OAI211_X1 U14819 ( .C1(n6954), .C2(n7233), .A(n14818), .B(n12384), .ZN(
        n12585) );
  OAI21_X1 U14820 ( .B1(n7233), .B2(n15989), .A(n12585), .ZN(n12191) );
  XNOR2_X1 U14821 ( .A(n12189), .B(n14341), .ZN(n12190) );
  AOI22_X1 U14822 ( .A1(n14376), .A2(n14415), .B1(n14413), .B2(n14086), .ZN(
        n12302) );
  OAI21_X1 U14823 ( .B1(n12190), .B2(n8640), .A(n12302), .ZN(n12586) );
  AOI211_X1 U14824 ( .C1(n12589), .C2(n15993), .A(n12191), .B(n12586), .ZN(
        n12194) );
  NAND2_X1 U14825 ( .A1(n16008), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n12192) );
  OAI21_X1 U14826 ( .B1(n12194), .B2(n16008), .A(n12192), .ZN(P2_U3507) );
  NAND2_X1 U14827 ( .A1(n16002), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n12193) );
  OAI21_X1 U14828 ( .B1(n12194), .B2(n16002), .A(n12193), .ZN(P2_U3454) );
  NAND2_X1 U14829 ( .A1(n12197), .A2(n15853), .ZN(n12198) );
  OR2_X1 U14830 ( .A1(n15780), .A2(n12199), .ZN(n12200) );
  NOR2_X1 U14831 ( .A1(n15869), .A2(n12201), .ZN(n12202) );
  XNOR2_X1 U14832 ( .A(n12360), .B(n12359), .ZN(n12205) );
  NAND2_X1 U14833 ( .A1(n15093), .A2(n15500), .ZN(n12204) );
  NAND2_X1 U14834 ( .A1(n15095), .A2(n15521), .ZN(n12203) );
  NAND2_X1 U14835 ( .A1(n12204), .A2(n12203), .ZN(n12513) );
  AOI21_X1 U14836 ( .B1(n12205), .B2(n15611), .A(n12513), .ZN(n15664) );
  AOI211_X1 U14837 ( .C1(n15662), .C2(n12342), .A(n15608), .B(n12367), .ZN(
        n15661) );
  INV_X1 U14838 ( .A(n15662), .ZN(n12210) );
  INV_X1 U14839 ( .A(n12515), .ZN(n12208) );
  AOI22_X1 U14840 ( .A1(n6556), .A2(P1_REG2_REG_9__SCAN_IN), .B1(n12208), .B2(
        n15525), .ZN(n12209) );
  OAI21_X1 U14841 ( .B1(n15807), .B2(n12210), .A(n12209), .ZN(n12218) );
  OR2_X1 U14842 ( .A1(n15097), .A2(n15853), .ZN(n12213) );
  OR2_X1 U14843 ( .A1(n15780), .A2(n15096), .ZN(n12214) );
  OR2_X1 U14844 ( .A1(n15869), .A2(n15095), .ZN(n12216) );
  XNOR2_X1 U14845 ( .A(n12358), .B(n12359), .ZN(n15665) );
  NOR2_X1 U14846 ( .A1(n15665), .A2(n15535), .ZN(n12217) );
  AOI211_X1 U14847 ( .C1(n15661), .C2(n15812), .A(n12218), .B(n12217), .ZN(
        n12219) );
  OAI21_X1 U14848 ( .B1(n6556), .B2(n15664), .A(n12219), .ZN(P1_U3284) );
  NAND2_X1 U14849 ( .A1(n12221), .A2(n12220), .ZN(n12607) );
  INV_X1 U14850 ( .A(n12607), .ZN(n12608) );
  XNOR2_X1 U14851 ( .A(n14417), .B(n8585), .ZN(n14337) );
  XNOR2_X1 U14852 ( .A(n12608), .B(n14337), .ZN(n15986) );
  XOR2_X1 U14853 ( .A(n12615), .B(n14337), .Z(n12223) );
  AOI21_X1 U14854 ( .B1(n12223), .B2(n14675), .A(n12222), .ZN(n15985) );
  MUX2_X1 U14855 ( .A(n12224), .B(n15985), .S(n6548), .Z(n12229) );
  AOI211_X1 U14856 ( .C1(n15983), .C2(n12225), .A(n14717), .B(n6730), .ZN(
        n15982) );
  OAI22_X1 U14857 ( .A1(n14698), .A2(n8585), .B1(n14736), .B2(n12226), .ZN(
        n12227) );
  AOI21_X1 U14858 ( .B1(n15982), .B2(n14703), .A(n12227), .ZN(n12228) );
  OAI211_X1 U14859 ( .C1(n14742), .C2(n15986), .A(n12229), .B(n12228), .ZN(
        P2_U3260) );
  OAI21_X1 U14860 ( .B1(n12608), .B2(n12231), .A(n12230), .ZN(n12233) );
  INV_X1 U14861 ( .A(n12232), .ZN(n14339) );
  XNOR2_X1 U14862 ( .A(n12233), .B(n14339), .ZN(n15999) );
  XNOR2_X1 U14863 ( .A(n12234), .B(n14339), .ZN(n12237) );
  INV_X1 U14864 ( .A(n12235), .ZN(n12236) );
  AOI21_X1 U14865 ( .B1(n12237), .B2(n14675), .A(n12236), .ZN(n15997) );
  MUX2_X1 U14866 ( .A(n12238), .B(n15997), .S(n6548), .Z(n12244) );
  AOI211_X1 U14867 ( .C1(n15995), .C2(n6604), .A(n14717), .B(n6954), .ZN(
        n15994) );
  INV_X1 U14868 ( .A(n12239), .ZN(n12240) );
  OAI22_X1 U14869 ( .A1(n14698), .A2(n12241), .B1(n14736), .B2(n12240), .ZN(
        n12242) );
  AOI21_X1 U14870 ( .B1(n15994), .B2(n14703), .A(n12242), .ZN(n12243) );
  OAI211_X1 U14871 ( .C1(n14742), .C2(n15999), .A(n12244), .B(n12243), .ZN(
        P2_U3258) );
  XNOR2_X1 U14872 ( .A(n13887), .B(n11436), .ZN(n12484) );
  XNOR2_X1 U14873 ( .A(n12484), .B(n13504), .ZN(n12257) );
  XNOR2_X1 U14874 ( .A(n11436), .B(n12245), .ZN(n12280) );
  XNOR2_X1 U14875 ( .A(n12246), .B(n12957), .ZN(n12472) );
  INV_X1 U14876 ( .A(n12247), .ZN(n12248) );
  NAND2_X1 U14877 ( .A1(n12248), .A2(n12286), .ZN(n12282) );
  XNOR2_X1 U14878 ( .A(n11436), .B(n12274), .ZN(n12253) );
  INV_X1 U14879 ( .A(n12280), .ZN(n12249) );
  INV_X1 U14880 ( .A(n13507), .ZN(n12310) );
  NOR2_X1 U14881 ( .A1(n12249), .A2(n12310), .ZN(n12306) );
  INV_X1 U14882 ( .A(n12472), .ZN(n12250) );
  AOI21_X1 U14883 ( .B1(n12306), .B2(n6630), .A(n12250), .ZN(n12252) );
  AOI21_X1 U14884 ( .B1(n13506), .B2(n6630), .A(n12472), .ZN(n12251) );
  NAND2_X1 U14885 ( .A1(n12253), .A2(n13505), .ZN(n12254) );
  AOI21_X1 U14886 ( .B1(n12257), .B2(n12256), .A(n12486), .ZN(n12265) );
  NOR2_X1 U14887 ( .A1(n13271), .A2(n12258), .ZN(n12259) );
  AOI211_X1 U14888 ( .C1(n13269), .C2(n13505), .A(n12260), .B(n12259), .ZN(
        n12261) );
  OAI21_X1 U14889 ( .B1(n13276), .B2(n13887), .A(n12261), .ZN(n12262) );
  AOI21_X1 U14890 ( .B1(n12263), .B2(n13273), .A(n12262), .ZN(n12264) );
  OAI21_X1 U14891 ( .B1(n12265), .B2(n13264), .A(n12264), .ZN(P3_U3171) );
  XNOR2_X1 U14892 ( .A(n12266), .B(n13373), .ZN(n16091) );
  INV_X1 U14893 ( .A(n16091), .ZN(n12279) );
  OAI21_X1 U14894 ( .B1(n11868), .B2(n12268), .A(n12267), .ZN(n12269) );
  XNOR2_X1 U14895 ( .A(n12269), .B(n13373), .ZN(n12271) );
  AOI22_X1 U14896 ( .A1(n16049), .A2(n13506), .B1(n13504), .B2(n16046), .ZN(
        n12270) );
  OAI21_X1 U14897 ( .B1(n12271), .B2(n16034), .A(n12270), .ZN(n12272) );
  AOI21_X1 U14898 ( .B1(n16091), .B2(n16054), .A(n12272), .ZN(n16087) );
  MUX2_X1 U14899 ( .A(n12273), .B(n16087), .S(n9401), .Z(n12278) );
  NOR2_X1 U14900 ( .A1(n12274), .A2(n16055), .ZN(n16089) );
  INV_X1 U14901 ( .A(n12483), .ZN(n12275) );
  AOI22_X1 U14902 ( .A1(n12276), .A2(n16089), .B1(n16061), .B2(n12275), .ZN(
        n12277) );
  OAI211_X1 U14903 ( .C1(n12279), .C2(n12629), .A(n12278), .B(n12277), .ZN(
        P3_U3225) );
  XNOR2_X1 U14904 ( .A(n12280), .B(n13507), .ZN(n12284) );
  NAND2_X1 U14905 ( .A1(n6768), .A2(n12282), .ZN(n12283) );
  NOR2_X1 U14906 ( .A1(n12283), .A2(n12284), .ZN(n12307) );
  AOI211_X1 U14907 ( .C1(n12284), .C2(n12283), .A(n13264), .B(n12307), .ZN(
        n12285) );
  INV_X1 U14908 ( .A(n12285), .ZN(n12291) );
  INV_X1 U14909 ( .A(n13269), .ZN(n13249) );
  INV_X1 U14910 ( .A(n13506), .ZN(n12477) );
  OAI22_X1 U14911 ( .A1(n13249), .A2(n12286), .B1(n12477), .B2(n13271), .ZN(
        n12287) );
  AOI211_X1 U14912 ( .C1(n12289), .C2(n13261), .A(n12288), .B(n12287), .ZN(
        n12290) );
  OAI211_X1 U14913 ( .C1(n12292), .C2(n13226), .A(n12291), .B(n12290), .ZN(
        P3_U3179) );
  INV_X1 U14914 ( .A(n12293), .ZN(n12295) );
  OAI222_X1 U14915 ( .A1(P3_U3151), .A2(n12296), .B1(n13102), .B2(n12295), 
        .C1(n12294), .C2(n13962), .ZN(P3_U3270) );
  INV_X1 U14916 ( .A(n12298), .ZN(n12299) );
  AOI21_X1 U14917 ( .B1(n12297), .B2(n12300), .A(n12299), .ZN(n12305) );
  NAND2_X1 U14918 ( .A1(n14088), .A2(n12583), .ZN(n12301) );
  NAND2_X1 U14919 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(P2_U3088), .ZN(n14477) );
  OAI211_X1 U14920 ( .C1(n12302), .C2(n14090), .A(n12301), .B(n14477), .ZN(
        n12303) );
  AOI21_X1 U14921 ( .B1(n14154), .B2(n14101), .A(n12303), .ZN(n12304) );
  OAI21_X1 U14922 ( .B1(n12305), .B2(n14103), .A(n12304), .ZN(P2_U3193) );
  NOR2_X1 U14923 ( .A1(n12307), .A2(n12306), .ZN(n12473) );
  XNOR2_X1 U14924 ( .A(n12473), .B(n12472), .ZN(n12308) );
  NAND2_X1 U14925 ( .A1(n12308), .A2(n13243), .ZN(n12315) );
  OAI22_X1 U14926 ( .A1(n13249), .A2(n12310), .B1(n12309), .B2(n13271), .ZN(
        n12311) );
  AOI211_X1 U14927 ( .C1(n12313), .C2(n13261), .A(n12312), .B(n12311), .ZN(
        n12314) );
  OAI211_X1 U14928 ( .C1(n12316), .C2(n13226), .A(n12315), .B(n12314), .ZN(
        P3_U3153) );
  INV_X1 U14929 ( .A(n12317), .ZN(n12322) );
  AOI21_X1 U14930 ( .B1(P2_DATAO_REG_23__SCAN_IN), .B2(n15691), .A(n12318), 
        .ZN(n12319) );
  OAI21_X1 U14931 ( .B1(n12322), .B2(n15703), .A(n12319), .ZN(P1_U3332) );
  NOR2_X1 U14932 ( .A1(n12320), .A2(P2_U3088), .ZN(n14382) );
  AOI21_X1 U14933 ( .B1(P1_DATAO_REG_23__SCAN_IN), .B2(n14897), .A(n14382), 
        .ZN(n12321) );
  OAI21_X1 U14934 ( .B1(n12322), .B2(n14903), .A(n12321), .ZN(P2_U3304) );
  NOR2_X1 U14935 ( .A1(n12326), .A2(n12325), .ZN(n12323) );
  NAND2_X1 U14936 ( .A1(n12326), .A2(n12325), .ZN(n12327) );
  INV_X1 U14937 ( .A(P3_ADDR_REG_11__SCAN_IN), .ZN(n12330) );
  NAND2_X1 U14938 ( .A1(n12330), .A2(P1_ADDR_REG_11__SCAN_IN), .ZN(n12528) );
  NAND2_X1 U14939 ( .A1(n11368), .A2(P3_ADDR_REG_11__SCAN_IN), .ZN(n12331) );
  AND2_X1 U14940 ( .A1(n12528), .A2(n12331), .ZN(n12526) );
  XNOR2_X1 U14941 ( .A(n12527), .B(n12526), .ZN(n12332) );
  OAI21_X1 U14942 ( .B1(n12334), .B2(n6601), .A(P2_ADDR_REG_11__SCAN_IN), .ZN(
        n12335) );
  OAI21_X1 U14943 ( .B1(n6721), .B2(n6601), .A(n12335), .ZN(SUB_1596_U69) );
  XNOR2_X1 U14944 ( .A(n12336), .B(n7206), .ZN(n15873) );
  XNOR2_X1 U14945 ( .A(n12338), .B(n12337), .ZN(n12339) );
  AOI222_X1 U14946 ( .A1(n15611), .A2(n12339), .B1(n15094), .B2(n15500), .C1(
        n15096), .C2(n15521), .ZN(n15872) );
  MUX2_X1 U14947 ( .A(n11102), .B(n15872), .S(n15528), .Z(n12345) );
  AOI21_X1 U14948 ( .B1(n15785), .B2(n15869), .A(n15608), .ZN(n12341) );
  AND2_X1 U14949 ( .A1(n12342), .A2(n12341), .ZN(n15868) );
  OAI22_X1 U14950 ( .A1(n15807), .A2(n12207), .B1(n15804), .B2(n12414), .ZN(
        n12343) );
  AOI21_X1 U14951 ( .B1(n15868), .B2(n15812), .A(n12343), .ZN(n12344) );
  OAI211_X1 U14952 ( .C1(n15535), .C2(n15873), .A(n12345), .B(n12344), .ZN(
        P1_U3285) );
  INV_X1 U14953 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n12346) );
  OAI22_X1 U14954 ( .A1(n6548), .A2(n11157), .B1(n12346), .B2(n14736), .ZN(
        n12348) );
  NOR2_X1 U14955 ( .A1(n14698), .A2(n7166), .ZN(n12347) );
  AOI211_X1 U14956 ( .C1(n12349), .C2(n14703), .A(n12348), .B(n12347), .ZN(
        n12352) );
  NAND2_X1 U14957 ( .A1(n14723), .A2(n12350), .ZN(n12351) );
  OAI211_X1 U14958 ( .C1(n14719), .C2(n12353), .A(n12352), .B(n12351), .ZN(
        P2_U3263) );
  INV_X1 U14959 ( .A(n12354), .ZN(n12355) );
  OAI222_X1 U14960 ( .A1(n14914), .A2(n12356), .B1(P2_U3088), .B2(n14379), 
        .C1(n14903), .C2(n12355), .ZN(P2_U3305) );
  XNOR2_X1 U14961 ( .A(n12559), .B(n12363), .ZN(n12420) );
  NAND2_X1 U14962 ( .A1(n15662), .A2(n12413), .ZN(n12361) );
  INV_X1 U14963 ( .A(n12557), .ZN(n12364) );
  OAI21_X1 U14964 ( .B1(n12364), .B2(n12363), .A(n15611), .ZN(n12365) );
  NOR2_X1 U14965 ( .A1(n12557), .A2(n12558), .ZN(n12717) );
  NAND2_X1 U14966 ( .A1(n15094), .A2(n15521), .ZN(n12745) );
  OAI21_X1 U14967 ( .B1(n12365), .B2(n12717), .A(n12745), .ZN(n12422) );
  NAND2_X1 U14968 ( .A1(n12422), .A2(n15528), .ZN(n12373) );
  OAI22_X1 U14969 ( .A1(n15528), .A2(n12366), .B1(n12743), .B2(n15804), .ZN(
        n12371) );
  INV_X1 U14970 ( .A(n12560), .ZN(n12368) );
  OAI211_X1 U14971 ( .C1(n12367), .C2(n12368), .A(n12723), .B(n7132), .ZN(
        n12369) );
  NAND2_X1 U14972 ( .A1(n15092), .A2(n15500), .ZN(n12744) );
  AND2_X1 U14973 ( .A1(n12369), .A2(n12744), .ZN(n12419) );
  NOR2_X1 U14974 ( .A1(n12419), .A2(n15344), .ZN(n12370) );
  AOI211_X1 U14975 ( .C1(n15496), .C2(n12560), .A(n12371), .B(n12370), .ZN(
        n12372) );
  OAI211_X1 U14976 ( .C1(n12420), .C2(n15535), .A(n12373), .B(n12372), .ZN(
        P1_U3283) );
  OR2_X1 U14977 ( .A1(n12374), .A2(n12379), .ZN(n12375) );
  NAND2_X1 U14978 ( .A1(n12376), .A2(n12375), .ZN(n12389) );
  NAND2_X1 U14979 ( .A1(n14412), .A2(n14086), .ZN(n12378) );
  NAND2_X1 U14980 ( .A1(n14414), .A2(n14376), .ZN(n12377) );
  AND2_X1 U14981 ( .A1(n12378), .A2(n12377), .ZN(n12431) );
  XNOR2_X1 U14982 ( .A(n12380), .B(n12379), .ZN(n12381) );
  NAND2_X1 U14983 ( .A1(n12381), .A2(n14675), .ZN(n12382) );
  OAI211_X1 U14984 ( .C1(n12389), .C2(n10420), .A(n12431), .B(n12382), .ZN(
        n12390) );
  MUX2_X1 U14985 ( .A(P2_REG2_REG_9__SCAN_IN), .B(n12390), .S(n6548), .Z(
        n12383) );
  INV_X1 U14986 ( .A(n12383), .ZN(n12388) );
  AOI211_X1 U14987 ( .C1(n14159), .C2(n12384), .A(n14717), .B(n12464), .ZN(
        n12391) );
  INV_X1 U14988 ( .A(n14159), .ZN(n12436) );
  INV_X1 U14989 ( .A(n12433), .ZN(n12385) );
  OAI22_X1 U14990 ( .A1(n14698), .A2(n12436), .B1(n14736), .B2(n12385), .ZN(
        n12386) );
  AOI21_X1 U14991 ( .B1(n12391), .B2(n14703), .A(n12386), .ZN(n12387) );
  OAI211_X1 U14992 ( .C1(n12389), .C2(n14682), .A(n12388), .B(n12387), .ZN(
        P2_U3256) );
  INV_X1 U14993 ( .A(n12389), .ZN(n12392) );
  INV_X1 U14994 ( .A(n14846), .ZN(n14837) );
  AOI211_X1 U14995 ( .C1(n12392), .C2(n14837), .A(n12391), .B(n12390), .ZN(
        n12399) );
  INV_X1 U14996 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n12393) );
  OAI22_X1 U14997 ( .A1(n14840), .A2(n12436), .B1(n16011), .B2(n12393), .ZN(
        n12394) );
  INV_X1 U14998 ( .A(n12394), .ZN(n12395) );
  OAI21_X1 U14999 ( .B1(n12399), .B2(n16008), .A(n12395), .ZN(P2_U3508) );
  OAI22_X1 U15000 ( .A1(n14892), .A2(n12436), .B1(n16004), .B2(n12396), .ZN(
        n12397) );
  INV_X1 U15001 ( .A(n12397), .ZN(n12398) );
  OAI21_X1 U15002 ( .B1(n12399), .B2(n16002), .A(n12398), .ZN(P2_U3457) );
  INV_X1 U15003 ( .A(n12400), .ZN(n12401) );
  OR2_X1 U15004 ( .A1(n12400), .A2(n13390), .ZN(n12449) );
  OAI21_X1 U15005 ( .B1(n12401), .B2(n7550), .A(n12449), .ZN(n12402) );
  AOI222_X1 U15006 ( .A1(n12402), .A2(n16044), .B1(n13503), .B2(n16049), .C1(
        n13501), .C2(n16046), .ZN(n12444) );
  OAI21_X1 U15007 ( .B1(n12404), .B2(n13390), .A(n12403), .ZN(n12443) );
  INV_X1 U15008 ( .A(n13955), .ZN(n13943) );
  NAND2_X1 U15009 ( .A1(n12443), .A2(n13943), .ZN(n12406) );
  INV_X1 U15010 ( .A(n12859), .ZN(n12438) );
  AOI22_X1 U15011 ( .A1(n13953), .A2(n12438), .B1(P3_REG0_REG_11__SCAN_IN), 
        .B2(n16092), .ZN(n12405) );
  OAI211_X1 U15012 ( .C1(n16092), .C2(n12444), .A(n12406), .B(n12405), .ZN(
        P3_U3423) );
  INV_X1 U15013 ( .A(n12407), .ZN(n12408) );
  AOI21_X1 U15014 ( .B1(n12410), .B2(n7200), .A(n12408), .ZN(n12418) );
  NAND2_X1 U15015 ( .A1(n15062), .A2(n15096), .ZN(n12412) );
  OAI211_X1 U15016 ( .C1(n12413), .C2(n15065), .A(n12412), .B(n12411), .ZN(
        n12416) );
  NOR2_X1 U15017 ( .A1(n15077), .A2(n12414), .ZN(n12415) );
  AOI211_X1 U15018 ( .C1(n15068), .C2(n15869), .A(n12416), .B(n12415), .ZN(
        n12417) );
  OAI21_X1 U15019 ( .B1(n12418), .B2(n15070), .A(n12417), .ZN(P1_U3221) );
  NAND2_X1 U15020 ( .A1(n12560), .A2(n15870), .ZN(n12750) );
  OAI211_X1 U15021 ( .C1(n12420), .C2(n15874), .A(n12419), .B(n12750), .ZN(
        n12421) );
  NOR2_X1 U15022 ( .A1(n12422), .A2(n12421), .ZN(n12425) );
  NAND2_X1 U15023 ( .A1(n15884), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n12423) );
  OAI21_X1 U15024 ( .B1(n12425), .B2(n15884), .A(n12423), .ZN(P1_U3538) );
  NAND2_X1 U15025 ( .A1(n15876), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n12424) );
  OAI21_X1 U15026 ( .B1(n12425), .B2(n15876), .A(n12424), .ZN(P1_U3489) );
  OAI21_X1 U15027 ( .B1(n12428), .B2(n12427), .A(n12426), .ZN(n12429) );
  NAND2_X1 U15028 ( .A1(n12429), .A2(n14065), .ZN(n12435) );
  OAI21_X1 U15029 ( .B1(n14090), .B2(n12431), .A(n12430), .ZN(n12432) );
  AOI21_X1 U15030 ( .B1(n12433), .B2(n14088), .A(n12432), .ZN(n12434) );
  OAI211_X1 U15031 ( .C1(n12436), .C2(n14073), .A(n12435), .B(n12434), .ZN(
        P2_U3203) );
  INV_X1 U15032 ( .A(n12443), .ZN(n12442) );
  INV_X1 U15033 ( .A(n12437), .ZN(n12864) );
  AOI22_X1 U15034 ( .A1(n13814), .A2(n12438), .B1(n16061), .B2(n12864), .ZN(
        n12441) );
  MUX2_X1 U15035 ( .A(n12439), .B(n12444), .S(n9401), .Z(n12440) );
  OAI211_X1 U15036 ( .C1(n12442), .C2(n13824), .A(n12441), .B(n12440), .ZN(
        P3_U3222) );
  INV_X1 U15037 ( .A(n13883), .ZN(n13875) );
  NAND2_X1 U15038 ( .A1(n12443), .A2(n13875), .ZN(n12446) );
  MUX2_X1 U15039 ( .A(n12593), .B(n12444), .S(n16106), .Z(n12445) );
  OAI211_X1 U15040 ( .C1(n13860), .C2(n12859), .A(n12446), .B(n12445), .ZN(
        P3_U3470) );
  XNOR2_X1 U15041 ( .A(n12447), .B(n13323), .ZN(n12739) );
  AOI22_X1 U15042 ( .A1(n13953), .A2(n12886), .B1(P3_REG0_REG_12__SCAN_IN), 
        .B2(n16092), .ZN(n12455) );
  NAND2_X1 U15043 ( .A1(n12449), .A2(n12448), .ZN(n12450) );
  XNOR2_X1 U15044 ( .A(n12450), .B(n13323), .ZN(n12451) );
  NAND2_X1 U15045 ( .A1(n12451), .A2(n16044), .ZN(n12453) );
  AOI22_X1 U15046 ( .A1(n16049), .A2(n13502), .B1(n13500), .B2(n16046), .ZN(
        n12452) );
  NAND2_X1 U15047 ( .A1(n12453), .A2(n12452), .ZN(n12736) );
  NAND2_X1 U15048 ( .A1(n12736), .A2(n16094), .ZN(n12454) );
  OAI211_X1 U15049 ( .C1(n12739), .C2(n13955), .A(n12455), .B(n12454), .ZN(
        P3_U3426) );
  XNOR2_X1 U15050 ( .A(n12456), .B(n14344), .ZN(n12463) );
  OR2_X1 U15051 ( .A1(n12457), .A2(n14344), .ZN(n12458) );
  NAND2_X1 U15052 ( .A1(n12459), .A2(n12458), .ZN(n14845) );
  NAND2_X1 U15053 ( .A1(n14413), .A2(n14376), .ZN(n12461) );
  NAND2_X1 U15054 ( .A1(n14411), .A2(n14086), .ZN(n12460) );
  AND2_X1 U15055 ( .A1(n12461), .A2(n12460), .ZN(n12818) );
  OAI21_X1 U15056 ( .B1(n14845), .B2(n10420), .A(n12818), .ZN(n12462) );
  AOI21_X1 U15057 ( .B1(n12463), .B2(n14675), .A(n12462), .ZN(n14844) );
  INV_X1 U15058 ( .A(n12464), .ZN(n12466) );
  AOI211_X1 U15059 ( .C1(n14842), .C2(n12466), .A(n14717), .B(n12465), .ZN(
        n14841) );
  AOI22_X1 U15060 ( .A1(n14738), .A2(P2_REG2_REG_10__SCAN_IN), .B1(n12815), 
        .B2(n14713), .ZN(n12467) );
  OAI21_X1 U15061 ( .B1(n12468), .B2(n14698), .A(n12467), .ZN(n12470) );
  NOR2_X1 U15062 ( .A1(n14845), .A2(n14682), .ZN(n12469) );
  AOI211_X1 U15063 ( .C1(n14841), .C2(n14703), .A(n12470), .B(n12469), .ZN(
        n12471) );
  OAI21_X1 U15064 ( .B1(n14738), .B2(n14844), .A(n12471), .ZN(P2_U3255) );
  MUX2_X1 U15065 ( .A(n12477), .B(n12473), .S(n12472), .Z(n12474) );
  XNOR2_X1 U15066 ( .A(n12474), .B(n6630), .ZN(n12475) );
  NAND2_X1 U15067 ( .A1(n12475), .A2(n13243), .ZN(n12482) );
  INV_X1 U15068 ( .A(n13504), .ZN(n12476) );
  OAI22_X1 U15069 ( .A1(n13249), .A2(n12477), .B1(n12476), .B2(n13271), .ZN(
        n12478) );
  AOI211_X1 U15070 ( .C1(n12480), .C2(n13261), .A(n12479), .B(n12478), .ZN(
        n12481) );
  OAI211_X1 U15071 ( .C1(n12483), .C2(n13226), .A(n12482), .B(n12481), .ZN(
        P3_U3161) );
  XNOR2_X1 U15072 ( .A(n12735), .B(n11436), .ZN(n12853) );
  XNOR2_X1 U15073 ( .A(n12853), .B(n13503), .ZN(n12488) );
  NOR2_X1 U15074 ( .A1(n12484), .A2(n13504), .ZN(n12485) );
  OR2_X1 U15075 ( .A1(n12486), .A2(n12485), .ZN(n12487) );
  AOI211_X1 U15076 ( .C1(n12488), .C2(n12487), .A(n13264), .B(n6717), .ZN(
        n12496) );
  INV_X1 U15077 ( .A(n12489), .ZN(n12625) );
  NAND2_X1 U15078 ( .A1(n13273), .A2(n12625), .ZN(n12494) );
  AOI21_X1 U15079 ( .B1(n13269), .B2(n13504), .A(n12490), .ZN(n12493) );
  INV_X1 U15080 ( .A(n12735), .ZN(n12626) );
  NAND2_X1 U15081 ( .A1(n13261), .A2(n12626), .ZN(n12492) );
  NAND2_X1 U15082 ( .A1(n13247), .A2(n13502), .ZN(n12491) );
  NAND4_X1 U15083 ( .A1(n12494), .A2(n12493), .A3(n12492), .A4(n12491), .ZN(
        n12495) );
  OR2_X1 U15084 ( .A1(n12496), .A2(n12495), .ZN(P3_U3157) );
  XNOR2_X1 U15085 ( .A(n12497), .B(n7844), .ZN(n12630) );
  INV_X1 U15086 ( .A(n12630), .ZN(n12504) );
  AOI22_X1 U15087 ( .A1(n16046), .A2(n13502), .B1(n13504), .B2(n16049), .ZN(
        n12502) );
  OAI211_X1 U15088 ( .C1(n12500), .C2(n12499), .A(n12498), .B(n16044), .ZN(
        n12501) );
  OAI211_X1 U15089 ( .C1(n12630), .C2(n12503), .A(n12502), .B(n12501), .ZN(
        n12622) );
  AOI21_X1 U15090 ( .B1(n16090), .B2(n12504), .A(n12622), .ZN(n12732) );
  AOI22_X1 U15091 ( .A1(n13953), .A2(n12626), .B1(P3_REG0_REG_10__SCAN_IN), 
        .B2(n16092), .ZN(n12505) );
  OAI21_X1 U15092 ( .B1(n12732), .B2(n16092), .A(n12505), .ZN(P3_U3420) );
  INV_X1 U15093 ( .A(n12506), .ZN(n12508) );
  OAI222_X1 U15094 ( .A1(n12509), .A2(P3_U3151), .B1(n13102), .B2(n12508), 
        .C1(n12507), .C2(n13970), .ZN(P3_U3269) );
  OAI211_X1 U15095 ( .C1(n12512), .C2(n12511), .A(n12510), .B(n15072), .ZN(
        n12518) );
  AOI22_X1 U15096 ( .A1(n15080), .A2(n12513), .B1(P1_REG3_REG_9__SCAN_IN), 
        .B2(P1_U3086), .ZN(n12514) );
  OAI21_X1 U15097 ( .B1(n15077), .B2(n12515), .A(n12514), .ZN(n12516) );
  AOI21_X1 U15098 ( .B1(n15068), .B2(n15662), .A(n12516), .ZN(n12517) );
  NAND2_X1 U15099 ( .A1(n12518), .A2(n12517), .ZN(P1_U3231) );
  MUX2_X1 U15100 ( .A(n12519), .B(P2_REG2_REG_1__SCAN_IN), .S(n14719), .Z(
        n12523) );
  AOI22_X1 U15101 ( .A1(n14739), .A2(n14114), .B1(P2_REG3_REG_1__SCAN_IN), 
        .B2(n14713), .ZN(n12520) );
  OAI21_X1 U15102 ( .B1(n14721), .B2(n12521), .A(n12520), .ZN(n12522) );
  AOI211_X1 U15103 ( .C1(n14723), .C2(n12524), .A(n12523), .B(n12522), .ZN(
        n12525) );
  INV_X1 U15104 ( .A(n12525), .ZN(P2_U3264) );
  NAND2_X1 U15105 ( .A1(n12527), .A2(n12526), .ZN(n12529) );
  NAND2_X1 U15106 ( .A1(n12529), .A2(n12528), .ZN(n12845) );
  INV_X1 U15107 ( .A(n12845), .ZN(n12531) );
  XNOR2_X1 U15108 ( .A(n13517), .B(P1_ADDR_REG_12__SCAN_IN), .ZN(n12844) );
  INV_X1 U15109 ( .A(n12844), .ZN(n12530) );
  XNOR2_X1 U15110 ( .A(n12531), .B(n12530), .ZN(n12842) );
  XNOR2_X1 U15111 ( .A(n12842), .B(P2_ADDR_REG_12__SCAN_IN), .ZN(n12532) );
  XNOR2_X1 U15112 ( .A(n12843), .B(n12532), .ZN(SUB_1596_U68) );
  INV_X1 U15113 ( .A(n12533), .ZN(n12536) );
  AOI22_X1 U15114 ( .A1(n14739), .A2(n14136), .B1(n14713), .B2(n12534), .ZN(
        n12535) );
  OAI21_X1 U15115 ( .B1(n12536), .B2(n14721), .A(n12535), .ZN(n12539) );
  MUX2_X1 U15116 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n12537), .S(n6548), .Z(
        n12538) );
  AOI211_X1 U15117 ( .C1(n14723), .C2(n12540), .A(n12539), .B(n12538), .ZN(
        n12541) );
  INV_X1 U15118 ( .A(n12541), .ZN(P2_U3261) );
  OAI22_X1 U15119 ( .A1(n6548), .A2(n11159), .B1(P2_REG3_REG_3__SCAN_IN), .B2(
        n14736), .ZN(n12542) );
  AOI21_X1 U15120 ( .B1(n14739), .B2(n14129), .A(n12542), .ZN(n12543) );
  OAI21_X1 U15121 ( .B1(n14721), .B2(n12544), .A(n12543), .ZN(n12545) );
  AOI21_X1 U15122 ( .B1(n14723), .B2(n12546), .A(n12545), .ZN(n12547) );
  OAI21_X1 U15123 ( .B1(n14719), .B2(n12548), .A(n12547), .ZN(P2_U3262) );
  INV_X1 U15124 ( .A(n15428), .ZN(n15480) );
  AND2_X1 U15125 ( .A1(n12902), .A2(n12552), .ZN(n12551) );
  INV_X1 U15126 ( .A(n12549), .ZN(n12550) );
  INV_X1 U15127 ( .A(n12902), .ZN(n12726) );
  NAND2_X1 U15128 ( .A1(n12553), .A2(n12552), .ZN(n12554) );
  INV_X1 U15129 ( .A(n12553), .ZN(n12716) );
  XNOR2_X1 U15130 ( .A(n13024), .B(n13023), .ZN(n15655) );
  NAND2_X1 U15131 ( .A1(n12559), .A2(n12558), .ZN(n12562) );
  OR2_X1 U15132 ( .A1(n12560), .A2(n15093), .ZN(n12561) );
  NOR2_X1 U15133 ( .A1(n12902), .A2(n15092), .ZN(n12564) );
  NAND2_X1 U15134 ( .A1(n12902), .A2(n15092), .ZN(n12563) );
  OAI21_X1 U15135 ( .B1(n12566), .B2(n7175), .A(n13000), .ZN(n15652) );
  INV_X1 U15136 ( .A(n15651), .ZN(n14978) );
  INV_X1 U15137 ( .A(n12567), .ZN(n12724) );
  AOI211_X1 U15138 ( .C1(n15651), .C2(n12724), .A(n15608), .B(n15526), .ZN(
        n15649) );
  NAND2_X1 U15139 ( .A1(n15649), .A2(n15812), .ZN(n12574) );
  NAND2_X1 U15140 ( .A1(n15092), .A2(n15521), .ZN(n12570) );
  NAND2_X1 U15141 ( .A1(n15502), .A2(n15500), .ZN(n12569) );
  NAND2_X1 U15142 ( .A1(n12570), .A2(n12569), .ZN(n15650) );
  INV_X1 U15143 ( .A(n15650), .ZN(n12571) );
  OAI22_X1 U15144 ( .A1(n6556), .A2(n12571), .B1(n14973), .B2(n15804), .ZN(
        n12572) );
  AOI21_X1 U15145 ( .B1(P1_REG2_REG_12__SCAN_IN), .B2(n6556), .A(n12572), .ZN(
        n12573) );
  OAI211_X1 U15146 ( .C1(n14978), .C2(n15807), .A(n12574), .B(n12573), .ZN(
        n12575) );
  AOI21_X1 U15147 ( .B1(n15652), .B2(n15513), .A(n12575), .ZN(n12576) );
  OAI21_X1 U15148 ( .B1(n15480), .B2(n15655), .A(n12576), .ZN(P1_U3281) );
  INV_X1 U15149 ( .A(n12577), .ZN(n12581) );
  OAI222_X1 U15150 ( .A1(n12579), .A2(P1_U3086), .B1(n15703), .B2(n12581), 
        .C1(n12578), .C2(n13134), .ZN(P1_U3331) );
  OAI222_X1 U15151 ( .A1(P2_U3088), .A2(n12582), .B1(n14903), .B2(n12581), 
        .C1(n12580), .C2(n14914), .ZN(P2_U3303) );
  AOI22_X1 U15152 ( .A1(n14739), .A2(n14154), .B1(n14713), .B2(n12583), .ZN(
        n12584) );
  OAI21_X1 U15153 ( .B1(n12585), .B2(n14721), .A(n12584), .ZN(n12588) );
  MUX2_X1 U15154 ( .A(P2_REG2_REG_8__SCAN_IN), .B(n12586), .S(n6548), .Z(
        n12587) );
  AOI211_X1 U15155 ( .C1(n12589), .C2(n14723), .A(n12588), .B(n12587), .ZN(
        n12590) );
  INV_X1 U15156 ( .A(n12590), .ZN(P2_U3257) );
  INV_X1 U15157 ( .A(n13525), .ZN(n12591) );
  AOI21_X1 U15158 ( .B1(n12593), .B2(n12592), .A(n12591), .ZN(n12606) );
  OAI21_X1 U15159 ( .B1(P3_REG2_REG_11__SCAN_IN), .B2(n12595), .A(n12594), 
        .ZN(n12596) );
  NAND2_X1 U15160 ( .A1(n12596), .A2(n13583), .ZN(n12605) );
  OAI21_X1 U15161 ( .B1(n12599), .B2(n12598), .A(n12597), .ZN(n12603) );
  NAND2_X1 U15162 ( .A1(P3_U3151), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n12860)
         );
  NAND2_X1 U15163 ( .A1(n16012), .A2(P3_ADDR_REG_11__SCAN_IN), .ZN(n12600) );
  OAI211_X1 U15164 ( .C1(n13617), .C2(n12601), .A(n12860), .B(n12600), .ZN(
        n12602) );
  AOI21_X1 U15165 ( .B1(n12603), .B2(n13537), .A(n12602), .ZN(n12604) );
  OAI211_X1 U15166 ( .C1(n12606), .C2(n16015), .A(n12605), .B(n12604), .ZN(
        P3_U3193) );
  NOR2_X1 U15167 ( .A1(n12607), .A2(n8585), .ZN(n12609) );
  OAI22_X1 U15168 ( .A1(n12609), .A2(n14417), .B1(n12608), .B2(n15983), .ZN(
        n12610) );
  XNOR2_X1 U15169 ( .A(n12610), .B(n14335), .ZN(n15992) );
  OAI211_X1 U15170 ( .C1(n7900), .C2(n6730), .A(n6604), .B(n14818), .ZN(n15988) );
  AOI22_X1 U15171 ( .A1(n14739), .A2(n14148), .B1(n14713), .B2(n12611), .ZN(
        n12612) );
  OAI21_X1 U15172 ( .B1(n15988), .B2(n14721), .A(n12612), .ZN(n12620) );
  OAI21_X1 U15173 ( .B1(n12615), .B2(n12614), .A(n12613), .ZN(n12616) );
  XOR2_X1 U15174 ( .A(n14335), .B(n12616), .Z(n12618) );
  OAI21_X1 U15175 ( .B1(n12618), .B2(n8640), .A(n12617), .ZN(n15990) );
  MUX2_X1 U15176 ( .A(P2_REG2_REG_6__SCAN_IN), .B(n15990), .S(n6548), .Z(
        n12619) );
  AOI211_X1 U15177 ( .C1(n14723), .C2(n15992), .A(n12620), .B(n12619), .ZN(
        n12621) );
  INV_X1 U15178 ( .A(n12621), .ZN(P2_U3259) );
  INV_X1 U15179 ( .A(n12622), .ZN(n12623) );
  MUX2_X1 U15180 ( .A(n12624), .B(n12623), .S(n9401), .Z(n12628) );
  AOI22_X1 U15181 ( .A1(n13814), .A2(n12626), .B1(n16061), .B2(n12625), .ZN(
        n12627) );
  OAI211_X1 U15182 ( .C1(n12630), .C2(n12629), .A(n12628), .B(n12627), .ZN(
        P3_U3223) );
  XNOR2_X1 U15183 ( .A(n15205), .B(P1_REG1_REG_16__SCAN_IN), .ZN(n12638) );
  NAND2_X1 U15184 ( .A1(n12634), .A2(n12633), .ZN(n12635) );
  INV_X1 U15185 ( .A(n15199), .ZN(n12636) );
  AOI211_X1 U15186 ( .C1(n12638), .C2(n12637), .A(n15248), .B(n12636), .ZN(
        n12656) );
  INV_X1 U15187 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n12639) );
  OR2_X1 U15188 ( .A1(n15205), .A2(n12639), .ZN(n12641) );
  NAND2_X1 U15189 ( .A1(n15205), .A2(n12639), .ZN(n12640) );
  AND2_X1 U15190 ( .A1(n12641), .A2(n12640), .ZN(n12650) );
  NAND2_X1 U15191 ( .A1(n12643), .A2(n12642), .ZN(n12647) );
  OR2_X1 U15192 ( .A1(n12645), .A2(n12644), .ZN(n12646) );
  NAND2_X1 U15193 ( .A1(n12647), .A2(n12646), .ZN(n12649) );
  INV_X1 U15194 ( .A(n15207), .ZN(n12648) );
  AOI211_X1 U15195 ( .C1(n12650), .C2(n12649), .A(n15242), .B(n12648), .ZN(
        n12655) );
  INV_X1 U15196 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n15745) );
  NAND2_X1 U15197 ( .A1(n15223), .A2(n15205), .ZN(n12653) );
  NOR2_X1 U15198 ( .A1(n12651), .A2(P1_STATE_REG_SCAN_IN), .ZN(n14994) );
  INV_X1 U15199 ( .A(n14994), .ZN(n12652) );
  OAI211_X1 U15200 ( .C1(n15745), .C2(n15252), .A(n12653), .B(n12652), .ZN(
        n12654) );
  OR3_X1 U15201 ( .A1(n12656), .A2(n12655), .A3(n12654), .ZN(P1_U3259) );
  XNOR2_X1 U15202 ( .A(n14171), .B(n14411), .ZN(n14345) );
  XOR2_X1 U15203 ( .A(n12657), .B(n14345), .Z(n14833) );
  AND2_X1 U15204 ( .A1(n12659), .A2(n12658), .ZN(n12660) );
  NAND2_X1 U15205 ( .A1(n12660), .A2(n14345), .ZN(n12827) );
  OAI21_X1 U15206 ( .B1(n12660), .B2(n14345), .A(n12827), .ZN(n12662) );
  INV_X1 U15207 ( .A(n14410), .ZN(n14174) );
  OAI22_X1 U15208 ( .A1(n12661), .A2(n14095), .B1(n14174), .B2(n14096), .ZN(
        n12872) );
  AOI21_X1 U15209 ( .B1(n12662), .B2(n14675), .A(n12872), .ZN(n12663) );
  OAI21_X1 U15210 ( .B1(n14833), .B2(n10420), .A(n12663), .ZN(n14834) );
  NAND2_X1 U15211 ( .A1(n14834), .A2(n6548), .ZN(n12668) );
  INV_X1 U15212 ( .A(n12465), .ZN(n12664) );
  AOI211_X1 U15213 ( .C1(n14171), .C2(n12664), .A(n14717), .B(n7224), .ZN(
        n14835) );
  AOI22_X1 U15214 ( .A1(n14719), .A2(P2_REG2_REG_11__SCAN_IN), .B1(n12871), 
        .B2(n14713), .ZN(n12665) );
  OAI21_X1 U15215 ( .B1(n14893), .B2(n14698), .A(n12665), .ZN(n12666) );
  AOI21_X1 U15216 ( .B1(n14835), .B2(n14703), .A(n12666), .ZN(n12667) );
  OAI211_X1 U15217 ( .C1(n14833), .C2(n14682), .A(n12668), .B(n12667), .ZN(
        P2_U3254) );
  NAND2_X1 U15218 ( .A1(P2_U3088), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n14041)
         );
  OAI21_X1 U15219 ( .B1(n15919), .B2(n12685), .A(n14041), .ZN(n12677) );
  NAND2_X1 U15220 ( .A1(n12669), .A2(n12679), .ZN(n12670) );
  NAND2_X1 U15221 ( .A1(n12671), .A2(n12670), .ZN(n15931) );
  XNOR2_X1 U15222 ( .A(n15935), .B(n14815), .ZN(n15930) );
  NAND2_X1 U15223 ( .A1(n15931), .A2(n15930), .ZN(n15929) );
  NAND2_X1 U15224 ( .A1(n15935), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n12672) );
  NAND2_X1 U15225 ( .A1(n15929), .A2(n12672), .ZN(n12674) );
  INV_X1 U15226 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n14807) );
  XNOR2_X1 U15227 ( .A(n12803), .B(n14807), .ZN(n12673) );
  NAND2_X1 U15228 ( .A1(n12674), .A2(n12673), .ZN(n12805) );
  OAI211_X1 U15229 ( .C1(n12674), .C2(n12673), .A(n12805), .B(n15928), .ZN(
        n12675) );
  INV_X1 U15230 ( .A(n12675), .ZN(n12676) );
  AOI211_X1 U15231 ( .C1(n15899), .C2(P2_ADDR_REG_17__SCAN_IN), .A(n12677), 
        .B(n12676), .ZN(n12692) );
  NAND2_X1 U15232 ( .A1(n12678), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n12682) );
  NAND2_X1 U15233 ( .A1(n12680), .A2(n12679), .ZN(n12681) );
  NAND2_X1 U15234 ( .A1(n12682), .A2(n12681), .ZN(n15940) );
  OR2_X1 U15235 ( .A1(n15935), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n12683) );
  NAND2_X1 U15236 ( .A1(n15935), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n12686) );
  AND2_X1 U15237 ( .A1(n12683), .A2(n12686), .ZN(n15939) );
  INV_X1 U15238 ( .A(n15938), .ZN(n12690) );
  NAND2_X1 U15239 ( .A1(n12685), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n12684) );
  OAI211_X1 U15240 ( .C1(P2_REG2_REG_17__SCAN_IN), .C2(n12685), .A(n12686), 
        .B(n12684), .ZN(n12689) );
  NAND2_X1 U15241 ( .A1(n12803), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n12795) );
  OAI21_X1 U15242 ( .B1(n12803), .B2(P2_REG2_REG_17__SCAN_IN), .A(n12795), 
        .ZN(n12687) );
  INV_X1 U15243 ( .A(n12687), .ZN(n12688) );
  OAI211_X1 U15244 ( .C1(n12690), .C2(n12689), .A(n12796), .B(n15937), .ZN(
        n12691) );
  NAND2_X1 U15245 ( .A1(n12692), .A2(n12691), .ZN(P2_U3231) );
  INV_X1 U15246 ( .A(n12883), .ZN(n12693) );
  AOI22_X1 U15247 ( .A1(n13814), .A2(n12886), .B1(n16061), .B2(n12693), .ZN(
        n12697) );
  INV_X1 U15248 ( .A(n12736), .ZN(n12695) );
  MUX2_X1 U15249 ( .A(n12695), .B(n12694), .S(n16066), .Z(n12696) );
  OAI211_X1 U15250 ( .C1(n12739), .C2(n13824), .A(n12697), .B(n12696), .ZN(
        P3_U3221) );
  INV_X1 U15251 ( .A(n12700), .ZN(n13398) );
  XNOR2_X1 U15252 ( .A(n12698), .B(n13398), .ZN(n12715) );
  OAI211_X1 U15253 ( .C1(n12701), .C2(n12700), .A(n12699), .B(n16044), .ZN(
        n12703) );
  OR2_X1 U15254 ( .A1(n12934), .A2(n13815), .ZN(n12702) );
  OAI211_X1 U15255 ( .C1(n13816), .C2(n13817), .A(n12703), .B(n12702), .ZN(
        n12713) );
  OAI22_X1 U15256 ( .A1(n13223), .A2(n13918), .B1(n12704), .B2(n16094), .ZN(
        n12705) );
  AOI21_X1 U15257 ( .B1(n12713), .B2(n16094), .A(n12705), .ZN(n12706) );
  OAI21_X1 U15258 ( .B1(n12715), .B2(n13955), .A(n12706), .ZN(P3_U3429) );
  NOR2_X1 U15259 ( .A1(n13223), .A2(n13737), .ZN(n12709) );
  OAI22_X1 U15260 ( .A1(n9401), .A2(n13532), .B1(n13227), .B2(n12707), .ZN(
        n12708) );
  AOI211_X1 U15261 ( .C1(n12713), .C2(n9401), .A(n12709), .B(n12708), .ZN(
        n12710) );
  OAI21_X1 U15262 ( .B1(n12715), .B2(n13824), .A(n12710), .ZN(P3_U3220) );
  OAI22_X1 U15263 ( .A1(n13223), .A2(n13860), .B1(n16106), .B2(n12711), .ZN(
        n12712) );
  AOI21_X1 U15264 ( .B1(n12713), .B2(n16106), .A(n12712), .ZN(n12714) );
  OAI21_X1 U15265 ( .B1(n12715), .B2(n13883), .A(n12714), .ZN(P3_U3472) );
  NOR2_X1 U15266 ( .A1(n12717), .A2(n12716), .ZN(n12718) );
  XNOR2_X1 U15267 ( .A(n12718), .B(n12720), .ZN(n12719) );
  AOI222_X1 U15268 ( .A1(n15611), .A2(n12719), .B1(n15520), .B2(n15500), .C1(
        n15093), .C2(n15521), .ZN(n15660) );
  INV_X1 U15269 ( .A(n12720), .ZN(n12721) );
  XNOR2_X1 U15270 ( .A(n12722), .B(n12721), .ZN(n15656) );
  INV_X1 U15271 ( .A(n12723), .ZN(n12725) );
  OAI211_X1 U15272 ( .C1(n12726), .C2(n12725), .A(n12724), .B(n7132), .ZN(
        n15659) );
  OAI22_X1 U15273 ( .A1(n15528), .A2(n12727), .B1(n12907), .B2(n15804), .ZN(
        n12728) );
  AOI21_X1 U15274 ( .B1(n15496), .B2(n12902), .A(n12728), .ZN(n12729) );
  OAI21_X1 U15275 ( .B1(n15659), .B2(n15344), .A(n12729), .ZN(n12730) );
  AOI21_X1 U15276 ( .B1(n15656), .B2(n15513), .A(n12730), .ZN(n12731) );
  OAI21_X1 U15277 ( .B1(n15660), .B2(n6556), .A(n12731), .ZN(P1_U3282) );
  MUX2_X1 U15278 ( .A(n12733), .B(n12732), .S(n16106), .Z(n12734) );
  OAI21_X1 U15279 ( .B1(n13860), .B2(n12735), .A(n12734), .ZN(P3_U3469) );
  MUX2_X1 U15280 ( .A(n12736), .B(P3_REG1_REG_12__SCAN_IN), .S(n16103), .Z(
        n12737) );
  AOI21_X1 U15281 ( .B1(n13880), .B2(n12886), .A(n12737), .ZN(n12738) );
  OAI21_X1 U15282 ( .B1(n12739), .B2(n13883), .A(n12738), .ZN(P3_U3471) );
  OAI211_X1 U15283 ( .C1(n12742), .C2(n12741), .A(n12740), .B(n15072), .ZN(
        n12749) );
  INV_X1 U15284 ( .A(n12743), .ZN(n12747) );
  AND2_X1 U15285 ( .A1(P1_U3086), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n15177) );
  AOI21_X1 U15286 ( .B1(n12745), .B2(n12744), .A(n15025), .ZN(n12746) );
  AOI211_X1 U15287 ( .C1(n12747), .C2(n15061), .A(n15177), .B(n12746), .ZN(
        n12748) );
  OAI211_X1 U15288 ( .C1(n12751), .C2(n12750), .A(n12749), .B(n12748), .ZN(
        P1_U3217) );
  XNOR2_X1 U15289 ( .A(n12752), .B(n14350), .ZN(n12783) );
  INV_X1 U15290 ( .A(n12783), .ZN(n12764) );
  INV_X1 U15291 ( .A(n14350), .ZN(n12753) );
  XNOR2_X1 U15292 ( .A(n12754), .B(n12753), .ZN(n12755) );
  NAND2_X1 U15293 ( .A1(n12755), .A2(n14675), .ZN(n12758) );
  NAND2_X1 U15294 ( .A1(n14408), .A2(n14086), .ZN(n12757) );
  NAND2_X1 U15295 ( .A1(n14410), .A2(n14376), .ZN(n12756) );
  AND2_X1 U15296 ( .A1(n12757), .A2(n12756), .ZN(n12926) );
  NAND2_X1 U15297 ( .A1(n12758), .A2(n12926), .ZN(n12782) );
  INV_X1 U15298 ( .A(n12917), .ZN(n12759) );
  AOI211_X1 U15299 ( .C1(n14191), .C2(n12834), .A(n14717), .B(n12759), .ZN(
        n12781) );
  NAND2_X1 U15300 ( .A1(n12781), .A2(n14703), .ZN(n12761) );
  AOI22_X1 U15301 ( .A1(n14719), .A2(P2_REG2_REG_13__SCAN_IN), .B1(n12929), 
        .B2(n14713), .ZN(n12760) );
  OAI211_X1 U15302 ( .C1(n6951), .C2(n14698), .A(n12761), .B(n12760), .ZN(
        n12762) );
  AOI21_X1 U15303 ( .B1(n6548), .B2(n12782), .A(n12762), .ZN(n12763) );
  OAI21_X1 U15304 ( .B1(n14742), .B2(n12764), .A(n12763), .ZN(P2_U3252) );
  XNOR2_X1 U15305 ( .A(n12765), .B(n13402), .ZN(n12780) );
  OAI211_X1 U15306 ( .C1(n12767), .C2(n13402), .A(n12766), .B(n16044), .ZN(
        n12769) );
  AOI22_X1 U15307 ( .A1(n16046), .A2(n13498), .B1(n13500), .B2(n16049), .ZN(
        n12768) );
  NAND2_X1 U15308 ( .A1(n12769), .A2(n12768), .ZN(n12777) );
  OAI22_X1 U15309 ( .A1(n13404), .A2(n13918), .B1(n12770), .B2(n16094), .ZN(
        n12771) );
  AOI21_X1 U15310 ( .B1(n12777), .B2(n16094), .A(n12771), .ZN(n12772) );
  OAI21_X1 U15311 ( .B1(n12780), .B2(n13955), .A(n12772), .ZN(P3_U3432) );
  AOI22_X1 U15312 ( .A1(n16066), .A2(P3_REG2_REG_14__SCAN_IN), .B1(n16061), 
        .B2(n13156), .ZN(n12773) );
  OAI21_X1 U15313 ( .B1(n13404), .B2(n13737), .A(n12773), .ZN(n12774) );
  AOI21_X1 U15314 ( .B1(n12777), .B2(n9401), .A(n12774), .ZN(n12775) );
  OAI21_X1 U15315 ( .B1(n12780), .B2(n13824), .A(n12775), .ZN(P3_U3219) );
  INV_X1 U15316 ( .A(n13404), .ZN(n12776) );
  AOI22_X1 U15317 ( .A1(n12776), .A2(n13880), .B1(P3_REG1_REG_14__SCAN_IN), 
        .B2(n16103), .ZN(n12779) );
  NAND2_X1 U15318 ( .A1(n12777), .A2(n16106), .ZN(n12778) );
  OAI211_X1 U15319 ( .C1(n12780), .C2(n13883), .A(n12779), .B(n12778), .ZN(
        P3_U3473) );
  AOI211_X1 U15320 ( .C1(n12783), .C2(n15993), .A(n12782), .B(n12781), .ZN(
        n12788) );
  AOI22_X1 U15321 ( .A1(n14191), .A2(n12784), .B1(P2_REG1_REG_13__SCAN_IN), 
        .B2(n16008), .ZN(n12785) );
  OAI21_X1 U15322 ( .B1(n12788), .B2(n16008), .A(n12785), .ZN(P2_U3512) );
  INV_X1 U15323 ( .A(n14892), .ZN(n12786) );
  AOI22_X1 U15324 ( .A1(n14191), .A2(n12786), .B1(P2_REG0_REG_13__SCAN_IN), 
        .B2(n16002), .ZN(n12787) );
  OAI21_X1 U15325 ( .B1(n12788), .B2(n16002), .A(n12787), .ZN(P2_U3469) );
  INV_X1 U15326 ( .A(n12789), .ZN(n12793) );
  OAI222_X1 U15327 ( .A1(n14914), .A2(n12791), .B1(n14903), .B2(n12793), .C1(
        P2_U3088), .C2(n12790), .ZN(P2_U3302) );
  OAI222_X1 U15328 ( .A1(P1_U3086), .A2(n12794), .B1(n15703), .B2(n12793), 
        .C1(n12792), .C2(n15700), .ZN(P1_U3330) );
  NAND2_X1 U15329 ( .A1(n12797), .A2(n12806), .ZN(n12798) );
  NAND2_X1 U15330 ( .A1(n14497), .A2(n12798), .ZN(n12800) );
  INV_X1 U15331 ( .A(n14498), .ZN(n12799) );
  AOI21_X1 U15332 ( .B1(P2_REG2_REG_18__SCAN_IN), .B2(n12800), .A(n12799), 
        .ZN(n12814) );
  NAND2_X1 U15333 ( .A1(P2_U3088), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n14077)
         );
  OAI21_X1 U15334 ( .B1(n15919), .B2(n12801), .A(n14077), .ZN(n12802) );
  AOI21_X1 U15335 ( .B1(P2_ADDR_REG_18__SCAN_IN), .B2(n15899), .A(n12802), 
        .ZN(n12813) );
  NAND2_X1 U15336 ( .A1(n12803), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n12804) );
  NAND2_X1 U15337 ( .A1(n12805), .A2(n12804), .ZN(n12807) );
  NAND2_X1 U15338 ( .A1(n12807), .A2(n12806), .ZN(n14494) );
  OR2_X1 U15339 ( .A1(n12807), .A2(n12806), .ZN(n12808) );
  NAND2_X1 U15340 ( .A1(n14494), .A2(n12808), .ZN(n12810) );
  INV_X1 U15341 ( .A(n12810), .ZN(n12811) );
  INV_X1 U15342 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n12809) );
  OR2_X1 U15343 ( .A1(n12810), .A2(n12809), .ZN(n14495) );
  OAI211_X1 U15344 ( .C1(n12811), .C2(P2_REG1_REG_18__SCAN_IN), .A(n15928), 
        .B(n14495), .ZN(n12812) );
  OAI211_X1 U15345 ( .C1(n12814), .C2(n14504), .A(n12813), .B(n12812), .ZN(
        P2_U3232) );
  NAND2_X1 U15346 ( .A1(n14088), .A2(n12815), .ZN(n12817) );
  OAI211_X1 U15347 ( .C1(n12818), .C2(n14090), .A(n12817), .B(n12816), .ZN(
        n12823) );
  XNOR2_X1 U15348 ( .A(n12820), .B(n12819), .ZN(n12821) );
  NOR2_X1 U15349 ( .A1(n12821), .A2(n14103), .ZN(n12822) );
  AOI211_X1 U15350 ( .C1(n14842), .C2(n14101), .A(n12823), .B(n12822), .ZN(
        n12824) );
  INV_X1 U15351 ( .A(n12824), .ZN(P2_U3189) );
  INV_X1 U15352 ( .A(n10420), .ZN(n12833) );
  XNOR2_X1 U15353 ( .A(n14829), .B(n14410), .ZN(n14348) );
  XNOR2_X1 U15354 ( .A(n12825), .B(n14348), .ZN(n12838) );
  NAND2_X1 U15355 ( .A1(n12827), .A2(n12826), .ZN(n12828) );
  XOR2_X1 U15356 ( .A(n14348), .B(n12828), .Z(n12831) );
  NAND2_X1 U15357 ( .A1(n14411), .A2(n14376), .ZN(n12830) );
  NAND2_X1 U15358 ( .A1(n14409), .A2(n14086), .ZN(n12829) );
  AND2_X1 U15359 ( .A1(n12830), .A2(n12829), .ZN(n12894) );
  OAI21_X1 U15360 ( .B1(n12831), .B2(n8640), .A(n12894), .ZN(n12832) );
  AOI21_X1 U15361 ( .B1(n12833), .B2(n12838), .A(n12832), .ZN(n14831) );
  INV_X1 U15362 ( .A(n12834), .ZN(n12835) );
  AOI211_X1 U15363 ( .C1(n14829), .C2(n12836), .A(n14717), .B(n12835), .ZN(
        n14828) );
  AOI22_X1 U15364 ( .A1(n14738), .A2(P2_REG2_REG_12__SCAN_IN), .B1(n12896), 
        .B2(n14713), .ZN(n12837) );
  OAI21_X1 U15365 ( .B1(n14173), .B2(n14698), .A(n12837), .ZN(n12840) );
  INV_X1 U15366 ( .A(n12838), .ZN(n14832) );
  NOR2_X1 U15367 ( .A1(n14832), .A2(n14682), .ZN(n12839) );
  AOI211_X1 U15368 ( .C1(n14828), .C2(n14703), .A(n12840), .B(n12839), .ZN(
        n12841) );
  OAI21_X1 U15369 ( .B1(n14831), .B2(n14719), .A(n12841), .ZN(P2_U3253) );
  NAND2_X1 U15370 ( .A1(n12846), .A2(P3_ADDR_REG_12__SCAN_IN), .ZN(n12847) );
  INV_X1 U15371 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n12849) );
  NAND2_X1 U15372 ( .A1(n12849), .A2(P3_ADDR_REG_13__SCAN_IN), .ZN(n15715) );
  NAND2_X1 U15373 ( .A1(P1_ADDR_REG_13__SCAN_IN), .A2(n12850), .ZN(n15713) );
  AND2_X1 U15374 ( .A1(n15715), .A2(n15713), .ZN(n12851) );
  XNOR2_X1 U15375 ( .A(n15714), .B(n12851), .ZN(n15710) );
  XNOR2_X1 U15376 ( .A(n15710), .B(P2_ADDR_REG_13__SCAN_IN), .ZN(n12852) );
  XNOR2_X1 U15377 ( .A(n15709), .B(n12852), .ZN(SUB_1596_U67) );
  XOR2_X1 U15378 ( .A(n11436), .B(n12859), .Z(n12854) );
  NAND2_X1 U15379 ( .A1(n12855), .A2(n12854), .ZN(n12879) );
  INV_X1 U15380 ( .A(n12880), .ZN(n12856) );
  NAND2_X1 U15381 ( .A1(n12879), .A2(n12856), .ZN(n12858) );
  XNOR2_X1 U15382 ( .A(n12858), .B(n12857), .ZN(n12866) );
  NOR2_X1 U15383 ( .A1(n12859), .A2(n13276), .ZN(n12863) );
  NAND2_X1 U15384 ( .A1(n13269), .A2(n13503), .ZN(n12861) );
  OAI211_X1 U15385 ( .C1(n12934), .C2(n13271), .A(n12861), .B(n12860), .ZN(
        n12862) );
  AOI211_X1 U15386 ( .C1(n12864), .C2(n13273), .A(n12863), .B(n12862), .ZN(
        n12865) );
  OAI21_X1 U15387 ( .B1(n12866), .B2(n13264), .A(n12865), .ZN(P3_U3176) );
  INV_X1 U15388 ( .A(n12867), .ZN(n12868) );
  AOI21_X1 U15389 ( .B1(n12870), .B2(n12869), .A(n12868), .ZN(n12878) );
  INV_X1 U15390 ( .A(n12871), .ZN(n12875) );
  NAND2_X1 U15391 ( .A1(n14097), .A2(n12872), .ZN(n12873) );
  OAI211_X1 U15392 ( .C1(n14099), .C2(n12875), .A(n12874), .B(n12873), .ZN(
        n12876) );
  AOI21_X1 U15393 ( .B1(n14171), .B2(n14101), .A(n12876), .ZN(n12877) );
  OAI21_X1 U15394 ( .B1(n12878), .B2(n14103), .A(n12877), .ZN(P2_U3208) );
  XNOR2_X1 U15395 ( .A(n12886), .B(n11436), .ZN(n12933) );
  XNOR2_X1 U15396 ( .A(n12933), .B(n12934), .ZN(n12881) );
  XNOR2_X1 U15397 ( .A(n12932), .B(n12881), .ZN(n12888) );
  NAND2_X1 U15398 ( .A1(n13269), .A2(n13502), .ZN(n12882) );
  NAND2_X1 U15399 ( .A1(P3_U3151), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n13516)
         );
  OAI211_X1 U15400 ( .C1(n12937), .C2(n13271), .A(n12882), .B(n13516), .ZN(
        n12885) );
  NOR2_X1 U15401 ( .A1(n13226), .A2(n12883), .ZN(n12884) );
  AOI211_X1 U15402 ( .C1(n12886), .C2(n13261), .A(n12885), .B(n12884), .ZN(
        n12887) );
  OAI21_X1 U15403 ( .B1(n12888), .B2(n13264), .A(n12887), .ZN(P3_U3164) );
  OAI21_X1 U15404 ( .B1(n12891), .B2(n12890), .A(n12889), .ZN(n12892) );
  NAND2_X1 U15405 ( .A1(n12892), .A2(n14065), .ZN(n12898) );
  OAI21_X1 U15406 ( .B1(n14090), .B2(n12894), .A(n12893), .ZN(n12895) );
  AOI21_X1 U15407 ( .B1(n12896), .B2(n14088), .A(n12895), .ZN(n12897) );
  OAI211_X1 U15408 ( .C1(n14173), .C2(n14073), .A(n12898), .B(n12897), .ZN(
        P2_U3196) );
  INV_X1 U15409 ( .A(n14969), .ZN(n12899) );
  AOI21_X1 U15410 ( .B1(n12901), .B2(n12900), .A(n12899), .ZN(n12912) );
  NAND2_X1 U15411 ( .A1(n12902), .A2(n15870), .ZN(n15657) );
  INV_X1 U15412 ( .A(n15657), .ZN(n12909) );
  OAI22_X1 U15413 ( .A1(n15056), .A2(n12904), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n12903), .ZN(n12905) );
  AOI21_X1 U15414 ( .B1(n15053), .B2(n15520), .A(n12905), .ZN(n12906) );
  OAI21_X1 U15415 ( .B1(n15077), .B2(n12907), .A(n12906), .ZN(n12908) );
  AOI21_X1 U15416 ( .B1(n12910), .B2(n12909), .A(n12908), .ZN(n12911) );
  OAI21_X1 U15417 ( .B1(n12912), .B2(n15070), .A(n12911), .ZN(P1_U3236) );
  XNOR2_X1 U15418 ( .A(n12913), .B(n14328), .ZN(n12915) );
  AOI22_X1 U15419 ( .A1(n14407), .A2(n14086), .B1(n14409), .B2(n14376), .ZN(
        n13983) );
  INV_X1 U15420 ( .A(n13983), .ZN(n12914) );
  AOI21_X1 U15421 ( .B1(n12915), .B2(n14675), .A(n12914), .ZN(n14826) );
  XNOR2_X1 U15422 ( .A(n12916), .B(n14328), .ZN(n14827) );
  INV_X1 U15423 ( .A(n14827), .ZN(n12923) );
  INV_X1 U15424 ( .A(n14824), .ZN(n14187) );
  NAND2_X1 U15425 ( .A1(n12917), .A2(n14824), .ZN(n12918) );
  NAND2_X1 U15426 ( .A1(n12918), .A2(n14818), .ZN(n12919) );
  NOR2_X1 U15427 ( .A1(n14730), .A2(n12919), .ZN(n14823) );
  NAND2_X1 U15428 ( .A1(n14823), .A2(n14703), .ZN(n12921) );
  AOI22_X1 U15429 ( .A1(n14719), .A2(P2_REG2_REG_14__SCAN_IN), .B1(n13985), 
        .B2(n14713), .ZN(n12920) );
  OAI211_X1 U15430 ( .C1(n14187), .C2(n14698), .A(n12921), .B(n12920), .ZN(
        n12922) );
  AOI21_X1 U15431 ( .B1(n12923), .B2(n14723), .A(n12922), .ZN(n12924) );
  OAI21_X1 U15432 ( .B1(n14738), .B2(n14826), .A(n12924), .ZN(P2_U3251) );
  XNOR2_X1 U15433 ( .A(n13974), .B(n13973), .ZN(n12931) );
  OAI22_X1 U15434 ( .A1(n14090), .A2(n12926), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n12925), .ZN(n12928) );
  NOR2_X1 U15435 ( .A1(n6951), .A2(n14073), .ZN(n12927) );
  AOI211_X1 U15436 ( .C1(n14088), .C2(n12929), .A(n12928), .B(n12927), .ZN(
        n12930) );
  OAI21_X1 U15437 ( .B1(n12931), .B2(n14103), .A(n12930), .ZN(P2_U3206) );
  OAI21_X1 U15438 ( .B1(n12934), .B2(n12933), .A(n12932), .ZN(n12935) );
  XNOR2_X1 U15439 ( .A(n13223), .B(n11436), .ZN(n13220) );
  NOR2_X1 U15440 ( .A1(n13220), .A2(n13500), .ZN(n12938) );
  INV_X1 U15441 ( .A(n13220), .ZN(n12936) );
  XNOR2_X1 U15442 ( .A(n13404), .B(n11436), .ZN(n12939) );
  XNOR2_X1 U15443 ( .A(n12939), .B(n13499), .ZN(n13152) );
  INV_X1 U15444 ( .A(n12939), .ZN(n12940) );
  XNOR2_X1 U15445 ( .A(n13952), .B(n11436), .ZN(n12941) );
  XNOR2_X1 U15446 ( .A(n12941), .B(n13804), .ZN(n13265) );
  INV_X1 U15447 ( .A(n12941), .ZN(n12942) );
  XNOR2_X1 U15448 ( .A(n13942), .B(n11436), .ZN(n13187) );
  NOR2_X1 U15449 ( .A1(n13187), .A2(n13818), .ZN(n12943) );
  NAND2_X1 U15450 ( .A1(n13187), .A2(n13818), .ZN(n12944) );
  XNOR2_X1 U15451 ( .A(n13939), .B(n11436), .ZN(n12946) );
  XNOR2_X1 U15452 ( .A(n12946), .B(n13805), .ZN(n13194) );
  INV_X1 U15453 ( .A(n13194), .ZN(n12945) );
  INV_X1 U15454 ( .A(n12946), .ZN(n12947) );
  NAND2_X1 U15455 ( .A1(n12947), .A2(n13774), .ZN(n12948) );
  XNOR2_X1 U15456 ( .A(n13868), .B(n11436), .ZN(n12949) );
  XNOR2_X1 U15457 ( .A(n12949), .B(n13496), .ZN(n13245) );
  INV_X1 U15458 ( .A(n12949), .ZN(n12950) );
  NAND2_X1 U15459 ( .A1(n12950), .A2(n13496), .ZN(n12951) );
  NAND2_X1 U15460 ( .A1(n13244), .A2(n12951), .ZN(n13166) );
  XNOR2_X1 U15461 ( .A(n13172), .B(n6554), .ZN(n12952) );
  XNOR2_X1 U15462 ( .A(n12952), .B(n13748), .ZN(n13165) );
  NAND2_X1 U15463 ( .A1(n13166), .A2(n13165), .ZN(n13164) );
  NAND2_X1 U15464 ( .A1(n12952), .A2(n13775), .ZN(n12953) );
  XNOR2_X1 U15465 ( .A(n13922), .B(n11436), .ZN(n12954) );
  XNOR2_X1 U15466 ( .A(n12954), .B(n13495), .ZN(n13213) );
  INV_X1 U15467 ( .A(n12954), .ZN(n12955) );
  NAND2_X1 U15468 ( .A1(n12955), .A2(n13495), .ZN(n12956) );
  XNOR2_X1 U15469 ( .A(n13734), .B(n11436), .ZN(n12958) );
  XNOR2_X1 U15470 ( .A(n12958), .B(n13749), .ZN(n13175) );
  XNOR2_X1 U15471 ( .A(n13911), .B(n11436), .ZN(n13234) );
  INV_X1 U15472 ( .A(n12958), .ZN(n12959) );
  NOR2_X1 U15473 ( .A1(n12959), .A2(n13721), .ZN(n13232) );
  AOI21_X1 U15474 ( .B1(n13733), .B2(n13234), .A(n13232), .ZN(n12960) );
  INV_X1 U15475 ( .A(n13234), .ZN(n12961) );
  NAND2_X1 U15476 ( .A1(n12961), .A2(n13705), .ZN(n12962) );
  XNOR2_X1 U15477 ( .A(n13899), .B(n11436), .ZN(n13206) );
  XNOR2_X1 U15478 ( .A(n13850), .B(n11436), .ZN(n12964) );
  OAI22_X1 U15479 ( .A1(n13206), .A2(n13683), .B1(n13444), .B2(n12964), .ZN(
        n12968) );
  INV_X1 U15480 ( .A(n12964), .ZN(n13204) );
  OAI21_X1 U15481 ( .B1(n13204), .B2(n13722), .A(n7128), .ZN(n12966) );
  NOR2_X1 U15482 ( .A1(n7128), .A2(n13722), .ZN(n12965) );
  AOI22_X1 U15483 ( .A1(n13206), .A2(n12966), .B1(n12965), .B2(n12964), .ZN(
        n12967) );
  XNOR2_X1 U15484 ( .A(n13841), .B(n6554), .ZN(n12973) );
  XNOR2_X1 U15485 ( .A(n12973), .B(n6947), .ZN(n13254) );
  XNOR2_X1 U15486 ( .A(n13836), .B(n11436), .ZN(n12969) );
  NAND2_X1 U15487 ( .A1(n12969), .A2(n13684), .ZN(n12974) );
  INV_X1 U15488 ( .A(n12974), .ZN(n12970) );
  XNOR2_X1 U15489 ( .A(n12969), .B(n13494), .ZN(n13257) );
  AND2_X1 U15490 ( .A1(n13254), .A2(n12972), .ZN(n12971) );
  INV_X1 U15491 ( .A(n12972), .ZN(n12976) );
  NAND2_X1 U15492 ( .A1(n12973), .A2(n13209), .ZN(n13256) );
  AND2_X1 U15493 ( .A1(n13256), .A2(n12974), .ZN(n12975) );
  XNOR2_X1 U15494 ( .A(n13460), .B(n11436), .ZN(n13136) );
  XNOR2_X1 U15495 ( .A(n13136), .B(n13666), .ZN(n13138) );
  XOR2_X1 U15496 ( .A(n13139), .B(n13138), .Z(n12982) );
  AOI22_X1 U15497 ( .A1(n13658), .A2(n13273), .B1(P3_REG3_REG_27__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12978) );
  NAND2_X1 U15498 ( .A1(n13494), .A2(n13269), .ZN(n12977) );
  OAI211_X1 U15499 ( .C1(n12979), .C2(n13271), .A(n12978), .B(n12977), .ZN(
        n12980) );
  AOI21_X1 U15500 ( .B1(n13460), .B2(n13261), .A(n12980), .ZN(n12981) );
  OAI21_X1 U15501 ( .B1(n12982), .B2(n13264), .A(n12981), .ZN(P3_U3154) );
  INV_X1 U15502 ( .A(n12983), .ZN(n12985) );
  OAI222_X1 U15503 ( .A1(n12986), .A2(P3_U3151), .B1(n13102), .B2(n12985), 
        .C1(n12984), .C2(n13970), .ZN(P3_U3271) );
  AOI21_X2 U15504 ( .B1(n13133), .B2(n13125), .A(n7982), .ZN(n14511) );
  OAI211_X1 U15505 ( .C1(n14511), .C2(n12987), .A(n14818), .B(n13129), .ZN(
        n14515) );
  NAND2_X1 U15506 ( .A1(n12988), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n12992) );
  NAND2_X1 U15507 ( .A1(n8643), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n12991) );
  NAND2_X1 U15508 ( .A1(n12989), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n12990) );
  OR2_X1 U15509 ( .A1(n14317), .A2(n12993), .ZN(n14507) );
  NAND2_X1 U15510 ( .A1(n14515), .A2(n14507), .ZN(n12996) );
  INV_X1 U15511 ( .A(n12994), .ZN(n12995) );
  OAI21_X1 U15512 ( .B1(n14511), .B2(n14892), .A(n12995), .ZN(P2_U3497) );
  INV_X1 U15513 ( .A(n12997), .ZN(n12998) );
  OAI21_X1 U15514 ( .B1(n14511), .B2(n14840), .A(n12998), .ZN(P2_U3529) );
  OR2_X1 U15515 ( .A1(n15651), .A2(n15520), .ZN(n12999) );
  OR2_X1 U15516 ( .A1(n15645), .A2(n15502), .ZN(n13001) );
  NAND2_X1 U15517 ( .A1(n15639), .A2(n15091), .ZN(n15482) );
  NAND2_X1 U15518 ( .A1(n15481), .A2(n13002), .ZN(n13005) );
  OR2_X1 U15519 ( .A1(n15628), .A2(n15090), .ZN(n13006) );
  NAND2_X1 U15520 ( .A1(n15622), .A2(n15089), .ZN(n13007) );
  OR2_X1 U15521 ( .A1(n15622), .A2(n15089), .ZN(n13008) );
  OR2_X1 U15522 ( .A1(n15605), .A2(n15088), .ZN(n15382) );
  NAND2_X1 U15523 ( .A1(n13039), .A2(n15382), .ZN(n15371) );
  NOR2_X1 U15524 ( .A1(n15597), .A2(n15363), .ZN(n13014) );
  NOR2_X1 U15525 ( .A1(n15371), .A2(n13014), .ZN(n13013) );
  NAND2_X1 U15526 ( .A1(n15602), .A2(n15421), .ZN(n15384) );
  NAND2_X1 U15527 ( .A1(n15385), .A2(n15384), .ZN(n15375) );
  INV_X1 U15528 ( .A(n13014), .ZN(n15373) );
  AOI21_X1 U15529 ( .B1(n15375), .B2(n15373), .A(n15374), .ZN(n13015) );
  NAND2_X1 U15530 ( .A1(n13016), .A2(n13015), .ZN(n15378) );
  NAND2_X1 U15531 ( .A1(n15370), .A2(n15391), .ZN(n13017) );
  NAND2_X1 U15532 ( .A1(n15586), .A2(n15362), .ZN(n13018) );
  NAND2_X1 U15533 ( .A1(n15578), .A2(n13045), .ZN(n13020) );
  NAND2_X1 U15534 ( .A1(n15318), .A2(n15330), .ZN(n13022) );
  NAND2_X2 U15535 ( .A1(n15308), .A2(n13022), .ZN(n15288) );
  INV_X1 U15536 ( .A(n15532), .ZN(n13026) );
  OR2_X1 U15537 ( .A1(n15645), .A2(n13027), .ZN(n13028) );
  INV_X1 U15538 ( .A(n15485), .ZN(n13031) );
  NAND2_X1 U15539 ( .A1(n15628), .A2(n15076), .ZN(n13034) );
  INV_X1 U15540 ( .A(n15450), .ZN(n13035) );
  OR2_X1 U15541 ( .A1(n15622), .A2(n15432), .ZN(n13036) );
  INV_X1 U15542 ( .A(n15419), .ZN(n14952) );
  OR2_X1 U15543 ( .A1(n15616), .A2(n14952), .ZN(n13037) );
  INV_X1 U15544 ( .A(n15374), .ZN(n15361) );
  NAND2_X1 U15545 ( .A1(n15318), .A2(n13043), .ZN(n15292) );
  NAND2_X1 U15546 ( .A1(n15341), .A2(n13045), .ZN(n13044) );
  NAND2_X1 U15547 ( .A1(n15586), .A2(n15332), .ZN(n15305) );
  AND2_X1 U15548 ( .A1(n13044), .A2(n15305), .ZN(n15289) );
  INV_X1 U15549 ( .A(n15293), .ZN(n13051) );
  OAI21_X1 U15550 ( .B1(n15586), .B2(n15332), .A(n13045), .ZN(n13047) );
  AND2_X1 U15551 ( .A1(n15306), .A2(n15362), .ZN(n13046) );
  AOI22_X1 U15552 ( .A1(n15578), .A2(n13047), .B1(n15356), .B2(n13046), .ZN(
        n13048) );
  AND2_X1 U15553 ( .A1(n15311), .A2(n13048), .ZN(n15290) );
  INV_X1 U15554 ( .A(n15292), .ZN(n13049) );
  OAI22_X1 U15555 ( .A1(n14927), .A2(n15516), .B1(n13055), .B2(n15431), .ZN(
        n13056) );
  INV_X1 U15556 ( .A(n13056), .ZN(n13057) );
  INV_X1 U15557 ( .A(n15639), .ZN(n15511) );
  INV_X1 U15558 ( .A(n15622), .ZN(n15459) );
  INV_X1 U15559 ( .A(n15616), .ZN(n15444) );
  NAND2_X1 U15560 ( .A1(n15392), .A2(n15370), .ZN(n15365) );
  NOR2_X2 U15561 ( .A1(n15365), .A2(n15586), .ZN(n13058) );
  INV_X1 U15562 ( .A(n15277), .ZN(n13059) );
  NAND2_X1 U15563 ( .A1(n15558), .A2(n15812), .ZN(n13062) );
  INV_X1 U15564 ( .A(n13060), .ZN(n14924) );
  AOI22_X1 U15565 ( .A1(n14924), .A2(n15525), .B1(P1_REG2_REG_27__SCAN_IN), 
        .B2(n6556), .ZN(n13061) );
  OAI211_X1 U15566 ( .C1(n13087), .C2(n15807), .A(n13062), .B(n13061), .ZN(
        n13063) );
  AOI21_X1 U15567 ( .B1(n15557), .B2(n15813), .A(n13063), .ZN(n13064) );
  OAI21_X1 U15568 ( .B1(n15561), .B2(n6556), .A(n13064), .ZN(P1_U3266) );
  OR2_X1 U15569 ( .A1(n7122), .A2(n15297), .ZN(n15267) );
  NAND2_X1 U15570 ( .A1(n13065), .A2(n15267), .ZN(n13071) );
  NAND2_X1 U15571 ( .A1(n15553), .A2(n15085), .ZN(n13073) );
  INV_X1 U15572 ( .A(n13073), .ZN(n13069) );
  AOI21_X1 U15573 ( .B1(n13071), .B2(n13073), .A(n13067), .ZN(n13072) );
  AOI21_X1 U15574 ( .B1(n13067), .B2(n13073), .A(n13072), .ZN(n13074) );
  INV_X1 U15575 ( .A(n15280), .ZN(n13077) );
  AOI21_X1 U15576 ( .B1(n13077), .B2(n13076), .A(n15260), .ZN(n15549) );
  NOR3_X1 U15577 ( .A1(n13079), .A2(n13078), .A3(n15804), .ZN(n13083) );
  NOR2_X1 U15578 ( .A1(n15699), .A2(n13080), .ZN(n13081) );
  NOR2_X1 U15579 ( .A1(n15516), .A2(n13081), .ZN(n15255) );
  AOI22_X1 U15580 ( .A1(n15085), .A2(n15521), .B1(n15255), .B2(n15084), .ZN(
        n15546) );
  NOR2_X1 U15581 ( .A1(n15546), .A2(n6556), .ZN(n13082) );
  AOI211_X1 U15582 ( .C1(n6556), .C2(P1_REG2_REG_29__SCAN_IN), .A(n13083), .B(
        n13082), .ZN(n13084) );
  OAI21_X1 U15583 ( .B1(n15547), .B2(n15807), .A(n13084), .ZN(n13085) );
  AOI21_X1 U15584 ( .B1(n15549), .B2(n13086), .A(n13085), .ZN(n13090) );
  NAND2_X1 U15585 ( .A1(n15545), .A2(n15428), .ZN(n13089) );
  OAI211_X1 U15586 ( .C1(n15551), .C2(n15535), .A(n13090), .B(n13089), .ZN(
        P1_U3356) );
  OAI22_X1 U15587 ( .A1(n15056), .A2(n10123), .B1(n7219), .B2(n15065), .ZN(
        n13091) );
  AOI21_X1 U15588 ( .B1(P1_REG3_REG_2__SCAN_IN), .B2(n13092), .A(n13091), .ZN(
        n13098) );
  OAI21_X1 U15589 ( .B1(n13095), .B2(n13094), .A(n13093), .ZN(n13096) );
  NAND2_X1 U15590 ( .A1(n13096), .A2(n15072), .ZN(n13097) );
  OAI211_X1 U15591 ( .C1(n15834), .C2(n15083), .A(n13098), .B(n13097), .ZN(
        P1_U3237) );
  NAND2_X1 U15592 ( .A1(n15694), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n13099) );
  INV_X1 U15593 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n14900) );
  XNOR2_X1 U15594 ( .A(n14900), .B(P2_DATAO_REG_30__SCAN_IN), .ZN(n13279) );
  XNOR2_X1 U15595 ( .A(n13280), .B(n13279), .ZN(n13295) );
  INV_X1 U15596 ( .A(n13295), .ZN(n13101) );
  OAI222_X1 U15597 ( .A1(n14914), .A2(n13105), .B1(n14917), .B2(n13104), .C1(
        n8584), .C2(P2_U3088), .ZN(P2_U3308) );
  INV_X1 U15598 ( .A(n14907), .ZN(n13107) );
  OAI222_X1 U15599 ( .A1(n15119), .A2(P1_U3086), .B1(n15703), .B2(n13107), 
        .C1(n13106), .C2(n13134), .ZN(P1_U3327) );
  INV_X1 U15600 ( .A(n13108), .ZN(n13110) );
  OAI222_X1 U15601 ( .A1(n13102), .A2(n13110), .B1(n13970), .B2(n13109), .C1(
        P3_U3151), .C2(n8892), .ZN(P3_U3268) );
  NAND2_X1 U15602 ( .A1(n14394), .A2(n13111), .ZN(n13113) );
  XNOR2_X1 U15603 ( .A(n13113), .B(n13112), .ZN(n13114) );
  XNOR2_X1 U15604 ( .A(n14519), .B(n13114), .ZN(n13115) );
  INV_X1 U15605 ( .A(n13115), .ZN(n13120) );
  AOI22_X1 U15606 ( .A1(n14517), .A2(n14088), .B1(P2_REG3_REG_28__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13117) );
  OAI21_X1 U15607 ( .B1(n13118), .B2(n14090), .A(n13117), .ZN(n13122) );
  NOR3_X1 U15608 ( .A1(n13120), .A2(n13119), .A3(n14103), .ZN(n13121) );
  AOI211_X1 U15609 ( .C1(n14519), .C2(n14101), .A(n13122), .B(n13121), .ZN(
        n13123) );
  NAND2_X1 U15610 ( .A1(n14895), .A2(n13125), .ZN(n13128) );
  NAND2_X1 U15611 ( .A1(n7193), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(n13127) );
  XNOR2_X1 U15612 ( .A(n13129), .B(n14849), .ZN(n13130) );
  NAND2_X1 U15613 ( .A1(n14510), .A2(n14507), .ZN(n14847) );
  OAI222_X1 U15614 ( .A1(P3_U3151), .A2(n8905), .B1(n13102), .B2(n13132), .C1(
        n13131), .C2(n13970), .ZN(P3_U3266) );
  INV_X1 U15615 ( .A(n13133), .ZN(n14901) );
  INV_X1 U15616 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n13278) );
  OAI222_X1 U15617 ( .A1(n15703), .A2(n14901), .B1(n13135), .B2(P1_U3086), 
        .C1(n13278), .C2(n13134), .ZN(P1_U3325) );
  AND2_X1 U15618 ( .A1(n13136), .A2(n13461), .ZN(n13137) );
  AOI21_X1 U15619 ( .B1(n13139), .B2(n13138), .A(n13137), .ZN(n13141) );
  XNOR2_X1 U15620 ( .A(n13469), .B(n6554), .ZN(n13140) );
  XNOR2_X1 U15621 ( .A(n13141), .B(n13140), .ZN(n13147) );
  AOI22_X1 U15622 ( .A1(n13652), .A2(n13273), .B1(P3_REG3_REG_28__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13143) );
  NAND2_X1 U15623 ( .A1(n13666), .A2(n13269), .ZN(n13142) );
  OAI211_X1 U15624 ( .C1(n13300), .C2(n13271), .A(n13143), .B(n13142), .ZN(
        n13144) );
  AOI21_X1 U15625 ( .B1(n13145), .B2(n13261), .A(n13144), .ZN(n13146) );
  OAI21_X1 U15626 ( .B1(n13147), .B2(n13264), .A(n13146), .ZN(P3_U3160) );
  INV_X1 U15627 ( .A(n13148), .ZN(n13150) );
  OAI222_X1 U15628 ( .A1(n13102), .A2(n13150), .B1(n13970), .B2(n13149), .C1(
        P3_U3151), .C2(n11431), .ZN(P3_U3274) );
  AOI21_X1 U15629 ( .B1(n13152), .B2(n13151), .A(n6719), .ZN(n13158) );
  NAND2_X1 U15630 ( .A1(n13269), .A2(n13500), .ZN(n13153) );
  NAND2_X1 U15631 ( .A1(P3_U3151), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n13554)
         );
  OAI211_X1 U15632 ( .C1(n13804), .C2(n13271), .A(n13153), .B(n13554), .ZN(
        n13155) );
  NOR2_X1 U15633 ( .A1(n13404), .A2(n13276), .ZN(n13154) );
  AOI211_X1 U15634 ( .C1(n13156), .C2(n13273), .A(n13155), .B(n13154), .ZN(
        n13157) );
  OAI21_X1 U15635 ( .B1(n13158), .B2(n13264), .A(n13157), .ZN(P3_U3155) );
  XNOR2_X1 U15636 ( .A(n13205), .B(n13444), .ZN(n13163) );
  AOI22_X1 U15637 ( .A1(n13705), .A2(n13269), .B1(P3_REG3_REG_23__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13160) );
  NAND2_X1 U15638 ( .A1(n13712), .A2(n13273), .ZN(n13159) );
  OAI211_X1 U15639 ( .C1(n13683), .C2(n13271), .A(n13160), .B(n13159), .ZN(
        n13161) );
  AOI21_X1 U15640 ( .B1(n13850), .B2(n13261), .A(n13161), .ZN(n13162) );
  OAI21_X1 U15641 ( .B1(n13163), .B2(n13264), .A(n13162), .ZN(P3_U3156) );
  OAI211_X1 U15642 ( .C1(n13166), .C2(n13165), .A(n13164), .B(n13243), .ZN(
        n13171) );
  NAND2_X1 U15643 ( .A1(n13496), .A2(n13269), .ZN(n13168) );
  OAI211_X1 U15644 ( .C1(n13761), .C2(n13271), .A(n13168), .B(n13167), .ZN(
        n13169) );
  AOI21_X1 U15645 ( .B1(n13757), .B2(n13273), .A(n13169), .ZN(n13170) );
  OAI211_X1 U15646 ( .C1(n13276), .C2(n13172), .A(n13171), .B(n13170), .ZN(
        P3_U3159) );
  INV_X1 U15647 ( .A(n13173), .ZN(n13233) );
  AOI21_X1 U15648 ( .B1(n13175), .B2(n13174), .A(n13233), .ZN(n13180) );
  AOI22_X1 U15649 ( .A1(n13495), .A2(n13269), .B1(P3_REG3_REG_21__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13177) );
  NAND2_X1 U15650 ( .A1(n13735), .A2(n13273), .ZN(n13176) );
  OAI211_X1 U15651 ( .C1(n13733), .C2(n13271), .A(n13177), .B(n13176), .ZN(
        n13178) );
  AOI21_X1 U15652 ( .B1(n13734), .B2(n13261), .A(n13178), .ZN(n13179) );
  OAI21_X1 U15653 ( .B1(n13180), .B2(n13264), .A(n13179), .ZN(P3_U3163) );
  XOR2_X1 U15654 ( .A(n13254), .B(n13255), .Z(n13185) );
  AOI22_X1 U15655 ( .A1(n7128), .A2(n13269), .B1(P3_REG3_REG_25__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13182) );
  NAND2_X1 U15656 ( .A1(n13688), .A2(n13273), .ZN(n13181) );
  OAI211_X1 U15657 ( .C1(n13684), .C2(n13271), .A(n13182), .B(n13181), .ZN(
        n13183) );
  AOI21_X1 U15658 ( .B1(n13841), .B2(n13261), .A(n13183), .ZN(n13184) );
  OAI21_X1 U15659 ( .B1(n13185), .B2(n13264), .A(n13184), .ZN(P3_U3165) );
  XNOR2_X1 U15660 ( .A(n13187), .B(n13497), .ZN(n13188) );
  XNOR2_X1 U15661 ( .A(n13186), .B(n13188), .ZN(n13193) );
  NAND2_X1 U15662 ( .A1(n13269), .A2(n13498), .ZN(n13189) );
  NAND2_X1 U15663 ( .A1(P3_U3151), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n13593)
         );
  OAI211_X1 U15664 ( .C1(n13805), .C2(n13271), .A(n13189), .B(n13593), .ZN(
        n13190) );
  AOI21_X1 U15665 ( .B1(n13799), .B2(n13273), .A(n13190), .ZN(n13192) );
  NAND2_X1 U15666 ( .A1(n13942), .A2(n13261), .ZN(n13191) );
  OAI211_X1 U15667 ( .C1(n13193), .C2(n13264), .A(n13192), .B(n13191), .ZN(
        P3_U3166) );
  INV_X1 U15668 ( .A(n13939), .ZN(n13202) );
  AOI21_X1 U15669 ( .B1(n13195), .B2(n13194), .A(n13264), .ZN(n13197) );
  NAND2_X1 U15670 ( .A1(n13197), .A2(n13196), .ZN(n13201) );
  NAND2_X1 U15671 ( .A1(n13269), .A2(n13497), .ZN(n13198) );
  NAND2_X1 U15672 ( .A1(P3_U3151), .A2(P3_REG3_REG_17__SCAN_IN), .ZN(n13615)
         );
  OAI211_X1 U15673 ( .C1(n13791), .C2(n13271), .A(n13198), .B(n13615), .ZN(
        n13199) );
  AOI21_X1 U15674 ( .B1(n13785), .B2(n13273), .A(n13199), .ZN(n13200) );
  OAI211_X1 U15675 ( .C1(n13202), .C2(n13276), .A(n13201), .B(n13200), .ZN(
        P3_U3168) );
  AOI22_X1 U15676 ( .A1(n13722), .A2(n13269), .B1(P3_REG3_REG_24__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13208) );
  NAND2_X1 U15677 ( .A1(n13695), .A2(n13273), .ZN(n13207) );
  OAI211_X1 U15678 ( .C1(n13209), .C2(n13271), .A(n13208), .B(n13207), .ZN(
        n13210) );
  AOI21_X1 U15679 ( .B1(n13899), .B2(n13261), .A(n13210), .ZN(n13211) );
  INV_X1 U15680 ( .A(n13922), .ZN(n13219) );
  OAI211_X1 U15681 ( .C1(n13214), .C2(n13213), .A(n13212), .B(n13243), .ZN(
        n13218) );
  AOI22_X1 U15682 ( .A1(n13721), .A2(n13247), .B1(P3_REG3_REG_20__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13215) );
  OAI21_X1 U15683 ( .B1(n13748), .B2(n13249), .A(n13215), .ZN(n13216) );
  AOI21_X1 U15684 ( .B1(n13743), .B2(n13273), .A(n13216), .ZN(n13217) );
  OAI211_X1 U15685 ( .C1(n13219), .C2(n13276), .A(n13218), .B(n13217), .ZN(
        P3_U3173) );
  XNOR2_X1 U15686 ( .A(n13220), .B(n13500), .ZN(n13221) );
  XNOR2_X1 U15687 ( .A(n13222), .B(n13221), .ZN(n13231) );
  INV_X1 U15688 ( .A(n13223), .ZN(n13229) );
  AND2_X1 U15689 ( .A1(P3_U3151), .A2(P3_REG3_REG_13__SCAN_IN), .ZN(n13540) );
  NOR2_X1 U15690 ( .A1(n13271), .A2(n13816), .ZN(n13224) );
  AOI211_X1 U15691 ( .C1(n13269), .C2(n13501), .A(n13540), .B(n13224), .ZN(
        n13225) );
  OAI21_X1 U15692 ( .B1(n13227), .B2(n13226), .A(n13225), .ZN(n13228) );
  AOI21_X1 U15693 ( .B1(n13229), .B2(n13261), .A(n13228), .ZN(n13230) );
  OAI21_X1 U15694 ( .B1(n13231), .B2(n13264), .A(n13230), .ZN(P3_U3174) );
  NOR2_X1 U15695 ( .A1(n13233), .A2(n13232), .ZN(n13236) );
  XNOR2_X1 U15696 ( .A(n13234), .B(n13705), .ZN(n13235) );
  XNOR2_X1 U15697 ( .A(n13236), .B(n13235), .ZN(n13242) );
  INV_X1 U15698 ( .A(P3_REG3_REG_22__SCAN_IN), .ZN(n13237) );
  OAI22_X1 U15699 ( .A1(n13749), .A2(n13249), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n13237), .ZN(n13239) );
  NOR2_X1 U15700 ( .A1(n13444), .A2(n13271), .ZN(n13238) );
  AOI211_X1 U15701 ( .C1(n13718), .C2(n13273), .A(n13239), .B(n13238), .ZN(
        n13241) );
  NAND2_X1 U15702 ( .A1(n13911), .A2(n13261), .ZN(n13240) );
  OAI211_X1 U15703 ( .C1(n13242), .C2(n13264), .A(n13241), .B(n13240), .ZN(
        P3_U3175) );
  INV_X1 U15704 ( .A(n13868), .ZN(n13253) );
  OAI211_X1 U15705 ( .C1(n13246), .C2(n13245), .A(n13244), .B(n13243), .ZN(
        n13252) );
  NAND2_X1 U15706 ( .A1(n13775), .A2(n13247), .ZN(n13248) );
  NAND2_X1 U15707 ( .A1(P3_U3151), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n13634)
         );
  OAI211_X1 U15708 ( .C1(n13249), .C2(n13805), .A(n13248), .B(n13634), .ZN(
        n13250) );
  AOI21_X1 U15709 ( .B1(n13778), .B2(n13273), .A(n13250), .ZN(n13251) );
  OAI211_X1 U15710 ( .C1(n13253), .C2(n13276), .A(n13252), .B(n13251), .ZN(
        P3_U3178) );
  AOI22_X1 U15711 ( .A1(n6947), .A2(n13269), .B1(P3_REG3_REG_26__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13259) );
  NAND2_X1 U15712 ( .A1(n13670), .A2(n13273), .ZN(n13258) );
  OAI211_X1 U15713 ( .C1(n13461), .C2(n13271), .A(n13259), .B(n13258), .ZN(
        n13260) );
  AOI21_X1 U15714 ( .B1(n13836), .B2(n13261), .A(n13260), .ZN(n13262) );
  OAI21_X1 U15715 ( .B1(n13263), .B2(n13264), .A(n13262), .ZN(P3_U3180) );
  INV_X1 U15716 ( .A(n13952), .ZN(n13277) );
  AOI21_X1 U15717 ( .B1(n13266), .B2(n13265), .A(n13264), .ZN(n13268) );
  NAND2_X1 U15718 ( .A1(n13268), .A2(n13267), .ZN(n13275) );
  NAND2_X1 U15719 ( .A1(n13269), .A2(n13499), .ZN(n13270) );
  NAND2_X1 U15720 ( .A1(P3_U3151), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n13574)
         );
  OAI211_X1 U15721 ( .C1(n13818), .C2(n13271), .A(n13270), .B(n13574), .ZN(
        n13272) );
  AOI21_X1 U15722 ( .B1(n13813), .B2(n13273), .A(n13272), .ZN(n13274) );
  OAI211_X1 U15723 ( .C1(n13277), .C2(n13276), .A(n13275), .B(n13274), .ZN(
        P3_U3181) );
  XNOR2_X1 U15724 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(P2_DATAO_REG_31__SCAN_IN), 
        .ZN(n13281) );
  NAND2_X1 U15725 ( .A1(n13967), .A2(n6564), .ZN(n13284) );
  OR2_X1 U15726 ( .A1(n6568), .A2(n13963), .ZN(n13283) );
  INV_X1 U15727 ( .A(n13825), .ZN(n13890) );
  INV_X1 U15728 ( .A(P3_REG1_REG_31__SCAN_IN), .ZN(n13827) );
  NAND2_X1 U15729 ( .A1(n13285), .A2(P3_REG0_REG_31__SCAN_IN), .ZN(n13287) );
  INV_X1 U15730 ( .A(P3_REG2_REG_31__SCAN_IN), .ZN(n13649) );
  OR2_X1 U15731 ( .A1(n9311), .A2(n13649), .ZN(n13286) );
  OAI211_X1 U15732 ( .C1(n7094), .C2(n13827), .A(n13287), .B(n13286), .ZN(
        n13288) );
  INV_X1 U15733 ( .A(n13288), .ZN(n13289) );
  INV_X1 U15734 ( .A(n13491), .ZN(n13297) );
  NOR2_X1 U15735 ( .A1(n6569), .A2(n13291), .ZN(n13293) );
  INV_X1 U15736 ( .A(n13893), .ZN(n13296) );
  OAI21_X1 U15737 ( .B1(n13474), .B2(n13309), .A(n13825), .ZN(n13298) );
  INV_X1 U15738 ( .A(n13298), .ZN(n13305) );
  INV_X1 U15739 ( .A(n13300), .ZN(n13492) );
  NOR4_X1 U15740 ( .A1(n13474), .A2(n13301), .A3(n13309), .A4(n13492), .ZN(
        n13303) );
  AOI21_X1 U15741 ( .B1(n13893), .B2(n13472), .A(n13825), .ZN(n13302) );
  NOR2_X1 U15742 ( .A1(n13303), .A2(n13302), .ZN(n13304) );
  XNOR2_X1 U15743 ( .A(n13307), .B(n13306), .ZN(n13484) );
  INV_X1 U15744 ( .A(n13308), .ZN(n13483) );
  AND2_X1 U15745 ( .A1(n13825), .A2(n13309), .ZN(n13477) );
  INV_X1 U15746 ( .A(n13310), .ZN(n13455) );
  INV_X1 U15747 ( .A(n13696), .ZN(n13331) );
  INV_X1 U15748 ( .A(n13313), .ZN(n13362) );
  NAND4_X1 U15749 ( .A1(n13314), .A2(n16027), .A3(n13362), .A4(n13370), .ZN(
        n13320) );
  INV_X1 U15750 ( .A(n16052), .ZN(n13318) );
  NAND4_X1 U15751 ( .A1(n13318), .A2(n13317), .A3(n13316), .A4(n13315), .ZN(
        n13319) );
  NOR3_X1 U15752 ( .A1(n13320), .A2(n13319), .A3(n13373), .ZN(n13321) );
  NAND4_X1 U15753 ( .A1(n13321), .A2(n7844), .A3(n13381), .A4(n13390), .ZN(
        n13322) );
  NOR2_X1 U15754 ( .A1(n13323), .A2(n13322), .ZN(n13324) );
  AND4_X1 U15755 ( .A1(n13797), .A2(n13398), .A3(n13324), .A4(n7547), .ZN(
        n13326) );
  NAND4_X1 U15756 ( .A1(n13770), .A2(n13788), .A3(n13326), .A4(n13325), .ZN(
        n13327) );
  OR3_X1 U15757 ( .A1(n13720), .A2(n9209), .A3(n13327), .ZN(n13328) );
  OR4_X1 U15758 ( .A1(n9236), .A2(n13710), .A3(n13329), .A4(n13328), .ZN(
        n13330) );
  NAND2_X1 U15759 ( .A1(n13335), .A2(n13333), .ZN(n13334) );
  NAND2_X1 U15760 ( .A1(n13334), .A2(n13450), .ZN(n13337) );
  NAND3_X1 U15761 ( .A1(n13342), .A2(n13335), .A3(n13487), .ZN(n13336) );
  NAND2_X1 U15762 ( .A1(n13337), .A2(n13336), .ZN(n13341) );
  NAND2_X1 U15763 ( .A1(n13354), .A2(n13338), .ZN(n13346) );
  INV_X1 U15764 ( .A(n13346), .ZN(n13344) );
  NAND2_X1 U15765 ( .A1(n13339), .A2(n11431), .ZN(n13340) );
  INV_X1 U15766 ( .A(n13342), .ZN(n13343) );
  OAI21_X1 U15767 ( .B1(n9402), .B2(n13450), .A(n13351), .ZN(n13345) );
  INV_X1 U15768 ( .A(n13345), .ZN(n13350) );
  NAND2_X1 U15769 ( .A1(n13346), .A2(n13450), .ZN(n13348) );
  NAND2_X1 U15770 ( .A1(n13348), .A2(n13347), .ZN(n13349) );
  NAND2_X1 U15771 ( .A1(n13352), .A2(n13468), .ZN(n13353) );
  NOR2_X1 U15772 ( .A1(n13354), .A2(n13450), .ZN(n13356) );
  NOR2_X1 U15773 ( .A1(n13356), .A2(n13355), .ZN(n13357) );
  NAND3_X1 U15774 ( .A1(n13363), .A2(n13362), .A3(n13358), .ZN(n13360) );
  NAND3_X1 U15775 ( .A1(n13360), .A2(n13359), .A3(n13365), .ZN(n13369) );
  NAND3_X1 U15776 ( .A1(n13363), .A2(n13362), .A3(n13361), .ZN(n13367) );
  AND2_X1 U15777 ( .A1(n13372), .A2(n13364), .ZN(n13366) );
  AOI21_X1 U15778 ( .B1(n13367), .B2(n13366), .A(n7565), .ZN(n13368) );
  MUX2_X1 U15779 ( .A(n13369), .B(n13368), .S(n13450), .Z(n13371) );
  OAI211_X1 U15780 ( .C1(n13372), .C2(n13450), .A(n13371), .B(n13370), .ZN(
        n13377) );
  MUX2_X1 U15781 ( .A(n13375), .B(n13374), .S(n13450), .Z(n13376) );
  NAND3_X1 U15782 ( .A1(n13377), .A2(n7251), .A3(n13376), .ZN(n13382) );
  MUX2_X1 U15783 ( .A(n13379), .B(n13378), .S(n13468), .Z(n13380) );
  NAND3_X1 U15784 ( .A1(n13382), .A2(n13381), .A3(n13380), .ZN(n13386) );
  MUX2_X1 U15785 ( .A(n7556), .B(n13384), .S(n13468), .Z(n13385) );
  MUX2_X1 U15786 ( .A(n13388), .B(n13387), .S(n13450), .Z(n13389) );
  NAND2_X1 U15787 ( .A1(n13396), .A2(n13391), .ZN(n13394) );
  NAND2_X1 U15788 ( .A1(n13395), .A2(n13392), .ZN(n13393) );
  MUX2_X1 U15789 ( .A(n13394), .B(n13393), .S(n13468), .Z(n13399) );
  MUX2_X1 U15790 ( .A(n13396), .B(n13395), .S(n13450), .Z(n13397) );
  MUX2_X1 U15791 ( .A(n13401), .B(n13400), .S(n13468), .Z(n13403) );
  AND2_X1 U15792 ( .A1(n13404), .A2(n13499), .ZN(n13406) );
  MUX2_X1 U15793 ( .A(n13406), .B(n13405), .S(n13450), .Z(n13407) );
  OR3_X1 U15794 ( .A1(n13409), .A2(n13408), .A3(n13407), .ZN(n13413) );
  OAI21_X1 U15795 ( .B1(n13804), .B2(n13952), .A(n13410), .ZN(n13411) );
  INV_X1 U15796 ( .A(n13415), .ZN(n13412) );
  AOI21_X1 U15797 ( .B1(n13415), .B2(n13414), .A(n13450), .ZN(n13416) );
  INV_X1 U15798 ( .A(n13417), .ZN(n13418) );
  AOI21_X1 U15799 ( .B1(n13423), .B2(n13418), .A(n13450), .ZN(n13419) );
  NAND2_X1 U15800 ( .A1(n13420), .A2(n13419), .ZN(n13422) );
  INV_X1 U15801 ( .A(n13770), .ZN(n13426) );
  NAND2_X1 U15802 ( .A1(n13423), .A2(n13450), .ZN(n13424) );
  MUX2_X1 U15803 ( .A(n13428), .B(n13427), .S(n13468), .Z(n13429) );
  NAND3_X1 U15804 ( .A1(n13430), .A2(n13745), .A3(n13429), .ZN(n13434) );
  MUX2_X1 U15805 ( .A(n13432), .B(n13431), .S(n13468), .Z(n13433) );
  NAND3_X1 U15806 ( .A1(n13434), .A2(n13731), .A3(n13433), .ZN(n13439) );
  MUX2_X1 U15807 ( .A(n13436), .B(n13435), .S(n13450), .Z(n13437) );
  NAND3_X1 U15808 ( .A1(n13439), .A2(n13438), .A3(n13437), .ZN(n13443) );
  MUX2_X1 U15809 ( .A(n13441), .B(n13440), .S(n13450), .Z(n13442) );
  NAND3_X1 U15810 ( .A1(n13443), .A2(n13704), .A3(n13442), .ZN(n13446) );
  NAND3_X1 U15811 ( .A1(n13850), .A2(n13444), .A3(n13468), .ZN(n13445) );
  NAND2_X1 U15812 ( .A1(n13446), .A2(n13445), .ZN(n13447) );
  NAND2_X1 U15813 ( .A1(n13448), .A2(n13450), .ZN(n13449) );
  MUX2_X1 U15814 ( .A(n13453), .B(n13452), .S(n13468), .Z(n13454) );
  MUX2_X1 U15815 ( .A(n13456), .B(n13455), .S(n13468), .Z(n13457) );
  NAND2_X1 U15816 ( .A1(n13459), .A2(n13458), .ZN(n13467) );
  INV_X1 U15817 ( .A(n13462), .ZN(n13463) );
  AOI21_X1 U15818 ( .B1(n13468), .B2(n13464), .A(n13463), .ZN(n13465) );
  NAND2_X1 U15819 ( .A1(n13466), .A2(n13465), .ZN(n13473) );
  INV_X1 U15820 ( .A(n13467), .ZN(n13470) );
  NAND3_X1 U15821 ( .A1(n13470), .A2(n13469), .A3(n13468), .ZN(n13471) );
  NAND3_X1 U15822 ( .A1(n13473), .A2(n13472), .A3(n13471), .ZN(n13476) );
  NAND3_X1 U15823 ( .A1(n13476), .A2(n13475), .A3(n7329), .ZN(n13478) );
  NOR3_X1 U15824 ( .A1(n13486), .A2(n13485), .A3(n8808), .ZN(n13489) );
  OAI21_X1 U15825 ( .B1(n13490), .B2(n13487), .A(P3_B_REG_SCAN_IN), .ZN(n13488) );
  MUX2_X1 U15826 ( .A(n13646), .B(P3_DATAO_REG_31__SCAN_IN), .S(n13510), .Z(
        P3_U3522) );
  MUX2_X1 U15827 ( .A(n13491), .B(P3_DATAO_REG_30__SCAN_IN), .S(n13510), .Z(
        P3_U3521) );
  MUX2_X1 U15828 ( .A(P3_DATAO_REG_29__SCAN_IN), .B(n13492), .S(P3_U3897), .Z(
        P3_U3520) );
  MUX2_X1 U15829 ( .A(P3_DATAO_REG_28__SCAN_IN), .B(n13493), .S(P3_U3897), .Z(
        P3_U3519) );
  MUX2_X1 U15830 ( .A(n13666), .B(P3_DATAO_REG_27__SCAN_IN), .S(n13510), .Z(
        P3_U3518) );
  MUX2_X1 U15831 ( .A(n13494), .B(P3_DATAO_REG_26__SCAN_IN), .S(n13510), .Z(
        P3_U3517) );
  MUX2_X1 U15832 ( .A(P3_DATAO_REG_25__SCAN_IN), .B(n6947), .S(P3_U3897), .Z(
        P3_U3516) );
  MUX2_X1 U15833 ( .A(P3_DATAO_REG_24__SCAN_IN), .B(n7128), .S(P3_U3897), .Z(
        P3_U3515) );
  MUX2_X1 U15834 ( .A(n13705), .B(P3_DATAO_REG_22__SCAN_IN), .S(n13510), .Z(
        P3_U3513) );
  MUX2_X1 U15835 ( .A(P3_DATAO_REG_21__SCAN_IN), .B(n13721), .S(P3_U3897), .Z(
        P3_U3512) );
  MUX2_X1 U15836 ( .A(P3_DATAO_REG_20__SCAN_IN), .B(n13495), .S(P3_U3897), .Z(
        P3_U3511) );
  MUX2_X1 U15837 ( .A(n13775), .B(P3_DATAO_REG_19__SCAN_IN), .S(n13510), .Z(
        P3_U3510) );
  MUX2_X1 U15838 ( .A(P3_DATAO_REG_18__SCAN_IN), .B(n13496), .S(P3_U3897), .Z(
        P3_U3509) );
  MUX2_X1 U15839 ( .A(P3_DATAO_REG_16__SCAN_IN), .B(n13497), .S(P3_U3897), .Z(
        P3_U3507) );
  MUX2_X1 U15840 ( .A(n13498), .B(P3_DATAO_REG_15__SCAN_IN), .S(n13510), .Z(
        P3_U3506) );
  MUX2_X1 U15841 ( .A(P3_DATAO_REG_14__SCAN_IN), .B(n13499), .S(P3_U3897), .Z(
        P3_U3505) );
  MUX2_X1 U15842 ( .A(n13500), .B(P3_DATAO_REG_13__SCAN_IN), .S(n13510), .Z(
        P3_U3504) );
  MUX2_X1 U15843 ( .A(P3_DATAO_REG_12__SCAN_IN), .B(n13501), .S(P3_U3897), .Z(
        P3_U3503) );
  MUX2_X1 U15844 ( .A(n13502), .B(P3_DATAO_REG_11__SCAN_IN), .S(n13510), .Z(
        P3_U3502) );
  MUX2_X1 U15845 ( .A(n13503), .B(P3_DATAO_REG_10__SCAN_IN), .S(n13510), .Z(
        P3_U3501) );
  MUX2_X1 U15846 ( .A(n13504), .B(P3_DATAO_REG_9__SCAN_IN), .S(n13510), .Z(
        P3_U3500) );
  MUX2_X1 U15847 ( .A(n13505), .B(P3_DATAO_REG_8__SCAN_IN), .S(n13510), .Z(
        P3_U3499) );
  MUX2_X1 U15848 ( .A(n13506), .B(P3_DATAO_REG_7__SCAN_IN), .S(n13510), .Z(
        P3_U3498) );
  MUX2_X1 U15849 ( .A(n13507), .B(P3_DATAO_REG_6__SCAN_IN), .S(n13510), .Z(
        P3_U3497) );
  MUX2_X1 U15850 ( .A(n13508), .B(P3_DATAO_REG_5__SCAN_IN), .S(n13510), .Z(
        P3_U3496) );
  MUX2_X1 U15851 ( .A(n13509), .B(P3_DATAO_REG_4__SCAN_IN), .S(n13510), .Z(
        P3_U3495) );
  MUX2_X1 U15852 ( .A(n16031), .B(P3_DATAO_REG_3__SCAN_IN), .S(n13510), .Z(
        P3_U3494) );
  MUX2_X1 U15853 ( .A(n16047), .B(P3_DATAO_REG_2__SCAN_IN), .S(n13510), .Z(
        P3_U3493) );
  MUX2_X1 U15854 ( .A(n16048), .B(P3_DATAO_REG_0__SCAN_IN), .S(n13510), .Z(
        P3_U3491) );
  OAI21_X1 U15855 ( .B1(n13513), .B2(n13512), .A(n13511), .ZN(n13514) );
  NAND2_X1 U15856 ( .A1(n13514), .A2(n13583), .ZN(n13529) );
  OAI21_X1 U15857 ( .B1(n16024), .B2(n13517), .A(n13516), .ZN(n13522) );
  INV_X1 U15858 ( .A(n13536), .ZN(n13518) );
  AOI211_X1 U15859 ( .C1(n13520), .C2(n13519), .A(n16013), .B(n13518), .ZN(
        n13521) );
  AOI211_X1 U15860 ( .C1(n16021), .C2(n6904), .A(n13522), .B(n13521), .ZN(
        n13528) );
  AND3_X1 U15861 ( .A1(n13525), .A2(n13524), .A3(n13523), .ZN(n13526) );
  NAND3_X1 U15862 ( .A1(n13529), .A2(n13528), .A3(n13527), .ZN(P3_U3194) );
  INV_X1 U15863 ( .A(n13552), .ZN(n13530) );
  AOI21_X1 U15864 ( .B1(n13532), .B2(n13531), .A(n13530), .ZN(n13547) );
  OAI21_X1 U15865 ( .B1(P3_REG1_REG_13__SCAN_IN), .B2(n13533), .A(n6906), .ZN(
        n13545) );
  INV_X1 U15866 ( .A(n13558), .ZN(n13539) );
  AOI21_X1 U15867 ( .B1(n13536), .B2(n13535), .A(n13534), .ZN(n13538) );
  OAI21_X1 U15868 ( .B1(n13539), .B2(n13538), .A(n13537), .ZN(n13542) );
  AOI21_X1 U15869 ( .B1(n16012), .B2(P3_ADDR_REG_13__SCAN_IN), .A(n13540), 
        .ZN(n13541) );
  OAI211_X1 U15870 ( .C1(n13617), .C2(n13543), .A(n13542), .B(n13541), .ZN(
        n13544) );
  AOI21_X1 U15871 ( .B1(n13545), .B2(n13631), .A(n13544), .ZN(n13546) );
  OAI21_X1 U15872 ( .B1(n13547), .B2(n16014), .A(n13546), .ZN(P3_U3195) );
  INV_X1 U15873 ( .A(n13548), .ZN(n13550) );
  NOR2_X1 U15874 ( .A1(n13550), .A2(n13549), .ZN(n13553) );
  AOI21_X1 U15875 ( .B1(n13553), .B2(n13552), .A(n13551), .ZN(n13571) );
  INV_X1 U15876 ( .A(P3_ADDR_REG_14__SCAN_IN), .ZN(n13555) );
  OAI21_X1 U15877 ( .B1(n16024), .B2(n13555), .A(n13554), .ZN(n13561) );
  AOI21_X1 U15878 ( .B1(n13558), .B2(n13557), .A(n13556), .ZN(n13559) );
  NOR3_X1 U15879 ( .A1(n6716), .A2(n13559), .A3(n16013), .ZN(n13560) );
  AOI211_X1 U15880 ( .C1(n16021), .C2(n13562), .A(n13561), .B(n13560), .ZN(
        n13570) );
  INV_X1 U15881 ( .A(n13563), .ZN(n13568) );
  NOR3_X1 U15882 ( .A1(n13566), .A2(n13565), .A3(n13564), .ZN(n13567) );
  OAI21_X1 U15883 ( .B1(n13568), .B2(n13567), .A(n13631), .ZN(n13569) );
  OAI211_X1 U15884 ( .C1(n13571), .C2(n16014), .A(n13570), .B(n13569), .ZN(
        P3_U3196) );
  AOI21_X1 U15885 ( .B1(n13879), .B2(n13573), .A(n13572), .ZN(n13587) );
  INV_X1 U15886 ( .A(P3_ADDR_REG_15__SCAN_IN), .ZN(n13575) );
  OAI21_X1 U15887 ( .B1(n16024), .B2(n13575), .A(n13574), .ZN(n13581) );
  AOI21_X1 U15888 ( .B1(n13578), .B2(n13577), .A(n13576), .ZN(n13579) );
  NOR2_X1 U15889 ( .A1(n13579), .A2(n16013), .ZN(n13580) );
  AOI211_X1 U15890 ( .C1(n16021), .C2(n13582), .A(n13581), .B(n13580), .ZN(
        n13586) );
  OAI21_X1 U15891 ( .B1(n6694), .B2(P3_REG2_REG_15__SCAN_IN), .A(n13591), .ZN(
        n13584) );
  NAND2_X1 U15892 ( .A1(n13584), .A2(n13583), .ZN(n13585) );
  OAI211_X1 U15893 ( .C1(n13587), .C2(n16015), .A(n13586), .B(n13585), .ZN(
        P3_U3197) );
  NOR2_X1 U15894 ( .A1(n6991), .A2(n13589), .ZN(n13592) );
  AOI21_X1 U15895 ( .B1(n13592), .B2(n13591), .A(n6555), .ZN(n13609) );
  INV_X1 U15896 ( .A(P3_ADDR_REG_16__SCAN_IN), .ZN(n15735) );
  OAI21_X1 U15897 ( .B1(n16024), .B2(n15735), .A(n13593), .ZN(n13600) );
  NOR2_X1 U15898 ( .A1(n13595), .A2(n7434), .ZN(n13596) );
  XNOR2_X1 U15899 ( .A(n13597), .B(n13596), .ZN(n13598) );
  NOR2_X1 U15900 ( .A1(n13598), .A2(n16013), .ZN(n13599) );
  AOI211_X1 U15901 ( .C1(n16021), .C2(n13601), .A(n13600), .B(n13599), .ZN(
        n13608) );
  INV_X1 U15902 ( .A(n13602), .ZN(n13606) );
  NOR3_X1 U15903 ( .A1(n13572), .A2(n13604), .A3(n13603), .ZN(n13605) );
  OAI21_X1 U15904 ( .B1(n13606), .B2(n13605), .A(n13631), .ZN(n13607) );
  OAI211_X1 U15905 ( .C1(n13609), .C2(n16014), .A(n13608), .B(n13607), .ZN(
        P3_U3198) );
  INV_X1 U15906 ( .A(n13625), .ZN(n13610) );
  AOI21_X1 U15907 ( .B1(n7652), .B2(n13611), .A(n13610), .ZN(n13622) );
  AOI211_X1 U15908 ( .C1(n13613), .C2(n13612), .A(n16013), .B(n6653), .ZN(
        n13619) );
  NAND2_X1 U15909 ( .A1(n16012), .A2(P3_ADDR_REG_17__SCAN_IN), .ZN(n13614) );
  OAI211_X1 U15910 ( .C1(n13617), .C2(n13616), .A(n13615), .B(n13614), .ZN(
        n13618) );
  AOI211_X1 U15911 ( .C1(n13620), .C2(n13631), .A(n13619), .B(n13618), .ZN(
        n13621) );
  OAI21_X1 U15912 ( .B1(n13622), .B2(n16014), .A(n13621), .ZN(P3_U3199) );
  AND3_X1 U15913 ( .A1(n13630), .A2(n13629), .A3(n13628), .ZN(n13632) );
  OAI21_X1 U15914 ( .B1(n13633), .B2(n13632), .A(n13631), .ZN(n13643) );
  INV_X1 U15915 ( .A(P3_ADDR_REG_18__SCAN_IN), .ZN(n15759) );
  OAI21_X1 U15916 ( .B1(n16024), .B2(n15759), .A(n13634), .ZN(n13640) );
  AOI21_X1 U15917 ( .B1(n13637), .B2(n13636), .A(n13635), .ZN(n13638) );
  NOR2_X1 U15918 ( .A1(n13638), .A2(n16013), .ZN(n13639) );
  AOI211_X1 U15919 ( .C1(n16021), .C2(n13641), .A(n13640), .B(n13639), .ZN(
        n13642) );
  OAI211_X1 U15920 ( .C1(n13644), .C2(n16014), .A(n13643), .B(n13642), .ZN(
        P3_U3200) );
  NAND2_X1 U15921 ( .A1(n13825), .A2(n13814), .ZN(n13648) );
  AOI21_X1 U15922 ( .B1(n13888), .B2(n9401), .A(n13647), .ZN(n13651) );
  OAI211_X1 U15923 ( .C1(n13649), .C2(n9401), .A(n13648), .B(n13651), .ZN(
        P3_U3202) );
  NAND2_X1 U15924 ( .A1(n16066), .A2(P3_REG2_REG_30__SCAN_IN), .ZN(n13650) );
  OAI211_X1 U15925 ( .C1(n13893), .C2(n13737), .A(n13651), .B(n13650), .ZN(
        P3_U3203) );
  AOI22_X1 U15926 ( .A1(n13652), .A2(n16061), .B1(n16066), .B2(
        P3_REG2_REG_28__SCAN_IN), .ZN(n13653) );
  OAI21_X1 U15927 ( .B1(n13832), .B2(n13737), .A(n13653), .ZN(n13654) );
  AOI21_X1 U15928 ( .B1(n13655), .B2(n9427), .A(n13654), .ZN(n13656) );
  OAI21_X1 U15929 ( .B1(n16066), .B2(n6663), .A(n13656), .ZN(P3_U3205) );
  INV_X1 U15930 ( .A(n13657), .ZN(n13663) );
  AOI22_X1 U15931 ( .A1(n13658), .A2(n16061), .B1(n16066), .B2(
        P3_REG2_REG_27__SCAN_IN), .ZN(n13659) );
  OAI21_X1 U15932 ( .B1(n13835), .B2(n13737), .A(n13659), .ZN(n13660) );
  AOI21_X1 U15933 ( .B1(n13661), .B2(n16062), .A(n13660), .ZN(n13662) );
  OAI21_X1 U15934 ( .B1(n13663), .B2(n16066), .A(n13662), .ZN(P3_U3206) );
  XNOR2_X1 U15935 ( .A(n13664), .B(n13665), .ZN(n13667) );
  AOI222_X1 U15936 ( .A1(n6947), .A2(n16049), .B1(n16044), .B2(n13667), .C1(
        n13666), .C2(n16046), .ZN(n13838) );
  XNOR2_X1 U15937 ( .A(n13668), .B(n13669), .ZN(n13837) );
  INV_X1 U15938 ( .A(n13836), .ZN(n13672) );
  AOI22_X1 U15939 ( .A1(n13670), .A2(n16061), .B1(n16066), .B2(
        P3_REG2_REG_26__SCAN_IN), .ZN(n13671) );
  OAI21_X1 U15940 ( .B1(n13672), .B2(n13737), .A(n13671), .ZN(n13673) );
  AOI21_X1 U15941 ( .B1(n13837), .B2(n9427), .A(n13673), .ZN(n13674) );
  OAI21_X1 U15942 ( .B1(n16066), .B2(n13838), .A(n13674), .ZN(P3_U3207) );
  AND2_X1 U15943 ( .A1(n13708), .A2(n13675), .ZN(n13694) );
  NAND2_X1 U15944 ( .A1(n13694), .A2(n13696), .ZN(n13693) );
  NAND2_X1 U15945 ( .A1(n13693), .A2(n13676), .ZN(n13678) );
  XNOR2_X1 U15946 ( .A(n13678), .B(n13677), .ZN(n13898) );
  NAND2_X1 U15947 ( .A1(n13680), .A2(n13679), .ZN(n13681) );
  NAND3_X1 U15948 ( .A1(n13682), .A2(n16044), .A3(n13681), .ZN(n13687) );
  OAI22_X1 U15949 ( .A1(n13684), .A2(n13817), .B1(n13683), .B2(n13815), .ZN(
        n13685) );
  INV_X1 U15950 ( .A(n13685), .ZN(n13686) );
  NAND2_X1 U15951 ( .A1(n13687), .A2(n13686), .ZN(n13840) );
  NAND2_X1 U15952 ( .A1(n13841), .A2(n13814), .ZN(n13690) );
  AOI22_X1 U15953 ( .A1(n13688), .A2(n16061), .B1(n16066), .B2(
        P3_REG2_REG_25__SCAN_IN), .ZN(n13689) );
  NAND2_X1 U15954 ( .A1(n13690), .A2(n13689), .ZN(n13691) );
  AOI21_X1 U15955 ( .B1(n13840), .B2(n9401), .A(n13691), .ZN(n13692) );
  OAI21_X1 U15956 ( .B1(n13898), .B2(n13824), .A(n13692), .ZN(P3_U3208) );
  OAI21_X1 U15957 ( .B1(n13694), .B2(n13696), .A(n13693), .ZN(n13900) );
  INV_X1 U15958 ( .A(n13900), .ZN(n13702) );
  AOI22_X1 U15959 ( .A1(n13899), .A2(n13814), .B1(n16061), .B2(n13695), .ZN(
        n13701) );
  XNOR2_X1 U15960 ( .A(n13697), .B(n13696), .ZN(n13698) );
  AOI222_X1 U15961 ( .A1(n13722), .A2(n16049), .B1(n16044), .B2(n13698), .C1(
        n6947), .C2(n16046), .ZN(n13901) );
  MUX2_X1 U15962 ( .A(n13699), .B(n13901), .S(n9401), .Z(n13700) );
  OAI211_X1 U15963 ( .C1(n13702), .C2(n13824), .A(n13701), .B(n13700), .ZN(
        P3_U3209) );
  XNOR2_X1 U15964 ( .A(n13703), .B(n13704), .ZN(n13706) );
  AOI222_X1 U15965 ( .A1(n13706), .A2(n16044), .B1(n7128), .B2(n16046), .C1(
        n13705), .C2(n16049), .ZN(n13848) );
  INV_X1 U15966 ( .A(n13707), .ZN(n13711) );
  INV_X1 U15967 ( .A(n13708), .ZN(n13709) );
  AOI21_X1 U15968 ( .B1(n13711), .B2(n13710), .A(n13709), .ZN(n13847) );
  INV_X1 U15969 ( .A(n13850), .ZN(n13714) );
  AOI22_X1 U15970 ( .A1(n13712), .A2(n16061), .B1(n16066), .B2(
        P3_REG2_REG_23__SCAN_IN), .ZN(n13713) );
  OAI21_X1 U15971 ( .B1(n13714), .B2(n13737), .A(n13713), .ZN(n13715) );
  AOI21_X1 U15972 ( .B1(n13847), .B2(n9427), .A(n13715), .ZN(n13716) );
  OAI21_X1 U15973 ( .B1(n16066), .B2(n13848), .A(n13716), .ZN(P3_U3210) );
  XNOR2_X1 U15974 ( .A(n13717), .B(n13720), .ZN(n13914) );
  AOI22_X1 U15975 ( .A1(n13911), .A2(n13814), .B1(n16061), .B2(n13718), .ZN(
        n13726) );
  INV_X1 U15976 ( .A(P3_REG2_REG_22__SCAN_IN), .ZN(n13724) );
  XNOR2_X1 U15977 ( .A(n13719), .B(n13720), .ZN(n13723) );
  AOI222_X1 U15978 ( .A1(n13723), .A2(n16044), .B1(n13722), .B2(n16046), .C1(
        n13721), .C2(n16049), .ZN(n13909) );
  MUX2_X1 U15979 ( .A(n13724), .B(n13909), .S(n9401), .Z(n13725) );
  OAI211_X1 U15980 ( .C1(n13914), .C2(n13824), .A(n13726), .B(n13725), .ZN(
        P3_U3211) );
  XNOR2_X1 U15981 ( .A(n13727), .B(n9236), .ZN(n13857) );
  INV_X1 U15982 ( .A(n13857), .ZN(n13740) );
  INV_X1 U15983 ( .A(n13728), .ZN(n13729) );
  AOI21_X1 U15984 ( .B1(n13731), .B2(n13730), .A(n13729), .ZN(n13732) );
  OAI222_X1 U15985 ( .A1(n13817), .A2(n13733), .B1(n13815), .B2(n13761), .C1(
        n13732), .C2(n16034), .ZN(n13856) );
  INV_X1 U15986 ( .A(n13734), .ZN(n13919) );
  AOI22_X1 U15987 ( .A1(n13735), .A2(n16061), .B1(n16066), .B2(
        P3_REG2_REG_21__SCAN_IN), .ZN(n13736) );
  OAI21_X1 U15988 ( .B1(n13919), .B2(n13737), .A(n13736), .ZN(n13738) );
  AOI21_X1 U15989 ( .B1(n13856), .B2(n9401), .A(n13738), .ZN(n13739) );
  OAI21_X1 U15990 ( .B1(n13740), .B2(n13824), .A(n13739), .ZN(P3_U3212) );
  OAI21_X1 U15991 ( .B1(n13742), .B2(n13745), .A(n13741), .ZN(n13925) );
  AOI22_X1 U15992 ( .A1(n13922), .A2(n13814), .B1(n16061), .B2(n13743), .ZN(
        n13754) );
  INV_X1 U15993 ( .A(P3_REG2_REG_20__SCAN_IN), .ZN(n13752) );
  INV_X1 U15994 ( .A(n13744), .ZN(n13746) );
  AOI21_X1 U15995 ( .B1(n13746), .B2(n13745), .A(n16034), .ZN(n13751) );
  OAI22_X1 U15996 ( .A1(n13749), .A2(n13817), .B1(n13748), .B2(n13815), .ZN(
        n13750) );
  AOI21_X1 U15997 ( .B1(n13751), .B2(n6559), .A(n13750), .ZN(n13920) );
  MUX2_X1 U15998 ( .A(n13752), .B(n13920), .S(n9401), .Z(n13753) );
  OAI211_X1 U15999 ( .C1(n13925), .C2(n13824), .A(n13754), .B(n13753), .ZN(
        P3_U3213) );
  NAND2_X1 U16000 ( .A1(n13767), .A2(n13755), .ZN(n13756) );
  XNOR2_X1 U16001 ( .A(n13756), .B(n13758), .ZN(n13931) );
  AOI22_X1 U16002 ( .A1(n13929), .A2(n13814), .B1(n16061), .B2(n13757), .ZN(
        n13766) );
  INV_X1 U16003 ( .A(P3_REG2_REG_19__SCAN_IN), .ZN(n13764) );
  AOI21_X1 U16004 ( .B1(n13759), .B2(n13758), .A(n16034), .ZN(n13763) );
  OAI22_X1 U16005 ( .A1(n13761), .A2(n13817), .B1(n13791), .B2(n13815), .ZN(
        n13762) );
  AOI21_X1 U16006 ( .B1(n13763), .B2(n13760), .A(n13762), .ZN(n13926) );
  MUX2_X1 U16007 ( .A(n13764), .B(n13926), .S(n9401), .Z(n13765) );
  OAI211_X1 U16008 ( .C1(n13931), .C2(n13824), .A(n13766), .B(n13765), .ZN(
        P3_U3214) );
  OAI21_X1 U16009 ( .B1(n13768), .B2(n13770), .A(n13767), .ZN(n13935) );
  NAND2_X1 U16010 ( .A1(n13771), .A2(n13770), .ZN(n13772) );
  NAND2_X1 U16011 ( .A1(n13769), .A2(n13772), .ZN(n13773) );
  NAND2_X1 U16012 ( .A1(n13773), .A2(n16044), .ZN(n13777) );
  AOI22_X1 U16013 ( .A1(n13775), .A2(n16046), .B1(n16049), .B2(n13774), .ZN(
        n13776) );
  NAND2_X1 U16014 ( .A1(n13777), .A2(n13776), .ZN(n13867) );
  NAND2_X1 U16015 ( .A1(n13868), .A2(n13814), .ZN(n13780) );
  AOI22_X1 U16016 ( .A1(n16066), .A2(P3_REG2_REG_18__SCAN_IN), .B1(n16061), 
        .B2(n13778), .ZN(n13779) );
  NAND2_X1 U16017 ( .A1(n13780), .A2(n13779), .ZN(n13781) );
  AOI21_X1 U16018 ( .B1(n13867), .B2(n9401), .A(n13781), .ZN(n13782) );
  OAI21_X1 U16019 ( .B1(n13935), .B2(n13824), .A(n13782), .ZN(P3_U3215) );
  XNOR2_X1 U16020 ( .A(n13784), .B(n13783), .ZN(n13941) );
  AOI22_X1 U16021 ( .A1(n13939), .A2(n13814), .B1(n16061), .B2(n13785), .ZN(
        n13795) );
  NAND3_X1 U16022 ( .A1(n13786), .A2(n13788), .A3(n13787), .ZN(n13789) );
  AND3_X1 U16023 ( .A1(n13790), .A2(n16044), .A3(n13789), .ZN(n13793) );
  OAI22_X1 U16024 ( .A1(n13791), .A2(n13817), .B1(n13818), .B2(n13815), .ZN(
        n13792) );
  NOR2_X1 U16025 ( .A1(n13793), .A2(n13792), .ZN(n13936) );
  MUX2_X1 U16026 ( .A(n7652), .B(n13936), .S(n9401), .Z(n13794) );
  OAI211_X1 U16027 ( .C1(n13941), .C2(n13824), .A(n13795), .B(n13794), .ZN(
        P3_U3216) );
  OAI21_X1 U16028 ( .B1(n13798), .B2(n13797), .A(n13796), .ZN(n13944) );
  INV_X1 U16029 ( .A(n13944), .ZN(n13811) );
  AOI22_X1 U16030 ( .A1(n13942), .A2(n13814), .B1(n16061), .B2(n13799), .ZN(
        n13810) );
  NOR2_X1 U16031 ( .A1(n13802), .A2(n7040), .ZN(n13803) );
  AOI21_X1 U16032 ( .B1(n13800), .B2(n13803), .A(n16034), .ZN(n13807) );
  OAI22_X1 U16033 ( .A1(n13805), .A2(n13817), .B1(n13804), .B2(n13815), .ZN(
        n13806) );
  AOI21_X1 U16034 ( .B1(n13786), .B2(n13807), .A(n13806), .ZN(n13945) );
  MUX2_X1 U16035 ( .A(n13808), .B(n13945), .S(n9401), .Z(n13809) );
  OAI211_X1 U16036 ( .C1(n13811), .C2(n13824), .A(n13810), .B(n13809), .ZN(
        P3_U3217) );
  XNOR2_X1 U16037 ( .A(n13812), .B(n7547), .ZN(n13956) );
  AOI22_X1 U16038 ( .A1(n13952), .A2(n13814), .B1(n16061), .B2(n13813), .ZN(
        n13823) );
  AOI21_X1 U16039 ( .B1(n6587), .B2(n7547), .A(n16034), .ZN(n13820) );
  OAI22_X1 U16040 ( .A1(n13818), .A2(n13817), .B1(n13816), .B2(n13815), .ZN(
        n13819) );
  AOI21_X1 U16041 ( .B1(n13820), .B2(n13800), .A(n13819), .ZN(n13949) );
  MUX2_X1 U16042 ( .A(n13821), .B(n13949), .S(n9401), .Z(n13822) );
  OAI211_X1 U16043 ( .C1(n13956), .C2(n13824), .A(n13823), .B(n13822), .ZN(
        P3_U3218) );
  NAND2_X1 U16044 ( .A1(n13825), .A2(n13880), .ZN(n13826) );
  NAND2_X1 U16045 ( .A1(n13888), .A2(n16106), .ZN(n13829) );
  OAI211_X1 U16046 ( .C1(n16106), .C2(n13827), .A(n13826), .B(n13829), .ZN(
        P3_U3490) );
  NAND2_X1 U16047 ( .A1(n16103), .A2(P3_REG1_REG_30__SCAN_IN), .ZN(n13828) );
  OAI211_X1 U16048 ( .C1(n13893), .C2(n13860), .A(n13829), .B(n13828), .ZN(
        P3_U3489) );
  OAI21_X1 U16049 ( .B1(n13832), .B2(n13860), .A(n13831), .ZN(P3_U3487) );
  AOI22_X1 U16050 ( .A1(n13837), .A2(n16070), .B1(n13869), .B2(n13836), .ZN(
        n13839) );
  NAND2_X1 U16051 ( .A1(n13839), .A2(n13838), .ZN(n13894) );
  MUX2_X1 U16052 ( .A(P3_REG1_REG_26__SCAN_IN), .B(n13894), .S(n16106), .Z(
        P3_U3485) );
  AOI21_X1 U16053 ( .B1(n13869), .B2(n13841), .A(n13840), .ZN(n13895) );
  MUX2_X1 U16054 ( .A(n13842), .B(n13895), .S(n16106), .Z(n13843) );
  OAI21_X1 U16055 ( .B1(n13898), .B2(n13883), .A(n13843), .ZN(P3_U3484) );
  AOI22_X1 U16056 ( .A1(n13900), .A2(n13875), .B1(n13880), .B2(n13899), .ZN(
        n13846) );
  MUX2_X1 U16057 ( .A(n13844), .B(n13901), .S(n16106), .Z(n13845) );
  NAND2_X1 U16058 ( .A1(n13846), .A2(n13845), .ZN(P3_U3483) );
  INV_X1 U16059 ( .A(n13847), .ZN(n13908) );
  INV_X1 U16060 ( .A(n13848), .ZN(n13849) );
  AOI21_X1 U16061 ( .B1(n13869), .B2(n13850), .A(n13849), .ZN(n13905) );
  MUX2_X1 U16062 ( .A(n13851), .B(n13905), .S(n16106), .Z(n13852) );
  OAI21_X1 U16063 ( .B1(n13908), .B2(n13883), .A(n13852), .ZN(P3_U3482) );
  MUX2_X1 U16064 ( .A(n13853), .B(n13909), .S(n16106), .Z(n13855) );
  NAND2_X1 U16065 ( .A1(n13911), .A2(n13880), .ZN(n13854) );
  OAI211_X1 U16066 ( .C1(n13914), .C2(n13883), .A(n13855), .B(n13854), .ZN(
        P3_U3481) );
  AOI21_X1 U16067 ( .B1(n13857), .B2(n16070), .A(n13856), .ZN(n13915) );
  MUX2_X1 U16068 ( .A(n13858), .B(n13915), .S(n16106), .Z(n13859) );
  OAI21_X1 U16069 ( .B1(n13919), .B2(n13860), .A(n13859), .ZN(P3_U3480) );
  MUX2_X1 U16070 ( .A(n13861), .B(n13920), .S(n16106), .Z(n13863) );
  NAND2_X1 U16071 ( .A1(n13922), .A2(n13880), .ZN(n13862) );
  OAI211_X1 U16072 ( .C1(n13925), .C2(n13883), .A(n13863), .B(n13862), .ZN(
        P3_U3479) );
  MUX2_X1 U16073 ( .A(n13864), .B(n13926), .S(n16106), .Z(n13866) );
  NAND2_X1 U16074 ( .A1(n13929), .A2(n13880), .ZN(n13865) );
  OAI211_X1 U16075 ( .C1(n13931), .C2(n13883), .A(n13866), .B(n13865), .ZN(
        P3_U3478) );
  AOI21_X1 U16076 ( .B1(n13869), .B2(n13868), .A(n13867), .ZN(n13932) );
  MUX2_X1 U16077 ( .A(n13870), .B(n13932), .S(n16106), .Z(n13871) );
  OAI21_X1 U16078 ( .B1(n13935), .B2(n13883), .A(n13871), .ZN(P3_U3477) );
  MUX2_X1 U16079 ( .A(n13872), .B(n13936), .S(n16106), .Z(n13874) );
  NAND2_X1 U16080 ( .A1(n13939), .A2(n13880), .ZN(n13873) );
  OAI211_X1 U16081 ( .C1(n13941), .C2(n13883), .A(n13874), .B(n13873), .ZN(
        P3_U3476) );
  AOI22_X1 U16082 ( .A1(n13944), .A2(n13875), .B1(n13880), .B2(n13942), .ZN(
        n13878) );
  MUX2_X1 U16083 ( .A(n13876), .B(n13945), .S(n16106), .Z(n13877) );
  NAND2_X1 U16084 ( .A1(n13878), .A2(n13877), .ZN(P3_U3475) );
  MUX2_X1 U16085 ( .A(n13879), .B(n13949), .S(n16106), .Z(n13882) );
  NAND2_X1 U16086 ( .A1(n13952), .A2(n13880), .ZN(n13881) );
  OAI211_X1 U16087 ( .C1(n13956), .C2(n13883), .A(n13882), .B(n13881), .ZN(
        P3_U3474) );
  NAND2_X1 U16088 ( .A1(n13884), .A2(n16070), .ZN(n13886) );
  OAI211_X1 U16089 ( .C1(n16055), .C2(n13887), .A(n13886), .B(n13885), .ZN(
        n13957) );
  MUX2_X1 U16090 ( .A(P3_REG1_REG_9__SCAN_IN), .B(n13957), .S(n16106), .Z(
        P3_U3468) );
  NAND2_X1 U16091 ( .A1(n16092), .A2(P3_REG0_REG_31__SCAN_IN), .ZN(n13889) );
  NAND2_X1 U16092 ( .A1(n13888), .A2(n16094), .ZN(n13892) );
  OAI211_X1 U16093 ( .C1(n13890), .C2(n13918), .A(n13889), .B(n13892), .ZN(
        P3_U3458) );
  NAND2_X1 U16094 ( .A1(n16092), .A2(P3_REG0_REG_30__SCAN_IN), .ZN(n13891) );
  OAI211_X1 U16095 ( .C1(n13893), .C2(n13918), .A(n13892), .B(n13891), .ZN(
        P3_U3457) );
  MUX2_X1 U16096 ( .A(P3_REG0_REG_26__SCAN_IN), .B(n13894), .S(n16094), .Z(
        P3_U3453) );
  INV_X1 U16097 ( .A(P3_REG0_REG_25__SCAN_IN), .ZN(n13896) );
  MUX2_X1 U16098 ( .A(n13896), .B(n13895), .S(n16094), .Z(n13897) );
  OAI21_X1 U16099 ( .B1(n13898), .B2(n13955), .A(n13897), .ZN(P3_U3452) );
  AOI22_X1 U16100 ( .A1(n13900), .A2(n13943), .B1(n13953), .B2(n13899), .ZN(
        n13904) );
  INV_X1 U16101 ( .A(P3_REG0_REG_24__SCAN_IN), .ZN(n13902) );
  MUX2_X1 U16102 ( .A(n13902), .B(n13901), .S(n16094), .Z(n13903) );
  NAND2_X1 U16103 ( .A1(n13904), .A2(n13903), .ZN(P3_U3451) );
  MUX2_X1 U16104 ( .A(n13906), .B(n13905), .S(n16094), .Z(n13907) );
  OAI21_X1 U16105 ( .B1(n13908), .B2(n13955), .A(n13907), .ZN(P3_U3450) );
  INV_X1 U16106 ( .A(P3_REG0_REG_22__SCAN_IN), .ZN(n13910) );
  MUX2_X1 U16107 ( .A(n13910), .B(n13909), .S(n16094), .Z(n13913) );
  NAND2_X1 U16108 ( .A1(n13911), .A2(n13953), .ZN(n13912) );
  OAI211_X1 U16109 ( .C1(n13914), .C2(n13955), .A(n13913), .B(n13912), .ZN(
        P3_U3449) );
  INV_X1 U16110 ( .A(P3_REG0_REG_21__SCAN_IN), .ZN(n13916) );
  MUX2_X1 U16111 ( .A(n13916), .B(n13915), .S(n16094), .Z(n13917) );
  OAI21_X1 U16112 ( .B1(n13919), .B2(n13918), .A(n13917), .ZN(P3_U3448) );
  INV_X1 U16113 ( .A(P3_REG0_REG_20__SCAN_IN), .ZN(n13921) );
  MUX2_X1 U16114 ( .A(n13921), .B(n13920), .S(n16094), .Z(n13924) );
  NAND2_X1 U16115 ( .A1(n13922), .A2(n13953), .ZN(n13923) );
  OAI211_X1 U16116 ( .C1(n13925), .C2(n13955), .A(n13924), .B(n13923), .ZN(
        P3_U3447) );
  INV_X1 U16117 ( .A(n13926), .ZN(n13927) );
  MUX2_X1 U16118 ( .A(P3_REG0_REG_19__SCAN_IN), .B(n13927), .S(n16094), .Z(
        n13928) );
  AOI21_X1 U16119 ( .B1(n13953), .B2(n13929), .A(n13928), .ZN(n13930) );
  OAI21_X1 U16120 ( .B1(n13931), .B2(n13955), .A(n13930), .ZN(P3_U3446) );
  INV_X1 U16121 ( .A(P3_REG0_REG_18__SCAN_IN), .ZN(n13933) );
  MUX2_X1 U16122 ( .A(n13933), .B(n13932), .S(n16094), .Z(n13934) );
  OAI21_X1 U16123 ( .B1(n13935), .B2(n13955), .A(n13934), .ZN(P3_U3444) );
  INV_X1 U16124 ( .A(n13936), .ZN(n13937) );
  MUX2_X1 U16125 ( .A(P3_REG0_REG_17__SCAN_IN), .B(n13937), .S(n16094), .Z(
        n13938) );
  AOI21_X1 U16126 ( .B1(n13953), .B2(n13939), .A(n13938), .ZN(n13940) );
  OAI21_X1 U16127 ( .B1(n13941), .B2(n13955), .A(n13940), .ZN(P3_U3441) );
  AOI22_X1 U16128 ( .A1(n13944), .A2(n13943), .B1(n13953), .B2(n13942), .ZN(
        n13948) );
  INV_X1 U16129 ( .A(P3_REG0_REG_16__SCAN_IN), .ZN(n13946) );
  MUX2_X1 U16130 ( .A(n13946), .B(n13945), .S(n16094), .Z(n13947) );
  NAND2_X1 U16131 ( .A1(n13948), .A2(n13947), .ZN(P3_U3438) );
  INV_X1 U16132 ( .A(n13949), .ZN(n13950) );
  MUX2_X1 U16133 ( .A(P3_REG0_REG_15__SCAN_IN), .B(n13950), .S(n16094), .Z(
        n13951) );
  AOI21_X1 U16134 ( .B1(n13953), .B2(n13952), .A(n13951), .ZN(n13954) );
  OAI21_X1 U16135 ( .B1(n13956), .B2(n13955), .A(n13954), .ZN(P3_U3435) );
  MUX2_X1 U16136 ( .A(P3_REG0_REG_9__SCAN_IN), .B(n13957), .S(n16094), .Z(
        P3_U3417) );
  MUX2_X1 U16137 ( .A(n13958), .B(P3_D_REG_1__SCAN_IN), .S(n13959), .Z(
        P3_U3377) );
  MUX2_X1 U16138 ( .A(n7478), .B(P3_D_REG_0__SCAN_IN), .S(n13959), .Z(P3_U3376) );
  NAND3_X1 U16139 ( .A1(n13961), .A2(P3_IR_REG_31__SCAN_IN), .A3(
        P3_STATE_REG_SCAN_IN), .ZN(n13964) );
  OAI22_X1 U16140 ( .A1(n13960), .A2(n13964), .B1(n13963), .B2(n13962), .ZN(
        n13965) );
  AOI21_X1 U16141 ( .B1(n13967), .B2(n13966), .A(n13965), .ZN(n13968) );
  INV_X1 U16142 ( .A(n13968), .ZN(P3_U3264) );
  INV_X1 U16143 ( .A(n13969), .ZN(n13972) );
  OR2_X1 U16144 ( .A1(n13974), .A2(n13973), .ZN(n13977) );
  AND2_X1 U16145 ( .A1(n13977), .A2(n13975), .ZN(n13979) );
  NAND2_X1 U16146 ( .A1(n13977), .A2(n13976), .ZN(n13978) );
  OAI21_X1 U16147 ( .B1(n13980), .B2(n13979), .A(n13978), .ZN(n13981) );
  NAND2_X1 U16148 ( .A1(n13981), .A2(n14065), .ZN(n13987) );
  OAI21_X1 U16149 ( .B1(n14090), .B2(n13983), .A(n13982), .ZN(n13984) );
  AOI21_X1 U16150 ( .B1(n13985), .B2(n14088), .A(n13984), .ZN(n13986) );
  OAI211_X1 U16151 ( .C1(n14187), .C2(n14073), .A(n13987), .B(n13986), .ZN(
        P2_U3187) );
  INV_X1 U16152 ( .A(n13988), .ZN(n13989) );
  NOR2_X1 U16153 ( .A1(n13989), .A2(n14063), .ZN(n14064) );
  NOR2_X1 U16154 ( .A1(n14064), .A2(n13990), .ZN(n13994) );
  XNOR2_X1 U16155 ( .A(n13992), .B(n13991), .ZN(n13993) );
  XNOR2_X1 U16156 ( .A(n13994), .B(n13993), .ZN(n14000) );
  AND2_X1 U16157 ( .A1(n14400), .A2(n14376), .ZN(n13995) );
  AOI21_X1 U16158 ( .B1(n14398), .B2(n14086), .A(n13995), .ZN(n14585) );
  INV_X1 U16159 ( .A(n14598), .ZN(n13996) );
  AOI22_X1 U16160 ( .A1(n13996), .A2(n14088), .B1(P2_REG3_REG_23__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13997) );
  OAI21_X1 U16161 ( .B1(n14585), .B2(n14090), .A(n13997), .ZN(n13998) );
  AOI21_X1 U16162 ( .B1(n14600), .B2(n14101), .A(n13998), .ZN(n13999) );
  OAI21_X1 U16163 ( .B1(n14000), .B2(n14103), .A(n13999), .ZN(P2_U3188) );
  NAND2_X1 U16164 ( .A1(n14002), .A2(n14001), .ZN(n14004) );
  XOR2_X1 U16165 ( .A(n14004), .B(n14003), .Z(n14008) );
  AOI22_X1 U16166 ( .A1(n14402), .A2(n14086), .B1(n14376), .B2(n14404), .ZN(
        n14659) );
  NAND2_X1 U16167 ( .A1(P2_U3088), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n14493)
         );
  NAND2_X1 U16168 ( .A1(n14088), .A2(n14661), .ZN(n14005) );
  OAI211_X1 U16169 ( .C1(n14659), .C2(n14090), .A(n14493), .B(n14005), .ZN(
        n14006) );
  AOI21_X1 U16170 ( .B1(n7907), .B2(n14101), .A(n14006), .ZN(n14007) );
  OAI21_X1 U16171 ( .B1(n14008), .B2(n14103), .A(n14007), .ZN(P2_U3191) );
  OAI211_X1 U16172 ( .C1(n14011), .C2(n14010), .A(n14009), .B(n14065), .ZN(
        n14016) );
  INV_X1 U16173 ( .A(n14012), .ZN(n14631) );
  AOI22_X1 U16174 ( .A1(n14400), .A2(n14086), .B1(n14376), .B2(n14402), .ZN(
        n14624) );
  OAI22_X1 U16175 ( .A1(n14624), .A2(n14090), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n14013), .ZN(n14014) );
  AOI21_X1 U16176 ( .B1(n14631), .B2(n14088), .A(n14014), .ZN(n14015) );
  OAI211_X1 U16177 ( .C1(n7905), .C2(n14073), .A(n14016), .B(n14015), .ZN(
        P2_U3195) );
  INV_X1 U16178 ( .A(n14562), .ZN(n14860) );
  OAI211_X1 U16179 ( .C1(n14019), .C2(n14018), .A(n14017), .B(n14065), .ZN(
        n14024) );
  OAI22_X1 U16180 ( .A1(n14266), .A2(n14096), .B1(n14261), .B2(n14095), .ZN(
        n14557) );
  INV_X1 U16181 ( .A(n14563), .ZN(n14021) );
  OAI22_X1 U16182 ( .A1(n14021), .A2(n14099), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n14020), .ZN(n14022) );
  AOI21_X1 U16183 ( .B1(n14557), .B2(n14097), .A(n14022), .ZN(n14023) );
  OAI211_X1 U16184 ( .C1(n14860), .C2(n14073), .A(n14024), .B(n14023), .ZN(
        P2_U3197) );
  NOR2_X1 U16185 ( .A1(n14026), .A2(n14025), .ZN(n14031) );
  XNOR2_X1 U16186 ( .A(n14027), .B(n14028), .ZN(n14094) );
  AOI22_X1 U16187 ( .A1(n14094), .A2(n14093), .B1(n14027), .B2(n14029), .ZN(
        n14030) );
  XOR2_X1 U16188 ( .A(n14031), .B(n14030), .Z(n14036) );
  NOR2_X1 U16189 ( .A1(n14099), .A2(n14707), .ZN(n14034) );
  AND2_X1 U16190 ( .A1(n14407), .A2(n14376), .ZN(n14032) );
  AOI21_X1 U16191 ( .B1(n14405), .B2(n14086), .A(n14032), .ZN(n14810) );
  OAI22_X1 U16192 ( .A1(n14810), .A2(n14090), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n15927), .ZN(n14033) );
  AOI211_X1 U16193 ( .C1(n14809), .C2(n14101), .A(n14034), .B(n14033), .ZN(
        n14035) );
  OAI21_X1 U16194 ( .B1(n14036), .B2(n14103), .A(n14035), .ZN(P2_U3198) );
  INV_X1 U16195 ( .A(n14038), .ZN(n14039) );
  AOI21_X1 U16196 ( .B1(n14037), .B2(n14040), .A(n14039), .ZN(n14045) );
  NOR2_X1 U16197 ( .A1(n14099), .A2(n14699), .ZN(n14043) );
  AOI22_X1 U16198 ( .A1(n14404), .A2(n14086), .B1(n14376), .B2(n14406), .ZN(
        n14689) );
  OAI21_X1 U16199 ( .B1(n14689), .B2(n14090), .A(n14041), .ZN(n14042) );
  AOI211_X1 U16200 ( .C1(n14697), .C2(n14101), .A(n14043), .B(n14042), .ZN(
        n14044) );
  OAI21_X1 U16201 ( .B1(n14045), .B2(n14103), .A(n14044), .ZN(P2_U3200) );
  OAI211_X1 U16202 ( .C1(n14048), .C2(n14047), .A(n14046), .B(n14065), .ZN(
        n14054) );
  NAND2_X1 U16203 ( .A1(n14397), .A2(n14086), .ZN(n14050) );
  NAND2_X1 U16204 ( .A1(n14399), .A2(n14376), .ZN(n14049) );
  NAND2_X1 U16205 ( .A1(n14050), .A2(n14049), .ZN(n14570) );
  OAI22_X1 U16206 ( .A1(n14574), .A2(n14099), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n14051), .ZN(n14052) );
  AOI21_X1 U16207 ( .B1(n14570), .B2(n14097), .A(n14052), .ZN(n14053) );
  OAI211_X1 U16208 ( .C1(n6952), .C2(n14073), .A(n14054), .B(n14053), .ZN(
        P2_U3201) );
  INV_X1 U16209 ( .A(n14055), .ZN(n14056) );
  AOI21_X1 U16210 ( .B1(n14058), .B2(n14057), .A(n14056), .ZN(n14062) );
  OAI22_X1 U16211 ( .A1(n14068), .A2(n14096), .B1(n14076), .B2(n14095), .ZN(
        n14650) );
  AOI22_X1 U16212 ( .A1(n14650), .A2(n14097), .B1(P2_REG3_REG_20__SCAN_IN), 
        .B2(P2_U3088), .ZN(n14059) );
  OAI21_X1 U16213 ( .B1(n14641), .B2(n14099), .A(n14059), .ZN(n14060) );
  AOI21_X1 U16214 ( .B1(n14790), .B2(n14101), .A(n14060), .ZN(n14061) );
  OAI21_X1 U16215 ( .B1(n14062), .B2(n14103), .A(n14061), .ZN(P2_U3205) );
  INV_X1 U16216 ( .A(n14063), .ZN(n14067) );
  INV_X1 U16217 ( .A(n14064), .ZN(n14066) );
  OAI211_X1 U16218 ( .C1(n13988), .C2(n14067), .A(n14066), .B(n14065), .ZN(
        n14072) );
  OAI22_X1 U16219 ( .A1(n14254), .A2(n14096), .B1(n14068), .B2(n14095), .ZN(
        n14606) );
  OAI22_X1 U16220 ( .A1(n14616), .A2(n14099), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n14069), .ZN(n14070) );
  AOI21_X1 U16221 ( .B1(n14606), .B2(n14097), .A(n14070), .ZN(n14071) );
  OAI211_X1 U16222 ( .C1(n14869), .C2(n14073), .A(n14072), .B(n14071), .ZN(
        P2_U3207) );
  XNOR2_X1 U16223 ( .A(n14074), .B(n14075), .ZN(n14081) );
  OAI22_X1 U16224 ( .A1(n14076), .A2(n14096), .B1(n14204), .B2(n14095), .ZN(
        n14673) );
  NAND2_X1 U16225 ( .A1(n14673), .A2(n14097), .ZN(n14078) );
  OAI211_X1 U16226 ( .C1(n14099), .C2(n14678), .A(n14078), .B(n14077), .ZN(
        n14079) );
  AOI21_X1 U16227 ( .B1(n14800), .B2(n14101), .A(n14079), .ZN(n14080) );
  OAI21_X1 U16228 ( .B1(n14081), .B2(n14103), .A(n14080), .ZN(P2_U3210) );
  AND2_X1 U16229 ( .A1(n14397), .A2(n14376), .ZN(n14085) );
  AOI21_X1 U16230 ( .B1(n14395), .B2(n14086), .A(n14085), .ZN(n14543) );
  INV_X1 U16231 ( .A(n14087), .ZN(n14548) );
  AOI22_X1 U16232 ( .A1(n14548), .A2(n14088), .B1(P2_REG3_REG_26__SCAN_IN), 
        .B2(P2_U3088), .ZN(n14089) );
  OAI21_X1 U16233 ( .B1(n14543), .B2(n14090), .A(n14089), .ZN(n14091) );
  AOI21_X1 U16234 ( .B1(n14549), .B2(n14101), .A(n14091), .ZN(n14092) );
  XNOR2_X1 U16235 ( .A(n14094), .B(n14093), .ZN(n14104) );
  OAI22_X1 U16236 ( .A1(n14178), .A2(n14096), .B1(n14188), .B2(n14095), .ZN(
        n14728) );
  AOI22_X1 U16237 ( .A1(n14097), .A2(n14728), .B1(P2_REG3_REG_15__SCAN_IN), 
        .B2(P2_U3088), .ZN(n14098) );
  OAI21_X1 U16238 ( .B1(n14099), .B2(n14735), .A(n14098), .ZN(n14100) );
  AOI21_X1 U16239 ( .B1(n14817), .B2(n14101), .A(n14100), .ZN(n14102) );
  OAI21_X1 U16240 ( .B1(n14104), .B2(n14103), .A(n14102), .ZN(P2_U3213) );
  MUX2_X1 U16241 ( .A(n14399), .B(n14600), .S(n14267), .Z(n14256) );
  INV_X1 U16242 ( .A(n14256), .ZN(n14260) );
  NAND2_X1 U16243 ( .A1(n14108), .A2(n14265), .ZN(n14109) );
  OAI211_X1 U16244 ( .C1(n14110), .C2(n14323), .A(n14421), .B(n14265), .ZN(
        n14111) );
  NAND2_X1 U16245 ( .A1(n14112), .A2(n14111), .ZN(n14117) );
  MUX2_X1 U16246 ( .A(n8040), .B(n14114), .S(n14265), .Z(n14113) );
  INV_X1 U16247 ( .A(n14113), .ZN(n14116) );
  MUX2_X1 U16248 ( .A(n14114), .B(n8040), .S(n14265), .Z(n14115) );
  OAI21_X1 U16249 ( .B1(n14117), .B2(n14116), .A(n14115), .ZN(n14119) );
  NAND2_X1 U16250 ( .A1(n14117), .A2(n14116), .ZN(n14118) );
  NAND2_X1 U16251 ( .A1(n14119), .A2(n14118), .ZN(n14123) );
  MUX2_X1 U16252 ( .A(n14120), .B(n14420), .S(n14265), .Z(n14124) );
  NAND2_X1 U16253 ( .A1(n14123), .A2(n14124), .ZN(n14122) );
  MUX2_X1 U16254 ( .A(n14420), .B(n14120), .S(n14265), .Z(n14121) );
  NAND2_X1 U16255 ( .A1(n14122), .A2(n14121), .ZN(n14128) );
  INV_X1 U16256 ( .A(n14123), .ZN(n14126) );
  INV_X1 U16257 ( .A(n14124), .ZN(n14125) );
  NAND2_X1 U16258 ( .A1(n14128), .A2(n14127), .ZN(n14132) );
  MUX2_X1 U16259 ( .A(n14419), .B(n14129), .S(n14267), .Z(n14133) );
  NAND2_X1 U16260 ( .A1(n14132), .A2(n14133), .ZN(n14131) );
  MUX2_X1 U16261 ( .A(n14129), .B(n14419), .S(n14265), .Z(n14130) );
  INV_X1 U16262 ( .A(n14132), .ZN(n14135) );
  INV_X1 U16263 ( .A(n14133), .ZN(n14134) );
  MUX2_X1 U16264 ( .A(n14136), .B(n14418), .S(n14265), .Z(n14138) );
  MUX2_X1 U16265 ( .A(n14418), .B(n14136), .S(n14265), .Z(n14137) );
  INV_X1 U16266 ( .A(n14138), .ZN(n14139) );
  MUX2_X1 U16267 ( .A(n14417), .B(n15983), .S(n14267), .Z(n14143) );
  MUX2_X1 U16268 ( .A(n15983), .B(n14417), .S(n14267), .Z(n14140) );
  NAND2_X1 U16269 ( .A1(n14141), .A2(n14140), .ZN(n14147) );
  INV_X1 U16270 ( .A(n14142), .ZN(n14145) );
  INV_X1 U16271 ( .A(n14143), .ZN(n14144) );
  NAND2_X1 U16272 ( .A1(n14145), .A2(n14144), .ZN(n14146) );
  MUX2_X1 U16273 ( .A(n14148), .B(n14416), .S(n14265), .Z(n14150) );
  MUX2_X1 U16274 ( .A(n14416), .B(n14148), .S(n14265), .Z(n14149) );
  INV_X1 U16275 ( .A(n14150), .ZN(n14151) );
  MUX2_X1 U16276 ( .A(n14415), .B(n15995), .S(n14265), .Z(n14153) );
  MUX2_X1 U16277 ( .A(n14415), .B(n15995), .S(n14263), .Z(n14152) );
  MUX2_X1 U16278 ( .A(n14414), .B(n14154), .S(n14316), .Z(n14157) );
  MUX2_X1 U16279 ( .A(n14414), .B(n14154), .S(n14265), .Z(n14155) );
  INV_X1 U16280 ( .A(n14157), .ZN(n14158) );
  MUX2_X1 U16281 ( .A(n14413), .B(n14159), .S(n14238), .Z(n14163) );
  MUX2_X1 U16282 ( .A(n14413), .B(n14159), .S(n14316), .Z(n14160) );
  NAND2_X1 U16283 ( .A1(n14161), .A2(n14160), .ZN(n14167) );
  INV_X1 U16284 ( .A(n14162), .ZN(n14165) );
  INV_X1 U16285 ( .A(n14163), .ZN(n14164) );
  NAND2_X1 U16286 ( .A1(n14165), .A2(n14164), .ZN(n14166) );
  MUX2_X1 U16287 ( .A(n14412), .B(n14842), .S(n14316), .Z(n14169) );
  MUX2_X1 U16288 ( .A(n14412), .B(n14842), .S(n14238), .Z(n14168) );
  MUX2_X1 U16289 ( .A(n14411), .B(n14171), .S(n14238), .Z(n14170) );
  MUX2_X1 U16290 ( .A(n14411), .B(n14171), .S(n14263), .Z(n14172) );
  MUX2_X1 U16291 ( .A(n14174), .B(n14173), .S(n14238), .Z(n14193) );
  MUX2_X1 U16292 ( .A(n14410), .B(n14829), .S(n14263), .Z(n14192) );
  NAND2_X1 U16293 ( .A1(n14193), .A2(n14192), .ZN(n14175) );
  MUX2_X1 U16294 ( .A(n14407), .B(n14817), .S(n14238), .Z(n14206) );
  NAND2_X1 U16295 ( .A1(n14207), .A2(n14206), .ZN(n14186) );
  INV_X1 U16296 ( .A(n14265), .ZN(n14263) );
  NAND2_X1 U16297 ( .A1(n14216), .A2(n14405), .ZN(n14179) );
  NAND2_X1 U16298 ( .A1(n14178), .A2(n14263), .ZN(n14181) );
  AOI21_X1 U16299 ( .B1(n14179), .B2(n14181), .A(n14882), .ZN(n14185) );
  NAND2_X1 U16300 ( .A1(n14216), .A2(n14204), .ZN(n14180) );
  OR2_X1 U16301 ( .A1(n14809), .A2(n14316), .ZN(n14211) );
  AOI21_X1 U16302 ( .B1(n14180), .B2(n14211), .A(n14697), .ZN(n14184) );
  NAND2_X1 U16303 ( .A1(n14405), .A2(n14267), .ZN(n14213) );
  OR2_X1 U16304 ( .A1(n14809), .A2(n14213), .ZN(n14183) );
  INV_X1 U16305 ( .A(n14181), .ZN(n14205) );
  NAND2_X1 U16306 ( .A1(n14204), .A2(n14205), .ZN(n14182) );
  NAND2_X1 U16307 ( .A1(n14183), .A2(n14182), .ZN(n14215) );
  OR3_X1 U16308 ( .A1(n14185), .A2(n14184), .A3(n14215), .ZN(n14210) );
  NAND2_X1 U16309 ( .A1(n14186), .A2(n14210), .ZN(n14203) );
  MUX2_X1 U16310 ( .A(n14188), .B(n14187), .S(n14263), .Z(n14199) );
  MUX2_X1 U16311 ( .A(n14408), .B(n14824), .S(n14238), .Z(n14198) );
  AND2_X1 U16312 ( .A1(n14199), .A2(n14198), .ZN(n14189) );
  MUX2_X1 U16313 ( .A(n14190), .B(n6951), .S(n14263), .Z(n14223) );
  MUX2_X1 U16314 ( .A(n14409), .B(n14191), .S(n14238), .Z(n14222) );
  INV_X1 U16315 ( .A(n14192), .ZN(n14195) );
  INV_X1 U16316 ( .A(n14193), .ZN(n14194) );
  AOI22_X1 U16317 ( .A1(n14223), .A2(n14222), .B1(n14195), .B2(n14194), .ZN(
        n14196) );
  INV_X1 U16318 ( .A(n14198), .ZN(n14201) );
  INV_X1 U16319 ( .A(n14199), .ZN(n14200) );
  NAND2_X1 U16320 ( .A1(n14201), .A2(n14200), .ZN(n14202) );
  NOR2_X1 U16321 ( .A1(n14203), .A2(n14202), .ZN(n14221) );
  AOI22_X1 U16322 ( .A1(n14216), .A2(n14205), .B1(n14204), .B2(n14263), .ZN(
        n14219) );
  INV_X1 U16323 ( .A(n14206), .ZN(n14209) );
  INV_X1 U16324 ( .A(n14207), .ZN(n14208) );
  INV_X1 U16325 ( .A(n14211), .ZN(n14212) );
  NAND2_X1 U16326 ( .A1(n14216), .A2(n14212), .ZN(n14214) );
  NAND2_X1 U16327 ( .A1(n14214), .A2(n14213), .ZN(n14217) );
  AOI22_X1 U16328 ( .A1(n14217), .A2(n14882), .B1(n14216), .B2(n14215), .ZN(
        n14218) );
  NOR2_X1 U16329 ( .A1(n14221), .A2(n14220), .ZN(n14228) );
  INV_X1 U16330 ( .A(n14222), .ZN(n14225) );
  INV_X1 U16331 ( .A(n14223), .ZN(n14224) );
  NAND3_X1 U16332 ( .A1(n14226), .A2(n14225), .A3(n14224), .ZN(n14227) );
  MUX2_X1 U16333 ( .A(n14404), .B(n14800), .S(n14263), .Z(n14229) );
  MUX2_X1 U16334 ( .A(n14404), .B(n14800), .S(n14238), .Z(n14230) );
  MUX2_X1 U16335 ( .A(n14403), .B(n7907), .S(n14238), .Z(n14234) );
  NAND2_X1 U16336 ( .A1(n14235), .A2(n14234), .ZN(n14233) );
  MUX2_X1 U16337 ( .A(n14403), .B(n7907), .S(n14263), .Z(n14232) );
  NAND2_X1 U16338 ( .A1(n14233), .A2(n14232), .ZN(n14237) );
  MUX2_X1 U16339 ( .A(n14402), .B(n14790), .S(n14263), .Z(n14241) );
  MUX2_X1 U16340 ( .A(n14402), .B(n14790), .S(n14238), .Z(n14239) );
  INV_X1 U16341 ( .A(n14241), .ZN(n14242) );
  MUX2_X1 U16342 ( .A(n14401), .B(n14628), .S(n14267), .Z(n14245) );
  MUX2_X1 U16343 ( .A(n14401), .B(n14628), .S(n14263), .Z(n14243) );
  NAND2_X1 U16344 ( .A1(n14244), .A2(n14243), .ZN(n14247) );
  AND2_X1 U16345 ( .A1(n14247), .A2(n14246), .ZN(n14251) );
  MUX2_X1 U16346 ( .A(n14869), .B(n14248), .S(n14267), .Z(n14250) );
  MUX2_X1 U16347 ( .A(n14400), .B(n14618), .S(n14267), .Z(n14249) );
  NAND2_X1 U16348 ( .A1(n14253), .A2(n14252), .ZN(n14257) );
  INV_X1 U16349 ( .A(n14257), .ZN(n14259) );
  MUX2_X1 U16350 ( .A(n14865), .B(n14254), .S(n14267), .Z(n14255) );
  AOI21_X1 U16351 ( .B1(n14257), .B2(n14256), .A(n14255), .ZN(n14258) );
  MUX2_X1 U16352 ( .A(n14769), .B(n14398), .S(n14263), .Z(n14277) );
  MUX2_X1 U16353 ( .A(n6952), .B(n14261), .S(n14238), .Z(n14278) );
  MUX2_X1 U16354 ( .A(n14262), .B(n14860), .S(n14238), .Z(n14282) );
  MUX2_X1 U16355 ( .A(n14562), .B(n14397), .S(n14267), .Z(n14281) );
  MUX2_X1 U16356 ( .A(n14395), .B(n14749), .S(n14267), .Z(n14288) );
  MUX2_X1 U16357 ( .A(n14396), .B(n14549), .S(n14267), .Z(n14284) );
  AOI22_X1 U16358 ( .A1(n14290), .A2(n14288), .B1(n14285), .B2(n14284), .ZN(
        n14283) );
  OAI21_X1 U16359 ( .B1(n14282), .B2(n14281), .A(n14283), .ZN(n14279) );
  NOR2_X1 U16360 ( .A1(n14317), .A2(n14263), .ZN(n14274) );
  INV_X1 U16361 ( .A(n14383), .ZN(n14269) );
  NOR2_X1 U16362 ( .A1(n14269), .A2(n14379), .ZN(n14369) );
  NOR3_X1 U16363 ( .A1(n14274), .A2(n14369), .A3(n14270), .ZN(n14271) );
  OAI22_X1 U16364 ( .A1(n14511), .A2(n14238), .B1(n14326), .B2(n14271), .ZN(
        n14309) );
  MUX2_X1 U16365 ( .A(n14326), .B(n14511), .S(n14238), .Z(n14308) );
  INV_X1 U16366 ( .A(n14393), .ZN(n14273) );
  MUX2_X1 U16367 ( .A(n14273), .B(n14272), .S(n14238), .Z(n14300) );
  MUX2_X1 U16368 ( .A(n14744), .B(n14393), .S(n14238), .Z(n14299) );
  AOI22_X1 U16369 ( .A1(n14309), .A2(n14308), .B1(n14300), .B2(n14299), .ZN(
        n14276) );
  MUX2_X1 U16370 ( .A(n14274), .B(n14317), .S(n14318), .Z(n14275) );
  NOR2_X1 U16371 ( .A1(n14276), .A2(n14275), .ZN(n14314) );
  NOR3_X1 U16372 ( .A1(n14279), .A2(n14278), .A3(n14277), .ZN(n14298) );
  INV_X1 U16373 ( .A(n14394), .ZN(n14280) );
  MUX2_X1 U16374 ( .A(n14280), .B(n14853), .S(n14263), .Z(n14302) );
  MUX2_X1 U16375 ( .A(n14394), .B(n14519), .S(n14238), .Z(n14301) );
  NAND3_X1 U16376 ( .A1(n14283), .A2(n14282), .A3(n14281), .ZN(n14296) );
  INV_X1 U16377 ( .A(n14284), .ZN(n14287) );
  INV_X1 U16378 ( .A(n14285), .ZN(n14286) );
  NAND2_X1 U16379 ( .A1(n14287), .A2(n14286), .ZN(n14289) );
  NAND2_X1 U16380 ( .A1(n14290), .A2(n14289), .ZN(n14294) );
  INV_X1 U16381 ( .A(n14288), .ZN(n14293) );
  INV_X1 U16382 ( .A(n14289), .ZN(n14292) );
  INV_X1 U16383 ( .A(n14290), .ZN(n14291) );
  AOI22_X1 U16384 ( .A1(n14294), .A2(n14293), .B1(n14292), .B2(n14291), .ZN(
        n14295) );
  OAI211_X1 U16385 ( .C1(n14302), .C2(n14301), .A(n14296), .B(n14295), .ZN(
        n14297) );
  INV_X1 U16386 ( .A(n14299), .ZN(n14307) );
  INV_X1 U16387 ( .A(n14300), .ZN(n14306) );
  INV_X1 U16388 ( .A(n14301), .ZN(n14304) );
  INV_X1 U16389 ( .A(n14302), .ZN(n14303) );
  INV_X1 U16390 ( .A(n14317), .ZN(n14391) );
  XNOR2_X1 U16391 ( .A(n14318), .B(n14391), .ZN(n14366) );
  OAI21_X1 U16392 ( .B1(n14304), .B2(n14303), .A(n14366), .ZN(n14305) );
  AOI21_X1 U16393 ( .B1(n14307), .B2(n14306), .A(n14305), .ZN(n14313) );
  INV_X1 U16394 ( .A(n14308), .ZN(n14311) );
  INV_X1 U16395 ( .A(n14309), .ZN(n14310) );
  NAND3_X1 U16396 ( .A1(n14849), .A2(n14316), .A3(n14391), .ZN(n14320) );
  NAND3_X1 U16397 ( .A1(n14318), .A2(n14317), .A3(n14238), .ZN(n14319) );
  INV_X1 U16398 ( .A(n14374), .ZN(n14325) );
  OAI22_X1 U16399 ( .A1(n14323), .A2(n7741), .B1(n14322), .B2(n14321), .ZN(
        n14324) );
  INV_X1 U16400 ( .A(n14511), .ZN(n14327) );
  INV_X1 U16401 ( .A(n14326), .ZN(n14392) );
  XNOR2_X1 U16402 ( .A(n14327), .B(n14392), .ZN(n14365) );
  INV_X1 U16403 ( .A(n14328), .ZN(n14352) );
  NOR2_X1 U16404 ( .A1(n14330), .A2(n14329), .ZN(n14334) );
  NAND4_X1 U16405 ( .A1(n14334), .A2(n14333), .A3(n14332), .A4(n14331), .ZN(
        n14336) );
  NOR2_X1 U16406 ( .A1(n14336), .A2(n14335), .ZN(n14342) );
  NOR2_X1 U16407 ( .A1(n14338), .A2(n14337), .ZN(n14340) );
  NAND4_X1 U16408 ( .A1(n14342), .A2(n14341), .A3(n14340), .A4(n14339), .ZN(
        n14343) );
  NOR2_X1 U16409 ( .A1(n14344), .A2(n14343), .ZN(n14347) );
  NAND4_X1 U16410 ( .A1(n14348), .A2(n14347), .A3(n14346), .A4(n14345), .ZN(
        n14349) );
  NOR2_X1 U16411 ( .A1(n14350), .A2(n14349), .ZN(n14351) );
  XNOR2_X1 U16412 ( .A(n14809), .B(n14406), .ZN(n14716) );
  NAND4_X1 U16413 ( .A1(n14352), .A2(n14351), .A3(n14695), .A4(n14716), .ZN(
        n14355) );
  NAND2_X1 U16414 ( .A1(n14671), .A2(n14353), .ZN(n14354) );
  NOR3_X1 U16415 ( .A1(n14604), .A2(n14355), .A3(n14354), .ZN(n14356) );
  NAND4_X1 U16416 ( .A1(n14356), .A2(n14657), .A3(n14626), .A4(n14646), .ZN(
        n14359) );
  NOR2_X1 U16417 ( .A1(n14359), .A2(n14592), .ZN(n14360) );
  NAND4_X1 U16418 ( .A1(n14545), .A2(n14360), .A3(n14569), .A4(n14560), .ZN(
        n14361) );
  NOR3_X1 U16419 ( .A1(n14362), .A2(n8539), .A3(n14361), .ZN(n14364) );
  NAND4_X1 U16420 ( .A1(n14366), .A2(n14365), .A3(n14364), .A4(n14363), .ZN(
        n14368) );
  OR2_X1 U16421 ( .A1(n14368), .A2(n8584), .ZN(n14367) );
  NAND2_X1 U16422 ( .A1(n14368), .A2(n8584), .ZN(n14385) );
  NAND2_X1 U16423 ( .A1(n14387), .A2(n14385), .ZN(n14371) );
  INV_X1 U16424 ( .A(n14369), .ZN(n14370) );
  OAI211_X1 U16425 ( .C1(n14372), .C2(n8584), .A(n14371), .B(n14370), .ZN(
        n14373) );
  NAND3_X1 U16426 ( .A1(n14374), .A2(n14382), .A3(n14373), .ZN(n14390) );
  NAND4_X1 U16427 ( .A1(n15981), .A2(n14377), .A3(n14376), .A4(n14375), .ZN(
        n14381) );
  AOI21_X1 U16428 ( .B1(n14382), .B2(n14379), .A(n14378), .ZN(n14380) );
  NAND2_X1 U16429 ( .A1(n14381), .A2(n14380), .ZN(n14389) );
  INV_X1 U16430 ( .A(n14382), .ZN(n14384) );
  NOR2_X1 U16431 ( .A1(n14384), .A2(n14383), .ZN(n14386) );
  NAND3_X1 U16432 ( .A1(n14387), .A2(n14386), .A3(n14385), .ZN(n14388) );
  MUX2_X1 U16433 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(n14391), .S(n15887), .Z(
        P2_U3562) );
  MUX2_X1 U16434 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(n14392), .S(n15887), .Z(
        P2_U3561) );
  MUX2_X1 U16435 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(n14393), .S(n15887), .Z(
        P2_U3560) );
  MUX2_X1 U16436 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(n14394), .S(n15887), .Z(
        P2_U3559) );
  MUX2_X1 U16437 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n14395), .S(n15887), .Z(
        P2_U3558) );
  MUX2_X1 U16438 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(n14396), .S(n15887), .Z(
        P2_U3557) );
  MUX2_X1 U16439 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n14397), .S(n15887), .Z(
        P2_U3556) );
  MUX2_X1 U16440 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(n14398), .S(n15887), .Z(
        P2_U3555) );
  MUX2_X1 U16441 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(n14399), .S(n15887), .Z(
        P2_U3554) );
  MUX2_X1 U16442 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n14400), .S(n15887), .Z(
        P2_U3553) );
  MUX2_X1 U16443 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n14401), .S(n15887), .Z(
        P2_U3552) );
  MUX2_X1 U16444 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n14402), .S(n15887), .Z(
        P2_U3551) );
  MUX2_X1 U16445 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n14403), .S(n15887), .Z(
        P2_U3550) );
  MUX2_X1 U16446 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(n14404), .S(n15887), .Z(
        P2_U3549) );
  MUX2_X1 U16447 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n14405), .S(n15887), .Z(
        P2_U3548) );
  MUX2_X1 U16448 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n14406), .S(n15887), .Z(
        P2_U3547) );
  MUX2_X1 U16449 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(n14407), .S(n15887), .Z(
        P2_U3546) );
  MUX2_X1 U16450 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(n14408), .S(n15887), .Z(
        P2_U3545) );
  MUX2_X1 U16451 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(n14409), .S(n15887), .Z(
        P2_U3544) );
  MUX2_X1 U16452 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(n14410), .S(n15887), .Z(
        P2_U3543) );
  MUX2_X1 U16453 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(n14411), .S(n15887), .Z(
        P2_U3542) );
  MUX2_X1 U16454 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(n14412), .S(n15887), .Z(
        P2_U3541) );
  MUX2_X1 U16455 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(n14413), .S(P2_U3947), .Z(
        P2_U3540) );
  MUX2_X1 U16456 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(n14414), .S(P2_U3947), .Z(
        P2_U3539) );
  MUX2_X1 U16457 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(n14415), .S(P2_U3947), .Z(
        P2_U3538) );
  MUX2_X1 U16458 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(n14416), .S(n15887), .Z(
        P2_U3537) );
  MUX2_X1 U16459 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(n14417), .S(P2_U3947), .Z(
        P2_U3536) );
  MUX2_X1 U16460 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(n14418), .S(P2_U3947), .Z(
        P2_U3535) );
  MUX2_X1 U16461 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(n14419), .S(P2_U3947), .Z(
        P2_U3534) );
  MUX2_X1 U16462 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(n14420), .S(P2_U3947), .Z(
        P2_U3533) );
  MUX2_X1 U16463 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(n8040), .S(P2_U3947), .Z(
        P2_U3532) );
  MUX2_X1 U16464 ( .A(P2_DATAO_REG_0__SCAN_IN), .B(n14421), .S(P2_U3947), .Z(
        P2_U3531) );
  NOR2_X1 U16465 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8057), .ZN(n14424) );
  NOR2_X1 U16466 ( .A1(n15944), .A2(n14422), .ZN(n14423) );
  AOI211_X1 U16467 ( .C1(n15936), .C2(n14428), .A(n14424), .B(n14423), .ZN(
        n14434) );
  OAI211_X1 U16468 ( .C1(n14427), .C2(n14426), .A(n15928), .B(n14425), .ZN(
        n14433) );
  MUX2_X1 U16469 ( .A(n11159), .B(P2_REG2_REG_3__SCAN_IN), .S(n14428), .Z(
        n14429) );
  NAND3_X1 U16470 ( .A1(n15907), .A2(n14430), .A3(n14429), .ZN(n14431) );
  NAND3_X1 U16471 ( .A1(n15937), .A2(n14443), .A3(n14431), .ZN(n14432) );
  NAND3_X1 U16472 ( .A1(n14434), .A2(n14433), .A3(n14432), .ZN(P2_U3217) );
  INV_X1 U16473 ( .A(n14435), .ZN(n14436) );
  AOI21_X1 U16474 ( .B1(n15936), .B2(n14440), .A(n14436), .ZN(n14448) );
  OAI211_X1 U16475 ( .C1(n14439), .C2(n14438), .A(n15928), .B(n14437), .ZN(
        n14447) );
  MUX2_X1 U16476 ( .A(n11162), .B(P2_REG2_REG_4__SCAN_IN), .S(n14440), .Z(
        n14441) );
  NAND3_X1 U16477 ( .A1(n14443), .A2(n14442), .A3(n14441), .ZN(n14444) );
  NAND3_X1 U16478 ( .A1(n15937), .A2(n14454), .A3(n14444), .ZN(n14446) );
  NAND2_X1 U16479 ( .A1(n15899), .A2(P2_ADDR_REG_4__SCAN_IN), .ZN(n14445) );
  NAND4_X1 U16480 ( .A1(n14448), .A2(n14447), .A3(n14446), .A4(n14445), .ZN(
        P2_U3218) );
  INV_X1 U16481 ( .A(n14449), .ZN(n14450) );
  AOI21_X1 U16482 ( .B1(n15936), .B2(n14451), .A(n14450), .ZN(n14463) );
  NAND2_X1 U16483 ( .A1(n15899), .A2(P2_ADDR_REG_5__SCAN_IN), .ZN(n14462) );
  MUX2_X1 U16484 ( .A(n12224), .B(P2_REG2_REG_5__SCAN_IN), .S(n14451), .Z(
        n14452) );
  NAND3_X1 U16485 ( .A1(n14454), .A2(n14453), .A3(n14452), .ZN(n14455) );
  NAND3_X1 U16486 ( .A1(n15937), .A2(n14456), .A3(n14455), .ZN(n14461) );
  OAI211_X1 U16487 ( .C1(n14459), .C2(n14458), .A(n15928), .B(n14457), .ZN(
        n14460) );
  NAND4_X1 U16488 ( .A1(n14463), .A2(n14462), .A3(n14461), .A4(n14460), .ZN(
        P2_U3219) );
  NOR2_X1 U16489 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8143), .ZN(n14466) );
  NOR2_X1 U16490 ( .A1(n15944), .A2(n14464), .ZN(n14465) );
  AOI211_X1 U16491 ( .C1(n15936), .C2(n14470), .A(n14466), .B(n14465), .ZN(
        n14476) );
  OAI211_X1 U16492 ( .C1(n14469), .C2(n14468), .A(n15928), .B(n14467), .ZN(
        n14475) );
  MUX2_X1 U16493 ( .A(n12238), .B(P2_REG2_REG_7__SCAN_IN), .S(n14470), .Z(
        n14471) );
  NAND3_X1 U16494 ( .A1(n15921), .A2(n14472), .A3(n14471), .ZN(n14473) );
  NAND3_X1 U16495 ( .A1(n15937), .A2(n14487), .A3(n14473), .ZN(n14474) );
  NAND3_X1 U16496 ( .A1(n14476), .A2(n14475), .A3(n14474), .ZN(P2_U3221) );
  INV_X1 U16497 ( .A(n14477), .ZN(n14480) );
  NOR2_X1 U16498 ( .A1(n15944), .A2(n14478), .ZN(n14479) );
  AOI211_X1 U16499 ( .C1(n15936), .C2(n14484), .A(n14480), .B(n14479), .ZN(
        n14492) );
  OAI211_X1 U16500 ( .C1(n14483), .C2(n14482), .A(n15928), .B(n14481), .ZN(
        n14491) );
  MUX2_X1 U16501 ( .A(n11170), .B(P2_REG2_REG_8__SCAN_IN), .S(n14484), .Z(
        n14485) );
  NAND3_X1 U16502 ( .A1(n14487), .A2(n14486), .A3(n14485), .ZN(n14488) );
  NAND3_X1 U16503 ( .A1(n15937), .A2(n14489), .A3(n14488), .ZN(n14490) );
  NAND3_X1 U16504 ( .A1(n14492), .A2(n14491), .A3(n14490), .ZN(P2_U3222) );
  INV_X1 U16505 ( .A(n14493), .ZN(n14506) );
  NAND2_X1 U16506 ( .A1(n14495), .A2(n14494), .ZN(n14496) );
  XNOR2_X1 U16507 ( .A(n14496), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n14503) );
  INV_X1 U16508 ( .A(n14503), .ZN(n14502) );
  NAND2_X1 U16509 ( .A1(n14498), .A2(n14497), .ZN(n14500) );
  XNOR2_X1 U16510 ( .A(n14500), .B(n14499), .ZN(n14505) );
  NAND2_X1 U16511 ( .A1(n14505), .A2(n15937), .ZN(n14501) );
  NOR2_X1 U16512 ( .A1(n14719), .A2(n14507), .ZN(n14513) );
  NOR2_X1 U16513 ( .A1(n14849), .A2(n14698), .ZN(n14508) );
  AOI211_X1 U16514 ( .C1(P2_REG2_REG_31__SCAN_IN), .C2(n14719), .A(n14513), 
        .B(n14508), .ZN(n14509) );
  OAI21_X1 U16515 ( .B1(n14721), .B2(n14510), .A(n14509), .ZN(P2_U3234) );
  NOR2_X1 U16516 ( .A1(n14511), .A2(n14698), .ZN(n14512) );
  AOI211_X1 U16517 ( .C1(n14719), .C2(P2_REG2_REG_30__SCAN_IN), .A(n14513), 
        .B(n14512), .ZN(n14514) );
  OAI21_X1 U16518 ( .B1(n14721), .B2(n14515), .A(n14514), .ZN(P2_U3235) );
  AOI21_X1 U16519 ( .B1(n14517), .B2(n14713), .A(n14516), .ZN(n14525) );
  INV_X1 U16520 ( .A(n14518), .ZN(n14523) );
  AOI22_X1 U16521 ( .A1(n14519), .A2(n14739), .B1(P2_REG2_REG_28__SCAN_IN), 
        .B2(n14738), .ZN(n14520) );
  OAI21_X1 U16522 ( .B1(n14521), .B2(n14721), .A(n14520), .ZN(n14522) );
  AOI21_X1 U16523 ( .B1(n14523), .B2(n14723), .A(n14522), .ZN(n14524) );
  OAI21_X1 U16524 ( .B1(n14525), .B2(n14738), .A(n14524), .ZN(P2_U3237) );
  XNOR2_X1 U16525 ( .A(n14526), .B(n14536), .ZN(n14527) );
  NAND2_X1 U16526 ( .A1(n14527), .A2(n14675), .ZN(n14529) );
  OAI211_X1 U16527 ( .C1(n14546), .C2(n14531), .A(n14818), .B(n14530), .ZN(
        n14750) );
  AOI22_X1 U16528 ( .A1(n14532), .A2(n14713), .B1(P2_REG2_REG_27__SCAN_IN), 
        .B2(n14738), .ZN(n14534) );
  NAND2_X1 U16529 ( .A1(n14749), .A2(n14739), .ZN(n14533) );
  OAI211_X1 U16530 ( .C1(n14750), .C2(n14721), .A(n14534), .B(n14533), .ZN(
        n14539) );
  NAND2_X1 U16531 ( .A1(n14537), .A2(n14536), .ZN(n14748) );
  AND3_X1 U16532 ( .A1(n14535), .A2(n14723), .A3(n14748), .ZN(n14538) );
  AOI211_X1 U16533 ( .C1(n14754), .C2(n6548), .A(n14539), .B(n14538), .ZN(
        n14540) );
  INV_X1 U16534 ( .A(n14540), .ZN(P2_U3238) );
  XNOR2_X1 U16535 ( .A(n14541), .B(n14545), .ZN(n14542) );
  NAND2_X1 U16536 ( .A1(n14542), .A2(n14675), .ZN(n14544) );
  NAND2_X1 U16537 ( .A1(n14544), .A2(n14543), .ZN(n14761) );
  INV_X1 U16538 ( .A(n14761), .ZN(n14554) );
  OAI21_X1 U16539 ( .B1(n14561), .B2(n14759), .A(n14818), .ZN(n14547) );
  AOI22_X1 U16540 ( .A1(n14548), .A2(n14713), .B1(P2_REG2_REG_26__SCAN_IN), 
        .B2(n14738), .ZN(n14551) );
  NAND2_X1 U16541 ( .A1(n14549), .A2(n14739), .ZN(n14550) );
  OAI211_X1 U16542 ( .C1(n14758), .C2(n14721), .A(n14551), .B(n14550), .ZN(
        n14552) );
  AOI21_X1 U16543 ( .B1(n14757), .B2(n14723), .A(n14552), .ZN(n14553) );
  OAI21_X1 U16544 ( .B1(n14554), .B2(n14738), .A(n14553), .ZN(P2_U3239) );
  OAI21_X1 U16545 ( .B1(n14556), .B2(n14560), .A(n14555), .ZN(n14558) );
  AOI21_X1 U16546 ( .B1(n14558), .B2(n14675), .A(n14557), .ZN(n14762) );
  XNOR2_X1 U16547 ( .A(n14559), .B(n14560), .ZN(n14765) );
  AOI211_X1 U16548 ( .C1(n14562), .C2(n14572), .A(n14717), .B(n14561), .ZN(
        n14764) );
  NAND2_X1 U16549 ( .A1(n14764), .A2(n14703), .ZN(n14565) );
  AOI22_X1 U16550 ( .A1(n14563), .A2(n14713), .B1(P2_REG2_REG_25__SCAN_IN), 
        .B2(n14738), .ZN(n14564) );
  OAI211_X1 U16551 ( .C1(n14860), .C2(n14698), .A(n14565), .B(n14564), .ZN(
        n14566) );
  AOI21_X1 U16552 ( .B1(n14723), .B2(n14765), .A(n14566), .ZN(n14567) );
  OAI21_X1 U16553 ( .B1(n14762), .B2(n14738), .A(n14567), .ZN(P2_U3240) );
  XNOR2_X1 U16554 ( .A(n14568), .B(n14569), .ZN(n14571) );
  AOI21_X1 U16555 ( .B1(n14571), .B2(n14675), .A(n14570), .ZN(n14771) );
  INV_X1 U16556 ( .A(n14572), .ZN(n14573) );
  AOI211_X1 U16557 ( .C1(n14769), .C2(n14596), .A(n14717), .B(n14573), .ZN(
        n14768) );
  INV_X1 U16558 ( .A(n14574), .ZN(n14575) );
  AOI22_X1 U16559 ( .A1(n14575), .A2(n14713), .B1(P2_REG2_REG_24__SCAN_IN), 
        .B2(n14738), .ZN(n14576) );
  OAI21_X1 U16560 ( .B1(n6952), .B2(n14698), .A(n14576), .ZN(n14582) );
  OR2_X1 U16561 ( .A1(n14578), .A2(n14577), .ZN(n14579) );
  NAND2_X1 U16562 ( .A1(n14580), .A2(n14579), .ZN(n14772) );
  NOR2_X1 U16563 ( .A1(n14772), .A2(n14742), .ZN(n14581) );
  AOI211_X1 U16564 ( .C1(n14768), .C2(n14703), .A(n14582), .B(n14581), .ZN(
        n14583) );
  OAI21_X1 U16565 ( .B1(n14719), .B2(n14771), .A(n14583), .ZN(P2_U3241) );
  XNOR2_X1 U16566 ( .A(n14584), .B(n14592), .ZN(n14587) );
  INV_X1 U16567 ( .A(n14585), .ZN(n14586) );
  AOI21_X1 U16568 ( .B1(n14587), .B2(n14675), .A(n14586), .ZN(n14775) );
  NAND2_X1 U16569 ( .A1(n14589), .A2(n14588), .ZN(n14610) );
  INV_X1 U16570 ( .A(n14604), .ZN(n14609) );
  INV_X1 U16571 ( .A(n14590), .ZN(n14591) );
  NAND2_X1 U16572 ( .A1(n14612), .A2(n14591), .ZN(n14594) );
  INV_X1 U16573 ( .A(n14592), .ZN(n14593) );
  XNOR2_X1 U16574 ( .A(n14594), .B(n14593), .ZN(n14773) );
  OAI211_X1 U16575 ( .C1(n14595), .C2(n14865), .A(n14818), .B(n14596), .ZN(
        n14774) );
  INV_X1 U16576 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n14597) );
  OAI22_X1 U16577 ( .A1(n14598), .A2(n14736), .B1(n14597), .B2(n6548), .ZN(
        n14599) );
  AOI21_X1 U16578 ( .B1(n14600), .B2(n14739), .A(n14599), .ZN(n14601) );
  OAI21_X1 U16579 ( .B1(n14774), .B2(n14721), .A(n14601), .ZN(n14602) );
  AOI21_X1 U16580 ( .B1(n14773), .B2(n14723), .A(n14602), .ZN(n14603) );
  OAI21_X1 U16581 ( .B1(n14719), .B2(n14775), .A(n14603), .ZN(P2_U3242) );
  AOI21_X1 U16582 ( .B1(n14605), .B2(n14604), .A(n8640), .ZN(n14608) );
  AOI21_X1 U16583 ( .B1(n14608), .B2(n14607), .A(n14606), .ZN(n14780) );
  NAND2_X1 U16584 ( .A1(n14610), .A2(n14609), .ZN(n14611) );
  NAND2_X1 U16585 ( .A1(n14612), .A2(n14611), .ZN(n14781) );
  INV_X1 U16586 ( .A(n14781), .ZN(n14621) );
  OAI21_X1 U16587 ( .B1(n6610), .B2(n14869), .A(n14818), .ZN(n14613) );
  OR2_X1 U16588 ( .A1(n14613), .A2(n14595), .ZN(n14779) );
  INV_X1 U16589 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n14615) );
  OAI22_X1 U16590 ( .A1(n14616), .A2(n14736), .B1(n14615), .B2(n6548), .ZN(
        n14617) );
  AOI21_X1 U16591 ( .B1(n14618), .B2(n14739), .A(n14617), .ZN(n14619) );
  OAI21_X1 U16592 ( .B1(n14779), .B2(n14721), .A(n14619), .ZN(n14620) );
  AOI21_X1 U16593 ( .B1(n14621), .B2(n14723), .A(n14620), .ZN(n14622) );
  OAI21_X1 U16594 ( .B1(n14719), .B2(n14780), .A(n14622), .ZN(P2_U3243) );
  XOR2_X1 U16595 ( .A(n14623), .B(n14626), .Z(n14625) );
  OAI21_X1 U16596 ( .B1(n14625), .B2(n8640), .A(n14624), .ZN(n14784) );
  INV_X1 U16597 ( .A(n14784), .ZN(n14636) );
  XNOR2_X1 U16598 ( .A(n14627), .B(n14626), .ZN(n14786) );
  NAND2_X1 U16599 ( .A1(n14639), .A2(n14628), .ZN(n14629) );
  NAND2_X1 U16600 ( .A1(n14629), .A2(n14818), .ZN(n14630) );
  NOR2_X1 U16601 ( .A1(n6610), .A2(n14630), .ZN(n14785) );
  NAND2_X1 U16602 ( .A1(n14785), .A2(n14703), .ZN(n14633) );
  AOI22_X1 U16603 ( .A1(n14631), .A2(n14713), .B1(n14719), .B2(
        P2_REG2_REG_21__SCAN_IN), .ZN(n14632) );
  OAI211_X1 U16604 ( .C1(n7905), .C2(n14698), .A(n14633), .B(n14632), .ZN(
        n14634) );
  AOI21_X1 U16605 ( .B1(n14786), .B2(n14723), .A(n14634), .ZN(n14635) );
  OAI21_X1 U16606 ( .B1(n14636), .B2(n14719), .A(n14635), .ZN(P2_U3244) );
  XNOR2_X1 U16607 ( .A(n14637), .B(n14646), .ZN(n14793) );
  INV_X1 U16608 ( .A(n14639), .ZN(n14640) );
  AOI211_X1 U16609 ( .C1(n14790), .C2(n14638), .A(n14717), .B(n14640), .ZN(
        n14789) );
  INV_X1 U16610 ( .A(n14790), .ZN(n14644) );
  INV_X1 U16611 ( .A(n14641), .ZN(n14642) );
  AOI22_X1 U16612 ( .A1(P2_REG2_REG_20__SCAN_IN), .A2(n14719), .B1(n14642), 
        .B2(n14713), .ZN(n14643) );
  OAI21_X1 U16613 ( .B1(n14644), .B2(n14698), .A(n14643), .ZN(n14653) );
  NAND3_X1 U16614 ( .A1(n14645), .A2(n7666), .A3(n14647), .ZN(n14648) );
  AOI21_X1 U16615 ( .B1(n14649), .B2(n14648), .A(n8640), .ZN(n14651) );
  NOR2_X1 U16616 ( .A1(n14651), .A2(n14650), .ZN(n14792) );
  NOR2_X1 U16617 ( .A1(n14792), .A2(n14719), .ZN(n14652) );
  AOI211_X1 U16618 ( .C1(n14789), .C2(n14703), .A(n14653), .B(n14652), .ZN(
        n14654) );
  OAI21_X1 U16619 ( .B1(n14742), .B2(n14793), .A(n14654), .ZN(P2_U3245) );
  XOR2_X1 U16620 ( .A(n14655), .B(n14657), .Z(n14796) );
  INV_X1 U16621 ( .A(n14796), .ZN(n14666) );
  OAI21_X1 U16622 ( .B1(n14657), .B2(n14656), .A(n14645), .ZN(n14658) );
  AND2_X1 U16623 ( .A1(n14658), .A2(n14675), .ZN(n14795) );
  OAI211_X1 U16624 ( .C1(n14877), .C2(n14676), .A(n14638), .B(n14818), .ZN(
        n14660) );
  NAND2_X1 U16625 ( .A1(n14660), .A2(n14659), .ZN(n14794) );
  NAND2_X1 U16626 ( .A1(n14794), .A2(n14703), .ZN(n14663) );
  AOI22_X1 U16627 ( .A1(n14719), .A2(P2_REG2_REG_19__SCAN_IN), .B1(n14661), 
        .B2(n14713), .ZN(n14662) );
  OAI211_X1 U16628 ( .C1(n14877), .C2(n14698), .A(n14663), .B(n14662), .ZN(
        n14664) );
  AOI21_X1 U16629 ( .B1(n14795), .B2(n6548), .A(n14664), .ZN(n14665) );
  OAI21_X1 U16630 ( .B1(n14666), .B2(n14742), .A(n14665), .ZN(P2_U3246) );
  XNOR2_X1 U16631 ( .A(n14667), .B(n14671), .ZN(n14674) );
  INV_X1 U16632 ( .A(n14668), .ZN(n14669) );
  AOI21_X1 U16633 ( .B1(n14671), .B2(n14670), .A(n14669), .ZN(n14803) );
  NOR2_X1 U16634 ( .A1(n14803), .A2(n10420), .ZN(n14672) );
  AOI211_X1 U16635 ( .C1(n14675), .C2(n14674), .A(n14673), .B(n14672), .ZN(
        n14802) );
  INV_X1 U16636 ( .A(n14696), .ZN(n14677) );
  AOI211_X1 U16637 ( .C1(n14800), .C2(n14677), .A(n14717), .B(n14676), .ZN(
        n14799) );
  INV_X1 U16638 ( .A(n14678), .ZN(n14679) );
  AOI22_X1 U16639 ( .A1(n14719), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n14679), 
        .B2(n14713), .ZN(n14680) );
  OAI21_X1 U16640 ( .B1(n14681), .B2(n14698), .A(n14680), .ZN(n14684) );
  NOR2_X1 U16641 ( .A1(n14803), .A2(n14682), .ZN(n14683) );
  AOI211_X1 U16642 ( .C1(n14799), .C2(n14703), .A(n14684), .B(n14683), .ZN(
        n14685) );
  OAI21_X1 U16643 ( .B1(n14802), .B2(n14719), .A(n14685), .ZN(P2_U3247) );
  NOR2_X1 U16644 ( .A1(n6574), .A2(n14686), .ZN(n14709) );
  INV_X1 U16645 ( .A(n14716), .ZN(n14708) );
  OAI21_X1 U16646 ( .B1(n14709), .B2(n14708), .A(n14687), .ZN(n14688) );
  XNOR2_X1 U16647 ( .A(n14688), .B(n14695), .ZN(n14690) );
  OAI21_X1 U16648 ( .B1(n14690), .B2(n8640), .A(n14689), .ZN(n14804) );
  INV_X1 U16649 ( .A(n14804), .ZN(n14706) );
  NAND2_X1 U16650 ( .A1(n14692), .A2(n14691), .ZN(n14715) );
  NOR2_X1 U16651 ( .A1(n14715), .A2(n14716), .ZN(n14714) );
  NOR2_X1 U16652 ( .A1(n14714), .A2(n14693), .ZN(n14694) );
  XOR2_X1 U16653 ( .A(n14695), .B(n14694), .Z(n14806) );
  NAND2_X1 U16654 ( .A1(n14806), .A2(n14723), .ZN(n14705) );
  AOI211_X1 U16655 ( .C1(n14697), .C2(n7989), .A(n14717), .B(n14696), .ZN(
        n14805) );
  NOR2_X1 U16656 ( .A1(n14882), .A2(n14698), .ZN(n14702) );
  INV_X1 U16657 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n14700) );
  OAI22_X1 U16658 ( .A1(n6548), .A2(n14700), .B1(n14699), .B2(n14736), .ZN(
        n14701) );
  AOI211_X1 U16659 ( .C1(n14805), .C2(n14703), .A(n14702), .B(n14701), .ZN(
        n14704) );
  OAI211_X1 U16660 ( .C1(n14738), .C2(n14706), .A(n14705), .B(n14704), .ZN(
        P2_U3248) );
  INV_X1 U16661 ( .A(n14707), .ZN(n14712) );
  INV_X1 U16662 ( .A(n14810), .ZN(n14711) );
  XNOR2_X1 U16663 ( .A(n14709), .B(n14708), .ZN(n14710) );
  NOR2_X1 U16664 ( .A1(n14710), .A2(n8640), .ZN(n14812) );
  AOI211_X1 U16665 ( .C1(n14713), .C2(n14712), .A(n14711), .B(n14812), .ZN(
        n14725) );
  AOI21_X1 U16666 ( .B1(n14716), .B2(n14715), .A(n14714), .ZN(n14814) );
  AOI21_X1 U16667 ( .B1(n14731), .B2(n14809), .A(n14717), .ZN(n14718) );
  NAND2_X1 U16668 ( .A1(n14718), .A2(n7989), .ZN(n14811) );
  AOI22_X1 U16669 ( .A1(n14809), .A2(n14739), .B1(n14719), .B2(
        P2_REG2_REG_16__SCAN_IN), .ZN(n14720) );
  OAI21_X1 U16670 ( .B1(n14811), .B2(n14721), .A(n14720), .ZN(n14722) );
  AOI21_X1 U16671 ( .B1(n14814), .B2(n14723), .A(n14722), .ZN(n14724) );
  OAI21_X1 U16672 ( .B1(n14725), .B2(n14738), .A(n14724), .ZN(P2_U3249) );
  XNOR2_X1 U16673 ( .A(n14726), .B(n8306), .ZN(n14822) );
  AOI211_X1 U16674 ( .C1(n8306), .C2(n14727), .A(n8640), .B(n6574), .ZN(n14729) );
  NOR2_X1 U16675 ( .A1(n14729), .A2(n14728), .ZN(n14821) );
  INV_X1 U16676 ( .A(n14730), .ZN(n14732) );
  AOI21_X1 U16677 ( .B1(n14817), .B2(n14732), .A(n7115), .ZN(n14819) );
  NAND2_X1 U16678 ( .A1(n14819), .A2(n14733), .ZN(n14734) );
  OAI211_X1 U16679 ( .C1(n14736), .C2(n14735), .A(n14821), .B(n14734), .ZN(
        n14737) );
  NAND2_X1 U16680 ( .A1(n14737), .A2(n6548), .ZN(n14741) );
  AOI22_X1 U16681 ( .A1(n14817), .A2(n14739), .B1(P2_REG2_REG_15__SCAN_IN), 
        .B2(n14738), .ZN(n14740) );
  OAI211_X1 U16682 ( .C1(n14822), .C2(n14742), .A(n14741), .B(n14740), .ZN(
        P2_U3250) );
  MUX2_X1 U16683 ( .A(P2_REG1_REG_29__SCAN_IN), .B(n14850), .S(n16011), .Z(
        P2_U3528) );
  INV_X1 U16684 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n14755) );
  NAND3_X1 U16685 ( .A1(n14535), .A2(n14748), .A3(n15993), .ZN(n14752) );
  NAND2_X1 U16686 ( .A1(n14749), .A2(n15996), .ZN(n14751) );
  NAND3_X1 U16687 ( .A1(n14752), .A2(n14751), .A3(n14750), .ZN(n14753) );
  MUX2_X1 U16688 ( .A(n14755), .B(n14854), .S(n16011), .Z(n14756) );
  INV_X1 U16689 ( .A(n14756), .ZN(P2_U3526) );
  OAI21_X1 U16690 ( .B1(n14759), .B2(n15989), .A(n14758), .ZN(n14760) );
  MUX2_X1 U16691 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n14856), .S(n16011), .Z(
        P2_U3525) );
  INV_X1 U16692 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n14766) );
  INV_X1 U16693 ( .A(n14762), .ZN(n14763) );
  MUX2_X1 U16694 ( .A(n14766), .B(n14857), .S(n16011), .Z(n14767) );
  OAI21_X1 U16695 ( .B1(n14860), .B2(n14840), .A(n14767), .ZN(P2_U3524) );
  AOI21_X1 U16696 ( .B1(n15996), .B2(n14769), .A(n14768), .ZN(n14770) );
  OAI211_X1 U16697 ( .C1(n16000), .C2(n14772), .A(n14771), .B(n14770), .ZN(
        n14861) );
  MUX2_X1 U16698 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n14861), .S(n16011), .Z(
        P2_U3523) );
  NAND2_X1 U16699 ( .A1(n14773), .A2(n15993), .ZN(n14776) );
  NAND3_X1 U16700 ( .A1(n14776), .A2(n14775), .A3(n14774), .ZN(n14862) );
  MUX2_X1 U16701 ( .A(n14862), .B(P2_REG1_REG_23__SCAN_IN), .S(n16008), .Z(
        n14777) );
  INV_X1 U16702 ( .A(n14777), .ZN(n14778) );
  OAI21_X1 U16703 ( .B1(n14865), .B2(n14840), .A(n14778), .ZN(P2_U3522) );
  OAI211_X1 U16704 ( .C1(n14781), .C2(n16000), .A(n14780), .B(n14779), .ZN(
        n14866) );
  MUX2_X1 U16705 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n14866), .S(n16011), .Z(
        n14782) );
  INV_X1 U16706 ( .A(n14782), .ZN(n14783) );
  OAI21_X1 U16707 ( .B1(n14869), .B2(n14840), .A(n14783), .ZN(P2_U3521) );
  AOI211_X1 U16708 ( .C1(n15993), .C2(n14786), .A(n14785), .B(n14784), .ZN(
        n14870) );
  MUX2_X1 U16709 ( .A(n14787), .B(n14870), .S(n16011), .Z(n14788) );
  OAI21_X1 U16710 ( .B1(n7905), .B2(n14840), .A(n14788), .ZN(P2_U3520) );
  AOI21_X1 U16711 ( .B1(n15996), .B2(n14790), .A(n14789), .ZN(n14791) );
  OAI211_X1 U16712 ( .C1(n14793), .C2(n16000), .A(n14792), .B(n14791), .ZN(
        n14873) );
  MUX2_X1 U16713 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n14873), .S(n16011), .Z(
        P2_U3519) );
  INV_X1 U16714 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n14797) );
  AOI211_X1 U16715 ( .C1(n14796), .C2(n15993), .A(n14795), .B(n14794), .ZN(
        n14874) );
  MUX2_X1 U16716 ( .A(n14797), .B(n14874), .S(n16011), .Z(n14798) );
  OAI21_X1 U16717 ( .B1(n14877), .B2(n14840), .A(n14798), .ZN(P2_U3518) );
  AOI21_X1 U16718 ( .B1(n15996), .B2(n14800), .A(n14799), .ZN(n14801) );
  OAI211_X1 U16719 ( .C1(n14803), .C2(n14846), .A(n14802), .B(n14801), .ZN(
        n14878) );
  MUX2_X1 U16720 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n14878), .S(n16011), .Z(
        P2_U3517) );
  AOI211_X1 U16721 ( .C1(n14806), .C2(n15993), .A(n14805), .B(n14804), .ZN(
        n14879) );
  MUX2_X1 U16722 ( .A(n14807), .B(n14879), .S(n16011), .Z(n14808) );
  OAI21_X1 U16723 ( .B1(n14882), .B2(n14840), .A(n14808), .ZN(P2_U3516) );
  NAND2_X1 U16724 ( .A1(n14811), .A2(n14810), .ZN(n14813) );
  AOI211_X1 U16725 ( .C1(n14814), .C2(n15993), .A(n14813), .B(n14812), .ZN(
        n14883) );
  MUX2_X1 U16726 ( .A(n14815), .B(n14883), .S(n16011), .Z(n14816) );
  OAI21_X1 U16727 ( .B1(n7114), .B2(n14840), .A(n14816), .ZN(P2_U3515) );
  AOI22_X1 U16728 ( .A1(n14819), .A2(n14818), .B1(n15996), .B2(n14817), .ZN(
        n14820) );
  OAI211_X1 U16729 ( .C1(n16000), .C2(n14822), .A(n14821), .B(n14820), .ZN(
        n14886) );
  MUX2_X1 U16730 ( .A(P2_REG1_REG_15__SCAN_IN), .B(n14886), .S(n16011), .Z(
        P2_U3514) );
  AOI21_X1 U16731 ( .B1(n15996), .B2(n14824), .A(n14823), .ZN(n14825) );
  OAI211_X1 U16732 ( .C1(n14827), .C2(n16000), .A(n14826), .B(n14825), .ZN(
        n14887) );
  MUX2_X1 U16733 ( .A(P2_REG1_REG_14__SCAN_IN), .B(n14887), .S(n16011), .Z(
        P2_U3513) );
  AOI21_X1 U16734 ( .B1(n15996), .B2(n14829), .A(n14828), .ZN(n14830) );
  OAI211_X1 U16735 ( .C1(n14832), .C2(n14846), .A(n14831), .B(n14830), .ZN(
        n14888) );
  MUX2_X1 U16736 ( .A(P2_REG1_REG_12__SCAN_IN), .B(n14888), .S(n16011), .Z(
        P2_U3511) );
  INV_X1 U16737 ( .A(n14833), .ZN(n14836) );
  AOI211_X1 U16738 ( .C1(n14837), .C2(n14836), .A(n14835), .B(n14834), .ZN(
        n14889) );
  MUX2_X1 U16739 ( .A(n14838), .B(n14889), .S(n16011), .Z(n14839) );
  OAI21_X1 U16740 ( .B1(n14893), .B2(n14840), .A(n14839), .ZN(P2_U3510) );
  AOI21_X1 U16741 ( .B1(n15996), .B2(n14842), .A(n14841), .ZN(n14843) );
  OAI211_X1 U16742 ( .C1(n14846), .C2(n14845), .A(n14844), .B(n14843), .ZN(
        n14894) );
  MUX2_X1 U16743 ( .A(P2_REG1_REG_10__SCAN_IN), .B(n14894), .S(n16011), .Z(
        P2_U3509) );
  OAI21_X1 U16744 ( .B1(n14849), .B2(n14892), .A(n14848), .ZN(P2_U3498) );
  MUX2_X1 U16745 ( .A(P2_REG0_REG_29__SCAN_IN), .B(n14850), .S(n16004), .Z(
        P2_U3496) );
  MUX2_X1 U16746 ( .A(n14856), .B(P2_REG0_REG_26__SCAN_IN), .S(n16002), .Z(
        P2_U3493) );
  MUX2_X1 U16747 ( .A(n14858), .B(n14857), .S(n16004), .Z(n14859) );
  OAI21_X1 U16748 ( .B1(n14860), .B2(n14892), .A(n14859), .ZN(P2_U3492) );
  MUX2_X1 U16749 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n14861), .S(n16004), .Z(
        P2_U3491) );
  MUX2_X1 U16750 ( .A(n14862), .B(P2_REG0_REG_23__SCAN_IN), .S(n16002), .Z(
        n14863) );
  INV_X1 U16751 ( .A(n14863), .ZN(n14864) );
  OAI21_X1 U16752 ( .B1(n14865), .B2(n14892), .A(n14864), .ZN(P2_U3490) );
  MUX2_X1 U16753 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n14866), .S(n16004), .Z(
        n14867) );
  INV_X1 U16754 ( .A(n14867), .ZN(n14868) );
  OAI21_X1 U16755 ( .B1(n14869), .B2(n14892), .A(n14868), .ZN(P2_U3489) );
  INV_X1 U16756 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n14871) );
  MUX2_X1 U16757 ( .A(n14871), .B(n14870), .S(n16004), .Z(n14872) );
  OAI21_X1 U16758 ( .B1(n7905), .B2(n14892), .A(n14872), .ZN(P2_U3488) );
  MUX2_X1 U16759 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n14873), .S(n16004), .Z(
        P2_U3487) );
  INV_X1 U16760 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n14875) );
  MUX2_X1 U16761 ( .A(n14875), .B(n14874), .S(n16004), .Z(n14876) );
  OAI21_X1 U16762 ( .B1(n14877), .B2(n14892), .A(n14876), .ZN(P2_U3486) );
  MUX2_X1 U16763 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n14878), .S(n16004), .Z(
        P2_U3484) );
  INV_X1 U16764 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n14880) );
  MUX2_X1 U16765 ( .A(n14880), .B(n14879), .S(n16004), .Z(n14881) );
  OAI21_X1 U16766 ( .B1(n14882), .B2(n14892), .A(n14881), .ZN(P2_U3481) );
  MUX2_X1 U16767 ( .A(n14884), .B(n14883), .S(n16004), .Z(n14885) );
  OAI21_X1 U16768 ( .B1(n7114), .B2(n14892), .A(n14885), .ZN(P2_U3478) );
  MUX2_X1 U16769 ( .A(P2_REG0_REG_15__SCAN_IN), .B(n14886), .S(n16004), .Z(
        P2_U3475) );
  MUX2_X1 U16770 ( .A(P2_REG0_REG_14__SCAN_IN), .B(n14887), .S(n16004), .Z(
        P2_U3472) );
  MUX2_X1 U16771 ( .A(P2_REG0_REG_12__SCAN_IN), .B(n14888), .S(n16004), .Z(
        P2_U3466) );
  MUX2_X1 U16772 ( .A(n14890), .B(n14889), .S(n16004), .Z(n14891) );
  OAI21_X1 U16773 ( .B1(n14893), .B2(n14892), .A(n14891), .ZN(P2_U3463) );
  MUX2_X1 U16774 ( .A(P2_REG0_REG_10__SCAN_IN), .B(n14894), .S(n16004), .Z(
        P2_U3460) );
  INV_X1 U16775 ( .A(n14895), .ZN(n15693) );
  NOR4_X1 U16776 ( .A1(n7310), .A2(P2_IR_REG_30__SCAN_IN), .A3(n8006), .A4(
        P2_U3088), .ZN(n14896) );
  AOI21_X1 U16777 ( .B1(n14897), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n14896), 
        .ZN(n14898) );
  OAI21_X1 U16778 ( .B1(n15693), .B2(n14917), .A(n14898), .ZN(P2_U3296) );
  OAI222_X1 U16779 ( .A1(n14917), .A2(n14901), .B1(P2_U3088), .B2(n14899), 
        .C1(n14900), .C2(n14914), .ZN(P2_U3297) );
  INV_X1 U16780 ( .A(n14902), .ZN(n15695) );
  OAI222_X1 U16781 ( .A1(n14914), .A2(n14905), .B1(P2_U3088), .B2(n14904), 
        .C1(n14903), .C2(n15695), .ZN(P2_U3298) );
  NAND2_X1 U16782 ( .A1(n14907), .A2(n14906), .ZN(n14909) );
  OAI211_X1 U16783 ( .C1(n14914), .C2(n14910), .A(n14909), .B(n14908), .ZN(
        P2_U3299) );
  INV_X1 U16784 ( .A(n14911), .ZN(n15698) );
  OAI222_X1 U16785 ( .A1(n14914), .A2(n14913), .B1(n14917), .B2(n15698), .C1(
        n14912), .C2(P2_U3088), .ZN(P2_U3300) );
  INV_X1 U16786 ( .A(n14915), .ZN(n15702) );
  INV_X1 U16787 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n14916) );
  OAI222_X1 U16788 ( .A1(P2_U3088), .A2(n14918), .B1(n14917), .B2(n15702), 
        .C1(n14916), .C2(n14914), .ZN(P2_U3301) );
  INV_X1 U16789 ( .A(n14920), .ZN(n14921) );
  MUX2_X1 U16790 ( .A(n14921), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3327) );
  XNOR2_X1 U16791 ( .A(n14923), .B(n14922), .ZN(n14930) );
  AOI22_X1 U16792 ( .A1(n14924), .A2(n15061), .B1(P1_REG3_REG_27__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14926) );
  NAND2_X1 U16793 ( .A1(n15086), .A2(n15062), .ZN(n14925) );
  OAI211_X1 U16794 ( .C1(n14927), .C2(n15065), .A(n14926), .B(n14925), .ZN(
        n14928) );
  AOI21_X1 U16795 ( .B1(n7122), .B2(n15068), .A(n14928), .ZN(n14929) );
  OAI21_X1 U16796 ( .B1(n14930), .B2(n15070), .A(n14929), .ZN(P1_U3214) );
  INV_X1 U16797 ( .A(n14931), .ZN(n14932) );
  AOI21_X1 U16798 ( .B1(n14934), .B2(n14933), .A(n14932), .ZN(n14940) );
  NOR2_X1 U16799 ( .A1(n14935), .A2(P1_STATE_REG_SCAN_IN), .ZN(n15190) );
  AOI21_X1 U16800 ( .B1(n15062), .B2(n15502), .A(n15190), .ZN(n14937) );
  NAND2_X1 U16801 ( .A1(n15061), .A2(n15508), .ZN(n14936) );
  OAI211_X1 U16802 ( .C1(n14993), .C2(n15065), .A(n14937), .B(n14936), .ZN(
        n14938) );
  AOI21_X1 U16803 ( .B1(n15639), .B2(n15068), .A(n14938), .ZN(n14939) );
  OAI21_X1 U16804 ( .B1(n14940), .B2(n15070), .A(n14939), .ZN(P1_U3215) );
  XOR2_X1 U16805 ( .A(n14942), .B(n14941), .Z(n14948) );
  NAND2_X1 U16806 ( .A1(n15306), .A2(n15500), .ZN(n14944) );
  NAND2_X1 U16807 ( .A1(n15087), .A2(n15521), .ZN(n14943) );
  AND2_X1 U16808 ( .A1(n14944), .A2(n14943), .ZN(n15583) );
  AOI22_X1 U16809 ( .A1(n15349), .A2(n15061), .B1(P1_REG3_REG_23__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14945) );
  OAI21_X1 U16810 ( .B1(n15583), .B2(n15025), .A(n14945), .ZN(n14946) );
  AOI21_X1 U16811 ( .B1(n15586), .B2(n15068), .A(n14946), .ZN(n14947) );
  OAI21_X1 U16812 ( .B1(n14948), .B2(n15070), .A(n14947), .ZN(P1_U3216) );
  OAI211_X1 U16813 ( .C1(n14951), .C2(n14950), .A(n14949), .B(n15072), .ZN(
        n14956) );
  NOR2_X1 U16814 ( .A1(n15077), .A2(n15422), .ZN(n14954) );
  NAND2_X1 U16815 ( .A1(P1_U3086), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n15251)
         );
  OAI21_X1 U16816 ( .B1(n15056), .B2(n14952), .A(n15251), .ZN(n14953) );
  AOI211_X1 U16817 ( .C1(n15053), .C2(n15421), .A(n14954), .B(n14953), .ZN(
        n14955) );
  OAI211_X1 U16818 ( .C1(n7456), .C2(n15083), .A(n14956), .B(n14955), .ZN(
        P1_U3219) );
  INV_X1 U16819 ( .A(n14957), .ZN(n14958) );
  AOI21_X1 U16820 ( .B1(n14960), .B2(n14959), .A(n14958), .ZN(n14966) );
  OAI22_X1 U16821 ( .A1(n15390), .A2(n15056), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14961), .ZN(n14962) );
  AOI21_X1 U16822 ( .B1(n15087), .B2(n15053), .A(n14962), .ZN(n14963) );
  OAI21_X1 U16823 ( .B1(n15077), .B2(n15394), .A(n14963), .ZN(n14964) );
  AOI21_X1 U16824 ( .B1(n15597), .B2(n15068), .A(n14964), .ZN(n14965) );
  OAI21_X1 U16825 ( .B1(n14966), .B2(n15070), .A(n14965), .ZN(P1_U3223) );
  AND2_X1 U16826 ( .A1(n14969), .A2(n14967), .ZN(n14972) );
  NAND2_X1 U16827 ( .A1(n14969), .A2(n14968), .ZN(n14970) );
  OAI211_X1 U16828 ( .C1(n14972), .C2(n14971), .A(n14970), .B(n15072), .ZN(
        n14977) );
  NOR2_X1 U16829 ( .A1(n15077), .A2(n14973), .ZN(n14974) );
  AOI211_X1 U16830 ( .C1(n15080), .C2(n15650), .A(n14975), .B(n14974), .ZN(
        n14976) );
  OAI211_X1 U16831 ( .C1(n14978), .C2(n15083), .A(n14977), .B(n14976), .ZN(
        P1_U3224) );
  AOI22_X1 U16832 ( .A1(n15086), .A2(n15500), .B1(n15521), .B2(n15306), .ZN(
        n15570) );
  NOR2_X1 U16833 ( .A1(n15570), .A2(n15025), .ZN(n14983) );
  OAI22_X1 U16834 ( .A1(n15314), .A2(n15077), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14981), .ZN(n14982) );
  AOI211_X1 U16835 ( .C1(n15318), .C2(n15068), .A(n14983), .B(n14982), .ZN(
        n14984) );
  XNOR2_X1 U16836 ( .A(n14986), .B(n14985), .ZN(n14992) );
  XNOR2_X1 U16837 ( .A(n14989), .B(n14987), .ZN(n15075) );
  INV_X1 U16838 ( .A(n14988), .ZN(n15074) );
  NAND2_X1 U16839 ( .A1(n15075), .A2(n15074), .ZN(n15073) );
  OAI21_X1 U16840 ( .B1(n14990), .B2(n14989), .A(n15073), .ZN(n14991) );
  NOR2_X1 U16841 ( .A1(n14991), .A2(n14992), .ZN(n15002) );
  AOI21_X1 U16842 ( .B1(n14992), .B2(n14991), .A(n15002), .ZN(n14998) );
  OAI22_X1 U16843 ( .A1(n15432), .A2(n15516), .B1(n14993), .B2(n15431), .ZN(
        n15627) );
  AOI21_X1 U16844 ( .B1(n15627), .B2(n15080), .A(n14994), .ZN(n14995) );
  OAI21_X1 U16845 ( .B1(n15077), .B2(n15472), .A(n14995), .ZN(n14996) );
  AOI21_X1 U16846 ( .B1(n15628), .B2(n15068), .A(n14996), .ZN(n14997) );
  OAI21_X1 U16847 ( .B1(n14998), .B2(n15070), .A(n14997), .ZN(P1_U3226) );
  INV_X1 U16848 ( .A(n14999), .ZN(n15001) );
  NOR3_X1 U16849 ( .A1(n15002), .A2(n15001), .A3(n15000), .ZN(n15005) );
  INV_X1 U16850 ( .A(n15003), .ZN(n15004) );
  OAI21_X1 U16851 ( .B1(n15005), .B2(n15004), .A(n15072), .ZN(n15010) );
  INV_X1 U16852 ( .A(n15457), .ZN(n15008) );
  AND2_X1 U16853 ( .A1(n15090), .A2(n15521), .ZN(n15006) );
  AOI21_X1 U16854 ( .B1(n15419), .B2(n15500), .A(n15006), .ZN(n15452) );
  NAND2_X1 U16855 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n15203)
         );
  OAI21_X1 U16856 ( .B1(n15452), .B2(n15025), .A(n15203), .ZN(n15007) );
  AOI21_X1 U16857 ( .B1(n15008), .B2(n15061), .A(n15007), .ZN(n15009) );
  OAI211_X1 U16858 ( .C1(n15459), .C2(n15083), .A(n15010), .B(n15009), .ZN(
        P1_U3228) );
  XOR2_X1 U16859 ( .A(n15011), .B(n15012), .Z(n15018) );
  NAND2_X1 U16860 ( .A1(n15330), .A2(n15053), .ZN(n15015) );
  INV_X1 U16861 ( .A(n15013), .ZN(n15340) );
  AOI22_X1 U16862 ( .A1(n15340), .A2(n15061), .B1(P1_REG3_REG_24__SCAN_IN), 
        .B2(P1_U3086), .ZN(n15014) );
  OAI211_X1 U16863 ( .C1(n15332), .C2(n15056), .A(n15015), .B(n15014), .ZN(
        n15016) );
  AOI21_X1 U16864 ( .B1(n15341), .B2(n15068), .A(n15016), .ZN(n15017) );
  OAI21_X1 U16865 ( .B1(n15018), .B2(n15070), .A(n15017), .ZN(P1_U3229) );
  OAI211_X1 U16866 ( .C1(n15021), .C2(n15020), .A(n15019), .B(n15072), .ZN(
        n15028) );
  INV_X1 U16867 ( .A(n15022), .ZN(n15410) );
  AND2_X1 U16868 ( .A1(n15088), .A2(n15521), .ZN(n15023) );
  AOI21_X1 U16869 ( .B1(n15363), .B2(n15500), .A(n15023), .ZN(n15406) );
  OAI22_X1 U16870 ( .A1(n15406), .A2(n15025), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n15024), .ZN(n15026) );
  AOI21_X1 U16871 ( .B1(n15410), .B2(n15061), .A(n15026), .ZN(n15027) );
  OAI211_X1 U16872 ( .C1(n7457), .C2(n15083), .A(n15028), .B(n15027), .ZN(
        P1_U3233) );
  AND2_X1 U16873 ( .A1(n15030), .A2(n15029), .ZN(n15033) );
  OAI211_X1 U16874 ( .C1(n15033), .C2(n15032), .A(n15031), .B(n15072), .ZN(
        n15039) );
  INV_X1 U16875 ( .A(n15034), .ZN(n15524) );
  NAND2_X1 U16876 ( .A1(n15062), .A2(n15520), .ZN(n15036) );
  OAI211_X1 U16877 ( .C1(n15517), .C2(n15065), .A(n15036), .B(n15035), .ZN(
        n15037) );
  AOI21_X1 U16878 ( .B1(n15524), .B2(n15061), .A(n15037), .ZN(n15038) );
  OAI211_X1 U16879 ( .C1(n15530), .C2(n15083), .A(n15039), .B(n15038), .ZN(
        P1_U3234) );
  OAI21_X1 U16880 ( .B1(n15042), .B2(n15041), .A(n15040), .ZN(n15043) );
  NAND2_X1 U16881 ( .A1(n15043), .A2(n15072), .ZN(n15049) );
  OAI22_X1 U16882 ( .A1(n15045), .A2(n15056), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n15044), .ZN(n15047) );
  NOR2_X1 U16883 ( .A1(n15332), .A2(n15065), .ZN(n15046) );
  AOI211_X1 U16884 ( .C1(n15368), .C2(n15061), .A(n15047), .B(n15046), .ZN(
        n15048) );
  OAI211_X1 U16885 ( .C1(n15083), .C2(n15370), .A(n15049), .B(n15048), .ZN(
        P1_U3235) );
  XOR2_X1 U16886 ( .A(n15050), .B(n15051), .Z(n15059) );
  NOR2_X1 U16887 ( .A1(n15052), .A2(P1_STATE_REG_SCAN_IN), .ZN(n15222) );
  AOI21_X1 U16888 ( .B1(n15088), .B2(n15053), .A(n15222), .ZN(n15055) );
  NAND2_X1 U16889 ( .A1(n15061), .A2(n15442), .ZN(n15054) );
  OAI211_X1 U16890 ( .C1(n15432), .C2(n15056), .A(n15055), .B(n15054), .ZN(
        n15057) );
  AOI21_X1 U16891 ( .B1(n15616), .B2(n15068), .A(n15057), .ZN(n15058) );
  OAI21_X1 U16892 ( .B1(n15059), .B2(n15070), .A(n15058), .ZN(P1_U3238) );
  AOI22_X1 U16893 ( .A1(n15298), .A2(n15061), .B1(P1_REG3_REG_26__SCAN_IN), 
        .B2(P1_U3086), .ZN(n15064) );
  NAND2_X1 U16894 ( .A1(n15330), .A2(n15062), .ZN(n15063) );
  OAI211_X1 U16895 ( .C1(n15066), .C2(n15065), .A(n15064), .B(n15063), .ZN(
        n15067) );
  AOI21_X1 U16896 ( .B1(n15301), .B2(n15068), .A(n15067), .ZN(n15069) );
  OAI21_X1 U16897 ( .B1(n15071), .B2(n15070), .A(n15069), .ZN(P1_U3240) );
  OAI211_X1 U16898 ( .C1(n15075), .C2(n15074), .A(n15073), .B(n15072), .ZN(
        n15082) );
  OAI22_X1 U16899 ( .A1(n15076), .A2(n15516), .B1(n15517), .B2(n15431), .ZN(
        n15487) );
  NOR2_X1 U16900 ( .A1(n15077), .A2(n15492), .ZN(n15078) );
  AOI211_X1 U16901 ( .C1(n15080), .C2(n15487), .A(n15079), .B(n15078), .ZN(
        n15081) );
  OAI211_X1 U16902 ( .C1(n6801), .C2(n15083), .A(n15082), .B(n15081), .ZN(
        P1_U3241) );
  MUX2_X1 U16903 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(n15256), .S(P1_U4016), .Z(
        P1_U3591) );
  MUX2_X1 U16904 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n15084), .S(P1_U4016), .Z(
        P1_U3590) );
  MUX2_X1 U16905 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n15272), .S(P1_U4016), .Z(
        P1_U3589) );
  MUX2_X1 U16906 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n15085), .S(P1_U4016), .Z(
        P1_U3588) );
  MUX2_X1 U16907 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n15297), .S(P1_U4016), .Z(
        P1_U3587) );
  MUX2_X1 U16908 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n15086), .S(P1_U4016), .Z(
        P1_U3586) );
  MUX2_X1 U16909 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n15330), .S(P1_U4016), .Z(
        P1_U3585) );
  MUX2_X1 U16910 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n15306), .S(P1_U4016), .Z(
        P1_U3584) );
  MUX2_X1 U16911 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n15362), .S(P1_U4016), .Z(
        P1_U3583) );
  MUX2_X1 U16912 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n15087), .S(P1_U4016), .Z(
        P1_U3582) );
  MUX2_X1 U16913 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n15363), .S(P1_U4016), .Z(
        P1_U3581) );
  MUX2_X1 U16914 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n15421), .S(n6547), .Z(
        P1_U3580) );
  MUX2_X1 U16915 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n15088), .S(n6547), .Z(
        P1_U3579) );
  MUX2_X1 U16916 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n15419), .S(n6547), .Z(
        P1_U3578) );
  MUX2_X1 U16917 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n15089), .S(n6547), .Z(
        P1_U3577) );
  MUX2_X1 U16918 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n15090), .S(n6547), .Z(
        P1_U3576) );
  MUX2_X1 U16919 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n15501), .S(n6547), .Z(
        P1_U3575) );
  MUX2_X1 U16920 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n15091), .S(n6547), .Z(
        P1_U3574) );
  MUX2_X1 U16921 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n15502), .S(n6547), .Z(
        P1_U3573) );
  MUX2_X1 U16922 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n15520), .S(n6547), .Z(
        P1_U3572) );
  MUX2_X1 U16923 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n15092), .S(n6547), .Z(
        P1_U3571) );
  MUX2_X1 U16924 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n15093), .S(n6547), .Z(
        P1_U3570) );
  MUX2_X1 U16925 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n15094), .S(n6547), .Z(
        P1_U3569) );
  MUX2_X1 U16926 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n15095), .S(n6547), .Z(
        P1_U3568) );
  MUX2_X1 U16927 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n15096), .S(n6547), .Z(
        P1_U3567) );
  MUX2_X1 U16928 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n15097), .S(n6547), .Z(
        P1_U3566) );
  MUX2_X1 U16929 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n15098), .S(n6547), .Z(
        P1_U3565) );
  MUX2_X1 U16930 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n15795), .S(n6547), .Z(
        P1_U3564) );
  MUX2_X1 U16931 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n15099), .S(P1_U4016), .Z(
        P1_U3563) );
  MUX2_X1 U16932 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n10144), .S(P1_U4016), .Z(
        P1_U3562) );
  MUX2_X1 U16933 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n10118), .S(P1_U4016), .Z(
        P1_U3561) );
  MUX2_X1 U16934 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(n7136), .S(P1_U4016), .Z(
        P1_U3560) );
  OAI22_X1 U16935 ( .A1(n15252), .A2(n15101), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n15100), .ZN(n15102) );
  AOI21_X1 U16936 ( .B1(n15223), .B2(n15103), .A(n15102), .ZN(n15111) );
  OAI211_X1 U16937 ( .C1(n15105), .C2(n15112), .A(n15244), .B(n15104), .ZN(
        n15110) );
  OAI211_X1 U16938 ( .C1(n15108), .C2(n15107), .A(n15218), .B(n15106), .ZN(
        n15109) );
  NAND3_X1 U16939 ( .A1(n15111), .A2(n15110), .A3(n15109), .ZN(P1_U3244) );
  INV_X1 U16940 ( .A(n15112), .ZN(n15114) );
  MUX2_X1 U16941 ( .A(n15115), .B(n15114), .S(n15113), .Z(n15120) );
  NAND2_X1 U16942 ( .A1(n15116), .A2(n7444), .ZN(n15117) );
  OAI211_X1 U16943 ( .C1(n15120), .C2(n15119), .A(n6547), .B(n15117), .ZN(
        n15159) );
  OAI22_X1 U16944 ( .A1(n15252), .A2(n15122), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n15121), .ZN(n15123) );
  AOI21_X1 U16945 ( .B1(n15223), .B2(n15124), .A(n15123), .ZN(n15133) );
  OAI211_X1 U16946 ( .C1(n15127), .C2(n15126), .A(n15218), .B(n15125), .ZN(
        n15132) );
  OAI211_X1 U16947 ( .C1(n15130), .C2(n15129), .A(n15244), .B(n15128), .ZN(
        n15131) );
  NAND4_X1 U16948 ( .A1(n15159), .A2(n15133), .A3(n15132), .A4(n15131), .ZN(
        P1_U3245) );
  NAND2_X1 U16949 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_U3086), .ZN(n15134) );
  OAI21_X1 U16950 ( .B1(n15252), .B2(n10629), .A(n15134), .ZN(n15135) );
  AOI21_X1 U16951 ( .B1(n15223), .B2(n15136), .A(n15135), .ZN(n15145) );
  OAI211_X1 U16952 ( .C1(n15139), .C2(n15138), .A(n15218), .B(n15137), .ZN(
        n15144) );
  OAI211_X1 U16953 ( .C1(n15142), .C2(n15141), .A(n15244), .B(n15140), .ZN(
        n15143) );
  NAND3_X1 U16954 ( .A1(n15145), .A2(n15144), .A3(n15143), .ZN(P1_U3246) );
  NOR2_X1 U16955 ( .A1(n15246), .A2(n15146), .ZN(n15147) );
  AOI211_X1 U16956 ( .C1(n15149), .C2(P1_ADDR_REG_4__SCAN_IN), .A(n15148), .B(
        n15147), .ZN(n15158) );
  OAI211_X1 U16957 ( .C1(n15152), .C2(n15151), .A(n15244), .B(n15150), .ZN(
        n15157) );
  OAI211_X1 U16958 ( .C1(n15155), .C2(n15154), .A(n15218), .B(n15153), .ZN(
        n15156) );
  NAND4_X1 U16959 ( .A1(n15159), .A2(n15158), .A3(n15157), .A4(n15156), .ZN(
        P1_U3247) );
  NAND2_X1 U16960 ( .A1(P1_REG3_REG_7__SCAN_IN), .A2(P1_U3086), .ZN(n15160) );
  OAI21_X1 U16961 ( .B1(n15252), .B2(n15161), .A(n15160), .ZN(n15162) );
  AOI21_X1 U16962 ( .B1(n15223), .B2(n15163), .A(n15162), .ZN(n15172) );
  OAI211_X1 U16963 ( .C1(n15166), .C2(n15165), .A(n15244), .B(n15164), .ZN(
        n15171) );
  OAI211_X1 U16964 ( .C1(n15169), .C2(n15168), .A(n15218), .B(n15167), .ZN(
        n15170) );
  NAND3_X1 U16965 ( .A1(n15172), .A2(n15171), .A3(n15170), .ZN(P1_U3250) );
  OAI211_X1 U16966 ( .C1(n15175), .C2(n15174), .A(n15173), .B(n15218), .ZN(
        n15184) );
  NOR2_X1 U16967 ( .A1(n15252), .A2(n12012), .ZN(n15176) );
  AOI211_X1 U16968 ( .C1(n15223), .C2(n15178), .A(n15177), .B(n15176), .ZN(
        n15183) );
  OAI211_X1 U16969 ( .C1(n15181), .C2(n15180), .A(n15179), .B(n15244), .ZN(
        n15182) );
  NAND3_X1 U16970 ( .A1(n15184), .A2(n15183), .A3(n15182), .ZN(P1_U3253) );
  OAI21_X1 U16971 ( .B1(n15187), .B2(n15186), .A(n15185), .ZN(n15188) );
  NAND2_X1 U16972 ( .A1(n15188), .A2(n15218), .ZN(n15197) );
  INV_X1 U16973 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n15725) );
  NOR2_X1 U16974 ( .A1(n15252), .A2(n15725), .ZN(n15189) );
  AOI211_X1 U16975 ( .C1(n15223), .C2(n15191), .A(n15190), .B(n15189), .ZN(
        n15196) );
  OAI211_X1 U16976 ( .C1(n15194), .C2(n15193), .A(n15192), .B(n15244), .ZN(
        n15195) );
  NAND3_X1 U16977 ( .A1(n15197), .A2(n15196), .A3(n15195), .ZN(P1_U3257) );
  NAND2_X1 U16978 ( .A1(n15205), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n15198) );
  NAND2_X1 U16979 ( .A1(n15199), .A2(n15198), .ZN(n15202) );
  INV_X1 U16980 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n15200) );
  XNOR2_X1 U16981 ( .A(n15224), .B(n15200), .ZN(n15201) );
  NAND2_X1 U16982 ( .A1(n15202), .A2(n15201), .ZN(n15216) );
  OAI211_X1 U16983 ( .C1(n15202), .C2(n15201), .A(n15216), .B(n15218), .ZN(
        n15214) );
  INV_X1 U16984 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n15756) );
  OAI21_X1 U16985 ( .B1(n15252), .B2(n15756), .A(n15203), .ZN(n15204) );
  AOI21_X1 U16986 ( .B1(n15223), .B2(n15224), .A(n15204), .ZN(n15213) );
  NAND2_X1 U16987 ( .A1(n15205), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n15206) );
  NAND2_X1 U16988 ( .A1(n15207), .A2(n15206), .ZN(n15211) );
  INV_X1 U16989 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n15209) );
  NAND2_X1 U16990 ( .A1(n15224), .A2(n15209), .ZN(n15208) );
  OAI21_X1 U16991 ( .B1(n15224), .B2(n15209), .A(n15208), .ZN(n15210) );
  NAND2_X1 U16992 ( .A1(n15211), .A2(n15210), .ZN(n15226) );
  OAI211_X1 U16993 ( .C1(n15211), .C2(n15210), .A(n15226), .B(n15244), .ZN(
        n15212) );
  NAND3_X1 U16994 ( .A1(n15214), .A2(n15213), .A3(n15212), .ZN(P1_U3260) );
  NAND2_X1 U16995 ( .A1(n15224), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n15215) );
  NAND2_X1 U16996 ( .A1(n15217), .A2(n15227), .ZN(n15235) );
  OAI211_X1 U16997 ( .C1(n15219), .C2(P1_REG1_REG_18__SCAN_IN), .A(n15236), 
        .B(n15218), .ZN(n15234) );
  INV_X1 U16998 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n15220) );
  NOR2_X1 U16999 ( .A1(n15252), .A2(n15220), .ZN(n15221) );
  AOI211_X1 U17000 ( .C1(n15227), .C2(n15223), .A(n15222), .B(n15221), .ZN(
        n15233) );
  NAND2_X1 U17001 ( .A1(n15224), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n15225) );
  NAND2_X1 U17002 ( .A1(n15226), .A2(n15225), .ZN(n15228) );
  NAND2_X1 U17003 ( .A1(n15228), .A2(n15227), .ZN(n15239) );
  OR2_X1 U17004 ( .A1(n15228), .A2(n15227), .ZN(n15229) );
  NAND2_X1 U17005 ( .A1(n15239), .A2(n15229), .ZN(n15230) );
  INV_X1 U17006 ( .A(n15230), .ZN(n15231) );
  OR2_X1 U17007 ( .A1(n15230), .A2(n9747), .ZN(n15240) );
  OAI211_X1 U17008 ( .C1(n15231), .C2(P1_REG2_REG_18__SCAN_IN), .A(n15244), 
        .B(n15240), .ZN(n15232) );
  NAND3_X1 U17009 ( .A1(n15234), .A2(n15233), .A3(n15232), .ZN(P1_U3261) );
  NAND2_X1 U17010 ( .A1(n15236), .A2(n15235), .ZN(n15238) );
  XNOR2_X1 U17011 ( .A(n15238), .B(n15237), .ZN(n15249) );
  INV_X1 U17012 ( .A(n15249), .ZN(n15243) );
  NAND2_X1 U17013 ( .A1(n15240), .A2(n15239), .ZN(n15241) );
  XNOR2_X1 U17014 ( .A(n15241), .B(P1_REG2_REG_19__SCAN_IN), .ZN(n15245) );
  NAND2_X1 U17015 ( .A1(n15245), .A2(n15244), .ZN(n15247) );
  INV_X1 U17016 ( .A(n15265), .ZN(n15544) );
  NAND2_X1 U17017 ( .A1(n15544), .A2(n15260), .ZN(n15253) );
  NOR2_X1 U17018 ( .A1(n15528), .A2(n15254), .ZN(n15257) );
  NAND2_X1 U17019 ( .A1(n15256), .A2(n15255), .ZN(n15542) );
  NOR2_X1 U17020 ( .A1(n6556), .A2(n15542), .ZN(n15263) );
  AOI211_X1 U17021 ( .C1(n15258), .C2(n15496), .A(n15257), .B(n15263), .ZN(
        n15259) );
  OAI21_X1 U17022 ( .B1(n15540), .B2(n15344), .A(n15259), .ZN(P1_U3263) );
  XNOR2_X1 U17023 ( .A(n15260), .B(n15265), .ZN(n15261) );
  NAND2_X1 U17024 ( .A1(n15261), .A2(n7132), .ZN(n15543) );
  NOR2_X1 U17025 ( .A1(n15528), .A2(n15262), .ZN(n15264) );
  AOI211_X1 U17026 ( .C1(n15265), .C2(n15496), .A(n15264), .B(n15263), .ZN(
        n15266) );
  OAI21_X1 U17027 ( .B1(n15543), .B2(n15344), .A(n15266), .ZN(P1_U3264) );
  XNOR2_X1 U17028 ( .A(n15268), .B(n15269), .ZN(n15556) );
  NAND2_X1 U17029 ( .A1(n15272), .A2(n15500), .ZN(n15274) );
  INV_X1 U17030 ( .A(n15555), .ZN(n15286) );
  NAND2_X1 U17031 ( .A1(n15553), .A2(n15277), .ZN(n15278) );
  NAND2_X1 U17032 ( .A1(n15278), .A2(n7132), .ZN(n15279) );
  NOR2_X1 U17033 ( .A1(n15280), .A2(n15279), .ZN(n15552) );
  NAND2_X1 U17034 ( .A1(n15552), .A2(n15812), .ZN(n15283) );
  AOI22_X1 U17035 ( .A1(n15281), .A2(n15525), .B1(P1_REG2_REG_28__SCAN_IN), 
        .B2(n6556), .ZN(n15282) );
  OAI211_X1 U17036 ( .C1(n15284), .C2(n15807), .A(n15283), .B(n15282), .ZN(
        n15285) );
  AOI21_X1 U17037 ( .B1(n15286), .B2(n15528), .A(n15285), .ZN(n15287) );
  OAI21_X1 U17038 ( .B1(n15556), .B2(n15535), .A(n15287), .ZN(P1_U3265) );
  XNOR2_X1 U17039 ( .A(n15288), .B(n15293), .ZN(n15569) );
  INV_X1 U17040 ( .A(n15289), .ZN(n15291) );
  OAI21_X1 U17041 ( .B1(n15352), .B2(n15291), .A(n15290), .ZN(n15294) );
  NAND3_X1 U17042 ( .A1(n15294), .A2(n15293), .A3(n15292), .ZN(n15296) );
  NAND2_X1 U17043 ( .A1(n15296), .A2(n15295), .ZN(n15567) );
  OAI211_X1 U17044 ( .C1(n15312), .C2(n15565), .A(n7132), .B(n6625), .ZN(
        n15564) );
  AOI22_X1 U17045 ( .A1(n15297), .A2(n15500), .B1(n15521), .B2(n15330), .ZN(
        n15563) );
  AOI22_X1 U17046 ( .A1(n15298), .A2(n15525), .B1(P1_REG2_REG_26__SCAN_IN), 
        .B2(n6556), .ZN(n15299) );
  OAI21_X1 U17047 ( .B1(n15563), .B2(n6556), .A(n15299), .ZN(n15300) );
  AOI21_X1 U17048 ( .B1(n15301), .B2(n15496), .A(n15300), .ZN(n15302) );
  OAI21_X1 U17049 ( .B1(n15564), .B2(n15344), .A(n15302), .ZN(n15303) );
  AOI21_X1 U17050 ( .B1(n15567), .B2(n15428), .A(n15303), .ZN(n15304) );
  OAI21_X1 U17051 ( .B1(n15569), .B2(n15535), .A(n15304), .ZN(P1_U3267) );
  NAND2_X1 U17052 ( .A1(n15350), .A2(n15305), .ZN(n15322) );
  INV_X1 U17053 ( .A(n15308), .ZN(n15309) );
  AOI21_X1 U17054 ( .B1(n15311), .B2(n15310), .A(n15309), .ZN(n15574) );
  INV_X1 U17055 ( .A(n15312), .ZN(n15313) );
  OAI211_X1 U17056 ( .C1(n15572), .C2(n15338), .A(n15313), .B(n7132), .ZN(
        n15571) );
  INV_X1 U17057 ( .A(n15314), .ZN(n15315) );
  AOI22_X1 U17058 ( .A1(n15315), .A2(n15525), .B1(P1_REG2_REG_25__SCAN_IN), 
        .B2(n6556), .ZN(n15316) );
  OAI21_X1 U17059 ( .B1(n15570), .B2(n6556), .A(n15316), .ZN(n15317) );
  AOI21_X1 U17060 ( .B1(n15318), .B2(n15496), .A(n15317), .ZN(n15319) );
  OAI21_X1 U17061 ( .B1(n15571), .B2(n15344), .A(n15319), .ZN(n15320) );
  AOI21_X1 U17062 ( .B1(n15574), .B2(n15513), .A(n15320), .ZN(n15321) );
  OAI21_X1 U17063 ( .B1(n15576), .B2(n15480), .A(n15321), .ZN(P1_U3268) );
  NAND2_X1 U17064 ( .A1(n15322), .A2(n13019), .ZN(n15323) );
  NAND2_X1 U17065 ( .A1(n15323), .A2(n15611), .ZN(n15324) );
  OR2_X1 U17066 ( .A1(n15325), .A2(n15324), .ZN(n15335) );
  NAND2_X1 U17067 ( .A1(n15327), .A2(n15326), .ZN(n15328) );
  NAND2_X1 U17068 ( .A1(n15329), .A2(n15328), .ZN(n15580) );
  NAND2_X1 U17069 ( .A1(n15330), .A2(n15500), .ZN(n15331) );
  OAI21_X1 U17070 ( .B1(n15332), .B2(n15431), .A(n15331), .ZN(n15333) );
  AOI21_X1 U17071 ( .B1(n15580), .B2(n15850), .A(n15333), .ZN(n15334) );
  NAND2_X1 U17072 ( .A1(n15336), .A2(n15341), .ZN(n15337) );
  NAND2_X1 U17073 ( .A1(n15337), .A2(n7132), .ZN(n15339) );
  OR2_X1 U17074 ( .A1(n15339), .A2(n15338), .ZN(n15577) );
  AOI22_X1 U17075 ( .A1(n15340), .A2(n15525), .B1(P1_REG2_REG_24__SCAN_IN), 
        .B2(n6556), .ZN(n15343) );
  NAND2_X1 U17076 ( .A1(n15341), .A2(n15496), .ZN(n15342) );
  OAI211_X1 U17077 ( .C1(n15577), .C2(n15344), .A(n15343), .B(n15342), .ZN(
        n15345) );
  AOI21_X1 U17078 ( .B1(n15580), .B2(n15813), .A(n15345), .ZN(n15346) );
  OAI21_X1 U17079 ( .B1(n15582), .B2(n6556), .A(n15346), .ZN(P1_U3269) );
  OAI21_X1 U17080 ( .B1(n7984), .B2(n15348), .A(n15347), .ZN(n15589) );
  INV_X1 U17081 ( .A(n15349), .ZN(n15354) );
  OAI21_X1 U17082 ( .B1(n15352), .B2(n15351), .A(n15350), .ZN(n15353) );
  NAND2_X1 U17083 ( .A1(n15353), .A2(n15611), .ZN(n15588) );
  OAI211_X1 U17084 ( .C1(n15804), .C2(n15354), .A(n15588), .B(n15583), .ZN(
        n15355) );
  NAND2_X1 U17085 ( .A1(n15355), .A2(n15528), .ZN(n15359) );
  AOI211_X1 U17086 ( .C1(n15586), .C2(n15365), .A(n15608), .B(n13058), .ZN(
        n15584) );
  OAI22_X1 U17087 ( .A1(n15356), .A2(n15807), .B1(n11015), .B2(n15528), .ZN(
        n15357) );
  AOI21_X1 U17088 ( .B1(n15584), .B2(n15812), .A(n15357), .ZN(n15358) );
  OAI211_X1 U17089 ( .C1(n15589), .C2(n15535), .A(n15359), .B(n15358), .ZN(
        P1_U3270) );
  XNOR2_X1 U17090 ( .A(n15360), .B(n15361), .ZN(n15364) );
  AOI222_X1 U17091 ( .A1(n15611), .A2(n15364), .B1(n15363), .B2(n15521), .C1(
        n15362), .C2(n15500), .ZN(n15593) );
  INV_X1 U17092 ( .A(n15392), .ZN(n15367) );
  INV_X1 U17093 ( .A(n15365), .ZN(n15366) );
  AOI211_X1 U17094 ( .C1(n15591), .C2(n15367), .A(n15608), .B(n15366), .ZN(
        n15590) );
  AOI22_X1 U17095 ( .A1(n15368), .A2(n15525), .B1(P1_REG2_REG_22__SCAN_IN), 
        .B2(n6556), .ZN(n15369) );
  OAI21_X1 U17096 ( .B1(n15370), .B2(n15807), .A(n15369), .ZN(n15380) );
  INV_X1 U17097 ( .A(n15383), .ZN(n15372) );
  NOR2_X1 U17098 ( .A1(n15372), .A2(n15371), .ZN(n15376) );
  OAI211_X1 U17099 ( .C1(n15376), .C2(n15375), .A(n15374), .B(n15373), .ZN(
        n15377) );
  AND2_X1 U17100 ( .A1(n15378), .A2(n15377), .ZN(n15594) );
  NOR2_X1 U17101 ( .A1(n15594), .A2(n15535), .ZN(n15379) );
  AOI211_X1 U17102 ( .C1(n15590), .C2(n15812), .A(n15380), .B(n15379), .ZN(
        n15381) );
  OAI21_X1 U17103 ( .B1(n15593), .B2(n6556), .A(n15381), .ZN(P1_U3271) );
  NAND2_X1 U17104 ( .A1(n15383), .A2(n15382), .ZN(n15400) );
  NAND2_X1 U17105 ( .A1(n15402), .A2(n15384), .ZN(n15386) );
  XNOR2_X1 U17106 ( .A(n15386), .B(n15385), .ZN(n15599) );
  XNOR2_X1 U17107 ( .A(n15388), .B(n15387), .ZN(n15389) );
  OAI222_X1 U17108 ( .A1(n15516), .A2(n15391), .B1(n15431), .B2(n15390), .C1(
        n15389), .C2(n15826), .ZN(n15595) );
  NAND2_X1 U17109 ( .A1(n15595), .A2(n15528), .ZN(n15399) );
  AOI211_X1 U17110 ( .C1(n15597), .C2(n15408), .A(n15608), .B(n15392), .ZN(
        n15596) );
  NOR2_X1 U17111 ( .A1(n15393), .A2(n15807), .ZN(n15397) );
  OAI22_X1 U17112 ( .A1(n15395), .A2(n15528), .B1(n15394), .B2(n15804), .ZN(
        n15396) );
  AOI211_X1 U17113 ( .C1(n15596), .C2(n15812), .A(n15397), .B(n15396), .ZN(
        n15398) );
  OAI211_X1 U17114 ( .C1(n15599), .C2(n15535), .A(n15399), .B(n15398), .ZN(
        P1_U3272) );
  NAND2_X1 U17115 ( .A1(n15400), .A2(n15404), .ZN(n15401) );
  NAND2_X1 U17116 ( .A1(n15402), .A2(n15401), .ZN(n15604) );
  OAI211_X1 U17117 ( .C1(n15405), .C2(n15404), .A(n15403), .B(n15611), .ZN(
        n15407) );
  NAND2_X1 U17118 ( .A1(n15407), .A2(n15406), .ZN(n15600) );
  NAND2_X1 U17119 ( .A1(n15600), .A2(n15528), .ZN(n15414) );
  INV_X1 U17120 ( .A(n15408), .ZN(n15409) );
  AOI211_X1 U17121 ( .C1(n15602), .C2(n15418), .A(n15608), .B(n15409), .ZN(
        n15601) );
  AOI22_X1 U17122 ( .A1(n15410), .A2(n15525), .B1(n6556), .B2(
        P1_REG2_REG_20__SCAN_IN), .ZN(n15411) );
  OAI21_X1 U17123 ( .B1(n7457), .B2(n15807), .A(n15411), .ZN(n15412) );
  AOI21_X1 U17124 ( .B1(n15601), .B2(n15812), .A(n15412), .ZN(n15413) );
  OAI211_X1 U17125 ( .C1(n15604), .C2(n15535), .A(n15414), .B(n15413), .ZN(
        P1_U3273) );
  XNOR2_X1 U17126 ( .A(n15415), .B(n15416), .ZN(n15614) );
  XNOR2_X1 U17127 ( .A(n15417), .B(n15416), .ZN(n15612) );
  OAI21_X1 U17128 ( .B1(n6612), .B2(n7456), .A(n15418), .ZN(n15609) );
  AND2_X1 U17129 ( .A1(n15419), .A2(n15521), .ZN(n15420) );
  AOI21_X1 U17130 ( .B1(n15421), .B2(n15500), .A(n15420), .ZN(n15607) );
  OAI22_X1 U17131 ( .A1(n15607), .A2(n6556), .B1(n15422), .B2(n15804), .ZN(
        n15424) );
  NOR2_X1 U17132 ( .A1(n7456), .A2(n15807), .ZN(n15423) );
  AOI211_X1 U17133 ( .C1(n6556), .C2(P1_REG2_REG_19__SCAN_IN), .A(n15424), .B(
        n15423), .ZN(n15425) );
  OAI21_X1 U17134 ( .B1(n15426), .B2(n15609), .A(n15425), .ZN(n15427) );
  AOI21_X1 U17135 ( .B1(n15612), .B2(n15428), .A(n15427), .ZN(n15429) );
  OAI21_X1 U17136 ( .B1(n15614), .B2(n15535), .A(n15429), .ZN(P1_U3274) );
  XOR2_X1 U17137 ( .A(n15430), .B(n15434), .Z(n15439) );
  OAI22_X1 U17138 ( .A1(n15433), .A2(n15516), .B1(n15432), .B2(n15431), .ZN(
        n15438) );
  XNOR2_X1 U17139 ( .A(n15435), .B(n15434), .ZN(n15619) );
  NOR2_X1 U17140 ( .A1(n15619), .A2(n15436), .ZN(n15437) );
  AOI211_X1 U17141 ( .C1(n15439), .C2(n15611), .A(n15438), .B(n15437), .ZN(
        n15618) );
  INV_X1 U17142 ( .A(n15440), .ZN(n15441) );
  AOI211_X1 U17143 ( .C1(n15616), .C2(n15441), .A(n15608), .B(n6612), .ZN(
        n15615) );
  AOI22_X1 U17144 ( .A1(n6556), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n15442), 
        .B2(n15525), .ZN(n15443) );
  OAI21_X1 U17145 ( .B1(n15444), .B2(n15807), .A(n15443), .ZN(n15447) );
  NOR2_X1 U17146 ( .A1(n15619), .A2(n15445), .ZN(n15446) );
  AOI211_X1 U17147 ( .C1(n15615), .C2(n15812), .A(n15447), .B(n15446), .ZN(
        n15448) );
  OAI21_X1 U17148 ( .B1(n15618), .B2(n6556), .A(n15448), .ZN(P1_U3275) );
  XOR2_X1 U17149 ( .A(n15449), .B(n15450), .Z(n15625) );
  AOI21_X1 U17150 ( .B1(n15451), .B2(n15450), .A(n15826), .ZN(n15455) );
  INV_X1 U17151 ( .A(n15452), .ZN(n15453) );
  AOI21_X1 U17152 ( .B1(n15455), .B2(n15454), .A(n15453), .ZN(n15624) );
  NAND2_X1 U17153 ( .A1(n6556), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n15456) );
  OAI21_X1 U17154 ( .B1(n15804), .B2(n15457), .A(n15456), .ZN(n15458) );
  AOI21_X1 U17155 ( .B1(n15622), .B2(n15496), .A(n15458), .ZN(n15462) );
  OAI21_X1 U17156 ( .B1(n15471), .B2(n15459), .A(n7132), .ZN(n15460) );
  NOR2_X1 U17157 ( .A1(n15460), .A2(n15440), .ZN(n15621) );
  NAND2_X1 U17158 ( .A1(n15621), .A2(n15812), .ZN(n15461) );
  OAI211_X1 U17159 ( .C1(n15624), .C2(n6556), .A(n15462), .B(n15461), .ZN(
        n15463) );
  INV_X1 U17160 ( .A(n15463), .ZN(n15464) );
  OAI21_X1 U17161 ( .B1(n15535), .B2(n15625), .A(n15464), .ZN(P1_U3276) );
  XOR2_X1 U17162 ( .A(n15465), .B(n15467), .Z(n15632) );
  OAI21_X1 U17163 ( .B1(n15468), .B2(n15467), .A(n15466), .ZN(n15629) );
  NAND2_X1 U17164 ( .A1(n15490), .A2(n15628), .ZN(n15469) );
  NAND2_X1 U17165 ( .A1(n15469), .A2(n7132), .ZN(n15470) );
  NOR2_X1 U17166 ( .A1(n15471), .A2(n15470), .ZN(n15626) );
  NAND2_X1 U17167 ( .A1(n15626), .A2(n15812), .ZN(n15476) );
  INV_X1 U17168 ( .A(n15627), .ZN(n15473) );
  OAI22_X1 U17169 ( .A1(n15473), .A2(n6556), .B1(n15472), .B2(n15804), .ZN(
        n15474) );
  AOI21_X1 U17170 ( .B1(P1_REG2_REG_16__SCAN_IN), .B2(n6556), .A(n15474), .ZN(
        n15475) );
  OAI211_X1 U17171 ( .C1(n15477), .C2(n15807), .A(n15476), .B(n15475), .ZN(
        n15478) );
  AOI21_X1 U17172 ( .B1(n15629), .B2(n15513), .A(n15478), .ZN(n15479) );
  OAI21_X1 U17173 ( .B1(n15632), .B2(n15480), .A(n15479), .ZN(P1_U3277) );
  INV_X1 U17174 ( .A(n15481), .ZN(n15506) );
  NAND2_X1 U17175 ( .A1(n15506), .A2(n15505), .ZN(n15504) );
  NAND2_X1 U17176 ( .A1(n15504), .A2(n15482), .ZN(n15483) );
  XNOR2_X1 U17177 ( .A(n15483), .B(n15485), .ZN(n15637) );
  XNOR2_X1 U17178 ( .A(n15486), .B(n15485), .ZN(n15488) );
  AOI21_X1 U17179 ( .B1(n15488), .B2(n15611), .A(n15487), .ZN(n15636) );
  INV_X1 U17180 ( .A(n15636), .ZN(n15495) );
  INV_X1 U17181 ( .A(n15490), .ZN(n15491) );
  AOI21_X1 U17182 ( .B1(n15633), .B2(n15489), .A(n15491), .ZN(n15634) );
  INV_X1 U17183 ( .A(n15634), .ZN(n15493) );
  OAI22_X1 U17184 ( .A1(n15493), .A2(n11835), .B1(n15492), .B2(n15804), .ZN(
        n15494) );
  OAI21_X1 U17185 ( .B1(n15495), .B2(n15494), .A(n15528), .ZN(n15498) );
  AOI22_X1 U17186 ( .A1(n15633), .A2(n15496), .B1(P1_REG2_REG_15__SCAN_IN), 
        .B2(n6556), .ZN(n15497) );
  OAI211_X1 U17187 ( .C1(n15637), .C2(n15535), .A(n15498), .B(n15497), .ZN(
        P1_U3278) );
  XNOR2_X1 U17188 ( .A(n15499), .B(n15505), .ZN(n15503) );
  AOI222_X1 U17189 ( .A1(n15611), .A2(n15503), .B1(n15502), .B2(n15521), .C1(
        n15501), .C2(n15500), .ZN(n15641) );
  OAI21_X1 U17190 ( .B1(n15506), .B2(n15505), .A(n15504), .ZN(n15642) );
  INV_X1 U17191 ( .A(n15642), .ZN(n15514) );
  OR2_X1 U17192 ( .A1(n15511), .A2(n15527), .ZN(n15507) );
  AND3_X1 U17193 ( .A1(n15489), .A2(n15507), .A3(n7132), .ZN(n15638) );
  NAND2_X1 U17194 ( .A1(n15638), .A2(n15812), .ZN(n15510) );
  AOI22_X1 U17195 ( .A1(n6556), .A2(P1_REG2_REG_14__SCAN_IN), .B1(n15508), 
        .B2(n15525), .ZN(n15509) );
  OAI211_X1 U17196 ( .C1(n15511), .C2(n15807), .A(n15510), .B(n15509), .ZN(
        n15512) );
  AOI21_X1 U17197 ( .B1(n15514), .B2(n15513), .A(n15512), .ZN(n15515) );
  OAI21_X1 U17198 ( .B1(n15641), .B2(n6556), .A(n15515), .ZN(P1_U3279) );
  NOR2_X1 U17199 ( .A1(n15517), .A2(n15516), .ZN(n15644) );
  XNOR2_X1 U17200 ( .A(n15519), .B(n15532), .ZN(n15522) );
  AOI22_X1 U17201 ( .A1(n15522), .A2(n15611), .B1(n15521), .B2(n15520), .ZN(
        n15646) );
  INV_X1 U17202 ( .A(n15646), .ZN(n15523) );
  AOI211_X1 U17203 ( .C1(n15525), .C2(n15524), .A(n15644), .B(n15523), .ZN(
        n15539) );
  AOI211_X1 U17204 ( .C1(n15645), .C2(n12568), .A(n15608), .B(n15527), .ZN(
        n15643) );
  OAI22_X1 U17205 ( .A1(n15530), .A2(n15807), .B1(n15529), .B2(n15528), .ZN(
        n15537) );
  OAI21_X1 U17206 ( .B1(n15533), .B2(n15532), .A(n15531), .ZN(n15534) );
  INV_X1 U17207 ( .A(n15534), .ZN(n15648) );
  NOR2_X1 U17208 ( .A1(n15648), .A2(n15535), .ZN(n15536) );
  AOI211_X1 U17209 ( .C1(n15643), .C2(n15812), .A(n15537), .B(n15536), .ZN(
        n15538) );
  OAI21_X1 U17210 ( .B1(n15539), .B2(n6556), .A(n15538), .ZN(P1_U3280) );
  OAI211_X1 U17211 ( .C1(n15844), .C2(n15544), .A(n15543), .B(n15542), .ZN(
        n15667) );
  MUX2_X1 U17212 ( .A(n15667), .B(P1_REG1_REG_30__SCAN_IN), .S(n15884), .Z(
        P1_U3558) );
  OAI21_X1 U17213 ( .B1(n15547), .B2(n15844), .A(n15546), .ZN(n15548) );
  AOI21_X1 U17214 ( .B1(n15870), .B2(n15553), .A(n15552), .ZN(n15554) );
  INV_X1 U17215 ( .A(n15557), .ZN(n15562) );
  AOI21_X1 U17216 ( .B1(n15870), .B2(n7122), .A(n15558), .ZN(n15560) );
  OAI211_X1 U17217 ( .C1(n15844), .C2(n15565), .A(n15564), .B(n15563), .ZN(
        n15566) );
  AOI21_X1 U17218 ( .B1(n15567), .B2(n15611), .A(n15566), .ZN(n15568) );
  OAI21_X1 U17219 ( .B1(n15874), .B2(n15569), .A(n15568), .ZN(n15671) );
  MUX2_X1 U17220 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n15671), .S(n15886), .Z(
        P1_U3554) );
  INV_X1 U17221 ( .A(n15874), .ZN(n15865) );
  OAI211_X1 U17222 ( .C1(n15844), .C2(n15572), .A(n15571), .B(n15570), .ZN(
        n15573) );
  AOI21_X1 U17223 ( .B1(n15574), .B2(n15865), .A(n15573), .ZN(n15575) );
  OAI21_X1 U17224 ( .B1(n15576), .B2(n15826), .A(n15575), .ZN(n15672) );
  MUX2_X1 U17225 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n15672), .S(n15886), .Z(
        P1_U3553) );
  INV_X1 U17226 ( .A(n15620), .ZN(n15851) );
  OAI21_X1 U17227 ( .B1(n15844), .B2(n15578), .A(n15577), .ZN(n15579) );
  AOI21_X1 U17228 ( .B1(n15580), .B2(n15851), .A(n15579), .ZN(n15581) );
  NAND2_X1 U17229 ( .A1(n15582), .A2(n15581), .ZN(n15673) );
  MUX2_X1 U17230 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n15673), .S(n15886), .Z(
        P1_U3552) );
  INV_X1 U17231 ( .A(n15583), .ZN(n15585) );
  AOI211_X1 U17232 ( .C1(n15870), .C2(n15586), .A(n15585), .B(n15584), .ZN(
        n15587) );
  OAI211_X1 U17233 ( .C1(n15874), .C2(n15589), .A(n15588), .B(n15587), .ZN(
        n15674) );
  MUX2_X1 U17234 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n15674), .S(n15886), .Z(
        P1_U3551) );
  AOI21_X1 U17235 ( .B1(n15591), .B2(n15870), .A(n15590), .ZN(n15592) );
  OAI211_X1 U17236 ( .C1(n15874), .C2(n15594), .A(n15593), .B(n15592), .ZN(
        n15675) );
  MUX2_X1 U17237 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n15675), .S(n15886), .Z(
        P1_U3550) );
  AOI211_X1 U17238 ( .C1(n15870), .C2(n15597), .A(n15596), .B(n15595), .ZN(
        n15598) );
  OAI21_X1 U17239 ( .B1(n15874), .B2(n15599), .A(n15598), .ZN(n15676) );
  MUX2_X1 U17240 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n15676), .S(n15886), .Z(
        P1_U3549) );
  AOI211_X1 U17241 ( .C1(n15870), .C2(n15602), .A(n15601), .B(n15600), .ZN(
        n15603) );
  OAI21_X1 U17242 ( .B1(n15874), .B2(n15604), .A(n15603), .ZN(n15677) );
  MUX2_X1 U17243 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n15677), .S(n15886), .Z(
        P1_U3548) );
  NAND2_X1 U17244 ( .A1(n15605), .A2(n15870), .ZN(n15606) );
  OAI211_X1 U17245 ( .C1(n15609), .C2(n15608), .A(n15607), .B(n15606), .ZN(
        n15610) );
  AOI21_X1 U17246 ( .B1(n15612), .B2(n15611), .A(n15610), .ZN(n15613) );
  OAI21_X1 U17247 ( .B1(n15874), .B2(n15614), .A(n15613), .ZN(n15678) );
  MUX2_X1 U17248 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n15678), .S(n15886), .Z(
        P1_U3547) );
  AOI21_X1 U17249 ( .B1(n15870), .B2(n15616), .A(n15615), .ZN(n15617) );
  OAI211_X1 U17250 ( .C1(n15620), .C2(n15619), .A(n15618), .B(n15617), .ZN(
        n15679) );
  MUX2_X1 U17251 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n15679), .S(n15886), .Z(
        P1_U3546) );
  AOI21_X1 U17252 ( .B1(n15870), .B2(n15622), .A(n15621), .ZN(n15623) );
  OAI211_X1 U17253 ( .C1(n15625), .C2(n15874), .A(n15624), .B(n15623), .ZN(
        n15680) );
  MUX2_X1 U17254 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n15680), .S(n15886), .Z(
        P1_U3545) );
  AOI211_X1 U17255 ( .C1(n15870), .C2(n15628), .A(n15627), .B(n15626), .ZN(
        n15631) );
  NAND2_X1 U17256 ( .A1(n15629), .A2(n15865), .ZN(n15630) );
  OAI211_X1 U17257 ( .C1(n15632), .C2(n15826), .A(n15631), .B(n15630), .ZN(
        n15681) );
  MUX2_X1 U17258 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n15681), .S(n15886), .Z(
        P1_U3544) );
  AOI22_X1 U17259 ( .A1(n15634), .A2(n7132), .B1(n15870), .B2(n15633), .ZN(
        n15635) );
  OAI211_X1 U17260 ( .C1(n15637), .C2(n15874), .A(n15636), .B(n15635), .ZN(
        n15682) );
  MUX2_X1 U17261 ( .A(P1_REG1_REG_15__SCAN_IN), .B(n15682), .S(n15886), .Z(
        P1_U3543) );
  AOI21_X1 U17262 ( .B1(n15870), .B2(n15639), .A(n15638), .ZN(n15640) );
  OAI211_X1 U17263 ( .C1(n15874), .C2(n15642), .A(n15641), .B(n15640), .ZN(
        n15683) );
  MUX2_X1 U17264 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n15683), .S(n15886), .Z(
        P1_U3542) );
  AOI211_X1 U17265 ( .C1(n15870), .C2(n15645), .A(n15644), .B(n15643), .ZN(
        n15647) );
  OAI211_X1 U17266 ( .C1(n15874), .C2(n15648), .A(n15647), .B(n15646), .ZN(
        n15684) );
  MUX2_X1 U17267 ( .A(P1_REG1_REG_13__SCAN_IN), .B(n15684), .S(n15886), .Z(
        P1_U3541) );
  AOI211_X1 U17268 ( .C1(n15870), .C2(n15651), .A(n15650), .B(n15649), .ZN(
        n15654) );
  NAND2_X1 U17269 ( .A1(n15652), .A2(n15865), .ZN(n15653) );
  OAI211_X1 U17270 ( .C1(n15826), .C2(n15655), .A(n15654), .B(n15653), .ZN(
        n15685) );
  MUX2_X1 U17271 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n15685), .S(n15886), .Z(
        P1_U3540) );
  NAND2_X1 U17272 ( .A1(n15656), .A2(n15865), .ZN(n15658) );
  NAND4_X1 U17273 ( .A1(n15660), .A2(n15659), .A3(n15658), .A4(n15657), .ZN(
        n15686) );
  MUX2_X1 U17274 ( .A(P1_REG1_REG_11__SCAN_IN), .B(n15686), .S(n15886), .Z(
        P1_U3539) );
  AOI21_X1 U17275 ( .B1(n15870), .B2(n15662), .A(n15661), .ZN(n15663) );
  OAI211_X1 U17276 ( .C1(n15874), .C2(n15665), .A(n15664), .B(n15663), .ZN(
        n15687) );
  MUX2_X1 U17277 ( .A(P1_REG1_REG_9__SCAN_IN), .B(n15687), .S(n15886), .Z(
        P1_U3537) );
  MUX2_X1 U17278 ( .A(n15667), .B(P1_REG0_REG_30__SCAN_IN), .S(n15876), .Z(
        P1_U3526) );
  MUX2_X1 U17279 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n15669), .S(n15877), .Z(
        P1_U3524) );
  MUX2_X1 U17280 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n15671), .S(n15877), .Z(
        P1_U3522) );
  MUX2_X1 U17281 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n15672), .S(n15877), .Z(
        P1_U3521) );
  MUX2_X1 U17282 ( .A(n15673), .B(P1_REG0_REG_24__SCAN_IN), .S(n15876), .Z(
        P1_U3520) );
  MUX2_X1 U17283 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n15674), .S(n15877), .Z(
        P1_U3519) );
  MUX2_X1 U17284 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n15675), .S(n15877), .Z(
        P1_U3518) );
  MUX2_X1 U17285 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n15676), .S(n15877), .Z(
        P1_U3517) );
  MUX2_X1 U17286 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n15677), .S(n15877), .Z(
        P1_U3516) );
  MUX2_X1 U17287 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n15678), .S(n15877), .Z(
        P1_U3515) );
  MUX2_X1 U17288 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n15679), .S(n15877), .Z(
        P1_U3513) );
  MUX2_X1 U17289 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n15680), .S(n15877), .Z(
        P1_U3510) );
  MUX2_X1 U17290 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n15681), .S(n15877), .Z(
        P1_U3507) );
  MUX2_X1 U17291 ( .A(P1_REG0_REG_15__SCAN_IN), .B(n15682), .S(n15877), .Z(
        P1_U3504) );
  MUX2_X1 U17292 ( .A(P1_REG0_REG_14__SCAN_IN), .B(n15683), .S(n15877), .Z(
        P1_U3501) );
  MUX2_X1 U17293 ( .A(P1_REG0_REG_13__SCAN_IN), .B(n15684), .S(n15877), .Z(
        P1_U3498) );
  MUX2_X1 U17294 ( .A(P1_REG0_REG_12__SCAN_IN), .B(n15685), .S(n15877), .Z(
        P1_U3495) );
  MUX2_X1 U17295 ( .A(P1_REG0_REG_11__SCAN_IN), .B(n15686), .S(n15877), .Z(
        P1_U3492) );
  MUX2_X1 U17296 ( .A(P1_REG0_REG_9__SCAN_IN), .B(n15687), .S(n15877), .Z(
        P1_U3486) );
  NOR4_X1 U17297 ( .A1(n15689), .A2(P1_IR_REG_30__SCAN_IN), .A3(P1_U3086), 
        .A4(n9447), .ZN(n15690) );
  AOI21_X1 U17298 ( .B1(n15691), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n15690), 
        .ZN(n15692) );
  OAI21_X1 U17299 ( .B1(n15693), .B2(n15703), .A(n15692), .ZN(P1_U3324) );
  OAI222_X1 U17300 ( .A1(n15699), .A2(P1_U3086), .B1(n15703), .B2(n15698), 
        .C1(n15697), .C2(n15700), .ZN(P1_U3328) );
  OAI222_X1 U17301 ( .A1(n15704), .A2(P1_U3086), .B1(n15703), .B2(n15702), 
        .C1(n15701), .C2(n15700), .ZN(P1_U3329) );
  MUX2_X1 U17302 ( .A(n15706), .B(n15705), .S(P1_STATE_REG_SCAN_IN), .Z(
        P1_U3333) );
  MUX2_X1 U17303 ( .A(n15707), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  XOR2_X1 U17304 ( .A(P2_ADDR_REG_0__SCAN_IN), .B(n15708), .Z(SUB_1596_U53) );
  INV_X1 U17305 ( .A(n15710), .ZN(n15712) );
  NAND2_X1 U17306 ( .A1(n15714), .A2(n15713), .ZN(n15716) );
  NAND2_X1 U17307 ( .A1(n15716), .A2(n15715), .ZN(n15727) );
  XNOR2_X1 U17308 ( .A(n15725), .B(P3_ADDR_REG_14__SCAN_IN), .ZN(n15726) );
  INV_X1 U17309 ( .A(n15726), .ZN(n15717) );
  XNOR2_X1 U17310 ( .A(n15727), .B(n15717), .ZN(n15721) );
  XNOR2_X1 U17311 ( .A(n15721), .B(P2_ADDR_REG_14__SCAN_IN), .ZN(n15718) );
  XNOR2_X1 U17312 ( .A(n15720), .B(n15718), .ZN(SUB_1596_U66) );
  INV_X1 U17313 ( .A(n15721), .ZN(n15723) );
  INV_X1 U17314 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n15722) );
  OAI22_X1 U17315 ( .A1(n15727), .A2(n15726), .B1(P3_ADDR_REG_14__SCAN_IN), 
        .B2(n15725), .ZN(n15731) );
  XNOR2_X1 U17316 ( .A(P3_ADDR_REG_15__SCAN_IN), .B(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n15728) );
  XNOR2_X1 U17317 ( .A(n15731), .B(n15728), .ZN(n15739) );
  XOR2_X1 U17318 ( .A(P2_ADDR_REG_15__SCAN_IN), .B(n15739), .Z(n15729) );
  XNOR2_X1 U17319 ( .A(n15736), .B(n15729), .ZN(SUB_1596_U65) );
  NOR2_X1 U17320 ( .A1(P3_ADDR_REG_15__SCAN_IN), .A2(n15732), .ZN(n15730) );
  OR2_X1 U17321 ( .A1(n15731), .A2(n15730), .ZN(n15734) );
  NAND2_X1 U17322 ( .A1(n15732), .A2(P3_ADDR_REG_15__SCAN_IN), .ZN(n15733) );
  NAND2_X1 U17323 ( .A1(n15734), .A2(n15733), .ZN(n15744) );
  XNOR2_X1 U17324 ( .A(n15744), .B(P1_ADDR_REG_16__SCAN_IN), .ZN(n15746) );
  XNOR2_X1 U17325 ( .A(n15746), .B(n15735), .ZN(n15738) );
  OAI211_X1 U17326 ( .C1(n15740), .C2(n15739), .A(n15738), .B(n15737), .ZN(
        n15742) );
  NAND2_X1 U17327 ( .A1(n6850), .A2(n15742), .ZN(n15741) );
  XNOR2_X1 U17328 ( .A(n15741), .B(P2_ADDR_REG_16__SCAN_IN), .ZN(SUB_1596_U64)
         );
  NAND2_X1 U17329 ( .A1(n15745), .A2(n15744), .ZN(n15748) );
  NAND2_X1 U17330 ( .A1(P3_ADDR_REG_16__SCAN_IN), .A2(n15746), .ZN(n15747) );
  NAND2_X1 U17331 ( .A1(n15748), .A2(n15747), .ZN(n15755) );
  XNOR2_X1 U17332 ( .A(n15755), .B(P1_ADDR_REG_17__SCAN_IN), .ZN(n15754) );
  XNOR2_X1 U17333 ( .A(n15754), .B(P3_ADDR_REG_17__SCAN_IN), .ZN(n15749) );
  INV_X1 U17334 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n15752) );
  XNOR2_X1 U17335 ( .A(n15753), .B(n15752), .ZN(SUB_1596_U63) );
  INV_X1 U17336 ( .A(n15749), .ZN(n15750) );
  NAND2_X1 U17337 ( .A1(n15754), .A2(P3_ADDR_REG_17__SCAN_IN), .ZN(n15758) );
  NAND2_X1 U17338 ( .A1(n15756), .A2(n15755), .ZN(n15757) );
  NAND2_X1 U17339 ( .A1(n15758), .A2(n15757), .ZN(n15763) );
  NAND2_X1 U17340 ( .A1(n15220), .A2(P3_ADDR_REG_18__SCAN_IN), .ZN(n15761) );
  NAND2_X1 U17341 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(n15759), .ZN(n15760) );
  NAND2_X1 U17342 ( .A1(n15761), .A2(n15760), .ZN(n15762) );
  NOR2_X1 U17343 ( .A1(n15763), .A2(n15762), .ZN(n15766) );
  AOI21_X1 U17344 ( .B1(n15763), .B2(n15762), .A(n15766), .ZN(n15764) );
  INV_X1 U17345 ( .A(n15766), .ZN(n15767) );
  OAI21_X1 U17346 ( .B1(P3_ADDR_REG_18__SCAN_IN), .B2(n15220), .A(n15767), 
        .ZN(n15771) );
  XNOR2_X1 U17347 ( .A(P2_ADDR_REG_19__SCAN_IN), .B(P1_ADDR_REG_19__SCAN_IN), 
        .ZN(n15769) );
  XNOR2_X1 U17348 ( .A(n15769), .B(n15768), .ZN(n15770) );
  XNOR2_X1 U17349 ( .A(n15771), .B(n15770), .ZN(n15772) );
  AOI21_X1 U17350 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(
        P3_WR_REG_SCAN_IN), .ZN(n15773) );
  OAI21_X1 U17351 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(n15773), 
        .ZN(U28) );
  AOI21_X1 U17352 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(
        P3_RD_REG_SCAN_IN), .ZN(n15774) );
  OAI21_X1 U17353 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(n15774), 
        .ZN(U29) );
  XNOR2_X1 U17354 ( .A(n15775), .B(n15776), .ZN(n15866) );
  INV_X1 U17355 ( .A(n15861), .ZN(n15779) );
  XNOR2_X1 U17356 ( .A(n15777), .B(n15776), .ZN(n15778) );
  NOR2_X1 U17357 ( .A1(n15778), .A2(n15826), .ZN(n15863) );
  AOI211_X1 U17358 ( .C1(n15850), .C2(n15866), .A(n15779), .B(n15863), .ZN(
        n15791) );
  INV_X1 U17359 ( .A(n15780), .ZN(n15786) );
  NOR2_X1 U17360 ( .A1(n15804), .A2(n15781), .ZN(n15782) );
  AOI21_X1 U17361 ( .B1(n6556), .B2(P1_REG2_REG_7__SCAN_IN), .A(n15782), .ZN(
        n15783) );
  OAI21_X1 U17362 ( .B1(n15807), .B2(n15786), .A(n15783), .ZN(n15784) );
  INV_X1 U17363 ( .A(n15784), .ZN(n15790) );
  INV_X1 U17364 ( .A(n12206), .ZN(n15787) );
  OAI211_X1 U17365 ( .C1(n15787), .C2(n15786), .A(n7132), .B(n15785), .ZN(
        n15862) );
  INV_X1 U17366 ( .A(n15862), .ZN(n15788) );
  AOI22_X1 U17367 ( .A1(n15866), .A2(n15813), .B1(n15812), .B2(n15788), .ZN(
        n15789) );
  OAI211_X1 U17368 ( .C1(n6556), .C2(n15791), .A(n15790), .B(n15789), .ZN(
        P1_U3286) );
  OAI21_X1 U17369 ( .B1(n12027), .B2(n15793), .A(n15792), .ZN(n15794) );
  OAI21_X1 U17370 ( .B1(n15796), .B2(n15795), .A(n15794), .ZN(n15797) );
  XOR2_X1 U17371 ( .A(n15799), .B(n15797), .Z(n15848) );
  XOR2_X1 U17372 ( .A(n15798), .B(n15799), .Z(n15801) );
  OAI21_X1 U17373 ( .B1(n15801), .B2(n15826), .A(n15800), .ZN(n15802) );
  AOI21_X1 U17374 ( .B1(n15848), .B2(n15850), .A(n15802), .ZN(n15845) );
  NOR2_X1 U17375 ( .A1(n15804), .A2(n15803), .ZN(n15805) );
  AOI21_X1 U17376 ( .B1(n6556), .B2(P1_REG2_REG_5__SCAN_IN), .A(n15805), .ZN(
        n15806) );
  OAI21_X1 U17377 ( .B1(n15807), .B2(n15843), .A(n15806), .ZN(n15808) );
  INV_X1 U17378 ( .A(n15808), .ZN(n15815) );
  OAI211_X1 U17379 ( .C1(n15843), .C2(n6605), .A(n7447), .B(n7132), .ZN(n15842) );
  INV_X1 U17380 ( .A(n15842), .ZN(n15811) );
  AOI22_X1 U17381 ( .A1(n15848), .A2(n15813), .B1(n15812), .B2(n15811), .ZN(
        n15814) );
  OAI211_X1 U17382 ( .C1(n6556), .C2(n15845), .A(n15815), .B(n15814), .ZN(
        P1_U3288) );
  AND2_X1 U17383 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n15821), .ZN(P1_U3294) );
  INV_X1 U17384 ( .A(n15821), .ZN(n15823) );
  NOR2_X1 U17385 ( .A1(n15823), .A2(n15816), .ZN(P1_U3295) );
  AND2_X1 U17386 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n15821), .ZN(P1_U3296) );
  AND2_X1 U17387 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n15821), .ZN(P1_U3297) );
  NOR2_X1 U17388 ( .A1(n15823), .A2(n15817), .ZN(P1_U3298) );
  AND2_X1 U17389 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n15821), .ZN(P1_U3299) );
  AND2_X1 U17390 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n15821), .ZN(P1_U3300) );
  AND2_X1 U17391 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n15821), .ZN(P1_U3301) );
  AND2_X1 U17392 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n15821), .ZN(P1_U3302) );
  AND2_X1 U17393 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n15821), .ZN(P1_U3303) );
  NOR2_X1 U17394 ( .A1(n15823), .A2(n15818), .ZN(P1_U3304) );
  AND2_X1 U17395 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n15821), .ZN(P1_U3305) );
  AND2_X1 U17396 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n15821), .ZN(P1_U3306) );
  AND2_X1 U17397 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n15821), .ZN(P1_U3307) );
  AND2_X1 U17398 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n15821), .ZN(P1_U3308) );
  NOR2_X1 U17399 ( .A1(n15823), .A2(n15819), .ZN(P1_U3309) );
  AND2_X1 U17400 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n15821), .ZN(P1_U3310) );
  AND2_X1 U17401 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n15821), .ZN(P1_U3311) );
  AND2_X1 U17402 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n15821), .ZN(P1_U3312) );
  AND2_X1 U17403 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n15821), .ZN(P1_U3313) );
  AND2_X1 U17404 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n15821), .ZN(P1_U3314) );
  NOR2_X1 U17405 ( .A1(n15823), .A2(n15820), .ZN(P1_U3315) );
  AND2_X1 U17406 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n15821), .ZN(P1_U3316) );
  AND2_X1 U17407 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n15821), .ZN(P1_U3317) );
  AND2_X1 U17408 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n15821), .ZN(P1_U3318) );
  AND2_X1 U17409 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n15821), .ZN(P1_U3319) );
  AND2_X1 U17410 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n15821), .ZN(P1_U3320) );
  AND2_X1 U17411 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n15821), .ZN(P1_U3321) );
  AND2_X1 U17412 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n15821), .ZN(P1_U3322) );
  NOR2_X1 U17413 ( .A1(n15823), .A2(n15822), .ZN(P1_U3323) );
  INV_X1 U17414 ( .A(n15824), .ZN(n15829) );
  AOI21_X1 U17415 ( .B1(n15874), .B2(n15826), .A(n15825), .ZN(n15827) );
  AOI211_X1 U17416 ( .C1(n7137), .C2(n15829), .A(n15828), .B(n15827), .ZN(
        n15878) );
  INV_X1 U17417 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n15830) );
  AOI22_X1 U17418 ( .A1(n15877), .A2(n15878), .B1(n15830), .B2(n15876), .ZN(
        P1_U3459) );
  NAND2_X1 U17419 ( .A1(n15831), .A2(n15851), .ZN(n15833) );
  OAI211_X1 U17420 ( .C1(n15844), .C2(n15834), .A(n15833), .B(n15832), .ZN(
        n15835) );
  NOR2_X1 U17421 ( .A1(n15836), .A2(n15835), .ZN(n15879) );
  AOI22_X1 U17422 ( .A1(n15877), .A2(n15879), .B1(n9507), .B2(n15876), .ZN(
        P1_U3465) );
  OAI21_X1 U17423 ( .B1(n15844), .B2(n7220), .A(n15837), .ZN(n15840) );
  INV_X1 U17424 ( .A(n15838), .ZN(n15839) );
  AOI211_X1 U17425 ( .C1(n15851), .C2(n15841), .A(n15840), .B(n15839), .ZN(
        n15880) );
  AOI22_X1 U17426 ( .A1(n15877), .A2(n15880), .B1(n9525), .B2(n15876), .ZN(
        P1_U3468) );
  OAI21_X1 U17427 ( .B1(n15844), .B2(n15843), .A(n15842), .ZN(n15847) );
  INV_X1 U17428 ( .A(n15845), .ZN(n15846) );
  AOI211_X1 U17429 ( .C1(n15851), .C2(n15848), .A(n15847), .B(n15846), .ZN(
        n15881) );
  INV_X1 U17430 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n15849) );
  AOI22_X1 U17431 ( .A1(n15877), .A2(n15881), .B1(n15849), .B2(n15876), .ZN(
        P1_U3474) );
  NAND2_X1 U17432 ( .A1(n15852), .A2(n15850), .ZN(n15857) );
  NAND2_X1 U17433 ( .A1(n15852), .A2(n15851), .ZN(n15856) );
  NAND2_X1 U17434 ( .A1(n15870), .A2(n15853), .ZN(n15854) );
  AND4_X1 U17435 ( .A1(n15857), .A2(n15856), .A3(n15855), .A4(n15854), .ZN(
        n15858) );
  AND2_X1 U17436 ( .A1(n15859), .A2(n15858), .ZN(n15882) );
  AOI22_X1 U17437 ( .A1(n15877), .A2(n15882), .B1(n9575), .B2(n15876), .ZN(
        P1_U3477) );
  NAND3_X1 U17438 ( .A1(n15862), .A2(n15861), .A3(n15860), .ZN(n15864) );
  AOI211_X1 U17439 ( .C1(n15866), .C2(n15865), .A(n15864), .B(n15863), .ZN(
        n15883) );
  INV_X1 U17440 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n15867) );
  AOI22_X1 U17441 ( .A1(n15877), .A2(n15883), .B1(n15867), .B2(n15876), .ZN(
        P1_U3480) );
  AOI21_X1 U17442 ( .B1(n15870), .B2(n15869), .A(n15868), .ZN(n15871) );
  OAI211_X1 U17443 ( .C1(n15874), .C2(n15873), .A(n15872), .B(n15871), .ZN(
        n15875) );
  INV_X1 U17444 ( .A(n15875), .ZN(n15885) );
  AOI22_X1 U17445 ( .A1(n15877), .A2(n15885), .B1(n9611), .B2(n15876), .ZN(
        P1_U3483) );
  AOI22_X1 U17446 ( .A1(n15886), .A2(n15878), .B1(n10725), .B2(n15884), .ZN(
        P1_U3528) );
  AOI22_X1 U17447 ( .A1(n15886), .A2(n15879), .B1(n9508), .B2(n15884), .ZN(
        P1_U3530) );
  AOI22_X1 U17448 ( .A1(n15886), .A2(n15880), .B1(n11064), .B2(n15884), .ZN(
        P1_U3531) );
  AOI22_X1 U17449 ( .A1(n15886), .A2(n15881), .B1(n9560), .B2(n15884), .ZN(
        P1_U3533) );
  AOI22_X1 U17450 ( .A1(n15886), .A2(n15882), .B1(n11091), .B2(n15884), .ZN(
        P1_U3534) );
  AOI22_X1 U17451 ( .A1(n15886), .A2(n15883), .B1(n9593), .B2(n15884), .ZN(
        P1_U3535) );
  AOI22_X1 U17452 ( .A1(n15886), .A2(n15885), .B1(n9607), .B2(n15884), .ZN(
        P1_U3536) );
  NOR2_X1 U17453 ( .A1(n15899), .A2(n15887), .ZN(P2_U3087) );
  AOI22_X1 U17454 ( .A1(n15899), .A2(P2_ADDR_REG_1__SCAN_IN), .B1(
        P2_REG3_REG_1__SCAN_IN), .B2(P2_U3088), .ZN(n15898) );
  XNOR2_X1 U17455 ( .A(n15889), .B(n15888), .ZN(n15890) );
  OR2_X1 U17456 ( .A1(n15904), .A2(n15890), .ZN(n15892) );
  OR2_X1 U17457 ( .A1(n15919), .A2(n8035), .ZN(n15891) );
  AND2_X1 U17458 ( .A1(n15892), .A2(n15891), .ZN(n15897) );
  OAI211_X1 U17459 ( .C1(n15895), .C2(n15894), .A(n15937), .B(n15893), .ZN(
        n15896) );
  NAND3_X1 U17460 ( .A1(n15898), .A2(n15897), .A3(n15896), .ZN(P2_U3215) );
  AOI22_X1 U17461 ( .A1(n15899), .A2(P2_ADDR_REG_2__SCAN_IN), .B1(
        P2_REG3_REG_2__SCAN_IN), .B2(P2_U3088), .ZN(n15912) );
  OAI21_X1 U17462 ( .B1(n15902), .B2(n15901), .A(n15900), .ZN(n15903) );
  OR2_X1 U17463 ( .A1(n15904), .A2(n15903), .ZN(n15906) );
  OR2_X1 U17464 ( .A1(n15919), .A2(n8053), .ZN(n15905) );
  AND2_X1 U17465 ( .A1(n15906), .A2(n15905), .ZN(n15911) );
  OAI211_X1 U17466 ( .C1(n15909), .C2(n15908), .A(n15937), .B(n15907), .ZN(
        n15910) );
  NAND3_X1 U17467 ( .A1(n15912), .A2(n15911), .A3(n15910), .ZN(P2_U3216) );
  INV_X1 U17468 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n15926) );
  OAI211_X1 U17469 ( .C1(n15915), .C2(n15914), .A(n15928), .B(n15913), .ZN(
        n15917) );
  OAI211_X1 U17470 ( .C1(n15919), .C2(n15918), .A(n15917), .B(n15916), .ZN(
        n15920) );
  INV_X1 U17471 ( .A(n15920), .ZN(n15925) );
  OAI211_X1 U17472 ( .C1(n15923), .C2(n15922), .A(n15937), .B(n15921), .ZN(
        n15924) );
  OAI211_X1 U17473 ( .C1(n15944), .C2(n15926), .A(n15925), .B(n15924), .ZN(
        P2_U3220) );
  NOR2_X1 U17474 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n15927), .ZN(n15934) );
  OAI211_X1 U17475 ( .C1(n15931), .C2(n15930), .A(n15929), .B(n15928), .ZN(
        n15932) );
  INV_X1 U17476 ( .A(n15932), .ZN(n15933) );
  AOI211_X1 U17477 ( .C1(n15936), .C2(n15935), .A(n15934), .B(n15933), .ZN(
        n15942) );
  OAI211_X1 U17478 ( .C1(n15940), .C2(n15939), .A(n15938), .B(n15937), .ZN(
        n15941) );
  OAI211_X1 U17479 ( .C1(n15944), .C2(n15943), .A(n15942), .B(n15941), .ZN(
        P2_U3230) );
  INV_X1 U17480 ( .A(n15981), .ZN(n15979) );
  INV_X1 U17481 ( .A(P2_D_REG_31__SCAN_IN), .ZN(n15946) );
  NOR2_X1 U17482 ( .A1(n15977), .A2(n15946), .ZN(P2_U3266) );
  NOR2_X1 U17483 ( .A1(n15977), .A2(n15947), .ZN(P2_U3267) );
  NOR2_X1 U17484 ( .A1(n15977), .A2(n15948), .ZN(P2_U3268) );
  INV_X1 U17485 ( .A(P2_D_REG_28__SCAN_IN), .ZN(n15949) );
  NOR2_X1 U17486 ( .A1(n15977), .A2(n15949), .ZN(P2_U3269) );
  INV_X1 U17487 ( .A(P2_D_REG_27__SCAN_IN), .ZN(n15950) );
  NOR2_X1 U17488 ( .A1(n15960), .A2(n15950), .ZN(P2_U3270) );
  NOR2_X1 U17489 ( .A1(n15960), .A2(n15951), .ZN(P2_U3271) );
  INV_X1 U17490 ( .A(P2_D_REG_25__SCAN_IN), .ZN(n15952) );
  NOR2_X1 U17491 ( .A1(n15960), .A2(n15952), .ZN(P2_U3272) );
  INV_X1 U17492 ( .A(P2_D_REG_24__SCAN_IN), .ZN(n15953) );
  NOR2_X1 U17493 ( .A1(n15960), .A2(n15953), .ZN(P2_U3273) );
  INV_X1 U17494 ( .A(P2_D_REG_23__SCAN_IN), .ZN(n15954) );
  NOR2_X1 U17495 ( .A1(n15960), .A2(n15954), .ZN(P2_U3274) );
  INV_X1 U17496 ( .A(P2_D_REG_22__SCAN_IN), .ZN(n15955) );
  NOR2_X1 U17497 ( .A1(n15960), .A2(n15955), .ZN(P2_U3275) );
  INV_X1 U17498 ( .A(P2_D_REG_21__SCAN_IN), .ZN(n15956) );
  NOR2_X1 U17499 ( .A1(n15960), .A2(n15956), .ZN(P2_U3276) );
  INV_X1 U17500 ( .A(P2_D_REG_20__SCAN_IN), .ZN(n15957) );
  NOR2_X1 U17501 ( .A1(n15960), .A2(n15957), .ZN(P2_U3277) );
  INV_X1 U17502 ( .A(P2_D_REG_19__SCAN_IN), .ZN(n15958) );
  NOR2_X1 U17503 ( .A1(n15960), .A2(n15958), .ZN(P2_U3278) );
  INV_X1 U17504 ( .A(P2_D_REG_18__SCAN_IN), .ZN(n15959) );
  NOR2_X1 U17505 ( .A1(n15960), .A2(n15959), .ZN(P2_U3279) );
  INV_X1 U17506 ( .A(P2_D_REG_17__SCAN_IN), .ZN(n15961) );
  NOR2_X1 U17507 ( .A1(n15977), .A2(n15961), .ZN(P2_U3280) );
  INV_X1 U17508 ( .A(P2_D_REG_16__SCAN_IN), .ZN(n15962) );
  NOR2_X1 U17509 ( .A1(n15977), .A2(n15962), .ZN(P2_U3281) );
  INV_X1 U17510 ( .A(P2_D_REG_15__SCAN_IN), .ZN(n15963) );
  NOR2_X1 U17511 ( .A1(n15977), .A2(n15963), .ZN(P2_U3282) );
  INV_X1 U17512 ( .A(P2_D_REG_14__SCAN_IN), .ZN(n15964) );
  NOR2_X1 U17513 ( .A1(n15977), .A2(n15964), .ZN(P2_U3283) );
  INV_X1 U17514 ( .A(P2_D_REG_13__SCAN_IN), .ZN(n15965) );
  NOR2_X1 U17515 ( .A1(n15977), .A2(n15965), .ZN(P2_U3284) );
  INV_X1 U17516 ( .A(P2_D_REG_12__SCAN_IN), .ZN(n15966) );
  NOR2_X1 U17517 ( .A1(n15977), .A2(n15966), .ZN(P2_U3285) );
  NOR2_X1 U17518 ( .A1(n15977), .A2(n15967), .ZN(P2_U3286) );
  INV_X1 U17519 ( .A(P2_D_REG_10__SCAN_IN), .ZN(n15968) );
  NOR2_X1 U17520 ( .A1(n15977), .A2(n15968), .ZN(P2_U3287) );
  INV_X1 U17521 ( .A(P2_D_REG_9__SCAN_IN), .ZN(n15969) );
  NOR2_X1 U17522 ( .A1(n15977), .A2(n15969), .ZN(P2_U3288) );
  INV_X1 U17523 ( .A(P2_D_REG_8__SCAN_IN), .ZN(n15970) );
  NOR2_X1 U17524 ( .A1(n15977), .A2(n15970), .ZN(P2_U3289) );
  INV_X1 U17525 ( .A(P2_D_REG_7__SCAN_IN), .ZN(n15971) );
  NOR2_X1 U17526 ( .A1(n15977), .A2(n15971), .ZN(P2_U3290) );
  INV_X1 U17527 ( .A(P2_D_REG_6__SCAN_IN), .ZN(n15972) );
  NOR2_X1 U17528 ( .A1(n15977), .A2(n15972), .ZN(P2_U3291) );
  INV_X1 U17529 ( .A(P2_D_REG_5__SCAN_IN), .ZN(n15973) );
  NOR2_X1 U17530 ( .A1(n15977), .A2(n15973), .ZN(P2_U3292) );
  NOR2_X1 U17531 ( .A1(n15977), .A2(n15974), .ZN(P2_U3293) );
  INV_X1 U17532 ( .A(P2_D_REG_3__SCAN_IN), .ZN(n15975) );
  NOR2_X1 U17533 ( .A1(n15977), .A2(n15975), .ZN(P2_U3294) );
  INV_X1 U17534 ( .A(P2_D_REG_2__SCAN_IN), .ZN(n15976) );
  NOR2_X1 U17535 ( .A1(n15977), .A2(n15976), .ZN(P2_U3295) );
  MUX2_X1 U17536 ( .A(P2_D_REG_0__SCAN_IN), .B(n15978), .S(n15977), .Z(
        P2_U3416) );
  AOI22_X1 U17537 ( .A1(n15981), .A2(n15980), .B1(n8682), .B2(n15979), .ZN(
        P2_U3417) );
  AOI21_X1 U17538 ( .B1(n15996), .B2(n15983), .A(n15982), .ZN(n15984) );
  OAI211_X1 U17539 ( .C1(n15986), .C2(n16000), .A(n15985), .B(n15984), .ZN(
        n15987) );
  INV_X1 U17540 ( .A(n15987), .ZN(n16006) );
  AOI22_X1 U17541 ( .A1(n16004), .A2(n16006), .B1(n8118), .B2(n16002), .ZN(
        P2_U3445) );
  OAI21_X1 U17542 ( .B1(n7900), .B2(n15989), .A(n15988), .ZN(n15991) );
  AOI211_X1 U17543 ( .C1(n15993), .C2(n15992), .A(n15991), .B(n15990), .ZN(
        n16007) );
  AOI22_X1 U17544 ( .A1(n16004), .A2(n16007), .B1(n8109), .B2(n16002), .ZN(
        P2_U3448) );
  AOI21_X1 U17545 ( .B1(n15996), .B2(n15995), .A(n15994), .ZN(n15998) );
  OAI211_X1 U17546 ( .C1(n16000), .C2(n15999), .A(n15998), .B(n15997), .ZN(
        n16001) );
  INV_X1 U17547 ( .A(n16001), .ZN(n16010) );
  INV_X1 U17548 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n16003) );
  AOI22_X1 U17549 ( .A1(n16004), .A2(n16010), .B1(n16003), .B2(n16002), .ZN(
        P2_U3451) );
  AOI22_X1 U17550 ( .A1(n16011), .A2(n16006), .B1(n16005), .B2(n16008), .ZN(
        P2_U3504) );
  AOI22_X1 U17551 ( .A1(n16011), .A2(n16007), .B1(n11138), .B2(n16008), .ZN(
        P2_U3505) );
  AOI22_X1 U17552 ( .A1(n16011), .A2(n16010), .B1(n16009), .B2(n16008), .ZN(
        P2_U3506) );
  NOR2_X1 U17553 ( .A1(P3_U3897), .A2(n16012), .ZN(P3_U3150) );
  NAND3_X1 U17554 ( .A1(n16015), .A2(n16014), .A3(n16013), .ZN(n16019) );
  OAI21_X1 U17555 ( .B1(P3_IR_REG_0__SCAN_IN), .B2(n16017), .A(n16016), .ZN(
        n16018) );
  NAND2_X1 U17556 ( .A1(n16019), .A2(n16018), .ZN(n16023) );
  AOI22_X1 U17557 ( .A1(n16021), .A2(P3_IR_REG_0__SCAN_IN), .B1(
        P3_REG3_REG_0__SCAN_IN), .B2(P3_U3151), .ZN(n16022) );
  OAI211_X1 U17558 ( .C1(n10608), .C2(n16024), .A(n16023), .B(n16022), .ZN(
        P3_U3182) );
  XNOR2_X1 U17559 ( .A(n16027), .B(n16025), .ZN(n16035) );
  OR2_X1 U17560 ( .A1(n16027), .A2(n16026), .ZN(n16028) );
  NAND2_X1 U17561 ( .A1(n16029), .A2(n16028), .ZN(n16073) );
  NAND2_X1 U17562 ( .A1(n16073), .A2(n16054), .ZN(n16033) );
  AOI22_X1 U17563 ( .A1(n16046), .A2(n16031), .B1(n7149), .B2(n16049), .ZN(
        n16032) );
  OAI211_X1 U17564 ( .C1(n16035), .C2(n16034), .A(n16033), .B(n16032), .ZN(
        n16071) );
  INV_X1 U17565 ( .A(n16073), .ZN(n16040) );
  NOR2_X1 U17566 ( .A1(n16036), .A2(n16055), .ZN(n16072) );
  INV_X1 U17567 ( .A(n16072), .ZN(n16037) );
  OAI22_X1 U17568 ( .A1(n16040), .A2(n16039), .B1(n16038), .B2(n16037), .ZN(
        n16041) );
  AOI211_X1 U17569 ( .C1(P3_REG3_REG_2__SCAN_IN), .C2(n16061), .A(n16071), .B(
        n16041), .ZN(n16042) );
  AOI22_X1 U17570 ( .A1(n16066), .A2(n7654), .B1(n16042), .B2(n9401), .ZN(
        P3_U3231) );
  XNOR2_X1 U17571 ( .A(n16052), .B(n16043), .ZN(n16045) );
  NAND2_X1 U17572 ( .A1(n16045), .A2(n16044), .ZN(n16051) );
  AOI22_X1 U17573 ( .A1(n16049), .A2(n16048), .B1(n16047), .B2(n16046), .ZN(
        n16050) );
  NAND2_X1 U17574 ( .A1(n16051), .A2(n16050), .ZN(n16067) );
  INV_X1 U17575 ( .A(n16067), .ZN(n16060) );
  XNOR2_X1 U17576 ( .A(n16052), .B(n16053), .ZN(n16069) );
  NAND2_X1 U17577 ( .A1(n16069), .A2(n16054), .ZN(n16059) );
  NOR2_X1 U17578 ( .A1(n16056), .A2(n16055), .ZN(n16068) );
  NAND2_X1 U17579 ( .A1(n16068), .A2(n16057), .ZN(n16058) );
  AND3_X1 U17580 ( .A1(n16060), .A2(n16059), .A3(n16058), .ZN(n16065) );
  AOI22_X1 U17581 ( .A1(n16062), .A2(n16069), .B1(P3_REG3_REG_1__SCAN_IN), 
        .B2(n16061), .ZN(n16063) );
  OAI221_X1 U17582 ( .B1(n16066), .B2(n16065), .C1(n9401), .C2(n16064), .A(
        n16063), .ZN(P3_U3232) );
  AOI211_X1 U17583 ( .C1(n16070), .C2(n16069), .A(n16068), .B(n16067), .ZN(
        n16096) );
  AOI22_X1 U17584 ( .A1(n16094), .A2(n16096), .B1(n7172), .B2(n16092), .ZN(
        P3_U3393) );
  AOI211_X1 U17585 ( .C1(n16090), .C2(n16073), .A(n16072), .B(n16071), .ZN(
        n16074) );
  INV_X1 U17586 ( .A(n16074), .ZN(n16097) );
  OAI22_X1 U17587 ( .A1(n16092), .A2(n16097), .B1(P3_REG0_REG_2__SCAN_IN), 
        .B2(n16094), .ZN(n16075) );
  INV_X1 U17588 ( .A(n16075), .ZN(P3_U3396) );
  INV_X1 U17589 ( .A(n16076), .ZN(n16079) );
  AND2_X1 U17590 ( .A1(n16077), .A2(n16090), .ZN(n16078) );
  NOR3_X1 U17591 ( .A1(n16080), .A2(n16079), .A3(n16078), .ZN(n16100) );
  INV_X1 U17592 ( .A(P3_REG0_REG_5__SCAN_IN), .ZN(n16081) );
  AOI22_X1 U17593 ( .A1(n16094), .A2(n16100), .B1(n16081), .B2(n16092), .ZN(
        P3_U3405) );
  INV_X1 U17594 ( .A(n16082), .ZN(n16083) );
  AOI211_X1 U17595 ( .C1(n16085), .C2(n16090), .A(n16084), .B(n16083), .ZN(
        n16102) );
  INV_X1 U17596 ( .A(P3_REG0_REG_7__SCAN_IN), .ZN(n16086) );
  AOI22_X1 U17597 ( .A1(n16094), .A2(n16102), .B1(n16086), .B2(n16092), .ZN(
        P3_U3411) );
  INV_X1 U17598 ( .A(n16087), .ZN(n16088) );
  AOI211_X1 U17599 ( .C1(n16091), .C2(n16090), .A(n16089), .B(n16088), .ZN(
        n16105) );
  INV_X1 U17600 ( .A(P3_REG0_REG_8__SCAN_IN), .ZN(n16093) );
  AOI22_X1 U17601 ( .A1(n16094), .A2(n16105), .B1(n16093), .B2(n16092), .ZN(
        P3_U3414) );
  AOI22_X1 U17602 ( .A1(n16106), .A2(n16096), .B1(n16095), .B2(n16103), .ZN(
        P3_U3460) );
  OAI22_X1 U17603 ( .A1(n16103), .A2(n16097), .B1(P3_REG1_REG_2__SCAN_IN), 
        .B2(n16106), .ZN(n16098) );
  INV_X1 U17604 ( .A(n16098), .ZN(P3_U3461) );
  AOI22_X1 U17605 ( .A1(n16106), .A2(n16100), .B1(n16099), .B2(n16103), .ZN(
        P3_U3464) );
  AOI22_X1 U17606 ( .A1(n16106), .A2(n16102), .B1(n16101), .B2(n16103), .ZN(
        P3_U3466) );
  AOI22_X1 U17607 ( .A1(n16106), .A2(n16105), .B1(n16104), .B2(n16103), .ZN(
        P3_U3467) );
  BUF_X1 U12132 ( .A(n9451), .Z(n13135) );
  CLKBUF_X3 U9963 ( .A(n8071), .Z(n8553) );
  INV_X1 U10645 ( .A(n8141), .ZN(n8521) );
  CLKBUF_X2 U7303 ( .A(n13292), .Z(n6569) );
  CLKBUF_X2 U7328 ( .A(n8809), .Z(n8895) );
  CLKBUF_X1 U7355 ( .A(n8554), .Z(n8643) );
  NAND2_X1 U7366 ( .A1(n8008), .A2(n14904), .ZN(n8376) );
  NAND2_X1 U7367 ( .A1(n13135), .A2(n9450), .ZN(n9526) );
  CLKBUF_X2 U7392 ( .A(n13294), .Z(n6564) );
  BUF_X2 U7524 ( .A(n9526), .Z(n6553) );
  OR3_X1 U8041 ( .A1(n9459), .A2(n9447), .A3(n9444), .ZN(n7792) );
  CLKBUF_X1 U9189 ( .A(n15960), .Z(n15977) );
endmodule

