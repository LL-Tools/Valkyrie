

module b21_C_lock ( keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, 
        keyinput_5, keyinput_6, keyinput_7, keyinput_8, keyinput_9, 
        keyinput_10, keyinput_11, keyinput_12, keyinput_13, keyinput_14, 
        keyinput_15, keyinput_16, keyinput_17, keyinput_18, keyinput_19, 
        keyinput_20, keyinput_21, keyinput_22, keyinput_23, keyinput_24, 
        keyinput_25, keyinput_26, keyinput_27, keyinput_28, keyinput_29, 
        keyinput_30, keyinput_31, keyinput_32, keyinput_33, keyinput_34, 
        keyinput_35, keyinput_36, keyinput_37, keyinput_38, keyinput_39, 
        keyinput_40, keyinput_41, keyinput_42, keyinput_43, keyinput_44, 
        keyinput_45, keyinput_46, keyinput_47, keyinput_48, keyinput_49, 
        keyinput_50, keyinput_51, keyinput_52, keyinput_53, keyinput_54, 
        keyinput_55, keyinput_56, keyinput_57, keyinput_58, keyinput_59, 
        keyinput_60, keyinput_61, keyinput_62, keyinput_63, keyinput_64, 
        keyinput_65, keyinput_66, keyinput_67, keyinput_68, keyinput_69, 
        keyinput_70, keyinput_71, keyinput_72, keyinput_73, keyinput_74, 
        keyinput_75, keyinput_76, keyinput_77, keyinput_78, keyinput_79, 
        keyinput_80, keyinput_81, keyinput_82, keyinput_83, keyinput_84, 
        keyinput_85, keyinput_86, keyinput_87, keyinput_88, keyinput_89, 
        keyinput_90, keyinput_91, keyinput_92, keyinput_93, keyinput_94, 
        keyinput_95, keyinput_96, keyinput_97, keyinput_98, keyinput_99, 
        keyinput_100, keyinput_101, keyinput_102, keyinput_103, keyinput_104, 
        keyinput_105, keyinput_106, keyinput_107, keyinput_108, keyinput_109, 
        keyinput_110, keyinput_111, keyinput_112, keyinput_113, keyinput_114, 
        keyinput_115, keyinput_116, keyinput_117, keyinput_118, keyinput_119, 
        keyinput_120, keyinput_121, keyinput_122, keyinput_123, keyinput_124, 
        keyinput_125, keyinput_126, keyinput_127, P2_WR_REG_SCAN_IN, SI_31_, 
        SI_30_, SI_29_, SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, 
        SI_21_, SI_20_, SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, 
        SI_12_, SI_11_, SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, 
        SI_3_, SI_2_, SI_1_, SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, 
        P2_REG3_REG_7__SCAN_IN, P2_REG3_REG_27__SCAN_IN, 
        P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_23__SCAN_IN, 
        P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_3__SCAN_IN, 
        P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_28__SCAN_IN, 
        P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_1__SCAN_IN, 
        P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_12__SCAN_IN, 
        P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_16__SCAN_IN, 
        P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_17__SCAN_IN, 
        P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_4__SCAN_IN, 
        P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, 
        P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, 
        P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, 
        P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, 
        P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, 
        P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, 
        P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, 
        P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, 
        P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, 
        P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, 
        P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, 
        P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, 
        P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, 
        P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, 
        P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, 
        P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, 
        P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, 
        P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, 
        P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, 
        P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, 
        P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, 
        P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, 
        P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, 
        P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, 
        P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, 
        ADD_1071_U57, ADD_1071_U58, ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, 
        ADD_1071_U62, ADD_1071_U63, ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, 
        ADD_1071_U50, ADD_1071_U51, ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, 
        ADD_1071_U5, ADD_1071_U46, U126, U123, P1_U3353, P1_U3352, P1_U3351, 
        P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, 
        P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, 
        P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, 
        P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, 
        P1_U3322, P1_U3440, P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, 
        P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, 
        P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, 
        P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, 
        P1_U3296, P1_U3295, P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, 
        P1_U3460, P1_U3463, P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, 
        P1_U3481, P1_U3484, P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, 
        P1_U3502, P1_U3505, P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, 
        P1_U3514, P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, 
        P1_U3521, P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, 
        P1_U3528, P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, 
        P1_U3535, P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, 
        P1_U3542, P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, 
        P1_U3549, P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, 
        P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, 
        P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, 
        P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, 
        P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, 
        P1_U3355, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, 
        P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, 
        P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, 
        P1_U3242, P1_U3241, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, 
        P1_U3560, P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, 
        P1_U3567, P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, 
        P1_U3574, P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, 
        P1_U3581, P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, 
        P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, 
        P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, 
        P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, 
        P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, 
        P1_U3211, P1_U3084, P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, 
        P2_U3355, P2_U3354, P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, 
        P2_U3348, P2_U3347, P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, 
        P2_U3341, P2_U3340, P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, 
        P2_U3334, P2_U3333, P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, 
        P2_U3327, P2_U3437, P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, 
        P2_U3322, P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, 
        P2_U3315, P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, 
        P2_U3308, P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, 
        P2_U3301, P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, 
        P2_U3457, P2_U3460, P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, 
        P2_U3478, P2_U3481, P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, 
        P2_U3499, P2_U3502, P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, 
        P2_U3511, P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, 
        P2_U3518, P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, 
        P2_U3525, P2_U3526, P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, 
        P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, 
        P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, 
        P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, 
        P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, 
        P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, 
        P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, 
        P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, 
        P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, 
        P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, 
        P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, 
        P2_U3246, P2_U3245, P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, 
        P2_U3557, P2_U3558, P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, 
        P2_U3564, P2_U3565, P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, 
        P2_U3571, P2_U3572, P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, 
        P2_U3578, P2_U3579, P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, 
        P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, 
        P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, 
        P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, 
        P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, 
        P2_U3215, P2_U3152, P2_U3151, P2_U3966 );
  input keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, keyinput_5,
         keyinput_6, keyinput_7, keyinput_8, keyinput_9, keyinput_10,
         keyinput_11, keyinput_12, keyinput_13, keyinput_14, keyinput_15,
         keyinput_16, keyinput_17, keyinput_18, keyinput_19, keyinput_20,
         keyinput_21, keyinput_22, keyinput_23, keyinput_24, keyinput_25,
         keyinput_26, keyinput_27, keyinput_28, keyinput_29, keyinput_30,
         keyinput_31, keyinput_32, keyinput_33, keyinput_34, keyinput_35,
         keyinput_36, keyinput_37, keyinput_38, keyinput_39, keyinput_40,
         keyinput_41, keyinput_42, keyinput_43, keyinput_44, keyinput_45,
         keyinput_46, keyinput_47, keyinput_48, keyinput_49, keyinput_50,
         keyinput_51, keyinput_52, keyinput_53, keyinput_54, keyinput_55,
         keyinput_56, keyinput_57, keyinput_58, keyinput_59, keyinput_60,
         keyinput_61, keyinput_62, keyinput_63, keyinput_64, keyinput_65,
         keyinput_66, keyinput_67, keyinput_68, keyinput_69, keyinput_70,
         keyinput_71, keyinput_72, keyinput_73, keyinput_74, keyinput_75,
         keyinput_76, keyinput_77, keyinput_78, keyinput_79, keyinput_80,
         keyinput_81, keyinput_82, keyinput_83, keyinput_84, keyinput_85,
         keyinput_86, keyinput_87, keyinput_88, keyinput_89, keyinput_90,
         keyinput_91, keyinput_92, keyinput_93, keyinput_94, keyinput_95,
         keyinput_96, keyinput_97, keyinput_98, keyinput_99, keyinput_100,
         keyinput_101, keyinput_102, keyinput_103, keyinput_104, keyinput_105,
         keyinput_106, keyinput_107, keyinput_108, keyinput_109, keyinput_110,
         keyinput_111, keyinput_112, keyinput_113, keyinput_114, keyinput_115,
         keyinput_116, keyinput_117, keyinput_118, keyinput_119, keyinput_120,
         keyinput_121, keyinput_122, keyinput_123, keyinput_124, keyinput_125,
         keyinput_126, keyinput_127, P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_,
         SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_,
         SI_20_, SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_,
         SI_12_, SI_11_, SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_,
         SI_3_, SI_2_, SI_1_, SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN,
         P2_REG3_REG_7__SCAN_IN, P2_REG3_REG_27__SCAN_IN,
         P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_23__SCAN_IN,
         P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_3__SCAN_IN,
         P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_28__SCAN_IN,
         P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_1__SCAN_IN,
         P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_12__SCAN_IN,
         P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_16__SCAN_IN,
         P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_17__SCAN_IN,
         P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_4__SCAN_IN,
         P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN,
         P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN,
         P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN,
         P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN,
         P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN,
         P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN,
         P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN,
         P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN,
         P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN,
         P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN,
         P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN,
         P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN,
         P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN,
         P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN,
         P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN,
         P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN,
         P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN,
         P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN,
         P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN,
         P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN,
         P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN,
         P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN,
         P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN,
         P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN,
         P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN,
         P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN,
         P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN,
         P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN,
         P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN,
         P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN,
         P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN,
         P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN,
         P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN,
         P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN,
         P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN,
         P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN,
         P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN,
         P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN,
         P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN,
         P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN,
         P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN,
         P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN,
         P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN,
         P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN,
         P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN,
         P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN,
         P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN,
         P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN,
         P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN,
         P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN,
         P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN,
         P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN,
         P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN,
         P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN,
         P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN,
         P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN,
         P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN,
         P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN,
         P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN,
         P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN,
         P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN,
         P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN,
         P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN,
         P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN,
         P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN,
         P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN,
         P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN,
         P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN,
         P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN,
         P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN,
         P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN,
         P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN,
         P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN,
         P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN,
         P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN,
         P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN,
         P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN,
         P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN,
         P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN,
         P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN,
         P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN,
         P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN,
         P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN,
         P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN,
         P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN,
         P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN,
         P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN,
         P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN,
         P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN,
         P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN,
         P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN,
         P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN,
         P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN,
         P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN,
         P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN,
         P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN,
         P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN,
         P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN,
         P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN,
         P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN,
         P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN,
         P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN,
         P1_REG3_REG_4__SCAN_IN, P1_REG3_REG_24__SCAN_IN,
         P1_REG3_REG_17__SCAN_IN, P1_REG3_REG_5__SCAN_IN,
         P1_REG3_REG_16__SCAN_IN, P1_REG3_REG_25__SCAN_IN,
         P1_REG3_REG_12__SCAN_IN, P1_REG3_REG_21__SCAN_IN,
         P1_REG3_REG_1__SCAN_IN, P1_REG3_REG_8__SCAN_IN,
         P1_REG3_REG_28__SCAN_IN, P1_REG3_REG_19__SCAN_IN,
         P1_REG3_REG_3__SCAN_IN, P1_REG3_REG_10__SCAN_IN,
         P1_REG3_REG_23__SCAN_IN, P1_REG3_REG_14__SCAN_IN,
         P1_REG3_REG_27__SCAN_IN, P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN,
         P1_RD_REG_SCAN_IN, P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN,
         P2_IR_REG_1__SCAN_IN, P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN,
         P2_IR_REG_4__SCAN_IN, P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN,
         P2_IR_REG_7__SCAN_IN, P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN,
         P2_IR_REG_10__SCAN_IN, P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN,
         P2_IR_REG_13__SCAN_IN, P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN,
         P2_IR_REG_16__SCAN_IN, P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN,
         P2_IR_REG_19__SCAN_IN, P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN,
         P2_IR_REG_22__SCAN_IN, P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN,
         P2_IR_REG_25__SCAN_IN, P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN,
         P2_IR_REG_28__SCAN_IN, P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN,
         P2_IR_REG_31__SCAN_IN, P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN,
         P2_D_REG_2__SCAN_IN, P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN,
         P2_D_REG_5__SCAN_IN, P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN,
         P2_D_REG_8__SCAN_IN, P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN,
         P2_D_REG_11__SCAN_IN, P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN,
         P2_D_REG_14__SCAN_IN, P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN,
         P2_D_REG_17__SCAN_IN, P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN,
         P2_D_REG_20__SCAN_IN, P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN,
         P2_D_REG_23__SCAN_IN, P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN,
         P2_D_REG_26__SCAN_IN, P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN,
         P2_D_REG_29__SCAN_IN, P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN,
         P2_REG0_REG_0__SCAN_IN, P2_REG0_REG_1__SCAN_IN,
         P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN,
         P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN,
         P2_REG0_REG_6__SCAN_IN, P2_REG0_REG_7__SCAN_IN,
         P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN,
         P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN,
         P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN,
         P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN,
         P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN,
         P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN,
         P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN,
         P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN,
         P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN,
         P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN,
         P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN,
         P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN,
         P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN,
         P2_REG1_REG_2__SCAN_IN, P2_REG1_REG_3__SCAN_IN,
         P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN,
         P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN,
         P2_REG1_REG_8__SCAN_IN, P2_REG1_REG_9__SCAN_IN,
         P2_REG1_REG_10__SCAN_IN, P2_REG1_REG_11__SCAN_IN,
         P2_REG1_REG_12__SCAN_IN, P2_REG1_REG_13__SCAN_IN,
         P2_REG1_REG_14__SCAN_IN, P2_REG1_REG_15__SCAN_IN,
         P2_REG1_REG_16__SCAN_IN, P2_REG1_REG_17__SCAN_IN,
         P2_REG1_REG_18__SCAN_IN, P2_REG1_REG_19__SCAN_IN,
         P2_REG1_REG_20__SCAN_IN, P2_REG1_REG_21__SCAN_IN,
         P2_REG1_REG_22__SCAN_IN, P2_REG1_REG_23__SCAN_IN,
         P2_REG1_REG_24__SCAN_IN, P2_REG1_REG_25__SCAN_IN,
         P2_REG1_REG_26__SCAN_IN, P2_REG1_REG_27__SCAN_IN,
         P2_REG1_REG_28__SCAN_IN, P2_REG1_REG_29__SCAN_IN,
         P2_REG1_REG_30__SCAN_IN, P2_REG1_REG_31__SCAN_IN,
         P2_REG2_REG_0__SCAN_IN, P2_REG2_REG_1__SCAN_IN,
         P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN,
         P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN,
         P2_REG2_REG_6__SCAN_IN, P2_REG2_REG_7__SCAN_IN,
         P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN,
         P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN,
         P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN,
         P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN,
         P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN,
         P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN,
         P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN,
         P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN,
         P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN,
         P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN,
         P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN,
         P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN,
         P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN,
         P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN,
         P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN,
         P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN,
         P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN,
         P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN,
         P2_ADDR_REG_7__SCAN_IN, P2_ADDR_REG_6__SCAN_IN,
         P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN,
         P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN,
         P2_ADDR_REG_1__SCAN_IN, P2_ADDR_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN;
  output ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, ADD_1071_U57, ADD_1071_U58,
         ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, ADD_1071_U62, ADD_1071_U63,
         ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, ADD_1071_U50, ADD_1071_U51,
         ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, ADD_1071_U5, ADD_1071_U46,
         U126, U123, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349,
         P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342,
         P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335,
         P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328,
         P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, P1_U3322, P1_U3440,
         P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316,
         P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309,
         P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302,
         P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295,
         P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, P1_U3460, P1_U3463,
         P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, P1_U3481, P1_U3484,
         P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, P1_U3502, P1_U3505,
         P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515,
         P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522,
         P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529,
         P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536,
         P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543,
         P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550,
         P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, P1_U3290, P1_U3289,
         P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282,
         P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275,
         P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268,
         P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, P1_U3355, P1_U3262,
         P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255,
         P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248,
         P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3242, P1_U3241,
         P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561,
         P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568,
         P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575,
         P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582,
         P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, P1_U3239, P1_U3238,
         P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231,
         P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224,
         P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217,
         P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, P1_U3084,
         P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, P2_U3355, P2_U3354,
         P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, P2_U3348, P2_U3347,
         P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, P2_U3341, P2_U3340,
         P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, P2_U3334, P2_U3333,
         P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, P2_U3327, P2_U3437,
         P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321,
         P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314,
         P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307,
         P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300,
         P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, P2_U3457, P2_U3460,
         P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481,
         P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, P2_U3499, P2_U3502,
         P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512,
         P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519,
         P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526,
         P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, P2_U3532, P2_U3533,
         P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540,
         P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547,
         P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, P2_U3295, P2_U3294,
         P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287,
         P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280,
         P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273,
         P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266,
         P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259,
         P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252,
         P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245,
         P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558,
         P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, P2_U3564, P2_U3565,
         P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, P2_U3571, P2_U3572,
         P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, P2_U3578, P2_U3579,
         P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, P2_U3243, P2_U3242,
         P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235,
         P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228,
         P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221,
         P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3152,
         P2_U3151, P2_U3966;
  wire   n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864,
         n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874,
         n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884,
         n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894,
         n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904,
         n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914,
         n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924,
         n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934,
         n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944,
         n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954,
         n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964,
         n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974,
         n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984,
         n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994,
         n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004,
         n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014,
         n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024,
         n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034,
         n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044,
         n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054,
         n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064,
         n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074,
         n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084,
         n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094,
         n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104,
         n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114,
         n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124,
         n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134,
         n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144,
         n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154,
         n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164,
         n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174,
         n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184,
         n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194,
         n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204,
         n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214,
         n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224,
         n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234,
         n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244,
         n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254,
         n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264,
         n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274,
         n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284,
         n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294,
         n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304,
         n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314,
         n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324,
         n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334,
         n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344,
         n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354,
         n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364,
         n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374,
         n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384,
         n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394,
         n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404,
         n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414,
         n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424,
         n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434,
         n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444,
         n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454,
         n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464,
         n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474,
         n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484,
         n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494,
         n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504,
         n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514,
         n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524,
         n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534,
         n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544,
         n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554,
         n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564,
         n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574,
         n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584,
         n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594,
         n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604,
         n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614,
         n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624,
         n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634,
         n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644,
         n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654,
         n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664,
         n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674,
         n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684,
         n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694,
         n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704,
         n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714,
         n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724,
         n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734,
         n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744,
         n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754,
         n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764,
         n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774,
         n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784,
         n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794,
         n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804,
         n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814,
         n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824,
         n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834,
         n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844,
         n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854,
         n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864,
         n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874,
         n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884,
         n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894,
         n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904,
         n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914,
         n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924,
         n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934,
         n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944,
         n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954,
         n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964,
         n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974,
         n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984,
         n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994,
         n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004,
         n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014,
         n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024,
         n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034,
         n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044,
         n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054,
         n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064,
         n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074,
         n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084,
         n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094,
         n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104,
         n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114,
         n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124,
         n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134,
         n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144,
         n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154,
         n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164,
         n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174,
         n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184,
         n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194,
         n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204,
         n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214,
         n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224,
         n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234,
         n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244,
         n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254,
         n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264,
         n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274,
         n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284,
         n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294,
         n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304,
         n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314,
         n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324,
         n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334,
         n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344,
         n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354,
         n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364,
         n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374,
         n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384,
         n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394,
         n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404,
         n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414,
         n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424,
         n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434,
         n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444,
         n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454,
         n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464,
         n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474,
         n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484,
         n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494,
         n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504,
         n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514,
         n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524,
         n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534,
         n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544,
         n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554,
         n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564,
         n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574,
         n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584,
         n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594,
         n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604,
         n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614,
         n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624,
         n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634,
         n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644,
         n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654,
         n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664,
         n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674,
         n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684,
         n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694,
         n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704,
         n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714,
         n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724,
         n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734,
         n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744,
         n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754,
         n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764,
         n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774,
         n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784,
         n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794,
         n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804,
         n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814,
         n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824,
         n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834,
         n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844,
         n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854,
         n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864,
         n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874,
         n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884,
         n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894,
         n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904,
         n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914,
         n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924,
         n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934,
         n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944,
         n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954,
         n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964,
         n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974,
         n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984,
         n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994,
         n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004,
         n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014,
         n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024,
         n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034,
         n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044,
         n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054,
         n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064,
         n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074,
         n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084,
         n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094,
         n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104,
         n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114,
         n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124,
         n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134,
         n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144,
         n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154,
         n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164,
         n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174,
         n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184,
         n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194,
         n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204,
         n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214,
         n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224,
         n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234,
         n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244,
         n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254,
         n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264,
         n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274,
         n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284,
         n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294,
         n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304,
         n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314,
         n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324,
         n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334,
         n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344,
         n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354,
         n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364,
         n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374,
         n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384,
         n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394,
         n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404,
         n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414,
         n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424,
         n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434,
         n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444,
         n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454,
         n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464,
         n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474,
         n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484,
         n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494,
         n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504,
         n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514,
         n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524,
         n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534,
         n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544,
         n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554,
         n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564,
         n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574,
         n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584,
         n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594,
         n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604,
         n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614,
         n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624,
         n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634,
         n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644,
         n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654,
         n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664,
         n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674,
         n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684,
         n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694,
         n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704,
         n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714,
         n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724,
         n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734,
         n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744,
         n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754,
         n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764,
         n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774,
         n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784,
         n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794,
         n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804,
         n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814,
         n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824,
         n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834,
         n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844,
         n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854,
         n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864,
         n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874,
         n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884,
         n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894,
         n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904,
         n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914,
         n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924,
         n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934,
         n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944,
         n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954,
         n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964,
         n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974,
         n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984,
         n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994,
         n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004,
         n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014,
         n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024,
         n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034,
         n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044,
         n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054,
         n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064,
         n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074,
         n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084,
         n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094,
         n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104,
         n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114,
         n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124,
         n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134,
         n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144,
         n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154,
         n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164,
         n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174,
         n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184,
         n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194,
         n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204,
         n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214,
         n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224,
         n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234,
         n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244,
         n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254,
         n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264,
         n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274,
         n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284,
         n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294,
         n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304,
         n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314,
         n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324,
         n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334,
         n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344,
         n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354,
         n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364,
         n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374,
         n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384,
         n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394,
         n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404,
         n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414,
         n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424,
         n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434,
         n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444,
         n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454,
         n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464,
         n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474,
         n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484,
         n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494,
         n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504,
         n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514,
         n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524,
         n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534,
         n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544,
         n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554,
         n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564,
         n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574,
         n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584,
         n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594,
         n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604,
         n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614,
         n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624,
         n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634,
         n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644,
         n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654,
         n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664,
         n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674,
         n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684,
         n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694,
         n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704,
         n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714,
         n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724,
         n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734,
         n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744,
         n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754,
         n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764,
         n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774,
         n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784,
         n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794,
         n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804,
         n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814,
         n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824,
         n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834,
         n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844,
         n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854,
         n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864,
         n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874,
         n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884,
         n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894,
         n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904,
         n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914,
         n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924,
         n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934,
         n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944,
         n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954,
         n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964,
         n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974,
         n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984,
         n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994,
         n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004,
         n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014,
         n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024,
         n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034,
         n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044,
         n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054,
         n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064,
         n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074,
         n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084,
         n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094,
         n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104,
         n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114,
         n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124,
         n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134,
         n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144,
         n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154,
         n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164,
         n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174,
         n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184,
         n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194,
         n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204,
         n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214,
         n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224,
         n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234,
         n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244,
         n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254,
         n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264,
         n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274,
         n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284,
         n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294,
         n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304,
         n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314,
         n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324,
         n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334,
         n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344,
         n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354,
         n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364,
         n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374,
         n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384,
         n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394,
         n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404,
         n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414,
         n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424,
         n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434,
         n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444,
         n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454,
         n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464,
         n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474,
         n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484,
         n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494,
         n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504,
         n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514,
         n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524,
         n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534,
         n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544,
         n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554,
         n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564,
         n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574,
         n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584,
         n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594,
         n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604,
         n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614,
         n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624,
         n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634,
         n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644,
         n9645, n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655,
         n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665,
         n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675,
         n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685,
         n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695,
         n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705,
         n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715,
         n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725,
         n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735,
         n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745,
         n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755,
         n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765,
         n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775,
         n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785,
         n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795,
         n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805,
         n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815,
         n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825,
         n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835,
         n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845,
         n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855,
         n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865,
         n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875,
         n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885,
         n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895,
         n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905,
         n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915,
         n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925,
         n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935,
         n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945,
         n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955,
         n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965,
         n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975,
         n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985,
         n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995,
         n9996, n9997, n9998, n9999, n10000, n10001, n10002, n10003, n10004,
         n10005, n10006, n10007, n10008, n10009, n10010, n10011, n10012,
         n10013, n10014, n10015, n10016, n10017, n10018, n10019, n10020,
         n10021, n10022, n10023, n10024, n10025, n10026, n10027, n10028,
         n10029, n10030, n10031, n10032, n10033, n10034, n10035, n10036,
         n10037, n10038, n10039, n10040, n10041, n10042, n10043, n10044,
         n10045, n10046, n10047, n10048, n10049, n10050, n10051, n10052,
         n10053, n10054, n10055, n10056, n10057, n10058, n10059, n10060,
         n10061, n10062, n10063, n10064, n10065, n10066, n10067, n10068,
         n10069, n10070, n10071, n10072, n10073, n10074, n10075, n10076,
         n10077, n10078, n10079, n10080, n10081, n10082, n10083, n10084,
         n10085, n10086, n10087, n10088, n10089, n10090, n10091, n10092,
         n10093, n10094, n10095, n10096, n10097, n10098, n10099, n10100,
         n10101, n10102, n10103, n10104, n10105, n10106, n10107, n10108,
         n10109, n10110, n10111, n10112, n10113, n10114, n10115, n10116,
         n10117, n10118, n10119, n10120, n10121, n10122, n10123, n10124,
         n10125, n10126, n10127, n10128, n10129, n10130, n10131, n10132,
         n10133, n10134, n10135, n10136, n10137, n10138, n10139, n10140,
         n10141, n10142, n10143, n10144, n10145, n10146, n10147, n10148,
         n10149, n10150, n10151, n10152, n10153, n10154, n10155, n10156,
         n10157, n10158, n10159, n10160, n10161, n10162, n10163, n10164,
         n10165, n10166, n10167, n10168, n10169, n10170, n10171, n10172,
         n10173, n10174, n10175, n10176, n10177, n10178, n10179, n10180,
         n10181, n10182, n10183, n10184, n10185, n10186, n10187, n10188,
         n10189, n10190, n10191, n10192, n10193, n10194, n10195, n10196,
         n10197, n10198, n10199, n10200, n10201, n10202, n10203, n10204,
         n10205, n10206, n10207, n10208, n10209, n10210, n10211, n10212,
         n10213, n10214, n10215, n10216, n10217, n10218, n10219, n10220,
         n10221, n10222, n10223, n10224, n10225, n10226, n10227, n10228,
         n10229, n10230, n10231, n10232, n10233, n10234, n10235, n10236,
         n10237, n10238, n10239, n10240, n10241, n10242, n10243, n10244,
         n10245, n10246, n10247, n10248, n10249, n10250, n10251, n10252,
         n10253, n10254, n10255, n10256, n10257, n10258, n10259, n10260,
         n10261, n10262, n10263, n10264, n10265, n10266, n10267, n10268,
         n10269, n10270, n10271, n10272, n10273, n10274, n10275, n10276,
         n10277, n10278, n10279, n10280, n10281, n10282, n10283, n10284,
         n10285, n10286, n10287, n10288, n10289, n10290, n10291, n10292,
         n10293, n10294, n10295, n10296, n10297, n10298, n10299, n10300,
         n10301, n10302, n10303, n10304, n10305, n10306, n10307, n10308,
         n10309, n10310, n10311, n10312, n10313, n10314, n10315, n10316,
         n10317, n10318, n10319, n10320, n10321, n10322, n10323, n10324,
         n10325, n10326, n10327, n10328, n10329, n10330, n10331, n10332,
         n10333, n10334, n10335, n10336, n10337, n10338, n10339, n10340,
         n10341, n10342, n10343, n10344, n10345, n10346, n10347, n10348,
         n10349, n10350, n10351, n10352, n10353, n10354, n10355, n10356,
         n10357, n10358, n10359, n10360, n10361, n10362, n10363, n10364,
         n10365, n10366, n10367, n10368, n10369, n10370, n10371, n10372,
         n10373, n10374, n10375, n10376, n10377, n10378, n10379, n10380,
         n10381, n10382, n10383, n10384, n10385, n10386, n10387, n10388,
         n10389, n10390, n10391, n10392, n10393, n10394, n10395, n10396,
         n10397, n10398, n10399, n10400, n10401, n10402, n10403, n10404,
         n10405, n10406, n10407, n10408, n10409, n10410, n10411, n10412,
         n10413, n10414, n10415, n10416, n10417, n10418, n10419, n10420,
         n10421, n10422, n10423, n10424, n10425, n10426, n10427, n10428,
         n10429, n10430, n10431, n10432, n10433, n10434, n10435, n10436,
         n10437, n10438, n10439, n10440, n10441, n10442, n10443, n10444,
         n10445, n10446, n10447, n10448, n10449, n10450, n10451, n10452,
         n10453, n10454, n10455, n10456, n10457, n10458, n10459, n10460,
         n10461, n10462, n10463, n10464, n10465, n10466, n10467, n10468,
         n10469, n10470, n10471, n10472, n10473, n10474, n10475, n10476,
         n10477, n10478, n10479, n10480, n10481, n10482, n10483, n10484,
         n10485, n10486, n10487, n10488, n10489, n10490, n10491, n10492,
         n10493, n10494, n10495, n10496, n10497, n10498, n10499, n10500,
         n10501, n10502, n10503, n10504, n10505, n10506, n10507, n10508,
         n10509, n10510, n10511, n10512, n10513, n10514, n10515, n10516,
         n10517, n10518, n10519, n10520, n10521, n10522, n10523, n10524,
         n10525, n10526, n10527, n10528, n10529, n10530, n10531, n10532,
         n10533, n10534, n10535, n10536, n10537, n10538, n10539, n10540,
         n10541, n10542, n10543, n10544, n10545, n10546, n10547, n10548,
         n10549, n10550, n10551, n10552, n10553, n10554, n10555, n10556,
         n10557, n10558, n10559, n10560, n10561, n10562, n10563, n10564,
         n10565, n10566, n10567, n10568, n10569, n10570, n10571, n10572,
         n10573, n10574, n10575, n10576, n10577, n10578, n10579, n10580,
         n10581, n10582, n10583, n10584, n10585, n10586, n10587, n10588,
         n10589, n10590, n10591, n10592, n10593, n10594, n10595, n10596,
         n10597, n10598, n10599, n10600, n10601, n10602, n10603, n10604,
         n10605, n10606, n10607, n10608, n10609, n10610, n10611, n10612,
         n10613, n10614, n10615, n10616, n10617, n10618, n10619, n10620,
         n10621, n10622, n10623, n10624, n10625, n10626, n10627, n10628,
         n10629, n10630, n10631, n10632, n10633, n10634, n10635, n10636,
         n10637, n10638, n10639, n10640, n10641, n10642, n10643, n10644,
         n10645, n10646;

  INV_X2 U4920 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3152) );
  INV_X1 U4921 ( .A(n8931), .ZN(n8933) );
  INV_X1 U4922 ( .A(n8932), .ZN(n5116) );
  INV_X2 U4924 ( .A(n5474), .ZN(n5975) );
  OAI21_X1 U4925 ( .B1(n8696), .B2(n4945), .A(n4942), .ZN(n8705) );
  OR3_X1 U4926 ( .A1(n8819), .A2(n6510), .A3(n9300), .ZN(n8749) );
  INV_X1 U4927 ( .A(n6305), .ZN(n8212) );
  INV_X1 U4928 ( .A(n6564), .ZN(n8727) );
  NOR2_X2 U4929 ( .A1(n10004), .A2(n10189), .ZN(n9963) );
  NAND2_X1 U4930 ( .A1(n6509), .A2(n9300), .ZN(n8825) );
  INV_X1 U4931 ( .A(n7247), .ZN(n6519) );
  NOR2_X1 U4933 ( .A1(n8251), .A2(n7084), .ZN(n4874) );
  OAI211_X1 U4934 ( .C1(n6683), .C2(n6567), .A(n6566), .B(n6565), .ZN(n10529)
         );
  NAND2_X1 U4935 ( .A1(n5888), .A2(n5887), .ZN(n6322) );
  XNOR2_X1 U4936 ( .A(n5841), .B(P1_IR_REG_22__SCAN_IN), .ZN(n8497) );
  AOI21_X1 U4937 ( .B1(n8525), .B2(n6282), .A(n8518), .ZN(n10176) );
  OAI21_X2 U4938 ( .B1(n8851), .B2(n8850), .A(n8849), .ZN(n8977) );
  AOI21_X2 U4939 ( .B1(n10434), .B2(P1_REG2_REG_9__SCAN_IN), .A(n10438), .ZN(
        n9933) );
  NOR2_X2 U4940 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5442) );
  OAI222_X1 U4941 ( .A1(P2_U3152), .A2(n6509), .B1(n8039), .B2(n6411), .C1(
        n8001), .C2(n8230), .ZN(P2_U3338) );
  NAND2_X4 U4942 ( .A1(n7212), .A2(n6511), .ZN(n8931) );
  AOI21_X2 U4943 ( .B1(n7106), .B2(P2_REG2_REG_9__SCAN_IN), .A(n6758), .ZN(
        n6748) );
  AOI21_X2 U4944 ( .B1(n10123), .B2(n10119), .A(n8388), .ZN(n10035) );
  AOI21_X2 U4945 ( .B1(n6063), .B2(P1_REG2_REG_16__SCAN_IN), .A(n7474), .ZN(
        n7756) );
  AOI21_X2 U4946 ( .B1(n9935), .B2(P1_REG2_REG_10__SCAN_IN), .A(n9931), .ZN(
        n8082) );
  INV_X1 U4947 ( .A(n9740), .ZN(n6621) );
  INV_X2 U4948 ( .A(n6585), .ZN(n8145) );
  INV_X1 U4949 ( .A(n8055), .ZN(n6879) );
  NAND4_X1 U4950 ( .A1(n5491), .A2(n5490), .A3(n5489), .A4(n5488), .ZN(n9881)
         );
  INV_X4 U4951 ( .A(n8208), .ZN(n6216) );
  NAND2_X2 U4952 ( .A1(n6322), .A2(n6281), .ZN(n8208) );
  CLKBUF_X2 U4953 ( .A(n5455), .Z(n5487) );
  INV_X1 U4954 ( .A(n8497), .ZN(n5945) );
  NAND2_X1 U4955 ( .A1(n5845), .A2(n5844), .ZN(n8440) );
  INV_X1 U4956 ( .A(n8329), .ZN(n8486) );
  AOI21_X1 U4957 ( .B1(n8331), .B2(n8330), .A(n8486), .ZN(n8448) );
  AOI211_X1 U4958 ( .C1(n10097), .C2(n10174), .A(n8528), .B(n8527), .ZN(n8529)
         );
  NAND2_X1 U4959 ( .A1(n9812), .A2(n9813), .ZN(n9811) );
  INV_X1 U4960 ( .A(n8525), .ZN(n10177) );
  XNOR2_X1 U4961 ( .A(n5944), .B(n8361), .ZN(n10172) );
  OAI21_X1 U4962 ( .B1(n8508), .B2(n10240), .A(n4975), .ZN(n4974) );
  AND2_X1 U4963 ( .A1(n8512), .A2(n8511), .ZN(n8525) );
  XNOR2_X1 U4964 ( .A(n4977), .B(n5082), .ZN(n8508) );
  NAND2_X1 U4965 ( .A1(n9803), .A2(n9804), .ZN(n9802) );
  AOI21_X1 U4966 ( .B1(n7855), .B2(P2_REG2_REG_16__SCAN_IN), .A(n7832), .ZN(
        n7835) );
  AOI21_X1 U4967 ( .B1(n5903), .B2(n5246), .A(n5902), .ZN(n6920) );
  NAND2_X1 U4968 ( .A1(n6314), .A2(n6313), .ZN(n6592) );
  NAND2_X1 U4969 ( .A1(n5504), .A2(n8461), .ZN(n6901) );
  NAND2_X1 U4970 ( .A1(n5583), .A2(n5582), .ZN(n7287) );
  AND2_X1 U4971 ( .A1(n5518), .A2(n5517), .ZN(n10574) );
  AND2_X2 U4972 ( .A1(n5950), .A2(n10145), .ZN(n10088) );
  INV_X1 U4973 ( .A(n10549), .ZN(n6890) );
  XNOR2_X1 U4974 ( .A(n6283), .B(n8145), .ZN(n6299) );
  NAND2_X1 U4975 ( .A1(n5543), .A2(n5542), .ZN(n5578) );
  AND3_X1 U4976 ( .A1(n5501), .A2(n5500), .A3(n5499), .ZN(n10549) );
  INV_X1 U4977 ( .A(n8057), .ZN(n10519) );
  OAI211_X1 U4978 ( .C1(n5474), .C2(n6527), .A(n5484), .B(n5483), .ZN(n9740)
         );
  NAND2_X2 U4979 ( .A1(n6408), .A2(n6338), .ZN(n9300) );
  AND2_X1 U4980 ( .A1(n5462), .A2(n5461), .ZN(n6303) );
  AND4_X1 U4981 ( .A1(n6539), .A2(n6538), .A3(n6537), .A4(n6536), .ZN(n9321)
         );
  AND2_X2 U4982 ( .A1(n5471), .A2(n6550), .ZN(n5775) );
  OR2_X2 U4983 ( .A1(n6627), .A2(n6211), .ZN(n6305) );
  OAI21_X1 U4984 ( .B1(n4960), .B2(n4961), .A(n5260), .ZN(n5493) );
  INV_X1 U4985 ( .A(n6562), .ZN(n7997) );
  AND2_X2 U4986 ( .A1(n8040), .A2(n8038), .ZN(n6554) );
  INV_X1 U4987 ( .A(n5456), .ZN(n5485) );
  XNOR2_X1 U4988 ( .A(n5869), .B(P1_IR_REG_26__SCAN_IN), .ZN(n5887) );
  NAND2_X1 U4989 ( .A1(n9706), .A2(n6377), .ZN(n8038) );
  AND2_X2 U4990 ( .A1(n10323), .A2(n8025), .ZN(n5476) );
  OR2_X1 U4991 ( .A1(n8440), .A2(n8329), .ZN(n6212) );
  INV_X1 U4992 ( .A(n6210), .ZN(n8491) );
  INV_X1 U4993 ( .A(n5368), .ZN(n8025) );
  XNOR2_X1 U4994 ( .A(n5365), .B(n5364), .ZN(n5369) );
  AND2_X1 U4995 ( .A1(n5344), .A2(n5346), .ZN(n5339) );
  NAND2_X1 U4996 ( .A1(n5363), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5367) );
  OR2_X1 U4997 ( .A1(n6372), .A2(n6162), .ZN(n6233) );
  AND2_X1 U4998 ( .A1(n6232), .A2(n6231), .ZN(n6372) );
  XNOR2_X1 U4999 ( .A(n5415), .B(n5414), .ZN(n9951) );
  NAND2_X2 U5000 ( .A1(n6483), .A2(P1_U3084), .ZN(n6276) );
  AND2_X1 U5001 ( .A1(n5250), .A2(n5249), .ZN(n5251) );
  INV_X2 U5002 ( .A(n6550), .ZN(n6110) );
  INV_X2 U5003 ( .A(n6550), .ZN(n6483) );
  INV_X1 U5004 ( .A(n6124), .ZN(n5186) );
  INV_X2 U5005 ( .A(n5270), .ZN(n6550) );
  NAND2_X2 U5006 ( .A1(n4919), .A2(n4917), .ZN(n5270) );
  BUF_X1 U5007 ( .A(n10478), .Z(n4856) );
  AND4_X1 U5008 ( .A1(n5331), .A2(n5330), .A3(n5329), .A4(n5328), .ZN(n5336)
         );
  AND4_X1 U5009 ( .A1(n5334), .A2(n5333), .A3(n5332), .A4(n5512), .ZN(n5335)
         );
  NOR2_X1 U5010 ( .A1(P1_IR_REG_11__SCAN_IN), .A2(P1_IR_REG_7__SCAN_IN), .ZN(
        n5329) );
  NOR2_X1 U5011 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_4__SCAN_IN), .ZN(
        n5328) );
  NOR2_X1 U5012 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(P1_IR_REG_6__SCAN_IN), .ZN(
        n5330) );
  NOR2_X1 U5013 ( .A1(P1_IR_REG_14__SCAN_IN), .A2(P1_IR_REG_18__SCAN_IN), .ZN(
        n5333) );
  NOR2_X1 U5014 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(P1_IR_REG_21__SCAN_IN), .ZN(
        n5338) );
  NOR2_X1 U5015 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(P1_IR_REG_15__SCAN_IN), .ZN(
        n5332) );
  NOR2_X1 U5016 ( .A1(P1_IR_REG_2__SCAN_IN), .A2(P1_IR_REG_3__SCAN_IN), .ZN(
        n5327) );
  INV_X1 U5017 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n5512) );
  NOR2_X2 U5018 ( .A1(n6217), .A2(n6348), .ZN(n6344) );
  CLKBUF_X1 U5019 ( .A(n5851), .Z(n4855) );
  OAI211_X1 U5020 ( .C1(n5487), .C2(P1_REG3_REG_3__SCAN_IN), .A(n4893), .B(
        n5480), .ZN(n8055) );
  XNOR2_X1 U5021 ( .A(n6111), .B(P2_IR_REG_1__SCAN_IN), .ZN(n10478) );
  AOI21_X2 U5022 ( .B1(n7759), .B2(P1_REG2_REG_17__SCAN_IN), .A(n7754), .ZN(
        n6059) );
  NAND2_X2 U5023 ( .A1(n6683), .A2(n6483), .ZN(n6562) );
  AND2_X1 U5024 ( .A1(n5471), .A2(n6550), .ZN(n4857) );
  AND2_X1 U5025 ( .A1(n5471), .A2(n6550), .ZN(n4858) );
  NAND2_X1 U5026 ( .A1(n4978), .A2(n5923), .ZN(n5925) );
  INV_X1 U5027 ( .A(n10067), .ZN(n4978) );
  OAI21_X1 U5028 ( .B1(n8753), .B2(n8752), .A(n8751), .ZN(n8794) );
  AOI21_X1 U5029 ( .B1(n4948), .B2(n4868), .A(n4947), .ZN(n8752) );
  NAND2_X1 U5030 ( .A1(n5140), .A2(n5619), .ZN(n4971) );
  NOR2_X2 U5031 ( .A1(n9164), .A2(n9374), .ZN(n9137) );
  NAND2_X1 U5032 ( .A1(n6683), .A2(n6550), .ZN(n6564) );
  NAND2_X2 U5033 ( .A1(n6492), .A2(n8824), .ZN(n6683) );
  NOR2_X1 U5034 ( .A1(n5221), .A2(P1_IR_REG_23__SCAN_IN), .ZN(n5005) );
  OR2_X1 U5035 ( .A1(n8606), .A2(n8605), .ZN(n8619) );
  OR2_X1 U5036 ( .A1(n5149), .A2(n5148), .ZN(n4950) );
  OR2_X1 U5037 ( .A1(n8714), .A2(n8746), .ZN(n5148) );
  AOI21_X1 U5038 ( .B1(n5151), .B2(n8757), .A(n5150), .ZN(n5149) );
  OR2_X1 U5039 ( .A1(n9379), .A2(n9185), .ZN(n8808) );
  OR2_X1 U5040 ( .A1(n9426), .A2(n8837), .ZN(n8656) );
  OR2_X1 U5041 ( .A1(n9437), .A2(n7970), .ZN(n8576) );
  XNOR2_X1 U5042 ( .A(n9432), .B(n9003), .ZN(n9294) );
  NAND2_X1 U5043 ( .A1(n6008), .A2(n5189), .ZN(n5188) );
  INV_X1 U5044 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n5189) );
  NAND2_X1 U5045 ( .A1(n6118), .A2(n6007), .ZN(n6124) );
  AND2_X1 U5046 ( .A1(n6587), .A2(n6588), .ZN(n6593) );
  XOR2_X1 U5047 ( .A(n6586), .B(n8195), .Z(n6595) );
  OAI22_X1 U5048 ( .A1(n6904), .A2(n8208), .B1(n6664), .B2(n6627), .ZN(n6586)
         );
  AND2_X1 U5049 ( .A1(n8326), .A2(n9867), .ZN(n8483) );
  NAND2_X1 U5050 ( .A1(n5073), .A2(n5077), .ZN(n8510) );
  INV_X1 U5051 ( .A(n5078), .ZN(n5077) );
  OAI22_X1 U5052 ( .A1(n8473), .A2(n5079), .B1(n9722), .B2(n9871), .ZN(n5078)
         );
  OR2_X1 U5053 ( .A1(n9722), .A2(n9971), .ZN(n8429) );
  OR2_X1 U5054 ( .A1(n10189), .A2(n10001), .ZN(n8426) );
  NAND2_X1 U5055 ( .A1(n5925), .A2(n4887), .ZN(n5929) );
  NOR2_X1 U5056 ( .A1(n4982), .A2(n4981), .ZN(n4980) );
  NAND2_X1 U5057 ( .A1(n5092), .A2(n10057), .ZN(n4981) );
  NOR2_X1 U5058 ( .A1(n10158), .A2(n5090), .ZN(n4982) );
  NAND2_X1 U5059 ( .A1(n4864), .A2(n8239), .ZN(n5092) );
  NAND2_X1 U5060 ( .A1(n4897), .A2(n5864), .ZN(n5112) );
  OAI21_X1 U5061 ( .B1(n5376), .B2(n4902), .A(n5152), .ZN(n5756) );
  AOI21_X1 U5062 ( .B1(n5737), .B2(n5153), .A(n4907), .ZN(n5152) );
  OAI21_X1 U5063 ( .B1(n5412), .B2(n5411), .A(n5316), .ZN(n5398) );
  XNOR2_X1 U5064 ( .A(n5307), .B(SI_16_), .ZN(n5686) );
  XNOR2_X1 U5065 ( .A(n5298), .B(SI_13_), .ZN(n5638) );
  AND2_X1 U5066 ( .A1(n5283), .A2(n5540), .ZN(n5282) );
  INV_X1 U5067 ( .A(n6509), .ZN(n8762) );
  AND2_X1 U5068 ( .A1(n6980), .A2(n8819), .ZN(n8755) );
  OAI211_X1 U5069 ( .C1(n8822), .C2(n8823), .A(n4865), .B(n4931), .ZN(n4930)
         );
  NAND2_X1 U5070 ( .A1(n8820), .A2(n8819), .ZN(n4931) );
  AND2_X1 U5071 ( .A1(n6510), .A2(n8813), .ZN(n6499) );
  NAND2_X1 U5072 ( .A1(n8536), .A2(n8535), .ZN(n9106) );
  AND2_X1 U5073 ( .A1(n8741), .A2(n8740), .ZN(n9173) );
  OR2_X1 U5074 ( .A1(n9391), .A2(n9219), .ZN(n9181) );
  NAND2_X1 U5075 ( .A1(n9123), .A2(n9219), .ZN(n5049) );
  OR2_X1 U5076 ( .A1(n8566), .A2(n9469), .ZN(n6607) );
  AOI21_X1 U5077 ( .B1(n7662), .B2(n7661), .A(n7660), .ZN(n7915) );
  NOR2_X1 U5078 ( .A1(n9032), .A2(n10633), .ZN(n7660) );
  INV_X1 U5079 ( .A(n6683), .ZN(n7996) );
  NAND2_X1 U5080 ( .A1(n8731), .A2(n8730), .ZN(n9374) );
  INV_X1 U5081 ( .A(n6226), .ZN(n6017) );
  NAND2_X1 U5082 ( .A1(n8497), .A2(n8453), .ZN(n6003) );
  OAI21_X1 U5083 ( .B1(n8053), .B2(n8054), .A(n6308), .ZN(n9737) );
  OR2_X1 U5084 ( .A1(n5728), .A2(n5418), .ZN(n5420) );
  NAND2_X1 U5085 ( .A1(n9857), .A2(n5210), .ZN(n5208) );
  NAND2_X1 U5086 ( .A1(n9811), .A2(n5211), .ZN(n5209) );
  AND2_X1 U5087 ( .A1(n9857), .A2(n5212), .ZN(n5211) );
  INV_X1 U5088 ( .A(n5478), .ZN(n5830) );
  INV_X1 U5089 ( .A(n5476), .ZN(n5421) );
  NAND2_X1 U5090 ( .A1(n10323), .A2(n5368), .ZN(n5455) );
  NAND2_X1 U5091 ( .A1(n5994), .A2(n5071), .ZN(n8514) );
  NOR2_X1 U5092 ( .A1(n5910), .A2(n5088), .ZN(n5087) );
  NAND2_X1 U5093 ( .A1(n5342), .A2(n5341), .ZN(n5343) );
  INV_X1 U5094 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n5346) );
  NAND2_X1 U5095 ( .A1(n5162), .A2(n5160), .ZN(n5702) );
  NAND2_X1 U5096 ( .A1(n5654), .A2(n5301), .ZN(n5658) );
  AND2_X1 U5097 ( .A1(n5300), .A2(n5653), .ZN(n5301) );
  AND2_X1 U5098 ( .A1(n4971), .A2(n4970), .ZN(n5622) );
  INV_X1 U5099 ( .A(n5257), .ZN(n5167) );
  INV_X2 U5100 ( .A(n5471), .ZN(n10408) );
  MUX2_X1 U5101 ( .A(n8595), .B(n8594), .S(n8749), .Z(n8596) );
  MUX2_X1 U5102 ( .A(n8623), .B(n8622), .S(n8749), .Z(n8626) );
  INV_X1 U5103 ( .A(n4941), .ZN(n4938) );
  AOI21_X1 U5104 ( .B1(n4946), .B2(n4944), .A(n4943), .ZN(n4942) );
  INV_X1 U5105 ( .A(n4946), .ZN(n4945) );
  INV_X1 U5106 ( .A(n9181), .ZN(n4943) );
  NAND2_X1 U5107 ( .A1(n5159), .A2(n5156), .ZN(n8694) );
  NAND2_X1 U5108 ( .A1(n8804), .A2(n4881), .ZN(n5159) );
  NAND2_X1 U5109 ( .A1(n8758), .A2(n5157), .ZN(n5156) );
  OAI21_X1 U5110 ( .B1(n5151), .B2(n4894), .A(n5147), .ZN(n5146) );
  NAND2_X1 U5111 ( .A1(n7908), .A2(n9294), .ZN(n7916) );
  OR2_X1 U5112 ( .A1(n7587), .A2(n7767), .ZN(n8608) );
  AND2_X1 U5113 ( .A1(n5186), .A2(n5187), .ZN(n6010) );
  INV_X1 U5114 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n6008) );
  INV_X1 U5115 ( .A(n7133), .ZN(n5206) );
  OR2_X1 U5116 ( .A1(n6835), .A2(n5206), .ZN(n5205) );
  INV_X1 U5117 ( .A(n7335), .ZN(n5203) );
  OR2_X1 U5118 ( .A1(n5083), .A2(n5080), .ZN(n5079) );
  INV_X1 U5119 ( .A(n5941), .ZN(n5080) );
  NAND2_X1 U5120 ( .A1(n6923), .A2(n6915), .ZN(n8369) );
  OR2_X1 U5121 ( .A1(n5273), .A2(n5272), .ZN(n5279) );
  INV_X1 U5122 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n4929) );
  INV_X1 U5123 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n4921) );
  INV_X1 U5124 ( .A(P1_RD_REG_SCAN_IN), .ZN(n4920) );
  NAND2_X1 U5125 ( .A1(n5116), .A2(n9040), .ZN(n6531) );
  OAI211_X1 U5126 ( .C1(n5181), .C2(n8818), .A(n5178), .B(n8817), .ZN(n8821)
         );
  OAI211_X1 U5127 ( .C1(n5180), .C2(n9130), .A(n8791), .B(n5179), .ZN(n5178)
         );
  INV_X1 U5128 ( .A(n8038), .ZN(n5168) );
  NOR2_X1 U5129 ( .A1(n5043), .A2(n8807), .ZN(n5042) );
  NOR2_X1 U5130 ( .A1(n5045), .A2(n8807), .ZN(n5041) );
  NAND2_X1 U5131 ( .A1(n9394), .A2(n9206), .ZN(n8758) );
  OR2_X1 U5132 ( .A1(n9394), .A2(n9206), .ZN(n8804) );
  AND2_X1 U5133 ( .A1(n8800), .A2(n5174), .ZN(n5173) );
  NAND2_X1 U5134 ( .A1(n5175), .A2(n8574), .ZN(n5174) );
  INV_X1 U5135 ( .A(n8575), .ZN(n5175) );
  INV_X1 U5136 ( .A(n8574), .ZN(n5176) );
  NOR2_X1 U5137 ( .A1(n9278), .A2(n5064), .ZN(n5061) );
  NOR2_X1 U5138 ( .A1(n7897), .A2(n5196), .ZN(n5195) );
  INV_X1 U5139 ( .A(n8630), .ZN(n5196) );
  NOR2_X1 U5140 ( .A1(n7897), .A2(n5193), .ZN(n5192) );
  NAND2_X1 U5141 ( .A1(n8630), .A2(n8629), .ZN(n5193) );
  NAND2_X1 U5142 ( .A1(n6393), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n7715) );
  OR2_X1 U5143 ( .A1(n7424), .A2(n9556), .ZN(n7626) );
  NOR3_X1 U5144 ( .A1(n7568), .A2(n5033), .A3(n7225), .ZN(n5032) );
  INV_X1 U5145 ( .A(n7387), .ZN(n5033) );
  AND2_X1 U5146 ( .A1(n8608), .A2(n8617), .ZN(n8770) );
  NOR2_X1 U5147 ( .A1(n7386), .A2(n6979), .ZN(n4984) );
  NOR2_X1 U5148 ( .A1(n9039), .A2(n6519), .ZN(n8593) );
  INV_X1 U5149 ( .A(n10529), .ZN(n6959) );
  NAND2_X1 U5150 ( .A1(n7257), .A2(n8761), .ZN(n7256) );
  NAND2_X1 U5151 ( .A1(n7259), .A2(n10529), .ZN(n8584) );
  AOI21_X1 U5152 ( .B1(n7941), .B2(n8576), .A(n7940), .ZN(n9295) );
  NOR2_X1 U5153 ( .A1(n6460), .A2(n7585), .ZN(n6471) );
  AND2_X1 U5154 ( .A1(n7360), .A2(n6459), .ZN(n6460) );
  AND2_X1 U5155 ( .A1(n6006), .A2(n6005), .ZN(n6118) );
  NOR2_X1 U5156 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_2__SCAN_IN), .ZN(
        n6006) );
  NOR2_X1 U5157 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_3__SCAN_IN), .ZN(
        n6005) );
  NAND2_X1 U5158 ( .A1(n5216), .A2(n9831), .ZN(n5215) );
  NOR2_X1 U5159 ( .A1(n5217), .A2(n5011), .ZN(n5010) );
  INV_X1 U5160 ( .A(n9831), .ZN(n5217) );
  NAND2_X1 U5161 ( .A1(n5010), .A2(n8148), .ZN(n5007) );
  XNOR2_X1 U5162 ( .A(n6309), .B(n8145), .ZN(n6310) );
  OR2_X1 U5163 ( .A1(n9757), .A2(n5012), .ZN(n5011) );
  INV_X1 U5164 ( .A(n8151), .ZN(n5012) );
  NAND2_X1 U5165 ( .A1(n6322), .A2(n6212), .ZN(n6627) );
  AOI21_X1 U5166 ( .B1(n8437), .B2(n8436), .A(n8435), .ZN(n8449) );
  INV_X1 U5167 ( .A(n8440), .ZN(n8453) );
  NAND2_X1 U5168 ( .A1(n5836), .A2(n9869), .ZN(n8314) );
  NOR2_X1 U5169 ( .A1(n8509), .A2(n5082), .ZN(n5068) );
  OR2_X1 U5170 ( .A1(n10075), .A2(n8155), .ZN(n5922) );
  NOR2_X1 U5171 ( .A1(n10155), .A2(n10237), .ZN(n5024) );
  OR2_X1 U5172 ( .A1(n10237), .A2(n8110), .ZN(n8416) );
  OR2_X1 U5173 ( .A1(n7809), .A2(n7878), .ZN(n8414) );
  OR2_X1 U5174 ( .A1(n10263), .A2(n7603), .ZN(n8404) );
  NOR2_X1 U5175 ( .A1(n10047), .A2(n10197), .ZN(n10017) );
  NOR2_X1 U5176 ( .A1(n6896), .A2(n5901), .ZN(n5902) );
  OR2_X1 U5177 ( .A1(n5960), .A2(n5959), .ZN(n5965) );
  XNOR2_X1 U5178 ( .A(n5960), .B(n5959), .ZN(n5958) );
  OR2_X1 U5179 ( .A1(n5810), .A2(n5809), .ZN(n5812) );
  OAI21_X1 U5180 ( .B1(n5756), .B2(n5755), .A(n5754), .ZN(n5774) );
  AOI21_X1 U5181 ( .B1(n5398), .B2(n5397), .A(n5318), .ZN(n5385) );
  OAI21_X1 U5182 ( .B1(n5674), .B2(n4967), .A(n4912), .ZN(n5412) );
  NOR2_X1 U5183 ( .A1(n4886), .A2(n4913), .ZN(n4912) );
  INV_X1 U5184 ( .A(n4964), .ZN(n4913) );
  NOR2_X1 U5185 ( .A1(n5700), .A2(n5161), .ZN(n5160) );
  INV_X1 U5186 ( .A(n5163), .ZN(n5161) );
  NOR2_X1 U5187 ( .A1(n5686), .A2(n5166), .ZN(n5165) );
  INV_X1 U5188 ( .A(n5306), .ZN(n5166) );
  OAI21_X1 U5189 ( .B1(n5270), .B2(n4956), .A(n4955), .ZN(n4954) );
  NAND2_X1 U5190 ( .A1(n5270), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n4955) );
  INV_X1 U5191 ( .A(n5465), .ZN(n5254) );
  NAND2_X1 U5192 ( .A1(n5270), .A2(n5248), .ZN(n5249) );
  INV_X1 U5193 ( .A(n4969), .ZN(n5250) );
  OAI21_X1 U5194 ( .B1(n5270), .B2(P1_DATAO_REG_0__SCAN_IN), .A(SI_0_), .ZN(
        n4969) );
  OR3_X1 U5195 ( .A1(n7206), .A2(n7585), .A3(n7360), .ZN(n6229) );
  AND2_X1 U5196 ( .A1(n7706), .A2(n5134), .ZN(n5133) );
  NAND2_X1 U5197 ( .A1(n7618), .A2(n7620), .ZN(n5134) );
  NAND2_X1 U5198 ( .A1(n6391), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n7117) );
  INV_X1 U5199 ( .A(n7048), .ZN(n6391) );
  INV_X1 U5200 ( .A(n8929), .ZN(n5123) );
  NOR2_X1 U5201 ( .A1(n9009), .A2(n5128), .ZN(n5127) );
  INV_X1 U5202 ( .A(n8888), .ZN(n5128) );
  INV_X1 U5203 ( .A(n5125), .ZN(n5124) );
  OAI21_X1 U5204 ( .B1(n9009), .B2(n5126), .A(n8891), .ZN(n5125) );
  NAND2_X1 U5205 ( .A1(n8964), .A2(n8888), .ZN(n5126) );
  OR2_X1 U5206 ( .A1(n6991), .A2(n6990), .ZN(n7048) );
  OR2_X1 U5207 ( .A1(n7305), .A2(n7304), .ZN(n7424) );
  OR2_X1 U5208 ( .A1(n8675), .A2(n9575), .ZN(n8685) );
  NAND2_X1 U5209 ( .A1(n6574), .A2(n5114), .ZN(n6717) );
  INV_X1 U5210 ( .A(n6715), .ZN(n5114) );
  NAND2_X1 U5211 ( .A1(n6568), .A2(n4875), .ZN(n8906) );
  INV_X1 U5212 ( .A(n8531), .ZN(n6568) );
  OR2_X1 U5213 ( .A1(n7117), .A2(n7116), .ZN(n7162) );
  NAND2_X1 U5214 ( .A1(n6392), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n7305) );
  INV_X1 U5215 ( .A(n7162), .ZN(n6392) );
  AND2_X1 U5216 ( .A1(n6488), .A2(n10362), .ZN(n6491) );
  INV_X1 U5217 ( .A(n6499), .ZN(n6981) );
  INV_X1 U5218 ( .A(n6491), .ZN(n6580) );
  OAI21_X1 U5219 ( .B1(n6238), .B2(P2_IR_REG_21__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n6237) );
  NAND2_X1 U5220 ( .A1(n8543), .A2(n8542), .ZN(n9113) );
  NAND2_X1 U5221 ( .A1(n9137), .A2(n9370), .ZN(n9138) );
  AND2_X1 U5222 ( .A1(n8807), .A2(n8806), .ZN(n5184) );
  NAND2_X1 U5223 ( .A1(n9200), .A2(n8805), .ZN(n5185) );
  NAND2_X1 U5224 ( .A1(n9163), .A2(n9169), .ZN(n9164) );
  INV_X1 U5225 ( .A(n5046), .ZN(n5045) );
  OAI21_X1 U5226 ( .B1(n9182), .B2(n5049), .A(n5047), .ZN(n5046) );
  NAND2_X1 U5227 ( .A1(n5048), .A2(n9172), .ZN(n5047) );
  NAND2_X1 U5228 ( .A1(n5044), .A2(n9124), .ZN(n5043) );
  INV_X1 U5229 ( .A(n9182), .ZN(n5044) );
  AND2_X1 U5230 ( .A1(n8726), .A2(n8725), .ZN(n9185) );
  OR2_X1 U5231 ( .A1(n9166), .A2(n7303), .ZN(n8726) );
  AND2_X1 U5232 ( .A1(n8756), .A2(n8806), .ZN(n9182) );
  NAND2_X1 U5233 ( .A1(n9231), .A2(n4915), .ZN(n9221) );
  AND2_X1 U5234 ( .A1(n8803), .A2(n8802), .ZN(n4915) );
  NAND2_X1 U5235 ( .A1(n5058), .A2(n5056), .ZN(n9237) );
  INV_X1 U5236 ( .A(n5057), .ZN(n5056) );
  OAI22_X1 U5237 ( .A1(n9120), .A2(n9119), .B1(n9404), .B2(n9280), .ZN(n5057)
         );
  OR2_X1 U5238 ( .A1(n9404), .A2(n8957), .ZN(n9230) );
  AND2_X1 U5239 ( .A1(n8759), .A2(n8802), .ZN(n9236) );
  NAND2_X1 U5240 ( .A1(n9230), .A2(n8691), .ZN(n9254) );
  NAND2_X1 U5241 ( .A1(n9414), .A2(n5061), .ZN(n5062) );
  OR2_X1 U5242 ( .A1(n6981), .A2(n6707), .ZN(n9318) );
  NAND2_X1 U5243 ( .A1(n10565), .A2(n7032), .ZN(n5055) );
  OAI21_X1 U5244 ( .B1(n7237), .B2(n6964), .A(n6963), .ZN(n7376) );
  INV_X1 U5245 ( .A(n9345), .ZN(n9320) );
  NAND2_X1 U5246 ( .A1(n9042), .A2(n10513), .ZN(n9338) );
  NOR2_X1 U5247 ( .A1(n9370), .A2(n10625), .ZN(n4990) );
  OR2_X1 U5248 ( .A1(n10501), .A2(n8762), .ZN(n10637) );
  INV_X1 U5249 ( .A(n10637), .ZN(n10511) );
  INV_X1 U5250 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n6162) );
  INV_X1 U5251 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n6371) );
  INV_X1 U5252 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n4996) );
  XNOR2_X1 U5253 ( .A(n6239), .B(P2_IR_REG_21__SCAN_IN), .ZN(n8813) );
  NAND2_X1 U5254 ( .A1(n6335), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6337) );
  NAND2_X1 U5255 ( .A1(n6337), .A2(n6336), .ZN(n6408) );
  AND3_X1 U5256 ( .A1(n6174), .A2(n6177), .A3(n6014), .ZN(n6015) );
  AND2_X1 U5257 ( .A1(n6179), .A2(n6195), .ZN(n7738) );
  NAND2_X1 U5258 ( .A1(n9727), .A2(n9726), .ZN(n9725) );
  NAND2_X1 U5259 ( .A1(n5003), .A2(n6314), .ZN(n5002) );
  AND2_X1 U5260 ( .A1(n6313), .A2(n6596), .ZN(n5003) );
  AND2_X1 U5261 ( .A1(n6595), .A2(n6594), .ZN(n6591) );
  OR2_X1 U5262 ( .A1(n5747), .A2(n9816), .ZN(n5760) );
  NAND2_X1 U5263 ( .A1(n5358), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n5403) );
  OR2_X1 U5264 ( .A1(n5403), .A2(n5391), .ZN(n5393) );
  AOI21_X1 U5265 ( .B1(n8328), .B2(n8327), .A(n8483), .ZN(n8330) );
  AND2_X1 U5266 ( .A1(n8486), .A2(n9951), .ZN(n6210) );
  NAND2_X1 U5267 ( .A1(n5485), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n5450) );
  AND2_X1 U5268 ( .A1(n9963), .A2(n5016), .ZN(n9958) );
  NOR2_X1 U5269 ( .A1(n10169), .A2(n5017), .ZN(n5016) );
  INV_X1 U5270 ( .A(n5018), .ZN(n5017) );
  INV_X1 U5271 ( .A(n10169), .ZN(n5836) );
  AOI21_X1 U5272 ( .B1(n8522), .B2(n5446), .A(n5821), .ZN(n9717) );
  AND2_X1 U5273 ( .A1(n5807), .A2(n5806), .ZN(n9971) );
  NAND2_X1 U5274 ( .A1(n9963), .A2(n9969), .ZN(n9964) );
  AND2_X1 U5275 ( .A1(n5767), .A2(n5766), .ZN(n10001) );
  OR2_X1 U5276 ( .A1(n5931), .A2(n5930), .ZN(n5932) );
  NAND2_X1 U5277 ( .A1(n5928), .A2(n4980), .ZN(n5933) );
  NOR3_X1 U5278 ( .A1(n7872), .A2(n5023), .A3(n10109), .ZN(n10108) );
  OR2_X1 U5279 ( .A1(n5094), .A2(n4864), .ZN(n10122) );
  AND2_X1 U5280 ( .A1(n8286), .A2(n8372), .ZN(n10157) );
  NOR2_X1 U5281 ( .A1(n7872), .A2(n10237), .ZN(n10151) );
  AND2_X1 U5282 ( .A1(n8414), .A2(n8376), .ZN(n8352) );
  NAND2_X1 U5283 ( .A1(n7600), .A2(n5915), .ZN(n7689) );
  NAND2_X1 U5284 ( .A1(n5914), .A2(n5085), .ZN(n7600) );
  NOR2_X1 U5285 ( .A1(n8351), .A2(n5086), .ZN(n5085) );
  INV_X1 U5286 ( .A(n5913), .ZN(n5086) );
  NOR2_X1 U5287 ( .A1(n7608), .A2(n10254), .ZN(n7697) );
  NAND2_X1 U5288 ( .A1(n6947), .A2(n5906), .ZN(n7085) );
  OR2_X1 U5289 ( .A1(n5571), .A2(n7147), .ZN(n5586) );
  AND2_X1 U5290 ( .A1(n8400), .A2(n8247), .ZN(n8344) );
  NAND2_X1 U5291 ( .A1(n5539), .A2(n5108), .ZN(n6921) );
  NAND2_X1 U5292 ( .A1(n5350), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n5550) );
  AND4_X1 U5293 ( .A1(n5556), .A2(n5555), .A3(n5554), .A4(n5553), .ZN(n7150)
         );
  INV_X1 U5294 ( .A(n6629), .ZN(n6923) );
  INV_X1 U5295 ( .A(n10141), .ZN(n10103) );
  INV_X1 U5296 ( .A(n10143), .ZN(n10101) );
  INV_X1 U5297 ( .A(n10140), .ZN(n9997) );
  AND2_X1 U5298 ( .A1(n6217), .A2(n6453), .ZN(n6343) );
  NAND2_X1 U5299 ( .A1(n5977), .A2(n5976), .ZN(n8233) );
  NAND2_X1 U5300 ( .A1(n5746), .A2(n5745), .ZN(n10007) );
  NAND2_X1 U5301 ( .A1(n5611), .A2(n5610), .ZN(n10268) );
  OR2_X1 U5302 ( .A1(n6451), .A2(n8329), .ZN(n10591) );
  INV_X1 U5303 ( .A(n10595), .ZN(n10240) );
  NOR2_X1 U5304 ( .A1(n4892), .A2(n5112), .ZN(n5111) );
  OR2_X1 U5305 ( .A1(n5958), .A2(n9597), .ZN(n5971) );
  INV_X1 U5306 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n5364) );
  NAND2_X1 U5307 ( .A1(n5201), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5365) );
  NAND2_X1 U5308 ( .A1(n5863), .A2(n5110), .ZN(n5345) );
  INV_X1 U5309 ( .A(n5112), .ZN(n5110) );
  NAND2_X1 U5310 ( .A1(n5388), .A2(n5323), .ZN(n5376) );
  XNOR2_X1 U5311 ( .A(n5376), .B(n5375), .ZN(n8671) );
  INV_X1 U5312 ( .A(n5309), .ZN(n4968) );
  NAND2_X1 U5313 ( .A1(n5164), .A2(n9619), .ZN(n5163) );
  INV_X1 U5314 ( .A(n5307), .ZN(n5164) );
  NAND2_X1 U5315 ( .A1(n5674), .A2(n5165), .ZN(n5162) );
  XNOR2_X1 U5316 ( .A(n5687), .B(n5686), .ZN(n7854) );
  NAND2_X1 U5317 ( .A1(n5622), .A2(n5295), .ZN(n5639) );
  NAND2_X1 U5318 ( .A1(n4923), .A2(n5141), .ZN(n5140) );
  AOI21_X1 U5319 ( .B1(n5144), .B2(n5143), .A(n5142), .ZN(n5141) );
  INV_X1 U5320 ( .A(n5291), .ZN(n5142) );
  NAND2_X1 U5321 ( .A1(n5285), .A2(n4885), .ZN(n5145) );
  NAND2_X1 U5322 ( .A1(n5255), .A2(n5254), .ZN(n5467) );
  NAND2_X1 U5323 ( .A1(n8665), .A2(n8664), .ZN(n9409) );
  NAND2_X1 U5324 ( .A1(n7418), .A2(n7417), .ZN(n10633) );
  NAND2_X1 U5325 ( .A1(n7925), .A2(n7924), .ZN(n9426) );
  AND2_X1 U5326 ( .A1(n6406), .A2(n6405), .ZN(n9219) );
  XNOR2_X1 U5327 ( .A(n6237), .B(P2_IR_REG_22__SCAN_IN), .ZN(n6510) );
  INV_X1 U5328 ( .A(n4930), .ZN(n4934) );
  NOR2_X1 U5329 ( .A1(n8762), .A2(n8755), .ZN(n5138) );
  INV_X1 U5330 ( .A(n9206), .ZN(n9233) );
  INV_X1 U5331 ( .A(n9300), .ZN(n9103) );
  INV_X1 U5332 ( .A(n9365), .ZN(n9112) );
  NAND2_X1 U5333 ( .A1(n9151), .A2(n9173), .ZN(n9125) );
  NAND2_X1 U5334 ( .A1(n7907), .A2(n7906), .ZN(n9432) );
  OR2_X1 U5335 ( .A1(n7905), .A2(n6564), .ZN(n7907) );
  AND2_X1 U5336 ( .A1(n7206), .A2(n7585), .ZN(n10465) );
  XNOR2_X1 U5337 ( .A(n6235), .B(n6231), .ZN(n8824) );
  NAND2_X1 U5338 ( .A1(n6234), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6235) );
  AND2_X1 U5339 ( .A1(n5208), .A2(n8201), .ZN(n5207) );
  NAND2_X1 U5340 ( .A1(n8200), .A2(n8199), .ZN(n8201) );
  NAND2_X1 U5341 ( .A1(n5798), .A2(n5797), .ZN(n9722) );
  NAND2_X1 U5342 ( .A1(n5663), .A2(n5662), .ZN(n8271) );
  OR2_X1 U5343 ( .A1(n7711), .A2(n5474), .ZN(n5663) );
  NAND2_X1 U5344 ( .A1(n4857), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n5484) );
  AOI21_X1 U5345 ( .B1(n5001), .B2(n5000), .A(n9853), .ZN(n4999) );
  NOR2_X1 U5346 ( .A1(n9857), .A2(n5210), .ZN(n5000) );
  NAND2_X1 U5347 ( .A1(n9811), .A2(n5212), .ZN(n5001) );
  INV_X1 U5348 ( .A(n9783), .ZN(n9858) );
  INV_X1 U5349 ( .A(n9971), .ZN(n9871) );
  AND2_X1 U5350 ( .A1(n6091), .A2(n6090), .ZN(n10443) );
  NAND2_X1 U5351 ( .A1(n5076), .A2(n5941), .ZN(n4977) );
  NAND2_X1 U5352 ( .A1(n5075), .A2(n5083), .ZN(n5076) );
  NAND2_X1 U5353 ( .A1(n5723), .A2(n5722), .ZN(n10133) );
  INV_X1 U5354 ( .A(n8333), .ZN(n10279) );
  NAND2_X1 U5355 ( .A1(n5471), .A2(n5029), .ZN(n5028) );
  OR2_X1 U5356 ( .A1(n5471), .A2(n6114), .ZN(n5445) );
  OAI21_X1 U5357 ( .B1(n6541), .B2(n6550), .A(n5030), .ZN(n5029) );
  NOR2_X1 U5358 ( .A1(n7523), .A2(n7522), .ZN(n10392) );
  NOR2_X1 U5359 ( .A1(n10390), .A2(n10389), .ZN(n7522) );
  NAND2_X1 U5360 ( .A1(n8627), .A2(n4957), .ZN(n8633) );
  AOI21_X1 U5361 ( .B1(n4959), .B2(n8746), .A(n4958), .ZN(n4957) );
  OAI21_X1 U5362 ( .B1(n8626), .B2(n8625), .A(n8624), .ZN(n8627) );
  OAI21_X1 U5363 ( .B1(n4869), .B2(n8746), .A(n8776), .ZN(n4958) );
  AOI21_X1 U5364 ( .B1(n8694), .B2(n8695), .A(n9394), .ZN(n4946) );
  INV_X1 U5365 ( .A(n8694), .ZN(n4944) );
  NOR2_X1 U5366 ( .A1(n5158), .A2(n8746), .ZN(n5157) );
  INV_X1 U5367 ( .A(n8802), .ZN(n5158) );
  NAND2_X1 U5368 ( .A1(n4938), .A2(n8666), .ZN(n4937) );
  NAND2_X1 U5369 ( .A1(n4940), .A2(n8666), .ZN(n4936) );
  OAI21_X1 U5370 ( .B1(n8696), .B2(n8695), .A(n8694), .ZN(n8697) );
  INV_X1 U5371 ( .A(n8805), .ZN(n5150) );
  NOR2_X1 U5372 ( .A1(n8713), .A2(n8749), .ZN(n5147) );
  AND2_X1 U5373 ( .A1(n8233), .A2(n8232), .ZN(n8318) );
  NOR2_X1 U5374 ( .A1(n5183), .A2(n8811), .ZN(n5182) );
  NOR2_X1 U5375 ( .A1(n5081), .A2(n9987), .ZN(n5074) );
  NAND2_X1 U5376 ( .A1(n5082), .A2(n5941), .ZN(n5081) );
  OR2_X1 U5377 ( .A1(n10157), .A2(n5091), .ZN(n5090) );
  INV_X1 U5378 ( .A(n8239), .ZN(n5091) );
  OAI21_X1 U5379 ( .B1(n5827), .B2(n5826), .A(n5825), .ZN(n5960) );
  INV_X1 U5380 ( .A(n5737), .ZN(n5154) );
  INV_X1 U5381 ( .A(n5326), .ZN(n5153) );
  AOI21_X1 U5382 ( .B1(n4966), .B2(n4968), .A(n4965), .ZN(n4964) );
  INV_X1 U5383 ( .A(n5313), .ZN(n4965) );
  INV_X1 U5384 ( .A(n5165), .ZN(n4914) );
  NAND2_X1 U5385 ( .A1(n6530), .A2(n6532), .ZN(n6573) );
  AND2_X1 U5386 ( .A1(n8810), .A2(n8811), .ZN(n9127) );
  INV_X1 U5387 ( .A(n9254), .ZN(n9120) );
  NOR2_X1 U5388 ( .A1(n5060), .A2(n9120), .ZN(n5059) );
  INV_X1 U5389 ( .A(n5061), .ZN(n5060) );
  NAND2_X1 U5390 ( .A1(n6397), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n8675) );
  INV_X1 U5391 ( .A(n8009), .ZN(n6397) );
  NAND2_X1 U5392 ( .A1(n9273), .A2(n9117), .ZN(n4993) );
  OR2_X1 U5393 ( .A1(n8004), .A2(n9557), .ZN(n8009) );
  NAND2_X1 U5394 ( .A1(n6396), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n8004) );
  INV_X1 U5395 ( .A(n7945), .ZN(n6396) );
  OR2_X1 U5396 ( .A1(n7927), .A2(n7926), .ZN(n7945) );
  NAND2_X1 U5397 ( .A1(n6395), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n7927) );
  INV_X1 U5398 ( .A(n7858), .ZN(n6395) );
  OR2_X1 U5399 ( .A1(n7793), .A2(n7792), .ZN(n7858) );
  AND2_X1 U5400 ( .A1(n8638), .A2(n8639), .ZN(n8778) );
  AND2_X1 U5401 ( .A1(n8634), .A2(n8635), .ZN(n8777) );
  NOR2_X1 U5402 ( .A1(n7571), .A2(n10633), .ZN(n4998) );
  NAND2_X1 U5403 ( .A1(n8046), .A2(n4866), .ZN(n4985) );
  NOR2_X1 U5404 ( .A1(n7060), .A2(n10582), .ZN(n5051) );
  AND2_X1 U5405 ( .A1(n5055), .A2(n4898), .ZN(n5053) );
  NAND2_X1 U5406 ( .A1(n9347), .A2(n6959), .ZN(n8585) );
  NAND2_X1 U5407 ( .A1(n6509), .A2(n8813), .ZN(n7212) );
  NOR2_X1 U5408 ( .A1(n9394), .A2(n9240), .ZN(n9196) );
  OAI21_X1 U5409 ( .B1(P2_D_REG_1__SCAN_IN), .B2(n10361), .A(n10360), .ZN(
        n7208) );
  NOR2_X1 U5410 ( .A1(n7002), .A2(n7001), .ZN(n7210) );
  AND2_X1 U5411 ( .A1(n4900), .A2(n5136), .ZN(n5135) );
  INV_X1 U5412 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n6333) );
  NOR2_X1 U5413 ( .A1(P2_IR_REG_16__SCAN_IN), .A2(P2_IR_REG_17__SCAN_IN), .ZN(
        n5136) );
  AND2_X1 U5414 ( .A1(n6013), .A2(n6022), .ZN(n6163) );
  INV_X1 U5415 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n6177) );
  NAND2_X1 U5416 ( .A1(n6010), .A2(n6009), .ZN(n6137) );
  NAND2_X1 U5417 ( .A1(n5204), .A2(n5202), .ZN(n7343) );
  AOI21_X1 U5418 ( .B1(n4879), .B2(n5206), .A(n5203), .ZN(n5202) );
  NOR2_X1 U5419 ( .A1(n9722), .A2(n10182), .ZN(n5020) );
  NOR2_X1 U5420 ( .A1(n10173), .A2(n5019), .ZN(n5018) );
  INV_X1 U5421 ( .A(n5020), .ZN(n5019) );
  OR2_X1 U5422 ( .A1(n5927), .A2(n5926), .ZN(n5928) );
  NAND2_X1 U5423 ( .A1(n5024), .A2(n10223), .ZN(n5023) );
  OAI21_X1 U5424 ( .B1(n7481), .B2(n5637), .A(n8377), .ZN(n7602) );
  INV_X1 U5425 ( .A(n5909), .ZN(n5088) );
  NAND2_X1 U5426 ( .A1(n7192), .A2(n8253), .ZN(n7191) );
  AND2_X1 U5427 ( .A1(n5025), .A2(n6886), .ZN(n7091) );
  AND2_X1 U5428 ( .A1(n4860), .A2(n5026), .ZN(n5025) );
  NAND2_X1 U5429 ( .A1(n10046), .A2(n10053), .ZN(n10047) );
  NAND2_X1 U5430 ( .A1(n5222), .A2(n5338), .ZN(n5221) );
  INV_X1 U5431 ( .A(n5223), .ZN(n5222) );
  INV_X1 U5432 ( .A(n5345), .ZN(n5344) );
  AND2_X1 U5433 ( .A1(n5811), .A2(n5796), .ZN(n5808) );
  OAI21_X1 U5434 ( .B1(n5774), .B2(n5773), .A(n5772), .ZN(n5788) );
  INV_X1 U5435 ( .A(SI_23_), .ZN(n9590) );
  INV_X1 U5436 ( .A(n5221), .ZN(n5004) );
  NAND2_X1 U5437 ( .A1(n5414), .A2(n5224), .ZN(n5223) );
  INV_X1 U5438 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n5224) );
  NAND2_X1 U5439 ( .A1(n4926), .A2(n4925), .ZN(n5283) );
  NAND2_X1 U5440 ( .A1(n4925), .A2(n5542), .ZN(n4924) );
  INV_X1 U5441 ( .A(n5592), .ZN(n5143) );
  INV_X1 U5442 ( .A(SI_11_), .ZN(n9584) );
  OR2_X1 U5443 ( .A1(n5608), .A2(P1_IR_REG_10__SCAN_IN), .ZN(n5623) );
  NAND2_X1 U5444 ( .A1(n5283), .A2(n4924), .ZN(n5284) );
  XNOR2_X1 U5445 ( .A(n5286), .B(n9624), .ZN(n5592) );
  OR2_X1 U5446 ( .A1(n5276), .A2(n5275), .ZN(n5579) );
  AND2_X1 U5447 ( .A1(n5557), .A2(n5279), .ZN(n5577) );
  AND2_X1 U5448 ( .A1(n5563), .A2(n5562), .ZN(n5594) );
  NAND2_X1 U5449 ( .A1(n4927), .A2(SI_7_), .ZN(n5558) );
  OAI21_X1 U5450 ( .B1(n4927), .B2(SI_7_), .A(n5558), .ZN(n5544) );
  INV_X1 U5451 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n4922) );
  XNOR2_X1 U5452 ( .A(n6532), .B(n6531), .ZN(n8908) );
  AND2_X1 U5453 ( .A1(n5232), .A2(n7156), .ZN(n5129) );
  NAND2_X1 U5454 ( .A1(n6718), .A2(n6576), .ZN(n6577) );
  NAND2_X1 U5455 ( .A1(n5115), .A2(n6573), .ZN(n6715) );
  INV_X1 U5456 ( .A(n8908), .ZN(n5115) );
  NOR2_X1 U5457 ( .A1(n6580), .A2(n8825), .ZN(n8920) );
  NAND2_X1 U5458 ( .A1(n6577), .A2(n6578), .ZN(n7026) );
  AND4_X1 U5459 ( .A1(n7863), .A2(n7862), .A3(n7861), .A4(n7860), .ZN(n9003)
         );
  AND4_X1 U5460 ( .A1(n7053), .A2(n7052), .A3(n7051), .A4(n7050), .ZN(n7767)
         );
  NOR2_X1 U5461 ( .A1(n6142), .A2(n5137), .ZN(n6013) );
  INV_X1 U5462 ( .A(n5197), .ZN(n5137) );
  AOI21_X1 U5463 ( .B1(P2_REG2_REG_12__SCAN_IN), .B2(n7416), .A(n6844), .ZN(
        n6847) );
  NAND2_X1 U5464 ( .A1(n9157), .A2(n8809), .ZN(n9130) );
  AND2_X1 U5465 ( .A1(n8561), .A2(n8560), .ZN(n9155) );
  XNOR2_X1 U5466 ( .A(n9374), .B(n9173), .ZN(n9153) );
  NAND2_X1 U5467 ( .A1(n5038), .A2(n5037), .ZN(n9148) );
  NOR2_X1 U5468 ( .A1(n5041), .A2(n4904), .ZN(n5037) );
  NOR2_X1 U5469 ( .A1(n9197), .A2(n9386), .ZN(n9163) );
  AND2_X1 U5470 ( .A1(n8872), .A2(n9121), .ZN(n9122) );
  NAND2_X1 U5471 ( .A1(n9239), .A2(n9244), .ZN(n9240) );
  NAND2_X1 U5472 ( .A1(n4916), .A2(n4877), .ZN(n9231) );
  OAI21_X1 U5473 ( .B1(n8032), .B2(n5176), .A(n5173), .ZN(n4916) );
  OR2_X1 U5474 ( .A1(n9416), .A2(n9118), .ZN(n9275) );
  NAND2_X1 U5475 ( .A1(n8027), .A2(n8030), .ZN(n8019) );
  NOR2_X1 U5476 ( .A1(n8019), .A2(n9416), .ZN(n9266) );
  NAND2_X1 U5477 ( .A1(n5172), .A2(n8574), .ZN(n8801) );
  NAND2_X1 U5478 ( .A1(n8032), .A2(n8575), .ZN(n5172) );
  AND2_X1 U5479 ( .A1(n9298), .A2(n7939), .ZN(n8027) );
  INV_X1 U5480 ( .A(n9294), .ZN(n9290) );
  NAND2_X1 U5481 ( .A1(n7904), .A2(n7917), .ZN(n9288) );
  NAND2_X1 U5482 ( .A1(n5194), .A2(n5191), .ZN(n7941) );
  NOR2_X1 U5483 ( .A1(n4888), .A2(n5192), .ZN(n5191) );
  AND4_X1 U5484 ( .A1(n7720), .A2(n7719), .A3(n7718), .A4(n7717), .ZN(n7884)
         );
  NAND2_X1 U5485 ( .A1(n4998), .A2(n4997), .ZN(n7819) );
  NAND2_X1 U5486 ( .A1(n5190), .A2(n8630), .ZN(n7986) );
  OR2_X1 U5487 ( .A1(n7654), .A2(n8629), .ZN(n5190) );
  AND4_X1 U5488 ( .A1(n7631), .A2(n7630), .A3(n7629), .A4(n7628), .ZN(n7818)
         );
  AND4_X1 U5489 ( .A1(n7310), .A2(n7309), .A3(n7308), .A4(n7307), .ZN(n7657)
         );
  AND4_X1 U5490 ( .A1(n7167), .A2(n7166), .A3(n7165), .A4(n7164), .ZN(n7768)
         );
  INV_X1 U5491 ( .A(n4998), .ZN(n7664) );
  NAND2_X1 U5492 ( .A1(n5034), .A2(n5031), .ZN(n7662) );
  NOR2_X1 U5493 ( .A1(n4883), .A2(n5032), .ZN(n5031) );
  INV_X1 U5494 ( .A(n7568), .ZN(n5035) );
  AND2_X1 U5495 ( .A1(n8628), .A2(n7655), .ZN(n8776) );
  NOR2_X1 U5496 ( .A1(n4985), .A2(n7563), .ZN(n7775) );
  NAND2_X1 U5497 ( .A1(n7388), .A2(n7387), .ZN(n7569) );
  NAND2_X1 U5498 ( .A1(n7394), .A2(n7393), .ZN(n7763) );
  NAND2_X1 U5499 ( .A1(n8046), .A2(n7280), .ZN(n7230) );
  NAND2_X1 U5500 ( .A1(n8046), .A2(n4984), .ZN(n7399) );
  NAND2_X1 U5501 ( .A1(n7227), .A2(n8769), .ZN(n7394) );
  OR2_X1 U5502 ( .A1(n7223), .A2(n8769), .ZN(n7388) );
  OAI21_X1 U5503 ( .B1(n5054), .B2(n5052), .A(n5050), .ZN(n7222) );
  INV_X1 U5504 ( .A(n5053), .ZN(n5052) );
  AOI21_X1 U5505 ( .B1(n4859), .B2(n5053), .A(n5051), .ZN(n5050) );
  INV_X1 U5506 ( .A(n7376), .ZN(n5054) );
  AND2_X1 U5507 ( .A1(n8610), .A2(n8618), .ZN(n8768) );
  AND2_X1 U5508 ( .A1(n8044), .A2(n10582), .ZN(n8046) );
  AND3_X1 U5509 ( .A1(n10527), .A2(n6519), .A3(n4994), .ZN(n8044) );
  NOR2_X1 U5510 ( .A1(n8904), .A2(n7381), .ZN(n4994) );
  NOR2_X1 U5511 ( .A1(n8593), .A2(n5171), .ZN(n5170) );
  INV_X1 U5512 ( .A(n8589), .ZN(n5171) );
  NAND2_X1 U5513 ( .A1(n10527), .A2(n10539), .ZN(n7254) );
  NAND2_X1 U5514 ( .A1(n7256), .A2(n8589), .ZN(n7243) );
  AND2_X1 U5515 ( .A1(n5234), .A2(n6561), .ZN(n7259) );
  AND2_X1 U5516 ( .A1(n8584), .A2(n8585), .ZN(n9316) );
  INV_X1 U5517 ( .A(n9318), .ZN(n9346) );
  AND2_X1 U5518 ( .A1(n6499), .A2(n6707), .ZN(n9345) );
  AND2_X1 U5519 ( .A1(n6471), .A2(n10463), .ZN(n6472) );
  NAND2_X1 U5520 ( .A1(n7047), .A2(n7046), .ZN(n7386) );
  INV_X1 U5521 ( .A(n10625), .ZN(n10632) );
  AND3_X1 U5522 ( .A1(n7210), .A2(n7208), .A3(n7003), .ZN(n7080) );
  NAND2_X1 U5523 ( .A1(n6372), .A2(n6371), .ZN(n6374) );
  INV_X1 U5524 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n6023) );
  NOR2_X1 U5525 ( .A1(n6124), .A2(n5188), .ZN(n6132) );
  NAND2_X1 U5526 ( .A1(n6834), .A2(n6835), .ZN(n7134) );
  INV_X1 U5527 ( .A(n8197), .ZN(n8200) );
  NAND2_X1 U5528 ( .A1(n5008), .A2(n5006), .ZN(n8179) );
  AND2_X1 U5529 ( .A1(n5007), .A2(n5214), .ZN(n5006) );
  AND2_X1 U5530 ( .A1(n5215), .A2(n9833), .ZN(n5214) );
  NAND2_X1 U5531 ( .A1(n8176), .A2(n8177), .ZN(n9727) );
  INV_X1 U5532 ( .A(n8179), .ZN(n8176) );
  INV_X1 U5533 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n5598) );
  OR2_X1 U5534 ( .A1(n8185), .A2(n8184), .ZN(n8186) );
  NAND2_X1 U5535 ( .A1(n5219), .A2(n4905), .ZN(n9791) );
  NAND2_X1 U5536 ( .A1(n8105), .A2(n8104), .ZN(n5218) );
  NAND2_X1 U5537 ( .A1(n8106), .A2(n5220), .ZN(n5219) );
  OR2_X1 U5538 ( .A1(n8105), .A2(n8104), .ZN(n5220) );
  NAND2_X1 U5539 ( .A1(n9791), .A2(n8116), .ZN(n9803) );
  INV_X1 U5540 ( .A(n5381), .ZN(n5360) );
  XNOR2_X1 U5541 ( .A(n6317), .B(n8145), .ZN(n6587) );
  NAND2_X1 U5542 ( .A1(n6316), .A2(n6315), .ZN(n6317) );
  NAND2_X1 U5543 ( .A1(n8138), .A2(n8139), .ZN(n9748) );
  NAND2_X1 U5544 ( .A1(n8162), .A2(n9756), .ZN(n9830) );
  NAND2_X1 U5545 ( .A1(n5013), .A2(n5009), .ZN(n8162) );
  INV_X1 U5546 ( .A(n5011), .ZN(n5009) );
  NAND2_X1 U5547 ( .A1(n5357), .A2(n5356), .ZN(n5728) );
  NAND2_X1 U5548 ( .A1(n5002), .A2(n4889), .ZN(n6639) );
  INV_X1 U5549 ( .A(n9780), .ZN(n5210) );
  NOR2_X1 U5550 ( .A1(n9779), .A2(n5213), .ZN(n5212) );
  INV_X1 U5551 ( .A(n8186), .ZN(n5213) );
  AND2_X1 U5552 ( .A1(n8485), .A2(n8484), .ZN(n8490) );
  AND3_X1 U5553 ( .A1(n5396), .A2(n5395), .A3(n5394), .ZN(n8155) );
  AND4_X1 U5554 ( .A1(n5604), .A2(n5603), .A3(n5602), .A4(n5601), .ZN(n7352)
         );
  OR2_X1 U5555 ( .A1(n5421), .A2(n6884), .ZN(n5491) );
  OR2_X1 U5556 ( .A1(n5456), .A2(n5431), .ZN(n5432) );
  AOI21_X1 U5557 ( .B1(n6105), .B2(P1_REG2_REG_3__SCAN_IN), .A(n6099), .ZN(
        n9893) );
  AOI21_X1 U5558 ( .B1(P1_REG2_REG_6__SCAN_IN), .B2(n10431), .A(n10427), .ZN(
        n9906) );
  OR2_X1 U5559 ( .A1(n5675), .A2(P1_IR_REG_14__SCAN_IN), .ZN(n5688) );
  OR2_X1 U5560 ( .A1(n6322), .A2(n6002), .ZN(n6093) );
  OR2_X1 U5561 ( .A1(n5816), .A2(n5815), .ZN(n5951) );
  NAND2_X1 U5562 ( .A1(n9963), .A2(n5018), .ZN(n8520) );
  AOI21_X1 U5563 ( .B1(n5071), .B2(n5082), .A(n5070), .ZN(n5069) );
  NOR2_X1 U5564 ( .A1(n8509), .A2(n8429), .ZN(n5070) );
  NOR2_X1 U5565 ( .A1(n5084), .A2(n5942), .ZN(n5083) );
  INV_X1 U5566 ( .A(n5940), .ZN(n5084) );
  INV_X1 U5567 ( .A(n5102), .ZN(n5101) );
  AOI21_X1 U5568 ( .B1(n5102), .B2(n5100), .A(n5099), .ZN(n5098) );
  INV_X1 U5569 ( .A(n5768), .ZN(n5100) );
  AOI21_X1 U5570 ( .B1(n5768), .B2(n9995), .A(n5103), .ZN(n5102) );
  INV_X1 U5571 ( .A(n8426), .ZN(n5103) );
  NAND2_X1 U5572 ( .A1(n9996), .A2(n5768), .ZN(n5097) );
  NAND2_X1 U5573 ( .A1(n9999), .A2(n5768), .ZN(n9986) );
  OR2_X1 U5574 ( .A1(n9996), .A2(n9995), .ZN(n9999) );
  NAND2_X1 U5575 ( .A1(n5922), .A2(n5921), .ZN(n10067) );
  AND4_X1 U5576 ( .A1(n5732), .A2(n5731), .A3(n5730), .A4(n5729), .ZN(n10102)
         );
  NOR2_X1 U5577 ( .A1(n7872), .A2(n5022), .ZN(n10149) );
  INV_X1 U5578 ( .A(n5024), .ZN(n5022) );
  OAI21_X1 U5579 ( .B1(n10138), .B2(n8355), .A(n8286), .ZN(n10123) );
  NAND2_X1 U5580 ( .A1(n5355), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n5693) );
  INV_X1 U5581 ( .A(n5680), .ZN(n5355) );
  AND4_X1 U5582 ( .A1(n5715), .A2(n5714), .A3(n5713), .A4(n5712), .ZN(n9795)
         );
  OAI21_X1 U5583 ( .B1(n7806), .B2(n5113), .A(n8376), .ZN(n7877) );
  INV_X1 U5584 ( .A(n8414), .ZN(n5113) );
  AND4_X1 U5585 ( .A1(n5698), .A2(n5697), .A3(n5696), .A4(n5695), .ZN(n8110)
         );
  NAND2_X1 U5586 ( .A1(n5671), .A2(n8409), .ZN(n7806) );
  OR2_X1 U5587 ( .A1(n7691), .A2(n7690), .ZN(n5671) );
  NAND2_X1 U5588 ( .A1(n7697), .A2(n10249), .ZN(n7808) );
  AND4_X1 U5589 ( .A1(n5652), .A2(n5651), .A3(n5650), .A4(n5649), .ZN(n7693)
         );
  AND4_X1 U5590 ( .A1(n5685), .A2(n5684), .A3(n5683), .A4(n5682), .ZN(n7878)
         );
  AND4_X1 U5591 ( .A1(n5636), .A2(n5635), .A3(n5634), .A4(n5633), .ZN(n7603)
         );
  AND4_X1 U5592 ( .A1(n5670), .A2(n5669), .A3(n5668), .A4(n5667), .ZN(n8275)
         );
  INV_X1 U5593 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n6360) );
  OR2_X1 U5594 ( .A1(n5630), .A2(n6360), .ZN(n5646) );
  NAND2_X1 U5595 ( .A1(n5015), .A2(n5014), .ZN(n7608) );
  OAI21_X1 U5596 ( .B1(n7317), .B2(n8383), .A(n8403), .ZN(n7481) );
  NAND2_X1 U5597 ( .A1(n5353), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n5630) );
  INV_X1 U5598 ( .A(n5613), .ZN(n5353) );
  NAND2_X1 U5599 ( .A1(n7190), .A2(n8347), .ZN(n5089) );
  NAND2_X1 U5600 ( .A1(n7191), .A2(n8380), .ZN(n7317) );
  INV_X1 U5601 ( .A(n5586), .ZN(n5352) );
  INV_X1 U5602 ( .A(n5105), .ZN(n5104) );
  OAI21_X1 U5603 ( .B1(n5108), .B2(n5106), .A(n8400), .ZN(n5105) );
  OR2_X1 U5604 ( .A1(n8385), .A2(n5107), .ZN(n5106) );
  NAND2_X1 U5605 ( .A1(n5351), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n5571) );
  AND2_X1 U5606 ( .A1(n5539), .A2(n8463), .ZN(n6922) );
  AND4_X1 U5607 ( .A1(n5576), .A2(n5575), .A3(n5574), .A4(n5573), .ZN(n7181)
         );
  AND4_X1 U5608 ( .A1(n5528), .A2(n5527), .A3(n5526), .A4(n5525), .ZN(n6904)
         );
  AND2_X1 U5609 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .ZN(n5519) );
  AND2_X1 U5610 ( .A1(n6902), .A2(n6900), .ZN(n8339) );
  AND2_X1 U5611 ( .A1(n6886), .A2(n6664), .ZN(n6911) );
  NOR2_X1 U5612 ( .A1(n6885), .A2(n6890), .ZN(n6886) );
  NAND2_X1 U5613 ( .A1(n6621), .A2(n8055), .ZN(n6875) );
  NAND2_X1 U5614 ( .A1(n5475), .A2(n8456), .ZN(n6877) );
  NOR2_X1 U5615 ( .A1(n6278), .A2(n6453), .ZN(n6866) );
  NAND2_X1 U5616 ( .A1(n5963), .A2(n5962), .ZN(n8333) );
  NAND2_X1 U5617 ( .A1(n5829), .A2(n5828), .ZN(n10169) );
  NAND2_X1 U5618 ( .A1(n5417), .A2(n5416), .ZN(n10109) );
  OR2_X1 U5619 ( .A1(n8319), .A2(n8329), .ZN(n10273) );
  NAND2_X1 U5620 ( .A1(n6550), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n5030) );
  AND2_X1 U5621 ( .A1(n5992), .A2(n8491), .ZN(n10269) );
  XNOR2_X1 U5622 ( .A(n5961), .B(n5967), .ZN(n8540) );
  NAND2_X1 U5623 ( .A1(n5971), .A2(n5965), .ZN(n5961) );
  XNOR2_X1 U5624 ( .A(n5958), .B(SI_29_), .ZN(n8550) );
  XNOR2_X1 U5625 ( .A(n5827), .B(n5826), .ZN(n8728) );
  NAND2_X1 U5626 ( .A1(n5868), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5869) );
  NAND2_X1 U5627 ( .A1(n5859), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5861) );
  INV_X1 U5628 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n5864) );
  XNOR2_X1 U5629 ( .A(n5756), .B(n5744), .ZN(n8562) );
  AND2_X1 U5630 ( .A1(n5296), .A2(n5295), .ZN(n5155) );
  INV_X1 U5631 ( .A(n5638), .ZN(n5296) );
  XNOR2_X1 U5632 ( .A(n4951), .B(n4880), .ZN(n7105) );
  AOI21_X1 U5633 ( .B1(n5578), .B2(n5577), .A(n4952), .ZN(n4951) );
  INV_X1 U5634 ( .A(n5579), .ZN(n4952) );
  OR2_X1 U5635 ( .A1(n5594), .A2(n10319), .ZN(n5566) );
  NAND2_X1 U5636 ( .A1(n5243), .A2(n4962), .ZN(n4961) );
  OR2_X1 U5637 ( .A1(n5254), .A2(n4963), .ZN(n4962) );
  AND2_X1 U5638 ( .A1(n5265), .A2(n5264), .ZN(n5492) );
  NAND2_X1 U5639 ( .A1(n5256), .A2(n4953), .ZN(n5465) );
  OR2_X1 U5640 ( .A1(n4954), .A2(SI_2_), .ZN(n4953) );
  OR2_X1 U5641 ( .A1(n6229), .A2(P2_U3152), .ZN(n6478) );
  NAND2_X1 U5642 ( .A1(n5121), .A2(n5124), .ZN(n8930) );
  NAND2_X1 U5643 ( .A1(n8718), .A2(n8717), .ZN(n9379) );
  AND4_X1 U5644 ( .A1(n7429), .A2(n7428), .A3(n7427), .A4(n7426), .ZN(n7825)
         );
  AOI21_X1 U5645 ( .B1(n5133), .B2(n5131), .A(n4867), .ZN(n5130) );
  INV_X1 U5646 ( .A(n5133), .ZN(n5132) );
  NAND2_X1 U5647 ( .A1(n7713), .A2(n7712), .ZN(n9446) );
  NAND2_X1 U5648 ( .A1(n7999), .A2(n7998), .ZN(n9422) );
  OAI21_X1 U5649 ( .B1(n5124), .B2(n5123), .A(n4906), .ZN(n5122) );
  OR2_X2 U5650 ( .A1(n5066), .A2(n5065), .ZN(n9352) );
  AND3_X1 U5651 ( .A1(n8679), .A2(n8678), .A3(n8677), .ZN(n8957) );
  AND2_X1 U5652 ( .A1(n8573), .A2(n8572), .ZN(n9206) );
  NAND2_X1 U5653 ( .A1(n7857), .A2(n7856), .ZN(n9437) );
  NAND2_X1 U5654 ( .A1(n7854), .A2(n8727), .ZN(n7857) );
  AND2_X1 U5655 ( .A1(n8920), .A2(n9345), .ZN(n8947) );
  AND4_X1 U5656 ( .A1(n6996), .A2(n6995), .A3(n6994), .A4(n6993), .ZN(n7390)
         );
  AND4_X1 U5657 ( .A1(n7122), .A2(n7121), .A3(n7120), .A4(n7119), .ZN(n7562)
         );
  NAND2_X1 U5658 ( .A1(n8674), .A2(n8673), .ZN(n9404) );
  NAND2_X1 U5659 ( .A1(n6479), .A2(n6669), .ZN(n8949) );
  NAND2_X1 U5660 ( .A1(n8830), .A2(n6553), .ZN(n8531) );
  AND2_X1 U5661 ( .A1(n8920), .A2(n9346), .ZN(n9005) );
  INV_X1 U5662 ( .A(n5119), .ZN(n5118) );
  OAI21_X1 U5663 ( .B1(n6578), .B2(n5120), .A(n7028), .ZN(n5119) );
  NAND2_X1 U5664 ( .A1(n7026), .A2(n7025), .ZN(n7027) );
  AND2_X1 U5665 ( .A1(n6490), .A2(n9304), .ZN(n8937) );
  INV_X1 U5666 ( .A(n8050), .ZN(n10582) );
  NOR2_X1 U5667 ( .A1(n6580), .A2(n6579), .ZN(n8941) );
  NAND2_X1 U5668 ( .A1(n8962), .A2(n8888), .ZN(n9010) );
  AND4_X1 U5669 ( .A1(n7798), .A2(n7797), .A3(n7796), .A4(n7795), .ZN(n7970)
         );
  NAND2_X1 U5670 ( .A1(n7791), .A2(n7790), .ZN(n9441) );
  INV_X1 U5671 ( .A(n8937), .ZN(n9017) );
  INV_X1 U5672 ( .A(n8957), .ZN(n9280) );
  INV_X1 U5673 ( .A(n7259), .ZN(n9347) );
  INV_X1 U5674 ( .A(n9022), .ZN(n9041) );
  AOI21_X1 U5675 ( .B1(n10492), .B2(P2_REG2_REG_2__SCAN_IN), .A(n10488), .ZN(
        n6794) );
  AOI21_X1 U5676 ( .B1(n6695), .B2(P2_REG2_REG_5__SCAN_IN), .A(n6804), .ZN(
        n6771) );
  AOI21_X1 U5677 ( .B1(n6970), .B2(P2_REG2_REG_7__SCAN_IN), .A(n6780), .ZN(
        n6736) );
  NAND2_X1 U5678 ( .A1(n6241), .A2(n6240), .ZN(n10486) );
  NOR2_X1 U5679 ( .A1(n9073), .A2(n9072), .ZN(n9089) );
  AND2_X1 U5680 ( .A1(n6708), .A2(n6492), .ZN(n10493) );
  INV_X1 U5681 ( .A(n9113), .ZN(n9368) );
  NOR2_X1 U5682 ( .A1(n9113), .A2(n9136), .ZN(n4995) );
  NAND2_X1 U5683 ( .A1(n5185), .A2(n8806), .ZN(n9170) );
  NAND2_X1 U5684 ( .A1(n5039), .A2(n5045), .ZN(n9162) );
  INV_X1 U5685 ( .A(n5043), .ZN(n5040) );
  AND2_X1 U5686 ( .A1(n8719), .A2(n6608), .ZN(n9188) );
  INV_X1 U5687 ( .A(n5049), .ZN(n5036) );
  NAND2_X1 U5688 ( .A1(n8701), .A2(n8700), .ZN(n9391) );
  AND2_X1 U5689 ( .A1(n5062), .A2(n9119), .ZN(n9248) );
  NAND2_X1 U5690 ( .A1(n9414), .A2(n5063), .ZN(n9265) );
  INV_X1 U5691 ( .A(n9422), .ZN(n8030) );
  NAND2_X1 U5692 ( .A1(n9307), .A2(n7216), .ZN(n9272) );
  OAI21_X1 U5693 ( .B1(n7376), .B2(n4859), .A(n5055), .ZN(n8041) );
  INV_X1 U5694 ( .A(n9285), .ZN(n9337) );
  OR2_X1 U5695 ( .A1(n6562), .A2(n6515), .ZN(n6518) );
  OR2_X1 U5696 ( .A1(n6562), .A2(n4956), .ZN(n6566) );
  AND2_X1 U5697 ( .A1(n10362), .A2(n6489), .ZN(n9350) );
  OR2_X1 U5698 ( .A1(n9352), .A2(n9351), .ZN(n10510) );
  INV_X1 U5699 ( .A(n9139), .ZN(n9353) );
  INV_X1 U5700 ( .A(n9272), .ZN(n9336) );
  NAND2_X1 U5701 ( .A1(n9363), .A2(n9362), .ZN(n9456) );
  NAND2_X1 U5702 ( .A1(n9359), .A2(n10511), .ZN(n9363) );
  OR2_X1 U5703 ( .A1(n9371), .A2(n10637), .ZN(n4991) );
  NOR2_X1 U5704 ( .A1(n9372), .A2(n4990), .ZN(n4989) );
  AND2_X2 U5705 ( .A1(n7080), .A2(n7209), .ZN(n10646) );
  NOR2_X1 U5706 ( .A1(n6230), .A2(P2_U3152), .ZN(n10464) );
  AND2_X1 U5707 ( .A1(n5199), .A2(n6231), .ZN(n5198) );
  AND2_X1 U5708 ( .A1(n6371), .A2(n5200), .ZN(n5199) );
  INV_X1 U5709 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n5200) );
  NAND2_X1 U5710 ( .A1(n6035), .A2(n6234), .ZN(n7585) );
  XNOR2_X1 U5711 ( .A(n6021), .B(n6024), .ZN(n7206) );
  NAND2_X1 U5712 ( .A1(n6020), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6021) );
  NAND2_X1 U5713 ( .A1(n6039), .A2(n6023), .ZN(n6020) );
  INV_X1 U5714 ( .A(n8813), .ZN(n8819) );
  OR2_X1 U5715 ( .A1(n6337), .A2(n6336), .ZN(n6338) );
  NAND2_X1 U5716 ( .A1(n6017), .A2(n6016), .ZN(n6243) );
  CLKBUF_X1 U5717 ( .A(n9737), .Z(n9738) );
  OR2_X1 U5718 ( .A1(n9714), .A2(n8216), .ZN(n8206) );
  AND3_X1 U5719 ( .A1(n5408), .A2(n5407), .A3(n5406), .ZN(n10104) );
  NAND2_X1 U5720 ( .A1(n5390), .A2(n5389), .ZN(n10075) );
  NAND2_X1 U5721 ( .A1(n5691), .A2(n5690), .ZN(n10237) );
  NAND2_X1 U5722 ( .A1(n5400), .A2(n5399), .ZN(n10213) );
  NAND2_X1 U5723 ( .A1(n5378), .A2(n5377), .ZN(n10205) );
  INV_X1 U5724 ( .A(n9860), .ZN(n9848) );
  NAND2_X1 U5725 ( .A1(n5678), .A2(n5677), .ZN(n7809) );
  OR2_X1 U5726 ( .A1(n7789), .A2(n5474), .ZN(n5678) );
  CLKBUF_X1 U5727 ( .A(n9851), .Z(n9837) );
  INV_X1 U5728 ( .A(n8446), .ZN(n8447) );
  INV_X1 U5729 ( .A(n10001), .ZN(n9872) );
  NAND2_X1 U5730 ( .A1(n5753), .A2(n5752), .ZN(n10026) );
  INV_X1 U5731 ( .A(n8155), .ZN(n10094) );
  NAND4_X1 U5732 ( .A1(n5510), .A2(n5509), .A3(n5508), .A4(n5507), .ZN(n6629)
         );
  OR2_X1 U5733 ( .A1(n6093), .A2(P1_U3084), .ZN(n9883) );
  NAND2_X1 U5734 ( .A1(n5446), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n5449) );
  NOR2_X1 U5735 ( .A1(n8077), .A2(n8078), .ZN(n6365) );
  NOR2_X1 U5736 ( .A1(n6056), .A2(n7364), .ZN(n7476) );
  AOI21_X1 U5737 ( .B1(n5858), .B2(n10140), .A(n5857), .ZN(n10171) );
  INV_X1 U5738 ( .A(n5856), .ZN(n5857) );
  AOI22_X1 U5739 ( .A1(n9870), .A2(n10143), .B1(n5982), .B2(n9868), .ZN(n5856)
         );
  NAND2_X1 U5740 ( .A1(n5758), .A2(n5757), .ZN(n10189) );
  NAND2_X1 U5741 ( .A1(n5349), .A2(n5348), .ZN(n10197) );
  NAND2_X1 U5742 ( .A1(n5093), .A2(n5096), .ZN(n10120) );
  INV_X1 U5743 ( .A(n5094), .ZN(n5093) );
  NAND2_X1 U5744 ( .A1(n7688), .A2(n5916), .ZN(n7805) );
  NAND2_X1 U5745 ( .A1(n5914), .A2(n5913), .ZN(n7598) );
  NAND2_X1 U5746 ( .A1(n5643), .A2(n5642), .ZN(n10254) );
  NAND2_X1 U5747 ( .A1(n6921), .A2(n8384), .ZN(n6950) );
  NAND2_X1 U5748 ( .A1(n6918), .A2(n5904), .ZN(n6949) );
  NAND2_X1 U5749 ( .A1(n10148), .A2(n6205), .ZN(n10115) );
  INV_X1 U5750 ( .A(n9951), .ZN(n10019) );
  OR2_X1 U5751 ( .A1(n10405), .A2(n5988), .ZN(n10145) );
  INV_X1 U5752 ( .A(n10115), .ZN(n10156) );
  AND2_X1 U5753 ( .A1(n10148), .A2(n6452), .ZN(n10097) );
  INV_X2 U5754 ( .A(n10607), .ZN(n10608) );
  INV_X1 U5755 ( .A(n8233), .ZN(n8326) );
  INV_X1 U5756 ( .A(n8100), .ZN(n5985) );
  AND2_X1 U5757 ( .A1(n10165), .A2(n10164), .ZN(n10277) );
  INV_X1 U5758 ( .A(n4974), .ZN(n10178) );
  NOR2_X1 U5759 ( .A1(n8506), .A2(n4976), .ZN(n4975) );
  AND2_X1 U5760 ( .A1(n8501), .A2(n5984), .ZN(n4976) );
  INV_X1 U5761 ( .A(n10007), .ZN(n10287) );
  INV_X2 U5762 ( .A(n10609), .ZN(n10612) );
  AND2_X1 U5763 ( .A1(n5111), .A2(n5366), .ZN(n5109) );
  AOI21_X1 U5764 ( .B1(n5971), .B2(n5970), .A(n5241), .ZN(n5974) );
  NAND2_X1 U5765 ( .A1(n5345), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5347) );
  NAND2_X1 U5766 ( .A1(n4979), .A2(n5388), .ZN(n8662) );
  OAI21_X1 U5767 ( .B1(n5162), .B2(n4968), .A(n4966), .ZN(n5719) );
  NAND2_X1 U5768 ( .A1(n5702), .A2(n5309), .ZN(n5717) );
  NAND2_X1 U5769 ( .A1(n5162), .A2(n5163), .ZN(n5701) );
  NAND2_X1 U5770 ( .A1(n4973), .A2(n4972), .ZN(n5620) );
  INV_X1 U5771 ( .A(n5140), .ZN(n4973) );
  NAND2_X1 U5772 ( .A1(n5145), .A2(n5144), .ZN(n5607) );
  AND2_X1 U5773 ( .A1(n5529), .A2(n5498), .ZN(n9895) );
  NAND2_X1 U5774 ( .A1(n5467), .A2(n5256), .ZN(n5481) );
  NOR2_X1 U5775 ( .A1(n7526), .A2(n7525), .ZN(n10394) );
  NOR2_X1 U5776 ( .A1(n10392), .A2(n10391), .ZN(n7525) );
  OR2_X1 U5777 ( .A1(n8828), .A2(n8827), .ZN(n5177) );
  NAND2_X1 U5778 ( .A1(n4988), .A2(n4986), .ZN(P2_U3549) );
  OR2_X1 U5779 ( .A1(n10642), .A2(n4987), .ZN(n4986) );
  NAND2_X1 U5780 ( .A1(n9458), .A2(n10642), .ZN(n4988) );
  INV_X1 U5781 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n4987) );
  NAND2_X1 U5782 ( .A1(n9856), .A2(n4999), .ZN(n9865) );
  AND2_X1 U5783 ( .A1(n9038), .A2(n7381), .ZN(n4859) );
  AND2_X1 U5784 ( .A1(n4863), .A2(n5027), .ZN(n4860) );
  AND3_X1 U5785 ( .A1(n5197), .A2(n5187), .A3(n4996), .ZN(n4861) );
  AND2_X1 U5786 ( .A1(n8313), .A2(n8431), .ZN(n8509) );
  OR2_X1 U5787 ( .A1(n5286), .A2(SI_10_), .ZN(n4862) );
  OR2_X1 U5788 ( .A1(n9136), .A2(n9155), .ZN(n8810) );
  AND2_X1 U5789 ( .A1(n6664), .A2(n10574), .ZN(n4863) );
  NAND2_X1 U5790 ( .A1(n5095), .A2(n5096), .ZN(n4864) );
  OR2_X1 U5791 ( .A1(n8821), .A2(n5116), .ZN(n4865) );
  OR2_X1 U5792 ( .A1(n5413), .A2(P1_IR_REG_19__SCAN_IN), .ZN(n5846) );
  AND2_X1 U5793 ( .A1(n4984), .A2(n4983), .ZN(n4866) );
  AND2_X1 U5794 ( .A1(n7710), .A2(n7709), .ZN(n4867) );
  AND2_X1 U5795 ( .A1(n6614), .A2(n6613), .ZN(n9172) );
  AND2_X1 U5796 ( .A1(n9127), .A2(n4891), .ZN(n4868) );
  AND2_X1 U5797 ( .A1(n8615), .A2(n8614), .ZN(n4869) );
  AND2_X1 U5798 ( .A1(n4862), .A2(n5290), .ZN(n5144) );
  INV_X1 U5799 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n6016) );
  AND2_X1 U5800 ( .A1(n5917), .A2(n5916), .ZN(n4870) );
  AND2_X1 U5801 ( .A1(n5905), .A2(n5904), .ZN(n4871) );
  AND2_X1 U5802 ( .A1(n8128), .A2(n8124), .ZN(n4872) );
  INV_X1 U5803 ( .A(n7138), .ZN(n5026) );
  NAND2_X1 U5804 ( .A1(n6886), .A2(n4863), .ZN(n6910) );
  AND2_X1 U5805 ( .A1(n5002), .A2(n4878), .ZN(n4873) );
  INV_X2 U5806 ( .A(n6535), .ZN(n6560) );
  OR2_X1 U5807 ( .A1(n9821), .A2(n8148), .ZN(n5013) );
  XOR2_X1 U5808 ( .A(n6569), .B(n6570), .Z(n4875) );
  NAND4_X1 U5809 ( .A1(n5450), .A2(n5449), .A3(n5448), .A4(n5447), .ZN(n6217)
         );
  NOR2_X1 U5810 ( .A1(n10158), .A2(n10157), .ZN(n5094) );
  NAND2_X1 U5811 ( .A1(n10122), .A2(n8239), .ZN(n10056) );
  AND4_X1 U5812 ( .A1(n5005), .A2(n5335), .A3(n5336), .A4(n5337), .ZN(n5863)
         );
  OR2_X1 U5813 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n4876) );
  AND2_X1 U5814 ( .A1(n8797), .A2(n8798), .ZN(n4877) );
  OR2_X1 U5815 ( .A1(n6595), .A2(n6594), .ZN(n4878) );
  INV_X1 U5816 ( .A(n7563), .ZN(n10614) );
  NAND2_X1 U5817 ( .A1(n5863), .A2(n5864), .ZN(n5859) );
  NAND2_X1 U5818 ( .A1(n5186), .A2(n6008), .ZN(n6123) );
  INV_X1 U5819 ( .A(n8904), .ZN(n10539) );
  OR2_X1 U5820 ( .A1(n9409), .A2(n9024), .ZN(n9119) );
  OAI21_X1 U5821 ( .B1(n9994), .B2(n5939), .A(n5938), .ZN(n9978) );
  AND2_X1 U5822 ( .A1(n7325), .A2(n5205), .ZN(n4879) );
  NAND2_X1 U5823 ( .A1(n8142), .A2(n9747), .ZN(n9821) );
  NAND2_X1 U5824 ( .A1(n5075), .A2(n5940), .ZN(n9962) );
  NAND2_X1 U5825 ( .A1(n5013), .A2(n8151), .ZN(n9755) );
  NAND2_X1 U5826 ( .A1(n9811), .A2(n8186), .ZN(n9778) );
  XOR2_X1 U5827 ( .A(n5277), .B(SI_9_), .Z(n4880) );
  NAND2_X1 U5828 ( .A1(n8553), .A2(n8552), .ZN(n9136) );
  AND2_X1 U5829 ( .A1(n8759), .A2(n8746), .ZN(n4881) );
  AND2_X1 U5830 ( .A1(n6972), .A2(n6971), .ZN(n7280) );
  AND2_X1 U5831 ( .A1(n9830), .A2(n9831), .ZN(n4882) );
  AND2_X1 U5832 ( .A1(n8429), .A2(n8430), .ZN(n8473) );
  INV_X1 U5833 ( .A(n8473), .ZN(n5082) );
  NAND2_X1 U5834 ( .A1(n5711), .A2(n5710), .ZN(n10155) );
  NOR2_X1 U5835 ( .A1(n7567), .A2(n7566), .ZN(n4883) );
  NAND2_X1 U5836 ( .A1(n5777), .A2(n5776), .ZN(n10182) );
  AND2_X1 U5837 ( .A1(n5097), .A2(n5102), .ZN(n4884) );
  AND4_X1 U5838 ( .A1(n6526), .A2(n6525), .A3(n6524), .A4(n6523), .ZN(n9319)
         );
  AND2_X1 U5839 ( .A1(n5284), .A2(n5592), .ZN(n4885) );
  INV_X1 U5840 ( .A(n10173), .ZN(n8524) );
  NAND2_X1 U5841 ( .A1(n5814), .A2(n5813), .ZN(n10173) );
  NAND2_X1 U5842 ( .A1(n9963), .A2(n5020), .ZN(n5021) );
  AND2_X1 U5843 ( .A1(n4966), .A2(n4914), .ZN(n4886) );
  NAND2_X1 U5844 ( .A1(n10060), .A2(n5923), .ZN(n4887) );
  NAND2_X1 U5845 ( .A1(n8644), .A2(n7896), .ZN(n4888) );
  AND2_X1 U5846 ( .A1(n4878), .A2(n6637), .ZN(n4889) );
  NAND2_X1 U5847 ( .A1(n9231), .A2(n8802), .ZN(n4890) );
  AND2_X1 U5848 ( .A1(n8745), .A2(n8744), .ZN(n4891) );
  NAND2_X1 U5849 ( .A1(n8564), .A2(n8563), .ZN(n9394) );
  AND2_X1 U5850 ( .A1(n8408), .A2(n8378), .ZN(n8351) );
  NAND2_X1 U5851 ( .A1(n5346), .A2(n5340), .ZN(n4892) );
  INV_X1 U5852 ( .A(n4967), .ZN(n4966) );
  OAI21_X1 U5853 ( .B1(n5160), .B2(n4968), .A(n5716), .ZN(n4967) );
  INV_X1 U5854 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n10319) );
  AND2_X1 U5855 ( .A1(n5231), .A2(n5479), .ZN(n4893) );
  NAND2_X1 U5856 ( .A1(n8806), .A2(n8757), .ZN(n4894) );
  OR2_X1 U5857 ( .A1(n5413), .A2(n5223), .ZN(n4895) );
  NAND2_X1 U5858 ( .A1(n5145), .A2(n4862), .ZN(n4896) );
  AND2_X1 U5859 ( .A1(n8427), .A2(n8432), .ZN(n9970) );
  INV_X1 U5860 ( .A(n9970), .ZN(n5099) );
  INV_X1 U5861 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n6009) );
  AND3_X1 U5862 ( .A1(n6487), .A2(n6486), .A3(n6485), .ZN(n10565) );
  INV_X1 U5863 ( .A(n4940), .ZN(n4939) );
  OAI21_X1 U5864 ( .B1(n5227), .B2(n4941), .A(n8661), .ZN(n4940) );
  NOR2_X1 U5865 ( .A1(P1_IR_REG_26__SCAN_IN), .A2(P1_IR_REG_25__SCAN_IN), .ZN(
        n4897) );
  OR2_X1 U5866 ( .A1(n7021), .A2(n8050), .ZN(n4898) );
  NAND2_X1 U5867 ( .A1(n8808), .A2(n8742), .ZN(n9171) );
  INV_X1 U5868 ( .A(n9171), .ZN(n8807) );
  AND2_X1 U5869 ( .A1(n5285), .A2(n5284), .ZN(n4899) );
  AND2_X1 U5870 ( .A1(n6025), .A2(n6333), .ZN(n4900) );
  OR2_X1 U5871 ( .A1(n9409), .A2(n9256), .ZN(n4901) );
  AND2_X1 U5872 ( .A1(n5733), .A2(n8374), .ZN(n10119) );
  INV_X1 U5873 ( .A(n10119), .ZN(n5095) );
  INV_X1 U5874 ( .A(n7025), .ZN(n5120) );
  INV_X1 U5875 ( .A(n5072), .ZN(n5071) );
  NAND2_X1 U5876 ( .A1(n8509), .A2(n8429), .ZN(n5072) );
  INV_X1 U5877 ( .A(n8810), .ZN(n5183) );
  INV_X1 U5878 ( .A(n5256), .ZN(n4963) );
  NAND2_X1 U5879 ( .A1(n4954), .A2(SI_2_), .ZN(n5256) );
  NAND2_X1 U5880 ( .A1(n8684), .A2(n8683), .ZN(n8872) );
  NAND2_X1 U5881 ( .A1(n7979), .A2(n7984), .ZN(n7936) );
  NAND2_X1 U5882 ( .A1(n7157), .A2(n7156), .ZN(n7405) );
  XNOR2_X1 U5883 ( .A(n5974), .B(n5973), .ZN(n9704) );
  NAND2_X1 U5884 ( .A1(n7134), .A2(n7133), .ZN(n7326) );
  INV_X1 U5885 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n4956) );
  OR2_X1 U5886 ( .A1(n5375), .A2(n5154), .ZN(n4902) );
  NAND2_X1 U5887 ( .A1(n7803), .A2(n5918), .ZN(n7871) );
  NAND2_X1 U5888 ( .A1(n5089), .A2(n5909), .ZN(n7315) );
  INV_X1 U5889 ( .A(n8384), .ZN(n5107) );
  NAND2_X1 U5890 ( .A1(n8003), .A2(n8002), .ZN(n9416) );
  NAND2_X1 U5891 ( .A1(n8712), .A2(n8711), .ZN(n9386) );
  INV_X1 U5892 ( .A(n9386), .ZN(n5048) );
  OR2_X1 U5893 ( .A1(n7872), .A2(n5023), .ZN(n4903) );
  NAND2_X1 U5894 ( .A1(n5219), .A2(n5218), .ZN(n9790) );
  NOR3_X1 U5895 ( .A1(n8019), .A2(n9404), .A3(n4993), .ZN(n9239) );
  NAND2_X1 U5896 ( .A1(n9802), .A2(n4872), .ZN(n9840) );
  INV_X1 U5897 ( .A(n5949), .ZN(n7872) );
  NOR2_X1 U5898 ( .A1(n7808), .A2(n7809), .ZN(n5949) );
  INV_X1 U5899 ( .A(n6010), .ZN(n6142) );
  INV_X1 U5900 ( .A(n10046), .ZN(n10074) );
  NOR2_X1 U5901 ( .A1(n10083), .A2(n10075), .ZN(n10046) );
  AND2_X1 U5902 ( .A1(n9169), .A2(n9185), .ZN(n4904) );
  INV_X1 U5903 ( .A(n5064), .ZN(n5063) );
  AND2_X1 U5904 ( .A1(n8115), .A2(n5218), .ZN(n4905) );
  INV_X1 U5905 ( .A(n4992), .ZN(n9267) );
  NOR2_X1 U5906 ( .A1(n8019), .A2(n4993), .ZN(n4992) );
  NAND2_X1 U5907 ( .A1(n8928), .A2(n8927), .ZN(n4906) );
  AND2_X1 U5908 ( .A1(n5740), .A2(n9590), .ZN(n4907) );
  AND2_X1 U5909 ( .A1(n5127), .A2(n8929), .ZN(n4908) );
  INV_X1 U5910 ( .A(P2_RD_REG_SCAN_IN), .ZN(n4918) );
  AND2_X1 U5911 ( .A1(n6886), .A2(n4860), .ZN(n4909) );
  AOI21_X1 U5912 ( .B1(n7372), .B2(n8764), .A(n6986), .ZN(n8042) );
  OAI21_X1 U5913 ( .B1(n7085), .B2(n5908), .A(n5907), .ZN(n7190) );
  INV_X1 U5914 ( .A(n7620), .ZN(n5131) );
  INV_X1 U5915 ( .A(n9756), .ZN(n5216) );
  INV_X1 U5916 ( .A(n5015), .ZN(n7486) );
  NOR2_X1 U5917 ( .A1(n7197), .A2(n10268), .ZN(n5015) );
  NAND4_X1 U5918 ( .A1(n5004), .A2(n5336), .A3(n5335), .A4(n5337), .ZN(n4910)
         );
  AND2_X1 U5919 ( .A1(n8812), .A2(n8813), .ZN(n4911) );
  XNOR2_X1 U5920 ( .A(n5347), .B(n5346), .ZN(n5851) );
  INV_X1 U5921 ( .A(n7016), .ZN(n5027) );
  AND2_X1 U5922 ( .A1(n5445), .A2(n5028), .ZN(n6347) );
  NAND2_X1 U5923 ( .A1(n7624), .A2(n7623), .ZN(n9451) );
  INV_X1 U5924 ( .A(n9451), .ZN(n4997) );
  NAND2_X1 U5925 ( .A1(n7108), .A2(n7107), .ZN(n7587) );
  INV_X1 U5926 ( .A(n7587), .ZN(n4983) );
  NAND2_X1 U5927 ( .A1(n5343), .A2(n5363), .ZN(n5850) );
  INV_X1 U5928 ( .A(n9853), .ZN(n9855) );
  NAND2_X1 U5929 ( .A1(n6223), .A2(n6324), .ZN(n9853) );
  NAND2_X1 U5930 ( .A1(n5629), .A2(n5628), .ZN(n10263) );
  INV_X1 U5931 ( .A(n10263), .ZN(n5014) );
  XNOR2_X1 U5932 ( .A(n6233), .B(n6371), .ZN(n6492) );
  INV_X1 U5933 ( .A(n5369), .ZN(n10323) );
  AND2_X1 U5934 ( .A1(n6232), .A2(n5198), .ZN(n6376) );
  NAND3_X1 U5935 ( .A1(n4918), .A2(P2_ADDR_REG_19__SCAN_IN), .A3(
        P1_ADDR_REG_19__SCAN_IN), .ZN(n4917) );
  NAND3_X1 U5936 ( .A1(n4922), .A2(n4921), .A3(n4920), .ZN(n4919) );
  NAND3_X1 U5937 ( .A1(n5144), .A2(n4924), .A3(n5283), .ZN(n4923) );
  NAND2_X1 U5938 ( .A1(n5235), .A2(n5280), .ZN(n4925) );
  NAND2_X1 U5939 ( .A1(n5577), .A2(n5280), .ZN(n4926) );
  OAI21_X1 U5940 ( .B1(n6550), .B2(n4929), .A(n4928), .ZN(n4927) );
  NAND2_X1 U5941 ( .A1(n6550), .A2(P1_DATAO_REG_7__SCAN_IN), .ZN(n4928) );
  NAND2_X1 U5942 ( .A1(n4932), .A2(n5177), .ZN(P2_U3244) );
  NAND2_X1 U5943 ( .A1(n4933), .A2(n6236), .ZN(n4932) );
  NAND2_X1 U5944 ( .A1(n4935), .A2(n4934), .ZN(n4933) );
  NAND2_X1 U5945 ( .A1(n5139), .A2(n5138), .ZN(n4935) );
  OAI21_X1 U5946 ( .B1(n8658), .B2(n4941), .A(n4939), .ZN(n8668) );
  OAI21_X1 U5947 ( .B1(n8658), .B2(n4937), .A(n4936), .ZN(n5238) );
  NAND2_X1 U5948 ( .A1(n9274), .A2(n8659), .ZN(n4941) );
  NAND2_X1 U5949 ( .A1(n8705), .A2(n8746), .ZN(n8702) );
  NAND3_X1 U5950 ( .A1(n8814), .A2(n8747), .A3(n8748), .ZN(n4947) );
  NAND3_X1 U5951 ( .A1(n4949), .A2(n9147), .A3(n8743), .ZN(n4948) );
  NAND3_X1 U5952 ( .A1(n4950), .A2(n5146), .A3(n8807), .ZN(n4949) );
  NAND3_X1 U5953 ( .A1(n8613), .A2(n8611), .A3(n8612), .ZN(n4959) );
  NOR2_X1 U5954 ( .A1(n5255), .A2(n4963), .ZN(n4960) );
  NAND3_X1 U5955 ( .A1(n4971), .A2(n5155), .A3(n4970), .ZN(n5654) );
  NAND4_X1 U5956 ( .A1(n5144), .A2(n5619), .A3(n5282), .A4(n5541), .ZN(n4970)
         );
  NAND2_X1 U5957 ( .A1(n5282), .A2(n5541), .ZN(n5285) );
  NAND3_X1 U5958 ( .A1(n5144), .A2(n5282), .A3(n5541), .ZN(n4972) );
  NAND3_X1 U5959 ( .A1(n4979), .A2(n5388), .A3(n5975), .ZN(n5390) );
  NAND2_X1 U5960 ( .A1(n5385), .A2(n5322), .ZN(n5388) );
  NAND2_X1 U5961 ( .A1(n5387), .A2(n5386), .ZN(n4979) );
  INV_X1 U5962 ( .A(n4985), .ZN(n7773) );
  NAND3_X1 U5963 ( .A1(n4991), .A2(n9373), .A3(n4989), .ZN(n9458) );
  NAND3_X1 U5964 ( .A1(n10527), .A2(n6519), .A3(n10539), .ZN(n7377) );
  NAND2_X1 U5965 ( .A1(n9137), .A2(n4995), .ZN(n9365) );
  NAND3_X1 U5966 ( .A1(n9364), .A2(n10511), .A3(n9365), .ZN(n9367) );
  NAND4_X1 U5967 ( .A1(n6032), .A2(n5186), .A3(n5197), .A4(n5187), .ZN(n6036)
         );
  NAND3_X1 U5968 ( .A1(n6032), .A2(n5186), .A3(n4861), .ZN(n6034) );
  NOR2_X2 U5969 ( .A1(n7819), .A2(n9446), .ZN(n7979) );
  AND3_X2 U5970 ( .A1(n8509), .A2(n8310), .A3(n8309), .ZN(n8315) );
  MUX2_X1 U5971 ( .A(n8268), .B(n8267), .S(n8319), .Z(n8279) );
  AOI21_X1 U5972 ( .B1(n8323), .B2(n8322), .A(n8321), .ZN(n8328) );
  NAND2_X1 U5973 ( .A1(n8448), .A2(n8447), .ZN(n8489) );
  NAND2_X1 U5974 ( .A1(n6903), .A2(n6902), .ZN(n8367) );
  INV_X1 U5975 ( .A(n8324), .ZN(n8331) );
  INV_X1 U5976 ( .A(n9352), .ZN(n10513) );
  OAI22_X1 U5977 ( .A1(n6562), .A2(n6540), .B1(n6542), .B2(n6683), .ZN(n5066)
         );
  AOI21_X2 U5978 ( .B1(P1_REG2_REG_14__SCAN_IN), .B2(n6939), .A(n6935), .ZN(
        n6055) );
  XNOR2_X2 U5979 ( .A(n5469), .B(P1_IR_REG_2__SCAN_IN), .ZN(n6269) );
  NAND2_X1 U5980 ( .A1(n8708), .A2(n8707), .ZN(n5151) );
  XNOR2_X1 U5981 ( .A(n8794), .B(n8754), .ZN(n5139) );
  NOR2_X1 U5982 ( .A1(n6564), .A2(n6541), .ZN(n5065) );
  NOR2_X4 U5983 ( .A1(n10510), .A2(n10529), .ZN(n10527) );
  NAND3_X1 U5984 ( .A1(n5337), .A2(n5336), .A3(n5335), .ZN(n5413) );
  NAND2_X1 U5985 ( .A1(n9821), .A2(n5010), .ZN(n5008) );
  NAND2_X2 U5986 ( .A1(n5850), .A2(n5851), .ZN(n5471) );
  INV_X1 U5987 ( .A(n5021), .ZN(n8519) );
  NAND2_X2 U5988 ( .A1(n5471), .A2(n6483), .ZN(n5474) );
  NAND3_X1 U5989 ( .A1(n7223), .A2(n7387), .A3(n5035), .ZN(n5034) );
  INV_X1 U5990 ( .A(n7223), .ZN(n7224) );
  NAND2_X1 U5991 ( .A1(n9193), .A2(n5042), .ZN(n5038) );
  NAND2_X1 U5992 ( .A1(n9193), .A2(n5040), .ZN(n5039) );
  AOI21_X1 U5993 ( .B1(n9193), .B2(n9124), .A(n5036), .ZN(n9180) );
  NAND2_X1 U5994 ( .A1(n9414), .A2(n5059), .ZN(n5058) );
  INV_X1 U5995 ( .A(n5062), .ZN(n9264) );
  NOR2_X1 U5996 ( .A1(n9117), .A2(n9118), .ZN(n5064) );
  NAND2_X1 U5997 ( .A1(n5995), .A2(n5068), .ZN(n5067) );
  NAND2_X1 U5998 ( .A1(n5995), .A2(n8473), .ZN(n5994) );
  OAI211_X1 U5999 ( .C1(n5995), .C2(n5072), .A(n5069), .B(n5067), .ZN(n8515)
         );
  NAND2_X1 U6000 ( .A1(n9978), .A2(n5074), .ZN(n5073) );
  NAND2_X1 U6001 ( .A1(n9978), .A2(n9984), .ZN(n5075) );
  NAND2_X1 U6002 ( .A1(n7688), .A2(n4870), .ZN(n7803) );
  NAND2_X1 U6003 ( .A1(n5089), .A2(n5087), .ZN(n5912) );
  NAND2_X1 U6004 ( .A1(n6918), .A2(n4871), .ZN(n6947) );
  OR2_X1 U6005 ( .A1(n10155), .A2(n10126), .ZN(n5096) );
  OAI21_X1 U6006 ( .B1(n9996), .B2(n5101), .A(n5098), .ZN(n9973) );
  OAI21_X1 U6007 ( .B1(n5539), .B2(n5106), .A(n5104), .ZN(n7086) );
  AND2_X1 U6008 ( .A1(n8342), .A2(n8463), .ZN(n5108) );
  NAND2_X1 U6009 ( .A1(n5863), .A2(n5111), .ZN(n5363) );
  NAND2_X1 U6010 ( .A1(n5863), .A2(n5109), .ZN(n5201) );
  NAND2_X1 U6011 ( .A1(n8457), .A2(n8456), .ZN(n6860) );
  NAND2_X1 U6012 ( .A1(n9882), .A2(n10519), .ZN(n8457) );
  INV_X1 U6013 ( .A(n6303), .ZN(n9882) );
  NAND2_X1 U6014 ( .A1(n5117), .A2(n5118), .ZN(n7038) );
  NAND3_X1 U6015 ( .A1(n6576), .A2(n6718), .A3(n7025), .ZN(n5117) );
  NAND2_X1 U6016 ( .A1(n8965), .A2(n5127), .ZN(n5121) );
  AOI21_X1 U6017 ( .B1(n8965), .B2(n4908), .A(n5122), .ZN(n8946) );
  OR2_X1 U6018 ( .A1(n8965), .A2(n8964), .ZN(n8962) );
  NAND2_X1 U6019 ( .A1(n7157), .A2(n5129), .ZN(n7414) );
  NAND2_X1 U6020 ( .A1(n7115), .A2(n7114), .ZN(n7157) );
  OAI21_X1 U6021 ( .B1(n7619), .B2(n5132), .A(n5130), .ZN(n7783) );
  OAI21_X1 U6022 ( .B1(n7619), .B2(n7618), .A(n7620), .ZN(n7707) );
  NAND2_X1 U6023 ( .A1(n6017), .A2(n5136), .ZN(n6272) );
  NAND2_X1 U6024 ( .A1(n6017), .A2(n5135), .ZN(n6238) );
  OAI21_X1 U6025 ( .B1(n5376), .B2(n5375), .A(n5326), .ZN(n5738) );
  NAND2_X1 U6026 ( .A1(n5674), .A2(n5306), .ZN(n5687) );
  NAND2_X1 U6027 ( .A1(n5167), .A2(n5258), .ZN(n5259) );
  MUX2_X1 U6028 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(P1_DATAO_REG_3__SCAN_IN), 
        .S(n6550), .Z(n5257) );
  NAND2_X1 U6029 ( .A1(n8040), .A2(n5168), .ZN(n6535) );
  AND2_X2 U6030 ( .A1(n6378), .A2(n5168), .ZN(n6556) );
  NAND2_X1 U6031 ( .A1(n7256), .A2(n5170), .ZN(n5169) );
  NAND2_X1 U6032 ( .A1(n5169), .A2(n8595), .ZN(n7372) );
  AOI21_X1 U6033 ( .B1(n9130), .B2(n8811), .A(n5183), .ZN(n8815) );
  AOI21_X1 U6034 ( .B1(n5182), .B2(n8814), .A(n4911), .ZN(n5179) );
  NAND2_X1 U6035 ( .A1(n8810), .A2(n8814), .ZN(n5180) );
  NAND2_X1 U6036 ( .A1(n8816), .A2(n9368), .ZN(n5181) );
  NAND2_X1 U6037 ( .A1(n5185), .A2(n5184), .ZN(n9175) );
  NOR2_X2 U6038 ( .A1(n5188), .A2(P2_IR_REG_7__SCAN_IN), .ZN(n5187) );
  NAND2_X1 U6039 ( .A1(n7654), .A2(n5195), .ZN(n5194) );
  NOR2_X2 U6040 ( .A1(n6012), .A2(P2_IR_REG_8__SCAN_IN), .ZN(n5197) );
  NAND2_X1 U6041 ( .A1(n6834), .A2(n4879), .ZN(n5204) );
  AND2_X1 U6042 ( .A1(n5209), .A2(n5208), .ZN(n9856) );
  NAND2_X1 U6043 ( .A1(n5209), .A2(n5207), .ZN(n9716) );
  NAND2_X1 U6044 ( .A1(n9802), .A2(n8124), .ZN(n8131) );
  NAND2_X1 U6045 ( .A1(n8825), .A2(n8755), .ZN(n10625) );
  NAND2_X1 U6046 ( .A1(n8977), .A2(n8856), .ZN(n8986) );
  OAI21_X1 U6047 ( .B1(n7059), .B2(n7058), .A(n7043), .ZN(n7104) );
  OAI21_X2 U6048 ( .B1(n7086), .B2(n8251), .A(n8379), .ZN(n7192) );
  OR2_X1 U6049 ( .A1(n6376), .A2(n6162), .ZN(n6373) );
  INV_X1 U6050 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n5513) );
  INV_X1 U6051 ( .A(n6554), .ZN(n8737) );
  OR2_X1 U6052 ( .A1(n5478), .A2(n10410), .ZN(n5448) );
  OR2_X1 U6053 ( .A1(n5455), .A2(n5454), .ZN(n5458) );
  OR2_X1 U6054 ( .A1(n5455), .A2(n6651), .ZN(n5433) );
  INV_X1 U6055 ( .A(n5455), .ZN(n5446) );
  OR2_X1 U6056 ( .A1(n9966), .A2(n5487), .ZN(n5786) );
  NAND2_X1 U6057 ( .A1(n6303), .A2(n8057), .ZN(n8456) );
  XNOR2_X1 U6058 ( .A(n6310), .B(n6311), .ZN(n9736) );
  NAND2_X1 U6059 ( .A1(n9725), .A2(n9729), .ZN(n9812) );
  OAI21_X1 U6060 ( .B1(n6592), .B2(n6593), .A(n6591), .ZN(n6638) );
  NOR2_X1 U6061 ( .A1(n5478), .A2(n5459), .ZN(n5460) );
  OAI22_X1 U6062 ( .A1(n6303), .A2(n8208), .B1(n10519), .B2(n6627), .ZN(n6304)
         );
  OR3_X1 U6063 ( .A1(P1_IR_REG_2__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .A3(
        P1_IR_REG_0__SCAN_IN), .ZN(n5225) );
  INV_X1 U6064 ( .A(n9963), .ZN(n9979) );
  AND2_X1 U6065 ( .A1(n8844), .A2(n8843), .ZN(n5226) );
  AND2_X1 U6066 ( .A1(n8657), .A2(n8784), .ZN(n5227) );
  INV_X1 U6067 ( .A(n10591), .ZN(n5984) );
  OR2_X1 U6068 ( .A1(n10171), .A2(n10088), .ZN(n5228) );
  AND2_X1 U6069 ( .A1(n6545), .A2(n6553), .ZN(n5229) );
  OR2_X1 U6070 ( .A1(n8326), .A2(n10246), .ZN(n5230) );
  NAND2_X1 U6071 ( .A1(n5476), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n5231) );
  NOR2_X1 U6072 ( .A1(n7407), .A2(n7409), .ZN(n5232) );
  AND2_X1 U6073 ( .A1(n7412), .A2(n7411), .ZN(n5233) );
  AND3_X1 U6074 ( .A1(n6559), .A2(n6558), .A3(n6557), .ZN(n5234) );
  NAND2_X1 U6075 ( .A1(n5579), .A2(n4880), .ZN(n5235) );
  NOR2_X1 U6076 ( .A1(n7409), .A2(n7408), .ZN(n5236) );
  NOR2_X1 U6077 ( .A1(n8848), .A2(n8914), .ZN(n5237) );
  OR2_X1 U6078 ( .A1(n10181), .A2(n10311), .ZN(n5239) );
  OR2_X1 U6079 ( .A1(n8524), .A2(n9717), .ZN(n5240) );
  NOR2_X1 U6080 ( .A1(n5969), .A2(n5968), .ZN(n5241) );
  AND2_X1 U6081 ( .A1(n5306), .A2(n5305), .ZN(n5242) );
  AND2_X1 U6082 ( .A1(n5260), .A2(n5259), .ZN(n5243) );
  NOR2_X1 U6083 ( .A1(n7913), .A2(n7912), .ZN(n5244) );
  INV_X1 U6084 ( .A(n6556), .ZN(n7303) );
  AND4_X1 U6085 ( .A1(n7932), .A2(n7931), .A3(n7930), .A4(n7929), .ZN(n8837)
         );
  AND2_X1 U6086 ( .A1(n8369), .A2(n6902), .ZN(n5245) );
  NOR2_X1 U6087 ( .A1(n8339), .A2(n5901), .ZN(n5246) );
  OR2_X1 U6088 ( .A1(n8668), .A2(n9119), .ZN(n8669) );
  INV_X1 U6089 ( .A(SI_9_), .ZN(n9507) );
  INV_X1 U6090 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n6007) );
  INV_X1 U6091 ( .A(n7626), .ZN(n6393) );
  INV_X1 U6092 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n6174) );
  OAI22_X1 U6093 ( .A1(n6879), .A2(n8208), .B1(n6621), .B2(n6627), .ZN(n6309)
         );
  INV_X1 U6094 ( .A(n8130), .ZN(n8128) );
  NOR2_X1 U6095 ( .A1(n6593), .A2(n6595), .ZN(n6596) );
  INV_X1 U6096 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n5340) );
  OR2_X1 U6097 ( .A1(n7287), .A2(n9879), .ZN(n5907) );
  OR2_X1 U6098 ( .A1(n6544), .A2(n6543), .ZN(n6545) );
  OR2_X1 U6099 ( .A1(n6607), .A2(n9689), .ZN(n8719) );
  INV_X1 U6100 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n6022) );
  INV_X1 U6101 ( .A(n5665), .ZN(n5354) );
  INV_X1 U6102 ( .A(n6212), .ZN(n6281) );
  INV_X1 U6103 ( .A(n9793), .ZN(n8115) );
  INV_X1 U6104 ( .A(n5420), .ZN(n5358) );
  AOI22_X1 U6105 ( .A1(n7334), .A2(n7333), .B1(n7332), .B2(n7331), .ZN(n7335)
         );
  INV_X1 U6106 ( .A(n5726), .ZN(n5357) );
  INV_X2 U6107 ( .A(n6627), .ZN(n8207) );
  INV_X1 U6108 ( .A(n5393), .ZN(n5359) );
  NAND2_X1 U6109 ( .A1(n5340), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5341) );
  OR2_X1 U6110 ( .A1(n5760), .A2(n5759), .ZN(n5779) );
  OR2_X1 U6111 ( .A1(n10015), .A2(n5935), .ZN(n5937) );
  OR2_X1 U6112 ( .A1(n10254), .A2(n7693), .ZN(n8408) );
  INV_X1 U6113 ( .A(n5550), .ZN(n5351) );
  AND2_X1 U6114 ( .A1(n5965), .A2(n5966), .ZN(n5970) );
  INV_X1 U6115 ( .A(SI_12_), .ZN(n9583) );
  INV_X1 U6116 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n6990) );
  INV_X1 U6117 ( .A(n9127), .ZN(n9128) );
  NAND2_X1 U6118 ( .A1(n5354), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n5680) );
  OR2_X1 U6119 ( .A1(n5599), .A2(n5598), .ZN(n5613) );
  INV_X1 U6120 ( .A(n8198), .ZN(n8199) );
  AND2_X1 U6121 ( .A1(n6215), .A2(n6214), .ZN(n6221) );
  OR2_X1 U6122 ( .A1(n5646), .A2(n5645), .ZN(n5665) );
  AND2_X1 U6123 ( .A1(n6302), .A2(n6301), .ZN(n8053) );
  NAND2_X1 U6124 ( .A1(n5778), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n5801) );
  NAND2_X1 U6125 ( .A1(n5359), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n5381) );
  NAND2_X1 U6126 ( .A1(n5485), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n5457) );
  AND2_X1 U6127 ( .A1(n6081), .A2(n6080), .ZN(n6942) );
  NAND2_X1 U6128 ( .A1(n5360), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n5747) );
  OR2_X1 U6129 ( .A1(n10155), .A2(n9795), .ZN(n8286) );
  OR2_X1 U6130 ( .A1(n5693), .A2(n5692), .ZN(n5726) );
  NAND2_X1 U6131 ( .A1(n5352), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n5599) );
  NAND2_X1 U6132 ( .A1(n5519), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n5523) );
  OR2_X1 U6133 ( .A1(n5688), .A2(P1_IR_REG_15__SCAN_IN), .ZN(n5689) );
  NAND2_X1 U6134 ( .A1(n5292), .A2(SI_12_), .ZN(n5295) );
  INV_X1 U6135 ( .A(SI_10_), .ZN(n9624) );
  NOR2_X1 U6136 ( .A1(n5545), .A2(P1_IR_REG_6__SCAN_IN), .ZN(n5563) );
  NAND2_X1 U6137 ( .A1(n6237), .A2(n6018), .ZN(n6019) );
  NOR2_X1 U6138 ( .A1(n5236), .A2(n5233), .ZN(n7413) );
  NOR2_X1 U6139 ( .A1(n5226), .A2(n5237), .ZN(n8849) );
  NAND2_X1 U6140 ( .A1(n8986), .A2(n8870), .ZN(n8987) );
  INV_X1 U6141 ( .A(n9037), .ZN(n7220) );
  INV_X1 U6142 ( .A(n9005), .ZN(n9011) );
  AND2_X1 U6143 ( .A1(n6478), .A2(n8829), .ZN(n6669) );
  INV_X1 U6144 ( .A(n9163), .ZN(n9186) );
  INV_X1 U6145 ( .A(n9239), .ZN(n9249) );
  NAND2_X1 U6146 ( .A1(n7939), .A2(n8837), .ZN(n8015) );
  OR2_X1 U6147 ( .A1(n7919), .A2(n7918), .ZN(n7920) );
  OR2_X1 U6148 ( .A1(n7569), .A2(n8770), .ZN(n7642) );
  AND2_X1 U6149 ( .A1(n8599), .A2(n8598), .ZN(n8764) );
  INV_X1 U6150 ( .A(n9307), .ZN(n9223) );
  INV_X1 U6151 ( .A(n8777), .ZN(n7892) );
  AND2_X1 U6152 ( .A1(n8823), .A2(n8754), .ZN(n9253) );
  NOR2_X1 U6153 ( .A1(n8217), .A2(n9853), .ZN(n8218) );
  NAND2_X1 U6154 ( .A1(n6287), .A2(n6286), .ZN(n6297) );
  OR2_X1 U6155 ( .A1(n7923), .A2(n5474), .ZN(n5723) );
  OR2_X1 U6156 ( .A1(n6325), .A2(n10405), .ZN(n6222) );
  AND2_X1 U6157 ( .A1(n5951), .A2(n5817), .ZN(n8522) );
  INV_X1 U6158 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n7147) );
  OR2_X1 U6159 ( .A1(n6077), .A2(n8085), .ZN(n8091) );
  AND2_X1 U6160 ( .A1(n8389), .A2(n10063), .ZN(n10099) );
  OR2_X1 U6161 ( .A1(n10591), .A2(n9951), .ZN(n5988) );
  OR2_X1 U6162 ( .A1(n5471), .A2(n5470), .ZN(n5472) );
  INV_X1 U6163 ( .A(n10164), .ZN(n5983) );
  OR2_X1 U6164 ( .A1(n7905), .A2(n5474), .ZN(n5711) );
  INV_X1 U6165 ( .A(n6600), .ZN(n6664) );
  AND2_X1 U6166 ( .A1(n5313), .A2(n5312), .ZN(n5716) );
  AND2_X1 U6167 ( .A1(n5295), .A2(n5294), .ZN(n5619) );
  AND2_X1 U6168 ( .A1(n5269), .A2(n5268), .ZN(n5531) );
  NAND2_X1 U6169 ( .A1(n6019), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6039) );
  INV_X1 U6170 ( .A(n8942), .ZN(n8943) );
  INV_X1 U6171 ( .A(n10565), .ZN(n7381) );
  AND3_X1 U6172 ( .A1(n8539), .A2(n8538), .A3(n8537), .ZN(n8812) );
  AND3_X1 U6173 ( .A1(n8008), .A2(n8007), .A3(n8006), .ZN(n9118) );
  INV_X1 U6174 ( .A(n10493), .ZN(n10467) );
  INV_X1 U6175 ( .A(n10468), .ZN(n10495) );
  INV_X1 U6176 ( .A(n9153), .ZN(n9147) );
  INV_X1 U6177 ( .A(n9124), .ZN(n9202) );
  AND2_X1 U6178 ( .A1(n8574), .A2(n8575), .ZN(n8784) );
  AND2_X1 U6179 ( .A1(n7642), .A2(n7641), .ZN(n7762) );
  INV_X1 U6180 ( .A(n9350), .ZN(n9304) );
  INV_X1 U6181 ( .A(n9253), .ZN(n9340) );
  INV_X1 U6182 ( .A(n9354), .ZN(n9307) );
  NOR2_X1 U6183 ( .A1(n10465), .A2(n6472), .ZN(n7079) );
  INV_X1 U6184 ( .A(n10639), .ZN(n10556) );
  AND2_X1 U6185 ( .A1(n6475), .A2(n6509), .ZN(n10619) );
  NAND2_X1 U6186 ( .A1(n9302), .A2(n7591), .ZN(n10639) );
  AND2_X1 U6187 ( .A1(n6229), .A2(n10464), .ZN(n10362) );
  INV_X1 U6188 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n6024) );
  INV_X1 U6189 ( .A(n9846), .ZN(n9863) );
  INV_X1 U6190 ( .A(n10425), .ZN(n10457) );
  INV_X1 U6191 ( .A(n9952), .ZN(n10459) );
  AND2_X1 U6192 ( .A1(n5850), .A2(n8325), .ZN(n10141) );
  INV_X1 U6193 ( .A(n6894), .ZN(n8244) );
  AND2_X1 U6194 ( .A1(n5885), .A2(n10318), .ZN(n6198) );
  OR2_X1 U6195 ( .A1(n6282), .A2(n10603), .ZN(n10595) );
  AND2_X1 U6196 ( .A1(n10403), .A2(n5990), .ZN(n5999) );
  INV_X1 U6197 ( .A(n5880), .ZN(n10317) );
  AND2_X1 U6198 ( .A1(n7005), .A2(P1_STATE_REG_SCAN_IN), .ZN(n5892) );
  AND2_X1 U6199 ( .A1(n5709), .A2(n5720), .ZN(n7759) );
  AND2_X1 U6200 ( .A1(n5627), .A2(n5640), .ZN(n6368) );
  AND2_X1 U6201 ( .A1(n5567), .A2(n5580), .ZN(n9922) );
  INV_X1 U6202 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n7493) );
  NOR2_X1 U6203 ( .A1(n10377), .A2(n7501), .ZN(n7502) );
  NOR2_X1 U6204 ( .A1(n10388), .A2(n10387), .ZN(n7519) );
  XNOR2_X1 U6205 ( .A(n6039), .B(P2_IR_REG_23__SCAN_IN), .ZN(n6230) );
  INV_X1 U6206 ( .A(n8949), .ZN(n9013) );
  INV_X1 U6207 ( .A(n8947), .ZN(n9014) );
  INV_X1 U6208 ( .A(n8941), .ZN(n9019) );
  INV_X1 U6209 ( .A(P2_U3966), .ZN(n9022) );
  NAND3_X1 U6210 ( .A1(n6708), .A2(n6707), .A3(n9107), .ZN(n10487) );
  INV_X1 U6211 ( .A(n9106), .ZN(n9360) );
  AND2_X1 U6212 ( .A1(n9293), .A2(n9292), .ZN(n9435) );
  AND2_X1 U6213 ( .A1(n7217), .A2(n9304), .ZN(n9354) );
  NAND2_X1 U6214 ( .A1(n9307), .A2(n7213), .ZN(n9285) );
  INV_X1 U6215 ( .A(n10642), .ZN(n10641) );
  AND2_X2 U6216 ( .A1(n7080), .A2(n7079), .ZN(n10642) );
  INV_X1 U6217 ( .A(n10646), .ZN(n10643) );
  NAND2_X1 U6218 ( .A1(n10362), .A2(n10361), .ZN(n10462) );
  INV_X1 U6219 ( .A(n6510), .ZN(n6980) );
  INV_X1 U6220 ( .A(n6273), .ZN(n8230) );
  NAND2_X1 U6221 ( .A1(n8489), .A2(n8488), .ZN(n8500) );
  NAND2_X1 U6222 ( .A1(n5786), .A2(n5785), .ZN(n9988) );
  OR2_X1 U6223 ( .A1(P1_U3083), .A2(n6094), .ZN(n10425) );
  INV_X1 U6224 ( .A(n10097), .ZN(n10152) );
  AND2_X1 U6225 ( .A1(n7607), .A2(n7606), .ZN(n10260) );
  NAND2_X1 U6226 ( .A1(n5999), .A2(n6198), .ZN(n10607) );
  INV_X1 U6227 ( .A(n10155), .ZN(n10306) );
  NAND2_X1 U6228 ( .A1(n5999), .A2(n5998), .ZN(n10609) );
  NOR2_X1 U6229 ( .A1(n10317), .A2(n10405), .ZN(n10345) );
  NAND2_X1 U6230 ( .A1(n6322), .A2(n5892), .ZN(n10405) );
  NOR2_X1 U6231 ( .A1(n7520), .A2(n7519), .ZN(n10390) );
  NOR2_X2 U6232 ( .A1(n6478), .A2(n6230), .ZN(P2_U3966) );
  INV_X1 U6233 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n5247) );
  INV_X1 U6234 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n5248) );
  NAND2_X1 U6235 ( .A1(n5251), .A2(SI_1_), .ZN(n5463) );
  INV_X1 U6236 ( .A(n5251), .ZN(n5252) );
  INV_X1 U6237 ( .A(SI_1_), .ZN(n9638) );
  NAND2_X1 U6238 ( .A1(n5252), .A2(n9638), .ZN(n5253) );
  AND2_X1 U6239 ( .A1(n5463), .A2(n5253), .ZN(n5436) );
  MUX2_X1 U6240 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .S(n5270), .Z(n5437) );
  NAND2_X1 U6241 ( .A1(n5436), .A2(n5437), .ZN(n5464) );
  NAND2_X1 U6242 ( .A1(n5464), .A2(n5463), .ZN(n5255) );
  NAND2_X1 U6243 ( .A1(n5257), .A2(SI_3_), .ZN(n5260) );
  INV_X1 U6244 ( .A(SI_3_), .ZN(n5258) );
  MUX2_X1 U6245 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(P2_DATAO_REG_4__SCAN_IN), 
        .S(n6110), .Z(n5261) );
  NAND2_X1 U6246 ( .A1(n5261), .A2(SI_4_), .ZN(n5265) );
  INV_X1 U6247 ( .A(n5261), .ZN(n5263) );
  INV_X1 U6248 ( .A(SI_4_), .ZN(n5262) );
  NAND2_X1 U6249 ( .A1(n5263), .A2(n5262), .ZN(n5264) );
  NAND2_X1 U6250 ( .A1(n5493), .A2(n5492), .ZN(n5495) );
  NAND2_X1 U6251 ( .A1(n5495), .A2(n5265), .ZN(n5532) );
  MUX2_X1 U6252 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(P2_DATAO_REG_5__SCAN_IN), 
        .S(n6110), .Z(n5266) );
  NAND2_X1 U6253 ( .A1(n5266), .A2(SI_5_), .ZN(n5269) );
  INV_X1 U6254 ( .A(n5266), .ZN(n5267) );
  INV_X1 U6255 ( .A(SI_5_), .ZN(n9627) );
  NAND2_X1 U6256 ( .A1(n5267), .A2(n9627), .ZN(n5268) );
  NAND2_X1 U6257 ( .A1(n5532), .A2(n5531), .ZN(n5534) );
  NAND2_X1 U6258 ( .A1(n5534), .A2(n5269), .ZN(n5541) );
  MUX2_X1 U6259 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(P2_DATAO_REG_8__SCAN_IN), 
        .S(n5270), .Z(n5271) );
  NAND2_X1 U6260 ( .A1(n5271), .A2(SI_8_), .ZN(n5274) );
  INV_X1 U6261 ( .A(n5274), .ZN(n5273) );
  OAI21_X1 U6262 ( .B1(n5271), .B2(SI_8_), .A(n5274), .ZN(n5560) );
  INV_X1 U6263 ( .A(n5560), .ZN(n5272) );
  INV_X1 U6264 ( .A(n5279), .ZN(n5276) );
  AND2_X1 U6265 ( .A1(n5558), .A2(n5274), .ZN(n5275) );
  MUX2_X1 U6266 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(P2_DATAO_REG_9__SCAN_IN), 
        .S(n6110), .Z(n5277) );
  INV_X1 U6267 ( .A(n5277), .ZN(n5278) );
  NAND2_X1 U6268 ( .A1(n5278), .A2(n9507), .ZN(n5280) );
  INV_X1 U6269 ( .A(n5544), .ZN(n5557) );
  MUX2_X1 U6270 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .S(n6110), .Z(n5281) );
  NAND2_X1 U6271 ( .A1(n5281), .A2(SI_6_), .ZN(n5542) );
  OAI21_X1 U6272 ( .B1(n5281), .B2(SI_6_), .A(n5542), .ZN(n5511) );
  INV_X1 U6273 ( .A(n5511), .ZN(n5540) );
  MUX2_X1 U6274 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(P2_DATAO_REG_10__SCAN_IN), 
        .S(n6483), .Z(n5286) );
  MUX2_X1 U6275 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(P2_DATAO_REG_11__SCAN_IN), 
        .S(n6110), .Z(n5287) );
  NAND2_X1 U6276 ( .A1(n5287), .A2(SI_11_), .ZN(n5291) );
  INV_X1 U6277 ( .A(n5287), .ZN(n5288) );
  NAND2_X1 U6278 ( .A1(n5288), .A2(n9584), .ZN(n5289) );
  NAND2_X1 U6279 ( .A1(n5291), .A2(n5289), .ZN(n5605) );
  INV_X1 U6280 ( .A(n5605), .ZN(n5290) );
  MUX2_X1 U6281 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(P2_DATAO_REG_12__SCAN_IN), 
        .S(n6110), .Z(n5292) );
  INV_X1 U6282 ( .A(n5292), .ZN(n5293) );
  NAND2_X1 U6283 ( .A1(n5293), .A2(n9583), .ZN(n5294) );
  MUX2_X1 U6284 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(P2_DATAO_REG_13__SCAN_IN), 
        .S(n6110), .Z(n5298) );
  MUX2_X1 U6285 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(P2_DATAO_REG_14__SCAN_IN), 
        .S(n6110), .Z(n5297) );
  NAND2_X1 U6286 ( .A1(n5297), .A2(SI_14_), .ZN(n5302) );
  OAI21_X1 U6287 ( .B1(n5297), .B2(SI_14_), .A(n5302), .ZN(n5655) );
  INV_X1 U6288 ( .A(n5655), .ZN(n5300) );
  INV_X1 U6289 ( .A(n5298), .ZN(n5299) );
  INV_X1 U6290 ( .A(SI_13_), .ZN(n9475) );
  NAND2_X1 U6291 ( .A1(n5299), .A2(n9475), .ZN(n5653) );
  NAND2_X1 U6292 ( .A1(n5658), .A2(n5302), .ZN(n5672) );
  MUX2_X1 U6293 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(P2_DATAO_REG_15__SCAN_IN), 
        .S(n6110), .Z(n5303) );
  NAND2_X1 U6294 ( .A1(n5303), .A2(SI_15_), .ZN(n5306) );
  INV_X1 U6295 ( .A(n5303), .ZN(n5304) );
  INV_X1 U6296 ( .A(SI_15_), .ZN(n9586) );
  NAND2_X1 U6297 ( .A1(n5304), .A2(n9586), .ZN(n5305) );
  NAND2_X1 U6298 ( .A1(n5672), .A2(n5242), .ZN(n5674) );
  MUX2_X1 U6299 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(P2_DATAO_REG_16__SCAN_IN), 
        .S(n6110), .Z(n5307) );
  MUX2_X1 U6300 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(P2_DATAO_REG_17__SCAN_IN), 
        .S(n6483), .Z(n5308) );
  NAND2_X1 U6301 ( .A1(n5308), .A2(SI_17_), .ZN(n5309) );
  OAI21_X1 U6302 ( .B1(n5308), .B2(SI_17_), .A(n5309), .ZN(n5700) );
  MUX2_X1 U6303 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .S(n6483), .Z(n5310) );
  NAND2_X1 U6304 ( .A1(n5310), .A2(SI_18_), .ZN(n5313) );
  INV_X1 U6305 ( .A(n5310), .ZN(n5311) );
  INV_X1 U6306 ( .A(SI_18_), .ZN(n9612) );
  NAND2_X1 U6307 ( .A1(n5311), .A2(n9612), .ZN(n5312) );
  MUX2_X1 U6308 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(P2_DATAO_REG_19__SCAN_IN), 
        .S(n6483), .Z(n5314) );
  XNOR2_X1 U6309 ( .A(n5314), .B(SI_19_), .ZN(n5411) );
  INV_X1 U6310 ( .A(n5314), .ZN(n5315) );
  INV_X1 U6311 ( .A(SI_19_), .ZN(n9493) );
  NAND2_X1 U6312 ( .A1(n5315), .A2(n9493), .ZN(n5316) );
  MUX2_X1 U6313 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(P2_DATAO_REG_20__SCAN_IN), 
        .S(n6483), .Z(n5317) );
  INV_X1 U6314 ( .A(SI_20_), .ZN(n9477) );
  XNOR2_X1 U6315 ( .A(n5317), .B(n9477), .ZN(n5397) );
  NOR2_X1 U6316 ( .A1(n5317), .A2(SI_20_), .ZN(n5318) );
  MUX2_X1 U6317 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(P2_DATAO_REG_21__SCAN_IN), 
        .S(n6110), .Z(n5319) );
  NAND2_X1 U6318 ( .A1(n5319), .A2(SI_21_), .ZN(n5323) );
  INV_X1 U6319 ( .A(n5319), .ZN(n5320) );
  INV_X1 U6320 ( .A(SI_21_), .ZN(n9588) );
  NAND2_X1 U6321 ( .A1(n5320), .A2(n9588), .ZN(n5321) );
  NAND2_X1 U6322 ( .A1(n5323), .A2(n5321), .ZN(n5386) );
  INV_X1 U6323 ( .A(n5386), .ZN(n5322) );
  MUX2_X1 U6324 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(P2_DATAO_REG_22__SCAN_IN), 
        .S(n6483), .Z(n5324) );
  XNOR2_X1 U6325 ( .A(n5324), .B(SI_22_), .ZN(n5375) );
  INV_X1 U6326 ( .A(n5324), .ZN(n5325) );
  INV_X1 U6327 ( .A(SI_22_), .ZN(n9593) );
  NAND2_X1 U6328 ( .A1(n5325), .A2(n9593), .ZN(n5326) );
  MUX2_X1 U6329 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(P2_DATAO_REG_23__SCAN_IN), 
        .S(n6483), .Z(n5739) );
  XNOR2_X1 U6330 ( .A(n5739), .B(n9590), .ZN(n5737) );
  XNOR2_X1 U6331 ( .A(n5738), .B(n5737), .ZN(n8681) );
  NAND2_X1 U6332 ( .A1(n5442), .A2(n5327), .ZN(n5515) );
  INV_X1 U6333 ( .A(n5515), .ZN(n5337) );
  NOR2_X1 U6334 ( .A1(P1_IR_REG_17__SCAN_IN), .A2(P1_IR_REG_12__SCAN_IN), .ZN(
        n5331) );
  NOR2_X1 U6335 ( .A1(P1_IR_REG_16__SCAN_IN), .A2(P1_IR_REG_13__SCAN_IN), .ZN(
        n5334) );
  OAI21_X1 U6336 ( .B1(n5339), .B2(n10319), .A(P1_IR_REG_28__SCAN_IN), .ZN(
        n5342) );
  NAND2_X1 U6337 ( .A1(n8681), .A2(n5975), .ZN(n5349) );
  NAND2_X1 U6338 ( .A1(n5775), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n5348) );
  INV_X1 U6339 ( .A(n5523), .ZN(n5350) );
  INV_X1 U6340 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n5645) );
  INV_X1 U6341 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n5692) );
  AND2_X1 U6342 ( .A1(P1_REG3_REG_18__SCAN_IN), .A2(P1_REG3_REG_17__SCAN_IN), 
        .ZN(n5356) );
  INV_X1 U6343 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n5418) );
  INV_X1 U6344 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n5391) );
  INV_X1 U6345 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n5361) );
  NAND2_X1 U6346 ( .A1(n5381), .A2(n5361), .ZN(n5362) );
  NAND2_X1 U6347 ( .A1(n5747), .A2(n5362), .ZN(n10018) );
  INV_X1 U6348 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n5366) );
  XNOR2_X2 U6349 ( .A(n5367), .B(P1_IR_REG_29__SCAN_IN), .ZN(n5368) );
  OR2_X1 U6350 ( .A1(n10018), .A2(n5487), .ZN(n5374) );
  INV_X1 U6351 ( .A(P1_REG0_REG_23__SCAN_IN), .ZN(n10289) );
  NAND2_X2 U6352 ( .A1(n8025), .A2(n5369), .ZN(n5456) );
  NAND2_X1 U6353 ( .A1(n5476), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n5371) );
  NAND2_X2 U6354 ( .A1(n5369), .A2(n5368), .ZN(n5478) );
  NAND2_X1 U6355 ( .A1(n5830), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n5370) );
  OAI211_X1 U6356 ( .C1(n10289), .C2(n5456), .A(n5371), .B(n5370), .ZN(n5372)
         );
  INV_X1 U6357 ( .A(n5372), .ZN(n5373) );
  NAND2_X1 U6358 ( .A1(n5374), .A2(n5373), .ZN(n10043) );
  XNOR2_X1 U6359 ( .A(n10197), .B(n10043), .ZN(n10024) );
  NAND2_X1 U6360 ( .A1(n8671), .A2(n5975), .ZN(n5378) );
  NAND2_X1 U6361 ( .A1(n5775), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n5377) );
  INV_X1 U6362 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n5384) );
  INV_X1 U6363 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n5379) );
  NAND2_X1 U6364 ( .A1(n5393), .A2(n5379), .ZN(n5380) );
  NAND2_X1 U6365 ( .A1(n5381), .A2(n5380), .ZN(n10049) );
  OR2_X1 U6366 ( .A1(n10049), .A2(n5487), .ZN(n5383) );
  AOI22_X1 U6367 ( .A1(n5978), .A2(P1_REG0_REG_22__SCAN_IN), .B1(n5476), .B2(
        P1_REG2_REG_22__SCAN_IN), .ZN(n5382) );
  OAI211_X1 U6368 ( .C1(n5478), .C2(n5384), .A(n5383), .B(n5382), .ZN(n10071)
         );
  INV_X1 U6369 ( .A(n10071), .ZN(n5429) );
  OR2_X1 U6370 ( .A1(n10205), .A2(n5429), .ZN(n8396) );
  INV_X1 U6371 ( .A(n8396), .ZN(n5430) );
  INV_X1 U6372 ( .A(n5385), .ZN(n5387) );
  NAND2_X1 U6373 ( .A1(n5775), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n5389) );
  NAND2_X1 U6374 ( .A1(n5403), .A2(n5391), .ZN(n5392) );
  AND2_X1 U6375 ( .A1(n5393), .A2(n5392), .ZN(n10076) );
  NAND2_X1 U6376 ( .A1(n10076), .A2(n5446), .ZN(n5396) );
  AOI22_X1 U6377 ( .A1(n5978), .A2(P1_REG0_REG_21__SCAN_IN), .B1(n5476), .B2(
        P1_REG2_REG_21__SCAN_IN), .ZN(n5395) );
  NAND2_X1 U6378 ( .A1(n5830), .A2(P1_REG1_REG_21__SCAN_IN), .ZN(n5394) );
  XNOR2_X1 U6379 ( .A(n5398), .B(n5397), .ZN(n8000) );
  NAND2_X1 U6380 ( .A1(n8000), .A2(n5975), .ZN(n5400) );
  NAND2_X1 U6381 ( .A1(n5775), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n5399) );
  INV_X1 U6382 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n5401) );
  NAND2_X1 U6383 ( .A1(n5420), .A2(n5401), .ZN(n5402) );
  NAND2_X1 U6384 ( .A1(n5403), .A2(n5402), .ZN(n10086) );
  OR2_X1 U6385 ( .A1(n10086), .A2(n5487), .ZN(n5408) );
  NAND2_X1 U6386 ( .A1(n5978), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n5405) );
  NAND2_X1 U6387 ( .A1(n5476), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n5404) );
  AND2_X1 U6388 ( .A1(n5405), .A2(n5404), .ZN(n5407) );
  NAND2_X1 U6389 ( .A1(n5830), .A2(P1_REG1_REG_20__SCAN_IN), .ZN(n5406) );
  OR2_X1 U6390 ( .A1(n10213), .A2(n10104), .ZN(n10065) );
  AND2_X1 U6391 ( .A1(n5922), .A2(n10065), .ZN(n8391) );
  NAND2_X1 U6392 ( .A1(n10075), .A2(n8155), .ZN(n5921) );
  INV_X1 U6393 ( .A(n5921), .ZN(n5409) );
  OR2_X1 U6394 ( .A1(n8391), .A2(n5409), .ZN(n8293) );
  INV_X1 U6395 ( .A(n8293), .ZN(n5428) );
  NAND2_X1 U6396 ( .A1(n10213), .A2(n10104), .ZN(n5924) );
  INV_X1 U6397 ( .A(n5924), .ZN(n10066) );
  NAND2_X1 U6398 ( .A1(n5922), .A2(n10066), .ZN(n5410) );
  AND2_X1 U6399 ( .A1(n5410), .A2(n5921), .ZN(n8393) );
  XNOR2_X1 U6400 ( .A(n5412), .B(n5411), .ZN(n7995) );
  NAND2_X1 U6401 ( .A1(n7995), .A2(n5975), .ZN(n5417) );
  NAND2_X1 U6402 ( .A1(n5413), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5415) );
  INV_X1 U6403 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n5414) );
  AOI22_X1 U6404 ( .A1(n5775), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n10019), 
        .B2(n10408), .ZN(n5416) );
  NAND2_X1 U6405 ( .A1(n5728), .A2(n5418), .ZN(n5419) );
  AND2_X1 U6406 ( .A1(n5420), .A2(n5419), .ZN(n10112) );
  NAND2_X1 U6407 ( .A1(n10112), .A2(n5446), .ZN(n5426) );
  NAND2_X1 U6408 ( .A1(n5978), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n5425) );
  INV_X1 U6409 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n5422) );
  OR2_X1 U6410 ( .A1(n5421), .A2(n5422), .ZN(n5424) );
  NAND2_X1 U6411 ( .A1(n5830), .A2(P1_REG1_REG_19__SCAN_IN), .ZN(n5423) );
  NAND4_X1 U6412 ( .A1(n5426), .A2(n5425), .A3(n5424), .A4(n5423), .ZN(n10125)
         );
  INV_X1 U6413 ( .A(n10125), .ZN(n9845) );
  NAND2_X1 U6414 ( .A1(n10109), .A2(n9845), .ZN(n10063) );
  AND2_X1 U6415 ( .A1(n8393), .A2(n10063), .ZN(n5427) );
  OR2_X1 U6416 ( .A1(n5428), .A2(n5427), .ZN(n10037) );
  NAND2_X1 U6417 ( .A1(n10205), .A2(n5429), .ZN(n8392) );
  NAND2_X1 U6418 ( .A1(n8396), .A2(n8392), .ZN(n10033) );
  INV_X1 U6419 ( .A(n10033), .ZN(n10041) );
  AND2_X1 U6420 ( .A1(n10037), .A2(n10041), .ZN(n10038) );
  OR2_X1 U6421 ( .A1(n5430), .A2(n10038), .ZN(n10021) );
  AND2_X1 U6422 ( .A1(n10024), .A2(n10021), .ZN(n5736) );
  NAND2_X1 U6423 ( .A1(n5476), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n5435) );
  INV_X1 U6424 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n6350) );
  OR2_X1 U6425 ( .A1(n5478), .A2(n6350), .ZN(n5434) );
  INV_X1 U6426 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n6651) );
  INV_X1 U6427 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n5431) );
  NAND4_X2 U6428 ( .A1(n5435), .A2(n5434), .A3(n5433), .A4(n5432), .ZN(n6277)
         );
  INV_X1 U6429 ( .A(n5436), .ZN(n5439) );
  INV_X1 U6430 ( .A(n5437), .ZN(n5438) );
  NAND2_X1 U6431 ( .A1(n5439), .A2(n5438), .ZN(n5440) );
  NAND2_X1 U6432 ( .A1(n5464), .A2(n5440), .ZN(n6541) );
  NAND2_X1 U6433 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5441) );
  MUX2_X1 U6434 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5441), .S(
        P1_IR_REG_1__SCAN_IN), .Z(n5444) );
  INV_X1 U6435 ( .A(n5442), .ZN(n5443) );
  NAND2_X1 U6436 ( .A1(n5444), .A2(n5443), .ZN(n6114) );
  XNOR2_X2 U6437 ( .A(n6277), .B(n6347), .ZN(n5895) );
  INV_X1 U6438 ( .A(n5895), .ZN(n6345) );
  INV_X1 U6439 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n10410) );
  NAND2_X1 U6440 ( .A1(n5476), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n5447) );
  NAND2_X1 U6441 ( .A1(n6483), .A2(SI_0_), .ZN(n5451) );
  XNOR2_X1 U6442 ( .A(n5451), .B(P2_DATAO_REG_0__SCAN_IN), .ZN(n10327) );
  MUX2_X1 U6443 ( .A(P1_IR_REG_0__SCAN_IN), .B(n10327), .S(n5471), .Z(n6453)
         );
  INV_X1 U6444 ( .A(n6453), .ZN(n6348) );
  NAND2_X1 U6445 ( .A1(n6345), .A2(n6344), .ZN(n5453) );
  INV_X1 U6446 ( .A(n6277), .ZN(n6861) );
  INV_X1 U6447 ( .A(n6347), .ZN(n6278) );
  NAND2_X1 U6448 ( .A1(n6861), .A2(n6278), .ZN(n5452) );
  NAND2_X1 U6449 ( .A1(n5453), .A2(n5452), .ZN(n8460) );
  INV_X1 U6450 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n5454) );
  AND2_X1 U6451 ( .A1(n5458), .A2(n5457), .ZN(n5462) );
  INV_X1 U6452 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n5459) );
  AOI21_X1 U6453 ( .B1(P1_REG2_REG_2__SCAN_IN), .B2(n5476), .A(n5460), .ZN(
        n5461) );
  AND2_X1 U6454 ( .A1(n5464), .A2(n5463), .ZN(n5466) );
  NAND2_X1 U6455 ( .A1(n5466), .A2(n5465), .ZN(n5468) );
  NAND2_X1 U6456 ( .A1(n5468), .A2(n5467), .ZN(n6563) );
  NAND2_X1 U6457 ( .A1(n4858), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n5473) );
  OR2_X1 U6458 ( .A1(n5442), .A2(n10319), .ZN(n5469) );
  INV_X1 U6459 ( .A(n6269), .ZN(n5470) );
  OAI211_X2 U6460 ( .C1(n5474), .C2(n6563), .A(n5473), .B(n5472), .ZN(n8057)
         );
  INV_X1 U6461 ( .A(n6860), .ZN(n8338) );
  NAND2_X1 U6462 ( .A1(n8460), .A2(n8338), .ZN(n5475) );
  NAND2_X1 U6463 ( .A1(n5485), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n5480) );
  INV_X1 U6464 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n5477) );
  OR2_X1 U6465 ( .A1(n5478), .A2(n5477), .ZN(n5479) );
  XNOR2_X1 U6466 ( .A(n5481), .B(n5243), .ZN(n6527) );
  NAND2_X1 U6467 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(n5225), .ZN(n5482) );
  XNOR2_X1 U6468 ( .A(n5482), .B(P1_IR_REG_3__SCAN_IN), .ZN(n6105) );
  NAND2_X1 U6469 ( .A1(n10408), .A2(n6105), .ZN(n5483) );
  INV_X1 U6470 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n6884) );
  NAND2_X1 U6471 ( .A1(n5485), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n5490) );
  INV_X1 U6472 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n5486) );
  OR2_X1 U6473 ( .A1(n5478), .A2(n5486), .ZN(n5489) );
  XNOR2_X1 U6474 ( .A(P1_REG3_REG_3__SCAN_IN), .B(P1_REG3_REG_4__SCAN_IN), 
        .ZN(n6883) );
  OR2_X1 U6475 ( .A1(n5487), .A2(n6883), .ZN(n5488) );
  OR2_X1 U6476 ( .A1(n5493), .A2(n5492), .ZN(n5494) );
  NAND2_X1 U6477 ( .A1(n5495), .A2(n5494), .ZN(n6516) );
  INV_X1 U6478 ( .A(n6516), .ZN(n5496) );
  NAND2_X1 U6479 ( .A1(n5975), .A2(n5496), .ZN(n5501) );
  NAND2_X1 U6480 ( .A1(n5775), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n5500) );
  NAND2_X1 U6481 ( .A1(n5515), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5497) );
  NAND2_X1 U6482 ( .A1(n5497), .A2(n5513), .ZN(n5529) );
  OR2_X1 U6483 ( .A1(n5497), .A2(n5513), .ZN(n5498) );
  NAND2_X1 U6484 ( .A1(n10408), .A2(n9895), .ZN(n5499) );
  NAND2_X1 U6485 ( .A1(n9881), .A2(n10549), .ZN(n5502) );
  AND2_X1 U6486 ( .A1(n6875), .A2(n5502), .ZN(n8458) );
  NAND2_X1 U6487 ( .A1(n6877), .A2(n8458), .ZN(n5504) );
  NAND2_X1 U6488 ( .A1(n6879), .A2(n9740), .ZN(n5898) );
  INV_X1 U6489 ( .A(n5898), .ZN(n6876) );
  NOR2_X1 U6490 ( .A1(n9881), .A2(n10549), .ZN(n5503) );
  AOI21_X1 U6491 ( .B1(n8458), .B2(n6876), .A(n5503), .ZN(n8461) );
  INV_X1 U6492 ( .A(n6901), .ZN(n5537) );
  NAND2_X1 U6493 ( .A1(n5978), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n5510) );
  INV_X1 U6494 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n6909) );
  OR2_X1 U6495 ( .A1(n5421), .A2(n6909), .ZN(n5509) );
  INV_X1 U6496 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n6643) );
  NAND2_X1 U6497 ( .A1(n5523), .A2(n6643), .ZN(n5505) );
  NAND2_X1 U6498 ( .A1(n5550), .A2(n5505), .ZN(n6908) );
  OR2_X1 U6499 ( .A1(n5487), .A2(n6908), .ZN(n5508) );
  INV_X1 U6500 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n5506) );
  OR2_X1 U6501 ( .A1(n5478), .A2(n5506), .ZN(n5507) );
  XNOR2_X1 U6502 ( .A(n5541), .B(n5511), .ZN(n6966) );
  NAND2_X1 U6503 ( .A1(n6966), .A2(n5975), .ZN(n5518) );
  NAND2_X1 U6504 ( .A1(n5513), .A2(n5512), .ZN(n5514) );
  OR2_X1 U6505 ( .A1(n5515), .A2(n5514), .ZN(n5545) );
  NAND2_X1 U6506 ( .A1(n5545), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5516) );
  XNOR2_X1 U6507 ( .A(n5516), .B(P1_IR_REG_6__SCAN_IN), .ZN(n10431) );
  AOI22_X1 U6508 ( .A1(n5775), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n10408), .B2(
        n10431), .ZN(n5517) );
  INV_X1 U6509 ( .A(n10574), .ZN(n6915) );
  NAND2_X1 U6510 ( .A1(n5978), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n5528) );
  INV_X1 U6511 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n6444) );
  OR2_X1 U6512 ( .A1(n5421), .A2(n6444), .ZN(n5527) );
  INV_X1 U6513 ( .A(n5519), .ZN(n5521) );
  INV_X1 U6514 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n5520) );
  NAND2_X1 U6515 ( .A1(n5521), .A2(n5520), .ZN(n5522) );
  NAND2_X1 U6516 ( .A1(n5523), .A2(n5522), .ZN(n6601) );
  OR2_X1 U6517 ( .A1(n5487), .A2(n6601), .ZN(n5526) );
  INV_X1 U6518 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n5524) );
  OR2_X1 U6519 ( .A1(n5478), .A2(n5524), .ZN(n5525) );
  NAND2_X1 U6520 ( .A1(n5529), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5530) );
  XNOR2_X1 U6521 ( .A(n5530), .B(P1_IR_REG_5__SCAN_IN), .ZN(n6189) );
  AOI22_X1 U6522 ( .A1(n5775), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n10408), .B2(
        n6189), .ZN(n5536) );
  OR2_X1 U6523 ( .A1(n5532), .A2(n5531), .ZN(n5533) );
  NAND2_X1 U6524 ( .A1(n5534), .A2(n5533), .ZN(n6482) );
  OR2_X1 U6525 ( .A1(n5474), .A2(n6482), .ZN(n5535) );
  NAND2_X1 U6526 ( .A1(n5536), .A2(n5535), .ZN(n6600) );
  NAND2_X1 U6527 ( .A1(n6904), .A2(n6600), .ZN(n6902) );
  NAND2_X1 U6528 ( .A1(n5537), .A2(n5245), .ZN(n5539) );
  NAND2_X1 U6529 ( .A1(n10574), .A2(n6629), .ZN(n8241) );
  INV_X1 U6530 ( .A(n6904), .ZN(n9880) );
  NAND2_X1 U6531 ( .A1(n9880), .A2(n6664), .ZN(n6900) );
  NAND2_X1 U6532 ( .A1(n8241), .A2(n6900), .ZN(n5538) );
  NAND2_X1 U6533 ( .A1(n5538), .A2(n8369), .ZN(n8463) );
  NAND2_X1 U6534 ( .A1(n5541), .A2(n5540), .ZN(n5543) );
  XNOR2_X1 U6535 ( .A(n5578), .B(n5544), .ZN(n6969) );
  NAND2_X1 U6536 ( .A1(n6969), .A2(n5975), .ZN(n5548) );
  OR2_X1 U6537 ( .A1(n5563), .A2(n10319), .ZN(n5546) );
  XNOR2_X1 U6538 ( .A(n5546), .B(P1_IR_REG_7__SCAN_IN), .ZN(n9908) );
  AOI22_X1 U6539 ( .A1(n5775), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n10408), .B2(
        n9908), .ZN(n5547) );
  NAND2_X2 U6540 ( .A1(n5548), .A2(n5547), .ZN(n7016) );
  NAND2_X1 U6541 ( .A1(n5978), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n5556) );
  INV_X1 U6542 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n6929) );
  OR2_X1 U6543 ( .A1(n5421), .A2(n6929), .ZN(n5555) );
  INV_X1 U6544 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n5549) );
  NAND2_X1 U6545 ( .A1(n5550), .A2(n5549), .ZN(n5551) );
  NAND2_X1 U6546 ( .A1(n5571), .A2(n5551), .ZN(n6928) );
  OR2_X1 U6547 ( .A1(n5487), .A2(n6928), .ZN(n5554) );
  INV_X1 U6548 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n5552) );
  OR2_X1 U6549 ( .A1(n5478), .A2(n5552), .ZN(n5553) );
  OR2_X1 U6550 ( .A1(n7016), .A2(n7150), .ZN(n8462) );
  NAND2_X1 U6551 ( .A1(n7016), .A2(n7150), .ZN(n8384) );
  NAND2_X1 U6552 ( .A1(n8462), .A2(n8384), .ZN(n6919) );
  INV_X1 U6553 ( .A(n6919), .ZN(n8342) );
  NAND2_X1 U6554 ( .A1(n5578), .A2(n5557), .ZN(n5559) );
  NAND2_X1 U6555 ( .A1(n5559), .A2(n5558), .ZN(n5561) );
  XNOR2_X1 U6556 ( .A(n5561), .B(n5560), .ZN(n7044) );
  NAND2_X1 U6557 ( .A1(n7044), .A2(n5975), .ZN(n5569) );
  INV_X1 U6558 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n5562) );
  INV_X1 U6559 ( .A(n5566), .ZN(n5564) );
  NAND2_X1 U6560 ( .A1(n5564), .A2(P1_IR_REG_8__SCAN_IN), .ZN(n5567) );
  INV_X1 U6561 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n5565) );
  NAND2_X1 U6562 ( .A1(n5566), .A2(n5565), .ZN(n5580) );
  AOI22_X1 U6563 ( .A1(n5775), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n10408), .B2(
        n9922), .ZN(n5568) );
  NAND2_X1 U6564 ( .A1(n5569), .A2(n5568), .ZN(n7138) );
  NAND2_X1 U6565 ( .A1(n5978), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n5576) );
  INV_X1 U6566 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n6952) );
  OR2_X1 U6567 ( .A1(n5421), .A2(n6952), .ZN(n5575) );
  INV_X1 U6568 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n5570) );
  OR2_X1 U6569 ( .A1(n5478), .A2(n5570), .ZN(n5574) );
  NAND2_X1 U6570 ( .A1(n5571), .A2(n7147), .ZN(n5572) );
  NAND2_X1 U6571 ( .A1(n5586), .A2(n5572), .ZN(n7146) );
  OR2_X1 U6572 ( .A1(n5487), .A2(n7146), .ZN(n5573) );
  NAND2_X1 U6573 ( .A1(n7138), .A2(n7181), .ZN(n8247) );
  INV_X1 U6574 ( .A(n8247), .ZN(n8385) );
  OR2_X1 U6575 ( .A1(n7138), .A2(n7181), .ZN(n8400) );
  NAND2_X1 U6576 ( .A1(n7105), .A2(n5975), .ZN(n5583) );
  NAND2_X1 U6577 ( .A1(n5580), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5581) );
  XNOR2_X1 U6578 ( .A(n5581), .B(P1_IR_REG_9__SCAN_IN), .ZN(n10434) );
  AOI22_X1 U6579 ( .A1(n5775), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n10408), .B2(
        n10434), .ZN(n5582) );
  INV_X1 U6580 ( .A(n7287), .ZN(n7093) );
  NAND2_X1 U6581 ( .A1(n5476), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n5591) );
  NAND2_X1 U6582 ( .A1(n5978), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n5590) );
  INV_X1 U6583 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n5584) );
  OR2_X1 U6584 ( .A1(n5478), .A2(n5584), .ZN(n5589) );
  INV_X1 U6585 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n5585) );
  NAND2_X1 U6586 ( .A1(n5586), .A2(n5585), .ZN(n5587) );
  NAND2_X1 U6587 ( .A1(n5599), .A2(n5587), .ZN(n7184) );
  OR2_X1 U6588 ( .A1(n5487), .A2(n7184), .ZN(n5588) );
  NAND4_X1 U6589 ( .A1(n5591), .A2(n5590), .A3(n5589), .A4(n5588), .ZN(n9879)
         );
  AND2_X1 U6590 ( .A1(n7093), .A2(n9879), .ZN(n8251) );
  INV_X1 U6591 ( .A(n9879), .ZN(n8068) );
  NAND2_X1 U6592 ( .A1(n7287), .A2(n8068), .ZN(n8379) );
  XNOR2_X1 U6593 ( .A(n4899), .B(n5592), .ZN(n7158) );
  NAND2_X1 U6594 ( .A1(n7158), .A2(n5975), .ZN(n5597) );
  NOR2_X1 U6595 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_8__SCAN_IN), .ZN(
        n5593) );
  NAND2_X1 U6596 ( .A1(n5594), .A2(n5593), .ZN(n5608) );
  NAND2_X1 U6597 ( .A1(n5608), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5595) );
  XNOR2_X1 U6598 ( .A(n5595), .B(P1_IR_REG_10__SCAN_IN), .ZN(n9935) );
  AOI22_X1 U6599 ( .A1(n5775), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n10408), 
        .B2(n9935), .ZN(n5596) );
  NAND2_X1 U6600 ( .A1(n5597), .A2(n5596), .ZN(n8074) );
  NAND2_X1 U6601 ( .A1(n5978), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n5604) );
  INV_X1 U6602 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n7199) );
  OR2_X1 U6603 ( .A1(n5421), .A2(n7199), .ZN(n5603) );
  NAND2_X1 U6604 ( .A1(n5599), .A2(n5598), .ZN(n5600) );
  NAND2_X1 U6605 ( .A1(n5613), .A2(n5600), .ZN(n8072) );
  OR2_X1 U6606 ( .A1(n5487), .A2(n8072), .ZN(n5602) );
  INV_X1 U6607 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n6064) );
  OR2_X1 U6608 ( .A1(n5478), .A2(n6064), .ZN(n5601) );
  OR2_X1 U6609 ( .A1(n8074), .A2(n7352), .ZN(n8401) );
  NAND2_X1 U6610 ( .A1(n8074), .A2(n7352), .ZN(n8380) );
  NAND2_X1 U6611 ( .A1(n8401), .A2(n8380), .ZN(n8347) );
  INV_X1 U6612 ( .A(n8347), .ZN(n8253) );
  NAND2_X1 U6613 ( .A1(n4896), .A2(n5605), .ZN(n5606) );
  NAND2_X1 U6614 ( .A1(n5607), .A2(n5606), .ZN(n7299) );
  OR2_X1 U6615 ( .A1(n7299), .A2(n5474), .ZN(n5611) );
  NAND2_X1 U6616 ( .A1(n5623), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5609) );
  XNOR2_X1 U6617 ( .A(n5609), .B(P1_IR_REG_11__SCAN_IN), .ZN(n8090) );
  AOI22_X1 U6618 ( .A1(n5775), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n10408), 
        .B2(n8090), .ZN(n5610) );
  NAND2_X1 U6619 ( .A1(n5830), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n5618) );
  NAND2_X1 U6620 ( .A1(n5978), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n5617) );
  INV_X1 U6621 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n5612) );
  NAND2_X1 U6622 ( .A1(n5613), .A2(n5612), .ZN(n5614) );
  NAND2_X1 U6623 ( .A1(n5630), .A2(n5614), .ZN(n7350) );
  OR2_X1 U6624 ( .A1(n5487), .A2(n7350), .ZN(n5616) );
  INV_X1 U6625 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n8081) );
  OR2_X1 U6626 ( .A1(n5421), .A2(n8081), .ZN(n5615) );
  NAND4_X1 U6627 ( .A1(n5618), .A2(n5617), .A3(n5616), .A4(n5615), .ZN(n9877)
         );
  INV_X1 U6628 ( .A(n9877), .ZN(n9770) );
  AND2_X1 U6629 ( .A1(n10268), .A2(n9770), .ZN(n8383) );
  OR2_X1 U6630 ( .A1(n10268), .A2(n9770), .ZN(n8403) );
  OR2_X1 U6631 ( .A1(n5620), .A2(n5619), .ZN(n5621) );
  NAND2_X1 U6632 ( .A1(n5622), .A2(n5621), .ZN(n7415) );
  OR2_X1 U6633 ( .A1(n7415), .A2(n5474), .ZN(n5629) );
  NOR2_X1 U6634 ( .A1(n5623), .A2(P1_IR_REG_11__SCAN_IN), .ZN(n5660) );
  OR2_X1 U6635 ( .A1(n5660), .A2(n10319), .ZN(n5626) );
  INV_X1 U6636 ( .A(n5626), .ZN(n5624) );
  NAND2_X1 U6637 ( .A1(n5624), .A2(P1_IR_REG_12__SCAN_IN), .ZN(n5627) );
  INV_X1 U6638 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n5625) );
  NAND2_X1 U6639 ( .A1(n5626), .A2(n5625), .ZN(n5640) );
  AOI22_X1 U6640 ( .A1(n5775), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n10408), 
        .B2(n6368), .ZN(n5628) );
  NAND2_X1 U6641 ( .A1(n5476), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n5636) );
  INV_X1 U6642 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n6078) );
  OR2_X1 U6643 ( .A1(n5478), .A2(n6078), .ZN(n5635) );
  NAND2_X1 U6644 ( .A1(n5630), .A2(n6360), .ZN(n5631) );
  NAND2_X1 U6645 ( .A1(n5646), .A2(n5631), .ZN(n9774) );
  OR2_X1 U6646 ( .A1(n5487), .A2(n9774), .ZN(n5634) );
  INV_X1 U6647 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n5632) );
  OR2_X1 U6648 ( .A1(n5456), .A2(n5632), .ZN(n5633) );
  INV_X1 U6649 ( .A(n8404), .ZN(n5637) );
  NAND2_X1 U6650 ( .A1(n10263), .A2(n7603), .ZN(n8377) );
  XNOR2_X1 U6651 ( .A(n5639), .B(n5638), .ZN(n7621) );
  NAND2_X1 U6652 ( .A1(n7621), .A2(n5975), .ZN(n5643) );
  NAND2_X1 U6653 ( .A1(n5640), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5641) );
  XNOR2_X1 U6654 ( .A(n5641), .B(P1_IR_REG_13__SCAN_IN), .ZN(n6416) );
  AOI22_X1 U6655 ( .A1(n5775), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n10408), 
        .B2(n6416), .ZN(n5642) );
  NAND2_X1 U6656 ( .A1(n5476), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n5652) );
  INV_X1 U6657 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n5644) );
  OR2_X1 U6658 ( .A1(n5478), .A2(n5644), .ZN(n5651) );
  NAND2_X1 U6659 ( .A1(n5646), .A2(n5645), .ZN(n5647) );
  NAND2_X1 U6660 ( .A1(n5665), .A2(n5647), .ZN(n7611) );
  OR2_X1 U6661 ( .A1(n5487), .A2(n7611), .ZN(n5650) );
  INV_X1 U6662 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n5648) );
  OR2_X1 U6663 ( .A1(n5456), .A2(n5648), .ZN(n5649) );
  NAND2_X1 U6664 ( .A1(n10254), .A2(n7693), .ZN(n8378) );
  NAND2_X1 U6665 ( .A1(n7602), .A2(n8351), .ZN(n7601) );
  NAND2_X1 U6666 ( .A1(n7601), .A2(n8378), .ZN(n7691) );
  NAND2_X1 U6667 ( .A1(n5654), .A2(n5653), .ZN(n5656) );
  NAND2_X1 U6668 ( .A1(n5656), .A2(n5655), .ZN(n5657) );
  NAND2_X1 U6669 ( .A1(n5658), .A2(n5657), .ZN(n7711) );
  NOR2_X1 U6670 ( .A1(P1_IR_REG_12__SCAN_IN), .A2(P1_IR_REG_13__SCAN_IN), .ZN(
        n5659) );
  NAND2_X1 U6671 ( .A1(n5660), .A2(n5659), .ZN(n5675) );
  NAND2_X1 U6672 ( .A1(n5675), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5661) );
  XNOR2_X1 U6673 ( .A(n5661), .B(P1_IR_REG_14__SCAN_IN), .ZN(n6939) );
  AOI22_X1 U6674 ( .A1(n5775), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n10408), 
        .B2(n6939), .ZN(n5662) );
  NAND2_X1 U6675 ( .A1(n5978), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n5670) );
  INV_X1 U6676 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n7699) );
  OR2_X1 U6677 ( .A1(n5421), .A2(n7699), .ZN(n5669) );
  INV_X1 U6678 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n5664) );
  NAND2_X1 U6679 ( .A1(n5665), .A2(n5664), .ZN(n5666) );
  NAND2_X1 U6680 ( .A1(n5680), .A2(n5666), .ZN(n7698) );
  OR2_X1 U6681 ( .A1(n5487), .A2(n7698), .ZN(n5668) );
  INV_X1 U6682 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n6082) );
  OR2_X1 U6683 ( .A1(n5478), .A2(n6082), .ZN(n5667) );
  XNOR2_X1 U6684 ( .A(n8271), .B(n8275), .ZN(n7690) );
  OR2_X1 U6685 ( .A1(n8271), .A2(n8275), .ZN(n8409) );
  OR2_X1 U6686 ( .A1(n5672), .A2(n5242), .ZN(n5673) );
  NAND2_X1 U6687 ( .A1(n5674), .A2(n5673), .ZN(n7789) );
  NAND2_X1 U6688 ( .A1(n5688), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5676) );
  XNOR2_X1 U6689 ( .A(n5676), .B(P1_IR_REG_15__SCAN_IN), .ZN(n7369) );
  AOI22_X1 U6690 ( .A1(n5775), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n10408), 
        .B2(n7369), .ZN(n5677) );
  NAND2_X1 U6691 ( .A1(n5978), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n5685) );
  INV_X1 U6692 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n7365) );
  OR2_X1 U6693 ( .A1(n5421), .A2(n7365), .ZN(n5684) );
  INV_X1 U6694 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n5679) );
  NAND2_X1 U6695 ( .A1(n5680), .A2(n5679), .ZN(n5681) );
  NAND2_X1 U6696 ( .A1(n5693), .A2(n5681), .ZN(n7810) );
  OR2_X1 U6697 ( .A1(n5487), .A2(n7810), .ZN(n5683) );
  INV_X1 U6698 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n10244) );
  OR2_X1 U6699 ( .A1(n5478), .A2(n10244), .ZN(n5682) );
  NAND2_X1 U6700 ( .A1(n7809), .A2(n7878), .ZN(n8376) );
  NAND2_X1 U6701 ( .A1(n7854), .A2(n5975), .ZN(n5691) );
  NAND2_X1 U6702 ( .A1(n5689), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5705) );
  XNOR2_X1 U6703 ( .A(n5705), .B(P1_IR_REG_16__SCAN_IN), .ZN(n6063) );
  AOI22_X1 U6704 ( .A1(n5775), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n10408), 
        .B2(n6063), .ZN(n5690) );
  NAND2_X1 U6705 ( .A1(n5978), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n5698) );
  INV_X1 U6706 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n7874) );
  OR2_X1 U6707 ( .A1(n5421), .A2(n7874), .ZN(n5697) );
  NAND2_X1 U6708 ( .A1(n5693), .A2(n5692), .ZN(n5694) );
  NAND2_X1 U6709 ( .A1(n5726), .A2(n5694), .ZN(n9798) );
  OR2_X1 U6710 ( .A1(n5487), .A2(n9798), .ZN(n5696) );
  INV_X1 U6711 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n6085) );
  OR2_X1 U6712 ( .A1(n5478), .A2(n6085), .ZN(n5695) );
  NAND2_X1 U6713 ( .A1(n7877), .A2(n8416), .ZN(n5699) );
  NAND2_X1 U6714 ( .A1(n10237), .A2(n8110), .ZN(n8371) );
  NAND2_X1 U6715 ( .A1(n5699), .A2(n8371), .ZN(n10138) );
  NAND2_X1 U6716 ( .A1(n5701), .A2(n5700), .ZN(n5703) );
  NAND2_X1 U6717 ( .A1(n5703), .A2(n5702), .ZN(n7905) );
  INV_X1 U6718 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n5704) );
  AOI21_X1 U6719 ( .B1(n5705), .B2(n5704), .A(n10319), .ZN(n5706) );
  NAND2_X1 U6720 ( .A1(n5706), .A2(P1_IR_REG_17__SCAN_IN), .ZN(n5709) );
  INV_X1 U6721 ( .A(n5706), .ZN(n5708) );
  INV_X1 U6722 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n5707) );
  NAND2_X1 U6723 ( .A1(n5708), .A2(n5707), .ZN(n5720) );
  AOI22_X1 U6724 ( .A1(n5775), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n7759), .B2(
        n10408), .ZN(n5710) );
  NAND2_X1 U6725 ( .A1(n5476), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n5715) );
  INV_X1 U6726 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n10233) );
  OR2_X1 U6727 ( .A1(n5478), .A2(n10233), .ZN(n5714) );
  INV_X1 U6728 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n5725) );
  XNOR2_X1 U6729 ( .A(n5726), .B(n5725), .ZN(n10146) );
  OR2_X1 U6730 ( .A1(n5487), .A2(n10146), .ZN(n5713) );
  INV_X1 U6731 ( .A(P1_REG0_REG_17__SCAN_IN), .ZN(n10304) );
  OR2_X1 U6732 ( .A1(n5456), .A2(n10304), .ZN(n5712) );
  NAND2_X1 U6733 ( .A1(n10155), .A2(n9795), .ZN(n8372) );
  INV_X1 U6734 ( .A(n10157), .ZN(n8355) );
  OR2_X1 U6735 ( .A1(n5717), .A2(n5716), .ZN(n5718) );
  NAND2_X1 U6736 ( .A1(n5719), .A2(n5718), .ZN(n7923) );
  NAND2_X1 U6737 ( .A1(n5720), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5721) );
  XNOR2_X1 U6738 ( .A(n5721), .B(P1_IR_REG_18__SCAN_IN), .ZN(n9946) );
  AOI22_X1 U6739 ( .A1(n9946), .A2(n10408), .B1(n5775), .B2(
        P2_DATAO_REG_18__SCAN_IN), .ZN(n5722) );
  NAND2_X1 U6740 ( .A1(n5978), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n5732) );
  INV_X1 U6741 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n10131) );
  OR2_X1 U6742 ( .A1(n5421), .A2(n10131), .ZN(n5731) );
  INV_X1 U6743 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n5724) );
  OAI21_X1 U6744 ( .B1(n5726), .B2(n5725), .A(n5724), .ZN(n5727) );
  NAND2_X1 U6745 ( .A1(n5728), .A2(n5727), .ZN(n10130) );
  OR2_X1 U6746 ( .A1(n5487), .A2(n10130), .ZN(n5730) );
  INV_X1 U6747 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n6061) );
  OR2_X1 U6748 ( .A1(n5478), .A2(n6061), .ZN(n5729) );
  OR2_X1 U6749 ( .A1(n10133), .A2(n10102), .ZN(n5733) );
  NAND2_X1 U6750 ( .A1(n10133), .A2(n10102), .ZN(n8374) );
  NAND2_X1 U6751 ( .A1(n5733), .A2(n8286), .ZN(n5734) );
  AND2_X1 U6752 ( .A1(n5734), .A2(n8374), .ZN(n8388) );
  OR2_X1 U6753 ( .A1(n10109), .A2(n9845), .ZN(n8389) );
  AND2_X1 U6754 ( .A1(n10099), .A2(n8293), .ZN(n10036) );
  AND2_X1 U6755 ( .A1(n10036), .A2(n8396), .ZN(n5735) );
  NAND2_X1 U6756 ( .A1(n10035), .A2(n5735), .ZN(n10022) );
  NAND2_X1 U6757 ( .A1(n5736), .A2(n10022), .ZN(n10023) );
  INV_X1 U6758 ( .A(n10043), .ZN(n10000) );
  OR2_X1 U6759 ( .A1(n10197), .A2(n10000), .ZN(n8238) );
  NAND2_X1 U6760 ( .A1(n10023), .A2(n8238), .ZN(n9996) );
  INV_X1 U6761 ( .A(n5739), .ZN(n5740) );
  MUX2_X1 U6762 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(P2_DATAO_REG_24__SCAN_IN), 
        .S(n6483), .Z(n5741) );
  NAND2_X1 U6763 ( .A1(n5741), .A2(SI_24_), .ZN(n5754) );
  INV_X1 U6764 ( .A(n5741), .ZN(n5742) );
  INV_X1 U6765 ( .A(SI_24_), .ZN(n9591) );
  NAND2_X1 U6766 ( .A1(n5742), .A2(n9591), .ZN(n5743) );
  NAND2_X1 U6767 ( .A1(n5754), .A2(n5743), .ZN(n5755) );
  INV_X1 U6768 ( .A(n5755), .ZN(n5744) );
  NAND2_X1 U6769 ( .A1(n8562), .A2(n5975), .ZN(n5746) );
  NAND2_X1 U6770 ( .A1(n5775), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n5745) );
  INV_X1 U6771 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n9816) );
  NAND2_X1 U6772 ( .A1(n5747), .A2(n9816), .ZN(n5748) );
  NAND2_X1 U6773 ( .A1(n5760), .A2(n5748), .ZN(n10008) );
  OR2_X1 U6774 ( .A1(n10008), .A2(n5487), .ZN(n5753) );
  INV_X1 U6775 ( .A(P1_REG0_REG_24__SCAN_IN), .ZN(n10285) );
  NAND2_X1 U6776 ( .A1(n5476), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n5750) );
  NAND2_X1 U6777 ( .A1(n5830), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n5749) );
  OAI211_X1 U6778 ( .C1(n10285), .C2(n5456), .A(n5750), .B(n5749), .ZN(n5751)
         );
  INV_X1 U6779 ( .A(n5751), .ZN(n5752) );
  INV_X1 U6780 ( .A(n10026), .ZN(n8237) );
  XNOR2_X1 U6781 ( .A(n10007), .B(n8237), .ZN(n9995) );
  MUX2_X1 U6782 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(P2_DATAO_REG_25__SCAN_IN), 
        .S(n6483), .Z(n5769) );
  XNOR2_X1 U6783 ( .A(n5769), .B(SI_25_), .ZN(n5773) );
  XNOR2_X1 U6784 ( .A(n5774), .B(n5773), .ZN(n8698) );
  NAND2_X1 U6785 ( .A1(n8698), .A2(n5975), .ZN(n5758) );
  NAND2_X1 U6786 ( .A1(n5775), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n5757) );
  INV_X1 U6787 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n5759) );
  NAND2_X1 U6788 ( .A1(n5760), .A2(n5759), .ZN(n5761) );
  AND2_X1 U6789 ( .A1(n5779), .A2(n5761), .ZN(n9980) );
  NAND2_X1 U6790 ( .A1(n9980), .A2(n5446), .ZN(n5767) );
  INV_X1 U6791 ( .A(P1_REG0_REG_25__SCAN_IN), .ZN(n5764) );
  NAND2_X1 U6792 ( .A1(n5830), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n5763) );
  NAND2_X1 U6793 ( .A1(n5476), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n5762) );
  OAI211_X1 U6794 ( .C1(n5456), .C2(n5764), .A(n5763), .B(n5762), .ZN(n5765)
         );
  INV_X1 U6795 ( .A(n5765), .ZN(n5766) );
  NAND2_X1 U6796 ( .A1(n10189), .A2(n10001), .ZN(n8423) );
  NAND2_X1 U6797 ( .A1(n8426), .A2(n8423), .ZN(n9984) );
  AND2_X1 U6798 ( .A1(n10007), .A2(n8237), .ZN(n9983) );
  NOR2_X1 U6799 ( .A1(n9984), .A2(n9983), .ZN(n5768) );
  INV_X1 U6800 ( .A(n5769), .ZN(n5771) );
  INV_X1 U6801 ( .A(SI_25_), .ZN(n5770) );
  NAND2_X1 U6802 ( .A1(n5771), .A2(n5770), .ZN(n5772) );
  MUX2_X1 U6803 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(P2_DATAO_REG_26__SCAN_IN), 
        .S(n6110), .Z(n5789) );
  INV_X1 U6804 ( .A(SI_26_), .ZN(n9604) );
  XNOR2_X1 U6805 ( .A(n5789), .B(n9604), .ZN(n5787) );
  XNOR2_X1 U6806 ( .A(n5788), .B(n5787), .ZN(n8709) );
  NAND2_X1 U6807 ( .A1(n8709), .A2(n5975), .ZN(n5777) );
  NAND2_X1 U6808 ( .A1(n5775), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n5776) );
  INV_X1 U6809 ( .A(n5779), .ZN(n5778) );
  INV_X1 U6810 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n9859) );
  NAND2_X1 U6811 ( .A1(n5779), .A2(n9859), .ZN(n5780) );
  NAND2_X1 U6812 ( .A1(n5801), .A2(n5780), .ZN(n9966) );
  INV_X1 U6813 ( .A(P1_REG0_REG_26__SCAN_IN), .ZN(n5783) );
  NAND2_X1 U6814 ( .A1(n5830), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n5782) );
  NAND2_X1 U6815 ( .A1(n5476), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n5781) );
  OAI211_X1 U6816 ( .C1(n5456), .C2(n5783), .A(n5782), .B(n5781), .ZN(n5784)
         );
  INV_X1 U6817 ( .A(n5784), .ZN(n5785) );
  INV_X1 U6818 ( .A(n9988), .ZN(n9786) );
  OR2_X1 U6819 ( .A1(n10182), .A2(n9786), .ZN(n8427) );
  NAND2_X1 U6820 ( .A1(n10182), .A2(n9786), .ZN(n8432) );
  NAND2_X1 U6821 ( .A1(n9973), .A2(n8427), .ZN(n5995) );
  NAND2_X1 U6822 ( .A1(n5788), .A2(n5787), .ZN(n5792) );
  INV_X1 U6823 ( .A(n5789), .ZN(n5790) );
  NAND2_X1 U6824 ( .A1(n5790), .A2(n9604), .ZN(n5791) );
  NAND2_X1 U6825 ( .A1(n5792), .A2(n5791), .ZN(n5810) );
  MUX2_X1 U6826 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(P2_DATAO_REG_27__SCAN_IN), 
        .S(n6483), .Z(n5793) );
  NAND2_X1 U6827 ( .A1(n5793), .A2(SI_27_), .ZN(n5811) );
  INV_X1 U6828 ( .A(n5793), .ZN(n5795) );
  INV_X1 U6829 ( .A(SI_27_), .ZN(n5794) );
  NAND2_X1 U6830 ( .A1(n5795), .A2(n5794), .ZN(n5796) );
  XNOR2_X1 U6831 ( .A(n5810), .B(n5808), .ZN(n8715) );
  NAND2_X1 U6832 ( .A1(n8715), .A2(n5975), .ZN(n5798) );
  NAND2_X1 U6833 ( .A1(n5775), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n5797) );
  INV_X1 U6834 ( .A(n5801), .ZN(n5799) );
  NAND2_X1 U6835 ( .A1(n5799), .A2(P1_REG3_REG_27__SCAN_IN), .ZN(n5816) );
  INV_X1 U6836 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n5800) );
  NAND2_X1 U6837 ( .A1(n5801), .A2(n5800), .ZN(n5802) );
  NAND2_X1 U6838 ( .A1(n5816), .A2(n5802), .ZN(n8502) );
  OR2_X1 U6839 ( .A1(n8502), .A2(n5487), .ZN(n5807) );
  INV_X1 U6840 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n6000) );
  NAND2_X1 U6841 ( .A1(n5476), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n5804) );
  NAND2_X1 U6842 ( .A1(n5830), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n5803) );
  OAI211_X1 U6843 ( .C1(n6000), .C2(n5456), .A(n5804), .B(n5803), .ZN(n5805)
         );
  INV_X1 U6844 ( .A(n5805), .ZN(n5806) );
  NAND2_X1 U6845 ( .A1(n9722), .A2(n9971), .ZN(n8430) );
  INV_X1 U6846 ( .A(n5808), .ZN(n5809) );
  NAND2_X1 U6847 ( .A1(n5812), .A2(n5811), .ZN(n5827) );
  MUX2_X1 U6848 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(P2_DATAO_REG_28__SCAN_IN), 
        .S(n6483), .Z(n5822) );
  XNOR2_X1 U6849 ( .A(n5822), .B(SI_28_), .ZN(n5826) );
  NAND2_X1 U6850 ( .A1(n8728), .A2(n5975), .ZN(n5814) );
  NAND2_X1 U6851 ( .A1(n5775), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n5813) );
  INV_X1 U6852 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n5815) );
  NAND2_X1 U6853 ( .A1(n5816), .A2(n5815), .ZN(n5817) );
  INV_X1 U6854 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n5820) );
  NAND2_X1 U6855 ( .A1(n5476), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n5819) );
  NAND2_X1 U6856 ( .A1(n5830), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n5818) );
  OAI211_X1 U6857 ( .C1(n5456), .C2(n5820), .A(n5819), .B(n5818), .ZN(n5821)
         );
  OR2_X1 U6858 ( .A1(n10173), .A2(n9717), .ZN(n8313) );
  NAND2_X1 U6859 ( .A1(n10173), .A2(n9717), .ZN(n8431) );
  INV_X1 U6860 ( .A(n8509), .ZN(n8513) );
  NAND2_X1 U6861 ( .A1(n8514), .A2(n8431), .ZN(n5839) );
  INV_X1 U6862 ( .A(n5822), .ZN(n5824) );
  INV_X1 U6863 ( .A(SI_28_), .ZN(n5823) );
  NAND2_X1 U6864 ( .A1(n5824), .A2(n5823), .ZN(n5825) );
  INV_X1 U6865 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n8551) );
  INV_X1 U6866 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n8024) );
  MUX2_X1 U6867 ( .A(n8551), .B(n8024), .S(n6483), .Z(n5959) );
  NAND2_X1 U6868 ( .A1(n8550), .A2(n5975), .ZN(n5829) );
  NAND2_X1 U6869 ( .A1(n5775), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n5828) );
  INV_X1 U6870 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n5833) );
  NAND2_X1 U6871 ( .A1(n5476), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n5832) );
  NAND2_X1 U6872 ( .A1(n5830), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n5831) );
  OAI211_X1 U6873 ( .C1(n5833), .C2(n5456), .A(n5832), .B(n5831), .ZN(n5834)
         );
  INV_X1 U6874 ( .A(n5834), .ZN(n5835) );
  OAI21_X1 U6875 ( .B1(n5951), .B2(n5487), .A(n5835), .ZN(n9869) );
  INV_X1 U6876 ( .A(n9869), .ZN(n5837) );
  NAND2_X1 U6877 ( .A1(n10169), .A2(n5837), .ZN(n8434) );
  NAND2_X1 U6878 ( .A1(n8314), .A2(n8434), .ZN(n8361) );
  INV_X1 U6879 ( .A(n8361), .ZN(n5838) );
  XNOR2_X1 U6880 ( .A(n5839), .B(n5838), .ZN(n5858) );
  NAND2_X1 U6881 ( .A1(n4895), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5842) );
  INV_X1 U6882 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n5840) );
  NAND2_X1 U6883 ( .A1(n5842), .A2(n5840), .ZN(n5844) );
  NAND2_X1 U6884 ( .A1(n5844), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5841) );
  NAND2_X1 U6885 ( .A1(n8497), .A2(n10019), .ZN(n5849) );
  INV_X1 U6886 ( .A(n5842), .ZN(n5843) );
  NAND2_X1 U6887 ( .A1(n5843), .A2(P1_IR_REG_21__SCAN_IN), .ZN(n5845) );
  NAND2_X1 U6888 ( .A1(n5846), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5847) );
  XNOR2_X1 U6889 ( .A(n5847), .B(P1_IR_REG_20__SCAN_IN), .ZN(n8329) );
  OR2_X1 U6890 ( .A1(n8440), .A2(n8486), .ZN(n5848) );
  NAND2_X1 U6891 ( .A1(n5849), .A2(n5848), .ZN(n10140) );
  INV_X1 U6892 ( .A(n9717), .ZN(n9870) );
  NOR2_X2 U6893 ( .A1(n5850), .A2(n6003), .ZN(n10143) );
  INV_X1 U6894 ( .A(n6003), .ZN(n8325) );
  INV_X1 U6895 ( .A(P1_B_REG_SCAN_IN), .ZN(n5852) );
  OR2_X1 U6896 ( .A1(n4855), .A2(n5852), .ZN(n5853) );
  AND2_X1 U6897 ( .A1(n10141), .A2(n5853), .ZN(n5982) );
  INV_X1 U6898 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n10166) );
  NAND2_X1 U6899 ( .A1(n5476), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n5855) );
  NAND2_X1 U6900 ( .A1(n5978), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n5854) );
  OAI211_X1 U6901 ( .C1(n5478), .C2(n10166), .A(n5855), .B(n5854), .ZN(n9868)
         );
  INV_X1 U6902 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n5860) );
  NAND2_X1 U6903 ( .A1(n5861), .A2(n5860), .ZN(n5868) );
  OR2_X1 U6904 ( .A1(n5861), .A2(n5860), .ZN(n5862) );
  NAND2_X1 U6905 ( .A1(n5868), .A2(n5862), .ZN(n5886) );
  NAND2_X1 U6906 ( .A1(n5886), .A2(P1_B_REG_SCAN_IN), .ZN(n5867) );
  INV_X1 U6907 ( .A(n5863), .ZN(n5890) );
  NAND2_X1 U6908 ( .A1(n5890), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5865) );
  XNOR2_X1 U6909 ( .A(n5865), .B(n5864), .ZN(n7189) );
  INV_X1 U6910 ( .A(n7189), .ZN(n5866) );
  MUX2_X1 U6911 ( .A(n5867), .B(P1_B_REG_SCAN_IN), .S(n5866), .Z(n5870) );
  NAND2_X1 U6912 ( .A1(n5870), .A2(n5887), .ZN(n5880) );
  INV_X1 U6913 ( .A(n5886), .ZN(n5871) );
  OAI22_X1 U6914 ( .A1(n5880), .A2(P1_D_REG_1__SCAN_IN), .B1(n5887), .B2(n5871), .ZN(n5987) );
  INV_X1 U6915 ( .A(n5987), .ZN(n5883) );
  NOR4_X1 U6916 ( .A1(P1_D_REG_15__SCAN_IN), .A2(P1_D_REG_14__SCAN_IN), .A3(
        P1_D_REG_13__SCAN_IN), .A4(P1_D_REG_12__SCAN_IN), .ZN(n5875) );
  NOR4_X1 U6917 ( .A1(P1_D_REG_17__SCAN_IN), .A2(P1_D_REG_19__SCAN_IN), .A3(
        P1_D_REG_18__SCAN_IN), .A4(P1_D_REG_16__SCAN_IN), .ZN(n5874) );
  NOR4_X1 U6918 ( .A1(P1_D_REG_7__SCAN_IN), .A2(P1_D_REG_6__SCAN_IN), .A3(
        P1_D_REG_5__SCAN_IN), .A4(P1_D_REG_2__SCAN_IN), .ZN(n5873) );
  NOR4_X1 U6919 ( .A1(P1_D_REG_11__SCAN_IN), .A2(P1_D_REG_10__SCAN_IN), .A3(
        P1_D_REG_9__SCAN_IN), .A4(P1_D_REG_8__SCAN_IN), .ZN(n5872) );
  NAND4_X1 U6920 ( .A1(n5875), .A2(n5874), .A3(n5873), .A4(n5872), .ZN(n5882)
         );
  NOR2_X1 U6921 ( .A1(P1_D_REG_31__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .ZN(
        n5879) );
  NOR4_X1 U6922 ( .A1(P1_D_REG_4__SCAN_IN), .A2(P1_D_REG_3__SCAN_IN), .A3(
        P1_D_REG_29__SCAN_IN), .A4(P1_D_REG_28__SCAN_IN), .ZN(n5878) );
  NOR4_X1 U6923 ( .A1(P1_D_REG_23__SCAN_IN), .A2(P1_D_REG_22__SCAN_IN), .A3(
        P1_D_REG_21__SCAN_IN), .A4(P1_D_REG_20__SCAN_IN), .ZN(n5877) );
  NOR4_X1 U6924 ( .A1(P1_D_REG_27__SCAN_IN), .A2(P1_D_REG_26__SCAN_IN), .A3(
        P1_D_REG_25__SCAN_IN), .A4(P1_D_REG_24__SCAN_IN), .ZN(n5876) );
  NAND4_X1 U6925 ( .A1(n5879), .A2(n5878), .A3(n5877), .A4(n5876), .ZN(n5881)
         );
  OAI21_X1 U6926 ( .B1(n5882), .B2(n5881), .A(n10317), .ZN(n5989) );
  AND2_X1 U6927 ( .A1(n5883), .A2(n5989), .ZN(n6199) );
  INV_X1 U6928 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n5884) );
  NAND2_X1 U6929 ( .A1(n10317), .A2(n5884), .ZN(n5885) );
  INV_X1 U6930 ( .A(n5887), .ZN(n7539) );
  NAND2_X1 U6931 ( .A1(n7539), .A2(n7189), .ZN(n10318) );
  NOR2_X1 U6932 ( .A1(n5886), .A2(n7189), .ZN(n5888) );
  NAND2_X1 U6933 ( .A1(n4910), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5889) );
  MUX2_X1 U6934 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5889), .S(
        P1_IR_REG_23__SCAN_IN), .Z(n5891) );
  NAND2_X1 U6935 ( .A1(n5891), .A2(n5890), .ZN(n7005) );
  OR2_X1 U6936 ( .A1(n6003), .A2(n6210), .ZN(n6321) );
  INV_X1 U6937 ( .A(n6321), .ZN(n5893) );
  OR2_X1 U6938 ( .A1(n10405), .A2(n5893), .ZN(n6202) );
  NOR2_X1 U6939 ( .A1(n6198), .A2(n6202), .ZN(n5894) );
  NAND2_X1 U6940 ( .A1(n6199), .A2(n5894), .ZN(n5950) );
  NAND2_X1 U6941 ( .A1(n5945), .A2(n8440), .ZN(n6451) );
  NAND2_X1 U6942 ( .A1(n6343), .A2(n5895), .ZN(n6342) );
  NAND2_X1 U6943 ( .A1(n6277), .A2(n6278), .ZN(n5896) );
  AND2_X1 U6944 ( .A1(n6342), .A2(n5896), .ZN(n6859) );
  NAND2_X1 U6945 ( .A1(n6859), .A2(n6860), .ZN(n6858) );
  NAND2_X1 U6946 ( .A1(n6303), .A2(n10519), .ZN(n5897) );
  NAND2_X1 U6947 ( .A1(n6858), .A2(n5897), .ZN(n6426) );
  NAND2_X1 U6948 ( .A1(n5898), .A2(n6875), .ZN(n8335) );
  NAND2_X1 U6949 ( .A1(n6426), .A2(n8335), .ZN(n6425) );
  NAND2_X1 U6950 ( .A1(n6879), .A2(n6621), .ZN(n5899) );
  NAND2_X1 U6951 ( .A1(n6425), .A2(n5899), .ZN(n6874) );
  XNOR2_X1 U6952 ( .A(n9881), .B(n10549), .ZN(n8341) );
  NAND2_X1 U6953 ( .A1(n6874), .A2(n8341), .ZN(n6873) );
  INV_X1 U6954 ( .A(n9881), .ZN(n6439) );
  NAND2_X1 U6955 ( .A1(n6439), .A2(n10549), .ZN(n5900) );
  NAND2_X1 U6956 ( .A1(n6873), .A2(n5900), .ZN(n6443) );
  INV_X1 U6957 ( .A(n6443), .ZN(n5903) );
  AND2_X1 U6958 ( .A1(n10574), .A2(n6923), .ZN(n5901) );
  NAND2_X1 U6959 ( .A1(n9880), .A2(n6600), .ZN(n6895) );
  NAND2_X1 U6960 ( .A1(n8369), .A2(n8241), .ZN(n6894) );
  AND2_X1 U6961 ( .A1(n6895), .A2(n6894), .ZN(n6896) );
  NAND2_X1 U6962 ( .A1(n6920), .A2(n6919), .ZN(n6918) );
  INV_X1 U6963 ( .A(n7150), .ZN(n6831) );
  OR2_X1 U6964 ( .A1(n7016), .A2(n6831), .ZN(n5904) );
  INV_X1 U6965 ( .A(n8344), .ZN(n5905) );
  INV_X1 U6966 ( .A(n7181), .ZN(n7087) );
  NAND2_X1 U6967 ( .A1(n7138), .A2(n7087), .ZN(n5906) );
  AND2_X1 U6968 ( .A1(n7287), .A2(n9879), .ZN(n5908) );
  INV_X1 U6969 ( .A(n7352), .ZN(n9878) );
  OR2_X1 U6970 ( .A1(n8074), .A2(n9878), .ZN(n5909) );
  NOR2_X1 U6971 ( .A1(n10268), .A2(n9877), .ZN(n5910) );
  NAND2_X1 U6972 ( .A1(n10268), .A2(n9877), .ZN(n5911) );
  NAND2_X1 U6973 ( .A1(n5912), .A2(n5911), .ZN(n7479) );
  NAND2_X1 U6974 ( .A1(n8404), .A2(n8377), .ZN(n8348) );
  NAND2_X1 U6975 ( .A1(n7479), .A2(n8348), .ZN(n5914) );
  INV_X1 U6976 ( .A(n7603), .ZN(n9876) );
  NAND2_X1 U6977 ( .A1(n10263), .A2(n9876), .ZN(n5913) );
  INV_X1 U6978 ( .A(n7693), .ZN(n9875) );
  OR2_X1 U6979 ( .A1(n10254), .A2(n9875), .ZN(n5915) );
  NAND2_X1 U6980 ( .A1(n7689), .A2(n7690), .ZN(n7688) );
  INV_X1 U6981 ( .A(n8275), .ZN(n9874) );
  OR2_X1 U6982 ( .A1(n8271), .A2(n9874), .ZN(n5916) );
  INV_X1 U6983 ( .A(n8352), .ZN(n5917) );
  INV_X1 U6984 ( .A(n7878), .ZN(n9873) );
  NAND2_X1 U6985 ( .A1(n7809), .A2(n9873), .ZN(n5918) );
  NAND2_X1 U6986 ( .A1(n8416), .A2(n8371), .ZN(n8354) );
  NAND2_X1 U6987 ( .A1(n7871), .A2(n8354), .ZN(n5920) );
  INV_X1 U6988 ( .A(n8110), .ZN(n10144) );
  NAND2_X1 U6989 ( .A1(n10237), .A2(n10144), .ZN(n5919) );
  NAND2_X1 U6990 ( .A1(n5920), .A2(n5919), .ZN(n10158) );
  INV_X1 U6991 ( .A(n9795), .ZN(n10126) );
  INV_X1 U6992 ( .A(n10102), .ZN(n10142) );
  NAND2_X1 U6993 ( .A1(n10133), .A2(n10142), .ZN(n8239) );
  OR2_X1 U6994 ( .A1(n10109), .A2(n10125), .ZN(n10057) );
  NAND2_X1 U6995 ( .A1(n10075), .A2(n10094), .ZN(n5923) );
  INV_X1 U6996 ( .A(n10104), .ZN(n10070) );
  NAND2_X1 U6997 ( .A1(n10213), .A2(n10070), .ZN(n10060) );
  INV_X1 U6998 ( .A(n5929), .ZN(n5927) );
  NAND2_X1 U6999 ( .A1(n10065), .A2(n5924), .ZN(n10092) );
  AND2_X1 U7000 ( .A1(n10092), .A2(n5925), .ZN(n5926) );
  INV_X1 U7001 ( .A(n5928), .ZN(n5931) );
  NAND2_X1 U7002 ( .A1(n10109), .A2(n10125), .ZN(n10058) );
  AND2_X1 U7003 ( .A1(n10058), .A2(n5929), .ZN(n5930) );
  NAND2_X1 U7004 ( .A1(n5933), .A2(n5932), .ZN(n10034) );
  AND2_X1 U7005 ( .A1(n10205), .A2(n10071), .ZN(n5934) );
  OAI22_X1 U7006 ( .A1(n10034), .A2(n5934), .B1(n10071), .B2(n10205), .ZN(
        n10015) );
  NOR2_X1 U7007 ( .A1(n10197), .A2(n10043), .ZN(n5935) );
  NAND2_X1 U7008 ( .A1(n10197), .A2(n10043), .ZN(n5936) );
  NAND2_X1 U7009 ( .A1(n5937), .A2(n5936), .ZN(n9994) );
  AND2_X1 U7010 ( .A1(n10007), .A2(n10026), .ZN(n5939) );
  OR2_X1 U7011 ( .A1(n10007), .A2(n10026), .ZN(n5938) );
  OR2_X1 U7012 ( .A1(n10189), .A2(n9872), .ZN(n5940) );
  NOR2_X1 U7013 ( .A1(n10182), .A2(n9988), .ZN(n5942) );
  NAND2_X1 U7014 ( .A1(n10182), .A2(n9988), .ZN(n5941) );
  INV_X1 U7015 ( .A(n8510), .ZN(n5943) );
  NAND2_X1 U7016 ( .A1(n5943), .A2(n8513), .ZN(n8512) );
  NAND2_X1 U7017 ( .A1(n8512), .A2(n5240), .ZN(n5944) );
  INV_X2 U7018 ( .A(n10088), .ZN(n10148) );
  OR2_X1 U7019 ( .A1(n6003), .A2(n8491), .ZN(n6203) );
  AND2_X2 U7020 ( .A1(n6203), .A2(n6451), .ZN(n6248) );
  OAI21_X1 U7021 ( .B1(n5945), .B2(n10019), .A(n8491), .ZN(n5946) );
  AND2_X4 U7022 ( .A1(n6248), .A2(n5946), .ZN(n6282) );
  NOR2_X1 U7023 ( .A1(n6212), .A2(n9951), .ZN(n6616) );
  OR2_X1 U7024 ( .A1(n6282), .A2(n6616), .ZN(n5947) );
  NAND2_X1 U7025 ( .A1(n10148), .A2(n5947), .ZN(n10137) );
  INV_X1 U7026 ( .A(n10213), .ZN(n10090) );
  NAND2_X1 U7027 ( .A1(n6866), .A2(n10519), .ZN(n6430) );
  OR2_X1 U7028 ( .A1(n6430), .A2(n9740), .ZN(n6885) );
  INV_X1 U7029 ( .A(n8074), .ZN(n10601) );
  AND2_X1 U7030 ( .A1(n10601), .A2(n7093), .ZN(n5948) );
  NAND2_X1 U7031 ( .A1(n7091), .A2(n5948), .ZN(n7197) );
  INV_X1 U7032 ( .A(n8271), .ZN(n10249) );
  INV_X1 U7033 ( .A(n10133), .ZN(n10223) );
  NAND2_X1 U7034 ( .A1(n10090), .A2(n10108), .ZN(n10083) );
  NAND2_X1 U7035 ( .A1(n10287), .A2(n10017), .ZN(n10004) );
  AOI211_X1 U7036 ( .C1(n10169), .C2(n8520), .A(n10591), .B(n9958), .ZN(n10168) );
  NOR2_X1 U7037 ( .A1(n5950), .A2(n10019), .ZN(n10110) );
  NOR2_X1 U7038 ( .A1(n6451), .A2(n8486), .ZN(n6205) );
  INV_X1 U7039 ( .A(n5951), .ZN(n5952) );
  INV_X1 U7040 ( .A(n10145), .ZN(n10111) );
  AOI22_X1 U7041 ( .A1(n5952), .A2(n10111), .B1(P1_REG2_REG_29__SCAN_IN), .B2(
        n10088), .ZN(n5953) );
  OAI21_X1 U7042 ( .B1(n5836), .B2(n10115), .A(n5953), .ZN(n5954) );
  AOI21_X1 U7043 ( .B1(n10168), .B2(n10110), .A(n5954), .ZN(n5955) );
  OAI21_X1 U7044 ( .B1(n10172), .B2(n10137), .A(n5955), .ZN(n5956) );
  INV_X1 U7045 ( .A(n5956), .ZN(n5957) );
  NAND2_X1 U7046 ( .A1(n5228), .A2(n5957), .ZN(P1_U3355) );
  INV_X1 U7047 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n5991) );
  INV_X1 U7048 ( .A(SI_29_), .ZN(n9597) );
  MUX2_X1 U7049 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(P2_DATAO_REG_30__SCAN_IN), 
        .S(n6110), .Z(n5964) );
  XNOR2_X1 U7050 ( .A(n5964), .B(SI_30_), .ZN(n5967) );
  NAND2_X1 U7051 ( .A1(n8540), .A2(n5975), .ZN(n5963) );
  NAND2_X1 U7052 ( .A1(n5775), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n5962) );
  NAND2_X1 U7053 ( .A1(n10279), .A2(n9958), .ZN(n10162) );
  NAND2_X1 U7054 ( .A1(n5964), .A2(SI_30_), .ZN(n5966) );
  INV_X1 U7055 ( .A(n5966), .ZN(n5969) );
  INV_X1 U7056 ( .A(n5967), .ZN(n5968) );
  MUX2_X1 U7057 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(P2_DATAO_REG_31__SCAN_IN), 
        .S(n6483), .Z(n5972) );
  XNOR2_X1 U7058 ( .A(n5972), .B(SI_31_), .ZN(n5973) );
  NAND2_X1 U7059 ( .A1(n9704), .A2(n5975), .ZN(n5977) );
  NAND2_X1 U7060 ( .A1(n5775), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(n5976) );
  XNOR2_X1 U7061 ( .A(n10162), .B(n8233), .ZN(n8100) );
  NAND2_X1 U7062 ( .A1(n5476), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n5981) );
  NAND2_X1 U7063 ( .A1(n5978), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n5980) );
  OR2_X1 U7064 ( .A1(n5478), .A2(n5991), .ZN(n5979) );
  AND3_X1 U7065 ( .A1(n5981), .A2(n5980), .A3(n5979), .ZN(n8232) );
  INV_X1 U7066 ( .A(n8232), .ZN(n9867) );
  NAND2_X1 U7067 ( .A1(n9867), .A2(n5982), .ZN(n10164) );
  AOI21_X1 U7068 ( .B1(n5985), .B2(n5984), .A(n5983), .ZN(n8062) );
  INV_X1 U7069 ( .A(n10405), .ZN(n5986) );
  AND2_X1 U7070 ( .A1(n5987), .A2(n5986), .ZN(n10403) );
  AND3_X1 U7071 ( .A1(n5989), .A2(n5988), .A3(n6321), .ZN(n5990) );
  MUX2_X1 U7072 ( .A(n5991), .B(n8062), .S(n10608), .Z(n5993) );
  INV_X1 U7073 ( .A(n6451), .ZN(n5992) );
  NAND2_X1 U7074 ( .A1(n10608), .A2(n10269), .ZN(n10246) );
  NAND2_X1 U7075 ( .A1(n5993), .A2(n5230), .ZN(P1_U3554) );
  AOI21_X1 U7076 ( .B1(n9722), .B2(n9964), .A(n8519), .ZN(n8501) );
  OAI211_X1 U7077 ( .C1(n5995), .C2(n8473), .A(n5994), .B(n10140), .ZN(n5997)
         );
  NAND2_X1 U7078 ( .A1(n9988), .A2(n10143), .ZN(n5996) );
  OAI211_X1 U7079 ( .C1(n9717), .C2(n10103), .A(n5997), .B(n5996), .ZN(n8506)
         );
  NAND2_X1 U7080 ( .A1(n5945), .A2(n10019), .ZN(n8319) );
  INV_X1 U7081 ( .A(n10273), .ZN(n10603) );
  INV_X1 U7082 ( .A(n6198), .ZN(n5998) );
  MUX2_X1 U7083 ( .A(n6000), .B(n10178), .S(n10612), .Z(n6001) );
  INV_X1 U7084 ( .A(n9722), .ZN(n10181) );
  NAND2_X1 U7085 ( .A1(n10612), .A2(n10269), .ZN(n10311) );
  NAND2_X1 U7086 ( .A1(n6001), .A2(n5239), .ZN(P1_U3518) );
  INV_X1 U7087 ( .A(n7005), .ZN(n6002) );
  OR2_X1 U7088 ( .A1(n6003), .A2(n6002), .ZN(n6004) );
  NAND2_X1 U7089 ( .A1(n6093), .A2(n6004), .ZN(n6089) );
  OAI21_X1 U7090 ( .B1(n6089), .B2(n10408), .A(P1_STATE_REG_SCAN_IN), .ZN(
        P1_U3083) );
  INV_X1 U7091 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n6138) );
  INV_X1 U7092 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n6150) );
  INV_X1 U7093 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n6011) );
  NAND3_X1 U7094 ( .A1(n6138), .A2(n6150), .A3(n6011), .ZN(n6012) );
  INV_X1 U7095 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n6014) );
  NAND2_X1 U7096 ( .A1(n6163), .A2(n6015), .ZN(n6226) );
  NOR2_X1 U7097 ( .A1(P2_IR_REG_20__SCAN_IN), .A2(P2_IR_REG_19__SCAN_IN), .ZN(
        n6025) );
  INV_X1 U7098 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n6018) );
  NAND4_X1 U7099 ( .A1(n6025), .A2(n6024), .A3(n6023), .A4(n6022), .ZN(n6031)
         );
  NOR2_X1 U7100 ( .A1(P2_IR_REG_22__SCAN_IN), .A2(P2_IR_REG_21__SCAN_IN), .ZN(
        n6029) );
  NOR2_X1 U7101 ( .A1(P2_IR_REG_17__SCAN_IN), .A2(P2_IR_REG_18__SCAN_IN), .ZN(
        n6028) );
  NOR2_X1 U7102 ( .A1(P2_IR_REG_16__SCAN_IN), .A2(P2_IR_REG_15__SCAN_IN), .ZN(
        n6027) );
  NOR2_X1 U7103 ( .A1(P2_IR_REG_13__SCAN_IN), .A2(P2_IR_REG_14__SCAN_IN), .ZN(
        n6026) );
  NAND4_X1 U7104 ( .A1(n6029), .A2(n6028), .A3(n6027), .A4(n6026), .ZN(n6030)
         );
  NOR2_X1 U7105 ( .A1(n6031), .A2(n6030), .ZN(n6032) );
  NAND2_X1 U7106 ( .A1(n6034), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6033) );
  MUX2_X1 U7107 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6033), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n6035) );
  NOR2_X2 U7108 ( .A1(n6034), .A2(P2_IR_REG_26__SCAN_IN), .ZN(n6232) );
  INV_X1 U7109 ( .A(n6232), .ZN(n6234) );
  NAND2_X1 U7110 ( .A1(n6036), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6037) );
  MUX2_X1 U7111 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6037), .S(
        P2_IR_REG_25__SCAN_IN), .Z(n6038) );
  NAND2_X1 U7112 ( .A1(n6038), .A2(n6034), .ZN(n7360) );
  INV_X2 U7113 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3084) );
  INV_X2 U7114 ( .A(n9883), .ZN(P1_U4006) );
  NOR2_X1 U7115 ( .A1(n9946), .A2(n10131), .ZN(n6040) );
  AOI21_X1 U7116 ( .B1(n9946), .B2(n10131), .A(n6040), .ZN(n6060) );
  NOR2_X1 U7117 ( .A1(n8090), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n8079) );
  NAND2_X1 U7118 ( .A1(n10434), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n6041) );
  OAI21_X1 U7119 ( .B1(n10434), .B2(P1_REG2_REG_9__SCAN_IN), .A(n6041), .ZN(
        n10439) );
  NOR2_X1 U7120 ( .A1(P1_REG2_REG_8__SCAN_IN), .A2(n9922), .ZN(n6042) );
  AOI21_X1 U7121 ( .B1(n9922), .B2(P1_REG2_REG_8__SCAN_IN), .A(n6042), .ZN(
        n9920) );
  NAND2_X1 U7122 ( .A1(n10431), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n6043) );
  OAI21_X1 U7123 ( .B1(n10431), .B2(P1_REG2_REG_6__SCAN_IN), .A(n6043), .ZN(
        n10428) );
  NOR2_X1 U7124 ( .A1(P1_REG2_REG_5__SCAN_IN), .A2(n6189), .ZN(n6044) );
  AOI21_X1 U7125 ( .B1(n6189), .B2(P1_REG2_REG_5__SCAN_IN), .A(n6044), .ZN(
        n6186) );
  INV_X1 U7126 ( .A(n6114), .ZN(n10458) );
  NAND2_X1 U7127 ( .A1(P1_REG2_REG_1__SCAN_IN), .A2(n10458), .ZN(n6045) );
  OAI21_X1 U7128 ( .B1(n10458), .B2(P1_REG2_REG_1__SCAN_IN), .A(n6045), .ZN(
        n10453) );
  NAND2_X1 U7129 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n10454) );
  NOR2_X1 U7130 ( .A1(n10453), .A2(n10454), .ZN(n10452) );
  AOI21_X1 U7131 ( .B1(n10458), .B2(P1_REG2_REG_1__SCAN_IN), .A(n10452), .ZN(
        n6266) );
  NAND2_X1 U7132 ( .A1(P1_REG2_REG_2__SCAN_IN), .A2(n6269), .ZN(n6046) );
  OAI21_X1 U7133 ( .B1(n6269), .B2(P1_REG2_REG_2__SCAN_IN), .A(n6046), .ZN(
        n6265) );
  NOR2_X1 U7134 ( .A1(n6266), .A2(n6265), .ZN(n6264) );
  AOI21_X1 U7135 ( .B1(n6269), .B2(P1_REG2_REG_2__SCAN_IN), .A(n6264), .ZN(
        n6101) );
  NAND2_X1 U7136 ( .A1(P1_REG2_REG_3__SCAN_IN), .A2(n6105), .ZN(n6047) );
  OAI21_X1 U7137 ( .B1(n6105), .B2(P1_REG2_REG_3__SCAN_IN), .A(n6047), .ZN(
        n6100) );
  NOR2_X1 U7138 ( .A1(n6101), .A2(n6100), .ZN(n6099) );
  NOR2_X1 U7139 ( .A1(n9895), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n6048) );
  AOI21_X1 U7140 ( .B1(P1_REG2_REG_4__SCAN_IN), .B2(n9895), .A(n6048), .ZN(
        n9892) );
  NAND2_X1 U7141 ( .A1(n9893), .A2(n9892), .ZN(n9891) );
  OAI21_X1 U7142 ( .B1(n9895), .B2(P1_REG2_REG_4__SCAN_IN), .A(n9891), .ZN(
        n6187) );
  NAND2_X1 U7143 ( .A1(n6186), .A2(n6187), .ZN(n6185) );
  OAI21_X1 U7144 ( .B1(n6189), .B2(P1_REG2_REG_5__SCAN_IN), .A(n6185), .ZN(
        n10429) );
  NOR2_X1 U7145 ( .A1(n10428), .A2(n10429), .ZN(n10427) );
  NOR2_X1 U7146 ( .A1(n9908), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n6049) );
  AOI21_X1 U7147 ( .B1(P1_REG2_REG_7__SCAN_IN), .B2(n9908), .A(n6049), .ZN(
        n9905) );
  NAND2_X1 U7148 ( .A1(n9906), .A2(n9905), .ZN(n9904) );
  OAI21_X1 U7149 ( .B1(n9908), .B2(P1_REG2_REG_7__SCAN_IN), .A(n9904), .ZN(
        n9919) );
  NAND2_X1 U7150 ( .A1(n9920), .A2(n9919), .ZN(n9918) );
  OAI21_X1 U7151 ( .B1(P1_REG2_REG_8__SCAN_IN), .B2(n9922), .A(n9918), .ZN(
        n10440) );
  NOR2_X1 U7152 ( .A1(n10439), .A2(n10440), .ZN(n10438) );
  MUX2_X1 U7153 ( .A(P1_REG2_REG_10__SCAN_IN), .B(n7199), .S(n9935), .Z(n6050)
         );
  INV_X1 U7154 ( .A(n6050), .ZN(n9932) );
  NOR2_X1 U7155 ( .A1(n9933), .A2(n9932), .ZN(n9931) );
  NOR2_X1 U7156 ( .A1(n8079), .A2(n8082), .ZN(n8077) );
  AND2_X1 U7157 ( .A1(n8090), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n8078) );
  OR2_X1 U7158 ( .A1(n6368), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n6052) );
  NAND2_X1 U7159 ( .A1(P1_REG2_REG_12__SCAN_IN), .A2(n6368), .ZN(n6051) );
  NAND2_X1 U7160 ( .A1(n6052), .A2(n6051), .ZN(n6364) );
  NOR2_X1 U7161 ( .A1(n6365), .A2(n6364), .ZN(n6363) );
  AOI21_X1 U7162 ( .B1(n6368), .B2(P1_REG2_REG_12__SCAN_IN), .A(n6363), .ZN(
        n6414) );
  NAND2_X1 U7163 ( .A1(P1_REG2_REG_13__SCAN_IN), .A2(n6416), .ZN(n6053) );
  OAI21_X1 U7164 ( .B1(n6416), .B2(P1_REG2_REG_13__SCAN_IN), .A(n6053), .ZN(
        n6413) );
  NOR2_X1 U7165 ( .A1(n6414), .A2(n6413), .ZN(n6412) );
  AOI21_X1 U7166 ( .B1(n6416), .B2(P1_REG2_REG_13__SCAN_IN), .A(n6412), .ZN(
        n6937) );
  MUX2_X1 U7167 ( .A(P1_REG2_REG_14__SCAN_IN), .B(n7699), .S(n6939), .Z(n6054)
         );
  INV_X1 U7168 ( .A(n6054), .ZN(n6936) );
  NOR2_X1 U7169 ( .A1(n6937), .A2(n6936), .ZN(n6935) );
  INV_X1 U7170 ( .A(n7369), .ZN(n6194) );
  NOR2_X1 U7171 ( .A1(n6055), .A2(n6194), .ZN(n6056) );
  XNOR2_X1 U7172 ( .A(n6194), .B(n6055), .ZN(n7366) );
  NOR2_X1 U7173 ( .A1(n7365), .A2(n7366), .ZN(n7364) );
  NAND2_X1 U7174 ( .A1(P1_REG2_REG_16__SCAN_IN), .A2(n6063), .ZN(n6057) );
  OAI21_X1 U7175 ( .B1(n6063), .B2(P1_REG2_REG_16__SCAN_IN), .A(n6057), .ZN(
        n7475) );
  NOR2_X1 U7176 ( .A1(n7476), .A2(n7475), .ZN(n7474) );
  NAND2_X1 U7177 ( .A1(n7759), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n6058) );
  OAI21_X1 U7178 ( .B1(n7759), .B2(P1_REG2_REG_17__SCAN_IN), .A(n6058), .ZN(
        n7755) );
  NOR2_X1 U7179 ( .A1(n7756), .A2(n7755), .ZN(n7754) );
  NOR2_X1 U7180 ( .A1(n6059), .A2(n6060), .ZN(n9945) );
  NOR2_X1 U7181 ( .A1(n6089), .A2(P1_U3084), .ZN(n10411) );
  INV_X1 U7182 ( .A(n4855), .ZN(n10407) );
  NAND2_X1 U7183 ( .A1(n10411), .A2(n10407), .ZN(n8083) );
  OR2_X1 U7184 ( .A1(n8083), .A2(n5850), .ZN(n10451) );
  AOI211_X1 U7185 ( .C1(n6060), .C2(n6059), .A(n9945), .B(n10451), .ZN(n6098)
         );
  INV_X1 U7186 ( .A(n5850), .ZN(n6253) );
  OR2_X1 U7187 ( .A1(n8083), .A2(n6253), .ZN(n9952) );
  INV_X1 U7188 ( .A(n9946), .ZN(n6062) );
  NOR2_X1 U7189 ( .A1(n9952), .A2(n6062), .ZN(n6097) );
  NAND2_X1 U7190 ( .A1(n6062), .A2(n6061), .ZN(n9942) );
  OAI21_X1 U7191 ( .B1(n6062), .B2(n6061), .A(n9942), .ZN(n6088) );
  INV_X1 U7192 ( .A(n7759), .ZN(n6086) );
  XNOR2_X1 U7193 ( .A(n7759), .B(n10233), .ZN(n7751) );
  INV_X1 U7194 ( .A(n6063), .ZN(n7473) );
  XOR2_X1 U7195 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n6063), .Z(n7468) );
  INV_X1 U7196 ( .A(n6939), .ZN(n6171) );
  OR2_X1 U7197 ( .A1(n6416), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n6081) );
  INV_X1 U7198 ( .A(n6368), .ZN(n6079) );
  OR2_X1 U7199 ( .A1(n9935), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n6074) );
  MUX2_X1 U7200 ( .A(P1_REG1_REG_10__SCAN_IN), .B(n6064), .S(n9935), .Z(n9928)
         );
  INV_X1 U7201 ( .A(n10434), .ZN(n6145) );
  AOI22_X1 U7202 ( .A1(n10434), .A2(P1_REG1_REG_9__SCAN_IN), .B1(n5584), .B2(
        n6145), .ZN(n10437) );
  NOR2_X1 U7203 ( .A1(P1_REG1_REG_8__SCAN_IN), .A2(n9922), .ZN(n6065) );
  AOI21_X1 U7204 ( .B1(n9922), .B2(P1_REG1_REG_8__SCAN_IN), .A(n6065), .ZN(
        n9915) );
  NAND2_X1 U7205 ( .A1(P1_REG1_REG_5__SCAN_IN), .A2(n6189), .ZN(n6066) );
  OAI21_X1 U7206 ( .B1(n6189), .B2(P1_REG1_REG_5__SCAN_IN), .A(n6066), .ZN(
        n6182) );
  INV_X1 U7207 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n10415) );
  XNOR2_X1 U7208 ( .A(n6114), .B(n6350), .ZN(n10449) );
  NOR3_X1 U7209 ( .A1(n10415), .A2(n10410), .A3(n10449), .ZN(n10448) );
  AOI21_X1 U7210 ( .B1(n10458), .B2(P1_REG1_REG_1__SCAN_IN), .A(n10448), .ZN(
        n6261) );
  NAND2_X1 U7211 ( .A1(P1_REG1_REG_2__SCAN_IN), .A2(n6269), .ZN(n6067) );
  OAI21_X1 U7212 ( .B1(P1_REG1_REG_2__SCAN_IN), .B2(n6269), .A(n6067), .ZN(
        n6260) );
  NOR2_X1 U7213 ( .A1(n6261), .A2(n6260), .ZN(n6259) );
  AND2_X1 U7214 ( .A1(n6269), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n6068) );
  NOR2_X1 U7215 ( .A1(n6259), .A2(n6068), .ZN(n6104) );
  NAND2_X1 U7216 ( .A1(P1_REG1_REG_3__SCAN_IN), .A2(n6105), .ZN(n6069) );
  OAI21_X1 U7217 ( .B1(n6105), .B2(P1_REG1_REG_3__SCAN_IN), .A(n6069), .ZN(
        n6103) );
  NOR2_X1 U7218 ( .A1(n6104), .A2(n6103), .ZN(n6102) );
  AOI21_X1 U7219 ( .B1(n6105), .B2(P1_REG1_REG_3__SCAN_IN), .A(n6102), .ZN(
        n9886) );
  NOR2_X1 U7220 ( .A1(n9895), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n6070) );
  AOI21_X1 U7221 ( .B1(P1_REG1_REG_4__SCAN_IN), .B2(n9895), .A(n6070), .ZN(
        n9885) );
  NAND2_X1 U7222 ( .A1(n9886), .A2(n9885), .ZN(n9884) );
  OAI21_X1 U7223 ( .B1(P1_REG1_REG_4__SCAN_IN), .B2(n9895), .A(n9884), .ZN(
        n6183) );
  NOR2_X1 U7224 ( .A1(n6182), .A2(n6183), .ZN(n6181) );
  AOI21_X1 U7225 ( .B1(n6189), .B2(P1_REG1_REG_5__SCAN_IN), .A(n6181), .ZN(
        n10420) );
  OR2_X1 U7226 ( .A1(n10431), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n6072) );
  NAND2_X1 U7227 ( .A1(n10431), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n6071) );
  NAND2_X1 U7228 ( .A1(n6072), .A2(n6071), .ZN(n10419) );
  NOR2_X1 U7229 ( .A1(n10420), .A2(n10419), .ZN(n10418) );
  AOI21_X1 U7230 ( .B1(P1_REG1_REG_6__SCAN_IN), .B2(n10431), .A(n10418), .ZN(
        n9901) );
  NOR2_X1 U7231 ( .A1(n9908), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n6073) );
  AOI21_X1 U7232 ( .B1(P1_REG1_REG_7__SCAN_IN), .B2(n9908), .A(n6073), .ZN(
        n9900) );
  NAND2_X1 U7233 ( .A1(n9901), .A2(n9900), .ZN(n9899) );
  OAI21_X1 U7234 ( .B1(n9908), .B2(P1_REG1_REG_7__SCAN_IN), .A(n9899), .ZN(
        n9914) );
  NAND2_X1 U7235 ( .A1(n9915), .A2(n9914), .ZN(n9913) );
  OAI21_X1 U7236 ( .B1(P1_REG1_REG_8__SCAN_IN), .B2(n9922), .A(n9913), .ZN(
        n10436) );
  NAND2_X1 U7237 ( .A1(n10437), .A2(n10436), .ZN(n10435) );
  OAI21_X1 U7238 ( .B1(P1_REG1_REG_9__SCAN_IN), .B2(n10434), .A(n10435), .ZN(
        n9929) );
  NAND2_X1 U7239 ( .A1(n9928), .A2(n9929), .ZN(n9927) );
  NAND2_X1 U7240 ( .A1(n6074), .A2(n9927), .ZN(n8092) );
  INV_X1 U7241 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n6076) );
  NAND2_X1 U7242 ( .A1(n8092), .A2(n6076), .ZN(n6075) );
  AND2_X1 U7243 ( .A1(n6075), .A2(n8090), .ZN(n6077) );
  NOR2_X1 U7244 ( .A1(n8092), .A2(n6076), .ZN(n8085) );
  XNOR2_X1 U7245 ( .A(n6368), .B(P1_REG1_REG_12__SCAN_IN), .ZN(n6356) );
  NOR2_X1 U7246 ( .A1(n8091), .A2(n6356), .ZN(n6357) );
  AOI21_X1 U7247 ( .B1(n6079), .B2(n6078), .A(n6357), .ZN(n6418) );
  XNOR2_X1 U7248 ( .A(n6416), .B(P1_REG1_REG_13__SCAN_IN), .ZN(n6419) );
  NOR2_X1 U7249 ( .A1(n6418), .A2(n6419), .ZN(n6417) );
  INV_X1 U7250 ( .A(n6417), .ZN(n6080) );
  XNOR2_X1 U7251 ( .A(n6939), .B(P1_REG1_REG_14__SCAN_IN), .ZN(n6941) );
  NOR2_X1 U7252 ( .A1(n6942), .A2(n6941), .ZN(n6940) );
  AOI21_X1 U7253 ( .B1(n6171), .B2(n6082), .A(n6940), .ZN(n6083) );
  NAND2_X1 U7254 ( .A1(n7369), .A2(n6083), .ZN(n6084) );
  XNOR2_X1 U7255 ( .A(n6194), .B(n6083), .ZN(n7362) );
  NAND2_X1 U7256 ( .A1(P1_REG1_REG_15__SCAN_IN), .A2(n7362), .ZN(n7361) );
  NAND2_X1 U7257 ( .A1(n6084), .A2(n7361), .ZN(n7469) );
  NAND2_X1 U7258 ( .A1(n7468), .A2(n7469), .ZN(n7467) );
  OAI21_X1 U7259 ( .B1(n7473), .B2(n6085), .A(n7467), .ZN(n7750) );
  NAND2_X1 U7260 ( .A1(n7751), .A2(n7750), .ZN(n7749) );
  OAI21_X1 U7261 ( .B1(n6086), .B2(n10233), .A(n7749), .ZN(n6087) );
  NOR2_X1 U7262 ( .A1(n6087), .A2(n6088), .ZN(n9940) );
  AOI21_X1 U7263 ( .B1(n6088), .B2(n6087), .A(n9940), .ZN(n6092) );
  NOR2_X1 U7264 ( .A1(n5850), .A2(P1_U3084), .ZN(n7726) );
  AND2_X1 U7265 ( .A1(n7726), .A2(n4855), .ZN(n6091) );
  INV_X1 U7266 ( .A(n6089), .ZN(n6090) );
  INV_X1 U7267 ( .A(n10443), .ZN(n10447) );
  NOR2_X1 U7268 ( .A1(n6092), .A2(n10447), .ZN(n6096) );
  INV_X1 U7269 ( .A(n6093), .ZN(n6094) );
  INV_X1 U7270 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n10402) );
  NAND2_X1 U7271 ( .A1(P1_U3084), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n9844) );
  OAI21_X1 U7272 ( .B1(n10425), .B2(n10402), .A(n9844), .ZN(n6095) );
  OR4_X1 U7273 ( .A1(n6098), .A2(n6097), .A3(n6096), .A4(n6095), .ZN(P1_U3259)
         );
  INV_X1 U7274 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n6618) );
  NOR2_X1 U7275 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6618), .ZN(n9741) );
  AOI211_X1 U7276 ( .C1(n6101), .C2(n6100), .A(n6099), .B(n10451), .ZN(n6108)
         );
  AOI211_X1 U7277 ( .C1(n6104), .C2(n6103), .A(n6102), .B(n10447), .ZN(n6107)
         );
  INV_X1 U7278 ( .A(n6105), .ZN(n6120) );
  INV_X1 U7279 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n7492) );
  OAI22_X1 U7280 ( .A1(n9952), .A2(n6120), .B1(n10425), .B2(n7492), .ZN(n6106)
         );
  OR4_X1 U7281 ( .A1(n9741), .A2(n6108), .A3(n6107), .A4(n6106), .ZN(P1_U3244)
         );
  NOR2_X2 U7282 ( .A1(n6483), .A2(P1_STATE_REG_SCAN_IN), .ZN(n10324) );
  AOI22_X1 U7283 ( .A1(n10324), .A2(P2_DATAO_REG_2__SCAN_IN), .B1(n6269), .B2(
        P1_STATE_REG_SCAN_IN), .ZN(n6109) );
  OAI21_X1 U7284 ( .B1(n6563), .B2(n6276), .A(n6109), .ZN(P1_U3351) );
  NAND2_X1 U7285 ( .A1(n6483), .A2(P2_U3152), .ZN(n9710) );
  INV_X1 U7286 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n6540) );
  NOR2_X1 U7287 ( .A1(n6110), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9705) );
  INV_X2 U7288 ( .A(n9705), .ZN(n8039) );
  NAND2_X1 U7289 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n6111) );
  INV_X1 U7290 ( .A(n4856), .ZN(n6542) );
  OAI222_X1 U7291 ( .A1(n9710), .A2(n6540), .B1(n8039), .B2(n6541), .C1(
        P2_U3152), .C2(n6542), .ZN(P2_U3357) );
  NAND2_X1 U7292 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(n4876), .ZN(n6112) );
  XNOR2_X1 U7293 ( .A(n6112), .B(P2_IR_REG_2__SCAN_IN), .ZN(n10492) );
  INV_X1 U7294 ( .A(n10492), .ZN(n6567) );
  OAI222_X1 U7295 ( .A1(n9710), .A2(n4956), .B1(n8039), .B2(n6563), .C1(
        P2_U3152), .C2(n6567), .ZN(P2_U3356) );
  INV_X1 U7296 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n6113) );
  INV_X1 U7297 ( .A(n10324), .ZN(n8101) );
  OAI222_X1 U7298 ( .A1(n6276), .A2(n6541), .B1(n6114), .B2(P1_U3084), .C1(
        n6113), .C2(n8101), .ZN(P1_U3352) );
  OAI21_X1 U7299 ( .B1(P2_IR_REG_2__SCAN_IN), .B2(n4876), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n6116) );
  INV_X1 U7300 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n6115) );
  XNOR2_X1 U7301 ( .A(n6116), .B(n6115), .ZN(n6801) );
  INV_X1 U7302 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n6173) );
  OAI222_X1 U7303 ( .A1(n6801), .A2(P2_U3152), .B1(n8039), .B2(n6527), .C1(
        n9710), .C2(n6173), .ZN(P2_U3355) );
  AOI22_X1 U7304 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n9895), .B1(n10324), .B2(
        P2_DATAO_REG_4__SCAN_IN), .ZN(n6117) );
  OAI21_X1 U7305 ( .B1(n6516), .B2(n6276), .A(n6117), .ZN(P1_U3349) );
  INV_X1 U7306 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n6515) );
  OR2_X1 U7307 ( .A1(n6118), .A2(n6162), .ZN(n6119) );
  XNOR2_X1 U7308 ( .A(n6119), .B(P2_IR_REG_4__SCAN_IN), .ZN(n6693) );
  INV_X1 U7309 ( .A(n6693), .ZN(n6825) );
  OAI222_X1 U7310 ( .A1(n9710), .A2(n6515), .B1(n8039), .B2(n6516), .C1(
        P2_U3152), .C2(n6825), .ZN(P2_U3354) );
  INV_X1 U7311 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n6121) );
  OAI222_X1 U7312 ( .A1(n8101), .A2(n6121), .B1(n6276), .B2(n6527), .C1(
        P1_U3084), .C2(n6120), .ZN(P1_U3350) );
  AOI22_X1 U7313 ( .A1(n6189), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_5__SCAN_IN), .B2(n10324), .ZN(n6122) );
  OAI21_X1 U7314 ( .B1(n6482), .B2(n6276), .A(n6122), .ZN(P1_U3348) );
  NAND2_X1 U7315 ( .A1(n6124), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6125) );
  MUX2_X1 U7316 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6125), .S(
        P2_IR_REG_5__SCAN_IN), .Z(n6126) );
  AND2_X1 U7317 ( .A1(n6123), .A2(n6126), .ZN(n6695) );
  INV_X1 U7318 ( .A(n6695), .ZN(n6813) );
  INV_X1 U7319 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n6484) );
  INV_X1 U7320 ( .A(n9710), .ZN(n6273) );
  OAI222_X1 U7321 ( .A1(P2_U3152), .A2(n6813), .B1(n8039), .B2(n6482), .C1(
        n6484), .C2(n8230), .ZN(P2_U3353) );
  INV_X1 U7322 ( .A(n6966), .ZN(n6129) );
  AOI22_X1 U7323 ( .A1(n10431), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_6__SCAN_IN), .B2(n10324), .ZN(n6127) );
  OAI21_X1 U7324 ( .B1(n6129), .B2(n6276), .A(n6127), .ZN(P1_U3347) );
  NAND2_X1 U7325 ( .A1(n6123), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6128) );
  XNOR2_X1 U7326 ( .A(n6128), .B(P2_IR_REG_6__SCAN_IN), .ZN(n6965) );
  INV_X1 U7327 ( .A(n6965), .ZN(n6777) );
  INV_X1 U7328 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n6160) );
  OAI222_X1 U7329 ( .A1(n6777), .A2(P2_U3152), .B1(n8039), .B2(n6129), .C1(
        n9710), .C2(n6160), .ZN(P2_U3352) );
  INV_X1 U7330 ( .A(n6969), .ZN(n6134) );
  AOI22_X1 U7331 ( .A1(n9908), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_7__SCAN_IN), .B2(n10324), .ZN(n6130) );
  OAI21_X1 U7332 ( .B1(n6134), .B2(n6276), .A(n6130), .ZN(P1_U3346) );
  INV_X1 U7333 ( .A(n7158), .ZN(n6141) );
  AOI22_X1 U7334 ( .A1(n9935), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n10324), .ZN(n6131) );
  OAI21_X1 U7335 ( .B1(n6141), .B2(n6276), .A(n6131), .ZN(P1_U3343) );
  OR2_X1 U7336 ( .A1(n6132), .A2(n6162), .ZN(n6133) );
  XNOR2_X1 U7337 ( .A(n6133), .B(P2_IR_REG_7__SCAN_IN), .ZN(n6970) );
  INV_X1 U7338 ( .A(n6970), .ZN(n6789) );
  INV_X1 U7339 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n6169) );
  OAI222_X1 U7340 ( .A1(n6789), .A2(P2_U3152), .B1(n8039), .B2(n6134), .C1(
        n9710), .C2(n6169), .ZN(P2_U3351) );
  INV_X1 U7341 ( .A(n7044), .ZN(n6144) );
  AOI22_X1 U7342 ( .A1(n9922), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(n10324), .ZN(n6135) );
  OAI21_X1 U7343 ( .B1(n6144), .B2(n6276), .A(n6135), .ZN(P1_U3345) );
  INV_X1 U7344 ( .A(n8090), .ZN(n8086) );
  INV_X1 U7345 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n6136) );
  OAI222_X1 U7346 ( .A1(n6276), .A2(n7299), .B1(n8086), .B2(P1_U3084), .C1(
        n6136), .C2(n8101), .ZN(P1_U3342) );
  NAND2_X1 U7347 ( .A1(n6137), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6147) );
  NAND2_X1 U7348 ( .A1(n6147), .A2(n6138), .ZN(n6139) );
  NAND2_X1 U7349 ( .A1(n6139), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6151) );
  XNOR2_X1 U7350 ( .A(n6151), .B(P2_IR_REG_10__SCAN_IN), .ZN(n7159) );
  INV_X1 U7351 ( .A(n7159), .ZN(n6755) );
  INV_X1 U7352 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n6140) );
  OAI222_X1 U7353 ( .A1(P2_U3152), .A2(n6755), .B1(n8039), .B2(n6141), .C1(
        n6140), .C2(n8230), .ZN(P2_U3348) );
  NAND2_X1 U7354 ( .A1(n6142), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6143) );
  XNOR2_X1 U7355 ( .A(n6143), .B(P2_IR_REG_8__SCAN_IN), .ZN(n7045) );
  INV_X1 U7356 ( .A(n7045), .ZN(n6743) );
  INV_X1 U7357 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n6167) );
  OAI222_X1 U7358 ( .A1(n6743), .A2(P2_U3152), .B1(n8039), .B2(n6144), .C1(
        n9710), .C2(n6167), .ZN(P2_U3350) );
  INV_X1 U7359 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n6146) );
  INV_X1 U7360 ( .A(n7105), .ZN(n6149) );
  OAI222_X1 U7361 ( .A1(n8101), .A2(n6146), .B1(n6276), .B2(n6149), .C1(
        P1_U3084), .C2(n6145), .ZN(P1_U3344) );
  XNOR2_X1 U7362 ( .A(n6147), .B(P2_IR_REG_9__SCAN_IN), .ZN(n7106) );
  INV_X1 U7363 ( .A(n7106), .ZN(n6766) );
  INV_X1 U7364 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n6148) );
  OAI222_X1 U7365 ( .A1(n6766), .A2(P2_U3152), .B1(n8039), .B2(n6149), .C1(
        n6148), .C2(n8230), .ZN(P2_U3349) );
  NAND2_X1 U7366 ( .A1(n6151), .A2(n6150), .ZN(n6152) );
  NAND2_X1 U7367 ( .A1(n6152), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6153) );
  XNOR2_X1 U7368 ( .A(n6153), .B(P2_IR_REG_11__SCAN_IN), .ZN(n9048) );
  INV_X1 U7369 ( .A(n9048), .ZN(n6679) );
  INV_X1 U7370 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n6154) );
  OAI222_X1 U7371 ( .A1(P2_U3152), .A2(n6679), .B1(n8039), .B2(n7299), .C1(
        n6154), .C2(n8230), .ZN(P2_U3347) );
  AOI22_X1 U7372 ( .A1(n6368), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(n10324), .ZN(n6155) );
  OAI21_X1 U7373 ( .B1(n7415), .B2(n6276), .A(n6155), .ZN(P1_U3341) );
  OR2_X1 U7374 ( .A1(n6013), .A2(n6162), .ZN(n6156) );
  XNOR2_X1 U7375 ( .A(n6156), .B(P2_IR_REG_12__SCAN_IN), .ZN(n7416) );
  INV_X1 U7376 ( .A(n7416), .ZN(n6850) );
  INV_X1 U7377 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n6157) );
  OAI222_X1 U7378 ( .A1(P2_U3152), .A2(n6850), .B1(n8039), .B2(n7415), .C1(
        n6157), .C2(n8230), .ZN(P2_U3346) );
  NAND2_X1 U7379 ( .A1(n6217), .A2(P1_U4006), .ZN(n6158) );
  OAI21_X1 U7380 ( .B1(P1_U4006), .B2(n5247), .A(n6158), .ZN(P1_U3555) );
  NAND2_X1 U7381 ( .A1(n6629), .A2(P1_U4006), .ZN(n6159) );
  OAI21_X1 U7382 ( .B1(P1_U4006), .B2(n6160), .A(n6159), .ZN(P1_U3561) );
  INV_X1 U7383 ( .A(n7621), .ZN(n6165) );
  AOI22_X1 U7384 ( .A1(n6416), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n10324), .ZN(n6161) );
  OAI21_X1 U7385 ( .B1(n6165), .B2(n6276), .A(n6161), .ZN(P1_U3340) );
  OR2_X1 U7386 ( .A1(n6163), .A2(n6162), .ZN(n6175) );
  XNOR2_X1 U7387 ( .A(n6175), .B(P2_IR_REG_13__SCAN_IN), .ZN(n7622) );
  INV_X1 U7388 ( .A(n7622), .ZN(n7067) );
  INV_X1 U7389 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n6164) );
  OAI222_X1 U7390 ( .A1(n7067), .A2(P2_U3152), .B1(n8039), .B2(n6165), .C1(
        n6164), .C2(n8230), .ZN(P2_U3345) );
  NAND2_X1 U7391 ( .A1(n7087), .A2(P1_U4006), .ZN(n6166) );
  OAI21_X1 U7392 ( .B1(P1_U4006), .B2(n6167), .A(n6166), .ZN(P1_U3563) );
  NAND2_X1 U7393 ( .A1(n6831), .A2(P1_U4006), .ZN(n6168) );
  OAI21_X1 U7394 ( .B1(P1_U4006), .B2(n6169), .A(n6168), .ZN(P1_U3562) );
  INV_X1 U7395 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n6170) );
  OAI222_X1 U7396 ( .A1(n6276), .A2(n7711), .B1(n6171), .B2(P1_U3084), .C1(
        n6170), .C2(n8101), .ZN(P1_U3339) );
  NAND2_X1 U7397 ( .A1(n8055), .A2(P1_U4006), .ZN(n6172) );
  OAI21_X1 U7398 ( .B1(P1_U4006), .B2(n6173), .A(n6172), .ZN(P1_U3558) );
  NAND2_X1 U7399 ( .A1(n6175), .A2(n6174), .ZN(n6176) );
  NAND2_X1 U7400 ( .A1(n6176), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6178) );
  OR2_X1 U7401 ( .A1(n6178), .A2(n6177), .ZN(n6179) );
  NAND2_X1 U7402 ( .A1(n6178), .A2(n6177), .ZN(n6195) );
  INV_X1 U7403 ( .A(n7738), .ZN(n7730) );
  INV_X1 U7404 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n6180) );
  OAI222_X1 U7405 ( .A1(P2_U3152), .A2(n7730), .B1(n8039), .B2(n7711), .C1(
        n6180), .C2(n8230), .ZN(P2_U3344) );
  INV_X1 U7406 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n6192) );
  AOI211_X1 U7407 ( .C1(n6183), .C2(n6182), .A(n6181), .B(n10447), .ZN(n6184)
         );
  AND2_X1 U7408 ( .A1(P1_U3084), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n6603) );
  NOR2_X1 U7409 ( .A1(n6184), .A2(n6603), .ZN(n6191) );
  INV_X1 U7410 ( .A(n10451), .ZN(n9955) );
  OAI21_X1 U7411 ( .B1(n6187), .B2(n6186), .A(n6185), .ZN(n6188) );
  AOI22_X1 U7412 ( .A1(n6189), .A2(n10459), .B1(n9955), .B2(n6188), .ZN(n6190)
         );
  OAI211_X1 U7413 ( .C1(n6192), .C2(n10425), .A(n6191), .B(n6190), .ZN(
        P1_U3246) );
  INV_X1 U7414 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n6193) );
  OAI222_X1 U7415 ( .A1(n6276), .A2(n7789), .B1(n6194), .B2(P1_U3084), .C1(
        n6193), .C2(n8101), .ZN(P1_U3338) );
  NAND2_X1 U7416 ( .A1(n6195), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6196) );
  XNOR2_X1 U7417 ( .A(n6196), .B(P2_IR_REG_15__SCAN_IN), .ZN(n9064) );
  INV_X1 U7418 ( .A(n9064), .ZN(n7739) );
  INV_X1 U7419 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n6197) );
  OAI222_X1 U7420 ( .A1(P2_U3152), .A2(n7739), .B1(n8039), .B2(n7789), .C1(
        n6197), .C2(n8230), .ZN(P2_U3343) );
  NAND2_X1 U7421 ( .A1(n6199), .A2(n6198), .ZN(n6325) );
  INV_X1 U7422 ( .A(n6205), .ZN(n6200) );
  OAI21_X1 U7423 ( .B1(n6222), .B2(n6200), .A(n10145), .ZN(n9851) );
  INV_X1 U7424 ( .A(n9851), .ZN(n9866) );
  NOR2_X1 U7425 ( .A1(n10405), .A2(n8491), .ZN(n8494) );
  INV_X1 U7426 ( .A(n8494), .ZN(n6201) );
  NOR2_X1 U7427 ( .A1(n6325), .A2(n6201), .ZN(n6291) );
  NAND2_X1 U7428 ( .A1(n6291), .A2(n10141), .ZN(n9846) );
  INV_X1 U7429 ( .A(n6325), .ZN(n6209) );
  INV_X1 U7430 ( .A(n6202), .ZN(n6208) );
  INV_X1 U7431 ( .A(n6203), .ZN(n6204) );
  NOR2_X1 U7432 ( .A1(n6205), .A2(n6204), .ZN(n6206) );
  NOR2_X1 U7433 ( .A1(n10405), .A2(n6206), .ZN(n6207) );
  NAND2_X1 U7434 ( .A1(n6325), .A2(n6207), .ZN(n6327) );
  OAI211_X1 U7435 ( .C1(n6209), .C2(n10269), .A(n6208), .B(n6327), .ZN(n8056)
         );
  AOI22_X1 U7436 ( .A1(n9863), .A2(n6277), .B1(n8056), .B2(
        P1_REG3_REG_0__SCAN_IN), .ZN(n6225) );
  AND2_X1 U7437 ( .A1(n5945), .A2(n6210), .ZN(n6211) );
  NAND2_X1 U7438 ( .A1(n6217), .A2(n8212), .ZN(n6215) );
  NOR2_X1 U7439 ( .A1(n6322), .A2(n10415), .ZN(n6213) );
  AOI21_X1 U7440 ( .B1(n6453), .B2(n6216), .A(n6213), .ZN(n6214) );
  NAND2_X1 U7441 ( .A1(n6217), .A2(n6216), .ZN(n6220) );
  NOR2_X1 U7442 ( .A1(n6322), .A2(n10410), .ZN(n6218) );
  AOI21_X1 U7443 ( .B1(n6453), .B2(n8207), .A(n6218), .ZN(n6219) );
  NAND2_X1 U7444 ( .A1(n6220), .A2(n6219), .ZN(n6284) );
  NAND2_X1 U7445 ( .A1(n6221), .A2(n6284), .ZN(n6287) );
  OAI21_X1 U7446 ( .B1(n6221), .B2(n6284), .A(n6287), .ZN(n6255) );
  INV_X1 U7447 ( .A(n6222), .ZN(n6223) );
  NOR2_X1 U7448 ( .A1(n10269), .A2(n8325), .ZN(n6324) );
  NAND2_X1 U7449 ( .A1(n6255), .A2(n9855), .ZN(n6224) );
  OAI211_X1 U7450 ( .C1(n9866), .C2(n6348), .A(n6225), .B(n6224), .ZN(P1_U3230) );
  INV_X1 U7451 ( .A(n7854), .ZN(n6246) );
  NAND2_X1 U7452 ( .A1(n6226), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6227) );
  XNOR2_X1 U7453 ( .A(n6227), .B(P2_IR_REG_16__SCAN_IN), .ZN(n7855) );
  AOI22_X1 U7454 ( .A1(n7855), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_16__SCAN_IN), .B2(n6273), .ZN(n6228) );
  OAI21_X1 U7455 ( .B1(n6246), .B2(n8039), .A(n6228), .ZN(P2_U3342) );
  NAND2_X1 U7456 ( .A1(n6230), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8829) );
  INV_X1 U7457 ( .A(n8829), .ZN(n6236) );
  INV_X1 U7458 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n6231) );
  OAI21_X1 U7459 ( .B1(n10362), .B2(n6236), .A(n7996), .ZN(n6241) );
  NAND2_X1 U7460 ( .A1(n6238), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6239) );
  NAND2_X1 U7461 ( .A1(n10362), .A2(n6499), .ZN(n6240) );
  NOR2_X1 U7462 ( .A1(n10486), .A2(P2_U3966), .ZN(P2_U3151) );
  AOI22_X1 U7463 ( .A1(n7759), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n10324), .ZN(n6242) );
  OAI21_X1 U7464 ( .B1(n7905), .B2(n6276), .A(n6242), .ZN(P1_U3336) );
  NAND2_X1 U7465 ( .A1(n6243), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6244) );
  XNOR2_X1 U7466 ( .A(n6244), .B(P2_IR_REG_17__SCAN_IN), .ZN(n9076) );
  AOI22_X1 U7467 ( .A1(n9076), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_17__SCAN_IN), .B2(n6273), .ZN(n6245) );
  OAI21_X1 U7468 ( .B1(n7905), .B2(n8039), .A(n6245), .ZN(P2_U3341) );
  INV_X1 U7469 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n6247) );
  OAI222_X1 U7470 ( .A1(n8101), .A2(n6247), .B1(n6276), .B2(n6246), .C1(
        P1_U3084), .C2(n7473), .ZN(P1_U3337) );
  INV_X1 U7471 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n6251) );
  AND2_X1 U7472 ( .A1(n6217), .A2(n6348), .ZN(n8451) );
  NOR2_X1 U7473 ( .A1(n8451), .A2(n6344), .ZN(n8336) );
  INV_X1 U7474 ( .A(n8336), .ZN(n6249) );
  AOI22_X1 U7475 ( .A1(n6249), .A2(n6248), .B1(n10141), .B2(n6277), .ZN(n6448)
         );
  OAI21_X1 U7476 ( .B1(n6348), .B2(n6451), .A(n6448), .ZN(n10275) );
  NAND2_X1 U7477 ( .A1(n10275), .A2(n10612), .ZN(n6250) );
  OAI21_X1 U7478 ( .B1(n10612), .B2(n6251), .A(n6250), .ZN(P1_U3454) );
  OR2_X1 U7479 ( .A1(n4855), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n6252) );
  NAND2_X1 U7480 ( .A1(n6253), .A2(n6252), .ZN(n6254) );
  INV_X1 U7481 ( .A(n6254), .ZN(n10406) );
  AND2_X1 U7482 ( .A1(n10406), .A2(P1_IR_REG_0__SCAN_IN), .ZN(n10409) );
  NOR2_X1 U7483 ( .A1(n6255), .A2(n6254), .ZN(n6256) );
  MUX2_X1 U7484 ( .A(n10409), .B(n6256), .S(n4855), .Z(n6257) );
  INV_X1 U7485 ( .A(n6257), .ZN(n6258) );
  OAI211_X1 U7486 ( .C1(P1_IR_REG_0__SCAN_IN), .C2(n10406), .A(n6258), .B(
        P1_U4006), .ZN(n9898) );
  AOI21_X1 U7487 ( .B1(n6261), .B2(n6260), .A(n6259), .ZN(n6262) );
  AOI22_X1 U7488 ( .A1(n10443), .A2(n6262), .B1(P1_REG3_REG_2__SCAN_IN), .B2(
        P1_U3084), .ZN(n6263) );
  OAI21_X1 U7489 ( .B1(n10425), .B2(n7493), .A(n6263), .ZN(n6268) );
  AOI211_X1 U7490 ( .C1(n6266), .C2(n6265), .A(n6264), .B(n10451), .ZN(n6267)
         );
  AOI211_X1 U7491 ( .C1(n10459), .C2(n6269), .A(n6268), .B(n6267), .ZN(n6270)
         );
  NAND2_X1 U7492 ( .A1(n9898), .A2(n6270), .ZN(P1_U3243) );
  INV_X1 U7493 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n7205) );
  NAND2_X1 U7494 ( .A1(n10026), .A2(P1_U4006), .ZN(n6271) );
  OAI21_X1 U7495 ( .B1(n7205), .B2(P1_U4006), .A(n6271), .ZN(P1_U3579) );
  NAND2_X1 U7496 ( .A1(n6272), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6334) );
  XNOR2_X1 U7497 ( .A(n6334), .B(P2_IR_REG_18__SCAN_IN), .ZN(n9088) );
  AOI22_X1 U7498 ( .A1(n9088), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_18__SCAN_IN), .B2(n6273), .ZN(n6274) );
  OAI21_X1 U7499 ( .B1(n7923), .B2(n8039), .A(n6274), .ZN(P2_U3340) );
  AOI22_X1 U7500 ( .A1(n9946), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n10324), .ZN(n6275) );
  OAI21_X1 U7501 ( .B1(n7923), .B2(n6276), .A(n6275), .ZN(P1_U3335) );
  NAND2_X1 U7502 ( .A1(n6277), .A2(n6216), .ZN(n6280) );
  NAND2_X1 U7503 ( .A1(n6278), .A2(n8207), .ZN(n6279) );
  NAND2_X1 U7504 ( .A1(n6280), .A2(n6279), .ZN(n6283) );
  OR2_X2 U7505 ( .A1(n6282), .A2(n6281), .ZN(n6585) );
  INV_X1 U7506 ( .A(n6284), .ZN(n6285) );
  NAND2_X1 U7507 ( .A1(n6285), .A2(n8195), .ZN(n6286) );
  NAND2_X1 U7508 ( .A1(n6277), .A2(n8212), .ZN(n6289) );
  NAND2_X1 U7509 ( .A1(n6278), .A2(n6216), .ZN(n6288) );
  NAND2_X1 U7510 ( .A1(n6289), .A2(n6288), .ZN(n6295) );
  INV_X1 U7511 ( .A(n6295), .ZN(n6300) );
  XNOR2_X1 U7512 ( .A(n6297), .B(n6300), .ZN(n6290) );
  XNOR2_X1 U7513 ( .A(n6299), .B(n6290), .ZN(n6294) );
  NAND2_X1 U7514 ( .A1(n6291), .A2(n10143), .ZN(n9860) );
  AOI22_X1 U7515 ( .A1(n9863), .A2(n9882), .B1(n9848), .B2(n6217), .ZN(n6293)
         );
  AOI22_X1 U7516 ( .A1(n6278), .A2(n9837), .B1(n8056), .B2(
        P1_REG3_REG_1__SCAN_IN), .ZN(n6292) );
  OAI211_X1 U7517 ( .C1(n6294), .C2(n9853), .A(n6293), .B(n6292), .ZN(P1_U3220) );
  INV_X1 U7518 ( .A(n6299), .ZN(n6296) );
  NAND2_X1 U7519 ( .A1(n6296), .A2(n6295), .ZN(n6298) );
  NAND2_X1 U7520 ( .A1(n6298), .A2(n6297), .ZN(n6302) );
  NAND2_X1 U7521 ( .A1(n6300), .A2(n6299), .ZN(n6301) );
  XNOR2_X1 U7522 ( .A(n6304), .B(n8195), .ZN(n6307) );
  OAI22_X1 U7523 ( .A1(n6303), .A2(n6305), .B1(n10519), .B2(n8208), .ZN(n6306)
         );
  XNOR2_X1 U7524 ( .A(n6307), .B(n6306), .ZN(n8054) );
  OR2_X1 U7525 ( .A1(n6307), .A2(n6306), .ZN(n6308) );
  OAI22_X1 U7526 ( .A1(n6879), .A2(n6305), .B1(n6621), .B2(n8208), .ZN(n6311)
         );
  NAND2_X1 U7527 ( .A1(n9737), .A2(n9736), .ZN(n6314) );
  INV_X1 U7528 ( .A(n6310), .ZN(n6312) );
  OR2_X1 U7529 ( .A1(n6312), .A2(n6311), .ZN(n6313) );
  NAND2_X1 U7530 ( .A1(n9881), .A2(n6216), .ZN(n6316) );
  NAND2_X1 U7531 ( .A1(n6890), .A2(n8207), .ZN(n6315) );
  NAND2_X1 U7532 ( .A1(n9881), .A2(n8212), .ZN(n6319) );
  NAND2_X1 U7533 ( .A1(n6890), .A2(n6216), .ZN(n6318) );
  AND2_X1 U7534 ( .A1(n6319), .A2(n6318), .ZN(n6588) );
  XNOR2_X1 U7535 ( .A(n6587), .B(n6588), .ZN(n6320) );
  XNOR2_X1 U7536 ( .A(n6592), .B(n6320), .ZN(n6332) );
  AOI22_X1 U7537 ( .A1(n9863), .A2(n9880), .B1(n9837), .B2(n6890), .ZN(n6331)
         );
  AND2_X1 U7538 ( .A1(P1_U3084), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n9889) );
  NAND3_X1 U7539 ( .A1(n6322), .A2(n7005), .A3(n6321), .ZN(n6323) );
  AOI21_X1 U7540 ( .B1(n6325), .B2(n6324), .A(n6323), .ZN(n6326) );
  OR2_X1 U7541 ( .A1(n6326), .A2(P1_U3084), .ZN(n6328) );
  NAND2_X1 U7542 ( .A1(n6328), .A2(n6327), .ZN(n9783) );
  NOR2_X1 U7543 ( .A1(n9858), .A2(n6883), .ZN(n6329) );
  AOI211_X1 U7544 ( .C1(n9848), .C2(n8055), .A(n9889), .B(n6329), .ZN(n6330)
         );
  OAI211_X1 U7545 ( .C1(n6332), .C2(n9853), .A(n6331), .B(n6330), .ZN(P1_U3228) );
  NAND2_X1 U7546 ( .A1(n6334), .A2(n6333), .ZN(n6335) );
  INV_X1 U7547 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n6336) );
  INV_X1 U7548 ( .A(n7995), .ZN(n6340) );
  INV_X1 U7549 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n6339) );
  OAI222_X1 U7550 ( .A1(n9300), .A2(P2_U3152), .B1(n8039), .B2(n6340), .C1(
        n6339), .C2(n8230), .ZN(P2_U3339) );
  INV_X1 U7551 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n6341) );
  OAI222_X1 U7552 ( .A1(n8101), .A2(n6341), .B1(n6276), .B2(n6340), .C1(n9951), 
        .C2(P1_U3084), .ZN(P1_U3334) );
  OAI21_X1 U7553 ( .B1(n5895), .B2(n6343), .A(n6342), .ZN(n6657) );
  XNOR2_X1 U7554 ( .A(n6345), .B(n6344), .ZN(n6346) );
  AOI222_X1 U7555 ( .A1(n6217), .A2(n10143), .B1(n9882), .B2(n10141), .C1(
        n10140), .C2(n6346), .ZN(n6650) );
  OAI21_X1 U7556 ( .B1(n6347), .B2(n6348), .A(n5984), .ZN(n6349) );
  OR2_X1 U7557 ( .A1(n6349), .A2(n6866), .ZN(n6652) );
  OAI211_X1 U7558 ( .C1(n10240), .C2(n6657), .A(n6650), .B(n6652), .ZN(n6354)
         );
  OAI22_X1 U7559 ( .A1(n10246), .A2(n6347), .B1(n10608), .B2(n6350), .ZN(n6351) );
  AOI21_X1 U7560 ( .B1(n6354), .B2(n10608), .A(n6351), .ZN(n6352) );
  INV_X1 U7561 ( .A(n6352), .ZN(P1_U3524) );
  OAI22_X1 U7562 ( .A1(n10311), .A2(n6347), .B1(n10612), .B2(n5431), .ZN(n6353) );
  AOI21_X1 U7563 ( .B1(n6354), .B2(n10612), .A(n6353), .ZN(n6355) );
  INV_X1 U7564 ( .A(n6355), .ZN(P1_U3457) );
  INV_X1 U7565 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n7518) );
  NAND2_X1 U7566 ( .A1(n6356), .A2(n8091), .ZN(n6359) );
  INV_X1 U7567 ( .A(n6357), .ZN(n6358) );
  NAND2_X1 U7568 ( .A1(n6359), .A2(n6358), .ZN(n6361) );
  NOR2_X1 U7569 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6360), .ZN(n9772) );
  AOI21_X1 U7570 ( .B1(n10443), .B2(n6361), .A(n9772), .ZN(n6362) );
  OAI21_X1 U7571 ( .B1(n10425), .B2(n7518), .A(n6362), .ZN(n6367) );
  AOI211_X1 U7572 ( .C1(n6365), .C2(n6364), .A(n6363), .B(n10451), .ZN(n6366)
         );
  AOI211_X1 U7573 ( .C1(n10459), .C2(n6368), .A(n6367), .B(n6366), .ZN(n6369)
         );
  INV_X1 U7574 ( .A(n6369), .ZN(P1_U3253) );
  INV_X1 U7575 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n6370) );
  OAI222_X1 U7576 ( .A1(n6276), .A2(n8662), .B1(n8440), .B2(P1_U3084), .C1(
        n6370), .C2(n8101), .ZN(P1_U3332) );
  INV_X1 U7577 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n6388) );
  XNOR2_X1 U7578 ( .A(n6373), .B(P2_IR_REG_30__SCAN_IN), .ZN(n6378) );
  NAND2_X1 U7579 ( .A1(n6374), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6375) );
  MUX2_X1 U7580 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6375), .S(
        P2_IR_REG_29__SCAN_IN), .Z(n6377) );
  INV_X1 U7581 ( .A(n6376), .ZN(n9706) );
  AND2_X2 U7582 ( .A1(n6378), .A2(n8038), .ZN(n6555) );
  NAND2_X1 U7583 ( .A1(n6555), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n6386) );
  INV_X1 U7584 ( .A(n6378), .ZN(n8040) );
  NAND2_X1 U7585 ( .A1(n6560), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n6385) );
  NAND2_X1 U7586 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n6493) );
  INV_X1 U7587 ( .A(n6493), .ZN(n6379) );
  NAND2_X1 U7588 ( .A1(n6379), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n6481) );
  INV_X1 U7589 ( .A(n6481), .ZN(n6380) );
  NAND2_X1 U7590 ( .A1(n6380), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n6973) );
  INV_X1 U7591 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n6381) );
  NAND2_X1 U7592 ( .A1(n6481), .A2(n6381), .ZN(n6382) );
  AND2_X1 U7593 ( .A1(n6973), .A2(n6382), .ZN(n8047) );
  NAND2_X1 U7594 ( .A1(n6556), .A2(n8047), .ZN(n6384) );
  NAND2_X1 U7595 ( .A1(n6554), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n6383) );
  NAND4_X1 U7596 ( .A1(n6386), .A2(n6385), .A3(n6384), .A4(n6383), .ZN(n7021)
         );
  NAND2_X1 U7597 ( .A1(P2_U3966), .A2(n7021), .ZN(n6387) );
  OAI21_X1 U7598 ( .B1(n9041), .B2(n6388), .A(n6387), .ZN(P2_U3558) );
  INV_X1 U7599 ( .A(n8000), .ZN(n6411) );
  INV_X1 U7600 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n6389) );
  OAI222_X1 U7601 ( .A1(n6276), .A2(n6411), .B1(P1_U3084), .B2(n8486), .C1(
        n6389), .C2(n8101), .ZN(P1_U3333) );
  INV_X1 U7602 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n7358) );
  INV_X1 U7603 ( .A(n6973), .ZN(n6390) );
  NAND2_X1 U7604 ( .A1(n6390), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n6991) );
  INV_X1 U7605 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n7116) );
  INV_X1 U7606 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n7304) );
  INV_X1 U7607 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n9556) );
  INV_X1 U7608 ( .A(n7715), .ZN(n6394) );
  NAND2_X1 U7609 ( .A1(n6394), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n7793) );
  INV_X1 U7610 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n7792) );
  INV_X1 U7611 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n7926) );
  INV_X1 U7612 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n9557) );
  INV_X1 U7613 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n9575) );
  INV_X1 U7614 ( .A(n8685), .ZN(n6399) );
  AND2_X1 U7615 ( .A1(P2_REG3_REG_24__SCAN_IN), .A2(P2_REG3_REG_23__SCAN_IN), 
        .ZN(n6398) );
  NAND2_X1 U7616 ( .A1(n6399), .A2(n6398), .ZN(n8566) );
  INV_X1 U7617 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n9469) );
  NAND2_X1 U7618 ( .A1(n8566), .A2(n9469), .ZN(n6400) );
  NAND2_X1 U7619 ( .A1(n6607), .A2(n6400), .ZN(n9194) );
  OR2_X1 U7620 ( .A1(n9194), .A2(n7303), .ZN(n6406) );
  INV_X1 U7621 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n6403) );
  NAND2_X1 U7622 ( .A1(n6560), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n6402) );
  NAND2_X1 U7623 ( .A1(n6555), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n6401) );
  OAI211_X1 U7624 ( .C1(n8737), .C2(n6403), .A(n6402), .B(n6401), .ZN(n6404)
         );
  INV_X1 U7625 ( .A(n6404), .ZN(n6405) );
  INV_X1 U7626 ( .A(n9219), .ZN(n8882) );
  NAND2_X1 U7627 ( .A1(n8882), .A2(P2_U3966), .ZN(n6407) );
  OAI21_X1 U7628 ( .B1(n7358), .B2(n9041), .A(n6407), .ZN(P2_U3577) );
  INV_X1 U7629 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n8663) );
  OAI222_X1 U7630 ( .A1(P2_U3152), .A2(n8819), .B1(n8039), .B2(n8662), .C1(
        n8663), .C2(n8230), .ZN(P2_U3337) );
  NAND2_X1 U7631 ( .A1(n6408), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6410) );
  INV_X1 U7632 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n6409) );
  XNOR2_X2 U7633 ( .A(n6410), .B(n6409), .ZN(n6509) );
  INV_X1 U7634 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n8001) );
  INV_X1 U7635 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n6424) );
  AOI211_X1 U7636 ( .C1(n6414), .C2(n6413), .A(n6412), .B(n10451), .ZN(n6415)
         );
  AOI21_X1 U7637 ( .B1(n10459), .B2(n6416), .A(n6415), .ZN(n6423) );
  AOI21_X1 U7638 ( .B1(n6419), .B2(n6418), .A(n6417), .ZN(n6420) );
  NAND2_X1 U7639 ( .A1(P1_U3084), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n7461) );
  OAI21_X1 U7640 ( .B1(n10447), .B2(n6420), .A(n7461), .ZN(n6421) );
  INV_X1 U7641 ( .A(n6421), .ZN(n6422) );
  OAI211_X1 U7642 ( .C1(n6424), .C2(n10425), .A(n6423), .B(n6422), .ZN(
        P1_U3254) );
  OAI21_X1 U7643 ( .B1(n6426), .B2(n8335), .A(n6425), .ZN(n6623) );
  INV_X1 U7644 ( .A(n6623), .ZN(n6433) );
  OAI22_X1 U7645 ( .A1(n6439), .A2(n10103), .B1(n6303), .B2(n10101), .ZN(n6429) );
  XNOR2_X1 U7646 ( .A(n6877), .B(n8335), .ZN(n6427) );
  NOR2_X1 U7647 ( .A1(n6427), .A2(n9997), .ZN(n6428) );
  AOI211_X1 U7648 ( .C1(n6282), .C2(n6623), .A(n6429), .B(n6428), .ZN(n6625)
         );
  INV_X1 U7649 ( .A(n6885), .ZN(n6431) );
  AOI21_X1 U7650 ( .B1(n9740), .B2(n6430), .A(n6431), .ZN(n6617) );
  AOI22_X1 U7651 ( .A1(n6617), .A2(n5984), .B1(n10269), .B2(n9740), .ZN(n6432)
         );
  OAI211_X1 U7652 ( .C1(n6433), .C2(n10273), .A(n6625), .B(n6432), .ZN(n6435)
         );
  NAND2_X1 U7653 ( .A1(n6435), .A2(n10608), .ZN(n6434) );
  OAI21_X1 U7654 ( .B1(n10608), .B2(n5477), .A(n6434), .ZN(P1_U3526) );
  INV_X1 U7655 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n6437) );
  NAND2_X1 U7656 ( .A1(n6435), .A2(n10612), .ZN(n6436) );
  OAI21_X1 U7657 ( .B1(n10612), .B2(n6437), .A(n6436), .ZN(P1_U3463) );
  OAI21_X1 U7658 ( .B1(n6886), .B2(n6664), .A(n5984), .ZN(n6438) );
  NOR2_X1 U7659 ( .A1(n6438), .A2(n6911), .ZN(n6659) );
  NOR2_X1 U7660 ( .A1(n10145), .A2(n6601), .ZN(n6441) );
  XOR2_X1 U7661 ( .A(n6901), .B(n8339), .Z(n6440) );
  OAI222_X1 U7662 ( .A1(n10103), .A2(n6923), .B1(n6440), .B2(n9997), .C1(
        n10101), .C2(n6439), .ZN(n6658) );
  AOI211_X1 U7663 ( .C1(n6659), .C2(n9951), .A(n6441), .B(n6658), .ZN(n6447)
         );
  OR2_X1 U7664 ( .A1(n6443), .A2(n8339), .ZN(n6897) );
  INV_X1 U7665 ( .A(n6897), .ZN(n6442) );
  AOI21_X1 U7666 ( .B1(n8339), .B2(n6443), .A(n6442), .ZN(n6660) );
  INV_X1 U7667 ( .A(n10137), .ZN(n10159) );
  OAI22_X1 U7668 ( .A1(n10115), .A2(n6664), .B1(n10148), .B2(n6444), .ZN(n6445) );
  AOI21_X1 U7669 ( .B1(n6660), .B2(n10159), .A(n6445), .ZN(n6446) );
  OAI21_X1 U7670 ( .B1(n6447), .B2(n10088), .A(n6446), .ZN(P1_U3286) );
  INV_X1 U7671 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n6456) );
  INV_X1 U7672 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n6449) );
  OAI21_X1 U7673 ( .B1(n6449), .B2(n10145), .A(n6448), .ZN(n6450) );
  NAND2_X1 U7674 ( .A1(n6450), .A2(n10148), .ZN(n6455) );
  NOR2_X1 U7675 ( .A1(n6451), .A2(n8491), .ZN(n6452) );
  OAI21_X1 U7676 ( .B1(n10156), .B2(n10097), .A(n6453), .ZN(n6454) );
  OAI211_X1 U7677 ( .C1(n6456), .C2(n10148), .A(n6455), .B(n6454), .ZN(
        P1_U3291) );
  INV_X1 U7678 ( .A(n7206), .ZN(n6458) );
  INV_X1 U7679 ( .A(P2_B_REG_SCAN_IN), .ZN(n6457) );
  AOI22_X1 U7680 ( .A1(P2_B_REG_SCAN_IN), .A2(n6458), .B1(n7206), .B2(n6457), 
        .ZN(n6459) );
  INV_X1 U7681 ( .A(n6471), .ZN(n10361) );
  NAND2_X1 U7682 ( .A1(n7360), .A2(n7585), .ZN(n10360) );
  NOR4_X1 U7683 ( .A1(P2_D_REG_23__SCAN_IN), .A2(P2_D_REG_22__SCAN_IN), .A3(
        P2_D_REG_21__SCAN_IN), .A4(P2_D_REG_20__SCAN_IN), .ZN(n6469) );
  OR4_X1 U7684 ( .A1(P2_D_REG_31__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        P2_D_REG_29__SCAN_IN), .A4(P2_D_REG_28__SCAN_IN), .ZN(n6466) );
  NOR4_X1 U7685 ( .A1(P2_D_REG_15__SCAN_IN), .A2(P2_D_REG_14__SCAN_IN), .A3(
        P2_D_REG_13__SCAN_IN), .A4(P2_D_REG_12__SCAN_IN), .ZN(n6464) );
  NOR4_X1 U7686 ( .A1(P2_D_REG_17__SCAN_IN), .A2(P2_D_REG_19__SCAN_IN), .A3(
        P2_D_REG_18__SCAN_IN), .A4(P2_D_REG_16__SCAN_IN), .ZN(n6463) );
  NOR4_X1 U7687 ( .A1(P2_D_REG_7__SCAN_IN), .A2(P2_D_REG_6__SCAN_IN), .A3(
        P2_D_REG_5__SCAN_IN), .A4(P2_D_REG_2__SCAN_IN), .ZN(n6462) );
  NOR4_X1 U7688 ( .A1(P2_D_REG_11__SCAN_IN), .A2(P2_D_REG_10__SCAN_IN), .A3(
        P2_D_REG_9__SCAN_IN), .A4(P2_D_REG_8__SCAN_IN), .ZN(n6461) );
  NAND4_X1 U7689 ( .A1(n6464), .A2(n6463), .A3(n6462), .A4(n6461), .ZN(n6465)
         );
  NOR4_X1 U7690 ( .A1(P2_D_REG_4__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .A3(
        n6466), .A4(n6465), .ZN(n6468) );
  NOR4_X1 U7691 ( .A1(P2_D_REG_27__SCAN_IN), .A2(P2_D_REG_26__SCAN_IN), .A3(
        P2_D_REG_25__SCAN_IN), .A4(P2_D_REG_24__SCAN_IN), .ZN(n6467) );
  NAND3_X1 U7692 ( .A1(n6469), .A2(n6468), .A3(n6467), .ZN(n6470) );
  AND2_X1 U7693 ( .A1(n6470), .A2(n6471), .ZN(n7002) );
  INV_X1 U7694 ( .A(n7002), .ZN(n6473) );
  INV_X1 U7695 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n10463) );
  NAND2_X1 U7696 ( .A1(n6473), .A2(n7079), .ZN(n6474) );
  NOR2_X1 U7697 ( .A1(n7208), .A2(n6474), .ZN(n6488) );
  INV_X1 U7698 ( .A(n6488), .ZN(n6476) );
  AND2_X1 U7699 ( .A1(n6980), .A2(n9103), .ZN(n6475) );
  NAND2_X1 U7700 ( .A1(n10619), .A2(n8819), .ZN(n7003) );
  NAND2_X1 U7701 ( .A1(n6476), .A2(n7003), .ZN(n6477) );
  NAND2_X1 U7702 ( .A1(n8825), .A2(n6499), .ZN(n7000) );
  NAND2_X1 U7703 ( .A1(n6477), .A2(n7000), .ZN(n6727) );
  NAND2_X1 U7704 ( .A1(n6727), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6479) );
  INV_X1 U7705 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n9668) );
  NAND2_X1 U7706 ( .A1(n6493), .A2(n9668), .ZN(n6480) );
  AND2_X1 U7707 ( .A1(n6481), .A2(n6480), .ZN(n7380) );
  INV_X1 U7708 ( .A(n7380), .ZN(n6584) );
  OR2_X1 U7709 ( .A1(n6564), .A2(n6482), .ZN(n6487) );
  OR2_X1 U7710 ( .A1(n6562), .A2(n6484), .ZN(n6486) );
  OR2_X1 U7711 ( .A1(n6683), .A2(n6813), .ZN(n6485) );
  AND2_X1 U7712 ( .A1(n8762), .A2(n8755), .ZN(n7216) );
  NAND2_X1 U7713 ( .A1(n6491), .A2(n7216), .ZN(n6490) );
  INV_X1 U7714 ( .A(n7003), .ZN(n6489) );
  INV_X1 U7715 ( .A(n8920), .ZN(n6502) );
  INV_X1 U7716 ( .A(n6492), .ZN(n6707) );
  NAND2_X1 U7717 ( .A1(n7021), .A2(n9346), .ZN(n6501) );
  NAND2_X1 U7718 ( .A1(n6555), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n6498) );
  INV_X1 U7719 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n9677) );
  INV_X1 U7720 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n9578) );
  NAND2_X1 U7721 ( .A1(n9677), .A2(n9578), .ZN(n6494) );
  AND2_X1 U7722 ( .A1(n6494), .A2(n6493), .ZN(n7242) );
  NAND2_X1 U7723 ( .A1(n6556), .A2(n7242), .ZN(n6497) );
  NAND2_X1 U7724 ( .A1(n6560), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n6496) );
  NAND2_X1 U7725 ( .A1(n6554), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n6495) );
  NAND4_X1 U7726 ( .A1(n6498), .A2(n6497), .A3(n6496), .A4(n6495), .ZN(n9039)
         );
  NAND2_X1 U7727 ( .A1(n9039), .A2(n9345), .ZN(n6500) );
  AND2_X1 U7728 ( .A1(n6501), .A2(n6500), .ZN(n7373) );
  OAI22_X1 U7729 ( .A1(n6502), .A2(n7373), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9668), .ZN(n6503) );
  AOI21_X1 U7730 ( .B1(n7381), .B2(n9017), .A(n6503), .ZN(n6583) );
  INV_X1 U7731 ( .A(n8825), .ZN(n6504) );
  AND2_X4 U7732 ( .A1(n6504), .A2(n8755), .ZN(n8932) );
  NAND2_X1 U7733 ( .A1(n6554), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n6508) );
  NAND2_X1 U7734 ( .A1(n6556), .A2(n7380), .ZN(n6507) );
  NAND2_X1 U7735 ( .A1(n6560), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n6506) );
  NAND2_X1 U7736 ( .A1(n6555), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n6505) );
  NAND4_X1 U7737 ( .A1(n6508), .A2(n6507), .A3(n6506), .A4(n6505), .ZN(n9038)
         );
  NAND2_X1 U7738 ( .A1(n5116), .A2(n9038), .ZN(n6513) );
  NAND2_X1 U7739 ( .A1(n6510), .A2(n9300), .ZN(n6511) );
  XNOR2_X1 U7740 ( .A(n8931), .B(n10565), .ZN(n6512) );
  NAND2_X1 U7741 ( .A1(n6513), .A2(n6512), .ZN(n7025) );
  OR2_X1 U7742 ( .A1(n6513), .A2(n6512), .ZN(n6514) );
  AND2_X1 U7743 ( .A1(n7025), .A2(n6514), .ZN(n6578) );
  NAND2_X1 U7744 ( .A1(n5116), .A2(n9039), .ZN(n6521) );
  OR2_X1 U7745 ( .A1(n6564), .A2(n6516), .ZN(n6517) );
  OAI211_X1 U7746 ( .C1(n6683), .C2(n6825), .A(n6518), .B(n6517), .ZN(n7247)
         );
  XNOR2_X1 U7747 ( .A(n8931), .B(n6519), .ZN(n6520) );
  NAND2_X1 U7748 ( .A1(n6521), .A2(n6520), .ZN(n6533) );
  OR2_X1 U7749 ( .A1(n6521), .A2(n6520), .ZN(n6522) );
  NAND2_X1 U7750 ( .A1(n6533), .A2(n6522), .ZN(n6720) );
  NAND2_X1 U7751 ( .A1(n6555), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n6526) );
  NAND2_X1 U7752 ( .A1(n6560), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n6525) );
  NAND2_X1 U7753 ( .A1(n6554), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n6524) );
  NAND2_X1 U7754 ( .A1(n6556), .A2(n9578), .ZN(n6523) );
  INV_X1 U7755 ( .A(n6531), .ZN(n6530) );
  OR2_X1 U7756 ( .A1(n6562), .A2(n6173), .ZN(n6529) );
  OR2_X1 U7757 ( .A1(n6564), .A2(n6527), .ZN(n6528) );
  OAI211_X1 U7758 ( .C1(n6683), .C2(n6801), .A(n6529), .B(n6528), .ZN(n8904)
         );
  XNOR2_X1 U7759 ( .A(n8931), .B(n8904), .ZN(n6532) );
  AND2_X1 U7760 ( .A1(n6717), .A2(n6533), .ZN(n6576) );
  INV_X1 U7761 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n6534) );
  OR2_X1 U7762 ( .A1(n6535), .A2(n6534), .ZN(n6539) );
  NAND2_X1 U7763 ( .A1(n6554), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n6538) );
  NAND2_X1 U7764 ( .A1(n6555), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n6537) );
  NAND2_X1 U7765 ( .A1(n6556), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n6536) );
  OR2_X1 U7766 ( .A1(n9321), .A2(n8932), .ZN(n6544) );
  XNOR2_X1 U7767 ( .A(n8931), .B(n10513), .ZN(n6543) );
  NAND2_X1 U7768 ( .A1(n6544), .A2(n6543), .ZN(n6553) );
  NAND2_X1 U7769 ( .A1(n6555), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n6549) );
  NAND2_X1 U7770 ( .A1(n6560), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n6548) );
  NAND2_X1 U7771 ( .A1(n6556), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n6547) );
  NAND2_X1 U7772 ( .A1(n6554), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n6546) );
  NAND4_X1 U7773 ( .A1(n6549), .A2(n6548), .A3(n6547), .A4(n6546), .ZN(n9344)
         );
  NAND2_X1 U7774 ( .A1(n6550), .A2(SI_0_), .ZN(n6551) );
  XNOR2_X1 U7775 ( .A(n6551), .B(P1_DATAO_REG_0__SCAN_IN), .ZN(n9712) );
  MUX2_X1 U7776 ( .A(P2_IR_REG_0__SCAN_IN), .B(n9712), .S(n6683), .Z(n9351) );
  AND2_X1 U7777 ( .A1(n9344), .A2(n9351), .ZN(n9333) );
  NOR2_X1 U7778 ( .A1(n8931), .A2(n9351), .ZN(n6552) );
  AOI21_X1 U7779 ( .B1(n5116), .B2(n9333), .A(n6552), .ZN(n8831) );
  NAND2_X1 U7780 ( .A1(n5229), .A2(n8831), .ZN(n8830) );
  NAND2_X1 U7781 ( .A1(n6554), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n6559) );
  NAND2_X1 U7782 ( .A1(n6555), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n6558) );
  NAND2_X1 U7783 ( .A1(n6556), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n6557) );
  NAND2_X1 U7784 ( .A1(n6560), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n6561) );
  OR2_X1 U7785 ( .A1(n7259), .A2(n8932), .ZN(n6569) );
  OR2_X1 U7786 ( .A1(n6564), .A2(n6563), .ZN(n6565) );
  XNOR2_X1 U7787 ( .A(n8931), .B(n6959), .ZN(n6570) );
  INV_X1 U7788 ( .A(n6569), .ZN(n6572) );
  INV_X1 U7789 ( .A(n6570), .ZN(n6571) );
  NAND2_X1 U7790 ( .A1(n6572), .A2(n6571), .ZN(n8905) );
  AND2_X1 U7791 ( .A1(n8905), .A2(n6573), .ZN(n6714) );
  INV_X1 U7792 ( .A(n6720), .ZN(n6574) );
  AND2_X1 U7793 ( .A1(n6714), .A2(n6574), .ZN(n6575) );
  NAND2_X1 U7794 ( .A1(n8906), .A2(n6575), .ZN(n6718) );
  OAI21_X1 U7795 ( .B1(n6578), .B2(n6577), .A(n7026), .ZN(n6581) );
  NAND2_X1 U7796 ( .A1(n10625), .A2(n6981), .ZN(n6579) );
  NAND2_X1 U7797 ( .A1(n6581), .A2(n8941), .ZN(n6582) );
  OAI211_X1 U7798 ( .C1(n9013), .C2(n6584), .A(n6583), .B(n6582), .ZN(P2_U3229) );
  INV_X1 U7799 ( .A(n6587), .ZN(n6590) );
  INV_X1 U7800 ( .A(n6588), .ZN(n6589) );
  NAND2_X1 U7801 ( .A1(n6590), .A2(n6589), .ZN(n6594) );
  NAND2_X1 U7802 ( .A1(n6638), .A2(n4873), .ZN(n6599) );
  OR2_X1 U7803 ( .A1(n6904), .A2(n6305), .ZN(n6598) );
  NAND2_X1 U7804 ( .A1(n6600), .A2(n6216), .ZN(n6597) );
  AND2_X1 U7805 ( .A1(n6598), .A2(n6597), .ZN(n6637) );
  XNOR2_X1 U7806 ( .A(n6599), .B(n6637), .ZN(n6606) );
  AOI22_X1 U7807 ( .A1(n9863), .A2(n6629), .B1(n9837), .B2(n6600), .ZN(n6605)
         );
  NOR2_X1 U7808 ( .A1(n9858), .A2(n6601), .ZN(n6602) );
  AOI211_X1 U7809 ( .C1(n9848), .C2(n9881), .A(n6603), .B(n6602), .ZN(n6604)
         );
  OAI211_X1 U7810 ( .C1(n6606), .C2(n9853), .A(n6605), .B(n6604), .ZN(P1_U3225) );
  INV_X1 U7811 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n7540) );
  INV_X1 U7812 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n9689) );
  NAND2_X1 U7813 ( .A1(n6607), .A2(n9689), .ZN(n6608) );
  NAND2_X1 U7814 ( .A1(n9188), .A2(n6556), .ZN(n6614) );
  INV_X1 U7815 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n6611) );
  NAND2_X1 U7816 ( .A1(n6560), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n6610) );
  NAND2_X1 U7817 ( .A1(n6555), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n6609) );
  OAI211_X1 U7818 ( .C1(n8737), .C2(n6611), .A(n6610), .B(n6609), .ZN(n6612)
         );
  INV_X1 U7819 ( .A(n6612), .ZN(n6613) );
  INV_X1 U7820 ( .A(n9172), .ZN(n9203) );
  NAND2_X1 U7821 ( .A1(n9203), .A2(n9041), .ZN(n6615) );
  OAI21_X1 U7822 ( .B1(n7540), .B2(P2_U3966), .A(n6615), .ZN(P2_U3578) );
  NAND2_X1 U7823 ( .A1(n10148), .A2(n6616), .ZN(n8526) );
  INV_X1 U7824 ( .A(n8526), .ZN(n7616) );
  NAND2_X1 U7825 ( .A1(n6617), .A2(n10097), .ZN(n6620) );
  AOI22_X1 U7826 ( .A1(n10088), .A2(P1_REG2_REG_3__SCAN_IN), .B1(n10111), .B2(
        n6618), .ZN(n6619) );
  OAI211_X1 U7827 ( .C1(n6621), .C2(n10115), .A(n6620), .B(n6619), .ZN(n6622)
         );
  AOI21_X1 U7828 ( .B1(n6623), .B2(n7616), .A(n6622), .ZN(n6624) );
  OAI21_X1 U7829 ( .B1(n6625), .B2(n10088), .A(n6624), .ZN(P1_U3288) );
  NAND2_X1 U7830 ( .A1(n6629), .A2(n6216), .ZN(n6626) );
  OAI21_X1 U7831 ( .B1(n10574), .B2(n6627), .A(n6626), .ZN(n6628) );
  XNOR2_X1 U7832 ( .A(n6628), .B(n8145), .ZN(n6632) );
  OR2_X1 U7833 ( .A1(n10574), .A2(n8208), .ZN(n6631) );
  NAND2_X1 U7834 ( .A1(n6629), .A2(n8212), .ZN(n6630) );
  AND2_X1 U7835 ( .A1(n6631), .A2(n6630), .ZN(n6633) );
  NAND2_X1 U7836 ( .A1(n6632), .A2(n6633), .ZN(n6832) );
  INV_X1 U7837 ( .A(n6632), .ZN(n6635) );
  INV_X1 U7838 ( .A(n6633), .ZN(n6634) );
  NAND2_X1 U7839 ( .A1(n6635), .A2(n6634), .ZN(n6636) );
  AND2_X1 U7840 ( .A1(n6832), .A2(n6636), .ZN(n6641) );
  NAND2_X1 U7841 ( .A1(n6639), .A2(n6638), .ZN(n6640) );
  NAND2_X1 U7842 ( .A1(n6640), .A2(n6641), .ZN(n6833) );
  OAI21_X1 U7843 ( .B1(n6641), .B2(n6640), .A(n6833), .ZN(n6642) );
  NAND2_X1 U7844 ( .A1(n6642), .A2(n9855), .ZN(n6648) );
  INV_X1 U7845 ( .A(n6908), .ZN(n6646) );
  NOR2_X1 U7846 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6643), .ZN(n10421) );
  AOI21_X1 U7847 ( .B1(n9863), .B2(n6831), .A(n10421), .ZN(n6644) );
  OAI21_X1 U7848 ( .B1(n6904), .B2(n9860), .A(n6644), .ZN(n6645) );
  AOI21_X1 U7849 ( .B1(n6646), .B2(n9783), .A(n6645), .ZN(n6647) );
  OAI211_X1 U7850 ( .C1(n10574), .C2(n9866), .A(n6648), .B(n6647), .ZN(
        P1_U3237) );
  NAND2_X1 U7851 ( .A1(n9041), .A2(n9344), .ZN(n6649) );
  OAI21_X1 U7852 ( .B1(P2_U3966), .B2(n5248), .A(n6649), .ZN(P2_U3552) );
  INV_X1 U7853 ( .A(n6650), .ZN(n6654) );
  OAI22_X1 U7854 ( .A1(n6652), .A2(n10019), .B1(n10145), .B2(n6651), .ZN(n6653) );
  OAI21_X1 U7855 ( .B1(n6654), .B2(n6653), .A(n10148), .ZN(n6656) );
  AOI22_X1 U7856 ( .A1(n10156), .A2(n6278), .B1(P1_REG2_REG_1__SCAN_IN), .B2(
        n10088), .ZN(n6655) );
  OAI211_X1 U7857 ( .C1(n10137), .C2(n6657), .A(n6656), .B(n6655), .ZN(
        P1_U3290) );
  AOI211_X1 U7858 ( .C1(n6660), .C2(n10595), .A(n6659), .B(n6658), .ZN(n6667)
         );
  INV_X1 U7859 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n6661) );
  OAI22_X1 U7860 ( .A1(n10311), .A2(n6664), .B1(n10612), .B2(n6661), .ZN(n6662) );
  INV_X1 U7861 ( .A(n6662), .ZN(n6663) );
  OAI21_X1 U7862 ( .B1(n6667), .B2(n10609), .A(n6663), .ZN(P1_U3469) );
  OAI22_X1 U7863 ( .A1(n10246), .A2(n6664), .B1(n10608), .B2(n5524), .ZN(n6665) );
  INV_X1 U7864 ( .A(n6665), .ZN(n6666) );
  OAI21_X1 U7865 ( .B1(n6667), .B2(n10607), .A(n6666), .ZN(P1_U3528) );
  NAND2_X1 U7866 ( .A1(n10362), .A2(n6981), .ZN(n6668) );
  NAND2_X1 U7867 ( .A1(n6669), .A2(n6668), .ZN(n6685) );
  NAND2_X1 U7868 ( .A1(n6685), .A2(n6683), .ZN(n6670) );
  NAND2_X1 U7869 ( .A1(n6670), .A2(n9022), .ZN(n6708) );
  INV_X1 U7870 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n10629) );
  MUX2_X1 U7871 ( .A(P2_REG1_REG_11__SCAN_IN), .B(n10629), .S(n9048), .Z(n9050) );
  INV_X1 U7872 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n10620) );
  MUX2_X1 U7873 ( .A(P2_REG1_REG_10__SCAN_IN), .B(n10620), .S(n7159), .Z(n6751) );
  INV_X1 U7874 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n7594) );
  MUX2_X1 U7875 ( .A(P2_REG1_REG_9__SCAN_IN), .B(n7594), .S(n7106), .Z(n6762)
         );
  INV_X1 U7876 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n7272) );
  MUX2_X1 U7877 ( .A(P2_REG1_REG_8__SCAN_IN), .B(n7272), .S(n7045), .Z(n6739)
         );
  INV_X1 U7878 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n6678) );
  MUX2_X1 U7879 ( .A(P2_REG1_REG_7__SCAN_IN), .B(n6678), .S(n6970), .Z(n6785)
         );
  INV_X1 U7880 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n10588) );
  MUX2_X1 U7881 ( .A(P2_REG1_REG_6__SCAN_IN), .B(n10588), .S(n6965), .Z(n6773)
         );
  NAND2_X1 U7882 ( .A1(n6695), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n6677) );
  INV_X1 U7883 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n6671) );
  MUX2_X1 U7884 ( .A(P2_REG1_REG_5__SCAN_IN), .B(n6671), .S(n6695), .Z(n6809)
         );
  NAND2_X1 U7885 ( .A1(n6693), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n6676) );
  INV_X1 U7886 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n6672) );
  MUX2_X1 U7887 ( .A(P2_REG1_REG_4__SCAN_IN), .B(n6672), .S(n6693), .Z(n6822)
         );
  INV_X1 U7888 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n10546) );
  MUX2_X1 U7889 ( .A(n10546), .B(P2_REG1_REG_3__SCAN_IN), .S(n6801), .Z(n6797)
         );
  NAND2_X1 U7890 ( .A1(n10492), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n6675) );
  INV_X1 U7891 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n6673) );
  MUX2_X1 U7892 ( .A(P2_REG1_REG_2__SCAN_IN), .B(n6673), .S(n10492), .Z(n10496) );
  NAND2_X1 U7893 ( .A1(n4856), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n6674) );
  MUX2_X1 U7894 ( .A(P2_REG1_REG_1__SCAN_IN), .B(n6534), .S(n4856), .Z(n10481)
         );
  NAND3_X1 U7895 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), 
        .A3(n10481), .ZN(n10480) );
  NAND2_X1 U7896 ( .A1(n6674), .A2(n10480), .ZN(n10497) );
  NAND2_X1 U7897 ( .A1(n10496), .A2(n10497), .ZN(n10494) );
  NAND2_X1 U7898 ( .A1(n6675), .A2(n10494), .ZN(n6798) );
  NAND2_X1 U7899 ( .A1(n6797), .A2(n6798), .ZN(n6796) );
  OAI21_X1 U7900 ( .B1(n6801), .B2(n10546), .A(n6796), .ZN(n6821) );
  NAND2_X1 U7901 ( .A1(n6822), .A2(n6821), .ZN(n6820) );
  NAND2_X1 U7902 ( .A1(n6676), .A2(n6820), .ZN(n6810) );
  NAND2_X1 U7903 ( .A1(n6809), .A2(n6810), .ZN(n6808) );
  NAND2_X1 U7904 ( .A1(n6677), .A2(n6808), .ZN(n6774) );
  NAND2_X1 U7905 ( .A1(n6773), .A2(n6774), .ZN(n6772) );
  OAI21_X1 U7906 ( .B1(n6777), .B2(n10588), .A(n6772), .ZN(n6786) );
  NAND2_X1 U7907 ( .A1(n6785), .A2(n6786), .ZN(n6784) );
  OAI21_X1 U7908 ( .B1(n6789), .B2(n6678), .A(n6784), .ZN(n6740) );
  NAND2_X1 U7909 ( .A1(n6739), .A2(n6740), .ZN(n6738) );
  OAI21_X1 U7910 ( .B1(n6743), .B2(n7272), .A(n6738), .ZN(n6763) );
  NAND2_X1 U7911 ( .A1(n6762), .A2(n6763), .ZN(n6761) );
  OAI21_X1 U7912 ( .B1(n6766), .B2(n7594), .A(n6761), .ZN(n6752) );
  NAND2_X1 U7913 ( .A1(n6751), .A2(n6752), .ZN(n6750) );
  OAI21_X1 U7914 ( .B1(n6755), .B2(n10620), .A(n6750), .ZN(n9051) );
  NAND2_X1 U7915 ( .A1(n9050), .A2(n9051), .ZN(n9049) );
  OAI21_X1 U7916 ( .B1(n6679), .B2(n10629), .A(n9049), .ZN(n6682) );
  INV_X1 U7917 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n6680) );
  MUX2_X1 U7918 ( .A(n6680), .B(P2_REG1_REG_12__SCAN_IN), .S(n7416), .Z(n6681)
         );
  NOR2_X1 U7919 ( .A1(n6681), .A2(n6682), .ZN(n6849) );
  AOI21_X1 U7920 ( .B1(n6682), .B2(n6681), .A(n6849), .ZN(n6687) );
  AND2_X1 U7921 ( .A1(n6683), .A2(n8824), .ZN(n6684) );
  NAND2_X1 U7922 ( .A1(n6685), .A2(n6684), .ZN(n10468) );
  NOR2_X1 U7923 ( .A1(n7304), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7430) );
  AOI21_X1 U7924 ( .B1(n10486), .B2(P2_ADDR_REG_12__SCAN_IN), .A(n7430), .ZN(
        n6686) );
  OAI21_X1 U7925 ( .B1(n6687), .B2(n10468), .A(n6686), .ZN(n6712) );
  INV_X1 U7926 ( .A(n6801), .ZN(n6691) );
  NAND2_X1 U7927 ( .A1(n10478), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n6688) );
  OAI21_X1 U7928 ( .B1(n4856), .B2(P2_REG2_REG_1__SCAN_IN), .A(n6688), .ZN(
        n10475) );
  NAND2_X1 U7929 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), 
        .ZN(n10476) );
  NOR2_X1 U7930 ( .A1(n10475), .A2(n10476), .ZN(n10474) );
  AOI21_X1 U7931 ( .B1(n4856), .B2(P2_REG2_REG_1__SCAN_IN), .A(n10474), .ZN(
        n10490) );
  NAND2_X1 U7932 ( .A1(n10492), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n6689) );
  OAI21_X1 U7933 ( .B1(n10492), .B2(P2_REG2_REG_2__SCAN_IN), .A(n6689), .ZN(
        n10489) );
  NOR2_X1 U7934 ( .A1(n10490), .A2(n10489), .ZN(n10488) );
  INV_X1 U7935 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n6690) );
  MUX2_X1 U7936 ( .A(P2_REG2_REG_3__SCAN_IN), .B(n6690), .S(n6801), .Z(n6793)
         );
  NOR2_X1 U7937 ( .A1(n6794), .A2(n6793), .ZN(n6792) );
  AOI21_X1 U7938 ( .B1(n6691), .B2(P2_REG2_REG_3__SCAN_IN), .A(n6792), .ZN(
        n6818) );
  NAND2_X1 U7939 ( .A1(n6693), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n6692) );
  OAI21_X1 U7940 ( .B1(n6693), .B2(P2_REG2_REG_4__SCAN_IN), .A(n6692), .ZN(
        n6817) );
  NOR2_X1 U7941 ( .A1(n6818), .A2(n6817), .ZN(n6816) );
  AOI21_X1 U7942 ( .B1(n6693), .B2(P2_REG2_REG_4__SCAN_IN), .A(n6816), .ZN(
        n6806) );
  NAND2_X1 U7943 ( .A1(n6695), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n6694) );
  OAI21_X1 U7944 ( .B1(n6695), .B2(P2_REG2_REG_5__SCAN_IN), .A(n6694), .ZN(
        n6805) );
  NOR2_X1 U7945 ( .A1(n6806), .A2(n6805), .ZN(n6804) );
  INV_X1 U7946 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n6696) );
  MUX2_X1 U7947 ( .A(P2_REG2_REG_6__SCAN_IN), .B(n6696), .S(n6965), .Z(n6697)
         );
  INV_X1 U7948 ( .A(n6697), .ZN(n6770) );
  NOR2_X1 U7949 ( .A1(n6771), .A2(n6770), .ZN(n6769) );
  AOI21_X1 U7950 ( .B1(n6965), .B2(P2_REG2_REG_6__SCAN_IN), .A(n6769), .ZN(
        n6782) );
  INV_X1 U7951 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n6698) );
  MUX2_X1 U7952 ( .A(P2_REG2_REG_7__SCAN_IN), .B(n6698), .S(n6970), .Z(n6699)
         );
  INV_X1 U7953 ( .A(n6699), .ZN(n6781) );
  NOR2_X1 U7954 ( .A1(n6782), .A2(n6781), .ZN(n6780) );
  INV_X1 U7955 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n6700) );
  MUX2_X1 U7956 ( .A(P2_REG2_REG_8__SCAN_IN), .B(n6700), .S(n7045), .Z(n6701)
         );
  INV_X1 U7957 ( .A(n6701), .ZN(n6735) );
  NOR2_X1 U7958 ( .A1(n6736), .A2(n6735), .ZN(n6734) );
  AOI21_X1 U7959 ( .B1(n7045), .B2(P2_REG2_REG_8__SCAN_IN), .A(n6734), .ZN(
        n6760) );
  NAND2_X1 U7960 ( .A1(n7106), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n6702) );
  OAI21_X1 U7961 ( .B1(n7106), .B2(P2_REG2_REG_9__SCAN_IN), .A(n6702), .ZN(
        n6759) );
  NOR2_X1 U7962 ( .A1(n6760), .A2(n6759), .ZN(n6758) );
  INV_X1 U7963 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n6703) );
  MUX2_X1 U7964 ( .A(P2_REG2_REG_10__SCAN_IN), .B(n6703), .S(n7159), .Z(n6704)
         );
  INV_X1 U7965 ( .A(n6704), .ZN(n6747) );
  NOR2_X1 U7966 ( .A1(n6748), .A2(n6747), .ZN(n6746) );
  AOI21_X1 U7967 ( .B1(n7159), .B2(P2_REG2_REG_10__SCAN_IN), .A(n6746), .ZN(
        n9044) );
  INV_X1 U7968 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n6705) );
  MUX2_X1 U7969 ( .A(P2_REG2_REG_11__SCAN_IN), .B(n6705), .S(n9048), .Z(n9045)
         );
  NAND2_X1 U7970 ( .A1(n9044), .A2(n9045), .ZN(n9043) );
  OAI21_X1 U7971 ( .B1(n9048), .B2(P2_REG2_REG_11__SCAN_IN), .A(n9043), .ZN(
        n6710) );
  NAND2_X1 U7972 ( .A1(n7416), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n6706) );
  OAI21_X1 U7973 ( .B1(n7416), .B2(P2_REG2_REG_12__SCAN_IN), .A(n6706), .ZN(
        n6709) );
  NOR2_X1 U7974 ( .A1(n6709), .A2(n6710), .ZN(n6844) );
  INV_X1 U7975 ( .A(n8824), .ZN(n9107) );
  AOI211_X1 U7976 ( .C1(n6710), .C2(n6709), .A(n6844), .B(n10487), .ZN(n6711)
         );
  AOI211_X1 U7977 ( .C1(n10493), .C2(n7416), .A(n6712), .B(n6711), .ZN(n6713)
         );
  INV_X1 U7978 ( .A(n6713), .ZN(P2_U3257) );
  NAND2_X1 U7979 ( .A1(n8906), .A2(n6714), .ZN(n6716) );
  AND2_X1 U7980 ( .A1(n6716), .A2(n6715), .ZN(n6721) );
  NAND2_X1 U7981 ( .A1(n6718), .A2(n6717), .ZN(n6719) );
  AOI21_X1 U7982 ( .B1(n6721), .B2(n6720), .A(n6719), .ZN(n6726) );
  NOR2_X1 U7983 ( .A1(n9677), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6819) );
  INV_X1 U7984 ( .A(n6819), .ZN(n6722) );
  OAI21_X1 U7985 ( .B1(n8937), .B2(n6519), .A(n6722), .ZN(n6723) );
  AOI21_X1 U7986 ( .B1(n7242), .B2(n8949), .A(n6723), .ZN(n6725) );
  INV_X1 U7987 ( .A(n9319), .ZN(n9040) );
  AOI22_X1 U7988 ( .A1(n9005), .A2(n9038), .B1(n8947), .B2(n9040), .ZN(n6724)
         );
  OAI211_X1 U7989 ( .C1(n6726), .C2(n9019), .A(n6725), .B(n6724), .ZN(P2_U3232) );
  INV_X1 U7990 ( .A(n10362), .ZN(n8826) );
  NOR2_X1 U7991 ( .A1(n6727), .A2(n8826), .ZN(n8530) );
  INV_X1 U7992 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n6731) );
  INV_X1 U7993 ( .A(n9321), .ZN(n9042) );
  AOI22_X1 U7994 ( .A1(n9351), .A2(n9017), .B1(n9005), .B2(n9042), .ZN(n6730)
         );
  INV_X1 U7995 ( .A(n9344), .ZN(n8836) );
  NAND2_X1 U7996 ( .A1(n8836), .A2(n9351), .ZN(n6984) );
  INV_X1 U7997 ( .A(n6984), .ZN(n9339) );
  INV_X1 U7998 ( .A(n9351), .ZN(n10502) );
  NAND2_X1 U7999 ( .A1(n9344), .A2(n10502), .ZN(n8578) );
  INV_X1 U8000 ( .A(n8578), .ZN(n7207) );
  MUX2_X1 U8001 ( .A(n7207), .B(n9351), .S(n8932), .Z(n6728) );
  OAI21_X1 U8002 ( .B1(n9339), .B2(n6728), .A(n8941), .ZN(n6729) );
  OAI211_X1 U8003 ( .C1(n8530), .C2(n6731), .A(n6730), .B(n6729), .ZN(P2_U3234) );
  INV_X1 U8004 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n6732) );
  INV_X1 U8005 ( .A(n8671), .ZN(n6733) );
  OAI222_X1 U8006 ( .A1(n8101), .A2(n6732), .B1(n6276), .B2(n6733), .C1(
        P1_U3084), .C2(n5945), .ZN(P1_U3331) );
  INV_X1 U8007 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n8672) );
  OAI222_X1 U8008 ( .A1(n6980), .A2(P2_U3152), .B1(n8039), .B2(n6733), .C1(
        n8672), .C2(n8230), .ZN(P2_U3336) );
  AOI211_X1 U8009 ( .C1(n6736), .C2(n6735), .A(n6734), .B(n10487), .ZN(n6745)
         );
  NOR2_X1 U8010 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6990), .ZN(n6737) );
  AOI21_X1 U8011 ( .B1(n10486), .B2(P2_ADDR_REG_8__SCAN_IN), .A(n6737), .ZN(
        n6742) );
  OAI211_X1 U8012 ( .C1(n6740), .C2(n6739), .A(n10495), .B(n6738), .ZN(n6741)
         );
  OAI211_X1 U8013 ( .C1(n10467), .C2(n6743), .A(n6742), .B(n6741), .ZN(n6744)
         );
  OR2_X1 U8014 ( .A1(n6745), .A2(n6744), .ZN(P2_U3253) );
  AOI211_X1 U8015 ( .C1(n6748), .C2(n6747), .A(n6746), .B(n10487), .ZN(n6757)
         );
  NOR2_X1 U8016 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7116), .ZN(n6749) );
  AOI21_X1 U8017 ( .B1(n10486), .B2(P2_ADDR_REG_10__SCAN_IN), .A(n6749), .ZN(
        n6754) );
  OAI211_X1 U8018 ( .C1(n6752), .C2(n6751), .A(n10495), .B(n6750), .ZN(n6753)
         );
  OAI211_X1 U8019 ( .C1(n10467), .C2(n6755), .A(n6754), .B(n6753), .ZN(n6756)
         );
  OR2_X1 U8020 ( .A1(n6757), .A2(n6756), .ZN(P2_U3255) );
  AOI211_X1 U8021 ( .C1(n6760), .C2(n6759), .A(n6758), .B(n10487), .ZN(n6768)
         );
  INV_X1 U8022 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n9679) );
  NOR2_X1 U8023 ( .A1(n9679), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7123) );
  AOI21_X1 U8024 ( .B1(n10486), .B2(P2_ADDR_REG_9__SCAN_IN), .A(n7123), .ZN(
        n6765) );
  OAI211_X1 U8025 ( .C1(n6763), .C2(n6762), .A(n10495), .B(n6761), .ZN(n6764)
         );
  OAI211_X1 U8026 ( .C1(n10467), .C2(n6766), .A(n6765), .B(n6764), .ZN(n6767)
         );
  OR2_X1 U8027 ( .A1(n6768), .A2(n6767), .ZN(P2_U3254) );
  AOI211_X1 U8028 ( .C1(n6771), .C2(n6770), .A(n6769), .B(n10487), .ZN(n6779)
         );
  NOR2_X1 U8029 ( .A1(n6381), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7029) );
  AOI21_X1 U8030 ( .B1(n10486), .B2(P2_ADDR_REG_6__SCAN_IN), .A(n7029), .ZN(
        n6776) );
  OAI211_X1 U8031 ( .C1(n6774), .C2(n6773), .A(n10495), .B(n6772), .ZN(n6775)
         );
  OAI211_X1 U8032 ( .C1(n10467), .C2(n6777), .A(n6776), .B(n6775), .ZN(n6778)
         );
  OR2_X1 U8033 ( .A1(n6779), .A2(n6778), .ZN(P2_U3251) );
  AOI211_X1 U8034 ( .C1(n6782), .C2(n6781), .A(n6780), .B(n10487), .ZN(n6791)
         );
  INV_X1 U8035 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n9649) );
  NOR2_X1 U8036 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9649), .ZN(n6783) );
  AOI21_X1 U8037 ( .B1(n10486), .B2(P2_ADDR_REG_7__SCAN_IN), .A(n6783), .ZN(
        n6788) );
  OAI211_X1 U8038 ( .C1(n6786), .C2(n6785), .A(n10495), .B(n6784), .ZN(n6787)
         );
  OAI211_X1 U8039 ( .C1(n10467), .C2(n6789), .A(n6788), .B(n6787), .ZN(n6790)
         );
  OR2_X1 U8040 ( .A1(n6791), .A2(n6790), .ZN(P2_U3252) );
  AOI211_X1 U8041 ( .C1(n6794), .C2(n6793), .A(n6792), .B(n10487), .ZN(n6803)
         );
  NOR2_X1 U8042 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9578), .ZN(n6795) );
  AOI21_X1 U8043 ( .B1(n10486), .B2(P2_ADDR_REG_3__SCAN_IN), .A(n6795), .ZN(
        n6800) );
  OAI211_X1 U8044 ( .C1(n6798), .C2(n6797), .A(n10495), .B(n6796), .ZN(n6799)
         );
  OAI211_X1 U8045 ( .C1(n10467), .C2(n6801), .A(n6800), .B(n6799), .ZN(n6802)
         );
  OR2_X1 U8046 ( .A1(n6803), .A2(n6802), .ZN(P2_U3248) );
  AOI211_X1 U8047 ( .C1(n6806), .C2(n6805), .A(n6804), .B(n10487), .ZN(n6815)
         );
  NOR2_X1 U8048 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9668), .ZN(n6807) );
  AOI21_X1 U8049 ( .B1(n10486), .B2(P2_ADDR_REG_5__SCAN_IN), .A(n6807), .ZN(
        n6812) );
  OAI211_X1 U8050 ( .C1(n6810), .C2(n6809), .A(n10495), .B(n6808), .ZN(n6811)
         );
  OAI211_X1 U8051 ( .C1(n10467), .C2(n6813), .A(n6812), .B(n6811), .ZN(n6814)
         );
  OR2_X1 U8052 ( .A1(n6815), .A2(n6814), .ZN(P2_U3250) );
  AOI211_X1 U8053 ( .C1(n6818), .C2(n6817), .A(n6816), .B(n10487), .ZN(n6827)
         );
  AOI21_X1 U8054 ( .B1(n10486), .B2(P2_ADDR_REG_4__SCAN_IN), .A(n6819), .ZN(
        n6824) );
  OAI211_X1 U8055 ( .C1(n6822), .C2(n6821), .A(n10495), .B(n6820), .ZN(n6823)
         );
  OAI211_X1 U8056 ( .C1(n10467), .C2(n6825), .A(n6824), .B(n6823), .ZN(n6826)
         );
  OR2_X1 U8057 ( .A1(n6827), .A2(n6826), .ZN(P2_U3249) );
  NAND2_X1 U8058 ( .A1(n7016), .A2(n8207), .ZN(n6829) );
  OR2_X1 U8059 ( .A1(n7150), .A2(n8208), .ZN(n6828) );
  NAND2_X1 U8060 ( .A1(n6829), .A2(n6828), .ZN(n6830) );
  XNOR2_X1 U8061 ( .A(n6830), .B(n8195), .ZN(n7130) );
  AOI22_X1 U8062 ( .A1(n7016), .A2(n6216), .B1(n6831), .B2(n8212), .ZN(n7131)
         );
  XNOR2_X1 U8063 ( .A(n7130), .B(n7131), .ZN(n6835) );
  NAND2_X1 U8064 ( .A1(n6833), .A2(n6832), .ZN(n6834) );
  OAI21_X1 U8065 ( .B1(n6835), .B2(n6834), .A(n7134), .ZN(n6836) );
  NAND2_X1 U8066 ( .A1(n6836), .A2(n9855), .ZN(n6843) );
  INV_X1 U8067 ( .A(n6928), .ZN(n6841) );
  OR2_X1 U8068 ( .A1(n9846), .A2(n7181), .ZN(n6838) );
  AND2_X1 U8069 ( .A1(P1_U3084), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n9903) );
  INV_X1 U8070 ( .A(n9903), .ZN(n6837) );
  OAI211_X1 U8071 ( .C1(n9860), .C2(n6923), .A(n6838), .B(n6837), .ZN(n6840)
         );
  NOR2_X1 U8072 ( .A1(n9866), .A2(n5027), .ZN(n6839) );
  AOI211_X1 U8073 ( .C1(n6841), .C2(n9783), .A(n6840), .B(n6839), .ZN(n6842)
         );
  NAND2_X1 U8074 ( .A1(n6843), .A2(n6842), .ZN(P1_U3211) );
  INV_X1 U8075 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n6845) );
  AOI22_X1 U8076 ( .A1(n7622), .A2(P2_REG2_REG_13__SCAN_IN), .B1(n6845), .B2(
        n7067), .ZN(n6846) );
  NAND2_X1 U8077 ( .A1(n6847), .A2(n6846), .ZN(n7071) );
  OAI21_X1 U8078 ( .B1(n6847), .B2(n6846), .A(n7071), .ZN(n6856) );
  INV_X1 U8079 ( .A(n10487), .ZN(n10466) );
  INV_X1 U8080 ( .A(n10486), .ZN(n9080) );
  INV_X1 U8081 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n7521) );
  NAND2_X1 U8082 ( .A1(n10493), .A2(n7622), .ZN(n6848) );
  NAND2_X1 U8083 ( .A1(P2_REG3_REG_13__SCAN_IN), .A2(P2_U3152), .ZN(n7632) );
  OAI211_X1 U8084 ( .C1(n9080), .C2(n7521), .A(n6848), .B(n7632), .ZN(n6855)
         );
  AOI21_X1 U8085 ( .B1(n6850), .B2(n6680), .A(n6849), .ZN(n6852) );
  INV_X1 U8086 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n7066) );
  AOI22_X1 U8087 ( .A1(n7622), .A2(n7066), .B1(P2_REG1_REG_13__SCAN_IN), .B2(
        n7067), .ZN(n6851) );
  NOR2_X1 U8088 ( .A1(n6852), .A2(n6851), .ZN(n7065) );
  AOI21_X1 U8089 ( .B1(n6852), .B2(n6851), .A(n7065), .ZN(n6853) );
  NOR2_X1 U8090 ( .A1(n6853), .A2(n10468), .ZN(n6854) );
  AOI211_X1 U8091 ( .C1(n6856), .C2(n10466), .A(n6855), .B(n6854), .ZN(n6857)
         );
  INV_X1 U8092 ( .A(n6857), .ZN(P2_U3258) );
  OAI21_X1 U8093 ( .B1(n6859), .B2(n6860), .A(n6858), .ZN(n10523) );
  INV_X1 U8094 ( .A(n10523), .ZN(n6872) );
  XNOR2_X1 U8095 ( .A(n6860), .B(n8460), .ZN(n6864) );
  OAI22_X1 U8096 ( .A1(n6861), .A2(n10101), .B1(n6879), .B2(n10103), .ZN(n6862) );
  AOI21_X1 U8097 ( .B1(n10523), .B2(n6282), .A(n6862), .ZN(n6863) );
  OAI21_X1 U8098 ( .B1(n9997), .B2(n6864), .A(n6863), .ZN(n10521) );
  NAND2_X1 U8099 ( .A1(n10521), .A2(n10148), .ZN(n6871) );
  INV_X1 U8100 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n6865) );
  OAI22_X1 U8101 ( .A1(n10148), .A2(n6865), .B1(n5454), .B2(n10145), .ZN(n6869) );
  OR2_X1 U8102 ( .A1(n6866), .A2(n10519), .ZN(n6867) );
  NAND2_X1 U8103 ( .A1(n6430), .A2(n6867), .ZN(n10520) );
  NOR2_X1 U8104 ( .A1(n10152), .A2(n10520), .ZN(n6868) );
  AOI211_X1 U8105 ( .C1(n10156), .C2(n8057), .A(n6869), .B(n6868), .ZN(n6870)
         );
  OAI211_X1 U8106 ( .C1(n6872), .C2(n8526), .A(n6871), .B(n6870), .ZN(P1_U3289) );
  OAI21_X1 U8107 ( .B1(n6874), .B2(n8341), .A(n6873), .ZN(n10553) );
  INV_X1 U8108 ( .A(n10553), .ZN(n6893) );
  OAI21_X1 U8109 ( .B1(n6877), .B2(n6876), .A(n6875), .ZN(n6878) );
  XOR2_X1 U8110 ( .A(n8341), .B(n6878), .Z(n6882) );
  OAI22_X1 U8111 ( .A1(n6879), .A2(n10101), .B1(n6904), .B2(n10103), .ZN(n6880) );
  AOI21_X1 U8112 ( .B1(n10553), .B2(n6282), .A(n6880), .ZN(n6881) );
  OAI21_X1 U8113 ( .B1(n9997), .B2(n6882), .A(n6881), .ZN(n10551) );
  NAND2_X1 U8114 ( .A1(n10551), .A2(n10148), .ZN(n6892) );
  OAI22_X1 U8115 ( .A1(n10148), .A2(n6884), .B1(n6883), .B2(n10145), .ZN(n6889) );
  AND2_X1 U8116 ( .A1(n6885), .A2(n6890), .ZN(n6887) );
  OR2_X1 U8117 ( .A1(n6887), .A2(n6886), .ZN(n10550) );
  NOR2_X1 U8118 ( .A1(n10550), .A2(n10152), .ZN(n6888) );
  AOI211_X1 U8119 ( .C1(n10156), .C2(n6890), .A(n6889), .B(n6888), .ZN(n6891)
         );
  OAI211_X1 U8120 ( .C1(n6893), .C2(n8526), .A(n6892), .B(n6891), .ZN(P1_U3287) );
  NAND2_X1 U8121 ( .A1(n6897), .A2(n6895), .ZN(n6899) );
  AND2_X1 U8122 ( .A1(n6897), .A2(n6896), .ZN(n6898) );
  AOI21_X1 U8123 ( .B1(n8244), .B2(n6899), .A(n6898), .ZN(n10573) );
  INV_X1 U8124 ( .A(n6282), .ZN(n6927) );
  NAND2_X1 U8125 ( .A1(n6901), .A2(n6900), .ZN(n6903) );
  XNOR2_X1 U8126 ( .A(n8367), .B(n8244), .ZN(n6906) );
  OAI22_X1 U8127 ( .A1(n6904), .A2(n10101), .B1(n7150), .B2(n10103), .ZN(n6905) );
  AOI21_X1 U8128 ( .B1(n6906), .B2(n10140), .A(n6905), .ZN(n6907) );
  OAI21_X1 U8129 ( .B1(n10573), .B2(n6927), .A(n6907), .ZN(n10576) );
  NAND2_X1 U8130 ( .A1(n10576), .A2(n10148), .ZN(n6917) );
  OAI22_X1 U8131 ( .A1(n10148), .A2(n6909), .B1(n6908), .B2(n10145), .ZN(n6914) );
  OR2_X1 U8132 ( .A1(n6911), .A2(n10574), .ZN(n6912) );
  NAND2_X1 U8133 ( .A1(n6910), .A2(n6912), .ZN(n10575) );
  NOR2_X1 U8134 ( .A1(n10575), .A2(n10152), .ZN(n6913) );
  AOI211_X1 U8135 ( .C1(n10156), .C2(n6915), .A(n6914), .B(n6913), .ZN(n6916)
         );
  OAI211_X1 U8136 ( .C1(n10573), .C2(n8526), .A(n6917), .B(n6916), .ZN(
        P1_U3285) );
  OAI21_X1 U8137 ( .B1(n6920), .B2(n6919), .A(n6918), .ZN(n7010) );
  INV_X1 U8138 ( .A(n7010), .ZN(n6934) );
  OAI21_X1 U8139 ( .B1(n8342), .B2(n6922), .A(n6921), .ZN(n6925) );
  OAI22_X1 U8140 ( .A1(n6923), .A2(n10101), .B1(n7181), .B2(n10103), .ZN(n6924) );
  AOI21_X1 U8141 ( .B1(n6925), .B2(n10140), .A(n6924), .ZN(n6926) );
  OAI21_X1 U8142 ( .B1(n6934), .B2(n6927), .A(n6926), .ZN(n7008) );
  NAND2_X1 U8143 ( .A1(n7008), .A2(n10148), .ZN(n6933) );
  AOI211_X1 U8144 ( .C1(n7016), .C2(n6910), .A(n10591), .B(n4909), .ZN(n7009)
         );
  NOR2_X1 U8145 ( .A1(n5027), .A2(n10115), .ZN(n6931) );
  OAI22_X1 U8146 ( .A1(n10148), .A2(n6929), .B1(n6928), .B2(n10145), .ZN(n6930) );
  AOI211_X1 U8147 ( .C1(n7009), .C2(n10110), .A(n6931), .B(n6930), .ZN(n6932)
         );
  OAI211_X1 U8148 ( .C1(n6934), .C2(n8526), .A(n6933), .B(n6932), .ZN(P1_U3284) );
  INV_X1 U8149 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n7524) );
  AOI211_X1 U8150 ( .C1(n6937), .C2(n6936), .A(n6935), .B(n10451), .ZN(n6938)
         );
  AOI21_X1 U8151 ( .B1(n10459), .B2(n6939), .A(n6938), .ZN(n6946) );
  AOI21_X1 U8152 ( .B1(n6942), .B2(n6941), .A(n6940), .ZN(n6943) );
  NAND2_X1 U8153 ( .A1(P1_U3084), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n7552) );
  OAI21_X1 U8154 ( .B1(n10447), .B2(n6943), .A(n7552), .ZN(n6944) );
  INV_X1 U8155 ( .A(n6944), .ZN(n6945) );
  OAI211_X1 U8156 ( .C1(n7524), .C2(n10425), .A(n6946), .B(n6945), .ZN(
        P1_U3255) );
  INV_X1 U8157 ( .A(n6947), .ZN(n6948) );
  AOI21_X1 U8158 ( .B1(n8344), .B2(n6949), .A(n6948), .ZN(n10596) );
  INV_X1 U8159 ( .A(n10596), .ZN(n6957) );
  XOR2_X1 U8160 ( .A(n8344), .B(n6950), .Z(n6951) );
  OAI222_X1 U8161 ( .A1(n10103), .A2(n8068), .B1(n6951), .B2(n9997), .C1(
        n10101), .C2(n7150), .ZN(n10594) );
  INV_X1 U8162 ( .A(n7091), .ZN(n7092) );
  OAI21_X1 U8163 ( .B1(n5026), .B2(n4909), .A(n7092), .ZN(n10592) );
  OAI22_X1 U8164 ( .A1(n10148), .A2(n6952), .B1(n7146), .B2(n10145), .ZN(n6953) );
  AOI21_X1 U8165 ( .B1(n7138), .B2(n10156), .A(n6953), .ZN(n6954) );
  OAI21_X1 U8166 ( .B1(n10592), .B2(n10152), .A(n6954), .ZN(n6955) );
  AOI21_X1 U8167 ( .B1(n10594), .B2(n10148), .A(n6955), .ZN(n6956) );
  OAI21_X1 U8168 ( .B1(n6957), .B2(n10137), .A(n6956), .ZN(P1_U3283) );
  NAND2_X1 U8169 ( .A1(n9321), .A2(n9352), .ZN(n8579) );
  NAND2_X1 U8170 ( .A1(n9338), .A2(n8579), .ZN(n9332) );
  NAND2_X1 U8171 ( .A1(n9332), .A2(n9333), .ZN(n9335) );
  NAND2_X1 U8172 ( .A1(n9042), .A2(n9352), .ZN(n6958) );
  NAND2_X1 U8173 ( .A1(n9335), .A2(n6958), .ZN(n9312) );
  NAND2_X1 U8174 ( .A1(n7259), .A2(n6959), .ZN(n6960) );
  OAI21_X1 U8175 ( .B1(n9312), .B2(n9316), .A(n6960), .ZN(n7250) );
  NAND2_X1 U8176 ( .A1(n9319), .A2(n8904), .ZN(n8589) );
  NAND2_X1 U8177 ( .A1(n9040), .A2(n10539), .ZN(n8588) );
  NAND2_X1 U8178 ( .A1(n8589), .A2(n8588), .ZN(n7251) );
  NAND2_X1 U8179 ( .A1(n7250), .A2(n7251), .ZN(n6962) );
  NAND2_X1 U8180 ( .A1(n9319), .A2(n10539), .ZN(n6961) );
  NAND2_X1 U8181 ( .A1(n6962), .A2(n6961), .ZN(n7237) );
  NOR2_X1 U8182 ( .A1(n9039), .A2(n7247), .ZN(n6964) );
  NAND2_X1 U8183 ( .A1(n9039), .A2(n7247), .ZN(n6963) );
  INV_X1 U8184 ( .A(n9038), .ZN(n7032) );
  AOI22_X1 U8185 ( .A1(n7997), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n7996), .B2(
        n6965), .ZN(n6968) );
  NAND2_X1 U8186 ( .A1(n6966), .A2(n8727), .ZN(n6967) );
  NAND2_X1 U8187 ( .A1(n6968), .A2(n6967), .ZN(n8050) );
  INV_X1 U8188 ( .A(n7021), .ZN(n7060) );
  NAND2_X1 U8189 ( .A1(n6969), .A2(n8727), .ZN(n6972) );
  AOI22_X1 U8190 ( .A1(n7997), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n7996), .B2(
        n6970), .ZN(n6971) );
  NAND2_X1 U8191 ( .A1(n6555), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n6978) );
  NAND2_X1 U8192 ( .A1(n6560), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n6977) );
  NAND2_X1 U8193 ( .A1(n6973), .A2(n9649), .ZN(n6974) );
  AND2_X1 U8194 ( .A1(n6991), .A2(n6974), .ZN(n7277) );
  NAND2_X1 U8195 ( .A1(n6556), .A2(n7277), .ZN(n6976) );
  NAND2_X1 U8196 ( .A1(n6554), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n6975) );
  NAND4_X1 U8197 ( .A1(n6978), .A2(n6977), .A3(n6976), .A4(n6975), .ZN(n9037)
         );
  NAND2_X1 U8198 ( .A1(n7280), .A2(n9037), .ZN(n8610) );
  INV_X1 U8199 ( .A(n7280), .ZN(n6979) );
  NAND2_X1 U8200 ( .A1(n7220), .A2(n6979), .ZN(n8618) );
  XNOR2_X1 U8201 ( .A(n7222), .B(n8768), .ZN(n7284) );
  NAND2_X1 U8202 ( .A1(n7212), .A2(n6980), .ZN(n6983) );
  AND2_X1 U8203 ( .A1(n6981), .A2(n9300), .ZN(n6982) );
  NAND2_X1 U8204 ( .A1(n6983), .A2(n6982), .ZN(n9302) );
  INV_X1 U8205 ( .A(n10619), .ZN(n7591) );
  OAI21_X1 U8206 ( .B1(n8046), .B2(n7280), .A(n7230), .ZN(n7276) );
  INV_X1 U8207 ( .A(n8755), .ZN(n10501) );
  OAI22_X1 U8208 ( .A1(n7276), .A2(n10637), .B1(n7280), .B2(n10625), .ZN(n6999) );
  NAND2_X1 U8209 ( .A1(n6984), .A2(n8579), .ZN(n9343) );
  NAND2_X1 U8210 ( .A1(n9343), .A2(n9338), .ZN(n9317) );
  INV_X1 U8211 ( .A(n8585), .ZN(n6985) );
  OAI21_X1 U8212 ( .B1(n9317), .B2(n6985), .A(n8584), .ZN(n7257) );
  INV_X1 U8213 ( .A(n7251), .ZN(n8761) );
  NAND2_X1 U8214 ( .A1(n9039), .A2(n6519), .ZN(n8595) );
  NAND2_X1 U8215 ( .A1(n7032), .A2(n7381), .ZN(n8599) );
  NAND2_X1 U8216 ( .A1(n9038), .A2(n10565), .ZN(n8598) );
  INV_X1 U8217 ( .A(n8598), .ZN(n6986) );
  NAND2_X1 U8218 ( .A1(n7021), .A2(n10582), .ZN(n8602) );
  NAND2_X1 U8219 ( .A1(n8042), .A2(n8602), .ZN(n6987) );
  NAND2_X1 U8220 ( .A1(n7060), .A2(n8050), .ZN(n8603) );
  NAND2_X1 U8221 ( .A1(n6987), .A2(n8603), .ZN(n6988) );
  NAND2_X1 U8222 ( .A1(n6988), .A2(n8768), .ZN(n7226) );
  OAI21_X1 U8223 ( .B1(n8768), .B2(n6988), .A(n7226), .ZN(n6989) );
  OR2_X1 U8224 ( .A1(n6509), .A2(n8819), .ZN(n8823) );
  NAND2_X1 U8225 ( .A1(n6510), .A2(n9103), .ZN(n8754) );
  NAND2_X1 U8226 ( .A1(n6989), .A2(n9340), .ZN(n6998) );
  NAND2_X1 U8227 ( .A1(n6560), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n6996) );
  NAND2_X1 U8228 ( .A1(n6991), .A2(n6990), .ZN(n6992) );
  AND2_X1 U8229 ( .A1(n7048), .A2(n6992), .ZN(n7231) );
  NAND2_X1 U8230 ( .A1(n6556), .A2(n7231), .ZN(n6995) );
  NAND2_X1 U8231 ( .A1(n6555), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n6994) );
  NAND2_X1 U8232 ( .A1(n6554), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n6993) );
  INV_X1 U8233 ( .A(n7390), .ZN(n9036) );
  AOI22_X1 U8234 ( .A1(n9036), .A2(n9346), .B1(n9345), .B2(n7021), .ZN(n6997)
         );
  NAND2_X1 U8235 ( .A1(n6998), .A2(n6997), .ZN(n7281) );
  AOI211_X1 U8236 ( .C1(n7284), .C2(n10639), .A(n6999), .B(n7281), .ZN(n7081)
         );
  NAND2_X1 U8237 ( .A1(n10362), .A2(n7000), .ZN(n7001) );
  NAND2_X1 U8238 ( .A1(n10641), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n7004) );
  OAI21_X1 U8239 ( .B1(n7081), .B2(n10641), .A(n7004), .ZN(P2_U3527) );
  INV_X1 U8240 ( .A(n8681), .ZN(n7007) );
  NOR2_X1 U8241 ( .A1(n7005), .A2(P1_U3084), .ZN(n8493) );
  AOI21_X1 U8242 ( .B1(P2_DATAO_REG_23__SCAN_IN), .B2(n10324), .A(n8493), .ZN(
        n7006) );
  OAI21_X1 U8243 ( .B1(n7007), .B2(n6276), .A(n7006), .ZN(P1_U3330) );
  AOI211_X1 U8244 ( .C1(n10603), .C2(n7010), .A(n7009), .B(n7008), .ZN(n7019)
         );
  INV_X1 U8245 ( .A(n10311), .ZN(n7013) );
  INV_X1 U8246 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n7011) );
  NOR2_X1 U8247 ( .A1(n10612), .A2(n7011), .ZN(n7012) );
  AOI21_X1 U8248 ( .B1(n7013), .B2(n7016), .A(n7012), .ZN(n7014) );
  OAI21_X1 U8249 ( .B1(n7019), .B2(n10609), .A(n7014), .ZN(P1_U3475) );
  INV_X1 U8250 ( .A(n10246), .ZN(n7017) );
  NOR2_X1 U8251 ( .A1(n10608), .A2(n5552), .ZN(n7015) );
  AOI21_X1 U8252 ( .B1(n7017), .B2(n7016), .A(n7015), .ZN(n7018) );
  OAI21_X1 U8253 ( .B1(n7019), .B2(n10607), .A(n7018), .ZN(P1_U3530) );
  INV_X1 U8254 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n8682) );
  NAND2_X1 U8255 ( .A1(n8681), .A2(n9705), .ZN(n7020) );
  OAI211_X1 U8256 ( .C1(n8682), .C2(n9710), .A(n7020), .B(n8829), .ZN(P2_U3335) );
  NAND2_X1 U8257 ( .A1(n5116), .A2(n7021), .ZN(n7023) );
  XNOR2_X1 U8258 ( .A(n8933), .B(n8050), .ZN(n7022) );
  NAND2_X1 U8259 ( .A1(n7023), .A2(n7022), .ZN(n7037) );
  OR2_X1 U8260 ( .A1(n7023), .A2(n7022), .ZN(n7024) );
  AND2_X1 U8261 ( .A1(n7037), .A2(n7024), .ZN(n7028) );
  OAI21_X1 U8262 ( .B1(n7028), .B2(n7027), .A(n7038), .ZN(n7035) );
  INV_X1 U8263 ( .A(n7029), .ZN(n7031) );
  NAND2_X1 U8264 ( .A1(n8949), .A2(n8047), .ZN(n7030) );
  OAI211_X1 U8265 ( .C1(n8937), .C2(n10582), .A(n7031), .B(n7030), .ZN(n7034)
         );
  OAI22_X1 U8266 ( .A1(n7032), .A2(n9014), .B1(n9011), .B2(n7220), .ZN(n7033)
         );
  AOI211_X1 U8267 ( .C1(n8941), .C2(n7035), .A(n7034), .B(n7033), .ZN(n7036)
         );
  INV_X1 U8268 ( .A(n7036), .ZN(P2_U3241) );
  NAND2_X1 U8269 ( .A1(n7038), .A2(n7037), .ZN(n7059) );
  XNOR2_X1 U8270 ( .A(n7280), .B(n8931), .ZN(n7039) );
  NAND2_X1 U8271 ( .A1(n5116), .A2(n9037), .ZN(n7040) );
  XNOR2_X1 U8272 ( .A(n7039), .B(n7040), .ZN(n7058) );
  INV_X1 U8273 ( .A(n7039), .ZN(n7042) );
  INV_X1 U8274 ( .A(n7040), .ZN(n7041) );
  NAND2_X1 U8275 ( .A1(n7042), .A2(n7041), .ZN(n7043) );
  NAND2_X1 U8276 ( .A1(n7044), .A2(n8727), .ZN(n7047) );
  AOI22_X1 U8277 ( .A1(n7997), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n7996), .B2(
        n7045), .ZN(n7046) );
  XNOR2_X1 U8278 ( .A(n7386), .B(n8933), .ZN(n7099) );
  NOR2_X1 U8279 ( .A1(n7390), .A2(n8932), .ZN(n7100) );
  XNOR2_X1 U8280 ( .A(n7099), .B(n7100), .ZN(n7103) );
  XNOR2_X1 U8281 ( .A(n7104), .B(n7103), .ZN(n7057) );
  INV_X1 U8282 ( .A(n7386), .ZN(n7233) );
  OAI22_X1 U8283 ( .A1(n8937), .A2(n7233), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n6990), .ZN(n7055) );
  NAND2_X1 U8284 ( .A1(n7048), .A2(n9679), .ZN(n7049) );
  AND2_X1 U8285 ( .A1(n7117), .A2(n7049), .ZN(n7400) );
  NAND2_X1 U8286 ( .A1(n6556), .A2(n7400), .ZN(n7053) );
  NAND2_X1 U8287 ( .A1(n6560), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n7052) );
  NAND2_X1 U8288 ( .A1(n6554), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n7051) );
  NAND2_X1 U8289 ( .A1(n6555), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n7050) );
  OAI22_X1 U8290 ( .A1(n7220), .A2(n9014), .B1(n9011), .B2(n7767), .ZN(n7054)
         );
  AOI211_X1 U8291 ( .C1(n7231), .C2(n8949), .A(n7055), .B(n7054), .ZN(n7056)
         );
  OAI21_X1 U8292 ( .B1(n9019), .B2(n7057), .A(n7056), .ZN(P2_U3223) );
  XNOR2_X1 U8293 ( .A(n7059), .B(n7058), .ZN(n7064) );
  OAI22_X1 U8294 ( .A1(n8937), .A2(n7280), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9649), .ZN(n7062) );
  OAI22_X1 U8295 ( .A1(n7060), .A2(n9014), .B1(n9011), .B2(n7390), .ZN(n7061)
         );
  AOI211_X1 U8296 ( .C1(n7277), .C2(n8949), .A(n7062), .B(n7061), .ZN(n7063)
         );
  OAI21_X1 U8297 ( .B1(n7064), .B2(n9019), .A(n7063), .ZN(P2_U3215) );
  AOI21_X1 U8298 ( .B1(n7067), .B2(n7066), .A(n7065), .ZN(n7069) );
  INV_X1 U8299 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n7729) );
  AOI22_X1 U8300 ( .A1(n7738), .A2(n7729), .B1(P2_REG1_REG_14__SCAN_IN), .B2(
        n7730), .ZN(n7068) );
  NOR2_X1 U8301 ( .A1(n7069), .A2(n7068), .ZN(n7728) );
  AOI21_X1 U8302 ( .B1(n7069), .B2(n7068), .A(n7728), .ZN(n7078) );
  NOR2_X1 U8303 ( .A1(n7738), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n7070) );
  AOI21_X1 U8304 ( .B1(P2_REG2_REG_14__SCAN_IN), .B2(n7738), .A(n7070), .ZN(
        n7073) );
  OAI21_X1 U8305 ( .B1(n7622), .B2(P2_REG2_REG_13__SCAN_IN), .A(n7071), .ZN(
        n7072) );
  NAND2_X1 U8306 ( .A1(n7073), .A2(n7072), .ZN(n7737) );
  OAI21_X1 U8307 ( .B1(n7073), .B2(n7072), .A(n7737), .ZN(n7076) );
  NAND2_X1 U8308 ( .A1(P2_U3152), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n7721) );
  NAND2_X1 U8309 ( .A1(n10486), .A2(P2_ADDR_REG_14__SCAN_IN), .ZN(n7074) );
  OAI211_X1 U8310 ( .C1(n10467), .C2(n7730), .A(n7721), .B(n7074), .ZN(n7075)
         );
  AOI21_X1 U8311 ( .B1(n7076), .B2(n10466), .A(n7075), .ZN(n7077) );
  OAI21_X1 U8312 ( .B1(n7078), .B2(n10468), .A(n7077), .ZN(P2_U3259) );
  INV_X1 U8313 ( .A(n7079), .ZN(n7209) );
  INV_X1 U8314 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n7083) );
  OR2_X1 U8315 ( .A1(n7081), .A2(n10643), .ZN(n7082) );
  OAI21_X1 U8316 ( .B1(n10646), .B2(n7083), .A(n7082), .ZN(P2_U3472) );
  INV_X1 U8317 ( .A(n8379), .ZN(n7084) );
  XNOR2_X1 U8318 ( .A(n7085), .B(n4874), .ZN(n7286) );
  XNOR2_X1 U8319 ( .A(n7086), .B(n4874), .ZN(n7089) );
  AOI22_X1 U8320 ( .A1(n10143), .A2(n7087), .B1(n9878), .B2(n10141), .ZN(n7088) );
  OAI21_X1 U8321 ( .B1(n7089), .B2(n9997), .A(n7088), .ZN(n7090) );
  AOI21_X1 U8322 ( .B1(n7286), .B2(n6282), .A(n7090), .ZN(n7290) );
  AND2_X1 U8323 ( .A1(n7091), .A2(n7093), .ZN(n7198) );
  AOI21_X1 U8324 ( .B1(n7287), .B2(n7092), .A(n7198), .ZN(n7288) );
  NOR2_X1 U8325 ( .A1(n7093), .A2(n10115), .ZN(n7096) );
  INV_X1 U8326 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n7094) );
  OAI22_X1 U8327 ( .A1(n10148), .A2(n7094), .B1(n7184), .B2(n10145), .ZN(n7095) );
  AOI211_X1 U8328 ( .C1(n7288), .C2(n10097), .A(n7096), .B(n7095), .ZN(n7098)
         );
  NAND2_X1 U8329 ( .A1(n7286), .A2(n7616), .ZN(n7097) );
  OAI211_X1 U8330 ( .C1(n7290), .C2(n10088), .A(n7098), .B(n7097), .ZN(
        P1_U3282) );
  INV_X1 U8331 ( .A(n7099), .ZN(n7101) );
  AND2_X1 U8332 ( .A1(n7101), .A2(n7100), .ZN(n7102) );
  AOI21_X1 U8333 ( .B1(n7104), .B2(n7103), .A(n7102), .ZN(n7115) );
  NAND2_X1 U8334 ( .A1(n7105), .A2(n8727), .ZN(n7108) );
  AOI22_X1 U8335 ( .A1(n7997), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n7996), .B2(
        n7106), .ZN(n7107) );
  XNOR2_X1 U8336 ( .A(n7587), .B(n8933), .ZN(n7109) );
  OR2_X1 U8337 ( .A1(n7767), .A2(n8932), .ZN(n7110) );
  NAND2_X1 U8338 ( .A1(n7109), .A2(n7110), .ZN(n7156) );
  INV_X1 U8339 ( .A(n7109), .ZN(n7112) );
  INV_X1 U8340 ( .A(n7110), .ZN(n7111) );
  NAND2_X1 U8341 ( .A1(n7112), .A2(n7111), .ZN(n7113) );
  AND2_X1 U8342 ( .A1(n7156), .A2(n7113), .ZN(n7114) );
  OAI21_X1 U8343 ( .B1(n7115), .B2(n7114), .A(n7157), .ZN(n7128) );
  NAND2_X1 U8344 ( .A1(n7117), .A2(n7116), .ZN(n7118) );
  AND2_X1 U8345 ( .A1(n7162), .A2(n7118), .ZN(n7776) );
  NAND2_X1 U8346 ( .A1(n6556), .A2(n7776), .ZN(n7122) );
  NAND2_X1 U8347 ( .A1(n6560), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n7121) );
  NAND2_X1 U8348 ( .A1(n6554), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n7120) );
  NAND2_X1 U8349 ( .A1(n6555), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n7119) );
  OAI22_X1 U8350 ( .A1(n7390), .A2(n9014), .B1(n9011), .B2(n7562), .ZN(n7127)
         );
  INV_X1 U8351 ( .A(n7123), .ZN(n7125) );
  NAND2_X1 U8352 ( .A1(n8949), .A2(n7400), .ZN(n7124) );
  OAI211_X1 U8353 ( .C1(n8937), .C2(n4983), .A(n7125), .B(n7124), .ZN(n7126)
         );
  AOI211_X1 U8354 ( .C1(n7128), .C2(n8941), .A(n7127), .B(n7126), .ZN(n7129)
         );
  INV_X1 U8355 ( .A(n7129), .ZN(P2_U3233) );
  INV_X1 U8356 ( .A(n7130), .ZN(n7132) );
  NAND2_X1 U8357 ( .A1(n7132), .A2(n7131), .ZN(n7133) );
  INV_X1 U8358 ( .A(n7326), .ZN(n7137) );
  NAND2_X1 U8359 ( .A1(n7138), .A2(n6216), .ZN(n7136) );
  OR2_X1 U8360 ( .A1(n7181), .A2(n6305), .ZN(n7135) );
  NAND2_X1 U8361 ( .A1(n7136), .A2(n7135), .ZN(n7329) );
  NAND2_X1 U8362 ( .A1(n7137), .A2(n7329), .ZN(n7143) );
  NAND2_X1 U8363 ( .A1(n7138), .A2(n8207), .ZN(n7140) );
  OR2_X1 U8364 ( .A1(n7181), .A2(n8208), .ZN(n7139) );
  NAND2_X1 U8365 ( .A1(n7140), .A2(n7139), .ZN(n7141) );
  XNOR2_X1 U8366 ( .A(n7141), .B(n8195), .ZN(n7327) );
  INV_X1 U8367 ( .A(n7327), .ZN(n7332) );
  NAND2_X1 U8368 ( .A1(n7143), .A2(n7332), .ZN(n7173) );
  INV_X1 U8369 ( .A(n7173), .ZN(n7145) );
  INV_X1 U8370 ( .A(n7329), .ZN(n7142) );
  NAND2_X1 U8371 ( .A1(n7326), .A2(n7142), .ZN(n7172) );
  AOI21_X1 U8372 ( .B1(n7143), .B2(n7172), .A(n7332), .ZN(n7144) );
  AOI21_X1 U8373 ( .B1(n7145), .B2(n7172), .A(n7144), .ZN(n7155) );
  INV_X1 U8374 ( .A(n7146), .ZN(n7153) );
  OR2_X1 U8375 ( .A1(n9846), .A2(n8068), .ZN(n7149) );
  NOR2_X1 U8376 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7147), .ZN(n9917) );
  INV_X1 U8377 ( .A(n9917), .ZN(n7148) );
  OAI211_X1 U8378 ( .C1(n9860), .C2(n7150), .A(n7149), .B(n7148), .ZN(n7152)
         );
  NOR2_X1 U8379 ( .A1(n5026), .A2(n9866), .ZN(n7151) );
  AOI211_X1 U8380 ( .C1(n7153), .C2(n9783), .A(n7152), .B(n7151), .ZN(n7154)
         );
  OAI21_X1 U8381 ( .B1(n7155), .B2(n9853), .A(n7154), .ZN(P1_U3219) );
  NAND2_X1 U8382 ( .A1(n7158), .A2(n8727), .ZN(n7161) );
  AOI22_X1 U8383 ( .A1(n7997), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n7996), .B2(
        n7159), .ZN(n7160) );
  NAND2_X1 U8384 ( .A1(n7161), .A2(n7160), .ZN(n7563) );
  XNOR2_X1 U8385 ( .A(n7563), .B(n8931), .ZN(n7297) );
  NOR2_X1 U8386 ( .A1(n7562), .A2(n8932), .ZN(n7296) );
  XNOR2_X1 U8387 ( .A(n7297), .B(n7296), .ZN(n7407) );
  XNOR2_X1 U8388 ( .A(n7405), .B(n7407), .ZN(n7171) );
  OAI22_X1 U8389 ( .A1(n8937), .A2(n10614), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7116), .ZN(n7169) );
  INV_X1 U8390 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n9561) );
  NAND2_X1 U8391 ( .A1(n7162), .A2(n9561), .ZN(n7163) );
  AND2_X1 U8392 ( .A1(n7305), .A2(n7163), .ZN(n7645) );
  NAND2_X1 U8393 ( .A1(n6556), .A2(n7645), .ZN(n7167) );
  NAND2_X1 U8394 ( .A1(n6560), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n7166) );
  NAND2_X1 U8395 ( .A1(n6554), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n7165) );
  NAND2_X1 U8396 ( .A1(n6555), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n7164) );
  OAI22_X1 U8397 ( .A1(n7767), .A2(n9014), .B1(n9011), .B2(n7768), .ZN(n7168)
         );
  AOI211_X1 U8398 ( .C1(n7776), .C2(n8949), .A(n7169), .B(n7168), .ZN(n7170)
         );
  OAI21_X1 U8399 ( .B1(n7171), .B2(n9019), .A(n7170), .ZN(P2_U3219) );
  NAND2_X1 U8400 ( .A1(n7173), .A2(n7172), .ZN(n7180) );
  NAND2_X1 U8401 ( .A1(n7287), .A2(n8207), .ZN(n7175) );
  NAND2_X1 U8402 ( .A1(n9879), .A2(n6216), .ZN(n7174) );
  NAND2_X1 U8403 ( .A1(n7175), .A2(n7174), .ZN(n7176) );
  XNOR2_X1 U8404 ( .A(n7176), .B(n8195), .ZN(n7328) );
  NAND2_X1 U8405 ( .A1(n7287), .A2(n6216), .ZN(n7178) );
  NAND2_X1 U8406 ( .A1(n9879), .A2(n8212), .ZN(n7177) );
  NAND2_X1 U8407 ( .A1(n7178), .A2(n7177), .ZN(n7330) );
  XNOR2_X1 U8408 ( .A(n7328), .B(n7330), .ZN(n7179) );
  XNOR2_X1 U8409 ( .A(n7180), .B(n7179), .ZN(n7187) );
  AND2_X1 U8410 ( .A1(P1_U3084), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n10442) );
  NOR2_X1 U8411 ( .A1(n9860), .A2(n7181), .ZN(n7182) );
  AOI211_X1 U8412 ( .C1(n9863), .C2(n9878), .A(n10442), .B(n7182), .ZN(n7183)
         );
  OAI21_X1 U8413 ( .B1(n9858), .B2(n7184), .A(n7183), .ZN(n7185) );
  AOI21_X1 U8414 ( .B1(n7287), .B2(n9837), .A(n7185), .ZN(n7186) );
  OAI21_X1 U8415 ( .B1(n7187), .B2(n9853), .A(n7186), .ZN(P1_U3229) );
  INV_X1 U8416 ( .A(n8562), .ZN(n7204) );
  INV_X1 U8417 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n7188) );
  OAI222_X1 U8418 ( .A1(n6276), .A2(n7204), .B1(P1_U3084), .B2(n7189), .C1(
        n7188), .C2(n8101), .ZN(P1_U3329) );
  XNOR2_X1 U8419 ( .A(n7190), .B(n8347), .ZN(n10604) );
  OAI21_X1 U8420 ( .B1(n8253), .B2(n7192), .A(n7191), .ZN(n7193) );
  NAND2_X1 U8421 ( .A1(n7193), .A2(n10140), .ZN(n7195) );
  AOI22_X1 U8422 ( .A1(n10143), .A2(n9879), .B1(n9877), .B2(n10141), .ZN(n7194) );
  NAND2_X1 U8423 ( .A1(n7195), .A2(n7194), .ZN(n7196) );
  AOI21_X1 U8424 ( .B1(n10604), .B2(n6282), .A(n7196), .ZN(n10606) );
  OAI211_X1 U8425 ( .C1(n7198), .C2(n10601), .A(n5984), .B(n7197), .ZN(n10599)
         );
  INV_X1 U8426 ( .A(n10110), .ZN(n7702) );
  OAI22_X1 U8427 ( .A1(n10148), .A2(n7199), .B1(n8072), .B2(n10145), .ZN(n7200) );
  AOI21_X1 U8428 ( .B1(n8074), .B2(n10156), .A(n7200), .ZN(n7201) );
  OAI21_X1 U8429 ( .B1(n10599), .B2(n7702), .A(n7201), .ZN(n7202) );
  AOI21_X1 U8430 ( .B1(n10604), .B2(n7616), .A(n7202), .ZN(n7203) );
  OAI21_X1 U8431 ( .B1(n10606), .B2(n10088), .A(n7203), .ZN(P1_U3281) );
  OAI222_X1 U8432 ( .A1(P2_U3152), .A2(n7206), .B1(n9710), .B2(n7205), .C1(
        n7204), .C2(n8039), .ZN(P2_U3334) );
  NOR2_X1 U8433 ( .A1(n9339), .A2(n7207), .ZN(n10503) );
  INV_X1 U8434 ( .A(n7208), .ZN(n7211) );
  NAND3_X1 U8435 ( .A1(n7211), .A2(n7210), .A3(n7209), .ZN(n7217) );
  OR2_X1 U8436 ( .A1(n7212), .A2(n9300), .ZN(n7252) );
  NAND2_X1 U8437 ( .A1(n9302), .A2(n7252), .ZN(n7213) );
  OAI22_X1 U8438 ( .A1(n10503), .A2(n9253), .B1(n9321), .B2(n9318), .ZN(n10505) );
  AOI21_X1 U8439 ( .B1(P2_REG3_REG_0__SCAN_IN), .B2(n9350), .A(n10505), .ZN(
        n7214) );
  NOR2_X1 U8440 ( .A1(n9223), .A2(n7214), .ZN(n7215) );
  AOI21_X1 U8441 ( .B1(n9354), .B2(P2_REG2_REG_0__SCAN_IN), .A(n7215), .ZN(
        n7219) );
  OR2_X1 U8442 ( .A1(n7217), .A2(n5116), .ZN(n9139) );
  OAI21_X1 U8443 ( .B1(n9336), .B2(n9353), .A(n9351), .ZN(n7218) );
  OAI211_X1 U8444 ( .C1(n10503), .C2(n9285), .A(n7219), .B(n7218), .ZN(
        P2_U3296) );
  NAND2_X1 U8445 ( .A1(n7280), .A2(n7220), .ZN(n7221) );
  OAI21_X1 U8446 ( .B1(n7222), .B2(n8768), .A(n7221), .ZN(n7223) );
  OR2_X1 U8447 ( .A1(n7386), .A2(n7390), .ZN(n8620) );
  NAND2_X1 U8448 ( .A1(n7386), .A2(n7390), .ZN(n8616) );
  NAND2_X1 U8449 ( .A1(n8620), .A2(n8616), .ZN(n7225) );
  OAI21_X1 U8450 ( .B1(n7224), .B2(n7225), .A(n7388), .ZN(n7270) );
  INV_X1 U8451 ( .A(n7225), .ZN(n8769) );
  NAND2_X1 U8452 ( .A1(n7226), .A2(n8618), .ZN(n7227) );
  OAI21_X1 U8453 ( .B1(n8769), .B2(n7227), .A(n7394), .ZN(n7228) );
  INV_X1 U8454 ( .A(n7767), .ZN(n9035) );
  AOI222_X1 U8455 ( .A1(n9340), .A2(n7228), .B1(n9035), .B2(n9346), .C1(n9037), 
        .C2(n9345), .ZN(n7269) );
  MUX2_X1 U8456 ( .A(n6700), .B(n7269), .S(n9307), .Z(n7236) );
  INV_X1 U8457 ( .A(n7399), .ZN(n7229) );
  AOI211_X1 U8458 ( .C1(n7386), .C2(n7230), .A(n10637), .B(n7229), .ZN(n7267)
         );
  NOR2_X1 U8459 ( .A1(n9223), .A2(n9103), .ZN(n9187) );
  INV_X1 U8460 ( .A(n7231), .ZN(n7232) );
  OAI22_X1 U8461 ( .A1(n9272), .A2(n7233), .B1(n9304), .B2(n7232), .ZN(n7234)
         );
  AOI21_X1 U8462 ( .B1(n7267), .B2(n9187), .A(n7234), .ZN(n7235) );
  OAI211_X1 U8463 ( .C1(n9285), .C2(n7270), .A(n7236), .B(n7235), .ZN(P2_U3288) );
  XNOR2_X1 U8464 ( .A(n9039), .B(n6519), .ZN(n8767) );
  INV_X1 U8465 ( .A(n8767), .ZN(n8591) );
  XNOR2_X1 U8466 ( .A(n7237), .B(n8591), .ZN(n10557) );
  NAND2_X1 U8467 ( .A1(n7254), .A2(n7247), .ZN(n7238) );
  NAND2_X1 U8468 ( .A1(n7377), .A2(n7238), .ZN(n10558) );
  NOR2_X1 U8469 ( .A1(n9139), .A2(n10558), .ZN(n7241) );
  INV_X1 U8470 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n7239) );
  NOR2_X1 U8471 ( .A1(n9307), .A2(n7239), .ZN(n7240) );
  AOI211_X1 U8472 ( .C1(n9350), .C2(n7242), .A(n7241), .B(n7240), .ZN(n7249)
         );
  XNOR2_X1 U8473 ( .A(n7243), .B(n8591), .ZN(n7244) );
  NAND2_X1 U8474 ( .A1(n7244), .A2(n9340), .ZN(n7246) );
  AOI22_X1 U8475 ( .A1(n9040), .A2(n9345), .B1(n9346), .B2(n9038), .ZN(n7245)
         );
  NAND2_X1 U8476 ( .A1(n7246), .A2(n7245), .ZN(n10560) );
  AOI22_X1 U8477 ( .A1(n9336), .A2(n7247), .B1(n9307), .B2(n10560), .ZN(n7248)
         );
  OAI211_X1 U8478 ( .C1(n9285), .C2(n10557), .A(n7249), .B(n7248), .ZN(
        P2_U3292) );
  XNOR2_X1 U8479 ( .A(n7251), .B(n7250), .ZN(n10538) );
  INV_X1 U8480 ( .A(n10538), .ZN(n7266) );
  OR2_X1 U8481 ( .A1(n9354), .A2(n7252), .ZN(n9311) );
  OR2_X1 U8482 ( .A1(n10527), .A2(n10539), .ZN(n7253) );
  NAND2_X1 U8483 ( .A1(n7254), .A2(n7253), .ZN(n10540) );
  OAI22_X1 U8484 ( .A1(n9139), .A2(n10540), .B1(P2_REG3_REG_3__SCAN_IN), .B2(
        n9304), .ZN(n7255) );
  AOI21_X1 U8485 ( .B1(n9354), .B2(P2_REG2_REG_3__SCAN_IN), .A(n7255), .ZN(
        n7265) );
  INV_X1 U8486 ( .A(n9302), .ZN(n9314) );
  NAND2_X1 U8487 ( .A1(n10538), .A2(n9314), .ZN(n7263) );
  OAI21_X1 U8488 ( .B1(n8761), .B2(n7257), .A(n7256), .ZN(n7261) );
  NAND2_X1 U8489 ( .A1(n9039), .A2(n9346), .ZN(n7258) );
  OAI21_X1 U8490 ( .B1(n7259), .B2(n9320), .A(n7258), .ZN(n7260) );
  AOI21_X1 U8491 ( .B1(n7261), .B2(n9340), .A(n7260), .ZN(n7262) );
  NAND2_X1 U8492 ( .A1(n7263), .A2(n7262), .ZN(n10545) );
  AOI22_X1 U8493 ( .A1(n9336), .A2(n8904), .B1(n9307), .B2(n10545), .ZN(n7264)
         );
  OAI211_X1 U8494 ( .C1(n7266), .C2(n9311), .A(n7265), .B(n7264), .ZN(P2_U3293) );
  AOI21_X1 U8495 ( .B1(n10632), .B2(n7386), .A(n7267), .ZN(n7268) );
  OAI211_X1 U8496 ( .C1(n10556), .C2(n7270), .A(n7269), .B(n7268), .ZN(n7273)
         );
  NAND2_X1 U8497 ( .A1(n7273), .A2(n10642), .ZN(n7271) );
  OAI21_X1 U8498 ( .B1(n10642), .B2(n7272), .A(n7271), .ZN(P2_U3528) );
  INV_X1 U8499 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n7275) );
  NAND2_X1 U8500 ( .A1(n7273), .A2(n10646), .ZN(n7274) );
  OAI21_X1 U8501 ( .B1(n10646), .B2(n7275), .A(n7274), .ZN(P2_U3475) );
  INV_X1 U8502 ( .A(n7276), .ZN(n7278) );
  AOI22_X1 U8503 ( .A1(n9353), .A2(n7278), .B1(n7277), .B2(n9350), .ZN(n7279)
         );
  OAI21_X1 U8504 ( .B1(n7280), .B2(n9272), .A(n7279), .ZN(n7283) );
  MUX2_X1 U8505 ( .A(P2_REG2_REG_7__SCAN_IN), .B(n7281), .S(n9307), .Z(n7282)
         );
  AOI211_X1 U8506 ( .C1(n7284), .C2(n9337), .A(n7283), .B(n7282), .ZN(n7285)
         );
  INV_X1 U8507 ( .A(n7285), .ZN(P2_U3289) );
  INV_X1 U8508 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n7293) );
  INV_X1 U8509 ( .A(n7286), .ZN(n7291) );
  AOI22_X1 U8510 ( .A1(n7288), .A2(n5984), .B1(n10269), .B2(n7287), .ZN(n7289)
         );
  OAI211_X1 U8511 ( .C1(n10273), .C2(n7291), .A(n7290), .B(n7289), .ZN(n7294)
         );
  NAND2_X1 U8512 ( .A1(n7294), .A2(n10612), .ZN(n7292) );
  OAI21_X1 U8513 ( .B1(n10612), .B2(n7293), .A(n7292), .ZN(P1_U3481) );
  NAND2_X1 U8514 ( .A1(n7294), .A2(n10608), .ZN(n7295) );
  OAI21_X1 U8515 ( .B1(n10608), .B2(n5584), .A(n7295), .ZN(P1_U3532) );
  OR2_X1 U8516 ( .A1(n7405), .A2(n7407), .ZN(n7298) );
  NAND2_X1 U8517 ( .A1(n7297), .A2(n7296), .ZN(n7408) );
  NAND2_X1 U8518 ( .A1(n7298), .A2(n7408), .ZN(n7302) );
  OR2_X1 U8519 ( .A1(n7299), .A2(n6564), .ZN(n7301) );
  AOI22_X1 U8520 ( .A1(n7997), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n7996), .B2(
        n9048), .ZN(n7300) );
  NAND2_X1 U8521 ( .A1(n7301), .A2(n7300), .ZN(n7651) );
  XNOR2_X1 U8522 ( .A(n7651), .B(n8933), .ZN(n7410) );
  NOR2_X1 U8523 ( .A1(n7768), .A2(n8932), .ZN(n7411) );
  XNOR2_X1 U8524 ( .A(n7410), .B(n7411), .ZN(n7406) );
  XNOR2_X1 U8525 ( .A(n7302), .B(n7406), .ZN(n7314) );
  INV_X1 U8526 ( .A(n7651), .ZN(n10626) );
  OAI22_X1 U8527 ( .A1(n8937), .A2(n10626), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9561), .ZN(n7312) );
  NAND2_X1 U8528 ( .A1(n7305), .A2(n7304), .ZN(n7306) );
  AND2_X1 U8529 ( .A1(n7424), .A2(n7306), .ZN(n7573) );
  NAND2_X1 U8530 ( .A1(n6556), .A2(n7573), .ZN(n7310) );
  NAND2_X1 U8531 ( .A1(n6560), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n7309) );
  NAND2_X1 U8532 ( .A1(n6554), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n7308) );
  NAND2_X1 U8533 ( .A1(n6555), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n7307) );
  OAI22_X1 U8534 ( .A1(n7562), .A2(n9014), .B1(n9011), .B2(n7657), .ZN(n7311)
         );
  AOI211_X1 U8535 ( .C1(n7645), .C2(n8949), .A(n7312), .B(n7311), .ZN(n7313)
         );
  OAI21_X1 U8536 ( .B1(n7314), .B2(n9019), .A(n7313), .ZN(P2_U3238) );
  INV_X1 U8537 ( .A(n8383), .ZN(n7316) );
  AND2_X1 U8538 ( .A1(n7316), .A2(n8403), .ZN(n8256) );
  INV_X1 U8539 ( .A(n8256), .ZN(n8346) );
  XNOR2_X1 U8540 ( .A(n7315), .B(n8346), .ZN(n10267) );
  XNOR2_X1 U8541 ( .A(n7317), .B(n8346), .ZN(n7319) );
  AOI22_X1 U8542 ( .A1(n10143), .A2(n9878), .B1(n9876), .B2(n10141), .ZN(n7318) );
  OAI21_X1 U8543 ( .B1(n7319), .B2(n9997), .A(n7318), .ZN(n7320) );
  AOI21_X1 U8544 ( .B1(n10267), .B2(n6282), .A(n7320), .ZN(n10272) );
  AOI21_X1 U8545 ( .B1(n10268), .B2(n7197), .A(n5015), .ZN(n10270) );
  INV_X1 U8546 ( .A(n10268), .ZN(n7357) );
  NOR2_X1 U8547 ( .A1(n7357), .A2(n10115), .ZN(n7322) );
  OAI22_X1 U8548 ( .A1(n10148), .A2(n8081), .B1(n7350), .B2(n10145), .ZN(n7321) );
  AOI211_X1 U8549 ( .C1(n10270), .C2(n10097), .A(n7322), .B(n7321), .ZN(n7324)
         );
  NAND2_X1 U8550 ( .A1(n10267), .A2(n7616), .ZN(n7323) );
  OAI211_X1 U8551 ( .C1(n10272), .C2(n10088), .A(n7324), .B(n7323), .ZN(
        P1_U3280) );
  AOI22_X1 U8552 ( .A1(n7328), .A2(n7330), .B1(n7329), .B2(n7327), .ZN(n7325)
         );
  OAI21_X1 U8553 ( .B1(n7327), .B2(n7329), .A(n7330), .ZN(n7334) );
  INV_X1 U8554 ( .A(n7328), .ZN(n7333) );
  NOR2_X1 U8555 ( .A1(n7330), .A2(n7329), .ZN(n7331) );
  INV_X1 U8556 ( .A(n7343), .ZN(n7340) );
  NAND2_X1 U8557 ( .A1(n8074), .A2(n8207), .ZN(n7337) );
  OR2_X1 U8558 ( .A1(n7352), .A2(n8208), .ZN(n7336) );
  NAND2_X1 U8559 ( .A1(n7337), .A2(n7336), .ZN(n7338) );
  XNOR2_X1 U8560 ( .A(n7338), .B(n8145), .ZN(n7342) );
  INV_X1 U8561 ( .A(n7342), .ZN(n7339) );
  NAND2_X1 U8562 ( .A1(n7340), .A2(n7339), .ZN(n8065) );
  NOR2_X1 U8563 ( .A1(n7352), .A2(n6305), .ZN(n7341) );
  AOI21_X1 U8564 ( .B1(n8074), .B2(n6216), .A(n7341), .ZN(n8066) );
  NAND2_X1 U8565 ( .A1(n8065), .A2(n8066), .ZN(n7442) );
  NAND2_X1 U8566 ( .A1(n7343), .A2(n7342), .ZN(n8064) );
  AND2_X1 U8567 ( .A1(n7442), .A2(n8064), .ZN(n7349) );
  NAND2_X1 U8568 ( .A1(n10268), .A2(n8207), .ZN(n7345) );
  NAND2_X1 U8569 ( .A1(n9877), .A2(n6216), .ZN(n7344) );
  NAND2_X1 U8570 ( .A1(n7345), .A2(n7344), .ZN(n7346) );
  XNOR2_X1 U8571 ( .A(n7346), .B(n8195), .ZN(n7446) );
  AND2_X1 U8572 ( .A1(n9877), .A2(n8212), .ZN(n7347) );
  AOI21_X1 U8573 ( .B1(n10268), .B2(n6216), .A(n7347), .ZN(n7444) );
  XNOR2_X1 U8574 ( .A(n7446), .B(n7444), .ZN(n7440) );
  AND2_X1 U8575 ( .A1(n8064), .A2(n7440), .ZN(n7348) );
  NAND2_X1 U8576 ( .A1(n7348), .A2(n7442), .ZN(n9767) );
  OAI211_X1 U8577 ( .C1(n7349), .C2(n7440), .A(n9855), .B(n9767), .ZN(n7356)
         );
  INV_X1 U8578 ( .A(n7350), .ZN(n7354) );
  AND2_X1 U8579 ( .A1(P1_U3084), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n8089) );
  AOI21_X1 U8580 ( .B1(n9863), .B2(n9876), .A(n8089), .ZN(n7351) );
  OAI21_X1 U8581 ( .B1(n7352), .B2(n9860), .A(n7351), .ZN(n7353) );
  AOI21_X1 U8582 ( .B1(n7354), .B2(n9783), .A(n7353), .ZN(n7355) );
  OAI211_X1 U8583 ( .C1(n7357), .C2(n9866), .A(n7356), .B(n7355), .ZN(P1_U3234) );
  INV_X1 U8584 ( .A(n8698), .ZN(n7359) );
  OAI222_X1 U8585 ( .A1(P1_U3084), .A2(n5886), .B1(n6276), .B2(n7359), .C1(
        n8101), .C2(n7358), .ZN(P1_U3328) );
  INV_X1 U8586 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n8699) );
  OAI222_X1 U8587 ( .A1(P2_U3152), .A2(n7360), .B1(n8039), .B2(n7359), .C1(
        n8699), .C2(n8230), .ZN(P2_U3333) );
  INV_X1 U8588 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n7527) );
  NAND2_X1 U8589 ( .A1(P1_U3084), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n7682) );
  OAI211_X1 U8590 ( .C1(P1_REG1_REG_15__SCAN_IN), .C2(n7362), .A(n10443), .B(
        n7361), .ZN(n7363) );
  OAI211_X1 U8591 ( .C1(n10425), .C2(n7527), .A(n7682), .B(n7363), .ZN(n7368)
         );
  AOI211_X1 U8592 ( .C1(n7366), .C2(n7365), .A(n7364), .B(n10451), .ZN(n7367)
         );
  AOI211_X1 U8593 ( .C1(n10459), .C2(n7369), .A(n7368), .B(n7367), .ZN(n7370)
         );
  INV_X1 U8594 ( .A(n7370), .ZN(P1_U3256) );
  INV_X1 U8595 ( .A(n8764), .ZN(n7371) );
  XNOR2_X1 U8596 ( .A(n7372), .B(n7371), .ZN(n7375) );
  INV_X1 U8597 ( .A(n7373), .ZN(n7374) );
  AOI21_X1 U8598 ( .B1(n7375), .B2(n9340), .A(n7374), .ZN(n10570) );
  XNOR2_X1 U8599 ( .A(n7376), .B(n8764), .ZN(n10567) );
  INV_X1 U8600 ( .A(n9187), .ZN(n7648) );
  NAND2_X1 U8601 ( .A1(n7377), .A2(n7381), .ZN(n7378) );
  NAND2_X1 U8602 ( .A1(n7378), .A2(n10511), .ZN(n7379) );
  OR2_X1 U8603 ( .A1(n7379), .A2(n8044), .ZN(n10564) );
  AOI22_X1 U8604 ( .A1(n9354), .A2(P2_REG2_REG_5__SCAN_IN), .B1(n7380), .B2(
        n9350), .ZN(n7383) );
  NAND2_X1 U8605 ( .A1(n9336), .A2(n7381), .ZN(n7382) );
  OAI211_X1 U8606 ( .C1(n7648), .C2(n10564), .A(n7383), .B(n7382), .ZN(n7384)
         );
  AOI21_X1 U8607 ( .B1(n9337), .B2(n10567), .A(n7384), .ZN(n7385) );
  OAI21_X1 U8608 ( .B1(n9223), .B2(n10570), .A(n7385), .ZN(P2_U3291) );
  NAND2_X1 U8609 ( .A1(n7386), .A2(n9036), .ZN(n7387) );
  INV_X1 U8610 ( .A(n7569), .ZN(n7389) );
  NAND2_X1 U8611 ( .A1(n7587), .A2(n7767), .ZN(n8617) );
  INV_X1 U8612 ( .A(n8770), .ZN(n7392) );
  OAI21_X1 U8613 ( .B1(n7389), .B2(n7392), .A(n7642), .ZN(n7586) );
  OAI22_X1 U8614 ( .A1(n7562), .A2(n9318), .B1(n7390), .B2(n9320), .ZN(n7398)
         );
  INV_X1 U8615 ( .A(n8616), .ZN(n7391) );
  NOR2_X1 U8616 ( .A1(n7392), .A2(n7391), .ZN(n7393) );
  INV_X1 U8617 ( .A(n7763), .ZN(n7396) );
  AOI21_X1 U8618 ( .B1(n7394), .B2(n8616), .A(n8770), .ZN(n7395) );
  NOR3_X1 U8619 ( .A1(n7396), .A2(n7395), .A3(n9253), .ZN(n7397) );
  AOI211_X1 U8620 ( .C1(n9314), .C2(n7586), .A(n7398), .B(n7397), .ZN(n7590)
         );
  INV_X1 U8621 ( .A(n9311), .ZN(n9313) );
  AOI21_X1 U8622 ( .B1(n7587), .B2(n7399), .A(n7773), .ZN(n7588) );
  NAND2_X1 U8623 ( .A1(n7588), .A2(n9353), .ZN(n7402) );
  AOI22_X1 U8624 ( .A1(n9354), .A2(P2_REG2_REG_9__SCAN_IN), .B1(n7400), .B2(
        n9350), .ZN(n7401) );
  OAI211_X1 U8625 ( .C1(n4983), .C2(n9272), .A(n7402), .B(n7401), .ZN(n7403)
         );
  AOI21_X1 U8626 ( .B1(n7586), .B2(n9313), .A(n7403), .ZN(n7404) );
  OAI21_X1 U8627 ( .B1(n7590), .B2(n9354), .A(n7404), .ZN(P2_U3287) );
  INV_X1 U8628 ( .A(n7406), .ZN(n7409) );
  INV_X1 U8629 ( .A(n7410), .ZN(n7412) );
  NAND2_X1 U8630 ( .A1(n7414), .A2(n7413), .ZN(n7619) );
  OR2_X1 U8631 ( .A1(n7415), .A2(n6564), .ZN(n7418) );
  AOI22_X1 U8632 ( .A1(n7997), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n7996), .B2(
        n7416), .ZN(n7417) );
  XNOR2_X1 U8633 ( .A(n10633), .B(n8931), .ZN(n7422) );
  INV_X1 U8634 ( .A(n7422), .ZN(n7420) );
  NOR2_X1 U8635 ( .A1(n7657), .A2(n8932), .ZN(n7421) );
  INV_X1 U8636 ( .A(n7421), .ZN(n7419) );
  NAND2_X1 U8637 ( .A1(n7420), .A2(n7419), .ZN(n7620) );
  AND2_X1 U8638 ( .A1(n7422), .A2(n7421), .ZN(n7618) );
  NOR2_X1 U8639 ( .A1(n5131), .A2(n7618), .ZN(n7423) );
  XNOR2_X1 U8640 ( .A(n7619), .B(n7423), .ZN(n7435) );
  INV_X1 U8641 ( .A(n7768), .ZN(n9033) );
  AOI22_X1 U8642 ( .A1(n8947), .A2(n9033), .B1(n7573), .B2(n8949), .ZN(n7434)
         );
  NAND2_X1 U8643 ( .A1(n7424), .A2(n9556), .ZN(n7425) );
  AND2_X1 U8644 ( .A1(n7626), .A2(n7425), .ZN(n7666) );
  NAND2_X1 U8645 ( .A1(n6556), .A2(n7666), .ZN(n7429) );
  NAND2_X1 U8646 ( .A1(n6560), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n7428) );
  NAND2_X1 U8647 ( .A1(n6554), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n7427) );
  NAND2_X1 U8648 ( .A1(n6555), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n7426) );
  INV_X1 U8649 ( .A(n7430), .ZN(n7431) );
  OAI21_X1 U8650 ( .B1(n9011), .B2(n7825), .A(n7431), .ZN(n7432) );
  AOI21_X1 U8651 ( .B1(n10633), .B2(n9017), .A(n7432), .ZN(n7433) );
  OAI211_X1 U8652 ( .C1(n7435), .C2(n9019), .A(n7434), .B(n7433), .ZN(P2_U3226) );
  NAND2_X1 U8653 ( .A1(n10263), .A2(n8207), .ZN(n7437) );
  OR2_X1 U8654 ( .A1(n7603), .A2(n8208), .ZN(n7436) );
  NAND2_X1 U8655 ( .A1(n7437), .A2(n7436), .ZN(n7438) );
  XNOR2_X1 U8656 ( .A(n7438), .B(n8145), .ZN(n7447) );
  NOR2_X1 U8657 ( .A1(n7603), .A2(n6305), .ZN(n7439) );
  AOI21_X1 U8658 ( .B1(n10263), .B2(n6216), .A(n7439), .ZN(n7448) );
  NAND2_X1 U8659 ( .A1(n7447), .A2(n7448), .ZN(n9764) );
  AND2_X1 U8660 ( .A1(n9764), .A2(n7440), .ZN(n7441) );
  AND2_X1 U8661 ( .A1(n7441), .A2(n8064), .ZN(n7443) );
  NAND2_X1 U8662 ( .A1(n7443), .A2(n7442), .ZN(n7454) );
  INV_X1 U8663 ( .A(n9764), .ZN(n7452) );
  INV_X1 U8664 ( .A(n7444), .ZN(n7445) );
  NAND2_X1 U8665 ( .A1(n7446), .A2(n7445), .ZN(n9766) );
  INV_X1 U8666 ( .A(n7447), .ZN(n7450) );
  INV_X1 U8667 ( .A(n7448), .ZN(n7449) );
  NAND2_X1 U8668 ( .A1(n7450), .A2(n7449), .ZN(n9765) );
  AND2_X1 U8669 ( .A1(n9766), .A2(n9765), .ZN(n7451) );
  OR2_X1 U8670 ( .A1(n7452), .A2(n7451), .ZN(n7453) );
  NAND2_X1 U8671 ( .A1(n7454), .A2(n7453), .ZN(n7543) );
  NAND2_X1 U8672 ( .A1(n10254), .A2(n6216), .ZN(n7456) );
  OR2_X1 U8673 ( .A1(n7693), .A2(n6305), .ZN(n7455) );
  NAND2_X1 U8674 ( .A1(n7456), .A2(n7455), .ZN(n7541) );
  NAND2_X1 U8675 ( .A1(n10254), .A2(n8207), .ZN(n7458) );
  OR2_X1 U8676 ( .A1(n7693), .A2(n8208), .ZN(n7457) );
  NAND2_X1 U8677 ( .A1(n7458), .A2(n7457), .ZN(n7459) );
  XNOR2_X1 U8678 ( .A(n7459), .B(n8195), .ZN(n7542) );
  XOR2_X1 U8679 ( .A(n7541), .B(n7542), .Z(n7460) );
  XNOR2_X1 U8680 ( .A(n7543), .B(n7460), .ZN(n7466) );
  OAI21_X1 U8681 ( .B1(n9860), .B2(n7603), .A(n7461), .ZN(n7462) );
  AOI21_X1 U8682 ( .B1(n9863), .B2(n9874), .A(n7462), .ZN(n7463) );
  OAI21_X1 U8683 ( .B1(n9858), .B2(n7611), .A(n7463), .ZN(n7464) );
  AOI21_X1 U8684 ( .B1(n10254), .B2(n9837), .A(n7464), .ZN(n7465) );
  OAI21_X1 U8685 ( .B1(n7466), .B2(n9853), .A(n7465), .ZN(P1_U3232) );
  OAI211_X1 U8686 ( .C1(n7469), .C2(n7468), .A(n10443), .B(n7467), .ZN(n7472)
         );
  INV_X1 U8687 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n7530) );
  NAND2_X1 U8688 ( .A1(P1_U3084), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n9794) );
  OAI21_X1 U8689 ( .B1(n10425), .B2(n7530), .A(n9794), .ZN(n7470) );
  INV_X1 U8690 ( .A(n7470), .ZN(n7471) );
  OAI211_X1 U8691 ( .C1(n7473), .C2(n9952), .A(n7472), .B(n7471), .ZN(n7478)
         );
  AOI211_X1 U8692 ( .C1(n7476), .C2(n7475), .A(n7474), .B(n10451), .ZN(n7477)
         );
  OR2_X1 U8693 ( .A1(n7478), .A2(n7477), .ZN(P1_U3257) );
  INV_X1 U8694 ( .A(n8348), .ZN(n7480) );
  XNOR2_X1 U8695 ( .A(n7479), .B(n7480), .ZN(n10261) );
  XOR2_X1 U8696 ( .A(n7481), .B(n8348), .Z(n7483) );
  AOI22_X1 U8697 ( .A1(n9875), .A2(n10141), .B1(n10143), .B2(n9877), .ZN(n7482) );
  OAI21_X1 U8698 ( .B1(n7483), .B2(n9997), .A(n7482), .ZN(n7484) );
  AOI21_X1 U8699 ( .B1(n10261), .B2(n6282), .A(n7484), .ZN(n10265) );
  INV_X1 U8700 ( .A(n7608), .ZN(n7485) );
  AOI211_X1 U8701 ( .C1(n10263), .C2(n7486), .A(n10591), .B(n7485), .ZN(n10262) );
  NOR2_X1 U8702 ( .A1(n5014), .A2(n10115), .ZN(n7489) );
  INV_X1 U8703 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n7487) );
  OAI22_X1 U8704 ( .A1(n10148), .A2(n7487), .B1(n9774), .B2(n10145), .ZN(n7488) );
  AOI211_X1 U8705 ( .C1(n10262), .C2(n10110), .A(n7489), .B(n7488), .ZN(n7491)
         );
  NAND2_X1 U8706 ( .A1(n10261), .A2(n7616), .ZN(n7490) );
  OAI211_X1 U8707 ( .C1(n10265), .C2(n10088), .A(n7491), .B(n7490), .ZN(
        P1_U3279) );
  NOR2_X1 U8708 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n7534) );
  NOR2_X1 U8709 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n7532) );
  NOR2_X1 U8710 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n7529) );
  NOR2_X1 U8711 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n7526) );
  NOR2_X1 U8712 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n7523) );
  NOR2_X1 U8713 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n7520) );
  NAND2_X1 U8714 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(P1_ADDR_REG_11__SCAN_IN), 
        .ZN(n7517) );
  XOR2_X1 U8715 ( .A(P2_ADDR_REG_11__SCAN_IN), .B(P1_ADDR_REG_11__SCAN_IN), 
        .Z(n10386) );
  NAND2_X1 U8716 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(P1_ADDR_REG_10__SCAN_IN), 
        .ZN(n7515) );
  XOR2_X1 U8717 ( .A(P2_ADDR_REG_10__SCAN_IN), .B(P1_ADDR_REG_10__SCAN_IN), 
        .Z(n10384) );
  NOR2_X1 U8718 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n7499) );
  INV_X1 U8719 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n9887) );
  XOR2_X1 U8720 ( .A(n9887), .B(P2_ADDR_REG_4__SCAN_IN), .Z(n10375) );
  NAND2_X1 U8721 ( .A1(P2_ADDR_REG_3__SCAN_IN), .A2(P1_ADDR_REG_3__SCAN_IN), 
        .ZN(n7497) );
  XNOR2_X1 U8722 ( .A(P2_ADDR_REG_3__SCAN_IN), .B(n7492), .ZN(n10373) );
  NAND2_X1 U8723 ( .A1(P1_ADDR_REG_2__SCAN_IN), .A2(P2_ADDR_REG_2__SCAN_IN), 
        .ZN(n7495) );
  XNOR2_X1 U8724 ( .A(n7493), .B(P2_ADDR_REG_2__SCAN_IN), .ZN(n10371) );
  AOI21_X1 U8725 ( .B1(P2_ADDR_REG_0__SCAN_IN), .B2(P1_ADDR_REG_0__SCAN_IN), 
        .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n10365) );
  INV_X1 U8726 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n10369) );
  NAND3_X1 U8727 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .A3(P1_ADDR_REG_0__SCAN_IN), .ZN(n10367) );
  OAI21_X1 U8728 ( .B1(n10365), .B2(n10369), .A(n10367), .ZN(n10370) );
  NAND2_X1 U8729 ( .A1(n10371), .A2(n10370), .ZN(n7494) );
  NAND2_X1 U8730 ( .A1(n7495), .A2(n7494), .ZN(n10372) );
  NAND2_X1 U8731 ( .A1(n10373), .A2(n10372), .ZN(n7496) );
  NAND2_X1 U8732 ( .A1(n7497), .A2(n7496), .ZN(n10374) );
  NOR2_X1 U8733 ( .A1(n10375), .A2(n10374), .ZN(n7498) );
  NOR2_X1 U8734 ( .A1(n7499), .A2(n7498), .ZN(n7500) );
  NOR2_X1 U8735 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n7500), .ZN(n10377) );
  AND2_X1 U8736 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n7500), .ZN(n10376) );
  NOR2_X1 U8737 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n10376), .ZN(n7501) );
  NAND2_X1 U8738 ( .A1(P1_ADDR_REG_6__SCAN_IN), .A2(n7502), .ZN(n7504) );
  XOR2_X1 U8739 ( .A(P1_ADDR_REG_6__SCAN_IN), .B(n7502), .Z(n10379) );
  NAND2_X1 U8740 ( .A1(P2_ADDR_REG_6__SCAN_IN), .A2(n10379), .ZN(n7503) );
  NAND2_X1 U8741 ( .A1(n7504), .A2(n7503), .ZN(n7505) );
  NAND2_X1 U8742 ( .A1(P1_ADDR_REG_7__SCAN_IN), .A2(n7505), .ZN(n7507) );
  XOR2_X1 U8743 ( .A(P1_ADDR_REG_7__SCAN_IN), .B(n7505), .Z(n10380) );
  NAND2_X1 U8744 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(n10380), .ZN(n7506) );
  NAND2_X1 U8745 ( .A1(n7507), .A2(n7506), .ZN(n7508) );
  NAND2_X1 U8746 ( .A1(P1_ADDR_REG_8__SCAN_IN), .A2(n7508), .ZN(n7510) );
  XOR2_X1 U8747 ( .A(P1_ADDR_REG_8__SCAN_IN), .B(n7508), .Z(n10381) );
  NAND2_X1 U8748 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(n10381), .ZN(n7509) );
  NAND2_X1 U8749 ( .A1(n7510), .A2(n7509), .ZN(n7511) );
  NAND2_X1 U8750 ( .A1(P1_ADDR_REG_9__SCAN_IN), .A2(n7511), .ZN(n7513) );
  XOR2_X1 U8751 ( .A(P1_ADDR_REG_9__SCAN_IN), .B(n7511), .Z(n10382) );
  NAND2_X1 U8752 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(n10382), .ZN(n7512) );
  NAND2_X1 U8753 ( .A1(n7513), .A2(n7512), .ZN(n10383) );
  NAND2_X1 U8754 ( .A1(n10384), .A2(n10383), .ZN(n7514) );
  NAND2_X1 U8755 ( .A1(n7515), .A2(n7514), .ZN(n10385) );
  NAND2_X1 U8756 ( .A1(n10386), .A2(n10385), .ZN(n7516) );
  NAND2_X1 U8757 ( .A1(n7517), .A2(n7516), .ZN(n10388) );
  XOR2_X1 U8758 ( .A(P2_ADDR_REG_12__SCAN_IN), .B(n7518), .Z(n10387) );
  XOR2_X1 U8759 ( .A(n7521), .B(P1_ADDR_REG_13__SCAN_IN), .Z(n10389) );
  XOR2_X1 U8760 ( .A(P2_ADDR_REG_14__SCAN_IN), .B(n7524), .Z(n10391) );
  XOR2_X1 U8761 ( .A(P2_ADDR_REG_15__SCAN_IN), .B(n7527), .Z(n10393) );
  NOR2_X1 U8762 ( .A1(n10394), .A2(n10393), .ZN(n7528) );
  NOR2_X1 U8763 ( .A1(n7529), .A2(n7528), .ZN(n10396) );
  XOR2_X1 U8764 ( .A(P2_ADDR_REG_16__SCAN_IN), .B(n7530), .Z(n10395) );
  NOR2_X1 U8765 ( .A1(n10396), .A2(n10395), .ZN(n7531) );
  NOR2_X1 U8766 ( .A1(n7532), .A2(n7531), .ZN(n10398) );
  INV_X1 U8767 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n7753) );
  XOR2_X1 U8768 ( .A(P2_ADDR_REG_17__SCAN_IN), .B(n7753), .Z(n10397) );
  NOR2_X1 U8769 ( .A1(n10398), .A2(n10397), .ZN(n7533) );
  NOR2_X1 U8770 ( .A1(n7534), .A2(n7533), .ZN(n7535) );
  AND2_X1 U8771 ( .A1(P2_ADDR_REG_18__SCAN_IN), .A2(n7535), .ZN(n10399) );
  NOR2_X1 U8772 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(n10399), .ZN(n7536) );
  NOR2_X1 U8773 ( .A1(P2_ADDR_REG_18__SCAN_IN), .A2(n7535), .ZN(n10400) );
  NOR2_X1 U8774 ( .A1(n7536), .A2(n10400), .ZN(n7538) );
  XNOR2_X1 U8775 ( .A(P1_ADDR_REG_19__SCAN_IN), .B(P2_ADDR_REG_19__SCAN_IN), 
        .ZN(n7537) );
  XNOR2_X1 U8776 ( .A(n7538), .B(n7537), .ZN(ADD_1071_U4) );
  INV_X1 U8777 ( .A(n8709), .ZN(n7584) );
  OAI222_X1 U8778 ( .A1(n6276), .A2(n7584), .B1(n8101), .B2(n7540), .C1(n7539), 
        .C2(P1_U3084), .ZN(P1_U3327) );
  OAI21_X1 U8779 ( .B1(n7543), .B2(n7542), .A(n7541), .ZN(n7545) );
  NAND2_X1 U8780 ( .A1(n7543), .A2(n7542), .ZN(n7544) );
  NAND2_X1 U8781 ( .A1(n7545), .A2(n7544), .ZN(n7673) );
  NAND2_X1 U8782 ( .A1(n8271), .A2(n6216), .ZN(n7547) );
  OR2_X1 U8783 ( .A1(n8275), .A2(n6305), .ZN(n7546) );
  NAND2_X1 U8784 ( .A1(n7547), .A2(n7546), .ZN(n7672) );
  NAND2_X1 U8785 ( .A1(n8271), .A2(n8207), .ZN(n7549) );
  OR2_X1 U8786 ( .A1(n8275), .A2(n8208), .ZN(n7548) );
  NAND2_X1 U8787 ( .A1(n7549), .A2(n7548), .ZN(n7550) );
  XNOR2_X1 U8788 ( .A(n7550), .B(n6585), .ZN(n7671) );
  XOR2_X1 U8789 ( .A(n7672), .B(n7671), .Z(n7551) );
  XNOR2_X1 U8790 ( .A(n7673), .B(n7551), .ZN(n7557) );
  OAI21_X1 U8791 ( .B1(n9860), .B2(n7693), .A(n7552), .ZN(n7553) );
  AOI21_X1 U8792 ( .B1(n9863), .B2(n9873), .A(n7553), .ZN(n7554) );
  OAI21_X1 U8793 ( .B1(n9858), .B2(n7698), .A(n7554), .ZN(n7555) );
  AOI21_X1 U8794 ( .B1(n8271), .B2(n9837), .A(n7555), .ZN(n7556) );
  OAI21_X1 U8795 ( .B1(n7557), .B2(n9853), .A(n7556), .ZN(P1_U3213) );
  NAND2_X1 U8796 ( .A1(n7651), .A2(n9033), .ZN(n7559) );
  INV_X1 U8797 ( .A(n7559), .ZN(n7558) );
  OR2_X1 U8798 ( .A1(n7651), .A2(n7768), .ZN(n8615) );
  NAND2_X1 U8799 ( .A1(n7651), .A2(n7768), .ZN(n8611) );
  NAND2_X1 U8800 ( .A1(n8615), .A2(n8611), .ZN(n8772) );
  OR2_X1 U8801 ( .A1(n7558), .A2(n8772), .ZN(n7564) );
  INV_X1 U8802 ( .A(n7564), .ZN(n7561) );
  INV_X1 U8803 ( .A(n7562), .ZN(n9034) );
  NAND2_X1 U8804 ( .A1(n7563), .A2(n9034), .ZN(n7643) );
  AND2_X1 U8805 ( .A1(n7643), .A2(n7559), .ZN(n7560) );
  NOR2_X1 U8806 ( .A1(n7561), .A2(n7560), .ZN(n7567) );
  OR2_X1 U8807 ( .A1(n8770), .A2(n7567), .ZN(n7568) );
  OR2_X1 U8808 ( .A1(n7563), .A2(n7562), .ZN(n8614) );
  NAND2_X1 U8809 ( .A1(n7563), .A2(n7562), .ZN(n8612) );
  NAND2_X1 U8810 ( .A1(n8614), .A2(n8612), .ZN(n8773) );
  AND2_X1 U8811 ( .A1(n8773), .A2(n7564), .ZN(n7565) );
  OR2_X1 U8812 ( .A1(n7587), .A2(n9035), .ZN(n7641) );
  AND2_X1 U8813 ( .A1(n7565), .A2(n7641), .ZN(n7566) );
  INV_X1 U8814 ( .A(n7662), .ZN(n7570) );
  OR2_X1 U8815 ( .A1(n10633), .A2(n7657), .ZN(n8628) );
  NAND2_X1 U8816 ( .A1(n10633), .A2(n7657), .ZN(n7655) );
  XNOR2_X1 U8817 ( .A(n7570), .B(n8776), .ZN(n10640) );
  NAND2_X1 U8818 ( .A1(n7775), .A2(n10626), .ZN(n7571) );
  NAND2_X1 U8819 ( .A1(n7571), .A2(n10633), .ZN(n7572) );
  NAND2_X1 U8820 ( .A1(n7664), .A2(n7572), .ZN(n10636) );
  AOI22_X1 U8821 ( .A1(n9354), .A2(P2_REG2_REG_12__SCAN_IN), .B1(n7573), .B2(
        n9350), .ZN(n7575) );
  NAND2_X1 U8822 ( .A1(n9336), .A2(n10633), .ZN(n7574) );
  OAI211_X1 U8823 ( .C1(n10636), .C2(n9139), .A(n7575), .B(n7574), .ZN(n7582)
         );
  INV_X1 U8824 ( .A(n8608), .ZN(n8625) );
  NOR2_X1 U8825 ( .A1(n8773), .A2(n8625), .ZN(n7576) );
  NAND2_X1 U8826 ( .A1(n7763), .A2(n7576), .ZN(n7765) );
  NAND2_X1 U8827 ( .A1(n7765), .A2(n8612), .ZN(n7654) );
  NAND2_X1 U8828 ( .A1(n7654), .A2(n8615), .ZN(n7577) );
  NAND2_X1 U8829 ( .A1(n7577), .A2(n8611), .ZN(n7578) );
  XNOR2_X1 U8830 ( .A(n7578), .B(n8776), .ZN(n7580) );
  OAI22_X1 U8831 ( .A1(n7825), .A2(n9318), .B1(n7768), .B2(n9320), .ZN(n7579)
         );
  AOI21_X1 U8832 ( .B1(n7580), .B2(n9340), .A(n7579), .ZN(n10635) );
  NOR2_X1 U8833 ( .A1(n10635), .A2(n9354), .ZN(n7581) );
  AOI211_X1 U8834 ( .C1(n10640), .C2(n9337), .A(n7582), .B(n7581), .ZN(n7583)
         );
  INV_X1 U8835 ( .A(n7583), .ZN(P2_U3284) );
  INV_X1 U8836 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n8710) );
  OAI222_X1 U8837 ( .A1(n7585), .A2(P2_U3152), .B1(n8039), .B2(n7584), .C1(
        n8710), .C2(n9710), .ZN(P2_U3332) );
  INV_X1 U8838 ( .A(n7586), .ZN(n7592) );
  AOI22_X1 U8839 ( .A1(n7588), .A2(n10511), .B1(n10632), .B2(n7587), .ZN(n7589) );
  OAI211_X1 U8840 ( .C1(n7592), .C2(n7591), .A(n7590), .B(n7589), .ZN(n7595)
         );
  NAND2_X1 U8841 ( .A1(n7595), .A2(n10642), .ZN(n7593) );
  OAI21_X1 U8842 ( .B1(n10642), .B2(n7594), .A(n7593), .ZN(P2_U3529) );
  INV_X1 U8843 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n7597) );
  NAND2_X1 U8844 ( .A1(n7595), .A2(n10646), .ZN(n7596) );
  OAI21_X1 U8845 ( .B1(n10646), .B2(n7597), .A(n7596), .ZN(P2_U3478) );
  NAND2_X1 U8846 ( .A1(n7598), .A2(n8351), .ZN(n7599) );
  NAND2_X1 U8847 ( .A1(n7600), .A2(n7599), .ZN(n10258) );
  NAND2_X1 U8848 ( .A1(n10258), .A2(n6282), .ZN(n7607) );
  OAI21_X1 U8849 ( .B1(n8351), .B2(n7602), .A(n7601), .ZN(n7605) );
  OAI22_X1 U8850 ( .A1(n8275), .A2(n10103), .B1(n7603), .B2(n10101), .ZN(n7604) );
  AOI21_X1 U8851 ( .B1(n7605), .B2(n10140), .A(n7604), .ZN(n7606) );
  INV_X1 U8852 ( .A(n7697), .ZN(n7610) );
  NAND2_X1 U8853 ( .A1(n7608), .A2(n10254), .ZN(n7609) );
  NAND2_X1 U8854 ( .A1(n7610), .A2(n7609), .ZN(n10256) );
  INV_X1 U8855 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n7612) );
  OAI22_X1 U8856 ( .A1(n10148), .A2(n7612), .B1(n7611), .B2(n10145), .ZN(n7613) );
  AOI21_X1 U8857 ( .B1(n10254), .B2(n10156), .A(n7613), .ZN(n7614) );
  OAI21_X1 U8858 ( .B1(n10256), .B2(n10152), .A(n7614), .ZN(n7615) );
  AOI21_X1 U8859 ( .B1(n10258), .B2(n7616), .A(n7615), .ZN(n7617) );
  OAI21_X1 U8860 ( .B1(n10260), .B2(n10088), .A(n7617), .ZN(P1_U3278) );
  NAND2_X1 U8861 ( .A1(n7621), .A2(n8727), .ZN(n7624) );
  AOI22_X1 U8862 ( .A1(n7997), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n7996), .B2(
        n7622), .ZN(n7623) );
  XNOR2_X1 U8863 ( .A(n9451), .B(n8933), .ZN(n7710) );
  NOR2_X1 U8864 ( .A1(n7825), .A2(n8932), .ZN(n7708) );
  XNOR2_X1 U8865 ( .A(n7710), .B(n7708), .ZN(n7706) );
  XNOR2_X1 U8866 ( .A(n7707), .B(n7706), .ZN(n7637) );
  INV_X1 U8867 ( .A(n7657), .ZN(n9032) );
  AOI22_X1 U8868 ( .A1(n8947), .A2(n9032), .B1(n7666), .B2(n8949), .ZN(n7635)
         );
  INV_X1 U8869 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n7625) );
  NAND2_X1 U8870 ( .A1(n7626), .A2(n7625), .ZN(n7627) );
  AND2_X1 U8871 ( .A1(n7715), .A2(n7627), .ZN(n7820) );
  NAND2_X1 U8872 ( .A1(n6556), .A2(n7820), .ZN(n7631) );
  NAND2_X1 U8873 ( .A1(n6560), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n7630) );
  NAND2_X1 U8874 ( .A1(n6554), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n7629) );
  NAND2_X1 U8875 ( .A1(n6555), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n7628) );
  INV_X1 U8876 ( .A(n7818), .ZN(n9030) );
  INV_X1 U8877 ( .A(n7632), .ZN(n7633) );
  AOI21_X1 U8878 ( .B1(n9005), .B2(n9030), .A(n7633), .ZN(n7634) );
  OAI211_X1 U8879 ( .C1(n4997), .C2(n8937), .A(n7635), .B(n7634), .ZN(n7636)
         );
  AOI21_X1 U8880 ( .B1(n7637), .B2(n8941), .A(n7636), .ZN(n7638) );
  INV_X1 U8881 ( .A(n7638), .ZN(P2_U3236) );
  INV_X1 U8882 ( .A(n8772), .ZN(n7639) );
  XNOR2_X1 U8883 ( .A(n7654), .B(n7639), .ZN(n7640) );
  NAND2_X1 U8884 ( .A1(n7640), .A2(n9340), .ZN(n10624) );
  NAND2_X1 U8885 ( .A1(n7762), .A2(n8773), .ZN(n7761) );
  NAND2_X1 U8886 ( .A1(n7761), .A2(n7643), .ZN(n7644) );
  XOR2_X1 U8887 ( .A(n8772), .B(n7644), .Z(n10628) );
  NAND2_X1 U8888 ( .A1(n10628), .A2(n9337), .ZN(n7653) );
  INV_X1 U8889 ( .A(n7645), .ZN(n7646) );
  OAI22_X1 U8890 ( .A1(n9307), .A2(n6705), .B1(n7646), .B2(n9304), .ZN(n7650)
         );
  XNOR2_X1 U8891 ( .A(n7775), .B(n7651), .ZN(n7647) );
  AOI222_X1 U8892 ( .A1(n9034), .A2(n9345), .B1(n10511), .B2(n7647), .C1(n9032), .C2(n9346), .ZN(n10623) );
  NOR2_X1 U8893 ( .A1(n10623), .A2(n7648), .ZN(n7649) );
  AOI211_X1 U8894 ( .C1(n9336), .C2(n7651), .A(n7650), .B(n7649), .ZN(n7652)
         );
  OAI211_X1 U8895 ( .C1(n9354), .C2(n10624), .A(n7653), .B(n7652), .ZN(
        P2_U3285) );
  NAND2_X1 U8896 ( .A1(n7655), .A2(n8611), .ZN(n8629) );
  NAND2_X1 U8897 ( .A1(n8628), .A2(n8615), .ZN(n7656) );
  NAND2_X1 U8898 ( .A1(n7656), .A2(n7655), .ZN(n8630) );
  OR2_X1 U8899 ( .A1(n9451), .A2(n7825), .ZN(n8634) );
  NAND2_X1 U8900 ( .A1(n9451), .A2(n7825), .ZN(n8635) );
  XNOR2_X1 U8901 ( .A(n7986), .B(n7892), .ZN(n7659) );
  OAI22_X1 U8902 ( .A1(n7818), .A2(n9318), .B1(n7657), .B2(n9320), .ZN(n7658)
         );
  AOI21_X1 U8903 ( .B1(n7659), .B2(n9340), .A(n7658), .ZN(n9454) );
  INV_X1 U8904 ( .A(n8776), .ZN(n7661) );
  INV_X1 U8905 ( .A(n7915), .ZN(n7663) );
  OR2_X1 U8906 ( .A1(n7663), .A2(n8777), .ZN(n7817) );
  OAI21_X1 U8907 ( .B1(n7915), .B2(n7892), .A(n7817), .ZN(n9455) );
  OR2_X1 U8908 ( .A1(n9455), .A2(n9285), .ZN(n7670) );
  NAND2_X1 U8909 ( .A1(n7664), .A2(n9451), .ZN(n7665) );
  AND2_X1 U8910 ( .A1(n7819), .A2(n7665), .ZN(n9452) );
  AOI22_X1 U8911 ( .A1(n9354), .A2(P2_REG2_REG_13__SCAN_IN), .B1(n7666), .B2(
        n9350), .ZN(n7667) );
  OAI21_X1 U8912 ( .B1(n4997), .B2(n9272), .A(n7667), .ZN(n7668) );
  AOI21_X1 U8913 ( .B1(n9452), .B2(n9353), .A(n7668), .ZN(n7669) );
  OAI211_X1 U8914 ( .C1(n9223), .C2(n9454), .A(n7670), .B(n7669), .ZN(P2_U3283) );
  OAI21_X1 U8915 ( .B1(n7673), .B2(n7672), .A(n7671), .ZN(n7675) );
  NAND2_X1 U8916 ( .A1(n7673), .A2(n7672), .ZN(n7674) );
  NAND2_X1 U8917 ( .A1(n7675), .A2(n7674), .ZN(n8106) );
  NAND2_X1 U8918 ( .A1(n7809), .A2(n6216), .ZN(n7677) );
  OR2_X1 U8919 ( .A1(n7878), .A2(n6305), .ZN(n7676) );
  NAND2_X1 U8920 ( .A1(n7677), .A2(n7676), .ZN(n8104) );
  NAND2_X1 U8921 ( .A1(n7809), .A2(n8207), .ZN(n7679) );
  OR2_X1 U8922 ( .A1(n7878), .A2(n8208), .ZN(n7678) );
  NAND2_X1 U8923 ( .A1(n7679), .A2(n7678), .ZN(n7680) );
  XNOR2_X1 U8924 ( .A(n7680), .B(n8195), .ZN(n8105) );
  XOR2_X1 U8925 ( .A(n8104), .B(n8105), .Z(n7681) );
  XNOR2_X1 U8926 ( .A(n8106), .B(n7681), .ZN(n7687) );
  OAI21_X1 U8927 ( .B1(n9860), .B2(n8275), .A(n7682), .ZN(n7683) );
  AOI21_X1 U8928 ( .B1(n9863), .B2(n10144), .A(n7683), .ZN(n7684) );
  OAI21_X1 U8929 ( .B1(n9858), .B2(n7810), .A(n7684), .ZN(n7685) );
  AOI21_X1 U8930 ( .B1(n7809), .B2(n9837), .A(n7685), .ZN(n7686) );
  OAI21_X1 U8931 ( .B1(n7687), .B2(n9853), .A(n7686), .ZN(P1_U3239) );
  INV_X1 U8932 ( .A(n8715), .ZN(n8103) );
  INV_X1 U8933 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n8716) );
  OAI222_X1 U8934 ( .A1(P2_U3152), .A2(n8824), .B1(n8039), .B2(n8103), .C1(
        n8716), .C2(n8230), .ZN(P2_U3331) );
  OAI21_X1 U8935 ( .B1(n7689), .B2(n7690), .A(n7688), .ZN(n10247) );
  INV_X1 U8936 ( .A(n10247), .ZN(n7705) );
  INV_X1 U8937 ( .A(n7690), .ZN(n8349) );
  XNOR2_X1 U8938 ( .A(n7691), .B(n8349), .ZN(n7692) );
  NAND2_X1 U8939 ( .A1(n7692), .A2(n10140), .ZN(n7696) );
  OAI22_X1 U8940 ( .A1(n7878), .A2(n10103), .B1(n7693), .B2(n10101), .ZN(n7694) );
  INV_X1 U8941 ( .A(n7694), .ZN(n7695) );
  NAND2_X1 U8942 ( .A1(n7696), .A2(n7695), .ZN(n10251) );
  OAI211_X1 U8943 ( .C1(n7697), .C2(n10249), .A(n5984), .B(n7808), .ZN(n10248)
         );
  OAI22_X1 U8944 ( .A1(n10148), .A2(n7699), .B1(n7698), .B2(n10145), .ZN(n7700) );
  AOI21_X1 U8945 ( .B1(n8271), .B2(n10156), .A(n7700), .ZN(n7701) );
  OAI21_X1 U8946 ( .B1(n10248), .B2(n7702), .A(n7701), .ZN(n7703) );
  AOI21_X1 U8947 ( .B1(n10251), .B2(n10148), .A(n7703), .ZN(n7704) );
  OAI21_X1 U8948 ( .B1(n7705), .B2(n10137), .A(n7704), .ZN(P1_U3277) );
  INV_X1 U8949 ( .A(n7708), .ZN(n7709) );
  OR2_X1 U8950 ( .A1(n7711), .A2(n6564), .ZN(n7713) );
  AOI22_X1 U8951 ( .A1(n7997), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n7996), .B2(
        n7738), .ZN(n7712) );
  XNOR2_X1 U8952 ( .A(n9446), .B(n8933), .ZN(n7786) );
  NOR2_X1 U8953 ( .A1(n7818), .A2(n8932), .ZN(n7784) );
  XNOR2_X1 U8954 ( .A(n7786), .B(n7784), .ZN(n7782) );
  XOR2_X1 U8955 ( .A(n7783), .B(n7782), .Z(n7725) );
  NAND2_X1 U8956 ( .A1(n6554), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n7720) );
  INV_X1 U8957 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n7714) );
  NAND2_X1 U8958 ( .A1(n7715), .A2(n7714), .ZN(n7716) );
  AND2_X1 U8959 ( .A1(n7793), .A2(n7716), .ZN(n7982) );
  NAND2_X1 U8960 ( .A1(n6556), .A2(n7982), .ZN(n7719) );
  NAND2_X1 U8961 ( .A1(n6560), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n7718) );
  NAND2_X1 U8962 ( .A1(n6555), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n7717) );
  INV_X1 U8963 ( .A(n7884), .ZN(n9029) );
  AOI22_X1 U8964 ( .A1(n9005), .A2(n9029), .B1(n7820), .B2(n8949), .ZN(n7722)
         );
  OAI211_X1 U8965 ( .C1(n9014), .C2(n7825), .A(n7722), .B(n7721), .ZN(n7723)
         );
  AOI21_X1 U8966 ( .B1(n9446), .B2(n9017), .A(n7723), .ZN(n7724) );
  OAI21_X1 U8967 ( .B1(n7725), .B2(n9019), .A(n7724), .ZN(P2_U3217) );
  INV_X1 U8968 ( .A(n8728), .ZN(n8231) );
  AOI21_X1 U8969 ( .B1(n10324), .B2(P2_DATAO_REG_28__SCAN_IN), .A(n7726), .ZN(
        n7727) );
  OAI21_X1 U8970 ( .B1(n8231), .B2(n6276), .A(n7727), .ZN(P1_U3325) );
  AOI21_X1 U8971 ( .B1(n7730), .B2(n7729), .A(n7728), .ZN(n7731) );
  NAND2_X1 U8972 ( .A1(n9064), .A2(n7731), .ZN(n7732) );
  XNOR2_X1 U8973 ( .A(n7731), .B(n7739), .ZN(n9061) );
  NAND2_X1 U8974 ( .A1(P2_REG1_REG_15__SCAN_IN), .A2(n9061), .ZN(n9060) );
  NAND2_X1 U8975 ( .A1(n7732), .A2(n9060), .ZN(n7734) );
  XNOR2_X1 U8976 ( .A(n7855), .B(P2_REG1_REG_16__SCAN_IN), .ZN(n7733) );
  NOR2_X1 U8977 ( .A1(n7734), .A2(n7733), .ZN(n7837) );
  AOI21_X1 U8978 ( .B1(n7734), .B2(n7733), .A(n7837), .ZN(n7748) );
  NOR2_X1 U8979 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7792), .ZN(n7735) );
  AOI21_X1 U8980 ( .B1(n10486), .B2(P2_ADDR_REG_16__SCAN_IN), .A(n7735), .ZN(
        n7736) );
  INV_X1 U8981 ( .A(n7736), .ZN(n7746) );
  OAI21_X1 U8982 ( .B1(n7738), .B2(P2_REG2_REG_14__SCAN_IN), .A(n7737), .ZN(
        n7740) );
  NAND2_X1 U8983 ( .A1(n7739), .A2(n7740), .ZN(n7741) );
  XNOR2_X1 U8984 ( .A(n7740), .B(n9064), .ZN(n9058) );
  INV_X1 U8985 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n9057) );
  NAND2_X1 U8986 ( .A1(n9058), .A2(n9057), .ZN(n9056) );
  NAND2_X1 U8987 ( .A1(n7741), .A2(n9056), .ZN(n7744) );
  NAND2_X1 U8988 ( .A1(n7855), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n7742) );
  OAI21_X1 U8989 ( .B1(n7855), .B2(P2_REG2_REG_16__SCAN_IN), .A(n7742), .ZN(
        n7743) );
  NOR2_X1 U8990 ( .A1(n7744), .A2(n7743), .ZN(n7832) );
  AOI211_X1 U8991 ( .C1(n7744), .C2(n7743), .A(n7832), .B(n10487), .ZN(n7745)
         );
  AOI211_X1 U8992 ( .C1(n10493), .C2(n7855), .A(n7746), .B(n7745), .ZN(n7747)
         );
  OAI21_X1 U8993 ( .B1(n7748), .B2(n10468), .A(n7747), .ZN(P2_U3261) );
  OAI211_X1 U8994 ( .C1(n7751), .C2(n7750), .A(n7749), .B(n10443), .ZN(n7752)
         );
  NAND2_X1 U8995 ( .A1(P1_U3084), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n9806) );
  OAI211_X1 U8996 ( .C1(n7753), .C2(n10425), .A(n7752), .B(n9806), .ZN(n7758)
         );
  AOI211_X1 U8997 ( .C1(n7756), .C2(n7755), .A(n7754), .B(n10451), .ZN(n7757)
         );
  AOI211_X1 U8998 ( .C1(n10459), .C2(n7759), .A(n7758), .B(n7757), .ZN(n7760)
         );
  INV_X1 U8999 ( .A(n7760), .ZN(P1_U3258) );
  OAI21_X1 U9000 ( .B1(n7762), .B2(n8773), .A(n7761), .ZN(n10613) );
  NAND2_X1 U9001 ( .A1(n7763), .A2(n8608), .ZN(n7764) );
  NAND2_X1 U9002 ( .A1(n7764), .A2(n8773), .ZN(n7766) );
  NAND2_X1 U9003 ( .A1(n7766), .A2(n7765), .ZN(n7770) );
  OAI22_X1 U9004 ( .A1(n7768), .A2(n9318), .B1(n7767), .B2(n9320), .ZN(n7769)
         );
  AOI21_X1 U9005 ( .B1(n7770), .B2(n9340), .A(n7769), .ZN(n7771) );
  OAI21_X1 U9006 ( .B1(n10613), .B2(n9302), .A(n7771), .ZN(n10616) );
  MUX2_X1 U9007 ( .A(P2_REG2_REG_10__SCAN_IN), .B(n10616), .S(n9307), .Z(n7772) );
  INV_X1 U9008 ( .A(n7772), .ZN(n7781) );
  NOR2_X1 U9009 ( .A1(n7773), .A2(n10614), .ZN(n7774) );
  OR2_X1 U9010 ( .A1(n7775), .A2(n7774), .ZN(n10615) );
  INV_X1 U9011 ( .A(n10615), .ZN(n7779) );
  INV_X1 U9012 ( .A(n7776), .ZN(n7777) );
  OAI22_X1 U9013 ( .A1(n9272), .A2(n10614), .B1(n9304), .B2(n7777), .ZN(n7778)
         );
  AOI21_X1 U9014 ( .B1(n7779), .B2(n9353), .A(n7778), .ZN(n7780) );
  OAI211_X1 U9015 ( .C1(n10613), .C2(n9311), .A(n7781), .B(n7780), .ZN(
        P2_U3286) );
  NAND2_X1 U9016 ( .A1(n7783), .A2(n7782), .ZN(n7788) );
  INV_X1 U9017 ( .A(n7784), .ZN(n7785) );
  NAND2_X1 U9018 ( .A1(n7786), .A2(n7785), .ZN(n7787) );
  NAND2_X1 U9019 ( .A1(n7788), .A2(n7787), .ZN(n7848) );
  OR2_X1 U9020 ( .A1(n7789), .A2(n6564), .ZN(n7791) );
  AOI22_X1 U9021 ( .A1(n7997), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n7996), .B2(
        n9064), .ZN(n7790) );
  XNOR2_X1 U9022 ( .A(n9441), .B(n8933), .ZN(n7851) );
  NOR2_X1 U9023 ( .A1(n7884), .A2(n8932), .ZN(n7849) );
  XNOR2_X1 U9024 ( .A(n7851), .B(n7849), .ZN(n7847) );
  XOR2_X1 U9025 ( .A(n7848), .B(n7847), .Z(n7802) );
  NAND2_X1 U9026 ( .A1(n7793), .A2(n7792), .ZN(n7794) );
  AND2_X1 U9027 ( .A1(n7858), .A2(n7794), .ZN(n7889) );
  NAND2_X1 U9028 ( .A1(n6556), .A2(n7889), .ZN(n7798) );
  NAND2_X1 U9029 ( .A1(n6560), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n7797) );
  NAND2_X1 U9030 ( .A1(n6554), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n7796) );
  NAND2_X1 U9031 ( .A1(n6555), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n7795) );
  AOI22_X1 U9032 ( .A1(n8947), .A2(n9030), .B1(n7982), .B2(n8949), .ZN(n7799)
         );
  NAND2_X1 U9033 ( .A1(P2_REG3_REG_15__SCAN_IN), .A2(P2_U3152), .ZN(n9062) );
  OAI211_X1 U9034 ( .C1(n9011), .C2(n7970), .A(n7799), .B(n9062), .ZN(n7800)
         );
  AOI21_X1 U9035 ( .B1(n9441), .B2(n9017), .A(n7800), .ZN(n7801) );
  OAI21_X1 U9036 ( .B1(n7802), .B2(n9019), .A(n7801), .ZN(P2_U3243) );
  INV_X1 U9037 ( .A(n7803), .ZN(n7804) );
  AOI21_X1 U9038 ( .B1(n8352), .B2(n7805), .A(n7804), .ZN(n10243) );
  INV_X1 U9039 ( .A(n10243), .ZN(n7816) );
  XNOR2_X1 U9040 ( .A(n7806), .B(n8352), .ZN(n7807) );
  OAI222_X1 U9041 ( .A1(n10103), .A2(n8110), .B1(n10101), .B2(n8275), .C1(
        n9997), .C2(n7807), .ZN(n10241) );
  INV_X1 U9042 ( .A(n7809), .ZN(n10312) );
  AOI211_X1 U9043 ( .C1(n7809), .C2(n7808), .A(n10591), .B(n5949), .ZN(n10242)
         );
  NAND2_X1 U9044 ( .A1(n10242), .A2(n10110), .ZN(n7813) );
  INV_X1 U9045 ( .A(n7810), .ZN(n7811) );
  AOI22_X1 U9046 ( .A1(n10088), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n7811), .B2(
        n10111), .ZN(n7812) );
  OAI211_X1 U9047 ( .C1(n10312), .C2(n10115), .A(n7813), .B(n7812), .ZN(n7814)
         );
  AOI21_X1 U9048 ( .B1(n10241), .B2(n10148), .A(n7814), .ZN(n7815) );
  OAI21_X1 U9049 ( .B1(n7816), .B2(n10137), .A(n7815), .ZN(P1_U3276) );
  INV_X1 U9050 ( .A(n7825), .ZN(n9031) );
  NAND2_X1 U9051 ( .A1(n9451), .A2(n9031), .ZN(n7910) );
  NAND2_X1 U9052 ( .A1(n7817), .A2(n7910), .ZN(n7882) );
  OR2_X1 U9053 ( .A1(n9446), .A2(n7818), .ZN(n8638) );
  NAND2_X1 U9054 ( .A1(n9446), .A2(n7818), .ZN(n8639) );
  INV_X1 U9055 ( .A(n8778), .ZN(n7911) );
  XNOR2_X1 U9056 ( .A(n7882), .B(n7911), .ZN(n9450) );
  AOI21_X1 U9057 ( .B1(n9446), .B2(n7819), .A(n7979), .ZN(n9447) );
  INV_X1 U9058 ( .A(n9446), .ZN(n7822) );
  AOI22_X1 U9059 ( .A1(n9223), .A2(P2_REG2_REG_14__SCAN_IN), .B1(n7820), .B2(
        n9350), .ZN(n7821) );
  OAI21_X1 U9060 ( .B1(n7822), .B2(n9272), .A(n7821), .ZN(n7830) );
  OR2_X1 U9061 ( .A1(n7986), .A2(n7892), .ZN(n7824) );
  NAND2_X1 U9062 ( .A1(n7824), .A2(n8635), .ZN(n7823) );
  AOI21_X1 U9063 ( .B1(n7823), .B2(n7911), .A(n9253), .ZN(n7828) );
  AND2_X1 U9064 ( .A1(n8778), .A2(n8635), .ZN(n7893) );
  NAND2_X1 U9065 ( .A1(n7824), .A2(n7893), .ZN(n7827) );
  OAI22_X1 U9066 ( .A1(n7884), .A2(n9318), .B1(n7825), .B2(n9320), .ZN(n7826)
         );
  AOI21_X1 U9067 ( .B1(n7828), .B2(n7827), .A(n7826), .ZN(n9449) );
  NOR2_X1 U9068 ( .A1(n9449), .A2(n9354), .ZN(n7829) );
  AOI211_X1 U9069 ( .C1(n9447), .C2(n9353), .A(n7830), .B(n7829), .ZN(n7831)
         );
  OAI21_X1 U9070 ( .B1(n9450), .B2(n9285), .A(n7831), .ZN(P2_U3282) );
  NAND2_X1 U9071 ( .A1(n9076), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n7833) );
  OAI21_X1 U9072 ( .B1(n9076), .B2(P2_REG2_REG_17__SCAN_IN), .A(n7833), .ZN(
        n7834) );
  NOR2_X1 U9073 ( .A1(n7835), .A2(n7834), .ZN(n9070) );
  AOI211_X1 U9074 ( .C1(n7835), .C2(n7834), .A(n9070), .B(n10487), .ZN(n7846)
         );
  INV_X1 U9075 ( .A(n9076), .ZN(n7844) );
  INV_X1 U9076 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n9671) );
  NOR2_X1 U9077 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9671), .ZN(n7836) );
  AOI21_X1 U9078 ( .B1(n10486), .B2(P2_ADDR_REG_17__SCAN_IN), .A(n7836), .ZN(
        n7843) );
  XOR2_X1 U9079 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n9076), .Z(n7841) );
  OR2_X1 U9080 ( .A1(n7855), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n7839) );
  INV_X1 U9081 ( .A(n7837), .ZN(n7838) );
  AND2_X1 U9082 ( .A1(n7839), .A2(n7838), .ZN(n7840) );
  NAND2_X1 U9083 ( .A1(n7841), .A2(n7840), .ZN(n9074) );
  OAI211_X1 U9084 ( .C1(n7841), .C2(n7840), .A(n10495), .B(n9074), .ZN(n7842)
         );
  OAI211_X1 U9085 ( .C1(n10467), .C2(n7844), .A(n7843), .B(n7842), .ZN(n7845)
         );
  OR2_X1 U9086 ( .A1(n7846), .A2(n7845), .ZN(P2_U3262) );
  NAND2_X1 U9087 ( .A1(n7848), .A2(n7847), .ZN(n7853) );
  INV_X1 U9088 ( .A(n7849), .ZN(n7850) );
  NAND2_X1 U9089 ( .A1(n7851), .A2(n7850), .ZN(n7852) );
  NAND2_X1 U9090 ( .A1(n7853), .A2(n7852), .ZN(n7957) );
  AOI22_X1 U9091 ( .A1(n7997), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n7996), .B2(
        n7855), .ZN(n7856) );
  XNOR2_X1 U9092 ( .A(n9437), .B(n8933), .ZN(n7960) );
  NOR2_X1 U9093 ( .A1(n7970), .A2(n8932), .ZN(n7958) );
  XNOR2_X1 U9094 ( .A(n7960), .B(n7958), .ZN(n7956) );
  XOR2_X1 U9095 ( .A(n7957), .B(n7956), .Z(n7870) );
  INV_X1 U9096 ( .A(n7889), .ZN(n7867) );
  OR2_X1 U9097 ( .A1(n7884), .A2(n9320), .ZN(n7865) );
  NAND2_X1 U9098 ( .A1(n6554), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n7863) );
  NAND2_X1 U9099 ( .A1(n7858), .A2(n9671), .ZN(n7859) );
  AND2_X1 U9100 ( .A1(n7927), .A2(n7859), .ZN(n7969) );
  NAND2_X1 U9101 ( .A1(n6556), .A2(n7969), .ZN(n7862) );
  NAND2_X1 U9102 ( .A1(n6560), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n7861) );
  NAND2_X1 U9103 ( .A1(n6555), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n7860) );
  OR2_X1 U9104 ( .A1(n9003), .A2(n9318), .ZN(n7864) );
  NAND2_X1 U9105 ( .A1(n7865), .A2(n7864), .ZN(n7898) );
  AOI22_X1 U9106 ( .A1(n8920), .A2(n7898), .B1(P2_REG3_REG_16__SCAN_IN), .B2(
        P2_U3152), .ZN(n7866) );
  OAI21_X1 U9107 ( .B1(n9013), .B2(n7867), .A(n7866), .ZN(n7868) );
  AOI21_X1 U9108 ( .B1(n9437), .B2(n9017), .A(n7868), .ZN(n7869) );
  OAI21_X1 U9109 ( .B1(n7870), .B2(n9019), .A(n7869), .ZN(P2_U3228) );
  XNOR2_X1 U9110 ( .A(n7871), .B(n8354), .ZN(n10239) );
  AOI211_X1 U9111 ( .C1(n10237), .C2(n7872), .A(n10591), .B(n10151), .ZN(
        n10236) );
  INV_X1 U9112 ( .A(n10237), .ZN(n7873) );
  NOR2_X1 U9113 ( .A1(n7873), .A2(n10115), .ZN(n7876) );
  OAI22_X1 U9114 ( .A1(n10148), .A2(n7874), .B1(n9798), .B2(n10145), .ZN(n7875) );
  AOI211_X1 U9115 ( .C1(n10236), .C2(n10110), .A(n7876), .B(n7875), .ZN(n7881)
         );
  XNOR2_X1 U9116 ( .A(n7877), .B(n8354), .ZN(n7879) );
  OAI222_X1 U9117 ( .A1(n10103), .A2(n9795), .B1(n7879), .B2(n9997), .C1(
        n10101), .C2(n7878), .ZN(n10235) );
  NAND2_X1 U9118 ( .A1(n10235), .A2(n10148), .ZN(n7880) );
  OAI211_X1 U9119 ( .C1(n10239), .C2(n10137), .A(n7881), .B(n7880), .ZN(
        P1_U3275) );
  OR2_X1 U9120 ( .A1(n7882), .A2(n8778), .ZN(n7883) );
  OR2_X1 U9121 ( .A1(n9446), .A2(n9030), .ZN(n7909) );
  NAND2_X1 U9122 ( .A1(n7883), .A2(n7909), .ZN(n9287) );
  OR2_X1 U9123 ( .A1(n9441), .A2(n7884), .ZN(n8643) );
  NAND2_X1 U9124 ( .A1(n9441), .A2(n7884), .ZN(n8644) );
  NAND2_X1 U9125 ( .A1(n8643), .A2(n8644), .ZN(n8780) );
  NAND2_X1 U9126 ( .A1(n9287), .A2(n8780), .ZN(n7977) );
  OR2_X1 U9127 ( .A1(n9441), .A2(n9029), .ZN(n7885) );
  AND2_X1 U9128 ( .A1(n7977), .A2(n7885), .ZN(n7887) );
  NAND2_X1 U9129 ( .A1(n9437), .A2(n7970), .ZN(n8577) );
  NAND2_X1 U9130 ( .A1(n8576), .A2(n8577), .ZN(n8781) );
  AND2_X1 U9131 ( .A1(n8781), .A2(n7885), .ZN(n7903) );
  NAND2_X1 U9132 ( .A1(n7977), .A2(n7903), .ZN(n7886) );
  OAI21_X1 U9133 ( .B1(n7887), .B2(n8781), .A(n7886), .ZN(n9440) );
  INV_X1 U9134 ( .A(n9441), .ZN(n7984) );
  OR2_X1 U9135 ( .A1(n7936), .A2(n9437), .ZN(n9299) );
  INV_X1 U9136 ( .A(n9299), .ZN(n7888) );
  AOI211_X1 U9137 ( .C1(n9437), .C2(n7936), .A(n10637), .B(n7888), .ZN(n9436)
         );
  INV_X1 U9138 ( .A(n9437), .ZN(n7891) );
  AOI22_X1 U9139 ( .A1(n9223), .A2(P2_REG2_REG_16__SCAN_IN), .B1(n7889), .B2(
        n9350), .ZN(n7890) );
  OAI21_X1 U9140 ( .B1(n7891), .B2(n9272), .A(n7890), .ZN(n7901) );
  INV_X1 U9141 ( .A(n8638), .ZN(n7894) );
  OR2_X1 U9142 ( .A1(n7892), .A2(n7894), .ZN(n7985) );
  INV_X1 U9143 ( .A(n8643), .ZN(n7895) );
  OR2_X1 U9144 ( .A1(n7985), .A2(n7895), .ZN(n7897) );
  OR2_X1 U9145 ( .A1(n7894), .A2(n7893), .ZN(n7987) );
  OR2_X1 U9146 ( .A1(n7895), .A2(n7987), .ZN(n7896) );
  INV_X1 U9147 ( .A(n8781), .ZN(n8647) );
  XNOR2_X1 U9148 ( .A(n7941), .B(n8647), .ZN(n7899) );
  AOI21_X1 U9149 ( .B1(n7899), .B2(n9340), .A(n7898), .ZN(n9439) );
  NOR2_X1 U9150 ( .A1(n9439), .A2(n9354), .ZN(n7900) );
  AOI211_X1 U9151 ( .C1(n9436), .C2(n9187), .A(n7901), .B(n7900), .ZN(n7902)
         );
  OAI21_X1 U9152 ( .B1(n9440), .B2(n9285), .A(n7902), .ZN(P2_U3280) );
  INV_X1 U9153 ( .A(n7903), .ZN(n7904) );
  INV_X1 U9154 ( .A(n7970), .ZN(n9028) );
  NAND2_X1 U9155 ( .A1(n9437), .A2(n9028), .ZN(n7917) );
  INV_X1 U9156 ( .A(n9288), .ZN(n7908) );
  AOI22_X1 U9157 ( .A1(n7997), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n7996), .B2(
        n9076), .ZN(n7906) );
  NAND2_X1 U9158 ( .A1(n7909), .A2(n7916), .ZN(n7913) );
  NOR2_X1 U9159 ( .A1(n8777), .A2(n7913), .ZN(n7914) );
  AND2_X1 U9160 ( .A1(n7911), .A2(n7910), .ZN(n7912) );
  AOI21_X1 U9161 ( .B1(n7915), .B2(n7914), .A(n5244), .ZN(n7921) );
  INV_X1 U9162 ( .A(n7916), .ZN(n7919) );
  AND2_X1 U9163 ( .A1(n8780), .A2(n7917), .ZN(n9286) );
  AND2_X1 U9164 ( .A1(n9286), .A2(n9294), .ZN(n7918) );
  NAND2_X1 U9165 ( .A1(n7921), .A2(n7920), .ZN(n9293) );
  INV_X1 U9166 ( .A(n9003), .ZN(n9027) );
  OR2_X1 U9167 ( .A1(n9432), .A2(n9027), .ZN(n7922) );
  NAND2_X1 U9168 ( .A1(n9293), .A2(n7922), .ZN(n7933) );
  OR2_X1 U9169 ( .A1(n7923), .A2(n6564), .ZN(n7925) );
  AOI22_X1 U9170 ( .A1(n7997), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n7996), .B2(
        n9088), .ZN(n7924) );
  NAND2_X1 U9171 ( .A1(n7927), .A2(n7926), .ZN(n7928) );
  AND2_X1 U9172 ( .A1(n7945), .A2(n7928), .ZN(n9001) );
  NAND2_X1 U9173 ( .A1(n6556), .A2(n9001), .ZN(n7932) );
  NAND2_X1 U9174 ( .A1(n6560), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n7931) );
  NAND2_X1 U9175 ( .A1(n6555), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n7930) );
  NAND2_X1 U9176 ( .A1(n6554), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n7929) );
  NAND2_X1 U9177 ( .A1(n9426), .A2(n8837), .ZN(n8655) );
  NAND2_X1 U9178 ( .A1(n8656), .A2(n8655), .ZN(n8782) );
  NAND2_X1 U9179 ( .A1(n7933), .A2(n8782), .ZN(n8016) );
  OAI21_X1 U9180 ( .B1(n7933), .B2(n8782), .A(n8016), .ZN(n7934) );
  INV_X1 U9181 ( .A(n7934), .ZN(n9430) );
  OR2_X1 U9182 ( .A1(n9432), .A2(n9437), .ZN(n7935) );
  NOR2_X2 U9183 ( .A1(n7936), .A2(n7935), .ZN(n9298) );
  INV_X1 U9184 ( .A(n9298), .ZN(n7937) );
  INV_X1 U9185 ( .A(n9426), .ZN(n7939) );
  AOI21_X1 U9186 ( .B1(n9426), .B2(n7937), .A(n8027), .ZN(n9427) );
  AOI22_X1 U9187 ( .A1(n9223), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n9001), .B2(
        n9350), .ZN(n7938) );
  OAI21_X1 U9188 ( .B1(n7939), .B2(n9272), .A(n7938), .ZN(n7954) );
  INV_X1 U9189 ( .A(n8577), .ZN(n7940) );
  NAND2_X1 U9190 ( .A1(n9295), .A2(n9290), .ZN(n7943) );
  OR2_X1 U9191 ( .A1(n9432), .A2(n9003), .ZN(n7942) );
  NAND2_X1 U9192 ( .A1(n7943), .A2(n7942), .ZN(n7944) );
  INV_X1 U9193 ( .A(n8782), .ZN(n8653) );
  NAND2_X1 U9194 ( .A1(n7944), .A2(n8653), .ZN(n7994) );
  OAI211_X1 U9195 ( .C1(n7944), .C2(n8653), .A(n7994), .B(n9340), .ZN(n7952)
         );
  INV_X1 U9196 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n9532) );
  NAND2_X1 U9197 ( .A1(n7945), .A2(n9532), .ZN(n7946) );
  AND2_X1 U9198 ( .A1(n8004), .A2(n7946), .ZN(n8918) );
  NAND2_X1 U9199 ( .A1(n8918), .A2(n6556), .ZN(n7950) );
  NAND2_X1 U9200 ( .A1(n6554), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n7949) );
  NAND2_X1 U9201 ( .A1(n6555), .A2(P2_REG2_REG_19__SCAN_IN), .ZN(n7948) );
  NAND2_X1 U9202 ( .A1(n6560), .A2(P2_REG1_REG_19__SCAN_IN), .ZN(n7947) );
  NAND4_X1 U9203 ( .A1(n7950), .A2(n7949), .A3(n7948), .A4(n7947), .ZN(n9025)
         );
  AOI22_X1 U9204 ( .A1(n9027), .A2(n9345), .B1(n9346), .B2(n9025), .ZN(n7951)
         );
  AND2_X1 U9205 ( .A1(n7952), .A2(n7951), .ZN(n9429) );
  NOR2_X1 U9206 ( .A1(n9429), .A2(n9223), .ZN(n7953) );
  AOI211_X1 U9207 ( .C1(n9427), .C2(n9353), .A(n7954), .B(n7953), .ZN(n7955)
         );
  OAI21_X1 U9208 ( .B1(n9430), .B2(n9285), .A(n7955), .ZN(P2_U3278) );
  NAND2_X1 U9209 ( .A1(n7957), .A2(n7956), .ZN(n7962) );
  INV_X1 U9210 ( .A(n7958), .ZN(n7959) );
  NAND2_X1 U9211 ( .A1(n7960), .A2(n7959), .ZN(n7961) );
  NAND2_X1 U9212 ( .A1(n7962), .A2(n7961), .ZN(n8851) );
  XNOR2_X1 U9213 ( .A(n9432), .B(n8933), .ZN(n7963) );
  OR2_X1 U9214 ( .A1(n9003), .A2(n8932), .ZN(n7964) );
  AND2_X1 U9215 ( .A1(n7963), .A2(n7964), .ZN(n8996) );
  INV_X1 U9216 ( .A(n8996), .ZN(n7967) );
  INV_X1 U9217 ( .A(n7963), .ZN(n7966) );
  INV_X1 U9218 ( .A(n7964), .ZN(n7965) );
  NAND2_X1 U9219 ( .A1(n7966), .A2(n7965), .ZN(n8997) );
  NAND2_X1 U9220 ( .A1(n7967), .A2(n8997), .ZN(n7968) );
  XNOR2_X1 U9221 ( .A(n8851), .B(n7968), .ZN(n7976) );
  INV_X1 U9222 ( .A(n7969), .ZN(n9305) );
  OR2_X1 U9223 ( .A1(n7970), .A2(n9320), .ZN(n7972) );
  OR2_X1 U9224 ( .A1(n8837), .A2(n9318), .ZN(n7971) );
  NAND2_X1 U9225 ( .A1(n7972), .A2(n7971), .ZN(n9296) );
  AOI22_X1 U9226 ( .A1(n8920), .A2(n9296), .B1(P2_REG3_REG_17__SCAN_IN), .B2(
        P2_U3152), .ZN(n7973) );
  OAI21_X1 U9227 ( .B1(n9013), .B2(n9305), .A(n7973), .ZN(n7974) );
  AOI21_X1 U9228 ( .B1(n9432), .B2(n9017), .A(n7974), .ZN(n7975) );
  OAI21_X1 U9229 ( .B1(n7976), .B2(n9019), .A(n7975), .ZN(P2_U3230) );
  OAI21_X1 U9230 ( .B1(n9287), .B2(n8780), .A(n7977), .ZN(n7978) );
  INV_X1 U9231 ( .A(n7978), .ZN(n9445) );
  INV_X1 U9232 ( .A(n7979), .ZN(n7981) );
  INV_X1 U9233 ( .A(n7936), .ZN(n7980) );
  AOI21_X1 U9234 ( .B1(n9441), .B2(n7981), .A(n7980), .ZN(n9442) );
  AOI22_X1 U9235 ( .A1(n9223), .A2(P2_REG2_REG_15__SCAN_IN), .B1(n7982), .B2(
        n9350), .ZN(n7983) );
  OAI21_X1 U9236 ( .B1(n7984), .B2(n9272), .A(n7983), .ZN(n7992) );
  OR2_X1 U9237 ( .A1(n7986), .A2(n7985), .ZN(n7988) );
  AND2_X1 U9238 ( .A1(n7988), .A2(n7987), .ZN(n7989) );
  XNOR2_X1 U9239 ( .A(n7989), .B(n8780), .ZN(n7990) );
  AOI222_X1 U9240 ( .A1(n9340), .A2(n7990), .B1(n9028), .B2(n9346), .C1(n9030), 
        .C2(n9345), .ZN(n9444) );
  NOR2_X1 U9241 ( .A1(n9444), .A2(n9223), .ZN(n7991) );
  AOI211_X1 U9242 ( .C1(n9442), .C2(n9353), .A(n7992), .B(n7991), .ZN(n7993)
         );
  OAI21_X1 U9243 ( .B1(n9445), .B2(n9285), .A(n7993), .ZN(P2_U3281) );
  NAND2_X1 U9244 ( .A1(n7994), .A2(n8656), .ZN(n8032) );
  NAND2_X1 U9245 ( .A1(n7995), .A2(n8727), .ZN(n7999) );
  AOI22_X1 U9246 ( .A1(n7997), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n9103), .B2(
        n7996), .ZN(n7998) );
  INV_X1 U9247 ( .A(n9025), .ZN(n8980) );
  NAND2_X1 U9248 ( .A1(n9422), .A2(n8980), .ZN(n8575) );
  OR2_X1 U9249 ( .A1(n9422), .A2(n8980), .ZN(n8574) );
  NAND2_X1 U9250 ( .A1(n8000), .A2(n8727), .ZN(n8003) );
  OR2_X1 U9251 ( .A1(n6562), .A2(n8001), .ZN(n8002) );
  NAND2_X1 U9252 ( .A1(n8004), .A2(n9557), .ZN(n8005) );
  AND2_X1 U9253 ( .A1(n8009), .A2(n8005), .ZN(n8978) );
  NAND2_X1 U9254 ( .A1(n8978), .A2(n6556), .ZN(n8008) );
  AOI22_X1 U9255 ( .A1(n6554), .A2(P2_REG0_REG_20__SCAN_IN), .B1(n6555), .B2(
        P2_REG2_REG_20__SCAN_IN), .ZN(n8007) );
  NAND2_X1 U9256 ( .A1(n6560), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n8006) );
  NAND2_X1 U9257 ( .A1(n9416), .A2(n9118), .ZN(n8660) );
  NAND2_X1 U9258 ( .A1(n9275), .A2(n8660), .ZN(n8786) );
  XNOR2_X1 U9259 ( .A(n8801), .B(n8786), .ZN(n8014) );
  INV_X1 U9260 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n8013) );
  INV_X1 U9261 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n9540) );
  NAND2_X1 U9262 ( .A1(n8009), .A2(n9540), .ZN(n8010) );
  NAND2_X1 U9263 ( .A1(n8675), .A2(n8010), .ZN(n9269) );
  OR2_X1 U9264 ( .A1(n9269), .A2(n7303), .ZN(n8012) );
  AOI22_X1 U9265 ( .A1(n6554), .A2(P2_REG0_REG_21__SCAN_IN), .B1(n6555), .B2(
        P2_REG2_REG_21__SCAN_IN), .ZN(n8011) );
  OAI211_X1 U9266 ( .C1(n6535), .C2(n8013), .A(n8012), .B(n8011), .ZN(n9024)
         );
  AOI222_X1 U9267 ( .A1(n9340), .A2(n8014), .B1(n9024), .B2(n9346), .C1(n9025), 
        .C2(n9345), .ZN(n9419) );
  INV_X1 U9268 ( .A(n8837), .ZN(n9026) );
  NAND2_X1 U9269 ( .A1(n8016), .A2(n8015), .ZN(n8026) );
  NAND2_X1 U9270 ( .A1(n9422), .A2(n9025), .ZN(n8017) );
  AOI22_X1 U9271 ( .A1(n8026), .A2(n8017), .B1(n8030), .B2(n8980), .ZN(n8018)
         );
  OR2_X1 U9272 ( .A1(n8018), .A2(n8786), .ZN(n9415) );
  NAND2_X1 U9273 ( .A1(n8018), .A2(n8786), .ZN(n9414) );
  NAND3_X1 U9274 ( .A1(n9415), .A2(n9414), .A3(n9337), .ZN(n8023) );
  AOI21_X1 U9275 ( .B1(n9416), .B2(n8019), .A(n9266), .ZN(n9417) );
  INV_X1 U9276 ( .A(n9416), .ZN(n9117) );
  AOI22_X1 U9277 ( .A1(n9354), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n8978), .B2(
        n9350), .ZN(n8020) );
  OAI21_X1 U9278 ( .B1(n9117), .B2(n9272), .A(n8020), .ZN(n8021) );
  AOI21_X1 U9279 ( .B1(n9417), .B2(n9353), .A(n8021), .ZN(n8022) );
  OAI211_X1 U9280 ( .C1(n9354), .C2(n9419), .A(n8023), .B(n8022), .ZN(P2_U3276) );
  INV_X1 U9281 ( .A(n8550), .ZN(n8037) );
  OAI222_X1 U9282 ( .A1(n6276), .A2(n8037), .B1(n8025), .B2(P1_U3084), .C1(
        n8024), .C2(n8101), .ZN(P1_U3324) );
  XNOR2_X1 U9283 ( .A(n8026), .B(n8784), .ZN(n9425) );
  XNOR2_X1 U9284 ( .A(n8030), .B(n8027), .ZN(n8028) );
  NOR2_X1 U9285 ( .A1(n8028), .A2(n10637), .ZN(n9421) );
  AOI22_X1 U9286 ( .A1(n9223), .A2(P2_REG2_REG_19__SCAN_IN), .B1(n8918), .B2(
        n9350), .ZN(n8029) );
  OAI21_X1 U9287 ( .B1(n8030), .B2(n9272), .A(n8029), .ZN(n8035) );
  INV_X1 U9288 ( .A(n8784), .ZN(n8031) );
  XNOR2_X1 U9289 ( .A(n8032), .B(n8031), .ZN(n8033) );
  OAI22_X1 U9290 ( .A1(n9118), .A2(n9318), .B1(n8837), .B2(n9320), .ZN(n8919)
         );
  AOI21_X1 U9291 ( .B1(n8033), .B2(n9340), .A(n8919), .ZN(n9424) );
  NOR2_X1 U9292 ( .A1(n9424), .A2(n9354), .ZN(n8034) );
  AOI211_X1 U9293 ( .C1(n9421), .C2(n9187), .A(n8035), .B(n8034), .ZN(n8036)
         );
  OAI21_X1 U9294 ( .B1(n9425), .B2(n9285), .A(n8036), .ZN(P2_U3277) );
  OAI222_X1 U9295 ( .A1(P2_U3152), .A2(n8038), .B1(n8039), .B2(n8037), .C1(
        n8551), .C2(n9710), .ZN(P2_U3329) );
  INV_X1 U9296 ( .A(n8540), .ZN(n10326) );
  INV_X1 U9297 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n8541) );
  OAI222_X1 U9298 ( .A1(n8040), .A2(P2_U3152), .B1(n8039), .B2(n10326), .C1(
        n8541), .C2(n9710), .ZN(P2_U3328) );
  NAND2_X1 U9299 ( .A1(n8603), .A2(n8602), .ZN(n8766) );
  XOR2_X1 U9300 ( .A(n8766), .B(n8041), .Z(n10581) );
  XOR2_X1 U9301 ( .A(n8766), .B(n8042), .Z(n8043) );
  AOI222_X1 U9302 ( .A1(n9340), .A2(n8043), .B1(n9037), .B2(n9346), .C1(n9038), 
        .C2(n9345), .ZN(n10584) );
  MUX2_X1 U9303 ( .A(n6696), .B(n10584), .S(n9307), .Z(n8052) );
  NOR2_X1 U9304 ( .A1(n8044), .A2(n10582), .ZN(n8045) );
  OR2_X1 U9305 ( .A1(n8046), .A2(n8045), .ZN(n10583) );
  INV_X1 U9306 ( .A(n8047), .ZN(n8048) );
  OAI22_X1 U9307 ( .A1(n9139), .A2(n10583), .B1(n8048), .B2(n9304), .ZN(n8049)
         );
  AOI21_X1 U9308 ( .B1(n9336), .B2(n8050), .A(n8049), .ZN(n8051) );
  OAI211_X1 U9309 ( .C1(n10581), .C2(n9285), .A(n8052), .B(n8051), .ZN(
        P2_U3290) );
  XOR2_X1 U9310 ( .A(n8053), .B(n8054), .Z(n8060) );
  AOI22_X1 U9311 ( .A1(n9863), .A2(n8055), .B1(n9848), .B2(n6277), .ZN(n8059)
         );
  AOI22_X1 U9312 ( .A1(n8057), .A2(n9837), .B1(n8056), .B2(
        P1_REG3_REG_2__SCAN_IN), .ZN(n8058) );
  OAI211_X1 U9313 ( .C1(n8060), .C2(n9853), .A(n8059), .B(n8058), .ZN(P1_U3235) );
  INV_X1 U9314 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n8061) );
  MUX2_X1 U9315 ( .A(n8062), .B(n8061), .S(n10609), .Z(n8063) );
  OAI21_X1 U9316 ( .B1(n8326), .B2(n10311), .A(n8063), .ZN(P1_U3522) );
  NAND2_X1 U9317 ( .A1(n8065), .A2(n8064), .ZN(n8067) );
  XNOR2_X1 U9318 ( .A(n8067), .B(n8066), .ZN(n8076) );
  NAND2_X1 U9319 ( .A1(P1_U3084), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n9938) );
  INV_X1 U9320 ( .A(n9938), .ZN(n8070) );
  NOR2_X1 U9321 ( .A1(n9860), .A2(n8068), .ZN(n8069) );
  AOI211_X1 U9322 ( .C1(n9863), .C2(n9877), .A(n8070), .B(n8069), .ZN(n8071)
         );
  OAI21_X1 U9323 ( .B1(n9858), .B2(n8072), .A(n8071), .ZN(n8073) );
  AOI21_X1 U9324 ( .B1(n8074), .B2(n9851), .A(n8073), .ZN(n8075) );
  OAI21_X1 U9325 ( .B1(n8076), .B2(n9853), .A(n8075), .ZN(P1_U3215) );
  AOI211_X1 U9326 ( .C1(n8082), .C2(n8079), .A(n8078), .B(n8077), .ZN(n8080)
         );
  INV_X1 U9327 ( .A(n8080), .ZN(n8097) );
  NOR3_X1 U9328 ( .A1(n8083), .A2(n8082), .A3(n8081), .ZN(n8084) );
  AOI21_X1 U9329 ( .B1(n8085), .B2(n10443), .A(n8084), .ZN(n8087) );
  AOI21_X1 U9330 ( .B1(n8087), .B2(n9952), .A(n8086), .ZN(n8088) );
  AOI211_X1 U9331 ( .C1(n10457), .C2(P1_ADDR_REG_11__SCAN_IN), .A(n8089), .B(
        n8088), .ZN(n8096) );
  NOR2_X1 U9332 ( .A1(n8090), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n8093) );
  AOI21_X1 U9333 ( .B1(n8093), .B2(n8092), .A(n8091), .ZN(n8094) );
  NAND2_X1 U9334 ( .A1(n8094), .A2(n10443), .ZN(n8095) );
  OAI211_X1 U9335 ( .C1(n8097), .C2(n10451), .A(n8096), .B(n8095), .ZN(
        P1_U3252) );
  NOR2_X1 U9336 ( .A1(n10164), .A2(n10088), .ZN(n9959) );
  NOR2_X1 U9337 ( .A1(n8326), .A2(n10115), .ZN(n8098) );
  AOI211_X1 U9338 ( .C1(n10088), .C2(P1_REG2_REG_31__SCAN_IN), .A(n9959), .B(
        n8098), .ZN(n8099) );
  OAI21_X1 U9339 ( .B1(n8100), .B2(n10152), .A(n8099), .ZN(P1_U3261) );
  INV_X1 U9340 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n8102) );
  OAI222_X1 U9341 ( .A1(n6276), .A2(n8103), .B1(n4855), .B2(P1_U3084), .C1(
        n8102), .C2(n8101), .ZN(P1_U3326) );
  NAND2_X1 U9342 ( .A1(n10237), .A2(n8207), .ZN(n8108) );
  OR2_X1 U9343 ( .A1(n8110), .A2(n8208), .ZN(n8107) );
  NAND2_X1 U9344 ( .A1(n8108), .A2(n8107), .ZN(n8109) );
  XNOR2_X1 U9345 ( .A(n8109), .B(n8145), .ZN(n8113) );
  NOR2_X1 U9346 ( .A1(n8110), .A2(n6305), .ZN(n8111) );
  AOI21_X1 U9347 ( .B1(n10237), .B2(n6216), .A(n8111), .ZN(n8112) );
  NAND2_X1 U9348 ( .A1(n8113), .A2(n8112), .ZN(n8116) );
  OR2_X1 U9349 ( .A1(n8113), .A2(n8112), .ZN(n8114) );
  NAND2_X1 U9350 ( .A1(n8116), .A2(n8114), .ZN(n9793) );
  NAND2_X1 U9351 ( .A1(n10155), .A2(n8207), .ZN(n8118) );
  NAND2_X1 U9352 ( .A1(n10126), .A2(n6216), .ZN(n8117) );
  NAND2_X1 U9353 ( .A1(n8118), .A2(n8117), .ZN(n8119) );
  XNOR2_X1 U9354 ( .A(n8119), .B(n8195), .ZN(n8121) );
  NOR2_X1 U9355 ( .A1(n9795), .A2(n6305), .ZN(n8120) );
  AOI21_X1 U9356 ( .B1(n10155), .B2(n6216), .A(n8120), .ZN(n8122) );
  XNOR2_X1 U9357 ( .A(n8121), .B(n8122), .ZN(n9804) );
  INV_X1 U9358 ( .A(n8121), .ZN(n8123) );
  NAND2_X1 U9359 ( .A1(n8123), .A2(n8122), .ZN(n8124) );
  NAND2_X1 U9360 ( .A1(n10133), .A2(n8207), .ZN(n8126) );
  OR2_X1 U9361 ( .A1(n10102), .A2(n8208), .ZN(n8125) );
  NAND2_X1 U9362 ( .A1(n8126), .A2(n8125), .ZN(n8127) );
  XNOR2_X1 U9363 ( .A(n8127), .B(n8145), .ZN(n8130) );
  NOR2_X1 U9364 ( .A1(n10102), .A2(n6305), .ZN(n8129) );
  AOI21_X1 U9365 ( .B1(n10133), .B2(n6216), .A(n8129), .ZN(n9842) );
  NAND2_X1 U9366 ( .A1(n9840), .A2(n9842), .ZN(n8132) );
  NAND2_X1 U9367 ( .A1(n8131), .A2(n8130), .ZN(n9841) );
  NAND2_X1 U9368 ( .A1(n8132), .A2(n9841), .ZN(n9746) );
  NAND2_X1 U9369 ( .A1(n10109), .A2(n8207), .ZN(n8134) );
  NAND2_X1 U9370 ( .A1(n10125), .A2(n6216), .ZN(n8133) );
  NAND2_X1 U9371 ( .A1(n8134), .A2(n8133), .ZN(n8135) );
  XNOR2_X1 U9372 ( .A(n8135), .B(n8195), .ZN(n8138) );
  NAND2_X1 U9373 ( .A1(n10109), .A2(n6216), .ZN(n8137) );
  NAND2_X1 U9374 ( .A1(n10125), .A2(n8212), .ZN(n8136) );
  NAND2_X1 U9375 ( .A1(n8137), .A2(n8136), .ZN(n8139) );
  NAND2_X1 U9376 ( .A1(n9746), .A2(n9748), .ZN(n8142) );
  INV_X1 U9377 ( .A(n8138), .ZN(n8141) );
  INV_X1 U9378 ( .A(n8139), .ZN(n8140) );
  NAND2_X1 U9379 ( .A1(n8141), .A2(n8140), .ZN(n9747) );
  NAND2_X1 U9380 ( .A1(n10213), .A2(n8207), .ZN(n8144) );
  NAND2_X1 U9381 ( .A1(n10070), .A2(n6216), .ZN(n8143) );
  NAND2_X1 U9382 ( .A1(n8144), .A2(n8143), .ZN(n8146) );
  XNOR2_X1 U9383 ( .A(n8146), .B(n8145), .ZN(n9823) );
  NOR2_X1 U9384 ( .A1(n10104), .A2(n6305), .ZN(n8147) );
  AOI21_X1 U9385 ( .B1(n10213), .B2(n6216), .A(n8147), .ZN(n9822) );
  AND2_X1 U9386 ( .A1(n9823), .A2(n9822), .ZN(n8148) );
  INV_X1 U9387 ( .A(n9823), .ZN(n8150) );
  INV_X1 U9388 ( .A(n9822), .ZN(n8149) );
  NAND2_X1 U9389 ( .A1(n8150), .A2(n8149), .ZN(n8151) );
  NAND2_X1 U9390 ( .A1(n10075), .A2(n8207), .ZN(n8153) );
  OR2_X1 U9391 ( .A1(n8155), .A2(n8208), .ZN(n8152) );
  NAND2_X1 U9392 ( .A1(n8153), .A2(n8152), .ZN(n8154) );
  XNOR2_X1 U9393 ( .A(n8154), .B(n6585), .ZN(n8158) );
  NAND2_X1 U9394 ( .A1(n10075), .A2(n6216), .ZN(n8157) );
  OR2_X1 U9395 ( .A1(n8155), .A2(n6305), .ZN(n8156) );
  NAND2_X1 U9396 ( .A1(n8157), .A2(n8156), .ZN(n8159) );
  AND2_X1 U9397 ( .A1(n8158), .A2(n8159), .ZN(n9757) );
  INV_X1 U9398 ( .A(n8158), .ZN(n8161) );
  INV_X1 U9399 ( .A(n8159), .ZN(n8160) );
  NAND2_X1 U9400 ( .A1(n8161), .A2(n8160), .ZN(n9756) );
  NAND2_X1 U9401 ( .A1(n10205), .A2(n8207), .ZN(n8164) );
  NAND2_X1 U9402 ( .A1(n10071), .A2(n6216), .ZN(n8163) );
  NAND2_X1 U9403 ( .A1(n8164), .A2(n8163), .ZN(n8165) );
  XNOR2_X1 U9404 ( .A(n8165), .B(n6585), .ZN(n8168) );
  NAND2_X1 U9405 ( .A1(n10205), .A2(n6216), .ZN(n8167) );
  NAND2_X1 U9406 ( .A1(n10071), .A2(n8212), .ZN(n8166) );
  NAND2_X1 U9407 ( .A1(n8167), .A2(n8166), .ZN(n8169) );
  NAND2_X1 U9408 ( .A1(n8168), .A2(n8169), .ZN(n9831) );
  INV_X1 U9409 ( .A(n8168), .ZN(n8171) );
  INV_X1 U9410 ( .A(n8169), .ZN(n8170) );
  NAND2_X1 U9411 ( .A1(n8171), .A2(n8170), .ZN(n9833) );
  NAND2_X1 U9412 ( .A1(n10197), .A2(n8207), .ZN(n8173) );
  NAND2_X1 U9413 ( .A1(n10043), .A2(n6216), .ZN(n8172) );
  NAND2_X1 U9414 ( .A1(n8173), .A2(n8172), .ZN(n8174) );
  XNOR2_X1 U9415 ( .A(n8174), .B(n8195), .ZN(n8177) );
  AND2_X1 U9416 ( .A1(n10043), .A2(n8212), .ZN(n8175) );
  AOI21_X1 U9417 ( .B1(n10197), .B2(n6216), .A(n8175), .ZN(n9726) );
  INV_X1 U9418 ( .A(n8177), .ZN(n8178) );
  NAND2_X1 U9419 ( .A1(n8179), .A2(n8178), .ZN(n9729) );
  NAND2_X1 U9420 ( .A1(n10007), .A2(n8207), .ZN(n8181) );
  NAND2_X1 U9421 ( .A1(n10026), .A2(n6216), .ZN(n8180) );
  NAND2_X1 U9422 ( .A1(n8181), .A2(n8180), .ZN(n8182) );
  XNOR2_X1 U9423 ( .A(n8182), .B(n8195), .ZN(n8185) );
  AOI22_X1 U9424 ( .A1(n10007), .A2(n6216), .B1(n8212), .B2(n10026), .ZN(n8183) );
  XNOR2_X1 U9425 ( .A(n8185), .B(n8183), .ZN(n9813) );
  INV_X1 U9426 ( .A(n8183), .ZN(n8184) );
  NAND2_X1 U9427 ( .A1(n10189), .A2(n8207), .ZN(n8188) );
  NAND2_X1 U9428 ( .A1(n9872), .A2(n6216), .ZN(n8187) );
  NAND2_X1 U9429 ( .A1(n8188), .A2(n8187), .ZN(n8189) );
  XNOR2_X1 U9430 ( .A(n8189), .B(n8195), .ZN(n8193) );
  NAND2_X1 U9431 ( .A1(n10189), .A2(n6216), .ZN(n8191) );
  NAND2_X1 U9432 ( .A1(n9872), .A2(n8212), .ZN(n8190) );
  NAND2_X1 U9433 ( .A1(n8191), .A2(n8190), .ZN(n8192) );
  NOR2_X1 U9434 ( .A1(n8193), .A2(n8192), .ZN(n9779) );
  NAND2_X1 U9435 ( .A1(n8193), .A2(n8192), .ZN(n9780) );
  AND2_X1 U9436 ( .A1(n9988), .A2(n8212), .ZN(n8194) );
  AOI21_X1 U9437 ( .B1(n10182), .B2(n6216), .A(n8194), .ZN(n8198) );
  AOI22_X1 U9438 ( .A1(n10182), .A2(n8207), .B1(n6216), .B2(n9988), .ZN(n8196)
         );
  XNOR2_X1 U9439 ( .A(n8196), .B(n8195), .ZN(n8197) );
  XOR2_X1 U9440 ( .A(n8198), .B(n8197), .Z(n9857) );
  NAND2_X1 U9441 ( .A1(n9722), .A2(n8207), .ZN(n8203) );
  NAND2_X1 U9442 ( .A1(n9871), .A2(n6216), .ZN(n8202) );
  NAND2_X1 U9443 ( .A1(n8203), .A2(n8202), .ZN(n8204) );
  XNOR2_X1 U9444 ( .A(n8204), .B(n6585), .ZN(n9714) );
  NOR2_X1 U9445 ( .A1(n9971), .A2(n6305), .ZN(n8205) );
  AOI21_X1 U9446 ( .B1(n9722), .B2(n6216), .A(n8205), .ZN(n9713) );
  INV_X1 U9447 ( .A(n9713), .ZN(n8216) );
  NAND2_X1 U9448 ( .A1(n9716), .A2(n8206), .ZN(n8229) );
  NAND2_X1 U9449 ( .A1(n10173), .A2(n8207), .ZN(n8210) );
  OR2_X1 U9450 ( .A1(n9717), .A2(n8208), .ZN(n8209) );
  NAND2_X1 U9451 ( .A1(n8210), .A2(n8209), .ZN(n8211) );
  XNOR2_X1 U9452 ( .A(n8211), .B(n6585), .ZN(n8214) );
  AOI22_X1 U9453 ( .A1(n10173), .A2(n6216), .B1(n8212), .B2(n9870), .ZN(n8213)
         );
  XNOR2_X1 U9454 ( .A(n8214), .B(n8213), .ZN(n8223) );
  INV_X1 U9455 ( .A(n8223), .ZN(n8215) );
  NAND2_X1 U9456 ( .A1(n8215), .A2(n9855), .ZN(n8228) );
  NAND2_X1 U9457 ( .A1(n9714), .A2(n8216), .ZN(n8222) );
  INV_X1 U9458 ( .A(n8222), .ZN(n8217) );
  AND2_X1 U9459 ( .A1(n8223), .A2(n8218), .ZN(n8219) );
  NAND2_X1 U9460 ( .A1(n8229), .A2(n8219), .ZN(n8227) );
  AOI22_X1 U9461 ( .A1(n8522), .A2(n9783), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3084), .ZN(n8221) );
  NAND2_X1 U9462 ( .A1(n9869), .A2(n9863), .ZN(n8220) );
  OAI211_X1 U9463 ( .C1(n9971), .C2(n9860), .A(n8221), .B(n8220), .ZN(n8225)
         );
  NOR3_X1 U9464 ( .A1(n8223), .A2(n9853), .A3(n8222), .ZN(n8224) );
  AOI211_X1 U9465 ( .C1(n10173), .C2(n9837), .A(n8225), .B(n8224), .ZN(n8226)
         );
  OAI211_X1 U9466 ( .C1(n8229), .C2(n8228), .A(n8227), .B(n8226), .ZN(P1_U3218) );
  INV_X1 U9467 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n8729) );
  OAI222_X1 U9468 ( .A1(n6492), .A2(P2_U3152), .B1(n8039), .B2(n8231), .C1(
        n8729), .C2(n8230), .ZN(P2_U3330) );
  INV_X1 U9469 ( .A(n9868), .ZN(n8332) );
  NOR2_X1 U9470 ( .A1(n8333), .A2(n8332), .ZN(n8362) );
  NAND2_X1 U9471 ( .A1(n8362), .A2(n8233), .ZN(n8234) );
  INV_X1 U9472 ( .A(n8318), .ZN(n8364) );
  NAND2_X1 U9473 ( .A1(n8234), .A2(n8364), .ZN(n8366) );
  NAND2_X1 U9474 ( .A1(n9868), .A2(n9867), .ZN(n8235) );
  NAND2_X1 U9475 ( .A1(n8333), .A2(n8235), .ZN(n8438) );
  INV_X1 U9476 ( .A(n8438), .ZN(n8236) );
  NOR2_X1 U9477 ( .A1(n8366), .A2(n8236), .ZN(n8323) );
  INV_X1 U9478 ( .A(n8319), .ZN(n8300) );
  MUX2_X1 U9479 ( .A(n8430), .B(n8429), .S(n8300), .Z(n8310) );
  MUX2_X1 U9480 ( .A(n8432), .B(n8427), .S(n8319), .Z(n8308) );
  MUX2_X1 U9481 ( .A(n8423), .B(n8426), .S(n8300), .Z(n8306) );
  OR2_X1 U9482 ( .A1(n10007), .A2(n8237), .ZN(n8301) );
  NAND2_X1 U9483 ( .A1(n8301), .A2(n8238), .ZN(n8425) );
  NAND2_X1 U9484 ( .A1(n8425), .A2(n8300), .ZN(n8299) );
  MUX2_X1 U9485 ( .A(n10133), .B(n10142), .S(n8319), .Z(n8240) );
  NAND2_X1 U9486 ( .A1(n8240), .A2(n8239), .ZN(n8290) );
  XNOR2_X1 U9487 ( .A(n8367), .B(n8319), .ZN(n8245) );
  NAND2_X1 U9488 ( .A1(n8462), .A2(n8241), .ZN(n8368) );
  NAND2_X1 U9489 ( .A1(n8384), .A2(n8369), .ZN(n8242) );
  MUX2_X1 U9490 ( .A(n8368), .B(n8242), .S(n8319), .Z(n8243) );
  AOI21_X1 U9491 ( .B1(n8245), .B2(n8244), .A(n8243), .ZN(n8250) );
  MUX2_X1 U9492 ( .A(n8384), .B(n8462), .S(n8319), .Z(n8246) );
  NAND2_X1 U9493 ( .A1(n8344), .A2(n8246), .ZN(n8249) );
  MUX2_X1 U9494 ( .A(n8247), .B(n8400), .S(n8300), .Z(n8248) );
  OAI211_X1 U9495 ( .C1(n8250), .C2(n8249), .A(n4874), .B(n8248), .ZN(n8254)
         );
  INV_X1 U9496 ( .A(n8251), .ZN(n8402) );
  MUX2_X1 U9497 ( .A(n8379), .B(n8402), .S(n8319), .Z(n8252) );
  NAND3_X1 U9498 ( .A1(n8254), .A2(n8253), .A3(n8252), .ZN(n8257) );
  MUX2_X1 U9499 ( .A(n8380), .B(n8401), .S(n8300), .Z(n8255) );
  NAND3_X1 U9500 ( .A1(n8257), .A2(n8256), .A3(n8255), .ZN(n8261) );
  INV_X1 U9501 ( .A(n8403), .ZN(n8258) );
  MUX2_X1 U9502 ( .A(n8383), .B(n8258), .S(n8319), .Z(n8259) );
  NOR2_X1 U9503 ( .A1(n8348), .A2(n8259), .ZN(n8260) );
  NAND2_X1 U9504 ( .A1(n8261), .A2(n8260), .ZN(n8270) );
  NAND2_X1 U9505 ( .A1(n8270), .A2(n8377), .ZN(n8263) );
  AND2_X1 U9506 ( .A1(n8408), .A2(n8319), .ZN(n8262) );
  NAND2_X1 U9507 ( .A1(n8263), .A2(n8262), .ZN(n8274) );
  AND2_X1 U9508 ( .A1(n8271), .A2(n9874), .ZN(n8264) );
  NAND2_X1 U9509 ( .A1(n8274), .A2(n8264), .ZN(n8266) );
  NAND2_X1 U9510 ( .A1(n8266), .A2(n9874), .ZN(n8268) );
  INV_X1 U9511 ( .A(n8378), .ZN(n8265) );
  AOI22_X1 U9512 ( .A1(n8266), .A2(n8271), .B1(n8265), .B2(n8409), .ZN(n8267)
         );
  NAND2_X1 U9513 ( .A1(n8378), .A2(n8300), .ZN(n8269) );
  AOI21_X1 U9514 ( .B1(n8270), .B2(n8404), .A(n8269), .ZN(n8273) );
  NOR2_X1 U9515 ( .A1(n8408), .A2(n8319), .ZN(n8272) );
  NAND2_X1 U9516 ( .A1(n8271), .A2(n8275), .ZN(n8375) );
  OAI21_X1 U9517 ( .B1(n8273), .B2(n8272), .A(n8375), .ZN(n8278) );
  INV_X1 U9518 ( .A(n8274), .ZN(n8276) );
  NAND2_X1 U9519 ( .A1(n8276), .A2(n8275), .ZN(n8277) );
  NAND4_X1 U9520 ( .A1(n8279), .A2(n8352), .A3(n8278), .A4(n8277), .ZN(n8282)
         );
  INV_X1 U9521 ( .A(n8354), .ZN(n8281) );
  MUX2_X1 U9522 ( .A(n8414), .B(n8376), .S(n8300), .Z(n8280) );
  NAND3_X1 U9523 ( .A1(n8282), .A2(n8281), .A3(n8280), .ZN(n8284) );
  MUX2_X1 U9524 ( .A(n8371), .B(n8416), .S(n8300), .Z(n8283) );
  NAND2_X1 U9525 ( .A1(n8284), .A2(n8283), .ZN(n8285) );
  NAND2_X1 U9526 ( .A1(n8285), .A2(n10157), .ZN(n8288) );
  MUX2_X1 U9527 ( .A(n8286), .B(n8372), .S(n8319), .Z(n8287) );
  NAND3_X1 U9528 ( .A1(n8288), .A2(n10119), .A3(n8287), .ZN(n8289) );
  NAND3_X1 U9529 ( .A1(n10099), .A2(n8290), .A3(n8289), .ZN(n8292) );
  MUX2_X1 U9530 ( .A(n10063), .B(n8389), .S(n8300), .Z(n8291) );
  AND2_X1 U9531 ( .A1(n8292), .A2(n8291), .ZN(n8295) );
  OR2_X1 U9532 ( .A1(n10067), .A2(n10092), .ZN(n8334) );
  MUX2_X1 U9533 ( .A(n8293), .B(n8393), .S(n8319), .Z(n8294) );
  OAI211_X1 U9534 ( .C1(n8295), .C2(n8334), .A(n8294), .B(n10041), .ZN(n8297)
         );
  MUX2_X1 U9535 ( .A(n8392), .B(n8396), .S(n8319), .Z(n8296) );
  NAND3_X1 U9536 ( .A1(n8297), .A2(n10024), .A3(n8296), .ZN(n8298) );
  AOI21_X1 U9537 ( .B1(n8299), .B2(n8298), .A(n9983), .ZN(n8304) );
  INV_X1 U9538 ( .A(n9983), .ZN(n8422) );
  NAND2_X1 U9539 ( .A1(n10197), .A2(n10000), .ZN(n8424) );
  AOI21_X1 U9540 ( .B1(n8422), .B2(n8424), .A(n8300), .ZN(n8303) );
  INV_X1 U9541 ( .A(n9984), .ZN(n9987) );
  OR2_X1 U9542 ( .A1(n8301), .A2(n8300), .ZN(n8302) );
  OAI211_X1 U9543 ( .C1(n8304), .C2(n8303), .A(n9987), .B(n8302), .ZN(n8305)
         );
  NAND3_X1 U9544 ( .A1(n9970), .A2(n8306), .A3(n8305), .ZN(n8307) );
  NAND3_X1 U9545 ( .A1(n8473), .A2(n8308), .A3(n8307), .ZN(n8309) );
  INV_X1 U9546 ( .A(n8315), .ZN(n8311) );
  NAND3_X1 U9547 ( .A1(n8434), .A2(n8431), .A3(n8311), .ZN(n8312) );
  NAND2_X1 U9548 ( .A1(n8312), .A2(n8314), .ZN(n8317) );
  NAND2_X1 U9549 ( .A1(n8314), .A2(n8313), .ZN(n8479) );
  OAI21_X1 U9550 ( .B1(n8479), .B2(n8315), .A(n8434), .ZN(n8316) );
  MUX2_X1 U9551 ( .A(n8317), .B(n8316), .S(n8319), .Z(n8322) );
  NOR2_X1 U9552 ( .A1(n8318), .A2(n8438), .ZN(n8320) );
  MUX2_X1 U9553 ( .A(n8366), .B(n8320), .S(n8319), .Z(n8321) );
  AOI21_X1 U9554 ( .B1(n8453), .B2(n5945), .A(n8328), .ZN(n8324) );
  NAND2_X1 U9555 ( .A1(n8325), .A2(n10019), .ZN(n8327) );
  AND2_X1 U9556 ( .A1(n8333), .A2(n8332), .ZN(n8476) );
  INV_X1 U9557 ( .A(n10024), .ZN(n10016) );
  INV_X1 U9558 ( .A(n8334), .ZN(n8357) );
  INV_X1 U9559 ( .A(n8335), .ZN(n8337) );
  NAND4_X1 U9560 ( .A1(n8339), .A2(n8338), .A3(n8337), .A4(n8336), .ZN(n8340)
         );
  NOR4_X1 U9561 ( .A1(n5895), .A2(n8341), .A3(n8340), .A4(n6894), .ZN(n8343)
         );
  NAND4_X1 U9562 ( .A1(n4874), .A2(n8344), .A3(n8343), .A4(n8342), .ZN(n8345)
         );
  NOR4_X1 U9563 ( .A1(n8348), .A2(n8347), .A3(n8346), .A4(n8345), .ZN(n8350)
         );
  NAND4_X1 U9564 ( .A1(n8352), .A2(n8351), .A3(n8350), .A4(n8349), .ZN(n8353)
         );
  NOR4_X1 U9565 ( .A1(n5095), .A2(n8355), .A3(n8354), .A4(n8353), .ZN(n8356)
         );
  NAND4_X1 U9566 ( .A1(n8357), .A2(n10041), .A3(n10099), .A4(n8356), .ZN(n8358) );
  NOR4_X1 U9567 ( .A1(n9984), .A2(n10016), .A3(n9995), .A4(n8358), .ZN(n8359)
         );
  NAND4_X1 U9568 ( .A1(n8509), .A2(n8473), .A3(n9970), .A4(n8359), .ZN(n8360)
         );
  NOR4_X1 U9569 ( .A1(n8483), .A2(n8476), .A3(n8361), .A4(n8360), .ZN(n8365)
         );
  INV_X1 U9570 ( .A(n8362), .ZN(n8363) );
  AND2_X1 U9571 ( .A1(n8364), .A2(n8363), .ZN(n8480) );
  AOI21_X1 U9572 ( .B1(n8365), .B2(n8480), .A(n8453), .ZN(n8445) );
  INV_X1 U9573 ( .A(n8366), .ZN(n8442) );
  INV_X1 U9574 ( .A(n8367), .ZN(n8370) );
  AOI21_X1 U9575 ( .B1(n8370), .B2(n8369), .A(n8368), .ZN(n8420) );
  NAND3_X1 U9576 ( .A1(n8393), .A2(n8392), .A3(n10063), .ZN(n8419) );
  AND2_X1 U9577 ( .A1(n8372), .A2(n8371), .ZN(n8373) );
  NAND2_X1 U9578 ( .A1(n8374), .A2(n8373), .ZN(n8417) );
  NAND2_X1 U9579 ( .A1(n8376), .A2(n8375), .ZN(n8399) );
  NAND2_X1 U9580 ( .A1(n8378), .A2(n8377), .ZN(n8411) );
  NAND2_X1 U9581 ( .A1(n8380), .A2(n8379), .ZN(n8381) );
  AND2_X1 U9582 ( .A1(n8381), .A2(n8401), .ZN(n8382) );
  OR2_X1 U9583 ( .A1(n8383), .A2(n8382), .ZN(n8406) );
  OR3_X1 U9584 ( .A1(n8406), .A2(n8385), .A3(n5107), .ZN(n8386) );
  OR3_X1 U9585 ( .A1(n8399), .A2(n8411), .A3(n8386), .ZN(n8387) );
  OR3_X1 U9586 ( .A1(n8419), .A2(n8417), .A3(n8387), .ZN(n8469) );
  INV_X1 U9587 ( .A(n8388), .ZN(n8390) );
  AND2_X1 U9588 ( .A1(n8390), .A2(n8389), .ZN(n8397) );
  INV_X1 U9589 ( .A(n8391), .ZN(n8394) );
  NAND3_X1 U9590 ( .A1(n8394), .A2(n8393), .A3(n8392), .ZN(n8395) );
  OAI211_X1 U9591 ( .C1(n8419), .C2(n8397), .A(n8396), .B(n8395), .ZN(n8398)
         );
  NOR2_X1 U9592 ( .A1(n8425), .A2(n8398), .ZN(n8450) );
  INV_X1 U9593 ( .A(n8399), .ZN(n8413) );
  AND3_X1 U9594 ( .A1(n8402), .A2(n8401), .A3(n8400), .ZN(n8405) );
  OAI211_X1 U9595 ( .C1(n8406), .C2(n8405), .A(n8404), .B(n8403), .ZN(n8407)
         );
  INV_X1 U9596 ( .A(n8407), .ZN(n8410) );
  OAI211_X1 U9597 ( .C1(n8411), .C2(n8410), .A(n8409), .B(n8408), .ZN(n8412)
         );
  NAND2_X1 U9598 ( .A1(n8413), .A2(n8412), .ZN(n8415) );
  AND3_X1 U9599 ( .A1(n8416), .A2(n8415), .A3(n8414), .ZN(n8418) );
  OR3_X1 U9600 ( .A1(n8419), .A2(n8418), .A3(n8417), .ZN(n8467) );
  OAI211_X1 U9601 ( .C1(n8420), .C2(n8469), .A(n8450), .B(n8467), .ZN(n8421)
         );
  INV_X1 U9602 ( .A(n8421), .ZN(n8428) );
  OAI211_X1 U9603 ( .C1(n8425), .C2(n8424), .A(n8423), .B(n8422), .ZN(n8474)
         );
  AND2_X1 U9604 ( .A1(n8427), .A2(n8426), .ZN(n8472) );
  OAI211_X1 U9605 ( .C1(n8428), .C2(n8474), .A(n8429), .B(n8472), .ZN(n8439)
         );
  INV_X1 U9606 ( .A(n8479), .ZN(n8437) );
  INV_X1 U9607 ( .A(n8429), .ZN(n8433) );
  OAI211_X1 U9608 ( .C1(n8433), .C2(n8432), .A(n8431), .B(n8430), .ZN(n8436)
         );
  INV_X1 U9609 ( .A(n8434), .ZN(n8435) );
  OAI211_X1 U9610 ( .C1(n8479), .C2(n8439), .A(n8449), .B(n8438), .ZN(n8441)
         );
  AOI211_X1 U9611 ( .C1(n8442), .C2(n8441), .A(n8440), .B(n8483), .ZN(n8443)
         );
  NOR2_X1 U9612 ( .A1(n8445), .A2(n8443), .ZN(n8444) );
  MUX2_X1 U9613 ( .A(n8445), .B(n8444), .S(n9951), .Z(n8446) );
  INV_X1 U9614 ( .A(n8449), .ZN(n8482) );
  INV_X1 U9615 ( .A(n8450), .ZN(n8471) );
  INV_X1 U9616 ( .A(n8451), .ZN(n8454) );
  NAND2_X1 U9617 ( .A1(n6277), .A2(n6347), .ZN(n8452) );
  NAND3_X1 U9618 ( .A1(n8454), .A2(n8453), .A3(n8452), .ZN(n8455) );
  NAND2_X1 U9619 ( .A1(n8456), .A2(n8455), .ZN(n8459) );
  OAI211_X1 U9620 ( .C1(n8460), .C2(n8459), .A(n8458), .B(n8457), .ZN(n8466)
         );
  AND2_X1 U9621 ( .A1(n8461), .A2(n5245), .ZN(n8465) );
  NAND2_X1 U9622 ( .A1(n8463), .A2(n8462), .ZN(n8464) );
  AOI21_X1 U9623 ( .B1(n8466), .B2(n8465), .A(n8464), .ZN(n8468) );
  OAI21_X1 U9624 ( .B1(n8469), .B2(n8468), .A(n8467), .ZN(n8470) );
  NOR2_X1 U9625 ( .A1(n8471), .A2(n8470), .ZN(n8475) );
  OAI211_X1 U9626 ( .C1(n8475), .C2(n8474), .A(n8473), .B(n8472), .ZN(n8478)
         );
  INV_X1 U9627 ( .A(n8476), .ZN(n8477) );
  OAI21_X1 U9628 ( .B1(n8479), .B2(n8478), .A(n8477), .ZN(n8481) );
  OAI21_X1 U9629 ( .B1(n8482), .B2(n8481), .A(n8480), .ZN(n8485) );
  INV_X1 U9630 ( .A(n8483), .ZN(n8484) );
  NOR2_X1 U9631 ( .A1(n8490), .A2(n9951), .ZN(n8487) );
  NAND2_X1 U9632 ( .A1(n8487), .A2(n8486), .ZN(n8488) );
  INV_X1 U9633 ( .A(n8490), .ZN(n8492) );
  OAI21_X1 U9634 ( .B1(n8492), .B2(n8491), .A(n8493), .ZN(n8499) );
  INV_X1 U9635 ( .A(n8493), .ZN(n8496) );
  NAND3_X1 U9636 ( .A1(n8494), .A2(n10407), .A3(n10143), .ZN(n8495) );
  OAI211_X1 U9637 ( .C1(n8497), .C2(n8496), .A(n8495), .B(P1_B_REG_SCAN_IN), 
        .ZN(n8498) );
  OAI21_X1 U9638 ( .B1(n8500), .B2(n8499), .A(n8498), .ZN(P1_U3240) );
  NAND2_X1 U9639 ( .A1(n8501), .A2(n10097), .ZN(n8504) );
  INV_X1 U9640 ( .A(n8502), .ZN(n9718) );
  AOI22_X1 U9641 ( .A1(n9718), .A2(n10111), .B1(P1_REG2_REG_27__SCAN_IN), .B2(
        n10088), .ZN(n8503) );
  OAI211_X1 U9642 ( .C1(n10181), .C2(n10115), .A(n8504), .B(n8503), .ZN(n8505)
         );
  AOI21_X1 U9643 ( .B1(n8506), .B2(n10148), .A(n8505), .ZN(n8507) );
  OAI21_X1 U9644 ( .B1(n8508), .B2(n10137), .A(n8507), .ZN(P1_U3264) );
  NAND2_X1 U9645 ( .A1(n8510), .A2(n8509), .ZN(n8511) );
  NAND2_X1 U9646 ( .A1(n8515), .A2(n10140), .ZN(n8517) );
  AOI22_X1 U9647 ( .A1(n9869), .A2(n10141), .B1(n9871), .B2(n10143), .ZN(n8516) );
  NAND2_X1 U9648 ( .A1(n8517), .A2(n8516), .ZN(n8518) );
  INV_X1 U9649 ( .A(n8520), .ZN(n8521) );
  AOI21_X1 U9650 ( .B1(n10173), .B2(n5021), .A(n8521), .ZN(n10174) );
  AOI22_X1 U9651 ( .A1(n8522), .A2(n10111), .B1(P1_REG2_REG_28__SCAN_IN), .B2(
        n10088), .ZN(n8523) );
  OAI21_X1 U9652 ( .B1(n8524), .B2(n10115), .A(n8523), .ZN(n8528) );
  NOR2_X1 U9653 ( .A1(n10177), .A2(n8526), .ZN(n8527) );
  OAI21_X1 U9654 ( .B1(n10176), .B2(n10088), .A(n8529), .ZN(P1_U3263) );
  AOI22_X1 U9655 ( .A1(n10529), .A2(n9017), .B1(n9005), .B2(n9040), .ZN(n8534)
         );
  INV_X1 U9656 ( .A(n8530), .ZN(n8833) );
  XNOR2_X1 U9657 ( .A(n8531), .B(n4875), .ZN(n8532) );
  AOI22_X1 U9658 ( .A1(n8833), .A2(P2_REG3_REG_2__SCAN_IN), .B1(n8941), .B2(
        n8532), .ZN(n8533) );
  OAI211_X1 U9659 ( .C1(n9321), .C2(n9014), .A(n8534), .B(n8533), .ZN(P2_U3239) );
  NAND2_X1 U9660 ( .A1(n9704), .A2(n8727), .ZN(n8536) );
  INV_X1 U9661 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n9711) );
  OR2_X1 U9662 ( .A1(n6562), .A2(n9711), .ZN(n8535) );
  NAND2_X1 U9663 ( .A1(n6560), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n8539) );
  NAND2_X1 U9664 ( .A1(n6555), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n8538) );
  NAND2_X1 U9665 ( .A1(n6554), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n8537) );
  OR2_X1 U9666 ( .A1(n9106), .A2(n8812), .ZN(n8547) );
  NAND2_X1 U9667 ( .A1(n8540), .A2(n8727), .ZN(n8543) );
  OR2_X1 U9668 ( .A1(n6562), .A2(n8541), .ZN(n8542) );
  INV_X1 U9669 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n8546) );
  NAND2_X1 U9670 ( .A1(n6560), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n8545) );
  NAND2_X1 U9671 ( .A1(n6555), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n8544) );
  OAI211_X1 U9672 ( .C1(n8737), .C2(n8546), .A(n8545), .B(n8544), .ZN(n9131)
         );
  INV_X1 U9673 ( .A(n9131), .ZN(n8548) );
  NAND2_X1 U9674 ( .A1(n9113), .A2(n8548), .ZN(n8748) );
  NAND2_X1 U9675 ( .A1(n8547), .A2(n8748), .ZN(n8818) );
  OR2_X1 U9676 ( .A1(n9113), .A2(n8548), .ZN(n8814) );
  NAND2_X1 U9677 ( .A1(n9106), .A2(n8812), .ZN(n8817) );
  NAND2_X1 U9678 ( .A1(n8814), .A2(n8817), .ZN(n8549) );
  MUX2_X1 U9679 ( .A(n8818), .B(n8549), .S(n8749), .Z(n8753) );
  NAND2_X1 U9680 ( .A1(n8550), .A2(n8727), .ZN(n8553) );
  OR2_X1 U9681 ( .A1(n6562), .A2(n8551), .ZN(n8552) );
  INV_X1 U9682 ( .A(n8719), .ZN(n8554) );
  NAND2_X1 U9683 ( .A1(n8554), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n8733) );
  INV_X1 U9684 ( .A(n8733), .ZN(n8555) );
  NAND2_X1 U9685 ( .A1(n8555), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n9140) );
  OR2_X1 U9686 ( .A1(n9140), .A2(n7303), .ZN(n8561) );
  INV_X1 U9687 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n8558) );
  NAND2_X1 U9688 ( .A1(n6560), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n8557) );
  NAND2_X1 U9689 ( .A1(n6555), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n8556) );
  OAI211_X1 U9690 ( .C1(n8737), .C2(n8558), .A(n8557), .B(n8556), .ZN(n8559)
         );
  INV_X1 U9691 ( .A(n8559), .ZN(n8560) );
  NAND2_X1 U9692 ( .A1(n9136), .A2(n9155), .ZN(n8811) );
  NAND2_X1 U9693 ( .A1(n8562), .A2(n8727), .ZN(n8564) );
  OR2_X1 U9694 ( .A1(n6562), .A2(n7205), .ZN(n8563) );
  INV_X1 U9695 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n8565) );
  INV_X1 U9696 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n9674) );
  OAI21_X1 U9697 ( .B1(n8685), .B2(n8565), .A(n9674), .ZN(n8567) );
  NAND2_X1 U9698 ( .A1(n8567), .A2(n8566), .ZN(n9214) );
  OR2_X1 U9699 ( .A1(n9214), .A2(n7303), .ZN(n8573) );
  INV_X1 U9700 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n8570) );
  NAND2_X1 U9701 ( .A1(n6560), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n8569) );
  NAND2_X1 U9702 ( .A1(n6555), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n8568) );
  OAI211_X1 U9703 ( .C1(n8737), .C2(n8570), .A(n8569), .B(n8568), .ZN(n8571)
         );
  INV_X1 U9704 ( .A(n8571), .ZN(n8572) );
  INV_X1 U9705 ( .A(n8804), .ZN(n8704) );
  INV_X1 U9706 ( .A(n8786), .ZN(n9274) );
  MUX2_X1 U9707 ( .A(n8575), .B(n8574), .S(n8749), .Z(n8659) );
  INV_X1 U9708 ( .A(n8749), .ZN(n8746) );
  MUX2_X1 U9709 ( .A(n8577), .B(n8576), .S(n8746), .Z(n8649) );
  AND2_X1 U9710 ( .A1(n9338), .A2(n8578), .ZN(n8763) );
  INV_X1 U9711 ( .A(n8763), .ZN(n8580) );
  AND2_X1 U9712 ( .A1(n8580), .A2(n8579), .ZN(n8582) );
  OAI21_X1 U9713 ( .B1(n8819), .B2(n8580), .A(n9317), .ZN(n8581) );
  MUX2_X1 U9714 ( .A(n8582), .B(n8581), .S(n8749), .Z(n8583) );
  NAND2_X1 U9715 ( .A1(n8583), .A2(n9316), .ZN(n8587) );
  MUX2_X1 U9716 ( .A(n8585), .B(n8584), .S(n8749), .Z(n8586) );
  NAND3_X1 U9717 ( .A1(n8587), .A2(n8761), .A3(n8586), .ZN(n8592) );
  MUX2_X1 U9718 ( .A(n8589), .B(n8588), .S(n8749), .Z(n8590) );
  NAND3_X1 U9719 ( .A1(n8592), .A2(n8591), .A3(n8590), .ZN(n8597) );
  INV_X1 U9720 ( .A(n8593), .ZN(n8594) );
  NAND3_X1 U9721 ( .A1(n8597), .A2(n8764), .A3(n8596), .ZN(n8601) );
  MUX2_X1 U9722 ( .A(n8599), .B(n8598), .S(n8749), .Z(n8600) );
  AOI21_X1 U9723 ( .B1(n8601), .B2(n8600), .A(n8766), .ZN(n8606) );
  MUX2_X1 U9724 ( .A(n8603), .B(n8602), .S(n8749), .Z(n8604) );
  NAND2_X1 U9725 ( .A1(n8604), .A2(n8768), .ZN(n8605) );
  AND2_X1 U9726 ( .A1(n8612), .A2(n8617), .ZN(n8607) );
  MUX2_X1 U9727 ( .A(n8608), .B(n8607), .S(n8749), .Z(n8609) );
  AND2_X1 U9728 ( .A1(n8609), .A2(n8614), .ZN(n8624) );
  NAND4_X1 U9729 ( .A1(n8619), .A2(n8769), .A3(n8624), .A4(n8610), .ZN(n8613)
         );
  NAND2_X1 U9730 ( .A1(n8617), .A2(n8616), .ZN(n8623) );
  NAND3_X1 U9731 ( .A1(n8619), .A2(n8769), .A3(n8618), .ZN(n8621) );
  NAND2_X1 U9732 ( .A1(n8621), .A2(n8620), .ZN(n8622) );
  NAND2_X1 U9733 ( .A1(n8629), .A2(n8628), .ZN(n8631) );
  MUX2_X1 U9734 ( .A(n8631), .B(n8630), .S(n8746), .Z(n8632) );
  NAND3_X1 U9735 ( .A1(n8633), .A2(n8777), .A3(n8632), .ZN(n8637) );
  MUX2_X1 U9736 ( .A(n8635), .B(n8634), .S(n8749), .Z(n8636) );
  NAND3_X1 U9737 ( .A1(n8637), .A2(n8778), .A3(n8636), .ZN(n8642) );
  INV_X1 U9738 ( .A(n8780), .ZN(n8641) );
  MUX2_X1 U9739 ( .A(n8639), .B(n8638), .S(n8746), .Z(n8640) );
  NAND3_X1 U9740 ( .A1(n8642), .A2(n8641), .A3(n8640), .ZN(n8646) );
  MUX2_X1 U9741 ( .A(n8644), .B(n8643), .S(n8749), .Z(n8645) );
  NAND3_X1 U9742 ( .A1(n8647), .A2(n8646), .A3(n8645), .ZN(n8648) );
  NAND3_X1 U9743 ( .A1(n9290), .A2(n8649), .A3(n8648), .ZN(n8654) );
  OR2_X1 U9744 ( .A1(n9003), .A2(n8746), .ZN(n8651) );
  NAND2_X1 U9745 ( .A1(n9003), .A2(n8746), .ZN(n8650) );
  MUX2_X1 U9746 ( .A(n8651), .B(n8650), .S(n9432), .Z(n8652) );
  NAND3_X1 U9747 ( .A1(n8654), .A2(n8653), .A3(n8652), .ZN(n8658) );
  MUX2_X1 U9748 ( .A(n8656), .B(n8655), .S(n8749), .Z(n8657) );
  MUX2_X1 U9749 ( .A(n8660), .B(n9275), .S(n8746), .Z(n8661) );
  OR2_X1 U9750 ( .A1(n8662), .A2(n6564), .ZN(n8665) );
  OR2_X1 U9751 ( .A1(n6562), .A2(n8663), .ZN(n8664) );
  NAND2_X1 U9752 ( .A1(n9409), .A2(n9024), .ZN(n8760) );
  INV_X1 U9753 ( .A(n8760), .ZN(n8666) );
  MUX2_X1 U9754 ( .A(n9024), .B(n9409), .S(n8746), .Z(n8667) );
  INV_X1 U9755 ( .A(n8667), .ZN(n8670) );
  OAI21_X1 U9756 ( .B1(n5238), .B2(n8670), .A(n8669), .ZN(n8680) );
  NAND2_X1 U9757 ( .A1(n8671), .A2(n8727), .ZN(n8674) );
  OR2_X1 U9758 ( .A1(n6562), .A2(n8672), .ZN(n8673) );
  NAND2_X1 U9759 ( .A1(n8675), .A2(n9575), .ZN(n8676) );
  AND2_X1 U9760 ( .A1(n8685), .A2(n8676), .ZN(n9250) );
  NAND2_X1 U9761 ( .A1(n9250), .A2(n6556), .ZN(n8679) );
  AOI22_X1 U9762 ( .A1(n6554), .A2(P2_REG0_REG_22__SCAN_IN), .B1(n6555), .B2(
        P2_REG2_REG_22__SCAN_IN), .ZN(n8678) );
  NAND2_X1 U9763 ( .A1(n6560), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n8677) );
  NAND2_X1 U9764 ( .A1(n9404), .A2(n8957), .ZN(n8691) );
  NAND2_X1 U9765 ( .A1(n8680), .A2(n9120), .ZN(n8690) );
  NAND2_X1 U9766 ( .A1(n8681), .A2(n8727), .ZN(n8684) );
  OR2_X1 U9767 ( .A1(n6562), .A2(n8682), .ZN(n8683) );
  XNOR2_X1 U9768 ( .A(n8685), .B(P2_REG3_REG_23__SCAN_IN), .ZN(n9242) );
  INV_X1 U9769 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n8688) );
  NAND2_X1 U9770 ( .A1(n6560), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n8687) );
  NAND2_X1 U9771 ( .A1(n6555), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n8686) );
  OAI211_X1 U9772 ( .C1(n8737), .C2(n8688), .A(n8687), .B(n8686), .ZN(n8689)
         );
  AOI21_X1 U9773 ( .B1(n9242), .B2(n6556), .A(n8689), .ZN(n9257) );
  NAND2_X1 U9774 ( .A1(n8872), .A2(n9257), .ZN(n8802) );
  NAND2_X1 U9775 ( .A1(n8690), .A2(n8802), .ZN(n8696) );
  INV_X1 U9776 ( .A(n8691), .ZN(n8693) );
  OR2_X1 U9777 ( .A1(n8872), .A2(n9257), .ZN(n8759) );
  NAND2_X1 U9778 ( .A1(n8759), .A2(n9230), .ZN(n8692) );
  MUX2_X1 U9779 ( .A(n8693), .B(n8692), .S(n8749), .Z(n8695) );
  INV_X1 U9780 ( .A(n8697), .ZN(n8703) );
  INV_X1 U9781 ( .A(n9394), .ZN(n9217) );
  NAND2_X1 U9782 ( .A1(n8698), .A2(n8727), .ZN(n8701) );
  OR2_X1 U9783 ( .A1(n6562), .A2(n8699), .ZN(n8700) );
  OAI21_X1 U9784 ( .B1(n8704), .B2(n8703), .A(n8702), .ZN(n8708) );
  INV_X1 U9785 ( .A(n8705), .ZN(n8706) );
  NAND3_X1 U9786 ( .A1(n8706), .A2(n9206), .A3(n8746), .ZN(n8707) );
  NAND2_X1 U9787 ( .A1(n8709), .A2(n8727), .ZN(n8712) );
  OR2_X1 U9788 ( .A1(n6562), .A2(n8710), .ZN(n8711) );
  NAND2_X1 U9789 ( .A1(n9386), .A2(n9172), .ZN(n8806) );
  NAND2_X1 U9790 ( .A1(n9391), .A2(n9219), .ZN(n8757) );
  OR2_X1 U9791 ( .A1(n9386), .A2(n9172), .ZN(n8756) );
  INV_X1 U9792 ( .A(n8756), .ZN(n8713) );
  AND2_X1 U9793 ( .A1(n8756), .A2(n9181), .ZN(n8805) );
  INV_X1 U9794 ( .A(n8806), .ZN(n8714) );
  NAND2_X1 U9795 ( .A1(n8715), .A2(n8727), .ZN(n8718) );
  OR2_X1 U9796 ( .A1(n6562), .A2(n8716), .ZN(n8717) );
  INV_X1 U9797 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n9651) );
  NAND2_X1 U9798 ( .A1(n8719), .A2(n9651), .ZN(n8720) );
  NAND2_X1 U9799 ( .A1(n8733), .A2(n8720), .ZN(n9166) );
  INV_X1 U9800 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n8723) );
  NAND2_X1 U9801 ( .A1(n6560), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n8722) );
  NAND2_X1 U9802 ( .A1(n6555), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n8721) );
  OAI211_X1 U9803 ( .C1(n8737), .C2(n8723), .A(n8722), .B(n8721), .ZN(n8724)
         );
  INV_X1 U9804 ( .A(n8724), .ZN(n8725) );
  NAND2_X1 U9805 ( .A1(n9379), .A2(n9185), .ZN(n8742) );
  NAND2_X1 U9806 ( .A1(n8728), .A2(n8727), .ZN(n8731) );
  OR2_X1 U9807 ( .A1(n6562), .A2(n8729), .ZN(n8730) );
  INV_X1 U9808 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n8732) );
  NAND2_X1 U9809 ( .A1(n8733), .A2(n8732), .ZN(n8734) );
  NAND2_X1 U9810 ( .A1(n9140), .A2(n8734), .ZN(n8948) );
  OR2_X1 U9811 ( .A1(n8948), .A2(n7303), .ZN(n8741) );
  INV_X1 U9812 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n8738) );
  NAND2_X1 U9813 ( .A1(n6560), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n8736) );
  NAND2_X1 U9814 ( .A1(n6555), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n8735) );
  OAI211_X1 U9815 ( .C1(n8738), .C2(n8737), .A(n8736), .B(n8735), .ZN(n8739)
         );
  INV_X1 U9816 ( .A(n8739), .ZN(n8740) );
  MUX2_X1 U9817 ( .A(n8808), .B(n8742), .S(n8749), .Z(n8743) );
  OR3_X1 U9818 ( .A1(n9374), .A2(n9173), .A3(n8746), .ZN(n8745) );
  NAND3_X1 U9819 ( .A1(n9374), .A2(n9173), .A3(n8746), .ZN(n8744) );
  MUX2_X1 U9820 ( .A(n8811), .B(n8810), .S(n8746), .Z(n8747) );
  INV_X1 U9821 ( .A(n8812), .ZN(n9109) );
  MUX2_X1 U9822 ( .A(n9106), .B(n9109), .S(n8749), .Z(n8750) );
  OAI21_X1 U9823 ( .B1(n9360), .B2(n8812), .A(n8750), .ZN(n8751) );
  INV_X1 U9824 ( .A(n8818), .ZN(n8791) );
  NAND2_X1 U9825 ( .A1(n9181), .A2(n8757), .ZN(n9124) );
  NAND2_X1 U9826 ( .A1(n8804), .A2(n8758), .ZN(n9218) );
  INV_X1 U9827 ( .A(n9218), .ZN(n8803) );
  INV_X1 U9828 ( .A(n9236), .ZN(n8787) );
  NAND2_X1 U9829 ( .A1(n9119), .A2(n8760), .ZN(n9278) );
  NAND4_X1 U9830 ( .A1(n8764), .A2(n8763), .A3(n8762), .A4(n8761), .ZN(n8765)
         );
  NAND2_X1 U9831 ( .A1(n9317), .A2(n9316), .ZN(n9315) );
  NOR4_X1 U9832 ( .A1(n8767), .A2(n8766), .A3(n8765), .A4(n9315), .ZN(n8771)
         );
  NAND4_X1 U9833 ( .A1(n8771), .A2(n8770), .A3(n8769), .A4(n8768), .ZN(n8774)
         );
  NOR3_X1 U9834 ( .A1(n8774), .A2(n8773), .A3(n8772), .ZN(n8775) );
  NAND4_X1 U9835 ( .A1(n8778), .A2(n8777), .A3(n8776), .A4(n8775), .ZN(n8779)
         );
  NOR4_X1 U9836 ( .A1(n8782), .A2(n8781), .A3(n8780), .A4(n8779), .ZN(n8783)
         );
  NAND4_X1 U9837 ( .A1(n9278), .A2(n8784), .A3(n8783), .A4(n9290), .ZN(n8785)
         );
  NOR4_X1 U9838 ( .A1(n8787), .A2(n9254), .A3(n8786), .A4(n8785), .ZN(n8788)
         );
  NAND4_X1 U9839 ( .A1(n9182), .A2(n9202), .A3(n8803), .A4(n8788), .ZN(n8789)
         );
  NOR4_X1 U9840 ( .A1(n9128), .A2(n9153), .A3(n9171), .A4(n8789), .ZN(n8790)
         );
  NAND4_X1 U9841 ( .A1(n8791), .A2(n8790), .A3(n8814), .A4(n8817), .ZN(n8792)
         );
  XNOR2_X1 U9842 ( .A(n8792), .B(n9300), .ZN(n8793) );
  AOI21_X1 U9843 ( .B1(n6509), .B2(n8794), .A(n8793), .ZN(n8820) );
  AND2_X1 U9844 ( .A1(n9236), .A2(n9230), .ZN(n8798) );
  INV_X1 U9845 ( .A(n9024), .ZN(n9256) );
  NAND2_X1 U9846 ( .A1(n9409), .A2(n9256), .ZN(n8799) );
  INV_X1 U9847 ( .A(n8799), .ZN(n8796) );
  AND2_X1 U9848 ( .A1(n4901), .A2(n9275), .ZN(n8795) );
  OR2_X1 U9849 ( .A1(n8796), .A2(n8795), .ZN(n9228) );
  OR2_X1 U9850 ( .A1(n9254), .A2(n9228), .ZN(n8797) );
  AND2_X1 U9851 ( .A1(n9274), .A2(n8799), .ZN(n9227) );
  AND2_X1 U9852 ( .A1(n9227), .A2(n9120), .ZN(n8800) );
  NAND2_X1 U9853 ( .A1(n9221), .A2(n8804), .ZN(n9201) );
  NAND2_X1 U9854 ( .A1(n9201), .A2(n9202), .ZN(n9200) );
  NAND2_X1 U9855 ( .A1(n9175), .A2(n8808), .ZN(n9152) );
  NAND2_X1 U9856 ( .A1(n9152), .A2(n9147), .ZN(n9157) );
  OR2_X1 U9857 ( .A1(n9374), .A2(n9173), .ZN(n8809) );
  INV_X1 U9858 ( .A(n8815), .ZN(n8816) );
  XNOR2_X1 U9859 ( .A(n8821), .B(n9300), .ZN(n8822) );
  NOR4_X1 U9860 ( .A1(n8826), .A2(n8825), .A3(n8824), .A4(n9320), .ZN(n8828)
         );
  OAI21_X1 U9861 ( .B1(n8829), .B2(n6510), .A(P2_B_REG_SCAN_IN), .ZN(n8827) );
  AOI22_X1 U9862 ( .A1(n9352), .A2(n9017), .B1(n9005), .B2(n9347), .ZN(n8835)
         );
  OAI21_X1 U9863 ( .B1(n8831), .B2(n5229), .A(n8830), .ZN(n8832) );
  AOI22_X1 U9864 ( .A1(n8833), .A2(P2_REG3_REG_1__SCAN_IN), .B1(n8941), .B2(
        n8832), .ZN(n8834) );
  OAI211_X1 U9865 ( .C1(n8836), .C2(n9014), .A(n8835), .B(n8834), .ZN(P2_U3224) );
  XNOR2_X1 U9866 ( .A(n9426), .B(n8933), .ZN(n8840) );
  INV_X1 U9867 ( .A(n8840), .ZN(n8838) );
  NOR2_X1 U9868 ( .A1(n8837), .A2(n8932), .ZN(n8839) );
  NAND2_X1 U9869 ( .A1(n8838), .A2(n8839), .ZN(n8845) );
  INV_X1 U9870 ( .A(n8845), .ZN(n8841) );
  XNOR2_X1 U9871 ( .A(n8840), .B(n8839), .ZN(n8999) );
  NOR2_X1 U9872 ( .A1(n8841), .A2(n8999), .ZN(n8847) );
  OR2_X1 U9873 ( .A1(n8996), .A2(n8847), .ZN(n8913) );
  XNOR2_X1 U9874 ( .A(n9422), .B(n8931), .ZN(n8844) );
  NAND2_X1 U9875 ( .A1(n5116), .A2(n9025), .ZN(n8842) );
  XNOR2_X1 U9876 ( .A(n8844), .B(n8842), .ZN(n8916) );
  INV_X1 U9877 ( .A(n8916), .ZN(n8848) );
  OR2_X1 U9878 ( .A1(n8913), .A2(n8848), .ZN(n8850) );
  INV_X1 U9879 ( .A(n8842), .ZN(n8843) );
  AND2_X1 U9880 ( .A1(n8997), .A2(n8845), .ZN(n8846) );
  OR2_X1 U9881 ( .A1(n8847), .A2(n8846), .ZN(n8914) );
  XNOR2_X1 U9882 ( .A(n9416), .B(n8933), .ZN(n8858) );
  NOR2_X1 U9883 ( .A1(n9118), .A2(n8932), .ZN(n8859) );
  XNOR2_X1 U9884 ( .A(n8858), .B(n8859), .ZN(n8976) );
  XNOR2_X1 U9885 ( .A(n9409), .B(n8931), .ZN(n8854) );
  NAND2_X1 U9886 ( .A1(n9024), .A2(n5116), .ZN(n8853) );
  INV_X1 U9887 ( .A(n8853), .ZN(n8852) );
  NAND2_X1 U9888 ( .A1(n8854), .A2(n8852), .ZN(n8861) );
  INV_X1 U9889 ( .A(n8861), .ZN(n8855) );
  XNOR2_X1 U9890 ( .A(n8854), .B(n8853), .ZN(n8955) );
  OR2_X1 U9891 ( .A1(n8855), .A2(n8955), .ZN(n8857) );
  AND2_X1 U9892 ( .A1(n8976), .A2(n8857), .ZN(n8856) );
  INV_X1 U9893 ( .A(n8857), .ZN(n8863) );
  INV_X1 U9894 ( .A(n8858), .ZN(n8860) );
  NAND2_X1 U9895 ( .A1(n8860), .A2(n8859), .ZN(n8953) );
  AND2_X1 U9896 ( .A1(n8953), .A2(n8861), .ZN(n8862) );
  OR2_X1 U9897 ( .A1(n8863), .A2(n8862), .ZN(n8985) );
  XNOR2_X1 U9898 ( .A(n9404), .B(n8933), .ZN(n8864) );
  OR2_X1 U9899 ( .A1(n8957), .A2(n8932), .ZN(n8865) );
  NAND2_X1 U9900 ( .A1(n8864), .A2(n8865), .ZN(n8871) );
  INV_X1 U9901 ( .A(n8864), .ZN(n8867) );
  INV_X1 U9902 ( .A(n8865), .ZN(n8866) );
  NAND2_X1 U9903 ( .A1(n8867), .A2(n8866), .ZN(n8868) );
  NAND2_X1 U9904 ( .A1(n8871), .A2(n8868), .ZN(n8989) );
  INV_X1 U9905 ( .A(n8989), .ZN(n8869) );
  AND2_X1 U9906 ( .A1(n8985), .A2(n8869), .ZN(n8870) );
  NAND2_X1 U9907 ( .A1(n8987), .A2(n8871), .ZN(n8875) );
  XNOR2_X1 U9908 ( .A(n8872), .B(n8931), .ZN(n8873) );
  XNOR2_X1 U9909 ( .A(n8875), .B(n8873), .ZN(n8898) );
  OR2_X1 U9910 ( .A1(n9257), .A2(n8932), .ZN(n8897) );
  NAND2_X1 U9911 ( .A1(n8898), .A2(n8897), .ZN(n8896) );
  INV_X1 U9912 ( .A(n8873), .ZN(n8874) );
  NAND2_X1 U9913 ( .A1(n8875), .A2(n8874), .ZN(n8876) );
  NAND2_X1 U9914 ( .A1(n8896), .A2(n8876), .ZN(n8879) );
  XNOR2_X1 U9915 ( .A(n9394), .B(n8931), .ZN(n8877) );
  XNOR2_X1 U9916 ( .A(n8879), .B(n8877), .ZN(n8970) );
  NOR2_X1 U9917 ( .A1(n9206), .A2(n8932), .ZN(n8971) );
  NAND2_X1 U9918 ( .A1(n8970), .A2(n8971), .ZN(n8881) );
  INV_X1 U9919 ( .A(n8877), .ZN(n8878) );
  OR2_X1 U9920 ( .A1(n8879), .A2(n8878), .ZN(n8880) );
  NAND2_X1 U9921 ( .A1(n8881), .A2(n8880), .ZN(n8965) );
  XNOR2_X1 U9922 ( .A(n9391), .B(n8933), .ZN(n8883) );
  NAND2_X1 U9923 ( .A1(n8882), .A2(n5116), .ZN(n8884) );
  NAND2_X1 U9924 ( .A1(n8883), .A2(n8884), .ZN(n8888) );
  INV_X1 U9925 ( .A(n8883), .ZN(n8886) );
  INV_X1 U9926 ( .A(n8884), .ZN(n8885) );
  NAND2_X1 U9927 ( .A1(n8886), .A2(n8885), .ZN(n8887) );
  NAND2_X1 U9928 ( .A1(n8888), .A2(n8887), .ZN(n8964) );
  XNOR2_X1 U9929 ( .A(n9386), .B(n8931), .ZN(n8890) );
  NOR2_X1 U9930 ( .A1(n9172), .A2(n8932), .ZN(n8889) );
  XNOR2_X1 U9931 ( .A(n8890), .B(n8889), .ZN(n9009) );
  NAND2_X1 U9932 ( .A1(n8890), .A2(n8889), .ZN(n8891) );
  XNOR2_X1 U9933 ( .A(n9379), .B(n8933), .ZN(n8926) );
  NOR2_X1 U9934 ( .A1(n9185), .A2(n8932), .ZN(n8927) );
  XNOR2_X1 U9935 ( .A(n8926), .B(n8927), .ZN(n8929) );
  XNOR2_X1 U9936 ( .A(n8930), .B(n8929), .ZN(n8895) );
  OAI22_X1 U9937 ( .A1(n9011), .A2(n9173), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9651), .ZN(n8893) );
  OAI22_X1 U9938 ( .A1(n9014), .A2(n9172), .B1(n9013), .B2(n9166), .ZN(n8892)
         );
  AOI211_X1 U9939 ( .C1(n9379), .C2(n9017), .A(n8893), .B(n8892), .ZN(n8894)
         );
  OAI21_X1 U9940 ( .B1(n8895), .B2(n9019), .A(n8894), .ZN(P2_U3216) );
  OAI21_X1 U9941 ( .B1(n8898), .B2(n8897), .A(n8896), .ZN(n8902) );
  INV_X1 U9942 ( .A(n8872), .ZN(n9244) );
  AOI22_X1 U9943 ( .A1(n9005), .A2(n9233), .B1(P2_REG3_REG_23__SCAN_IN), .B2(
        P2_U3152), .ZN(n8900) );
  AOI22_X1 U9944 ( .A1(n8947), .A2(n9280), .B1(n9242), .B2(n8949), .ZN(n8899)
         );
  OAI211_X1 U9945 ( .C1(n9244), .C2(n8937), .A(n8900), .B(n8899), .ZN(n8901)
         );
  AOI21_X1 U9946 ( .B1(n8902), .B2(n8941), .A(n8901), .ZN(n8903) );
  INV_X1 U9947 ( .A(n8903), .ZN(P2_U3218) );
  AOI22_X1 U9948 ( .A1(n8904), .A2(n9017), .B1(n9005), .B2(n9039), .ZN(n8912)
         );
  NAND2_X1 U9949 ( .A1(n8906), .A2(n8905), .ZN(n8907) );
  XOR2_X1 U9950 ( .A(n8908), .B(n8907), .Z(n8909) );
  AOI22_X1 U9951 ( .A1(n8947), .A2(n9347), .B1(n8909), .B2(n8941), .ZN(n8911)
         );
  MUX2_X1 U9952 ( .A(P2_STATE_REG_SCAN_IN), .B(n9013), .S(n9578), .Z(n8910) );
  NAND3_X1 U9953 ( .A1(n8912), .A2(n8911), .A3(n8910), .ZN(P2_U3220) );
  OR2_X1 U9954 ( .A1(n8851), .A2(n8913), .ZN(n8915) );
  NAND2_X1 U9955 ( .A1(n8915), .A2(n8914), .ZN(n8917) );
  XNOR2_X1 U9956 ( .A(n8917), .B(n8916), .ZN(n8925) );
  INV_X1 U9957 ( .A(n8918), .ZN(n8922) );
  NOR2_X1 U9958 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9532), .ZN(n9099) );
  AOI21_X1 U9959 ( .B1(n8920), .B2(n8919), .A(n9099), .ZN(n8921) );
  OAI21_X1 U9960 ( .B1(n9013), .B2(n8922), .A(n8921), .ZN(n8923) );
  AOI21_X1 U9961 ( .B1(n9422), .B2(n9017), .A(n8923), .ZN(n8924) );
  OAI21_X1 U9962 ( .B1(n8925), .B2(n9019), .A(n8924), .ZN(P2_U3221) );
  INV_X1 U9963 ( .A(n8926), .ZN(n8928) );
  INV_X1 U9964 ( .A(n9374), .ZN(n9151) );
  NOR2_X1 U9965 ( .A1(n8932), .A2(n8931), .ZN(n8935) );
  NAND2_X1 U9966 ( .A1(n9173), .A2(n8933), .ZN(n8934) );
  OAI21_X1 U9967 ( .B1(n9173), .B2(n8935), .A(n8934), .ZN(n8939) );
  NOR3_X1 U9968 ( .A1(n9151), .A2(n9017), .A3(n8939), .ZN(n8936) );
  AOI21_X1 U9969 ( .B1(n9151), .B2(n8939), .A(n8936), .ZN(n8945) );
  NAND3_X1 U9970 ( .A1(n9374), .A2(n8937), .A3(n8939), .ZN(n8938) );
  OAI21_X1 U9971 ( .B1(n9374), .B2(n8939), .A(n8938), .ZN(n8940) );
  NAND2_X1 U9972 ( .A1(n8946), .A2(n8940), .ZN(n8944) );
  AOI21_X1 U9973 ( .B1(n9374), .B2(n9017), .A(n8941), .ZN(n8942) );
  OAI211_X1 U9974 ( .C1(n8946), .C2(n8945), .A(n8944), .B(n8943), .ZN(n8952)
         );
  INV_X1 U9975 ( .A(n9185), .ZN(n9023) );
  AOI22_X1 U9976 ( .A1(n8947), .A2(n9023), .B1(P2_REG3_REG_28__SCAN_IN), .B2(
        P2_U3152), .ZN(n8951) );
  INV_X1 U9977 ( .A(n9155), .ZN(n9021) );
  INV_X1 U9978 ( .A(n8948), .ZN(n9149) );
  AOI22_X1 U9979 ( .A1(n9005), .A2(n9021), .B1(n9149), .B2(n8949), .ZN(n8950)
         );
  NAND3_X1 U9980 ( .A1(n8952), .A2(n8951), .A3(n8950), .ZN(P2_U3222) );
  NAND2_X1 U9981 ( .A1(n8977), .A2(n8976), .ZN(n8954) );
  NAND2_X1 U9982 ( .A1(n8954), .A2(n8953), .ZN(n8956) );
  XNOR2_X1 U9983 ( .A(n8956), .B(n8955), .ZN(n8961) );
  OAI22_X1 U9984 ( .A1(n9011), .A2(n8957), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9540), .ZN(n8959) );
  OAI22_X1 U9985 ( .A1(n9014), .A2(n9118), .B1(n9013), .B2(n9269), .ZN(n8958)
         );
  AOI211_X1 U9986 ( .C1(n9409), .C2(n9017), .A(n8959), .B(n8958), .ZN(n8960)
         );
  OAI21_X1 U9987 ( .B1(n8961), .B2(n9019), .A(n8960), .ZN(P2_U3225) );
  INV_X1 U9988 ( .A(n8962), .ZN(n8963) );
  AOI21_X1 U9989 ( .B1(n8965), .B2(n8964), .A(n8963), .ZN(n8969) );
  OAI22_X1 U9990 ( .A1(n9011), .A2(n9172), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9469), .ZN(n8967) );
  OAI22_X1 U9991 ( .A1(n9014), .A2(n9206), .B1(n9013), .B2(n9194), .ZN(n8966)
         );
  AOI211_X1 U9992 ( .C1(n9391), .C2(n9017), .A(n8967), .B(n8966), .ZN(n8968)
         );
  OAI21_X1 U9993 ( .B1(n8969), .B2(n9019), .A(n8968), .ZN(P2_U3227) );
  XNOR2_X1 U9994 ( .A(n8970), .B(n8971), .ZN(n8975) );
  OAI22_X1 U9995 ( .A1(n9011), .A2(n9219), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9674), .ZN(n8973) );
  OAI22_X1 U9996 ( .A1(n9014), .A2(n9257), .B1(n9013), .B2(n9214), .ZN(n8972)
         );
  AOI211_X1 U9997 ( .C1(n9394), .C2(n9017), .A(n8973), .B(n8972), .ZN(n8974)
         );
  OAI21_X1 U9998 ( .B1(n8975), .B2(n9019), .A(n8974), .ZN(P2_U3231) );
  XNOR2_X1 U9999 ( .A(n8977), .B(n8976), .ZN(n8984) );
  OAI22_X1 U10000 ( .A1(n9011), .A2(n9256), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9557), .ZN(n8982) );
  INV_X1 U10001 ( .A(n8978), .ZN(n8979) );
  OAI22_X1 U10002 ( .A1(n9014), .A2(n8980), .B1(n9013), .B2(n8979), .ZN(n8981)
         );
  AOI211_X1 U10003 ( .C1(n9416), .C2(n9017), .A(n8982), .B(n8981), .ZN(n8983)
         );
  OAI21_X1 U10004 ( .B1(n8984), .B2(n9019), .A(n8983), .ZN(P2_U3235) );
  NAND2_X1 U10005 ( .A1(n8986), .A2(n8985), .ZN(n8990) );
  INV_X1 U10006 ( .A(n8987), .ZN(n8988) );
  AOI21_X1 U10007 ( .B1(n8990), .B2(n8989), .A(n8988), .ZN(n8995) );
  OAI22_X1 U10008 ( .A1(n9011), .A2(n9257), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9575), .ZN(n8993) );
  INV_X1 U10009 ( .A(n9250), .ZN(n8991) );
  OAI22_X1 U10010 ( .A1(n9014), .A2(n9256), .B1(n9013), .B2(n8991), .ZN(n8992)
         );
  AOI211_X1 U10011 ( .C1(n9404), .C2(n9017), .A(n8993), .B(n8992), .ZN(n8994)
         );
  OAI21_X1 U10012 ( .B1(n8995), .B2(n9019), .A(n8994), .ZN(P2_U3237) );
  OR2_X1 U10013 ( .A1(n8851), .A2(n8996), .ZN(n8998) );
  NAND2_X1 U10014 ( .A1(n8998), .A2(n8997), .ZN(n9000) );
  XNOR2_X1 U10015 ( .A(n9000), .B(n8999), .ZN(n9008) );
  AND2_X1 U10016 ( .A1(P2_U3152), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n9082) );
  INV_X1 U10017 ( .A(n9001), .ZN(n9002) );
  OAI22_X1 U10018 ( .A1(n9014), .A2(n9003), .B1(n9013), .B2(n9002), .ZN(n9004)
         );
  AOI211_X1 U10019 ( .C1(n9005), .C2(n9025), .A(n9082), .B(n9004), .ZN(n9007)
         );
  NAND2_X1 U10020 ( .A1(n9426), .A2(n9017), .ZN(n9006) );
  OAI211_X1 U10021 ( .C1(n9008), .C2(n9019), .A(n9007), .B(n9006), .ZN(
        P2_U3240) );
  XNOR2_X1 U10022 ( .A(n9010), .B(n9009), .ZN(n9020) );
  OAI22_X1 U10023 ( .A1(n9011), .A2(n9185), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9689), .ZN(n9016) );
  INV_X1 U10024 ( .A(n9188), .ZN(n9012) );
  OAI22_X1 U10025 ( .A1(n9014), .A2(n9219), .B1(n9013), .B2(n9012), .ZN(n9015)
         );
  AOI211_X1 U10026 ( .C1(n9386), .C2(n9017), .A(n9016), .B(n9015), .ZN(n9018)
         );
  OAI21_X1 U10027 ( .B1(n9020), .B2(n9019), .A(n9018), .ZN(P2_U3242) );
  MUX2_X1 U10028 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(n9109), .S(n9041), .Z(
        P2_U3583) );
  MUX2_X1 U10029 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(n9131), .S(n9041), .Z(
        P2_U3582) );
  MUX2_X1 U10030 ( .A(n9021), .B(P2_DATAO_REG_29__SCAN_IN), .S(n9022), .Z(
        P2_U3581) );
  INV_X1 U10031 ( .A(n9173), .ZN(n9133) );
  MUX2_X1 U10032 ( .A(n9133), .B(P2_DATAO_REG_28__SCAN_IN), .S(n9022), .Z(
        P2_U3580) );
  MUX2_X1 U10033 ( .A(n9023), .B(P2_DATAO_REG_27__SCAN_IN), .S(n9022), .Z(
        P2_U3579) );
  MUX2_X1 U10034 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(n9233), .S(n9041), .Z(
        P2_U3576) );
  INV_X1 U10035 ( .A(n9257), .ZN(n9121) );
  MUX2_X1 U10036 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(n9121), .S(P2_U3966), .Z(
        P2_U3575) );
  MUX2_X1 U10037 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n9280), .S(P2_U3966), .Z(
        P2_U3574) );
  MUX2_X1 U10038 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n9024), .S(P2_U3966), .Z(
        P2_U3573) );
  INV_X1 U10039 ( .A(n9118), .ZN(n9281) );
  MUX2_X1 U10040 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n9281), .S(P2_U3966), .Z(
        P2_U3572) );
  MUX2_X1 U10041 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n9025), .S(P2_U3966), .Z(
        P2_U3571) );
  MUX2_X1 U10042 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(n9026), .S(P2_U3966), .Z(
        P2_U3570) );
  MUX2_X1 U10043 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n9027), .S(P2_U3966), .Z(
        P2_U3569) );
  MUX2_X1 U10044 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n9028), .S(P2_U3966), .Z(
        P2_U3568) );
  MUX2_X1 U10045 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(n9029), .S(P2_U3966), .Z(
        P2_U3567) );
  MUX2_X1 U10046 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(n9030), .S(n9041), .Z(
        P2_U3566) );
  MUX2_X1 U10047 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(n9031), .S(n9041), .Z(
        P2_U3565) );
  MUX2_X1 U10048 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(n9032), .S(n9041), .Z(
        P2_U3564) );
  MUX2_X1 U10049 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(n9033), .S(n9041), .Z(
        P2_U3563) );
  MUX2_X1 U10050 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(n9034), .S(n9041), .Z(
        P2_U3562) );
  MUX2_X1 U10051 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(n9035), .S(n9041), .Z(
        P2_U3561) );
  MUX2_X1 U10052 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(n9036), .S(n9041), .Z(
        P2_U3560) );
  MUX2_X1 U10053 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(n9037), .S(n9041), .Z(
        P2_U3559) );
  MUX2_X1 U10054 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(n9038), .S(n9041), .Z(
        P2_U3557) );
  MUX2_X1 U10055 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(n9039), .S(n9041), .Z(
        P2_U3556) );
  MUX2_X1 U10056 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(n9040), .S(n9041), .Z(
        P2_U3555) );
  MUX2_X1 U10057 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(n9347), .S(n9041), .Z(
        P2_U3554) );
  MUX2_X1 U10058 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(n9042), .S(n9041), .Z(
        P2_U3553) );
  OAI21_X1 U10059 ( .B1(n9045), .B2(n9044), .A(n9043), .ZN(n9046) );
  NAND2_X1 U10060 ( .A1(n10466), .A2(n9046), .ZN(n9055) );
  NOR2_X1 U10061 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9561), .ZN(n9047) );
  AOI21_X1 U10062 ( .B1(n10486), .B2(P2_ADDR_REG_11__SCAN_IN), .A(n9047), .ZN(
        n9054) );
  NAND2_X1 U10063 ( .A1(n10493), .A2(n9048), .ZN(n9053) );
  OAI211_X1 U10064 ( .C1(n9051), .C2(n9050), .A(n10495), .B(n9049), .ZN(n9052)
         );
  NAND4_X1 U10065 ( .A1(n9055), .A2(n9054), .A3(n9053), .A4(n9052), .ZN(
        P2_U3256) );
  OAI21_X1 U10066 ( .B1(n9058), .B2(n9057), .A(n9056), .ZN(n9059) );
  NAND2_X1 U10067 ( .A1(n9059), .A2(n10466), .ZN(n9068) );
  OAI211_X1 U10068 ( .C1(n9061), .C2(P2_REG1_REG_15__SCAN_IN), .A(n10495), .B(
        n9060), .ZN(n9067) );
  INV_X1 U10069 ( .A(n9062), .ZN(n9063) );
  AOI21_X1 U10070 ( .B1(n10486), .B2(P2_ADDR_REG_15__SCAN_IN), .A(n9063), .ZN(
        n9066) );
  NAND2_X1 U10071 ( .A1(n10493), .A2(n9064), .ZN(n9065) );
  NAND4_X1 U10072 ( .A1(n9068), .A2(n9067), .A3(n9066), .A4(n9065), .ZN(
        P2_U3260) );
  INV_X1 U10073 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n9069) );
  MUX2_X1 U10074 ( .A(n9069), .B(P2_REG2_REG_18__SCAN_IN), .S(n9088), .Z(n9073) );
  AOI21_X1 U10075 ( .B1(n9076), .B2(P2_REG2_REG_17__SCAN_IN), .A(n9070), .ZN(
        n9071) );
  INV_X1 U10076 ( .A(n9071), .ZN(n9072) );
  AOI21_X1 U10077 ( .B1(n9073), .B2(n9072), .A(n9089), .ZN(n9086) );
  NOR2_X1 U10078 ( .A1(n9088), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n9094) );
  AOI21_X1 U10079 ( .B1(n9088), .B2(P2_REG1_REG_18__SCAN_IN), .A(n9094), .ZN(
        n9078) );
  INV_X1 U10080 ( .A(n9074), .ZN(n9075) );
  AOI21_X1 U10081 ( .B1(n9076), .B2(P2_REG1_REG_17__SCAN_IN), .A(n9075), .ZN(
        n9077) );
  NAND2_X1 U10082 ( .A1(n9078), .A2(n9077), .ZN(n9096) );
  OAI21_X1 U10083 ( .B1(n9078), .B2(n9077), .A(n9096), .ZN(n9083) );
  INV_X1 U10084 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n9079) );
  NOR2_X1 U10085 ( .A1(n9080), .A2(n9079), .ZN(n9081) );
  AOI211_X1 U10086 ( .C1(n10495), .C2(n9083), .A(n9082), .B(n9081), .ZN(n9085)
         );
  NAND2_X1 U10087 ( .A1(n10493), .A2(n9088), .ZN(n9084) );
  OAI211_X1 U10088 ( .C1(n9086), .C2(n10487), .A(n9085), .B(n9084), .ZN(
        P2_U3263) );
  INV_X1 U10089 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n9087) );
  MUX2_X1 U10090 ( .A(P2_REG2_REG_19__SCAN_IN), .B(n9087), .S(n9300), .Z(n9092) );
  INV_X1 U10091 ( .A(n9088), .ZN(n9090) );
  AOI21_X1 U10092 ( .B1(n9069), .B2(n9090), .A(n9089), .ZN(n9091) );
  XOR2_X1 U10093 ( .A(n9092), .B(n9091), .Z(n9105) );
  INV_X1 U10094 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n9093) );
  MUX2_X1 U10095 ( .A(n9093), .B(P2_REG1_REG_19__SCAN_IN), .S(n9300), .Z(n9098) );
  INV_X1 U10096 ( .A(n9094), .ZN(n9095) );
  NAND2_X1 U10097 ( .A1(n9096), .A2(n9095), .ZN(n9097) );
  XOR2_X1 U10098 ( .A(n9098), .B(n9097), .Z(n9101) );
  AOI21_X1 U10099 ( .B1(n10486), .B2(P2_ADDR_REG_19__SCAN_IN), .A(n9099), .ZN(
        n9100) );
  OAI21_X1 U10100 ( .B1(n10468), .B2(n9101), .A(n9100), .ZN(n9102) );
  AOI21_X1 U10101 ( .B1(n9103), .B2(n10493), .A(n9102), .ZN(n9104) );
  OAI21_X1 U10102 ( .B1(n9105), .B2(n10487), .A(n9104), .ZN(P2_U3264) );
  INV_X1 U10103 ( .A(n9391), .ZN(n9123) );
  INV_X1 U10104 ( .A(n9409), .ZN(n9273) );
  NAND2_X1 U10105 ( .A1(n9123), .A2(n9196), .ZN(n9197) );
  XNOR2_X1 U10106 ( .A(n9112), .B(n9106), .ZN(n9359) );
  NAND2_X1 U10107 ( .A1(n9359), .A2(n9353), .ZN(n9111) );
  AND2_X1 U10108 ( .A1(n9107), .A2(P2_B_REG_SCAN_IN), .ZN(n9108) );
  NOR2_X1 U10109 ( .A1(n9318), .A2(n9108), .ZN(n9132) );
  NAND2_X1 U10110 ( .A1(n9109), .A2(n9132), .ZN(n9366) );
  NOR2_X1 U10111 ( .A1(n9223), .A2(n9366), .ZN(n9114) );
  AOI21_X1 U10112 ( .B1(n9354), .B2(P2_REG2_REG_31__SCAN_IN), .A(n9114), .ZN(
        n9110) );
  OAI211_X1 U10113 ( .C1(n9360), .C2(n9272), .A(n9111), .B(n9110), .ZN(
        P2_U3265) );
  NAND2_X1 U10114 ( .A1(n9138), .A2(n9113), .ZN(n9364) );
  NAND3_X1 U10115 ( .A1(n9365), .A2(n9353), .A3(n9364), .ZN(n9116) );
  AOI21_X1 U10116 ( .B1(n9223), .B2(P2_REG2_REG_30__SCAN_IN), .A(n9114), .ZN(
        n9115) );
  OAI211_X1 U10117 ( .C1(n9368), .C2(n9272), .A(n9116), .B(n9115), .ZN(
        P2_U3266) );
  NOR2_X1 U10118 ( .A1(n9237), .A2(n9236), .ZN(n9235) );
  NOR2_X1 U10119 ( .A1(n9235), .A2(n9122), .ZN(n9212) );
  NAND2_X1 U10120 ( .A1(n9212), .A2(n9218), .ZN(n9211) );
  OAI21_X1 U10121 ( .B1(n9394), .B2(n9233), .A(n9211), .ZN(n9193) );
  INV_X1 U10122 ( .A(n9379), .ZN(n9169) );
  NAND2_X1 U10123 ( .A1(n9148), .A2(n9153), .ZN(n9126) );
  NAND2_X1 U10124 ( .A1(n9126), .A2(n9125), .ZN(n9129) );
  XNOR2_X1 U10125 ( .A(n9129), .B(n9128), .ZN(n9369) );
  INV_X1 U10126 ( .A(n9369), .ZN(n9146) );
  XOR2_X1 U10127 ( .A(n9128), .B(n9130), .Z(n9135) );
  AOI22_X1 U10128 ( .A1(n9133), .A2(n9345), .B1(n9132), .B2(n9131), .ZN(n9134)
         );
  OAI21_X1 U10129 ( .B1(n9135), .B2(n9253), .A(n9134), .ZN(n9372) );
  INV_X1 U10130 ( .A(n9136), .ZN(n9370) );
  OAI21_X1 U10131 ( .B1(n9370), .B2(n9137), .A(n9138), .ZN(n9371) );
  NOR2_X1 U10132 ( .A1(n9371), .A2(n9139), .ZN(n9144) );
  INV_X1 U10133 ( .A(n9140), .ZN(n9141) );
  AOI22_X1 U10134 ( .A1(n9354), .A2(P2_REG2_REG_29__SCAN_IN), .B1(n9141), .B2(
        n9350), .ZN(n9142) );
  OAI21_X1 U10135 ( .B1(n9370), .B2(n9272), .A(n9142), .ZN(n9143) );
  AOI211_X1 U10136 ( .C1(n9372), .C2(n9307), .A(n9144), .B(n9143), .ZN(n9145)
         );
  OAI21_X1 U10137 ( .B1(n9146), .B2(n9285), .A(n9145), .ZN(P2_U3267) );
  XNOR2_X1 U10138 ( .A(n9148), .B(n9147), .ZN(n9378) );
  AOI21_X1 U10139 ( .B1(n9374), .B2(n9164), .A(n9137), .ZN(n9375) );
  AOI22_X1 U10140 ( .A1(n9223), .A2(P2_REG2_REG_28__SCAN_IN), .B1(n9149), .B2(
        n9350), .ZN(n9150) );
  OAI21_X1 U10141 ( .B1(n9151), .B2(n9272), .A(n9150), .ZN(n9160) );
  INV_X1 U10142 ( .A(n9152), .ZN(n9154) );
  AOI21_X1 U10143 ( .B1(n9154), .B2(n9153), .A(n9253), .ZN(n9158) );
  OAI22_X1 U10144 ( .A1(n9155), .A2(n9318), .B1(n9185), .B2(n9320), .ZN(n9156)
         );
  AOI21_X1 U10145 ( .B1(n9158), .B2(n9157), .A(n9156), .ZN(n9377) );
  NOR2_X1 U10146 ( .A1(n9377), .A2(n9223), .ZN(n9159) );
  AOI211_X1 U10147 ( .C1(n9353), .C2(n9375), .A(n9160), .B(n9159), .ZN(n9161)
         );
  OAI21_X1 U10148 ( .B1(n9378), .B2(n9285), .A(n9161), .ZN(P2_U3268) );
  XOR2_X1 U10149 ( .A(n9171), .B(n9162), .Z(n9383) );
  INV_X1 U10150 ( .A(n9164), .ZN(n9165) );
  AOI21_X1 U10151 ( .B1(n9379), .B2(n9186), .A(n9165), .ZN(n9380) );
  INV_X1 U10152 ( .A(n9166), .ZN(n9167) );
  AOI22_X1 U10153 ( .A1(n9223), .A2(P2_REG2_REG_27__SCAN_IN), .B1(n9167), .B2(
        n9350), .ZN(n9168) );
  OAI21_X1 U10154 ( .B1(n9169), .B2(n9272), .A(n9168), .ZN(n9178) );
  AOI21_X1 U10155 ( .B1(n9170), .B2(n9171), .A(n9253), .ZN(n9176) );
  OAI22_X1 U10156 ( .A1(n9173), .A2(n9318), .B1(n9172), .B2(n9320), .ZN(n9174)
         );
  AOI21_X1 U10157 ( .B1(n9176), .B2(n9175), .A(n9174), .ZN(n9382) );
  NOR2_X1 U10158 ( .A1(n9382), .A2(n9223), .ZN(n9177) );
  AOI211_X1 U10159 ( .C1(n9353), .C2(n9380), .A(n9178), .B(n9177), .ZN(n9179)
         );
  OAI21_X1 U10160 ( .B1(n9383), .B2(n9285), .A(n9179), .ZN(P2_U3269) );
  XOR2_X1 U10161 ( .A(n9182), .B(n9180), .Z(n9388) );
  NAND2_X1 U10162 ( .A1(n9200), .A2(n9181), .ZN(n9183) );
  XNOR2_X1 U10163 ( .A(n9183), .B(n9182), .ZN(n9184) );
  OAI222_X1 U10164 ( .A1(n9318), .A2(n9185), .B1(n9320), .B2(n9219), .C1(n9253), .C2(n9184), .ZN(n9384) );
  AOI211_X1 U10165 ( .C1(n9386), .C2(n9197), .A(n10637), .B(n9163), .ZN(n9385)
         );
  NAND2_X1 U10166 ( .A1(n9385), .A2(n9187), .ZN(n9190) );
  AOI22_X1 U10167 ( .A1(n9223), .A2(P2_REG2_REG_26__SCAN_IN), .B1(n9188), .B2(
        n9350), .ZN(n9189) );
  OAI211_X1 U10168 ( .C1(n5048), .C2(n9272), .A(n9190), .B(n9189), .ZN(n9191)
         );
  AOI21_X1 U10169 ( .B1(n9384), .B2(n9307), .A(n9191), .ZN(n9192) );
  OAI21_X1 U10170 ( .B1(n9388), .B2(n9285), .A(n9192), .ZN(P2_U3270) );
  XNOR2_X1 U10171 ( .A(n9193), .B(n9202), .ZN(n9393) );
  INV_X1 U10172 ( .A(P2_REG2_REG_25__SCAN_IN), .ZN(n9195) );
  OAI22_X1 U10173 ( .A1(n9307), .A2(n9195), .B1(n9194), .B2(n9304), .ZN(n9209)
         );
  INV_X1 U10174 ( .A(n9196), .ZN(n9199) );
  INV_X1 U10175 ( .A(n9197), .ZN(n9198) );
  AOI211_X1 U10176 ( .C1(n9391), .C2(n9199), .A(n10637), .B(n9198), .ZN(n9390)
         );
  OAI211_X1 U10177 ( .C1(n9202), .C2(n9201), .A(n9200), .B(n9340), .ZN(n9205)
         );
  NAND2_X1 U10178 ( .A1(n9203), .A2(n9346), .ZN(n9204) );
  OAI211_X1 U10179 ( .C1(n9206), .C2(n9320), .A(n9205), .B(n9204), .ZN(n9389)
         );
  AOI21_X1 U10180 ( .B1(n9390), .B2(n9300), .A(n9389), .ZN(n9207) );
  NOR2_X1 U10181 ( .A1(n9207), .A2(n9223), .ZN(n9208) );
  AOI211_X1 U10182 ( .C1(n9336), .C2(n9391), .A(n9209), .B(n9208), .ZN(n9210)
         );
  OAI21_X1 U10183 ( .B1(n9393), .B2(n9285), .A(n9210), .ZN(P2_U3271) );
  OAI21_X1 U10184 ( .B1(n9212), .B2(n9218), .A(n9211), .ZN(n9213) );
  INV_X1 U10185 ( .A(n9213), .ZN(n9398) );
  XNOR2_X1 U10186 ( .A(n9240), .B(n9217), .ZN(n9395) );
  INV_X1 U10187 ( .A(n9214), .ZN(n9215) );
  AOI22_X1 U10188 ( .A1(n9223), .A2(P2_REG2_REG_24__SCAN_IN), .B1(n9215), .B2(
        n9350), .ZN(n9216) );
  OAI21_X1 U10189 ( .B1(n9217), .B2(n9272), .A(n9216), .ZN(n9225) );
  AOI21_X1 U10190 ( .B1(n4890), .B2(n9218), .A(n9253), .ZN(n9222) );
  OAI22_X1 U10191 ( .A1(n9219), .A2(n9318), .B1(n9257), .B2(n9320), .ZN(n9220)
         );
  AOI21_X1 U10192 ( .B1(n9222), .B2(n9221), .A(n9220), .ZN(n9397) );
  NOR2_X1 U10193 ( .A1(n9397), .A2(n9223), .ZN(n9224) );
  AOI211_X1 U10194 ( .C1(n9395), .C2(n9353), .A(n9225), .B(n9224), .ZN(n9226)
         );
  OAI21_X1 U10195 ( .B1(n9398), .B2(n9285), .A(n9226), .ZN(P2_U3272) );
  NAND2_X1 U10196 ( .A1(n8801), .A2(n9227), .ZN(n9229) );
  AND2_X1 U10197 ( .A1(n9229), .A2(n9228), .ZN(n9255) );
  OR2_X1 U10198 ( .A1(n9255), .A2(n9254), .ZN(n9259) );
  AND2_X1 U10199 ( .A1(n9259), .A2(n9230), .ZN(n9232) );
  OAI21_X1 U10200 ( .B1(n9232), .B2(n9236), .A(n9231), .ZN(n9234) );
  AOI222_X1 U10201 ( .A1(n9340), .A2(n9234), .B1(n9233), .B2(n9346), .C1(n9280), .C2(n9345), .ZN(n9402) );
  INV_X1 U10202 ( .A(n9235), .ZN(n9238) );
  NAND2_X1 U10203 ( .A1(n9237), .A2(n9236), .ZN(n9399) );
  NAND3_X1 U10204 ( .A1(n9238), .A2(n9337), .A3(n9399), .ZN(n9247) );
  INV_X1 U10205 ( .A(n9240), .ZN(n9241) );
  AOI21_X1 U10206 ( .B1(n8872), .B2(n9249), .A(n9241), .ZN(n9400) );
  AOI22_X1 U10207 ( .A1(n9223), .A2(P2_REG2_REG_23__SCAN_IN), .B1(n9242), .B2(
        n9350), .ZN(n9243) );
  OAI21_X1 U10208 ( .B1(n9244), .B2(n9272), .A(n9243), .ZN(n9245) );
  AOI21_X1 U10209 ( .B1(n9400), .B2(n9353), .A(n9245), .ZN(n9246) );
  OAI211_X1 U10210 ( .C1(n9354), .C2(n9402), .A(n9247), .B(n9246), .ZN(
        P2_U3273) );
  XNOR2_X1 U10211 ( .A(n9248), .B(n9254), .ZN(n9408) );
  AOI21_X1 U10212 ( .B1(n9404), .B2(n9267), .A(n9239), .ZN(n9405) );
  INV_X1 U10213 ( .A(n9404), .ZN(n9252) );
  AOI22_X1 U10214 ( .A1(n9354), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n9250), .B2(
        n9350), .ZN(n9251) );
  OAI21_X1 U10215 ( .B1(n9252), .B2(n9272), .A(n9251), .ZN(n9262) );
  AOI21_X1 U10216 ( .B1(n9255), .B2(n9254), .A(n9253), .ZN(n9260) );
  OAI22_X1 U10217 ( .A1(n9257), .A2(n9318), .B1(n9256), .B2(n9320), .ZN(n9258)
         );
  AOI21_X1 U10218 ( .B1(n9260), .B2(n9259), .A(n9258), .ZN(n9407) );
  NOR2_X1 U10219 ( .A1(n9407), .A2(n9223), .ZN(n9261) );
  AOI211_X1 U10220 ( .C1(n9405), .C2(n9353), .A(n9262), .B(n9261), .ZN(n9263)
         );
  OAI21_X1 U10221 ( .B1(n9408), .B2(n9285), .A(n9263), .ZN(P2_U3274) );
  AOI21_X1 U10222 ( .B1(n9278), .B2(n9265), .A(n9264), .ZN(n9413) );
  INV_X1 U10223 ( .A(n9266), .ZN(n9268) );
  AOI21_X1 U10224 ( .B1(n9409), .B2(n9268), .A(n4992), .ZN(n9410) );
  INV_X1 U10225 ( .A(n9269), .ZN(n9270) );
  AOI22_X1 U10226 ( .A1(n9354), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n9270), .B2(
        n9350), .ZN(n9271) );
  OAI21_X1 U10227 ( .B1(n9273), .B2(n9272), .A(n9271), .ZN(n9283) );
  NAND2_X1 U10228 ( .A1(n8801), .A2(n9274), .ZN(n9276) );
  NAND2_X1 U10229 ( .A1(n9276), .A2(n9275), .ZN(n9277) );
  XOR2_X1 U10230 ( .A(n9278), .B(n9277), .Z(n9279) );
  AOI222_X1 U10231 ( .A1(n9281), .A2(n9345), .B1(n9280), .B2(n9346), .C1(n9340), .C2(n9279), .ZN(n9412) );
  NOR2_X1 U10232 ( .A1(n9412), .A2(n9354), .ZN(n9282) );
  AOI211_X1 U10233 ( .C1(n9410), .C2(n9353), .A(n9283), .B(n9282), .ZN(n9284)
         );
  OAI21_X1 U10234 ( .B1(n9413), .B2(n9285), .A(n9284), .ZN(P2_U3275) );
  NAND2_X1 U10235 ( .A1(n9287), .A2(n9286), .ZN(n9289) );
  AND2_X1 U10236 ( .A1(n9289), .A2(n9288), .ZN(n9291) );
  NAND2_X1 U10237 ( .A1(n9291), .A2(n9290), .ZN(n9292) );
  XNOR2_X1 U10238 ( .A(n9295), .B(n9294), .ZN(n9297) );
  AOI21_X1 U10239 ( .B1(n9297), .B2(n9340), .A(n9296), .ZN(n9434) );
  AOI211_X1 U10240 ( .C1(n9432), .C2(n9299), .A(n10637), .B(n9298), .ZN(n9431)
         );
  NAND2_X1 U10241 ( .A1(n9431), .A2(n9300), .ZN(n9301) );
  OAI211_X1 U10242 ( .C1(n9435), .C2(n9302), .A(n9434), .B(n9301), .ZN(n9303)
         );
  NAND2_X1 U10243 ( .A1(n9303), .A2(n9307), .ZN(n9310) );
  INV_X1 U10244 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n9306) );
  OAI22_X1 U10245 ( .A1(n9307), .A2(n9306), .B1(n9305), .B2(n9304), .ZN(n9308)
         );
  AOI21_X1 U10246 ( .B1(n9432), .B2(n9336), .A(n9308), .ZN(n9309) );
  OAI211_X1 U10247 ( .C1(n9435), .C2(n9311), .A(n9310), .B(n9309), .ZN(
        P2_U3279) );
  XNOR2_X1 U10248 ( .A(n9312), .B(n9316), .ZN(n10526) );
  AOI22_X1 U10249 ( .A1(n9313), .A2(n10526), .B1(n9336), .B2(n10529), .ZN(
        n9331) );
  NAND2_X1 U10250 ( .A1(n10526), .A2(n9314), .ZN(n9326) );
  OAI211_X1 U10251 ( .C1(n9317), .C2(n9316), .A(n9315), .B(n9340), .ZN(n9324)
         );
  OAI22_X1 U10252 ( .A1(n9321), .A2(n9320), .B1(n9319), .B2(n9318), .ZN(n9322)
         );
  INV_X1 U10253 ( .A(n9322), .ZN(n9323) );
  AND2_X1 U10254 ( .A1(n9324), .A2(n9323), .ZN(n9325) );
  NAND2_X1 U10255 ( .A1(n9326), .A2(n9325), .ZN(n10535) );
  AND2_X1 U10256 ( .A1(P2_REG3_REG_2__SCAN_IN), .A2(n9350), .ZN(n9327) );
  AOI21_X1 U10257 ( .B1(n9307), .B2(n10535), .A(n9327), .ZN(n9330) );
  AND2_X1 U10258 ( .A1(n10510), .A2(n10529), .ZN(n10528) );
  NOR2_X1 U10259 ( .A1(n10527), .A2(n10528), .ZN(n9328) );
  AOI22_X1 U10260 ( .A1(n9353), .A2(n9328), .B1(n9354), .B2(
        P2_REG2_REG_2__SCAN_IN), .ZN(n9329) );
  NAND3_X1 U10261 ( .A1(n9331), .A2(n9330), .A3(n9329), .ZN(P2_U3294) );
  OR2_X1 U10262 ( .A1(n9333), .A2(n9332), .ZN(n9334) );
  AND2_X1 U10263 ( .A1(n9335), .A2(n9334), .ZN(n10516) );
  AOI22_X1 U10264 ( .A1(n10516), .A2(n9337), .B1(n9336), .B2(n9352), .ZN(n9358) );
  INV_X1 U10265 ( .A(n9338), .ZN(n9342) );
  NAND2_X1 U10266 ( .A1(n9332), .A2(n9339), .ZN(n9341) );
  OAI211_X1 U10267 ( .C1(n9343), .C2(n9342), .A(n9341), .B(n9340), .ZN(n9349)
         );
  AOI22_X1 U10268 ( .A1(n9347), .A2(n9346), .B1(n9345), .B2(n9344), .ZN(n9348)
         );
  NAND2_X1 U10269 ( .A1(n9349), .A2(n9348), .ZN(n10514) );
  AOI22_X1 U10270 ( .A1(n9307), .A2(n10514), .B1(P2_REG3_REG_1__SCAN_IN), .B2(
        n9350), .ZN(n9357) );
  NAND2_X1 U10271 ( .A1(n9352), .A2(n9351), .ZN(n10509) );
  NAND3_X1 U10272 ( .A1(n9353), .A2(n10510), .A3(n10509), .ZN(n9356) );
  NAND2_X1 U10273 ( .A1(n9354), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n9355) );
  NAND4_X1 U10274 ( .A1(n9358), .A2(n9357), .A3(n9356), .A4(n9355), .ZN(
        P2_U3295) );
  OAI21_X1 U10275 ( .B1(n9360), .B2(n10625), .A(n9366), .ZN(n9361) );
  INV_X1 U10276 ( .A(n9361), .ZN(n9362) );
  MUX2_X1 U10277 ( .A(P2_REG1_REG_31__SCAN_IN), .B(n9456), .S(n10642), .Z(
        P2_U3551) );
  OAI211_X1 U10278 ( .C1(n9368), .C2(n10625), .A(n9367), .B(n9366), .ZN(n9457)
         );
  MUX2_X1 U10279 ( .A(P2_REG1_REG_30__SCAN_IN), .B(n9457), .S(n10642), .Z(
        P2_U3550) );
  NAND2_X1 U10280 ( .A1(n9369), .A2(n10639), .ZN(n9373) );
  AOI22_X1 U10281 ( .A1(n9375), .A2(n10511), .B1(n10632), .B2(n9374), .ZN(
        n9376) );
  OAI211_X1 U10282 ( .C1(n9378), .C2(n10556), .A(n9377), .B(n9376), .ZN(n9459)
         );
  MUX2_X1 U10283 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n9459), .S(n10642), .Z(
        P2_U3548) );
  AOI22_X1 U10284 ( .A1(n9380), .A2(n10511), .B1(n10632), .B2(n9379), .ZN(
        n9381) );
  OAI211_X1 U10285 ( .C1(n9383), .C2(n10556), .A(n9382), .B(n9381), .ZN(n9460)
         );
  MUX2_X1 U10286 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n9460), .S(n10642), .Z(
        P2_U3547) );
  AOI211_X1 U10287 ( .C1(n10632), .C2(n9386), .A(n9385), .B(n9384), .ZN(n9387)
         );
  OAI21_X1 U10288 ( .B1(n9388), .B2(n10556), .A(n9387), .ZN(n9461) );
  MUX2_X1 U10289 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n9461), .S(n10642), .Z(
        P2_U3546) );
  AOI211_X1 U10290 ( .C1(n10632), .C2(n9391), .A(n9390), .B(n9389), .ZN(n9392)
         );
  OAI21_X1 U10291 ( .B1(n9393), .B2(n10556), .A(n9392), .ZN(n9462) );
  MUX2_X1 U10292 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n9462), .S(n10642), .Z(
        P2_U3545) );
  AOI22_X1 U10293 ( .A1(n9395), .A2(n10511), .B1(n10632), .B2(n9394), .ZN(
        n9396) );
  OAI211_X1 U10294 ( .C1(n9398), .C2(n10556), .A(n9397), .B(n9396), .ZN(n9463)
         );
  MUX2_X1 U10295 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n9463), .S(n10642), .Z(
        P2_U3544) );
  NAND2_X1 U10296 ( .A1(n9399), .A2(n10639), .ZN(n9403) );
  AOI22_X1 U10297 ( .A1(n9400), .A2(n10511), .B1(n10632), .B2(n8872), .ZN(
        n9401) );
  OAI211_X1 U10298 ( .C1(n9235), .C2(n9403), .A(n9402), .B(n9401), .ZN(n9464)
         );
  MUX2_X1 U10299 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n9464), .S(n10642), .Z(
        P2_U3543) );
  AOI22_X1 U10300 ( .A1(n9405), .A2(n10511), .B1(n10632), .B2(n9404), .ZN(
        n9406) );
  OAI211_X1 U10301 ( .C1(n9408), .C2(n10556), .A(n9407), .B(n9406), .ZN(n9465)
         );
  MUX2_X1 U10302 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n9465), .S(n10642), .Z(
        P2_U3542) );
  AOI22_X1 U10303 ( .A1(n9410), .A2(n10511), .B1(n10632), .B2(n9409), .ZN(
        n9411) );
  OAI211_X1 U10304 ( .C1(n9413), .C2(n10556), .A(n9412), .B(n9411), .ZN(n9466)
         );
  MUX2_X1 U10305 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n9466), .S(n10642), .Z(
        P2_U3541) );
  NAND3_X1 U10306 ( .A1(n9415), .A2(n9414), .A3(n10639), .ZN(n9420) );
  AOI22_X1 U10307 ( .A1(n9417), .A2(n10511), .B1(n10632), .B2(n9416), .ZN(
        n9418) );
  NAND3_X1 U10308 ( .A1(n9420), .A2(n9419), .A3(n9418), .ZN(n9467) );
  MUX2_X1 U10309 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n9467), .S(n10642), .Z(
        P2_U3540) );
  AOI21_X1 U10310 ( .B1(n10632), .B2(n9422), .A(n9421), .ZN(n9423) );
  OAI211_X1 U10311 ( .C1(n9425), .C2(n10556), .A(n9424), .B(n9423), .ZN(n9695)
         );
  MUX2_X1 U10312 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n9695), .S(n10642), .Z(
        P2_U3539) );
  AOI22_X1 U10313 ( .A1(n9427), .A2(n10511), .B1(n10632), .B2(n9426), .ZN(
        n9428) );
  OAI211_X1 U10314 ( .C1(n9430), .C2(n10556), .A(n9429), .B(n9428), .ZN(n9698)
         );
  MUX2_X1 U10315 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n9698), .S(n10642), .Z(
        P2_U3538) );
  AOI21_X1 U10316 ( .B1(n10632), .B2(n9432), .A(n9431), .ZN(n9433) );
  OAI211_X1 U10317 ( .C1(n9435), .C2(n10556), .A(n9434), .B(n9433), .ZN(n9699)
         );
  MUX2_X1 U10318 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n9699), .S(n10642), .Z(
        P2_U3537) );
  AOI21_X1 U10319 ( .B1(n10632), .B2(n9437), .A(n9436), .ZN(n9438) );
  OAI211_X1 U10320 ( .C1(n9440), .C2(n10556), .A(n9439), .B(n9438), .ZN(n9700)
         );
  MUX2_X1 U10321 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n9700), .S(n10642), .Z(
        P2_U3536) );
  AOI22_X1 U10322 ( .A1(n9442), .A2(n10511), .B1(n10632), .B2(n9441), .ZN(
        n9443) );
  OAI211_X1 U10323 ( .C1(n9445), .C2(n10556), .A(n9444), .B(n9443), .ZN(n9701)
         );
  MUX2_X1 U10324 ( .A(P2_REG1_REG_15__SCAN_IN), .B(n9701), .S(n10642), .Z(
        P2_U3535) );
  AOI22_X1 U10325 ( .A1(n9447), .A2(n10511), .B1(n10632), .B2(n9446), .ZN(
        n9448) );
  OAI211_X1 U10326 ( .C1(n9450), .C2(n10556), .A(n9449), .B(n9448), .ZN(n9702)
         );
  MUX2_X1 U10327 ( .A(P2_REG1_REG_14__SCAN_IN), .B(n9702), .S(n10642), .Z(
        P2_U3534) );
  AOI22_X1 U10328 ( .A1(n9452), .A2(n10511), .B1(n10632), .B2(n9451), .ZN(
        n9453) );
  OAI211_X1 U10329 ( .C1(n9455), .C2(n10556), .A(n9454), .B(n9453), .ZN(n9703)
         );
  MUX2_X1 U10330 ( .A(P2_REG1_REG_13__SCAN_IN), .B(n9703), .S(n10642), .Z(
        P2_U3533) );
  MUX2_X1 U10331 ( .A(P2_REG0_REG_31__SCAN_IN), .B(n9456), .S(n10646), .Z(
        P2_U3519) );
  MUX2_X1 U10332 ( .A(P2_REG0_REG_30__SCAN_IN), .B(n9457), .S(n10646), .Z(
        P2_U3518) );
  MUX2_X1 U10333 ( .A(P2_REG0_REG_29__SCAN_IN), .B(n9458), .S(n10646), .Z(
        P2_U3517) );
  MUX2_X1 U10334 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n9459), .S(n10646), .Z(
        P2_U3516) );
  MUX2_X1 U10335 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n9460), .S(n10646), .Z(
        P2_U3515) );
  MUX2_X1 U10336 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n9461), .S(n10646), .Z(
        P2_U3514) );
  MUX2_X1 U10337 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n9462), .S(n10646), .Z(
        P2_U3513) );
  MUX2_X1 U10338 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n9463), .S(n10646), .Z(
        P2_U3512) );
  MUX2_X1 U10339 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n9464), .S(n10646), .Z(
        P2_U3511) );
  MUX2_X1 U10340 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n9465), .S(n10646), .Z(
        P2_U3510) );
  MUX2_X1 U10341 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n9466), .S(n10646), .Z(
        P2_U3509) );
  MUX2_X1 U10342 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n9467), .S(n10646), .Z(
        P2_U3508) );
  INV_X1 U10343 ( .A(keyinput_62), .ZN(n9568) );
  INV_X1 U10344 ( .A(keyinput_53), .ZN(n9553) );
  INV_X1 U10345 ( .A(keyinput_52), .ZN(n9551) );
  INV_X1 U10346 ( .A(keyinput_51), .ZN(n9549) );
  INV_X1 U10347 ( .A(keyinput_50), .ZN(n9547) );
  INV_X1 U10348 ( .A(keyinput_49), .ZN(n9545) );
  OAI22_X1 U10349 ( .A1(n9469), .A2(keyinput_47), .B1(P2_REG3_REG_16__SCAN_IN), 
        .B2(keyinput_48), .ZN(n9468) );
  AOI221_X1 U10350 ( .B1(n9469), .B2(keyinput_47), .C1(keyinput_48), .C2(
        P2_REG3_REG_16__SCAN_IN), .A(n9468), .ZN(n9542) );
  INV_X1 U10351 ( .A(keyinput_45), .ZN(n9539) );
  AOI22_X1 U10352 ( .A1(P2_REG3_REG_23__SCAN_IN), .A2(keyinput_38), .B1(
        P2_REG3_REG_14__SCAN_IN), .B2(keyinput_37), .ZN(n9470) );
  OAI221_X1 U10353 ( .B1(P2_REG3_REG_23__SCAN_IN), .B2(keyinput_38), .C1(
        P2_REG3_REG_14__SCAN_IN), .C2(keyinput_37), .A(n9470), .ZN(n9529) );
  INV_X1 U10354 ( .A(keyinput_36), .ZN(n9527) );
  INV_X1 U10355 ( .A(keyinput_35), .ZN(n9525) );
  INV_X1 U10356 ( .A(keyinput_34), .ZN(n9523) );
  INV_X1 U10357 ( .A(SI_0_), .ZN(n9472) );
  AOI22_X1 U10358 ( .A1(SI_1_), .A2(keyinput_31), .B1(n9472), .B2(keyinput_32), 
        .ZN(n9471) );
  OAI221_X1 U10359 ( .B1(SI_1_), .B2(keyinput_31), .C1(n9472), .C2(keyinput_32), .A(n9471), .ZN(n9520) );
  AOI22_X1 U10360 ( .A1(n9584), .A2(keyinput_21), .B1(n9583), .B2(keyinput_20), 
        .ZN(n9473) );
  OAI221_X1 U10361 ( .B1(n9584), .B2(keyinput_21), .C1(n9583), .C2(keyinput_20), .A(n9473), .ZN(n9504) );
  OAI22_X1 U10362 ( .A1(n9475), .A2(keyinput_19), .B1(SI_14_), .B2(keyinput_18), .ZN(n9474) );
  AOI221_X1 U10363 ( .B1(n9475), .B2(keyinput_19), .C1(keyinput_18), .C2(
        SI_14_), .A(n9474), .ZN(n9501) );
  INV_X1 U10364 ( .A(SI_16_), .ZN(n9619) );
  INV_X1 U10365 ( .A(keyinput_16), .ZN(n9499) );
  INV_X1 U10366 ( .A(SI_17_), .ZN(n9616) );
  INV_X1 U10367 ( .A(keyinput_15), .ZN(n9497) );
  INV_X1 U10368 ( .A(keyinput_14), .ZN(n9495) );
  OAI22_X1 U10369 ( .A1(n9588), .A2(keyinput_11), .B1(n9477), .B2(keyinput_12), 
        .ZN(n9476) );
  AOI221_X1 U10370 ( .B1(n9588), .B2(keyinput_11), .C1(keyinput_12), .C2(n9477), .A(n9476), .ZN(n9491) );
  OAI22_X1 U10371 ( .A1(SI_30_), .A2(keyinput_2), .B1(SI_29_), .B2(keyinput_3), 
        .ZN(n9478) );
  AOI221_X1 U10372 ( .B1(SI_30_), .B2(keyinput_2), .C1(keyinput_3), .C2(SI_29_), .A(n9478), .ZN(n9483) );
  AOI22_X1 U10373 ( .A1(P2_WR_REG_SCAN_IN), .A2(keyinput_0), .B1(SI_31_), .B2(
        keyinput_1), .ZN(n9479) );
  OAI221_X1 U10374 ( .B1(P2_WR_REG_SCAN_IN), .B2(keyinput_0), .C1(SI_31_), 
        .C2(keyinput_1), .A(n9479), .ZN(n9482) );
  AOI22_X1 U10375 ( .A1(SI_28_), .A2(keyinput_4), .B1(SI_27_), .B2(keyinput_5), 
        .ZN(n9480) );
  OAI221_X1 U10376 ( .B1(SI_28_), .B2(keyinput_4), .C1(SI_27_), .C2(keyinput_5), .A(n9480), .ZN(n9481) );
  AOI21_X1 U10377 ( .B1(n9483), .B2(n9482), .A(n9481), .ZN(n9489) );
  XOR2_X1 U10378 ( .A(n9604), .B(keyinput_6), .Z(n9488) );
  OAI22_X1 U10379 ( .A1(n9590), .A2(keyinput_9), .B1(keyinput_8), .B2(SI_24_), 
        .ZN(n9484) );
  AOI221_X1 U10380 ( .B1(n9590), .B2(keyinput_9), .C1(SI_24_), .C2(keyinput_8), 
        .A(n9484), .ZN(n9487) );
  OAI22_X1 U10381 ( .A1(SI_25_), .A2(keyinput_7), .B1(keyinput_10), .B2(SI_22_), .ZN(n9485) );
  AOI221_X1 U10382 ( .B1(SI_25_), .B2(keyinput_7), .C1(SI_22_), .C2(
        keyinput_10), .A(n9485), .ZN(n9486) );
  OAI211_X1 U10383 ( .C1(n9489), .C2(n9488), .A(n9487), .B(n9486), .ZN(n9490)
         );
  AOI22_X1 U10384 ( .A1(keyinput_13), .A2(n9493), .B1(n9491), .B2(n9490), .ZN(
        n9492) );
  OAI21_X1 U10385 ( .B1(n9493), .B2(keyinput_13), .A(n9492), .ZN(n9494) );
  OAI221_X1 U10386 ( .B1(SI_18_), .B2(n9495), .C1(n9612), .C2(keyinput_14), 
        .A(n9494), .ZN(n9496) );
  OAI221_X1 U10387 ( .B1(SI_17_), .B2(keyinput_15), .C1(n9616), .C2(n9497), 
        .A(n9496), .ZN(n9498) );
  OAI221_X1 U10388 ( .B1(SI_16_), .B2(keyinput_16), .C1(n9619), .C2(n9499), 
        .A(n9498), .ZN(n9500) );
  OAI211_X1 U10389 ( .C1(SI_15_), .C2(keyinput_17), .A(n9501), .B(n9500), .ZN(
        n9502) );
  AOI21_X1 U10390 ( .B1(SI_15_), .B2(keyinput_17), .A(n9502), .ZN(n9503) );
  OAI22_X1 U10391 ( .A1(n9504), .A2(n9503), .B1(keyinput_22), .B2(SI_10_), 
        .ZN(n9505) );
  AOI21_X1 U10392 ( .B1(keyinput_22), .B2(SI_10_), .A(n9505), .ZN(n9513) );
  INV_X1 U10393 ( .A(SI_8_), .ZN(n9581) );
  AOI22_X1 U10394 ( .A1(n9507), .A2(keyinput_23), .B1(keyinput_24), .B2(n9581), 
        .ZN(n9506) );
  OAI221_X1 U10395 ( .B1(n9507), .B2(keyinput_23), .C1(n9581), .C2(keyinput_24), .A(n9506), .ZN(n9512) );
  INV_X1 U10396 ( .A(SI_6_), .ZN(n9509) );
  OAI22_X1 U10397 ( .A1(n9509), .A2(keyinput_26), .B1(SI_7_), .B2(keyinput_25), 
        .ZN(n9508) );
  AOI221_X1 U10398 ( .B1(n9509), .B2(keyinput_26), .C1(keyinput_25), .C2(SI_7_), .A(n9508), .ZN(n9511) );
  XOR2_X1 U10399 ( .A(n9627), .B(keyinput_27), .Z(n9510) );
  OAI211_X1 U10400 ( .C1(n9513), .C2(n9512), .A(n9511), .B(n9510), .ZN(n9517)
         );
  XOR2_X1 U10401 ( .A(SI_2_), .B(keyinput_30), .Z(n9516) );
  OR2_X1 U10402 ( .A1(SI_4_), .A2(keyinput_28), .ZN(n9515) );
  XNOR2_X1 U10403 ( .A(SI_3_), .B(keyinput_29), .ZN(n9514) );
  NAND4_X1 U10404 ( .A1(n9517), .A2(n9516), .A3(n9515), .A4(n9514), .ZN(n9518)
         );
  AOI21_X1 U10405 ( .B1(SI_4_), .B2(keyinput_28), .A(n9518), .ZN(n9519) );
  OAI22_X1 U10406 ( .A1(n9520), .A2(n9519), .B1(keyinput_33), .B2(
        P2_RD_REG_SCAN_IN), .ZN(n9521) );
  AOI21_X1 U10407 ( .B1(keyinput_33), .B2(P2_RD_REG_SCAN_IN), .A(n9521), .ZN(
        n9522) );
  AOI221_X1 U10408 ( .B1(P2_STATE_REG_SCAN_IN), .B2(n9523), .C1(P2_U3152), 
        .C2(keyinput_34), .A(n9522), .ZN(n9524) );
  AOI221_X1 U10409 ( .B1(P2_REG3_REG_7__SCAN_IN), .B2(keyinput_35), .C1(n9649), 
        .C2(n9525), .A(n9524), .ZN(n9526) );
  AOI221_X1 U10410 ( .B1(P2_REG3_REG_27__SCAN_IN), .B2(keyinput_36), .C1(n9651), .C2(n9527), .A(n9526), .ZN(n9528) );
  OAI22_X1 U10411 ( .A1(keyinput_39), .A2(n7116), .B1(n9529), .B2(n9528), .ZN(
        n9530) );
  AOI21_X1 U10412 ( .B1(keyinput_39), .B2(n7116), .A(n9530), .ZN(n9537) );
  AOI22_X1 U10413 ( .A1(n9532), .A2(keyinput_41), .B1(n9578), .B2(keyinput_40), 
        .ZN(n9531) );
  OAI221_X1 U10414 ( .B1(n9532), .B2(keyinput_41), .C1(n9578), .C2(keyinput_40), .A(n9531), .ZN(n9536) );
  OAI22_X1 U10415 ( .A1(n6990), .A2(keyinput_43), .B1(P2_REG3_REG_1__SCAN_IN), 
        .B2(keyinput_44), .ZN(n9533) );
  AOI221_X1 U10416 ( .B1(n6990), .B2(keyinput_43), .C1(keyinput_44), .C2(
        P2_REG3_REG_1__SCAN_IN), .A(n9533), .ZN(n9535) );
  XNOR2_X1 U10417 ( .A(P2_REG3_REG_28__SCAN_IN), .B(keyinput_42), .ZN(n9534)
         );
  OAI211_X1 U10418 ( .C1(n9537), .C2(n9536), .A(n9535), .B(n9534), .ZN(n9538)
         );
  OAI221_X1 U10419 ( .B1(P2_REG3_REG_21__SCAN_IN), .B2(keyinput_45), .C1(n9540), .C2(n9539), .A(n9538), .ZN(n9541) );
  OAI211_X1 U10420 ( .C1(P2_REG3_REG_12__SCAN_IN), .C2(keyinput_46), .A(n9542), 
        .B(n9541), .ZN(n9543) );
  AOI21_X1 U10421 ( .B1(P2_REG3_REG_12__SCAN_IN), .B2(keyinput_46), .A(n9543), 
        .ZN(n9544) );
  AOI221_X1 U10422 ( .B1(P2_REG3_REG_5__SCAN_IN), .B2(keyinput_49), .C1(n9668), 
        .C2(n9545), .A(n9544), .ZN(n9546) );
  AOI221_X1 U10423 ( .B1(P2_REG3_REG_17__SCAN_IN), .B2(n9547), .C1(n9671), 
        .C2(keyinput_50), .A(n9546), .ZN(n9548) );
  AOI221_X1 U10424 ( .B1(P2_REG3_REG_24__SCAN_IN), .B2(n9549), .C1(n9674), 
        .C2(keyinput_51), .A(n9548), .ZN(n9550) );
  AOI221_X1 U10425 ( .B1(P2_REG3_REG_4__SCAN_IN), .B2(n9551), .C1(n9677), .C2(
        keyinput_52), .A(n9550), .ZN(n9552) );
  AOI221_X1 U10426 ( .B1(P2_REG3_REG_9__SCAN_IN), .B2(n9553), .C1(n9679), .C2(
        keyinput_53), .A(n9552), .ZN(n9554) );
  AOI21_X1 U10427 ( .B1(P2_REG3_REG_0__SCAN_IN), .B2(keyinput_54), .A(n9554), 
        .ZN(n9559) );
  AOI22_X1 U10428 ( .A1(n9557), .A2(keyinput_55), .B1(n9556), .B2(keyinput_56), 
        .ZN(n9555) );
  OAI221_X1 U10429 ( .B1(n9557), .B2(keyinput_55), .C1(n9556), .C2(keyinput_56), .A(n9555), .ZN(n9558) );
  AOI221_X1 U10430 ( .B1(P2_REG3_REG_0__SCAN_IN), .B2(n9559), .C1(keyinput_54), 
        .C2(n9559), .A(n9558), .ZN(n9566) );
  AOI22_X1 U10431 ( .A1(P2_REG3_REG_22__SCAN_IN), .A2(keyinput_57), .B1(n9561), 
        .B2(keyinput_58), .ZN(n9560) );
  OAI221_X1 U10432 ( .B1(P2_REG3_REG_22__SCAN_IN), .B2(keyinput_57), .C1(n9561), .C2(keyinput_58), .A(n9560), .ZN(n9565) );
  OAI22_X1 U10433 ( .A1(n6381), .A2(keyinput_61), .B1(P2_REG3_REG_18__SCAN_IN), 
        .B2(keyinput_60), .ZN(n9562) );
  AOI221_X1 U10434 ( .B1(n6381), .B2(keyinput_61), .C1(keyinput_60), .C2(
        P2_REG3_REG_18__SCAN_IN), .A(n9562), .ZN(n9564) );
  XNOR2_X1 U10435 ( .A(P2_REG3_REG_2__SCAN_IN), .B(keyinput_59), .ZN(n9563) );
  OAI211_X1 U10436 ( .C1(n9566), .C2(n9565), .A(n9564), .B(n9563), .ZN(n9567)
         );
  OAI221_X1 U10437 ( .B1(P2_REG3_REG_26__SCAN_IN), .B2(keyinput_62), .C1(n9689), .C2(n9568), .A(n9567), .ZN(n9570) );
  INV_X1 U10438 ( .A(keyinput_127), .ZN(n9571) );
  AOI21_X1 U10439 ( .B1(keyinput_63), .B2(n9570), .A(n9571), .ZN(n9573) );
  INV_X1 U10440 ( .A(keyinput_63), .ZN(n9569) );
  AOI21_X1 U10441 ( .B1(n9570), .B2(n9569), .A(P2_REG3_REG_15__SCAN_IN), .ZN(
        n9572) );
  AOI22_X1 U10442 ( .A1(n9573), .A2(P2_REG3_REG_15__SCAN_IN), .B1(n9572), .B2(
        n9571), .ZN(n9694) );
  AOI22_X1 U10443 ( .A1(P2_REG3_REG_11__SCAN_IN), .A2(keyinput_122), .B1(n9575), .B2(keyinput_121), .ZN(n9574) );
  OAI221_X1 U10444 ( .B1(P2_REG3_REG_11__SCAN_IN), .B2(keyinput_122), .C1(
        n9575), .C2(keyinput_121), .A(n9574), .ZN(n9686) );
  XNOR2_X1 U10445 ( .A(P2_REG3_REG_0__SCAN_IN), .B(keyinput_118), .ZN(n9684)
         );
  INV_X1 U10446 ( .A(keyinput_117), .ZN(n9680) );
  INV_X1 U10447 ( .A(keyinput_116), .ZN(n9676) );
  INV_X1 U10448 ( .A(keyinput_115), .ZN(n9673) );
  INV_X1 U10449 ( .A(keyinput_114), .ZN(n9670) );
  INV_X1 U10450 ( .A(keyinput_113), .ZN(n9667) );
  AOI22_X1 U10451 ( .A1(P2_REG3_REG_28__SCAN_IN), .A2(keyinput_106), .B1(
        P2_REG3_REG_8__SCAN_IN), .B2(keyinput_107), .ZN(n9576) );
  OAI221_X1 U10452 ( .B1(P2_REG3_REG_28__SCAN_IN), .B2(keyinput_106), .C1(
        P2_REG3_REG_8__SCAN_IN), .C2(keyinput_107), .A(n9576), .ZN(n9660) );
  OAI22_X1 U10453 ( .A1(n9578), .A2(keyinput_104), .B1(P2_REG3_REG_19__SCAN_IN), .B2(keyinput_105), .ZN(n9577) );
  AOI221_X1 U10454 ( .B1(n9578), .B2(keyinput_104), .C1(keyinput_105), .C2(
        P2_REG3_REG_19__SCAN_IN), .A(n9577), .ZN(n9657) );
  OAI22_X1 U10455 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(keyinput_101), .B1(
        keyinput_102), .B2(P2_REG3_REG_23__SCAN_IN), .ZN(n9579) );
  AOI221_X1 U10456 ( .B1(P2_REG3_REG_14__SCAN_IN), .B2(keyinput_101), .C1(
        P2_REG3_REG_23__SCAN_IN), .C2(keyinput_102), .A(n9579), .ZN(n9654) );
  INV_X1 U10457 ( .A(keyinput_100), .ZN(n9652) );
  INV_X1 U10458 ( .A(keyinput_99), .ZN(n9648) );
  INV_X1 U10459 ( .A(keyinput_98), .ZN(n9645) );
  OAI22_X1 U10460 ( .A1(n9581), .A2(keyinput_88), .B1(SI_9_), .B2(keyinput_87), 
        .ZN(n9580) );
  AOI221_X1 U10461 ( .B1(n9581), .B2(keyinput_88), .C1(keyinput_87), .C2(SI_9_), .A(n9580), .ZN(n9633) );
  AOI22_X1 U10462 ( .A1(n9584), .A2(keyinput_85), .B1(n9583), .B2(keyinput_84), 
        .ZN(n9582) );
  OAI221_X1 U10463 ( .B1(n9584), .B2(keyinput_85), .C1(n9583), .C2(keyinput_84), .A(n9582), .ZN(n9626) );
  OAI22_X1 U10464 ( .A1(n9586), .A2(keyinput_81), .B1(keyinput_82), .B2(SI_14_), .ZN(n9585) );
  AOI221_X1 U10465 ( .B1(n9586), .B2(keyinput_81), .C1(SI_14_), .C2(
        keyinput_82), .A(n9585), .ZN(n9621) );
  INV_X1 U10466 ( .A(keyinput_80), .ZN(n9618) );
  INV_X1 U10467 ( .A(keyinput_79), .ZN(n9615) );
  INV_X1 U10468 ( .A(keyinput_78), .ZN(n9613) );
  OAI22_X1 U10469 ( .A1(n9588), .A2(keyinput_75), .B1(keyinput_76), .B2(SI_20_), .ZN(n9587) );
  AOI221_X1 U10470 ( .B1(n9588), .B2(keyinput_75), .C1(SI_20_), .C2(
        keyinput_76), .A(n9587), .ZN(n9609) );
  OAI22_X1 U10471 ( .A1(n9591), .A2(keyinput_72), .B1(n9590), .B2(keyinput_73), 
        .ZN(n9589) );
  AOI221_X1 U10472 ( .B1(n9591), .B2(keyinput_72), .C1(keyinput_73), .C2(n9590), .A(n9589), .ZN(n9607) );
  OAI22_X1 U10473 ( .A1(n9593), .A2(keyinput_74), .B1(SI_25_), .B2(keyinput_71), .ZN(n9592) );
  AOI221_X1 U10474 ( .B1(n9593), .B2(keyinput_74), .C1(keyinput_71), .C2(
        SI_25_), .A(n9592), .ZN(n9606) );
  INV_X1 U10475 ( .A(keyinput_70), .ZN(n9603) );
  OAI22_X1 U10476 ( .A1(SI_31_), .A2(keyinput_65), .B1(keyinput_64), .B2(
        P2_WR_REG_SCAN_IN), .ZN(n9594) );
  AOI221_X1 U10477 ( .B1(SI_31_), .B2(keyinput_65), .C1(P2_WR_REG_SCAN_IN), 
        .C2(keyinput_64), .A(n9594), .ZN(n9601) );
  INV_X1 U10478 ( .A(SI_30_), .ZN(n9596) );
  AOI22_X1 U10479 ( .A1(n9597), .A2(keyinput_67), .B1(n9596), .B2(keyinput_66), 
        .ZN(n9595) );
  OAI221_X1 U10480 ( .B1(n9597), .B2(keyinput_67), .C1(n9596), .C2(keyinput_66), .A(n9595), .ZN(n9600) );
  OAI22_X1 U10481 ( .A1(SI_27_), .A2(keyinput_69), .B1(SI_28_), .B2(
        keyinput_68), .ZN(n9598) );
  AOI221_X1 U10482 ( .B1(SI_27_), .B2(keyinput_69), .C1(keyinput_68), .C2(
        SI_28_), .A(n9598), .ZN(n9599) );
  OAI21_X1 U10483 ( .B1(n9601), .B2(n9600), .A(n9599), .ZN(n9602) );
  OAI221_X1 U10484 ( .B1(SI_26_), .B2(keyinput_70), .C1(n9604), .C2(n9603), 
        .A(n9602), .ZN(n9605) );
  NAND3_X1 U10485 ( .A1(n9607), .A2(n9606), .A3(n9605), .ZN(n9608) );
  AOI22_X1 U10486 ( .A1(n9609), .A2(n9608), .B1(keyinput_77), .B2(SI_19_), 
        .ZN(n9610) );
  OAI21_X1 U10487 ( .B1(keyinput_77), .B2(SI_19_), .A(n9610), .ZN(n9611) );
  OAI221_X1 U10488 ( .B1(SI_18_), .B2(n9613), .C1(n9612), .C2(keyinput_78), 
        .A(n9611), .ZN(n9614) );
  OAI221_X1 U10489 ( .B1(SI_17_), .B2(keyinput_79), .C1(n9616), .C2(n9615), 
        .A(n9614), .ZN(n9617) );
  OAI221_X1 U10490 ( .B1(SI_16_), .B2(keyinput_80), .C1(n9619), .C2(n9618), 
        .A(n9617), .ZN(n9620) );
  OAI211_X1 U10491 ( .C1(SI_13_), .C2(keyinput_83), .A(n9621), .B(n9620), .ZN(
        n9622) );
  AOI21_X1 U10492 ( .B1(SI_13_), .B2(keyinput_83), .A(n9622), .ZN(n9625) );
  NAND2_X1 U10493 ( .A1(n9624), .A2(keyinput_86), .ZN(n9623) );
  OAI221_X1 U10494 ( .B1(n9626), .B2(n9625), .C1(n9624), .C2(keyinput_86), .A(
        n9623), .ZN(n9632) );
  XOR2_X1 U10495 ( .A(n9627), .B(keyinput_91), .Z(n9631) );
  INV_X1 U10496 ( .A(SI_7_), .ZN(n9629) );
  AOI22_X1 U10497 ( .A1(SI_6_), .A2(keyinput_90), .B1(n9629), .B2(keyinput_89), 
        .ZN(n9628) );
  OAI221_X1 U10498 ( .B1(SI_6_), .B2(keyinput_90), .C1(n9629), .C2(keyinput_89), .A(n9628), .ZN(n9630) );
  AOI211_X1 U10499 ( .C1(n9633), .C2(n9632), .A(n9631), .B(n9630), .ZN(n9637)
         );
  XOR2_X1 U10500 ( .A(SI_2_), .B(keyinput_94), .Z(n9636) );
  XNOR2_X1 U10501 ( .A(SI_3_), .B(keyinput_93), .ZN(n9635) );
  XNOR2_X1 U10502 ( .A(SI_4_), .B(keyinput_92), .ZN(n9634) );
  NOR4_X1 U10503 ( .A1(n9637), .A2(n9636), .A3(n9635), .A4(n9634), .ZN(n9641)
         );
  XNOR2_X1 U10504 ( .A(n9638), .B(keyinput_95), .ZN(n9640) );
  XNOR2_X1 U10505 ( .A(SI_0_), .B(keyinput_96), .ZN(n9639) );
  NOR3_X1 U10506 ( .A1(n9641), .A2(n9640), .A3(n9639), .ZN(n9642) );
  AOI21_X1 U10507 ( .B1(keyinput_97), .B2(n4918), .A(n9642), .ZN(n9643) );
  OAI21_X1 U10508 ( .B1(n4918), .B2(keyinput_97), .A(n9643), .ZN(n9644) );
  OAI221_X1 U10509 ( .B1(P2_STATE_REG_SCAN_IN), .B2(keyinput_98), .C1(P2_U3152), .C2(n9645), .A(n9644), .ZN(n9647) );
  OAI221_X1 U10510 ( .B1(P2_REG3_REG_7__SCAN_IN), .B2(keyinput_99), .C1(n9649), 
        .C2(n9648), .A(n9647), .ZN(n9650) );
  OAI221_X1 U10511 ( .B1(P2_REG3_REG_27__SCAN_IN), .B2(n9652), .C1(n9651), 
        .C2(keyinput_100), .A(n9650), .ZN(n9653) );
  AOI22_X1 U10512 ( .A1(n9654), .A2(n9653), .B1(keyinput_103), .B2(
        P2_REG3_REG_10__SCAN_IN), .ZN(n9655) );
  OAI21_X1 U10513 ( .B1(keyinput_103), .B2(P2_REG3_REG_10__SCAN_IN), .A(n9655), 
        .ZN(n9656) );
  AOI22_X1 U10514 ( .A1(n9657), .A2(n9656), .B1(P2_REG3_REG_1__SCAN_IN), .B2(
        keyinput_108), .ZN(n9658) );
  OAI21_X1 U10515 ( .B1(P2_REG3_REG_1__SCAN_IN), .B2(keyinput_108), .A(n9658), 
        .ZN(n9659) );
  OAI22_X1 U10516 ( .A1(n9660), .A2(n9659), .B1(keyinput_109), .B2(
        P2_REG3_REG_21__SCAN_IN), .ZN(n9661) );
  AOI21_X1 U10517 ( .B1(keyinput_109), .B2(P2_REG3_REG_21__SCAN_IN), .A(n9661), 
        .ZN(n9664) );
  AOI22_X1 U10518 ( .A1(n7304), .A2(keyinput_110), .B1(keyinput_112), .B2(
        n7792), .ZN(n9662) );
  OAI221_X1 U10519 ( .B1(n7304), .B2(keyinput_110), .C1(n7792), .C2(
        keyinput_112), .A(n9662), .ZN(n9663) );
  AOI211_X1 U10520 ( .C1(P2_REG3_REG_25__SCAN_IN), .C2(keyinput_111), .A(n9664), .B(n9663), .ZN(n9665) );
  OAI21_X1 U10521 ( .B1(P2_REG3_REG_25__SCAN_IN), .B2(keyinput_111), .A(n9665), 
        .ZN(n9666) );
  OAI221_X1 U10522 ( .B1(P2_REG3_REG_5__SCAN_IN), .B2(keyinput_113), .C1(n9668), .C2(n9667), .A(n9666), .ZN(n9669) );
  OAI221_X1 U10523 ( .B1(P2_REG3_REG_17__SCAN_IN), .B2(keyinput_114), .C1(
        n9671), .C2(n9670), .A(n9669), .ZN(n9672) );
  OAI221_X1 U10524 ( .B1(P2_REG3_REG_24__SCAN_IN), .B2(keyinput_115), .C1(
        n9674), .C2(n9673), .A(n9672), .ZN(n9675) );
  OAI221_X1 U10525 ( .B1(P2_REG3_REG_4__SCAN_IN), .B2(keyinput_116), .C1(n9677), .C2(n9676), .A(n9675), .ZN(n9678) );
  OAI221_X1 U10526 ( .B1(P2_REG3_REG_9__SCAN_IN), .B2(n9680), .C1(n9679), .C2(
        keyinput_117), .A(n9678), .ZN(n9683) );
  AOI22_X1 U10527 ( .A1(P2_REG3_REG_20__SCAN_IN), .A2(keyinput_119), .B1(
        P2_REG3_REG_13__SCAN_IN), .B2(keyinput_120), .ZN(n9681) );
  OAI221_X1 U10528 ( .B1(P2_REG3_REG_20__SCAN_IN), .B2(keyinput_119), .C1(
        P2_REG3_REG_13__SCAN_IN), .C2(keyinput_120), .A(n9681), .ZN(n9682) );
  AOI21_X1 U10529 ( .B1(n9684), .B2(n9683), .A(n9682), .ZN(n9685) );
  OAI22_X1 U10530 ( .A1(n9686), .A2(n9685), .B1(n6381), .B2(keyinput_125), 
        .ZN(n9687) );
  AOI21_X1 U10531 ( .B1(n6381), .B2(keyinput_125), .A(n9687), .ZN(n9692) );
  OAI22_X1 U10532 ( .A1(P2_REG3_REG_18__SCAN_IN), .A2(keyinput_124), .B1(
        P2_REG3_REG_2__SCAN_IN), .B2(keyinput_123), .ZN(n9688) );
  AOI221_X1 U10533 ( .B1(P2_REG3_REG_18__SCAN_IN), .B2(keyinput_124), .C1(
        keyinput_123), .C2(P2_REG3_REG_2__SCAN_IN), .A(n9688), .ZN(n9691) );
  XNOR2_X1 U10534 ( .A(n9689), .B(keyinput_126), .ZN(n9690) );
  AOI21_X1 U10535 ( .B1(n9692), .B2(n9691), .A(n9690), .ZN(n9693) );
  NOR2_X1 U10536 ( .A1(n9694), .A2(n9693), .ZN(n9697) );
  MUX2_X1 U10537 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n9695), .S(n10646), .Z(
        n9696) );
  XOR2_X1 U10538 ( .A(n9697), .B(n9696), .Z(P2_U3507) );
  MUX2_X1 U10539 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n9698), .S(n10646), .Z(
        P2_U3505) );
  MUX2_X1 U10540 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n9699), .S(n10646), .Z(
        P2_U3502) );
  MUX2_X1 U10541 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n9700), .S(n10646), .Z(
        P2_U3499) );
  MUX2_X1 U10542 ( .A(P2_REG0_REG_15__SCAN_IN), .B(n9701), .S(n10646), .Z(
        P2_U3496) );
  MUX2_X1 U10543 ( .A(P2_REG0_REG_14__SCAN_IN), .B(n9702), .S(n10646), .Z(
        P2_U3493) );
  MUX2_X1 U10544 ( .A(P2_REG0_REG_13__SCAN_IN), .B(n9703), .S(n10646), .Z(
        P2_U3490) );
  NAND2_X1 U10545 ( .A1(n9704), .A2(n9705), .ZN(n9709) );
  INV_X1 U10546 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n9707) );
  NAND4_X1 U10547 ( .A1(n6376), .A2(P2_STATE_REG_SCAN_IN), .A3(
        P2_IR_REG_31__SCAN_IN), .A4(n9707), .ZN(n9708) );
  OAI211_X1 U10548 ( .C1(n9711), .C2(n9710), .A(n9709), .B(n9708), .ZN(
        P2_U3327) );
  MUX2_X1 U10549 ( .A(n9712), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3358) );
  XNOR2_X1 U10550 ( .A(n9714), .B(n9713), .ZN(n9715) );
  XNOR2_X1 U10551 ( .A(n9716), .B(n9715), .ZN(n9724) );
  NOR2_X1 U10552 ( .A1(n9717), .A2(n9846), .ZN(n9721) );
  AOI22_X1 U10553 ( .A1(n9718), .A2(n9783), .B1(P1_REG3_REG_27__SCAN_IN), .B2(
        P1_U3084), .ZN(n9719) );
  OAI21_X1 U10554 ( .B1(n9786), .B2(n9860), .A(n9719), .ZN(n9720) );
  AOI211_X1 U10555 ( .C1(n9722), .C2(n9837), .A(n9721), .B(n9720), .ZN(n9723)
         );
  OAI21_X1 U10556 ( .B1(n9724), .B2(n9853), .A(n9723), .ZN(P1_U3212) );
  INV_X1 U10557 ( .A(n9725), .ZN(n9730) );
  AOI21_X1 U10558 ( .B1(n9727), .B2(n9729), .A(n9726), .ZN(n9728) );
  AOI21_X1 U10559 ( .B1(n9730), .B2(n9729), .A(n9728), .ZN(n9735) );
  NAND2_X1 U10560 ( .A1(n10026), .A2(n9863), .ZN(n9732) );
  AOI22_X1 U10561 ( .A1(n10071), .A2(n9848), .B1(P1_REG3_REG_23__SCAN_IN), 
        .B2(P1_U3084), .ZN(n9731) );
  OAI211_X1 U10562 ( .C1(n9858), .C2(n10018), .A(n9732), .B(n9731), .ZN(n9733)
         );
  AOI21_X1 U10563 ( .B1(n10197), .B2(n9851), .A(n9733), .ZN(n9734) );
  OAI21_X1 U10564 ( .B1(n9735), .B2(n9853), .A(n9734), .ZN(P1_U3214) );
  XNOR2_X1 U10565 ( .A(n9736), .B(n9738), .ZN(n9739) );
  NAND2_X1 U10566 ( .A1(n9739), .A2(n9855), .ZN(n9745) );
  AOI22_X1 U10567 ( .A1(n9848), .A2(n9882), .B1(n9837), .B2(n9740), .ZN(n9744)
         );
  AOI21_X1 U10568 ( .B1(n9863), .B2(n9881), .A(n9741), .ZN(n9743) );
  NAND2_X1 U10569 ( .A1(n9783), .A2(n6618), .ZN(n9742) );
  NAND4_X1 U10570 ( .A1(n9745), .A2(n9744), .A3(n9743), .A4(n9742), .ZN(
        P1_U3216) );
  NAND2_X1 U10571 ( .A1(n9748), .A2(n9747), .ZN(n9749) );
  XNOR2_X1 U10572 ( .A(n9746), .B(n9749), .ZN(n9754) );
  NAND2_X1 U10573 ( .A1(n9848), .A2(n10142), .ZN(n9750) );
  NAND2_X1 U10574 ( .A1(P1_U3084), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n9949) );
  OAI211_X1 U10575 ( .C1(n10104), .C2(n9846), .A(n9750), .B(n9949), .ZN(n9752)
         );
  INV_X1 U10576 ( .A(n10109), .ZN(n10301) );
  NOR2_X1 U10577 ( .A1(n10301), .A2(n9866), .ZN(n9751) );
  AOI211_X1 U10578 ( .C1(n10112), .C2(n9783), .A(n9752), .B(n9751), .ZN(n9753)
         );
  OAI21_X1 U10579 ( .B1(n9754), .B2(n9853), .A(n9753), .ZN(P1_U3217) );
  NOR2_X1 U10580 ( .A1(n5216), .A2(n9757), .ZN(n9758) );
  XNOR2_X1 U10581 ( .A(n9755), .B(n9758), .ZN(n9763) );
  AOI22_X1 U10582 ( .A1(n10071), .A2(n9863), .B1(P1_REG3_REG_21__SCAN_IN), 
        .B2(P1_U3084), .ZN(n9760) );
  NAND2_X1 U10583 ( .A1(n9783), .A2(n10076), .ZN(n9759) );
  OAI211_X1 U10584 ( .C1(n10104), .C2(n9860), .A(n9760), .B(n9759), .ZN(n9761)
         );
  AOI21_X1 U10585 ( .B1(n10075), .B2(n9851), .A(n9761), .ZN(n9762) );
  OAI21_X1 U10586 ( .B1(n9763), .B2(n9853), .A(n9762), .ZN(P1_U3221) );
  NAND2_X1 U10587 ( .A1(n9765), .A2(n9764), .ZN(n9769) );
  NAND2_X1 U10588 ( .A1(n9767), .A2(n9766), .ZN(n9768) );
  XOR2_X1 U10589 ( .A(n9769), .B(n9768), .Z(n9777) );
  NOR2_X1 U10590 ( .A1(n9860), .A2(n9770), .ZN(n9771) );
  AOI211_X1 U10591 ( .C1(n9863), .C2(n9875), .A(n9772), .B(n9771), .ZN(n9773)
         );
  OAI21_X1 U10592 ( .B1(n9858), .B2(n9774), .A(n9773), .ZN(n9775) );
  AOI21_X1 U10593 ( .B1(n10263), .B2(n9837), .A(n9775), .ZN(n9776) );
  OAI21_X1 U10594 ( .B1(n9777), .B2(n9853), .A(n9776), .ZN(P1_U3222) );
  INV_X1 U10595 ( .A(n9779), .ZN(n9781) );
  NAND2_X1 U10596 ( .A1(n9781), .A2(n9780), .ZN(n9782) );
  XNOR2_X1 U10597 ( .A(n9778), .B(n9782), .ZN(n9789) );
  AOI22_X1 U10598 ( .A1(n10026), .A2(n9848), .B1(P1_REG3_REG_25__SCAN_IN), 
        .B2(P1_U3084), .ZN(n9785) );
  NAND2_X1 U10599 ( .A1(n9980), .A2(n9783), .ZN(n9784) );
  OAI211_X1 U10600 ( .C1(n9786), .C2(n9846), .A(n9785), .B(n9784), .ZN(n9787)
         );
  AOI21_X1 U10601 ( .B1(n10189), .B2(n9851), .A(n9787), .ZN(n9788) );
  OAI21_X1 U10602 ( .B1(n9789), .B2(n9853), .A(n9788), .ZN(P1_U3223) );
  INV_X1 U10603 ( .A(n9791), .ZN(n9792) );
  AOI21_X1 U10604 ( .B1(n9790), .B2(n9793), .A(n9792), .ZN(n9801) );
  OAI21_X1 U10605 ( .B1(n9795), .B2(n9846), .A(n9794), .ZN(n9796) );
  AOI21_X1 U10606 ( .B1(n9848), .B2(n9873), .A(n9796), .ZN(n9797) );
  OAI21_X1 U10607 ( .B1(n9858), .B2(n9798), .A(n9797), .ZN(n9799) );
  AOI21_X1 U10608 ( .B1(n10237), .B2(n9837), .A(n9799), .ZN(n9800) );
  OAI21_X1 U10609 ( .B1(n9801), .B2(n9853), .A(n9800), .ZN(P1_U3224) );
  OAI21_X1 U10610 ( .B1(n9804), .B2(n9803), .A(n9802), .ZN(n9805) );
  NAND2_X1 U10611 ( .A1(n9805), .A2(n9855), .ZN(n9810) );
  OAI21_X1 U10612 ( .B1(n9846), .B2(n10102), .A(n9806), .ZN(n9808) );
  NOR2_X1 U10613 ( .A1(n9858), .A2(n10146), .ZN(n9807) );
  AOI211_X1 U10614 ( .C1(n9848), .C2(n10144), .A(n9808), .B(n9807), .ZN(n9809)
         );
  OAI211_X1 U10615 ( .C1(n10306), .C2(n9866), .A(n9810), .B(n9809), .ZN(
        P1_U3226) );
  OAI21_X1 U10616 ( .B1(n9813), .B2(n9812), .A(n9811), .ZN(n9814) );
  NAND2_X1 U10617 ( .A1(n9814), .A2(n9855), .ZN(n9820) );
  NOR2_X1 U10618 ( .A1(n10008), .A2(n9858), .ZN(n9818) );
  NAND2_X1 U10619 ( .A1(n10043), .A2(n9848), .ZN(n9815) );
  OAI21_X1 U10620 ( .B1(P1_STATE_REG_SCAN_IN), .B2(n9816), .A(n9815), .ZN(
        n9817) );
  AOI211_X1 U10621 ( .C1(n9872), .C2(n9863), .A(n9818), .B(n9817), .ZN(n9819)
         );
  OAI211_X1 U10622 ( .C1(n10287), .C2(n9866), .A(n9820), .B(n9819), .ZN(
        P1_U3227) );
  XNOR2_X1 U10623 ( .A(n9823), .B(n9822), .ZN(n9824) );
  XNOR2_X1 U10624 ( .A(n9821), .B(n9824), .ZN(n9829) );
  AOI22_X1 U10625 ( .A1(n10094), .A2(n9863), .B1(P1_REG3_REG_20__SCAN_IN), 
        .B2(P1_U3084), .ZN(n9826) );
  NAND2_X1 U10626 ( .A1(n9848), .A2(n10125), .ZN(n9825) );
  OAI211_X1 U10627 ( .C1(n9858), .C2(n10086), .A(n9826), .B(n9825), .ZN(n9827)
         );
  AOI21_X1 U10628 ( .B1(n10213), .B2(n9837), .A(n9827), .ZN(n9828) );
  OAI21_X1 U10629 ( .B1(n9829), .B2(n9853), .A(n9828), .ZN(P1_U3231) );
  AOI21_X1 U10630 ( .B1(n9833), .B2(n9831), .A(n9830), .ZN(n9832) );
  AOI21_X1 U10631 ( .B1(n4882), .B2(n9833), .A(n9832), .ZN(n9839) );
  AOI22_X1 U10632 ( .A1(n10094), .A2(n9848), .B1(P1_REG3_REG_22__SCAN_IN), 
        .B2(P1_U3084), .ZN(n9835) );
  NAND2_X1 U10633 ( .A1(n10043), .A2(n9863), .ZN(n9834) );
  OAI211_X1 U10634 ( .C1(n9858), .C2(n10049), .A(n9835), .B(n9834), .ZN(n9836)
         );
  AOI21_X1 U10635 ( .B1(n10205), .B2(n9837), .A(n9836), .ZN(n9838) );
  OAI21_X1 U10636 ( .B1(n9839), .B2(n9853), .A(n9838), .ZN(P1_U3233) );
  NAND2_X1 U10637 ( .A1(n9840), .A2(n9841), .ZN(n9843) );
  XNOR2_X1 U10638 ( .A(n9843), .B(n9842), .ZN(n9854) );
  OAI21_X1 U10639 ( .B1(n9846), .B2(n9845), .A(n9844), .ZN(n9847) );
  AOI21_X1 U10640 ( .B1(n9848), .B2(n10126), .A(n9847), .ZN(n9849) );
  OAI21_X1 U10641 ( .B1(n9858), .B2(n10130), .A(n9849), .ZN(n9850) );
  AOI21_X1 U10642 ( .B1(n10133), .B2(n9851), .A(n9850), .ZN(n9852) );
  OAI21_X1 U10643 ( .B1(n9854), .B2(n9853), .A(n9852), .ZN(P1_U3236) );
  INV_X1 U10644 ( .A(n10182), .ZN(n9969) );
  NOR2_X1 U10645 ( .A1(n9966), .A2(n9858), .ZN(n9862) );
  OAI22_X1 U10646 ( .A1(n10001), .A2(n9860), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9859), .ZN(n9861) );
  AOI211_X1 U10647 ( .C1(n9871), .C2(n9863), .A(n9862), .B(n9861), .ZN(n9864)
         );
  OAI211_X1 U10648 ( .C1(n9969), .C2(n9866), .A(n9865), .B(n9864), .ZN(
        P1_U3238) );
  MUX2_X1 U10649 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(n9867), .S(P1_U4006), .Z(
        P1_U3586) );
  MUX2_X1 U10650 ( .A(n9868), .B(P1_DATAO_REG_30__SCAN_IN), .S(n9883), .Z(
        P1_U3585) );
  MUX2_X1 U10651 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n9869), .S(P1_U4006), .Z(
        P1_U3584) );
  MUX2_X1 U10652 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n9870), .S(P1_U4006), .Z(
        P1_U3583) );
  MUX2_X1 U10653 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n9871), .S(P1_U4006), .Z(
        P1_U3582) );
  MUX2_X1 U10654 ( .A(n9988), .B(P1_DATAO_REG_26__SCAN_IN), .S(n9883), .Z(
        P1_U3581) );
  MUX2_X1 U10655 ( .A(n9872), .B(P1_DATAO_REG_25__SCAN_IN), .S(n9883), .Z(
        P1_U3580) );
  MUX2_X1 U10656 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n10043), .S(P1_U4006), .Z(
        P1_U3578) );
  MUX2_X1 U10657 ( .A(n10071), .B(P1_DATAO_REG_22__SCAN_IN), .S(n9883), .Z(
        P1_U3577) );
  MUX2_X1 U10658 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n10094), .S(P1_U4006), .Z(
        P1_U3576) );
  MUX2_X1 U10659 ( .A(n10070), .B(P1_DATAO_REG_20__SCAN_IN), .S(n9883), .Z(
        P1_U3575) );
  MUX2_X1 U10660 ( .A(n10125), .B(P1_DATAO_REG_19__SCAN_IN), .S(n9883), .Z(
        P1_U3574) );
  MUX2_X1 U10661 ( .A(n10142), .B(P1_DATAO_REG_18__SCAN_IN), .S(n9883), .Z(
        P1_U3573) );
  MUX2_X1 U10662 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n10126), .S(P1_U4006), .Z(
        P1_U3572) );
  MUX2_X1 U10663 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n10144), .S(P1_U4006), .Z(
        P1_U3571) );
  MUX2_X1 U10664 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n9873), .S(P1_U4006), .Z(
        P1_U3570) );
  MUX2_X1 U10665 ( .A(n9874), .B(P1_DATAO_REG_14__SCAN_IN), .S(n9883), .Z(
        P1_U3569) );
  MUX2_X1 U10666 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n9875), .S(P1_U4006), .Z(
        P1_U3568) );
  MUX2_X1 U10667 ( .A(n9876), .B(P1_DATAO_REG_12__SCAN_IN), .S(n9883), .Z(
        P1_U3567) );
  MUX2_X1 U10668 ( .A(n9877), .B(P1_DATAO_REG_11__SCAN_IN), .S(n9883), .Z(
        P1_U3566) );
  MUX2_X1 U10669 ( .A(n9878), .B(P1_DATAO_REG_10__SCAN_IN), .S(n9883), .Z(
        P1_U3565) );
  MUX2_X1 U10670 ( .A(n9879), .B(P1_DATAO_REG_9__SCAN_IN), .S(n9883), .Z(
        P1_U3564) );
  MUX2_X1 U10671 ( .A(n9880), .B(P1_DATAO_REG_5__SCAN_IN), .S(n9883), .Z(
        P1_U3560) );
  MUX2_X1 U10672 ( .A(n9881), .B(P1_DATAO_REG_4__SCAN_IN), .S(n9883), .Z(
        P1_U3559) );
  MUX2_X1 U10673 ( .A(n9882), .B(P1_DATAO_REG_2__SCAN_IN), .S(n9883), .Z(
        P1_U3557) );
  MUX2_X1 U10674 ( .A(n6277), .B(P1_DATAO_REG_1__SCAN_IN), .S(n9883), .Z(
        P1_U3556) );
  OAI21_X1 U10675 ( .B1(n9886), .B2(n9885), .A(n9884), .ZN(n9890) );
  NOR2_X1 U10676 ( .A1(n10425), .A2(n9887), .ZN(n9888) );
  AOI211_X1 U10677 ( .C1(n10443), .C2(n9890), .A(n9889), .B(n9888), .ZN(n9897)
         );
  OAI21_X1 U10678 ( .B1(n9893), .B2(n9892), .A(n9891), .ZN(n9894) );
  AOI22_X1 U10679 ( .A1(n9895), .A2(n10459), .B1(n9955), .B2(n9894), .ZN(n9896) );
  NAND3_X1 U10680 ( .A1(n9898), .A2(n9897), .A3(n9896), .ZN(P1_U3245) );
  OAI21_X1 U10681 ( .B1(n9901), .B2(n9900), .A(n9899), .ZN(n9902) );
  NAND2_X1 U10682 ( .A1(n9902), .A2(n10443), .ZN(n9912) );
  AOI21_X1 U10683 ( .B1(n10457), .B2(P1_ADDR_REG_7__SCAN_IN), .A(n9903), .ZN(
        n9911) );
  OAI21_X1 U10684 ( .B1(n9906), .B2(n9905), .A(n9904), .ZN(n9907) );
  NAND2_X1 U10685 ( .A1(n9907), .A2(n9955), .ZN(n9910) );
  NAND2_X1 U10686 ( .A1(n10459), .A2(n9908), .ZN(n9909) );
  NAND4_X1 U10687 ( .A1(n9912), .A2(n9911), .A3(n9910), .A4(n9909), .ZN(
        P1_U3248) );
  OAI21_X1 U10688 ( .B1(n9915), .B2(n9914), .A(n9913), .ZN(n9916) );
  NAND2_X1 U10689 ( .A1(n9916), .A2(n10443), .ZN(n9926) );
  AOI21_X1 U10690 ( .B1(n10457), .B2(P1_ADDR_REG_8__SCAN_IN), .A(n9917), .ZN(
        n9925) );
  OAI21_X1 U10691 ( .B1(n9920), .B2(n9919), .A(n9918), .ZN(n9921) );
  NAND2_X1 U10692 ( .A1(n9921), .A2(n9955), .ZN(n9924) );
  NAND2_X1 U10693 ( .A1(n10459), .A2(n9922), .ZN(n9923) );
  NAND4_X1 U10694 ( .A1(n9926), .A2(n9925), .A3(n9924), .A4(n9923), .ZN(
        P1_U3249) );
  OAI21_X1 U10695 ( .B1(n9929), .B2(n9928), .A(n9927), .ZN(n9930) );
  NAND2_X1 U10696 ( .A1(n9930), .A2(n10443), .ZN(n9939) );
  AOI211_X1 U10697 ( .C1(n9933), .C2(n9932), .A(n9931), .B(n10451), .ZN(n9934)
         );
  AOI21_X1 U10698 ( .B1(n10459), .B2(n9935), .A(n9934), .ZN(n9937) );
  NAND2_X1 U10699 ( .A1(n10457), .A2(P1_ADDR_REG_10__SCAN_IN), .ZN(n9936) );
  NAND4_X1 U10700 ( .A1(n9939), .A2(n9938), .A3(n9937), .A4(n9936), .ZN(
        P1_U3251) );
  INV_X1 U10701 ( .A(n9940), .ZN(n9941) );
  NAND2_X1 U10702 ( .A1(n9942), .A2(n9941), .ZN(n9944) );
  INV_X1 U10703 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n10221) );
  XNOR2_X1 U10704 ( .A(n9951), .B(n10221), .ZN(n9943) );
  XNOR2_X1 U10705 ( .A(n9944), .B(n9943), .ZN(n9957) );
  AOI21_X1 U10706 ( .B1(n9946), .B2(P1_REG2_REG_18__SCAN_IN), .A(n9945), .ZN(
        n9948) );
  MUX2_X1 U10707 ( .A(n5422), .B(P1_REG2_REG_19__SCAN_IN), .S(n9951), .Z(n9947) );
  XNOR2_X1 U10708 ( .A(n9948), .B(n9947), .ZN(n9954) );
  NAND2_X1 U10709 ( .A1(n10457), .A2(P1_ADDR_REG_19__SCAN_IN), .ZN(n9950) );
  OAI211_X1 U10710 ( .C1(n9952), .C2(n9951), .A(n9950), .B(n9949), .ZN(n9953)
         );
  AOI21_X1 U10711 ( .B1(n9955), .B2(n9954), .A(n9953), .ZN(n9956) );
  OAI21_X1 U10712 ( .B1(n10447), .B2(n9957), .A(n9956), .ZN(P1_U3260) );
  OR2_X1 U10713 ( .A1(n10279), .A2(n9958), .ZN(n10163) );
  NAND3_X1 U10714 ( .A1(n10163), .A2(n10162), .A3(n10097), .ZN(n9961) );
  AOI21_X1 U10715 ( .B1(n10088), .B2(P1_REG2_REG_30__SCAN_IN), .A(n9959), .ZN(
        n9960) );
  OAI211_X1 U10716 ( .C1(n10279), .C2(n10115), .A(n9961), .B(n9960), .ZN(
        P1_U3262) );
  XNOR2_X1 U10717 ( .A(n9962), .B(n9970), .ZN(n10186) );
  INV_X1 U10718 ( .A(n9964), .ZN(n9965) );
  AOI21_X1 U10719 ( .B1(n10182), .B2(n9979), .A(n9965), .ZN(n10183) );
  INV_X1 U10720 ( .A(n9966), .ZN(n9967) );
  AOI22_X1 U10721 ( .A1(n9967), .A2(n10111), .B1(P1_REG2_REG_26__SCAN_IN), 
        .B2(n10088), .ZN(n9968) );
  OAI21_X1 U10722 ( .B1(n9969), .B2(n10115), .A(n9968), .ZN(n9976) );
  AOI21_X1 U10723 ( .B1(n4884), .B2(n5099), .A(n9997), .ZN(n9974) );
  OAI22_X1 U10724 ( .A1(n9971), .A2(n10103), .B1(n10001), .B2(n10101), .ZN(
        n9972) );
  AOI21_X1 U10725 ( .B1(n9974), .B2(n9973), .A(n9972), .ZN(n10185) );
  NOR2_X1 U10726 ( .A1(n10185), .A2(n10088), .ZN(n9975) );
  AOI211_X1 U10727 ( .C1(n10097), .C2(n10183), .A(n9976), .B(n9975), .ZN(n9977) );
  OAI21_X1 U10728 ( .B1(n10186), .B2(n10137), .A(n9977), .ZN(P1_U3265) );
  XNOR2_X1 U10729 ( .A(n9978), .B(n9987), .ZN(n10191) );
  AOI22_X1 U10730 ( .A1(n10189), .A2(n10156), .B1(P1_REG2_REG_25__SCAN_IN), 
        .B2(n10088), .ZN(n9993) );
  AOI211_X1 U10731 ( .C1(n10189), .C2(n10004), .A(n10591), .B(n9963), .ZN(
        n10188) );
  INV_X1 U10732 ( .A(n10188), .ZN(n9982) );
  INV_X1 U10733 ( .A(n9980), .ZN(n9981) );
  OAI22_X1 U10734 ( .A1(n9982), .A2(n10019), .B1(n10145), .B2(n9981), .ZN(
        n9991) );
  AOI21_X1 U10735 ( .B1(n9984), .B2(n9983), .A(n9997), .ZN(n9985) );
  OAI211_X1 U10736 ( .C1(n9999), .C2(n9987), .A(n9986), .B(n9985), .ZN(n9990)
         );
  AOI22_X1 U10737 ( .A1(n9988), .A2(n10141), .B1(n10143), .B2(n10026), .ZN(
        n9989) );
  NAND2_X1 U10738 ( .A1(n9990), .A2(n9989), .ZN(n10187) );
  OAI21_X1 U10739 ( .B1(n9991), .B2(n10187), .A(n10148), .ZN(n9992) );
  OAI211_X1 U10740 ( .C1(n10191), .C2(n10137), .A(n9993), .B(n9992), .ZN(
        P1_U3266) );
  XOR2_X1 U10741 ( .A(n9995), .B(n9994), .Z(n10194) );
  INV_X1 U10742 ( .A(n10194), .ZN(n10014) );
  NAND2_X1 U10743 ( .A1(n9996), .A2(n9995), .ZN(n9998) );
  AOI21_X1 U10744 ( .B1(n9999), .B2(n9998), .A(n9997), .ZN(n10003) );
  OAI22_X1 U10745 ( .A1(n10001), .A2(n10103), .B1(n10000), .B2(n10101), .ZN(
        n10002) );
  OR2_X1 U10746 ( .A1(n10003), .A2(n10002), .ZN(n10192) );
  INV_X1 U10747 ( .A(n10017), .ZN(n10006) );
  INV_X1 U10748 ( .A(n10004), .ZN(n10005) );
  AOI211_X1 U10749 ( .C1(n10007), .C2(n10006), .A(n10591), .B(n10005), .ZN(
        n10193) );
  NAND2_X1 U10750 ( .A1(n10193), .A2(n10110), .ZN(n10011) );
  INV_X1 U10751 ( .A(n10008), .ZN(n10009) );
  AOI22_X1 U10752 ( .A1(n10009), .A2(n10111), .B1(P1_REG2_REG_24__SCAN_IN), 
        .B2(n10088), .ZN(n10010) );
  OAI211_X1 U10753 ( .C1(n10287), .C2(n10115), .A(n10011), .B(n10010), .ZN(
        n10012) );
  AOI21_X1 U10754 ( .B1(n10148), .B2(n10192), .A(n10012), .ZN(n10013) );
  OAI21_X1 U10755 ( .B1(n10014), .B2(n10137), .A(n10013), .ZN(P1_U3267) );
  XNOR2_X1 U10756 ( .A(n10015), .B(n10016), .ZN(n10200) );
  INV_X1 U10757 ( .A(n10200), .ZN(n10032) );
  AOI22_X1 U10758 ( .A1(n10197), .A2(n10156), .B1(P1_REG2_REG_23__SCAN_IN), 
        .B2(n10088), .ZN(n10031) );
  AOI211_X1 U10759 ( .C1(n10197), .C2(n10047), .A(n10591), .B(n10017), .ZN(
        n10199) );
  INV_X1 U10760 ( .A(n10199), .ZN(n10020) );
  OAI22_X1 U10761 ( .A1(n10020), .A2(n10019), .B1(n10145), .B2(n10018), .ZN(
        n10029) );
  AND2_X1 U10762 ( .A1(n10022), .A2(n10021), .ZN(n10025) );
  OAI211_X1 U10763 ( .C1(n10025), .C2(n10024), .A(n10023), .B(n10140), .ZN(
        n10028) );
  AOI22_X1 U10764 ( .A1(n10026), .A2(n10141), .B1(n10143), .B2(n10071), .ZN(
        n10027) );
  NAND2_X1 U10765 ( .A1(n10028), .A2(n10027), .ZN(n10198) );
  OAI21_X1 U10766 ( .B1(n10029), .B2(n10198), .A(n10148), .ZN(n10030) );
  OAI211_X1 U10767 ( .C1(n10032), .C2(n10137), .A(n10031), .B(n10030), .ZN(
        P1_U3268) );
  XNOR2_X1 U10768 ( .A(n10034), .B(n10033), .ZN(n10207) );
  NAND2_X1 U10769 ( .A1(n10035), .A2(n10036), .ZN(n10039) );
  AND2_X1 U10770 ( .A1(n10039), .A2(n10037), .ZN(n10042) );
  NAND2_X1 U10771 ( .A1(n10039), .A2(n10038), .ZN(n10040) );
  OAI211_X1 U10772 ( .C1(n10042), .C2(n10041), .A(n10040), .B(n10140), .ZN(
        n10045) );
  AOI22_X1 U10773 ( .A1(n10043), .A2(n10141), .B1(n10094), .B2(n10143), .ZN(
        n10044) );
  NAND2_X1 U10774 ( .A1(n10045), .A2(n10044), .ZN(n10203) );
  INV_X1 U10775 ( .A(n10205), .ZN(n10053) );
  INV_X1 U10776 ( .A(n10047), .ZN(n10048) );
  AOI211_X1 U10777 ( .C1(n10205), .C2(n10074), .A(n10591), .B(n10048), .ZN(
        n10204) );
  NAND2_X1 U10778 ( .A1(n10204), .A2(n10110), .ZN(n10052) );
  INV_X1 U10779 ( .A(n10049), .ZN(n10050) );
  AOI22_X1 U10780 ( .A1(n10050), .A2(n10111), .B1(P1_REG2_REG_22__SCAN_IN), 
        .B2(n10088), .ZN(n10051) );
  OAI211_X1 U10781 ( .C1(n10053), .C2(n10115), .A(n10052), .B(n10051), .ZN(
        n10054) );
  AOI21_X1 U10782 ( .B1(n10148), .B2(n10203), .A(n10054), .ZN(n10055) );
  OAI21_X1 U10783 ( .B1(n10207), .B2(n10137), .A(n10055), .ZN(P1_U3269) );
  NAND2_X1 U10784 ( .A1(n10056), .A2(n10057), .ZN(n10059) );
  NAND2_X1 U10785 ( .A1(n10059), .A2(n10058), .ZN(n10082) );
  NAND2_X1 U10786 ( .A1(n10082), .A2(n10092), .ZN(n10061) );
  NAND2_X1 U10787 ( .A1(n10061), .A2(n10060), .ZN(n10062) );
  XOR2_X1 U10788 ( .A(n10067), .B(n10062), .Z(n10210) );
  INV_X1 U10789 ( .A(n10210), .ZN(n10081) );
  NAND2_X1 U10790 ( .A1(n10035), .A2(n10099), .ZN(n10064) );
  NAND2_X1 U10791 ( .A1(n10064), .A2(n10063), .ZN(n10091) );
  OAI21_X1 U10792 ( .B1(n10091), .B2(n10066), .A(n10065), .ZN(n10068) );
  XNOR2_X1 U10793 ( .A(n10068), .B(n10067), .ZN(n10069) );
  NAND2_X1 U10794 ( .A1(n10069), .A2(n10140), .ZN(n10073) );
  AOI22_X1 U10795 ( .A1(n10071), .A2(n10141), .B1(n10143), .B2(n10070), .ZN(
        n10072) );
  NAND2_X1 U10796 ( .A1(n10073), .A2(n10072), .ZN(n10208) );
  INV_X1 U10797 ( .A(n10075), .ZN(n10296) );
  AOI211_X1 U10798 ( .C1(n10075), .C2(n10083), .A(n10591), .B(n10046), .ZN(
        n10209) );
  NAND2_X1 U10799 ( .A1(n10209), .A2(n10110), .ZN(n10078) );
  AOI22_X1 U10800 ( .A1(n10088), .A2(P1_REG2_REG_21__SCAN_IN), .B1(n10076), 
        .B2(n10111), .ZN(n10077) );
  OAI211_X1 U10801 ( .C1(n10296), .C2(n10115), .A(n10078), .B(n10077), .ZN(
        n10079) );
  AOI21_X1 U10802 ( .B1(n10208), .B2(n10148), .A(n10079), .ZN(n10080) );
  OAI21_X1 U10803 ( .B1(n10081), .B2(n10137), .A(n10080), .ZN(P1_U3270) );
  XNOR2_X1 U10804 ( .A(n10082), .B(n10092), .ZN(n10217) );
  INV_X1 U10805 ( .A(n10108), .ZN(n10085) );
  INV_X1 U10806 ( .A(n10083), .ZN(n10084) );
  AOI21_X1 U10807 ( .B1(n10213), .B2(n10085), .A(n10084), .ZN(n10214) );
  INV_X1 U10808 ( .A(n10086), .ZN(n10087) );
  AOI22_X1 U10809 ( .A1(n10088), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n10087), 
        .B2(n10111), .ZN(n10089) );
  OAI21_X1 U10810 ( .B1(n10090), .B2(n10115), .A(n10089), .ZN(n10096) );
  XOR2_X1 U10811 ( .A(n10092), .B(n10091), .Z(n10093) );
  AOI222_X1 U10812 ( .A1(n10125), .A2(n10143), .B1(n10094), .B2(n10141), .C1(
        n10140), .C2(n10093), .ZN(n10216) );
  NOR2_X1 U10813 ( .A1(n10216), .A2(n10088), .ZN(n10095) );
  AOI211_X1 U10814 ( .C1(n10214), .C2(n10097), .A(n10096), .B(n10095), .ZN(
        n10098) );
  OAI21_X1 U10815 ( .B1(n10137), .B2(n10217), .A(n10098), .ZN(P1_U3271) );
  XNOR2_X1 U10816 ( .A(n10056), .B(n10099), .ZN(n10220) );
  INV_X1 U10817 ( .A(n10220), .ZN(n10118) );
  XNOR2_X1 U10818 ( .A(n10035), .B(n10099), .ZN(n10100) );
  NAND2_X1 U10819 ( .A1(n10100), .A2(n10140), .ZN(n10107) );
  OAI22_X1 U10820 ( .A1(n10104), .A2(n10103), .B1(n10102), .B2(n10101), .ZN(
        n10105) );
  INV_X1 U10821 ( .A(n10105), .ZN(n10106) );
  NAND2_X1 U10822 ( .A1(n10107), .A2(n10106), .ZN(n10218) );
  AOI211_X1 U10823 ( .C1(n10109), .C2(n4903), .A(n10591), .B(n10108), .ZN(
        n10219) );
  NAND2_X1 U10824 ( .A1(n10219), .A2(n10110), .ZN(n10114) );
  AOI22_X1 U10825 ( .A1(n10088), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n10112), 
        .B2(n10111), .ZN(n10113) );
  OAI211_X1 U10826 ( .C1(n10301), .C2(n10115), .A(n10114), .B(n10113), .ZN(
        n10116) );
  AOI21_X1 U10827 ( .B1(n10218), .B2(n10148), .A(n10116), .ZN(n10117) );
  OAI21_X1 U10828 ( .B1(n10118), .B2(n10137), .A(n10117), .ZN(P1_U3272) );
  NAND2_X1 U10829 ( .A1(n10120), .A2(n10119), .ZN(n10121) );
  NAND2_X1 U10830 ( .A1(n10122), .A2(n10121), .ZN(n10228) );
  XNOR2_X1 U10831 ( .A(n10123), .B(n5095), .ZN(n10124) );
  NAND2_X1 U10832 ( .A1(n10124), .A2(n10140), .ZN(n10128) );
  AOI22_X1 U10833 ( .A1(n10126), .A2(n10143), .B1(n10141), .B2(n10125), .ZN(
        n10127) );
  NAND2_X1 U10834 ( .A1(n10128), .A2(n10127), .ZN(n10226) );
  OR2_X1 U10835 ( .A1(n10223), .A2(n10149), .ZN(n10129) );
  NAND2_X1 U10836 ( .A1(n10129), .A2(n4903), .ZN(n10224) );
  OAI22_X1 U10837 ( .A1(n10148), .A2(n10131), .B1(n10130), .B2(n10145), .ZN(
        n10132) );
  AOI21_X1 U10838 ( .B1(n10133), .B2(n10156), .A(n10132), .ZN(n10134) );
  OAI21_X1 U10839 ( .B1(n10224), .B2(n10152), .A(n10134), .ZN(n10135) );
  AOI21_X1 U10840 ( .B1(n10226), .B2(n10148), .A(n10135), .ZN(n10136) );
  OAI21_X1 U10841 ( .B1(n10228), .B2(n10137), .A(n10136), .ZN(P1_U3273) );
  XNOR2_X1 U10842 ( .A(n10138), .B(n10157), .ZN(n10139) );
  AOI222_X1 U10843 ( .A1(n10144), .A2(n10143), .B1(n10142), .B2(n10141), .C1(
        n10140), .C2(n10139), .ZN(n10229) );
  INV_X1 U10844 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n10147) );
  OAI22_X1 U10845 ( .A1(n10148), .A2(n10147), .B1(n10146), .B2(n10145), .ZN(
        n10154) );
  INV_X1 U10846 ( .A(n10149), .ZN(n10150) );
  OAI21_X1 U10847 ( .B1(n10306), .B2(n10151), .A(n10150), .ZN(n10230) );
  NOR2_X1 U10848 ( .A1(n10230), .A2(n10152), .ZN(n10153) );
  AOI211_X1 U10849 ( .C1(n10156), .C2(n10155), .A(n10154), .B(n10153), .ZN(
        n10161) );
  XNOR2_X1 U10850 ( .A(n10158), .B(n10157), .ZN(n10232) );
  NAND2_X1 U10851 ( .A1(n10232), .A2(n10159), .ZN(n10160) );
  OAI211_X1 U10852 ( .C1(n10229), .C2(n10088), .A(n10161), .B(n10160), .ZN(
        P1_U3274) );
  NAND3_X1 U10853 ( .A1(n10163), .A2(n10162), .A3(n5984), .ZN(n10165) );
  MUX2_X1 U10854 ( .A(n10166), .B(n10277), .S(n10608), .Z(n10167) );
  OAI21_X1 U10855 ( .B1(n10279), .B2(n10246), .A(n10167), .ZN(P1_U3553) );
  AOI21_X1 U10856 ( .B1(n10269), .B2(n10169), .A(n10168), .ZN(n10170) );
  OAI211_X1 U10857 ( .C1(n10172), .C2(n10240), .A(n10171), .B(n10170), .ZN(
        n10280) );
  MUX2_X1 U10858 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n10280), .S(n10608), .Z(
        P1_U3552) );
  AOI22_X1 U10859 ( .A1(n10174), .A2(n5984), .B1(n10269), .B2(n10173), .ZN(
        n10175) );
  OAI211_X1 U10860 ( .C1(n10273), .C2(n10177), .A(n10176), .B(n10175), .ZN(
        n10281) );
  MUX2_X1 U10861 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n10281), .S(n10608), .Z(
        P1_U3551) );
  INV_X1 U10862 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n10179) );
  MUX2_X1 U10863 ( .A(n10179), .B(n10178), .S(n10608), .Z(n10180) );
  OAI21_X1 U10864 ( .B1(n10181), .B2(n10246), .A(n10180), .ZN(P1_U3550) );
  AOI22_X1 U10865 ( .A1(n10183), .A2(n5984), .B1(n10269), .B2(n10182), .ZN(
        n10184) );
  OAI211_X1 U10866 ( .C1(n10186), .C2(n10240), .A(n10185), .B(n10184), .ZN(
        n10282) );
  MUX2_X1 U10867 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n10282), .S(n10608), .Z(
        P1_U3549) );
  AOI211_X1 U10868 ( .C1(n10269), .C2(n10189), .A(n10188), .B(n10187), .ZN(
        n10190) );
  OAI21_X1 U10869 ( .B1(n10191), .B2(n10240), .A(n10190), .ZN(n10283) );
  MUX2_X1 U10870 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n10283), .S(n10608), .Z(
        P1_U3548) );
  INV_X1 U10871 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n10195) );
  AOI211_X1 U10872 ( .C1(n10194), .C2(n10595), .A(n10193), .B(n10192), .ZN(
        n10284) );
  MUX2_X1 U10873 ( .A(n10195), .B(n10284), .S(n10608), .Z(n10196) );
  OAI21_X1 U10874 ( .B1(n10287), .B2(n10246), .A(n10196), .ZN(P1_U3547) );
  INV_X1 U10875 ( .A(n10197), .ZN(n10291) );
  INV_X1 U10876 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n10201) );
  AOI211_X1 U10877 ( .C1(n10200), .C2(n10595), .A(n10199), .B(n10198), .ZN(
        n10288) );
  MUX2_X1 U10878 ( .A(n10201), .B(n10288), .S(n10608), .Z(n10202) );
  OAI21_X1 U10879 ( .B1(n10291), .B2(n10246), .A(n10202), .ZN(P1_U3546) );
  AOI211_X1 U10880 ( .C1(n10269), .C2(n10205), .A(n10204), .B(n10203), .ZN(
        n10206) );
  OAI21_X1 U10881 ( .B1(n10207), .B2(n10240), .A(n10206), .ZN(n10292) );
  MUX2_X1 U10882 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n10292), .S(n10608), .Z(
        P1_U3545) );
  INV_X1 U10883 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n10211) );
  AOI211_X1 U10884 ( .C1(n10210), .C2(n10595), .A(n10209), .B(n10208), .ZN(
        n10293) );
  MUX2_X1 U10885 ( .A(n10211), .B(n10293), .S(n10608), .Z(n10212) );
  OAI21_X1 U10886 ( .B1(n10296), .B2(n10246), .A(n10212), .ZN(P1_U3544) );
  AOI22_X1 U10887 ( .A1(n10214), .A2(n5984), .B1(n10269), .B2(n10213), .ZN(
        n10215) );
  OAI211_X1 U10888 ( .C1(n10240), .C2(n10217), .A(n10216), .B(n10215), .ZN(
        n10297) );
  MUX2_X1 U10889 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n10297), .S(n10608), .Z(
        P1_U3543) );
  AOI211_X1 U10890 ( .C1(n10220), .C2(n10595), .A(n10219), .B(n10218), .ZN(
        n10298) );
  MUX2_X1 U10891 ( .A(n10221), .B(n10298), .S(n10608), .Z(n10222) );
  OAI21_X1 U10892 ( .B1(n10301), .B2(n10246), .A(n10222), .ZN(P1_U3542) );
  INV_X1 U10893 ( .A(n10269), .ZN(n10600) );
  OAI22_X1 U10894 ( .A1(n10224), .A2(n10591), .B1(n10223), .B2(n10600), .ZN(
        n10225) );
  NOR2_X1 U10895 ( .A1(n10226), .A2(n10225), .ZN(n10227) );
  OAI21_X1 U10896 ( .B1(n10228), .B2(n10240), .A(n10227), .ZN(n10302) );
  MUX2_X1 U10897 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n10302), .S(n10608), .Z(
        P1_U3541) );
  OAI21_X1 U10898 ( .B1(n10591), .B2(n10230), .A(n10229), .ZN(n10231) );
  AOI21_X1 U10899 ( .B1(n10232), .B2(n10595), .A(n10231), .ZN(n10303) );
  MUX2_X1 U10900 ( .A(n10233), .B(n10303), .S(n10608), .Z(n10234) );
  OAI21_X1 U10901 ( .B1(n10306), .B2(n10246), .A(n10234), .ZN(P1_U3540) );
  AOI211_X1 U10902 ( .C1(n10269), .C2(n10237), .A(n10236), .B(n10235), .ZN(
        n10238) );
  OAI21_X1 U10903 ( .B1(n10240), .B2(n10239), .A(n10238), .ZN(n10307) );
  MUX2_X1 U10904 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n10307), .S(n10608), .Z(
        P1_U3539) );
  AOI211_X1 U10905 ( .C1(n10243), .C2(n10595), .A(n10242), .B(n10241), .ZN(
        n10308) );
  MUX2_X1 U10906 ( .A(n10244), .B(n10308), .S(n10608), .Z(n10245) );
  OAI21_X1 U10907 ( .B1(n10312), .B2(n10246), .A(n10245), .ZN(P1_U3538) );
  NAND2_X1 U10908 ( .A1(n10247), .A2(n10595), .ZN(n10253) );
  OAI21_X1 U10909 ( .B1(n10249), .B2(n10600), .A(n10248), .ZN(n10250) );
  NOR2_X1 U10910 ( .A1(n10251), .A2(n10250), .ZN(n10252) );
  NAND2_X1 U10911 ( .A1(n10253), .A2(n10252), .ZN(n10313) );
  MUX2_X1 U10912 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n10313), .S(n10608), .Z(
        P1_U3537) );
  INV_X1 U10913 ( .A(n10254), .ZN(n10255) );
  OAI22_X1 U10914 ( .A1(n10256), .A2(n10591), .B1(n10255), .B2(n10600), .ZN(
        n10257) );
  AOI21_X1 U10915 ( .B1(n10258), .B2(n10603), .A(n10257), .ZN(n10259) );
  NAND2_X1 U10916 ( .A1(n10260), .A2(n10259), .ZN(n10314) );
  MUX2_X1 U10917 ( .A(P1_REG1_REG_13__SCAN_IN), .B(n10314), .S(n10608), .Z(
        P1_U3536) );
  INV_X1 U10918 ( .A(n10261), .ZN(n10266) );
  AOI21_X1 U10919 ( .B1(n10269), .B2(n10263), .A(n10262), .ZN(n10264) );
  OAI211_X1 U10920 ( .C1(n10273), .C2(n10266), .A(n10265), .B(n10264), .ZN(
        n10315) );
  MUX2_X1 U10921 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n10315), .S(n10608), .Z(
        P1_U3535) );
  INV_X1 U10922 ( .A(n10267), .ZN(n10274) );
  AOI22_X1 U10923 ( .A1(n10270), .A2(n5984), .B1(n10269), .B2(n10268), .ZN(
        n10271) );
  OAI211_X1 U10924 ( .C1(n10274), .C2(n10273), .A(n10272), .B(n10271), .ZN(
        n10316) );
  MUX2_X1 U10925 ( .A(P1_REG1_REG_11__SCAN_IN), .B(n10316), .S(n10608), .Z(
        P1_U3534) );
  MUX2_X1 U10926 ( .A(P1_REG1_REG_0__SCAN_IN), .B(n10275), .S(n10608), .Z(
        P1_U3523) );
  INV_X1 U10927 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n10276) );
  MUX2_X1 U10928 ( .A(n10277), .B(n10276), .S(n10609), .Z(n10278) );
  OAI21_X1 U10929 ( .B1(n10279), .B2(n10311), .A(n10278), .ZN(P1_U3521) );
  MUX2_X1 U10930 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n10280), .S(n10612), .Z(
        P1_U3520) );
  MUX2_X1 U10931 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n10281), .S(n10612), .Z(
        P1_U3519) );
  MUX2_X1 U10932 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n10282), .S(n10612), .Z(
        P1_U3517) );
  MUX2_X1 U10933 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n10283), .S(n10612), .Z(
        P1_U3516) );
  MUX2_X1 U10934 ( .A(n10285), .B(n10284), .S(n10612), .Z(n10286) );
  OAI21_X1 U10935 ( .B1(n10287), .B2(n10311), .A(n10286), .ZN(P1_U3515) );
  MUX2_X1 U10936 ( .A(n10289), .B(n10288), .S(n10612), .Z(n10290) );
  OAI21_X1 U10937 ( .B1(n10291), .B2(n10311), .A(n10290), .ZN(P1_U3514) );
  MUX2_X1 U10938 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n10292), .S(n10612), .Z(
        P1_U3513) );
  INV_X1 U10939 ( .A(P1_REG0_REG_21__SCAN_IN), .ZN(n10294) );
  MUX2_X1 U10940 ( .A(n10294), .B(n10293), .S(n10612), .Z(n10295) );
  OAI21_X1 U10941 ( .B1(n10296), .B2(n10311), .A(n10295), .ZN(P1_U3512) );
  MUX2_X1 U10942 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n10297), .S(n10612), .Z(
        P1_U3511) );
  INV_X1 U10943 ( .A(P1_REG0_REG_19__SCAN_IN), .ZN(n10299) );
  MUX2_X1 U10944 ( .A(n10299), .B(n10298), .S(n10612), .Z(n10300) );
  OAI21_X1 U10945 ( .B1(n10301), .B2(n10311), .A(n10300), .ZN(P1_U3510) );
  MUX2_X1 U10946 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n10302), .S(n10612), .Z(
        P1_U3508) );
  MUX2_X1 U10947 ( .A(n10304), .B(n10303), .S(n10612), .Z(n10305) );
  OAI21_X1 U10948 ( .B1(n10306), .B2(n10311), .A(n10305), .ZN(P1_U3505) );
  MUX2_X1 U10949 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n10307), .S(n10612), .Z(
        P1_U3502) );
  INV_X1 U10950 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n10309) );
  MUX2_X1 U10951 ( .A(n10309), .B(n10308), .S(n10612), .Z(n10310) );
  OAI21_X1 U10952 ( .B1(n10312), .B2(n10311), .A(n10310), .ZN(P1_U3499) );
  MUX2_X1 U10953 ( .A(P1_REG0_REG_14__SCAN_IN), .B(n10313), .S(n10612), .Z(
        P1_U3496) );
  MUX2_X1 U10954 ( .A(P1_REG0_REG_13__SCAN_IN), .B(n10314), .S(n10612), .Z(
        P1_U3493) );
  MUX2_X1 U10955 ( .A(P1_REG0_REG_12__SCAN_IN), .B(n10315), .S(n10612), .Z(
        P1_U3490) );
  MUX2_X1 U10956 ( .A(P1_REG0_REG_11__SCAN_IN), .B(n10316), .S(n10612), .Z(
        P1_U3487) );
  CLKBUF_X1 U10957 ( .A(n10345), .Z(n10359) );
  MUX2_X1 U10958 ( .A(P1_D_REG_0__SCAN_IN), .B(n10318), .S(n10359), .Z(
        P1_U3440) );
  INV_X1 U10959 ( .A(n9704), .ZN(n10322) );
  NOR4_X1 U10960 ( .A1(n5201), .A2(P1_IR_REG_30__SCAN_IN), .A3(P1_U3084), .A4(
        n10319), .ZN(n10320) );
  AOI21_X1 U10961 ( .B1(P2_DATAO_REG_31__SCAN_IN), .B2(n10324), .A(n10320), 
        .ZN(n10321) );
  OAI21_X1 U10962 ( .B1(n10322), .B2(n6276), .A(n10321), .ZN(P1_U3322) );
  AOI22_X1 U10963 ( .A1(n10323), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_30__SCAN_IN), .B2(n10324), .ZN(n10325) );
  OAI21_X1 U10964 ( .B1(n10326), .B2(n6276), .A(n10325), .ZN(P1_U3323) );
  MUX2_X1 U10965 ( .A(n10327), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3353) );
  INV_X1 U10966 ( .A(P1_D_REG_2__SCAN_IN), .ZN(n10328) );
  NOR2_X1 U10967 ( .A1(n10345), .A2(n10328), .ZN(P1_U3321) );
  INV_X1 U10968 ( .A(P1_D_REG_3__SCAN_IN), .ZN(n10329) );
  NOR2_X1 U10969 ( .A1(n10345), .A2(n10329), .ZN(P1_U3320) );
  INV_X1 U10970 ( .A(P1_D_REG_4__SCAN_IN), .ZN(n10330) );
  NOR2_X1 U10971 ( .A1(n10359), .A2(n10330), .ZN(P1_U3319) );
  INV_X1 U10972 ( .A(P1_D_REG_5__SCAN_IN), .ZN(n10331) );
  NOR2_X1 U10973 ( .A1(n10359), .A2(n10331), .ZN(P1_U3318) );
  INV_X1 U10974 ( .A(P1_D_REG_6__SCAN_IN), .ZN(n10332) );
  NOR2_X1 U10975 ( .A1(n10359), .A2(n10332), .ZN(P1_U3317) );
  INV_X1 U10976 ( .A(P1_D_REG_7__SCAN_IN), .ZN(n10333) );
  NOR2_X1 U10977 ( .A1(n10359), .A2(n10333), .ZN(P1_U3316) );
  INV_X1 U10978 ( .A(P1_D_REG_8__SCAN_IN), .ZN(n10334) );
  NOR2_X1 U10979 ( .A1(n10359), .A2(n10334), .ZN(P1_U3315) );
  INV_X1 U10980 ( .A(P1_D_REG_9__SCAN_IN), .ZN(n10335) );
  NOR2_X1 U10981 ( .A1(n10359), .A2(n10335), .ZN(P1_U3314) );
  INV_X1 U10982 ( .A(P1_D_REG_10__SCAN_IN), .ZN(n10336) );
  NOR2_X1 U10983 ( .A1(n10359), .A2(n10336), .ZN(P1_U3313) );
  INV_X1 U10984 ( .A(P1_D_REG_11__SCAN_IN), .ZN(n10337) );
  NOR2_X1 U10985 ( .A1(n10345), .A2(n10337), .ZN(P1_U3312) );
  INV_X1 U10986 ( .A(P1_D_REG_12__SCAN_IN), .ZN(n10338) );
  NOR2_X1 U10987 ( .A1(n10345), .A2(n10338), .ZN(P1_U3311) );
  INV_X1 U10988 ( .A(P1_D_REG_13__SCAN_IN), .ZN(n10339) );
  NOR2_X1 U10989 ( .A1(n10345), .A2(n10339), .ZN(P1_U3310) );
  INV_X1 U10990 ( .A(P1_D_REG_14__SCAN_IN), .ZN(n10340) );
  NOR2_X1 U10991 ( .A1(n10345), .A2(n10340), .ZN(P1_U3309) );
  INV_X1 U10992 ( .A(P1_D_REG_15__SCAN_IN), .ZN(n10341) );
  NOR2_X1 U10993 ( .A1(n10345), .A2(n10341), .ZN(P1_U3308) );
  INV_X1 U10994 ( .A(P1_D_REG_16__SCAN_IN), .ZN(n10342) );
  NOR2_X1 U10995 ( .A1(n10345), .A2(n10342), .ZN(P1_U3307) );
  INV_X1 U10996 ( .A(P1_D_REG_17__SCAN_IN), .ZN(n10343) );
  NOR2_X1 U10997 ( .A1(n10345), .A2(n10343), .ZN(P1_U3306) );
  INV_X1 U10998 ( .A(P1_D_REG_18__SCAN_IN), .ZN(n10344) );
  NOR2_X1 U10999 ( .A1(n10345), .A2(n10344), .ZN(P1_U3305) );
  INV_X1 U11000 ( .A(P1_D_REG_19__SCAN_IN), .ZN(n10346) );
  NOR2_X1 U11001 ( .A1(n10359), .A2(n10346), .ZN(P1_U3304) );
  INV_X1 U11002 ( .A(P1_D_REG_20__SCAN_IN), .ZN(n10347) );
  NOR2_X1 U11003 ( .A1(n10359), .A2(n10347), .ZN(P1_U3303) );
  INV_X1 U11004 ( .A(P1_D_REG_21__SCAN_IN), .ZN(n10348) );
  NOR2_X1 U11005 ( .A1(n10359), .A2(n10348), .ZN(P1_U3302) );
  INV_X1 U11006 ( .A(P1_D_REG_22__SCAN_IN), .ZN(n10349) );
  NOR2_X1 U11007 ( .A1(n10359), .A2(n10349), .ZN(P1_U3301) );
  INV_X1 U11008 ( .A(P1_D_REG_23__SCAN_IN), .ZN(n10350) );
  NOR2_X1 U11009 ( .A1(n10359), .A2(n10350), .ZN(P1_U3300) );
  INV_X1 U11010 ( .A(P1_D_REG_24__SCAN_IN), .ZN(n10351) );
  NOR2_X1 U11011 ( .A1(n10359), .A2(n10351), .ZN(P1_U3299) );
  INV_X1 U11012 ( .A(P1_D_REG_25__SCAN_IN), .ZN(n10352) );
  NOR2_X1 U11013 ( .A1(n10359), .A2(n10352), .ZN(P1_U3298) );
  INV_X1 U11014 ( .A(P1_D_REG_26__SCAN_IN), .ZN(n10353) );
  NOR2_X1 U11015 ( .A1(n10359), .A2(n10353), .ZN(P1_U3297) );
  INV_X1 U11016 ( .A(P1_D_REG_27__SCAN_IN), .ZN(n10354) );
  NOR2_X1 U11017 ( .A1(n10359), .A2(n10354), .ZN(P1_U3296) );
  INV_X1 U11018 ( .A(P1_D_REG_28__SCAN_IN), .ZN(n10355) );
  NOR2_X1 U11019 ( .A1(n10359), .A2(n10355), .ZN(P1_U3295) );
  INV_X1 U11020 ( .A(P1_D_REG_29__SCAN_IN), .ZN(n10356) );
  NOR2_X1 U11021 ( .A1(n10359), .A2(n10356), .ZN(P1_U3294) );
  INV_X1 U11022 ( .A(P1_D_REG_30__SCAN_IN), .ZN(n10357) );
  NOR2_X1 U11023 ( .A1(n10359), .A2(n10357), .ZN(P1_U3293) );
  INV_X1 U11024 ( .A(P1_D_REG_31__SCAN_IN), .ZN(n10358) );
  NOR2_X1 U11025 ( .A1(n10359), .A2(n10358), .ZN(P1_U3292) );
  INV_X1 U11026 ( .A(n10360), .ZN(n10364) );
  INV_X1 U11027 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n10363) );
  AOI22_X1 U11028 ( .A1(n10364), .A2(n10464), .B1(n10363), .B2(n10462), .ZN(
        P2_U3438) );
  AND2_X1 U11029 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n10462), .ZN(P2_U3326) );
  AND2_X1 U11030 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n10462), .ZN(P2_U3325) );
  AND2_X1 U11031 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n10462), .ZN(P2_U3324) );
  AND2_X1 U11032 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n10462), .ZN(P2_U3323) );
  AND2_X1 U11033 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n10462), .ZN(P2_U3322) );
  AND2_X1 U11034 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n10462), .ZN(P2_U3321) );
  AND2_X1 U11035 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n10462), .ZN(P2_U3320) );
  AND2_X1 U11036 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n10462), .ZN(P2_U3319) );
  AND2_X1 U11037 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n10462), .ZN(P2_U3318) );
  AND2_X1 U11038 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n10462), .ZN(P2_U3317) );
  AND2_X1 U11039 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n10462), .ZN(P2_U3316) );
  AND2_X1 U11040 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n10462), .ZN(P2_U3315) );
  AND2_X1 U11041 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n10462), .ZN(P2_U3314) );
  AND2_X1 U11042 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n10462), .ZN(P2_U3313) );
  AND2_X1 U11043 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n10462), .ZN(P2_U3312) );
  AND2_X1 U11044 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n10462), .ZN(P2_U3311) );
  AND2_X1 U11045 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n10462), .ZN(P2_U3310) );
  AND2_X1 U11046 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n10462), .ZN(P2_U3309) );
  AND2_X1 U11047 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n10462), .ZN(P2_U3308) );
  AND2_X1 U11048 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n10462), .ZN(P2_U3307) );
  AND2_X1 U11049 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n10462), .ZN(P2_U3306) );
  AND2_X1 U11050 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n10462), .ZN(P2_U3305) );
  AND2_X1 U11051 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n10462), .ZN(P2_U3304) );
  AND2_X1 U11052 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n10462), .ZN(P2_U3303) );
  AND2_X1 U11053 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n10462), .ZN(P2_U3302) );
  AND2_X1 U11054 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n10462), .ZN(P2_U3301) );
  AND2_X1 U11055 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n10462), .ZN(P2_U3300) );
  AND2_X1 U11056 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n10462), .ZN(P2_U3299) );
  AND2_X1 U11057 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n10462), .ZN(P2_U3298) );
  AND2_X1 U11058 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n10462), .ZN(P2_U3297) );
  XOR2_X1 U11059 ( .A(P2_ADDR_REG_0__SCAN_IN), .B(P1_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1071_U46) );
  INV_X1 U11060 ( .A(n10365), .ZN(n10366) );
  NAND2_X1 U11061 ( .A1(n10367), .A2(n10366), .ZN(n10368) );
  XOR2_X1 U11062 ( .A(n10369), .B(n10368), .Z(ADD_1071_U5) );
  XOR2_X1 U11063 ( .A(n10371), .B(n10370), .Z(ADD_1071_U54) );
  XOR2_X1 U11064 ( .A(n10373), .B(n10372), .Z(ADD_1071_U53) );
  XNOR2_X1 U11065 ( .A(n10375), .B(n10374), .ZN(ADD_1071_U52) );
  NOR2_X1 U11066 ( .A1(n10377), .A2(n10376), .ZN(n10378) );
  XOR2_X1 U11067 ( .A(P2_ADDR_REG_5__SCAN_IN), .B(n10378), .Z(ADD_1071_U51) );
  XOR2_X1 U11068 ( .A(P2_ADDR_REG_6__SCAN_IN), .B(n10379), .Z(ADD_1071_U50) );
  XOR2_X1 U11069 ( .A(P2_ADDR_REG_7__SCAN_IN), .B(n10380), .Z(ADD_1071_U49) );
  XOR2_X1 U11070 ( .A(P2_ADDR_REG_8__SCAN_IN), .B(n10381), .Z(ADD_1071_U48) );
  XOR2_X1 U11071 ( .A(P2_ADDR_REG_9__SCAN_IN), .B(n10382), .Z(ADD_1071_U47) );
  XOR2_X1 U11072 ( .A(n10384), .B(n10383), .Z(ADD_1071_U63) );
  XOR2_X1 U11073 ( .A(n10386), .B(n10385), .Z(ADD_1071_U62) );
  XNOR2_X1 U11074 ( .A(n10388), .B(n10387), .ZN(ADD_1071_U61) );
  XNOR2_X1 U11075 ( .A(n10390), .B(n10389), .ZN(ADD_1071_U60) );
  XNOR2_X1 U11076 ( .A(n10392), .B(n10391), .ZN(ADD_1071_U59) );
  XNOR2_X1 U11077 ( .A(n10394), .B(n10393), .ZN(ADD_1071_U58) );
  XNOR2_X1 U11078 ( .A(n10396), .B(n10395), .ZN(ADD_1071_U57) );
  XNOR2_X1 U11079 ( .A(n10398), .B(n10397), .ZN(ADD_1071_U56) );
  NOR2_X1 U11080 ( .A1(n10400), .A2(n10399), .ZN(n10401) );
  XNOR2_X1 U11081 ( .A(n10402), .B(n10401), .ZN(ADD_1071_U55) );
  INV_X1 U11082 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n10404) );
  AOI21_X1 U11083 ( .B1(n10405), .B2(n10404), .A(n10403), .ZN(P1_U3441) );
  OAI21_X1 U11084 ( .B1(n10407), .B2(P1_REG1_REG_0__SCAN_IN), .A(n10406), .ZN(
        n10414) );
  NOR2_X1 U11085 ( .A1(n10409), .A2(n10408), .ZN(n10412) );
  AOI22_X1 U11086 ( .A1(n10412), .A2(n10411), .B1(n10443), .B2(n10410), .ZN(
        n10413) );
  AOI21_X1 U11087 ( .B1(n10415), .B2(n10414), .A(n10413), .ZN(n10416) );
  AOI21_X1 U11088 ( .B1(n10457), .B2(P1_ADDR_REG_0__SCAN_IN), .A(n10416), .ZN(
        n10417) );
  OAI21_X1 U11089 ( .B1(P1_STATE_REG_SCAN_IN), .B2(n6449), .A(n10417), .ZN(
        P1_U3241) );
  INV_X1 U11090 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n10424) );
  AOI21_X1 U11091 ( .B1(n10420), .B2(n10419), .A(n10418), .ZN(n10422) );
  AOI21_X1 U11092 ( .B1(n10443), .B2(n10422), .A(n10421), .ZN(n10423) );
  OAI21_X1 U11093 ( .B1(n10425), .B2(n10424), .A(n10423), .ZN(n10426) );
  INV_X1 U11094 ( .A(n10426), .ZN(n10433) );
  AOI211_X1 U11095 ( .C1(n10429), .C2(n10428), .A(n10427), .B(n10451), .ZN(
        n10430) );
  AOI21_X1 U11096 ( .B1(n10459), .B2(n10431), .A(n10430), .ZN(n10432) );
  NAND2_X1 U11097 ( .A1(n10433), .A2(n10432), .ZN(P1_U3247) );
  AOI22_X1 U11098 ( .A1(n10459), .A2(n10434), .B1(n10457), .B2(
        P1_ADDR_REG_9__SCAN_IN), .ZN(n10446) );
  OAI21_X1 U11099 ( .B1(n10437), .B2(n10436), .A(n10435), .ZN(n10444) );
  AOI211_X1 U11100 ( .C1(n10440), .C2(n10439), .A(n10438), .B(n10451), .ZN(
        n10441) );
  AOI211_X1 U11101 ( .C1(n10444), .C2(n10443), .A(n10442), .B(n10441), .ZN(
        n10445) );
  NAND2_X1 U11102 ( .A1(n10446), .A2(n10445), .ZN(P1_U3250) );
  NAND2_X1 U11103 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), 
        .ZN(n10450) );
  AOI211_X1 U11104 ( .C1(n10450), .C2(n10449), .A(n10448), .B(n10447), .ZN(
        n10456) );
  AOI211_X1 U11105 ( .C1(n10454), .C2(n10453), .A(n10452), .B(n10451), .ZN(
        n10455) );
  AOI211_X1 U11106 ( .C1(P1_REG3_REG_1__SCAN_IN), .C2(P1_U3084), .A(n10456), 
        .B(n10455), .ZN(n10461) );
  AOI22_X1 U11107 ( .A1(n10459), .A2(n10458), .B1(n10457), .B2(
        P1_ADDR_REG_1__SCAN_IN), .ZN(n10460) );
  NAND2_X1 U11108 ( .A1(n10461), .A2(n10460), .ZN(P1_U3242) );
  AOI22_X1 U11109 ( .A1(n10465), .A2(n10464), .B1(n10463), .B2(n10462), .ZN(
        P2_U3437) );
  AOI22_X1 U11110 ( .A1(n10466), .A2(P2_REG2_REG_0__SCAN_IN), .B1(
        P2_REG1_REG_0__SCAN_IN), .B2(n10495), .ZN(n10473) );
  AOI22_X1 U11111 ( .A1(n10486), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3152), .ZN(n10472) );
  OAI21_X1 U11112 ( .B1(P2_REG1_REG_0__SCAN_IN), .B2(n10468), .A(n10467), .ZN(
        n10470) );
  NOR2_X1 U11113 ( .A1(n10487), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n10469) );
  OAI21_X1 U11114 ( .B1(n10470), .B2(n10469), .A(P2_IR_REG_0__SCAN_IN), .ZN(
        n10471) );
  OAI211_X1 U11115 ( .C1(P2_IR_REG_0__SCAN_IN), .C2(n10473), .A(n10472), .B(
        n10471), .ZN(P2_U3245) );
  AOI22_X1 U11116 ( .A1(n10486), .A2(P2_ADDR_REG_1__SCAN_IN), .B1(
        P2_REG3_REG_1__SCAN_IN), .B2(P2_U3152), .ZN(n10485) );
  AOI211_X1 U11117 ( .C1(n10476), .C2(n10475), .A(n10474), .B(n10487), .ZN(
        n10477) );
  AOI21_X1 U11118 ( .B1(n10493), .B2(n4856), .A(n10477), .ZN(n10484) );
  INV_X1 U11119 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n10479) );
  INV_X1 U11120 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n10506) );
  NOR2_X1 U11121 ( .A1(n10479), .A2(n10506), .ZN(n10482) );
  OAI211_X1 U11122 ( .C1(n10482), .C2(n10481), .A(n10495), .B(n10480), .ZN(
        n10483) );
  NAND3_X1 U11123 ( .A1(n10485), .A2(n10484), .A3(n10483), .ZN(P2_U3246) );
  AOI22_X1 U11124 ( .A1(n10486), .A2(P2_ADDR_REG_2__SCAN_IN), .B1(
        P2_REG3_REG_2__SCAN_IN), .B2(P2_U3152), .ZN(n10500) );
  AOI211_X1 U11125 ( .C1(n10490), .C2(n10489), .A(n10488), .B(n10487), .ZN(
        n10491) );
  AOI21_X1 U11126 ( .B1(n10493), .B2(n10492), .A(n10491), .ZN(n10499) );
  OAI211_X1 U11127 ( .C1(n10497), .C2(n10496), .A(n10495), .B(n10494), .ZN(
        n10498) );
  NAND3_X1 U11128 ( .A1(n10500), .A2(n10499), .A3(n10498), .ZN(P2_U3247) );
  XOR2_X1 U11129 ( .A(n4918), .B(P1_RD_REG_SCAN_IN), .Z(U126) );
  OAI22_X1 U11130 ( .A1(n10503), .A2(n10556), .B1(n10502), .B2(n10501), .ZN(
        n10504) );
  NOR2_X1 U11131 ( .A1(n10505), .A2(n10504), .ZN(n10508) );
  AOI22_X1 U11132 ( .A1(n10642), .A2(n10508), .B1(n10506), .B2(n10641), .ZN(
        P2_U3520) );
  INV_X1 U11133 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n10507) );
  AOI22_X1 U11134 ( .A1(n10646), .A2(n10508), .B1(n10507), .B2(n10643), .ZN(
        P2_U3451) );
  NAND3_X1 U11135 ( .A1(n10511), .A2(n10510), .A3(n10509), .ZN(n10512) );
  OAI21_X1 U11136 ( .B1(n10513), .B2(n10625), .A(n10512), .ZN(n10515) );
  AOI211_X1 U11137 ( .C1(n10516), .C2(n10639), .A(n10515), .B(n10514), .ZN(
        n10518) );
  AOI22_X1 U11138 ( .A1(n10642), .A2(n10518), .B1(n6534), .B2(n10641), .ZN(
        P2_U3521) );
  INV_X1 U11139 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n10517) );
  AOI22_X1 U11140 ( .A1(n10646), .A2(n10518), .B1(n10517), .B2(n10643), .ZN(
        P2_U3454) );
  OAI22_X1 U11141 ( .A1(n10520), .A2(n10591), .B1(n10519), .B2(n10600), .ZN(
        n10522) );
  AOI211_X1 U11142 ( .C1(n10603), .C2(n10523), .A(n10522), .B(n10521), .ZN(
        n10525) );
  AOI22_X1 U11143 ( .A1(n10608), .A2(n10525), .B1(n5459), .B2(n10607), .ZN(
        P1_U3525) );
  INV_X1 U11144 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n10524) );
  AOI22_X1 U11145 ( .A1(n10612), .A2(n10525), .B1(n10524), .B2(n10609), .ZN(
        P1_U3460) );
  NAND2_X1 U11146 ( .A1(n10526), .A2(n10619), .ZN(n10533) );
  INV_X1 U11147 ( .A(n10527), .ZN(n10531) );
  NOR2_X1 U11148 ( .A1(n10528), .A2(n10637), .ZN(n10530) );
  AOI22_X1 U11149 ( .A1(n10531), .A2(n10530), .B1(n10632), .B2(n10529), .ZN(
        n10532) );
  NAND2_X1 U11150 ( .A1(n10533), .A2(n10532), .ZN(n10534) );
  NOR2_X1 U11151 ( .A1(n10535), .A2(n10534), .ZN(n10537) );
  AOI22_X1 U11152 ( .A1(n10642), .A2(n10537), .B1(n6673), .B2(n10641), .ZN(
        P2_U3522) );
  INV_X1 U11153 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n10536) );
  AOI22_X1 U11154 ( .A1(n10646), .A2(n10537), .B1(n10536), .B2(n10643), .ZN(
        P2_U3457) );
  NAND2_X1 U11155 ( .A1(n10538), .A2(n10619), .ZN(n10543) );
  OAI22_X1 U11156 ( .A1(n10540), .A2(n10637), .B1(n10539), .B2(n10625), .ZN(
        n10541) );
  INV_X1 U11157 ( .A(n10541), .ZN(n10542) );
  NAND2_X1 U11158 ( .A1(n10543), .A2(n10542), .ZN(n10544) );
  NOR2_X1 U11159 ( .A1(n10545), .A2(n10544), .ZN(n10548) );
  AOI22_X1 U11160 ( .A1(n10642), .A2(n10548), .B1(n10546), .B2(n10641), .ZN(
        P2_U3523) );
  INV_X1 U11161 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n10547) );
  AOI22_X1 U11162 ( .A1(n10646), .A2(n10548), .B1(n10547), .B2(n10643), .ZN(
        P2_U3460) );
  OAI22_X1 U11163 ( .A1(n10550), .A2(n10591), .B1(n10549), .B2(n10600), .ZN(
        n10552) );
  AOI211_X1 U11164 ( .C1(n10603), .C2(n10553), .A(n10552), .B(n10551), .ZN(
        n10555) );
  AOI22_X1 U11165 ( .A1(n10608), .A2(n10555), .B1(n5486), .B2(n10607), .ZN(
        P1_U3527) );
  INV_X1 U11166 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n10554) );
  AOI22_X1 U11167 ( .A1(n10612), .A2(n10555), .B1(n10554), .B2(n10609), .ZN(
        P1_U3466) );
  NOR2_X1 U11168 ( .A1(n10557), .A2(n10556), .ZN(n10561) );
  OAI22_X1 U11169 ( .A1(n10558), .A2(n10637), .B1(n6519), .B2(n10625), .ZN(
        n10559) );
  NOR3_X1 U11170 ( .A1(n10561), .A2(n10560), .A3(n10559), .ZN(n10563) );
  AOI22_X1 U11171 ( .A1(n10642), .A2(n10563), .B1(n6672), .B2(n10641), .ZN(
        P2_U3524) );
  INV_X1 U11172 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n10562) );
  AOI22_X1 U11173 ( .A1(n10646), .A2(n10563), .B1(n10562), .B2(n10643), .ZN(
        P2_U3463) );
  OAI21_X1 U11174 ( .B1(n10565), .B2(n10625), .A(n10564), .ZN(n10566) );
  INV_X1 U11175 ( .A(n10566), .ZN(n10569) );
  NAND2_X1 U11176 ( .A1(n10567), .A2(n10639), .ZN(n10568) );
  AND3_X1 U11177 ( .A1(n10570), .A2(n10569), .A3(n10568), .ZN(n10572) );
  AOI22_X1 U11178 ( .A1(n10642), .A2(n10572), .B1(n6671), .B2(n10641), .ZN(
        P2_U3525) );
  INV_X1 U11179 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n10571) );
  AOI22_X1 U11180 ( .A1(n10646), .A2(n10572), .B1(n10571), .B2(n10643), .ZN(
        P2_U3466) );
  INV_X1 U11181 ( .A(n10573), .ZN(n10578) );
  OAI22_X1 U11182 ( .A1(n10575), .A2(n10591), .B1(n10574), .B2(n10600), .ZN(
        n10577) );
  AOI211_X1 U11183 ( .C1(n10603), .C2(n10578), .A(n10577), .B(n10576), .ZN(
        n10580) );
  AOI22_X1 U11184 ( .A1(n10608), .A2(n10580), .B1(n5506), .B2(n10607), .ZN(
        P1_U3529) );
  INV_X1 U11185 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n10579) );
  AOI22_X1 U11186 ( .A1(n10612), .A2(n10580), .B1(n10579), .B2(n10609), .ZN(
        P1_U3472) );
  INV_X1 U11187 ( .A(n10581), .ZN(n10587) );
  OAI22_X1 U11188 ( .A1(n10583), .A2(n10637), .B1(n10582), .B2(n10625), .ZN(
        n10586) );
  INV_X1 U11189 ( .A(n10584), .ZN(n10585) );
  AOI211_X1 U11190 ( .C1(n10639), .C2(n10587), .A(n10586), .B(n10585), .ZN(
        n10590) );
  AOI22_X1 U11191 ( .A1(n10642), .A2(n10590), .B1(n10588), .B2(n10641), .ZN(
        P2_U3526) );
  INV_X1 U11192 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n10589) );
  AOI22_X1 U11193 ( .A1(n10646), .A2(n10590), .B1(n10589), .B2(n10643), .ZN(
        P2_U3469) );
  OAI22_X1 U11194 ( .A1(n10592), .A2(n10591), .B1(n5026), .B2(n10600), .ZN(
        n10593) );
  AOI211_X1 U11195 ( .C1(n10596), .C2(n10595), .A(n10594), .B(n10593), .ZN(
        n10598) );
  AOI22_X1 U11196 ( .A1(n10608), .A2(n10598), .B1(n5570), .B2(n10607), .ZN(
        P1_U3531) );
  INV_X1 U11197 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n10597) );
  AOI22_X1 U11198 ( .A1(n10612), .A2(n10598), .B1(n10597), .B2(n10609), .ZN(
        P1_U3478) );
  OAI21_X1 U11199 ( .B1(n10601), .B2(n10600), .A(n10599), .ZN(n10602) );
  AOI21_X1 U11200 ( .B1(n10604), .B2(n10603), .A(n10602), .ZN(n10605) );
  AND2_X1 U11201 ( .A1(n10606), .A2(n10605), .ZN(n10611) );
  AOI22_X1 U11202 ( .A1(n10608), .A2(n10611), .B1(n6064), .B2(n10607), .ZN(
        P1_U3533) );
  INV_X1 U11203 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n10610) );
  AOI22_X1 U11204 ( .A1(n10612), .A2(n10611), .B1(n10610), .B2(n10609), .ZN(
        P1_U3484) );
  INV_X1 U11205 ( .A(n10613), .ZN(n10618) );
  OAI22_X1 U11206 ( .A1(n10615), .A2(n10637), .B1(n10614), .B2(n10625), .ZN(
        n10617) );
  AOI211_X1 U11207 ( .C1(n10619), .C2(n10618), .A(n10617), .B(n10616), .ZN(
        n10622) );
  AOI22_X1 U11208 ( .A1(n10642), .A2(n10622), .B1(n10620), .B2(n10641), .ZN(
        P2_U3530) );
  INV_X1 U11209 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n10621) );
  AOI22_X1 U11210 ( .A1(n10646), .A2(n10622), .B1(n10621), .B2(n10643), .ZN(
        P2_U3481) );
  OAI211_X1 U11211 ( .C1(n10626), .C2(n10625), .A(n10624), .B(n10623), .ZN(
        n10627) );
  AOI21_X1 U11212 ( .B1(n10628), .B2(n10639), .A(n10627), .ZN(n10631) );
  AOI22_X1 U11213 ( .A1(n10642), .A2(n10631), .B1(n10629), .B2(n10641), .ZN(
        P2_U3531) );
  INV_X1 U11214 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n10630) );
  AOI22_X1 U11215 ( .A1(n10646), .A2(n10631), .B1(n10630), .B2(n10643), .ZN(
        P2_U3484) );
  NAND2_X1 U11216 ( .A1(n10633), .A2(n10632), .ZN(n10634) );
  OAI211_X1 U11217 ( .C1(n10637), .C2(n10636), .A(n10635), .B(n10634), .ZN(
        n10638) );
  AOI21_X1 U11218 ( .B1(n10640), .B2(n10639), .A(n10638), .ZN(n10645) );
  AOI22_X1 U11219 ( .A1(n10642), .A2(n10645), .B1(n6680), .B2(n10641), .ZN(
        P2_U3532) );
  INV_X1 U11220 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n10644) );
  AOI22_X1 U11221 ( .A1(n10646), .A2(n10645), .B1(n10644), .B2(n10643), .ZN(
        P2_U3487) );
  XNOR2_X1 U11222 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  CLKBUF_X2 U4923 ( .A(n6585), .Z(n8195) );
  CLKBUF_X1 U4932 ( .A(n5485), .Z(n5978) );
endmodule

