

module b21_C_2inp_gates_syn ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, 
        P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, 
        P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, 
        P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, 
        P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, 
        P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, 
        P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, 
        P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, 
        P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, 
        P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, 
        P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, 
        P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, 
        P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, 
        P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, 
        P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, 
        P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, 
        P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, 
        P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, 
        P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, 
        P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, 
        P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, 
        P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, 
        P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, 
        P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, 
        P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, 
        ADD_1071_U57, ADD_1071_U58, ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, 
        ADD_1071_U62, ADD_1071_U63, ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, 
        ADD_1071_U50, ADD_1071_U51, ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, 
        ADD_1071_U5, ADD_1071_U46, U126, U123, P1_U3353, P1_U3352, P1_U3351, 
        P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, 
        P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, 
        P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, 
        P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, 
        P1_U3322, P1_U3440, P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, 
        P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, 
        P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, 
        P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, 
        P1_U3296, P1_U3295, P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, 
        P1_U3460, P1_U3463, P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, 
        P1_U3481, P1_U3484, P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, 
        P1_U3502, P1_U3505, P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, 
        P1_U3514, P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, 
        P1_U3521, P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, 
        P1_U3528, P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, 
        P1_U3535, P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, 
        P1_U3542, P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, 
        P1_U3549, P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, 
        P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, 
        P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, 
        P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, 
        P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, 
        P1_U3355, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, 
        P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, 
        P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, 
        P1_U3242, P1_U3241, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, 
        P1_U3560, P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, 
        P1_U3567, P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, 
        P1_U3574, P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, 
        P1_U3581, P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, 
        P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, 
        P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, 
        P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, 
        P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, 
        P1_U3211, P1_U3084, P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, 
        P2_U3355, P2_U3354, P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, 
        P2_U3348, P2_U3347, P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, 
        P2_U3341, P2_U3340, P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, 
        P2_U3334, P2_U3333, P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, 
        P2_U3327, P2_U3437, P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, 
        P2_U3322, P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, 
        P2_U3315, P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, 
        P2_U3308, P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, 
        P2_U3301, P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, 
        P2_U3457, P2_U3460, P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, 
        P2_U3478, P2_U3481, P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, 
        P2_U3499, P2_U3502, P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, 
        P2_U3511, P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, 
        P2_U3518, P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, 
        P2_U3525, P2_U3526, P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, 
        P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, 
        P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, 
        P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, 
        P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, 
        P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, 
        P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, 
        P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, 
        P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, 
        P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, 
        P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, 
        P2_U3246, P2_U3245, P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, 
        P2_U3557, P2_U3558, P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, 
        P2_U3564, P2_U3565, P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, 
        P2_U3571, P2_U3572, P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, 
        P2_U3578, P2_U3579, P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, 
        P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, 
        P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, 
        P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, 
        P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, 
        P2_U3215, P2_U3152, P2_U3151, P2_U3966, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN,
         P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN,
         P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN,
         P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN,
         P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN,
         P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN,
         P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN,
         P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN,
         P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN,
         P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN,
         P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN,
         P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN,
         P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN,
         P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN,
         P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN,
         P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN,
         P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN,
         P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN,
         P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN,
         P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN,
         P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN,
         P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63;
  output ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, ADD_1071_U57, ADD_1071_U58,
         ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, ADD_1071_U62, ADD_1071_U63,
         ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, ADD_1071_U50, ADD_1071_U51,
         ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, ADD_1071_U5, ADD_1071_U46,
         U126, U123, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349,
         P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342,
         P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335,
         P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328,
         P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, P1_U3322, P1_U3440,
         P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316,
         P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309,
         P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302,
         P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295,
         P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, P1_U3460, P1_U3463,
         P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, P1_U3481, P1_U3484,
         P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, P1_U3502, P1_U3505,
         P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515,
         P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522,
         P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529,
         P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536,
         P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543,
         P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550,
         P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, P1_U3290, P1_U3289,
         P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282,
         P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275,
         P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268,
         P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, P1_U3355, P1_U3262,
         P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255,
         P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248,
         P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3242, P1_U3241,
         P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561,
         P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568,
         P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575,
         P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582,
         P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, P1_U3239, P1_U3238,
         P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231,
         P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224,
         P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217,
         P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, P1_U3084,
         P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, P2_U3355, P2_U3354,
         P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, P2_U3348, P2_U3347,
         P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, P2_U3341, P2_U3340,
         P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, P2_U3334, P2_U3333,
         P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, P2_U3327, P2_U3437,
         P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321,
         P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314,
         P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307,
         P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300,
         P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, P2_U3457, P2_U3460,
         P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481,
         P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, P2_U3499, P2_U3502,
         P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512,
         P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519,
         P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526,
         P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, P2_U3532, P2_U3533,
         P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540,
         P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547,
         P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, P2_U3295, P2_U3294,
         P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287,
         P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280,
         P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273,
         P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266,
         P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259,
         P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252,
         P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245,
         P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558,
         P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, P2_U3564, P2_U3565,
         P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, P2_U3571, P2_U3572,
         P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, P2_U3578, P2_U3579,
         P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, P2_U3243, P2_U3242,
         P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235,
         P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228,
         P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221,
         P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3152,
         P2_U3151, P2_U3966;
  wire   n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267,
         n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277,
         n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287,
         n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297,
         n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307,
         n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317,
         n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327,
         n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337,
         n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347,
         n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357,
         n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367,
         n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377,
         n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387,
         n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397,
         n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407,
         n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417,
         n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427,
         n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437,
         n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447,
         n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457,
         n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467,
         n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477,
         n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487,
         n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497,
         n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507,
         n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517,
         n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527,
         n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537,
         n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547,
         n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557,
         n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567,
         n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577,
         n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587,
         n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597,
         n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607,
         n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617,
         n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627,
         n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637,
         n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647,
         n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657,
         n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667,
         n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677,
         n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687,
         n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697,
         n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707,
         n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717,
         n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727,
         n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737,
         n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747,
         n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757,
         n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767,
         n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777,
         n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787,
         n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797,
         n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807,
         n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817,
         n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827,
         n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837,
         n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847,
         n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857,
         n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867,
         n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877,
         n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887,
         n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897,
         n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907,
         n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917,
         n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927,
         n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937,
         n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947,
         n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957,
         n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967,
         n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977,
         n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987,
         n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997,
         n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007,
         n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017,
         n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027,
         n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037,
         n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047,
         n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057,
         n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067,
         n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077,
         n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087,
         n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097,
         n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107,
         n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117,
         n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127,
         n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137,
         n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147,
         n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157,
         n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167,
         n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177,
         n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187,
         n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197,
         n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207,
         n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217,
         n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227,
         n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237,
         n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247,
         n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257,
         n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267,
         n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277,
         n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287,
         n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297,
         n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307,
         n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317,
         n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327,
         n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337,
         n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347,
         n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357,
         n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367,
         n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377,
         n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387,
         n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397,
         n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407,
         n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417,
         n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427,
         n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437,
         n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447,
         n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457,
         n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467,
         n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477,
         n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487,
         n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497,
         n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507,
         n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517,
         n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527,
         n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537,
         n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547,
         n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557,
         n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567,
         n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577,
         n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587,
         n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597,
         n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607,
         n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617,
         n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627,
         n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637,
         n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647,
         n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657,
         n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667,
         n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677,
         n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687,
         n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697,
         n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707,
         n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717,
         n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727,
         n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737,
         n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747,
         n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757,
         n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767,
         n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777,
         n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787,
         n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797,
         n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807,
         n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817,
         n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827,
         n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837,
         n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847,
         n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857,
         n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867,
         n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877,
         n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887,
         n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897,
         n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907,
         n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917,
         n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927,
         n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937,
         n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947,
         n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957,
         n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967,
         n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977,
         n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987,
         n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997,
         n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007,
         n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017,
         n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027,
         n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037,
         n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047,
         n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057,
         n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067,
         n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077,
         n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087,
         n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097,
         n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107,
         n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117,
         n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127,
         n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137,
         n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147,
         n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157,
         n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167,
         n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177,
         n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187,
         n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197,
         n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207,
         n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217,
         n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227,
         n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237,
         n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247,
         n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257,
         n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267,
         n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277,
         n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287,
         n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297,
         n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307,
         n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317,
         n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327,
         n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337,
         n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347,
         n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357,
         n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367,
         n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377,
         n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387,
         n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397,
         n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407,
         n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417,
         n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427,
         n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437,
         n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447,
         n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457,
         n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467,
         n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477,
         n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487,
         n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497,
         n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507,
         n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517,
         n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527,
         n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537,
         n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547,
         n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557,
         n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567,
         n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577,
         n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587,
         n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597,
         n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607,
         n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617,
         n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627,
         n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637,
         n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647,
         n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657,
         n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667,
         n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677,
         n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687,
         n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697,
         n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707,
         n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717,
         n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727,
         n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737,
         n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747,
         n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757,
         n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767,
         n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777,
         n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787,
         n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797,
         n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807,
         n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817,
         n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827,
         n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837,
         n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847,
         n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857,
         n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867,
         n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877,
         n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887,
         n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897,
         n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907,
         n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917,
         n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927,
         n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937,
         n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947,
         n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957,
         n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967,
         n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977,
         n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987,
         n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997,
         n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007,
         n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017,
         n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027,
         n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037,
         n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047,
         n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057,
         n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067,
         n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077,
         n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087,
         n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097,
         n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107,
         n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117,
         n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127,
         n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137,
         n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147,
         n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157,
         n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167,
         n7168, n7169, n7170, n7171, n7172, n7173, n7175, n7176, n7177, n7178,
         n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188,
         n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198,
         n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208,
         n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218,
         n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228,
         n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238,
         n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248,
         n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258,
         n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268,
         n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278,
         n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288,
         n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298,
         n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308,
         n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318,
         n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328,
         n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338,
         n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348,
         n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358,
         n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368,
         n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378,
         n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388,
         n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398,
         n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408,
         n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418,
         n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428,
         n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438,
         n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448,
         n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458,
         n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468,
         n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478,
         n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488,
         n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498,
         n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508,
         n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518,
         n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528,
         n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538,
         n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548,
         n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558,
         n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568,
         n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578,
         n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588,
         n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598,
         n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608,
         n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618,
         n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628,
         n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638,
         n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648,
         n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658,
         n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668,
         n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678,
         n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688,
         n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698,
         n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708,
         n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718,
         n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728,
         n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738,
         n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748,
         n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758,
         n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768,
         n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778,
         n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788,
         n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798,
         n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808,
         n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818,
         n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828,
         n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838,
         n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848,
         n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858,
         n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868,
         n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878,
         n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888,
         n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898,
         n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908,
         n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918,
         n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928,
         n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938,
         n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948,
         n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958,
         n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968,
         n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978,
         n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988,
         n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998,
         n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008,
         n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018,
         n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028,
         n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038,
         n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048,
         n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058,
         n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068,
         n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078,
         n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088,
         n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098,
         n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108,
         n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118,
         n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128,
         n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138,
         n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148,
         n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158,
         n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168,
         n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178,
         n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188,
         n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198,
         n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208,
         n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218,
         n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228,
         n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238,
         n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248,
         n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258,
         n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268,
         n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278,
         n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288,
         n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298,
         n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308,
         n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318,
         n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328,
         n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338,
         n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348,
         n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358,
         n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368,
         n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378,
         n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388,
         n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398,
         n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408,
         n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418,
         n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428,
         n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438,
         n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448,
         n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458,
         n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468,
         n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478,
         n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488,
         n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498,
         n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508,
         n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518,
         n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528,
         n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538,
         n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548,
         n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558,
         n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568,
         n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578,
         n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588,
         n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598,
         n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608,
         n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618,
         n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628,
         n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638,
         n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648,
         n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658,
         n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668,
         n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678,
         n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688,
         n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698,
         n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708,
         n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718,
         n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728,
         n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738,
         n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748,
         n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758,
         n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768,
         n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778,
         n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788,
         n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798,
         n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808,
         n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818,
         n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828,
         n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838,
         n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848,
         n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858,
         n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868,
         n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878,
         n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888,
         n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898,
         n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908,
         n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918,
         n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928,
         n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938,
         n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948,
         n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958,
         n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968,
         n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978,
         n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988,
         n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998,
         n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008,
         n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018,
         n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028,
         n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038,
         n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048,
         n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058,
         n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068,
         n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078,
         n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088,
         n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098,
         n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108,
         n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118,
         n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128,
         n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138,
         n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148,
         n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158,
         n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168,
         n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178,
         n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188,
         n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198,
         n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208,
         n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218,
         n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228,
         n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238,
         n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248,
         n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258,
         n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268,
         n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278,
         n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288,
         n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298,
         n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308,
         n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318,
         n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328,
         n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338,
         n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348,
         n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358,
         n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368,
         n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378,
         n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388,
         n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398,
         n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408,
         n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418,
         n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428,
         n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438,
         n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448,
         n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458,
         n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468,
         n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478,
         n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488,
         n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498,
         n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508,
         n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518,
         n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528,
         n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538,
         n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548,
         n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558,
         n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568,
         n9569, n9570, n9571, n9572, n9573, n9574, n9576, n9577, n9578, n9579,
         n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589,
         n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599,
         n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609,
         n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619,
         n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629,
         n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639,
         n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649,
         n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659,
         n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669,
         n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679,
         n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689,
         n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699,
         n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709,
         n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719,
         n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729,
         n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739,
         n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749,
         n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759,
         n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769,
         n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779,
         n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789,
         n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799,
         n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809,
         n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819,
         n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829,
         n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839,
         n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849,
         n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859,
         n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869,
         n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879,
         n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889,
         n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899,
         n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909,
         n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919,
         n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929,
         n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939,
         n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949,
         n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959,
         n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969,
         n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979,
         n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989,
         n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999,
         n10000, n10001, n10002, n10003, n10004, n10005, n10006, n10007,
         n10008, n10009, n10010, n10011, n10012, n10013, n10014, n10015,
         n10016, n10017, n10018, n10019, n10020, n10021, n10022, n10023,
         n10024, n10025, n10026, n10027, n10028, n10029, n10030, n10031,
         n10032, n10033, n10034, n10035, n10036, n10037, n10038, n10039,
         n10040, n10041, n10042, n10043, n10044, n10045, n10046, n10047,
         n10048, n10049, n10050, n10051, n10052, n10053, n10054, n10055,
         n10056, n10057, n10058, n10059, n10060, n10061, n10062, n10063,
         n10064, n10065, n10066, n10067, n10068, n10069, n10070, n10071;

  INV_X1 U4763 ( .A(n4259), .ZN(n7690) );
  INV_X4 U4764 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3152) );
  BUF_X1 U4765 ( .A(n5850), .Z(n5856) );
  CLKBUF_X2 U4766 ( .A(n6003), .Z(n8824) );
  BUF_X2 U4767 ( .A(n6069), .Z(n6582) );
  BUF_X2 U4768 ( .A(n5062), .Z(n5474) );
  INV_X1 U4769 ( .A(n6584), .ZN(n6087) );
  INV_X1 U4770 ( .A(n6575), .ZN(n4392) );
  NOR2_X1 U4771 ( .A1(P1_IR_REG_6__SCAN_IN), .A2(P1_IR_REG_10__SCAN_IN), .ZN(
        n5918) );
  AND2_X1 U4772 ( .A1(P2_REG2_REG_8__SCAN_IN), .A2(n7292), .ZN(n4258) );
  NOR2_X1 U4773 ( .A1(n4258), .A2(n7291), .ZN(n7294) );
  NAND2_X2 U4775 ( .A1(n7763), .A2(n4401), .ZN(n7765) );
  OAI21_X1 U4776 ( .B1(n8084), .B2(P2_REG2_REG_14__SCAN_IN), .A(n8083), .ZN(
        n8104) );
  INV_X1 U4777 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n5205) );
  NOR2_X1 U4778 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P1_IR_REG_20__SCAN_IN), .ZN(
        n5928) );
  NOR2_X1 U4779 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_11__SCAN_IN), .ZN(
        n5916) );
  OR2_X1 U4780 ( .A1(n5749), .A2(P2_IR_REG_27__SCAN_IN), .ZN(n4982) );
  OR2_X1 U4781 ( .A1(n5752), .A2(n5590), .ZN(n5722) );
  INV_X2 U4782 ( .A(n6045), .ZN(n6499) );
  AND3_X1 U4783 ( .A1(n6259), .A2(n5920), .A3(n5919), .ZN(n5931) );
  AND3_X1 U4784 ( .A1(n5918), .A2(n5917), .A3(n5916), .ZN(n4878) );
  NOR2_X1 U4785 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_4__SCAN_IN), .ZN(
        n5914) );
  CLKBUF_X2 U4786 ( .A(n5771), .Z(n5850) );
  AND3_X1 U4787 ( .A1(n4972), .A2(n4971), .A3(n4970), .ZN(n5251) );
  OR2_X1 U4788 ( .A1(n9477), .A2(n7900), .ZN(n9050) );
  OR2_X1 U4789 ( .A1(n5968), .A2(n5960), .ZN(n5970) );
  NAND2_X1 U4791 ( .A1(n4999), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n5162) );
  INV_X1 U4792 ( .A(n7207), .ZN(n5587) );
  OR2_X1 U4793 ( .A1(n4264), .A2(n9222), .ZN(n6432) );
  INV_X1 U4794 ( .A(n9225), .ZN(n9466) );
  NAND2_X1 U4795 ( .A1(n5970), .A2(n5969), .ZN(n6640) );
  INV_X1 U4796 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n6472) );
  NOR2_X1 U4797 ( .A1(n8178), .A2(n8444), .ZN(n8172) );
  XNOR2_X1 U4798 ( .A(n4994), .B(P2_IR_REG_29__SCAN_IN), .ZN(n5002) );
  AND4_X1 U4799 ( .A1(n6095), .A2(n6094), .A3(n6093), .A4(n6092), .ZN(n7615)
         );
  AND2_X1 U4800 ( .A1(n6425), .A2(n6424), .ZN(n9225) );
  INV_X1 U4801 ( .A(n7354), .ZN(n9115) );
  INV_X2 U4802 ( .A(n9713), .ZN(n9716) );
  NAND2_X2 U4803 ( .A1(n9697), .A2(n7375), .ZN(n9713) );
  NAND2_X2 U4804 ( .A1(n7017), .A2(n7173), .ZN(n7116) );
  XNOR2_X2 U4806 ( .A(n9144), .B(n4420), .ZN(n7274) );
  NAND2_X2 U4807 ( .A1(n4266), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n5980) );
  NAND2_X2 U4808 ( .A1(n8421), .A2(n8434), .ZN(n5241) );
  OAI21_X2 U4809 ( .B1(n7739), .B2(n7745), .A(n5221), .ZN(n8421) );
  OR2_X1 U4810 ( .A1(n8239), .A2(n4995), .ZN(n5465) );
  NAND3_X1 U4811 ( .A1(n4815), .A2(n4814), .A3(n6943), .ZN(n7058) );
  NAND2_X2 U4812 ( .A1(n8883), .A2(n8882), .ZN(n8892) );
  INV_X2 U4813 ( .A(n5948), .ZN(n7856) );
  AOI21_X2 U4814 ( .B1(n8328), .B2(n8327), .A(n7833), .ZN(n8314) );
  INV_X2 U4815 ( .A(n5951), .ZN(n9570) );
  NAND2_X2 U4816 ( .A1(n7638), .A2(n5659), .ZN(n7739) );
  AOI21_X2 U4817 ( .B1(n5193), .B2(n5198), .A(n4381), .ZN(n5223) );
  NAND3_X2 U4818 ( .A1(n4553), .A2(n4552), .A3(n4556), .ZN(n7886) );
  OAI21_X2 U4819 ( .B1(n9414), .B2(n9413), .A(n8893), .ZN(n9394) );
  XNOR2_X2 U4820 ( .A(n5077), .B(P2_IR_REG_4__SCAN_IN), .ZN(n6832) );
  OR2_X4 U4821 ( .A1(n7478), .A2(n6541), .ZN(n4282) );
  XNOR2_X2 U4822 ( .A(n4879), .B(P1_IR_REG_30__SCAN_IN), .ZN(n5948) );
  XNOR2_X2 U4823 ( .A(n5058), .B(P2_IR_REG_2__SCAN_IN), .ZN(n6806) );
  XNOR2_X2 U4824 ( .A(n5556), .B(n5555), .ZN(n7207) );
  OAI22_X2 U4825 ( .A1(n7886), .A2(n7885), .B1(n9477), .B2(n9268), .ZN(n9233)
         );
  NAND2_X2 U4826 ( .A1(n4618), .A2(n5057), .ZN(n6737) );
  AND2_X1 U4827 ( .A1(n4462), .A2(n4460), .ZN(n4294) );
  NAND2_X1 U4828 ( .A1(n4259), .A2(n4406), .ZN(n7729) );
  OAI21_X1 U4829 ( .B1(n7335), .B2(n6083), .A(n7333), .ZN(n6086) );
  OAI211_X1 U4830 ( .C1(n7508), .C2(n9066), .A(n7507), .B(n7506), .ZN(n7583)
         );
  AND4_X1 U4831 ( .A1(n6382), .A2(n6381), .A3(n6380), .A4(n6379), .ZN(n8833)
         );
  NAND2_X1 U4832 ( .A1(n7184), .A2(n9846), .ZN(n7423) );
  NAND2_X1 U4833 ( .A1(n7247), .A2(n5625), .ZN(n7214) );
  OR2_X1 U4834 ( .A1(n6480), .A2(n6522), .ZN(n9101) );
  NAND2_X2 U4836 ( .A1(n7366), .A2(n8987), .ZN(n9058) );
  INV_X2 U4837 ( .A(n5722), .ZN(n5715) );
  NAND4_X1 U4838 ( .A1(n5055), .A2(n5054), .A3(n5053), .A4(n5052), .ZN(n8066)
         );
  INV_X8 U4839 ( .A(n4282), .ZN(n4260) );
  INV_X1 U4840 ( .A(n9689), .ZN(n4261) );
  XNOR2_X1 U4841 ( .A(n5943), .B(n5942), .ZN(n5975) );
  NAND2_X1 U4842 ( .A1(n5752), .A2(n5587), .ZN(n7029) );
  BUF_X2 U4843 ( .A(n5098), .Z(n5537) );
  NAND2_X1 U4844 ( .A1(n5925), .A2(n5941), .ZN(n9091) );
  INV_X2 U4845 ( .A(n7458), .ZN(n9690) );
  XNOR2_X1 U4847 ( .A(n5926), .B(n6473), .ZN(n8938) );
  NAND2_X1 U4848 ( .A1(n6575), .A2(P1_U3084), .ZN(n9576) );
  AND2_X2 U4849 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n6052) );
  OR2_X1 U4850 ( .A1(n4423), .A2(n8704), .ZN(n4422) );
  AND3_X1 U4851 ( .A1(n4521), .A2(n4584), .A3(n7852), .ZN(n4363) );
  AND2_X1 U4852 ( .A1(n4880), .A2(n4288), .ZN(n9205) );
  AOI21_X1 U4853 ( .B1(n8244), .B2(n4796), .A(n4793), .ZN(n8224) );
  NAND2_X1 U4854 ( .A1(n8259), .A2(n7836), .ZN(n8244) );
  NAND2_X1 U4855 ( .A1(n4741), .A2(n4747), .ZN(n8744) );
  NAND2_X1 U4856 ( .A1(n8247), .A2(n8246), .ZN(n8245) );
  NAND2_X1 U4857 ( .A1(n5528), .A2(n5527), .ZN(n8444) );
  OAI21_X1 U4858 ( .B1(n4294), .B2(n8997), .A(n9050), .ZN(n9240) );
  OR2_X1 U4859 ( .A1(n5827), .A2(n4828), .ZN(n4827) );
  NAND2_X1 U4860 ( .A1(n8694), .A2(n6291), .ZN(n8635) );
  AND2_X2 U4861 ( .A1(n8286), .A2(n4649), .ZN(n8225) );
  NAND2_X1 U4862 ( .A1(n8818), .A2(n8817), .ZN(n9198) );
  NAND2_X2 U4863 ( .A1(n6483), .A2(n6482), .ZN(n9455) );
  OR2_X2 U4864 ( .A1(n9466), .A2(n7901), .ZN(n9047) );
  AND2_X1 U4865 ( .A1(n4820), .A2(n7948), .ZN(n4816) );
  CLKBUF_X1 U4866 ( .A(n8392), .Z(n8435) );
  NOR2_X1 U4867 ( .A1(n9298), .A2(n4898), .ZN(n4897) );
  NAND2_X1 U4868 ( .A1(n6408), .A2(n6407), .ZN(n9472) );
  NAND2_X1 U4869 ( .A1(n4646), .A2(n4645), .ZN(n7747) );
  OR2_X2 U4870 ( .A1(n9487), .A2(n8652), .ZN(n9057) );
  OAI211_X2 U4871 ( .C1(n7446), .C2(n4833), .A(n4831), .B(n4830), .ZN(n7625)
         );
  INV_X1 U4872 ( .A(n7729), .ZN(n4646) );
  AND2_X1 U4873 ( .A1(n8942), .A2(n8981), .ZN(n9322) );
  OR2_X1 U4874 ( .A1(n7585), .A2(n4448), .ZN(n4450) );
  NAND2_X1 U4875 ( .A1(n6329), .A2(n6328), .ZN(n9498) );
  AND2_X1 U4876 ( .A1(n4449), .A2(n8874), .ZN(n4454) );
  AND2_X1 U4877 ( .A1(n5566), .A2(n5642), .ZN(n7646) );
  INV_X1 U4878 ( .A(n7897), .ZN(n9524) );
  NAND2_X1 U4879 ( .A1(n5284), .A2(n5283), .ZN(n8509) );
  NOR2_X1 U4880 ( .A1(n4616), .A2(n7716), .ZN(n4615) );
  NAND2_X1 U4881 ( .A1(n4822), .A2(n4310), .ZN(n7300) );
  NAND2_X1 U4882 ( .A1(n5159), .A2(n5158), .ZN(n8546) );
  NAND2_X1 U4883 ( .A1(n7515), .A2(n8868), .ZN(n7585) );
  AND2_X1 U4884 ( .A1(n5650), .A2(n7724), .ZN(n7694) );
  NAND2_X1 U4885 ( .A1(n5184), .A2(n5183), .ZN(n8529) );
  OR2_X1 U4886 ( .A1(n7469), .A2(n7468), .ZN(n4622) );
  INV_X1 U4887 ( .A(n8833), .ZN(n9287) );
  NAND2_X1 U4888 ( .A1(n6130), .A2(n6129), .ZN(n8720) );
  NAND2_X1 U4889 ( .A1(n5012), .A2(n5011), .ZN(n8540) );
  OAI21_X1 U4890 ( .B1(n7182), .B2(n5123), .A(n5635), .ZN(n5124) );
  NAND2_X1 U4891 ( .A1(n5285), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n5321) );
  INV_X2 U4892 ( .A(n9798), .ZN(n4262) );
  INV_X1 U4893 ( .A(n7423), .ZN(n4644) );
  AND2_X2 U4894 ( .A1(n8771), .A2(n9398), .ZN(n8808) );
  XNOR2_X1 U4895 ( .A(n5152), .B(n5151), .ZN(n6604) );
  NAND2_X1 U4896 ( .A1(n6115), .A2(n6114), .ZN(n7620) );
  INV_X4 U4897 ( .A(n6081), .ZN(n6497) );
  NAND2_X1 U4898 ( .A1(n6078), .A2(n6077), .ZN(n7358) );
  AOI21_X1 U4899 ( .B1(n7021), .B2(n5774), .A(n5761), .ZN(n6925) );
  INV_X1 U4900 ( .A(n7141), .ZN(n4407) );
  XNOR2_X1 U4901 ( .A(n5094), .B(n5093), .ZN(n6579) );
  NAND2_X1 U4902 ( .A1(n4445), .A2(n4446), .ZN(n4693) );
  INV_X2 U4903 ( .A(n5774), .ZN(n6869) );
  NAND2_X1 U4904 ( .A1(n4261), .A2(n6894), .ZN(n7484) );
  NAND2_X1 U4905 ( .A1(n4663), .A2(n4939), .ZN(n5088) );
  INV_X1 U4906 ( .A(n9114), .ZN(n9676) );
  NAND2_X1 U4907 ( .A1(n5032), .A2(n5031), .ZN(n7077) );
  NAND4_X1 U4908 ( .A1(n5087), .A2(n5086), .A3(n5085), .A4(n5084), .ZN(n8063)
         );
  INV_X1 U4909 ( .A(n6868), .ZN(n4263) );
  AND4_X1 U4910 ( .A1(n6075), .A2(n6074), .A3(n6073), .A4(n6072), .ZN(n7357)
         );
  NAND2_X1 U4911 ( .A1(n7478), .A2(n6506), .ZN(n6045) );
  NAND4_X1 U4912 ( .A1(n6059), .A2(n6058), .A3(n6057), .A4(n6056), .ZN(n9114)
         );
  NAND4_X1 U4913 ( .A1(n6018), .A2(n6017), .A3(n6016), .A4(n6015), .ZN(n9116)
         );
  BUF_X1 U4914 ( .A(n5554), .Z(n5755) );
  CLKBUF_X1 U4915 ( .A(n5586), .Z(n5752) );
  INV_X1 U4916 ( .A(n5102), .ZN(n4995) );
  CLKBUF_X3 U4917 ( .A(n6055), .Z(n6116) );
  NAND2_X2 U4918 ( .A1(n5948), .A2(n9570), .ZN(n6051) );
  MUX2_X1 U4919 ( .A(P1_IR_REG_0__SCAN_IN), .B(n9577), .S(n6640), .Z(n7458) );
  CLKBUF_X3 U4920 ( .A(n6053), .Z(n4264) );
  XNOR2_X1 U4921 ( .A(n5944), .B(n6474), .ZN(n9694) );
  NAND2_X2 U4922 ( .A1(P1_U3084), .A2(n4392), .ZN(n9572) );
  XNOR2_X1 U4923 ( .A(n4945), .B(SI_7_), .ZN(n5109) );
  NAND2_X1 U4924 ( .A1(n5948), .A2(n5951), .ZN(n6053) );
  NOR2_X1 U4925 ( .A1(n6731), .A2(n4314), .ZN(n6803) );
  XNOR2_X1 U4926 ( .A(n4992), .B(P2_IR_REG_30__SCAN_IN), .ZN(n7912) );
  OAI21_X1 U4927 ( .B1(n6277), .B2(n4775), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n5926) );
  XNOR2_X1 U4928 ( .A(n4943), .B(SI_6_), .ZN(n5093) );
  NAND2_X1 U4929 ( .A1(n5534), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5556) );
  NAND2_X2 U4930 ( .A1(n6575), .A2(P2_U3152), .ZN(n8583) );
  NAND2_X1 U4931 ( .A1(n6117), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n6152) );
  AND3_X1 U4932 ( .A1(n5555), .A2(n5558), .A3(n5738), .ZN(n4979) );
  AND2_X1 U4933 ( .A1(n4974), .A2(n4973), .ZN(n5279) );
  AND3_X1 U4934 ( .A1(n5961), .A2(n6513), .A3(n5927), .ZN(n4908) );
  INV_X4 U4935 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3084) );
  INV_X1 U4936 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n5558) );
  NOR2_X1 U4937 ( .A1(P1_IR_REG_16__SCAN_IN), .A2(P1_IR_REG_12__SCAN_IN), .ZN(
        n5920) );
  NOR2_X1 U4938 ( .A1(P1_IR_REG_2__SCAN_IN), .A2(P1_IR_REG_5__SCAN_IN), .ZN(
        n5913) );
  NOR2_X1 U4939 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5915) );
  NOR2_X1 U4940 ( .A1(P2_IR_REG_11__SCAN_IN), .A2(P2_IR_REG_15__SCAN_IN), .ZN(
        n4971) );
  INV_X1 U4941 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n5738) );
  NOR2_X1 U4942 ( .A1(P2_IR_REG_9__SCAN_IN), .A2(P2_IR_REG_8__SCAN_IN), .ZN(
        n4972) );
  NOR2_X1 U4943 ( .A1(P2_IR_REG_16__SCAN_IN), .A2(P2_IR_REG_6__SCAN_IN), .ZN(
        n4973) );
  NOR2_X2 U4944 ( .A1(P1_IR_REG_26__SCAN_IN), .A2(P1_IR_REG_25__SCAN_IN), .ZN(
        n6513) );
  NAND2_X2 U4945 ( .A1(n7448), .A2(n7447), .ZN(n7446) );
  AOI21_X2 U4946 ( .B1(n7725), .B2(n5172), .A(n5171), .ZN(n7639) );
  AND2_X2 U4947 ( .A1(n7388), .A2(n9762), .ZN(n7591) );
  AND3_X4 U4948 ( .A1(n5065), .A2(n5064), .A3(n5063), .ZN(n7124) );
  NOR2_X2 U4949 ( .A1(n5162), .A2(n4313), .ZN(n5013) );
  NAND2_X1 U4950 ( .A1(n8961), .A2(n4307), .ZN(n7596) );
  AOI22_X2 U4951 ( .A1(n8314), .A2(n7834), .B1(n8307), .B2(n8318), .ZN(n8295)
         );
  INV_X1 U4952 ( .A(n6640), .ZN(n4265) );
  MUX2_X2 U4953 ( .A(n8881), .B(n8880), .S(n8925), .Z(n8883) );
  OAI21_X1 U4954 ( .B1(n4865), .B2(n4583), .A(n8199), .ZN(n4582) );
  AOI21_X1 U4955 ( .B1(n4868), .B2(n7839), .A(n4866), .ZN(n4865) );
  INV_X1 U4956 ( .A(n6051), .ZN(n4266) );
  AND2_X2 U4957 ( .A1(n7258), .A2(n9842), .ZN(n7184) );
  AND2_X1 U4958 ( .A1(n7912), .A2(n8585), .ZN(n5098) );
  NAND2_X2 U4959 ( .A1(n6052), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n6090) );
  OAI21_X2 U4960 ( .B1(n5603), .B2(n7066), .A(n5607), .ZN(n7078) );
  NOR2_X4 U4961 ( .A1(n7439), .A2(n8552), .ZN(n7570) );
  INV_X1 U4962 ( .A(n7163), .ZN(n4647) );
  INV_X1 U4963 ( .A(n5526), .ZN(n5056) );
  XNOR2_X2 U4964 ( .A(n9205), .B(n9204), .ZN(n9465) );
  INV_X1 U4965 ( .A(n4566), .ZN(n4565) );
  OR2_X1 U4966 ( .A1(n6897), .A2(n6896), .ZN(n4446) );
  NOR2_X2 U4967 ( .A1(n6265), .A2(n9972), .ZN(n6282) );
  OR2_X2 U4968 ( .A1(n8430), .A2(n8512), .ZN(n4269) );
  NAND4_X4 U4969 ( .A1(n5983), .A2(n5982), .A3(n5981), .A4(n5980), .ZN(n6890)
         );
  NAND2_X1 U4970 ( .A1(n5549), .A2(n4392), .ZN(n5526) );
  NAND2_X1 U4971 ( .A1(n6893), .A2(n6894), .ZN(n8987) );
  OR2_X1 U4972 ( .A1(n6893), .A2(n6894), .ZN(n7366) );
  INV_X2 U4974 ( .A(n7162), .ZN(n9791) );
  NAND2_X1 U4975 ( .A1(n8064), .A2(n9829), .ZN(n7247) );
  NAND2_X1 U4976 ( .A1(n4407), .A2(n9829), .ZN(n7255) );
  OAI22_X2 U4977 ( .A1(n9393), .A2(n7874), .B1(n7897), .B2(n9418), .ZN(n9375)
         );
  NAND2_X1 U4978 ( .A1(n5951), .A2(n7856), .ZN(n6055) );
  NOR2_X2 U4979 ( .A1(n6311), .A2(n10029), .ZN(n6330) );
  OR2_X2 U4980 ( .A1(n6297), .A2(n6296), .ZN(n6311) );
  NAND2_X1 U4981 ( .A1(n8901), .A2(n4284), .ZN(n8907) );
  OR2_X1 U4982 ( .A1(n4690), .A2(n8915), .ZN(n4685) );
  NOR2_X1 U4983 ( .A1(n8923), .A2(n9011), .ZN(n8919) );
  INV_X1 U4984 ( .A(n5593), .ZN(n4870) );
  AND2_X1 U4985 ( .A1(n9089), .A2(n9433), .ZN(n8923) );
  OR2_X1 U4986 ( .A1(n8466), .A2(n7974), .ZN(n5593) );
  OAI21_X1 U4987 ( .B1(n5450), .B2(n5449), .A(n5448), .ZN(n5467) );
  AND2_X1 U4988 ( .A1(n5417), .A2(n5403), .ZN(n5415) );
  AND2_X1 U4989 ( .A1(n8476), .A2(n8266), .ZN(n7835) );
  OR2_X1 U4990 ( .A1(n6084), .A2(n7332), .ZN(n6085) );
  NOR2_X1 U4991 ( .A1(n9472), .A2(n7887), .ZN(n7888) );
  INV_X1 U4992 ( .A(n7884), .ZN(n4895) );
  NAND2_X1 U4993 ( .A1(n4883), .A2(n4882), .ZN(n9450) );
  AND2_X1 U4994 ( .A1(n9085), .A2(n4884), .ZN(n4882) );
  OR2_X1 U4995 ( .A1(n8907), .A2(n8906), .ZN(n4416) );
  NOR2_X1 U4996 ( .A1(n4388), .A2(n9308), .ZN(n4387) );
  NAND2_X1 U4997 ( .A1(n4390), .A2(n4389), .ZN(n4388) );
  INV_X1 U4998 ( .A(n9285), .ZN(n4389) );
  AND2_X1 U4999 ( .A1(n4333), .A2(n9298), .ZN(n4390) );
  NAND3_X1 U5000 ( .A1(n8919), .A2(n8920), .A3(n8918), .ZN(n8929) );
  NAND2_X1 U5001 ( .A1(n5308), .A2(n5307), .ZN(n5353) );
  INV_X1 U5002 ( .A(n5306), .ZN(n5307) );
  INV_X1 U5003 ( .A(n5204), .ZN(n4381) );
  NAND2_X1 U5004 ( .A1(n4948), .A2(n4947), .ZN(n5139) );
  NAND2_X1 U5005 ( .A1(n4507), .A2(n4506), .ZN(n4510) );
  NAND2_X1 U5006 ( .A1(n7625), .A2(n4505), .ZN(n4507) );
  AND2_X1 U5007 ( .A1(n7811), .A2(n4296), .ZN(n4505) );
  INV_X1 U5008 ( .A(n7766), .ZN(n4640) );
  OR2_X1 U5009 ( .A1(n8274), .A2(n7940), .ZN(n5700) );
  AND2_X1 U5010 ( .A1(n8282), .A2(n5695), .ZN(n4849) );
  NOR2_X1 U5011 ( .A1(n8498), .A2(n8502), .ZN(n4659) );
  OR2_X1 U5012 ( .A1(n8517), .A2(n8403), .ZN(n5669) );
  OR2_X1 U5013 ( .A1(n7751), .A2(n8424), .ZN(n7821) );
  OR2_X1 U5014 ( .A1(n8535), .A2(n7993), .ZN(n5170) );
  NAND2_X1 U5015 ( .A1(n4501), .A2(n7219), .ZN(n5633) );
  OR2_X1 U5016 ( .A1(n7219), .A2(n4501), .ZN(n5627) );
  AND2_X1 U5017 ( .A1(n5752), .A2(n5755), .ZN(n5885) );
  NAND2_X1 U5018 ( .A1(n4263), .A2(n4647), .ZN(n5567) );
  OR2_X1 U5019 ( .A1(n8189), .A2(n8203), .ZN(n5716) );
  INV_X1 U5020 ( .A(n6258), .ZN(n4729) );
  OR2_X1 U5021 ( .A1(n6290), .A2(n6289), .ZN(n6291) );
  NOR2_X1 U5022 ( .A1(n4600), .A2(n4597), .ZN(n4596) );
  INV_X1 U5023 ( .A(n4555), .ZN(n4554) );
  OAI21_X1 U5024 ( .B1(n4894), .B2(n4272), .A(n4325), .ZN(n4555) );
  NAND2_X1 U5025 ( .A1(n9309), .A2(n4463), .ZN(n4462) );
  AND2_X1 U5026 ( .A1(n9384), .A2(n4710), .ZN(n4709) );
  NOR2_X1 U5027 ( .A1(n8844), .A2(n4712), .ZN(n4711) );
  INV_X1 U5028 ( .A(n8951), .ZN(n4712) );
  AND2_X1 U5029 ( .A1(n7897), .A2(n9387), .ZN(n8845) );
  NAND2_X1 U5030 ( .A1(n5523), .A2(n5524), .ZN(n5544) );
  OAI21_X1 U5031 ( .B1(n5434), .B2(n5433), .A(n5432), .ZN(n5450) );
  AND2_X1 U5032 ( .A1(n4960), .A2(n4957), .ZN(n4909) );
  XNOR2_X1 U5033 ( .A(n4940), .B(SI_5_), .ZN(n5089) );
  NAND2_X1 U5034 ( .A1(n4329), .A2(n4848), .ZN(n4843) );
  NAND2_X1 U5035 ( .A1(n7957), .A2(n5815), .ZN(n4847) );
  NAND2_X1 U5036 ( .A1(n7980), .A2(n7981), .ZN(n5827) );
  BUF_X1 U5037 ( .A(n5045), .Z(n5080) );
  AOI21_X1 U5038 ( .B1(n8253), .B2(n5514), .A(n5447), .ZN(n7974) );
  AND2_X1 U5039 ( .A1(n7912), .A2(n5002), .ZN(n5102) );
  OR2_X1 U5040 ( .A1(n7764), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n4401) );
  AOI21_X1 U5041 ( .B1(n8161), .B2(n8167), .A(n5587), .ZN(n4632) );
  NOR2_X1 U5042 ( .A1(n8450), .A2(n8049), .ZN(n8182) );
  NAND2_X1 U5043 ( .A1(n4805), .A2(n4803), .ZN(n8259) );
  NOR2_X1 U5044 ( .A1(n4806), .A2(n4804), .ZN(n4803) );
  OR2_X1 U5045 ( .A1(n8482), .A2(n8322), .ZN(n4811) );
  OR2_X1 U5046 ( .A1(n8482), .A2(n7916), .ZN(n5695) );
  OR2_X1 U5047 ( .A1(n8347), .A2(n7983), .ZN(n4906) );
  NOR2_X1 U5048 ( .A1(n4786), .A2(n4783), .ZN(n4782) );
  OR2_X1 U5049 ( .A1(n8509), .A2(n8405), .ZN(n5597) );
  AND2_X1 U5050 ( .A1(n8512), .A2(n8426), .ZN(n7826) );
  NOR2_X1 U5051 ( .A1(n7743), .A2(n4802), .ZN(n4801) );
  INV_X1 U5052 ( .A(n7652), .ZN(n4802) );
  NAND2_X1 U5053 ( .A1(n7181), .A2(n4303), .ZN(n4498) );
  NAND2_X1 U5054 ( .A1(n4528), .A2(n7262), .ZN(n7213) );
  INV_X1 U5055 ( .A(n8063), .ZN(n4528) );
  INV_X1 U5056 ( .A(n8404), .ZN(n8425) );
  INV_X2 U5057 ( .A(n5549), .ZN(n5315) );
  NAND2_X1 U5058 ( .A1(n5716), .A2(n5717), .ZN(n8185) );
  NAND2_X1 U5059 ( .A1(n7025), .A2(n5875), .ZN(n8553) );
  NAND2_X1 U5060 ( .A1(n7200), .A2(n7199), .ZN(n4756) );
  INV_X1 U5061 ( .A(n4759), .ZN(n4440) );
  AND2_X1 U5062 ( .A1(n6085), .A2(n8732), .ZN(n4437) );
  NAND2_X1 U5063 ( .A1(n4758), .A2(n8732), .ZN(n4439) );
  OAI21_X1 U5064 ( .B1(n4268), .B2(n4759), .A(n4287), .ZN(n4758) );
  OAI21_X1 U5065 ( .B1(n4460), .B2(n9254), .A(n4458), .ZN(n9255) );
  NAND2_X1 U5066 ( .A1(n9309), .A2(n4459), .ZN(n4458) );
  NOR2_X1 U5067 ( .A1(n9254), .A2(n4464), .ZN(n4459) );
  OR2_X1 U5068 ( .A1(n9492), .A2(n7882), .ZN(n9283) );
  AOI21_X1 U5069 ( .B1(n4897), .B2(n7881), .A(n4312), .ZN(n4896) );
  AND2_X1 U5070 ( .A1(n9283), .A2(n9282), .ZN(n9298) );
  NAND2_X1 U5071 ( .A1(n4902), .A2(n4901), .ZN(n4900) );
  AOI21_X1 U5072 ( .B1(n4891), .B2(n4270), .A(n4315), .ZN(n4558) );
  OAI21_X1 U5073 ( .B1(n7664), .B2(n4274), .A(n4298), .ZN(n4546) );
  NOR2_X1 U5074 ( .A1(n9069), .A2(n4274), .ZN(n4547) );
  AND2_X1 U5075 ( .A1(n8939), .A2(n9574), .ZN(n9398) );
  INV_X1 U5076 ( .A(n9706), .ZN(n9416) );
  OR2_X1 U5077 ( .A1(n6890), .A2(n9692), .ZN(n6891) );
  AOI21_X1 U5078 ( .B1(n5975), .B2(n7478), .A(n9169), .ZN(n4724) );
  NAND2_X1 U5079 ( .A1(n6900), .A2(n8937), .ZN(n9706) );
  INV_X1 U5080 ( .A(n9396), .ZN(n9703) );
  AOI21_X1 U5081 ( .B1(n5968), .B2(n5967), .A(n5966), .ZN(n5969) );
  NAND2_X1 U5082 ( .A1(n9564), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4879) );
  NAND2_X1 U5083 ( .A1(n4444), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4443) );
  XNOR2_X1 U5084 ( .A(n5467), .B(n5466), .ZN(n7710) );
  INV_X1 U5085 ( .A(n4674), .ZN(n5416) );
  AOI21_X1 U5086 ( .B1(n4682), .B2(n4675), .A(n4678), .ZN(n4674) );
  NAND2_X1 U5087 ( .A1(n4682), .A2(n5376), .ZN(n5397) );
  OR2_X1 U5088 ( .A1(n6277), .A2(P1_IR_REG_18__SCAN_IN), .ZN(n6476) );
  NAND2_X1 U5089 ( .A1(n4880), .A2(n4302), .ZN(n4883) );
  NAND2_X1 U5090 ( .A1(n5728), .A2(n5568), .ZN(n4532) );
  INV_X1 U5091 ( .A(n7890), .ZN(n9228) );
  NAND2_X1 U5092 ( .A1(n9046), .A2(n9045), .ZN(n9447) );
  NAND2_X1 U5093 ( .A1(n5632), .A2(n4291), .ZN(n4536) );
  NOR2_X1 U5094 ( .A1(n9052), .A2(n4569), .ZN(n4568) );
  INV_X1 U5095 ( .A(n9057), .ZN(n4569) );
  NAND2_X1 U5096 ( .A1(n4416), .A2(n4414), .ZN(n4410) );
  NAND2_X1 U5097 ( .A1(n8843), .A2(n4565), .ZN(n8909) );
  AND2_X1 U5098 ( .A1(n4382), .A2(n4540), .ZN(n4539) );
  AND2_X1 U5099 ( .A1(n8282), .A2(n4322), .ZN(n4540) );
  NOR2_X1 U5100 ( .A1(n8466), .A2(n8274), .ZN(n4653) );
  AND2_X1 U5101 ( .A1(n9080), .A2(n4387), .ZN(n9081) );
  OAI21_X1 U5102 ( .B1(n8922), .B2(n8921), .A(n8929), .ZN(n8926) );
  AND2_X1 U5103 ( .A1(n4669), .A2(n5294), .ZN(n4273) );
  INV_X1 U5104 ( .A(n5271), .ZN(n4666) );
  INV_X1 U5105 ( .A(n5222), .ZN(n4671) );
  AND2_X1 U5106 ( .A1(n4909), .A2(n5141), .ZN(n4907) );
  INV_X1 U5107 ( .A(n4941), .ZN(n4573) );
  NAND3_X1 U5108 ( .A1(n4915), .A2(P1_ADDR_REG_19__SCAN_IN), .A3(
        P2_ADDR_REG_19__SCAN_IN), .ZN(n4488) );
  AND2_X1 U5109 ( .A1(n5853), .A2(n5852), .ZN(n5887) );
  NOR2_X1 U5110 ( .A1(n5592), .A2(n4858), .ZN(n4857) );
  NAND2_X1 U5111 ( .A1(n4862), .A2(n4859), .ZN(n4858) );
  NAND2_X1 U5112 ( .A1(n4860), .A2(n4346), .ZN(n4859) );
  NAND2_X1 U5113 ( .A1(n5719), .A2(n4863), .ZN(n4862) );
  INV_X1 U5114 ( .A(n5718), .ZN(n4379) );
  INV_X1 U5115 ( .A(n4642), .ZN(n4639) );
  AND2_X1 U5116 ( .A1(n4653), .A2(n4652), .ZN(n4651) );
  NOR2_X1 U5117 ( .A1(n5407), .A2(n5406), .ZN(n4398) );
  INV_X1 U5118 ( .A(n4849), .ZN(n4481) );
  NAND2_X1 U5119 ( .A1(n8350), .A2(n4874), .ZN(n4873) );
  INV_X1 U5120 ( .A(n5677), .ZN(n4874) );
  INV_X1 U5121 ( .A(n5690), .ZN(n4872) );
  OR2_X1 U5122 ( .A1(n8492), .A2(n7932), .ZN(n5690) );
  NAND2_X1 U5123 ( .A1(n7831), .A2(n4784), .ZN(n4783) );
  INV_X1 U5124 ( .A(n7829), .ZN(n4784) );
  OR2_X1 U5125 ( .A1(n8498), .A2(n8367), .ZN(n7831) );
  OR2_X1 U5126 ( .A1(n8529), .A2(n7741), .ZN(n5658) );
  OR2_X1 U5127 ( .A1(n8540), .A2(n7627), .ZN(n5650) );
  NAND2_X1 U5128 ( .A1(n7213), .A2(n7135), .ZN(n5614) );
  NAND2_X1 U5129 ( .A1(n8065), .A2(n9821), .ZN(n5623) );
  AOI21_X1 U5130 ( .B1(n4581), .B2(n4583), .A(n4580), .ZN(n4579) );
  NAND2_X1 U5131 ( .A1(n8286), .A2(n4653), .ZN(n8251) );
  NOR2_X1 U5132 ( .A1(n8282), .A2(n4809), .ZN(n4808) );
  INV_X1 U5133 ( .A(n4811), .ZN(n4809) );
  INV_X1 U5134 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n4970) );
  AND2_X1 U5135 ( .A1(n6399), .A2(n6398), .ZN(n6402) );
  NOR2_X1 U5136 ( .A1(n4283), .A2(n4739), .ZN(n4738) );
  INV_X1 U5137 ( .A(n6327), .ZN(n4739) );
  NOR2_X1 U5138 ( .A1(n4749), .A2(n4283), .ZN(n4748) );
  NAND2_X1 U5139 ( .A1(n8744), .A2(n6372), .ZN(n8600) );
  OAI21_X1 U5140 ( .B1(n4596), .B2(n4317), .A(n7231), .ZN(n4593) );
  INV_X1 U5141 ( .A(n4600), .ZN(n4598) );
  NAND2_X1 U5142 ( .A1(n9145), .A2(n9146), .ZN(n9147) );
  NAND2_X1 U5143 ( .A1(n9211), .A2(n4614), .ZN(n4613) );
  AND2_X1 U5144 ( .A1(n4461), .A2(n8950), .ZN(n4460) );
  NAND2_X1 U5145 ( .A1(n6345), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n6363) );
  NAND2_X1 U5146 ( .A1(n7870), .A2(n4549), .ZN(n4548) );
  NOR2_X1 U5147 ( .A1(n4886), .A2(n4320), .ZN(n4885) );
  INV_X1 U5148 ( .A(n7771), .ZN(n4549) );
  OR2_X1 U5149 ( .A1(n7513), .A2(n8760), .ZN(n8877) );
  OR2_X1 U5150 ( .A1(n7620), .A2(n8714), .ZN(n8871) );
  AND2_X1 U5151 ( .A1(n7385), .A2(n7384), .ZN(n7359) );
  OR2_X1 U5152 ( .A1(n7602), .A2(n9676), .ZN(n9016) );
  AND2_X1 U5153 ( .A1(n9016), .A2(n9018), .ZN(n9063) );
  AND2_X1 U5154 ( .A1(n9369), .A2(n9509), .ZN(n9353) );
  AND2_X1 U5155 ( .A1(n5484), .A2(n5473), .ZN(n5482) );
  AOI21_X1 U5156 ( .B1(n4680), .B2(n5395), .A(n4677), .ZN(n4676) );
  NAND2_X1 U5157 ( .A1(n4564), .A2(n5267), .ZN(n5243) );
  NAND2_X1 U5158 ( .A1(n5223), .A2(n5222), .ZN(n4564) );
  NAND2_X1 U5159 ( .A1(n5193), .A2(n5194), .ZN(n5174) );
  NAND2_X1 U5160 ( .A1(n4662), .A2(n4946), .ZN(n5126) );
  INV_X1 U5161 ( .A(n4826), .ZN(n4825) );
  OAI21_X1 U5162 ( .B1(n4828), .B2(n5826), .A(n5835), .ZN(n4826) );
  OR3_X1 U5163 ( .A1(n5490), .A2(n5489), .A3(n5488), .ZN(n5510) );
  NAND2_X1 U5164 ( .A1(n7029), .A2(n4492), .ZN(n4493) );
  NOR2_X1 U5165 ( .A1(n7017), .A2(n5755), .ZN(n4492) );
  INV_X1 U5166 ( .A(n4837), .ZN(n4832) );
  NAND2_X1 U5167 ( .A1(n5796), .A2(n5797), .ZN(n4837) );
  NAND2_X1 U5168 ( .A1(n4514), .A2(n4818), .ZN(n4820) );
  AOI21_X1 U5169 ( .B1(n5806), .B2(n5804), .A(n8030), .ZN(n4818) );
  NAND2_X1 U5170 ( .A1(n4510), .A2(n5806), .ZN(n4514) );
  NOR2_X1 U5171 ( .A1(n7131), .A2(n5766), .ZN(n5768) );
  INV_X1 U5172 ( .A(n5774), .ZN(n5766) );
  XNOR2_X1 U5173 ( .A(n5771), .B(n7077), .ZN(n5767) );
  NAND2_X1 U5174 ( .A1(n4843), .A2(n5822), .ZN(n4842) );
  AND2_X1 U5175 ( .A1(n4848), .A2(n5815), .ZN(n4845) );
  NAND2_X1 U5176 ( .A1(n5384), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n5407) );
  INV_X1 U5177 ( .A(n5385), .ZN(n5384) );
  NAND2_X1 U5178 ( .A1(n4829), .A2(n4520), .ZN(n4519) );
  INV_X1 U5179 ( .A(n7936), .ZN(n4520) );
  NAND3_X1 U5180 ( .A1(n5846), .A2(n5845), .A3(n4342), .ZN(n4518) );
  NAND2_X1 U5181 ( .A1(n4396), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n5260) );
  INV_X1 U5182 ( .A(n5234), .ZN(n4396) );
  AND2_X1 U5183 ( .A1(n5428), .A2(n5427), .ZN(n7940) );
  INV_X1 U5184 ( .A(n5537), .ZN(n5494) );
  AND4_X1 U5185 ( .A1(n5006), .A2(n5005), .A3(n5004), .A4(n5003), .ZN(n7993)
         );
  AND4_X2 U5186 ( .A1(n5037), .A2(n5036), .A3(n5035), .A4(n5034), .ZN(n6868)
         );
  NAND2_X1 U5187 ( .A1(n5262), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n5037) );
  OAI21_X1 U5188 ( .B1(n6737), .B2(P2_REG1_REG_1__SCAN_IN), .A(n4365), .ZN(
        n6725) );
  NAND2_X1 U5189 ( .A1(n6737), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n4365) );
  AND2_X1 U5190 ( .A1(n7467), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n4623) );
  AND2_X1 U5191 ( .A1(n7793), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n4642) );
  AND2_X1 U5192 ( .A1(n4641), .A2(n4640), .ZN(n7792) );
  INV_X1 U5193 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n4918) );
  NAND2_X1 U5195 ( .A1(n5509), .A2(n5508), .ZN(n8189) );
  NAND2_X1 U5196 ( .A1(n5487), .A2(n5486), .ZN(n8450) );
  NAND2_X1 U5197 ( .A1(n4789), .A2(n4790), .ZN(n8198) );
  AOI21_X1 U5198 ( .B1(n4793), .B2(n4866), .A(n4311), .ZN(n4790) );
  NAND2_X1 U5199 ( .A1(n8244), .A2(n4791), .ZN(n4789) );
  NAND2_X1 U5200 ( .A1(n5457), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n5490) );
  INV_X1 U5201 ( .A(n5459), .ZN(n5457) );
  NAND2_X1 U5202 ( .A1(n4398), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n5442) );
  OR2_X1 U5203 ( .A1(n5442), .A2(n5441), .ZN(n5459) );
  AOI21_X1 U5204 ( .B1(n4480), .B2(n4849), .A(n4323), .ZN(n4479) );
  INV_X1 U5205 ( .A(n5394), .ZN(n4480) );
  OR2_X1 U5206 ( .A1(n8320), .A2(n4481), .ZN(n4475) );
  OR2_X1 U5207 ( .A1(n8295), .A2(n8303), .ZN(n4810) );
  AND2_X1 U5208 ( .A1(n5695), .A2(n5685), .ZN(n8303) );
  NOR2_X1 U5209 ( .A1(n8487), .A2(n4656), .ZN(n4655) );
  INV_X1 U5210 ( .A(n4657), .ZN(n4656) );
  AND2_X1 U5211 ( .A1(n5689), .A2(n8334), .ZN(n8350) );
  AND2_X1 U5212 ( .A1(n7830), .A2(n8373), .ZN(n4788) );
  AND2_X1 U5213 ( .A1(n7830), .A2(n4787), .ZN(n4786) );
  INV_X1 U5214 ( .A(n7827), .ZN(n4787) );
  INV_X1 U5215 ( .A(n7830), .ZN(n8365) );
  OR2_X1 U5216 ( .A1(n8509), .A2(n8366), .ZN(n7827) );
  NAND2_X1 U5217 ( .A1(n8374), .A2(n8373), .ZN(n8372) );
  NAND2_X1 U5218 ( .A1(n8398), .A2(n7823), .ZN(n7824) );
  INV_X1 U5219 ( .A(n8393), .ZN(n7823) );
  AND3_X1 U5220 ( .A1(n5291), .A2(n5290), .A3(n5289), .ZN(n8405) );
  NAND2_X1 U5221 ( .A1(n8428), .A2(n8433), .ZN(n8430) );
  NAND2_X1 U5222 ( .A1(n5212), .A2(n5211), .ZN(n7751) );
  NOR2_X1 U5223 ( .A1(n4800), .A2(n4798), .ZN(n4797) );
  INV_X1 U5224 ( .A(n4500), .ZN(n4496) );
  INV_X1 U5225 ( .A(n5124), .ZN(n7415) );
  NAND2_X1 U5226 ( .A1(n9842), .A2(n4501), .ZN(n4500) );
  NAND2_X1 U5227 ( .A1(n6579), .A2(n5062), .ZN(n4482) );
  NOR2_X1 U5228 ( .A1(P2_IR_REG_28__SCAN_IN), .A2(P2_IR_REG_27__SCAN_IN), .ZN(
        n4877) );
  NAND2_X1 U5229 ( .A1(n4504), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4992) );
  NAND2_X1 U5230 ( .A1(n4327), .A2(n4275), .ZN(n4761) );
  INV_X1 U5231 ( .A(n6143), .ZN(n4764) );
  AND2_X1 U5232 ( .A1(n6502), .A2(n8794), .ZN(n6503) );
  NAND2_X1 U5233 ( .A1(n7103), .A2(n7105), .ZN(n7099) );
  NAND2_X1 U5234 ( .A1(n5993), .A2(n5992), .ZN(n7100) );
  INV_X1 U5235 ( .A(n8723), .ZN(n4751) );
  NOR2_X1 U5236 ( .A1(n6326), .A2(n4341), .ZN(n4749) );
  INV_X1 U5237 ( .A(n4429), .ZN(n4428) );
  OAI21_X1 U5238 ( .B1(n4431), .B2(n6273), .A(n8696), .ZN(n4429) );
  NOR2_X1 U5239 ( .A1(n4728), .A2(n4432), .ZN(n4431) );
  INV_X1 U5240 ( .A(n8687), .ZN(n4432) );
  AND2_X1 U5241 ( .A1(n5971), .A2(n4442), .ZN(n6970) );
  OR2_X1 U5242 ( .A1(n4441), .A2(n7323), .ZN(n4442) );
  NAND2_X1 U5243 ( .A1(n7106), .A2(n6499), .ZN(n4441) );
  NAND3_X1 U5244 ( .A1(n7099), .A2(n8768), .A3(n7100), .ZN(n8767) );
  NAND2_X1 U5245 ( .A1(n9694), .A2(n8938), .ZN(n6522) );
  OR2_X1 U5246 ( .A1(n6480), .A2(n4436), .ZN(n7319) );
  INV_X1 U5247 ( .A(n6522), .ZN(n4436) );
  OAI21_X1 U5248 ( .B1(n4756), .B2(n4285), .A(n4434), .ZN(n6084) );
  INV_X1 U5249 ( .A(n4435), .ZN(n4434) );
  OAI21_X1 U5250 ( .B1(n4754), .B2(n4285), .A(n4913), .ZN(n4435) );
  NAND2_X1 U5251 ( .A1(n6427), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n6486) );
  NOR2_X1 U5252 ( .A1(n4774), .A2(n4301), .ZN(n4773) );
  NOR2_X1 U5253 ( .A1(n8678), .A2(n6420), .ZN(n4774) );
  AND2_X1 U5254 ( .A1(n6509), .A2(n6751), .ZN(n6521) );
  NAND2_X1 U5255 ( .A1(n4732), .A2(n8592), .ZN(n4731) );
  INV_X1 U5256 ( .A(n6238), .ZN(n4732) );
  INV_X1 U5257 ( .A(n8592), .ZN(n4735) );
  NAND3_X1 U5258 ( .A1(n4439), .A2(n6225), .A3(n4438), .ZN(n6239) );
  AND2_X1 U5259 ( .A1(n9174), .A2(n8936), .ZN(n9090) );
  AND2_X1 U5260 ( .A1(n6303), .A2(n6302), .ZN(n8640) );
  OR2_X1 U5261 ( .A1(n6991), .A2(n6990), .ZN(n6988) );
  NAND2_X1 U5262 ( .A1(n6808), .A2(n4304), .ZN(n6986) );
  INV_X1 U5263 ( .A(n6983), .ZN(n4591) );
  OR2_X1 U5264 ( .A1(n6786), .A2(n6787), .ZN(n6784) );
  NOR2_X1 U5265 ( .A1(n7001), .A2(n7000), .ZN(n4602) );
  OR2_X1 U5266 ( .A1(n6884), .A2(n6883), .ZN(n7008) );
  XNOR2_X1 U5267 ( .A(n9147), .B(n4421), .ZN(n9611) );
  NAND2_X1 U5268 ( .A1(n8826), .A2(n8825), .ZN(n9179) );
  INV_X1 U5269 ( .A(n4702), .ZN(n4701) );
  AOI21_X1 U5270 ( .B1(n4684), .B2(n8999), .A(n8912), .ZN(n4702) );
  NAND2_X1 U5271 ( .A1(n9482), .A2(n9287), .ZN(n4556) );
  NAND2_X1 U5272 ( .A1(n4554), .A2(n4894), .ZN(n4553) );
  AND2_X1 U5273 ( .A1(n9050), .A2(n9049), .ZN(n9256) );
  NAND2_X1 U5274 ( .A1(n7887), .A2(n9398), .ZN(n4472) );
  INV_X1 U5275 ( .A(n4900), .ZN(n4898) );
  OR2_X1 U5276 ( .A1(n9307), .A2(n7881), .ZN(n4899) );
  NAND2_X1 U5277 ( .A1(n4706), .A2(n8981), .ZN(n4705) );
  NAND2_X1 U5278 ( .A1(n4708), .A2(n9322), .ZN(n4706) );
  NAND2_X1 U5279 ( .A1(n9385), .A2(n4709), .ZN(n4704) );
  NAND2_X1 U5280 ( .A1(n9385), .A2(n9384), .ZN(n4713) );
  NAND2_X1 U5281 ( .A1(n6264), .A2(n6263), .ZN(n9382) );
  INV_X1 U5282 ( .A(n9077), .ZN(n9384) );
  NAND2_X1 U5283 ( .A1(n7772), .A2(n7771), .ZN(n7871) );
  INV_X1 U5284 ( .A(n9397), .ZN(n8846) );
  NAND2_X1 U5285 ( .A1(n7512), .A2(n7511), .ZN(n7665) );
  AND2_X1 U5286 ( .A1(n7510), .A2(n4889), .ZN(n4888) );
  AND2_X1 U5287 ( .A1(n8877), .A2(n8879), .ZN(n9069) );
  NAND2_X1 U5288 ( .A1(n9015), .A2(n4413), .ZN(n4412) );
  OAI21_X1 U5289 ( .B1(n9450), .B2(n9449), .A(n4321), .ZN(n9451) );
  NOR2_X1 U5290 ( .A1(n9448), .A2(n4610), .ZN(n4609) );
  NAND2_X1 U5291 ( .A1(n6209), .A2(n6208), .ZN(n9533) );
  AND2_X1 U5292 ( .A1(n6750), .A2(n6522), .ZN(n9736) );
  OR2_X1 U5293 ( .A1(n6479), .A2(n6504), .ZN(n9754) );
  NAND2_X1 U5294 ( .A1(n6566), .A2(n6274), .ZN(n5985) );
  INV_X1 U5295 ( .A(n9736), .ZN(n9768) );
  INV_X1 U5296 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n5919) );
  XNOR2_X1 U5297 ( .A(n5483), .B(n5482), .ZN(n7808) );
  XNOR2_X1 U5298 ( .A(n5450), .B(n5449), .ZN(n7632) );
  NAND2_X1 U5299 ( .A1(n5360), .A2(n5359), .ZN(n5377) );
  NAND2_X1 U5300 ( .A1(n5922), .A2(n6474), .ZN(n4775) );
  XNOR2_X1 U5301 ( .A(n5330), .B(n5329), .ZN(n7206) );
  AND2_X1 U5302 ( .A1(n6164), .A2(n5931), .ZN(n5935) );
  NAND2_X1 U5303 ( .A1(n4667), .A2(n4669), .ZN(n5297) );
  NAND2_X1 U5304 ( .A1(n4668), .A2(n5271), .ZN(n4667) );
  XNOR2_X1 U5305 ( .A(n5174), .B(n5173), .ZN(n6758) );
  XNOR2_X1 U5306 ( .A(n5008), .B(n5007), .ZN(n6608) );
  XNOR2_X1 U5307 ( .A(n5155), .B(n4909), .ZN(n6610) );
  AND2_X1 U5308 ( .A1(n6042), .A2(n6060), .ZN(n6658) );
  XNOR2_X1 U5309 ( .A(n4589), .B(P1_IR_REG_3__SCAN_IN), .ZN(n6665) );
  NAND2_X1 U5310 ( .A1(n6019), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4589) );
  NOR2_X1 U5311 ( .A1(n9589), .A2(n9588), .ZN(n9590) );
  NAND2_X1 U5312 ( .A1(n9593), .A2(n9594), .ZN(n9595) );
  NAND2_X1 U5313 ( .A1(n4508), .A2(n4515), .ZN(n4511) );
  NAND2_X1 U5314 ( .A1(n5405), .A2(n5404), .ZN(n8476) );
  INV_X2 U5315 ( .A(n7077), .ZN(n9821) );
  INV_X1 U5316 ( .A(n8050), .ZN(n8204) );
  NAND2_X2 U5317 ( .A1(n5092), .A2(n5091), .ZN(n7262) );
  NAND2_X1 U5318 ( .A1(n6574), .A2(n5474), .ZN(n5092) );
  NAND2_X1 U5319 ( .A1(n5383), .A2(n5382), .ZN(n8482) );
  NAND2_X1 U5320 ( .A1(n7961), .A2(n8423), .ZN(n8039) );
  OR2_X1 U5321 ( .A1(n5884), .A2(n5876), .ZN(n8019) );
  NAND2_X1 U5322 ( .A1(n7091), .A2(n5778), .ZN(n7151) );
  NAND2_X1 U5323 ( .A1(n5883), .A2(n5874), .ZN(n8029) );
  AND2_X1 U5324 ( .A1(n5729), .A2(n7343), .ZN(n4531) );
  NOR4_X1 U5325 ( .A1(n5591), .A2(n5592), .A3(n8185), .A4(n5584), .ZN(n5585)
         );
  NAND2_X1 U5326 ( .A1(n7343), .A2(n4352), .ZN(n4533) );
  INV_X1 U5327 ( .A(n7916), .ZN(n8322) );
  AOI22_X1 U5328 ( .A1(n7463), .A2(n7462), .B1(n7467), .B2(
        P2_REG1_REG_9__SCAN_IN), .ZN(n7539) );
  OAI21_X1 U5329 ( .B1(n4631), .B2(n5325), .A(n4626), .ZN(n4625) );
  NAND2_X1 U5330 ( .A1(n4632), .A2(n5325), .ZN(n4626) );
  OAI21_X1 U5331 ( .B1(n4631), .B2(P2_REG2_REG_19__SCAN_IN), .A(n4629), .ZN(
        n4628) );
  NAND2_X1 U5332 ( .A1(n4632), .A2(P2_REG2_REG_19__SCAN_IN), .ZN(n4629) );
  AOI22_X1 U5333 ( .A1(n4632), .A2(n8163), .B1(n8169), .B2(n8163), .ZN(n4630)
         );
  NOR2_X1 U5334 ( .A1(n8171), .A2(n4918), .ZN(n4404) );
  NAND2_X1 U5335 ( .A1(n7710), .A2(n5474), .ZN(n5456) );
  NAND2_X1 U5336 ( .A1(n8237), .A2(n8236), .ZN(n8460) );
  NAND2_X1 U5337 ( .A1(n8244), .A2(n7837), .ZN(n4792) );
  NAND2_X1 U5338 ( .A1(n5557), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5559) );
  NAND2_X1 U5339 ( .A1(n6086), .A2(n6085), .ZN(n7496) );
  NAND2_X1 U5340 ( .A1(n6228), .A2(n6227), .ZN(n9530) );
  INV_X1 U5341 ( .A(n9265), .ZN(n9482) );
  INV_X1 U5342 ( .A(n9099), .ZN(n4358) );
  NAND2_X1 U5343 ( .A1(n8940), .A2(n4360), .ZN(n4359) );
  INV_X1 U5344 ( .A(n9104), .ZN(n4354) );
  INV_X1 U5345 ( .A(n8640), .ZN(n9363) );
  OR2_X1 U5346 ( .A1(n6584), .A2(n5978), .ZN(n5983) );
  NAND2_X1 U5347 ( .A1(n7010), .A2(n7009), .ZN(n7239) );
  AOI21_X1 U5348 ( .B1(n9171), .B2(P1_ADDR_REG_19__SCAN_IN), .A(n9170), .ZN(
        n4605) );
  NAND2_X1 U5349 ( .A1(n4608), .A2(n9166), .ZN(n4361) );
  OR2_X1 U5350 ( .A1(n9168), .A2(n9167), .ZN(n4608) );
  NAND2_X1 U5351 ( .A1(n4419), .A2(n4418), .ZN(n4606) );
  OR2_X1 U5352 ( .A1(n9165), .A2(n9163), .ZN(n4418) );
  NAND2_X1 U5353 ( .A1(n9168), .A2(n9648), .ZN(n4419) );
  OAI21_X1 U5354 ( .B1(n4721), .B2(n9416), .A(n9191), .ZN(n9441) );
  XNOR2_X1 U5355 ( .A(n9186), .B(n9447), .ZN(n4721) );
  AOI21_X1 U5356 ( .B1(n7908), .B2(n9706), .A(n7907), .ZN(n9458) );
  NAND2_X1 U5357 ( .A1(n7906), .A2(n7905), .ZN(n7907) );
  NAND2_X1 U5358 ( .A1(n7891), .A2(n9450), .ZN(n9460) );
  NAND2_X1 U5359 ( .A1(n4892), .A2(n7877), .ZN(n9337) );
  NAND2_X1 U5360 ( .A1(n6295), .A2(n6294), .ZN(n9357) );
  NAND2_X1 U5361 ( .A1(n5941), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5943) );
  NOR2_X1 U5362 ( .A1(n9602), .A2(n10063), .ZN(n9902) );
  OAI21_X1 U5363 ( .B1(P1_ADDR_REG_17__SCAN_IN), .B2(P2_ADDR_REG_17__SCAN_IN), 
        .A(n9879), .ZN(n10059) );
  NAND2_X1 U5364 ( .A1(n5567), .A2(n6870), .ZN(n5608) );
  NAND2_X1 U5365 ( .A1(n4529), .A2(n4527), .ZN(n5626) );
  NAND2_X1 U5366 ( .A1(n5614), .A2(n5715), .ZN(n4527) );
  NAND2_X1 U5367 ( .A1(n7214), .A2(n5722), .ZN(n4529) );
  AND2_X1 U5368 ( .A1(n8876), .A2(n8877), .ZN(n4417) );
  OAI21_X1 U5369 ( .B1(n4535), .B2(n4534), .A(n5639), .ZN(n5645) );
  NAND2_X1 U5370 ( .A1(n5138), .A2(n5636), .ZN(n4534) );
  AOI21_X1 U5371 ( .B1(n5631), .B2(n5630), .A(n4536), .ZN(n4535) );
  OR2_X1 U5372 ( .A1(n8838), .A2(n8925), .ZN(n8908) );
  AND2_X1 U5373 ( .A1(n8864), .A2(n8879), .ZN(n8954) );
  OAI21_X1 U5374 ( .B1(n8907), .B2(n8943), .A(n4567), .ZN(n4566) );
  AND2_X1 U5375 ( .A1(n8903), .A2(n4568), .ZN(n4567) );
  NOR2_X1 U5376 ( .A1(n8908), .A2(n4415), .ZN(n4414) );
  NAND2_X1 U5377 ( .A1(n9053), .A2(n8981), .ZN(n4415) );
  NAND2_X1 U5378 ( .A1(n8997), .A2(n9050), .ZN(n4684) );
  OR3_X1 U5379 ( .A1(n9078), .A2(n9077), .A3(n9361), .ZN(n9079) );
  INV_X1 U5380 ( .A(n5717), .ZN(n4863) );
  NAND2_X1 U5381 ( .A1(n4861), .A2(n5717), .ZN(n4860) );
  INV_X1 U5382 ( .A(n8444), .ZN(n4861) );
  NAND2_X1 U5383 ( .A1(n8246), .A2(n5702), .ZN(n4537) );
  OAI21_X1 U5384 ( .B1(n5684), .B2(n5715), .A(n4539), .ZN(n4538) );
  INV_X1 U5385 ( .A(n5710), .ZN(n4583) );
  INV_X1 U5386 ( .A(n7872), .ZN(n4886) );
  OR2_X1 U5387 ( .A1(n9455), .A2(n9189), .ZN(n8941) );
  AND2_X1 U5388 ( .A1(n4679), .A2(n5395), .ZN(n4673) );
  INV_X1 U5389 ( .A(n5415), .ZN(n4677) );
  NAND2_X1 U5390 ( .A1(n4681), .A2(n5376), .ZN(n4680) );
  INV_X1 U5391 ( .A(n5396), .ZN(n4681) );
  AND2_X1 U5392 ( .A1(n5359), .A2(n5373), .ZN(n4679) );
  NAND2_X1 U5393 ( .A1(n5225), .A2(SI_14_), .ZN(n5267) );
  OAI21_X1 U5394 ( .B1(n4921), .B2(n4587), .A(n4586), .ZN(n4938) );
  OAI211_X1 U5395 ( .C1(n4919), .C2(n4544), .A(n4542), .B(n4541), .ZN(n4935)
         );
  NAND2_X1 U5396 ( .A1(n4543), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n4542) );
  INV_X1 U5397 ( .A(P1_RD_REG_SCAN_IN), .ZN(n4916) );
  INV_X1 U5398 ( .A(P2_RD_REG_SCAN_IN), .ZN(n4915) );
  NAND2_X1 U5399 ( .A1(n4306), .A2(n7929), .ZN(n4828) );
  NOR2_X1 U5400 ( .A1(n5321), .A2(n5320), .ZN(n4397) );
  XNOR2_X1 U5401 ( .A(n4823), .B(n5771), .ZN(n4824) );
  XNOR2_X1 U5402 ( .A(n5771), .B(n7027), .ZN(n5763) );
  NAND2_X1 U5403 ( .A1(n4857), .A2(n4864), .ZN(n4856) );
  NOR2_X1 U5404 ( .A1(n5719), .A2(n4346), .ZN(n4864) );
  NAND2_X1 U5405 ( .A1(n5002), .A2(n4523), .ZN(n5045) );
  AND2_X1 U5406 ( .A1(n4796), .A2(n4866), .ZN(n4791) );
  NAND2_X1 U5407 ( .A1(n8245), .A2(n4868), .ZN(n4867) );
  NAND2_X1 U5408 ( .A1(n4397), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n5364) );
  AND2_X1 U5409 ( .A1(n4658), .A2(n4659), .ZN(n4657) );
  INV_X1 U5410 ( .A(n8398), .ZN(n5266) );
  NAND2_X1 U5411 ( .A1(n4498), .A2(n4500), .ZN(n4495) );
  NAND2_X1 U5412 ( .A1(n5735), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5749) );
  OR2_X1 U5413 ( .A1(n5181), .A2(P2_IR_REG_12__SCAN_IN), .ZN(n5182) );
  OR2_X1 U5414 ( .A1(n5142), .A2(P2_IR_REG_9__SCAN_IN), .ZN(n5156) );
  OR2_X1 U5415 ( .A1(n5255), .A2(P2_IR_REG_8__SCAN_IN), .ZN(n5142) );
  NOR2_X1 U5416 ( .A1(n4730), .A2(n6273), .ZN(n4430) );
  NAND2_X1 U5417 ( .A1(n4761), .A2(n4760), .ZN(n4759) );
  INV_X1 U5418 ( .A(n6195), .ZN(n4760) );
  NOR2_X1 U5419 ( .A1(n7400), .A2(n4755), .ZN(n4754) );
  INV_X1 U5420 ( .A(n6028), .ZN(n4755) );
  NOR2_X1 U5421 ( .A1(n6401), .A2(n6402), .ZN(n8677) );
  AND2_X1 U5422 ( .A1(n9083), .A2(n4279), .ZN(n9086) );
  AND2_X1 U5423 ( .A1(n9179), .A2(n8828), .ZN(n9011) );
  NAND2_X1 U5424 ( .A1(n8930), .A2(n9198), .ZN(n8931) );
  INV_X1 U5425 ( .A(n6051), .ZN(n6069) );
  INV_X1 U5426 ( .A(n9091), .ZN(n9043) );
  INV_X1 U5427 ( .A(n9105), .ZN(n9002) );
  NAND2_X1 U5428 ( .A1(n9455), .A2(n9189), .ZN(n9184) );
  OAI21_X1 U5429 ( .B1(n4701), .B2(n4699), .A(n9048), .ZN(n4698) );
  INV_X1 U5430 ( .A(n9047), .ZN(n4699) );
  AND2_X1 U5431 ( .A1(n8843), .A2(n9047), .ZN(n4700) );
  NOR2_X1 U5432 ( .A1(n9466), .A2(n9472), .ZN(n4614) );
  OR2_X1 U5433 ( .A1(n8838), .A2(n4465), .ZN(n4461) );
  AND2_X1 U5434 ( .A1(n7899), .A2(n8839), .ZN(n4465) );
  OR2_X1 U5435 ( .A1(n9357), .A2(n8640), .ZN(n8905) );
  INV_X1 U5436 ( .A(n4718), .ZN(n4716) );
  INV_X1 U5437 ( .A(n8967), .ZN(n4715) );
  NOR2_X1 U5438 ( .A1(n4720), .A2(n4719), .ZN(n4718) );
  INV_X1 U5439 ( .A(n8889), .ZN(n4719) );
  NAND2_X1 U5440 ( .A1(n4454), .A2(n4453), .ZN(n4452) );
  INV_X1 U5441 ( .A(n4455), .ZN(n4453) );
  NOR2_X1 U5442 ( .A1(n8860), .A2(n4456), .ZN(n4455) );
  INV_X1 U5443 ( .A(n8871), .ZN(n4456) );
  NAND2_X1 U5444 ( .A1(n4455), .A2(n7516), .ZN(n4449) );
  NOR2_X1 U5445 ( .A1(n7620), .A2(n8720), .ZN(n4617) );
  OR2_X1 U5446 ( .A1(n7363), .A2(n7615), .ZN(n8870) );
  NAND2_X1 U5447 ( .A1(n4693), .A2(n7368), .ZN(n8961) );
  AND2_X1 U5448 ( .A1(n8988), .A2(n8987), .ZN(n7367) );
  NOR2_X1 U5449 ( .A1(n9445), .A2(n9768), .ZN(n4610) );
  NAND2_X1 U5450 ( .A1(n8941), .A2(n9184), .ZN(n9085) );
  NAND2_X1 U5451 ( .A1(n9369), .A2(n4286), .ZN(n9331) );
  NAND2_X1 U5452 ( .A1(n8632), .A2(n7533), .ZN(n7672) );
  INV_X1 U5453 ( .A(n4680), .ZN(n4675) );
  NAND2_X1 U5454 ( .A1(n4664), .A2(n4665), .ZN(n5308) );
  AOI21_X1 U5455 ( .B1(n4273), .B2(n4666), .A(n4326), .ZN(n4665) );
  NAND2_X1 U5456 ( .A1(n5223), .A2(n4273), .ZN(n4664) );
  AND2_X1 U5457 ( .A1(n5277), .A2(n4670), .ZN(n4669) );
  AOI21_X1 U5458 ( .B1(n5276), .B2(n5275), .A(n5274), .ZN(n5277) );
  NAND2_X1 U5459 ( .A1(n4399), .A2(n4559), .ZN(n4683) );
  AND2_X1 U5460 ( .A1(n4907), .A2(n4560), .ZN(n4559) );
  NAND2_X1 U5461 ( .A1(n4572), .A2(n4571), .ZN(n5110) );
  AOI21_X1 U5462 ( .B1(n4942), .B2(n4573), .A(n4316), .ZN(n4571) );
  INV_X1 U5463 ( .A(n5039), .ZN(n4661) );
  NAND2_X1 U5464 ( .A1(n4490), .A2(P2_ADDR_REG_19__SCAN_IN), .ZN(n4920) );
  NAND2_X1 U5465 ( .A1(n4915), .A2(P1_ADDR_REG_19__SCAN_IN), .ZN(n4490) );
  NAND2_X1 U5466 ( .A1(n7988), .A2(n4512), .ZN(n4508) );
  NAND2_X1 U5467 ( .A1(n4513), .A2(n7623), .ZN(n4512) );
  INV_X1 U5468 ( .A(n4397), .ZN(n5339) );
  NOR2_X1 U5469 ( .A1(n7192), .A2(n5781), .ZN(n4821) );
  INV_X1 U5470 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n5000) );
  INV_X1 U5471 ( .A(n4398), .ZN(n5422) );
  NAND2_X1 U5472 ( .A1(n5841), .A2(n5840), .ZN(n7966) );
  NAND2_X1 U5473 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n5082) );
  INV_X1 U5474 ( .A(n5132), .ZN(n4999) );
  NAND2_X1 U5475 ( .A1(n5185), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n5214) );
  INV_X1 U5476 ( .A(n5187), .ZN(n5185) );
  OR2_X1 U5477 ( .A1(n5015), .A2(n5000), .ZN(n5187) );
  INV_X1 U5478 ( .A(n4347), .ZN(n4513) );
  NAND2_X1 U5479 ( .A1(n5013), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n5015) );
  OR2_X1 U5480 ( .A1(n9801), .A2(n5885), .ZN(n7015) );
  NAND2_X1 U5481 ( .A1(n4996), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n5100) );
  INV_X1 U5482 ( .A(n5082), .ZN(n4996) );
  NAND2_X1 U5483 ( .A1(n4997), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5116) );
  INV_X1 U5484 ( .A(n5100), .ZN(n4997) );
  OAI21_X1 U5485 ( .B1(n4267), .B2(n5587), .A(n4852), .ZN(n4851) );
  NAND2_X1 U5486 ( .A1(n4267), .A2(n4853), .ZN(n4852) );
  NAND2_X1 U5487 ( .A1(n4854), .A2(n7207), .ZN(n4853) );
  INV_X1 U5488 ( .A(n4857), .ZN(n4854) );
  NAND2_X1 U5489 ( .A1(n4267), .A2(n7207), .ZN(n4855) );
  NAND2_X1 U5490 ( .A1(n5723), .A2(n5720), .ZN(n5592) );
  AND2_X1 U5491 ( .A1(n5721), .A2(n4377), .ZN(n5726) );
  NOR2_X1 U5492 ( .A1(n4379), .A2(n4378), .ZN(n4377) );
  NAND2_X1 U5493 ( .A1(n5719), .A2(n5720), .ZN(n4378) );
  AND3_X1 U5494 ( .A1(n5265), .A2(n5264), .A3(n5263), .ZN(n7825) );
  OR2_X1 U5495 ( .A1(n5051), .A2(n5050), .ZN(n5052) );
  OAI22_X1 U5496 ( .A1(n8585), .A2(n4526), .B1(n5002), .B2(n4525), .ZN(n4522)
         );
  AND2_X1 U5497 ( .A1(n4622), .A2(n4621), .ZN(n7542) );
  NAND2_X1 U5498 ( .A1(n7541), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n4621) );
  NAND2_X1 U5499 ( .A1(n4633), .A2(n4635), .ZN(n8075) );
  INV_X1 U5500 ( .A(n4636), .ZN(n4635) );
  OAI21_X1 U5501 ( .B1(n4638), .B2(n4640), .A(n8073), .ZN(n4636) );
  NAND2_X1 U5502 ( .A1(n8106), .A2(n8107), .ZN(n8110) );
  AOI21_X1 U5503 ( .B1(n8091), .B2(n8090), .A(n8089), .ZN(n8098) );
  NOR2_X1 U5504 ( .A1(n8110), .A2(n8109), .ZN(n8127) );
  AND2_X1 U5505 ( .A1(n8121), .A2(n8120), .ZN(n8122) );
  NOR2_X1 U5506 ( .A1(n8146), .A2(n8145), .ZN(n8153) );
  INV_X1 U5507 ( .A(n8169), .ZN(n4631) );
  AND2_X1 U5508 ( .A1(n7839), .A2(n7837), .ZN(n4796) );
  NAND2_X1 U5509 ( .A1(n4794), .A2(n4308), .ZN(n4793) );
  NAND2_X1 U5510 ( .A1(n7839), .A2(n4795), .ZN(n4794) );
  INV_X1 U5511 ( .A(n7838), .ZN(n4795) );
  NOR2_X1 U5512 ( .A1(n8455), .A2(n4650), .ZN(n4649) );
  INV_X1 U5513 ( .A(n4651), .ZN(n4650) );
  NAND2_X1 U5514 ( .A1(n4867), .A2(n4865), .ZN(n8222) );
  NAND2_X1 U5515 ( .A1(n8245), .A2(n5593), .ZN(n8234) );
  NAND2_X1 U5516 ( .A1(n8234), .A2(n8235), .ZN(n8233) );
  NAND2_X1 U5517 ( .A1(n5593), .A2(n5594), .ZN(n7837) );
  AOI21_X1 U5518 ( .B1(n4479), .B2(n4481), .A(n4477), .ZN(n4476) );
  INV_X1 U5519 ( .A(n5700), .ZN(n4477) );
  INV_X1 U5520 ( .A(n7837), .ZN(n8246) );
  NAND2_X1 U5521 ( .A1(n8286), .A2(n8469), .ZN(n8270) );
  NAND2_X1 U5522 ( .A1(n8302), .A2(n4849), .ZN(n8279) );
  NAND2_X1 U5523 ( .A1(n8320), .A2(n5394), .ZN(n8302) );
  INV_X1 U5524 ( .A(n8337), .ZN(n8307) );
  INV_X1 U5525 ( .A(n4871), .ZN(n4491) );
  AOI21_X1 U5526 ( .B1(n4324), .B2(n5347), .A(n4872), .ZN(n4871) );
  INV_X1 U5527 ( .A(n8319), .ZN(n5372) );
  NAND2_X1 U5528 ( .A1(n8376), .A2(n4657), .ZN(n8329) );
  NAND2_X1 U5529 ( .A1(n8349), .A2(n8350), .ZN(n8348) );
  NAND2_X1 U5530 ( .A1(n8376), .A2(n4659), .ZN(n8343) );
  NAND2_X1 U5531 ( .A1(n8376), .A2(n8362), .ZN(n8357) );
  NAND2_X1 U5532 ( .A1(n4395), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n5287) );
  INV_X1 U5533 ( .A(n5260), .ZN(n4395) );
  NAND2_X1 U5534 ( .A1(n5673), .A2(n8385), .ZN(n8398) );
  AND4_X1 U5535 ( .A1(n5192), .A2(n5191), .A3(n5190), .A4(n5189), .ZN(n7741)
         );
  AND3_X1 U5536 ( .A1(n5240), .A2(n5239), .A3(n5238), .ZN(n8403) );
  NAND2_X1 U5537 ( .A1(n7732), .A2(n7652), .ZN(n7744) );
  AND2_X1 U5538 ( .A1(n5658), .A2(n5659), .ZN(n7743) );
  INV_X1 U5539 ( .A(n5170), .ZN(n5171) );
  AND2_X1 U5540 ( .A1(n5170), .A2(n5654), .ZN(n7735) );
  NAND2_X1 U5541 ( .A1(n7693), .A2(n7694), .ZN(n7725) );
  AND4_X1 U5542 ( .A1(n5019), .A2(n5018), .A3(n5017), .A4(n5016), .ZN(n7627)
         );
  NAND2_X1 U5543 ( .A1(n7415), .A2(n5138), .ZN(n7433) );
  INV_X1 U5544 ( .A(n7560), .ZN(n5138) );
  OAI211_X1 U5545 ( .C1(n7137), .C2(n5614), .A(n7225), .B(n5107), .ZN(n5108)
         );
  INV_X1 U5546 ( .A(n8423), .ZN(n8402) );
  NOR2_X2 U5547 ( .A1(n7255), .A2(n7262), .ZN(n7258) );
  INV_X1 U5548 ( .A(n7021), .ZN(n7022) );
  OR2_X1 U5549 ( .A1(n5873), .A2(n7207), .ZN(n7111) );
  NOR2_X1 U5550 ( .A1(n7850), .A2(n4585), .ZN(n4521) );
  INV_X1 U5551 ( .A(n7846), .ZN(n4585) );
  NAND2_X1 U5552 ( .A1(n7843), .A2(n9786), .ZN(n4584) );
  AND2_X1 U5553 ( .A1(n4810), .A2(n4808), .ZN(n8481) );
  NAND2_X1 U5554 ( .A1(n5317), .A2(n5316), .ZN(n8498) );
  INV_X1 U5555 ( .A(n7262), .ZN(n9835) );
  INV_X1 U5556 ( .A(n8553), .ZN(n9854) );
  AND2_X1 U5557 ( .A1(n5860), .A2(n5859), .ZN(n9800) );
  NAND2_X1 U5558 ( .A1(n6539), .A2(n9806), .ZN(n9801) );
  INV_X1 U5559 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n4876) );
  NAND2_X1 U5560 ( .A1(n5314), .A2(n4911), .ZN(n5735) );
  NOR2_X1 U5561 ( .A1(n5730), .A2(n5733), .ZN(n5737) );
  XNOR2_X1 U5562 ( .A(n5536), .B(P2_IR_REG_21__SCAN_IN), .ZN(n5554) );
  NAND2_X1 U5563 ( .A1(n5535), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5536) );
  CLKBUF_X1 U5564 ( .A(n5251), .Z(n5252) );
  NAND2_X1 U5565 ( .A1(n6210), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n6230) );
  NAND2_X1 U5566 ( .A1(n6388), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n6412) );
  INV_X1 U5567 ( .A(n6389), .ZN(n6388) );
  NAND2_X1 U5568 ( .A1(n6377), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n6389) );
  NAND2_X1 U5569 ( .A1(n4424), .A2(n8676), .ZN(n4423) );
  NAND2_X1 U5570 ( .A1(n4756), .A2(n4754), .ZN(n7397) );
  INV_X1 U5571 ( .A(n6107), .ZN(n4763) );
  NAND2_X1 U5572 ( .A1(n7496), .A2(n7495), .ZN(n4765) );
  AND2_X1 U5573 ( .A1(n6330), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n6345) );
  INV_X1 U5574 ( .A(n6363), .ZN(n6364) );
  NAND2_X1 U5575 ( .A1(n4737), .A2(n4745), .ZN(n8745) );
  NOR2_X1 U5576 ( .A1(n4748), .A2(n4746), .ZN(n4745) );
  OR2_X1 U5577 ( .A1(n4271), .A2(n4747), .ZN(n4746) );
  AOI22_X1 U5578 ( .A1(n4750), .A2(n4743), .B1(n4283), .B2(n4742), .ZN(n4741)
         );
  NOR2_X1 U5579 ( .A1(n4744), .A2(n4271), .ZN(n4743) );
  INV_X1 U5580 ( .A(n4749), .ZN(n4744) );
  NAND2_X1 U5581 ( .A1(n6282), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n6297) );
  AND2_X1 U5582 ( .A1(n9042), .A2(n4349), .ZN(n4360) );
  AND4_X1 U5583 ( .A1(n6395), .A2(n6394), .A3(n6393), .A4(n6392), .ZN(n7900)
         );
  AND2_X1 U5584 ( .A1(n6353), .A2(n6352), .ZN(n7882) );
  INV_X1 U5585 ( .A(n6116), .ZN(n6524) );
  AND4_X1 U5586 ( .A1(n6122), .A2(n6121), .A3(n6120), .A4(n6119), .ZN(n8714)
         );
  NAND2_X1 U5587 ( .A1(n6988), .A2(n6653), .ZN(n9133) );
  OR2_X1 U5588 ( .A1(n6705), .A2(n6706), .ZN(n6861) );
  NAND2_X1 U5589 ( .A1(n6999), .A2(n4601), .ZN(n4600) );
  OAI21_X1 U5590 ( .B1(n7001), .B2(n4594), .A(n4592), .ZN(n7278) );
  NAND2_X1 U5591 ( .A1(n4595), .A2(n7229), .ZN(n4594) );
  INV_X1 U5592 ( .A(n4593), .ZN(n4592) );
  INV_X1 U5593 ( .A(n4596), .ZN(n4595) );
  AOI21_X1 U5594 ( .B1(n9148), .B2(n9614), .A(n9610), .ZN(n9623) );
  NAND2_X1 U5595 ( .A1(n9628), .A2(n4588), .ZN(n9159) );
  NAND2_X1 U5596 ( .A1(n9626), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n4588) );
  NOR2_X1 U5597 ( .A1(n9194), .A2(n9179), .ZN(n9178) );
  OR2_X1 U5598 ( .A1(n9198), .A2(n9002), .ZN(n9046) );
  NAND2_X1 U5599 ( .A1(n9228), .A2(n9396), .ZN(n7906) );
  NAND2_X1 U5600 ( .A1(n9012), .A2(n9005), .ZN(n9212) );
  INV_X1 U5601 ( .A(n4694), .ZN(n9213) );
  OAI21_X1 U5602 ( .B1(n9266), .B2(n4696), .A(n4695), .ZN(n4694) );
  NAND2_X1 U5603 ( .A1(n4700), .A2(n8950), .ZN(n4696) );
  INV_X1 U5604 ( .A(n4698), .ZN(n4695) );
  NOR2_X1 U5605 ( .A1(n9248), .A2(n4612), .ZN(n9220) );
  INV_X1 U5606 ( .A(n4614), .ZN(n4612) );
  NOR2_X1 U5607 ( .A1(n9248), .A2(n9472), .ZN(n9234) );
  NAND2_X1 U5608 ( .A1(n9031), .A2(n8999), .ZN(n9239) );
  NAND2_X1 U5609 ( .A1(n4462), .A2(n4461), .ZN(n9266) );
  OR2_X1 U5610 ( .A1(n9055), .A2(n9054), .ZN(n9308) );
  AND2_X1 U5611 ( .A1(n8905), .A2(n8953), .ZN(n9342) );
  AND2_X1 U5612 ( .A1(n9343), .A2(n7877), .ZN(n4891) );
  OR2_X1 U5613 ( .A1(n9360), .A2(n4270), .ZN(n4892) );
  AND2_X1 U5614 ( .A1(n4713), .A2(n4711), .ZN(n9341) );
  AND2_X1 U5615 ( .A1(n4575), .A2(n6244), .ZN(n7897) );
  NAND2_X1 U5616 ( .A1(n6964), .A2(n6274), .ZN(n4575) );
  NAND2_X1 U5617 ( .A1(n4551), .A2(n7873), .ZN(n9393) );
  INV_X1 U5618 ( .A(n7870), .ZN(n4550) );
  NAND2_X1 U5619 ( .A1(n7774), .A2(n8965), .ZN(n7777) );
  NAND2_X1 U5620 ( .A1(n7667), .A2(n4718), .ZN(n7774) );
  NOR2_X2 U5621 ( .A1(n6184), .A2(n6183), .ZN(n6185) );
  NAND2_X1 U5622 ( .A1(n4276), .A2(n4450), .ZN(n7667) );
  NAND2_X1 U5623 ( .A1(n4451), .A2(n4454), .ZN(n7517) );
  NAND2_X1 U5624 ( .A1(n7585), .A2(n4455), .ZN(n4451) );
  INV_X1 U5625 ( .A(n4616), .ZN(n7533) );
  NAND2_X1 U5626 ( .A1(n7591), .A2(n9769), .ZN(n7590) );
  NAND2_X1 U5627 ( .A1(n4457), .A2(n8871), .ZN(n7528) );
  OR2_X1 U5628 ( .A1(n7585), .A2(n7516), .ZN(n4457) );
  NAND2_X1 U5629 ( .A1(n7582), .A2(n7509), .ZN(n7527) );
  NOR2_X2 U5630 ( .A1(n6090), .A2(n6089), .ZN(n6117) );
  NAND2_X1 U5631 ( .A1(P1_REG3_REG_6__SCAN_IN), .A2(P1_REG3_REG_7__SCAN_IN), 
        .ZN(n6089) );
  NAND2_X1 U5632 ( .A1(n7359), .A2(n9063), .ZN(n7361) );
  AND2_X1 U5633 ( .A1(n8870), .A2(n8868), .ZN(n9066) );
  NOR2_X1 U5634 ( .A1(n7601), .A2(n7358), .ZN(n7388) );
  INV_X1 U5635 ( .A(n9063), .ZN(n7606) );
  NAND2_X1 U5636 ( .A1(n4384), .A2(n4383), .ZN(n7601) );
  INV_X1 U5637 ( .A(n9668), .ZN(n4384) );
  NAND2_X1 U5638 ( .A1(n9014), .A2(n8988), .ZN(n9060) );
  NAND2_X1 U5639 ( .A1(n8821), .A2(n8820), .ZN(n9433) );
  NAND2_X1 U5640 ( .A1(n4691), .A2(n6386), .ZN(n9477) );
  NAND2_X1 U5641 ( .A1(n7474), .A2(n8822), .ZN(n4691) );
  NAND2_X1 U5642 ( .A1(n6044), .A2(n6043), .ZN(n9735) );
  XNOR2_X1 U5643 ( .A(n5544), .B(n5525), .ZN(n8823) );
  XNOR2_X1 U5644 ( .A(n5520), .B(n5506), .ZN(n8816) );
  XNOR2_X1 U5645 ( .A(n5501), .B(n5500), .ZN(n8586) );
  AND2_X1 U5646 ( .A1(n5940), .A2(n5939), .ZN(n6464) );
  XNOR2_X1 U5647 ( .A(n5434), .B(n5429), .ZN(n7474) );
  XNOR2_X1 U5648 ( .A(n5335), .B(n5358), .ZN(n7245) );
  INV_X1 U5649 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n5921) );
  OR2_X1 U5650 ( .A1(n6144), .A2(P1_IR_REG_9__SCAN_IN), .ZN(n6179) );
  OR2_X1 U5651 ( .A1(n6108), .A2(P1_IR_REG_7__SCAN_IN), .ZN(n6110) );
  NAND2_X1 U5652 ( .A1(n4574), .A2(n4941), .ZN(n5094) );
  OR2_X1 U5653 ( .A1(n6041), .A2(P1_IR_REG_4__SCAN_IN), .ZN(n6060) );
  XNOR2_X1 U5654 ( .A(n5088), .B(n5089), .ZN(n6574) );
  NAND2_X1 U5655 ( .A1(n6037), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6001) );
  NAND2_X1 U5656 ( .A1(n6001), .A2(n6000), .ZN(n6019) );
  NOR2_X1 U5657 ( .A1(n9591), .A2(n10055), .ZN(n9592) );
  NAND2_X1 U5658 ( .A1(n9596), .A2(n9597), .ZN(n9598) );
  NAND2_X1 U5659 ( .A1(n9211), .A2(n7890), .ZN(n4884) );
  AND2_X1 U5660 ( .A1(n5392), .A2(n5391), .ZN(n7916) );
  AND4_X1 U5661 ( .A1(n5149), .A2(n5148), .A3(n5147), .A4(n5146), .ZN(n7556)
         );
  NAND2_X1 U5662 ( .A1(n7922), .A2(n7921), .ZN(n7920) );
  NAND2_X1 U5663 ( .A1(n4844), .A2(n4843), .ZN(n7922) );
  NAND2_X1 U5664 ( .A1(n7958), .A2(n4845), .ZN(n4844) );
  NOR2_X1 U5665 ( .A1(n5896), .A2(n5895), .ZN(n5897) );
  AND2_X1 U5666 ( .A1(n5491), .A2(n5510), .ZN(n8210) );
  AND4_X1 U5667 ( .A1(n5122), .A2(n5121), .A3(n5120), .A4(n5119), .ZN(n7416)
         );
  NOR2_X1 U5668 ( .A1(n5771), .A2(n7162), .ZN(n5761) );
  NAND2_X1 U5669 ( .A1(n5362), .A2(n5361), .ZN(n8487) );
  NAND2_X1 U5670 ( .A1(n4838), .A2(n4837), .ZN(n4833) );
  OR2_X1 U5671 ( .A1(n6542), .A2(n4832), .ZN(n4831) );
  NAND2_X1 U5672 ( .A1(n4836), .A2(n4278), .ZN(n4830) );
  NAND2_X1 U5673 ( .A1(n5440), .A2(n5439), .ZN(n8466) );
  AND2_X1 U5674 ( .A1(n4817), .A2(n4820), .ZN(n7947) );
  OR2_X1 U5675 ( .A1(n5760), .A2(n9791), .ZN(n7165) );
  INV_X1 U5676 ( .A(n4840), .ZN(n4839) );
  OAI21_X1 U5677 ( .B1(n4842), .B2(n4845), .A(n4841), .ZN(n4840) );
  OR2_X1 U5678 ( .A1(n7921), .A2(n5821), .ZN(n4841) );
  XNOR2_X1 U5679 ( .A(n5825), .B(n5823), .ZN(n7981) );
  NAND2_X1 U5680 ( .A1(n7928), .A2(n7929), .ZN(n8001) );
  AND4_X1 U5681 ( .A1(n5168), .A2(n5167), .A3(n5166), .A4(n5165), .ZN(n7435)
         );
  NAND2_X1 U5682 ( .A1(n4834), .A2(n4838), .ZN(n6543) );
  NAND2_X1 U5683 ( .A1(n7446), .A2(n4835), .ZN(n4834) );
  INV_X1 U5684 ( .A(n8024), .ZN(n7961) );
  NAND2_X1 U5685 ( .A1(n4846), .A2(n5815), .ZN(n8012) );
  OR2_X1 U5686 ( .A1(n7958), .A2(n7957), .ZN(n4846) );
  INV_X1 U5687 ( .A(n8019), .ZN(n8033) );
  NOR2_X1 U5688 ( .A1(n8020), .A2(n4517), .ZN(n4516) );
  INV_X1 U5689 ( .A(n4519), .ZN(n4517) );
  NAND2_X1 U5690 ( .A1(n4518), .A2(n4519), .ZN(n8018) );
  NAND2_X1 U5691 ( .A1(n5232), .A2(n5231), .ZN(n8517) );
  INV_X1 U5692 ( .A(n8029), .ZN(n8041) );
  INV_X1 U5693 ( .A(n8219), .ZN(n8049) );
  NAND2_X1 U5694 ( .A1(n5481), .A2(n5480), .ZN(n8050) );
  INV_X1 U5695 ( .A(n7932), .ZN(n8351) );
  OR2_X1 U5696 ( .A1(n6713), .A2(n6540), .ZN(n8052) );
  INV_X1 U5697 ( .A(n7177), .ZN(n8064) );
  AND3_X1 U5698 ( .A1(n5022), .A2(n5021), .A3(n5020), .ZN(n5024) );
  NAND2_X1 U5699 ( .A1(n5118), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n5023) );
  NOR2_X1 U5700 ( .A1(n6717), .A2(n4364), .ZN(n6731) );
  NAND2_X1 U5701 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), 
        .ZN(n4364) );
  NOR2_X1 U5702 ( .A1(n6801), .A2(n4910), .ZN(n6734) );
  NOR2_X1 U5703 ( .A1(n6734), .A2(n6733), .ZN(n6762) );
  NOR2_X1 U5704 ( .A1(n6827), .A2(n4289), .ZN(n6766) );
  NOR2_X1 U5705 ( .A1(n6766), .A2(n6765), .ZN(n6843) );
  INV_X1 U5706 ( .A(n4622), .ZN(n7540) );
  OAI22_X1 U5707 ( .A1(n7539), .A2(n7538), .B1(n7537), .B2(n7536), .ZN(n7757)
         );
  NAND2_X1 U5708 ( .A1(n4637), .A2(n4634), .ZN(n8074) );
  INV_X1 U5709 ( .A(n7792), .ZN(n4637) );
  AND2_X1 U5710 ( .A1(n5229), .A2(n5210), .ZN(n8084) );
  NOR2_X1 U5711 ( .A1(n8127), .A2(n4400), .ZN(n8131) );
  AND2_X1 U5712 ( .A1(n8128), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n4400) );
  NOR2_X1 U5713 ( .A1(n8131), .A2(n8130), .ZN(n8146) );
  NAND2_X1 U5714 ( .A1(n4392), .A2(n5545), .ZN(n4391) );
  AND2_X1 U5715 ( .A1(n5459), .A2(n5443), .ZN(n8253) );
  AND2_X1 U5716 ( .A1(n4805), .A2(n4807), .ZN(n8260) );
  NAND2_X1 U5717 ( .A1(n4475), .A2(n4479), .ZN(n8264) );
  NAND2_X1 U5718 ( .A1(n4810), .A2(n4811), .ZN(n8283) );
  NOR2_X1 U5719 ( .A1(n4781), .A2(n4780), .ZN(n8342) );
  OR2_X1 U5720 ( .A1(n4786), .A2(n7829), .ZN(n4780) );
  INV_X1 U5721 ( .A(n4785), .ZN(n4781) );
  AND2_X1 U5722 ( .A1(n8383), .A2(n5597), .ZN(n8364) );
  NAND2_X1 U5723 ( .A1(n8372), .A2(n7827), .ZN(n8356) );
  NAND2_X1 U5724 ( .A1(n5258), .A2(n5257), .ZN(n8512) );
  INV_X1 U5725 ( .A(n8517), .ZN(n8433) );
  AND2_X1 U5726 ( .A1(n4799), .A2(n7742), .ZN(n7746) );
  OR2_X1 U5727 ( .A1(n7687), .A2(n7565), .ZN(n8550) );
  NAND2_X1 U5728 ( .A1(n4494), .A2(n4500), .ZN(n7411) );
  NAND2_X1 U5729 ( .A1(n4778), .A2(n4497), .ZN(n4494) );
  INV_X1 U5730 ( .A(n4498), .ZN(n4497) );
  NAND2_X1 U5731 ( .A1(n4778), .A2(n7181), .ZN(n7226) );
  NAND2_X1 U5732 ( .A1(n7179), .A2(n7178), .ZN(n4779) );
  AOI22_X1 U5733 ( .A1(n5056), .A2(P1_DATAO_REG_3__SCAN_IN), .B1(n5315), .B2(
        n6767), .ZN(n5032) );
  INV_X1 U5734 ( .A(n7124), .ZN(n7027) );
  AND2_X1 U5735 ( .A1(n9798), .A2(n7026), .ZN(n8414) );
  AND2_X1 U5736 ( .A1(n9798), .A2(n9787), .ZN(n8284) );
  XNOR2_X1 U5737 ( .A(n4812), .B(n7021), .ZN(n9809) );
  OR2_X1 U5738 ( .A1(n9801), .A2(n7111), .ZN(n8411) );
  INV_X1 U5739 ( .A(n8284), .ZN(n8436) );
  INV_X1 U5740 ( .A(n9870), .ZN(n9871) );
  INV_X1 U5741 ( .A(n8452), .ZN(n4376) );
  OAI21_X1 U5742 ( .B1(n8463), .B2(n8544), .A(n4385), .ZN(n8562) );
  NOR2_X1 U5743 ( .A1(n8460), .A2(n4290), .ZN(n4385) );
  AND2_X1 U5744 ( .A1(n8462), .A2(n8553), .ZN(n4486) );
  AND2_X1 U5745 ( .A1(n4877), .A2(n4503), .ZN(n4502) );
  INV_X1 U5746 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n9904) );
  INV_X1 U5747 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n6938) );
  INV_X1 U5748 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n6850) );
  INV_X1 U5749 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n6612) );
  INV_X1 U5750 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n6611) );
  INV_X1 U5751 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n6605) );
  INV_X1 U5752 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n6603) );
  XNOR2_X1 U5753 ( .A(n5096), .B(P2_IR_REG_6__SCAN_IN), .ZN(n6908) );
  NAND2_X1 U5754 ( .A1(n6437), .A2(n6436), .ZN(n9462) );
  NOR2_X1 U5755 ( .A1(n6239), .A2(n6238), .ZN(n8591) );
  NAND2_X1 U5756 ( .A1(n4757), .A2(n4761), .ZN(n8623) );
  NAND2_X1 U5757 ( .A1(n7496), .A2(n4268), .ZN(n4757) );
  NAND2_X1 U5758 ( .A1(n8767), .A2(n6013), .ZN(n7200) );
  AOI21_X1 U5759 ( .B1(n6421), .B2(n4773), .A(n4767), .ZN(n4766) );
  NAND2_X1 U5760 ( .A1(n4292), .A2(n4768), .ZN(n4767) );
  NAND2_X1 U5761 ( .A1(n4773), .A2(n8678), .ZN(n4768) );
  NAND2_X1 U5762 ( .A1(n6450), .A2(n4770), .ZN(n4769) );
  NAND2_X1 U5763 ( .A1(n6450), .A2(n4772), .ZN(n4771) );
  INV_X1 U5764 ( .A(n4773), .ZN(n4770) );
  AND2_X1 U5765 ( .A1(n4752), .A2(n4751), .ZN(n8648) );
  NAND2_X1 U5766 ( .A1(n4740), .A2(n4749), .ZN(n4752) );
  NAND2_X1 U5767 ( .A1(n4433), .A2(n4431), .ZN(n8686) );
  NAND2_X1 U5768 ( .A1(n4726), .A2(n4725), .ZN(n4433) );
  OAI21_X1 U5769 ( .B1(n4726), .B2(n4427), .A(n4426), .ZN(n8695) );
  INV_X1 U5770 ( .A(n4431), .ZN(n4427) );
  AOI21_X1 U5771 ( .B1(n4431), .B2(n4730), .A(n6273), .ZN(n4426) );
  INV_X1 U5772 ( .A(n9477), .ZN(n9253) );
  NAND2_X1 U5773 ( .A1(n4756), .A2(n6028), .ZN(n7399) );
  AND2_X1 U5774 ( .A1(n4740), .A2(n4753), .ZN(n8725) );
  AND4_X1 U5775 ( .A1(n6173), .A2(n6172), .A3(n6171), .A4(n6170), .ZN(n8737)
         );
  NAND2_X1 U5776 ( .A1(n6361), .A2(n6360), .ZN(n9487) );
  AND4_X1 U5777 ( .A1(n6158), .A2(n6157), .A3(n6156), .A4(n6155), .ZN(n8760)
         );
  NAND2_X1 U5778 ( .A1(n6486), .A2(n6429), .ZN(n9222) );
  AND2_X1 U5779 ( .A1(n6521), .A2(n6481), .ZN(n8794) );
  INV_X1 U5780 ( .A(n8794), .ZN(n8814) );
  AND2_X1 U5781 ( .A1(n6512), .A2(n6511), .ZN(n8810) );
  OAI21_X1 U5782 ( .B1(n6239), .B2(n4733), .A(n4731), .ZN(n4736) );
  AND2_X1 U5783 ( .A1(n8656), .A2(n9736), .ZN(n8812) );
  INV_X1 U5784 ( .A(n7901), .ZN(n9241) );
  INV_X1 U5785 ( .A(n7900), .ZN(n9268) );
  OR2_X1 U5786 ( .A1(n6623), .A2(P1_U3084), .ZN(n9117) );
  OR2_X1 U5787 ( .A1(n6055), .A2(n6637), .ZN(n5952) );
  OR2_X1 U5788 ( .A1(n6584), .A2(n5947), .ZN(n5955) );
  XNOR2_X1 U5789 ( .A(n4362), .B(P1_REG2_REG_2__SCAN_IN), .ZN(n9127) );
  NAND2_X1 U5790 ( .A1(n6808), .A2(n6666), .ZN(n6984) );
  AND2_X1 U5791 ( .A1(n6986), .A2(n4332), .ZN(n9139) );
  INV_X1 U5792 ( .A(n6668), .ZN(n4590) );
  NAND2_X1 U5793 ( .A1(n6986), .A2(n6668), .ZN(n9137) );
  NAND2_X1 U5794 ( .A1(n6784), .A2(n6657), .ZN(n6700) );
  NOR2_X1 U5795 ( .A1(n4602), .A2(n4600), .ZN(n7233) );
  NAND2_X1 U5796 ( .A1(n4599), .A2(n6999), .ZN(n7002) );
  AND2_X1 U5797 ( .A1(n7008), .A2(n7007), .ZN(n7010) );
  NAND2_X1 U5798 ( .A1(n9630), .A2(n9629), .ZN(n9628) );
  INV_X1 U5799 ( .A(n9159), .ZN(n9641) );
  INV_X1 U5800 ( .A(n9163), .ZN(n9659) );
  NAND2_X1 U5801 ( .A1(n9195), .A2(n9194), .ZN(n9444) );
  AND2_X1 U5802 ( .A1(n9193), .A2(n9737), .ZN(n9195) );
  NAND2_X1 U5803 ( .A1(n4697), .A2(n4701), .ZN(n9226) );
  NAND2_X1 U5804 ( .A1(n4294), .A2(n8843), .ZN(n4697) );
  AOI21_X1 U5805 ( .B1(n9257), .B2(n9706), .A(n4470), .ZN(n9479) );
  NAND2_X1 U5806 ( .A1(n4472), .A2(n4471), .ZN(n4470) );
  NAND2_X1 U5807 ( .A1(n9287), .A2(n9396), .ZN(n4471) );
  AND2_X1 U5808 ( .A1(n6374), .A2(n6373), .ZN(n9265) );
  AOI21_X1 U5809 ( .B1(n9307), .B2(n4272), .A(n4894), .ZN(n9259) );
  INV_X1 U5810 ( .A(n9487), .ZN(n9280) );
  NAND2_X1 U5811 ( .A1(n4893), .A2(n4896), .ZN(n9273) );
  NAND2_X1 U5812 ( .A1(n9307), .A2(n4897), .ZN(n4893) );
  NAND2_X1 U5813 ( .A1(n4899), .A2(n4900), .ZN(n9299) );
  NAND2_X1 U5814 ( .A1(n4899), .A2(n4897), .ZN(n9297) );
  NAND2_X1 U5815 ( .A1(n4704), .A2(n4707), .ZN(n9323) );
  NAND2_X1 U5816 ( .A1(n6310), .A2(n6309), .ZN(n9503) );
  NAND2_X1 U5817 ( .A1(n6281), .A2(n6280), .ZN(n9514) );
  AND2_X1 U5818 ( .A1(n4713), .A2(n8952), .ZN(n9362) );
  NAND2_X1 U5819 ( .A1(n4887), .A2(n7872), .ZN(n9412) );
  NAND2_X1 U5820 ( .A1(n7871), .A2(n7870), .ZN(n4887) );
  NAND2_X1 U5821 ( .A1(n6167), .A2(n6166), .ZN(n8657) );
  OAI21_X1 U5822 ( .B1(n7665), .B2(n9069), .A(n7664), .ZN(n7666) );
  NAND2_X1 U5823 ( .A1(n6182), .A2(n6181), .ZN(n7716) );
  NAND2_X1 U5824 ( .A1(n6147), .A2(n6146), .ZN(n7513) );
  NAND2_X1 U5825 ( .A1(n4446), .A2(n6898), .ZN(n7365) );
  OR2_X1 U5826 ( .A1(n9754), .A2(n6505), .ZN(n9697) );
  INV_X1 U5827 ( .A(n9785), .ZN(n9783) );
  INV_X1 U5828 ( .A(n9441), .ZN(n9454) );
  AND2_X1 U5829 ( .A1(n9458), .A2(n9457), .ZN(n9459) );
  OR3_X1 U5830 ( .A1(n9512), .A2(n9511), .A3(n9510), .ZN(n9556) );
  INV_X1 U5831 ( .A(n9776), .ZN(n9774) );
  AND2_X1 U5832 ( .A1(n5931), .A2(n5946), .ZN(n4723) );
  AND2_X1 U5833 ( .A1(n4908), .A2(n5945), .ZN(n4722) );
  INV_X1 U5834 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n6606) );
  INV_X1 U5835 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n6601) );
  OAI21_X1 U5836 ( .B1(n9875), .B2(n9583), .A(n9877), .ZN(n10066) );
  AND2_X1 U5837 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n9590), .ZN(n10054) );
  XNOR2_X1 U5838 ( .A(n9592), .B(n4375), .ZN(n10053) );
  XNOR2_X1 U5839 ( .A(n9595), .B(n4373), .ZN(n10057) );
  INV_X1 U5840 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n4373) );
  XNOR2_X1 U5841 ( .A(n9598), .B(n4374), .ZN(n10062) );
  NOR2_X1 U5842 ( .A1(n9900), .A2(n4348), .ZN(n9899) );
  NOR2_X1 U5843 ( .A1(n9899), .A2(n9898), .ZN(n9897) );
  AND2_X1 U5844 ( .A1(n4369), .A2(n4368), .ZN(n9896) );
  NAND2_X1 U5845 ( .A1(P1_ADDR_REG_11__SCAN_IN), .A2(P2_ADDR_REG_11__SCAN_IN), 
        .ZN(n4368) );
  INV_X1 U5846 ( .A(n9897), .ZN(n4369) );
  NAND2_X1 U5847 ( .A1(n9896), .A2(n9895), .ZN(n9894) );
  OAI21_X1 U5848 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(P1_ADDR_REG_12__SCAN_IN), 
        .A(n9894), .ZN(n9892) );
  NAND2_X1 U5849 ( .A1(n9892), .A2(n9893), .ZN(n9891) );
  NAND2_X1 U5850 ( .A1(n9891), .A2(n4366), .ZN(n9889) );
  NAND2_X1 U5851 ( .A1(n9997), .A2(n4367), .ZN(n4366) );
  INV_X1 U5852 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n4367) );
  OAI21_X1 U5853 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(P1_ADDR_REG_14__SCAN_IN), 
        .A(n9888), .ZN(n9886) );
  NAND2_X1 U5854 ( .A1(n9886), .A2(n9887), .ZN(n9885) );
  NAND2_X1 U5855 ( .A1(n9885), .A2(n4370), .ZN(n9883) );
  NAND2_X1 U5856 ( .A1(n4372), .A2(n4371), .ZN(n4370) );
  INV_X1 U5857 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n4372) );
  NAND2_X1 U5858 ( .A1(n4883), .A2(n4884), .ZN(n4881) );
  NAND2_X1 U5859 ( .A1(n7150), .A2(n5782), .ZN(n7193) );
  OR2_X1 U5860 ( .A1(n4532), .A2(n4533), .ZN(n4393) );
  NAND2_X1 U5861 ( .A1(n4532), .A2(n4531), .ZN(n4530) );
  AND2_X1 U5862 ( .A1(n5754), .A2(n5753), .ZN(n4394) );
  NOR2_X1 U5863 ( .A1(n4404), .A2(n4403), .ZN(n4402) );
  OAI211_X1 U5864 ( .C1(n4627), .C2(n8156), .A(n4624), .B(n4630), .ZN(n4405)
         );
  INV_X1 U5865 ( .A(n8170), .ZN(n4403) );
  NAND2_X1 U5866 ( .A1(n4485), .A2(n4483), .ZN(P2_U3514) );
  OR2_X1 U5867 ( .A1(n9862), .A2(n4484), .ZN(n4483) );
  NAND2_X1 U5868 ( .A1(n8562), .A2(n9862), .ZN(n4485) );
  INV_X1 U5869 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n4484) );
  OR2_X1 U5870 ( .A1(n9103), .A2(n9102), .ZN(n4411) );
  AOI21_X1 U5871 ( .B1(n4606), .B2(n9694), .A(n4604), .ZN(n4603) );
  NAND2_X1 U5872 ( .A1(n4361), .A2(n9169), .ZN(n4607) );
  INV_X1 U5873 ( .A(n4605), .ZN(n4604) );
  OAI21_X1 U5874 ( .B1(n9479), .B2(n9716), .A(n4467), .ZN(P1_U3267) );
  INV_X1 U5875 ( .A(n4468), .ZN(n4467) );
  OAI21_X1 U5876 ( .B1(n9480), .B2(n9431), .A(n4469), .ZN(n4468) );
  AOI21_X1 U5877 ( .B1(n9476), .B2(n9407), .A(n9258), .ZN(n4469) );
  OAI21_X1 U5878 ( .B1(P1_ADDR_REG_18__SCAN_IN), .B2(n9606), .A(n10058), .ZN(
        n9608) );
  AND2_X1 U5879 ( .A1(n4856), .A2(n5724), .ZN(n4267) );
  OAI21_X1 U5880 ( .B1(n4896), .B2(n4895), .A(n4319), .ZN(n4894) );
  AND2_X1 U5881 ( .A1(n4275), .A2(n7495), .ZN(n4268) );
  INV_X4 U5882 ( .A(n5051), .ZN(n5118) );
  AND2_X1 U5883 ( .A1(n9514), .A2(n9386), .ZN(n4270) );
  AND2_X1 U5884 ( .A1(n6359), .A2(n6358), .ZN(n4271) );
  AND2_X1 U5885 ( .A1(n4897), .A2(n7884), .ZN(n4272) );
  XNOR2_X1 U5886 ( .A(n8455), .B(n8050), .ZN(n8223) );
  INV_X1 U5887 ( .A(n8223), .ZN(n4866) );
  OAI21_X1 U5888 ( .B1(n4731), .B2(n4729), .A(n4318), .ZN(n4728) );
  AND2_X1 U5889 ( .A1(n7716), .A2(n9108), .ZN(n4274) );
  NOR2_X1 U5890 ( .A1(n6142), .A2(n8621), .ZN(n4275) );
  AND2_X1 U5891 ( .A1(n4452), .A2(n9069), .ZN(n4276) );
  AND4_X1 U5892 ( .A1(n8899), .A2(n8898), .A3(n8952), .A4(n8897), .ZN(n4277)
         );
  INV_X1 U5893 ( .A(n9498), .ZN(n4902) );
  AND2_X1 U5894 ( .A1(n4838), .A2(n4837), .ZN(n4278) );
  NAND2_X1 U5895 ( .A1(n9031), .A2(n9050), .ZN(n4703) );
  XNOR2_X1 U5896 ( .A(n4935), .B(SI_3_), .ZN(n5029) );
  AND3_X1 U5897 ( .A1(n9204), .A2(n9084), .A3(n4386), .ZN(n4279) );
  AND2_X1 U5898 ( .A1(n4857), .A2(n5587), .ZN(n4280) );
  AND2_X1 U5899 ( .A1(n4433), .A2(n4727), .ZN(n4281) );
  INV_X1 U5900 ( .A(n9324), .ZN(n4901) );
  INV_X1 U5901 ( .A(n8678), .ZN(n4772) );
  INV_X1 U5902 ( .A(n5045), .ZN(n5262) );
  AND2_X1 U5903 ( .A1(n6098), .A2(n4878), .ZN(n6164) );
  NAND2_X1 U5904 ( .A1(n4751), .A2(n8646), .ZN(n4283) );
  OR2_X1 U5905 ( .A1(n7912), .A2(n5002), .ZN(n5051) );
  INV_X1 U5906 ( .A(n4730), .ZN(n4725) );
  NAND2_X1 U5907 ( .A1(n4734), .A2(n6258), .ZN(n4730) );
  AND2_X1 U5908 ( .A1(n8900), .A2(n4570), .ZN(n4284) );
  NAND2_X1 U5909 ( .A1(n7307), .A2(n6068), .ZN(n4285) );
  AND2_X1 U5910 ( .A1(n9329), .A2(n9509), .ZN(n4286) );
  NAND2_X1 U5911 ( .A1(n6101), .A2(n6100), .ZN(n7363) );
  AND2_X1 U5912 ( .A1(n6206), .A2(n8731), .ZN(n4287) );
  INV_X1 U5913 ( .A(n5223), .ZN(n4668) );
  INV_X1 U5914 ( .A(n7839), .ZN(n8235) );
  NAND2_X1 U5915 ( .A1(n9466), .A2(n9241), .ZN(n4288) );
  NAND2_X1 U5916 ( .A1(n5827), .A2(n5826), .ZN(n7928) );
  INV_X1 U5917 ( .A(n8197), .ZN(n8199) );
  NAND2_X1 U5918 ( .A1(n5711), .A2(n5499), .ZN(n8197) );
  INV_X1 U5919 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n5946) );
  AND2_X1 U5920 ( .A1(n6832), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n4289) );
  OR2_X1 U5921 ( .A1(n8461), .A2(n4486), .ZN(n4290) );
  OR2_X1 U5922 ( .A1(n5633), .A2(n5722), .ZN(n4291) );
  NAND2_X1 U5923 ( .A1(n4482), .A2(n5097), .ZN(n7219) );
  AND3_X1 U5924 ( .A1(n6006), .A2(n6005), .A3(n6004), .ZN(n6894) );
  AND2_X1 U5925 ( .A1(n6450), .A2(n6503), .ZN(n4292) );
  AND2_X1 U5926 ( .A1(n6239), .A2(n6238), .ZN(n4293) );
  INV_X1 U5927 ( .A(n8914), .ZN(n4690) );
  AND2_X1 U5928 ( .A1(n5347), .A2(n4873), .ZN(n4295) );
  AND2_X1 U5929 ( .A1(n4515), .A2(n7623), .ZN(n4296) );
  NAND2_X1 U5930 ( .A1(n5241), .A2(n5669), .ZN(n8397) );
  NAND2_X1 U5931 ( .A1(n4518), .A2(n4516), .ZN(n8021) );
  AND2_X1 U5932 ( .A1(n9322), .A2(n4709), .ZN(n4297) );
  NAND2_X1 U5933 ( .A1(n4892), .A2(n4891), .ZN(n9336) );
  NAND2_X1 U5934 ( .A1(n5700), .A2(n5701), .ZN(n8261) );
  INV_X1 U5935 ( .A(n8261), .ZN(n4804) );
  OR2_X1 U5936 ( .A1(n7716), .A2(n9108), .ZN(n4298) );
  AND2_X1 U5937 ( .A1(n4885), .A2(n4548), .ZN(n4299) );
  OR2_X1 U5938 ( .A1(n8063), .A2(n7262), .ZN(n4300) );
  NAND2_X1 U5939 ( .A1(n5476), .A2(n5475), .ZN(n8455) );
  OR2_X1 U5940 ( .A1(n8790), .A2(n8791), .ZN(n4301) );
  XNOR2_X1 U5941 ( .A(n5295), .B(SI_17_), .ZN(n5294) );
  NAND2_X1 U5942 ( .A1(n8286), .A2(n4651), .ZN(n4654) );
  AND2_X1 U5943 ( .A1(n9212), .A2(n4288), .ZN(n4302) );
  AND2_X1 U5944 ( .A1(n7821), .A2(n5220), .ZN(n7745) );
  INV_X1 U5945 ( .A(n7745), .ZN(n4798) );
  NAND2_X1 U5946 ( .A1(n7219), .A2(n8062), .ZN(n4303) );
  INV_X1 U5947 ( .A(n8274), .ZN(n8469) );
  NAND2_X1 U5948 ( .A1(n5420), .A2(n5419), .ZN(n8274) );
  AND2_X1 U5949 ( .A1(n4591), .A2(n6666), .ZN(n4304) );
  INV_X1 U5950 ( .A(n4611), .ZN(n9206) );
  NOR2_X1 U5951 ( .A1(n9248), .A2(n4613), .ZN(n4611) );
  AND2_X1 U5952 ( .A1(n8365), .A2(n5597), .ZN(n4305) );
  OR2_X1 U5953 ( .A1(n8003), .A2(n5829), .ZN(n4306) );
  AND2_X1 U5954 ( .A1(n4412), .A2(n8991), .ZN(n4307) );
  OR2_X1 U5955 ( .A1(n8462), .A2(n8051), .ZN(n4308) );
  INV_X1 U5956 ( .A(n8502), .ZN(n8362) );
  NAND2_X1 U5957 ( .A1(n5301), .A2(n5300), .ZN(n8502) );
  INV_X1 U5958 ( .A(n5554), .ZN(n7173) );
  OR2_X1 U5959 ( .A1(n8462), .A2(n8218), .ZN(n8216) );
  INV_X1 U5960 ( .A(n8216), .ZN(n4869) );
  INV_X1 U5961 ( .A(n4762), .ZN(n8616) );
  NAND2_X1 U5962 ( .A1(n4765), .A2(n4763), .ZN(n4762) );
  AND2_X1 U5963 ( .A1(n5266), .A2(n5669), .ZN(n4309) );
  OR2_X1 U5964 ( .A1(n8450), .A2(n8219), .ZN(n5711) );
  INV_X1 U5965 ( .A(n5711), .ZN(n4580) );
  OR2_X1 U5966 ( .A1(n5786), .A2(n5785), .ZN(n4310) );
  AND2_X1 U5967 ( .A1(n8228), .A2(n8204), .ZN(n4311) );
  NOR2_X1 U5968 ( .A1(n7883), .A2(n7882), .ZN(n4312) );
  INV_X1 U5969 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n6275) );
  NAND2_X1 U5970 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(P2_REG3_REG_10__SCAN_IN), 
        .ZN(n4313) );
  AND2_X1 U5971 ( .A1(n6732), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n4314) );
  AND2_X1 U5972 ( .A1(n9357), .A2(n9363), .ZN(n4315) );
  INV_X1 U5973 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n4990) );
  AND2_X1 U5974 ( .A1(n4943), .A2(SI_6_), .ZN(n4316) );
  OR2_X1 U5975 ( .A1(n4598), .A2(n7232), .ZN(n4317) );
  NAND2_X1 U5976 ( .A1(n6257), .A2(n6256), .ZN(n4318) );
  NAND2_X1 U5977 ( .A1(n9487), .A2(n9293), .ZN(n4319) );
  AND2_X1 U5978 ( .A1(n9466), .A2(n7901), .ZN(n9003) );
  INV_X1 U5979 ( .A(n4464), .ZN(n4463) );
  NAND2_X1 U5980 ( .A1(n4466), .A2(n9053), .ZN(n4464) );
  AND2_X1 U5981 ( .A1(n9530), .A2(n9397), .ZN(n4320) );
  AND2_X1 U5982 ( .A1(n9444), .A2(n4609), .ZN(n4321) );
  OR2_X1 U5983 ( .A1(n5685), .A2(n5722), .ZN(n4322) );
  OR2_X1 U5984 ( .A1(n8261), .A2(n8262), .ZN(n4323) );
  AND2_X1 U5985 ( .A1(n4873), .A2(n4875), .ZN(n4324) );
  NAND2_X1 U5986 ( .A1(n9265), .A2(n8833), .ZN(n4325) );
  AND2_X1 U5987 ( .A1(n5296), .A2(SI_17_), .ZN(n4326) );
  INV_X1 U5988 ( .A(n4708), .ZN(n4707) );
  OAI21_X1 U5989 ( .B1(n4711), .B2(n8851), .A(n8953), .ZN(n4708) );
  INV_X1 U5990 ( .A(n9031), .ZN(n8912) );
  OR2_X1 U5991 ( .A1(n9472), .A2(n8796), .ZN(n9031) );
  OR2_X1 U5992 ( .A1(n4764), .A2(n6107), .ZN(n4327) );
  AND2_X1 U5993 ( .A1(n5007), .A2(n4960), .ZN(n4328) );
  NAND2_X1 U5994 ( .A1(n4847), .A2(n8011), .ZN(n4329) );
  NAND2_X1 U5995 ( .A1(n5794), .A2(n5795), .ZN(n4838) );
  INV_X1 U5996 ( .A(n4734), .ZN(n4733) );
  NAND2_X1 U5997 ( .A1(n6238), .A2(n4735), .ZN(n4734) );
  INV_X1 U5998 ( .A(n8851), .ZN(n4710) );
  NAND2_X1 U5999 ( .A1(n7513), .A2(n8760), .ZN(n8879) );
  INV_X1 U6000 ( .A(n8879), .ZN(n4720) );
  INV_X1 U6001 ( .A(n4836), .ZN(n4835) );
  OR2_X1 U6002 ( .A1(n6553), .A2(n5792), .ZN(n4836) );
  INV_X1 U6003 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n6933) );
  XNOR2_X1 U6004 ( .A(n8476), .B(n8266), .ZN(n8282) );
  INV_X1 U6005 ( .A(n5806), .ZN(n4819) );
  AND3_X1 U6006 ( .A1(n5667), .A2(n5666), .A3(n8434), .ZN(n4330) );
  AND3_X1 U6007 ( .A1(n4710), .A2(n8886), .A3(n8885), .ZN(n4331) );
  INV_X1 U6008 ( .A(n5395), .ZN(n4678) );
  AND2_X1 U6009 ( .A1(n9265), .A2(n9287), .ZN(n9052) );
  NOR2_X1 U6010 ( .A1(n9136), .A2(n4590), .ZN(n4332) );
  INV_X1 U6011 ( .A(n8838), .ZN(n4466) );
  OAI21_X1 U6012 ( .B1(n8948), .B2(n9282), .A(n9056), .ZN(n8838) );
  AND2_X1 U6013 ( .A1(n9322), .A2(n9342), .ZN(n4333) );
  NOR2_X1 U6014 ( .A1(n8451), .A2(n4904), .ZN(n4334) );
  AND2_X1 U6015 ( .A1(n7178), .A2(n4300), .ZN(n4335) );
  INV_X1 U6016 ( .A(n4807), .ZN(n4806) );
  AOI21_X1 U6017 ( .B1(n4808), .B2(n8303), .A(n7835), .ZN(n4807) );
  XNOR2_X1 U6018 ( .A(n5374), .B(SI_21_), .ZN(n5373) );
  AND2_X1 U6019 ( .A1(n6767), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n4336) );
  AND2_X1 U6020 ( .A1(n8302), .A2(n5695), .ZN(n4337) );
  AND2_X1 U6021 ( .A1(n4684), .A2(n8999), .ZN(n8904) );
  INV_X1 U6022 ( .A(n8904), .ZN(n4409) );
  AND2_X1 U6023 ( .A1(n4804), .A2(n5699), .ZN(n4338) );
  AND2_X1 U6024 ( .A1(n4286), .A2(n4902), .ZN(n4339) );
  AND2_X1 U6025 ( .A1(n4902), .A2(n9324), .ZN(n9055) );
  AND2_X1 U6026 ( .A1(n8890), .A2(n7773), .ZN(n8965) );
  INV_X1 U6027 ( .A(n8965), .ZN(n4717) );
  OR2_X1 U6028 ( .A1(n7694), .A2(n7646), .ZN(n4340) );
  NAND2_X1 U6029 ( .A1(n8441), .A2(n5551), .ZN(n5724) );
  INV_X1 U6030 ( .A(n5125), .ZN(n4951) );
  NAND2_X1 U6031 ( .A1(n5139), .A2(n4950), .ZN(n5125) );
  INV_X1 U6032 ( .A(n8938), .ZN(n6504) );
  INV_X1 U6033 ( .A(n6371), .ZN(n4747) );
  OR2_X1 U6034 ( .A1(n7351), .A2(n9116), .ZN(n9014) );
  INV_X1 U6035 ( .A(n9014), .ZN(n4413) );
  NAND2_X1 U6036 ( .A1(n7446), .A2(n5793), .ZN(n6552) );
  NAND2_X1 U6037 ( .A1(n5337), .A2(n5336), .ZN(n8492) );
  INV_X1 U6038 ( .A(n8492), .ZN(n4658) );
  AND2_X1 U6039 ( .A1(n6342), .A2(n6341), .ZN(n4341) );
  NAND2_X1 U6040 ( .A1(n6899), .A2(n9043), .ZN(n6480) );
  NAND2_X1 U6041 ( .A1(n5730), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5560) );
  OR2_X1 U6042 ( .A1(n7583), .A2(n9068), .ZN(n7582) );
  NAND2_X1 U6043 ( .A1(n5456), .A2(n5455), .ZN(n8462) );
  INV_X1 U6044 ( .A(n8462), .ZN(n4652) );
  NAND2_X1 U6045 ( .A1(n7936), .A2(n7937), .ZN(n4342) );
  NAND3_X1 U6046 ( .A1(n4967), .A2(n5205), .A3(n5208), .ZN(n5253) );
  INV_X1 U6047 ( .A(n4271), .ZN(n4742) );
  NOR2_X1 U6048 ( .A1(n7792), .A2(n4642), .ZN(n4343) );
  INV_X1 U6049 ( .A(n4728), .ZN(n4727) );
  NAND2_X1 U6050 ( .A1(n4439), .A2(n4438), .ZN(n4344) );
  INV_X1 U6051 ( .A(n7937), .ZN(n4829) );
  AND2_X1 U6052 ( .A1(n7667), .A2(n8879), .ZN(n4345) );
  INV_X1 U6053 ( .A(n7742), .ZN(n4800) );
  INV_X1 U6054 ( .A(n6326), .ZN(n4753) );
  INV_X1 U6055 ( .A(n5975), .ZN(n6899) );
  INV_X1 U6056 ( .A(n9614), .ZN(n4421) );
  INV_X1 U6057 ( .A(n7429), .ZN(n4643) );
  INV_X1 U6058 ( .A(n8540), .ZN(n4406) );
  AND2_X1 U6059 ( .A1(n7099), .A2(n7100), .ZN(n7102) );
  AND2_X1 U6060 ( .A1(n5551), .A2(n5755), .ZN(n4346) );
  NAND2_X1 U6061 ( .A1(n4989), .A2(n4988), .ZN(n8535) );
  INV_X1 U6062 ( .A(n8535), .ZN(n4645) );
  NAND2_X1 U6063 ( .A1(n7794), .A2(n4639), .ZN(n4638) );
  INV_X1 U6064 ( .A(n4638), .ZN(n4634) );
  OR2_X1 U6065 ( .A1(n5799), .A2(n5798), .ZN(n4347) );
  NAND2_X1 U6066 ( .A1(n7073), .A2(n9821), .ZN(n7141) );
  AND2_X1 U6067 ( .A1(P1_ADDR_REG_10__SCAN_IN), .A2(P2_ADDR_REG_10__SCAN_IN), 
        .ZN(n4348) );
  AND2_X1 U6068 ( .A1(n8939), .A2(n4912), .ZN(n4349) );
  NAND3_X1 U6069 ( .A1(n5314), .A2(n4911), .A3(n4876), .ZN(n4350) );
  AND2_X1 U6070 ( .A1(n6722), .A2(n4391), .ZN(n4351) );
  INV_X1 U6071 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n4525) );
  INV_X1 U6072 ( .A(n9155), .ZN(n4420) );
  INV_X1 U6073 ( .A(n7000), .ZN(n4597) );
  INV_X1 U6074 ( .A(n7912), .ZN(n4523) );
  NAND2_X1 U6075 ( .A1(n6063), .A2(n6062), .ZN(n7602) );
  INV_X1 U6076 ( .A(n7602), .ZN(n4383) );
  AND2_X1 U6077 ( .A1(n7029), .A2(n7116), .ZN(n4352) );
  INV_X1 U6078 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n4503) );
  INV_X1 U6079 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n4526) );
  INV_X1 U6080 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n4375) );
  INV_X1 U6081 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n4692) );
  INV_X1 U6082 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n4587) );
  INV_X1 U6083 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n4371) );
  INV_X1 U6084 ( .A(n4362), .ZN(n9124) );
  NAND2_X1 U6085 ( .A1(n6002), .A2(n6019), .ZN(n4362) );
  INV_X1 U6086 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n4544) );
  INV_X1 U6087 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n4374) );
  NAND2_X1 U6088 ( .A1(n4353), .A2(n4411), .ZN(P1_U3240) );
  OAI21_X1 U6089 ( .B1(n9100), .B2(n4357), .A(n4354), .ZN(n4353) );
  NAND2_X1 U6090 ( .A1(n5469), .A2(n5468), .ZN(n5483) );
  NAND2_X1 U6091 ( .A1(n5418), .A2(n5417), .ZN(n5434) );
  NOR4_X2 U6092 ( .A1(n8940), .A2(n6899), .A3(n9090), .A4(n8937), .ZN(n9100)
         );
  NAND2_X1 U6093 ( .A1(n4683), .A2(n4328), .ZN(n5193) );
  NAND3_X1 U6094 ( .A1(n4356), .A2(n8927), .A3(n4355), .ZN(n8935) );
  NAND2_X1 U6095 ( .A1(n8926), .A2(n9445), .ZN(n4355) );
  INV_X1 U6096 ( .A(n8924), .ZN(n4356) );
  NAND2_X1 U6097 ( .A1(n4359), .A2(n4358), .ZN(n4357) );
  NAND2_X2 U6098 ( .A1(n8178), .A2(n7847), .ZN(n8192) );
  OAI22_X2 U6099 ( .A1(n7058), .A2(n7059), .B1(n5770), .B2(n5769), .ZN(n6956)
         );
  NAND2_X1 U6100 ( .A1(n7651), .A2(n7650), .ZN(n7732) );
  NAND2_X1 U6101 ( .A1(n4817), .A2(n4816), .ZN(n7946) );
  NAND2_X1 U6102 ( .A1(n7176), .A2(n7175), .ZN(n7179) );
  NAND2_X1 U6103 ( .A1(n7832), .A2(n4906), .ZN(n8328) );
  OAI21_X1 U6104 ( .B1(n7647), .B2(n4340), .A(n7649), .ZN(n7734) );
  AOI21_X1 U6105 ( .B1(n8392), .B2(n8422), .A(n7824), .ZN(n8396) );
  NAND3_X1 U6106 ( .A1(n5314), .A2(n4502), .A3(n4911), .ZN(n4504) );
  NAND2_X1 U6107 ( .A1(n5271), .A2(n4671), .ZN(n4670) );
  NAND2_X1 U6108 ( .A1(n4921), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n4586) );
  INV_X4 U6109 ( .A(n4563), .ZN(n4921) );
  NAND2_X1 U6110 ( .A1(n4489), .A2(n4488), .ZN(n4563) );
  AND2_X1 U6111 ( .A1(n8910), .A2(n8911), .ZN(n4408) );
  INV_X1 U6112 ( .A(n6377), .ZN(n6376) );
  NAND2_X1 U6113 ( .A1(n8295), .A2(n4808), .ZN(n4805) );
  INV_X1 U6114 ( .A(n7163), .ZN(n4823) );
  NAND2_X1 U6115 ( .A1(n7272), .A2(n7271), .ZN(n9144) );
  NAND2_X1 U6116 ( .A1(n8374), .A2(n4788), .ZN(n4785) );
  XNOR2_X1 U6117 ( .A(n9153), .B(P1_REG2_REG_19__SCAN_IN), .ZN(n9168) );
  NAND2_X1 U6118 ( .A1(n4363), .A2(n7851), .ZN(n7855) );
  NAND2_X1 U6120 ( .A1(n7822), .A2(n7821), .ZN(n8392) );
  NOR2_X1 U6121 ( .A1(n8396), .A2(n7826), .ZN(n8374) );
  NAND2_X1 U6122 ( .A1(n4499), .A2(n7413), .ZN(n7558) );
  BUF_X8 U6123 ( .A(n4921), .Z(n6575) );
  NAND2_X1 U6124 ( .A1(n5125), .A2(n4953), .ZN(n4560) );
  INV_X1 U6125 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n4917) );
  AND2_X2 U6126 ( .A1(n6364), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n6377) );
  NAND2_X1 U6127 ( .A1(n6410), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n6428) );
  OAI21_X1 U6128 ( .B1(n8915), .B2(n8913), .A(n4690), .ZN(n4689) );
  AOI21_X1 U6129 ( .B1(n7799), .B2(n7798), .A(n7797), .ZN(n8069) );
  NOR2_X1 U6130 ( .A1(n8102), .A2(n8103), .ZN(n8119) );
  NOR2_X1 U6131 ( .A1(n8139), .A2(n8138), .ZN(n8159) );
  OAI21_X1 U6132 ( .B1(n7053), .B2(n7051), .A(n7050), .ZN(n7286) );
  NAND2_X1 U6133 ( .A1(n8928), .A2(n8827), .ZN(n9089) );
  NAND2_X1 U6134 ( .A1(n5485), .A2(n5484), .ZN(n5501) );
  NAND2_X1 U6135 ( .A1(n5505), .A2(n5504), .ZN(n5520) );
  NAND2_X1 U6136 ( .A1(n9433), .A2(n9173), .ZN(n8928) );
  NAND2_X1 U6137 ( .A1(n5126), .A2(n4953), .ZN(n4399) );
  NAND2_X1 U6138 ( .A1(n5501), .A2(n5500), .ZN(n5505) );
  NAND2_X1 U6139 ( .A1(n8086), .A2(n8085), .ZN(n8106) );
  NAND2_X1 U6140 ( .A1(n5483), .A2(n5482), .ZN(n5485) );
  NAND2_X1 U6141 ( .A1(n4799), .A2(n4797), .ZN(n7822) );
  OAI211_X1 U6142 ( .C1(n4778), .C2(n4496), .A(n7410), .B(n4495), .ZN(n4499)
         );
  OAI21_X1 U6143 ( .B1(n8842), .B2(n8841), .A(n8904), .ZN(n8910) );
  NAND3_X1 U6144 ( .A1(n8453), .A2(n4376), .A3(n4334), .ZN(n8560) );
  INV_X1 U6145 ( .A(n7129), .ZN(n7079) );
  NAND2_X1 U6146 ( .A1(n8222), .A2(n5710), .ZN(n8200) );
  NAND2_X1 U6147 ( .A1(n7639), .A2(n7743), .ZN(n7638) );
  INV_X1 U6148 ( .A(n8065), .ZN(n7131) );
  NAND2_X1 U6149 ( .A1(n5024), .A2(n5023), .ZN(n8065) );
  NAND2_X1 U6150 ( .A1(n4478), .A2(n4476), .ZN(n8247) );
  NAND2_X1 U6151 ( .A1(n6773), .A2(n6772), .ZN(n6839) );
  INV_X1 U6152 ( .A(n4628), .ZN(n4627) );
  NAND2_X2 U6153 ( .A1(n7880), .A2(n7879), .ZN(n9307) );
  NAND2_X1 U6154 ( .A1(n7353), .A2(n7352), .ZN(n9665) );
  NAND2_X1 U6155 ( .A1(n7350), .A2(n7349), .ZN(n7477) );
  AND2_X2 U6156 ( .A1(n6640), .A2(n4392), .ZN(n6274) );
  NAND2_X1 U6157 ( .A1(n4380), .A2(n4330), .ZN(n5671) );
  NAND2_X1 U6158 ( .A1(n5653), .A2(n5652), .ZN(n4380) );
  AOI21_X1 U6159 ( .B1(n5688), .B2(n5687), .A(n5686), .ZN(n5693) );
  NAND2_X1 U6160 ( .A1(n5675), .A2(n5676), .ZN(n5688) );
  AOI21_X1 U6161 ( .B1(n4538), .B2(n4338), .A(n4537), .ZN(n5705) );
  NAND4_X1 U6162 ( .A1(n5696), .A2(n5695), .A3(n5694), .A4(n5715), .ZN(n4382)
         );
  NOR2_X2 U6163 ( .A1(n7484), .A2(n9729), .ZN(n9667) );
  NAND2_X1 U6164 ( .A1(n4776), .A2(n7564), .ZN(n7647) );
  NOR2_X1 U6165 ( .A1(n7466), .A2(n4623), .ZN(n7469) );
  NOR2_X1 U6166 ( .A1(n6762), .A2(n4336), .ZN(n6829) );
  AOI21_X1 U6167 ( .B1(P2_REG2_REG_7__SCAN_IN), .B2(n7043), .A(n7042), .ZN(
        n7045) );
  NAND2_X1 U6168 ( .A1(n4683), .A2(n4960), .ZN(n5008) );
  NOR2_X1 U6169 ( .A1(n7045), .A2(n7044), .ZN(n7291) );
  NOR2_X1 U6170 ( .A1(n6803), .A2(n6802), .ZN(n6801) );
  NOR2_X1 U6171 ( .A1(n6829), .A2(n6828), .ZN(n6827) );
  NOR2_X1 U6172 ( .A1(n6906), .A2(n6905), .ZN(n7042) );
  NOR2_X1 U6173 ( .A1(n7294), .A2(n7293), .ZN(n7466) );
  NAND2_X1 U6174 ( .A1(n5140), .A2(n5139), .ZN(n5152) );
  NAND2_X1 U6175 ( .A1(n5154), .A2(n5153), .ZN(n5155) );
  OR3_X2 U6176 ( .A1(n9090), .A2(n9089), .A3(n9088), .ZN(n9092) );
  INV_X2 U6177 ( .A(n9085), .ZN(n4386) );
  OAI21_X1 U6178 ( .B1(n8819), .B2(n4392), .A(n4351), .ZN(n8175) );
  NAND2_X1 U6179 ( .A1(n5518), .A2(SI_29_), .ZN(n5524) );
  NAND3_X1 U6180 ( .A1(n4394), .A2(n4530), .A3(n4393), .ZN(P2_U3244) );
  NAND2_X1 U6181 ( .A1(n5467), .A2(n5466), .ZN(n5469) );
  AOI21_X1 U6182 ( .B1(n8878), .B2(n4417), .A(n4720), .ZN(n8880) );
  NAND2_X1 U6183 ( .A1(n4998), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n5132) );
  NAND2_X1 U6184 ( .A1(n4792), .A2(n7838), .ZN(n8232) );
  INV_X1 U6185 ( .A(n4582), .ZN(n4581) );
  INV_X1 U6186 ( .A(n5126), .ZN(n4576) );
  NAND2_X1 U6187 ( .A1(n6933), .A2(n5025), .ZN(n5057) );
  NAND2_X1 U6188 ( .A1(n7542), .A2(n7543), .ZN(n7763) );
  XNOR2_X1 U6189 ( .A(n8104), .B(n8099), .ZN(n8086) );
  NAND2_X1 U6190 ( .A1(n7765), .A2(n4634), .ZN(n4633) );
  OAI21_X1 U6191 ( .B1(P2_IR_REG_31__SCAN_IN), .B2(P2_IR_REG_1__SCAN_IN), .A(
        n4620), .ZN(n4619) );
  XNOR2_X1 U6192 ( .A(n8153), .B(n8151), .ZN(n8147) );
  NAND2_X1 U6193 ( .A1(n8147), .A2(n5304), .ZN(n8154) );
  INV_X1 U6194 ( .A(n4619), .ZN(n4618) );
  NAND2_X1 U6195 ( .A1(n4405), .A2(n4402), .ZN(P2_U3264) );
  NOR2_X4 U6197 ( .A1(n4269), .A2(n8509), .ZN(n8376) );
  OAI21_X1 U6198 ( .B1(n8896), .B2(n8895), .A(n8969), .ZN(n8897) );
  OAI211_X2 U6199 ( .C1(n4410), .C2(n4409), .A(n4408), .B(n8909), .ZN(n8915)
         );
  NAND2_X2 U6200 ( .A1(n5353), .A2(n5352), .ZN(n5360) );
  NAND2_X1 U6201 ( .A1(n4672), .A2(n4676), .ZN(n5418) );
  NAND3_X1 U6202 ( .A1(n4722), .A2(n4723), .A3(n6164), .ZN(n9564) );
  OAI21_X1 U6203 ( .B1(n8915), .B2(n8912), .A(n4690), .ZN(n4687) );
  NOR2_X1 U6204 ( .A1(n4277), .A2(n4331), .ZN(n4570) );
  NAND2_X2 U6205 ( .A1(n9115), .A2(n9682), .ZN(n9015) );
  NAND2_X1 U6206 ( .A1(n4607), .A2(n4603), .ZN(P1_U3260) );
  XNOR2_X2 U6207 ( .A(n5984), .B(P1_IR_REG_1__SCAN_IN), .ZN(n6659) );
  NAND2_X1 U6208 ( .A1(n8703), .A2(n4422), .ZN(n8705) );
  NAND2_X1 U6209 ( .A1(n4423), .A2(n8704), .ZN(n8703) );
  NAND2_X1 U6210 ( .A1(n8675), .A2(n8674), .ZN(n4424) );
  NAND2_X1 U6211 ( .A1(n4726), .A2(n4430), .ZN(n4425) );
  NAND2_X1 U6212 ( .A1(n4425), .A2(n4428), .ZN(n8694) );
  INV_X1 U6213 ( .A(n6084), .ZN(n7335) );
  NAND3_X1 U6214 ( .A1(n4440), .A2(n6086), .A3(n4437), .ZN(n4438) );
  OR2_X2 U6215 ( .A1(n7323), .A2(n6045), .ZN(n6397) );
  NAND2_X1 U6216 ( .A1(n6969), .A2(n6970), .ZN(n6968) );
  AND3_X2 U6217 ( .A1(n5915), .A2(n5914), .A3(n5913), .ZN(n6098) );
  XNOR2_X2 U6218 ( .A(n4443), .B(P1_IR_REG_29__SCAN_IN), .ZN(n5951) );
  NAND4_X1 U6219 ( .A1(n6164), .A2(n4908), .A3(n5945), .A4(n5931), .ZN(n4444)
         );
  AND2_X1 U6220 ( .A1(n6898), .A2(n7366), .ZN(n4445) );
  NAND2_X1 U6221 ( .A1(n4447), .A2(n4714), .ZN(n7775) );
  NAND3_X1 U6222 ( .A1(n4276), .A2(n8965), .A3(n4450), .ZN(n4447) );
  INV_X1 U6223 ( .A(n4454), .ZN(n4448) );
  AOI21_X1 U6224 ( .B1(n9309), .B2(n9053), .A(n9055), .ZN(n9281) );
  NAND2_X1 U6225 ( .A1(n4473), .A2(n4936), .ZN(n5074) );
  NAND2_X1 U6226 ( .A1(n5030), .A2(n4934), .ZN(n4473) );
  NAND2_X1 U6227 ( .A1(n4474), .A2(n4933), .ZN(n5030) );
  NAND2_X1 U6228 ( .A1(n4932), .A2(n5059), .ZN(n4474) );
  NAND2_X1 U6229 ( .A1(n8320), .A2(n4479), .ZN(n4478) );
  NAND2_X1 U6230 ( .A1(n4917), .A2(n4916), .ZN(n4487) );
  NAND2_X1 U6231 ( .A1(n4487), .A2(n4918), .ZN(n4919) );
  NAND3_X1 U6232 ( .A1(n4918), .A2(n4917), .A3(n4916), .ZN(n4489) );
  AOI21_X2 U6233 ( .B1(n8363), .B2(n4295), .A(n4491), .ZN(n8321) );
  NAND2_X2 U6234 ( .A1(n8383), .A2(n4305), .ZN(n8363) );
  NAND2_X2 U6235 ( .A1(n4493), .A2(n7020), .ZN(n5771) );
  INV_X2 U6236 ( .A(n8062), .ZN(n4501) );
  NAND3_X1 U6237 ( .A1(n5314), .A2(n4911), .A3(n4877), .ZN(n4993) );
  AND4_X4 U6238 ( .A1(n4975), .A2(n4983), .A3(n5251), .A4(n5279), .ZN(n5314)
         );
  NAND3_X1 U6239 ( .A1(n4508), .A2(n4515), .A3(n7811), .ZN(n4506) );
  NAND2_X1 U6240 ( .A1(n4511), .A2(n4509), .ZN(n7810) );
  NAND2_X1 U6241 ( .A1(n7625), .A2(n4296), .ZN(n4509) );
  INV_X1 U6242 ( .A(n4510), .ZN(n7809) );
  OAI21_X1 U6243 ( .B1(n7625), .B2(n4513), .A(n7623), .ZN(n7989) );
  NAND2_X1 U6244 ( .A1(n5800), .A2(n5801), .ZN(n4515) );
  NAND2_X1 U6245 ( .A1(n5846), .A2(n5845), .ZN(n7939) );
  NAND2_X1 U6246 ( .A1(n4522), .A2(n4523), .ZN(n4524) );
  NAND3_X1 U6247 ( .A1(n5047), .A2(n5046), .A3(n4524), .ZN(n5760) );
  OAI21_X2 U6248 ( .B1(n7958), .B2(n4842), .A(n4839), .ZN(n7980) );
  NAND2_X2 U6249 ( .A1(n7946), .A2(n5811), .ZN(n7958) );
  NAND2_X1 U6250 ( .A1(n9835), .A2(n8063), .ZN(n5625) );
  INV_X1 U6251 ( .A(n4920), .ZN(n4543) );
  NAND3_X1 U6252 ( .A1(n4919), .A2(n4920), .A3(P2_DATAO_REG_3__SCAN_IN), .ZN(
        n4541) );
  INV_X1 U6253 ( .A(n7665), .ZN(n4545) );
  AOI21_X1 U6254 ( .B1(n4547), .B2(n4545), .A(n4546), .ZN(n7707) );
  OAI21_X1 U6255 ( .B1(n7772), .B2(n4550), .A(n4299), .ZN(n4551) );
  NAND2_X1 U6256 ( .A1(n4554), .A2(n9307), .ZN(n4552) );
  INV_X1 U6257 ( .A(n7886), .ZN(n9246) );
  NAND2_X1 U6258 ( .A1(n9360), .A2(n4891), .ZN(n4557) );
  NAND2_X1 U6259 ( .A1(n4557), .A2(n4558), .ZN(n9321) );
  NAND2_X1 U6260 ( .A1(n4576), .A2(n4951), .ZN(n5140) );
  NAND2_X1 U6261 ( .A1(n4563), .A2(n4925), .ZN(n4930) );
  OAI211_X1 U6262 ( .C1(n4921), .C2(n6598), .A(n4931), .B(n4561), .ZN(n4932)
         );
  NAND2_X1 U6263 ( .A1(n4921), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n4561) );
  OAI211_X1 U6264 ( .C1(n4921), .C2(P2_DATAO_REG_2__SCAN_IN), .A(SI_2_), .B(
        n4562), .ZN(n4933) );
  NAND2_X1 U6265 ( .A1(n4921), .A2(n6561), .ZN(n4562) );
  MUX2_X1 U6266 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(P1_DATAO_REG_5__SCAN_IN), 
        .S(n4921), .Z(n4940) );
  MUX2_X1 U6267 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(P1_DATAO_REG_1__SCAN_IN), 
        .S(n4921), .Z(n5041) );
  MUX2_X1 U6268 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(P1_DATAO_REG_6__SCAN_IN), 
        .S(n4921), .Z(n4943) );
  MUX2_X1 U6269 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(P1_DATAO_REG_2__SCAN_IN), 
        .S(n4921), .Z(n5060) );
  MUX2_X1 U6270 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(P1_DATAO_REG_7__SCAN_IN), 
        .S(n6575), .Z(n4945) );
  MUX2_X1 U6271 ( .A(n6601), .B(n6603), .S(n4921), .Z(n4948) );
  MUX2_X1 U6272 ( .A(n5244), .B(n5245), .S(n4921), .Z(n5247) );
  MUX2_X1 U6273 ( .A(n6852), .B(n6796), .S(n4921), .Z(n5224) );
  MUX2_X1 U6274 ( .A(n6614), .B(n6611), .S(n6575), .Z(n4955) );
  MUX2_X1 U6275 ( .A(n6965), .B(n6967), .S(n6575), .Z(n5227) );
  MUX2_X1 U6276 ( .A(n4961), .B(n6612), .S(n6575), .Z(n4962) );
  MUX2_X1 U6277 ( .A(n6606), .B(n6605), .S(n6575), .Z(n4958) );
  MUX2_X1 U6278 ( .A(n5175), .B(n6850), .S(n6575), .Z(n5177) );
  MUX2_X1 U6279 ( .A(n6759), .B(n6761), .S(n6575), .Z(n4965) );
  MUX2_X1 U6280 ( .A(n5278), .B(n6938), .S(n6575), .Z(n5295) );
  MUX2_X1 U6281 ( .A(n7268), .B(n7246), .S(n6575), .Z(n5332) );
  MUX2_X1 U6282 ( .A(n7209), .B(n7208), .S(n6575), .Z(n5311) );
  MUX2_X1 U6283 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(P1_DATAO_REG_18__SCAN_IN), 
        .S(n6575), .Z(n5309) );
  MUX2_X1 U6284 ( .A(n7211), .B(n9904), .S(n6575), .Z(n5374) );
  MUX2_X1 U6285 ( .A(n7407), .B(n7409), .S(n6575), .Z(n5379) );
  MUX2_X1 U6286 ( .A(n5398), .B(n5399), .S(n6575), .Z(n5401) );
  MUX2_X1 U6287 ( .A(n7475), .B(n7494), .S(n6575), .Z(n5430) );
  MUX2_X1 U6288 ( .A(n7633), .B(n7637), .S(n6575), .Z(n5436) );
  MUX2_X1 U6289 ( .A(n7712), .B(n10015), .S(n6575), .Z(n5452) );
  MUX2_X1 U6290 ( .A(n10017), .B(n7820), .S(n6575), .Z(n5471) );
  MUX2_X1 U6291 ( .A(n9990), .B(n8588), .S(n6575), .Z(n5503) );
  MUX2_X1 U6292 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(P1_DATAO_REG_29__SCAN_IN), 
        .S(n6575), .Z(n5521) );
  NAND2_X1 U6293 ( .A1(n5088), .A2(n4577), .ZN(n4574) );
  NAND3_X1 U6294 ( .A1(n5088), .A2(n4577), .A3(n4942), .ZN(n4572) );
  INV_X1 U6295 ( .A(n5089), .ZN(n4577) );
  NAND2_X1 U6296 ( .A1(n4867), .A2(n4581), .ZN(n4578) );
  NAND2_X1 U6297 ( .A1(n4578), .A2(n4579), .ZN(n7842) );
  NAND2_X2 U6298 ( .A1(n8401), .A2(n5293), .ZN(n8383) );
  NAND2_X1 U6299 ( .A1(n4584), .A2(n7846), .ZN(n8194) );
  INV_X1 U6300 ( .A(n4602), .ZN(n4599) );
  INV_X1 U6301 ( .A(n7003), .ZN(n4601) );
  NAND2_X1 U6302 ( .A1(n7278), .A2(n7277), .ZN(n7279) );
  NOR2_X2 U6303 ( .A1(n9406), .A2(n9382), .ZN(n9377) );
  NAND2_X1 U6304 ( .A1(n9404), .A2(n7897), .ZN(n9406) );
  NOR2_X2 U6305 ( .A1(n9419), .A2(n9530), .ZN(n9404) );
  NAND2_X1 U6306 ( .A1(n7782), .A2(n8743), .ZN(n9419) );
  NOR3_X4 U6307 ( .A1(n9248), .A2(n9455), .A3(n4613), .ZN(n9192) );
  NAND2_X1 U6308 ( .A1(n9369), .A2(n4339), .ZN(n9315) );
  NAND2_X1 U6309 ( .A1(n4617), .A2(n7591), .ZN(n4616) );
  NAND2_X1 U6310 ( .A1(n4615), .A2(n8632), .ZN(n7702) );
  MUX2_X1 U6311 ( .A(P2_REG2_REG_1__SCAN_IN), .B(n6711), .S(n6737), .Z(n6717)
         );
  NAND3_X1 U6312 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .A3(
        P2_IR_REG_0__SCAN_IN), .ZN(n4620) );
  NAND2_X1 U6313 ( .A1(n8156), .A2(n4625), .ZN(n4624) );
  INV_X1 U6314 ( .A(n7765), .ZN(n4641) );
  AND2_X2 U6316 ( .A1(n7748), .A2(n8522), .ZN(n8428) );
  NOR2_X2 U6317 ( .A1(n7747), .A2(n8529), .ZN(n7748) );
  AND3_X2 U6318 ( .A1(n4647), .A2(n9791), .A3(n7124), .ZN(n7073) );
  OR2_X1 U6319 ( .A1(n7163), .A2(n7162), .ZN(n4648) );
  INV_X1 U6320 ( .A(n4648), .ZN(n7161) );
  INV_X1 U6321 ( .A(n4654), .ZN(n8238) );
  AND2_X2 U6322 ( .A1(n8376), .A2(n4655), .ZN(n8315) );
  NAND2_X1 U6323 ( .A1(n4660), .A2(n5958), .ZN(n5040) );
  NAND2_X1 U6324 ( .A1(n4921), .A2(n4661), .ZN(n4660) );
  NAND3_X1 U6325 ( .A1(n4919), .A2(n4920), .A3(n5038), .ZN(n5958) );
  XNOR2_X2 U6326 ( .A(n5028), .B(P2_IR_REG_3__SCAN_IN), .ZN(n6767) );
  AOI21_X1 U6327 ( .B1(P2_REG2_REG_5__SCAN_IN), .B2(n6844), .A(n6843), .ZN(
        n6846) );
  AOI21_X1 U6328 ( .B1(P2_REG2_REG_6__SCAN_IN), .B2(n6908), .A(n6904), .ZN(
        n6906) );
  NAND2_X1 U6329 ( .A1(n8075), .A2(n8076), .ZN(n8083) );
  NOR2_X1 U6330 ( .A1(n6846), .A2(n6845), .ZN(n6904) );
  AND2_X2 U6331 ( .A1(n6640), .A2(n6575), .ZN(n6003) );
  NAND2_X1 U6332 ( .A1(n5110), .A2(n4944), .ZN(n4662) );
  NAND2_X1 U6333 ( .A1(n5074), .A2(n4937), .ZN(n4663) );
  NAND2_X1 U6334 ( .A1(n5360), .A2(n4679), .ZN(n4682) );
  NAND2_X1 U6335 ( .A1(n5360), .A2(n4673), .ZN(n4672) );
  NAND4_X1 U6336 ( .A1(n4688), .A2(n4686), .A3(n9204), .A4(n4685), .ZN(n8917)
         );
  NAND3_X1 U6337 ( .A1(n4687), .A2(n9466), .A3(n8927), .ZN(n4686) );
  NAND3_X1 U6338 ( .A1(n4689), .A2(n8925), .A3(n9241), .ZN(n4688) );
  NAND2_X1 U6339 ( .A1(n4693), .A2(n8987), .ZN(n7479) );
  AOI21_X2 U6340 ( .B1(n9385), .B2(n4297), .A(n4705), .ZN(n9309) );
  AOI21_X1 U6341 ( .B1(n8965), .B2(n4716), .A(n4715), .ZN(n4714) );
  NAND2_X2 U6342 ( .A1(n9101), .A2(n4724), .ZN(n9710) );
  OR2_X2 U6343 ( .A1(n9091), .A2(n6504), .ZN(n7478) );
  INV_X1 U6344 ( .A(n6239), .ZN(n4726) );
  INV_X1 U6345 ( .A(n4736), .ZN(n8805) );
  NAND2_X1 U6346 ( .A1(n8635), .A2(n6327), .ZN(n4750) );
  NAND2_X1 U6347 ( .A1(n8635), .A2(n4738), .ZN(n4737) );
  CLKBUF_X1 U6348 ( .A(n4750), .Z(n4740) );
  OAI21_X1 U6349 ( .B1(n6421), .B2(n8678), .A(n4773), .ZN(n8793) );
  INV_X1 U6350 ( .A(n4766), .ZN(n6537) );
  OAI21_X1 U6351 ( .B1(n6421), .B2(n4771), .A(n4769), .ZN(n7863) );
  AOI21_X1 U6352 ( .B1(n6421), .B2(n6420), .A(n8678), .ZN(n8792) );
  NAND2_X1 U6353 ( .A1(n7558), .A2(n4777), .ZN(n4776) );
  AND2_X1 U6354 ( .A1(n7563), .A2(n7557), .ZN(n4777) );
  NAND2_X1 U6355 ( .A1(n7179), .A2(n4335), .ZN(n4778) );
  XNOR2_X1 U6356 ( .A(n4779), .B(n7250), .ZN(n9833) );
  NAND2_X1 U6357 ( .A1(n4785), .A2(n4782), .ZN(n7832) );
  NAND2_X1 U6358 ( .A1(n7732), .A2(n4801), .ZN(n4799) );
  NAND2_X1 U6359 ( .A1(n5567), .A2(n5609), .ZN(n4813) );
  NAND2_X1 U6360 ( .A1(n4813), .A2(n7022), .ZN(n7024) );
  CLKBUF_X1 U6361 ( .A(n4813), .Z(n4812) );
  NOR2_X1 U6362 ( .A1(n7066), .A2(n4812), .ZN(n5570) );
  XNOR2_X1 U6363 ( .A(n4812), .B(n7165), .ZN(n7167) );
  NAND2_X1 U6364 ( .A1(n5756), .A2(n6942), .ZN(n4815) );
  NAND3_X1 U6365 ( .A1(n6923), .A2(n6942), .A3(n6925), .ZN(n4814) );
  AOI21_X2 U6366 ( .B1(n6956), .B2(n6952), .A(n6954), .ZN(n7092) );
  NAND2_X1 U6367 ( .A1(n5807), .A2(n4819), .ZN(n4817) );
  NAND2_X1 U6368 ( .A1(n7809), .A2(n5805), .ZN(n8032) );
  NAND2_X1 U6369 ( .A1(n7150), .A2(n4821), .ZN(n4822) );
  NAND2_X1 U6370 ( .A1(n7151), .A2(n7152), .ZN(n7150) );
  INV_X1 U6371 ( .A(n4824), .ZN(n5758) );
  NAND2_X1 U6372 ( .A1(n5757), .A2(n4824), .ZN(n6944) );
  NAND2_X1 U6374 ( .A1(n5817), .A2(n5818), .ZN(n4848) );
  NAND3_X1 U6375 ( .A1(n6870), .A2(n5567), .A3(n5755), .ZN(n5604) );
  NAND2_X1 U6376 ( .A1(n5049), .A2(n5567), .ZN(n5603) );
  NAND2_X2 U6377 ( .A1(n5241), .A2(n4309), .ZN(n8401) );
  NAND2_X1 U6378 ( .A1(n5517), .A2(n4280), .ZN(n4850) );
  OAI211_X1 U6379 ( .C1(n5517), .C2(n4855), .A(n4851), .B(n4850), .ZN(n5565)
         );
  AOI21_X2 U6380 ( .B1(n8235), .B2(n4870), .A(n4869), .ZN(n4868) );
  INV_X1 U6381 ( .A(n8350), .ZN(n4875) );
  NAND2_X1 U6382 ( .A1(n8363), .A2(n5677), .ZN(n8349) );
  AND2_X1 U6383 ( .A1(n4878), .A2(n5927), .ZN(n5932) );
  NAND2_X1 U6384 ( .A1(n9219), .A2(n7889), .ZN(n4880) );
  NAND2_X1 U6385 ( .A1(n7583), .A2(n7509), .ZN(n4890) );
  NAND2_X1 U6386 ( .A1(n9068), .A2(n7509), .ZN(n4889) );
  NAND2_X1 U6387 ( .A1(n4890), .A2(n4888), .ZN(n7512) );
  NAND2_X1 U6388 ( .A1(n5924), .A2(n6472), .ZN(n5941) );
  INV_X1 U6389 ( .A(n8455), .ZN(n8228) );
  NAND2_X1 U6390 ( .A1(n5923), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5924) );
  NAND2_X1 U6391 ( .A1(n8225), .A2(n8209), .ZN(n8208) );
  INV_X1 U6392 ( .A(n5990), .ZN(n5993) );
  NAND2_X1 U6393 ( .A1(n5774), .A2(n4263), .ZN(n5757) );
  NAND2_X1 U6394 ( .A1(n5904), .A2(n5903), .ZN(n5905) );
  NAND2_X1 U6395 ( .A1(n5749), .A2(P2_IR_REG_28__SCAN_IN), .ZN(n4981) );
  OR2_X1 U6396 ( .A1(n8184), .A2(n7841), .ZN(n7851) );
  NAND2_X1 U6397 ( .A1(n6868), .A2(n7163), .ZN(n5609) );
  XNOR2_X1 U6398 ( .A(n5126), .B(n5125), .ZN(n6600) );
  AND2_X1 U6399 ( .A1(n7735), .A2(n7724), .ZN(n5172) );
  AND2_X2 U6400 ( .A1(n5549), .A2(n6575), .ZN(n5062) );
  NAND3_X2 U6401 ( .A1(n4982), .A2(n4981), .A3(n4980), .ZN(n5549) );
  AOI21_X2 U6402 ( .B1(n9233), .B2(n9239), .A(n7888), .ZN(n9219) );
  OR2_X1 U6403 ( .A1(n4264), .A2(n9122), .ZN(n5997) );
  OR2_X1 U6404 ( .A1(n6053), .A2(n9698), .ZN(n5982) );
  OR2_X1 U6405 ( .A1(n4264), .A2(n7892), .ZN(n6492) );
  OR2_X1 U6406 ( .A1(n4264), .A2(n9235), .ZN(n6416) );
  OR2_X1 U6407 ( .A1(n4264), .A2(n9250), .ZN(n6393) );
  OAI21_X1 U6408 ( .B1(n9313), .B2(n4264), .A(n6336), .ZN(n9324) );
  OAI21_X1 U6409 ( .B1(n9326), .B2(n4264), .A(n6316), .ZN(n9346) );
  AND2_X1 U6410 ( .A1(n5760), .A2(n7162), .ZN(n7021) );
  AOI22_X2 U6411 ( .A1(n7300), .A2(n7299), .B1(n5789), .B2(n5788), .ZN(n7448)
         );
  AND2_X1 U6412 ( .A1(n9446), .A2(n9759), .ZN(n4903) );
  AND2_X1 U6413 ( .A1(n8450), .A2(n8553), .ZN(n4904) );
  INV_X1 U6414 ( .A(n6397), .ZN(n6445) );
  AND2_X1 U6415 ( .A1(n4386), .A2(n9012), .ZN(n4905) );
  INV_X1 U6416 ( .A(n8796), .ZN(n7887) );
  INV_X1 U6417 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n5942) );
  AND2_X1 U6418 ( .A1(n6806), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n4910) );
  NAND2_X1 U6419 ( .A1(n5762), .A2(n5763), .ZN(n6942) );
  AND4_X2 U6420 ( .A1(n4979), .A2(n4978), .A3(n4977), .A4(n4976), .ZN(n4911)
         );
  INV_X1 U6421 ( .A(n8053), .ZN(n7828) );
  NOR2_X1 U6422 ( .A1(n8938), .A2(n9694), .ZN(n4912) );
  INV_X1 U6423 ( .A(n9862), .ZN(n9860) );
  OR2_X1 U6424 ( .A1(n7308), .A2(n7309), .ZN(n4913) );
  INV_X1 U6425 ( .A(n9472), .ZN(n9238) );
  OR3_X1 U6426 ( .A1(n8634), .A2(n8636), .A3(n8781), .ZN(n4914) );
  INV_X1 U6427 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n4967) );
  OR2_X1 U6428 ( .A1(n7363), .A2(n9112), .ZN(n7506) );
  AOI21_X1 U6429 ( .B1(n7902), .B2(n9012), .A(n4386), .ZN(n7903) );
  OR2_X1 U6430 ( .A1(n8444), .A2(n5550), .ZN(n5719) );
  AND2_X1 U6431 ( .A1(n8144), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n8145) );
  INV_X1 U6432 ( .A(n8164), .ZN(n8165) );
  INV_X1 U6433 ( .A(n7735), .ZN(n7650) );
  INV_X1 U6434 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n5026) );
  INV_X1 U6435 ( .A(n8925), .ZN(n8927) );
  OR2_X1 U6436 ( .A1(n9192), .A2(n9445), .ZN(n9193) );
  INV_X1 U6437 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n6183) );
  NOR2_X1 U6438 ( .A1(n5351), .A2(n5350), .ZN(n5352) );
  NOR2_X1 U6439 ( .A1(n5270), .A2(n5269), .ZN(n5271) );
  INV_X1 U6440 ( .A(n5109), .ZN(n4944) );
  INV_X1 U6441 ( .A(n5116), .ZN(n4998) );
  INV_X1 U6442 ( .A(n5850), .ZN(n5836) );
  NAND2_X1 U6443 ( .A1(n5759), .A2(n5758), .ZN(n6923) );
  OR2_X1 U6444 ( .A1(n9801), .A2(n5880), .ZN(n7014) );
  OR2_X1 U6445 ( .A1(n8072), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n8073) );
  INV_X1 U6446 ( .A(n5568), .ZN(n5588) );
  INV_X1 U6447 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n5313) );
  INV_X1 U6448 ( .A(n5991), .ZN(n5992) );
  INV_X1 U6449 ( .A(n8633), .ZN(n6325) );
  AND2_X1 U6450 ( .A1(n7318), .A2(n9563), .ZN(n6509) );
  INV_X1 U6451 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n9972) );
  INV_X1 U6452 ( .A(n9198), .ZN(n9445) );
  NAND2_X1 U6453 ( .A1(n5379), .A2(n5378), .ZN(n5395) );
  AOI21_X1 U6454 ( .B1(n5358), .B2(n5357), .A(n5356), .ZN(n5359) );
  INV_X1 U6455 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n5922) );
  AOI21_X1 U6456 ( .B1(n5203), .B2(n5202), .A(n5201), .ZN(n5204) );
  NAND2_X1 U6457 ( .A1(n4955), .A2(n4954), .ZN(n4960) );
  NAND2_X1 U6458 ( .A1(n5894), .A2(n5893), .ZN(n5895) );
  XNOR2_X1 U6459 ( .A(n5768), .B(n5767), .ZN(n7059) );
  OR2_X1 U6460 ( .A1(n5884), .A2(n7014), .ZN(n8024) );
  OAI21_X1 U6461 ( .B1(n6869), .B2(n5562), .A(n7343), .ZN(n5563) );
  OR2_X1 U6462 ( .A1(n8272), .A2(n4995), .ZN(n5428) );
  AND2_X1 U6463 ( .A1(n8492), .A2(n8351), .ZN(n7833) );
  NOR2_X1 U6464 ( .A1(n8502), .A2(n7828), .ZN(n7829) );
  INV_X1 U6465 ( .A(n8175), .ZN(n8441) );
  OR2_X1 U6466 ( .A1(n7019), .A2(n6719), .ZN(n8404) );
  AND2_X1 U6467 ( .A1(n6106), .A2(n6105), .ZN(n6107) );
  NAND2_X1 U6468 ( .A1(n4914), .A2(n6325), .ZN(n6326) );
  OR2_X1 U6469 ( .A1(n4264), .A2(n9208), .ZN(n6441) );
  OR2_X1 U6470 ( .A1(n6643), .A2(P1_U3084), .ZN(n6625) );
  INV_X1 U6471 ( .A(n9694), .ZN(n9169) );
  INV_X1 U6472 ( .A(n9462), .ZN(n9211) );
  NOR2_X1 U6473 ( .A1(n9253), .A2(n7900), .ZN(n7885) );
  INV_X1 U6474 ( .A(n9106), .ZN(n9417) );
  AND2_X1 U6475 ( .A1(n8894), .A2(n8966), .ZN(n9076) );
  INV_X1 U6476 ( .A(n9754), .ZN(n9737) );
  AND2_X1 U6477 ( .A1(n5468), .A2(n5454), .ZN(n5466) );
  NAND2_X1 U6478 ( .A1(n5395), .A2(n5381), .ZN(n5396) );
  XNOR2_X1 U6479 ( .A(n5309), .B(SI_18_), .ZN(n5306) );
  XNOR2_X1 U6480 ( .A(n5224), .B(SI_14_), .ZN(n5222) );
  XNOR2_X1 U6481 ( .A(n4962), .B(SI_11_), .ZN(n5007) );
  XNOR2_X1 U6482 ( .A(n5110), .B(n5109), .ZN(n6096) );
  NOR2_X1 U6483 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n10054), .ZN(n9591) );
  OAI21_X1 U6484 ( .B1(n8228), .B2(n8029), .A(n5909), .ZN(n5910) );
  AND2_X1 U6485 ( .A1(n6867), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8042) );
  AOI21_X1 U6486 ( .B1(n8188), .B2(n5514), .A(n5513), .ZN(n8203) );
  AND2_X1 U6487 ( .A1(n5346), .A2(n5345), .ZN(n7932) );
  AND2_X1 U6488 ( .A1(n6724), .A2(n6723), .ZN(n8167) );
  AND2_X1 U6489 ( .A1(n6720), .A2(n8589), .ZN(n8164) );
  AND2_X1 U6490 ( .A1(n5885), .A2(n6719), .ZN(n8423) );
  INV_X1 U6491 ( .A(n9792), .ZN(n8439) );
  INV_X1 U6492 ( .A(n8414), .ZN(n9793) );
  NAND2_X1 U6493 ( .A1(n5872), .A2(n5871), .ZN(n7115) );
  OR2_X1 U6494 ( .A1(n8396), .A2(n8395), .ZN(n8516) );
  INV_X1 U6495 ( .A(n9851), .ZN(n8544) );
  INV_X1 U6496 ( .A(n7115), .ZN(n7853) );
  AND4_X1 U6497 ( .A1(n6494), .A2(n6493), .A3(n6492), .A4(n6491), .ZN(n9189)
         );
  INV_X1 U6498 ( .A(n9620), .ZN(n9648) );
  AND2_X1 U6499 ( .A1(n9164), .A2(n9574), .ZN(n9627) );
  INV_X1 U6500 ( .A(n9433), .ZN(n9174) );
  AND2_X1 U6501 ( .A1(n8939), .A2(n6895), .ZN(n9396) );
  INV_X1 U6502 ( .A(n9354), .ZN(n9407) );
  AND2_X1 U6503 ( .A1(n9713), .A2(n9693), .ZN(n9426) );
  AND2_X1 U6504 ( .A1(n9710), .A2(n9740), .ZN(n9745) );
  INV_X1 U6505 ( .A(n9745), .ZN(n9759) );
  AND2_X1 U6506 ( .A1(n6756), .A2(n6755), .ZN(n6918) );
  INV_X1 U6507 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n6473) );
  INV_X1 U6508 ( .A(n8171), .ZN(n8088) );
  INV_X1 U6509 ( .A(n8042), .ZN(n8023) );
  NAND2_X1 U6510 ( .A1(n5414), .A2(n5413), .ZN(n8266) );
  OR2_X1 U6511 ( .A1(n7218), .A2(n5873), .ZN(n9792) );
  NAND2_X2 U6512 ( .A1(n7016), .A2(n8411), .ZN(n9798) );
  INV_X1 U6513 ( .A(n9871), .ZN(n9874) );
  NOR2_X2 U6514 ( .A1(n7854), .A2(n7115), .ZN(n9870) );
  INV_X1 U6515 ( .A(n9802), .ZN(n9903) );
  XNOR2_X1 U6516 ( .A(n5745), .B(n5732), .ZN(n7493) );
  INV_X1 U6517 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n6796) );
  INV_X1 U6518 ( .A(n9514), .ZN(n9368) );
  INV_X1 U6519 ( .A(n8812), .ZN(n8801) );
  INV_X1 U6520 ( .A(n9189), .ZN(n9214) );
  INV_X1 U6521 ( .A(n7882), .ZN(n9310) );
  INV_X1 U6522 ( .A(n9627), .ZN(n9654) );
  INV_X1 U6523 ( .A(n9426), .ZN(n9683) );
  AND2_X2 U6524 ( .A1(n6918), .A2(n9563), .ZN(n9785) );
  AND2_X2 U6525 ( .A1(n6918), .A2(n6917), .ZN(n9776) );
  OR2_X1 U6526 ( .A1(n9718), .A2(n9722), .ZN(n9720) );
  AND2_X1 U6527 ( .A1(n6471), .A2(n6470), .ZN(n9563) );
  INV_X1 U6528 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n6852) );
  INV_X1 U6529 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n6614) );
  NOR2_X1 U6530 ( .A1(n10065), .A2(n10064), .ZN(n10063) );
  NOR2_X1 U6531 ( .A1(n9902), .A2(n9901), .ZN(n9900) );
  INV_X1 U6532 ( .A(n5029), .ZN(n4934) );
  NOR2_X1 U6533 ( .A1(P2_DATAO_REG_1__SCAN_IN), .A2(SI_1_), .ZN(n4924) );
  AND2_X1 U6534 ( .A1(SI_0_), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n5038) );
  INV_X1 U6535 ( .A(n5038), .ZN(n4923) );
  NAND2_X1 U6536 ( .A1(P2_DATAO_REG_1__SCAN_IN), .A2(SI_1_), .ZN(n4922) );
  OAI21_X1 U6537 ( .B1(n4924), .B2(n4923), .A(n4922), .ZN(n4925) );
  NOR2_X1 U6538 ( .A1(SI_1_), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n4927) );
  NAND2_X1 U6539 ( .A1(SI_0_), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n5039) );
  NAND2_X1 U6540 ( .A1(SI_1_), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n4926) );
  OAI21_X1 U6541 ( .B1(n4927), .B2(n5039), .A(n4926), .ZN(n4928) );
  NAND2_X1 U6542 ( .A1(n4921), .A2(n4928), .ZN(n4929) );
  NAND2_X1 U6543 ( .A1(n4930), .A2(n4929), .ZN(n5059) );
  INV_X1 U6544 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n6561) );
  INV_X1 U6545 ( .A(SI_2_), .ZN(n4931) );
  INV_X1 U6546 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n6598) );
  NAND2_X1 U6547 ( .A1(n4935), .A2(SI_3_), .ZN(n4936) );
  XNOR2_X1 U6548 ( .A(n4938), .B(SI_4_), .ZN(n5075) );
  INV_X1 U6549 ( .A(n5075), .ZN(n4937) );
  NAND2_X1 U6550 ( .A1(n4938), .A2(SI_4_), .ZN(n4939) );
  NAND2_X1 U6551 ( .A1(n4940), .A2(SI_5_), .ZN(n4941) );
  INV_X1 U6552 ( .A(n5093), .ZN(n4942) );
  NAND2_X1 U6553 ( .A1(n4945), .A2(SI_7_), .ZN(n4946) );
  INV_X1 U6554 ( .A(SI_8_), .ZN(n4947) );
  INV_X1 U6555 ( .A(n4948), .ZN(n4949) );
  NAND2_X1 U6556 ( .A1(n4949), .A2(SI_8_), .ZN(n4950) );
  INV_X1 U6557 ( .A(SI_9_), .ZN(n4952) );
  NAND2_X1 U6558 ( .A1(n4958), .A2(n4952), .ZN(n5153) );
  AND2_X1 U6559 ( .A1(n5139), .A2(n5153), .ZN(n4953) );
  INV_X1 U6560 ( .A(SI_10_), .ZN(n4954) );
  INV_X1 U6561 ( .A(n4955), .ZN(n4956) );
  NAND2_X1 U6562 ( .A1(n4956), .A2(SI_10_), .ZN(n4957) );
  INV_X1 U6563 ( .A(n4958), .ZN(n4959) );
  NAND2_X1 U6564 ( .A1(n4959), .A2(SI_9_), .ZN(n5141) );
  INV_X1 U6565 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n4961) );
  INV_X1 U6566 ( .A(n4962), .ZN(n4963) );
  NAND2_X1 U6567 ( .A1(n4963), .A2(SI_11_), .ZN(n5194) );
  INV_X1 U6568 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n6761) );
  INV_X1 U6569 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n6759) );
  INV_X1 U6570 ( .A(SI_12_), .ZN(n4964) );
  NAND2_X1 U6571 ( .A1(n4965), .A2(n4964), .ZN(n5199) );
  INV_X1 U6572 ( .A(n4965), .ZN(n4966) );
  NAND2_X1 U6573 ( .A1(n4966), .A2(SI_12_), .ZN(n5195) );
  NAND2_X1 U6574 ( .A1(n5199), .A2(n5195), .ZN(n5173) );
  NOR2_X2 U6576 ( .A1(n5253), .A2(P2_IR_REG_17__SCAN_IN), .ZN(n4975) );
  NOR2_X2 U6577 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_3__SCAN_IN), .ZN(
        n4969) );
  NOR2_X2 U6578 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_4__SCAN_IN), .ZN(
        n4968) );
  AND3_X2 U6579 ( .A1(n4969), .A2(n4968), .A3(n5026), .ZN(n4983) );
  NOR2_X1 U6580 ( .A1(P2_IR_REG_7__SCAN_IN), .A2(P2_IR_REG_5__SCAN_IN), .ZN(
        n4974) );
  INV_X2 U6581 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n5555) );
  NOR2_X1 U6582 ( .A1(P2_IR_REG_26__SCAN_IN), .A2(P2_IR_REG_24__SCAN_IN), .ZN(
        n4978) );
  NOR2_X1 U6583 ( .A1(P2_IR_REG_22__SCAN_IN), .A2(P2_IR_REG_23__SCAN_IN), .ZN(
        n4977) );
  NOR2_X1 U6584 ( .A1(P2_IR_REG_21__SCAN_IN), .A2(P2_IR_REG_18__SCAN_IN), .ZN(
        n4976) );
  NAND2_X1 U6585 ( .A1(n4990), .A2(P2_IR_REG_27__SCAN_IN), .ZN(n4980) );
  NAND2_X1 U6586 ( .A1(n6758), .A2(n5474), .ZN(n4989) );
  INV_X1 U6587 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n4984) );
  NAND2_X1 U6588 ( .A1(n4983), .A2(n4984), .ZN(n5095) );
  NOR2_X1 U6589 ( .A1(n5095), .A2(P2_IR_REG_6__SCAN_IN), .ZN(n5111) );
  INV_X1 U6590 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n4985) );
  NAND2_X1 U6591 ( .A1(n5111), .A2(n4985), .ZN(n5255) );
  NOR2_X1 U6592 ( .A1(n5156), .A2(P2_IR_REG_10__SCAN_IN), .ZN(n5009) );
  INV_X1 U6593 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n4986) );
  NAND2_X1 U6594 ( .A1(n5009), .A2(n4986), .ZN(n5181) );
  NAND2_X1 U6595 ( .A1(n5181), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4987) );
  XNOR2_X1 U6596 ( .A(n4987), .B(P2_IR_REG_12__SCAN_IN), .ZN(n7793) );
  AOI22_X1 U6597 ( .A1(n7793), .A2(n5315), .B1(n5507), .B2(
        P1_DATAO_REG_12__SCAN_IN), .ZN(n4988) );
  INV_X1 U6598 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n4991) );
  NAND2_X1 U6599 ( .A1(n4993), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4994) );
  INV_X4 U6600 ( .A(n5080), .ZN(n5529) );
  NAND2_X1 U6601 ( .A1(n5529), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n5006) );
  NAND2_X1 U6602 ( .A1(n5118), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n5005) );
  INV_X4 U6603 ( .A(n4995), .ZN(n5514) );
  NAND2_X1 U6604 ( .A1(n5015), .A2(n5000), .ZN(n5001) );
  AND2_X1 U6605 ( .A1(n5187), .A2(n5001), .ZN(n7730) );
  NAND2_X1 U6606 ( .A1(n5514), .A2(n7730), .ZN(n5004) );
  INV_X1 U6607 ( .A(n5002), .ZN(n8585) );
  NAND2_X1 U6608 ( .A1(n5537), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n5003) );
  NAND2_X1 U6609 ( .A1(n8535), .A2(n7993), .ZN(n5654) );
  NAND2_X1 U6610 ( .A1(n6608), .A2(n5474), .ZN(n5012) );
  OR2_X1 U6611 ( .A1(n5009), .A2(n4991), .ZN(n5010) );
  XNOR2_X1 U6612 ( .A(n5010), .B(P2_IR_REG_11__SCAN_IN), .ZN(n7764) );
  AOI22_X1 U6613 ( .A1(n7764), .A2(n5315), .B1(n5507), .B2(
        P1_DATAO_REG_11__SCAN_IN), .ZN(n5011) );
  NAND2_X1 U6614 ( .A1(n5529), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n5019) );
  NAND2_X1 U6615 ( .A1(n5118), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n5018) );
  INV_X1 U6616 ( .A(n5013), .ZN(n5163) );
  INV_X1 U6617 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n6545) );
  NAND2_X1 U6618 ( .A1(n5163), .A2(n6545), .ZN(n5014) );
  AND2_X1 U6619 ( .A1(n5015), .A2(n5014), .ZN(n7691) );
  NAND2_X1 U6620 ( .A1(n5514), .A2(n7691), .ZN(n5017) );
  NAND2_X1 U6621 ( .A1(n5537), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n5016) );
  NAND2_X1 U6622 ( .A1(n8540), .A2(n7627), .ZN(n7724) );
  INV_X1 U6623 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n5068) );
  NAND2_X1 U6624 ( .A1(n5102), .A2(n5068), .ZN(n5022) );
  NAND2_X1 U6625 ( .A1(n5098), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n5021) );
  NAND2_X1 U6626 ( .A1(n5262), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n5020) );
  INV_X1 U6627 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n5025) );
  INV_X1 U6628 ( .A(n5057), .ZN(n5027) );
  NAND2_X1 U6629 ( .A1(n5027), .A2(n5026), .ZN(n5076) );
  NAND2_X1 U6630 ( .A1(n5076), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5028) );
  XNOR2_X1 U6631 ( .A(n5029), .B(n5030), .ZN(n6565) );
  NAND2_X1 U6632 ( .A1(n6565), .A2(n5062), .ZN(n5031) );
  NAND2_X1 U6633 ( .A1(n7131), .A2(n7077), .ZN(n5617) );
  NAND2_X1 U6634 ( .A1(n5617), .A2(n5623), .ZN(n7129) );
  NAND2_X1 U6635 ( .A1(n5102), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n5036) );
  INV_X1 U6636 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n5033) );
  OR2_X1 U6637 ( .A1(n5051), .A2(n5033), .ZN(n5035) );
  NAND2_X1 U6638 ( .A1(n5098), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n5034) );
  INV_X1 U6639 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n6567) );
  XNOR2_X1 U6640 ( .A(n5040), .B(SI_1_), .ZN(n5042) );
  XNOR2_X1 U6641 ( .A(n5042), .B(n5041), .ZN(n6566) );
  NAND2_X1 U6642 ( .A1(n5062), .A2(n6566), .ZN(n5044) );
  INV_X1 U6643 ( .A(n6737), .ZN(n6732) );
  NAND2_X1 U6644 ( .A1(n5315), .A2(n6732), .ZN(n5043) );
  OAI211_X2 U6645 ( .C1(n5526), .C2(n6567), .A(n5044), .B(n5043), .ZN(n7163)
         );
  NAND2_X1 U6646 ( .A1(n5102), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n5047) );
  NAND2_X1 U6647 ( .A1(n5098), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n5046) );
  NAND2_X1 U6648 ( .A1(n6575), .A2(SI_0_), .ZN(n5048) );
  XNOR2_X1 U6649 ( .A(n5048), .B(P1_DATAO_REG_0__SCAN_IN), .ZN(n8590) );
  MUX2_X1 U6650 ( .A(P2_IR_REG_0__SCAN_IN), .B(n8590), .S(n5549), .Z(n7162) );
  NAND2_X1 U6651 ( .A1(n5609), .A2(n7165), .ZN(n5049) );
  NAND2_X1 U6652 ( .A1(n5262), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n5055) );
  NAND2_X1 U6653 ( .A1(n5102), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n5054) );
  NAND2_X1 U6654 ( .A1(n5098), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n5053) );
  INV_X1 U6655 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n5050) );
  NAND2_X1 U6656 ( .A1(n5056), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n5065) );
  NAND2_X1 U6657 ( .A1(n5057), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5058) );
  NAND2_X1 U6658 ( .A1(n5315), .A2(n6806), .ZN(n5064) );
  XNOR2_X1 U6659 ( .A(n5059), .B(SI_2_), .ZN(n5061) );
  XNOR2_X1 U6660 ( .A(n5061), .B(n5060), .ZN(n6560) );
  NAND2_X1 U6661 ( .A1(n5062), .A2(n6560), .ZN(n5063) );
  OR2_X2 U6662 ( .A1(n8066), .A2(n7124), .ZN(n5607) );
  NAND2_X1 U6663 ( .A1(n8066), .A2(n7124), .ZN(n5610) );
  NAND2_X2 U6664 ( .A1(n5607), .A2(n5610), .ZN(n7066) );
  NAND2_X1 U6665 ( .A1(n7079), .A2(n7078), .ZN(n5066) );
  NAND2_X1 U6666 ( .A1(n5066), .A2(n5617), .ZN(n7137) );
  NAND2_X1 U6667 ( .A1(n5262), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n5073) );
  NAND2_X1 U6668 ( .A1(n5118), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n5072) );
  INV_X1 U6669 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n5067) );
  NAND2_X1 U6670 ( .A1(n5068), .A2(n5067), .ZN(n5069) );
  AND2_X1 U6671 ( .A1(n5069), .A2(n5082), .ZN(n7142) );
  NAND2_X1 U6672 ( .A1(n5514), .A2(n7142), .ZN(n5071) );
  NAND2_X1 U6673 ( .A1(n5537), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n5070) );
  AND4_X2 U6674 ( .A1(n5073), .A2(n5072), .A3(n5071), .A4(n5070), .ZN(n7177)
         );
  XNOR2_X1 U6675 ( .A(n5075), .B(n5074), .ZN(n6563) );
  NAND2_X1 U6676 ( .A1(n6563), .A2(n5062), .ZN(n5079) );
  OAI21_X1 U6677 ( .B1(n5076), .B2(P2_IR_REG_3__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5077) );
  AOI22_X1 U6678 ( .A1(n5056), .A2(P1_DATAO_REG_4__SCAN_IN), .B1(n5315), .B2(
        n6832), .ZN(n5078) );
  NAND2_X1 U6679 ( .A1(n5079), .A2(n5078), .ZN(n7145) );
  NAND2_X1 U6680 ( .A1(n7177), .A2(n7145), .ZN(n7135) );
  NAND2_X1 U6681 ( .A1(n5118), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n5087) );
  NAND2_X1 U6682 ( .A1(n5262), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n5086) );
  INV_X1 U6683 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n5081) );
  NAND2_X1 U6684 ( .A1(n5082), .A2(n5081), .ZN(n5083) );
  AND2_X1 U6685 ( .A1(n5100), .A2(n5083), .ZN(n7088) );
  NAND2_X1 U6686 ( .A1(n5514), .A2(n7088), .ZN(n5085) );
  NAND2_X1 U6687 ( .A1(n5537), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n5084) );
  OR2_X1 U6688 ( .A1(n4983), .A2(n4991), .ZN(n5090) );
  XNOR2_X1 U6689 ( .A(n5090), .B(P2_IR_REG_5__SCAN_IN), .ZN(n6844) );
  AOI22_X1 U6690 ( .A1(n5507), .A2(P1_DATAO_REG_5__SCAN_IN), .B1(n5315), .B2(
        n6844), .ZN(n5091) );
  NAND2_X1 U6691 ( .A1(n5095), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5096) );
  AOI22_X1 U6692 ( .A1(n5507), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n5315), .B2(
        n6908), .ZN(n5097) );
  NAND2_X1 U6693 ( .A1(n5529), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n5106) );
  NAND2_X1 U6694 ( .A1(n5098), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n5105) );
  INV_X1 U6695 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n5099) );
  NAND2_X1 U6696 ( .A1(n5100), .A2(n5099), .ZN(n5101) );
  AND2_X1 U6697 ( .A1(n5116), .A2(n5101), .ZN(n7221) );
  NAND2_X1 U6698 ( .A1(n5102), .A2(n7221), .ZN(n5104) );
  NAND2_X1 U6699 ( .A1(n5118), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n5103) );
  NAND4_X1 U6700 ( .A1(n5106), .A2(n5105), .A3(n5104), .A4(n5103), .ZN(n8062)
         );
  AND2_X2 U6701 ( .A1(n5627), .A2(n5633), .ZN(n7225) );
  NAND2_X1 U6702 ( .A1(n7214), .A2(n7213), .ZN(n5107) );
  NAND2_X1 U6703 ( .A1(n5108), .A2(n5633), .ZN(n7182) );
  NAND2_X1 U6704 ( .A1(n6096), .A2(n5474), .ZN(n5114) );
  OR2_X1 U6705 ( .A1(n5111), .A2(n4991), .ZN(n5112) );
  XNOR2_X1 U6706 ( .A(n5112), .B(P2_IR_REG_7__SCAN_IN), .ZN(n7043) );
  AOI22_X1 U6707 ( .A1(n5507), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n5315), .B2(
        n7043), .ZN(n5113) );
  NAND2_X1 U6708 ( .A1(n5114), .A2(n5113), .ZN(n7412) );
  NAND2_X1 U6709 ( .A1(n5529), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n5122) );
  NAND2_X1 U6710 ( .A1(n5537), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n5121) );
  INV_X1 U6711 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n5115) );
  NAND2_X1 U6712 ( .A1(n5116), .A2(n5115), .ZN(n5117) );
  AND2_X1 U6713 ( .A1(n5132), .A2(n5117), .ZN(n7196) );
  NAND2_X1 U6714 ( .A1(n5514), .A2(n7196), .ZN(n5120) );
  NAND2_X1 U6715 ( .A1(n5118), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n5119) );
  NAND2_X1 U6716 ( .A1(n7412), .A2(n7416), .ZN(n5634) );
  INV_X1 U6717 ( .A(n5634), .ZN(n5123) );
  OR2_X1 U6718 ( .A1(n7412), .A2(n7416), .ZN(n5635) );
  NAND2_X1 U6719 ( .A1(n6600), .A2(n5474), .ZN(n5130) );
  NAND2_X1 U6720 ( .A1(n5255), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5127) );
  MUX2_X1 U6721 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5127), .S(
        P2_IR_REG_8__SCAN_IN), .Z(n5128) );
  AND2_X1 U6722 ( .A1(n5128), .A2(n5142), .ZN(n7292) );
  AOI22_X1 U6723 ( .A1(n5507), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n7292), .B2(
        n5315), .ZN(n5129) );
  NAND2_X1 U6724 ( .A1(n5130), .A2(n5129), .ZN(n7429) );
  NAND2_X1 U6725 ( .A1(n5118), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n5137) );
  NAND2_X1 U6726 ( .A1(n5529), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n5136) );
  INV_X1 U6727 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n5131) );
  NAND2_X1 U6728 ( .A1(n5132), .A2(n5131), .ZN(n5133) );
  AND2_X1 U6729 ( .A1(n5162), .A2(n5133), .ZN(n7420) );
  NAND2_X1 U6730 ( .A1(n5514), .A2(n7420), .ZN(n5135) );
  NAND2_X1 U6731 ( .A1(n5537), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n5134) );
  NAND4_X1 U6732 ( .A1(n5137), .A2(n5136), .A3(n5135), .A4(n5134), .ZN(n8060)
         );
  INV_X1 U6733 ( .A(n8060), .ZN(n7452) );
  OR2_X1 U6734 ( .A1(n7429), .A2(n7452), .ZN(n5637) );
  NAND2_X1 U6735 ( .A1(n7429), .A2(n7452), .ZN(n7432) );
  NAND2_X1 U6736 ( .A1(n5637), .A2(n7432), .ZN(n7560) );
  AND2_X1 U6737 ( .A1(n5153), .A2(n5141), .ZN(n5151) );
  NAND2_X1 U6738 ( .A1(n6604), .A2(n5474), .ZN(n5145) );
  NAND2_X1 U6739 ( .A1(n5142), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5143) );
  XNOR2_X1 U6740 ( .A(n5143), .B(P2_IR_REG_9__SCAN_IN), .ZN(n7467) );
  AOI22_X1 U6741 ( .A1(n7467), .A2(n5315), .B1(n5507), .B2(
        P1_DATAO_REG_9__SCAN_IN), .ZN(n5144) );
  NAND2_X2 U6742 ( .A1(n5145), .A2(n5144), .ZN(n8552) );
  NAND2_X1 U6743 ( .A1(n5529), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n5149) );
  NAND2_X1 U6744 ( .A1(n5537), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n5148) );
  XNOR2_X1 U6745 ( .A(n5162), .B(P2_REG3_REG_9__SCAN_IN), .ZN(n7454) );
  NAND2_X1 U6746 ( .A1(n5514), .A2(n7454), .ZN(n5147) );
  NAND2_X1 U6747 ( .A1(n5118), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n5146) );
  NAND2_X1 U6748 ( .A1(n8552), .A2(n7556), .ZN(n5640) );
  AND2_X1 U6749 ( .A1(n5640), .A2(n7432), .ZN(n5150) );
  NAND2_X1 U6750 ( .A1(n7433), .A2(n5150), .ZN(n7554) );
  NAND2_X1 U6751 ( .A1(n5152), .A2(n5151), .ZN(n5154) );
  NAND2_X1 U6752 ( .A1(n6610), .A2(n5474), .ZN(n5159) );
  NAND2_X1 U6753 ( .A1(n5156), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5157) );
  XNOR2_X1 U6754 ( .A(n5157), .B(P2_IR_REG_10__SCAN_IN), .ZN(n7541) );
  AOI22_X1 U6755 ( .A1(n7541), .A2(n5315), .B1(n5507), .B2(
        P1_DATAO_REG_10__SCAN_IN), .ZN(n5158) );
  NAND2_X1 U6756 ( .A1(n5118), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n5168) );
  NAND2_X1 U6757 ( .A1(n5529), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n5167) );
  INV_X1 U6758 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n5161) );
  INV_X1 U6759 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n5160) );
  OAI21_X1 U6760 ( .B1(n5162), .B2(n5161), .A(n5160), .ZN(n5164) );
  AND2_X1 U6761 ( .A1(n5164), .A2(n5163), .ZN(n7572) );
  NAND2_X1 U6762 ( .A1(n5514), .A2(n7572), .ZN(n5166) );
  NAND2_X1 U6763 ( .A1(n5537), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n5165) );
  OR2_X1 U6764 ( .A1(n8546), .A2(n7435), .ZN(n5566) );
  OR2_X1 U6765 ( .A1(n8552), .A2(n7556), .ZN(n7553) );
  AND2_X1 U6766 ( .A1(n5566), .A2(n7553), .ZN(n5644) );
  NAND2_X1 U6767 ( .A1(n7554), .A2(n5644), .ZN(n5169) );
  NAND2_X1 U6768 ( .A1(n8546), .A2(n7435), .ZN(n5642) );
  NAND2_X1 U6769 ( .A1(n5169), .A2(n5642), .ZN(n7693) );
  OAI21_X1 U6770 ( .B1(n5174), .B2(n5173), .A(n5199), .ZN(n5180) );
  INV_X1 U6771 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n5175) );
  INV_X1 U6772 ( .A(SI_13_), .ZN(n5176) );
  NAND2_X1 U6773 ( .A1(n5177), .A2(n5176), .ZN(n5200) );
  INV_X1 U6774 ( .A(n5177), .ZN(n5178) );
  NAND2_X1 U6775 ( .A1(n5178), .A2(SI_13_), .ZN(n5179) );
  NAND2_X1 U6776 ( .A1(n5200), .A2(n5179), .ZN(n5197) );
  INV_X1 U6777 ( .A(n5197), .ZN(n5203) );
  XNOR2_X1 U6778 ( .A(n5180), .B(n5203), .ZN(n6793) );
  NAND2_X1 U6779 ( .A1(n6793), .A2(n5474), .ZN(n5184) );
  NAND2_X1 U6780 ( .A1(n5182), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5206) );
  XNOR2_X1 U6781 ( .A(n5206), .B(P2_IR_REG_13__SCAN_IN), .ZN(n8072) );
  AOI22_X1 U6782 ( .A1(n8072), .A2(n5315), .B1(n5507), .B2(
        P1_DATAO_REG_13__SCAN_IN), .ZN(n5183) );
  NAND2_X1 U6783 ( .A1(n5118), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n5192) );
  NAND2_X1 U6784 ( .A1(n5529), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n5191) );
  INV_X1 U6785 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n5186) );
  NAND2_X1 U6786 ( .A1(n5187), .A2(n5186), .ZN(n5188) );
  AND2_X1 U6787 ( .A1(n5214), .A2(n5188), .ZN(n7995) );
  NAND2_X1 U6788 ( .A1(n5514), .A2(n7995), .ZN(n5190) );
  NAND2_X1 U6789 ( .A1(n5537), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n5189) );
  NAND2_X1 U6790 ( .A1(n8529), .A2(n7741), .ZN(n5659) );
  NAND2_X1 U6791 ( .A1(n5195), .A2(n5194), .ZN(n5196) );
  NOR2_X1 U6792 ( .A1(n5197), .A2(n5196), .ZN(n5198) );
  INV_X1 U6793 ( .A(n5199), .ZN(n5202) );
  INV_X1 U6794 ( .A(n5200), .ZN(n5201) );
  XNOR2_X1 U6795 ( .A(n4668), .B(n5222), .ZN(n6795) );
  NAND2_X1 U6796 ( .A1(n6795), .A2(n5474), .ZN(n5212) );
  NAND2_X1 U6797 ( .A1(n5206), .A2(n5205), .ZN(n5207) );
  NAND2_X1 U6798 ( .A1(n5207), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5209) );
  NAND2_X1 U6799 ( .A1(n5209), .A2(n5208), .ZN(n5229) );
  OR2_X1 U6800 ( .A1(n5209), .A2(n5208), .ZN(n5210) );
  AOI22_X1 U6801 ( .A1(n8084), .A2(n5315), .B1(n5507), .B2(
        P1_DATAO_REG_14__SCAN_IN), .ZN(n5211) );
  INV_X1 U6802 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n5213) );
  OR2_X2 U6803 ( .A1(n5214), .A2(n5213), .ZN(n5234) );
  NAND2_X1 U6804 ( .A1(n5214), .A2(n5213), .ZN(n5215) );
  NAND2_X1 U6805 ( .A1(n5234), .A2(n5215), .ZN(n7813) );
  OR2_X1 U6806 ( .A1(n4995), .A2(n7813), .ZN(n5219) );
  NAND2_X1 U6807 ( .A1(n5118), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n5218) );
  NAND2_X1 U6808 ( .A1(n5529), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n5217) );
  NAND2_X1 U6809 ( .A1(n5537), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n5216) );
  NAND4_X1 U6810 ( .A1(n5219), .A2(n5218), .A3(n5217), .A4(n5216), .ZN(n8424)
         );
  NAND2_X1 U6811 ( .A1(n7751), .A2(n8424), .ZN(n5220) );
  INV_X1 U6812 ( .A(n8424), .ZN(n8038) );
  OR2_X1 U6813 ( .A1(n7751), .A2(n8038), .ZN(n5221) );
  INV_X1 U6814 ( .A(n5224), .ZN(n5225) );
  INV_X1 U6815 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n6967) );
  INV_X1 U6816 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n6965) );
  INV_X1 U6817 ( .A(SI_15_), .ZN(n5226) );
  NAND2_X1 U6818 ( .A1(n5227), .A2(n5226), .ZN(n5272) );
  INV_X1 U6819 ( .A(n5227), .ZN(n5228) );
  NAND2_X1 U6820 ( .A1(n5228), .A2(SI_15_), .ZN(n5268) );
  NAND2_X1 U6821 ( .A1(n5272), .A2(n5268), .ZN(n5242) );
  XNOR2_X1 U6822 ( .A(n5243), .B(n5242), .ZN(n6964) );
  NAND2_X1 U6823 ( .A1(n6964), .A2(n5474), .ZN(n5232) );
  NAND2_X1 U6824 ( .A1(n5229), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5230) );
  XNOR2_X1 U6825 ( .A(n5230), .B(P2_IR_REG_15__SCAN_IN), .ZN(n8099) );
  AOI22_X1 U6826 ( .A1(n8099), .A2(n5315), .B1(n5507), .B2(
        P1_DATAO_REG_15__SCAN_IN), .ZN(n5231) );
  INV_X1 U6827 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n5233) );
  NAND2_X1 U6828 ( .A1(n5234), .A2(n5233), .ZN(n5235) );
  AND2_X1 U6829 ( .A1(n5260), .A2(n5235), .ZN(n8431) );
  NAND2_X1 U6830 ( .A1(n8431), .A2(n5514), .ZN(n5240) );
  NAND2_X1 U6831 ( .A1(n5118), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n5237) );
  NAND2_X1 U6832 ( .A1(n5529), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n5236) );
  AND2_X1 U6833 ( .A1(n5237), .A2(n5236), .ZN(n5239) );
  NAND2_X1 U6834 ( .A1(n5537), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n5238) );
  NAND2_X1 U6835 ( .A1(n8517), .A2(n8403), .ZN(n5668) );
  NAND2_X1 U6836 ( .A1(n5669), .A2(n5668), .ZN(n8422) );
  INV_X1 U6837 ( .A(n8422), .ZN(n8434) );
  OAI21_X1 U6838 ( .B1(n5243), .B2(n5242), .A(n5272), .ZN(n5250) );
  INV_X1 U6839 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n5245) );
  INV_X1 U6840 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n5244) );
  INV_X1 U6841 ( .A(SI_16_), .ZN(n5246) );
  NAND2_X1 U6842 ( .A1(n5247), .A2(n5246), .ZN(n5273) );
  INV_X1 U6843 ( .A(n5247), .ZN(n5248) );
  NAND2_X1 U6844 ( .A1(n5248), .A2(SI_16_), .ZN(n5249) );
  NAND2_X1 U6845 ( .A1(n5273), .A2(n5249), .ZN(n5270) );
  INV_X1 U6846 ( .A(n5270), .ZN(n5276) );
  XNOR2_X1 U6847 ( .A(n5250), .B(n5276), .ZN(n6973) );
  NAND2_X1 U6848 ( .A1(n6973), .A2(n5474), .ZN(n5258) );
  INV_X1 U6849 ( .A(n5253), .ZN(n5254) );
  NAND2_X1 U6850 ( .A1(n5252), .A2(n5254), .ZN(n5281) );
  OAI21_X1 U6851 ( .B1(n5255), .B2(n5281), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n5256) );
  XNOR2_X1 U6852 ( .A(n5256), .B(P2_IR_REG_16__SCAN_IN), .ZN(n8128) );
  AOI22_X1 U6853 ( .A1(n8128), .A2(n5315), .B1(n5507), .B2(
        P1_DATAO_REG_16__SCAN_IN), .ZN(n5257) );
  INV_X1 U6854 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n5259) );
  NAND2_X1 U6855 ( .A1(n5260), .A2(n5259), .ZN(n5261) );
  NAND2_X1 U6856 ( .A1(n5287), .A2(n5261), .ZN(n8410) );
  OR2_X1 U6857 ( .A1(n8410), .A2(n4995), .ZN(n5265) );
  AOI22_X1 U6858 ( .A1(n5118), .A2(P2_REG0_REG_16__SCAN_IN), .B1(n5529), .B2(
        P2_REG1_REG_16__SCAN_IN), .ZN(n5264) );
  NAND2_X1 U6859 ( .A1(n5537), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n5263) );
  OR2_X1 U6860 ( .A1(n8512), .A2(n7825), .ZN(n5673) );
  NAND2_X1 U6861 ( .A1(n8512), .A2(n7825), .ZN(n8385) );
  INV_X1 U6862 ( .A(n8385), .ZN(n5292) );
  NAND2_X1 U6863 ( .A1(n5268), .A2(n5267), .ZN(n5269) );
  INV_X1 U6864 ( .A(n5272), .ZN(n5275) );
  INV_X1 U6865 ( .A(n5273), .ZN(n5274) );
  INV_X1 U6866 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n5278) );
  XNOR2_X1 U6867 ( .A(n5297), .B(n5294), .ZN(n6921) );
  NAND2_X1 U6868 ( .A1(n6921), .A2(n5474), .ZN(n5284) );
  NAND2_X1 U6869 ( .A1(n4983), .A2(n5279), .ZN(n5280) );
  OAI21_X1 U6870 ( .B1(n5281), .B2(n5280), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n5282) );
  XNOR2_X1 U6871 ( .A(n5282), .B(P2_IR_REG_17__SCAN_IN), .ZN(n8144) );
  AOI22_X1 U6872 ( .A1(n5507), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n5315), .B2(
        n8144), .ZN(n5283) );
  INV_X1 U6873 ( .A(n5287), .ZN(n5285) );
  INV_X1 U6874 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n5286) );
  NAND2_X1 U6875 ( .A1(n5287), .A2(n5286), .ZN(n5288) );
  NAND2_X1 U6876 ( .A1(n5321), .A2(n5288), .ZN(n8378) );
  OR2_X1 U6877 ( .A1(n8378), .A2(n4995), .ZN(n5291) );
  AOI22_X1 U6878 ( .A1(n5537), .A2(P2_REG2_REG_17__SCAN_IN), .B1(n5529), .B2(
        P2_REG1_REG_17__SCAN_IN), .ZN(n5290) );
  NAND2_X1 U6879 ( .A1(n5118), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n5289) );
  NAND2_X1 U6880 ( .A1(n8509), .A2(n8405), .ZN(n5598) );
  NAND2_X1 U6881 ( .A1(n5597), .A2(n5598), .ZN(n8373) );
  NOR2_X1 U6882 ( .A1(n5292), .A2(n8373), .ZN(n5293) );
  INV_X1 U6883 ( .A(n5295), .ZN(n5296) );
  XNOR2_X1 U6884 ( .A(n5308), .B(n5306), .ZN(n7097) );
  NAND2_X1 U6885 ( .A1(n7097), .A2(n5474), .ZN(n5301) );
  INV_X1 U6886 ( .A(n5314), .ZN(n5298) );
  NAND2_X1 U6887 ( .A1(n5298), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5299) );
  XNOR2_X1 U6888 ( .A(n5299), .B(P2_IR_REG_18__SCAN_IN), .ZN(n8151) );
  AOI22_X1 U6889 ( .A1(n5507), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n5315), .B2(
        n8151), .ZN(n5300) );
  XNOR2_X1 U6890 ( .A(n5321), .B(P2_REG3_REG_18__SCAN_IN), .ZN(n8360) );
  INV_X1 U6891 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n5304) );
  NAND2_X1 U6892 ( .A1(n5529), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n5303) );
  NAND2_X1 U6893 ( .A1(n5118), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n5302) );
  OAI211_X1 U6894 ( .C1(n5494), .C2(n5304), .A(n5303), .B(n5302), .ZN(n5305)
         );
  AOI21_X1 U6895 ( .B1(n8360), .B2(n5514), .A(n5305), .ZN(n8053) );
  OR2_X1 U6896 ( .A1(n8502), .A2(n8053), .ZN(n5687) );
  NAND2_X1 U6897 ( .A1(n8502), .A2(n8053), .ZN(n5677) );
  NAND2_X1 U6898 ( .A1(n5687), .A2(n5677), .ZN(n7830) );
  NAND2_X1 U6899 ( .A1(n5309), .A2(SI_18_), .ZN(n5348) );
  NAND2_X1 U6900 ( .A1(n5353), .A2(n5348), .ZN(n5330) );
  INV_X1 U6901 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n7208) );
  INV_X1 U6902 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n7209) );
  INV_X1 U6903 ( .A(SI_19_), .ZN(n5310) );
  NAND2_X1 U6904 ( .A1(n5311), .A2(n5310), .ZN(n5354) );
  INV_X1 U6905 ( .A(n5311), .ZN(n5312) );
  NAND2_X1 U6906 ( .A1(n5312), .A2(SI_19_), .ZN(n5349) );
  NAND2_X1 U6907 ( .A1(n5354), .A2(n5349), .ZN(n5329) );
  NAND2_X1 U6908 ( .A1(n7206), .A2(n5474), .ZN(n5317) );
  NAND2_X1 U6909 ( .A1(n5314), .A2(n5313), .ZN(n5534) );
  AOI22_X1 U6910 ( .A1(n5507), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n5315), .B2(
        n5587), .ZN(n5316) );
  INV_X1 U6911 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n5319) );
  INV_X1 U6912 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n5318) );
  OAI21_X1 U6913 ( .B1(n5321), .B2(n5319), .A(n5318), .ZN(n5322) );
  NAND2_X1 U6914 ( .A1(P2_REG3_REG_19__SCAN_IN), .A2(P2_REG3_REG_18__SCAN_IN), 
        .ZN(n5320) );
  AND2_X1 U6915 ( .A1(n5322), .A2(n5339), .ZN(n8345) );
  NAND2_X1 U6916 ( .A1(n8345), .A2(n5514), .ZN(n5328) );
  INV_X1 U6917 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n5325) );
  NAND2_X1 U6918 ( .A1(n5529), .A2(P2_REG1_REG_19__SCAN_IN), .ZN(n5324) );
  NAND2_X1 U6919 ( .A1(n5118), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n5323) );
  OAI211_X1 U6920 ( .C1(n5494), .C2(n5325), .A(n5324), .B(n5323), .ZN(n5326)
         );
  INV_X1 U6921 ( .A(n5326), .ZN(n5327) );
  NAND2_X1 U6922 ( .A1(n5328), .A2(n5327), .ZN(n8367) );
  INV_X1 U6923 ( .A(n8367), .ZN(n7983) );
  OR2_X1 U6924 ( .A1(n8498), .A2(n7983), .ZN(n5689) );
  NAND2_X1 U6925 ( .A1(n8498), .A2(n7983), .ZN(n8334) );
  OAI21_X1 U6926 ( .B1(n5330), .B2(n5329), .A(n5354), .ZN(n5335) );
  INV_X1 U6927 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n7246) );
  INV_X1 U6928 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n7268) );
  INV_X1 U6929 ( .A(SI_20_), .ZN(n5331) );
  NAND2_X1 U6930 ( .A1(n5332), .A2(n5331), .ZN(n5355) );
  INV_X1 U6931 ( .A(n5332), .ZN(n5333) );
  NAND2_X1 U6932 ( .A1(n5333), .A2(SI_20_), .ZN(n5334) );
  NAND2_X1 U6933 ( .A1(n5355), .A2(n5334), .ZN(n5351) );
  INV_X1 U6934 ( .A(n5351), .ZN(n5358) );
  NAND2_X1 U6935 ( .A1(n7245), .A2(n5474), .ZN(n5337) );
  NAND2_X1 U6936 ( .A1(n5507), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n5336) );
  INV_X1 U6937 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n5338) );
  NAND2_X1 U6938 ( .A1(n5339), .A2(n5338), .ZN(n5340) );
  NAND2_X1 U6939 ( .A1(n5364), .A2(n5340), .ZN(n8331) );
  OR2_X1 U6940 ( .A1(n8331), .A2(n4995), .ZN(n5346) );
  INV_X1 U6941 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n5343) );
  NAND2_X1 U6942 ( .A1(n5529), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n5342) );
  NAND2_X1 U6943 ( .A1(n5118), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n5341) );
  OAI211_X1 U6944 ( .C1(n5494), .C2(n5343), .A(n5342), .B(n5341), .ZN(n5344)
         );
  INV_X1 U6945 ( .A(n5344), .ZN(n5345) );
  NAND2_X1 U6946 ( .A1(n8492), .A2(n7932), .ZN(n5691) );
  NAND2_X1 U6947 ( .A1(n5690), .A2(n5691), .ZN(n8327) );
  INV_X1 U6948 ( .A(n8334), .ZN(n5686) );
  NOR2_X1 U6949 ( .A1(n8327), .A2(n5686), .ZN(n5347) );
  NAND2_X1 U6950 ( .A1(n5349), .A2(n5348), .ZN(n5350) );
  INV_X1 U6951 ( .A(n5354), .ZN(n5357) );
  INV_X1 U6952 ( .A(n5355), .ZN(n5356) );
  INV_X1 U6953 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n7211) );
  XNOR2_X1 U6954 ( .A(n5377), .B(n5373), .ZN(n7172) );
  NAND2_X1 U6955 ( .A1(n7172), .A2(n5474), .ZN(n5362) );
  NAND2_X1 U6956 ( .A1(n5507), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n5361) );
  INV_X1 U6957 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n5363) );
  OR2_X2 U6958 ( .A1(n5364), .A2(n5363), .ZN(n5385) );
  NAND2_X1 U6959 ( .A1(n5364), .A2(n5363), .ZN(n5365) );
  AND2_X1 U6960 ( .A1(n5385), .A2(n5365), .ZN(n8316) );
  NAND2_X1 U6961 ( .A1(n8316), .A2(n5514), .ZN(n5371) );
  INV_X1 U6962 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n5368) );
  NAND2_X1 U6963 ( .A1(n5118), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n5367) );
  NAND2_X1 U6964 ( .A1(n5529), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n5366) );
  OAI211_X1 U6965 ( .C1(n5368), .C2(n5494), .A(n5367), .B(n5366), .ZN(n5369)
         );
  INV_X1 U6966 ( .A(n5369), .ZN(n5370) );
  NAND2_X1 U6967 ( .A1(n5371), .A2(n5370), .ZN(n8337) );
  OR2_X1 U6968 ( .A1(n8487), .A2(n8307), .ZN(n5694) );
  NAND2_X1 U6969 ( .A1(n8487), .A2(n8307), .ZN(n8304) );
  NAND2_X1 U6970 ( .A1(n5694), .A2(n8304), .ZN(n8319) );
  NAND2_X2 U6971 ( .A1(n8321), .A2(n5372), .ZN(n8320) );
  INV_X1 U6972 ( .A(n5374), .ZN(n5375) );
  NAND2_X1 U6973 ( .A1(n5375), .A2(SI_21_), .ZN(n5376) );
  INV_X1 U6974 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n7409) );
  INV_X1 U6975 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n7407) );
  INV_X1 U6976 ( .A(SI_22_), .ZN(n5378) );
  INV_X1 U6977 ( .A(n5379), .ZN(n5380) );
  NAND2_X1 U6978 ( .A1(n5380), .A2(SI_22_), .ZN(n5381) );
  XNOR2_X1 U6979 ( .A(n5397), .B(n5396), .ZN(n7406) );
  NAND2_X1 U6980 ( .A1(n7406), .A2(n5474), .ZN(n5383) );
  NAND2_X1 U6981 ( .A1(n5507), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n5382) );
  INV_X1 U6982 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n10032) );
  NAND2_X1 U6983 ( .A1(n5385), .A2(n10032), .ZN(n5386) );
  NAND2_X1 U6984 ( .A1(n5407), .A2(n5386), .ZN(n8298) );
  OR2_X1 U6985 ( .A1(n8298), .A2(n4995), .ZN(n5392) );
  INV_X1 U6986 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n5389) );
  NAND2_X1 U6987 ( .A1(n5529), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n5388) );
  NAND2_X1 U6988 ( .A1(n5118), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n5387) );
  OAI211_X1 U6989 ( .C1(n5494), .C2(n5389), .A(n5388), .B(n5387), .ZN(n5390)
         );
  INV_X1 U6990 ( .A(n5390), .ZN(n5391) );
  NAND2_X1 U6991 ( .A1(n8482), .A2(n7916), .ZN(n5685) );
  INV_X1 U6992 ( .A(n8303), .ZN(n8294) );
  INV_X1 U6993 ( .A(n8304), .ZN(n5393) );
  NOR2_X1 U6994 ( .A1(n8294), .A2(n5393), .ZN(n5394) );
  INV_X1 U6995 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n5399) );
  INV_X1 U6996 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n5398) );
  INV_X1 U6997 ( .A(SI_23_), .ZN(n5400) );
  NAND2_X1 U6998 ( .A1(n5401), .A2(n5400), .ZN(n5417) );
  INV_X1 U6999 ( .A(n5401), .ZN(n5402) );
  NAND2_X1 U7000 ( .A1(n5402), .A2(SI_23_), .ZN(n5403) );
  XNOR2_X1 U7001 ( .A(n5416), .B(n5415), .ZN(n7342) );
  NAND2_X1 U7002 ( .A1(n7342), .A2(n5474), .ZN(n5405) );
  NAND2_X1 U7003 ( .A1(n5507), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n5404) );
  INV_X1 U7004 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n5406) );
  NAND2_X1 U7005 ( .A1(n5407), .A2(n5406), .ZN(n5408) );
  AND2_X1 U7006 ( .A1(n5422), .A2(n5408), .ZN(n8288) );
  NAND2_X1 U7007 ( .A1(n8288), .A2(n5514), .ZN(n5414) );
  INV_X1 U7008 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n5411) );
  NAND2_X1 U7009 ( .A1(n5118), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n5410) );
  NAND2_X1 U7010 ( .A1(n5529), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n5409) );
  OAI211_X1 U7011 ( .C1(n5411), .C2(n5494), .A(n5410), .B(n5409), .ZN(n5412)
         );
  INV_X1 U7012 ( .A(n5412), .ZN(n5413) );
  INV_X1 U7013 ( .A(n8282), .ZN(n5582) );
  INV_X1 U7014 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n7494) );
  INV_X1 U7015 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n7475) );
  XNOR2_X1 U7016 ( .A(n5430), .B(SI_24_), .ZN(n5429) );
  NAND2_X1 U7017 ( .A1(n7474), .A2(n5474), .ZN(n5420) );
  NAND2_X1 U7018 ( .A1(n5507), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n5419) );
  INV_X1 U7019 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n5421) );
  NAND2_X1 U7020 ( .A1(n5422), .A2(n5421), .ZN(n5423) );
  NAND2_X1 U7021 ( .A1(n5442), .A2(n5423), .ZN(n8272) );
  INV_X1 U7022 ( .A(P2_REG2_REG_24__SCAN_IN), .ZN(n8271) );
  NAND2_X1 U7023 ( .A1(n5529), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n5425) );
  NAND2_X1 U7024 ( .A1(n5118), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n5424) );
  OAI211_X1 U7025 ( .C1(n8271), .C2(n5494), .A(n5425), .B(n5424), .ZN(n5426)
         );
  INV_X1 U7026 ( .A(n5426), .ZN(n5427) );
  NAND2_X1 U7027 ( .A1(n8274), .A2(n7940), .ZN(n5701) );
  INV_X1 U7028 ( .A(n8266), .ZN(n8308) );
  AND2_X1 U7029 ( .A1(n8476), .A2(n8308), .ZN(n8262) );
  INV_X1 U7030 ( .A(n5429), .ZN(n5433) );
  INV_X1 U7031 ( .A(n5430), .ZN(n5431) );
  NAND2_X1 U7032 ( .A1(n5431), .A2(SI_24_), .ZN(n5432) );
  INV_X1 U7033 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n7637) );
  INV_X1 U7034 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n7633) );
  INV_X1 U7035 ( .A(SI_25_), .ZN(n5435) );
  NAND2_X1 U7036 ( .A1(n5436), .A2(n5435), .ZN(n5448) );
  INV_X1 U7037 ( .A(n5436), .ZN(n5437) );
  NAND2_X1 U7038 ( .A1(n5437), .A2(SI_25_), .ZN(n5438) );
  NAND2_X1 U7039 ( .A1(n5448), .A2(n5438), .ZN(n5449) );
  NAND2_X1 U7040 ( .A1(n7632), .A2(n5474), .ZN(n5440) );
  NAND2_X1 U7041 ( .A1(n5507), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n5439) );
  INV_X1 U7042 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n5441) );
  NAND2_X1 U7043 ( .A1(n5442), .A2(n5441), .ZN(n5443) );
  INV_X1 U7044 ( .A(P2_REG2_REG_25__SCAN_IN), .ZN(n5446) );
  NAND2_X1 U7045 ( .A1(n5118), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n5445) );
  NAND2_X1 U7046 ( .A1(n5529), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n5444) );
  OAI211_X1 U7047 ( .C1(n5446), .C2(n5494), .A(n5445), .B(n5444), .ZN(n5447)
         );
  NAND2_X1 U7048 ( .A1(n8466), .A2(n7974), .ZN(n5594) );
  INV_X1 U7049 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n10015) );
  INV_X1 U7050 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n7712) );
  INV_X1 U7051 ( .A(SI_26_), .ZN(n5451) );
  NAND2_X1 U7052 ( .A1(n5452), .A2(n5451), .ZN(n5468) );
  INV_X1 U7053 ( .A(n5452), .ZN(n5453) );
  NAND2_X1 U7054 ( .A1(n5453), .A2(SI_26_), .ZN(n5454) );
  NAND2_X1 U7055 ( .A1(n5507), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n5455) );
  INV_X1 U7056 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n5458) );
  NAND2_X1 U7057 ( .A1(n5459), .A2(n5458), .ZN(n5460) );
  NAND2_X1 U7058 ( .A1(n5490), .A2(n5460), .ZN(n8239) );
  INV_X1 U7059 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n9909) );
  NAND2_X1 U7060 ( .A1(n5118), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n5462) );
  NAND2_X1 U7061 ( .A1(n5529), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n5461) );
  OAI211_X1 U7062 ( .C1(n9909), .C2(n5494), .A(n5462), .B(n5461), .ZN(n5463)
         );
  INV_X1 U7063 ( .A(n5463), .ZN(n5464) );
  AND2_X2 U7064 ( .A1(n5465), .A2(n5464), .ZN(n8218) );
  NAND2_X1 U7065 ( .A1(n8462), .A2(n8218), .ZN(n5703) );
  NAND2_X2 U7066 ( .A1(n8216), .A2(n5703), .ZN(n7839) );
  INV_X1 U7067 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n7820) );
  INV_X1 U7068 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n10017) );
  INV_X1 U7069 ( .A(SI_27_), .ZN(n5470) );
  NAND2_X1 U7070 ( .A1(n5471), .A2(n5470), .ZN(n5484) );
  INV_X1 U7071 ( .A(n5471), .ZN(n5472) );
  NAND2_X1 U7072 ( .A1(n5472), .A2(SI_27_), .ZN(n5473) );
  NAND2_X1 U7073 ( .A1(n7808), .A2(n5474), .ZN(n5476) );
  NAND2_X1 U7074 ( .A1(n5507), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n5475) );
  XNOR2_X1 U7075 ( .A(n5490), .B(P2_REG3_REG_27__SCAN_IN), .ZN(n8226) );
  NAND2_X1 U7076 ( .A1(n8226), .A2(n5514), .ZN(n5481) );
  INV_X1 U7077 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n10003) );
  NAND2_X1 U7078 ( .A1(n5529), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n5478) );
  NAND2_X1 U7079 ( .A1(n5537), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n5477) );
  OAI211_X1 U7080 ( .C1(n5051), .C2(n10003), .A(n5478), .B(n5477), .ZN(n5479)
         );
  INV_X1 U7081 ( .A(n5479), .ZN(n5480) );
  OR2_X1 U7082 ( .A1(n8455), .A2(n8204), .ZN(n5710) );
  INV_X1 U7083 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n8588) );
  INV_X1 U7084 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n9990) );
  XNOR2_X1 U7085 ( .A(n5503), .B(SI_28_), .ZN(n5500) );
  NAND2_X1 U7086 ( .A1(n8586), .A2(n5474), .ZN(n5487) );
  NAND2_X1 U7087 ( .A1(n5507), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n5486) );
  INV_X1 U7088 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n5489) );
  INV_X1 U7089 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n5488) );
  OAI21_X1 U7090 ( .B1(n5490), .B2(n5489), .A(n5488), .ZN(n5491) );
  NAND2_X1 U7091 ( .A1(n8210), .A2(n5514), .ZN(n5498) );
  INV_X1 U7092 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n5495) );
  NAND2_X1 U7093 ( .A1(n5118), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n5493) );
  NAND2_X1 U7094 ( .A1(n5529), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n5492) );
  OAI211_X1 U7095 ( .C1(n5495), .C2(n5494), .A(n5493), .B(n5492), .ZN(n5496)
         );
  INV_X1 U7096 ( .A(n5496), .ZN(n5497) );
  AND2_X2 U7097 ( .A1(n5498), .A2(n5497), .ZN(n8219) );
  NAND2_X1 U7098 ( .A1(n8450), .A2(n8219), .ZN(n5499) );
  INV_X1 U7099 ( .A(n7842), .ZN(n5516) );
  INV_X1 U7100 ( .A(SI_28_), .ZN(n5502) );
  NAND2_X1 U7101 ( .A1(n5503), .A2(n5502), .ZN(n5504) );
  INV_X1 U7102 ( .A(SI_29_), .ZN(n5519) );
  XNOR2_X1 U7103 ( .A(n5521), .B(n5519), .ZN(n5506) );
  NAND2_X1 U7104 ( .A1(n8816), .A2(n5474), .ZN(n5509) );
  NAND2_X1 U7105 ( .A1(n5507), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n5508) );
  INV_X1 U7106 ( .A(n5510), .ZN(n8188) );
  INV_X1 U7107 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n9993) );
  NAND2_X1 U7108 ( .A1(n5118), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n5512) );
  NAND2_X1 U7109 ( .A1(n5537), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n5511) );
  OAI211_X1 U7110 ( .C1(n5080), .C2(n9993), .A(n5512), .B(n5511), .ZN(n5513)
         );
  NAND2_X1 U7111 ( .A1(n8189), .A2(n8203), .ZN(n5717) );
  INV_X1 U7112 ( .A(n8185), .ZN(n5515) );
  NAND2_X1 U7113 ( .A1(n5516), .A2(n5515), .ZN(n5517) );
  INV_X1 U7114 ( .A(n5520), .ZN(n5518) );
  NAND2_X1 U7115 ( .A1(n5520), .A2(n5519), .ZN(n5522) );
  NAND2_X1 U7116 ( .A1(n5522), .A2(n5521), .ZN(n5523) );
  MUX2_X1 U7117 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(P1_DATAO_REG_30__SCAN_IN), 
        .S(n6575), .Z(n5542) );
  XNOR2_X1 U7118 ( .A(n5542), .B(SI_30_), .ZN(n5525) );
  NAND2_X1 U7119 ( .A1(n8823), .A2(n5474), .ZN(n5528) );
  INV_X1 U7120 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n9963) );
  OR2_X1 U7121 ( .A1(n5526), .A2(n9963), .ZN(n5527) );
  NAND2_X1 U7122 ( .A1(n5529), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n5532) );
  NAND2_X1 U7123 ( .A1(n5537), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n5531) );
  NAND2_X1 U7124 ( .A1(n5118), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n5530) );
  AND3_X1 U7125 ( .A1(n5532), .A2(n5531), .A3(n5530), .ZN(n5551) );
  NAND2_X1 U7126 ( .A1(n5555), .A2(n5558), .ZN(n5533) );
  NOR2_X2 U7127 ( .A1(n5534), .A2(n5533), .ZN(n5553) );
  INV_X1 U7128 ( .A(n5553), .ZN(n5535) );
  INV_X1 U7129 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n9977) );
  NAND2_X1 U7130 ( .A1(n5118), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n5539) );
  NAND2_X1 U7131 ( .A1(n5537), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n5538) );
  OAI211_X1 U7132 ( .C1(n5080), .C2(n9977), .A(n5539), .B(n5538), .ZN(n8047)
         );
  INV_X1 U7133 ( .A(n8047), .ZN(n5550) );
  INV_X1 U7134 ( .A(n5542), .ZN(n5541) );
  INV_X1 U7135 ( .A(SI_30_), .ZN(n5540) );
  NOR2_X1 U7136 ( .A1(n5541), .A2(n5540), .ZN(n5543) );
  OAI22_X1 U7137 ( .A1(n5544), .A2(n5543), .B1(n5542), .B2(SI_30_), .ZN(n5548)
         );
  INV_X1 U7138 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n5545) );
  MUX2_X1 U7139 ( .A(n6693), .B(n5545), .S(n6575), .Z(n5546) );
  XNOR2_X1 U7140 ( .A(n5546), .B(SI_31_), .ZN(n5547) );
  XNOR2_X1 U7141 ( .A(n5548), .B(n5547), .ZN(n8819) );
  INV_X1 U7142 ( .A(n5551), .ZN(n8174) );
  NAND2_X1 U7143 ( .A1(n8175), .A2(n8174), .ZN(n5723) );
  NAND2_X1 U7144 ( .A1(n8444), .A2(n5550), .ZN(n5720) );
  INV_X1 U7145 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n5552) );
  NAND2_X1 U7146 ( .A1(n5553), .A2(n5552), .ZN(n5730) );
  XNOR2_X1 U7147 ( .A(n5560), .B(P2_IR_REG_22__SCAN_IN), .ZN(n5586) );
  NAND2_X1 U7148 ( .A1(n5556), .A2(n5555), .ZN(n5557) );
  XNOR2_X2 U7149 ( .A(n5559), .B(n5558), .ZN(n5568) );
  OR2_X4 U7150 ( .A1(n7116), .A2(n5588), .ZN(n5873) );
  OR2_X4 U7151 ( .A1(n5873), .A2(n5587), .ZN(n5774) );
  NAND2_X1 U7152 ( .A1(n5755), .A2(n5588), .ZN(n7028) );
  INV_X1 U7153 ( .A(n7028), .ZN(n5562) );
  INV_X1 U7154 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n5731) );
  NAND2_X1 U7155 ( .A1(n5560), .A2(n5731), .ZN(n5561) );
  NAND2_X1 U7156 ( .A1(n5561), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5743) );
  XNOR2_X1 U7157 ( .A(n5743), .B(P2_IR_REG_23__SCAN_IN), .ZN(n6540) );
  AND2_X1 U7158 ( .A1(n6540), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7343) );
  INV_X1 U7159 ( .A(n5563), .ZN(n5564) );
  NAND2_X1 U7160 ( .A1(n5565), .A2(n5564), .ZN(n5754) );
  NAND2_X1 U7161 ( .A1(n5724), .A2(n5719), .ZN(n5591) );
  INV_X1 U7162 ( .A(n8327), .ZN(n8335) );
  INV_X1 U7163 ( .A(n8373), .ZN(n8384) );
  NAND2_X1 U7164 ( .A1(n7553), .A2(n5640), .ZN(n7563) );
  NAND2_X1 U7165 ( .A1(n5635), .A2(n5634), .ZN(n7410) );
  INV_X1 U7166 ( .A(n7410), .ZN(n5632) );
  NAND2_X1 U7167 ( .A1(n7135), .A2(n7247), .ZN(n7175) );
  INV_X1 U7168 ( .A(n7175), .ZN(n7134) );
  NAND2_X1 U7169 ( .A1(n5760), .A2(n9791), .ZN(n6870) );
  NAND2_X1 U7170 ( .A1(n7165), .A2(n6870), .ZN(n9790) );
  NOR2_X1 U7171 ( .A1(n9790), .A2(n5568), .ZN(n5569) );
  NAND4_X1 U7172 ( .A1(n5570), .A2(n7134), .A3(n7079), .A4(n5569), .ZN(n5571)
         );
  NAND2_X1 U7173 ( .A1(n7213), .A2(n5625), .ZN(n7250) );
  NOR2_X1 U7174 ( .A1(n5571), .A2(n7250), .ZN(n5572) );
  NAND4_X1 U7175 ( .A1(n5138), .A2(n5632), .A3(n7225), .A4(n5572), .ZN(n5573)
         );
  NOR2_X1 U7176 ( .A1(n7563), .A2(n5573), .ZN(n5574) );
  NAND4_X1 U7177 ( .A1(n7735), .A2(n7646), .A3(n7694), .A4(n5574), .ZN(n5575)
         );
  NOR2_X1 U7178 ( .A1(n5575), .A2(n7745), .ZN(n5576) );
  NAND4_X1 U7179 ( .A1(n8384), .A2(n8434), .A3(n7743), .A4(n5576), .ZN(n5577)
         );
  NOR2_X1 U7180 ( .A1(n5577), .A2(n8398), .ZN(n5578) );
  NAND3_X1 U7181 ( .A1(n8350), .A2(n8365), .A3(n5578), .ZN(n5579) );
  NOR2_X1 U7182 ( .A1(n5579), .A2(n8319), .ZN(n5580) );
  NAND3_X1 U7183 ( .A1(n8303), .A2(n8335), .A3(n5580), .ZN(n5581) );
  NOR4_X1 U7184 ( .A1(n7837), .A2(n8261), .A3(n5582), .A4(n5581), .ZN(n5583)
         );
  NAND4_X1 U7185 ( .A1(n8199), .A2(n8235), .A3(n5583), .A4(n8223), .ZN(n5584)
         );
  XNOR2_X1 U7186 ( .A(n5585), .B(n5587), .ZN(n5589) );
  OAI22_X1 U7187 ( .A1(n5589), .A2(n5755), .B1(n5588), .B2(n7029), .ZN(n5729)
         );
  NAND2_X1 U7188 ( .A1(n5755), .A2(n5587), .ZN(n5590) );
  MUX2_X1 U7189 ( .A(n5592), .B(n5591), .S(n5722), .Z(n5727) );
  NAND2_X1 U7190 ( .A1(n8216), .A2(n5593), .ZN(n5596) );
  NAND2_X1 U7191 ( .A1(n8235), .A2(n5594), .ZN(n5595) );
  MUX2_X1 U7192 ( .A(n5596), .B(n5595), .S(n5722), .Z(n5706) );
  INV_X1 U7193 ( .A(n5597), .ZN(n5600) );
  OAI211_X1 U7194 ( .C1(n8373), .C2(n8385), .A(n5677), .B(n5598), .ZN(n5599)
         );
  MUX2_X1 U7195 ( .A(n5600), .B(n5599), .S(n5715), .Z(n5602) );
  INV_X1 U7196 ( .A(n5687), .ZN(n5601) );
  NOR2_X1 U7197 ( .A1(n5602), .A2(n5601), .ZN(n5676) );
  NAND2_X1 U7198 ( .A1(n5603), .A2(n5604), .ZN(n5605) );
  NAND2_X1 U7199 ( .A1(n5605), .A2(n5610), .ZN(n5606) );
  NAND2_X1 U7200 ( .A1(n5606), .A2(n5607), .ZN(n5613) );
  NAND3_X1 U7201 ( .A1(n5609), .A2(n5608), .A3(n5607), .ZN(n5611) );
  NAND2_X1 U7202 ( .A1(n5611), .A2(n5610), .ZN(n5612) );
  MUX2_X1 U7203 ( .A(n5613), .B(n5612), .S(n5715), .Z(n5616) );
  INV_X1 U7204 ( .A(n5626), .ZN(n5615) );
  NAND3_X1 U7205 ( .A1(n5616), .A2(n5615), .A3(n7079), .ZN(n5621) );
  AND2_X1 U7206 ( .A1(n7135), .A2(n5617), .ZN(n5618) );
  OAI211_X1 U7207 ( .C1(n5626), .C2(n5618), .A(n7213), .B(n5633), .ZN(n5619)
         );
  NAND2_X1 U7208 ( .A1(n5619), .A2(n5722), .ZN(n5620) );
  NAND2_X1 U7209 ( .A1(n5621), .A2(n5620), .ZN(n5622) );
  NAND2_X1 U7210 ( .A1(n5622), .A2(n5627), .ZN(n5631) );
  INV_X1 U7211 ( .A(n7214), .ZN(n5624) );
  AOI22_X1 U7212 ( .A1(n5626), .A2(n5625), .B1(n5624), .B2(n5623), .ZN(n5629)
         );
  INV_X1 U7213 ( .A(n5627), .ZN(n5628) );
  OAI21_X1 U7214 ( .B1(n5629), .B2(n5628), .A(n5715), .ZN(n5630) );
  MUX2_X1 U7215 ( .A(n5635), .B(n5634), .S(n5722), .Z(n5636) );
  MUX2_X1 U7216 ( .A(n7432), .B(n5637), .S(n5722), .Z(n5638) );
  AND2_X1 U7217 ( .A1(n5640), .A2(n5638), .ZN(n5639) );
  NAND2_X1 U7218 ( .A1(n5645), .A2(n5640), .ZN(n5641) );
  MUX2_X1 U7219 ( .A(n5715), .B(n5641), .S(n5644), .Z(n5649) );
  INV_X1 U7220 ( .A(n5642), .ZN(n5648) );
  NAND2_X1 U7221 ( .A1(n7724), .A2(n5642), .ZN(n5643) );
  AOI21_X1 U7222 ( .B1(n5645), .B2(n5644), .A(n5643), .ZN(n5646) );
  MUX2_X1 U7223 ( .A(n5646), .B(n5650), .S(n5722), .Z(n5647) );
  OAI21_X1 U7224 ( .B1(n5649), .B2(n5648), .A(n5647), .ZN(n5653) );
  MUX2_X1 U7225 ( .A(n5650), .B(n7724), .S(n5722), .Z(n5651) );
  AND4_X1 U7226 ( .A1(n7743), .A2(n4798), .A3(n7735), .A4(n5651), .ZN(n5652)
         );
  INV_X1 U7227 ( .A(n5659), .ZN(n5656) );
  NOR2_X1 U7228 ( .A1(n5654), .A2(n5722), .ZN(n5655) );
  AOI22_X1 U7229 ( .A1(n5656), .A2(n5715), .B1(n5658), .B2(n5655), .ZN(n5662)
         );
  OR2_X1 U7230 ( .A1(n7993), .A2(n5715), .ZN(n5657) );
  OAI22_X1 U7231 ( .A1(n5658), .A2(n5715), .B1(n8535), .B2(n5657), .ZN(n5660)
         );
  NAND2_X1 U7232 ( .A1(n5660), .A2(n5659), .ZN(n5661) );
  NAND2_X1 U7233 ( .A1(n5662), .A2(n5661), .ZN(n5663) );
  NAND2_X1 U7234 ( .A1(n5663), .A2(n4798), .ZN(n5667) );
  NAND2_X1 U7235 ( .A1(n8424), .A2(n5722), .ZN(n5665) );
  NAND2_X1 U7236 ( .A1(n8038), .A2(n5715), .ZN(n5664) );
  MUX2_X1 U7237 ( .A(n5665), .B(n5664), .S(n7751), .Z(n5666) );
  MUX2_X1 U7238 ( .A(n5669), .B(n5668), .S(n5722), .Z(n5670) );
  NAND3_X1 U7239 ( .A1(n5671), .A2(n5266), .A3(n5670), .ZN(n5672) );
  OAI21_X1 U7240 ( .B1(n5715), .B2(n5673), .A(n5672), .ZN(n5674) );
  NAND2_X1 U7241 ( .A1(n5674), .A2(n8384), .ZN(n5675) );
  NAND2_X1 U7242 ( .A1(n5688), .A2(n5677), .ZN(n5678) );
  NAND2_X1 U7243 ( .A1(n5678), .A2(n5689), .ZN(n5679) );
  NAND3_X1 U7244 ( .A1(n5679), .A2(n5691), .A3(n8334), .ZN(n5680) );
  NAND3_X1 U7245 ( .A1(n5680), .A2(n5690), .A3(n5694), .ZN(n5683) );
  AND2_X1 U7246 ( .A1(n5685), .A2(n8304), .ZN(n5682) );
  INV_X1 U7247 ( .A(n5695), .ZN(n5681) );
  AOI21_X1 U7248 ( .B1(n5683), .B2(n5682), .A(n5681), .ZN(n5684) );
  NAND2_X1 U7249 ( .A1(n5690), .A2(n5689), .ZN(n5692) );
  OAI211_X1 U7250 ( .C1(n5693), .C2(n5692), .A(n5691), .B(n8304), .ZN(n5696)
         );
  NAND2_X1 U7251 ( .A1(n8266), .A2(n5715), .ZN(n5698) );
  OR2_X1 U7252 ( .A1(n8266), .A2(n5715), .ZN(n5697) );
  MUX2_X1 U7253 ( .A(n5698), .B(n5697), .S(n8476), .Z(n5699) );
  MUX2_X1 U7254 ( .A(n5701), .B(n5700), .S(n5722), .Z(n5702) );
  MUX2_X1 U7255 ( .A(n8216), .B(n5703), .S(n5715), .Z(n5704) );
  OAI211_X1 U7256 ( .C1(n5706), .C2(n5705), .A(n8223), .B(n5704), .ZN(n5709)
         );
  AND2_X1 U7257 ( .A1(n8455), .A2(n8204), .ZN(n5707) );
  OAI21_X1 U7258 ( .B1(n8197), .B2(n5707), .A(n5722), .ZN(n5708) );
  AOI21_X1 U7259 ( .B1(n5709), .B2(n5708), .A(n4580), .ZN(n5714) );
  AOI21_X1 U7260 ( .B1(n5711), .B2(n5710), .A(n5722), .ZN(n5713) );
  NAND3_X1 U7261 ( .A1(n8450), .A2(n8219), .A3(n5715), .ZN(n5712) );
  OAI211_X1 U7262 ( .C1(n5714), .C2(n5713), .A(n5515), .B(n5712), .ZN(n5721)
         );
  MUX2_X1 U7263 ( .A(n5717), .B(n5716), .S(n5715), .Z(n5718) );
  MUX2_X1 U7264 ( .A(n5724), .B(n5723), .S(n5722), .Z(n5725) );
  OAI21_X1 U7265 ( .B1(n5727), .B2(n5726), .A(n5725), .ZN(n5728) );
  INV_X1 U7266 ( .A(n7343), .ZN(n6712) );
  INV_X1 U7267 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n5732) );
  INV_X1 U7268 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n5742) );
  NAND3_X1 U7269 ( .A1(n5732), .A2(n5731), .A3(n5742), .ZN(n5733) );
  NAND2_X1 U7270 ( .A1(n5737), .A2(n5738), .ZN(n5740) );
  NAND2_X1 U7271 ( .A1(n5740), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5734) );
  MUX2_X1 U7272 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5734), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n5736) );
  NAND2_X1 U7273 ( .A1(n5736), .A2(n5735), .ZN(n7711) );
  OR2_X1 U7274 ( .A1(n5737), .A2(n4991), .ZN(n5739) );
  MUX2_X1 U7275 ( .A(n5739), .B(P2_IR_REG_31__SCAN_IN), .S(n5738), .Z(n5741)
         );
  NAND2_X1 U7276 ( .A1(n5741), .A2(n5740), .ZN(n7635) );
  NOR2_X1 U7277 ( .A1(n7711), .A2(n7635), .ZN(n5747) );
  NAND2_X1 U7278 ( .A1(n5743), .A2(n5742), .ZN(n5744) );
  NAND2_X1 U7279 ( .A1(n5744), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5745) );
  INV_X1 U7280 ( .A(n7493), .ZN(n5746) );
  NAND2_X1 U7281 ( .A1(n5747), .A2(n5746), .ZN(n6539) );
  NOR2_X1 U7282 ( .A1(n6540), .A2(P2_U3152), .ZN(n9806) );
  NAND2_X1 U7283 ( .A1(n5568), .A2(n7207), .ZN(n5880) );
  INV_X1 U7284 ( .A(n7014), .ZN(n5750) );
  NAND2_X1 U7285 ( .A1(n4350), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5748) );
  XNOR2_X1 U7286 ( .A(n5748), .B(P2_IR_REG_28__SCAN_IN), .ZN(n6719) );
  XNOR2_X1 U7287 ( .A(n5749), .B(P2_IR_REG_27__SCAN_IN), .ZN(n7844) );
  NAND3_X1 U7288 ( .A1(n5750), .A2(n8423), .A3(n7844), .ZN(n5751) );
  OAI211_X1 U7289 ( .C1(n5752), .C2(n6712), .A(n5751), .B(P2_B_REG_SCAN_IN), 
        .ZN(n5753) );
  NAND2_X1 U7290 ( .A1(n5755), .A2(n5568), .ZN(n7020) );
  INV_X1 U7291 ( .A(n6944), .ZN(n5756) );
  AND2_X1 U7292 ( .A1(n8066), .A2(n5774), .ZN(n5762) );
  INV_X1 U7293 ( .A(n5757), .ZN(n5759) );
  INV_X1 U7294 ( .A(n5762), .ZN(n5765) );
  INV_X1 U7295 ( .A(n5763), .ZN(n5764) );
  NAND2_X1 U7296 ( .A1(n5765), .A2(n5764), .ZN(n6943) );
  INV_X1 U7297 ( .A(n5767), .ZN(n5770) );
  INV_X1 U7298 ( .A(n5768), .ZN(n5769) );
  OR2_X1 U7299 ( .A1(n7177), .A2(n6869), .ZN(n5773) );
  XNOR2_X1 U7300 ( .A(n5836), .B(n7145), .ZN(n5772) );
  NAND2_X1 U7301 ( .A1(n5773), .A2(n5772), .ZN(n6952) );
  NOR2_X1 U7302 ( .A1(n5773), .A2(n5772), .ZN(n6954) );
  AND2_X1 U7303 ( .A1(n8063), .A2(n5851), .ZN(n5776) );
  XNOR2_X1 U7304 ( .A(n7262), .B(n5850), .ZN(n5775) );
  NOR2_X1 U7305 ( .A1(n5775), .A2(n5776), .ZN(n5777) );
  AOI21_X1 U7306 ( .B1(n5776), .B2(n5775), .A(n5777), .ZN(n7093) );
  NAND2_X1 U7307 ( .A1(n7092), .A2(n7093), .ZN(n7091) );
  INV_X1 U7308 ( .A(n5777), .ZN(n5778) );
  AND2_X1 U7309 ( .A1(n8062), .A2(n5851), .ZN(n5780) );
  XNOR2_X1 U7310 ( .A(n7219), .B(n5850), .ZN(n5779) );
  NOR2_X1 U7311 ( .A1(n5779), .A2(n5780), .ZN(n5781) );
  AOI21_X1 U7312 ( .B1(n5780), .B2(n5779), .A(n5781), .ZN(n7152) );
  INV_X1 U7313 ( .A(n5781), .ZN(n5782) );
  XNOR2_X1 U7314 ( .A(n7412), .B(n5850), .ZN(n5783) );
  NOR2_X1 U7315 ( .A1(n7416), .A2(n6869), .ZN(n5784) );
  XNOR2_X1 U7316 ( .A(n5783), .B(n5784), .ZN(n7192) );
  INV_X1 U7317 ( .A(n5783), .ZN(n5786) );
  INV_X1 U7318 ( .A(n5784), .ZN(n5785) );
  XNOR2_X1 U7319 ( .A(n7429), .B(n5850), .ZN(n5788) );
  NAND2_X1 U7320 ( .A1(n8060), .A2(n5851), .ZN(n5787) );
  XNOR2_X1 U7321 ( .A(n5788), .B(n5787), .ZN(n7299) );
  INV_X1 U7322 ( .A(n5787), .ZN(n5789) );
  NOR2_X1 U7323 ( .A1(n7556), .A2(n6869), .ZN(n5791) );
  XNOR2_X1 U7324 ( .A(n8552), .B(n5850), .ZN(n5790) );
  NOR2_X1 U7325 ( .A1(n5790), .A2(n5791), .ZN(n5792) );
  AOI21_X1 U7326 ( .B1(n5791), .B2(n5790), .A(n5792), .ZN(n7447) );
  INV_X1 U7327 ( .A(n5792), .ZN(n5793) );
  XNOR2_X1 U7328 ( .A(n8546), .B(n5856), .ZN(n5794) );
  NOR2_X1 U7329 ( .A1(n7435), .A2(n6869), .ZN(n5795) );
  XNOR2_X1 U7330 ( .A(n5794), .B(n5795), .ZN(n6553) );
  NOR2_X1 U7331 ( .A1(n7627), .A2(n6869), .ZN(n5797) );
  XNOR2_X1 U7332 ( .A(n8540), .B(n5850), .ZN(n5796) );
  XOR2_X1 U7333 ( .A(n5797), .B(n5796), .Z(n6542) );
  XNOR2_X1 U7334 ( .A(n8535), .B(n5850), .ZN(n5799) );
  NOR2_X1 U7335 ( .A1(n7993), .A2(n6869), .ZN(n5798) );
  NAND2_X1 U7336 ( .A1(n5799), .A2(n5798), .ZN(n7623) );
  NOR2_X1 U7337 ( .A1(n7741), .A2(n6869), .ZN(n5801) );
  XNOR2_X1 U7338 ( .A(n8529), .B(n5850), .ZN(n5800) );
  XOR2_X1 U7339 ( .A(n5801), .B(n5800), .Z(n7988) );
  AND2_X1 U7340 ( .A1(n8424), .A2(n5851), .ZN(n5803) );
  XNOR2_X1 U7341 ( .A(n7751), .B(n5856), .ZN(n5802) );
  NOR2_X1 U7342 ( .A1(n5802), .A2(n5803), .ZN(n5804) );
  AOI21_X1 U7343 ( .B1(n5803), .B2(n5802), .A(n5804), .ZN(n7811) );
  INV_X1 U7344 ( .A(n5804), .ZN(n5805) );
  INV_X1 U7345 ( .A(n8032), .ZN(n5807) );
  XNOR2_X1 U7346 ( .A(n8433), .B(n5856), .ZN(n5806) );
  INV_X1 U7347 ( .A(n8403), .ZN(n8054) );
  NAND2_X1 U7348 ( .A1(n8054), .A2(n5851), .ZN(n8030) );
  NOR2_X1 U7349 ( .A1(n7825), .A2(n6869), .ZN(n5809) );
  XNOR2_X1 U7350 ( .A(n8512), .B(n5856), .ZN(n5808) );
  NOR2_X1 U7351 ( .A1(n5808), .A2(n5809), .ZN(n5810) );
  AOI21_X1 U7352 ( .B1(n5809), .B2(n5808), .A(n5810), .ZN(n7948) );
  INV_X1 U7353 ( .A(n5810), .ZN(n5811) );
  INV_X1 U7354 ( .A(n8405), .ZN(n8366) );
  NAND2_X1 U7355 ( .A1(n8366), .A2(n5851), .ZN(n5812) );
  XNOR2_X1 U7356 ( .A(n8509), .B(n5856), .ZN(n5814) );
  XOR2_X1 U7357 ( .A(n5812), .B(n5814), .Z(n7957) );
  INV_X1 U7358 ( .A(n5812), .ZN(n5813) );
  NAND2_X1 U7359 ( .A1(n5814), .A2(n5813), .ZN(n5815) );
  XNOR2_X1 U7360 ( .A(n8362), .B(n5856), .ZN(n5816) );
  NOR2_X1 U7361 ( .A1(n8053), .A2(n6869), .ZN(n5818) );
  XNOR2_X1 U7362 ( .A(n5816), .B(n5818), .ZN(n8011) );
  INV_X1 U7363 ( .A(n5816), .ZN(n5817) );
  AND2_X1 U7364 ( .A1(n8367), .A2(n5851), .ZN(n5820) );
  XNOR2_X1 U7365 ( .A(n8498), .B(n5856), .ZN(n5819) );
  NOR2_X1 U7366 ( .A1(n5819), .A2(n5820), .ZN(n5821) );
  AOI21_X1 U7367 ( .B1(n5820), .B2(n5819), .A(n5821), .ZN(n7921) );
  INV_X1 U7368 ( .A(n5821), .ZN(n5822) );
  XNOR2_X1 U7369 ( .A(n8492), .B(n5856), .ZN(n5825) );
  NAND2_X1 U7370 ( .A1(n8351), .A2(n5851), .ZN(n5823) );
  INV_X1 U7371 ( .A(n5823), .ZN(n5824) );
  NAND2_X1 U7372 ( .A1(n5825), .A2(n5824), .ZN(n5826) );
  XNOR2_X1 U7373 ( .A(n8487), .B(n5856), .ZN(n5830) );
  NAND2_X1 U7374 ( .A1(n8337), .A2(n5851), .ZN(n5831) );
  XNOR2_X1 U7375 ( .A(n5830), .B(n5831), .ZN(n7929) );
  XNOR2_X1 U7376 ( .A(n8482), .B(n5856), .ZN(n8003) );
  NOR2_X1 U7377 ( .A1(n7916), .A2(n6869), .ZN(n5829) );
  INV_X1 U7378 ( .A(n5831), .ZN(n5828) );
  NAND2_X1 U7379 ( .A1(n5830), .A2(n5828), .ZN(n8000) );
  INV_X1 U7380 ( .A(n5829), .ZN(n8002) );
  NAND2_X1 U7381 ( .A1(n8000), .A2(n8002), .ZN(n5834) );
  INV_X1 U7382 ( .A(n5830), .ZN(n5832) );
  NOR3_X1 U7383 ( .A1(n5832), .A2(n7916), .A3(n5831), .ZN(n5833) );
  AOI21_X1 U7384 ( .B1(n8003), .B2(n5834), .A(n5833), .ZN(n5835) );
  XNOR2_X1 U7385 ( .A(n8476), .B(n5836), .ZN(n5839) );
  XNOR2_X2 U7386 ( .A(n5841), .B(n5839), .ZN(n7969) );
  XNOR2_X1 U7387 ( .A(n8274), .B(n5850), .ZN(n7971) );
  INV_X1 U7388 ( .A(n7940), .ZN(n8280) );
  AND2_X1 U7389 ( .A1(n8266), .A2(n5851), .ZN(n7968) );
  OAI21_X1 U7390 ( .B1(n7971), .B2(n8280), .A(n7968), .ZN(n5837) );
  INV_X1 U7391 ( .A(n5837), .ZN(n5838) );
  NAND2_X1 U7392 ( .A1(n7969), .A2(n5838), .ZN(n5846) );
  INV_X1 U7393 ( .A(n5839), .ZN(n5840) );
  NOR2_X1 U7394 ( .A1(n7940), .A2(n6869), .ZN(n7970) );
  NOR2_X1 U7395 ( .A1(n7971), .A2(n7970), .ZN(n5843) );
  NAND2_X1 U7396 ( .A1(n7971), .A2(n7970), .ZN(n5842) );
  OAI21_X1 U7397 ( .B1(n7966), .B2(n5843), .A(n5842), .ZN(n5844) );
  INV_X1 U7398 ( .A(n5844), .ZN(n5845) );
  XNOR2_X1 U7399 ( .A(n8466), .B(n5856), .ZN(n7936) );
  NOR2_X1 U7400 ( .A1(n7974), .A2(n6869), .ZN(n7937) );
  XNOR2_X1 U7401 ( .A(n8462), .B(n5856), .ZN(n5848) );
  NOR2_X1 U7402 ( .A1(n8218), .A2(n6869), .ZN(n5847) );
  NAND2_X1 U7403 ( .A1(n5848), .A2(n5847), .ZN(n5849) );
  OAI21_X1 U7404 ( .B1(n5848), .B2(n5847), .A(n5849), .ZN(n8020) );
  NAND2_X1 U7405 ( .A1(n8021), .A2(n5849), .ZN(n5901) );
  XNOR2_X1 U7406 ( .A(n8455), .B(n5850), .ZN(n5853) );
  INV_X1 U7407 ( .A(n5853), .ZN(n5855) );
  AND2_X1 U7408 ( .A1(n8050), .A2(n5851), .ZN(n5852) );
  INV_X1 U7409 ( .A(n5852), .ZN(n5854) );
  AOI21_X1 U7410 ( .B1(n5855), .B2(n5854), .A(n5887), .ZN(n5902) );
  NAND2_X1 U7411 ( .A1(n5901), .A2(n5902), .ZN(n5906) );
  NOR2_X1 U7412 ( .A1(n8219), .A2(n6869), .ZN(n5857) );
  XNOR2_X1 U7413 ( .A(n5857), .B(n5856), .ZN(n5890) );
  INV_X1 U7414 ( .A(n5890), .ZN(n5879) );
  INV_X1 U7415 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n9805) );
  INV_X1 U7416 ( .A(n7711), .ZN(n5860) );
  XNOR2_X1 U7417 ( .A(n7493), .B(P2_B_REG_SCAN_IN), .ZN(n5858) );
  NAND2_X1 U7418 ( .A1(n7635), .A2(n5858), .ZN(n5859) );
  AND2_X1 U7419 ( .A1(n7711), .A2(n7635), .ZN(n9807) );
  AOI21_X1 U7420 ( .B1(n9805), .B2(n9800), .A(n9807), .ZN(n7114) );
  NOR4_X1 U7421 ( .A1(P2_D_REG_28__SCAN_IN), .A2(P2_D_REG_2__SCAN_IN), .A3(
        P2_D_REG_3__SCAN_IN), .A4(P2_D_REG_4__SCAN_IN), .ZN(n5869) );
  OR4_X1 U7422 ( .A1(P2_D_REG_10__SCAN_IN), .A2(P2_D_REG_14__SCAN_IN), .A3(
        P2_D_REG_19__SCAN_IN), .A4(P2_D_REG_29__SCAN_IN), .ZN(n5866) );
  NOR4_X1 U7423 ( .A1(P2_D_REG_15__SCAN_IN), .A2(P2_D_REG_16__SCAN_IN), .A3(
        P2_D_REG_17__SCAN_IN), .A4(P2_D_REG_18__SCAN_IN), .ZN(n5864) );
  NOR4_X1 U7424 ( .A1(P2_D_REG_12__SCAN_IN), .A2(P2_D_REG_9__SCAN_IN), .A3(
        P2_D_REG_11__SCAN_IN), .A4(P2_D_REG_13__SCAN_IN), .ZN(n5863) );
  NOR4_X1 U7425 ( .A1(P2_D_REG_24__SCAN_IN), .A2(P2_D_REG_25__SCAN_IN), .A3(
        P2_D_REG_26__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n5862) );
  NOR4_X1 U7426 ( .A1(P2_D_REG_20__SCAN_IN), .A2(P2_D_REG_21__SCAN_IN), .A3(
        P2_D_REG_22__SCAN_IN), .A4(P2_D_REG_23__SCAN_IN), .ZN(n5861) );
  NAND4_X1 U7427 ( .A1(n5864), .A2(n5863), .A3(n5862), .A4(n5861), .ZN(n5865)
         );
  NOR4_X1 U7428 ( .A1(P2_D_REG_27__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        n5866), .A4(n5865), .ZN(n5868) );
  NOR4_X1 U7429 ( .A1(P2_D_REG_5__SCAN_IN), .A2(P2_D_REG_6__SCAN_IN), .A3(
        P2_D_REG_7__SCAN_IN), .A4(P2_D_REG_8__SCAN_IN), .ZN(n5867) );
  NAND3_X1 U7430 ( .A1(n5869), .A2(n5868), .A3(n5867), .ZN(n5870) );
  NAND2_X1 U7431 ( .A1(n5870), .A2(n9800), .ZN(n7112) );
  AND2_X1 U7432 ( .A1(n7114), .A2(n7112), .ZN(n7035) );
  INV_X1 U7433 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n9803) );
  NAND2_X1 U7434 ( .A1(n9800), .A2(n9803), .ZN(n5872) );
  AND2_X1 U7435 ( .A1(n7493), .A2(n7711), .ZN(n9804) );
  INV_X1 U7436 ( .A(n9804), .ZN(n5871) );
  NAND2_X1 U7437 ( .A1(n7035), .A2(n7853), .ZN(n5884) );
  NAND2_X1 U7438 ( .A1(n5884), .A2(n7111), .ZN(n5883) );
  OR2_X1 U7439 ( .A1(n7116), .A2(n5568), .ZN(n7025) );
  OAI21_X1 U7440 ( .B1(n9801), .B2(n7025), .A(n8411), .ZN(n5874) );
  NAND2_X1 U7441 ( .A1(n8450), .A2(n8029), .ZN(n5891) );
  OR2_X1 U7442 ( .A1(n5891), .A2(n5890), .ZN(n5878) );
  NAND2_X1 U7443 ( .A1(n8450), .A2(n8041), .ZN(n5877) );
  OR2_X1 U7444 ( .A1(n7116), .A2(n7207), .ZN(n5875) );
  OR2_X1 U7445 ( .A1(n7015), .A2(n8553), .ZN(n5876) );
  NAND2_X1 U7446 ( .A1(n5877), .A2(n8019), .ZN(n5893) );
  OAI211_X1 U7447 ( .C1(n8450), .C2(n5879), .A(n5878), .B(n5893), .ZN(n5900)
         );
  AOI21_X1 U7448 ( .B1(n5885), .B2(n5880), .A(n6540), .ZN(n5881) );
  AND2_X1 U7449 ( .A1(n6539), .A2(n5881), .ZN(n5882) );
  NAND2_X1 U7450 ( .A1(n5883), .A2(n5882), .ZN(n6867) );
  INV_X1 U7451 ( .A(n8203), .ZN(n8048) );
  INV_X1 U7452 ( .A(n5885), .ZN(n7019) );
  NOR2_X2 U7453 ( .A1(n8024), .A2(n8404), .ZN(n8035) );
  AOI22_X1 U7454 ( .A1(n8048), .A2(n8035), .B1(P2_REG3_REG_28__SCAN_IN), .B2(
        P2_U3152), .ZN(n5886) );
  OAI21_X1 U7455 ( .B1(n8204), .B2(n8039), .A(n5886), .ZN(n5889) );
  INV_X1 U7456 ( .A(n5887), .ZN(n5894) );
  NOR2_X1 U7457 ( .A1(n5900), .A2(n5894), .ZN(n5888) );
  AOI211_X1 U7458 ( .C1(n8210), .C2(n8042), .A(n5889), .B(n5888), .ZN(n5899)
         );
  MUX2_X1 U7459 ( .A(n8450), .B(n5891), .S(n5890), .Z(n5892) );
  INV_X1 U7460 ( .A(n5892), .ZN(n5896) );
  NAND2_X1 U7461 ( .A1(n5906), .A2(n5897), .ZN(n5898) );
  OAI211_X1 U7462 ( .C1(n5906), .C2(n5900), .A(n5899), .B(n5898), .ZN(P2_U3222) );
  INV_X1 U7463 ( .A(n5901), .ZN(n5904) );
  INV_X1 U7464 ( .A(n5902), .ZN(n5903) );
  NAND3_X1 U7465 ( .A1(n5906), .A2(n8033), .A3(n5905), .ZN(n5912) );
  AOI22_X1 U7466 ( .A1(n8049), .A2(n8035), .B1(P2_REG3_REG_27__SCAN_IN), .B2(
        P2_U3152), .ZN(n5907) );
  OAI21_X1 U7467 ( .B1(n8218), .B2(n8039), .A(n5907), .ZN(n5908) );
  AOI21_X1 U7468 ( .B1(n8226), .B2(n8042), .A(n5908), .ZN(n5909) );
  INV_X1 U7469 ( .A(n5910), .ZN(n5911) );
  NAND2_X1 U7470 ( .A1(n5912), .A2(n5911), .ZN(P2_U3216) );
  NOR2_X2 U7472 ( .A1(P1_IR_REG_15__SCAN_IN), .A2(P1_IR_REG_14__SCAN_IN), .ZN(
        n6259) );
  NAND2_X1 U7473 ( .A1(n5935), .A2(n5921), .ZN(n6277) );
  NAND2_X1 U7474 ( .A1(n5926), .A2(n6473), .ZN(n5923) );
  OR2_X1 U7475 ( .A1(n5924), .A2(n6472), .ZN(n5925) );
  INV_X1 U7476 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n5927) );
  NOR2_X1 U7477 ( .A1(P1_IR_REG_18__SCAN_IN), .A2(P1_IR_REG_17__SCAN_IN), .ZN(
        n5930) );
  NOR2_X1 U7478 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(P1_IR_REG_23__SCAN_IN), .ZN(
        n5929) );
  AND4_X2 U7479 ( .A1(n5930), .A2(n5929), .A3(n5928), .A4(n6472), .ZN(n5945)
         );
  NAND4_X1 U7480 ( .A1(n5932), .A2(n5945), .A3(n5931), .A4(n6098), .ZN(n5968)
         );
  NAND2_X1 U7481 ( .A1(n5968), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6516) );
  INV_X1 U7482 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n5933) );
  NAND2_X1 U7483 ( .A1(n6516), .A2(n5933), .ZN(n5939) );
  NAND2_X1 U7484 ( .A1(n5939), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5934) );
  XNOR2_X1 U7485 ( .A(n5934), .B(P1_IR_REG_26__SCAN_IN), .ZN(n6468) );
  NAND2_X1 U7486 ( .A1(n5935), .A2(n5945), .ZN(n5936) );
  NAND2_X1 U7487 ( .A1(n5936), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5937) );
  XNOR2_X1 U7488 ( .A(n5937), .B(P1_IR_REG_24__SCAN_IN), .ZN(n6469) );
  INV_X1 U7489 ( .A(n6516), .ZN(n5938) );
  NAND2_X1 U7490 ( .A1(n5938), .A2(P1_IR_REG_25__SCAN_IN), .ZN(n5940) );
  NAND3_X1 U7491 ( .A1(n6468), .A2(n6469), .A3(n6464), .ZN(n6506) );
  NAND2_X1 U7492 ( .A1(n5975), .A2(n9091), .ZN(n6479) );
  NAND2_X1 U7493 ( .A1(n6476), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5944) );
  INV_X1 U7494 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n6474) );
  NOR2_X1 U7495 ( .A1(n6479), .A2(n6522), .ZN(n7323) );
  NOR2_X1 U7496 ( .A1(P1_IR_REG_28__SCAN_IN), .A2(P1_IR_REG_27__SCAN_IN), .ZN(
        n5961) );
  NAND2_X4 U7497 ( .A1(n7856), .A2(n9570), .ZN(n6584) );
  INV_X1 U7498 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n5947) );
  INV_X1 U7499 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n5949) );
  OR2_X1 U7500 ( .A1(n4264), .A2(n5949), .ZN(n5954) );
  INV_X1 U7501 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n5950) );
  OR2_X1 U7502 ( .A1(n6051), .A2(n5950), .ZN(n5953) );
  INV_X1 U7503 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n6637) );
  NAND4_X4 U7504 ( .A1(n5955), .A2(n5954), .A3(n5953), .A4(n5952), .ZN(n7106)
         );
  INV_X1 U7505 ( .A(n7106), .ZN(n9704) );
  INV_X1 U7506 ( .A(n6506), .ZN(n6541) );
  INV_X1 U7507 ( .A(SI_0_), .ZN(n5957) );
  INV_X1 U7508 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n5956) );
  OAI21_X1 U7509 ( .B1(n6575), .B2(n5957), .A(n5956), .ZN(n5959) );
  AND2_X1 U7510 ( .A1(n5959), .A2(n5958), .ZN(n9577) );
  NAND2_X1 U7511 ( .A1(n6513), .A2(P1_IR_REG_28__SCAN_IN), .ZN(n5960) );
  INV_X1 U7512 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n5963) );
  NAND2_X1 U7513 ( .A1(n5963), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5965) );
  INV_X1 U7514 ( .A(n5965), .ZN(n5967) );
  NAND2_X1 U7515 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_27__SCAN_IN), 
        .ZN(n6517) );
  INV_X1 U7516 ( .A(n5961), .ZN(n5962) );
  OAI21_X1 U7517 ( .B1(n6517), .B2(n5963), .A(n5962), .ZN(n5964) );
  OAI21_X1 U7518 ( .B1(n6513), .B2(n5965), .A(n5964), .ZN(n5966) );
  AOI22_X1 U7519 ( .A1(n4260), .A2(n7458), .B1(n6541), .B2(
        P1_IR_REG_0__SCAN_IN), .ZN(n5971) );
  NOR2_X1 U7520 ( .A1(n6506), .A2(n6637), .ZN(n5972) );
  AOI21_X1 U7521 ( .B1(n6499), .B2(n7458), .A(n5972), .ZN(n5974) );
  NAND2_X1 U7522 ( .A1(n4260), .A2(n7106), .ZN(n5973) );
  NAND2_X1 U7523 ( .A1(n5974), .A2(n5973), .ZN(n6969) );
  NAND2_X2 U7524 ( .A1(n9710), .A2(n7478), .ZN(n7322) );
  INV_X1 U7525 ( .A(n6969), .ZN(n5976) );
  NAND2_X1 U7526 ( .A1(n7322), .A2(n5976), .ZN(n5977) );
  NAND2_X1 U7527 ( .A1(n6968), .A2(n5977), .ZN(n5990) );
  INV_X1 U7528 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n5978) );
  INV_X1 U7529 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n9698) );
  INV_X1 U7530 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n5979) );
  OR2_X1 U7531 ( .A1(n6055), .A2(n5979), .ZN(n5981) );
  INV_X2 U7532 ( .A(n6640), .ZN(n6620) );
  NAND2_X1 U7533 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5984) );
  AOI22_X1 U7534 ( .A1(n6003), .A2(P2_DATAO_REG_1__SCAN_IN), .B1(n4265), .B2(
        n6659), .ZN(n5986) );
  AND2_X2 U7535 ( .A1(n5986), .A2(n5985), .ZN(n9724) );
  INV_X1 U7536 ( .A(n9724), .ZN(n9692) );
  AOI22_X1 U7537 ( .A1(n4260), .A2(n6890), .B1(n6499), .B2(n9692), .ZN(n5987)
         );
  XNOR2_X1 U7538 ( .A(n7322), .B(n5987), .ZN(n5991) );
  NAND2_X1 U7539 ( .A1(n5990), .A2(n5991), .ZN(n7103) );
  INV_X1 U7540 ( .A(n6890), .ZN(n8770) );
  OR2_X1 U7541 ( .A1(n6397), .A2(n8770), .ZN(n5989) );
  NAND2_X1 U7542 ( .A1(n4260), .A2(n9692), .ZN(n5988) );
  NAND2_X1 U7543 ( .A1(n5989), .A2(n5988), .ZN(n7105) );
  INV_X1 U7544 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n5994) );
  OR2_X1 U7545 ( .A1(n6584), .A2(n5994), .ZN(n5998) );
  INV_X1 U7546 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n9122) );
  INV_X1 U7547 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n6662) );
  OR2_X1 U7548 ( .A1(n6055), .A2(n6662), .ZN(n5996) );
  NAND2_X1 U7549 ( .A1(n6069), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n5995) );
  NAND2_X1 U7550 ( .A1(n6560), .A2(n6274), .ZN(n6006) );
  INV_X1 U7551 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n6978) );
  INV_X1 U7552 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n5999) );
  NAND2_X1 U7553 ( .A1(n6978), .A2(n5999), .ZN(n6037) );
  INV_X1 U7554 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n6000) );
  OR2_X1 U7555 ( .A1(n6001), .A2(n6000), .ZN(n6002) );
  NAND2_X1 U7556 ( .A1(n6620), .A2(n9124), .ZN(n6005) );
  NAND2_X1 U7557 ( .A1(n6003), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n6004) );
  INV_X1 U7558 ( .A(n6894), .ZN(n8774) );
  AOI22_X1 U7559 ( .A1(n4260), .A2(n6893), .B1(n6499), .B2(n8774), .ZN(n6007)
         );
  XNOR2_X1 U7560 ( .A(n7322), .B(n6007), .ZN(n6011) );
  INV_X1 U7561 ( .A(n6893), .ZN(n9701) );
  OR2_X1 U7562 ( .A1(n6397), .A2(n9701), .ZN(n6009) );
  NAND2_X1 U7563 ( .A1(n4260), .A2(n8774), .ZN(n6008) );
  NAND2_X1 U7564 ( .A1(n6009), .A2(n6008), .ZN(n6010) );
  XNOR2_X1 U7565 ( .A(n6011), .B(n6010), .ZN(n8768) );
  INV_X1 U7566 ( .A(n6010), .ZN(n6012) );
  NAND2_X1 U7567 ( .A1(n6012), .A2(n6011), .ZN(n6013) );
  NAND2_X1 U7568 ( .A1(n6069), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n6018) );
  OR2_X1 U7569 ( .A1(n4264), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n6017) );
  INV_X1 U7570 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n6014) );
  OR2_X1 U7571 ( .A1(n6584), .A2(n6014), .ZN(n6016) );
  INV_X1 U7572 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n6664) );
  OR2_X1 U7573 ( .A1(n6055), .A2(n6664), .ZN(n6015) );
  NAND2_X1 U7574 ( .A1(n6565), .A2(n6274), .ZN(n6021) );
  AOI22_X1 U7575 ( .A1(n6003), .A2(P2_DATAO_REG_3__SCAN_IN), .B1(n6620), .B2(
        n6665), .ZN(n6020) );
  AND2_X1 U7576 ( .A1(n6021), .A2(n6020), .ZN(n7351) );
  INV_X1 U7577 ( .A(n7351), .ZN(n9729) );
  AOI22_X1 U7578 ( .A1(n4260), .A2(n9116), .B1(n6499), .B2(n9729), .ZN(n6022)
         );
  XNOR2_X1 U7579 ( .A(n7322), .B(n6022), .ZN(n6026) );
  INV_X1 U7580 ( .A(n9116), .ZN(n9677) );
  OR2_X1 U7581 ( .A1(n6397), .A2(n9677), .ZN(n6024) );
  NAND2_X1 U7582 ( .A1(n4260), .A2(n9729), .ZN(n6023) );
  NAND2_X1 U7583 ( .A1(n6024), .A2(n6023), .ZN(n6025) );
  XNOR2_X1 U7584 ( .A(n6026), .B(n6025), .ZN(n7199) );
  INV_X1 U7585 ( .A(n6025), .ZN(n6027) );
  NAND2_X1 U7586 ( .A1(n6027), .A2(n6026), .ZN(n6028) );
  NAND2_X1 U7587 ( .A1(n6087), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n6036) );
  INV_X1 U7588 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n6667) );
  OR2_X1 U7589 ( .A1(n6116), .A2(n6667), .ZN(n6035) );
  INV_X1 U7590 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n6652) );
  OR2_X1 U7591 ( .A1(n6051), .A2(n6652), .ZN(n6034) );
  INV_X1 U7592 ( .A(n6052), .ZN(n6032) );
  INV_X1 U7593 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n6030) );
  INV_X1 U7594 ( .A(P1_REG3_REG_4__SCAN_IN), .ZN(n6029) );
  NAND2_X1 U7595 ( .A1(n6030), .A2(n6029), .ZN(n6031) );
  NAND2_X1 U7596 ( .A1(n6032), .A2(n6031), .ZN(n9681) );
  OR2_X1 U7597 ( .A1(n4264), .A2(n9681), .ZN(n6033) );
  AND4_X2 U7598 ( .A1(n6036), .A2(n6035), .A3(n6034), .A4(n6033), .ZN(n7354)
         );
  NAND2_X1 U7599 ( .A1(n6563), .A2(n6274), .ZN(n6044) );
  INV_X1 U7600 ( .A(n6037), .ZN(n6039) );
  NOR2_X1 U7601 ( .A1(P1_IR_REG_2__SCAN_IN), .A2(P1_IR_REG_3__SCAN_IN), .ZN(
        n6038) );
  NAND2_X1 U7602 ( .A1(n6039), .A2(n6038), .ZN(n6041) );
  NAND2_X1 U7603 ( .A1(n6041), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6040) );
  MUX2_X1 U7604 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6040), .S(
        P1_IR_REG_4__SCAN_IN), .Z(n6042) );
  AOI22_X1 U7605 ( .A1(n6003), .A2(P2_DATAO_REG_4__SCAN_IN), .B1(n6620), .B2(
        n6658), .ZN(n6043) );
  INV_X1 U7606 ( .A(n9735), .ZN(n9682) );
  OAI22_X1 U7607 ( .A1(n4282), .A2(n7354), .B1(n9682), .B2(n6045), .ZN(n6046)
         );
  XNOR2_X1 U7608 ( .A(n7322), .B(n6046), .ZN(n6050) );
  OR2_X1 U7609 ( .A1(n6397), .A2(n7354), .ZN(n6048) );
  NAND2_X1 U7610 ( .A1(n4260), .A2(n9735), .ZN(n6047) );
  NAND2_X1 U7611 ( .A1(n6048), .A2(n6047), .ZN(n6049) );
  XNOR2_X1 U7612 ( .A(n6050), .B(n6049), .ZN(n7400) );
  NAND2_X1 U7613 ( .A1(n6050), .A2(n6049), .ZN(n7307) );
  NAND2_X1 U7614 ( .A1(n6087), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n6059) );
  INV_X1 U7615 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n6654) );
  OR2_X1 U7616 ( .A1(n6051), .A2(n6654), .ZN(n6058) );
  OAI21_X1 U7617 ( .B1(n6052), .B2(P1_REG3_REG_5__SCAN_IN), .A(n6090), .ZN(
        n7603) );
  OR2_X1 U7618 ( .A1(n4264), .A2(n7603), .ZN(n6057) );
  INV_X1 U7619 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n6054) );
  OR2_X1 U7620 ( .A1(n6055), .A2(n6054), .ZN(n6056) );
  NAND2_X1 U7621 ( .A1(n6574), .A2(n6274), .ZN(n6063) );
  NAND2_X1 U7622 ( .A1(n6060), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6061) );
  XNOR2_X1 U7623 ( .A(n6061), .B(P1_IR_REG_5__SCAN_IN), .ZN(n9134) );
  AOI22_X1 U7624 ( .A1(n6003), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n6620), .B2(
        n9134), .ZN(n6062) );
  NAND2_X1 U7625 ( .A1(n6499), .A2(n7602), .ZN(n6064) );
  OAI21_X1 U7626 ( .B1(n4282), .B2(n9676), .A(n6064), .ZN(n6065) );
  XNOR2_X1 U7627 ( .A(n7322), .B(n6065), .ZN(n7308) );
  OR2_X1 U7628 ( .A1(n6397), .A2(n9676), .ZN(n6067) );
  NAND2_X1 U7629 ( .A1(n4260), .A2(n7602), .ZN(n6066) );
  NAND2_X1 U7630 ( .A1(n6067), .A2(n6066), .ZN(n7309) );
  NAND2_X1 U7631 ( .A1(n7308), .A2(n7309), .ZN(n6068) );
  NAND2_X1 U7632 ( .A1(n6582), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n6075) );
  INV_X1 U7633 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n6070) );
  OR2_X1 U7634 ( .A1(n6584), .A2(n6070), .ZN(n6074) );
  INV_X1 U7635 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n6071) );
  XNOR2_X1 U7636 ( .A(n6090), .B(n6071), .ZN(n7390) );
  OR2_X1 U7637 ( .A1(n4264), .A2(n7390), .ZN(n6073) );
  INV_X1 U7638 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n6669) );
  OR2_X1 U7639 ( .A1(n6116), .A2(n6669), .ZN(n6072) );
  OR2_X1 U7640 ( .A1(n6397), .A2(n7357), .ZN(n6080) );
  NAND2_X1 U7641 ( .A1(n6579), .A2(n6274), .ZN(n6078) );
  OR2_X1 U7642 ( .A1(n6098), .A2(n6275), .ZN(n6076) );
  XNOR2_X1 U7643 ( .A(n6076), .B(P1_IR_REG_6__SCAN_IN), .ZN(n6670) );
  AOI22_X1 U7644 ( .A1(n6003), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n6620), .B2(
        n6670), .ZN(n6077) );
  NAND2_X1 U7645 ( .A1(n7358), .A2(n4260), .ZN(n6079) );
  NAND2_X1 U7646 ( .A1(n6080), .A2(n6079), .ZN(n6083) );
  INV_X1 U7647 ( .A(n7357), .ZN(n9113) );
  AOI22_X1 U7648 ( .A1(n7358), .A2(n6499), .B1(n4260), .B2(n9113), .ZN(n6082)
         );
  INV_X2 U7649 ( .A(n7322), .ZN(n6081) );
  XOR2_X1 U7650 ( .A(n6082), .B(n6497), .Z(n7333) );
  INV_X1 U7651 ( .A(n6083), .ZN(n7332) );
  NAND2_X1 U7652 ( .A1(n6087), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n6095) );
  INV_X1 U7653 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n7377) );
  OR2_X1 U7654 ( .A1(n6051), .A2(n7377), .ZN(n6094) );
  INV_X1 U7655 ( .A(n6090), .ZN(n6088) );
  AOI21_X1 U7656 ( .B1(n6088), .B2(P1_REG3_REG_6__SCAN_IN), .A(
        P1_REG3_REG_7__SCAN_IN), .ZN(n6091) );
  OR2_X1 U7657 ( .A1(n6091), .A2(n6117), .ZN(n7500) );
  OR2_X1 U7658 ( .A1(n4264), .A2(n7500), .ZN(n6093) );
  INV_X1 U7659 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n6672) );
  OR2_X1 U7660 ( .A1(n6116), .A2(n6672), .ZN(n6092) );
  OR2_X1 U7661 ( .A1(n6397), .A2(n7615), .ZN(n6103) );
  NAND2_X1 U7662 ( .A1(n6096), .A2(n6274), .ZN(n6101) );
  INV_X1 U7663 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n6097) );
  NAND2_X1 U7664 ( .A1(n6098), .A2(n6097), .ZN(n6108) );
  NAND2_X1 U7665 ( .A1(n6108), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6099) );
  XNOR2_X1 U7666 ( .A(n6099), .B(P1_IR_REG_7__SCAN_IN), .ZN(n6671) );
  AOI22_X1 U7667 ( .A1(n6003), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n6620), .B2(
        n6671), .ZN(n6100) );
  NAND2_X1 U7668 ( .A1(n7363), .A2(n4260), .ZN(n6102) );
  NAND2_X1 U7669 ( .A1(n6103), .A2(n6102), .ZN(n6105) );
  INV_X1 U7670 ( .A(n7363), .ZN(n9762) );
  OAI22_X1 U7671 ( .A1(n9762), .A2(n6045), .B1(n7615), .B2(n4282), .ZN(n6104)
         );
  XNOR2_X1 U7672 ( .A(n6104), .B(n6497), .ZN(n6106) );
  XOR2_X1 U7673 ( .A(n6105), .B(n6106), .Z(n7495) );
  NAND2_X1 U7674 ( .A1(n6600), .A2(n6274), .ZN(n6115) );
  NAND2_X1 U7675 ( .A1(n6110), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6109) );
  MUX2_X1 U7676 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6109), .S(
        P1_IR_REG_8__SCAN_IN), .Z(n6113) );
  INV_X1 U7677 ( .A(n6110), .ZN(n6112) );
  INV_X1 U7678 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n6111) );
  NAND2_X1 U7679 ( .A1(n6112), .A2(n6111), .ZN(n6144) );
  NAND2_X1 U7680 ( .A1(n6113), .A2(n6144), .ZN(n6701) );
  INV_X1 U7681 ( .A(n6701), .ZN(n6678) );
  AOI22_X1 U7682 ( .A1(n6620), .A2(n6678), .B1(n8824), .B2(
        P2_DATAO_REG_8__SCAN_IN), .ZN(n6114) );
  NAND2_X1 U7683 ( .A1(n7620), .A2(n4260), .ZN(n6124) );
  NAND2_X1 U7684 ( .A1(n6087), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n6122) );
  INV_X1 U7685 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n6695) );
  OR2_X1 U7686 ( .A1(n6116), .A2(n6695), .ZN(n6121) );
  INV_X1 U7687 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n7589) );
  OR2_X1 U7688 ( .A1(n6051), .A2(n7589), .ZN(n6120) );
  OR2_X1 U7689 ( .A1(n6117), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n6118) );
  NAND2_X1 U7690 ( .A1(n6152), .A2(n6118), .ZN(n7618) );
  OR2_X1 U7691 ( .A1(n4264), .A2(n7618), .ZN(n6119) );
  OR2_X1 U7692 ( .A1(n6397), .A2(n8714), .ZN(n6123) );
  NAND2_X1 U7693 ( .A1(n6124), .A2(n6123), .ZN(n8613) );
  NAND2_X1 U7694 ( .A1(n7620), .A2(n6499), .ZN(n6126) );
  INV_X1 U7695 ( .A(n8714), .ZN(n9111) );
  NAND2_X1 U7696 ( .A1(n4260), .A2(n9111), .ZN(n6125) );
  NAND2_X1 U7697 ( .A1(n6126), .A2(n6125), .ZN(n6127) );
  XNOR2_X1 U7698 ( .A(n6127), .B(n6497), .ZN(n8612) );
  NAND2_X1 U7699 ( .A1(n6604), .A2(n8822), .ZN(n6130) );
  NAND2_X1 U7700 ( .A1(n6144), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6128) );
  XNOR2_X1 U7701 ( .A(n6128), .B(P1_IR_REG_9__SCAN_IN), .ZN(n6859) );
  AOI22_X1 U7702 ( .A1(n6859), .A2(n6620), .B1(n8824), .B2(
        P2_DATAO_REG_9__SCAN_IN), .ZN(n6129) );
  NAND2_X1 U7703 ( .A1(n8720), .A2(n6499), .ZN(n6137) );
  NAND2_X1 U7704 ( .A1(n6582), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n6135) );
  INV_X1 U7705 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n6855) );
  OR2_X1 U7706 ( .A1(n6116), .A2(n6855), .ZN(n6134) );
  INV_X1 U7707 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n6150) );
  XNOR2_X1 U7708 ( .A(n6152), .B(n6150), .ZN(n8718) );
  OR2_X1 U7709 ( .A1(n4264), .A2(n8718), .ZN(n6133) );
  INV_X1 U7710 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n6131) );
  OR2_X1 U7711 ( .A1(n6584), .A2(n6131), .ZN(n6132) );
  NAND4_X1 U7712 ( .A1(n6135), .A2(n6134), .A3(n6133), .A4(n6132), .ZN(n9110)
         );
  NAND2_X1 U7713 ( .A1(n4260), .A2(n9110), .ZN(n6136) );
  NAND2_X1 U7714 ( .A1(n6137), .A2(n6136), .ZN(n6138) );
  XNOR2_X1 U7715 ( .A(n6138), .B(n6081), .ZN(n6141) );
  INV_X1 U7716 ( .A(n9110), .ZN(n7518) );
  NOR2_X1 U7717 ( .A1(n6397), .A2(n7518), .ZN(n6139) );
  AOI21_X1 U7718 ( .B1(n8720), .B2(n4260), .A(n6139), .ZN(n6140) );
  NOR2_X1 U7719 ( .A1(n6141), .A2(n6140), .ZN(n8617) );
  AOI21_X1 U7720 ( .B1(n8613), .B2(n8612), .A(n8617), .ZN(n6143) );
  NOR3_X1 U7721 ( .A1(n8617), .A2(n8613), .A3(n8612), .ZN(n6142) );
  AND2_X1 U7722 ( .A1(n6141), .A2(n6140), .ZN(n8621) );
  NAND2_X1 U7723 ( .A1(n6610), .A2(n8822), .ZN(n6147) );
  NAND2_X1 U7724 ( .A1(n6179), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6145) );
  XNOR2_X1 U7725 ( .A(n6145), .B(P1_IR_REG_10__SCAN_IN), .ZN(n6880) );
  AOI22_X1 U7726 ( .A1(n6880), .A2(n6620), .B1(n8824), .B2(
        P2_DATAO_REG_10__SCAN_IN), .ZN(n6146) );
  NAND2_X1 U7727 ( .A1(n7513), .A2(n4260), .ZN(n6160) );
  NAND2_X1 U7728 ( .A1(n6582), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n6158) );
  INV_X1 U7729 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n6148) );
  OR2_X1 U7730 ( .A1(n6116), .A2(n6148), .ZN(n6157) );
  INV_X1 U7731 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n6149) );
  OAI21_X1 U7732 ( .B1(n6152), .B2(n6150), .A(n6149), .ZN(n6153) );
  NAND2_X1 U7733 ( .A1(P1_REG3_REG_9__SCAN_IN), .A2(P1_REG3_REG_10__SCAN_IN), 
        .ZN(n6151) );
  OR2_X2 U7734 ( .A1(n6152), .A2(n6151), .ZN(n6184) );
  NAND2_X1 U7735 ( .A1(n6153), .A2(n6184), .ZN(n8625) );
  OR2_X1 U7736 ( .A1(n4264), .A2(n8625), .ZN(n6156) );
  INV_X1 U7737 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n6154) );
  OR2_X1 U7738 ( .A1(n6584), .A2(n6154), .ZN(n6155) );
  OR2_X1 U7739 ( .A1(n6397), .A2(n8760), .ZN(n6159) );
  NAND2_X1 U7740 ( .A1(n6160), .A2(n6159), .ZN(n8618) );
  INV_X1 U7741 ( .A(n8618), .ZN(n6197) );
  NAND2_X1 U7742 ( .A1(n7513), .A2(n6499), .ZN(n6162) );
  INV_X1 U7743 ( .A(n8760), .ZN(n9109) );
  NAND2_X1 U7744 ( .A1(n4260), .A2(n9109), .ZN(n6161) );
  NAND2_X1 U7745 ( .A1(n6162), .A2(n6161), .ZN(n6163) );
  XNOR2_X1 U7746 ( .A(n6163), .B(n6497), .ZN(n8619) );
  INV_X1 U7747 ( .A(n8619), .ZN(n6198) );
  NAND2_X1 U7748 ( .A1(n6758), .A2(n8822), .ZN(n6167) );
  OR2_X1 U7749 ( .A1(n6164), .A2(n6275), .ZN(n6165) );
  XNOR2_X1 U7750 ( .A(n6165), .B(P1_IR_REG_12__SCAN_IN), .ZN(n7237) );
  AOI22_X1 U7751 ( .A1(n6003), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n6620), .B2(
        n7237), .ZN(n6166) );
  NAND2_X1 U7752 ( .A1(n8657), .A2(n6499), .ZN(n6175) );
  NAND2_X1 U7753 ( .A1(n6582), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n6173) );
  INV_X1 U7754 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n6168) );
  OR2_X1 U7755 ( .A1(n6584), .A2(n6168), .ZN(n6172) );
  AND2_X2 U7756 ( .A1(n6185), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n6210) );
  NOR2_X1 U7757 ( .A1(n6185), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n6169) );
  OR2_X1 U7758 ( .A1(n6210), .A2(n6169), .ZN(n8669) );
  OR2_X1 U7759 ( .A1(n4264), .A2(n8669), .ZN(n6171) );
  INV_X1 U7760 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n6997) );
  OR2_X1 U7761 ( .A1(n6116), .A2(n6997), .ZN(n6170) );
  INV_X1 U7762 ( .A(n8737), .ZN(n9107) );
  NAND2_X1 U7763 ( .A1(n4260), .A2(n9107), .ZN(n6174) );
  NAND2_X1 U7764 ( .A1(n6175), .A2(n6174), .ZN(n6176) );
  XNOR2_X1 U7765 ( .A(n6176), .B(n6497), .ZN(n6202) );
  NAND2_X1 U7766 ( .A1(n8657), .A2(n4260), .ZN(n6178) );
  OR2_X1 U7767 ( .A1(n6397), .A2(n8737), .ZN(n6177) );
  NAND2_X1 U7768 ( .A1(n6178), .A2(n6177), .ZN(n6203) );
  NAND2_X1 U7769 ( .A1(n6202), .A2(n6203), .ZN(n8660) );
  NAND2_X1 U7770 ( .A1(n6608), .A2(n8822), .ZN(n6182) );
  OAI21_X1 U7771 ( .B1(n6179), .B2(P1_IR_REG_10__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n6180) );
  XNOR2_X1 U7772 ( .A(n6180), .B(P1_IR_REG_11__SCAN_IN), .ZN(n7006) );
  AOI22_X1 U7773 ( .A1(n7006), .A2(n6620), .B1(n8824), .B2(
        P2_DATAO_REG_11__SCAN_IN), .ZN(n6181) );
  NAND2_X1 U7774 ( .A1(n7716), .A2(n6499), .ZN(n6192) );
  NAND2_X1 U7775 ( .A1(n6524), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n6190) );
  INV_X1 U7776 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n7671) );
  OR2_X1 U7777 ( .A1(n6051), .A2(n7671), .ZN(n6189) );
  AND2_X1 U7778 ( .A1(n6184), .A2(n6183), .ZN(n6186) );
  OR2_X1 U7779 ( .A1(n6186), .A2(n6185), .ZN(n8761) );
  OR2_X1 U7780 ( .A1(n4264), .A2(n8761), .ZN(n6188) );
  INV_X1 U7781 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n9938) );
  OR2_X1 U7782 ( .A1(n6584), .A2(n9938), .ZN(n6187) );
  NAND4_X1 U7783 ( .A1(n6190), .A2(n6189), .A3(n6188), .A4(n6187), .ZN(n9108)
         );
  NAND2_X1 U7784 ( .A1(n4260), .A2(n9108), .ZN(n6191) );
  NAND2_X1 U7785 ( .A1(n6192), .A2(n6191), .ZN(n6193) );
  XNOR2_X1 U7786 ( .A(n6193), .B(n6497), .ZN(n8659) );
  INV_X1 U7787 ( .A(n9108), .ZN(n8668) );
  NOR2_X1 U7788 ( .A1(n6397), .A2(n8668), .ZN(n6194) );
  AOI21_X1 U7789 ( .B1(n7716), .B2(n4260), .A(n6194), .ZN(n6196) );
  INV_X1 U7790 ( .A(n6196), .ZN(n8658) );
  NAND2_X1 U7791 ( .A1(n8659), .A2(n8658), .ZN(n8665) );
  OAI211_X1 U7792 ( .C1(n6197), .C2(n6198), .A(n8660), .B(n8665), .ZN(n6195)
         );
  NOR2_X1 U7793 ( .A1(n8619), .A2(n8618), .ZN(n8755) );
  NOR2_X1 U7794 ( .A1(n8755), .A2(n6196), .ZN(n6200) );
  NAND3_X1 U7795 ( .A1(n6198), .A2(n6197), .A3(n6196), .ZN(n6199) );
  OAI21_X1 U7796 ( .B1(n6200), .B2(n8659), .A(n6199), .ZN(n6201) );
  NAND2_X1 U7797 ( .A1(n6201), .A2(n8660), .ZN(n6206) );
  INV_X1 U7798 ( .A(n6202), .ZN(n6205) );
  INV_X1 U7799 ( .A(n6203), .ZN(n6204) );
  NAND2_X1 U7800 ( .A1(n6205), .A2(n6204), .ZN(n8731) );
  NAND2_X1 U7801 ( .A1(n6793), .A2(n6274), .ZN(n6209) );
  INV_X1 U7802 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n9910) );
  NAND2_X1 U7803 ( .A1(n6164), .A2(n9910), .ZN(n6226) );
  NAND2_X1 U7804 ( .A1(n6226), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6207) );
  XNOR2_X1 U7805 ( .A(n6207), .B(P1_IR_REG_13__SCAN_IN), .ZN(n7270) );
  AOI22_X1 U7806 ( .A1(n6003), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n7270), .B2(
        n6620), .ZN(n6208) );
  NAND2_X1 U7807 ( .A1(n9533), .A2(n6499), .ZN(n6219) );
  NAND2_X1 U7808 ( .A1(n6582), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n6217) );
  OR2_X1 U7809 ( .A1(n6210), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n6211) );
  NAND2_X1 U7810 ( .A1(n6230), .A2(n6211), .ZN(n8738) );
  OR2_X1 U7811 ( .A1(n4264), .A2(n8738), .ZN(n6216) );
  INV_X1 U7812 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n6212) );
  OR2_X1 U7813 ( .A1(n6584), .A2(n6212), .ZN(n6215) );
  INV_X1 U7814 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n6213) );
  OR2_X1 U7815 ( .A1(n6116), .A2(n6213), .ZN(n6214) );
  NAND4_X1 U7816 ( .A1(n6217), .A2(n6216), .A3(n6215), .A4(n6214), .ZN(n9106)
         );
  NAND2_X1 U7817 ( .A1(n4260), .A2(n9106), .ZN(n6218) );
  NAND2_X1 U7818 ( .A1(n6219), .A2(n6218), .ZN(n6220) );
  XNOR2_X1 U7819 ( .A(n6220), .B(n6497), .ZN(n6224) );
  NOR2_X1 U7820 ( .A1(n6397), .A2(n9417), .ZN(n6221) );
  AOI21_X1 U7821 ( .B1(n9533), .B2(n4260), .A(n6221), .ZN(n6222) );
  XNOR2_X1 U7822 ( .A(n6224), .B(n6222), .ZN(n8732) );
  INV_X1 U7823 ( .A(n6222), .ZN(n6223) );
  OR2_X1 U7824 ( .A1(n6224), .A2(n6223), .ZN(n6225) );
  NAND2_X1 U7825 ( .A1(n6795), .A2(n6274), .ZN(n6228) );
  OR2_X1 U7826 ( .A1(n6226), .A2(P1_IR_REG_13__SCAN_IN), .ZN(n6261) );
  NAND2_X1 U7827 ( .A1(n6261), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6241) );
  XNOR2_X1 U7828 ( .A(n6241), .B(P1_IR_REG_14__SCAN_IN), .ZN(n9155) );
  AOI22_X1 U7829 ( .A1(n9155), .A2(n6620), .B1(n8824), .B2(
        P2_DATAO_REG_14__SCAN_IN), .ZN(n6227) );
  INV_X1 U7830 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n6229) );
  OR2_X2 U7831 ( .A1(n6230), .A2(n6229), .ZN(n6246) );
  NAND2_X1 U7832 ( .A1(n6230), .A2(n6229), .ZN(n6231) );
  NAND2_X1 U7833 ( .A1(n6246), .A2(n6231), .ZN(n9424) );
  OR2_X1 U7834 ( .A1(n9424), .A2(n4264), .ZN(n6235) );
  INV_X1 U7835 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n7276) );
  OR2_X1 U7836 ( .A1(n6116), .A2(n7276), .ZN(n6234) );
  NAND2_X1 U7837 ( .A1(n6582), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n6233) );
  INV_X1 U7838 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n10006) );
  OR2_X1 U7839 ( .A1(n6584), .A2(n10006), .ZN(n6232) );
  NAND4_X1 U7840 ( .A1(n6235), .A2(n6234), .A3(n6233), .A4(n6232), .ZN(n9397)
         );
  AOI22_X1 U7841 ( .A1(n9530), .A2(n6499), .B1(n4260), .B2(n9397), .ZN(n6236)
         );
  XNOR2_X1 U7842 ( .A(n6236), .B(n6497), .ZN(n6238) );
  INV_X1 U7843 ( .A(n9530), .ZN(n6237) );
  OAI22_X1 U7844 ( .A1(n6237), .A2(n4282), .B1(n8846), .B2(n6397), .ZN(n8592)
         );
  INV_X1 U7845 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n6240) );
  NAND2_X1 U7846 ( .A1(n6241), .A2(n6240), .ZN(n6242) );
  NAND2_X1 U7847 ( .A1(n6242), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6243) );
  XNOR2_X1 U7848 ( .A(n6243), .B(P1_IR_REG_15__SCAN_IN), .ZN(n9614) );
  AOI22_X1 U7849 ( .A1(n9614), .A2(n6620), .B1(n8824), .B2(
        P2_DATAO_REG_15__SCAN_IN), .ZN(n6244) );
  NAND2_X1 U7850 ( .A1(n9524), .A2(n6499), .ZN(n6253) );
  INV_X1 U7851 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n6245) );
  OR2_X2 U7852 ( .A1(n6246), .A2(n6245), .ZN(n6265) );
  NAND2_X1 U7853 ( .A1(n6246), .A2(n6245), .ZN(n6247) );
  NAND2_X1 U7854 ( .A1(n6265), .A2(n6247), .ZN(n9401) );
  INV_X1 U7855 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n9157) );
  OR2_X1 U7856 ( .A1(n6116), .A2(n9157), .ZN(n6249) );
  INV_X1 U7857 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n9402) );
  OR2_X1 U7858 ( .A1(n6051), .A2(n9402), .ZN(n6248) );
  AND2_X1 U7859 ( .A1(n6249), .A2(n6248), .ZN(n6251) );
  NAND2_X1 U7860 ( .A1(n6087), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n6250) );
  OAI211_X1 U7861 ( .C1(n9401), .C2(n4264), .A(n6251), .B(n6250), .ZN(n9387)
         );
  NAND2_X1 U7862 ( .A1(n4260), .A2(n9387), .ZN(n6252) );
  NAND2_X1 U7863 ( .A1(n6253), .A2(n6252), .ZN(n6254) );
  XNOR2_X1 U7864 ( .A(n6254), .B(n6081), .ZN(n8803) );
  INV_X1 U7865 ( .A(n9387), .ZN(n9418) );
  NOR2_X1 U7866 ( .A1(n6397), .A2(n9418), .ZN(n6255) );
  AOI21_X1 U7867 ( .B1(n9524), .B2(n4260), .A(n6255), .ZN(n8802) );
  NAND2_X1 U7868 ( .A1(n8803), .A2(n8802), .ZN(n6258) );
  INV_X1 U7869 ( .A(n8803), .ZN(n6257) );
  INV_X1 U7870 ( .A(n8802), .ZN(n6256) );
  NAND2_X1 U7871 ( .A1(n6973), .A2(n8822), .ZN(n6264) );
  INV_X1 U7872 ( .A(n6259), .ZN(n6260) );
  OAI21_X1 U7873 ( .B1(n6261), .B2(n6260), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n6262) );
  XNOR2_X1 U7874 ( .A(n6262), .B(P1_IR_REG_16__SCAN_IN), .ZN(n9626) );
  AOI22_X1 U7875 ( .A1(n9626), .A2(n6620), .B1(n8824), .B2(
        P2_DATAO_REG_16__SCAN_IN), .ZN(n6263) );
  AND2_X1 U7876 ( .A1(n6265), .A2(n9972), .ZN(n6266) );
  OR2_X1 U7877 ( .A1(n6266), .A2(n6282), .ZN(n9379) );
  AOI22_X1 U7878 ( .A1(n6524), .A2(P1_REG1_REG_16__SCAN_IN), .B1(n6582), .B2(
        P1_REG2_REG_16__SCAN_IN), .ZN(n6268) );
  NAND2_X1 U7879 ( .A1(n6087), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n6267) );
  OAI211_X1 U7880 ( .C1(n9379), .C2(n4264), .A(n6268), .B(n6267), .ZN(n9399)
         );
  AOI22_X1 U7881 ( .A1(n9382), .A2(n6499), .B1(n4260), .B2(n9399), .ZN(n6269)
         );
  XOR2_X1 U7882 ( .A(n7322), .B(n6269), .Z(n6272) );
  INV_X1 U7883 ( .A(n9382), .ZN(n6270) );
  INV_X1 U7884 ( .A(n9399), .ZN(n8698) );
  OAI22_X1 U7885 ( .A1(n6270), .A2(n4282), .B1(n8698), .B2(n6397), .ZN(n6271)
         );
  NOR2_X1 U7886 ( .A1(n6272), .A2(n6271), .ZN(n6273) );
  AOI21_X1 U7887 ( .B1(n6272), .B2(n6271), .A(n6273), .ZN(n8687) );
  NAND2_X1 U7888 ( .A1(n6921), .A2(n6274), .ZN(n6281) );
  NOR2_X1 U7889 ( .A1(n5935), .A2(n6275), .ZN(n6276) );
  MUX2_X1 U7890 ( .A(n6275), .B(n6276), .S(P1_IR_REG_17__SCAN_IN), .Z(n6279)
         );
  INV_X1 U7891 ( .A(n6277), .ZN(n6278) );
  NOR2_X1 U7892 ( .A1(n6279), .A2(n6278), .ZN(n9158) );
  AOI22_X1 U7893 ( .A1(n9158), .A2(n6620), .B1(n8824), .B2(
        P2_DATAO_REG_17__SCAN_IN), .ZN(n6280) );
  OR2_X1 U7894 ( .A1(n6282), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n6283) );
  NAND2_X1 U7895 ( .A1(n6297), .A2(n6283), .ZN(n9365) );
  AOI22_X1 U7896 ( .A1(n6582), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n6087), .B2(
        P1_REG0_REG_17__SCAN_IN), .ZN(n6285) );
  NAND2_X1 U7897 ( .A1(n6524), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n6284) );
  OAI211_X1 U7898 ( .C1(n9365), .C2(n4264), .A(n6285), .B(n6284), .ZN(n9386)
         );
  INV_X1 U7899 ( .A(n9386), .ZN(n8784) );
  OAI22_X1 U7900 ( .A1(n9368), .A2(n4282), .B1(n8784), .B2(n6397), .ZN(n6289)
         );
  NAND2_X1 U7901 ( .A1(n9514), .A2(n6499), .ZN(n6287) );
  NAND2_X1 U7902 ( .A1(n9386), .A2(n4260), .ZN(n6286) );
  NAND2_X1 U7903 ( .A1(n6287), .A2(n6286), .ZN(n6288) );
  XNOR2_X1 U7904 ( .A(n6288), .B(n6497), .ZN(n6290) );
  XOR2_X1 U7905 ( .A(n6289), .B(n6290), .Z(n8696) );
  NAND2_X1 U7906 ( .A1(n7097), .A2(n8822), .ZN(n6295) );
  NAND2_X1 U7907 ( .A1(n6277), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6292) );
  MUX2_X1 U7908 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6292), .S(
        P1_IR_REG_18__SCAN_IN), .Z(n6293) );
  AND2_X1 U7909 ( .A1(n6476), .A2(n6293), .ZN(n9152) );
  AOI22_X1 U7910 ( .A1(n9152), .A2(n6620), .B1(n8824), .B2(
        P2_DATAO_REG_18__SCAN_IN), .ZN(n6294) );
  NAND2_X1 U7911 ( .A1(n9357), .A2(n4260), .ZN(n6305) );
  INV_X1 U7912 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n6296) );
  NAND2_X1 U7913 ( .A1(n6297), .A2(n6296), .ZN(n6298) );
  AND2_X1 U7914 ( .A1(n6311), .A2(n6298), .ZN(n9349) );
  INV_X1 U7915 ( .A(n4264), .ZN(n6347) );
  NAND2_X1 U7916 ( .A1(n9349), .A2(n6347), .ZN(n6303) );
  INV_X1 U7917 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n9161) );
  NAND2_X1 U7918 ( .A1(n6087), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n6300) );
  INV_X1 U7919 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n9351) );
  OR2_X1 U7920 ( .A1(n6051), .A2(n9351), .ZN(n6299) );
  OAI211_X1 U7921 ( .C1(n6116), .C2(n9161), .A(n6300), .B(n6299), .ZN(n6301)
         );
  INV_X1 U7922 ( .A(n6301), .ZN(n6302) );
  NAND2_X1 U7923 ( .A1(n9363), .A2(n6445), .ZN(n6304) );
  NAND2_X1 U7924 ( .A1(n6305), .A2(n6304), .ZN(n8781) );
  NAND2_X1 U7925 ( .A1(n9357), .A2(n6499), .ZN(n6307) );
  NAND2_X1 U7926 ( .A1(n9363), .A2(n4260), .ZN(n6306) );
  NAND2_X1 U7927 ( .A1(n6307), .A2(n6306), .ZN(n6308) );
  XNOR2_X1 U7928 ( .A(n6308), .B(n6497), .ZN(n8636) );
  NAND2_X1 U7929 ( .A1(n7206), .A2(n8822), .ZN(n6310) );
  AOI22_X1 U7930 ( .A1(n9169), .A2(n6620), .B1(n8824), .B2(
        P2_DATAO_REG_19__SCAN_IN), .ZN(n6309) );
  NAND2_X1 U7931 ( .A1(n9503), .A2(n6499), .ZN(n6318) );
  INV_X1 U7932 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n10029) );
  AND2_X1 U7933 ( .A1(n6311), .A2(n10029), .ZN(n6312) );
  OR2_X1 U7934 ( .A1(n6312), .A2(n6330), .ZN(n9326) );
  INV_X1 U7935 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n10033) );
  NAND2_X1 U7936 ( .A1(n6582), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n6314) );
  NAND2_X1 U7937 ( .A1(n6087), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n6313) );
  OAI211_X1 U7938 ( .C1(n6116), .C2(n10033), .A(n6314), .B(n6313), .ZN(n6315)
         );
  INV_X1 U7939 ( .A(n6315), .ZN(n6316) );
  NAND2_X1 U7940 ( .A1(n9346), .A2(n4260), .ZN(n6317) );
  NAND2_X1 U7941 ( .A1(n6318), .A2(n6317), .ZN(n6319) );
  XNOR2_X1 U7942 ( .A(n6319), .B(n6081), .ZN(n6321) );
  AND2_X1 U7943 ( .A1(n9346), .A2(n6445), .ZN(n6320) );
  AOI21_X1 U7944 ( .B1(n9503), .B2(n4260), .A(n6320), .ZN(n6322) );
  NOR2_X1 U7945 ( .A1(n6321), .A2(n6322), .ZN(n8634) );
  AOI21_X1 U7946 ( .B1(n8781), .B2(n8636), .A(n8634), .ZN(n6327) );
  INV_X1 U7947 ( .A(n6321), .ZN(n6324) );
  INV_X1 U7948 ( .A(n6322), .ZN(n6323) );
  NOR2_X1 U7949 ( .A1(n6324), .A2(n6323), .ZN(n8633) );
  NAND2_X1 U7950 ( .A1(n7245), .A2(n8822), .ZN(n6329) );
  NAND2_X1 U7951 ( .A1(n8824), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n6328) );
  NAND2_X1 U7952 ( .A1(n9498), .A2(n6499), .ZN(n6338) );
  NOR2_X1 U7953 ( .A1(n6330), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n6331) );
  OR2_X1 U7954 ( .A1(n6345), .A2(n6331), .ZN(n9313) );
  INV_X1 U7955 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n6334) );
  NAND2_X1 U7956 ( .A1(n6087), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n6333) );
  NAND2_X1 U7957 ( .A1(n6582), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n6332) );
  OAI211_X1 U7958 ( .C1(n6116), .C2(n6334), .A(n6333), .B(n6332), .ZN(n6335)
         );
  INV_X1 U7959 ( .A(n6335), .ZN(n6336) );
  NAND2_X1 U7960 ( .A1(n9324), .A2(n4260), .ZN(n6337) );
  NAND2_X1 U7961 ( .A1(n6338), .A2(n6337), .ZN(n6339) );
  XNOR2_X1 U7962 ( .A(n6339), .B(n6081), .ZN(n6342) );
  AND2_X1 U7963 ( .A1(n9324), .A2(n6445), .ZN(n6340) );
  AOI21_X1 U7964 ( .B1(n9498), .B2(n4260), .A(n6340), .ZN(n6341) );
  NOR2_X1 U7965 ( .A1(n6342), .A2(n6341), .ZN(n8723) );
  NAND2_X1 U7966 ( .A1(n7172), .A2(n8822), .ZN(n6344) );
  NAND2_X1 U7967 ( .A1(n8824), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n6343) );
  NAND2_X2 U7968 ( .A1(n6344), .A2(n6343), .ZN(n9492) );
  NAND2_X1 U7969 ( .A1(n9492), .A2(n6499), .ZN(n6355) );
  OR2_X1 U7970 ( .A1(n6345), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n6346) );
  AND2_X1 U7971 ( .A1(n6346), .A2(n6363), .ZN(n9292) );
  NAND2_X1 U7972 ( .A1(n9292), .A2(n6347), .ZN(n6353) );
  INV_X1 U7973 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n6350) );
  NAND2_X1 U7974 ( .A1(n6582), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n6349) );
  NAND2_X1 U7975 ( .A1(n6087), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n6348) );
  OAI211_X1 U7976 ( .C1(n6350), .C2(n6116), .A(n6349), .B(n6348), .ZN(n6351)
         );
  INV_X1 U7977 ( .A(n6351), .ZN(n6352) );
  NAND2_X1 U7978 ( .A1(n9310), .A2(n4260), .ZN(n6354) );
  NAND2_X1 U7979 ( .A1(n6355), .A2(n6354), .ZN(n6356) );
  XNOR2_X1 U7980 ( .A(n6356), .B(n6081), .ZN(n6359) );
  NOR2_X1 U7981 ( .A1(n7882), .A2(n6397), .ZN(n6357) );
  AOI21_X1 U7982 ( .B1(n9492), .B2(n4260), .A(n6357), .ZN(n6358) );
  OR2_X1 U7983 ( .A1(n6359), .A2(n6358), .ZN(n8646) );
  NAND2_X1 U7984 ( .A1(n7406), .A2(n8822), .ZN(n6361) );
  NAND2_X1 U7985 ( .A1(n8824), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n6360) );
  NAND2_X1 U7986 ( .A1(n6582), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n6369) );
  INV_X1 U7987 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n6362) );
  OR2_X1 U7988 ( .A1(n6116), .A2(n6362), .ZN(n6368) );
  OAI21_X1 U7989 ( .B1(P1_REG3_REG_22__SCAN_IN), .B2(n6364), .A(n6376), .ZN(
        n9276) );
  OR2_X1 U7990 ( .A1(n4264), .A2(n9276), .ZN(n6367) );
  INV_X1 U7991 ( .A(P1_REG0_REG_22__SCAN_IN), .ZN(n6365) );
  OR2_X1 U7992 ( .A1(n6584), .A2(n6365), .ZN(n6366) );
  AND4_X2 U7993 ( .A1(n6369), .A2(n6368), .A3(n6367), .A4(n6366), .ZN(n8652)
         );
  OAI22_X1 U7994 ( .A1(n9280), .A2(n4282), .B1(n8652), .B2(n6397), .ZN(n6371)
         );
  OAI22_X1 U7995 ( .A1(n9280), .A2(n6045), .B1(n8652), .B2(n4282), .ZN(n6370)
         );
  XOR2_X1 U7996 ( .A(n7322), .B(n6370), .Z(n8746) );
  NAND2_X1 U7997 ( .A1(n8745), .A2(n8746), .ZN(n6372) );
  NAND2_X1 U7998 ( .A1(n7342), .A2(n8822), .ZN(n6374) );
  NAND2_X1 U7999 ( .A1(n8824), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n6373) );
  OR2_X1 U8000 ( .A1(n9265), .A2(n4282), .ZN(n6384) );
  NAND2_X1 U8001 ( .A1(n6524), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n6382) );
  INV_X1 U8002 ( .A(P1_REG2_REG_23__SCAN_IN), .ZN(n6375) );
  OR2_X1 U8003 ( .A1(n6051), .A2(n6375), .ZN(n6381) );
  OAI21_X1 U8004 ( .B1(P1_REG3_REG_23__SCAN_IN), .B2(n6377), .A(n6389), .ZN(
        n9262) );
  OR2_X1 U8005 ( .A1(n4264), .A2(n9262), .ZN(n6380) );
  INV_X1 U8006 ( .A(P1_REG0_REG_23__SCAN_IN), .ZN(n6378) );
  OR2_X1 U8007 ( .A1(n6584), .A2(n6378), .ZN(n6379) );
  OR2_X1 U8008 ( .A1(n6397), .A2(n8833), .ZN(n6383) );
  NAND2_X1 U8009 ( .A1(n6384), .A2(n6383), .ZN(n8604) );
  OAI22_X1 U8010 ( .A1(n9265), .A2(n6045), .B1(n8833), .B2(n4282), .ZN(n6385)
         );
  XNOR2_X1 U8011 ( .A(n6385), .B(n6497), .ZN(n8602) );
  NAND2_X1 U8012 ( .A1(n8824), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n6386) );
  NAND2_X1 U8013 ( .A1(n6524), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n6395) );
  INV_X1 U8014 ( .A(P1_REG2_REG_24__SCAN_IN), .ZN(n6387) );
  OR2_X1 U8015 ( .A1(n6051), .A2(n6387), .ZN(n6394) );
  INV_X1 U8016 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n8706) );
  NAND2_X1 U8017 ( .A1(n6389), .A2(n8706), .ZN(n6390) );
  NAND2_X1 U8018 ( .A1(n6412), .A2(n6390), .ZN(n9250) );
  INV_X1 U8019 ( .A(P1_REG0_REG_24__SCAN_IN), .ZN(n6391) );
  OR2_X1 U8020 ( .A1(n6584), .A2(n6391), .ZN(n6392) );
  OAI22_X1 U8021 ( .A1(n9253), .A2(n6045), .B1(n7900), .B2(n4282), .ZN(n6396)
         );
  XNOR2_X1 U8022 ( .A(n6396), .B(n6081), .ZN(n6401) );
  OR2_X1 U8023 ( .A1(n9253), .A2(n4282), .ZN(n6399) );
  OR2_X1 U8024 ( .A1(n6397), .A2(n7900), .ZN(n6398) );
  AOI21_X1 U8025 ( .B1(n8604), .B2(n8602), .A(n8677), .ZN(n6400) );
  NAND2_X1 U8026 ( .A1(n8600), .A2(n6400), .ZN(n6421) );
  NOR2_X1 U8027 ( .A1(n8602), .A2(n8604), .ZN(n6406) );
  INV_X1 U8028 ( .A(n8677), .ZN(n6405) );
  INV_X1 U8029 ( .A(n6401), .ZN(n6404) );
  INV_X1 U8030 ( .A(n6402), .ZN(n6403) );
  NOR2_X1 U8031 ( .A1(n6404), .A2(n6403), .ZN(n8679) );
  AOI21_X1 U8032 ( .B1(n6406), .B2(n6405), .A(n8679), .ZN(n6420) );
  NAND2_X1 U8033 ( .A1(n7632), .A2(n8822), .ZN(n6408) );
  NAND2_X1 U8034 ( .A1(n8824), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n6407) );
  NAND2_X1 U8035 ( .A1(n6582), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n6418) );
  INV_X1 U8036 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n6409) );
  OR2_X1 U8037 ( .A1(n6116), .A2(n6409), .ZN(n6417) );
  INV_X1 U8038 ( .A(n6412), .ZN(n6410) );
  INV_X1 U8039 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n6411) );
  NAND2_X1 U8040 ( .A1(n6412), .A2(n6411), .ZN(n6413) );
  NAND2_X1 U8041 ( .A1(n6428), .A2(n6413), .ZN(n9235) );
  INV_X1 U8042 ( .A(P1_REG0_REG_25__SCAN_IN), .ZN(n6414) );
  OR2_X1 U8043 ( .A1(n6584), .A2(n6414), .ZN(n6415) );
  AND4_X2 U8044 ( .A1(n6418), .A2(n6417), .A3(n6416), .A4(n6415), .ZN(n8796)
         );
  OAI22_X1 U8045 ( .A1(n9238), .A2(n6045), .B1(n8796), .B2(n4282), .ZN(n6419)
         );
  XNOR2_X1 U8046 ( .A(n6419), .B(n6497), .ZN(n6423) );
  OAI22_X1 U8047 ( .A1(n9238), .A2(n4282), .B1(n8796), .B2(n6397), .ZN(n6422)
         );
  XNOR2_X1 U8048 ( .A(n6423), .B(n6422), .ZN(n8678) );
  NOR2_X1 U8049 ( .A1(n6423), .A2(n6422), .ZN(n8791) );
  NAND2_X1 U8050 ( .A1(n7710), .A2(n8822), .ZN(n6425) );
  NAND2_X1 U8051 ( .A1(n8824), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n6424) );
  NAND2_X1 U8052 ( .A1(n6524), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n6434) );
  INV_X1 U8053 ( .A(P1_REG2_REG_26__SCAN_IN), .ZN(n6426) );
  OR2_X1 U8054 ( .A1(n6051), .A2(n6426), .ZN(n6433) );
  INV_X1 U8055 ( .A(n6428), .ZN(n6427) );
  INV_X1 U8056 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n10036) );
  NAND2_X1 U8057 ( .A1(n6428), .A2(n10036), .ZN(n6429) );
  INV_X1 U8058 ( .A(P1_REG0_REG_26__SCAN_IN), .ZN(n6430) );
  OR2_X1 U8059 ( .A1(n6584), .A2(n6430), .ZN(n6431) );
  AND4_X2 U8060 ( .A1(n6434), .A2(n6433), .A3(n6432), .A4(n6431), .ZN(n7901)
         );
  OAI22_X1 U8061 ( .A1(n9225), .A2(n6045), .B1(n7901), .B2(n4282), .ZN(n6435)
         );
  XNOR2_X1 U8062 ( .A(n6435), .B(n6497), .ZN(n6449) );
  OAI22_X1 U8063 ( .A1(n9225), .A2(n4282), .B1(n7901), .B2(n6397), .ZN(n6448)
         );
  XNOR2_X1 U8064 ( .A(n6449), .B(n6448), .ZN(n8790) );
  NAND2_X1 U8065 ( .A1(n7808), .A2(n8822), .ZN(n6437) );
  NAND2_X1 U8066 ( .A1(n8824), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n6436) );
  NAND2_X1 U8067 ( .A1(n6524), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n6443) );
  INV_X1 U8068 ( .A(P1_REG2_REG_27__SCAN_IN), .ZN(n6438) );
  OR2_X1 U8069 ( .A1(n6051), .A2(n6438), .ZN(n6442) );
  INV_X1 U8070 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n7864) );
  XNOR2_X1 U8071 ( .A(n6486), .B(n7864), .ZN(n9208) );
  INV_X1 U8072 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n6439) );
  OR2_X1 U8073 ( .A1(n6584), .A2(n6439), .ZN(n6440) );
  AND4_X2 U8074 ( .A1(n6443), .A2(n6442), .A3(n6441), .A4(n6440), .ZN(n7890)
         );
  OAI22_X1 U8075 ( .A1(n9211), .A2(n6045), .B1(n7890), .B2(n4282), .ZN(n6444)
         );
  XOR2_X1 U8076 ( .A(n7322), .B(n6444), .Z(n6447) );
  AOI22_X1 U8077 ( .A1(n9462), .A2(n4260), .B1(n6445), .B2(n9228), .ZN(n6446)
         );
  NAND2_X1 U8078 ( .A1(n6447), .A2(n6446), .ZN(n6533) );
  OAI21_X1 U8079 ( .B1(n6447), .B2(n6446), .A(n6533), .ZN(n7859) );
  AND2_X1 U8080 ( .A1(n6449), .A2(n6448), .ZN(n7858) );
  NOR2_X1 U8081 ( .A1(n7859), .A2(n7858), .ZN(n6450) );
  INV_X1 U8082 ( .A(n6464), .ZN(n7634) );
  NAND2_X1 U8083 ( .A1(n7634), .A2(P1_B_REG_SCAN_IN), .ZN(n6451) );
  MUX2_X1 U8084 ( .A(n6451), .B(P1_B_REG_SCAN_IN), .S(n6469), .Z(n6452) );
  NAND2_X1 U8085 ( .A1(n6452), .A2(n6468), .ZN(n9717) );
  NOR4_X1 U8086 ( .A1(P1_D_REG_17__SCAN_IN), .A2(P1_D_REG_18__SCAN_IN), .A3(
        P1_D_REG_19__SCAN_IN), .A4(P1_D_REG_20__SCAN_IN), .ZN(n6456) );
  NOR4_X1 U8087 ( .A1(P1_D_REG_15__SCAN_IN), .A2(P1_D_REG_13__SCAN_IN), .A3(
        P1_D_REG_14__SCAN_IN), .A4(P1_D_REG_16__SCAN_IN), .ZN(n6455) );
  NOR4_X1 U8088 ( .A1(P1_D_REG_25__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n6454) );
  NOR4_X1 U8089 ( .A1(P1_D_REG_21__SCAN_IN), .A2(P1_D_REG_22__SCAN_IN), .A3(
        P1_D_REG_23__SCAN_IN), .A4(P1_D_REG_24__SCAN_IN), .ZN(n6453) );
  NAND4_X1 U8090 ( .A1(n6456), .A2(n6455), .A3(n6454), .A4(n6453), .ZN(n6462)
         );
  NOR2_X1 U8091 ( .A1(P1_D_REG_9__SCAN_IN), .A2(P1_D_REG_26__SCAN_IN), .ZN(
        n6460) );
  NOR4_X1 U8092 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        P1_D_REG_2__SCAN_IN), .A4(P1_D_REG_3__SCAN_IN), .ZN(n6459) );
  NOR4_X1 U8093 ( .A1(P1_D_REG_8__SCAN_IN), .A2(P1_D_REG_10__SCAN_IN), .A3(
        P1_D_REG_11__SCAN_IN), .A4(P1_D_REG_12__SCAN_IN), .ZN(n6458) );
  NOR4_X1 U8094 ( .A1(P1_D_REG_4__SCAN_IN), .A2(P1_D_REG_5__SCAN_IN), .A3(
        P1_D_REG_6__SCAN_IN), .A4(P1_D_REG_7__SCAN_IN), .ZN(n6457) );
  NAND4_X1 U8095 ( .A1(n6460), .A2(n6459), .A3(n6458), .A4(n6457), .ZN(n6461)
         );
  NOR2_X1 U8096 ( .A1(n6462), .A2(n6461), .ZN(n6463) );
  OR2_X1 U8097 ( .A1(n9717), .A2(n6463), .ZN(n6753) );
  INV_X1 U8098 ( .A(n6753), .ZN(n6467) );
  OR2_X1 U8099 ( .A1(n9717), .A2(P1_D_REG_1__SCAN_IN), .ZN(n6466) );
  OR2_X1 U8100 ( .A1(n6468), .A2(n6464), .ZN(n6465) );
  NAND2_X1 U8101 ( .A1(n6466), .A2(n6465), .ZN(n6752) );
  NOR2_X1 U8102 ( .A1(n6467), .A2(n6752), .ZN(n7318) );
  OR2_X1 U8103 ( .A1(n9717), .A2(P1_D_REG_0__SCAN_IN), .ZN(n6471) );
  INV_X1 U8104 ( .A(n6468), .ZN(n7714) );
  INV_X1 U8105 ( .A(n6469), .ZN(n7476) );
  NAND2_X1 U8106 ( .A1(n7714), .A2(n7476), .ZN(n6470) );
  NAND4_X1 U8107 ( .A1(n6474), .A2(n6473), .A3(n6472), .A4(n5942), .ZN(n6475)
         );
  OAI21_X1 U8108 ( .B1(n6476), .B2(n6475), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n6478) );
  INV_X1 U8109 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n6477) );
  XNOR2_X1 U8110 ( .A(n6478), .B(n6477), .ZN(n7345) );
  NAND3_X1 U8111 ( .A1(n7345), .A2(P1_STATE_REG_SCAN_IN), .A3(n6506), .ZN(
        n9722) );
  INV_X1 U8112 ( .A(n9722), .ZN(n6751) );
  INV_X1 U8113 ( .A(n6479), .ZN(n6750) );
  INV_X1 U8114 ( .A(n6480), .ZN(n8939) );
  NOR2_X1 U8115 ( .A1(n9736), .A2(n8939), .ZN(n6481) );
  NAND2_X1 U8116 ( .A1(n8586), .A2(n8822), .ZN(n6483) );
  NAND2_X1 U8117 ( .A1(n6003), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n6482) );
  NAND2_X1 U8118 ( .A1(n9455), .A2(n4260), .ZN(n6496) );
  NAND2_X1 U8119 ( .A1(n6582), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n6494) );
  INV_X1 U8120 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n6484) );
  OR2_X1 U8121 ( .A1(n6116), .A2(n6484), .ZN(n6493) );
  INV_X1 U8122 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n6485) );
  OAI21_X1 U8123 ( .B1(n6486), .B2(n7864), .A(n6485), .ZN(n6489) );
  INV_X1 U8124 ( .A(n6486), .ZN(n6488) );
  AND2_X1 U8125 ( .A1(P1_REG3_REG_27__SCAN_IN), .A2(P1_REG3_REG_28__SCAN_IN), 
        .ZN(n6487) );
  NAND2_X1 U8126 ( .A1(n6488), .A2(n6487), .ZN(n9196) );
  NAND2_X1 U8127 ( .A1(n6489), .A2(n9196), .ZN(n7892) );
  INV_X1 U8128 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n6490) );
  OR2_X1 U8129 ( .A1(n6584), .A2(n6490), .ZN(n6491) );
  OR2_X1 U8130 ( .A1(n6397), .A2(n9189), .ZN(n6495) );
  NAND2_X1 U8131 ( .A1(n6496), .A2(n6495), .ZN(n6498) );
  XNOR2_X1 U8132 ( .A(n6498), .B(n6497), .ZN(n6501) );
  AOI22_X1 U8133 ( .A1(n9455), .A2(n6499), .B1(n4260), .B2(n9214), .ZN(n6500)
         );
  XNOR2_X1 U8134 ( .A(n6501), .B(n6500), .ZN(n6502) );
  INV_X1 U8135 ( .A(n6502), .ZN(n6532) );
  NAND3_X1 U8136 ( .A1(n6533), .A2(n8794), .A3(n6532), .ZN(n6538) );
  INV_X1 U8137 ( .A(n6521), .ZN(n6523) );
  OR2_X1 U8138 ( .A1(n9722), .A2(n9694), .ZN(n6505) );
  NAND2_X1 U8139 ( .A1(n6523), .A2(n9697), .ZN(n8656) );
  AND2_X1 U8140 ( .A1(n7345), .A2(n6506), .ZN(n6507) );
  OAI211_X1 U8141 ( .C1(n9736), .C2(n6509), .A(n6507), .B(n7319), .ZN(n6508)
         );
  NAND2_X1 U8142 ( .A1(n6508), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6512) );
  NOR2_X1 U8143 ( .A1(n6479), .A2(n8938), .ZN(n9693) );
  INV_X1 U8144 ( .A(n6509), .ZN(n6510) );
  NAND3_X1 U8145 ( .A1(n9693), .A2(n6751), .A3(n6510), .ZN(n6511) );
  INV_X1 U8146 ( .A(n6513), .ZN(n6514) );
  NAND2_X1 U8147 ( .A1(n6514), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6515) );
  NAND2_X1 U8148 ( .A1(n6516), .A2(n6515), .ZN(n6622) );
  INV_X1 U8149 ( .A(n6517), .ZN(n6518) );
  OR2_X1 U8150 ( .A1(n6622), .A2(n6518), .ZN(n6519) );
  XNOR2_X1 U8151 ( .A(n6519), .B(P1_IR_REG_28__SCAN_IN), .ZN(n9574) );
  NOR2_X1 U8152 ( .A1(n9101), .A2(n9574), .ZN(n6520) );
  NAND2_X1 U8153 ( .A1(n6521), .A2(n6520), .ZN(n8806) );
  INV_X1 U8154 ( .A(n8806), .ZN(n8748) );
  AOI22_X1 U8155 ( .A1(n8748), .A2(n9228), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3084), .ZN(n6531) );
  NOR2_X1 U8156 ( .A1(n6523), .A2(n6522), .ZN(n8771) );
  NAND2_X1 U8157 ( .A1(n6524), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n6529) );
  NAND2_X1 U8158 ( .A1(n6582), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n6528) );
  OR2_X1 U8159 ( .A1(n4264), .A2(n9196), .ZN(n6527) );
  INV_X1 U8160 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n6525) );
  OR2_X1 U8161 ( .A1(n6584), .A2(n6525), .ZN(n6526) );
  NAND4_X1 U8162 ( .A1(n6529), .A2(n6528), .A3(n6527), .A4(n6526), .ZN(n9105)
         );
  NAND2_X1 U8163 ( .A1(n8808), .A2(n9105), .ZN(n6530) );
  OAI211_X1 U8164 ( .C1(n7892), .C2(n8810), .A(n6531), .B(n6530), .ZN(n6535)
         );
  NOR3_X1 U8165 ( .A1(n6533), .A2(n6532), .A3(n8814), .ZN(n6534) );
  AOI211_X1 U8166 ( .C1(n8812), .C2(n9455), .A(n6535), .B(n6534), .ZN(n6536)
         );
  OAI211_X1 U8167 ( .C1(n7863), .C2(n6538), .A(n6537), .B(n6536), .ZN(P1_U3218) );
  OR2_X1 U8168 ( .A1(n6539), .A2(P2_U3152), .ZN(n6713) );
  INV_X2 U8169 ( .A(n8052), .ZN(P2_U3966) );
  NAND2_X1 U8170 ( .A1(n6541), .A2(n7345), .ZN(n6623) );
  INV_X2 U8171 ( .A(n9117), .ZN(P1_U4006) );
  XNOR2_X1 U8172 ( .A(n6543), .B(n6542), .ZN(n6544) );
  NOR2_X1 U8173 ( .A1(n6544), .A2(n8019), .ZN(n6551) );
  NOR2_X1 U8174 ( .A1(n8029), .A2(n4406), .ZN(n6550) );
  AND2_X1 U8175 ( .A1(n8042), .A2(n7691), .ZN(n6549) );
  INV_X1 U8176 ( .A(n7993), .ZN(n8056) );
  NAND2_X1 U8177 ( .A1(n8035), .A2(n8056), .ZN(n6547) );
  NOR2_X1 U8178 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6545), .ZN(n7547) );
  INV_X1 U8179 ( .A(n7547), .ZN(n6546) );
  OAI211_X1 U8180 ( .C1(n8039), .C2(n7435), .A(n6547), .B(n6546), .ZN(n6548)
         );
  OR4_X1 U8181 ( .A1(n6551), .A2(n6550), .A3(n6549), .A4(n6548), .ZN(P2_U3238)
         );
  XNOR2_X1 U8182 ( .A(n6552), .B(n6553), .ZN(n6554) );
  NOR2_X1 U8183 ( .A1(n6554), .A2(n8019), .ZN(n6559) );
  INV_X1 U8184 ( .A(n8546), .ZN(n7575) );
  NOR2_X1 U8185 ( .A1(n8029), .A2(n7575), .ZN(n6558) );
  AND2_X1 U8186 ( .A1(n8042), .A2(n7572), .ZN(n6557) );
  INV_X1 U8187 ( .A(n7627), .ZN(n8057) );
  NAND2_X1 U8188 ( .A1(n8035), .A2(n8057), .ZN(n6555) );
  NAND2_X1 U8189 ( .A1(P2_U3152), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n7465) );
  OAI211_X1 U8190 ( .C1(n8039), .C2(n7556), .A(n6555), .B(n7465), .ZN(n6556)
         );
  OR4_X1 U8191 ( .A1(n6559), .A2(n6558), .A3(n6557), .A4(n6556), .ZN(P2_U3219)
         );
  INV_X1 U8192 ( .A(n6806), .ZN(n6562) );
  INV_X1 U8193 ( .A(n6560), .ZN(n6599) );
  NOR2_X1 U8194 ( .A1(n6575), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8581) );
  INV_X1 U8195 ( .A(n8581), .ZN(n8587) );
  OAI222_X1 U8196 ( .A1(n6562), .A2(P2_U3152), .B1(n8583), .B2(n6599), .C1(
        n6561), .C2(n8587), .ZN(P2_U3356) );
  INV_X1 U8197 ( .A(n6563), .ZN(n6595) );
  AOI22_X1 U8198 ( .A1(n6832), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_4__SCAN_IN), .B2(n8581), .ZN(n6564) );
  OAI21_X1 U8199 ( .B1(n6595), .B2(n8583), .A(n6564), .ZN(P2_U3354) );
  INV_X1 U8200 ( .A(n6565), .ZN(n6590) );
  INV_X1 U8201 ( .A(n6767), .ZN(n6745) );
  OAI222_X1 U8202 ( .A1(n8587), .A2(n4544), .B1(n8583), .B2(n6590), .C1(
        P2_U3152), .C2(n6745), .ZN(P2_U3355) );
  INV_X1 U8203 ( .A(n6566), .ZN(n6597) );
  OAI222_X1 U8204 ( .A1(n6737), .A2(P2_U3152), .B1(n8583), .B2(n6597), .C1(
        n6567), .C2(n8587), .ZN(P2_U3357) );
  NAND2_X1 U8205 ( .A1(n6582), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n6572) );
  INV_X1 U8206 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n6568) );
  OR2_X1 U8207 ( .A1(n6116), .A2(n6568), .ZN(n6571) );
  INV_X1 U8208 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n6569) );
  OR2_X1 U8209 ( .A1(n6584), .A2(n6569), .ZN(n6570) );
  AND3_X1 U8210 ( .A1(n6572), .A2(n6571), .A3(n6570), .ZN(n9187) );
  NAND2_X1 U8211 ( .A1(n9117), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n6573) );
  OAI21_X1 U8212 ( .B1(n9187), .B2(n9117), .A(n6573), .ZN(P1_U3585) );
  INV_X1 U8213 ( .A(n6574), .ZN(n6577) );
  INV_X1 U8214 ( .A(n9576), .ZN(n9566) );
  AOI22_X1 U8215 ( .A1(n9134), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_5__SCAN_IN), .B2(n9566), .ZN(n6576) );
  OAI21_X1 U8216 ( .B1(n6577), .B2(n9572), .A(n6576), .ZN(P1_U3348) );
  INV_X1 U8217 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n6578) );
  INV_X1 U8218 ( .A(n6844), .ZN(n6779) );
  OAI222_X1 U8219 ( .A1(n8587), .A2(n6578), .B1(n8583), .B2(n6577), .C1(
        P2_U3152), .C2(n6779), .ZN(P2_U3353) );
  INV_X1 U8220 ( .A(n6579), .ZN(n6594) );
  AOI22_X1 U8221 ( .A1(n6908), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_6__SCAN_IN), .B2(n8581), .ZN(n6580) );
  OAI21_X1 U8222 ( .B1(n6594), .B2(n8583), .A(n6580), .ZN(P2_U3352) );
  INV_X1 U8223 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n9944) );
  NAND2_X1 U8224 ( .A1(P1_U4006), .A2(n7106), .ZN(n6581) );
  OAI21_X1 U8225 ( .B1(P1_U4006), .B2(n9944), .A(n6581), .ZN(P1_U3555) );
  NAND2_X1 U8226 ( .A1(n6582), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n6587) );
  INV_X1 U8227 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n9962) );
  OR2_X1 U8228 ( .A1(n6116), .A2(n9962), .ZN(n6586) );
  INV_X1 U8229 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n6583) );
  OR2_X1 U8230 ( .A1(n6584), .A2(n6583), .ZN(n6585) );
  AND3_X1 U8231 ( .A1(n6587), .A2(n6586), .A3(n6585), .ZN(n9173) );
  INV_X1 U8232 ( .A(n9173), .ZN(n8936) );
  NAND2_X1 U8233 ( .A1(n8936), .A2(P1_U4006), .ZN(n6588) );
  OAI21_X1 U8234 ( .B1(P1_U4006), .B2(n5545), .A(n6588), .ZN(P1_U3586) );
  INV_X1 U8235 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n6589) );
  INV_X1 U8236 ( .A(n6096), .ZN(n6592) );
  INV_X1 U8237 ( .A(n7043), .ZN(n7047) );
  OAI222_X1 U8238 ( .A1(n8587), .A2(n6589), .B1(n8583), .B2(n6592), .C1(
        P2_U3152), .C2(n7047), .ZN(P2_U3351) );
  INV_X1 U8239 ( .A(n6665), .ZN(n6819) );
  OAI222_X1 U8240 ( .A1(n6819), .A2(P1_U3084), .B1(n9572), .B2(n6590), .C1(
        n4692), .C2(n9576), .ZN(P1_U3350) );
  INV_X1 U8241 ( .A(n6671), .ZN(n6789) );
  INV_X1 U8242 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n6591) );
  OAI222_X1 U8243 ( .A1(n6789), .A2(P1_U3084), .B1(n9572), .B2(n6592), .C1(
        n6591), .C2(n9576), .ZN(P1_U3346) );
  INV_X1 U8244 ( .A(n6670), .ZN(n6691) );
  INV_X1 U8245 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n6593) );
  OAI222_X1 U8246 ( .A1(n6691), .A2(P1_U3084), .B1(n9572), .B2(n6594), .C1(
        n6593), .C2(n9576), .ZN(P1_U3347) );
  INV_X1 U8247 ( .A(n6658), .ZN(n6993) );
  OAI222_X1 U8248 ( .A1(n6993), .A2(P1_U3084), .B1(n9572), .B2(n6595), .C1(
        n4587), .C2(n9576), .ZN(P1_U3349) );
  INV_X1 U8249 ( .A(n6659), .ZN(n6636) );
  INV_X1 U8250 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n6596) );
  OAI222_X1 U8251 ( .A1(P1_U3084), .A2(n6636), .B1(n9572), .B2(n6597), .C1(
        n6596), .C2(n9576), .ZN(P1_U3352) );
  OAI222_X1 U8252 ( .A1(P1_U3084), .A2(n4362), .B1(n9572), .B2(n6599), .C1(
        n6598), .C2(n9576), .ZN(P1_U3351) );
  INV_X1 U8253 ( .A(n6600), .ZN(n6602) );
  OAI222_X1 U8254 ( .A1(n6701), .A2(P1_U3084), .B1(n9572), .B2(n6602), .C1(
        n6601), .C2(n9576), .ZN(P1_U3345) );
  INV_X1 U8255 ( .A(n7292), .ZN(n7287) );
  OAI222_X1 U8256 ( .A1(n8587), .A2(n6603), .B1(n8583), .B2(n6602), .C1(
        P2_U3152), .C2(n7287), .ZN(P2_U3350) );
  INV_X1 U8257 ( .A(n6604), .ZN(n6607) );
  INV_X1 U8258 ( .A(n7467), .ZN(n7290) );
  OAI222_X1 U8259 ( .A1(n8583), .A2(n6607), .B1(n7290), .B2(P2_U3152), .C1(
        n6605), .C2(n8587), .ZN(P2_U3349) );
  INV_X1 U8260 ( .A(n6859), .ZN(n6856) );
  OAI222_X1 U8261 ( .A1(P1_U3084), .A2(n6856), .B1(n9572), .B2(n6607), .C1(
        n6606), .C2(n9576), .ZN(P1_U3344) );
  INV_X1 U8262 ( .A(n6608), .ZN(n6613) );
  AOI22_X1 U8263 ( .A1(n7006), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_11__SCAN_IN), .B2(n9566), .ZN(n6609) );
  OAI21_X1 U8264 ( .B1(n6613), .B2(n9572), .A(n6609), .ZN(P1_U3342) );
  INV_X1 U8265 ( .A(n6610), .ZN(n6615) );
  INV_X1 U8266 ( .A(n7541), .ZN(n7537) );
  OAI222_X1 U8267 ( .A1(n8583), .A2(n6615), .B1(n7537), .B2(P2_U3152), .C1(
        n6611), .C2(n8587), .ZN(P2_U3348) );
  INV_X1 U8268 ( .A(n7764), .ZN(n7545) );
  OAI222_X1 U8269 ( .A1(n8583), .A2(n6613), .B1(n7545), .B2(P2_U3152), .C1(
        n6612), .C2(n8587), .ZN(P2_U3347) );
  INV_X1 U8270 ( .A(n6880), .ZN(n6857) );
  OAI222_X1 U8271 ( .A1(P1_U3084), .A2(n6857), .B1(n9572), .B2(n6615), .C1(
        n6614), .C2(n9576), .ZN(P1_U3343) );
  OAI21_X1 U8272 ( .B1(n9801), .B2(n7019), .A(n6722), .ZN(n6617) );
  NAND2_X1 U8273 ( .A1(n9801), .A2(n6712), .ZN(n6616) );
  NAND2_X1 U8274 ( .A1(n6617), .A2(n6616), .ZN(n8171) );
  NOR2_X1 U8275 ( .A1(n8088), .A2(P2_U3966), .ZN(P2_U3151) );
  INV_X1 U8276 ( .A(n7345), .ZN(n6618) );
  OR2_X1 U8277 ( .A1(n6480), .A2(n6618), .ZN(n6619) );
  NAND2_X1 U8278 ( .A1(n6619), .A2(n6623), .ZN(n6643) );
  OR2_X1 U8279 ( .A1(n6643), .A2(n6620), .ZN(n6621) );
  NAND2_X1 U8280 ( .A1(n6621), .A2(P1_STATE_REG_SCAN_IN), .ZN(P1_U3083) );
  XNOR2_X1 U8281 ( .A(n6622), .B(P1_IR_REG_27__SCAN_IN), .ZN(n9172) );
  NOR2_X1 U8282 ( .A1(n6625), .A2(n9172), .ZN(n9164) );
  INV_X1 U8283 ( .A(P1_U3083), .ZN(n6624) );
  NAND2_X1 U8284 ( .A1(n6624), .A2(n6623), .ZN(n9662) );
  INV_X1 U8285 ( .A(n9662), .ZN(n9171) );
  INV_X1 U8286 ( .A(n6625), .ZN(n6627) );
  INV_X1 U8287 ( .A(n9172), .ZN(n6977) );
  NOR2_X1 U8288 ( .A1(n6977), .A2(n9574), .ZN(n6626) );
  NAND2_X1 U8289 ( .A1(n6627), .A2(n6626), .ZN(n9163) );
  MUX2_X1 U8290 ( .A(P1_REG1_REG_1__SCAN_IN), .B(n5979), .S(n6659), .Z(n6629)
         );
  AND2_X1 U8291 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(
        n6628) );
  NAND2_X1 U8292 ( .A1(n6629), .A2(n6628), .ZN(n6661) );
  OAI21_X1 U8293 ( .B1(n6629), .B2(n6628), .A(n6661), .ZN(n6630) );
  OAI22_X1 U8294 ( .A1(n9163), .A2(n6630), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9698), .ZN(n6631) );
  AOI21_X1 U8295 ( .B1(n9171), .B2(P1_ADDR_REG_1__SCAN_IN), .A(n6631), .ZN(
        n6635) );
  INV_X1 U8296 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n9715) );
  MUX2_X1 U8297 ( .A(P1_REG2_REG_1__SCAN_IN), .B(n9715), .S(n6659), .Z(n6633)
         );
  AND2_X1 U8298 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(
        n6632) );
  INV_X1 U8299 ( .A(n9574), .ZN(n6895) );
  NAND2_X1 U8300 ( .A1(n9164), .A2(n6895), .ZN(n9620) );
  NAND2_X1 U8301 ( .A1(n6633), .A2(n6632), .ZN(n6649) );
  OAI211_X1 U8302 ( .C1(n6633), .C2(n6632), .A(n9648), .B(n6649), .ZN(n6634)
         );
  OAI211_X1 U8303 ( .C1(n9654), .C2(n6636), .A(n6635), .B(n6634), .ZN(P1_U3242) );
  INV_X1 U8304 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n6647) );
  AOI21_X1 U8305 ( .B1(n9172), .B2(n6637), .A(P1_IR_REG_0__SCAN_IN), .ZN(n6639) );
  NOR2_X1 U8306 ( .A1(n9172), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n6638) );
  NOR2_X1 U8307 ( .A1(n6638), .A2(n9574), .ZN(n6980) );
  MUX2_X1 U8308 ( .A(P1_IR_REG_0__SCAN_IN), .B(n6639), .S(n6980), .Z(n6641) );
  NAND3_X1 U8309 ( .A1(n6641), .A2(P1_STATE_REG_SCAN_IN), .A3(n6640), .ZN(
        n6642) );
  NOR2_X1 U8310 ( .A1(n6643), .A2(n6642), .ZN(n6645) );
  NOR3_X1 U8311 ( .A1(n9163), .A2(P1_REG1_REG_0__SCAN_IN), .A3(n6978), .ZN(
        n6644) );
  AOI211_X1 U8312 ( .C1(P1_REG3_REG_0__SCAN_IN), .C2(P1_U3084), .A(n6645), .B(
        n6644), .ZN(n6646) );
  OAI21_X1 U8313 ( .B1(n9662), .B2(n6647), .A(n6646), .ZN(P1_U3241) );
  XNOR2_X1 U8314 ( .A(n6701), .B(P1_REG2_REG_8__SCAN_IN), .ZN(n6699) );
  MUX2_X1 U8315 ( .A(n6652), .B(P1_REG2_REG_4__SCAN_IN), .S(n6658), .Z(n6991)
         );
  NAND2_X1 U8316 ( .A1(n6659), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n6648) );
  NAND2_X1 U8317 ( .A1(n6649), .A2(n6648), .ZN(n9126) );
  INV_X1 U8318 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n7324) );
  NAND2_X1 U8319 ( .A1(n9126), .A2(n9127), .ZN(n9125) );
  NAND2_X1 U8320 ( .A1(n9124), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n6650) );
  NAND2_X1 U8321 ( .A1(n9125), .A2(n6650), .ZN(n6815) );
  INV_X1 U8322 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n7483) );
  XNOR2_X1 U8323 ( .A(n6665), .B(n7483), .ZN(n6816) );
  NAND2_X1 U8324 ( .A1(n6815), .A2(n6816), .ZN(n6814) );
  NAND2_X1 U8325 ( .A1(n6665), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n6651) );
  NAND2_X1 U8326 ( .A1(n6814), .A2(n6651), .ZN(n6990) );
  NAND2_X1 U8327 ( .A1(n6993), .A2(n6652), .ZN(n6653) );
  XNOR2_X1 U8328 ( .A(n9134), .B(n6654), .ZN(n9132) );
  NOR2_X1 U8329 ( .A1(n9134), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n6655) );
  AOI21_X1 U8330 ( .B1(n9133), .B2(n9132), .A(n6655), .ZN(n6687) );
  INV_X1 U8331 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n7391) );
  XNOR2_X1 U8332 ( .A(n6670), .B(n7391), .ZN(n6688) );
  NAND2_X1 U8333 ( .A1(n6687), .A2(n6688), .ZN(n6686) );
  NAND2_X1 U8334 ( .A1(n6670), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n6656) );
  NAND2_X1 U8335 ( .A1(n6686), .A2(n6656), .ZN(n6786) );
  XNOR2_X1 U8336 ( .A(n6671), .B(P1_REG2_REG_7__SCAN_IN), .ZN(n6787) );
  OR2_X1 U8337 ( .A1(n6671), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n6657) );
  XOR2_X1 U8338 ( .A(n6699), .B(n6700), .Z(n6680) );
  NAND2_X1 U8339 ( .A1(P1_U3084), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n7614) );
  OAI21_X1 U8340 ( .B1(n9662), .B2(n4374), .A(n7614), .ZN(n6677) );
  MUX2_X1 U8341 ( .A(P1_REG1_REG_8__SCAN_IN), .B(n6695), .S(n6701), .Z(n6674)
         );
  MUX2_X1 U8342 ( .A(n6667), .B(P1_REG1_REG_4__SCAN_IN), .S(n6658), .Z(n6983)
         );
  NAND2_X1 U8343 ( .A1(n6659), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n6660) );
  NAND2_X1 U8344 ( .A1(n6661), .A2(n6660), .ZN(n9119) );
  XNOR2_X1 U8345 ( .A(n9124), .B(n6662), .ZN(n9120) );
  NAND2_X1 U8346 ( .A1(n9119), .A2(n9120), .ZN(n9118) );
  NAND2_X1 U8347 ( .A1(n9124), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n6663) );
  NAND2_X1 U8348 ( .A1(n9118), .A2(n6663), .ZN(n6809) );
  XNOR2_X1 U8349 ( .A(n6665), .B(n6664), .ZN(n6810) );
  NAND2_X1 U8350 ( .A1(n6809), .A2(n6810), .ZN(n6808) );
  NAND2_X1 U8351 ( .A1(n6665), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n6666) );
  NAND2_X1 U8352 ( .A1(n6993), .A2(n6667), .ZN(n6668) );
  XNOR2_X1 U8353 ( .A(n9134), .B(P1_REG1_REG_5__SCAN_IN), .ZN(n9136) );
  AOI21_X1 U8354 ( .B1(n9134), .B2(P1_REG1_REG_5__SCAN_IN), .A(n9139), .ZN(
        n6682) );
  XNOR2_X1 U8355 ( .A(n6670), .B(n6669), .ZN(n6683) );
  NAND2_X1 U8356 ( .A1(n6682), .A2(n6683), .ZN(n6681) );
  OAI21_X1 U8357 ( .B1(P1_REG1_REG_6__SCAN_IN), .B2(n6670), .A(n6681), .ZN(
        n6782) );
  XNOR2_X1 U8358 ( .A(n6671), .B(n6672), .ZN(n6783) );
  AOI22_X1 U8359 ( .A1(n6782), .A2(n6783), .B1(n6672), .B2(n6789), .ZN(n6673)
         );
  NOR2_X1 U8360 ( .A1(n6673), .A2(n6674), .ZN(n6694) );
  AOI21_X1 U8361 ( .B1(n6674), .B2(n6673), .A(n6694), .ZN(n6675) );
  NOR2_X1 U8362 ( .A1(n6675), .A2(n9163), .ZN(n6676) );
  AOI211_X1 U8363 ( .C1(n9627), .C2(n6678), .A(n6677), .B(n6676), .ZN(n6679)
         );
  OAI21_X1 U8364 ( .B1(n9620), .B2(n6680), .A(n6679), .ZN(P1_U3249) );
  OAI21_X1 U8365 ( .B1(n6683), .B2(n6682), .A(n6681), .ZN(n6685) );
  AND2_X1 U8366 ( .A1(P1_U3084), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n7336) );
  NOR2_X1 U8367 ( .A1(n9662), .A2(n4375), .ZN(n6684) );
  AOI211_X1 U8368 ( .C1(n9659), .C2(n6685), .A(n7336), .B(n6684), .ZN(n6690)
         );
  OAI211_X1 U8369 ( .C1(n6688), .C2(n6687), .A(n9648), .B(n6686), .ZN(n6689)
         );
  OAI211_X1 U8370 ( .C1(n9654), .C2(n6691), .A(n6690), .B(n6689), .ZN(P1_U3247) );
  INV_X1 U8371 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n6693) );
  NAND2_X1 U8372 ( .A1(P2_U3966), .A2(n8174), .ZN(n6692) );
  OAI21_X1 U8373 ( .B1(P2_U3966), .B2(n6693), .A(n6692), .ZN(P2_U3583) );
  MUX2_X1 U8374 ( .A(n6855), .B(P1_REG1_REG_9__SCAN_IN), .S(n6859), .Z(n6697)
         );
  AOI21_X1 U8375 ( .B1(n6695), .B2(n6701), .A(n6694), .ZN(n6696) );
  NOR2_X1 U8376 ( .A1(n6696), .A2(n6697), .ZN(n6854) );
  AOI21_X1 U8377 ( .B1(n6697), .B2(n6696), .A(n6854), .ZN(n6710) );
  INV_X1 U8378 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n10065) );
  AND2_X1 U8379 ( .A1(P1_U3084), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n8716) );
  INV_X1 U8380 ( .A(n8716), .ZN(n6698) );
  OAI21_X1 U8381 ( .B1(n9662), .B2(n10065), .A(n6698), .ZN(n6708) );
  XNOR2_X1 U8382 ( .A(n6859), .B(P1_REG2_REG_9__SCAN_IN), .ZN(n6706) );
  NAND2_X1 U8383 ( .A1(n6700), .A2(n6699), .ZN(n6703) );
  NAND2_X1 U8384 ( .A1(n6701), .A2(n7589), .ZN(n6702) );
  NAND2_X1 U8385 ( .A1(n6703), .A2(n6702), .ZN(n6705) );
  INV_X1 U8386 ( .A(n6861), .ZN(n6704) );
  AOI211_X1 U8387 ( .C1(n6706), .C2(n6705), .A(n6704), .B(n9620), .ZN(n6707)
         );
  AOI211_X1 U8388 ( .C1(n9627), .C2(n6859), .A(n6708), .B(n6707), .ZN(n6709)
         );
  OAI21_X1 U8389 ( .B1(n6710), .B2(n9163), .A(n6709), .ZN(P1_U3250) );
  NAND2_X1 U8390 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), 
        .ZN(n6718) );
  INV_X1 U8391 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n6711) );
  INV_X1 U8392 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n9797) );
  AND2_X1 U8393 ( .A1(n6713), .A2(n6712), .ZN(n6714) );
  NAND2_X1 U8394 ( .A1(n6714), .A2(n7015), .ZN(n6724) );
  NAND2_X1 U8395 ( .A1(n6724), .A2(n6722), .ZN(n6715) );
  NAND2_X1 U8396 ( .A1(n8052), .A2(n6715), .ZN(n6720) );
  AND2_X1 U8397 ( .A1(n6719), .A2(n7844), .ZN(n6716) );
  NAND2_X1 U8398 ( .A1(n6720), .A2(n6716), .ZN(n8163) );
  AOI211_X1 U8399 ( .C1(n6718), .C2(n6717), .A(n6731), .B(n8163), .ZN(n6730)
         );
  INV_X1 U8400 ( .A(n6719), .ZN(n8589) );
  AOI22_X1 U8401 ( .A1(n8088), .A2(P2_ADDR_REG_1__SCAN_IN), .B1(
        P2_REG3_REG_1__SCAN_IN), .B2(P2_U3152), .ZN(n6728) );
  AND2_X1 U8402 ( .A1(P2_REG1_REG_0__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n6726) );
  INV_X1 U8403 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n6721) );
  INV_X1 U8404 ( .A(n7844), .ZN(n7819) );
  AND2_X1 U8405 ( .A1(n7819), .A2(n6722), .ZN(n6723) );
  NAND2_X1 U8406 ( .A1(n6725), .A2(n6726), .ZN(n6736) );
  OAI211_X1 U8407 ( .C1(n6726), .C2(n6725), .A(n8167), .B(n6736), .ZN(n6727)
         );
  OAI211_X1 U8408 ( .C1(n8165), .C2(n6737), .A(n6728), .B(n6727), .ZN(n6729)
         );
  OR2_X1 U8409 ( .A1(n6730), .A2(n6729), .ZN(P2_U3246) );
  XNOR2_X1 U8410 ( .A(n6806), .B(P2_REG2_REG_2__SCAN_IN), .ZN(n6802) );
  XNOR2_X1 U8411 ( .A(n6767), .B(P2_REG2_REG_3__SCAN_IN), .ZN(n6733) );
  AOI211_X1 U8412 ( .C1(n6734), .C2(n6733), .A(n6762), .B(n8163), .ZN(n6747)
         );
  AOI22_X1 U8413 ( .A1(n8088), .A2(P2_ADDR_REG_3__SCAN_IN), .B1(
        P2_REG3_REG_3__SCAN_IN), .B2(P2_U3152), .ZN(n6744) );
  INV_X1 U8414 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n6735) );
  MUX2_X1 U8415 ( .A(P2_REG1_REG_3__SCAN_IN), .B(n6735), .S(n6767), .Z(n6742)
         );
  OAI21_X1 U8416 ( .B1(n6721), .B2(n6737), .A(n6736), .ZN(n6798) );
  INV_X1 U8417 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n6738) );
  XNOR2_X1 U8418 ( .A(n6806), .B(n6738), .ZN(n6797) );
  NAND2_X1 U8419 ( .A1(n6798), .A2(n6797), .ZN(n6740) );
  NAND2_X1 U8420 ( .A1(n6806), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n6739) );
  NAND2_X1 U8421 ( .A1(n6740), .A2(n6739), .ZN(n6741) );
  NAND2_X1 U8422 ( .A1(n6741), .A2(n6742), .ZN(n6822) );
  OAI211_X1 U8423 ( .C1(n6742), .C2(n6741), .A(n8167), .B(n6822), .ZN(n6743)
         );
  OAI211_X1 U8424 ( .C1(n8165), .C2(n6745), .A(n6744), .B(n6743), .ZN(n6746)
         );
  OR2_X1 U8425 ( .A1(n6747), .A2(n6746), .ZN(P2_U3248) );
  INV_X1 U8426 ( .A(n9398), .ZN(n9702) );
  NOR2_X2 U8427 ( .A1(n7106), .A2(n9690), .ZN(n9699) );
  NAND2_X1 U8428 ( .A1(n7106), .A2(n9690), .ZN(n8986) );
  INV_X1 U8429 ( .A(n8986), .ZN(n6748) );
  OR2_X1 U8430 ( .A1(n9699), .A2(n6748), .ZN(n9059) );
  NAND3_X1 U8431 ( .A1(n9101), .A2(n9059), .A3(n6479), .ZN(n6749) );
  OAI21_X1 U8432 ( .B1(n9702), .B2(n8770), .A(n6749), .ZN(n7459) );
  AOI21_X1 U8433 ( .B1(n7458), .B2(n6750), .A(n7459), .ZN(n6920) );
  AND2_X1 U8434 ( .A1(n6752), .A2(n6751), .ZN(n9721) );
  AND2_X1 U8435 ( .A1(n9721), .A2(n6753), .ZN(n6754) );
  AND2_X1 U8436 ( .A1(n7319), .A2(n6754), .ZN(n6756) );
  OR2_X1 U8437 ( .A1(n9754), .A2(n9694), .ZN(n6755) );
  NAND2_X1 U8438 ( .A1(n9783), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n6757) );
  OAI21_X1 U8439 ( .B1(n6920), .B2(n9783), .A(n6757), .ZN(P1_U3523) );
  INV_X1 U8440 ( .A(n7237), .ZN(n6998) );
  INV_X1 U8441 ( .A(n6758), .ZN(n6760) );
  OAI222_X1 U8442 ( .A1(n6998), .A2(P1_U3084), .B1(n9572), .B2(n6760), .C1(
        n6759), .C2(n9576), .ZN(P1_U3341) );
  INV_X1 U8443 ( .A(n7793), .ZN(n7762) );
  OAI222_X1 U8444 ( .A1(n8587), .A2(n6761), .B1(n8583), .B2(n6760), .C1(
        P2_U3152), .C2(n7762), .ZN(P2_U3346) );
  INV_X1 U8445 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n6763) );
  MUX2_X1 U8446 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n6763), .S(n6832), .Z(n6764)
         );
  INV_X1 U8447 ( .A(n6764), .ZN(n6828) );
  XNOR2_X1 U8448 ( .A(n6844), .B(P2_REG2_REG_5__SCAN_IN), .ZN(n6765) );
  AOI211_X1 U8449 ( .C1(n6766), .C2(n6765), .A(n8163), .B(n6843), .ZN(n6781)
         );
  AND2_X1 U8450 ( .A1(P2_REG3_REG_5__SCAN_IN), .A2(P2_U3152), .ZN(n7090) );
  AOI21_X1 U8451 ( .B1(n8088), .B2(P2_ADDR_REG_5__SCAN_IN), .A(n7090), .ZN(
        n6778) );
  NAND2_X1 U8452 ( .A1(n6767), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n6821) );
  NAND2_X1 U8453 ( .A1(n6822), .A2(n6821), .ZN(n6770) );
  INV_X1 U8454 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n6768) );
  MUX2_X1 U8455 ( .A(P2_REG1_REG_4__SCAN_IN), .B(n6768), .S(n6832), .Z(n6769)
         );
  NAND2_X1 U8456 ( .A1(n6770), .A2(n6769), .ZN(n6824) );
  NAND2_X1 U8457 ( .A1(n6832), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n6775) );
  NAND2_X1 U8458 ( .A1(n6824), .A2(n6775), .ZN(n6773) );
  INV_X1 U8459 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n6771) );
  MUX2_X1 U8460 ( .A(P2_REG1_REG_5__SCAN_IN), .B(n6771), .S(n6844), .Z(n6772)
         );
  MUX2_X1 U8461 ( .A(n6771), .B(P2_REG1_REG_5__SCAN_IN), .S(n6844), .Z(n6774)
         );
  NAND3_X1 U8462 ( .A1(n6824), .A2(n6775), .A3(n6774), .ZN(n6776) );
  NAND3_X1 U8463 ( .A1(n8167), .A2(n6839), .A3(n6776), .ZN(n6777) );
  OAI211_X1 U8464 ( .C1(n8165), .C2(n6779), .A(n6778), .B(n6777), .ZN(n6780)
         );
  OR2_X1 U8465 ( .A1(n6781), .A2(n6780), .ZN(P2_U3250) );
  XOR2_X1 U8466 ( .A(n6783), .B(n6782), .Z(n6792) );
  AND2_X1 U8467 ( .A1(P1_U3084), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n7497) );
  INV_X1 U8468 ( .A(n6784), .ZN(n6785) );
  AOI21_X1 U8469 ( .B1(n6787), .B2(n6786), .A(n6785), .ZN(n6788) );
  OAI22_X1 U8470 ( .A1(n9654), .A2(n6789), .B1(n6788), .B2(n9620), .ZN(n6790)
         );
  AOI211_X1 U8471 ( .C1(n9171), .C2(P1_ADDR_REG_7__SCAN_IN), .A(n7497), .B(
        n6790), .ZN(n6791) );
  OAI21_X1 U8472 ( .B1(n9163), .B2(n6792), .A(n6791), .ZN(P1_U3248) );
  INV_X1 U8473 ( .A(n6793), .ZN(n6851) );
  AOI22_X1 U8474 ( .A1(n7270), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n9566), .ZN(n6794) );
  OAI21_X1 U8475 ( .B1(n6851), .B2(n9572), .A(n6794), .ZN(P1_U3340) );
  INV_X1 U8476 ( .A(n6795), .ZN(n6853) );
  INV_X1 U8477 ( .A(n8084), .ZN(n8091) );
  OAI222_X1 U8478 ( .A1(n8583), .A2(n6853), .B1(n8091), .B2(P2_U3152), .C1(
        n6796), .C2(n8587), .ZN(P2_U3344) );
  INV_X1 U8479 ( .A(n8167), .ZN(n8117) );
  XNOR2_X1 U8480 ( .A(n6798), .B(n6797), .ZN(n6800) );
  AOI22_X1 U8481 ( .A1(n8088), .A2(P2_ADDR_REG_2__SCAN_IN), .B1(
        P2_REG3_REG_2__SCAN_IN), .B2(P2_U3152), .ZN(n6799) );
  OAI21_X1 U8482 ( .B1(n8117), .B2(n6800), .A(n6799), .ZN(n6805) );
  AOI211_X1 U8483 ( .C1(n6803), .C2(n6802), .A(n6801), .B(n8163), .ZN(n6804)
         );
  AOI211_X1 U8484 ( .C1(n8164), .C2(n6806), .A(n6805), .B(n6804), .ZN(n6807)
         );
  INV_X1 U8485 ( .A(n6807), .ZN(P2_U3247) );
  NAND2_X1 U8486 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_U3084), .ZN(n7201) );
  INV_X1 U8487 ( .A(n7201), .ZN(n6813) );
  OAI211_X1 U8488 ( .C1(n6810), .C2(n6809), .A(n9659), .B(n6808), .ZN(n6811)
         );
  INV_X1 U8489 ( .A(n6811), .ZN(n6812) );
  AOI211_X1 U8490 ( .C1(P1_ADDR_REG_3__SCAN_IN), .C2(n9171), .A(n6813), .B(
        n6812), .ZN(n6818) );
  OAI211_X1 U8491 ( .C1(n6816), .C2(n6815), .A(n9648), .B(n6814), .ZN(n6817)
         );
  OAI211_X1 U8492 ( .C1(n9654), .C2(n6819), .A(n6818), .B(n6817), .ZN(P1_U3244) );
  INV_X1 U8493 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n6826) );
  MUX2_X1 U8494 ( .A(n6768), .B(P2_REG1_REG_4__SCAN_IN), .S(n6832), .Z(n6820)
         );
  NAND3_X1 U8495 ( .A1(n6822), .A2(n6821), .A3(n6820), .ZN(n6823) );
  NAND3_X1 U8496 ( .A1(n8167), .A2(n6824), .A3(n6823), .ZN(n6825) );
  NAND2_X1 U8497 ( .A1(P2_U3152), .A2(P2_REG3_REG_4__SCAN_IN), .ZN(n6959) );
  OAI211_X1 U8498 ( .C1(n8171), .C2(n6826), .A(n6825), .B(n6959), .ZN(n6831)
         );
  AOI211_X1 U8499 ( .C1(n6829), .C2(n6828), .A(n8163), .B(n6827), .ZN(n6830)
         );
  AOI211_X1 U8500 ( .C1(n8164), .C2(n6832), .A(n6831), .B(n6830), .ZN(n6833)
         );
  INV_X1 U8501 ( .A(n6833), .ZN(P2_U3249) );
  INV_X1 U8502 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n6842) );
  NAND2_X1 U8503 ( .A1(n6844), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n6838) );
  NAND2_X1 U8504 ( .A1(n6839), .A2(n6838), .ZN(n6836) );
  INV_X1 U8505 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n6834) );
  MUX2_X1 U8506 ( .A(P2_REG1_REG_6__SCAN_IN), .B(n6834), .S(n6908), .Z(n6835)
         );
  NAND2_X1 U8507 ( .A1(n6836), .A2(n6835), .ZN(n6911) );
  MUX2_X1 U8508 ( .A(n6834), .B(P2_REG1_REG_6__SCAN_IN), .S(n6908), .Z(n6837)
         );
  NAND3_X1 U8509 ( .A1(n6839), .A2(n6838), .A3(n6837), .ZN(n6840) );
  NAND3_X1 U8510 ( .A1(n8167), .A2(n6911), .A3(n6840), .ZN(n6841) );
  NAND2_X1 U8511 ( .A1(P2_U3152), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n7156) );
  OAI211_X1 U8512 ( .C1(n8171), .C2(n6842), .A(n6841), .B(n7156), .ZN(n6848)
         );
  XNOR2_X1 U8513 ( .A(n6908), .B(P2_REG2_REG_6__SCAN_IN), .ZN(n6845) );
  AOI211_X1 U8514 ( .C1(n6846), .C2(n6845), .A(n8163), .B(n6904), .ZN(n6847)
         );
  AOI211_X1 U8515 ( .C1(n8164), .C2(n6908), .A(n6848), .B(n6847), .ZN(n6849)
         );
  INV_X1 U8516 ( .A(n6849), .ZN(P2_U3251) );
  INV_X1 U8517 ( .A(n8072), .ZN(n7803) );
  OAI222_X1 U8518 ( .A1(n8583), .A2(n6851), .B1(n7803), .B2(P2_U3152), .C1(
        n6850), .C2(n8587), .ZN(P2_U3345) );
  OAI222_X1 U8519 ( .A1(P1_U3084), .A2(n4420), .B1(n9572), .B2(n6853), .C1(
        n6852), .C2(n9576), .ZN(P1_U3339) );
  XNOR2_X1 U8520 ( .A(n6880), .B(P1_REG1_REG_10__SCAN_IN), .ZN(n6876) );
  AOI21_X1 U8521 ( .B1(n6856), .B2(n6855), .A(n6854), .ZN(n6877) );
  XOR2_X1 U8522 ( .A(n6876), .B(n6877), .Z(n6866) );
  AND2_X1 U8523 ( .A1(P1_U3084), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n8626) );
  NOR2_X1 U8524 ( .A1(n9654), .A2(n6857), .ZN(n6858) );
  AOI211_X1 U8525 ( .C1(n9171), .C2(P1_ADDR_REG_10__SCAN_IN), .A(n8626), .B(
        n6858), .ZN(n6865) );
  INV_X1 U8526 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n7522) );
  XNOR2_X1 U8527 ( .A(n6880), .B(n7522), .ZN(n6863) );
  NAND2_X1 U8528 ( .A1(n6859), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n6860) );
  NAND2_X1 U8529 ( .A1(n6861), .A2(n6860), .ZN(n6862) );
  NAND2_X1 U8530 ( .A1(n6862), .A2(n6863), .ZN(n6882) );
  OAI211_X1 U8531 ( .C1(n6863), .C2(n6862), .A(n6882), .B(n9648), .ZN(n6864)
         );
  OAI211_X1 U8532 ( .C1(n6866), .C2(n9163), .A(n6865), .B(n6864), .ZN(P1_U3251) );
  NOR2_X1 U8533 ( .A1(n6867), .A2(P2_U3152), .ZN(n6951) );
  INV_X1 U8534 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n6875) );
  NOR2_X1 U8535 ( .A1(n6868), .A2(n8404), .ZN(n9788) );
  NOR2_X1 U8536 ( .A1(n8029), .A2(n9791), .ZN(n6873) );
  MUX2_X1 U8537 ( .A(n6870), .B(n9791), .S(n6869), .Z(n6871) );
  AOI21_X1 U8538 ( .B1(n7165), .B2(n6871), .A(n8019), .ZN(n6872) );
  AOI211_X1 U8539 ( .C1(n7961), .C2(n9788), .A(n6873), .B(n6872), .ZN(n6874)
         );
  OAI21_X1 U8540 ( .B1(n6951), .B2(n6875), .A(n6874), .ZN(P2_U3234) );
  OAI22_X1 U8541 ( .A1(n6877), .A2(n6876), .B1(P1_REG1_REG_10__SCAN_IN), .B2(
        n6880), .ZN(n7001) );
  NOR2_X1 U8542 ( .A1(n7006), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n7000) );
  NAND2_X1 U8543 ( .A1(n7006), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n6999) );
  NAND2_X1 U8544 ( .A1(n4597), .A2(n6999), .ZN(n6878) );
  XNOR2_X1 U8545 ( .A(n7001), .B(n6878), .ZN(n6889) );
  INV_X1 U8546 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n6879) );
  NAND2_X1 U8547 ( .A1(P1_U3084), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n8759) );
  OAI21_X1 U8548 ( .B1(n9662), .B2(n6879), .A(n8759), .ZN(n6887) );
  NAND2_X1 U8549 ( .A1(n6880), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n6881) );
  NAND2_X1 U8550 ( .A1(n6882), .A2(n6881), .ZN(n6884) );
  XNOR2_X1 U8551 ( .A(n7006), .B(P1_REG2_REG_11__SCAN_IN), .ZN(n6883) );
  NAND2_X1 U8552 ( .A1(n6884), .A2(n6883), .ZN(n6885) );
  AOI21_X1 U8553 ( .B1(n7008), .B2(n6885), .A(n9620), .ZN(n6886) );
  AOI211_X1 U8554 ( .C1(n9627), .C2(n7006), .A(n6887), .B(n6886), .ZN(n6888)
         );
  OAI21_X1 U8555 ( .B1(n6889), .B2(n9163), .A(n6888), .ZN(P1_U3252) );
  NAND2_X1 U8556 ( .A1(n5975), .A2(n9169), .ZN(n8925) );
  OR2_X1 U8557 ( .A1(n8925), .A2(n6504), .ZN(n9740) );
  XNOR2_X2 U8558 ( .A(n6890), .B(n9724), .ZN(n6896) );
  NAND2_X1 U8559 ( .A1(n7106), .A2(n7458), .ZN(n9688) );
  NAND2_X1 U8560 ( .A1(n6896), .A2(n9688), .ZN(n6892) );
  NAND2_X1 U8561 ( .A1(n6892), .A2(n6891), .ZN(n7348) );
  XNOR2_X1 U8562 ( .A(n7348), .B(n9058), .ZN(n7329) );
  NAND2_X1 U8563 ( .A1(n9724), .A2(n9690), .ZN(n9689) );
  OAI21_X1 U8564 ( .B1(n4261), .B2(n6894), .A(n7484), .ZN(n7327) );
  OAI22_X1 U8565 ( .A1(n9768), .A2(n6894), .B1(n7327), .B2(n9754), .ZN(n6902)
         );
  INV_X1 U8566 ( .A(n9699), .ZN(n6897) );
  OR2_X1 U8567 ( .A1(n6890), .A2(n9724), .ZN(n6898) );
  XNOR2_X1 U8568 ( .A(n7365), .B(n9058), .ZN(n6901) );
  NAND2_X1 U8569 ( .A1(n6899), .A2(n9169), .ZN(n6900) );
  OR2_X1 U8570 ( .A1(n9091), .A2(n8938), .ZN(n8937) );
  OAI222_X1 U8571 ( .A1(n9703), .A2(n8770), .B1(n9702), .B2(n9677), .C1(n6901), 
        .C2(n9416), .ZN(n7321) );
  AOI211_X1 U8572 ( .C1(n9759), .C2(n7329), .A(n6902), .B(n7321), .ZN(n9728)
         );
  NAND2_X1 U8573 ( .A1(n9783), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n6903) );
  OAI21_X1 U8574 ( .B1(n9728), .B2(n9783), .A(n6903), .ZN(P1_U3525) );
  XNOR2_X1 U8575 ( .A(n7043), .B(P2_REG2_REG_7__SCAN_IN), .ZN(n6905) );
  AOI211_X1 U8576 ( .C1(n6906), .C2(n6905), .A(n8163), .B(n7042), .ZN(n6907)
         );
  INV_X1 U8577 ( .A(n6907), .ZN(n6916) );
  NOR2_X1 U8578 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n5115), .ZN(n6914) );
  NAND2_X1 U8579 ( .A1(n6908), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n6910) );
  INV_X1 U8580 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n9868) );
  MUX2_X1 U8581 ( .A(n9868), .B(P2_REG1_REG_7__SCAN_IN), .S(n7043), .Z(n6909)
         );
  AOI21_X1 U8582 ( .B1(n6911), .B2(n6910), .A(n6909), .ZN(n7053) );
  AND3_X1 U8583 ( .A1(n6911), .A2(n6910), .A3(n6909), .ZN(n6912) );
  NOR3_X1 U8584 ( .A1(n8117), .A2(n7053), .A3(n6912), .ZN(n6913) );
  AOI211_X1 U8585 ( .C1(n8088), .C2(P2_ADDR_REG_7__SCAN_IN), .A(n6914), .B(
        n6913), .ZN(n6915) );
  OAI211_X1 U8586 ( .C1(n8165), .C2(n7047), .A(n6916), .B(n6915), .ZN(P2_U3252) );
  INV_X1 U8587 ( .A(n9563), .ZN(n6917) );
  OR2_X1 U8588 ( .A1(n9776), .A2(n5947), .ZN(n6919) );
  OAI21_X1 U8589 ( .B1(n6920), .B2(n9774), .A(n6919), .ZN(P1_U3454) );
  INV_X1 U8590 ( .A(n6921), .ZN(n6939) );
  AOI22_X1 U8591 ( .A1(n9158), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n9566), .ZN(n6922) );
  OAI21_X1 U8592 ( .B1(n6939), .B2(n9572), .A(n6922), .ZN(P1_U3336) );
  INV_X1 U8593 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n7168) );
  AND2_X1 U8594 ( .A1(n6944), .A2(n6923), .ZN(n6924) );
  NAND2_X1 U8595 ( .A1(n6924), .A2(n6925), .ZN(n6945) );
  OAI21_X1 U8596 ( .B1(n6925), .B2(n6924), .A(n6945), .ZN(n6928) );
  NAND2_X1 U8597 ( .A1(n8066), .A2(n8425), .ZN(n6927) );
  NAND2_X1 U8598 ( .A1(n5760), .A2(n8423), .ZN(n6926) );
  NAND2_X1 U8599 ( .A1(n6927), .A2(n6926), .ZN(n7166) );
  AOI22_X1 U8600 ( .A1(n8033), .A2(n6928), .B1(n7961), .B2(n7166), .ZN(n6930)
         );
  NAND2_X1 U8601 ( .A1(n8041), .A2(n7163), .ZN(n6929) );
  OAI211_X1 U8602 ( .C1(n6951), .C2(n7168), .A(n6930), .B(n6929), .ZN(P2_U3224) );
  NAND2_X1 U8603 ( .A1(n8167), .A2(n4526), .ZN(n6931) );
  OAI211_X1 U8604 ( .C1(P2_REG2_REG_0__SCAN_IN), .C2(n8163), .A(n8165), .B(
        n6931), .ZN(n6932) );
  INV_X1 U8605 ( .A(n6932), .ZN(n6935) );
  INV_X1 U8606 ( .A(n8163), .ZN(n8162) );
  AOI22_X1 U8607 ( .A1(n8162), .A2(P2_REG2_REG_0__SCAN_IN), .B1(
        P2_REG1_REG_0__SCAN_IN), .B2(n8167), .ZN(n6934) );
  MUX2_X1 U8608 ( .A(n6935), .B(n6934), .S(n6933), .Z(n6937) );
  AOI22_X1 U8609 ( .A1(n8088), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3152), .ZN(n6936) );
  NAND2_X1 U8610 ( .A1(n6937), .A2(n6936), .ZN(P2_U3245) );
  INV_X1 U8611 ( .A(n8144), .ZN(n8137) );
  OAI222_X1 U8612 ( .A1(n8583), .A2(n6939), .B1(n8137), .B2(P2_U3152), .C1(
        n6938), .C2(n8587), .ZN(P2_U3341) );
  INV_X1 U8613 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n7037) );
  OR2_X1 U8614 ( .A1(n7131), .A2(n8404), .ZN(n6941) );
  OR2_X1 U8615 ( .A1(n6868), .A2(n8402), .ZN(n6940) );
  NAND2_X1 U8616 ( .A1(n6941), .A2(n6940), .ZN(n7030) );
  AOI22_X1 U8617 ( .A1(n8041), .A2(n7027), .B1(n7961), .B2(n7030), .ZN(n6950)
         );
  NAND2_X1 U8618 ( .A1(n6942), .A2(n6943), .ZN(n6947) );
  NAND2_X1 U8619 ( .A1(n6945), .A2(n6944), .ZN(n6946) );
  XOR2_X1 U8620 ( .A(n6947), .B(n6946), .Z(n6948) );
  NAND2_X1 U8621 ( .A1(n8033), .A2(n6948), .ZN(n6949) );
  OAI211_X1 U8622 ( .C1(n6951), .C2(n7037), .A(n6950), .B(n6949), .ZN(P2_U3239) );
  INV_X1 U8623 ( .A(n6952), .ZN(n6953) );
  NOR2_X1 U8624 ( .A1(n6954), .A2(n6953), .ZN(n6955) );
  XNOR2_X1 U8625 ( .A(n6956), .B(n6955), .ZN(n6963) );
  OR2_X1 U8626 ( .A1(n7131), .A2(n8402), .ZN(n6958) );
  NAND2_X1 U8627 ( .A1(n8063), .A2(n8425), .ZN(n6957) );
  NAND2_X1 U8628 ( .A1(n6958), .A2(n6957), .ZN(n7138) );
  NAND2_X1 U8629 ( .A1(n7961), .A2(n7138), .ZN(n6960) );
  OAI211_X1 U8630 ( .C1(n8029), .C2(n9829), .A(n6960), .B(n6959), .ZN(n6961)
         );
  AOI21_X1 U8631 ( .B1(n7142), .B2(n8042), .A(n6961), .ZN(n6962) );
  OAI21_X1 U8632 ( .B1(n6963), .B2(n8019), .A(n6962), .ZN(P2_U3232) );
  INV_X1 U8633 ( .A(n6964), .ZN(n6966) );
  OAI222_X1 U8634 ( .A1(n4421), .A2(P1_U3084), .B1(n9572), .B2(n6966), .C1(
        n6965), .C2(n9576), .ZN(P1_U3338) );
  INV_X1 U8635 ( .A(n8099), .ZN(n8105) );
  OAI222_X1 U8636 ( .A1(n8587), .A2(n6967), .B1(n8583), .B2(n6966), .C1(
        P2_U3152), .C2(n8105), .ZN(P2_U3343) );
  OAI21_X1 U8637 ( .B1(n6970), .B2(n6969), .A(n6968), .ZN(n6979) );
  NAND2_X1 U8638 ( .A1(n6979), .A2(n8794), .ZN(n6972) );
  NAND2_X1 U8639 ( .A1(n8656), .A2(n7319), .ZN(n8773) );
  AOI22_X1 U8640 ( .A1(n8808), .A2(n6890), .B1(P1_REG3_REG_0__SCAN_IN), .B2(
        n8773), .ZN(n6971) );
  OAI211_X1 U8641 ( .C1(n8801), .C2(n9690), .A(n6972), .B(n6971), .ZN(P1_U3230) );
  INV_X1 U8642 ( .A(n6973), .ZN(n6976) );
  AOI22_X1 U8643 ( .A1(n9626), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(n9566), .ZN(n6974) );
  OAI21_X1 U8644 ( .B1(n6976), .B2(n9572), .A(n6974), .ZN(P1_U3337) );
  AOI22_X1 U8645 ( .A1(n8128), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_16__SCAN_IN), .B2(n8581), .ZN(n6975) );
  OAI21_X1 U8646 ( .B1(n6976), .B2(n8583), .A(n6975), .ZN(P2_U3342) );
  MUX2_X1 U8647 ( .A(n6979), .B(n6978), .S(n6977), .Z(n6981) );
  MUX2_X1 U8648 ( .A(P1_IR_REG_0__SCAN_IN), .B(n6981), .S(n6980), .Z(n6982) );
  NAND2_X1 U8649 ( .A1(n6982), .A2(P1_U4006), .ZN(n9131) );
  NAND2_X1 U8650 ( .A1(n6984), .A2(n6983), .ZN(n6985) );
  AND2_X1 U8651 ( .A1(n6986), .A2(n6985), .ZN(n6987) );
  NAND2_X1 U8652 ( .A1(P1_U3084), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n7401) );
  OAI21_X1 U8653 ( .B1(n9163), .B2(n6987), .A(n7401), .ZN(n6995) );
  INV_X1 U8654 ( .A(n6988), .ZN(n6989) );
  AOI21_X1 U8655 ( .B1(n6991), .B2(n6990), .A(n6989), .ZN(n6992) );
  OAI22_X1 U8656 ( .A1(n9654), .A2(n6993), .B1(n6992), .B2(n9620), .ZN(n6994)
         );
  AOI211_X1 U8657 ( .C1(n9171), .C2(P1_ADDR_REG_4__SCAN_IN), .A(n6995), .B(
        n6994), .ZN(n6996) );
  NAND2_X1 U8658 ( .A1(n9131), .A2(n6996), .ZN(P1_U3245) );
  NAND2_X1 U8659 ( .A1(n6998), .A2(n6997), .ZN(n7229) );
  OAI21_X1 U8660 ( .B1(n6998), .B2(n6997), .A(n7229), .ZN(n7003) );
  AOI21_X1 U8661 ( .B1(n7003), .B2(n7002), .A(n7233), .ZN(n7013) );
  INV_X1 U8662 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n7004) );
  NAND2_X1 U8663 ( .A1(P1_U3084), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n8667) );
  OAI21_X1 U8664 ( .B1(n9662), .B2(n7004), .A(n8667), .ZN(n7005) );
  AOI21_X1 U8665 ( .B1(n7237), .B2(n9627), .A(n7005), .ZN(n7012) );
  OR2_X1 U8666 ( .A1(n7006), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n7007) );
  INV_X1 U8667 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n7701) );
  XNOR2_X1 U8668 ( .A(n7237), .B(n7701), .ZN(n7009) );
  OAI211_X1 U8669 ( .C1(n7010), .C2(n7009), .A(n7239), .B(n9648), .ZN(n7011)
         );
  OAI211_X1 U8670 ( .C1(n7013), .C2(n9163), .A(n7012), .B(n7011), .ZN(P1_U3253) );
  INV_X1 U8671 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n7041) );
  NAND2_X1 U8672 ( .A1(n7015), .A2(n7014), .ZN(n7110) );
  AND2_X1 U8673 ( .A1(n7110), .A2(n7115), .ZN(n7033) );
  NAND2_X1 U8674 ( .A1(n7035), .A2(n7033), .ZN(n7016) );
  NAND2_X1 U8675 ( .A1(n7017), .A2(n7020), .ZN(n7018) );
  NAND3_X1 U8676 ( .A1(n7019), .A2(n7207), .A3(n7018), .ZN(n7566) );
  OR2_X1 U8677 ( .A1(n7020), .A2(n7207), .ZN(n7071) );
  NAND2_X1 U8678 ( .A1(n7566), .A2(n7071), .ZN(n9787) );
  NAND2_X1 U8679 ( .A1(n6868), .A2(n4823), .ZN(n7023) );
  NAND2_X1 U8680 ( .A1(n7024), .A2(n7023), .ZN(n7067) );
  XNOR2_X1 U8681 ( .A(n7067), .B(n7066), .ZN(n7127) );
  INV_X1 U8682 ( .A(n7025), .ZN(n7026) );
  AOI22_X1 U8683 ( .A1(n8284), .A2(n7127), .B1(n8414), .B2(n7027), .ZN(n7040)
         );
  XOR2_X1 U8684 ( .A(n5603), .B(n7066), .Z(n7032) );
  NAND2_X1 U8685 ( .A1(n7029), .A2(n7028), .ZN(n9786) );
  INV_X1 U8686 ( .A(n9786), .ZN(n8399) );
  INV_X1 U8687 ( .A(n7030), .ZN(n7031) );
  OAI21_X1 U8688 ( .B1(n7032), .B2(n8399), .A(n7031), .ZN(n7125) );
  AND2_X1 U8689 ( .A1(n7033), .A2(n7207), .ZN(n7034) );
  NAND2_X1 U8690 ( .A1(n7035), .A2(n7034), .ZN(n7218) );
  INV_X1 U8691 ( .A(n7073), .ZN(n7036) );
  INV_X1 U8692 ( .A(n5873), .ZN(n9811) );
  OAI211_X1 U8693 ( .C1(n7124), .C2(n7161), .A(n7036), .B(n9811), .ZN(n7123)
         );
  OAI22_X1 U8694 ( .A1(n7218), .A2(n7123), .B1(n7037), .B2(n8411), .ZN(n7038)
         );
  AOI21_X1 U8695 ( .B1(n9798), .B2(n7125), .A(n7038), .ZN(n7039) );
  OAI211_X1 U8696 ( .C1(n7041), .C2(n9798), .A(n7040), .B(n7039), .ZN(P2_U3294) );
  XNOR2_X1 U8697 ( .A(n7292), .B(P2_REG2_REG_8__SCAN_IN), .ZN(n7044) );
  AOI211_X1 U8698 ( .C1(n7045), .C2(n7044), .A(n8163), .B(n7291), .ZN(n7057)
         );
  NAND2_X1 U8699 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(P2_U3152), .ZN(n7301) );
  INV_X1 U8700 ( .A(n7301), .ZN(n7046) );
  AOI21_X1 U8701 ( .B1(n8088), .B2(P2_ADDR_REG_8__SCAN_IN), .A(n7046), .ZN(
        n7055) );
  INV_X1 U8702 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n9872) );
  MUX2_X1 U8703 ( .A(n9872), .B(P2_REG1_REG_8__SCAN_IN), .S(n7292), .Z(n7049)
         );
  NOR2_X1 U8704 ( .A1(n7047), .A2(n9868), .ZN(n7051) );
  INV_X1 U8705 ( .A(n7051), .ZN(n7048) );
  NAND2_X1 U8706 ( .A1(n7049), .A2(n7048), .ZN(n7052) );
  MUX2_X1 U8707 ( .A(P2_REG1_REG_8__SCAN_IN), .B(n9872), .S(n7292), .Z(n7050)
         );
  OAI211_X1 U8708 ( .C1(n7053), .C2(n7052), .A(n8167), .B(n7286), .ZN(n7054)
         );
  OAI211_X1 U8709 ( .C1(n8165), .C2(n7287), .A(n7055), .B(n7054), .ZN(n7056)
         );
  OR2_X1 U8710 ( .A1(n7057), .A2(n7056), .ZN(P2_U3253) );
  XOR2_X1 U8711 ( .A(n7059), .B(n7058), .Z(n7064) );
  OR2_X1 U8712 ( .A1(n7177), .A2(n8404), .ZN(n7061) );
  NAND2_X1 U8713 ( .A1(n8066), .A2(n8423), .ZN(n7060) );
  AND2_X1 U8714 ( .A1(n7061), .A2(n7060), .ZN(n7080) );
  OAI22_X1 U8715 ( .A1(n8029), .A2(n9821), .B1(n8024), .B2(n7080), .ZN(n7063)
         );
  MUX2_X1 U8716 ( .A(n8042), .B(P2_U3152), .S(P2_REG3_REG_3__SCAN_IN), .Z(
        n7062) );
  AOI211_X1 U8717 ( .C1(n8033), .C2(n7064), .A(n7063), .B(n7062), .ZN(n7065)
         );
  INV_X1 U8718 ( .A(n7065), .ZN(P2_U3220) );
  NAND2_X1 U8719 ( .A1(n7067), .A2(n7066), .ZN(n7070) );
  INV_X1 U8720 ( .A(n8066), .ZN(n7068) );
  NAND2_X1 U8721 ( .A1(n7068), .A2(n7124), .ZN(n7069) );
  NAND2_X1 U8722 ( .A1(n7070), .A2(n7069), .ZN(n7130) );
  XNOR2_X1 U8723 ( .A(n7130), .B(n7129), .ZN(n9819) );
  INV_X1 U8724 ( .A(n9819), .ZN(n7087) );
  INV_X1 U8725 ( .A(n7071), .ZN(n7072) );
  NAND2_X1 U8726 ( .A1(n9798), .A2(n7072), .ZN(n8418) );
  OAI211_X1 U8727 ( .C1(n7073), .C2(n9821), .A(n9811), .B(n7141), .ZN(n9820)
         );
  OAI22_X1 U8728 ( .A1(n7218), .A2(n9820), .B1(P2_REG3_REG_3__SCAN_IN), .B2(
        n8411), .ZN(n7076) );
  INV_X1 U8729 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n7074) );
  NOR2_X1 U8730 ( .A1(n9798), .A2(n7074), .ZN(n7075) );
  AOI211_X1 U8731 ( .C1(n8414), .C2(n7077), .A(n7076), .B(n7075), .ZN(n7086)
         );
  INV_X1 U8732 ( .A(n7566), .ZN(n8408) );
  NAND2_X1 U8733 ( .A1(n9819), .A2(n8408), .ZN(n7084) );
  XNOR2_X1 U8734 ( .A(n7078), .B(n7079), .ZN(n7082) );
  INV_X1 U8735 ( .A(n7080), .ZN(n7081) );
  AOI21_X1 U8736 ( .B1(n7082), .B2(n9786), .A(n7081), .ZN(n7083) );
  NAND2_X1 U8737 ( .A1(n7084), .A2(n7083), .ZN(n9823) );
  NAND2_X1 U8738 ( .A1(n9823), .A2(n9798), .ZN(n7085) );
  OAI211_X1 U8739 ( .C1(n7087), .C2(n8418), .A(n7086), .B(n7085), .ZN(P2_U3293) );
  INV_X1 U8740 ( .A(n7088), .ZN(n7259) );
  INV_X1 U8741 ( .A(n8035), .ZN(n7950) );
  OAI22_X1 U8742 ( .A1(n7950), .A2(n4501), .B1(n7177), .B2(n8039), .ZN(n7089)
         );
  AOI211_X1 U8743 ( .C1(n8041), .C2(n7262), .A(n7090), .B(n7089), .ZN(n7096)
         );
  OAI21_X1 U8744 ( .B1(n7093), .B2(n7092), .A(n7091), .ZN(n7094) );
  NAND2_X1 U8745 ( .A1(n7094), .A2(n8033), .ZN(n7095) );
  OAI211_X1 U8746 ( .C1(n8023), .C2(n7259), .A(n7096), .B(n7095), .ZN(P2_U3229) );
  INV_X1 U8747 ( .A(n7097), .ZN(n7149) );
  AOI22_X1 U8748 ( .A1(n8151), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_18__SCAN_IN), .B2(n8581), .ZN(n7098) );
  OAI21_X1 U8749 ( .B1(n7149), .B2(n8583), .A(n7098), .ZN(P2_U3340) );
  INV_X1 U8750 ( .A(n7099), .ZN(n7101) );
  NAND2_X1 U8751 ( .A1(n7101), .A2(n7100), .ZN(n7104) );
  AOI22_X1 U8752 ( .A1(n7105), .A2(n7104), .B1(n7102), .B2(n7103), .ZN(n7109)
         );
  AOI22_X1 U8753 ( .A1(n8808), .A2(n6893), .B1(n8748), .B2(n7106), .ZN(n7108)
         );
  AOI22_X1 U8754 ( .A1(n8812), .A2(n9692), .B1(n8773), .B2(
        P1_REG3_REG_1__SCAN_IN), .ZN(n7107) );
  OAI211_X1 U8755 ( .C1(n7109), .C2(n8814), .A(n7108), .B(n7107), .ZN(P1_U3220) );
  NAND3_X1 U8756 ( .A1(n7112), .A2(n7111), .A3(n7110), .ZN(n7113) );
  OR2_X1 U8757 ( .A1(n7114), .A2(n7113), .ZN(n7854) );
  NOR2_X1 U8758 ( .A1(n9791), .A2(n7116), .ZN(n7117) );
  NOR2_X1 U8759 ( .A1(n9788), .A2(n7117), .ZN(n7121) );
  NAND2_X1 U8760 ( .A1(n9790), .A2(n9786), .ZN(n7120) );
  AND2_X1 U8761 ( .A1(n5568), .A2(n5587), .ZN(n7118) );
  NAND2_X1 U8762 ( .A1(n7017), .A2(n7118), .ZN(n9818) );
  NAND2_X1 U8763 ( .A1(n7566), .A2(n9818), .ZN(n9851) );
  NAND2_X1 U8764 ( .A1(n9790), .A2(n9851), .ZN(n7119) );
  AND3_X1 U8765 ( .A1(n7121), .A2(n7120), .A3(n7119), .ZN(n9808) );
  NAND2_X1 U8766 ( .A1(n9871), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n7122) );
  OAI21_X1 U8767 ( .B1(n9871), .B2(n9808), .A(n7122), .ZN(P2_U3520) );
  OAI21_X1 U8768 ( .B1(n9854), .B2(n7124), .A(n7123), .ZN(n7126) );
  AOI211_X1 U8769 ( .C1(n9851), .C2(n7127), .A(n7126), .B(n7125), .ZN(n9817)
         );
  NAND2_X1 U8770 ( .A1(n9871), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n7128) );
  OAI21_X1 U8771 ( .B1(n9817), .B2(n9871), .A(n7128), .ZN(P2_U3522) );
  NAND2_X1 U8772 ( .A1(n7130), .A2(n7129), .ZN(n7133) );
  NAND2_X1 U8773 ( .A1(n7131), .A2(n9821), .ZN(n7132) );
  NAND2_X1 U8774 ( .A1(n7133), .A2(n7132), .ZN(n7176) );
  XNOR2_X1 U8775 ( .A(n7176), .B(n7134), .ZN(n9826) );
  INV_X1 U8776 ( .A(n7135), .ZN(n7136) );
  NOR2_X1 U8777 ( .A1(n7137), .A2(n7136), .ZN(n7249) );
  NAND2_X1 U8778 ( .A1(n7249), .A2(n7247), .ZN(n7140) );
  AOI21_X1 U8779 ( .B1(n7137), .B2(n7175), .A(n8399), .ZN(n7139) );
  AOI21_X1 U8780 ( .B1(n7140), .B2(n7139), .A(n7138), .ZN(n9828) );
  MUX2_X1 U8781 ( .A(n6763), .B(n9828), .S(n9798), .Z(n7147) );
  OAI211_X1 U8782 ( .C1(n4407), .C2(n9829), .A(n9811), .B(n7255), .ZN(n9827)
         );
  INV_X1 U8783 ( .A(n7142), .ZN(n7143) );
  OAI22_X1 U8784 ( .A1(n7218), .A2(n9827), .B1(n8411), .B2(n7143), .ZN(n7144)
         );
  AOI21_X1 U8785 ( .B1(n8414), .B2(n7145), .A(n7144), .ZN(n7146) );
  OAI211_X1 U8786 ( .C1(n9826), .C2(n8436), .A(n7147), .B(n7146), .ZN(P2_U3292) );
  INV_X1 U8787 ( .A(n9152), .ZN(n9653) );
  INV_X1 U8788 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n7148) );
  OAI222_X1 U8789 ( .A1(n9653), .A2(P1_U3084), .B1(n9572), .B2(n7149), .C1(
        n7148), .C2(n9576), .ZN(P1_U3335) );
  OAI21_X1 U8790 ( .B1(n7152), .B2(n7151), .A(n7150), .ZN(n7153) );
  NAND2_X1 U8791 ( .A1(n7153), .A2(n8033), .ZN(n7160) );
  INV_X1 U8792 ( .A(n7219), .ZN(n9842) );
  OR2_X1 U8793 ( .A1(n7416), .A2(n8404), .ZN(n7155) );
  NAND2_X1 U8794 ( .A1(n8063), .A2(n8423), .ZN(n7154) );
  NAND2_X1 U8795 ( .A1(n7155), .A2(n7154), .ZN(n7216) );
  NAND2_X1 U8796 ( .A1(n7961), .A2(n7216), .ZN(n7157) );
  OAI211_X1 U8797 ( .C1(n8029), .C2(n9842), .A(n7157), .B(n7156), .ZN(n7158)
         );
  AOI21_X1 U8798 ( .B1(n7221), .B2(n8042), .A(n7158), .ZN(n7159) );
  NAND2_X1 U8799 ( .A1(n7160), .A2(n7159), .ZN(P2_U3241) );
  OAI22_X1 U8800 ( .A1(n4823), .A2(n9793), .B1(n8436), .B2(n9809), .ZN(n7171)
         );
  NAND2_X1 U8801 ( .A1(n7163), .A2(n7162), .ZN(n9810) );
  NAND2_X1 U8802 ( .A1(n4648), .A2(n9810), .ZN(n7164) );
  OAI22_X1 U8803 ( .A1(n9792), .A2(n7164), .B1(n9798), .B2(n6711), .ZN(n7170)
         );
  AOI21_X1 U8804 ( .B1(n7167), .B2(n9786), .A(n7166), .ZN(n9813) );
  OAI22_X1 U8805 ( .A1(n4262), .A2(n9813), .B1(n8411), .B2(n7168), .ZN(n7169)
         );
  OR3_X1 U8806 ( .A1(n7171), .A2(n7170), .A3(n7169), .ZN(P2_U3295) );
  INV_X1 U8807 ( .A(n7172), .ZN(n7212) );
  OAI222_X1 U8808 ( .A1(n8583), .A2(n7212), .B1(P2_U3152), .B2(n7173), .C1(
        n9904), .C2(n8587), .ZN(P2_U3337) );
  NAND2_X1 U8809 ( .A1(n7177), .A2(n9829), .ZN(n7178) );
  INV_X1 U8810 ( .A(n7250), .ZN(n7180) );
  NAND2_X1 U8811 ( .A1(n7180), .A2(n7262), .ZN(n7181) );
  XNOR2_X1 U8812 ( .A(n7411), .B(n7410), .ZN(n9850) );
  INV_X1 U8813 ( .A(n9850), .ZN(n7191) );
  XNOR2_X1 U8814 ( .A(n7182), .B(n7410), .ZN(n7183) );
  OAI222_X1 U8815 ( .A1(n8404), .A2(n7452), .B1(n8402), .B2(n4501), .C1(n7183), 
        .C2(n8399), .ZN(n9848) );
  INV_X1 U8816 ( .A(n7412), .ZN(n9846) );
  OAI21_X1 U8817 ( .B1(n7184), .B2(n9846), .A(n7423), .ZN(n9847) );
  INV_X1 U8818 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n7186) );
  INV_X1 U8819 ( .A(n7196), .ZN(n7185) );
  OAI22_X1 U8820 ( .A1(n9798), .A2(n7186), .B1(n8411), .B2(n7185), .ZN(n7187)
         );
  AOI21_X1 U8821 ( .B1(n8414), .B2(n7412), .A(n7187), .ZN(n7188) );
  OAI21_X1 U8822 ( .B1(n9792), .B2(n9847), .A(n7188), .ZN(n7189) );
  AOI21_X1 U8823 ( .B1(n9848), .B2(n9798), .A(n7189), .ZN(n7190) );
  OAI21_X1 U8824 ( .B1(n7191), .B2(n8436), .A(n7190), .ZN(P2_U3289) );
  XNOR2_X1 U8825 ( .A(n7193), .B(n7192), .ZN(n7198) );
  OAI22_X1 U8826 ( .A1(n8029), .A2(n9846), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n5115), .ZN(n7195) );
  OAI22_X1 U8827 ( .A1(n7950), .A2(n7452), .B1(n4501), .B2(n8039), .ZN(n7194)
         );
  AOI211_X1 U8828 ( .C1(n7196), .C2(n8042), .A(n7195), .B(n7194), .ZN(n7197)
         );
  OAI21_X1 U8829 ( .B1(n7198), .B2(n8019), .A(n7197), .ZN(P2_U3215) );
  XOR2_X1 U8830 ( .A(n7200), .B(n7199), .Z(n7205) );
  OAI21_X1 U8831 ( .B1(n8806), .B2(n9701), .A(n7201), .ZN(n7203) );
  OAI22_X1 U8832 ( .A1(n7351), .A2(n8801), .B1(n8810), .B2(
        P1_REG3_REG_3__SCAN_IN), .ZN(n7202) );
  AOI211_X1 U8833 ( .C1(n8808), .C2(n9115), .A(n7203), .B(n7202), .ZN(n7204)
         );
  OAI21_X1 U8834 ( .B1(n7205), .B2(n8814), .A(n7204), .ZN(P1_U3216) );
  INV_X1 U8835 ( .A(n7206), .ZN(n7210) );
  OAI222_X1 U8836 ( .A1(n8587), .A2(n7208), .B1(n8583), .B2(n7210), .C1(n7207), 
        .C2(P2_U3152), .ZN(P2_U3339) );
  OAI222_X1 U8837 ( .A1(P1_U3084), .A2(n9694), .B1(n9572), .B2(n7210), .C1(
        n7209), .C2(n9576), .ZN(P1_U3334) );
  OAI222_X1 U8838 ( .A1(n9091), .A2(P1_U3084), .B1(n9572), .B2(n7212), .C1(
        n7211), .C2(n9576), .ZN(P1_U3332) );
  OAI21_X1 U8839 ( .B1(n7249), .B2(n7214), .A(n7213), .ZN(n7215) );
  XNOR2_X1 U8840 ( .A(n7215), .B(n7225), .ZN(n7217) );
  AOI21_X1 U8841 ( .B1(n7217), .B2(n9786), .A(n7216), .ZN(n9841) );
  INV_X1 U8842 ( .A(n7218), .ZN(n7645) );
  XNOR2_X1 U8843 ( .A(n7258), .B(n7219), .ZN(n7220) );
  NAND2_X1 U8844 ( .A1(n7220), .A2(n9811), .ZN(n9840) );
  INV_X1 U8845 ( .A(n9840), .ZN(n7224) );
  INV_X1 U8846 ( .A(n8411), .ZN(n9795) );
  AOI22_X1 U8847 ( .A1(n4262), .A2(P2_REG2_REG_6__SCAN_IN), .B1(n9795), .B2(
        n7221), .ZN(n7222) );
  OAI21_X1 U8848 ( .B1(n9793), .B2(n9842), .A(n7222), .ZN(n7223) );
  AOI21_X1 U8849 ( .B1(n7645), .B2(n7224), .A(n7223), .ZN(n7228) );
  XNOR2_X1 U8850 ( .A(n7226), .B(n7225), .ZN(n9844) );
  NAND2_X1 U8851 ( .A1(n9844), .A2(n8284), .ZN(n7227) );
  OAI211_X1 U8852 ( .C1(n9841), .C2(n4262), .A(n7228), .B(n7227), .ZN(P2_U3290) );
  INV_X1 U8853 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n9997) );
  NAND2_X1 U8854 ( .A1(P1_U3084), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n8736) );
  OAI21_X1 U8855 ( .B1(n9662), .B2(n9997), .A(n8736), .ZN(n7236) );
  INV_X1 U8856 ( .A(n7229), .ZN(n7232) );
  OR2_X1 U8857 ( .A1(n7270), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n7277) );
  NAND2_X1 U8858 ( .A1(n7270), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n7230) );
  AND2_X1 U8859 ( .A1(n7277), .A2(n7230), .ZN(n7231) );
  OR3_X1 U8860 ( .A1(n7233), .A2(n7232), .A3(n7231), .ZN(n7234) );
  AOI21_X1 U8861 ( .B1(n7278), .B2(n7234), .A(n9163), .ZN(n7235) );
  AOI211_X1 U8862 ( .C1(n9627), .C2(n7270), .A(n7236), .B(n7235), .ZN(n7244)
         );
  NAND2_X1 U8863 ( .A1(n7237), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n7238) );
  NAND2_X1 U8864 ( .A1(n7239), .A2(n7238), .ZN(n7242) );
  INV_X1 U8865 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n7240) );
  XNOR2_X1 U8866 ( .A(n7270), .B(n7240), .ZN(n7241) );
  NAND2_X1 U8867 ( .A1(n7242), .A2(n7241), .ZN(n7272) );
  OAI211_X1 U8868 ( .C1(n7242), .C2(n7241), .A(n7272), .B(n9648), .ZN(n7243)
         );
  NAND2_X1 U8869 ( .A1(n7244), .A2(n7243), .ZN(P1_U3254) );
  INV_X1 U8870 ( .A(n7245), .ZN(n7269) );
  OAI222_X1 U8871 ( .A1(n8583), .A2(n7269), .B1(P2_U3152), .B2(n5568), .C1(
        n7246), .C2(n8587), .ZN(P2_U3338) );
  INV_X1 U8872 ( .A(n9833), .ZN(n7267) );
  INV_X1 U8873 ( .A(n7247), .ZN(n7248) );
  OR2_X1 U8874 ( .A1(n7249), .A2(n7248), .ZN(n7251) );
  XNOR2_X1 U8875 ( .A(n7250), .B(n7251), .ZN(n7252) );
  NAND2_X1 U8876 ( .A1(n7252), .A2(n9786), .ZN(n7254) );
  AOI22_X1 U8877 ( .A1(n8064), .A2(n8423), .B1(n8425), .B2(n8062), .ZN(n7253)
         );
  NAND2_X1 U8878 ( .A1(n7254), .A2(n7253), .ZN(n9838) );
  NOR2_X1 U8879 ( .A1(n4262), .A2(n5587), .ZN(n8382) );
  INV_X1 U8880 ( .A(n8382), .ZN(n7264) );
  NAND2_X1 U8881 ( .A1(n7255), .A2(n7262), .ZN(n7256) );
  NAND2_X1 U8882 ( .A1(n7256), .A2(n9811), .ZN(n7257) );
  OR2_X1 U8883 ( .A1(n7258), .A2(n7257), .ZN(n9834) );
  INV_X1 U8884 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n7260) );
  OAI22_X1 U8885 ( .A1(n9798), .A2(n7260), .B1(n8411), .B2(n7259), .ZN(n7261)
         );
  AOI21_X1 U8886 ( .B1(n8414), .B2(n7262), .A(n7261), .ZN(n7263) );
  OAI21_X1 U8887 ( .B1(n7264), .B2(n9834), .A(n7263), .ZN(n7265) );
  AOI21_X1 U8888 ( .B1(n9798), .B2(n9838), .A(n7265), .ZN(n7266) );
  OAI21_X1 U8889 ( .B1(n7267), .B2(n8436), .A(n7266), .ZN(P2_U3291) );
  OAI222_X1 U8890 ( .A1(n8938), .A2(P1_U3084), .B1(n9572), .B2(n7269), .C1(
        n7268), .C2(n9576), .ZN(P1_U3333) );
  NAND2_X1 U8891 ( .A1(n7270), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n7271) );
  INV_X1 U8892 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n7273) );
  NAND2_X1 U8893 ( .A1(n7274), .A2(n7273), .ZN(n9145) );
  OAI21_X1 U8894 ( .B1(n7274), .B2(n7273), .A(n9145), .ZN(n7275) );
  INV_X1 U8895 ( .A(n7275), .ZN(n7285) );
  XNOR2_X1 U8896 ( .A(n9155), .B(n7276), .ZN(n7280) );
  NAND2_X1 U8897 ( .A1(n7279), .A2(n7280), .ZN(n9154) );
  OAI21_X1 U8898 ( .B1(n7280), .B2(n7279), .A(n9154), .ZN(n7283) );
  NAND2_X1 U8899 ( .A1(P1_U3084), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n8594) );
  NAND2_X1 U8900 ( .A1(n9171), .A2(P1_ADDR_REG_14__SCAN_IN), .ZN(n7281) );
  OAI211_X1 U8901 ( .C1(n9654), .C2(n4420), .A(n8594), .B(n7281), .ZN(n7282)
         );
  AOI21_X1 U8902 ( .B1(n7283), .B2(n9659), .A(n7282), .ZN(n7284) );
  OAI21_X1 U8903 ( .B1(n7285), .B2(n9620), .A(n7284), .ZN(P1_U3255) );
  XOR2_X1 U8904 ( .A(P2_REG1_REG_9__SCAN_IN), .B(n7467), .Z(n7462) );
  OAI21_X1 U8905 ( .B1(n9872), .B2(n7287), .A(n7286), .ZN(n7463) );
  XOR2_X1 U8906 ( .A(n7462), .B(n7463), .Z(n7297) );
  NAND2_X1 U8907 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(P2_U3152), .ZN(n7450) );
  INV_X1 U8908 ( .A(n7450), .ZN(n7288) );
  AOI21_X1 U8909 ( .B1(n8088), .B2(P2_ADDR_REG_9__SCAN_IN), .A(n7288), .ZN(
        n7289) );
  OAI21_X1 U8910 ( .B1(n8165), .B2(n7290), .A(n7289), .ZN(n7296) );
  XNOR2_X1 U8911 ( .A(n7467), .B(P2_REG2_REG_9__SCAN_IN), .ZN(n7293) );
  AOI211_X1 U8912 ( .C1(n7294), .C2(n7293), .A(n8163), .B(n7466), .ZN(n7295)
         );
  AOI211_X1 U8913 ( .C1(n8167), .C2(n7297), .A(n7296), .B(n7295), .ZN(n7298)
         );
  INV_X1 U8914 ( .A(n7298), .ZN(P2_U3254) );
  XNOR2_X1 U8915 ( .A(n7300), .B(n7299), .ZN(n7306) );
  INV_X1 U8916 ( .A(n7556), .ZN(n8059) );
  NAND2_X1 U8917 ( .A1(n8035), .A2(n8059), .ZN(n7302) );
  NAND2_X1 U8918 ( .A1(n7302), .A2(n7301), .ZN(n7304) );
  OAI22_X1 U8919 ( .A1(n8039), .A2(n7416), .B1(n4643), .B2(n8029), .ZN(n7303)
         );
  AOI211_X1 U8920 ( .C1(n7420), .C2(n8042), .A(n7304), .B(n7303), .ZN(n7305)
         );
  OAI21_X1 U8921 ( .B1(n7306), .B2(n8019), .A(n7305), .ZN(P2_U3223) );
  NAND2_X1 U8922 ( .A1(n7397), .A2(n7307), .ZN(n7311) );
  XOR2_X1 U8923 ( .A(n7309), .B(n7308), .Z(n7310) );
  XNOR2_X1 U8924 ( .A(n7311), .B(n7310), .ZN(n7316) );
  AND2_X1 U8925 ( .A1(n9736), .A2(n7602), .ZN(n9750) );
  AND2_X1 U8926 ( .A1(n9398), .A2(n9113), .ZN(n7597) );
  NAND2_X1 U8927 ( .A1(n8771), .A2(n7597), .ZN(n7312) );
  NAND2_X1 U8928 ( .A1(P1_U3084), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n9142) );
  OAI211_X1 U8929 ( .C1(n8806), .C2(n7354), .A(n7312), .B(n9142), .ZN(n7314)
         );
  NOR2_X1 U8930 ( .A1(n8810), .A2(n7603), .ZN(n7313) );
  AOI211_X1 U8931 ( .C1(n9750), .C2(n8656), .A(n7314), .B(n7313), .ZN(n7315)
         );
  OAI21_X1 U8932 ( .B1(n7316), .B2(n8814), .A(n7315), .ZN(P1_U3225) );
  NOR2_X1 U8933 ( .A1(n9563), .A2(n9722), .ZN(n7317) );
  AND2_X1 U8934 ( .A1(n7318), .A2(n7317), .ZN(n7320) );
  NAND2_X1 U8935 ( .A1(n7320), .A2(n7319), .ZN(n7375) );
  INV_X1 U8936 ( .A(n7321), .ZN(n7331) );
  NAND3_X1 U8937 ( .A1(n9713), .A2(n9101), .A3(n7322), .ZN(n9431) );
  INV_X1 U8938 ( .A(n9431), .ZN(n9391) );
  AND2_X1 U8939 ( .A1(n9713), .A2(n7323), .ZN(n9670) );
  INV_X1 U8940 ( .A(n9670), .ZN(n9177) );
  OAI22_X1 U8941 ( .A1(n9713), .A2(n7324), .B1(n9122), .B2(n9697), .ZN(n7325)
         );
  AOI21_X1 U8942 ( .B1(n9426), .B2(n8774), .A(n7325), .ZN(n7326) );
  OAI21_X1 U8943 ( .B1(n9177), .B2(n7327), .A(n7326), .ZN(n7328) );
  AOI21_X1 U8944 ( .B1(n9391), .B2(n7329), .A(n7328), .ZN(n7330) );
  OAI21_X1 U8945 ( .B1(n9716), .B2(n7331), .A(n7330), .ZN(P1_U3289) );
  XNOR2_X1 U8946 ( .A(n7333), .B(n7332), .ZN(n7334) );
  XNOR2_X1 U8947 ( .A(n7335), .B(n7334), .ZN(n7341) );
  AOI21_X1 U8948 ( .B1(n8748), .B2(n9114), .A(n7336), .ZN(n7338) );
  INV_X1 U8949 ( .A(n7615), .ZN(n9112) );
  NAND2_X1 U8950 ( .A1(n8808), .A2(n9112), .ZN(n7337) );
  OAI211_X1 U8951 ( .C1(n8810), .C2(n7390), .A(n7338), .B(n7337), .ZN(n7339)
         );
  AOI21_X1 U8952 ( .B1(n8812), .B2(n7358), .A(n7339), .ZN(n7340) );
  OAI21_X1 U8953 ( .B1(n7341), .B2(n8814), .A(n7340), .ZN(P1_U3237) );
  INV_X1 U8954 ( .A(n7342), .ZN(n7347) );
  AOI21_X1 U8955 ( .B1(P1_DATAO_REG_23__SCAN_IN), .B2(n8581), .A(n7343), .ZN(
        n7344) );
  OAI21_X1 U8956 ( .B1(n7347), .B2(n8583), .A(n7344), .ZN(P2_U3335) );
  OR2_X1 U8957 ( .A1(n7345), .A2(P1_U3084), .ZN(n9104) );
  NAND2_X1 U8958 ( .A1(n9566), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n7346) );
  OAI211_X1 U8959 ( .C1(n7347), .C2(n9572), .A(n9104), .B(n7346), .ZN(P1_U3330) );
  NAND2_X1 U8960 ( .A1(n7348), .A2(n9058), .ZN(n7350) );
  OR2_X1 U8961 ( .A1(n6893), .A2(n8774), .ZN(n7349) );
  NAND2_X1 U8962 ( .A1(n9116), .A2(n7351), .ZN(n8988) );
  NAND2_X1 U8963 ( .A1(n7477), .A2(n9060), .ZN(n7353) );
  OR2_X1 U8964 ( .A1(n9116), .A2(n9729), .ZN(n7352) );
  NAND2_X1 U8965 ( .A1(n7354), .A2(n9735), .ZN(n8991) );
  NAND2_X1 U8966 ( .A1(n8991), .A2(n9015), .ZN(n9675) );
  NAND2_X1 U8967 ( .A1(n9665), .A2(n9675), .ZN(n7356) );
  OR2_X1 U8968 ( .A1(n9735), .A2(n9115), .ZN(n7355) );
  NAND2_X1 U8969 ( .A1(n7356), .A2(n7355), .ZN(n7383) );
  OR2_X1 U8970 ( .A1(n7358), .A2(n7357), .ZN(n8861) );
  NAND2_X1 U8971 ( .A1(n7358), .A2(n7357), .ZN(n9019) );
  NAND2_X1 U8972 ( .A1(n8861), .A2(n9019), .ZN(n7385) );
  NAND2_X1 U8973 ( .A1(n7602), .A2(n9114), .ZN(n7384) );
  NAND2_X1 U8974 ( .A1(n7383), .A2(n7359), .ZN(n7508) );
  NAND2_X1 U8975 ( .A1(n7602), .A2(n9676), .ZN(n9018) );
  OR2_X1 U8976 ( .A1(n7358), .A2(n9113), .ZN(n7360) );
  NAND2_X1 U8977 ( .A1(n7361), .A2(n7360), .ZN(n7505) );
  INV_X1 U8978 ( .A(n7505), .ZN(n7362) );
  NAND2_X1 U8979 ( .A1(n7508), .A2(n7362), .ZN(n7364) );
  NAND2_X1 U8980 ( .A1(n7363), .A2(n7615), .ZN(n8868) );
  INV_X1 U8981 ( .A(n9066), .ZN(n7504) );
  XNOR2_X1 U8982 ( .A(n7364), .B(n7504), .ZN(n9760) );
  INV_X1 U8983 ( .A(n9760), .ZN(n7382) );
  AND2_X1 U8984 ( .A1(n9015), .A2(n7367), .ZN(n7368) );
  NAND2_X1 U8985 ( .A1(n7596), .A2(n9016), .ZN(n7369) );
  NAND2_X2 U8986 ( .A1(n7369), .A2(n9018), .ZN(n8867) );
  NAND2_X1 U8987 ( .A1(n8867), .A2(n8861), .ZN(n7370) );
  NAND2_X1 U8988 ( .A1(n7370), .A2(n9019), .ZN(n7371) );
  NAND2_X1 U8989 ( .A1(n7371), .A2(n9066), .ZN(n7515) );
  OAI21_X1 U8990 ( .B1(n9066), .B2(n7371), .A(n7515), .ZN(n7372) );
  NAND2_X1 U8991 ( .A1(n7372), .A2(n9706), .ZN(n7374) );
  AOI22_X1 U8992 ( .A1(n9396), .A2(n9113), .B1(n9398), .B2(n9111), .ZN(n7373)
         );
  NAND2_X1 U8993 ( .A1(n7374), .A2(n7373), .ZN(n9765) );
  OR2_X1 U8994 ( .A1(n7375), .A2(n9169), .ZN(n9422) );
  NAND2_X1 U8995 ( .A1(n9667), .A2(n9682), .ZN(n9668) );
  OAI21_X1 U8996 ( .B1(n7388), .B2(n9762), .A(n9737), .ZN(n7376) );
  OR2_X1 U8997 ( .A1(n7376), .A2(n7591), .ZN(n9761) );
  OAI22_X1 U8998 ( .A1(n9713), .A2(n7377), .B1(n7500), .B2(n9697), .ZN(n7378)
         );
  AOI21_X1 U8999 ( .B1(n9426), .B2(n7363), .A(n7378), .ZN(n7379) );
  OAI21_X1 U9000 ( .B1(n9422), .B2(n9761), .A(n7379), .ZN(n7380) );
  AOI21_X1 U9001 ( .B1(n9765), .B2(n9713), .A(n7380), .ZN(n7381) );
  OAI21_X1 U9002 ( .B1(n7382), .B2(n9431), .A(n7381), .ZN(P1_U3284) );
  INV_X1 U9003 ( .A(n7383), .ZN(n7607) );
  NAND2_X1 U9004 ( .A1(n7607), .A2(n7606), .ZN(n7608) );
  NAND2_X1 U9005 ( .A1(n7608), .A2(n7384), .ZN(n7386) );
  INV_X1 U9006 ( .A(n7385), .ZN(n8866) );
  XNOR2_X1 U9007 ( .A(n7386), .B(n8866), .ZN(n9758) );
  INV_X1 U9008 ( .A(n9758), .ZN(n7396) );
  XNOR2_X1 U9009 ( .A(n7385), .B(n8867), .ZN(n7387) );
  OAI222_X1 U9010 ( .A1(n9702), .A2(n7615), .B1(n9703), .B2(n9676), .C1(n7387), 
        .C2(n9416), .ZN(n9756) );
  AND2_X1 U9011 ( .A1(n7601), .A2(n7358), .ZN(n7389) );
  OR2_X1 U9012 ( .A1(n7389), .A2(n7388), .ZN(n9755) );
  OAI22_X1 U9013 ( .A1(n9713), .A2(n7391), .B1(n7390), .B2(n9697), .ZN(n7392)
         );
  AOI21_X1 U9014 ( .B1(n9426), .B2(n7358), .A(n7392), .ZN(n7393) );
  OAI21_X1 U9015 ( .B1(n9177), .B2(n9755), .A(n7393), .ZN(n7394) );
  AOI21_X1 U9016 ( .B1(n9756), .B2(n9713), .A(n7394), .ZN(n7395) );
  OAI21_X1 U9017 ( .B1(n9431), .B2(n7396), .A(n7395), .ZN(P1_U3285) );
  INV_X1 U9018 ( .A(n7397), .ZN(n7398) );
  AOI211_X1 U9019 ( .C1(n7400), .C2(n7399), .A(n8814), .B(n7398), .ZN(n7405)
         );
  NAND2_X1 U9020 ( .A1(n8808), .A2(n9114), .ZN(n7402) );
  OAI211_X1 U9021 ( .C1(n9677), .C2(n8806), .A(n7402), .B(n7401), .ZN(n7404)
         );
  OAI22_X1 U9022 ( .A1(n9682), .A2(n8801), .B1(n8810), .B2(n9681), .ZN(n7403)
         );
  OR3_X1 U9023 ( .A1(n7405), .A2(n7404), .A3(n7403), .ZN(P1_U3228) );
  INV_X1 U9024 ( .A(n7406), .ZN(n7408) );
  OAI222_X1 U9025 ( .A1(P1_U3084), .A2(n5975), .B1(n9572), .B2(n7408), .C1(
        n7407), .C2(n9576), .ZN(P1_U3331) );
  OAI222_X1 U9026 ( .A1(n8587), .A2(n7409), .B1(n8583), .B2(n7408), .C1(n7017), 
        .C2(P2_U3152), .ZN(P2_U3336) );
  INV_X1 U9027 ( .A(n7416), .ZN(n8061) );
  OR2_X1 U9028 ( .A1(n7412), .A2(n8061), .ZN(n7413) );
  NOR2_X1 U9029 ( .A1(n7558), .A2(n5138), .ZN(n7430) );
  AND2_X1 U9030 ( .A1(n7558), .A2(n5138), .ZN(n7414) );
  OR2_X1 U9031 ( .A1(n7430), .A2(n7414), .ZN(n9853) );
  OAI21_X1 U9032 ( .B1(n7415), .B2(n5138), .A(n7433), .ZN(n7418) );
  OAI22_X1 U9033 ( .A1(n7416), .A2(n8402), .B1(n7556), .B2(n8404), .ZN(n7417)
         );
  AOI21_X1 U9034 ( .B1(n7418), .B2(n9786), .A(n7417), .ZN(n7419) );
  OAI21_X1 U9035 ( .B1(n9853), .B2(n7566), .A(n7419), .ZN(n9856) );
  NAND2_X1 U9036 ( .A1(n9856), .A2(n9798), .ZN(n7428) );
  INV_X1 U9037 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n7422) );
  INV_X1 U9038 ( .A(n7420), .ZN(n7421) );
  OAI22_X1 U9039 ( .A1(n9798), .A2(n7422), .B1(n8411), .B2(n7421), .ZN(n7426)
         );
  NAND2_X1 U9040 ( .A1(n7423), .A2(n7429), .ZN(n7424) );
  NAND2_X1 U9041 ( .A1(n7439), .A2(n7424), .ZN(n9855) );
  NOR2_X1 U9042 ( .A1(n9792), .A2(n9855), .ZN(n7425) );
  AOI211_X1 U9043 ( .C1(n8414), .C2(n7429), .A(n7426), .B(n7425), .ZN(n7427)
         );
  OAI211_X1 U9044 ( .C1(n9853), .C2(n8418), .A(n7428), .B(n7427), .ZN(P2_U3288) );
  NAND2_X1 U9045 ( .A1(n7429), .A2(n8060), .ZN(n7557) );
  INV_X1 U9046 ( .A(n7557), .ZN(n7559) );
  NOR2_X1 U9047 ( .A1(n7430), .A2(n7559), .ZN(n7431) );
  XNOR2_X1 U9048 ( .A(n7431), .B(n7563), .ZN(n8551) );
  NAND2_X1 U9049 ( .A1(n7433), .A2(n7432), .ZN(n7434) );
  XNOR2_X1 U9050 ( .A(n7434), .B(n7563), .ZN(n7437) );
  INV_X1 U9051 ( .A(n7435), .ZN(n8058) );
  AOI22_X1 U9052 ( .A1(n8058), .A2(n8425), .B1(n8423), .B2(n8060), .ZN(n7436)
         );
  OAI21_X1 U9053 ( .B1(n7437), .B2(n8399), .A(n7436), .ZN(n7438) );
  AOI21_X1 U9054 ( .B1(n8551), .B2(n8408), .A(n7438), .ZN(n8556) );
  AOI21_X1 U9055 ( .B1(n8552), .B2(n7439), .A(n7570), .ZN(n8554) );
  INV_X1 U9056 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n7441) );
  INV_X1 U9057 ( .A(n7454), .ZN(n7440) );
  OAI22_X1 U9058 ( .A1(n9798), .A2(n7441), .B1(n8411), .B2(n7440), .ZN(n7443)
         );
  INV_X1 U9059 ( .A(n8552), .ZN(n7457) );
  NOR2_X1 U9060 ( .A1(n9793), .A2(n7457), .ZN(n7442) );
  AOI211_X1 U9061 ( .C1(n8554), .C2(n8439), .A(n7443), .B(n7442), .ZN(n7445)
         );
  INV_X1 U9062 ( .A(n8418), .ZN(n7578) );
  NAND2_X1 U9063 ( .A1(n8551), .A2(n7578), .ZN(n7444) );
  OAI211_X1 U9064 ( .C1(n8556), .C2(n4262), .A(n7445), .B(n7444), .ZN(P2_U3287) );
  OAI21_X1 U9065 ( .B1(n7448), .B2(n7447), .A(n7446), .ZN(n7449) );
  NAND2_X1 U9066 ( .A1(n7449), .A2(n8033), .ZN(n7456) );
  NAND2_X1 U9067 ( .A1(n8035), .A2(n8058), .ZN(n7451) );
  OAI211_X1 U9068 ( .C1(n7452), .C2(n8039), .A(n7451), .B(n7450), .ZN(n7453)
         );
  AOI21_X1 U9069 ( .B1(n7454), .B2(n8042), .A(n7453), .ZN(n7455) );
  OAI211_X1 U9070 ( .C1(n7457), .C2(n8029), .A(n7456), .B(n7455), .ZN(P2_U3233) );
  OAI21_X1 U9071 ( .B1(n9426), .B2(n9670), .A(n7458), .ZN(n7461) );
  INV_X1 U9072 ( .A(n9697), .ZN(n9277) );
  AOI22_X1 U9073 ( .A1(n7459), .A2(n9713), .B1(P1_REG3_REG_0__SCAN_IN), .B2(
        n9277), .ZN(n7460) );
  OAI211_X1 U9074 ( .C1(n5950), .C2(n9713), .A(n7461), .B(n7460), .ZN(P1_U3291) );
  XNOR2_X1 U9075 ( .A(n7541), .B(P2_REG1_REG_10__SCAN_IN), .ZN(n7538) );
  XOR2_X1 U9076 ( .A(n7538), .B(n7539), .Z(n7472) );
  NAND2_X1 U9077 ( .A1(n8088), .A2(P2_ADDR_REG_10__SCAN_IN), .ZN(n7464) );
  OAI211_X1 U9078 ( .C1(n8165), .C2(n7537), .A(n7465), .B(n7464), .ZN(n7471)
         );
  XNOR2_X1 U9079 ( .A(n7541), .B(P2_REG2_REG_10__SCAN_IN), .ZN(n7468) );
  AOI211_X1 U9080 ( .C1(n7469), .C2(n7468), .A(n8163), .B(n7540), .ZN(n7470)
         );
  AOI211_X1 U9081 ( .C1(n8167), .C2(n7472), .A(n7471), .B(n7470), .ZN(n7473)
         );
  INV_X1 U9082 ( .A(n7473), .ZN(P2_U3255) );
  INV_X1 U9083 ( .A(n7474), .ZN(n7492) );
  OAI222_X1 U9084 ( .A1(n7476), .A2(P1_U3084), .B1(n9572), .B2(n7492), .C1(
        n7475), .C2(n9576), .ZN(P1_U3329) );
  XNOR2_X1 U9085 ( .A(n7477), .B(n9060), .ZN(n9734) );
  INV_X1 U9086 ( .A(n9734), .ZN(n7491) );
  NOR2_X1 U9087 ( .A1(n7478), .A2(n9694), .ZN(n9712) );
  NAND2_X1 U9088 ( .A1(n9713), .A2(n9712), .ZN(n9666) );
  NOR2_X1 U9089 ( .A1(n7479), .A2(n9060), .ZN(n9673) );
  AOI21_X1 U9090 ( .B1(n7479), .B2(n9060), .A(n9673), .ZN(n7482) );
  AOI22_X1 U9091 ( .A1(n9398), .A2(n9115), .B1(n9396), .B2(n6893), .ZN(n7481)
         );
  INV_X1 U9092 ( .A(n9710), .ZN(n7781) );
  NAND2_X1 U9093 ( .A1(n9734), .A2(n7781), .ZN(n7480) );
  OAI211_X1 U9094 ( .C1(n7482), .C2(n9416), .A(n7481), .B(n7480), .ZN(n9732)
         );
  NAND2_X1 U9095 ( .A1(n9732), .A2(n9713), .ZN(n7490) );
  OAI22_X1 U9096 ( .A1(n9713), .A2(n7483), .B1(P1_REG3_REG_3__SCAN_IN), .B2(
        n9697), .ZN(n7488) );
  INV_X1 U9097 ( .A(n9667), .ZN(n7486) );
  NAND2_X1 U9098 ( .A1(n9729), .A2(n7484), .ZN(n7485) );
  NAND2_X1 U9099 ( .A1(n7486), .A2(n7485), .ZN(n9731) );
  NOR2_X1 U9100 ( .A1(n9177), .A2(n9731), .ZN(n7487) );
  AOI211_X1 U9101 ( .C1(n9426), .C2(n9729), .A(n7488), .B(n7487), .ZN(n7489)
         );
  OAI211_X1 U9102 ( .C1(n7491), .C2(n9666), .A(n7490), .B(n7489), .ZN(P1_U3288) );
  OAI222_X1 U9103 ( .A1(n8587), .A2(n7494), .B1(P2_U3152), .B2(n7493), .C1(
        n8583), .C2(n7492), .ZN(P2_U3334) );
  XNOR2_X1 U9104 ( .A(n7496), .B(n7495), .ZN(n7503) );
  AOI21_X1 U9105 ( .B1(n8748), .B2(n9113), .A(n7497), .ZN(n7499) );
  NAND2_X1 U9106 ( .A1(n8808), .A2(n9111), .ZN(n7498) );
  OAI211_X1 U9107 ( .C1(n8810), .C2(n7500), .A(n7499), .B(n7498), .ZN(n7501)
         );
  AOI21_X1 U9108 ( .B1(n8812), .B2(n7363), .A(n7501), .ZN(n7502) );
  OAI21_X1 U9109 ( .B1(n7503), .B2(n8814), .A(n7502), .ZN(P1_U3211) );
  NAND2_X1 U9110 ( .A1(n7505), .A2(n7504), .ZN(n7507) );
  NAND2_X1 U9111 ( .A1(n7620), .A2(n8714), .ZN(n8873) );
  AND2_X2 U9112 ( .A1(n8871), .A2(n8873), .ZN(n9068) );
  NAND2_X1 U9113 ( .A1(n7620), .A2(n9111), .ZN(n7509) );
  OR2_X1 U9114 ( .A1(n8720), .A2(n9110), .ZN(n7510) );
  NAND2_X1 U9115 ( .A1(n8720), .A2(n9110), .ZN(n7511) );
  INV_X1 U9116 ( .A(n9069), .ZN(n7514) );
  XNOR2_X1 U9117 ( .A(n7665), .B(n7514), .ZN(n7678) );
  INV_X1 U9118 ( .A(n9068), .ZN(n7516) );
  INV_X1 U9119 ( .A(n8720), .ZN(n7657) );
  AND2_X1 U9120 ( .A1(n7657), .A2(n9110), .ZN(n8860) );
  NAND2_X1 U9121 ( .A1(n8720), .A2(n7518), .ZN(n8874) );
  OAI21_X1 U9122 ( .B1(n9069), .B2(n7517), .A(n7667), .ZN(n7520) );
  OAI22_X1 U9123 ( .A1(n7518), .A2(n9703), .B1(n9702), .B2(n8668), .ZN(n7519)
         );
  AOI21_X1 U9124 ( .B1(n7520), .B2(n9706), .A(n7519), .ZN(n7521) );
  OAI21_X1 U9125 ( .B1(n9710), .B2(n7678), .A(n7521), .ZN(n7680) );
  NAND2_X1 U9126 ( .A1(n7680), .A2(n9713), .ZN(n7526) );
  OAI22_X1 U9127 ( .A1(n9713), .A2(n7522), .B1(n8625), .B2(n9697), .ZN(n7524)
         );
  INV_X1 U9128 ( .A(n7513), .ZN(n8632) );
  INV_X1 U9129 ( .A(n7620), .ZN(n9769) );
  OAI211_X1 U9130 ( .C1(n8632), .C2(n7533), .A(n9737), .B(n7672), .ZN(n7679)
         );
  NOR2_X1 U9131 ( .A1(n7679), .A2(n9422), .ZN(n7523) );
  AOI211_X1 U9132 ( .C1(n9426), .C2(n7513), .A(n7524), .B(n7523), .ZN(n7525)
         );
  OAI211_X1 U9133 ( .C1(n7678), .C2(n9666), .A(n7526), .B(n7525), .ZN(P1_U3281) );
  INV_X1 U9134 ( .A(n8874), .ZN(n8863) );
  NOR2_X1 U9135 ( .A1(n8860), .A2(n8863), .ZN(n9070) );
  XNOR2_X1 U9136 ( .A(n7527), .B(n9070), .ZN(n7532) );
  INV_X1 U9137 ( .A(n7532), .ZN(n7658) );
  XNOR2_X1 U9138 ( .A(n7528), .B(n9070), .ZN(n7530) );
  AOI22_X1 U9139 ( .A1(n9396), .A2(n9111), .B1(n9398), .B2(n9109), .ZN(n7529)
         );
  OAI21_X1 U9140 ( .B1(n7530), .B2(n9416), .A(n7529), .ZN(n7531) );
  AOI21_X1 U9141 ( .B1(n7781), .B2(n7532), .A(n7531), .ZN(n7663) );
  AOI21_X1 U9142 ( .B1(n8720), .B2(n7590), .A(n7533), .ZN(n7661) );
  AOI22_X1 U9143 ( .A1(n7661), .A2(n9737), .B1(n9736), .B2(n8720), .ZN(n7534)
         );
  OAI211_X1 U9144 ( .C1(n9740), .C2(n7658), .A(n7663), .B(n7534), .ZN(n7551)
         );
  NAND2_X1 U9145 ( .A1(n7551), .A2(n9785), .ZN(n7535) );
  OAI21_X1 U9146 ( .B1(n9785), .B2(n6855), .A(n7535), .ZN(P1_U3532) );
  INV_X1 U9147 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n7536) );
  XOR2_X1 U9148 ( .A(P2_REG1_REG_11__SCAN_IN), .B(n7764), .Z(n7756) );
  XNOR2_X1 U9149 ( .A(n7757), .B(n7756), .ZN(n7550) );
  XOR2_X1 U9150 ( .A(n7764), .B(P2_REG2_REG_11__SCAN_IN), .Z(n7543) );
  OAI21_X1 U9151 ( .B1(n7543), .B2(n7542), .A(n7763), .ZN(n7544) );
  NAND2_X1 U9152 ( .A1(n7544), .A2(n8162), .ZN(n7549) );
  NOR2_X1 U9153 ( .A1(n8165), .A2(n7545), .ZN(n7546) );
  AOI211_X1 U9154 ( .C1(n8088), .C2(P2_ADDR_REG_11__SCAN_IN), .A(n7547), .B(
        n7546), .ZN(n7548) );
  OAI211_X1 U9155 ( .C1(n7550), .C2(n8117), .A(n7549), .B(n7548), .ZN(P2_U3256) );
  NAND2_X1 U9156 ( .A1(n7551), .A2(n9776), .ZN(n7552) );
  OAI21_X1 U9157 ( .B1(n9776), .B2(n6131), .A(n7552), .ZN(P1_U3481) );
  NAND2_X1 U9158 ( .A1(n7554), .A2(n7553), .ZN(n7555) );
  XOR2_X1 U9159 ( .A(n7646), .B(n7555), .Z(n7569) );
  OAI22_X1 U9160 ( .A1(n7556), .A2(n8402), .B1(n7627), .B2(n8404), .ZN(n7568)
         );
  NOR2_X1 U9161 ( .A1(n7560), .A2(n7559), .ZN(n7562) );
  NOR2_X1 U9162 ( .A1(n8552), .A2(n8059), .ZN(n7561) );
  AOI21_X1 U9163 ( .B1(n7563), .B2(n7562), .A(n7561), .ZN(n7564) );
  NOR2_X1 U9164 ( .A1(n7647), .A2(n7646), .ZN(n7687) );
  AND2_X1 U9165 ( .A1(n7647), .A2(n7646), .ZN(n7565) );
  NOR2_X1 U9166 ( .A1(n8550), .A2(n7566), .ZN(n7567) );
  AOI211_X1 U9167 ( .C1(n9786), .C2(n7569), .A(n7568), .B(n7567), .ZN(n8549)
         );
  INV_X1 U9168 ( .A(n7570), .ZN(n7571) );
  AOI21_X1 U9169 ( .B1(n8546), .B2(n7571), .A(n4259), .ZN(n8547) );
  INV_X1 U9170 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n7574) );
  INV_X1 U9171 ( .A(n7572), .ZN(n7573) );
  OAI22_X1 U9172 ( .A1(n9798), .A2(n7574), .B1(n8411), .B2(n7573), .ZN(n7577)
         );
  NOR2_X1 U9173 ( .A1(n9793), .A2(n7575), .ZN(n7576) );
  AOI211_X1 U9174 ( .C1(n8547), .C2(n8439), .A(n7577), .B(n7576), .ZN(n7581)
         );
  INV_X1 U9175 ( .A(n8550), .ZN(n7579) );
  NAND2_X1 U9176 ( .A1(n7579), .A2(n7578), .ZN(n7580) );
  OAI211_X1 U9177 ( .C1(n8549), .C2(n4262), .A(n7581), .B(n7580), .ZN(P2_U3286) );
  NAND2_X1 U9178 ( .A1(n7583), .A2(n9068), .ZN(n7584) );
  NAND2_X1 U9179 ( .A1(n7582), .A2(n7584), .ZN(n9766) );
  XNOR2_X1 U9180 ( .A(n7585), .B(n9068), .ZN(n7586) );
  NAND2_X1 U9181 ( .A1(n7586), .A2(n9706), .ZN(n7588) );
  AOI22_X1 U9182 ( .A1(n9396), .A2(n9112), .B1(n9398), .B2(n9110), .ZN(n7587)
         );
  OAI211_X1 U9183 ( .C1(n9766), .C2(n9710), .A(n7588), .B(n7587), .ZN(n9770)
         );
  NAND2_X1 U9184 ( .A1(n9770), .A2(n9713), .ZN(n7595) );
  OAI22_X1 U9185 ( .A1(n9713), .A2(n7589), .B1(n7618), .B2(n9697), .ZN(n7593)
         );
  OAI211_X1 U9186 ( .C1(n9769), .C2(n7591), .A(n9737), .B(n7590), .ZN(n9767)
         );
  NAND2_X1 U9187 ( .A1(n9713), .A2(n9694), .ZN(n9354) );
  NOR2_X1 U9188 ( .A1(n9767), .A2(n9354), .ZN(n7592) );
  AOI211_X1 U9189 ( .C1(n9426), .C2(n7620), .A(n7593), .B(n7592), .ZN(n7594)
         );
  OAI211_X1 U9190 ( .C1(n9766), .C2(n9666), .A(n7595), .B(n7594), .ZN(P1_U3283) );
  XNOR2_X1 U9191 ( .A(n7596), .B(n7606), .ZN(n7599) );
  AOI21_X1 U9192 ( .B1(n9396), .B2(n9115), .A(n7597), .ZN(n7598) );
  OAI21_X1 U9193 ( .B1(n7599), .B2(n9416), .A(n7598), .ZN(n9748) );
  INV_X1 U9194 ( .A(n9748), .ZN(n7612) );
  NAND2_X1 U9195 ( .A1(n9668), .A2(n7602), .ZN(n7600) );
  AND3_X1 U9196 ( .A1(n9737), .A2(n7601), .A3(n7600), .ZN(n9749) );
  INV_X1 U9197 ( .A(n7603), .ZN(n7604) );
  AOI22_X1 U9198 ( .A1(n9716), .A2(P1_REG2_REG_5__SCAN_IN), .B1(n7604), .B2(
        n9277), .ZN(n7605) );
  OAI21_X1 U9199 ( .B1(n9683), .B2(n4383), .A(n7605), .ZN(n7610) );
  NOR2_X1 U9200 ( .A1(n7607), .A2(n7606), .ZN(n9747) );
  INV_X1 U9201 ( .A(n7608), .ZN(n9746) );
  NOR3_X1 U9202 ( .A1(n9747), .A2(n9746), .A3(n9431), .ZN(n7609) );
  AOI211_X1 U9203 ( .C1(n9749), .C2(n9407), .A(n7610), .B(n7609), .ZN(n7611)
         );
  OAI21_X1 U9204 ( .B1(n9716), .B2(n7612), .A(n7611), .ZN(P1_U3286) );
  XNOR2_X1 U9205 ( .A(n8612), .B(n8613), .ZN(n7613) );
  XNOR2_X1 U9206 ( .A(n8616), .B(n7613), .ZN(n7622) );
  OAI21_X1 U9207 ( .B1(n8806), .B2(n7615), .A(n7614), .ZN(n7616) );
  AOI21_X1 U9208 ( .B1(n8808), .B2(n9110), .A(n7616), .ZN(n7617) );
  OAI21_X1 U9209 ( .B1(n8810), .B2(n7618), .A(n7617), .ZN(n7619) );
  AOI21_X1 U9210 ( .B1(n8812), .B2(n7620), .A(n7619), .ZN(n7621) );
  OAI21_X1 U9211 ( .B1(n7622), .B2(n8814), .A(n7621), .ZN(P1_U3219) );
  NAND2_X1 U9212 ( .A1(n4347), .A2(n7623), .ZN(n7624) );
  XNOR2_X1 U9213 ( .A(n7625), .B(n7624), .ZN(n7631) );
  INV_X1 U9214 ( .A(n7741), .ZN(n8055) );
  NAND2_X1 U9215 ( .A1(n8035), .A2(n8055), .ZN(n7626) );
  NAND2_X1 U9216 ( .A1(P2_U3152), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n7761) );
  OAI211_X1 U9217 ( .C1(n8039), .C2(n7627), .A(n7626), .B(n7761), .ZN(n7628)
         );
  AOI21_X1 U9218 ( .B1(n7730), .B2(n8042), .A(n7628), .ZN(n7630) );
  NAND2_X1 U9219 ( .A1(n8041), .A2(n8535), .ZN(n7629) );
  OAI211_X1 U9220 ( .C1(n7631), .C2(n8019), .A(n7630), .B(n7629), .ZN(P2_U3226) );
  INV_X1 U9221 ( .A(n7632), .ZN(n7636) );
  OAI222_X1 U9222 ( .A1(P1_U3084), .A2(n7634), .B1(n9572), .B2(n7636), .C1(
        n7633), .C2(n9576), .ZN(P1_U3328) );
  OAI222_X1 U9223 ( .A1(n8587), .A2(n7637), .B1(n8583), .B2(n7636), .C1(n7635), 
        .C2(P2_U3152), .ZN(P2_U3333) );
  OAI21_X1 U9224 ( .B1(n7639), .B2(n7743), .A(n7638), .ZN(n7640) );
  AOI222_X1 U9225 ( .A1(n9786), .A2(n7640), .B1(n8424), .B2(n8425), .C1(n8056), 
        .C2(n8423), .ZN(n8534) );
  XNOR2_X1 U9226 ( .A(n7747), .B(n8529), .ZN(n7641) );
  NOR2_X1 U9227 ( .A1(n7641), .A2(n5873), .ZN(n8528) );
  INV_X1 U9228 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n7791) );
  NAND2_X1 U9229 ( .A1(n8529), .A2(n8414), .ZN(n7643) );
  NAND2_X1 U9230 ( .A1(n9795), .A2(n7995), .ZN(n7642) );
  OAI211_X1 U9231 ( .C1(n9798), .C2(n7791), .A(n7643), .B(n7642), .ZN(n7644)
         );
  AOI21_X1 U9232 ( .B1(n8528), .B2(n7645), .A(n7644), .ZN(n7654) );
  INV_X1 U9233 ( .A(n7694), .ZN(n7648) );
  AND2_X1 U9234 ( .A1(n8546), .A2(n8058), .ZN(n7686) );
  AOI22_X1 U9235 ( .A1(n7648), .A2(n7686), .B1(n8540), .B2(n8057), .ZN(n7649)
         );
  INV_X1 U9236 ( .A(n7734), .ZN(n7651) );
  OR2_X1 U9237 ( .A1(n8535), .A2(n8056), .ZN(n7652) );
  OR2_X1 U9238 ( .A1(n7744), .A2(n7743), .ZN(n8531) );
  NAND2_X1 U9239 ( .A1(n7744), .A2(n7743), .ZN(n8530) );
  NAND3_X1 U9240 ( .A1(n8531), .A2(n8530), .A3(n8284), .ZN(n7653) );
  OAI211_X1 U9241 ( .C1(n8534), .C2(n4262), .A(n7654), .B(n7653), .ZN(P2_U3283) );
  INV_X1 U9242 ( .A(n8718), .ZN(n7655) );
  AOI22_X1 U9243 ( .A1(n9716), .A2(P1_REG2_REG_9__SCAN_IN), .B1(n7655), .B2(
        n9277), .ZN(n7656) );
  OAI21_X1 U9244 ( .B1(n7657), .B2(n9683), .A(n7656), .ZN(n7660) );
  NOR2_X1 U9245 ( .A1(n7658), .A2(n9666), .ZN(n7659) );
  AOI211_X1 U9246 ( .C1(n7661), .C2(n9670), .A(n7660), .B(n7659), .ZN(n7662)
         );
  OAI21_X1 U9247 ( .B1(n9716), .B2(n7663), .A(n7662), .ZN(P1_U3282) );
  OR2_X1 U9248 ( .A1(n7513), .A2(n9109), .ZN(n7664) );
  XNOR2_X1 U9249 ( .A(n7716), .B(n9108), .ZN(n8882) );
  XNOR2_X1 U9250 ( .A(n7666), .B(n8882), .ZN(n7715) );
  INV_X1 U9251 ( .A(n8882), .ZN(n9071) );
  XNOR2_X1 U9252 ( .A(n4345), .B(n9071), .ZN(n7669) );
  OAI22_X1 U9253 ( .A1(n8760), .A2(n9703), .B1(n9702), .B2(n8737), .ZN(n7668)
         );
  AOI21_X1 U9254 ( .B1(n7669), .B2(n9706), .A(n7668), .ZN(n7670) );
  OAI21_X1 U9255 ( .B1(n9710), .B2(n7715), .A(n7670), .ZN(n7718) );
  NAND2_X1 U9256 ( .A1(n7718), .A2(n9713), .ZN(n7677) );
  OAI22_X1 U9257 ( .A1(n9713), .A2(n7671), .B1(n8761), .B2(n9697), .ZN(n7675)
         );
  NAND2_X1 U9258 ( .A1(n7672), .A2(n7716), .ZN(n7673) );
  NAND2_X1 U9259 ( .A1(n7702), .A2(n7673), .ZN(n7717) );
  NOR2_X1 U9260 ( .A1(n7717), .A2(n9177), .ZN(n7674) );
  AOI211_X1 U9261 ( .C1(n9426), .C2(n7716), .A(n7675), .B(n7674), .ZN(n7676)
         );
  OAI211_X1 U9262 ( .C1(n7715), .C2(n9666), .A(n7677), .B(n7676), .ZN(P1_U3280) );
  INV_X1 U9263 ( .A(n9740), .ZN(n9773) );
  INV_X1 U9264 ( .A(n7678), .ZN(n7682) );
  OAI21_X1 U9265 ( .B1(n8632), .B2(n9768), .A(n7679), .ZN(n7681) );
  AOI211_X1 U9266 ( .C1(n9773), .C2(n7682), .A(n7681), .B(n7680), .ZN(n7685)
         );
  NAND2_X1 U9267 ( .A1(n9774), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n7683) );
  OAI21_X1 U9268 ( .B1(n7685), .B2(n9774), .A(n7683), .ZN(P1_U3484) );
  NAND2_X1 U9269 ( .A1(n9783), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n7684) );
  OAI21_X1 U9270 ( .B1(n7685), .B2(n9783), .A(n7684), .ZN(P1_U3533) );
  NOR2_X1 U9271 ( .A1(n7687), .A2(n7686), .ZN(n7688) );
  XNOR2_X1 U9272 ( .A(n7688), .B(n7694), .ZN(n8545) );
  INV_X1 U9273 ( .A(n7729), .ZN(n7689) );
  AOI21_X1 U9274 ( .B1(n8540), .B2(n7690), .A(n7689), .ZN(n8541) );
  AOI22_X1 U9275 ( .A1(n4262), .A2(P2_REG2_REG_11__SCAN_IN), .B1(n9795), .B2(
        n7691), .ZN(n7692) );
  OAI21_X1 U9276 ( .B1(n9793), .B2(n4406), .A(n7692), .ZN(n7697) );
  OAI21_X1 U9277 ( .B1(n7694), .B2(n7693), .A(n7725), .ZN(n7695) );
  AOI222_X1 U9278 ( .A1(n9786), .A2(n7695), .B1(n8058), .B2(n8423), .C1(n8056), 
        .C2(n8425), .ZN(n8543) );
  NOR2_X1 U9279 ( .A1(n8543), .A2(n4262), .ZN(n7696) );
  AOI211_X1 U9280 ( .C1(n8541), .C2(n8439), .A(n7697), .B(n7696), .ZN(n7698)
         );
  OAI21_X1 U9281 ( .B1(n8436), .B2(n8545), .A(n7698), .ZN(P2_U3285) );
  NAND2_X1 U9282 ( .A1(n7716), .A2(n8668), .ZN(n8889) );
  OR2_X1 U9283 ( .A1(n7716), .A2(n8668), .ZN(n7773) );
  NAND2_X1 U9284 ( .A1(n7774), .A2(n7773), .ZN(n7699) );
  OR2_X1 U9285 ( .A1(n8657), .A2(n8737), .ZN(n8890) );
  NAND2_X1 U9286 ( .A1(n8657), .A2(n8737), .ZN(n8967) );
  NAND2_X1 U9287 ( .A1(n8890), .A2(n8967), .ZN(n9073) );
  XNOR2_X1 U9288 ( .A(n7699), .B(n9073), .ZN(n7700) );
  AOI222_X1 U9289 ( .A1(n9706), .A2(n7700), .B1(n9108), .B2(n9396), .C1(n9106), 
        .C2(n9398), .ZN(n9542) );
  OAI22_X1 U9290 ( .A1(n9713), .A2(n7701), .B1(n8669), .B2(n9697), .ZN(n7706)
         );
  INV_X1 U9291 ( .A(n8657), .ZN(n7704) );
  INV_X1 U9292 ( .A(n7702), .ZN(n7703) );
  NOR2_X2 U9293 ( .A1(n7702), .A2(n8657), .ZN(n7782) );
  INV_X1 U9294 ( .A(n7782), .ZN(n7784) );
  OAI211_X1 U9295 ( .C1(n7704), .C2(n7703), .A(n7784), .B(n9737), .ZN(n9539)
         );
  NOR2_X1 U9296 ( .A1(n9539), .A2(n9422), .ZN(n7705) );
  AOI211_X1 U9297 ( .C1(n9426), .C2(n8657), .A(n7706), .B(n7705), .ZN(n7709)
         );
  OR2_X1 U9298 ( .A1(n7707), .A2(n9073), .ZN(n9538) );
  NAND2_X1 U9299 ( .A1(n7707), .A2(n9073), .ZN(n7772) );
  NAND3_X1 U9300 ( .A1(n9538), .A2(n7772), .A3(n9391), .ZN(n7708) );
  OAI211_X1 U9301 ( .C1(n9542), .C2(n9716), .A(n7709), .B(n7708), .ZN(P1_U3279) );
  INV_X1 U9302 ( .A(n7710), .ZN(n7713) );
  OAI222_X1 U9303 ( .A1(n8583), .A2(n7713), .B1(P2_U3152), .B2(n7711), .C1(
        n10015), .C2(n8587), .ZN(P2_U3332) );
  OAI222_X1 U9304 ( .A1(n7714), .A2(P1_U3084), .B1(n9572), .B2(n7713), .C1(
        n7712), .C2(n9576), .ZN(P1_U3327) );
  INV_X1 U9305 ( .A(n7715), .ZN(n7720) );
  INV_X1 U9306 ( .A(n7716), .ZN(n8766) );
  OAI22_X1 U9307 ( .A1(n7717), .A2(n9754), .B1(n8766), .B2(n9768), .ZN(n7719)
         );
  AOI211_X1 U9308 ( .C1(n9773), .C2(n7720), .A(n7719), .B(n7718), .ZN(n7723)
         );
  NAND2_X1 U9309 ( .A1(n9783), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n7721) );
  OAI21_X1 U9310 ( .B1(n7723), .B2(n9783), .A(n7721), .ZN(P1_U3534) );
  NAND2_X1 U9311 ( .A1(n9774), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n7722) );
  OAI21_X1 U9312 ( .B1(n7723), .B2(n9774), .A(n7722), .ZN(P1_U3487) );
  NAND2_X1 U9313 ( .A1(n7725), .A2(n7724), .ZN(n7726) );
  XNOR2_X1 U9314 ( .A(n7726), .B(n7735), .ZN(n7727) );
  AOI222_X1 U9315 ( .A1(n9786), .A2(n7727), .B1(n8055), .B2(n8425), .C1(n8057), 
        .C2(n8423), .ZN(n8538) );
  INV_X1 U9316 ( .A(n7747), .ZN(n7728) );
  AOI21_X1 U9317 ( .B1(n8535), .B2(n7729), .A(n7728), .ZN(n8536) );
  AOI22_X1 U9318 ( .A1(n4262), .A2(P2_REG2_REG_12__SCAN_IN), .B1(n9795), .B2(
        n7730), .ZN(n7731) );
  OAI21_X1 U9319 ( .B1(n9793), .B2(n4645), .A(n7731), .ZN(n7737) );
  INV_X1 U9320 ( .A(n7732), .ZN(n7733) );
  AOI21_X1 U9321 ( .B1(n7735), .B2(n7734), .A(n7733), .ZN(n8539) );
  NOR2_X1 U9322 ( .A1(n8539), .A2(n8436), .ZN(n7736) );
  AOI211_X1 U9323 ( .C1(n8536), .C2(n8439), .A(n7737), .B(n7736), .ZN(n7738)
         );
  OAI21_X1 U9324 ( .B1(n4262), .B2(n8538), .A(n7738), .ZN(P2_U3284) );
  XNOR2_X1 U9325 ( .A(n7739), .B(n7745), .ZN(n7740) );
  OAI222_X1 U9326 ( .A1(n8402), .A2(n7741), .B1(n8404), .B2(n8403), .C1(n8399), 
        .C2(n7740), .ZN(n8524) );
  INV_X1 U9327 ( .A(n8524), .ZN(n7755) );
  NAND2_X1 U9328 ( .A1(n8529), .A2(n8055), .ZN(n7742) );
  OAI21_X1 U9329 ( .B1(n7746), .B2(n7745), .A(n7822), .ZN(n8526) );
  INV_X1 U9330 ( .A(n7751), .ZN(n8522) );
  NOR2_X1 U9331 ( .A1(n7748), .A2(n8522), .ZN(n7749) );
  OR2_X1 U9332 ( .A1(n8428), .A2(n7749), .ZN(n8523) );
  INV_X1 U9333 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n9976) );
  OAI22_X1 U9334 ( .A1(n9798), .A2(n9976), .B1(n8411), .B2(n7813), .ZN(n7750)
         );
  AOI21_X1 U9335 ( .B1(n8414), .B2(n7751), .A(n7750), .ZN(n7752) );
  OAI21_X1 U9336 ( .B1(n8523), .B2(n9792), .A(n7752), .ZN(n7753) );
  AOI21_X1 U9337 ( .B1(n8526), .B2(n8284), .A(n7753), .ZN(n7754) );
  OAI21_X1 U9338 ( .B1(n7755), .B2(n4262), .A(n7754), .ZN(P2_U3282) );
  NOR2_X1 U9339 ( .A1(n7793), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n7795) );
  AOI21_X1 U9340 ( .B1(P2_REG1_REG_12__SCAN_IN), .B2(n7793), .A(n7795), .ZN(
        n7759) );
  AOI22_X1 U9341 ( .A1(n7757), .A2(n7756), .B1(n7764), .B2(
        P2_REG1_REG_11__SCAN_IN), .ZN(n7758) );
  NAND2_X1 U9342 ( .A1(n7758), .A2(n7759), .ZN(n7799) );
  OAI21_X1 U9343 ( .B1(n7759), .B2(n7758), .A(n7799), .ZN(n7769) );
  NAND2_X1 U9344 ( .A1(n8088), .A2(P2_ADDR_REG_12__SCAN_IN), .ZN(n7760) );
  OAI211_X1 U9345 ( .C1(n8165), .C2(n7762), .A(n7761), .B(n7760), .ZN(n7768)
         );
  XNOR2_X1 U9346 ( .A(n7793), .B(P2_REG2_REG_12__SCAN_IN), .ZN(n7766) );
  AOI211_X1 U9347 ( .C1(n7766), .C2(n7765), .A(n8163), .B(n7792), .ZN(n7767)
         );
  AOI211_X1 U9348 ( .C1(n8167), .C2(n7769), .A(n7768), .B(n7767), .ZN(n7770)
         );
  INV_X1 U9349 ( .A(n7770), .ZN(P2_U3257) );
  NAND2_X1 U9350 ( .A1(n8657), .A2(n9107), .ZN(n7771) );
  OR2_X1 U9351 ( .A1(n9533), .A2(n9417), .ZN(n8894) );
  NAND2_X1 U9352 ( .A1(n9533), .A2(n9417), .ZN(n8966) );
  XNOR2_X1 U9353 ( .A(n7871), .B(n9076), .ZN(n7787) );
  OAI22_X1 U9354 ( .A1(n8846), .A2(n9702), .B1(n9703), .B2(n8737), .ZN(n7780)
         );
  NAND2_X1 U9355 ( .A1(n7775), .A2(n9076), .ZN(n7896) );
  INV_X1 U9356 ( .A(n9076), .ZN(n7776) );
  NAND3_X1 U9357 ( .A1(n7777), .A2(n8967), .A3(n7776), .ZN(n7778) );
  AOI21_X1 U9358 ( .B1(n7896), .B2(n7778), .A(n9416), .ZN(n7779) );
  AOI211_X1 U9359 ( .C1(n7787), .C2(n7781), .A(n7780), .B(n7779), .ZN(n9536)
         );
  INV_X1 U9360 ( .A(n9533), .ZN(n8743) );
  INV_X1 U9361 ( .A(n9419), .ZN(n7783) );
  AOI21_X1 U9362 ( .B1(n9533), .B2(n7784), .A(n7783), .ZN(n9534) );
  INV_X1 U9363 ( .A(n8738), .ZN(n7785) );
  AOI22_X1 U9364 ( .A1(n9716), .A2(P1_REG2_REG_13__SCAN_IN), .B1(n7785), .B2(
        n9277), .ZN(n7786) );
  OAI21_X1 U9365 ( .B1(n8743), .B2(n9683), .A(n7786), .ZN(n7789) );
  INV_X1 U9366 ( .A(n7787), .ZN(n9537) );
  NOR2_X1 U9367 ( .A1(n9537), .A2(n9666), .ZN(n7788) );
  AOI211_X1 U9368 ( .C1(n9534), .C2(n9670), .A(n7789), .B(n7788), .ZN(n7790)
         );
  OAI21_X1 U9369 ( .B1(n9716), .B2(n9536), .A(n7790), .ZN(P1_U3278) );
  XNOR2_X1 U9370 ( .A(n8072), .B(n7791), .ZN(n7794) );
  OAI21_X1 U9371 ( .B1(n7794), .B2(n4343), .A(n8074), .ZN(n7806) );
  INV_X1 U9372 ( .A(n7795), .ZN(n7798) );
  OR2_X1 U9373 ( .A1(n8072), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n8067) );
  NAND2_X1 U9374 ( .A1(n8072), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n7796) );
  NAND2_X1 U9375 ( .A1(n8067), .A2(n7796), .ZN(n7797) );
  INV_X1 U9376 ( .A(n8069), .ZN(n7801) );
  NAND3_X1 U9377 ( .A1(n7799), .A2(n7798), .A3(n7797), .ZN(n7800) );
  AOI21_X1 U9378 ( .B1(n7801), .B2(n7800), .A(n8117), .ZN(n7805) );
  NAND2_X1 U9379 ( .A1(P2_U3152), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n7991) );
  NAND2_X1 U9380 ( .A1(n8088), .A2(P2_ADDR_REG_13__SCAN_IN), .ZN(n7802) );
  OAI211_X1 U9381 ( .C1(n8165), .C2(n7803), .A(n7991), .B(n7802), .ZN(n7804)
         );
  AOI211_X1 U9382 ( .C1(n7806), .C2(n8162), .A(n7805), .B(n7804), .ZN(n7807)
         );
  INV_X1 U9383 ( .A(n7807), .ZN(P2_U3258) );
  INV_X1 U9384 ( .A(n7808), .ZN(n7818) );
  OAI222_X1 U9385 ( .A1(n9576), .A2(n10017), .B1(P1_U3084), .B2(n9172), .C1(
        n7818), .C2(n9572), .ZN(P1_U3326) );
  OAI21_X1 U9386 ( .B1(n7811), .B2(n7810), .A(n7809), .ZN(n7812) );
  NAND2_X1 U9387 ( .A1(n7812), .A2(n8033), .ZN(n7817) );
  INV_X1 U9388 ( .A(n8039), .ZN(n7953) );
  NOR2_X1 U9389 ( .A1(n8023), .A2(n7813), .ZN(n7815) );
  NAND2_X1 U9390 ( .A1(P2_U3152), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n8078) );
  OAI21_X1 U9391 ( .B1(n7950), .B2(n8403), .A(n8078), .ZN(n7814) );
  AOI211_X1 U9392 ( .C1(n7953), .C2(n8055), .A(n7815), .B(n7814), .ZN(n7816)
         );
  OAI211_X1 U9393 ( .C1(n8522), .C2(n8029), .A(n7817), .B(n7816), .ZN(P2_U3217) );
  OAI222_X1 U9394 ( .A1(n8587), .A2(n7820), .B1(n7819), .B2(P2_U3152), .C1(
        n8583), .C2(n7818), .ZN(P2_U3331) );
  NOR2_X1 U9395 ( .A1(n8517), .A2(n8054), .ZN(n8393) );
  INV_X1 U9396 ( .A(n7825), .ZN(n8426) );
  INV_X1 U9397 ( .A(n8498), .ZN(n8347) );
  NAND2_X1 U9398 ( .A1(n8487), .A2(n8337), .ZN(n7834) );
  INV_X1 U9399 ( .A(n8487), .ZN(n8318) );
  NAND2_X1 U9400 ( .A1(n8469), .A2(n7940), .ZN(n7836) );
  INV_X1 U9401 ( .A(n8466), .ZN(n8256) );
  NAND2_X1 U9402 ( .A1(n8256), .A2(n7974), .ZN(n7838) );
  INV_X1 U9403 ( .A(n8218), .ZN(n8051) );
  NAND2_X1 U9404 ( .A1(n8198), .A2(n8197), .ZN(n8184) );
  NOR3_X1 U9405 ( .A1(n8185), .A2(n8544), .A3(n8182), .ZN(n7840) );
  NAND2_X1 U9406 ( .A1(n8184), .A2(n7840), .ZN(n7852) );
  NAND2_X1 U9407 ( .A1(n8185), .A2(n9851), .ZN(n7841) );
  XNOR2_X1 U9408 ( .A(n7842), .B(n8185), .ZN(n7843) );
  AND2_X1 U9409 ( .A1(n7844), .A2(P2_B_REG_SCAN_IN), .ZN(n7845) );
  NOR2_X1 U9410 ( .A1(n8404), .A2(n7845), .ZN(n8173) );
  AOI22_X1 U9411 ( .A1(n8049), .A2(n8423), .B1(n8173), .B2(n8047), .ZN(n7846)
         );
  INV_X1 U9412 ( .A(n8482), .ZN(n8301) );
  AND2_X2 U9413 ( .A1(n8315), .A2(n8301), .ZN(n8296) );
  INV_X1 U9414 ( .A(n8476), .ZN(n8290) );
  INV_X1 U9415 ( .A(n8450), .ZN(n8209) );
  OR2_X2 U9416 ( .A1(n8208), .A2(n8189), .ZN(n8178) );
  NAND2_X1 U9417 ( .A1(n8208), .A2(n8189), .ZN(n7847) );
  NAND2_X1 U9418 ( .A1(n8189), .A2(n8553), .ZN(n7849) );
  NAND3_X1 U9419 ( .A1(n8185), .A2(n8182), .A3(n9851), .ZN(n7848) );
  OAI211_X1 U9420 ( .C1(n8192), .C2(n5873), .A(n7849), .B(n7848), .ZN(n7850)
         );
  NOR2_X4 U9421 ( .A1(n7854), .A2(n7853), .ZN(n9862) );
  MUX2_X1 U9422 ( .A(P2_REG0_REG_29__SCAN_IN), .B(n7855), .S(n9862), .Z(
        P2_U3517) );
  MUX2_X1 U9423 ( .A(n7855), .B(P2_REG1_REG_29__SCAN_IN), .S(n9871), .Z(
        P2_U3549) );
  INV_X1 U9424 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n7857) );
  INV_X1 U9425 ( .A(n8823), .ZN(n7913) );
  OAI222_X1 U9426 ( .A1(n9576), .A2(n7857), .B1(n9572), .B2(n7913), .C1(
        P1_U3084), .C2(n7856), .ZN(P1_U3323) );
  INV_X1 U9427 ( .A(n7858), .ZN(n7861) );
  INV_X1 U9428 ( .A(n7859), .ZN(n7860) );
  AOI21_X1 U9429 ( .B1(n8793), .B2(n7861), .A(n7860), .ZN(n7862) );
  OAI21_X1 U9430 ( .B1(n7863), .B2(n7862), .A(n8794), .ZN(n7869) );
  OAI22_X1 U9431 ( .A1(n8806), .A2(n7901), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n7864), .ZN(n7865) );
  AOI21_X1 U9432 ( .B1(n8808), .B2(n9214), .A(n7865), .ZN(n7866) );
  OAI21_X1 U9433 ( .B1(n9208), .B2(n8810), .A(n7866), .ZN(n7867) );
  AOI21_X1 U9434 ( .B1(n9462), .B2(n8812), .A(n7867), .ZN(n7868) );
  NAND2_X1 U9435 ( .A1(n7869), .A2(n7868), .ZN(P1_U3212) );
  OR2_X1 U9436 ( .A1(n9533), .A2(n9106), .ZN(n7870) );
  NAND2_X1 U9437 ( .A1(n9533), .A2(n9106), .ZN(n7872) );
  OR2_X1 U9438 ( .A1(n9530), .A2(n9397), .ZN(n7873) );
  NOR2_X1 U9439 ( .A1(n9524), .A2(n9387), .ZN(n7874) );
  OR2_X1 U9440 ( .A1(n9382), .A2(n8698), .ZN(n8858) );
  NAND2_X1 U9441 ( .A1(n9382), .A2(n8698), .ZN(n8952) );
  NAND2_X1 U9442 ( .A1(n8858), .A2(n8952), .ZN(n9077) );
  NAND2_X1 U9443 ( .A1(n9375), .A2(n9077), .ZN(n7876) );
  NAND2_X1 U9444 ( .A1(n9382), .A2(n9399), .ZN(n7875) );
  NAND2_X1 U9445 ( .A1(n7876), .A2(n7875), .ZN(n9360) );
  OR2_X1 U9446 ( .A1(n9514), .A2(n9386), .ZN(n7877) );
  NAND2_X1 U9447 ( .A1(n9357), .A2(n8640), .ZN(n8953) );
  OR2_X1 U9448 ( .A1(n9503), .A2(n9346), .ZN(n7878) );
  NAND2_X1 U9449 ( .A1(n9321), .A2(n7878), .ZN(n7880) );
  NAND2_X1 U9450 ( .A1(n9503), .A2(n9346), .ZN(n7879) );
  AND2_X1 U9451 ( .A1(n9498), .A2(n9324), .ZN(n7881) );
  NAND2_X1 U9452 ( .A1(n9492), .A2(n7882), .ZN(n9282) );
  INV_X1 U9453 ( .A(n9492), .ZN(n7883) );
  NAND2_X1 U9454 ( .A1(n9280), .A2(n8652), .ZN(n7884) );
  INV_X1 U9455 ( .A(n8652), .ZN(n9293) );
  NAND2_X1 U9456 ( .A1(n9472), .A2(n8796), .ZN(n8999) );
  NAND2_X1 U9457 ( .A1(n9225), .A2(n7901), .ZN(n7889) );
  OR2_X2 U9458 ( .A1(n9462), .A2(n7890), .ZN(n9012) );
  NAND2_X1 U9459 ( .A1(n9462), .A2(n7890), .ZN(n9005) );
  NAND2_X1 U9460 ( .A1(n4881), .A2(n4386), .ZN(n7891) );
  AND2_X2 U9461 ( .A1(n9377), .A2(n9368), .ZN(n9369) );
  INV_X1 U9462 ( .A(n9357), .ZN(n9509) );
  INV_X1 U9463 ( .A(n9503), .ZN(n9329) );
  NOR2_X2 U9464 ( .A1(n9315), .A2(n9492), .ZN(n9302) );
  AND2_X2 U9465 ( .A1(n9302), .A2(n9280), .ZN(n9274) );
  NAND2_X1 U9466 ( .A1(n9274), .A2(n9265), .ZN(n9247) );
  OR2_X2 U9467 ( .A1(n9247), .A2(n9477), .ZN(n9248) );
  AOI21_X1 U9468 ( .B1(n9455), .B2(n9206), .A(n9192), .ZN(n9456) );
  INV_X1 U9469 ( .A(n9455), .ZN(n7895) );
  INV_X1 U9470 ( .A(n7892), .ZN(n7893) );
  AOI22_X1 U9471 ( .A1(n9716), .A2(P1_REG2_REG_28__SCAN_IN), .B1(n7893), .B2(
        n9277), .ZN(n7894) );
  OAI21_X1 U9472 ( .B1(n7895), .B2(n9683), .A(n7894), .ZN(n7910) );
  NAND2_X1 U9473 ( .A1(n7896), .A2(n8966), .ZN(n9414) );
  XNOR2_X1 U9474 ( .A(n9530), .B(n8846), .ZN(n9413) );
  OR2_X1 U9475 ( .A1(n9530), .A2(n8846), .ZN(n8893) );
  NAND2_X1 U9476 ( .A1(n9524), .A2(n9418), .ZN(n8888) );
  OAI21_X2 U9477 ( .B1(n9394), .B2(n8845), .A(n8888), .ZN(n9385) );
  INV_X1 U9478 ( .A(n8952), .ZN(n8844) );
  NAND2_X1 U9479 ( .A1(n9514), .A2(n8784), .ZN(n8951) );
  OR2_X1 U9480 ( .A1(n9514), .A2(n8784), .ZN(n9339) );
  NAND2_X1 U9481 ( .A1(n8905), .A2(n9339), .ZN(n8851) );
  INV_X1 U9482 ( .A(n9346), .ZN(n7898) );
  OR2_X1 U9483 ( .A1(n9503), .A2(n7898), .ZN(n8942) );
  NAND2_X1 U9484 ( .A1(n9503), .A2(n7898), .ZN(n8981) );
  NAND2_X1 U9485 ( .A1(n9498), .A2(n4901), .ZN(n9053) );
  NAND2_X1 U9486 ( .A1(n9057), .A2(n9283), .ZN(n8948) );
  INV_X1 U9487 ( .A(n8948), .ZN(n7899) );
  NAND2_X1 U9488 ( .A1(n9487), .A2(n8652), .ZN(n9056) );
  NAND2_X1 U9489 ( .A1(n9477), .A2(n7900), .ZN(n9049) );
  NAND2_X1 U9490 ( .A1(n9482), .A2(n8833), .ZN(n9051) );
  NAND2_X1 U9491 ( .A1(n9049), .A2(n9051), .ZN(n8997) );
  INV_X2 U9492 ( .A(n9212), .ZN(n9204) );
  NAND2_X1 U9493 ( .A1(n9213), .A2(n9204), .ZN(n7902) );
  NAND2_X1 U9494 ( .A1(n7902), .A2(n4905), .ZN(n9185) );
  INV_X1 U9495 ( .A(n7903), .ZN(n7904) );
  NAND2_X1 U9496 ( .A1(n9185), .A2(n7904), .ZN(n7908) );
  NAND2_X1 U9497 ( .A1(n9105), .A2(n9398), .ZN(n7905) );
  NOR2_X1 U9498 ( .A1(n9458), .A2(n9716), .ZN(n7909) );
  AOI211_X1 U9499 ( .C1(n9456), .C2(n9670), .A(n7910), .B(n7909), .ZN(n7911)
         );
  OAI21_X1 U9500 ( .B1(n9460), .B2(n9431), .A(n7911), .ZN(P1_U3263) );
  OAI222_X1 U9501 ( .A1(n8587), .A2(n9963), .B1(n8583), .B2(n7913), .C1(n4523), 
        .C2(P2_U3152), .ZN(P2_U3328) );
  XNOR2_X1 U9502 ( .A(n7969), .B(n7968), .ZN(n7919) );
  AOI22_X1 U9503 ( .A1(n8280), .A2(n8035), .B1(P2_REG3_REG_23__SCAN_IN), .B2(
        P2_U3152), .ZN(n7915) );
  NAND2_X1 U9504 ( .A1(n8042), .A2(n8288), .ZN(n7914) );
  OAI211_X1 U9505 ( .C1(n7916), .C2(n8039), .A(n7915), .B(n7914), .ZN(n7917)
         );
  AOI21_X1 U9506 ( .B1(n8476), .B2(n8041), .A(n7917), .ZN(n7918) );
  OAI21_X1 U9507 ( .B1(n7919), .B2(n8019), .A(n7918), .ZN(P2_U3218) );
  OAI21_X1 U9508 ( .B1(n7922), .B2(n7921), .A(n7920), .ZN(n7923) );
  NAND2_X1 U9509 ( .A1(n7923), .A2(n8033), .ZN(n7927) );
  NAND2_X1 U9510 ( .A1(n8035), .A2(n8351), .ZN(n7924) );
  NAND2_X1 U9511 ( .A1(P2_U3152), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n8170) );
  OAI211_X1 U9512 ( .C1(n8039), .C2(n8053), .A(n7924), .B(n8170), .ZN(n7925)
         );
  AOI21_X1 U9513 ( .B1(n8345), .B2(n8042), .A(n7925), .ZN(n7926) );
  OAI211_X1 U9514 ( .C1(n8347), .C2(n8029), .A(n7927), .B(n7926), .ZN(P2_U3221) );
  XNOR2_X1 U9515 ( .A(n7928), .B(n7929), .ZN(n7935) );
  AOI22_X1 U9516 ( .A1(n8035), .A2(n8322), .B1(P2_REG3_REG_21__SCAN_IN), .B2(
        P2_U3152), .ZN(n7931) );
  NAND2_X1 U9517 ( .A1(n8042), .A2(n8316), .ZN(n7930) );
  OAI211_X1 U9518 ( .C1(n7932), .C2(n8039), .A(n7931), .B(n7930), .ZN(n7933)
         );
  AOI21_X1 U9519 ( .B1(n8487), .B2(n8041), .A(n7933), .ZN(n7934) );
  OAI21_X1 U9520 ( .B1(n7935), .B2(n8019), .A(n7934), .ZN(P2_U3225) );
  XOR2_X1 U9521 ( .A(n7937), .B(n7936), .Z(n7938) );
  XNOR2_X1 U9522 ( .A(n7939), .B(n7938), .ZN(n7945) );
  INV_X1 U9523 ( .A(n8253), .ZN(n7942) );
  OAI22_X1 U9524 ( .A1(n8218), .A2(n8404), .B1(n7940), .B2(n8402), .ZN(n8248)
         );
  AOI22_X1 U9525 ( .A1(n8248), .A2(n7961), .B1(P2_REG3_REG_25__SCAN_IN), .B2(
        P2_U3152), .ZN(n7941) );
  OAI21_X1 U9526 ( .B1(n7942), .B2(n8023), .A(n7941), .ZN(n7943) );
  AOI21_X1 U9527 ( .B1(n8466), .B2(n8041), .A(n7943), .ZN(n7944) );
  OAI21_X1 U9528 ( .B1(n7945), .B2(n8019), .A(n7944), .ZN(P2_U3227) );
  INV_X1 U9529 ( .A(n8512), .ZN(n7956) );
  OAI21_X1 U9530 ( .B1(n7948), .B2(n7947), .A(n7946), .ZN(n7949) );
  NAND2_X1 U9531 ( .A1(n7949), .A2(n8033), .ZN(n7955) );
  NOR2_X1 U9532 ( .A1(n8023), .A2(n8410), .ZN(n7952) );
  NAND2_X1 U9533 ( .A1(P2_U3152), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n8112) );
  OAI21_X1 U9534 ( .B1(n7950), .B2(n8405), .A(n8112), .ZN(n7951) );
  AOI211_X1 U9535 ( .C1(n7953), .C2(n8054), .A(n7952), .B(n7951), .ZN(n7954)
         );
  OAI211_X1 U9536 ( .C1(n7956), .C2(n8029), .A(n7955), .B(n7954), .ZN(P2_U3228) );
  XNOR2_X1 U9537 ( .A(n7958), .B(n7957), .ZN(n7965) );
  NAND2_X1 U9538 ( .A1(P2_U3152), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n8124) );
  OR2_X1 U9539 ( .A1(n8053), .A2(n8404), .ZN(n7960) );
  NAND2_X1 U9540 ( .A1(n8426), .A2(n8423), .ZN(n7959) );
  NAND2_X1 U9541 ( .A1(n7960), .A2(n7959), .ZN(n8386) );
  NAND2_X1 U9542 ( .A1(n7961), .A2(n8386), .ZN(n7962) );
  OAI211_X1 U9543 ( .C1(n8023), .C2(n8378), .A(n8124), .B(n7962), .ZN(n7963)
         );
  AOI21_X1 U9544 ( .B1(n8041), .B2(n8509), .A(n7963), .ZN(n7964) );
  OAI21_X1 U9545 ( .B1(n7965), .B2(n8019), .A(n7964), .ZN(P2_U3230) );
  INV_X1 U9546 ( .A(n7966), .ZN(n7967) );
  AOI21_X1 U9547 ( .B1(n7969), .B2(n7968), .A(n7967), .ZN(n7973) );
  XNOR2_X1 U9548 ( .A(n7971), .B(n7970), .ZN(n7972) );
  XNOR2_X1 U9549 ( .A(n7973), .B(n7972), .ZN(n7979) );
  NOR2_X1 U9550 ( .A1(n8023), .A2(n8272), .ZN(n7977) );
  INV_X1 U9551 ( .A(n7974), .ZN(n8267) );
  AOI22_X1 U9552 ( .A1(n8267), .A2(n8035), .B1(P2_REG3_REG_24__SCAN_IN), .B2(
        P2_U3152), .ZN(n7975) );
  OAI21_X1 U9553 ( .B1(n8308), .B2(n8039), .A(n7975), .ZN(n7976) );
  AOI211_X1 U9554 ( .C1(n8274), .C2(n8041), .A(n7977), .B(n7976), .ZN(n7978)
         );
  OAI21_X1 U9555 ( .B1(n7979), .B2(n8019), .A(n7978), .ZN(P2_U3231) );
  XNOR2_X1 U9556 ( .A(n7980), .B(n7981), .ZN(n7987) );
  NOR2_X1 U9557 ( .A1(n8023), .A2(n8331), .ZN(n7985) );
  AOI22_X1 U9558 ( .A1(n8035), .A2(n8337), .B1(P2_REG3_REG_20__SCAN_IN), .B2(
        P2_U3152), .ZN(n7982) );
  OAI21_X1 U9559 ( .B1(n7983), .B2(n8039), .A(n7982), .ZN(n7984) );
  AOI211_X1 U9560 ( .C1(n8492), .C2(n8041), .A(n7985), .B(n7984), .ZN(n7986)
         );
  OAI21_X1 U9561 ( .B1(n7987), .B2(n8019), .A(n7986), .ZN(P2_U3235) );
  XOR2_X1 U9562 ( .A(n7989), .B(n7988), .Z(n7990) );
  NAND2_X1 U9563 ( .A1(n7990), .A2(n8033), .ZN(n7999) );
  NAND2_X1 U9564 ( .A1(n8035), .A2(n8424), .ZN(n7992) );
  OAI211_X1 U9565 ( .C1(n8039), .C2(n7993), .A(n7992), .B(n7991), .ZN(n7994)
         );
  INV_X1 U9566 ( .A(n7994), .ZN(n7998) );
  NAND2_X1 U9567 ( .A1(n8529), .A2(n8041), .ZN(n7997) );
  NAND2_X1 U9568 ( .A1(n8042), .A2(n7995), .ZN(n7996) );
  NAND4_X1 U9569 ( .A1(n7999), .A2(n7998), .A3(n7997), .A4(n7996), .ZN(
        P2_U3236) );
  NAND2_X1 U9570 ( .A1(n8001), .A2(n8000), .ZN(n8005) );
  XNOR2_X1 U9571 ( .A(n8003), .B(n8002), .ZN(n8004) );
  XNOR2_X1 U9572 ( .A(n8005), .B(n8004), .ZN(n8010) );
  NOR2_X1 U9573 ( .A1(n8023), .A2(n8298), .ZN(n8008) );
  AOI22_X1 U9574 ( .A1(n8035), .A2(n8266), .B1(P2_REG3_REG_22__SCAN_IN), .B2(
        P2_U3152), .ZN(n8006) );
  OAI21_X1 U9575 ( .B1(n8307), .B2(n8039), .A(n8006), .ZN(n8007) );
  AOI211_X1 U9576 ( .C1(n8482), .C2(n8041), .A(n8008), .B(n8007), .ZN(n8009)
         );
  OAI21_X1 U9577 ( .B1(n8010), .B2(n8019), .A(n8009), .ZN(P2_U3237) );
  XNOR2_X1 U9578 ( .A(n8012), .B(n8011), .ZN(n8017) );
  NAND2_X1 U9579 ( .A1(n8035), .A2(n8367), .ZN(n8013) );
  NAND2_X1 U9580 ( .A1(P2_U3152), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n8141) );
  OAI211_X1 U9581 ( .C1(n8039), .C2(n8405), .A(n8013), .B(n8141), .ZN(n8015)
         );
  NOR2_X1 U9582 ( .A1(n8362), .A2(n8029), .ZN(n8014) );
  AOI211_X1 U9583 ( .C1(n8042), .C2(n8360), .A(n8015), .B(n8014), .ZN(n8016)
         );
  OAI21_X1 U9584 ( .B1(n8017), .B2(n8019), .A(n8016), .ZN(P2_U3240) );
  AOI21_X1 U9585 ( .B1(n8018), .B2(n8020), .A(n8019), .ZN(n8022) );
  NAND2_X1 U9586 ( .A1(n8022), .A2(n8021), .ZN(n8028) );
  NOR2_X1 U9587 ( .A1(n8023), .A2(n8239), .ZN(n8026) );
  AOI22_X1 U9588 ( .A1(n8050), .A2(n8425), .B1(n8267), .B2(n8423), .ZN(n8236)
         );
  NOR2_X1 U9589 ( .A1(n8236), .A2(n8024), .ZN(n8025) );
  AOI211_X1 U9590 ( .C1(P2_REG3_REG_26__SCAN_IN), .C2(P2_U3152), .A(n8026), 
        .B(n8025), .ZN(n8027) );
  OAI211_X1 U9591 ( .C1(n4652), .C2(n8029), .A(n8028), .B(n8027), .ZN(P2_U3242) );
  XNOR2_X1 U9592 ( .A(n4819), .B(n8030), .ZN(n8031) );
  XNOR2_X1 U9593 ( .A(n8032), .B(n8031), .ZN(n8034) );
  NAND2_X1 U9594 ( .A1(n8034), .A2(n8033), .ZN(n8046) );
  NAND2_X1 U9595 ( .A1(n8035), .A2(n8426), .ZN(n8037) );
  NAND2_X1 U9596 ( .A1(P2_U3152), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n8036) );
  OAI211_X1 U9597 ( .C1(n8039), .C2(n8038), .A(n8037), .B(n8036), .ZN(n8040)
         );
  INV_X1 U9598 ( .A(n8040), .ZN(n8045) );
  NAND2_X1 U9599 ( .A1(n8517), .A2(n8041), .ZN(n8044) );
  NAND2_X1 U9600 ( .A1(n8042), .A2(n8431), .ZN(n8043) );
  NAND4_X1 U9601 ( .A1(n8046), .A2(n8045), .A3(n8044), .A4(n8043), .ZN(
        P2_U3243) );
  MUX2_X1 U9602 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(n8047), .S(P2_U3966), .Z(
        P2_U3582) );
  MUX2_X1 U9603 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(n8048), .S(P2_U3966), .Z(
        P2_U3581) );
  MUX2_X1 U9604 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(n8049), .S(P2_U3966), .Z(
        P2_U3580) );
  MUX2_X1 U9605 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n8050), .S(P2_U3966), .Z(
        P2_U3579) );
  MUX2_X1 U9606 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(n8051), .S(P2_U3966), .Z(
        P2_U3578) );
  MUX2_X1 U9607 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n8267), .S(P2_U3966), .Z(
        P2_U3577) );
  MUX2_X1 U9608 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(n8280), .S(P2_U3966), .Z(
        P2_U3576) );
  MUX2_X1 U9609 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(n8266), .S(P2_U3966), .Z(
        P2_U3575) );
  MUX2_X1 U9610 ( .A(n8322), .B(P2_DATAO_REG_22__SCAN_IN), .S(n8052), .Z(
        P2_U3574) );
  MUX2_X1 U9611 ( .A(n8337), .B(P2_DATAO_REG_21__SCAN_IN), .S(n8052), .Z(
        P2_U3573) );
  MUX2_X1 U9612 ( .A(n8351), .B(P2_DATAO_REG_20__SCAN_IN), .S(n8052), .Z(
        P2_U3572) );
  MUX2_X1 U9613 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n8367), .S(P2_U3966), .Z(
        P2_U3571) );
  MUX2_X1 U9614 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(n7828), .S(P2_U3966), .Z(
        P2_U3570) );
  MUX2_X1 U9615 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n8366), .S(P2_U3966), .Z(
        P2_U3569) );
  MUX2_X1 U9616 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n8426), .S(P2_U3966), .Z(
        P2_U3568) );
  MUX2_X1 U9617 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(n8054), .S(P2_U3966), .Z(
        P2_U3567) );
  MUX2_X1 U9618 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(n8424), .S(P2_U3966), .Z(
        P2_U3566) );
  MUX2_X1 U9619 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(n8055), .S(P2_U3966), .Z(
        P2_U3565) );
  MUX2_X1 U9620 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(n8056), .S(P2_U3966), .Z(
        P2_U3564) );
  MUX2_X1 U9621 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(n8057), .S(P2_U3966), .Z(
        P2_U3563) );
  MUX2_X1 U9622 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(n8058), .S(P2_U3966), .Z(
        P2_U3562) );
  MUX2_X1 U9623 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(n8059), .S(P2_U3966), .Z(
        P2_U3561) );
  MUX2_X1 U9624 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(n8060), .S(P2_U3966), .Z(
        P2_U3560) );
  MUX2_X1 U9625 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(n8061), .S(P2_U3966), .Z(
        P2_U3559) );
  MUX2_X1 U9626 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(n8062), .S(P2_U3966), .Z(
        P2_U3558) );
  MUX2_X1 U9627 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(n8063), .S(P2_U3966), .Z(
        P2_U3557) );
  MUX2_X1 U9628 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(n8064), .S(P2_U3966), .Z(
        P2_U3556) );
  MUX2_X1 U9629 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(n8065), .S(P2_U3966), .Z(
        P2_U3555) );
  MUX2_X1 U9630 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(n8066), .S(P2_U3966), .Z(
        P2_U3554) );
  MUX2_X1 U9631 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(n4263), .S(P2_U3966), .Z(
        P2_U3553) );
  MUX2_X1 U9632 ( .A(P2_DATAO_REG_0__SCAN_IN), .B(n5760), .S(P2_U3966), .Z(
        P2_U3552) );
  INV_X1 U9633 ( .A(n8067), .ZN(n8068) );
  NOR2_X1 U9634 ( .A1(n8069), .A2(n8068), .ZN(n8071) );
  XNOR2_X1 U9635 ( .A(n8084), .B(P2_REG1_REG_14__SCAN_IN), .ZN(n8070) );
  NOR2_X1 U9636 ( .A1(n8071), .A2(n8070), .ZN(n8089) );
  AOI21_X1 U9637 ( .B1(n8071), .B2(n8070), .A(n8089), .ZN(n8082) );
  XNOR2_X1 U9638 ( .A(n8084), .B(n9976), .ZN(n8076) );
  OAI21_X1 U9639 ( .B1(n8076), .B2(n8075), .A(n8083), .ZN(n8077) );
  NAND2_X1 U9640 ( .A1(n8077), .A2(n8162), .ZN(n8081) );
  INV_X1 U9641 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n9964) );
  OAI21_X1 U9642 ( .B1(n8171), .B2(n9964), .A(n8078), .ZN(n8079) );
  AOI21_X1 U9643 ( .B1(n8164), .B2(n8084), .A(n8079), .ZN(n8080) );
  OAI211_X1 U9644 ( .C1(n8082), .C2(n8117), .A(n8081), .B(n8080), .ZN(P2_U3259) );
  INV_X1 U9645 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n8085) );
  OAI21_X1 U9646 ( .B1(n8086), .B2(n8085), .A(n8106), .ZN(n8096) );
  AND2_X1 U9647 ( .A1(P2_U3152), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n8087) );
  AOI21_X1 U9648 ( .B1(n8088), .B2(P2_ADDR_REG_15__SCAN_IN), .A(n8087), .ZN(
        n8094) );
  INV_X1 U9649 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n8090) );
  XNOR2_X1 U9650 ( .A(n8105), .B(n8098), .ZN(n8092) );
  NAND2_X1 U9651 ( .A1(P2_REG1_REG_15__SCAN_IN), .A2(n8092), .ZN(n8100) );
  OAI211_X1 U9652 ( .C1(n8092), .C2(P2_REG1_REG_15__SCAN_IN), .A(n8167), .B(
        n8100), .ZN(n8093) );
  OAI211_X1 U9653 ( .C1(n8165), .C2(n8105), .A(n8094), .B(n8093), .ZN(n8095)
         );
  AOI21_X1 U9654 ( .B1(n8162), .B2(n8096), .A(n8095), .ZN(n8097) );
  INV_X1 U9655 ( .A(n8097), .ZN(P2_U3260) );
  NAND2_X1 U9656 ( .A1(n8099), .A2(n8098), .ZN(n8101) );
  NAND2_X1 U9657 ( .A1(n8101), .A2(n8100), .ZN(n8103) );
  XNOR2_X1 U9658 ( .A(n8128), .B(P2_REG1_REG_16__SCAN_IN), .ZN(n8102) );
  AOI21_X1 U9659 ( .B1(n8103), .B2(n8102), .A(n8119), .ZN(n8118) );
  NAND2_X1 U9660 ( .A1(n8105), .A2(n8104), .ZN(n8107) );
  NAND2_X1 U9661 ( .A1(n8128), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n8108) );
  OAI21_X1 U9662 ( .B1(n8128), .B2(P2_REG2_REG_16__SCAN_IN), .A(n8108), .ZN(
        n8109) );
  AOI211_X1 U9663 ( .C1(n8110), .C2(n8109), .A(n8127), .B(n8163), .ZN(n8111)
         );
  INV_X1 U9664 ( .A(n8111), .ZN(n8116) );
  INV_X1 U9665 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n8113) );
  OAI21_X1 U9666 ( .B1(n8171), .B2(n8113), .A(n8112), .ZN(n8114) );
  AOI21_X1 U9667 ( .B1(n8164), .B2(n8128), .A(n8114), .ZN(n8115) );
  OAI211_X1 U9668 ( .C1(n8118), .C2(n8117), .A(n8116), .B(n8115), .ZN(P2_U3261) );
  INV_X1 U9669 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n8126) );
  INV_X1 U9670 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n9932) );
  XNOR2_X1 U9671 ( .A(n8144), .B(n9932), .ZN(n8123) );
  OR2_X1 U9672 ( .A1(n8128), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n8121) );
  INV_X1 U9673 ( .A(n8119), .ZN(n8120) );
  NAND2_X1 U9674 ( .A1(n8123), .A2(n8122), .ZN(n8136) );
  OAI211_X1 U9675 ( .C1(n8123), .C2(n8122), .A(n8167), .B(n8136), .ZN(n8125)
         );
  OAI211_X1 U9676 ( .C1(n8171), .C2(n8126), .A(n8125), .B(n8124), .ZN(n8133)
         );
  NAND2_X1 U9677 ( .A1(n8144), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n8129) );
  OAI21_X1 U9678 ( .B1(n8144), .B2(P2_REG2_REG_17__SCAN_IN), .A(n8129), .ZN(
        n8130) );
  AOI211_X1 U9679 ( .C1(n8131), .C2(n8130), .A(n8146), .B(n8163), .ZN(n8132)
         );
  AOI211_X1 U9680 ( .C1(n8164), .C2(n8144), .A(n8133), .B(n8132), .ZN(n8134)
         );
  INV_X1 U9681 ( .A(n8134), .ZN(P2_U3262) );
  INV_X1 U9682 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n10060) );
  OR2_X1 U9683 ( .A1(n8151), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n8157) );
  NAND2_X1 U9684 ( .A1(n8151), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n8135) );
  NAND2_X1 U9685 ( .A1(n8157), .A2(n8135), .ZN(n8139) );
  OAI21_X1 U9686 ( .B1(n9932), .B2(n8137), .A(n8136), .ZN(n8138) );
  AND2_X1 U9687 ( .A1(n8139), .A2(n8138), .ZN(n8140) );
  OAI21_X1 U9688 ( .B1(n8159), .B2(n8140), .A(n8167), .ZN(n8142) );
  OAI211_X1 U9689 ( .C1(n10060), .C2(n8171), .A(n8142), .B(n8141), .ZN(n8143)
         );
  AOI21_X1 U9690 ( .B1(n8151), .B2(n8164), .A(n8143), .ZN(n8150) );
  OAI21_X1 U9691 ( .B1(n8147), .B2(n5304), .A(n8154), .ZN(n8148) );
  NAND2_X1 U9692 ( .A1(n8162), .A2(n8148), .ZN(n8149) );
  NAND2_X1 U9693 ( .A1(n8150), .A2(n8149), .ZN(P2_U3263) );
  INV_X1 U9694 ( .A(n8151), .ZN(n8152) );
  NAND2_X1 U9695 ( .A1(n8153), .A2(n8152), .ZN(n8155) );
  NAND2_X1 U9696 ( .A1(n8155), .A2(n8154), .ZN(n8156) );
  INV_X1 U9697 ( .A(n8157), .ZN(n8158) );
  NOR2_X1 U9698 ( .A1(n8159), .A2(n8158), .ZN(n8160) );
  XNOR2_X1 U9699 ( .A(n8160), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n8168) );
  INV_X1 U9700 ( .A(n8168), .ZN(n8161) );
  NAND2_X1 U9701 ( .A1(n8165), .A2(n5587), .ZN(n8166) );
  AOI21_X1 U9702 ( .B1(n8168), .B2(n8167), .A(n8166), .ZN(n8169) );
  XNOR2_X1 U9703 ( .A(n8175), .B(n8172), .ZN(n8443) );
  NAND2_X1 U9704 ( .A1(n8174), .A2(n8173), .ZN(n8446) );
  NOR2_X1 U9705 ( .A1(n4262), .A2(n8446), .ZN(n8179) );
  NOR2_X1 U9706 ( .A1(n8175), .A2(n9793), .ZN(n8176) );
  AOI211_X1 U9707 ( .C1(n4262), .C2(P2_REG2_REG_31__SCAN_IN), .A(n8179), .B(
        n8176), .ZN(n8177) );
  OAI21_X1 U9708 ( .B1(n8443), .B2(n9792), .A(n8177), .ZN(P2_U3265) );
  XNOR2_X1 U9709 ( .A(n8178), .B(n8444), .ZN(n8447) );
  AOI21_X1 U9710 ( .B1(n4262), .B2(P2_REG2_REG_30__SCAN_IN), .A(n8179), .ZN(
        n8181) );
  NAND2_X1 U9711 ( .A1(n8444), .A2(n8414), .ZN(n8180) );
  OAI211_X1 U9712 ( .C1(n8447), .C2(n9792), .A(n8181), .B(n8180), .ZN(P2_U3266) );
  INV_X1 U9713 ( .A(n8182), .ZN(n8183) );
  NAND2_X1 U9714 ( .A1(n8184), .A2(n8183), .ZN(n8186) );
  XNOR2_X1 U9715 ( .A(n8186), .B(n8185), .ZN(n8187) );
  NAND2_X1 U9716 ( .A1(n8187), .A2(n8284), .ZN(n8196) );
  AOI22_X1 U9717 ( .A1(n8188), .A2(n9795), .B1(P2_REG2_REG_29__SCAN_IN), .B2(
        n4262), .ZN(n8191) );
  NAND2_X1 U9718 ( .A1(n8189), .A2(n8414), .ZN(n8190) );
  OAI211_X1 U9719 ( .C1(n8192), .C2(n9792), .A(n8191), .B(n8190), .ZN(n8193)
         );
  AOI21_X1 U9720 ( .B1(n8194), .B2(n9798), .A(n8193), .ZN(n8195) );
  NAND2_X1 U9721 ( .A1(n8196), .A2(n8195), .ZN(P2_U3267) );
  XNOR2_X1 U9722 ( .A(n8198), .B(n8197), .ZN(n8448) );
  INV_X1 U9723 ( .A(n8448), .ZN(n8215) );
  XNOR2_X1 U9724 ( .A(n8200), .B(n8197), .ZN(n8202) );
  INV_X1 U9725 ( .A(n8399), .ZN(n8201) );
  NAND2_X1 U9726 ( .A1(n8202), .A2(n8201), .ZN(n8207) );
  OAI22_X1 U9727 ( .A1(n8204), .A2(n8402), .B1(n8404), .B2(n8203), .ZN(n8205)
         );
  INV_X1 U9728 ( .A(n8205), .ZN(n8206) );
  NAND2_X1 U9729 ( .A1(n8207), .A2(n8206), .ZN(n8452) );
  OAI21_X1 U9730 ( .B1(n8225), .B2(n8209), .A(n8208), .ZN(n8449) );
  AOI22_X1 U9731 ( .A1(n8210), .A2(n9795), .B1(P2_REG2_REG_28__SCAN_IN), .B2(
        n4262), .ZN(n8212) );
  NAND2_X1 U9732 ( .A1(n8450), .A2(n8414), .ZN(n8211) );
  OAI211_X1 U9733 ( .C1(n8449), .C2(n9792), .A(n8212), .B(n8211), .ZN(n8213)
         );
  AOI21_X1 U9734 ( .B1(n8452), .B2(n9798), .A(n8213), .ZN(n8214) );
  OAI21_X1 U9735 ( .B1(n8215), .B2(n8436), .A(n8214), .ZN(P2_U3268) );
  NOR2_X1 U9736 ( .A1(n8223), .A2(n4869), .ZN(n8217) );
  AOI21_X1 U9737 ( .B1(n8233), .B2(n8217), .A(n8399), .ZN(n8221) );
  OAI22_X1 U9738 ( .A1(n8219), .A2(n8404), .B1(n8218), .B2(n8402), .ZN(n8220)
         );
  AOI21_X1 U9739 ( .B1(n8222), .B2(n8221), .A(n8220), .ZN(n8458) );
  XNOR2_X1 U9740 ( .A(n8224), .B(n8223), .ZN(n8454) );
  NAND2_X1 U9741 ( .A1(n8454), .A2(n8284), .ZN(n8231) );
  AOI21_X1 U9742 ( .B1(n8455), .B2(n4654), .A(n8225), .ZN(n8456) );
  AOI22_X1 U9743 ( .A1(n8226), .A2(n9795), .B1(P2_REG2_REG_27__SCAN_IN), .B2(
        n4262), .ZN(n8227) );
  OAI21_X1 U9744 ( .B1(n8228), .B2(n9793), .A(n8227), .ZN(n8229) );
  AOI21_X1 U9745 ( .B1(n8456), .B2(n8439), .A(n8229), .ZN(n8230) );
  OAI211_X1 U9746 ( .C1(n8458), .C2(n4262), .A(n8231), .B(n8230), .ZN(P2_U3269) );
  XNOR2_X1 U9747 ( .A(n8232), .B(n8235), .ZN(n8463) );
  AOI22_X1 U9748 ( .A1(n8462), .A2(n8414), .B1(n4262), .B2(
        P2_REG2_REG_26__SCAN_IN), .ZN(n8243) );
  OAI211_X1 U9749 ( .C1(n8235), .C2(n8234), .A(n8233), .B(n9786), .ZN(n8237)
         );
  AOI211_X1 U9750 ( .C1(n8462), .C2(n8251), .A(n5873), .B(n8238), .ZN(n8461)
         );
  INV_X1 U9751 ( .A(n8461), .ZN(n8240) );
  OAI22_X1 U9752 ( .A1(n8240), .A2(n5587), .B1(n8239), .B2(n8411), .ZN(n8241)
         );
  OAI21_X1 U9753 ( .B1(n8460), .B2(n8241), .A(n9798), .ZN(n8242) );
  OAI211_X1 U9754 ( .C1(n8463), .C2(n8436), .A(n8243), .B(n8242), .ZN(P2_U3270) );
  XNOR2_X1 U9755 ( .A(n8244), .B(n8246), .ZN(n8468) );
  OAI211_X1 U9756 ( .C1(n8247), .C2(n8246), .A(n8245), .B(n9786), .ZN(n8250)
         );
  INV_X1 U9757 ( .A(n8248), .ZN(n8249) );
  NAND2_X1 U9758 ( .A1(n8250), .A2(n8249), .ZN(n8464) );
  INV_X1 U9759 ( .A(n8251), .ZN(n8252) );
  AOI211_X1 U9760 ( .C1(n8466), .C2(n8270), .A(n5873), .B(n8252), .ZN(n8465)
         );
  NAND2_X1 U9761 ( .A1(n8465), .A2(n8382), .ZN(n8255) );
  AOI22_X1 U9762 ( .A1(n8253), .A2(n9795), .B1(P2_REG2_REG_25__SCAN_IN), .B2(
        n4262), .ZN(n8254) );
  OAI211_X1 U9763 ( .C1(n8256), .C2(n9793), .A(n8255), .B(n8254), .ZN(n8257)
         );
  AOI21_X1 U9764 ( .B1(n8464), .B2(n9798), .A(n8257), .ZN(n8258) );
  OAI21_X1 U9765 ( .B1(n8468), .B2(n8436), .A(n8258), .ZN(P2_U3271) );
  OAI21_X1 U9766 ( .B1(n8260), .B2(n8261), .A(n8259), .ZN(n8473) );
  INV_X1 U9767 ( .A(n8473), .ZN(n8278) );
  INV_X1 U9768 ( .A(n8279), .ZN(n8263) );
  OAI21_X1 U9769 ( .B1(n8263), .B2(n8262), .A(n8261), .ZN(n8265) );
  NAND3_X1 U9770 ( .A1(n8265), .A2(n9786), .A3(n8264), .ZN(n8269) );
  AOI22_X1 U9771 ( .A1(n8267), .A2(n8425), .B1(n8423), .B2(n8266), .ZN(n8268)
         );
  NAND2_X1 U9772 ( .A1(n8269), .A2(n8268), .ZN(n8472) );
  OAI21_X1 U9773 ( .B1(n8286), .B2(n8469), .A(n8270), .ZN(n8470) );
  OAI22_X1 U9774 ( .A1(n8411), .A2(n8272), .B1(n9798), .B2(n8271), .ZN(n8273)
         );
  AOI21_X1 U9775 ( .B1(n8274), .B2(n8414), .A(n8273), .ZN(n8275) );
  OAI21_X1 U9776 ( .B1(n8470), .B2(n9792), .A(n8275), .ZN(n8276) );
  AOI21_X1 U9777 ( .B1(n8472), .B2(n9798), .A(n8276), .ZN(n8277) );
  OAI21_X1 U9778 ( .B1(n8278), .B2(n8436), .A(n8277), .ZN(P2_U3272) );
  OAI21_X1 U9779 ( .B1(n4337), .B2(n8282), .A(n8279), .ZN(n8281) );
  AOI222_X1 U9780 ( .A1(n9786), .A2(n8281), .B1(n8322), .B2(n8423), .C1(n8280), 
        .C2(n8425), .ZN(n8479) );
  INV_X1 U9781 ( .A(n8481), .ZN(n8285) );
  NAND2_X1 U9782 ( .A1(n8283), .A2(n8282), .ZN(n8475) );
  NAND3_X1 U9783 ( .A1(n8285), .A2(n8284), .A3(n8475), .ZN(n8293) );
  INV_X1 U9784 ( .A(n8296), .ZN(n8287) );
  AOI21_X1 U9785 ( .B1(n8476), .B2(n8287), .A(n8286), .ZN(n8477) );
  AOI22_X1 U9786 ( .A1(n4262), .A2(P2_REG2_REG_23__SCAN_IN), .B1(n9795), .B2(
        n8288), .ZN(n8289) );
  OAI21_X1 U9787 ( .B1(n8290), .B2(n9793), .A(n8289), .ZN(n8291) );
  AOI21_X1 U9788 ( .B1(n8477), .B2(n8439), .A(n8291), .ZN(n8292) );
  OAI211_X1 U9789 ( .C1(n4262), .C2(n8479), .A(n8293), .B(n8292), .ZN(P2_U3273) );
  XNOR2_X1 U9790 ( .A(n8295), .B(n8294), .ZN(n8486) );
  INV_X1 U9791 ( .A(n8315), .ZN(n8297) );
  AOI21_X1 U9792 ( .B1(n8482), .B2(n8297), .A(n8296), .ZN(n8483) );
  INV_X1 U9793 ( .A(n8298), .ZN(n8299) );
  AOI22_X1 U9794 ( .A1(n4262), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n9795), .B2(
        n8299), .ZN(n8300) );
  OAI21_X1 U9795 ( .B1(n8301), .B2(n9793), .A(n8300), .ZN(n8312) );
  INV_X1 U9796 ( .A(n8302), .ZN(n8306) );
  AOI21_X1 U9797 ( .B1(n8320), .B2(n8304), .A(n8303), .ZN(n8305) );
  NOR3_X1 U9798 ( .A1(n8306), .A2(n8305), .A3(n8399), .ZN(n8310) );
  OAI22_X1 U9799 ( .A1(n8308), .A2(n8404), .B1(n8307), .B2(n8402), .ZN(n8309)
         );
  NOR2_X1 U9800 ( .A1(n8310), .A2(n8309), .ZN(n8485) );
  NOR2_X1 U9801 ( .A1(n8485), .A2(n4262), .ZN(n8311) );
  AOI211_X1 U9802 ( .C1(n8483), .C2(n8439), .A(n8312), .B(n8311), .ZN(n8313)
         );
  OAI21_X1 U9803 ( .B1(n8486), .B2(n8436), .A(n8313), .ZN(P2_U3274) );
  XOR2_X1 U9804 ( .A(n8314), .B(n8319), .Z(n8491) );
  AOI21_X1 U9805 ( .B1(n8487), .B2(n8329), .A(n8315), .ZN(n8488) );
  AOI22_X1 U9806 ( .A1(n4262), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n9795), .B2(
        n8316), .ZN(n8317) );
  OAI21_X1 U9807 ( .B1(n8318), .B2(n9793), .A(n8317), .ZN(n8325) );
  OAI21_X1 U9808 ( .B1(n8321), .B2(n5372), .A(n8320), .ZN(n8323) );
  AOI222_X1 U9809 ( .A1(n9786), .A2(n8323), .B1(n8322), .B2(n8425), .C1(n8351), 
        .C2(n8423), .ZN(n8490) );
  NOR2_X1 U9810 ( .A1(n8490), .A2(n4262), .ZN(n8324) );
  AOI211_X1 U9811 ( .C1(n8488), .C2(n8439), .A(n8325), .B(n8324), .ZN(n8326)
         );
  OAI21_X1 U9812 ( .B1(n8491), .B2(n8436), .A(n8326), .ZN(P2_U3275) );
  XNOR2_X1 U9813 ( .A(n8328), .B(n8327), .ZN(n8496) );
  INV_X1 U9814 ( .A(n8329), .ZN(n8330) );
  AOI21_X1 U9815 ( .B1(n8492), .B2(n8343), .A(n8330), .ZN(n8493) );
  INV_X1 U9816 ( .A(n8331), .ZN(n8332) );
  AOI22_X1 U9817 ( .A1(n4262), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n9795), .B2(
        n8332), .ZN(n8333) );
  OAI21_X1 U9818 ( .B1(n4658), .B2(n9793), .A(n8333), .ZN(n8340) );
  NAND2_X1 U9819 ( .A1(n8348), .A2(n8334), .ZN(n8336) );
  XNOR2_X1 U9820 ( .A(n8336), .B(n8335), .ZN(n8338) );
  AOI222_X1 U9821 ( .A1(n9786), .A2(n8338), .B1(n8367), .B2(n8423), .C1(n8337), 
        .C2(n8425), .ZN(n8495) );
  NOR2_X1 U9822 ( .A1(n8495), .A2(n4262), .ZN(n8339) );
  AOI211_X1 U9823 ( .C1(n8493), .C2(n8439), .A(n8340), .B(n8339), .ZN(n8341)
         );
  OAI21_X1 U9824 ( .B1(n8436), .B2(n8496), .A(n8341), .ZN(P2_U3276) );
  XOR2_X1 U9825 ( .A(n8342), .B(n8350), .Z(n8501) );
  INV_X1 U9826 ( .A(n8343), .ZN(n8344) );
  AOI211_X1 U9827 ( .C1(n8498), .C2(n8357), .A(n5873), .B(n8344), .ZN(n8497)
         );
  AOI22_X1 U9828 ( .A1(n4262), .A2(P2_REG2_REG_19__SCAN_IN), .B1(n9795), .B2(
        n8345), .ZN(n8346) );
  OAI21_X1 U9829 ( .B1(n8347), .B2(n9793), .A(n8346), .ZN(n8354) );
  OAI21_X1 U9830 ( .B1(n8350), .B2(n8349), .A(n8348), .ZN(n8352) );
  AOI222_X1 U9831 ( .A1(n9786), .A2(n8352), .B1(n8351), .B2(n8425), .C1(n7828), 
        .C2(n8423), .ZN(n8500) );
  NOR2_X1 U9832 ( .A1(n8500), .A2(n4262), .ZN(n8353) );
  AOI211_X1 U9833 ( .C1(n8497), .C2(n8382), .A(n8354), .B(n8353), .ZN(n8355)
         );
  OAI21_X1 U9834 ( .B1(n8501), .B2(n8436), .A(n8355), .ZN(P2_U3277) );
  XNOR2_X1 U9835 ( .A(n8356), .B(n8365), .ZN(n8506) );
  INV_X1 U9836 ( .A(n8376), .ZN(n8359) );
  INV_X1 U9837 ( .A(n8357), .ZN(n8358) );
  AOI21_X1 U9838 ( .B1(n8502), .B2(n8359), .A(n8358), .ZN(n8503) );
  AOI22_X1 U9839 ( .A1(n4262), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n9795), .B2(
        n8360), .ZN(n8361) );
  OAI21_X1 U9840 ( .B1(n8362), .B2(n9793), .A(n8361), .ZN(n8370) );
  OAI21_X1 U9841 ( .B1(n8365), .B2(n8364), .A(n8363), .ZN(n8368) );
  AOI222_X1 U9842 ( .A1(n9786), .A2(n8368), .B1(n8367), .B2(n8425), .C1(n8366), 
        .C2(n8423), .ZN(n8505) );
  NOR2_X1 U9843 ( .A1(n8505), .A2(n4262), .ZN(n8369) );
  AOI211_X1 U9844 ( .C1(n8503), .C2(n8439), .A(n8370), .B(n8369), .ZN(n8371)
         );
  OAI21_X1 U9845 ( .B1(n8506), .B2(n8436), .A(n8371), .ZN(P2_U3278) );
  OAI21_X1 U9846 ( .B1(n8374), .B2(n8373), .A(n8372), .ZN(n8375) );
  INV_X1 U9847 ( .A(n8375), .ZN(n8511) );
  AOI211_X1 U9848 ( .C1(n8509), .C2(n4269), .A(n5873), .B(n8376), .ZN(n8508)
         );
  INV_X1 U9849 ( .A(n8509), .ZN(n8377) );
  NOR2_X1 U9850 ( .A1(n8377), .A2(n9793), .ZN(n8381) );
  INV_X1 U9851 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n8379) );
  OAI22_X1 U9852 ( .A1(n9798), .A2(n8379), .B1(n8411), .B2(n8378), .ZN(n8380)
         );
  AOI211_X1 U9853 ( .C1(n8508), .C2(n8382), .A(n8381), .B(n8380), .ZN(n8391)
         );
  NAND2_X1 U9854 ( .A1(n8383), .A2(n9786), .ZN(n8389) );
  AOI21_X1 U9855 ( .B1(n8401), .B2(n8385), .A(n8384), .ZN(n8388) );
  INV_X1 U9856 ( .A(n8386), .ZN(n8387) );
  OAI21_X1 U9857 ( .B1(n8389), .B2(n8388), .A(n8387), .ZN(n8507) );
  NAND2_X1 U9858 ( .A1(n8507), .A2(n9798), .ZN(n8390) );
  OAI211_X1 U9859 ( .C1(n8511), .C2(n8436), .A(n8391), .B(n8390), .ZN(P2_U3279) );
  AOI21_X1 U9860 ( .B1(n8435), .B2(n8422), .A(n8393), .ZN(n8394) );
  NOR2_X1 U9861 ( .A1(n8394), .A2(n8398), .ZN(n8395) );
  INV_X1 U9862 ( .A(n8516), .ZN(n8409) );
  NAND2_X1 U9863 ( .A1(n8397), .A2(n8398), .ZN(n8400) );
  AOI21_X1 U9864 ( .B1(n8401), .B2(n8400), .A(n8399), .ZN(n8407) );
  OAI22_X1 U9865 ( .A1(n8405), .A2(n8404), .B1(n8403), .B2(n8402), .ZN(n8406)
         );
  AOI211_X1 U9866 ( .C1(n8409), .C2(n8408), .A(n8407), .B(n8406), .ZN(n8515)
         );
  INV_X1 U9867 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n8412) );
  OAI22_X1 U9868 ( .A1(n9798), .A2(n8412), .B1(n8411), .B2(n8410), .ZN(n8413)
         );
  AOI21_X1 U9869 ( .B1(n8512), .B2(n8414), .A(n8413), .ZN(n8417) );
  NAND2_X1 U9870 ( .A1(n8430), .A2(n8512), .ZN(n8415) );
  AND2_X1 U9871 ( .A1(n4269), .A2(n8415), .ZN(n8513) );
  NAND2_X1 U9872 ( .A1(n8513), .A2(n8439), .ZN(n8416) );
  OAI211_X1 U9873 ( .C1(n8516), .C2(n8418), .A(n8417), .B(n8416), .ZN(n8419)
         );
  INV_X1 U9874 ( .A(n8419), .ZN(n8420) );
  OAI21_X1 U9875 ( .B1(n8515), .B2(n4262), .A(n8420), .ZN(P2_U3280) );
  XNOR2_X1 U9876 ( .A(n8421), .B(n8422), .ZN(n8427) );
  AOI222_X1 U9877 ( .A1(n9786), .A2(n8427), .B1(n8426), .B2(n8425), .C1(n8424), 
        .C2(n8423), .ZN(n8520) );
  OR2_X1 U9878 ( .A1(n8428), .A2(n8433), .ZN(n8429) );
  AND2_X1 U9879 ( .A1(n8430), .A2(n8429), .ZN(n8518) );
  AOI22_X1 U9880 ( .A1(n4262), .A2(P2_REG2_REG_15__SCAN_IN), .B1(n9795), .B2(
        n8431), .ZN(n8432) );
  OAI21_X1 U9881 ( .B1(n8433), .B2(n9793), .A(n8432), .ZN(n8438) );
  XNOR2_X1 U9882 ( .A(n8435), .B(n8434), .ZN(n8521) );
  NOR2_X1 U9883 ( .A1(n8521), .A2(n8436), .ZN(n8437) );
  AOI211_X1 U9884 ( .C1(n8518), .C2(n8439), .A(n8438), .B(n8437), .ZN(n8440)
         );
  OAI21_X1 U9885 ( .B1(n4262), .B2(n8520), .A(n8440), .ZN(P2_U3281) );
  NAND2_X1 U9886 ( .A1(n8441), .A2(n8553), .ZN(n8442) );
  OAI211_X1 U9887 ( .C1(n8443), .C2(n5873), .A(n8442), .B(n8446), .ZN(n8558)
         );
  MUX2_X1 U9888 ( .A(P2_REG1_REG_31__SCAN_IN), .B(n8558), .S(n9870), .Z(
        P2_U3551) );
  NAND2_X1 U9889 ( .A1(n8444), .A2(n8553), .ZN(n8445) );
  OAI211_X1 U9890 ( .C1(n8447), .C2(n5873), .A(n8446), .B(n8445), .ZN(n8559)
         );
  MUX2_X1 U9891 ( .A(P2_REG1_REG_30__SCAN_IN), .B(n8559), .S(n9870), .Z(
        P2_U3550) );
  NAND2_X1 U9892 ( .A1(n8448), .A2(n9851), .ZN(n8453) );
  NOR2_X1 U9893 ( .A1(n8449), .A2(n5873), .ZN(n8451) );
  MUX2_X1 U9894 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n8560), .S(n9870), .Z(
        P2_U3548) );
  NAND2_X1 U9895 ( .A1(n8454), .A2(n9851), .ZN(n8459) );
  AOI22_X1 U9896 ( .A1(n8456), .A2(n9811), .B1(n8553), .B2(n8455), .ZN(n8457)
         );
  NAND3_X1 U9897 ( .A1(n8459), .A2(n8458), .A3(n8457), .ZN(n8561) );
  MUX2_X1 U9898 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n8561), .S(n9870), .Z(
        P2_U3547) );
  MUX2_X1 U9899 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n8562), .S(n9870), .Z(
        P2_U3546) );
  AOI211_X1 U9900 ( .C1(n8553), .C2(n8466), .A(n8465), .B(n8464), .ZN(n8467)
         );
  OAI21_X1 U9901 ( .B1(n8468), .B2(n8544), .A(n8467), .ZN(n8563) );
  MUX2_X1 U9902 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n8563), .S(n9870), .Z(
        P2_U3545) );
  OAI22_X1 U9903 ( .A1(n8470), .A2(n5873), .B1(n9854), .B2(n8469), .ZN(n8471)
         );
  AOI211_X1 U9904 ( .C1(n8473), .C2(n9851), .A(n8472), .B(n8471), .ZN(n8474)
         );
  INV_X1 U9905 ( .A(n8474), .ZN(n8564) );
  MUX2_X1 U9906 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n8564), .S(n9870), .Z(
        P2_U3544) );
  NAND2_X1 U9907 ( .A1(n8475), .A2(n9851), .ZN(n8480) );
  AOI22_X1 U9908 ( .A1(n8477), .A2(n9811), .B1(n8553), .B2(n8476), .ZN(n8478)
         );
  OAI211_X1 U9909 ( .C1(n8481), .C2(n8480), .A(n8479), .B(n8478), .ZN(n8565)
         );
  MUX2_X1 U9910 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n8565), .S(n9870), .Z(
        P2_U3543) );
  AOI22_X1 U9911 ( .A1(n8483), .A2(n9811), .B1(n8553), .B2(n8482), .ZN(n8484)
         );
  OAI211_X1 U9912 ( .C1(n8486), .C2(n8544), .A(n8485), .B(n8484), .ZN(n8566)
         );
  MUX2_X1 U9913 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n8566), .S(n9870), .Z(
        P2_U3542) );
  AOI22_X1 U9914 ( .A1(n8488), .A2(n9811), .B1(n8553), .B2(n8487), .ZN(n8489)
         );
  OAI211_X1 U9915 ( .C1(n8491), .C2(n8544), .A(n8490), .B(n8489), .ZN(n8567)
         );
  MUX2_X1 U9916 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n8567), .S(n9870), .Z(
        P2_U3541) );
  AOI22_X1 U9917 ( .A1(n8493), .A2(n9811), .B1(n8553), .B2(n8492), .ZN(n8494)
         );
  OAI211_X1 U9918 ( .C1(n8496), .C2(n8544), .A(n8495), .B(n8494), .ZN(n8568)
         );
  MUX2_X1 U9919 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n8568), .S(n9870), .Z(
        P2_U3540) );
  AOI21_X1 U9920 ( .B1(n8553), .B2(n8498), .A(n8497), .ZN(n8499) );
  OAI211_X1 U9921 ( .C1(n8501), .C2(n8544), .A(n8500), .B(n8499), .ZN(n8569)
         );
  MUX2_X1 U9922 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n8569), .S(n9874), .Z(
        P2_U3539) );
  AOI22_X1 U9923 ( .A1(n8503), .A2(n9811), .B1(n8553), .B2(n8502), .ZN(n8504)
         );
  OAI211_X1 U9924 ( .C1(n8506), .C2(n8544), .A(n8505), .B(n8504), .ZN(n8570)
         );
  MUX2_X1 U9925 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n8570), .S(n9874), .Z(
        P2_U3538) );
  AOI211_X1 U9926 ( .C1(n8553), .C2(n8509), .A(n8508), .B(n8507), .ZN(n8510)
         );
  OAI21_X1 U9927 ( .B1(n8511), .B2(n8544), .A(n8510), .ZN(n8571) );
  MUX2_X1 U9928 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n8571), .S(n9874), .Z(
        P2_U3537) );
  AOI22_X1 U9929 ( .A1(n8513), .A2(n9811), .B1(n8553), .B2(n8512), .ZN(n8514)
         );
  OAI211_X1 U9930 ( .C1(n9818), .C2(n8516), .A(n8515), .B(n8514), .ZN(n8572)
         );
  MUX2_X1 U9931 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n8572), .S(n9874), .Z(
        P2_U3536) );
  AOI22_X1 U9932 ( .A1(n8518), .A2(n9811), .B1(n8553), .B2(n8517), .ZN(n8519)
         );
  OAI211_X1 U9933 ( .C1(n8521), .C2(n8544), .A(n8520), .B(n8519), .ZN(n8573)
         );
  MUX2_X1 U9934 ( .A(P2_REG1_REG_15__SCAN_IN), .B(n8573), .S(n9874), .Z(
        P2_U3535) );
  OAI22_X1 U9935 ( .A1(n8523), .A2(n5873), .B1(n9854), .B2(n8522), .ZN(n8525)
         );
  AOI211_X1 U9936 ( .C1(n9851), .C2(n8526), .A(n8525), .B(n8524), .ZN(n8527)
         );
  INV_X1 U9937 ( .A(n8527), .ZN(n8574) );
  MUX2_X1 U9938 ( .A(P2_REG1_REG_14__SCAN_IN), .B(n8574), .S(n9874), .Z(
        P2_U3534) );
  AOI21_X1 U9939 ( .B1(n8553), .B2(n8529), .A(n8528), .ZN(n8533) );
  NAND3_X1 U9940 ( .A1(n8531), .A2(n9851), .A3(n8530), .ZN(n8532) );
  NAND3_X1 U9941 ( .A1(n8534), .A2(n8533), .A3(n8532), .ZN(n8575) );
  MUX2_X1 U9942 ( .A(P2_REG1_REG_13__SCAN_IN), .B(n8575), .S(n9874), .Z(
        P2_U3533) );
  AOI22_X1 U9943 ( .A1(n8536), .A2(n9811), .B1(n8553), .B2(n8535), .ZN(n8537)
         );
  OAI211_X1 U9944 ( .C1(n8539), .C2(n8544), .A(n8538), .B(n8537), .ZN(n8576)
         );
  MUX2_X1 U9945 ( .A(P2_REG1_REG_12__SCAN_IN), .B(n8576), .S(n9874), .Z(
        P2_U3532) );
  AOI22_X1 U9946 ( .A1(n8541), .A2(n9811), .B1(n8553), .B2(n8540), .ZN(n8542)
         );
  OAI211_X1 U9947 ( .C1(n8545), .C2(n8544), .A(n8543), .B(n8542), .ZN(n8577)
         );
  MUX2_X1 U9948 ( .A(P2_REG1_REG_11__SCAN_IN), .B(n8577), .S(n9874), .Z(
        P2_U3531) );
  AOI22_X1 U9949 ( .A1(n8547), .A2(n9811), .B1(n8553), .B2(n8546), .ZN(n8548)
         );
  OAI211_X1 U9950 ( .C1(n9818), .C2(n8550), .A(n8549), .B(n8548), .ZN(n8578)
         );
  MUX2_X1 U9951 ( .A(P2_REG1_REG_10__SCAN_IN), .B(n8578), .S(n9874), .Z(
        P2_U3530) );
  INV_X1 U9952 ( .A(n8551), .ZN(n8557) );
  AOI22_X1 U9953 ( .A1(n8554), .A2(n9811), .B1(n8553), .B2(n8552), .ZN(n8555)
         );
  OAI211_X1 U9954 ( .C1(n8557), .C2(n9818), .A(n8556), .B(n8555), .ZN(n8579)
         );
  MUX2_X1 U9955 ( .A(P2_REG1_REG_9__SCAN_IN), .B(n8579), .S(n9874), .Z(
        P2_U3529) );
  MUX2_X1 U9956 ( .A(P2_REG0_REG_31__SCAN_IN), .B(n8558), .S(n9862), .Z(
        P2_U3519) );
  MUX2_X1 U9957 ( .A(P2_REG0_REG_30__SCAN_IN), .B(n8559), .S(n9862), .Z(
        P2_U3518) );
  MUX2_X1 U9958 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n8560), .S(n9862), .Z(
        P2_U3516) );
  MUX2_X1 U9959 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n8561), .S(n9862), .Z(
        P2_U3515) );
  MUX2_X1 U9960 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n8563), .S(n9862), .Z(
        P2_U3513) );
  MUX2_X1 U9961 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n8564), .S(n9862), .Z(
        P2_U3512) );
  MUX2_X1 U9962 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n8565), .S(n9862), .Z(
        P2_U3511) );
  MUX2_X1 U9963 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n8566), .S(n9862), .Z(
        P2_U3510) );
  MUX2_X1 U9964 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n8567), .S(n9862), .Z(
        P2_U3509) );
  MUX2_X1 U9965 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n8568), .S(n9862), .Z(
        P2_U3508) );
  MUX2_X1 U9966 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n8569), .S(n9862), .Z(
        P2_U3507) );
  MUX2_X1 U9967 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n8570), .S(n9862), .Z(
        P2_U3505) );
  MUX2_X1 U9968 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n8571), .S(n9862), .Z(
        P2_U3502) );
  MUX2_X1 U9969 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n8572), .S(n9862), .Z(
        P2_U3499) );
  MUX2_X1 U9970 ( .A(P2_REG0_REG_15__SCAN_IN), .B(n8573), .S(n9862), .Z(
        P2_U3496) );
  MUX2_X1 U9971 ( .A(P2_REG0_REG_14__SCAN_IN), .B(n8574), .S(n9862), .Z(
        P2_U3493) );
  MUX2_X1 U9972 ( .A(P2_REG0_REG_13__SCAN_IN), .B(n8575), .S(n9862), .Z(
        P2_U3490) );
  MUX2_X1 U9973 ( .A(P2_REG0_REG_12__SCAN_IN), .B(n8576), .S(n9862), .Z(
        P2_U3487) );
  MUX2_X1 U9974 ( .A(P2_REG0_REG_11__SCAN_IN), .B(n8577), .S(n9862), .Z(
        P2_U3484) );
  MUX2_X1 U9975 ( .A(P2_REG0_REG_10__SCAN_IN), .B(n8578), .S(n9862), .Z(
        P2_U3481) );
  MUX2_X1 U9976 ( .A(P2_REG0_REG_9__SCAN_IN), .B(n8579), .S(n9862), .Z(
        P2_U3478) );
  INV_X1 U9977 ( .A(n8819), .ZN(n9568) );
  NOR4_X1 U9978 ( .A1(n4504), .A2(P2_IR_REG_30__SCAN_IN), .A3(n4991), .A4(
        P2_U3152), .ZN(n8580) );
  AOI21_X1 U9979 ( .B1(n8581), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n8580), .ZN(
        n8582) );
  OAI21_X1 U9980 ( .B1(n9568), .B2(n8583), .A(n8582), .ZN(P2_U3327) );
  INV_X1 U9981 ( .A(n8816), .ZN(n9571) );
  INV_X1 U9982 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n8584) );
  OAI222_X1 U9983 ( .A1(n8583), .A2(n9571), .B1(P2_U3152), .B2(n8585), .C1(
        n8584), .C2(n8587), .ZN(P2_U3329) );
  INV_X1 U9984 ( .A(n8586), .ZN(n9573) );
  OAI222_X1 U9985 ( .A1(n8589), .A2(P2_U3152), .B1(n8583), .B2(n9573), .C1(
        n8588), .C2(n8587), .ZN(P2_U3330) );
  MUX2_X1 U9986 ( .A(n8590), .B(P2_IR_REG_0__SCAN_IN), .S(P2_STATE_REG_SCAN_IN), .Z(P2_U3358) );
  NOR2_X1 U9987 ( .A1(n8591), .A2(n4293), .ZN(n8593) );
  XNOR2_X1 U9988 ( .A(n8593), .B(n8592), .ZN(n8599) );
  OAI21_X1 U9989 ( .B1(n8806), .B2(n9417), .A(n8594), .ZN(n8595) );
  AOI21_X1 U9990 ( .B1(n8808), .B2(n9387), .A(n8595), .ZN(n8596) );
  OAI21_X1 U9991 ( .B1(n8810), .B2(n9424), .A(n8596), .ZN(n8597) );
  AOI21_X1 U9992 ( .B1(n9530), .B2(n8812), .A(n8597), .ZN(n8598) );
  OAI21_X1 U9993 ( .B1(n8599), .B2(n8814), .A(n8598), .ZN(P1_U3213) );
  INV_X1 U9994 ( .A(n8600), .ZN(n8601) );
  NAND2_X1 U9995 ( .A1(n8601), .A2(n8602), .ZN(n8675) );
  INV_X1 U9996 ( .A(n8602), .ZN(n8603) );
  NAND2_X1 U9997 ( .A1(n8600), .A2(n8603), .ZN(n8676) );
  NAND2_X1 U9998 ( .A1(n8675), .A2(n8676), .ZN(n8605) );
  INV_X1 U9999 ( .A(n8604), .ZN(n8674) );
  XNOR2_X1 U10000 ( .A(n8605), .B(n8674), .ZN(n8611) );
  INV_X1 U10001 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n8606) );
  OAI22_X1 U10002 ( .A1(n8806), .A2(n8652), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8606), .ZN(n8607) );
  AOI21_X1 U10003 ( .B1(n8808), .B2(n9268), .A(n8607), .ZN(n8608) );
  OAI21_X1 U10004 ( .B1(n8810), .B2(n9262), .A(n8608), .ZN(n8609) );
  AOI21_X1 U10005 ( .B1(n9482), .B2(n8812), .A(n8609), .ZN(n8610) );
  OAI21_X1 U10006 ( .B1(n8611), .B2(n8814), .A(n8610), .ZN(P1_U3214) );
  INV_X1 U10007 ( .A(n8613), .ZN(n8615) );
  OAI21_X1 U10008 ( .B1(n4762), .B2(n8613), .A(n8612), .ZN(n8614) );
  OAI21_X1 U10009 ( .B1(n8616), .B2(n8615), .A(n8614), .ZN(n8712) );
  OR2_X1 U10010 ( .A1(n8621), .A2(n8617), .ZN(n8713) );
  NOR2_X1 U10011 ( .A1(n8712), .A2(n8713), .ZN(n8711) );
  XNOR2_X1 U10012 ( .A(n8619), .B(n8618), .ZN(n8622) );
  INV_X1 U10013 ( .A(n8622), .ZN(n8620) );
  NOR3_X1 U10014 ( .A1(n8711), .A2(n8621), .A3(n8620), .ZN(n8624) );
  NOR2_X1 U10015 ( .A1(n8623), .A2(n8622), .ZN(n8756) );
  OAI21_X1 U10016 ( .B1(n8624), .B2(n8756), .A(n8794), .ZN(n8631) );
  INV_X1 U10017 ( .A(n8625), .ZN(n8629) );
  INV_X1 U10018 ( .A(n8810), .ZN(n8787) );
  INV_X1 U10019 ( .A(n8808), .ZN(n8651) );
  AOI21_X1 U10020 ( .B1(n8748), .B2(n9110), .A(n8626), .ZN(n8627) );
  OAI21_X1 U10021 ( .B1(n8651), .B2(n8668), .A(n8627), .ZN(n8628) );
  AOI21_X1 U10022 ( .B1(n8629), .B2(n8787), .A(n8628), .ZN(n8630) );
  OAI211_X1 U10023 ( .C1(n8632), .C2(n8801), .A(n8631), .B(n8630), .ZN(
        P1_U3215) );
  NOR2_X1 U10024 ( .A1(n8634), .A2(n8633), .ZN(n8639) );
  INV_X1 U10025 ( .A(n8636), .ZN(n8637) );
  NAND2_X1 U10026 ( .A1(n8635), .A2(n8637), .ZN(n8778) );
  NOR2_X1 U10027 ( .A1(n8635), .A2(n8637), .ZN(n8780) );
  AOI21_X1 U10028 ( .B1(n8781), .B2(n8778), .A(n8780), .ZN(n8638) );
  XOR2_X1 U10029 ( .A(n8639), .B(n8638), .Z(n8645) );
  NOR2_X1 U10030 ( .A1(n10029), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9170) );
  NOR2_X1 U10031 ( .A1(n8806), .A2(n8640), .ZN(n8641) );
  AOI211_X1 U10032 ( .C1(n9324), .C2(n8808), .A(n9170), .B(n8641), .ZN(n8642)
         );
  OAI21_X1 U10033 ( .B1(n8810), .B2(n9326), .A(n8642), .ZN(n8643) );
  AOI21_X1 U10034 ( .B1(n9503), .B2(n8812), .A(n8643), .ZN(n8644) );
  OAI21_X1 U10035 ( .B1(n8645), .B2(n8814), .A(n8644), .ZN(P1_U3217) );
  NAND2_X1 U10036 ( .A1(n4742), .A2(n8646), .ZN(n8647) );
  XNOR2_X1 U10037 ( .A(n8648), .B(n8647), .ZN(n8655) );
  AOI22_X1 U10038 ( .A1(n9324), .A2(n8748), .B1(P1_REG3_REG_21__SCAN_IN), .B2(
        P1_U3084), .ZN(n8650) );
  NAND2_X1 U10039 ( .A1(n8787), .A2(n9292), .ZN(n8649) );
  OAI211_X1 U10040 ( .C1(n8652), .C2(n8651), .A(n8650), .B(n8649), .ZN(n8653)
         );
  AOI21_X1 U10041 ( .B1(n9492), .B2(n8812), .A(n8653), .ZN(n8654) );
  OAI21_X1 U10042 ( .B1(n8655), .B2(n8814), .A(n8654), .ZN(P1_U3221) );
  INV_X1 U10043 ( .A(n8656), .ZN(n8693) );
  NAND2_X1 U10044 ( .A1(n8657), .A2(n9736), .ZN(n9541) );
  XNOR2_X1 U10045 ( .A(n8659), .B(n8658), .ZN(n8754) );
  NOR3_X1 U10046 ( .A1(n8756), .A2(n8755), .A3(n8754), .ZN(n8662) );
  INV_X1 U10047 ( .A(n8665), .ZN(n8661) );
  NAND2_X1 U10048 ( .A1(n8660), .A2(n8731), .ZN(n8663) );
  NOR3_X1 U10049 ( .A1(n8662), .A2(n8661), .A3(n8663), .ZN(n8734) );
  INV_X1 U10050 ( .A(n8662), .ZN(n8758) );
  INV_X1 U10051 ( .A(n8663), .ZN(n8664) );
  AOI21_X1 U10052 ( .B1(n8758), .B2(n8665), .A(n8664), .ZN(n8666) );
  OAI21_X1 U10053 ( .B1(n8734), .B2(n8666), .A(n8794), .ZN(n8673) );
  OAI21_X1 U10054 ( .B1(n8806), .B2(n8668), .A(n8667), .ZN(n8671) );
  NOR2_X1 U10055 ( .A1(n8810), .A2(n8669), .ZN(n8670) );
  AOI211_X1 U10056 ( .C1(n8808), .C2(n9106), .A(n8671), .B(n8670), .ZN(n8672)
         );
  OAI211_X1 U10057 ( .C1(n8693), .C2(n9541), .A(n8673), .B(n8672), .ZN(
        P1_U3222) );
  NOR2_X1 U10058 ( .A1(n8677), .A2(n8679), .ZN(n8704) );
  NOR2_X1 U10059 ( .A1(n4772), .A2(n8679), .ZN(n8680) );
  AOI21_X1 U10060 ( .B1(n8703), .B2(n8680), .A(n8792), .ZN(n8685) );
  AOI22_X1 U10061 ( .A1(n8748), .A2(n9268), .B1(P1_REG3_REG_25__SCAN_IN), .B2(
        P1_U3084), .ZN(n8682) );
  NAND2_X1 U10062 ( .A1(n8808), .A2(n9241), .ZN(n8681) );
  OAI211_X1 U10063 ( .C1(n8810), .C2(n9235), .A(n8682), .B(n8681), .ZN(n8683)
         );
  AOI21_X1 U10064 ( .B1(n9472), .B2(n8812), .A(n8683), .ZN(n8684) );
  OAI21_X1 U10065 ( .B1(n8685), .B2(n8814), .A(n8684), .ZN(P1_U3223) );
  NAND2_X1 U10066 ( .A1(n9382), .A2(n9736), .ZN(n9520) );
  OAI21_X1 U10067 ( .B1(n4281), .B2(n8687), .A(n8686), .ZN(n8688) );
  NAND2_X1 U10068 ( .A1(n8688), .A2(n8794), .ZN(n8692) );
  NAND2_X1 U10069 ( .A1(P1_U3084), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n9619) );
  OAI21_X1 U10070 ( .B1(n8806), .B2(n9418), .A(n9619), .ZN(n8690) );
  NOR2_X1 U10071 ( .A1(n8810), .A2(n9379), .ZN(n8689) );
  AOI211_X1 U10072 ( .C1(n8808), .C2(n9386), .A(n8690), .B(n8689), .ZN(n8691)
         );
  OAI211_X1 U10073 ( .C1(n8693), .C2(n9520), .A(n8692), .B(n8691), .ZN(
        P1_U3224) );
  OAI21_X1 U10074 ( .B1(n8696), .B2(n8695), .A(n8694), .ZN(n8697) );
  NAND2_X1 U10075 ( .A1(n8697), .A2(n8794), .ZN(n8702) );
  NAND2_X1 U10076 ( .A1(P1_U3084), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n9638) );
  OAI21_X1 U10077 ( .B1(n8806), .B2(n8698), .A(n9638), .ZN(n8700) );
  NOR2_X1 U10078 ( .A1(n8810), .A2(n9365), .ZN(n8699) );
  AOI211_X1 U10079 ( .C1(n8808), .C2(n9363), .A(n8700), .B(n8699), .ZN(n8701)
         );
  OAI211_X1 U10080 ( .C1(n9368), .C2(n8801), .A(n8702), .B(n8701), .ZN(
        P1_U3226) );
  NAND2_X1 U10081 ( .A1(n8705), .A2(n8794), .ZN(n8710) );
  OAI22_X1 U10082 ( .A1(n8806), .A2(n8833), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8706), .ZN(n8708) );
  NOR2_X1 U10083 ( .A1(n9250), .A2(n8810), .ZN(n8707) );
  AOI211_X1 U10084 ( .C1(n8808), .C2(n7887), .A(n8708), .B(n8707), .ZN(n8709)
         );
  OAI211_X1 U10085 ( .C1(n9253), .C2(n8801), .A(n8710), .B(n8709), .ZN(
        P1_U3227) );
  AOI21_X1 U10086 ( .B1(n8713), .B2(n8712), .A(n8711), .ZN(n8722) );
  NOR2_X1 U10087 ( .A1(n8806), .A2(n8714), .ZN(n8715) );
  AOI211_X1 U10088 ( .C1(n8808), .C2(n9109), .A(n8716), .B(n8715), .ZN(n8717)
         );
  OAI21_X1 U10089 ( .B1(n8810), .B2(n8718), .A(n8717), .ZN(n8719) );
  AOI21_X1 U10090 ( .B1(n8812), .B2(n8720), .A(n8719), .ZN(n8721) );
  OAI21_X1 U10091 ( .B1(n8722), .B2(n8814), .A(n8721), .ZN(P1_U3229) );
  NOR2_X1 U10092 ( .A1(n8723), .A2(n4341), .ZN(n8724) );
  XNOR2_X1 U10093 ( .A(n8725), .B(n8724), .ZN(n8730) );
  NAND2_X1 U10094 ( .A1(n9310), .A2(n8808), .ZN(n8727) );
  AOI22_X1 U10095 ( .A1(n9346), .A2(n8748), .B1(P1_REG3_REG_20__SCAN_IN), .B2(
        P1_U3084), .ZN(n8726) );
  OAI211_X1 U10096 ( .C1(n8810), .C2(n9313), .A(n8727), .B(n8726), .ZN(n8728)
         );
  AOI21_X1 U10097 ( .B1(n9498), .B2(n8812), .A(n8728), .ZN(n8729) );
  OAI21_X1 U10098 ( .B1(n8730), .B2(n8814), .A(n8729), .ZN(P1_U3231) );
  INV_X1 U10099 ( .A(n8731), .ZN(n8733) );
  NOR3_X1 U10100 ( .A1(n8734), .A2(n8733), .A3(n8732), .ZN(n8735) );
  OAI21_X1 U10101 ( .B1(n8735), .B2(n4344), .A(n8794), .ZN(n8742) );
  OAI21_X1 U10102 ( .B1(n8806), .B2(n8737), .A(n8736), .ZN(n8740) );
  NOR2_X1 U10103 ( .A1(n8810), .A2(n8738), .ZN(n8739) );
  AOI211_X1 U10104 ( .C1(n8808), .C2(n9397), .A(n8740), .B(n8739), .ZN(n8741)
         );
  OAI211_X1 U10105 ( .C1(n8743), .C2(n8801), .A(n8742), .B(n8741), .ZN(
        P1_U3232) );
  NAND2_X1 U10106 ( .A1(n8745), .A2(n8744), .ZN(n8747) );
  XNOR2_X1 U10107 ( .A(n8747), .B(n8746), .ZN(n8753) );
  AOI22_X1 U10108 ( .A1(n9310), .A2(n8748), .B1(P1_REG3_REG_22__SCAN_IN), .B2(
        P1_U3084), .ZN(n8750) );
  NAND2_X1 U10109 ( .A1(n8808), .A2(n9287), .ZN(n8749) );
  OAI211_X1 U10110 ( .C1(n9276), .C2(n8810), .A(n8750), .B(n8749), .ZN(n8751)
         );
  AOI21_X1 U10111 ( .B1(n9487), .B2(n8812), .A(n8751), .ZN(n8752) );
  OAI21_X1 U10112 ( .B1(n8753), .B2(n8814), .A(n8752), .ZN(P1_U3233) );
  OAI21_X1 U10113 ( .B1(n8756), .B2(n8755), .A(n8754), .ZN(n8757) );
  NAND3_X1 U10114 ( .A1(n8758), .A2(n8794), .A3(n8757), .ZN(n8765) );
  OAI21_X1 U10115 ( .B1(n8806), .B2(n8760), .A(n8759), .ZN(n8763) );
  NOR2_X1 U10116 ( .A1(n8810), .A2(n8761), .ZN(n8762) );
  AOI211_X1 U10117 ( .C1(n8808), .C2(n9107), .A(n8763), .B(n8762), .ZN(n8764)
         );
  OAI211_X1 U10118 ( .C1(n8766), .C2(n8801), .A(n8765), .B(n8764), .ZN(
        P1_U3234) );
  OAI21_X1 U10119 ( .B1(n8768), .B2(n7102), .A(n8767), .ZN(n8769) );
  NAND2_X1 U10120 ( .A1(n8769), .A2(n8794), .ZN(n8777) );
  NOR2_X1 U10121 ( .A1(n9703), .A2(n8770), .ZN(n8772) );
  AOI22_X1 U10122 ( .A1(n8808), .A2(n9116), .B1(n8772), .B2(n8771), .ZN(n8776)
         );
  AOI22_X1 U10123 ( .A1(n8812), .A2(n8774), .B1(n8773), .B2(
        P1_REG3_REG_2__SCAN_IN), .ZN(n8775) );
  NAND3_X1 U10124 ( .A1(n8777), .A2(n8776), .A3(n8775), .ZN(P1_U3235) );
  INV_X1 U10125 ( .A(n8778), .ZN(n8779) );
  NOR2_X1 U10126 ( .A1(n8780), .A2(n8779), .ZN(n8782) );
  XNOR2_X1 U10127 ( .A(n8782), .B(n8781), .ZN(n8789) );
  NAND2_X1 U10128 ( .A1(n8808), .A2(n9346), .ZN(n8783) );
  NAND2_X1 U10129 ( .A1(P1_U3084), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n9652) );
  OAI211_X1 U10130 ( .C1(n8784), .C2(n8806), .A(n8783), .B(n9652), .ZN(n8786)
         );
  NOR2_X1 U10131 ( .A1(n9509), .A2(n8801), .ZN(n8785) );
  AOI211_X1 U10132 ( .C1(n9349), .C2(n8787), .A(n8786), .B(n8785), .ZN(n8788)
         );
  OAI21_X1 U10133 ( .B1(n8789), .B2(n8814), .A(n8788), .ZN(P1_U3236) );
  OAI21_X1 U10134 ( .B1(n8792), .B2(n8791), .A(n8790), .ZN(n8795) );
  NAND3_X1 U10135 ( .A1(n8795), .A2(n8794), .A3(n8793), .ZN(n8800) );
  OAI22_X1 U10136 ( .A1(n8806), .A2(n8796), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n10036), .ZN(n8798) );
  NOR2_X1 U10137 ( .A1(n9222), .A2(n8810), .ZN(n8797) );
  AOI211_X1 U10138 ( .C1(n8808), .C2(n9228), .A(n8798), .B(n8797), .ZN(n8799)
         );
  OAI211_X1 U10139 ( .C1(n9225), .C2(n8801), .A(n8800), .B(n8799), .ZN(
        P1_U3238) );
  XNOR2_X1 U10140 ( .A(n8803), .B(n8802), .ZN(n8804) );
  XNOR2_X1 U10141 ( .A(n8805), .B(n8804), .ZN(n8815) );
  NAND2_X1 U10142 ( .A1(P1_U3084), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n9609) );
  OAI21_X1 U10143 ( .B1(n8806), .B2(n8846), .A(n9609), .ZN(n8807) );
  AOI21_X1 U10144 ( .B1(n8808), .B2(n9399), .A(n8807), .ZN(n8809) );
  OAI21_X1 U10145 ( .B1(n8810), .B2(n9401), .A(n8809), .ZN(n8811) );
  AOI21_X1 U10146 ( .B1(n9524), .B2(n8812), .A(n8811), .ZN(n8813) );
  OAI21_X1 U10147 ( .B1(n8815), .B2(n8814), .A(n8813), .ZN(P1_U3239) );
  NAND2_X1 U10148 ( .A1(n8816), .A2(n8822), .ZN(n8818) );
  NAND2_X1 U10149 ( .A1(n6003), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n8817) );
  NOR2_X1 U10150 ( .A1(n9198), .A2(n9105), .ZN(n8922) );
  NAND2_X1 U10151 ( .A1(n8819), .A2(n8822), .ZN(n8821) );
  NAND2_X1 U10152 ( .A1(n6003), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(n8820) );
  NAND2_X1 U10153 ( .A1(n8823), .A2(n8822), .ZN(n8826) );
  NAND2_X1 U10154 ( .A1(n8824), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n8825) );
  OR2_X1 U10155 ( .A1(n9179), .A2(n9187), .ZN(n8827) );
  OR2_X1 U10156 ( .A1(n9173), .A2(n9187), .ZN(n8828) );
  INV_X1 U10157 ( .A(n8919), .ZN(n8921) );
  INV_X1 U10158 ( .A(n9003), .ZN(n9048) );
  OAI21_X1 U10159 ( .B1(n8912), .B2(n9241), .A(n9048), .ZN(n8830) );
  INV_X1 U10160 ( .A(n8999), .ZN(n8913) );
  OAI21_X1 U10161 ( .B1(n8913), .B2(n9466), .A(n9047), .ZN(n8829) );
  MUX2_X1 U10162 ( .A(n8830), .B(n8829), .S(n8925), .Z(n8914) );
  NOR2_X1 U10163 ( .A1(n9049), .A2(n8927), .ZN(n8837) );
  INV_X1 U10164 ( .A(n9283), .ZN(n8831) );
  OR2_X1 U10165 ( .A1(n8831), .A2(n9053), .ZN(n8832) );
  NAND3_X1 U10166 ( .A1(n8832), .A2(n9056), .A3(n9282), .ZN(n8984) );
  NAND3_X1 U10167 ( .A1(n8984), .A2(n8925), .A3(n9057), .ZN(n8835) );
  NAND2_X1 U10168 ( .A1(n8925), .A2(n8833), .ZN(n8834) );
  OAI22_X1 U10169 ( .A1(n9052), .A2(n8835), .B1(n9265), .B2(n8834), .ZN(n8836)
         );
  AND2_X1 U10170 ( .A1(n9031), .A2(n9050), .ZN(n8843) );
  OAI21_X1 U10171 ( .B1(n8837), .B2(n8836), .A(n8843), .ZN(n8911) );
  INV_X1 U10172 ( .A(n9055), .ZN(n8839) );
  AND3_X1 U10173 ( .A1(n8839), .A2(n9283), .A3(n9057), .ZN(n8840) );
  NOR2_X1 U10174 ( .A1(n8908), .A2(n8840), .ZN(n8842) );
  INV_X1 U10175 ( .A(n9052), .ZN(n8950) );
  AOI21_X1 U10176 ( .B1(n8950), .B2(n9050), .A(n8925), .ZN(n8841) );
  NAND2_X1 U10177 ( .A1(n8981), .A2(n8953), .ZN(n8943) );
  NAND2_X1 U10178 ( .A1(n9339), .A2(n8951), .ZN(n9361) );
  OAI21_X1 U10179 ( .B1(n8844), .B2(n9361), .A(n8925), .ZN(n8850) );
  INV_X1 U10180 ( .A(n8845), .ZN(n8859) );
  XNOR2_X1 U10181 ( .A(n9524), .B(n9418), .ZN(n9395) );
  NAND4_X1 U10182 ( .A1(n8859), .A2(n8858), .A3(n9395), .A4(n8925), .ZN(n8849)
         );
  NAND2_X1 U10183 ( .A1(n8859), .A2(n8858), .ZN(n8963) );
  NAND2_X1 U10184 ( .A1(n9530), .A2(n8846), .ZN(n8887) );
  AND2_X1 U10185 ( .A1(n8966), .A2(n8887), .ZN(n8847) );
  NAND2_X1 U10186 ( .A1(n8893), .A2(n8925), .ZN(n8856) );
  OR3_X1 U10187 ( .A1(n8963), .A2(n8847), .A3(n8856), .ZN(n8848) );
  NAND3_X1 U10188 ( .A1(n8850), .A2(n8849), .A3(n8848), .ZN(n8852) );
  NAND2_X1 U10189 ( .A1(n8852), .A2(n4710), .ZN(n8901) );
  AND2_X1 U10190 ( .A1(n8953), .A2(n8951), .ZN(n8899) );
  NAND4_X1 U10191 ( .A1(n8952), .A2(n9395), .A3(n8927), .A4(n8888), .ZN(n8854)
         );
  NAND2_X1 U10192 ( .A1(n9361), .A2(n8927), .ZN(n8853) );
  OAI211_X1 U10193 ( .C1(n8858), .C2(n8925), .A(n8854), .B(n8853), .ZN(n8855)
         );
  NAND2_X1 U10194 ( .A1(n8899), .A2(n8855), .ZN(n8900) );
  INV_X1 U10195 ( .A(n8856), .ZN(n8857) );
  AND4_X1 U10196 ( .A1(n8859), .A2(n8858), .A3(n8857), .A4(n8894), .ZN(n8886)
         );
  INV_X1 U10197 ( .A(n8860), .ZN(n8876) );
  NAND3_X1 U10198 ( .A1(n8876), .A2(n8877), .A3(n8871), .ZN(n8964) );
  OR2_X1 U10199 ( .A1(n8867), .A2(n7385), .ZN(n8862) );
  AND2_X1 U10200 ( .A1(n8861), .A2(n8870), .ZN(n8956) );
  NAND2_X1 U10201 ( .A1(n8873), .A2(n8868), .ZN(n8959) );
  AOI21_X1 U10202 ( .B1(n8862), .B2(n8956), .A(n8959), .ZN(n8865) );
  NAND2_X1 U10203 ( .A1(n8877), .A2(n8863), .ZN(n8864) );
  OAI21_X1 U10204 ( .B1(n8964), .B2(n8865), .A(n8954), .ZN(n8881) );
  NAND2_X1 U10205 ( .A1(n8867), .A2(n8866), .ZN(n8869) );
  NAND3_X1 U10206 ( .A1(n8869), .A2(n9019), .A3(n8868), .ZN(n8872) );
  NAND3_X1 U10207 ( .A1(n8872), .A2(n8871), .A3(n8870), .ZN(n8875) );
  NAND3_X1 U10208 ( .A1(n8875), .A2(n8874), .A3(n8873), .ZN(n8878) );
  NAND2_X1 U10209 ( .A1(n8892), .A2(n8965), .ZN(n8884) );
  NAND2_X1 U10210 ( .A1(n8884), .A2(n8967), .ZN(n8885) );
  NAND2_X1 U10211 ( .A1(n8888), .A2(n8887), .ZN(n8972) );
  NOR2_X1 U10212 ( .A1(n8972), .A2(n8925), .ZN(n8898) );
  AND2_X1 U10213 ( .A1(n8967), .A2(n8889), .ZN(n8955) );
  INV_X1 U10214 ( .A(n8890), .ZN(n8891) );
  AOI21_X1 U10215 ( .B1(n8892), .B2(n8955), .A(n8891), .ZN(n8896) );
  INV_X1 U10216 ( .A(n8966), .ZN(n8895) );
  AND2_X1 U10217 ( .A1(n8894), .A2(n8893), .ZN(n8969) );
  NAND3_X1 U10218 ( .A1(n9283), .A2(n8925), .A3(n8942), .ZN(n8902) );
  NOR2_X1 U10219 ( .A1(n9055), .A2(n8902), .ZN(n8903) );
  NAND2_X1 U10220 ( .A1(n8942), .A2(n8905), .ZN(n8906) );
  MUX2_X1 U10221 ( .A(n9012), .B(n9005), .S(n8925), .Z(n8916) );
  NAND3_X1 U10222 ( .A1(n8917), .A2(n4386), .A3(n8916), .ZN(n8920) );
  MUX2_X1 U10223 ( .A(n9184), .B(n8941), .S(n8925), .Z(n8918) );
  INV_X1 U10224 ( .A(n8923), .ZN(n9041) );
  OAI21_X1 U10225 ( .B1(n8929), .B2(n9002), .A(n9041), .ZN(n8924) );
  NAND2_X1 U10226 ( .A1(n8926), .A2(n9002), .ZN(n8933) );
  AOI21_X1 U10227 ( .B1(n9011), .B2(n8928), .A(n8927), .ZN(n8932) );
  INV_X1 U10228 ( .A(n8929), .ZN(n8930) );
  NAND3_X1 U10229 ( .A1(n8933), .A2(n8932), .A3(n8931), .ZN(n8934) );
  NAND2_X1 U10230 ( .A1(n8935), .A2(n8934), .ZN(n8940) );
  INV_X1 U10231 ( .A(n9090), .ZN(n9042) );
  AND2_X1 U10232 ( .A1(n9046), .A2(n8941), .ZN(n9037) );
  INV_X1 U10233 ( .A(n8942), .ZN(n8945) );
  NOR2_X1 U10234 ( .A1(n8943), .A2(n4710), .ZN(n8944) );
  OR3_X1 U10235 ( .A1(n9055), .A2(n8945), .A3(n8944), .ZN(n8947) );
  NAND2_X1 U10236 ( .A1(n8984), .A2(n9057), .ZN(n8946) );
  OAI21_X1 U10237 ( .B1(n8948), .B2(n8947), .A(n8946), .ZN(n8949) );
  AND2_X1 U10238 ( .A1(n8950), .A2(n8949), .ZN(n9013) );
  AND3_X1 U10239 ( .A1(n8953), .A2(n8952), .A3(n8951), .ZN(n8978) );
  INV_X1 U10240 ( .A(n8978), .ZN(n8980) );
  NAND3_X1 U10241 ( .A1(n8966), .A2(n8955), .A3(n8954), .ZN(n8971) );
  INV_X1 U10242 ( .A(n8956), .ZN(n9023) );
  INV_X1 U10243 ( .A(n9016), .ZN(n8957) );
  AND2_X1 U10244 ( .A1(n9019), .A2(n8957), .ZN(n8958) );
  OR2_X1 U10245 ( .A1(n9023), .A2(n8958), .ZN(n8993) );
  INV_X1 U10246 ( .A(n8959), .ZN(n8960) );
  OAI21_X1 U10247 ( .B1(n8993), .B2(n8961), .A(n8960), .ZN(n8962) );
  OR3_X1 U10248 ( .A1(n8971), .A2(n8972), .A3(n8962), .ZN(n8979) );
  INV_X1 U10249 ( .A(n8963), .ZN(n8976) );
  INV_X1 U10250 ( .A(n8964), .ZN(n8970) );
  NAND3_X1 U10251 ( .A1(n4717), .A2(n8967), .A3(n8966), .ZN(n8968) );
  OAI211_X1 U10252 ( .C1(n8971), .C2(n8970), .A(n8969), .B(n8968), .ZN(n8974)
         );
  INV_X1 U10253 ( .A(n8972), .ZN(n8973) );
  NAND2_X1 U10254 ( .A1(n8974), .A2(n8973), .ZN(n8975) );
  NAND2_X1 U10255 ( .A1(n8976), .A2(n8975), .ZN(n8977) );
  NAND2_X1 U10256 ( .A1(n8978), .A2(n8977), .ZN(n9025) );
  OAI21_X1 U10257 ( .B1(n8980), .B2(n8979), .A(n9025), .ZN(n8982) );
  NAND2_X1 U10258 ( .A1(n8982), .A2(n8981), .ZN(n8983) );
  NOR2_X1 U10259 ( .A1(n8984), .A2(n8983), .ZN(n9026) );
  NAND2_X1 U10260 ( .A1(n6890), .A2(n9724), .ZN(n8985) );
  NAND4_X1 U10261 ( .A1(n8987), .A2(n8986), .A3(n9043), .A4(n8985), .ZN(n8990)
         );
  NAND2_X1 U10262 ( .A1(n9015), .A2(n8988), .ZN(n8989) );
  AOI21_X1 U10263 ( .B1(n9014), .B2(n8990), .A(n8989), .ZN(n8995) );
  AND2_X1 U10264 ( .A1(n9018), .A2(n8991), .ZN(n8992) );
  NAND2_X1 U10265 ( .A1(n9019), .A2(n8992), .ZN(n9021) );
  INV_X1 U10266 ( .A(n8993), .ZN(n8994) );
  OAI211_X1 U10267 ( .C1(n8995), .C2(n9021), .A(n9025), .B(n8994), .ZN(n8996)
         );
  NAND2_X1 U10268 ( .A1(n9026), .A2(n8996), .ZN(n8998) );
  AOI21_X1 U10269 ( .B1(n9013), .B2(n8998), .A(n8997), .ZN(n9000) );
  OAI21_X1 U10270 ( .B1(n9000), .B2(n4703), .A(n8999), .ZN(n9001) );
  NAND4_X1 U10271 ( .A1(n9037), .A2(n9204), .A3(n9047), .A4(n9001), .ZN(n9008)
         );
  NAND2_X1 U10272 ( .A1(n9179), .A2(n9187), .ZN(n9087) );
  NAND2_X1 U10273 ( .A1(n9198), .A2(n9002), .ZN(n9045) );
  INV_X1 U10274 ( .A(n9037), .ZN(n9006) );
  NAND2_X1 U10275 ( .A1(n9012), .A2(n9003), .ZN(n9004) );
  AND3_X1 U10276 ( .A1(n9184), .A2(n9005), .A3(n9004), .ZN(n9033) );
  OR2_X1 U10277 ( .A1(n9006), .A2(n9033), .ZN(n9007) );
  AND4_X1 U10278 ( .A1(n9008), .A2(n9087), .A3(n9045), .A4(n9007), .ZN(n9009)
         );
  OAI21_X1 U10279 ( .B1(n9089), .B2(n9009), .A(n9042), .ZN(n9010) );
  XNOR2_X1 U10280 ( .A(n9010), .B(n9169), .ZN(n9098) );
  INV_X1 U10281 ( .A(n9011), .ZN(n9039) );
  INV_X1 U10282 ( .A(n9012), .ZN(n9035) );
  INV_X1 U10283 ( .A(n9013), .ZN(n9030) );
  NAND2_X1 U10284 ( .A1(n9016), .A2(n9015), .ZN(n9017) );
  NAND3_X1 U10285 ( .A1(n9019), .A2(n9018), .A3(n9017), .ZN(n9020) );
  OAI21_X1 U10286 ( .B1(n9021), .B2(n4413), .A(n9020), .ZN(n9022) );
  NOR2_X1 U10287 ( .A1(n9023), .A2(n9022), .ZN(n9024) );
  AND2_X1 U10288 ( .A1(n9025), .A2(n9024), .ZN(n9028) );
  INV_X1 U10289 ( .A(n9026), .ZN(n9027) );
  OAI21_X1 U10290 ( .B1(n9028), .B2(n9027), .A(n9050), .ZN(n9029) );
  NOR2_X1 U10291 ( .A1(n9030), .A2(n9029), .ZN(n9032) );
  OAI211_X1 U10292 ( .C1(n9032), .C2(n4409), .A(n9047), .B(n9031), .ZN(n9034)
         );
  OAI21_X1 U10293 ( .B1(n9035), .B2(n9034), .A(n9033), .ZN(n9036) );
  NAND2_X1 U10294 ( .A1(n9037), .A2(n9036), .ZN(n9038) );
  NAND3_X1 U10295 ( .A1(n9039), .A2(n9038), .A3(n9045), .ZN(n9040) );
  NAND2_X1 U10296 ( .A1(n9041), .A2(n9040), .ZN(n9044) );
  NAND3_X1 U10297 ( .A1(n9044), .A2(n9043), .A3(n9042), .ZN(n9093) );
  INV_X1 U10298 ( .A(n9447), .ZN(n9443) );
  NAND2_X1 U10299 ( .A1(n9048), .A2(n9047), .ZN(n9227) );
  INV_X1 U10300 ( .A(n9227), .ZN(n9084) );
  INV_X1 U10301 ( .A(n9051), .ZN(n9254) );
  NOR2_X1 U10302 ( .A1(n9052), .A2(n9254), .ZN(n9267) );
  INV_X1 U10303 ( .A(n9053), .ZN(n9054) );
  NAND2_X1 U10304 ( .A1(n9057), .A2(n9056), .ZN(n9285) );
  NOR3_X1 U10305 ( .A1(n9059), .A2(n6896), .A3(n9058), .ZN(n9062) );
  INV_X1 U10306 ( .A(n9675), .ZN(n9664) );
  INV_X1 U10307 ( .A(n9060), .ZN(n9061) );
  NAND4_X1 U10308 ( .A1(n9063), .A2(n9062), .A3(n9664), .A4(n9061), .ZN(n9064)
         );
  NOR2_X1 U10309 ( .A1(n9064), .A2(n7385), .ZN(n9065) );
  AND2_X1 U10310 ( .A1(n9066), .A2(n9065), .ZN(n9067) );
  NAND4_X1 U10311 ( .A1(n9070), .A2(n9069), .A3(n9068), .A4(n9067), .ZN(n9072)
         );
  NOR3_X1 U10312 ( .A1(n9073), .A2(n9072), .A3(n9071), .ZN(n9075) );
  INV_X1 U10313 ( .A(n9413), .ZN(n9074) );
  NAND3_X1 U10314 ( .A1(n9076), .A2(n9075), .A3(n9074), .ZN(n9078) );
  NOR2_X1 U10315 ( .A1(n9079), .A2(n9395), .ZN(n9080) );
  NAND3_X1 U10316 ( .A1(n9256), .A2(n9267), .A3(n9081), .ZN(n9082) );
  NOR2_X1 U10317 ( .A1(n9239), .A2(n9082), .ZN(n9083) );
  NAND3_X1 U10318 ( .A1(n9087), .A2(n9443), .A3(n9086), .ZN(n9088) );
  NAND2_X1 U10319 ( .A1(n9092), .A2(n9091), .ZN(n9094) );
  NAND4_X1 U10320 ( .A1(n9093), .A2(n6504), .A3(n9694), .A4(n9094), .ZN(n9097)
         );
  INV_X1 U10321 ( .A(n9094), .ZN(n9095) );
  NAND2_X1 U10322 ( .A1(n9095), .A2(n4912), .ZN(n9096) );
  OAI211_X1 U10323 ( .C1(n9098), .C2(n6504), .A(n9097), .B(n9096), .ZN(n9099)
         );
  NOR4_X1 U10324 ( .A1(n9101), .A2(n9574), .A3(n9172), .A4(n9722), .ZN(n9103)
         );
  OAI21_X1 U10325 ( .B1(n6899), .B2(n9104), .A(P1_B_REG_SCAN_IN), .ZN(n9102)
         );
  MUX2_X1 U10326 ( .A(n9105), .B(P1_DATAO_REG_29__SCAN_IN), .S(n9117), .Z(
        P1_U3584) );
  MUX2_X1 U10327 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n9214), .S(P1_U4006), .Z(
        P1_U3583) );
  MUX2_X1 U10328 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n9228), .S(P1_U4006), .Z(
        P1_U3582) );
  MUX2_X1 U10329 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n9241), .S(P1_U4006), .Z(
        P1_U3581) );
  MUX2_X1 U10330 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n7887), .S(P1_U4006), .Z(
        P1_U3580) );
  MUX2_X1 U10331 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n9268), .S(P1_U4006), .Z(
        P1_U3579) );
  MUX2_X1 U10332 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n9287), .S(P1_U4006), .Z(
        P1_U3578) );
  MUX2_X1 U10333 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n9293), .S(P1_U4006), .Z(
        P1_U3577) );
  MUX2_X1 U10334 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n9310), .S(P1_U4006), .Z(
        P1_U3576) );
  MUX2_X1 U10335 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n9324), .S(P1_U4006), .Z(
        P1_U3575) );
  MUX2_X1 U10336 ( .A(n9346), .B(P1_DATAO_REG_19__SCAN_IN), .S(n9117), .Z(
        P1_U3574) );
  MUX2_X1 U10337 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n9363), .S(P1_U4006), .Z(
        P1_U3573) );
  MUX2_X1 U10338 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n9386), .S(P1_U4006), .Z(
        P1_U3572) );
  MUX2_X1 U10339 ( .A(n9399), .B(P1_DATAO_REG_16__SCAN_IN), .S(n9117), .Z(
        P1_U3571) );
  MUX2_X1 U10340 ( .A(n9387), .B(P1_DATAO_REG_15__SCAN_IN), .S(n9117), .Z(
        P1_U3570) );
  MUX2_X1 U10341 ( .A(n9397), .B(P1_DATAO_REG_14__SCAN_IN), .S(n9117), .Z(
        P1_U3569) );
  MUX2_X1 U10342 ( .A(n9106), .B(P1_DATAO_REG_13__SCAN_IN), .S(n9117), .Z(
        P1_U3568) );
  MUX2_X1 U10343 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n9107), .S(P1_U4006), .Z(
        P1_U3567) );
  MUX2_X1 U10344 ( .A(n9108), .B(P1_DATAO_REG_11__SCAN_IN), .S(n9117), .Z(
        P1_U3566) );
  MUX2_X1 U10345 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n9109), .S(P1_U4006), .Z(
        P1_U3565) );
  MUX2_X1 U10346 ( .A(n9110), .B(P1_DATAO_REG_9__SCAN_IN), .S(n9117), .Z(
        P1_U3564) );
  MUX2_X1 U10347 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n9111), .S(P1_U4006), .Z(
        P1_U3563) );
  MUX2_X1 U10348 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n9112), .S(P1_U4006), .Z(
        P1_U3562) );
  MUX2_X1 U10349 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n9113), .S(P1_U4006), .Z(
        P1_U3561) );
  MUX2_X1 U10350 ( .A(n9114), .B(P1_DATAO_REG_5__SCAN_IN), .S(n9117), .Z(
        P1_U3560) );
  MUX2_X1 U10351 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n9115), .S(P1_U4006), .Z(
        P1_U3559) );
  MUX2_X1 U10352 ( .A(n9116), .B(P1_DATAO_REG_3__SCAN_IN), .S(n9117), .Z(
        P1_U3558) );
  MUX2_X1 U10353 ( .A(n6893), .B(P1_DATAO_REG_2__SCAN_IN), .S(n9117), .Z(
        P1_U3557) );
  MUX2_X1 U10354 ( .A(n6890), .B(P1_DATAO_REG_1__SCAN_IN), .S(n9117), .Z(
        P1_U3556) );
  OAI211_X1 U10355 ( .C1(n9120), .C2(n9119), .A(n9659), .B(n9118), .ZN(n9121)
         );
  OAI21_X1 U10356 ( .B1(P1_STATE_REG_SCAN_IN), .B2(n9122), .A(n9121), .ZN(
        n9123) );
  AOI21_X1 U10357 ( .B1(n9171), .B2(P1_ADDR_REG_2__SCAN_IN), .A(n9123), .ZN(
        n9130) );
  NAND2_X1 U10358 ( .A1(n9627), .A2(n9124), .ZN(n9129) );
  OAI211_X1 U10359 ( .C1(n9127), .C2(n9126), .A(n9648), .B(n9125), .ZN(n9128)
         );
  NAND4_X1 U10360 ( .A1(n9131), .A2(n9130), .A3(n9129), .A4(n9128), .ZN(
        P1_U3243) );
  XNOR2_X1 U10361 ( .A(n9133), .B(n9132), .ZN(n9135) );
  AOI22_X1 U10362 ( .A1(n9648), .A2(n9135), .B1(n9627), .B2(n9134), .ZN(n9143)
         );
  NAND2_X1 U10363 ( .A1(n9171), .A2(P1_ADDR_REG_5__SCAN_IN), .ZN(n9141) );
  AND2_X1 U10364 ( .A1(n9137), .A2(n9136), .ZN(n9138) );
  OR3_X1 U10365 ( .A1(n9163), .A2(n9139), .A3(n9138), .ZN(n9140) );
  NAND4_X1 U10366 ( .A1(n9143), .A2(n9142), .A3(n9141), .A4(n9140), .ZN(
        P1_U3246) );
  INV_X1 U10367 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n9366) );
  XNOR2_X1 U10368 ( .A(n9158), .B(n9366), .ZN(n9636) );
  NAND2_X1 U10369 ( .A1(n9626), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n9150) );
  OR2_X1 U10370 ( .A1(n9144), .A2(n9155), .ZN(n9146) );
  INV_X1 U10371 ( .A(n9147), .ZN(n9148) );
  NOR2_X1 U10372 ( .A1(n9611), .A2(n9402), .ZN(n9610) );
  OAI21_X1 U10373 ( .B1(n9626), .B2(P1_REG2_REG_16__SCAN_IN), .A(n9150), .ZN(
        n9622) );
  NOR2_X1 U10374 ( .A1(n9623), .A2(n9622), .ZN(n9621) );
  INV_X1 U10375 ( .A(n9621), .ZN(n9149) );
  NAND2_X1 U10376 ( .A1(n9150), .A2(n9149), .ZN(n9635) );
  NAND2_X1 U10377 ( .A1(n9636), .A2(n9635), .ZN(n9634) );
  NAND2_X1 U10378 ( .A1(n9158), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n9151) );
  NAND2_X1 U10379 ( .A1(n9634), .A2(n9151), .ZN(n9649) );
  MUX2_X1 U10380 ( .A(P1_REG2_REG_18__SCAN_IN), .B(n9351), .S(n9152), .Z(n9650) );
  AND2_X1 U10381 ( .A1(n9649), .A2(n9650), .ZN(n9646) );
  AOI21_X1 U10382 ( .B1(n9152), .B2(P1_REG2_REG_18__SCAN_IN), .A(n9646), .ZN(
        n9153) );
  INV_X1 U10383 ( .A(n9158), .ZN(n9639) );
  XNOR2_X1 U10384 ( .A(n9639), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n9642) );
  XOR2_X1 U10385 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n9626), .Z(n9629) );
  OAI21_X1 U10386 ( .B1(P1_REG1_REG_14__SCAN_IN), .B2(n9155), .A(n9154), .ZN(
        n9156) );
  XOR2_X1 U10387 ( .A(n9614), .B(n9156), .Z(n9615) );
  OAI22_X1 U10388 ( .A1(n9615), .A2(n9157), .B1(n4421), .B2(n9156), .ZN(n9630)
         );
  AOI22_X1 U10389 ( .A1(n9642), .A2(n9159), .B1(n9158), .B2(
        P1_REG1_REG_17__SCAN_IN), .ZN(n9657) );
  XNOR2_X1 U10390 ( .A(n9653), .B(P1_REG1_REG_18__SCAN_IN), .ZN(n9656) );
  AND2_X1 U10391 ( .A1(n9657), .A2(n9656), .ZN(n9160) );
  AOI21_X1 U10392 ( .B1(n9653), .B2(n9161), .A(n9160), .ZN(n9162) );
  XOR2_X1 U10393 ( .A(n9162), .B(n10033), .Z(n9165) );
  INV_X1 U10394 ( .A(n9164), .ZN(n9167) );
  AOI21_X1 U10395 ( .B1(n9165), .B2(n9659), .A(n9627), .ZN(n9166) );
  NAND2_X1 U10396 ( .A1(n9192), .A2(n9445), .ZN(n9194) );
  XNOR2_X1 U10397 ( .A(n9178), .B(n9174), .ZN(n9435) );
  INV_X1 U10398 ( .A(P1_B_REG_SCAN_IN), .ZN(n10035) );
  OAI21_X1 U10399 ( .B1(n9172), .B2(n10035), .A(n9398), .ZN(n9188) );
  NOR2_X1 U10400 ( .A1(n9188), .A2(n9173), .ZN(n9432) );
  INV_X1 U10401 ( .A(n9432), .ZN(n9438) );
  NOR2_X1 U10402 ( .A1(n9438), .A2(n9716), .ZN(n9180) );
  NOR2_X1 U10403 ( .A1(n9174), .A2(n9683), .ZN(n9175) );
  AOI211_X1 U10404 ( .C1(n9716), .C2(P1_REG2_REG_31__SCAN_IN), .A(n9180), .B(
        n9175), .ZN(n9176) );
  OAI21_X1 U10405 ( .B1(n9177), .B2(n9435), .A(n9176), .ZN(P1_U3261) );
  INV_X1 U10406 ( .A(n9179), .ZN(n9440) );
  INV_X1 U10407 ( .A(n9178), .ZN(n9437) );
  NAND2_X1 U10408 ( .A1(n9194), .A2(n9179), .ZN(n9436) );
  NAND3_X1 U10409 ( .A1(n9437), .A2(n9670), .A3(n9436), .ZN(n9182) );
  AOI21_X1 U10410 ( .B1(n9716), .B2(P1_REG2_REG_30__SCAN_IN), .A(n9180), .ZN(
        n9181) );
  OAI211_X1 U10411 ( .C1(n9440), .C2(n9683), .A(n9182), .B(n9181), .ZN(
        P1_U3262) );
  NAND2_X1 U10412 ( .A1(n9455), .A2(n9214), .ZN(n9446) );
  NAND2_X1 U10413 ( .A1(n9450), .A2(n9446), .ZN(n9183) );
  XNOR2_X1 U10414 ( .A(n9183), .B(n9447), .ZN(n9203) );
  NAND2_X1 U10415 ( .A1(n9185), .A2(n9184), .ZN(n9186) );
  OAI22_X1 U10416 ( .A1(n9189), .A2(n9703), .B1(n9188), .B2(n9187), .ZN(n9190)
         );
  INV_X1 U10417 ( .A(n9190), .ZN(n9191) );
  INV_X1 U10418 ( .A(n9196), .ZN(n9197) );
  AOI22_X1 U10419 ( .A1(n9716), .A2(P1_REG2_REG_29__SCAN_IN), .B1(n9197), .B2(
        n9277), .ZN(n9200) );
  NAND2_X1 U10420 ( .A1(n9198), .A2(n9426), .ZN(n9199) );
  OAI211_X1 U10421 ( .C1(n9444), .C2(n9354), .A(n9200), .B(n9199), .ZN(n9201)
         );
  AOI21_X1 U10422 ( .B1(n9441), .B2(n9713), .A(n9201), .ZN(n9202) );
  OAI21_X1 U10423 ( .B1(n9203), .B2(n9431), .A(n9202), .ZN(P1_U3355) );
  INV_X1 U10424 ( .A(n9220), .ZN(n9207) );
  AOI211_X1 U10425 ( .C1(n9462), .C2(n9207), .A(n9754), .B(n4611), .ZN(n9461)
         );
  INV_X1 U10426 ( .A(n9208), .ZN(n9209) );
  AOI22_X1 U10427 ( .A1(n9716), .A2(P1_REG2_REG_27__SCAN_IN), .B1(n9209), .B2(
        n9277), .ZN(n9210) );
  OAI21_X1 U10428 ( .B1(n9211), .B2(n9683), .A(n9210), .ZN(n9217) );
  XNOR2_X1 U10429 ( .A(n9213), .B(n9212), .ZN(n9215) );
  AOI222_X1 U10430 ( .A1(n9706), .A2(n9215), .B1(n9214), .B2(n9398), .C1(n9241), .C2(n9396), .ZN(n9464) );
  NOR2_X1 U10431 ( .A1(n9464), .A2(n9716), .ZN(n9216) );
  AOI211_X1 U10432 ( .C1(n9407), .C2(n9461), .A(n9217), .B(n9216), .ZN(n9218)
         );
  OAI21_X1 U10433 ( .B1(n9465), .B2(n9431), .A(n9218), .ZN(P1_U3264) );
  XNOR2_X1 U10434 ( .A(n9219), .B(n9227), .ZN(n9470) );
  INV_X1 U10435 ( .A(n9234), .ZN(n9221) );
  AOI21_X1 U10436 ( .B1(n9466), .B2(n9221), .A(n9220), .ZN(n9467) );
  INV_X1 U10437 ( .A(n9222), .ZN(n9223) );
  AOI22_X1 U10438 ( .A1(n9716), .A2(P1_REG2_REG_26__SCAN_IN), .B1(n9223), .B2(
        n9277), .ZN(n9224) );
  OAI21_X1 U10439 ( .B1(n9225), .B2(n9683), .A(n9224), .ZN(n9231) );
  XOR2_X1 U10440 ( .A(n9227), .B(n9226), .Z(n9229) );
  AOI222_X1 U10441 ( .A1(n9706), .A2(n9229), .B1(n7887), .B2(n9396), .C1(n9228), .C2(n9398), .ZN(n9469) );
  NOR2_X1 U10442 ( .A1(n9469), .A2(n9716), .ZN(n9230) );
  AOI211_X1 U10443 ( .C1(n9670), .C2(n9467), .A(n9231), .B(n9230), .ZN(n9232)
         );
  OAI21_X1 U10444 ( .B1(n9470), .B2(n9431), .A(n9232), .ZN(P1_U3265) );
  XOR2_X1 U10445 ( .A(n9239), .B(n9233), .Z(n9475) );
  AOI211_X1 U10446 ( .C1(n9472), .C2(n9248), .A(n9754), .B(n9234), .ZN(n9471)
         );
  INV_X1 U10447 ( .A(n9235), .ZN(n9236) );
  AOI22_X1 U10448 ( .A1(n9716), .A2(P1_REG2_REG_25__SCAN_IN), .B1(n9236), .B2(
        n9277), .ZN(n9237) );
  OAI21_X1 U10449 ( .B1(n9238), .B2(n9683), .A(n9237), .ZN(n9244) );
  XNOR2_X1 U10450 ( .A(n9240), .B(n9239), .ZN(n9242) );
  AOI222_X1 U10451 ( .A1(n9706), .A2(n9242), .B1(n9241), .B2(n9398), .C1(n9268), .C2(n9396), .ZN(n9474) );
  NOR2_X1 U10452 ( .A1(n9474), .A2(n9716), .ZN(n9243) );
  AOI211_X1 U10453 ( .C1(n9471), .C2(n9407), .A(n9244), .B(n9243), .ZN(n9245)
         );
  OAI21_X1 U10454 ( .B1(n9475), .B2(n9431), .A(n9245), .ZN(P1_U3266) );
  XNOR2_X1 U10455 ( .A(n9246), .B(n9256), .ZN(n9480) );
  INV_X1 U10456 ( .A(n9248), .ZN(n9249) );
  AOI211_X1 U10457 ( .C1(n9477), .C2(n9247), .A(n9754), .B(n9249), .ZN(n9476)
         );
  INV_X1 U10458 ( .A(n9250), .ZN(n9251) );
  AOI22_X1 U10459 ( .A1(n9716), .A2(P1_REG2_REG_24__SCAN_IN), .B1(n9251), .B2(
        n9277), .ZN(n9252) );
  OAI21_X1 U10460 ( .B1(n9253), .B2(n9683), .A(n9252), .ZN(n9258) );
  XOR2_X1 U10461 ( .A(n9256), .B(n9255), .Z(n9257) );
  XNOR2_X1 U10462 ( .A(n9259), .B(n9267), .ZN(n9485) );
  INV_X1 U10463 ( .A(n9274), .ZN(n9261) );
  INV_X1 U10464 ( .A(n9247), .ZN(n9260) );
  AOI211_X1 U10465 ( .C1(n9482), .C2(n9261), .A(n9754), .B(n9260), .ZN(n9481)
         );
  INV_X1 U10466 ( .A(n9262), .ZN(n9263) );
  AOI22_X1 U10467 ( .A1(n9716), .A2(P1_REG2_REG_23__SCAN_IN), .B1(n9263), .B2(
        n9277), .ZN(n9264) );
  OAI21_X1 U10468 ( .B1(n9265), .B2(n9683), .A(n9264), .ZN(n9271) );
  XOR2_X1 U10469 ( .A(n9267), .B(n9266), .Z(n9269) );
  AOI222_X1 U10470 ( .A1(n9706), .A2(n9269), .B1(n9268), .B2(n9398), .C1(n9293), .C2(n9396), .ZN(n9484) );
  NOR2_X1 U10471 ( .A1(n9484), .A2(n9716), .ZN(n9270) );
  AOI211_X1 U10472 ( .C1(n9481), .C2(n9407), .A(n9271), .B(n9270), .ZN(n9272)
         );
  OAI21_X1 U10473 ( .B1(n9431), .B2(n9485), .A(n9272), .ZN(P1_U3268) );
  XNOR2_X1 U10474 ( .A(n9273), .B(n9285), .ZN(n9490) );
  INV_X1 U10475 ( .A(n9302), .ZN(n9275) );
  AOI211_X1 U10476 ( .C1(n9487), .C2(n9275), .A(n9754), .B(n9274), .ZN(n9486)
         );
  INV_X1 U10477 ( .A(n9276), .ZN(n9278) );
  AOI22_X1 U10478 ( .A1(n9716), .A2(P1_REG2_REG_22__SCAN_IN), .B1(n9278), .B2(
        n9277), .ZN(n9279) );
  OAI21_X1 U10479 ( .B1(n9280), .B2(n9683), .A(n9279), .ZN(n9290) );
  INV_X1 U10480 ( .A(n9282), .ZN(n9284) );
  OAI21_X1 U10481 ( .B1(n9281), .B2(n9284), .A(n9283), .ZN(n9286) );
  XNOR2_X1 U10482 ( .A(n9286), .B(n9285), .ZN(n9288) );
  AOI222_X1 U10483 ( .A1(n9706), .A2(n9288), .B1(n9287), .B2(n9398), .C1(n9310), .C2(n9396), .ZN(n9489) );
  NOR2_X1 U10484 ( .A1(n9489), .A2(n9716), .ZN(n9289) );
  AOI211_X1 U10485 ( .C1(n9486), .C2(n9407), .A(n9290), .B(n9289), .ZN(n9291)
         );
  OAI21_X1 U10486 ( .B1(n9431), .B2(n9490), .A(n9291), .ZN(P1_U3269) );
  INV_X1 U10487 ( .A(n9292), .ZN(n9295) );
  XNOR2_X1 U10488 ( .A(n9281), .B(n9298), .ZN(n9294) );
  AOI222_X1 U10489 ( .A1(n9706), .A2(n9294), .B1(n9293), .B2(n9398), .C1(n9324), .C2(n9396), .ZN(n9496) );
  OAI21_X1 U10490 ( .B1(n9295), .B2(n9697), .A(n9496), .ZN(n9296) );
  NAND2_X1 U10491 ( .A1(n9296), .A2(n9713), .ZN(n9306) );
  AOI22_X1 U10492 ( .A1(n9492), .A2(n9426), .B1(P1_REG2_REG_21__SCAN_IN), .B2(
        n9716), .ZN(n9305) );
  NAND2_X1 U10493 ( .A1(n9299), .A2(n9298), .ZN(n9493) );
  NAND3_X1 U10494 ( .A1(n9297), .A2(n9493), .A3(n9391), .ZN(n9304) );
  NAND2_X1 U10495 ( .A1(n9315), .A2(n9492), .ZN(n9300) );
  NAND2_X1 U10496 ( .A1(n9300), .A2(n9737), .ZN(n9301) );
  NOR2_X1 U10497 ( .A1(n9302), .A2(n9301), .ZN(n9491) );
  NAND2_X1 U10498 ( .A1(n9491), .A2(n9407), .ZN(n9303) );
  NAND4_X1 U10499 ( .A1(n9306), .A2(n9305), .A3(n9304), .A4(n9303), .ZN(
        P1_U3270) );
  XNOR2_X1 U10500 ( .A(n9307), .B(n9308), .ZN(n9501) );
  XNOR2_X1 U10501 ( .A(n9309), .B(n9308), .ZN(n9311) );
  AOI222_X1 U10502 ( .A1(n9706), .A2(n9311), .B1(n9310), .B2(n9398), .C1(n9346), .C2(n9396), .ZN(n9500) );
  INV_X1 U10503 ( .A(P1_REG2_REG_20__SCAN_IN), .ZN(n9312) );
  OAI22_X1 U10504 ( .A1(n9313), .A2(n9697), .B1(n9312), .B2(n9713), .ZN(n9314)
         );
  AOI21_X1 U10505 ( .B1(n9498), .B2(n9426), .A(n9314), .ZN(n9318) );
  AOI21_X1 U10506 ( .B1(n9331), .B2(n9498), .A(n9754), .ZN(n9316) );
  AND2_X1 U10507 ( .A1(n9316), .A2(n9315), .ZN(n9497) );
  NAND2_X1 U10508 ( .A1(n9497), .A2(n9407), .ZN(n9317) );
  OAI211_X1 U10509 ( .C1(n9500), .C2(n9716), .A(n9318), .B(n9317), .ZN(n9319)
         );
  INV_X1 U10510 ( .A(n9319), .ZN(n9320) );
  OAI21_X1 U10511 ( .B1(n9431), .B2(n9501), .A(n9320), .ZN(P1_U3271) );
  XOR2_X1 U10512 ( .A(n9321), .B(n9322), .Z(n9506) );
  XNOR2_X1 U10513 ( .A(n9323), .B(n9322), .ZN(n9325) );
  AOI222_X1 U10514 ( .A1(n9706), .A2(n9325), .B1(n9324), .B2(n9398), .C1(n9363), .C2(n9396), .ZN(n9505) );
  INV_X1 U10515 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n9327) );
  OAI22_X1 U10516 ( .A1(n9713), .A2(n9327), .B1(n9326), .B2(n9697), .ZN(n9328)
         );
  AOI21_X1 U10517 ( .B1(n9503), .B2(n9426), .A(n9328), .ZN(n9333) );
  OR2_X1 U10518 ( .A1(n9353), .A2(n9329), .ZN(n9330) );
  AND3_X1 U10519 ( .A1(n9331), .A2(n9330), .A3(n9737), .ZN(n9502) );
  NAND2_X1 U10520 ( .A1(n9502), .A2(n9407), .ZN(n9332) );
  OAI211_X1 U10521 ( .C1(n9505), .C2(n9716), .A(n9333), .B(n9332), .ZN(n9334)
         );
  INV_X1 U10522 ( .A(n9334), .ZN(n9335) );
  OAI21_X1 U10523 ( .B1(n9431), .B2(n9506), .A(n9335), .ZN(P1_U3272) );
  NAND2_X1 U10524 ( .A1(n9337), .A2(n9342), .ZN(n9338) );
  NAND2_X1 U10525 ( .A1(n9336), .A2(n9338), .ZN(n9507) );
  INV_X1 U10526 ( .A(n9339), .ZN(n9340) );
  OR2_X1 U10527 ( .A1(n9341), .A2(n9340), .ZN(n9344) );
  INV_X1 U10528 ( .A(n9342), .ZN(n9343) );
  XNOR2_X1 U10529 ( .A(n9344), .B(n9343), .ZN(n9345) );
  NAND2_X1 U10530 ( .A1(n9345), .A2(n9706), .ZN(n9348) );
  AOI22_X1 U10531 ( .A1(n9346), .A2(n9398), .B1(n9396), .B2(n9386), .ZN(n9347)
         );
  NAND2_X1 U10532 ( .A1(n9348), .A2(n9347), .ZN(n9512) );
  NAND2_X1 U10533 ( .A1(n9512), .A2(n9713), .ZN(n9359) );
  INV_X1 U10534 ( .A(n9349), .ZN(n9350) );
  OAI22_X1 U10535 ( .A1(n9713), .A2(n9351), .B1(n9350), .B2(n9697), .ZN(n9356)
         );
  OAI21_X1 U10536 ( .B1(n9369), .B2(n9509), .A(n9737), .ZN(n9352) );
  OR2_X1 U10537 ( .A1(n9353), .A2(n9352), .ZN(n9508) );
  NOR2_X1 U10538 ( .A1(n9508), .A2(n9354), .ZN(n9355) );
  AOI211_X1 U10539 ( .C1(n9426), .C2(n9357), .A(n9356), .B(n9355), .ZN(n9358)
         );
  OAI211_X1 U10540 ( .C1(n9507), .C2(n9431), .A(n9359), .B(n9358), .ZN(
        P1_U3273) );
  XNOR2_X1 U10541 ( .A(n9360), .B(n9361), .ZN(n9517) );
  XNOR2_X1 U10542 ( .A(n9362), .B(n9361), .ZN(n9364) );
  AOI222_X1 U10543 ( .A1(n9706), .A2(n9364), .B1(n9363), .B2(n9398), .C1(n9399), .C2(n9396), .ZN(n9516) );
  OAI22_X1 U10544 ( .A1(n9713), .A2(n9366), .B1(n9365), .B2(n9697), .ZN(n9367)
         );
  AOI21_X1 U10545 ( .B1(n9514), .B2(n9426), .A(n9367), .ZN(n9372) );
  OAI21_X1 U10546 ( .B1(n9377), .B2(n9368), .A(n9737), .ZN(n9370) );
  NOR2_X1 U10547 ( .A1(n9370), .A2(n9369), .ZN(n9513) );
  NAND2_X1 U10548 ( .A1(n9513), .A2(n9407), .ZN(n9371) );
  OAI211_X1 U10549 ( .C1(n9516), .C2(n9716), .A(n9372), .B(n9371), .ZN(n9373)
         );
  INV_X1 U10550 ( .A(n9373), .ZN(n9374) );
  OAI21_X1 U10551 ( .B1(n9431), .B2(n9517), .A(n9374), .ZN(P1_U3274) );
  XNOR2_X1 U10552 ( .A(n9375), .B(n9384), .ZN(n9518) );
  NAND2_X1 U10553 ( .A1(n9406), .A2(n9382), .ZN(n9376) );
  NAND2_X1 U10554 ( .A1(n9376), .A2(n9737), .ZN(n9378) );
  OR2_X1 U10555 ( .A1(n9378), .A2(n9377), .ZN(n9519) );
  INV_X1 U10556 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n9380) );
  OAI22_X1 U10557 ( .A1(n9713), .A2(n9380), .B1(n9379), .B2(n9697), .ZN(n9381)
         );
  AOI21_X1 U10558 ( .B1(n9382), .B2(n9426), .A(n9381), .ZN(n9383) );
  OAI21_X1 U10559 ( .B1(n9519), .B2(n9422), .A(n9383), .ZN(n9390) );
  XNOR2_X1 U10560 ( .A(n9385), .B(n9384), .ZN(n9388) );
  AOI222_X1 U10561 ( .A1(n9706), .A2(n9388), .B1(n9387), .B2(n9396), .C1(n9386), .C2(n9398), .ZN(n9522) );
  NOR2_X1 U10562 ( .A1(n9522), .A2(n9716), .ZN(n9389) );
  AOI211_X1 U10563 ( .C1(n9518), .C2(n9391), .A(n9390), .B(n9389), .ZN(n9392)
         );
  INV_X1 U10564 ( .A(n9392), .ZN(P1_U3275) );
  XOR2_X1 U10565 ( .A(n9395), .B(n9393), .Z(n9527) );
  XNOR2_X1 U10566 ( .A(n9394), .B(n9395), .ZN(n9400) );
  AOI222_X1 U10567 ( .A1(n9706), .A2(n9400), .B1(n9399), .B2(n9398), .C1(n9397), .C2(n9396), .ZN(n9526) );
  OAI22_X1 U10568 ( .A1(n9713), .A2(n9402), .B1(n9401), .B2(n9697), .ZN(n9403)
         );
  AOI21_X1 U10569 ( .B1(n9524), .B2(n9426), .A(n9403), .ZN(n9409) );
  INV_X1 U10570 ( .A(n9404), .ZN(n9420) );
  AOI21_X1 U10571 ( .B1(n9420), .B2(n9524), .A(n9754), .ZN(n9405) );
  AND2_X1 U10572 ( .A1(n9406), .A2(n9405), .ZN(n9523) );
  NAND2_X1 U10573 ( .A1(n9523), .A2(n9407), .ZN(n9408) );
  OAI211_X1 U10574 ( .C1(n9526), .C2(n9716), .A(n9409), .B(n9408), .ZN(n9410)
         );
  INV_X1 U10575 ( .A(n9410), .ZN(n9411) );
  OAI21_X1 U10576 ( .B1(n9431), .B2(n9527), .A(n9411), .ZN(P1_U3276) );
  XNOR2_X1 U10577 ( .A(n9412), .B(n9413), .ZN(n9532) );
  XNOR2_X1 U10578 ( .A(n9414), .B(n9413), .ZN(n9415) );
  OAI222_X1 U10579 ( .A1(n9702), .A2(n9418), .B1(n9703), .B2(n9417), .C1(n9416), .C2(n9415), .ZN(n9528) );
  AOI21_X1 U10580 ( .B1(n9419), .B2(n9530), .A(n9754), .ZN(n9421) );
  AND2_X1 U10581 ( .A1(n9421), .A2(n9420), .ZN(n9529) );
  INV_X1 U10582 ( .A(n9422), .ZN(n9423) );
  NAND2_X1 U10583 ( .A1(n9529), .A2(n9423), .ZN(n9428) );
  OAI22_X1 U10584 ( .A1(n9713), .A2(n7273), .B1(n9424), .B2(n9697), .ZN(n9425)
         );
  AOI21_X1 U10585 ( .B1(n9530), .B2(n9426), .A(n9425), .ZN(n9427) );
  NAND2_X1 U10586 ( .A1(n9428), .A2(n9427), .ZN(n9429) );
  AOI21_X1 U10587 ( .B1(n9528), .B2(n9713), .A(n9429), .ZN(n9430) );
  OAI21_X1 U10588 ( .B1(n9532), .B2(n9431), .A(n9430), .ZN(P1_U3277) );
  AOI21_X1 U10589 ( .B1(n9433), .B2(n9736), .A(n9432), .ZN(n9434) );
  OAI21_X1 U10590 ( .B1(n9435), .B2(n9754), .A(n9434), .ZN(n9543) );
  MUX2_X1 U10591 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n9543), .S(n9785), .Z(
        P1_U3554) );
  NAND3_X1 U10592 ( .A1(n9437), .A2(n9737), .A3(n9436), .ZN(n9439) );
  OAI211_X1 U10593 ( .C1(n9440), .C2(n9768), .A(n9439), .B(n9438), .ZN(n9544)
         );
  MUX2_X1 U10594 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n9544), .S(n9785), .Z(
        P1_U3553) );
  AND2_X1 U10595 ( .A1(n9447), .A2(n4903), .ZN(n9442) );
  NAND2_X1 U10596 ( .A1(n9450), .A2(n9442), .ZN(n9453) );
  NAND2_X1 U10597 ( .A1(n9443), .A2(n9759), .ZN(n9449) );
  NOR3_X1 U10598 ( .A1(n9447), .A2(n9745), .A3(n9446), .ZN(n9448) );
  INV_X1 U10599 ( .A(n9451), .ZN(n9452) );
  NAND3_X1 U10600 ( .A1(n9454), .A2(n9453), .A3(n9452), .ZN(n9545) );
  MUX2_X1 U10601 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n9545), .S(n9785), .Z(
        P1_U3552) );
  AOI22_X1 U10602 ( .A1(n9456), .A2(n9737), .B1(n9736), .B2(n9455), .ZN(n9457)
         );
  OAI21_X1 U10603 ( .B1(n9460), .B2(n9745), .A(n9459), .ZN(n9546) );
  MUX2_X1 U10604 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n9546), .S(n9785), .Z(
        P1_U3551) );
  AOI21_X1 U10605 ( .B1(n9736), .B2(n9462), .A(n9461), .ZN(n9463) );
  OAI211_X1 U10606 ( .C1(n9465), .C2(n9745), .A(n9464), .B(n9463), .ZN(n9547)
         );
  MUX2_X1 U10607 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n9547), .S(n9785), .Z(
        P1_U3550) );
  AOI22_X1 U10608 ( .A1(n9467), .A2(n9737), .B1(n9736), .B2(n9466), .ZN(n9468)
         );
  OAI211_X1 U10609 ( .C1(n9470), .C2(n9745), .A(n9469), .B(n9468), .ZN(n9548)
         );
  MUX2_X1 U10610 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n9548), .S(n9785), .Z(
        P1_U3549) );
  AOI21_X1 U10611 ( .B1(n9736), .B2(n9472), .A(n9471), .ZN(n9473) );
  OAI211_X1 U10612 ( .C1(n9475), .C2(n9745), .A(n9474), .B(n9473), .ZN(n9549)
         );
  MUX2_X1 U10613 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n9549), .S(n9785), .Z(
        P1_U3548) );
  AOI21_X1 U10614 ( .B1(n9736), .B2(n9477), .A(n9476), .ZN(n9478) );
  OAI211_X1 U10615 ( .C1(n9745), .C2(n9480), .A(n9479), .B(n9478), .ZN(n9550)
         );
  MUX2_X1 U10616 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n9550), .S(n9785), .Z(
        P1_U3547) );
  AOI21_X1 U10617 ( .B1(n9736), .B2(n9482), .A(n9481), .ZN(n9483) );
  OAI211_X1 U10618 ( .C1(n9745), .C2(n9485), .A(n9484), .B(n9483), .ZN(n9551)
         );
  MUX2_X1 U10619 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n9551), .S(n9785), .Z(
        P1_U3546) );
  AOI21_X1 U10620 ( .B1(n9736), .B2(n9487), .A(n9486), .ZN(n9488) );
  OAI211_X1 U10621 ( .C1(n9745), .C2(n9490), .A(n9489), .B(n9488), .ZN(n9552)
         );
  MUX2_X1 U10622 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n9552), .S(n9785), .Z(
        P1_U3545) );
  AOI21_X1 U10623 ( .B1(n9736), .B2(n9492), .A(n9491), .ZN(n9495) );
  NAND3_X1 U10624 ( .A1(n9297), .A2(n9493), .A3(n9759), .ZN(n9494) );
  NAND3_X1 U10625 ( .A1(n9496), .A2(n9495), .A3(n9494), .ZN(n9553) );
  MUX2_X1 U10626 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n9553), .S(n9785), .Z(
        P1_U3544) );
  AOI21_X1 U10627 ( .B1(n9736), .B2(n9498), .A(n9497), .ZN(n9499) );
  OAI211_X1 U10628 ( .C1(n9745), .C2(n9501), .A(n9500), .B(n9499), .ZN(n9554)
         );
  MUX2_X1 U10629 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n9554), .S(n9785), .Z(
        P1_U3543) );
  AOI21_X1 U10630 ( .B1(n9736), .B2(n9503), .A(n9502), .ZN(n9504) );
  OAI211_X1 U10631 ( .C1(n9745), .C2(n9506), .A(n9505), .B(n9504), .ZN(n9555)
         );
  MUX2_X1 U10632 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n9555), .S(n9785), .Z(
        P1_U3542) );
  NOR2_X1 U10633 ( .A1(n9507), .A2(n9745), .ZN(n9511) );
  OAI21_X1 U10634 ( .B1(n9509), .B2(n9768), .A(n9508), .ZN(n9510) );
  MUX2_X1 U10635 ( .A(n9556), .B(P1_REG1_REG_18__SCAN_IN), .S(n9783), .Z(
        P1_U3541) );
  AOI21_X1 U10636 ( .B1(n9736), .B2(n9514), .A(n9513), .ZN(n9515) );
  OAI211_X1 U10637 ( .C1(n9745), .C2(n9517), .A(n9516), .B(n9515), .ZN(n9557)
         );
  MUX2_X1 U10638 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n9557), .S(n9785), .Z(
        P1_U3540) );
  NAND2_X1 U10639 ( .A1(n9518), .A2(n9759), .ZN(n9521) );
  NAND4_X1 U10640 ( .A1(n9522), .A2(n9521), .A3(n9520), .A4(n9519), .ZN(n9558)
         );
  MUX2_X1 U10641 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n9558), .S(n9785), .Z(
        P1_U3539) );
  AOI21_X1 U10642 ( .B1(n9736), .B2(n9524), .A(n9523), .ZN(n9525) );
  OAI211_X1 U10643 ( .C1(n9745), .C2(n9527), .A(n9526), .B(n9525), .ZN(n9559)
         );
  MUX2_X1 U10644 ( .A(P1_REG1_REG_15__SCAN_IN), .B(n9559), .S(n9785), .Z(
        P1_U3538) );
  AOI211_X1 U10645 ( .C1(n9736), .C2(n9530), .A(n9529), .B(n9528), .ZN(n9531)
         );
  OAI21_X1 U10646 ( .B1(n9745), .B2(n9532), .A(n9531), .ZN(n9560) );
  MUX2_X1 U10647 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n9560), .S(n9785), .Z(
        P1_U3537) );
  AOI22_X1 U10648 ( .A1(n9534), .A2(n9737), .B1(n9736), .B2(n9533), .ZN(n9535)
         );
  OAI211_X1 U10649 ( .C1(n9740), .C2(n9537), .A(n9536), .B(n9535), .ZN(n9561)
         );
  MUX2_X1 U10650 ( .A(P1_REG1_REG_13__SCAN_IN), .B(n9561), .S(n9785), .Z(
        P1_U3536) );
  NAND3_X1 U10651 ( .A1(n9538), .A2(n9759), .A3(n7772), .ZN(n9540) );
  NAND4_X1 U10652 ( .A1(n9542), .A2(n9541), .A3(n9540), .A4(n9539), .ZN(n9562)
         );
  MUX2_X1 U10653 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n9562), .S(n9785), .Z(
        P1_U3535) );
  MUX2_X1 U10654 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n9543), .S(n9776), .Z(
        P1_U3522) );
  MUX2_X1 U10655 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n9544), .S(n9776), .Z(
        P1_U3521) );
  MUX2_X1 U10656 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n9545), .S(n9776), .Z(
        P1_U3520) );
  MUX2_X1 U10657 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n9546), .S(n9776), .Z(
        P1_U3519) );
  MUX2_X1 U10658 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n9547), .S(n9776), .Z(
        P1_U3518) );
  MUX2_X1 U10659 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n9548), .S(n9776), .Z(
        P1_U3517) );
  MUX2_X1 U10660 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n9549), .S(n9776), .Z(
        P1_U3516) );
  MUX2_X1 U10661 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n9550), .S(n9776), .Z(
        P1_U3515) );
  MUX2_X1 U10662 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n9551), .S(n9776), .Z(
        P1_U3514) );
  MUX2_X1 U10663 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n9552), .S(n9776), .Z(
        P1_U3513) );
  MUX2_X1 U10664 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n9553), .S(n9776), .Z(
        P1_U3512) );
  MUX2_X1 U10665 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n9554), .S(n9776), .Z(
        P1_U3511) );
  MUX2_X1 U10666 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n9555), .S(n9776), .Z(
        P1_U3510) );
  MUX2_X1 U10667 ( .A(n9556), .B(P1_REG0_REG_18__SCAN_IN), .S(n9774), .Z(
        P1_U3508) );
  MUX2_X1 U10668 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n9557), .S(n9776), .Z(
        P1_U3505) );
  MUX2_X1 U10669 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n9558), .S(n9776), .Z(
        P1_U3502) );
  MUX2_X1 U10670 ( .A(P1_REG0_REG_15__SCAN_IN), .B(n9559), .S(n9776), .Z(
        P1_U3499) );
  MUX2_X1 U10671 ( .A(P1_REG0_REG_14__SCAN_IN), .B(n9560), .S(n9776), .Z(
        P1_U3496) );
  MUX2_X1 U10672 ( .A(P1_REG0_REG_13__SCAN_IN), .B(n9561), .S(n9776), .Z(
        P1_U3493) );
  MUX2_X1 U10673 ( .A(P1_REG0_REG_12__SCAN_IN), .B(n9562), .S(n9776), .Z(
        P1_U3490) );
  MUX2_X1 U10674 ( .A(n9563), .B(P1_D_REG_0__SCAN_IN), .S(n9722), .Z(P1_U3440)
         );
  NOR4_X1 U10675 ( .A1(n9564), .A2(P1_IR_REG_30__SCAN_IN), .A3(P1_U3084), .A4(
        n6275), .ZN(n9565) );
  AOI21_X1 U10676 ( .B1(n9566), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n9565), .ZN(
        n9567) );
  OAI21_X1 U10677 ( .B1(n9568), .B2(n9572), .A(n9567), .ZN(P1_U3322) );
  INV_X1 U10678 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n9569) );
  OAI222_X1 U10679 ( .A1(n9572), .A2(n9571), .B1(n9570), .B2(P1_U3084), .C1(
        n9569), .C2(n9576), .ZN(P1_U3324) );
  OAI222_X1 U10680 ( .A1(n9576), .A2(n9990), .B1(P1_U3084), .B2(n9574), .C1(
        n9573), .C2(n9572), .ZN(P1_U3325) );
  MUX2_X1 U10681 ( .A(n9577), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3353) );
  NOR2_X1 U10682 ( .A1(P1_ADDR_REG_17__SCAN_IN), .A2(P2_ADDR_REG_17__SCAN_IN), 
        .ZN(n9578) );
  AOI21_X1 U10683 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(P1_ADDR_REG_17__SCAN_IN), 
        .A(n9578), .ZN(n9881) );
  NOR2_X1 U10684 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n9579) );
  AOI21_X1 U10685 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(P2_ADDR_REG_16__SCAN_IN), 
        .A(n9579), .ZN(n9884) );
  NOR2_X1 U10686 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n9580) );
  AOI21_X1 U10687 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(P2_ADDR_REG_15__SCAN_IN), 
        .A(n9580), .ZN(n9887) );
  NOR2_X1 U10688 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n9581) );
  AOI21_X1 U10689 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(P2_ADDR_REG_14__SCAN_IN), 
        .A(n9581), .ZN(n9890) );
  NOR2_X1 U10690 ( .A1(P1_ADDR_REG_13__SCAN_IN), .A2(P2_ADDR_REG_13__SCAN_IN), 
        .ZN(n9582) );
  AOI21_X1 U10691 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(P1_ADDR_REG_13__SCAN_IN), 
        .A(n9582), .ZN(n9893) );
  NOR2_X1 U10692 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n9589) );
  XNOR2_X1 U10693 ( .A(P1_ADDR_REG_4__SCAN_IN), .B(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n10071) );
  NAND2_X1 U10694 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n9587) );
  XOR2_X1 U10695 ( .A(P1_ADDR_REG_3__SCAN_IN), .B(P2_ADDR_REG_3__SCAN_IN), .Z(
        n10069) );
  NAND2_X1 U10696 ( .A1(P2_ADDR_REG_2__SCAN_IN), .A2(P1_ADDR_REG_2__SCAN_IN), 
        .ZN(n9585) );
  XOR2_X1 U10697 ( .A(P2_ADDR_REG_2__SCAN_IN), .B(P1_ADDR_REG_2__SCAN_IN), .Z(
        n10067) );
  AOI21_X1 U10698 ( .B1(P2_ADDR_REG_0__SCAN_IN), .B2(P1_ADDR_REG_0__SCAN_IN), 
        .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n9875) );
  INV_X1 U10699 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n9583) );
  NAND3_X1 U10700 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .A3(P1_ADDR_REG_1__SCAN_IN), .ZN(n9877) );
  NAND2_X1 U10701 ( .A1(n10067), .A2(n10066), .ZN(n9584) );
  NAND2_X1 U10702 ( .A1(n9585), .A2(n9584), .ZN(n10068) );
  NAND2_X1 U10703 ( .A1(n10069), .A2(n10068), .ZN(n9586) );
  NAND2_X1 U10704 ( .A1(n9587), .A2(n9586), .ZN(n10070) );
  NOR2_X1 U10705 ( .A1(n10071), .A2(n10070), .ZN(n9588) );
  NOR2_X1 U10706 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n9590), .ZN(n10055) );
  NAND2_X1 U10707 ( .A1(n9592), .A2(P1_ADDR_REG_6__SCAN_IN), .ZN(n9594) );
  NAND2_X1 U10708 ( .A1(n10053), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n9593) );
  NAND2_X1 U10709 ( .A1(P1_ADDR_REG_7__SCAN_IN), .A2(n9595), .ZN(n9597) );
  NAND2_X1 U10710 ( .A1(n10057), .A2(P2_ADDR_REG_7__SCAN_IN), .ZN(n9596) );
  NAND2_X1 U10711 ( .A1(P1_ADDR_REG_8__SCAN_IN), .A2(n9598), .ZN(n9600) );
  NAND2_X1 U10712 ( .A1(n10062), .A2(P2_ADDR_REG_8__SCAN_IN), .ZN(n9599) );
  NAND2_X1 U10713 ( .A1(n9600), .A2(n9599), .ZN(n9601) );
  AND2_X1 U10714 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(n9601), .ZN(n9602) );
  XNOR2_X1 U10715 ( .A(P2_ADDR_REG_9__SCAN_IN), .B(n9601), .ZN(n10064) );
  NAND2_X1 U10716 ( .A1(P1_ADDR_REG_10__SCAN_IN), .A2(P2_ADDR_REG_10__SCAN_IN), 
        .ZN(n9603) );
  OAI21_X1 U10717 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(P2_ADDR_REG_10__SCAN_IN), 
        .A(n9603), .ZN(n9901) );
  NAND2_X1 U10718 ( .A1(P1_ADDR_REG_11__SCAN_IN), .A2(P2_ADDR_REG_11__SCAN_IN), 
        .ZN(n9604) );
  OAI21_X1 U10719 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(P2_ADDR_REG_11__SCAN_IN), 
        .A(n9604), .ZN(n9898) );
  NOR2_X1 U10720 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n9605) );
  AOI21_X1 U10721 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(P2_ADDR_REG_12__SCAN_IN), 
        .A(n9605), .ZN(n9895) );
  NAND2_X1 U10722 ( .A1(n9890), .A2(n9889), .ZN(n9888) );
  NAND2_X1 U10723 ( .A1(n9884), .A2(n9883), .ZN(n9882) );
  OAI21_X1 U10724 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(P1_ADDR_REG_16__SCAN_IN), 
        .A(n9882), .ZN(n9880) );
  NAND2_X1 U10725 ( .A1(n9881), .A2(n9880), .ZN(n9879) );
  NOR2_X1 U10726 ( .A1(n10060), .A2(n10059), .ZN(n9606) );
  NAND2_X1 U10727 ( .A1(n10060), .A2(n10059), .ZN(n10058) );
  XOR2_X1 U10728 ( .A(P1_ADDR_REG_19__SCAN_IN), .B(P2_ADDR_REG_19__SCAN_IN), 
        .Z(n9607) );
  XNOR2_X1 U10729 ( .A(n9608), .B(n9607), .ZN(ADD_1071_U4) );
  XNOR2_X1 U10730 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  XNOR2_X1 U10731 ( .A(P1_RD_REG_SCAN_IN), .B(P2_RD_REG_SCAN_IN), .ZN(U126) );
  INV_X1 U10732 ( .A(n9609), .ZN(n9613) );
  AOI211_X1 U10733 ( .C1(n9402), .C2(n9611), .A(n9620), .B(n9610), .ZN(n9612)
         );
  AOI211_X1 U10734 ( .C1(n9627), .C2(n9614), .A(n9613), .B(n9612), .ZN(n9618)
         );
  XNOR2_X1 U10735 ( .A(n9615), .B(P1_REG1_REG_15__SCAN_IN), .ZN(n9616) );
  NAND2_X1 U10736 ( .A1(n9616), .A2(n9659), .ZN(n9617) );
  OAI211_X1 U10737 ( .C1(n4371), .C2(n9662), .A(n9618), .B(n9617), .ZN(
        P1_U3256) );
  INV_X1 U10738 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n9633) );
  INV_X1 U10739 ( .A(n9619), .ZN(n9625) );
  AOI211_X1 U10740 ( .C1(n9623), .C2(n9622), .A(n9621), .B(n9620), .ZN(n9624)
         );
  AOI211_X1 U10741 ( .C1(n9627), .C2(n9626), .A(n9625), .B(n9624), .ZN(n9632)
         );
  OAI211_X1 U10742 ( .C1(n9630), .C2(n9629), .A(n9659), .B(n9628), .ZN(n9631)
         );
  OAI211_X1 U10743 ( .C1(n9633), .C2(n9662), .A(n9632), .B(n9631), .ZN(
        P1_U3257) );
  INV_X1 U10744 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n10030) );
  OAI211_X1 U10745 ( .C1(n9636), .C2(n9635), .A(n9648), .B(n9634), .ZN(n9637)
         );
  OAI211_X1 U10746 ( .C1(n9654), .C2(n9639), .A(n9638), .B(n9637), .ZN(n9640)
         );
  INV_X1 U10747 ( .A(n9640), .ZN(n9645) );
  XNOR2_X1 U10748 ( .A(n9642), .B(n9641), .ZN(n9643) );
  NAND2_X1 U10749 ( .A1(n9659), .A2(n9643), .ZN(n9644) );
  OAI211_X1 U10750 ( .C1(n10030), .C2(n9662), .A(n9645), .B(n9644), .ZN(
        P1_U3258) );
  INV_X1 U10751 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n9663) );
  INV_X1 U10752 ( .A(n9646), .ZN(n9647) );
  OAI211_X1 U10753 ( .C1(n9650), .C2(n9649), .A(n9648), .B(n9647), .ZN(n9651)
         );
  OAI211_X1 U10754 ( .C1(n9654), .C2(n9653), .A(n9652), .B(n9651), .ZN(n9655)
         );
  INV_X1 U10755 ( .A(n9655), .ZN(n9661) );
  XNOR2_X1 U10756 ( .A(n9657), .B(n9656), .ZN(n9658) );
  NAND2_X1 U10757 ( .A1(n9659), .A2(n9658), .ZN(n9660) );
  OAI211_X1 U10758 ( .C1(n9663), .C2(n9662), .A(n9661), .B(n9660), .ZN(
        P1_U3259) );
  XNOR2_X1 U10759 ( .A(n9665), .B(n9664), .ZN(n9741) );
  OR2_X1 U10760 ( .A1(n9741), .A2(n9666), .ZN(n9672) );
  OR2_X1 U10761 ( .A1(n9667), .A2(n9682), .ZN(n9669) );
  AND2_X1 U10762 ( .A1(n9669), .A2(n9668), .ZN(n9738) );
  NAND2_X1 U10763 ( .A1(n9670), .A2(n9738), .ZN(n9671) );
  AND2_X1 U10764 ( .A1(n9672), .A2(n9671), .ZN(n9687) );
  NOR2_X1 U10765 ( .A1(n9673), .A2(n4413), .ZN(n9674) );
  XNOR2_X1 U10766 ( .A(n9675), .B(n9674), .ZN(n9679) );
  OAI22_X1 U10767 ( .A1(n9677), .A2(n9703), .B1(n9702), .B2(n9676), .ZN(n9678)
         );
  AOI21_X1 U10768 ( .B1(n9679), .B2(n9706), .A(n9678), .ZN(n9680) );
  OAI21_X1 U10769 ( .B1(n9741), .B2(n9710), .A(n9680), .ZN(n9743) );
  MUX2_X1 U10770 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n9743), .S(n9713), .Z(n9685)
         );
  OAI22_X1 U10771 ( .A1(n9683), .A2(n9682), .B1(n9681), .B2(n9697), .ZN(n9684)
         );
  NOR2_X1 U10772 ( .A1(n9685), .A2(n9684), .ZN(n9686) );
  NAND2_X1 U10773 ( .A1(n9687), .A2(n9686), .ZN(P1_U3287) );
  INV_X1 U10774 ( .A(n6896), .ZN(n9700) );
  XNOR2_X1 U10775 ( .A(n9700), .B(n9688), .ZN(n9709) );
  INV_X1 U10776 ( .A(n9709), .ZN(n9727) );
  OAI21_X1 U10777 ( .B1(n9724), .B2(n9690), .A(n9689), .ZN(n9691) );
  OR2_X1 U10778 ( .A1(n9754), .A2(n9691), .ZN(n9723) );
  INV_X1 U10779 ( .A(n9723), .ZN(n9695) );
  AOI22_X1 U10780 ( .A1(n9695), .A2(n9694), .B1(n9693), .B2(n9692), .ZN(n9696)
         );
  OAI21_X1 U10781 ( .B1(n9698), .B2(n9697), .A(n9696), .ZN(n9711) );
  XNOR2_X1 U10782 ( .A(n9700), .B(n9699), .ZN(n9707) );
  OAI22_X1 U10783 ( .A1(n9704), .A2(n9703), .B1(n9702), .B2(n9701), .ZN(n9705)
         );
  AOI21_X1 U10784 ( .B1(n9707), .B2(n9706), .A(n9705), .ZN(n9708) );
  OAI21_X1 U10785 ( .B1(n9710), .B2(n9709), .A(n9708), .ZN(n9725) );
  AOI211_X1 U10786 ( .C1(n9712), .C2(n9727), .A(n9711), .B(n9725), .ZN(n9714)
         );
  AOI22_X1 U10787 ( .A1(n9716), .A2(n9715), .B1(n9714), .B2(n9713), .ZN(
        P1_U3290) );
  INV_X1 U10788 ( .A(n9717), .ZN(n9718) );
  AND2_X1 U10789 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n9720), .ZN(P1_U3292) );
  AND2_X1 U10790 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n9720), .ZN(P1_U3293) );
  AND2_X1 U10791 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n9720), .ZN(P1_U3294) );
  AND2_X1 U10792 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n9720), .ZN(P1_U3295) );
  AND2_X1 U10793 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n9720), .ZN(P1_U3296) );
  INV_X1 U10794 ( .A(n9720), .ZN(n9719) );
  INV_X1 U10795 ( .A(P1_D_REG_26__SCAN_IN), .ZN(n9960) );
  NOR2_X1 U10796 ( .A1(n9719), .A2(n9960), .ZN(P1_U3297) );
  AND2_X1 U10797 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n9720), .ZN(P1_U3298) );
  AND2_X1 U10798 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n9720), .ZN(P1_U3299) );
  AND2_X1 U10799 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n9720), .ZN(P1_U3300) );
  AND2_X1 U10800 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n9720), .ZN(P1_U3301) );
  AND2_X1 U10801 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n9720), .ZN(P1_U3302) );
  AND2_X1 U10802 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n9720), .ZN(P1_U3303) );
  AND2_X1 U10803 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n9720), .ZN(P1_U3304) );
  AND2_X1 U10804 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n9720), .ZN(P1_U3305) );
  AND2_X1 U10805 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n9720), .ZN(P1_U3306) );
  AND2_X1 U10806 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n9720), .ZN(P1_U3307) );
  AND2_X1 U10807 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n9720), .ZN(P1_U3308) );
  AND2_X1 U10808 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n9720), .ZN(P1_U3309) );
  AND2_X1 U10809 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n9720), .ZN(P1_U3310) );
  AND2_X1 U10810 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n9720), .ZN(P1_U3311) );
  AND2_X1 U10811 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n9720), .ZN(P1_U3312) );
  AND2_X1 U10812 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n9720), .ZN(P1_U3313) );
  INV_X1 U10813 ( .A(P1_D_REG_9__SCAN_IN), .ZN(n9933) );
  NOR2_X1 U10814 ( .A1(n9719), .A2(n9933), .ZN(P1_U3314) );
  AND2_X1 U10815 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n9720), .ZN(P1_U3315) );
  AND2_X1 U10816 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n9720), .ZN(P1_U3316) );
  AND2_X1 U10817 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n9720), .ZN(P1_U3317) );
  AND2_X1 U10818 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n9720), .ZN(P1_U3318) );
  AND2_X1 U10819 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n9720), .ZN(P1_U3319) );
  AND2_X1 U10820 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n9720), .ZN(P1_U3320) );
  AND2_X1 U10821 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n9720), .ZN(P1_U3321) );
  INV_X1 U10822 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n10025) );
  AOI21_X1 U10823 ( .B1(n9722), .B2(n10025), .A(n9721), .ZN(P1_U3441) );
  OAI21_X1 U10824 ( .B1(n9768), .B2(n9724), .A(n9723), .ZN(n9726) );
  AOI211_X1 U10825 ( .C1(n9773), .C2(n9727), .A(n9726), .B(n9725), .ZN(n9777)
         );
  AOI22_X1 U10826 ( .A1(n9776), .A2(n9777), .B1(n5978), .B2(n9774), .ZN(
        P1_U3457) );
  AOI22_X1 U10827 ( .A1(n9776), .A2(n9728), .B1(n5994), .B2(n9774), .ZN(
        P1_U3460) );
  NAND2_X1 U10828 ( .A1(n9736), .A2(n9729), .ZN(n9730) );
  OAI21_X1 U10829 ( .B1(n9731), .B2(n9754), .A(n9730), .ZN(n9733) );
  AOI211_X1 U10830 ( .C1(n9773), .C2(n9734), .A(n9733), .B(n9732), .ZN(n9778)
         );
  AOI22_X1 U10831 ( .A1(n9776), .A2(n9778), .B1(n6014), .B2(n9774), .ZN(
        P1_U3463) );
  AOI22_X1 U10832 ( .A1(n9738), .A2(n9737), .B1(n9736), .B2(n9735), .ZN(n9739)
         );
  OAI21_X1 U10833 ( .B1(n9741), .B2(n9740), .A(n9739), .ZN(n9742) );
  NOR2_X1 U10834 ( .A1(n9743), .A2(n9742), .ZN(n9779) );
  INV_X1 U10835 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n9744) );
  AOI22_X1 U10836 ( .A1(n9776), .A2(n9779), .B1(n9744), .B2(n9774), .ZN(
        P1_U3466) );
  NOR3_X1 U10837 ( .A1(n9747), .A2(n9746), .A3(n9745), .ZN(n9751) );
  NOR4_X1 U10838 ( .A1(n9751), .A2(n9750), .A3(n9749), .A4(n9748), .ZN(n9780)
         );
  INV_X1 U10839 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n9752) );
  AOI22_X1 U10840 ( .A1(n9776), .A2(n9780), .B1(n9752), .B2(n9774), .ZN(
        P1_U3469) );
  INV_X1 U10841 ( .A(n7358), .ZN(n9753) );
  OAI22_X1 U10842 ( .A1(n9755), .A2(n9754), .B1(n9753), .B2(n9768), .ZN(n9757)
         );
  AOI211_X1 U10843 ( .C1(n9758), .C2(n9759), .A(n9757), .B(n9756), .ZN(n9781)
         );
  AOI22_X1 U10844 ( .A1(n9776), .A2(n9781), .B1(n6070), .B2(n9774), .ZN(
        P1_U3472) );
  AND2_X1 U10845 ( .A1(n9760), .A2(n9759), .ZN(n9764) );
  OAI21_X1 U10846 ( .B1(n9762), .B2(n9768), .A(n9761), .ZN(n9763) );
  NOR3_X1 U10847 ( .A1(n9765), .A2(n9764), .A3(n9763), .ZN(n9782) );
  INV_X1 U10848 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n9974) );
  AOI22_X1 U10849 ( .A1(n9776), .A2(n9782), .B1(n9974), .B2(n9774), .ZN(
        P1_U3475) );
  INV_X1 U10850 ( .A(n9766), .ZN(n9772) );
  OAI21_X1 U10851 ( .B1(n9769), .B2(n9768), .A(n9767), .ZN(n9771) );
  AOI211_X1 U10852 ( .C1(n9773), .C2(n9772), .A(n9771), .B(n9770), .ZN(n9784)
         );
  INV_X1 U10853 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n9775) );
  AOI22_X1 U10854 ( .A1(n9776), .A2(n9784), .B1(n9775), .B2(n9774), .ZN(
        P1_U3478) );
  AOI22_X1 U10855 ( .A1(n9785), .A2(n9777), .B1(n5979), .B2(n9783), .ZN(
        P1_U3524) );
  AOI22_X1 U10856 ( .A1(n9785), .A2(n9778), .B1(n6664), .B2(n9783), .ZN(
        P1_U3526) );
  AOI22_X1 U10857 ( .A1(n9785), .A2(n9779), .B1(n6667), .B2(n9783), .ZN(
        P1_U3527) );
  AOI22_X1 U10858 ( .A1(n9785), .A2(n9780), .B1(n6054), .B2(n9783), .ZN(
        P1_U3528) );
  AOI22_X1 U10859 ( .A1(n9785), .A2(n9781), .B1(n6669), .B2(n9783), .ZN(
        P1_U3529) );
  AOI22_X1 U10860 ( .A1(n9785), .A2(n9782), .B1(n6672), .B2(n9783), .ZN(
        P1_U3530) );
  AOI22_X1 U10861 ( .A1(n9785), .A2(n9784), .B1(n6695), .B2(n9783), .ZN(
        P1_U3531) );
  OR2_X1 U10862 ( .A1(n9787), .A2(n9786), .ZN(n9789) );
  AOI21_X1 U10863 ( .B1(n9790), .B2(n9789), .A(n9788), .ZN(n9799) );
  AOI21_X1 U10864 ( .B1(n9793), .B2(n9792), .A(n9791), .ZN(n9794) );
  AOI21_X1 U10865 ( .B1(P2_REG3_REG_0__SCAN_IN), .B2(n9795), .A(n9794), .ZN(
        n9796) );
  OAI221_X1 U10866 ( .B1(n4262), .B2(n9799), .C1(n9798), .C2(n9797), .A(n9796), 
        .ZN(P2_U3296) );
  NOR2_X1 U10867 ( .A1(n9801), .A2(n9800), .ZN(n9802) );
  AND2_X1 U10868 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n9903), .ZN(P2_U3297) );
  AND2_X1 U10869 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n9903), .ZN(P2_U3298) );
  INV_X1 U10870 ( .A(P2_D_REG_29__SCAN_IN), .ZN(n9957) );
  NOR2_X1 U10871 ( .A1(n9802), .A2(n9957), .ZN(P2_U3299) );
  INV_X1 U10872 ( .A(P2_D_REG_28__SCAN_IN), .ZN(n10005) );
  NOR2_X1 U10873 ( .A1(n9802), .A2(n10005), .ZN(P2_U3300) );
  AND2_X1 U10874 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n9903), .ZN(P2_U3301) );
  AND2_X1 U10875 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n9903), .ZN(P2_U3302) );
  AND2_X1 U10876 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n9903), .ZN(P2_U3303) );
  AND2_X1 U10877 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n9903), .ZN(P2_U3304) );
  AND2_X1 U10878 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n9903), .ZN(P2_U3305) );
  AND2_X1 U10879 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n9903), .ZN(P2_U3306) );
  AND2_X1 U10880 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n9903), .ZN(P2_U3307) );
  AND2_X1 U10881 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n9903), .ZN(P2_U3308) );
  INV_X1 U10882 ( .A(P2_D_REG_19__SCAN_IN), .ZN(n9959) );
  NOR2_X1 U10883 ( .A1(n9802), .A2(n9959), .ZN(P2_U3309) );
  AND2_X1 U10884 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n9903), .ZN(P2_U3310) );
  AND2_X1 U10885 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n9903), .ZN(P2_U3311) );
  AND2_X1 U10886 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n9903), .ZN(P2_U3312) );
  AND2_X1 U10887 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n9903), .ZN(P2_U3313) );
  INV_X1 U10888 ( .A(P2_D_REG_14__SCAN_IN), .ZN(n9940) );
  NOR2_X1 U10889 ( .A1(n9802), .A2(n9940), .ZN(P2_U3314) );
  AND2_X1 U10890 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n9903), .ZN(P2_U3315) );
  AND2_X1 U10891 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n9903), .ZN(P2_U3316) );
  AND2_X1 U10892 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n9903), .ZN(P2_U3317) );
  AND2_X1 U10893 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n9903), .ZN(P2_U3319) );
  AND2_X1 U10894 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n9903), .ZN(P2_U3320) );
  AND2_X1 U10895 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n9903), .ZN(P2_U3321) );
  AND2_X1 U10896 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n9903), .ZN(P2_U3322) );
  AND2_X1 U10897 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n9903), .ZN(P2_U3323) );
  AND2_X1 U10898 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n9903), .ZN(P2_U3324) );
  AND2_X1 U10899 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n9903), .ZN(P2_U3325) );
  AND2_X1 U10900 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n9903), .ZN(P2_U3326) );
  AOI22_X1 U10901 ( .A1(n9804), .A2(n9806), .B1(n9803), .B2(n9903), .ZN(
        P2_U3437) );
  AOI22_X1 U10902 ( .A1(n9807), .A2(n9806), .B1(n9805), .B2(n9903), .ZN(
        P2_U3438) );
  AOI22_X1 U10903 ( .A1(n9862), .A2(n9808), .B1(n4525), .B2(n9860), .ZN(
        P2_U3451) );
  INV_X1 U10904 ( .A(n9809), .ZN(n9816) );
  NAND3_X1 U10905 ( .A1(n4648), .A2(n9811), .A3(n9810), .ZN(n9812) );
  OAI21_X1 U10906 ( .B1(n9854), .B2(n4823), .A(n9812), .ZN(n9815) );
  INV_X1 U10907 ( .A(n9813), .ZN(n9814) );
  AOI211_X1 U10908 ( .C1(n9851), .C2(n9816), .A(n9815), .B(n9814), .ZN(n9863)
         );
  AOI22_X1 U10909 ( .A1(n9862), .A2(n9863), .B1(n5033), .B2(n9860), .ZN(
        P2_U3454) );
  AOI22_X1 U10910 ( .A1(n9862), .A2(n9817), .B1(n5050), .B2(n9860), .ZN(
        P2_U3457) );
  INV_X1 U10911 ( .A(n9818), .ZN(n9859) );
  AND2_X1 U10912 ( .A1(n9819), .A2(n9859), .ZN(n9824) );
  OAI21_X1 U10913 ( .B1(n9854), .B2(n9821), .A(n9820), .ZN(n9822) );
  NOR3_X1 U10914 ( .A1(n9824), .A2(n9823), .A3(n9822), .ZN(n9864) );
  INV_X1 U10915 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n9825) );
  AOI22_X1 U10916 ( .A1(n9862), .A2(n9864), .B1(n9825), .B2(n9860), .ZN(
        P2_U3460) );
  INV_X1 U10917 ( .A(n9826), .ZN(n9831) );
  OAI211_X1 U10918 ( .C1(n9854), .C2(n9829), .A(n9828), .B(n9827), .ZN(n9830)
         );
  AOI21_X1 U10919 ( .B1(n9851), .B2(n9831), .A(n9830), .ZN(n9865) );
  INV_X1 U10920 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n9832) );
  AOI22_X1 U10921 ( .A1(n9862), .A2(n9865), .B1(n9832), .B2(n9860), .ZN(
        P2_U3463) );
  AND2_X1 U10922 ( .A1(n9833), .A2(n9851), .ZN(n9837) );
  OAI21_X1 U10923 ( .B1(n9854), .B2(n9835), .A(n9834), .ZN(n9836) );
  NOR3_X1 U10924 ( .A1(n9838), .A2(n9837), .A3(n9836), .ZN(n9866) );
  INV_X1 U10925 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n9839) );
  AOI22_X1 U10926 ( .A1(n9862), .A2(n9866), .B1(n9839), .B2(n9860), .ZN(
        P2_U3466) );
  OAI211_X1 U10927 ( .C1(n9854), .C2(n9842), .A(n9841), .B(n9840), .ZN(n9843)
         );
  AOI21_X1 U10928 ( .B1(n9844), .B2(n9851), .A(n9843), .ZN(n9867) );
  INV_X1 U10929 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n9845) );
  AOI22_X1 U10930 ( .A1(n9862), .A2(n9867), .B1(n9845), .B2(n9860), .ZN(
        P2_U3469) );
  OAI22_X1 U10931 ( .A1(n9847), .A2(n5873), .B1(n9854), .B2(n9846), .ZN(n9849)
         );
  AOI211_X1 U10932 ( .C1(n9851), .C2(n9850), .A(n9849), .B(n9848), .ZN(n9869)
         );
  INV_X1 U10933 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n9852) );
  AOI22_X1 U10934 ( .A1(n9862), .A2(n9869), .B1(n9852), .B2(n9860), .ZN(
        P2_U3472) );
  INV_X1 U10935 ( .A(n9853), .ZN(n9858) );
  OAI22_X1 U10936 ( .A1(n9855), .A2(n5873), .B1(n9854), .B2(n4643), .ZN(n9857)
         );
  AOI211_X1 U10937 ( .C1(n9859), .C2(n9858), .A(n9857), .B(n9856), .ZN(n9873)
         );
  INV_X1 U10938 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n9861) );
  AOI22_X1 U10939 ( .A1(n9862), .A2(n9873), .B1(n9861), .B2(n9860), .ZN(
        P2_U3475) );
  AOI22_X1 U10940 ( .A1(n9870), .A2(n9863), .B1(n6721), .B2(n9871), .ZN(
        P2_U3521) );
  AOI22_X1 U10941 ( .A1(n9870), .A2(n9864), .B1(n6735), .B2(n9871), .ZN(
        P2_U3523) );
  AOI22_X1 U10942 ( .A1(n9874), .A2(n9865), .B1(n6768), .B2(n9871), .ZN(
        P2_U3524) );
  AOI22_X1 U10943 ( .A1(n9870), .A2(n9866), .B1(n6771), .B2(n9871), .ZN(
        P2_U3525) );
  AOI22_X1 U10944 ( .A1(n9870), .A2(n9867), .B1(n6834), .B2(n9871), .ZN(
        P2_U3526) );
  AOI22_X1 U10945 ( .A1(n9870), .A2(n9869), .B1(n9868), .B2(n9871), .ZN(
        P2_U3527) );
  AOI22_X1 U10946 ( .A1(n9874), .A2(n9873), .B1(n9872), .B2(n9871), .ZN(
        P2_U3528) );
  INV_X1 U10947 ( .A(n9875), .ZN(n9876) );
  NAND2_X1 U10948 ( .A1(n9877), .A2(n9876), .ZN(n9878) );
  XNOR2_X1 U10949 ( .A(P2_ADDR_REG_1__SCAN_IN), .B(n9878), .ZN(ADD_1071_U5) );
  XOR2_X1 U10950 ( .A(P1_ADDR_REG_0__SCAN_IN), .B(P2_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1071_U46) );
  OAI21_X1 U10951 ( .B1(n9881), .B2(n9880), .A(n9879), .ZN(ADD_1071_U56) );
  OAI21_X1 U10952 ( .B1(n9884), .B2(n9883), .A(n9882), .ZN(ADD_1071_U57) );
  OAI21_X1 U10953 ( .B1(n9887), .B2(n9886), .A(n9885), .ZN(ADD_1071_U58) );
  OAI21_X1 U10954 ( .B1(n9890), .B2(n9889), .A(n9888), .ZN(ADD_1071_U59) );
  OAI21_X1 U10955 ( .B1(n9893), .B2(n9892), .A(n9891), .ZN(ADD_1071_U60) );
  OAI21_X1 U10956 ( .B1(n9896), .B2(n9895), .A(n9894), .ZN(ADD_1071_U61) );
  AOI21_X1 U10957 ( .B1(n9899), .B2(n9898), .A(n9897), .ZN(ADD_1071_U62) );
  AOI21_X1 U10958 ( .B1(n9902), .B2(n9901), .A(n9900), .ZN(ADD_1071_U63) );
  NAND2_X1 U10959 ( .A1(n9903), .A2(P2_D_REG_10__SCAN_IN), .ZN(n10052) );
  NAND4_X1 U10960 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .A3(P1_ADDR_REG_4__SCAN_IN), .A4(n10030), .ZN(n9908) );
  INV_X1 U10961 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n9945) );
  NAND4_X1 U10962 ( .A1(P2_IR_REG_4__SCAN_IN), .A2(P2_IR_REG_19__SCAN_IN), 
        .A3(P2_IR_REG_1__SCAN_IN), .A4(n9945), .ZN(n9907) );
  NAND4_X1 U10963 ( .A1(P1_REG0_REG_11__SCAN_IN), .A2(P1_D_REG_9__SCAN_IN), 
        .A3(P2_IR_REG_24__SCAN_IN), .A4(n8412), .ZN(n9906) );
  NAND4_X1 U10964 ( .A1(P1_REG1_REG_5__SCAN_IN), .A2(P2_D_REG_14__SCAN_IN), 
        .A3(n9904), .A4(n9932), .ZN(n9905) );
  NOR4_X1 U10965 ( .A1(n9908), .A2(n9907), .A3(n9906), .A4(n9905), .ZN(n10050)
         );
  NAND3_X1 U10966 ( .A1(P1_RD_REG_SCAN_IN), .A2(SI_6_), .A3(
        P2_REG1_REG_29__SCAN_IN), .ZN(n9930) );
  NOR4_X1 U10967 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n10006), .A3(n10003), .A4(
        n6771), .ZN(n9913) );
  NOR4_X1 U10968 ( .A1(P1_IR_REG_28__SCAN_IN), .A2(P2_REG0_REG_12__SCAN_IN), 
        .A3(n7377), .A4(n4525), .ZN(n9912) );
  NOR4_X1 U10969 ( .A1(n9910), .A2(n9909), .A3(P2_REG2_REG_13__SCAN_IN), .A4(
        P1_REG0_REG_7__SCAN_IN), .ZN(n9911) );
  NAND3_X1 U10970 ( .A1(n9913), .A2(n9912), .A3(n9911), .ZN(n9929) );
  NOR4_X1 U10971 ( .A1(P2_DATAO_REG_7__SCAN_IN), .A2(P1_REG0_REG_1__SCAN_IN), 
        .A3(P2_D_REG_29__SCAN_IN), .A4(n9963), .ZN(n9927) );
  NAND4_X1 U10972 ( .A1(P1_REG1_REG_31__SCAN_IN), .A2(n9972), .A3(n9976), .A4(
        n9977), .ZN(n9914) );
  OR4_X1 U10973 ( .A1(P2_REG3_REG_1__SCAN_IN), .A2(n4503), .A3(
        P1_DATAO_REG_0__SCAN_IN), .A4(n9914), .ZN(n9917) );
  NAND3_X1 U10974 ( .A1(P1_D_REG_26__SCAN_IN), .A2(P2_DATAO_REG_6__SCAN_IN), 
        .A3(P2_D_REG_19__SCAN_IN), .ZN(n9916) );
  INV_X1 U10975 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n9915) );
  NOR4_X1 U10976 ( .A1(n9917), .A2(n9916), .A3(P1_REG3_REG_8__SCAN_IN), .A4(
        n9915), .ZN(n9926) );
  NOR4_X1 U10977 ( .A1(P1_REG3_REG_19__SCAN_IN), .A2(P2_REG3_REG_22__SCAN_IN), 
        .A3(n10033), .A4(n5304), .ZN(n9925) );
  INV_X1 U10978 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n9918) );
  NAND4_X1 U10979 ( .A1(P2_DATAO_REG_27__SCAN_IN), .A2(P1_IR_REG_14__SCAN_IN), 
        .A3(P1_DATAO_REG_3__SCAN_IN), .A4(n9918), .ZN(n9920) );
  NAND3_X1 U10980 ( .A1(P1_IR_REG_25__SCAN_IN), .A2(P1_DATAO_REG_26__SCAN_IN), 
        .A3(n10025), .ZN(n9919) );
  NOR3_X1 U10981 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(n9920), .A3(n9919), .ZN(
        n9922) );
  INV_X1 U10982 ( .A(SI_3_), .ZN(n9921) );
  NAND3_X1 U10983 ( .A1(n9922), .A2(P1_IR_REG_30__SCAN_IN), .A3(n9921), .ZN(
        n9923) );
  NOR3_X1 U10984 ( .A1(n9923), .A2(n10035), .A3(n10036), .ZN(n9924) );
  NAND4_X1 U10985 ( .A1(n9927), .A2(n9926), .A3(n9925), .A4(n9924), .ZN(n9928)
         );
  NOR4_X1 U10986 ( .A1(P2_DATAO_REG_28__SCAN_IN), .A2(n9930), .A3(n9929), .A4(
        n9928), .ZN(n10049) );
  AOI22_X1 U10987 ( .A1(n6054), .A2(keyinput45), .B1(keyinput22), .B2(n9932), 
        .ZN(n9931) );
  OAI221_X1 U10988 ( .B1(n6054), .B2(keyinput45), .C1(n9932), .C2(keyinput22), 
        .A(n9931), .ZN(n9936) );
  XNOR2_X1 U10989 ( .A(n9933), .B(keyinput17), .ZN(n9935) );
  XOR2_X1 U10990 ( .A(P2_IR_REG_4__SCAN_IN), .B(keyinput5), .Z(n9934) );
  OR3_X1 U10991 ( .A1(n9936), .A2(n9935), .A3(n9934), .ZN(n9943) );
  AOI22_X1 U10992 ( .A1(n9938), .A2(keyinput18), .B1(keyinput52), .B2(n8412), 
        .ZN(n9937) );
  OAI221_X1 U10993 ( .B1(n9938), .B2(keyinput18), .C1(n8412), .C2(keyinput52), 
        .A(n9937), .ZN(n9942) );
  AOI22_X1 U10994 ( .A1(n9940), .A2(keyinput36), .B1(n5025), .B2(keyinput58), 
        .ZN(n9939) );
  OAI221_X1 U10995 ( .B1(n9940), .B2(keyinput36), .C1(n5025), .C2(keyinput58), 
        .A(n9939), .ZN(n9941) );
  NOR3_X1 U10996 ( .A1(n9943), .A2(n9942), .A3(n9941), .ZN(n9987) );
  XOR2_X1 U10997 ( .A(n9944), .B(keyinput27), .Z(n9949) );
  XOR2_X1 U10998 ( .A(n9945), .B(keyinput13), .Z(n9948) );
  XNOR2_X1 U10999 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(keyinput28), .ZN(n9947) );
  XNOR2_X1 U11000 ( .A(P2_IR_REG_29__SCAN_IN), .B(keyinput29), .ZN(n9946) );
  NAND4_X1 U11001 ( .A1(n9949), .A2(n9948), .A3(n9947), .A4(n9946), .ZN(n9955)
         );
  XNOR2_X1 U11002 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(keyinput53), .ZN(n9953)
         );
  XNOR2_X1 U11003 ( .A(P2_REG3_REG_1__SCAN_IN), .B(keyinput0), .ZN(n9952) );
  XNOR2_X1 U11004 ( .A(P2_REG0_REG_30__SCAN_IN), .B(keyinput3), .ZN(n9951) );
  XNOR2_X1 U11005 ( .A(P1_REG3_REG_8__SCAN_IN), .B(keyinput62), .ZN(n9950) );
  NAND4_X1 U11006 ( .A1(n9953), .A2(n9952), .A3(n9951), .A4(n9950), .ZN(n9954)
         );
  NOR2_X1 U11007 ( .A1(n9955), .A2(n9954), .ZN(n9986) );
  AOI22_X1 U11008 ( .A1(n5978), .A2(keyinput37), .B1(keyinput44), .B2(n9957), 
        .ZN(n9956) );
  OAI221_X1 U11009 ( .B1(n5978), .B2(keyinput37), .C1(n9957), .C2(keyinput44), 
        .A(n9956), .ZN(n9970) );
  AOI22_X1 U11010 ( .A1(n9960), .A2(keyinput32), .B1(keyinput23), .B2(n9959), 
        .ZN(n9958) );
  OAI221_X1 U11011 ( .B1(n9960), .B2(keyinput32), .C1(n9959), .C2(keyinput23), 
        .A(n9958), .ZN(n9969) );
  AOI22_X1 U11012 ( .A1(n9963), .A2(keyinput20), .B1(keyinput9), .B2(n9962), 
        .ZN(n9961) );
  OAI221_X1 U11013 ( .B1(n9963), .B2(keyinput20), .C1(n9962), .C2(keyinput9), 
        .A(n9961), .ZN(n9967) );
  XNOR2_X1 U11014 ( .A(n9964), .B(keyinput56), .ZN(n9966) );
  XOR2_X1 U11015 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(keyinput50), .Z(n9965) );
  OR3_X1 U11016 ( .A1(n9967), .A2(n9966), .A3(n9965), .ZN(n9968) );
  NOR3_X1 U11017 ( .A1(n9970), .A2(n9969), .A3(n9968), .ZN(n9985) );
  AOI22_X1 U11018 ( .A1(n9972), .A2(keyinput7), .B1(keyinput11), .B2(n5732), 
        .ZN(n9971) );
  OAI221_X1 U11019 ( .B1(n9972), .B2(keyinput7), .C1(n5732), .C2(keyinput11), 
        .A(n9971), .ZN(n9983) );
  AOI22_X1 U11020 ( .A1(n9974), .A2(keyinput16), .B1(keyinput40), .B2(n7791), 
        .ZN(n9973) );
  OAI221_X1 U11021 ( .B1(n9974), .B2(keyinput16), .C1(n7791), .C2(keyinput40), 
        .A(n9973), .ZN(n9982) );
  AOI22_X1 U11022 ( .A1(n9977), .A2(keyinput39), .B1(n9976), .B2(keyinput12), 
        .ZN(n9975) );
  OAI221_X1 U11023 ( .B1(n9977), .B2(keyinput39), .C1(n9976), .C2(keyinput12), 
        .A(n9975), .ZN(n9981) );
  XOR2_X1 U11024 ( .A(n9909), .B(keyinput30), .Z(n9979) );
  XNOR2_X1 U11025 ( .A(P1_IR_REG_12__SCAN_IN), .B(keyinput38), .ZN(n9978) );
  NAND2_X1 U11026 ( .A1(n9979), .A2(n9978), .ZN(n9980) );
  NOR4_X1 U11027 ( .A1(n9983), .A2(n9982), .A3(n9981), .A4(n9980), .ZN(n9984)
         );
  NAND4_X1 U11028 ( .A1(n9987), .A2(n9986), .A3(n9985), .A4(n9984), .ZN(n10048) );
  INV_X1 U11029 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n9989) );
  AOI22_X1 U11030 ( .A1(n9990), .A2(keyinput48), .B1(keyinput34), .B2(n9989), 
        .ZN(n9988) );
  OAI221_X1 U11031 ( .B1(n9990), .B2(keyinput48), .C1(n9989), .C2(keyinput34), 
        .A(n9988), .ZN(n10001) );
  INV_X1 U11032 ( .A(P1_RD_REG_SCAN_IN), .ZN(n9992) );
  AOI22_X1 U11033 ( .A1(n9993), .A2(keyinput15), .B1(n9992), .B2(keyinput10), 
        .ZN(n9991) );
  OAI221_X1 U11034 ( .B1(n9993), .B2(keyinput15), .C1(n9992), .C2(keyinput10), 
        .A(n9991), .ZN(n10000) );
  XOR2_X1 U11035 ( .A(n5555), .B(keyinput2), .Z(n9996) );
  XNOR2_X1 U11036 ( .A(SI_6_), .B(keyinput47), .ZN(n9995) );
  XNOR2_X1 U11037 ( .A(P2_REG3_REG_6__SCAN_IN), .B(keyinput19), .ZN(n9994) );
  NAND3_X1 U11038 ( .A1(n9996), .A2(n9995), .A3(n9994), .ZN(n9999) );
  XNOR2_X1 U11039 ( .A(n9997), .B(keyinput54), .ZN(n9998) );
  NOR4_X1 U11040 ( .A1(n10001), .A2(n10000), .A3(n9999), .A4(n9998), .ZN(
        n10046) );
  AOI22_X1 U11041 ( .A1(n6771), .A2(keyinput8), .B1(n10003), .B2(keyinput60), 
        .ZN(n10002) );
  OAI221_X1 U11042 ( .B1(n6771), .B2(keyinput8), .C1(n10003), .C2(keyinput60), 
        .A(n10002), .ZN(n10013) );
  AOI22_X1 U11043 ( .A1(n10006), .A2(keyinput49), .B1(keyinput59), .B2(n10005), 
        .ZN(n10004) );
  OAI221_X1 U11044 ( .B1(n10006), .B2(keyinput49), .C1(n10005), .C2(keyinput59), .A(n10004), .ZN(n10012) );
  AOI22_X1 U11045 ( .A1(n4525), .A2(keyinput46), .B1(n5963), .B2(keyinput31), 
        .ZN(n10007) );
  OAI221_X1 U11046 ( .B1(n4525), .B2(keyinput46), .C1(n5963), .C2(keyinput31), 
        .A(n10007), .ZN(n10011) );
  INV_X1 U11047 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n10009) );
  AOI22_X1 U11048 ( .A1(n10009), .A2(keyinput6), .B1(n7377), .B2(keyinput43), 
        .ZN(n10008) );
  OAI221_X1 U11049 ( .B1(n10009), .B2(keyinput6), .C1(n7377), .C2(keyinput43), 
        .A(n10008), .ZN(n10010) );
  NOR4_X1 U11050 ( .A1(n10013), .A2(n10012), .A3(n10011), .A4(n10010), .ZN(
        n10045) );
  INV_X1 U11051 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n10016) );
  AOI22_X1 U11052 ( .A1(n10016), .A2(keyinput4), .B1(n10015), .B2(keyinput21), 
        .ZN(n10014) );
  OAI221_X1 U11053 ( .B1(n10016), .B2(keyinput4), .C1(n10015), .C2(keyinput21), 
        .A(n10014), .ZN(n10020) );
  XNOR2_X1 U11054 ( .A(n10017), .B(keyinput14), .ZN(n10019) );
  XOR2_X1 U11055 ( .A(P2_REG0_REG_16__SCAN_IN), .B(keyinput57), .Z(n10018) );
  NOR3_X1 U11056 ( .A1(n10020), .A2(n10019), .A3(n10018), .ZN(n10024) );
  XNOR2_X1 U11057 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(keyinput33), .ZN(n10023)
         );
  XNOR2_X1 U11058 ( .A(P1_IR_REG_14__SCAN_IN), .B(keyinput24), .ZN(n10022) );
  XNOR2_X1 U11059 ( .A(P1_IR_REG_25__SCAN_IN), .B(keyinput61), .ZN(n10021) );
  NAND4_X1 U11060 ( .A1(n10024), .A2(n10023), .A3(n10022), .A4(n10021), .ZN(
        n10027) );
  XNOR2_X1 U11061 ( .A(n10025), .B(keyinput25), .ZN(n10026) );
  NOR2_X1 U11062 ( .A1(n10027), .A2(n10026), .ZN(n10044) );
  AOI22_X1 U11063 ( .A1(n10030), .A2(keyinput55), .B1(n10029), .B2(keyinput26), 
        .ZN(n10028) );
  OAI221_X1 U11064 ( .B1(n10030), .B2(keyinput55), .C1(n10029), .C2(keyinput26), .A(n10028), .ZN(n10042) );
  AOI22_X1 U11065 ( .A1(n10033), .A2(keyinput42), .B1(keyinput51), .B2(n10032), 
        .ZN(n10031) );
  OAI221_X1 U11066 ( .B1(n10033), .B2(keyinput42), .C1(n10032), .C2(keyinput51), .A(n10031), .ZN(n10041) );
  AOI22_X1 U11067 ( .A1(n10036), .A2(keyinput41), .B1(n10035), .B2(keyinput1), 
        .ZN(n10034) );
  OAI221_X1 U11068 ( .B1(n10036), .B2(keyinput41), .C1(n10035), .C2(keyinput1), 
        .A(n10034), .ZN(n10040) );
  XOR2_X1 U11069 ( .A(n5304), .B(keyinput63), .Z(n10038) );
  XNOR2_X1 U11070 ( .A(SI_3_), .B(keyinput35), .ZN(n10037) );
  NAND2_X1 U11071 ( .A1(n10038), .A2(n10037), .ZN(n10039) );
  NOR4_X1 U11072 ( .A1(n10042), .A2(n10041), .A3(n10040), .A4(n10039), .ZN(
        n10043) );
  NAND4_X1 U11073 ( .A1(n10046), .A2(n10045), .A3(n10044), .A4(n10043), .ZN(
        n10047) );
  AOI211_X1 U11074 ( .C1(n10050), .C2(n10049), .A(n10048), .B(n10047), .ZN(
        n10051) );
  XNOR2_X1 U11075 ( .A(n10052), .B(n10051), .ZN(P2_U3318) );
  XOR2_X1 U11076 ( .A(n10053), .B(P2_ADDR_REG_6__SCAN_IN), .Z(ADD_1071_U50) );
  NOR2_X1 U11077 ( .A1(n10055), .A2(n10054), .ZN(n10056) );
  XOR2_X1 U11078 ( .A(P1_ADDR_REG_5__SCAN_IN), .B(n10056), .Z(ADD_1071_U51) );
  XOR2_X1 U11079 ( .A(n10057), .B(P2_ADDR_REG_7__SCAN_IN), .Z(ADD_1071_U49) );
  OAI21_X1 U11080 ( .B1(n10060), .B2(n10059), .A(n10058), .ZN(n10061) );
  XNOR2_X1 U11081 ( .A(n10061), .B(P1_ADDR_REG_18__SCAN_IN), .ZN(ADD_1071_U55)
         );
  XOR2_X1 U11082 ( .A(n10062), .B(P2_ADDR_REG_8__SCAN_IN), .Z(ADD_1071_U48) );
  AOI21_X1 U11083 ( .B1(n10065), .B2(n10064), .A(n10063), .ZN(ADD_1071_U47) );
  XOR2_X1 U11084 ( .A(n10067), .B(n10066), .Z(ADD_1071_U54) );
  XOR2_X1 U11085 ( .A(n10068), .B(n10069), .Z(ADD_1071_U53) );
  XNOR2_X1 U11086 ( .A(n10071), .B(n10070), .ZN(ADD_1071_U52) );
  INV_X1 U6575 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n5208) );
  NAND4_X2 U4973 ( .A1(n5998), .A2(n5997), .A3(n5996), .A4(n5995), .ZN(n6893)
         );
  INV_X1 U4835 ( .A(n7145), .ZN(n9829) );
  BUF_X1 U4846 ( .A(n6274), .Z(n8822) );
  NAND2_X1 U6315 ( .A1(n4644), .A2(n4643), .ZN(n7439) );
  NAND2_X1 U6373 ( .A1(n4827), .A2(n4825), .ZN(n5841) );
  INV_X1 U4805 ( .A(n5586), .ZN(n7017) );
  NOR2_X1 U4774 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(P1_IR_REG_7__SCAN_IN), .ZN(
        n5917) );
  CLKBUF_X1 U4790 ( .A(n5549), .Z(n6722) );
  CLKBUF_X3 U5194 ( .A(n5056), .Z(n5507) );
  CLKBUF_X1 U6119 ( .A(n5774), .Z(n5851) );
  AND2_X2 U6196 ( .A1(n8296), .A2(n8290), .ZN(n8286) );
  AND2_X2 U7471 ( .A1(n7570), .A2(n7575), .ZN(n4259) );
endmodule

