

module b20_C_lock ( keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, 
        keyinput_5, keyinput_6, keyinput_7, keyinput_8, keyinput_9, 
        keyinput_10, keyinput_11, keyinput_12, keyinput_13, keyinput_14, 
        keyinput_15, keyinput_16, keyinput_17, keyinput_18, keyinput_19, 
        keyinput_20, keyinput_21, keyinput_22, keyinput_23, keyinput_24, 
        keyinput_25, keyinput_26, keyinput_27, keyinput_28, keyinput_29, 
        keyinput_30, keyinput_31, keyinput_32, keyinput_33, keyinput_34, 
        keyinput_35, keyinput_36, keyinput_37, keyinput_38, keyinput_39, 
        keyinput_40, keyinput_41, keyinput_42, keyinput_43, keyinput_44, 
        keyinput_45, keyinput_46, keyinput_47, keyinput_48, keyinput_49, 
        keyinput_50, keyinput_51, keyinput_52, keyinput_53, keyinput_54, 
        keyinput_55, keyinput_56, keyinput_57, keyinput_58, keyinput_59, 
        keyinput_60, keyinput_61, keyinput_62, keyinput_63, keyinput_64, 
        keyinput_65, keyinput_66, keyinput_67, keyinput_68, keyinput_69, 
        keyinput_70, keyinput_71, keyinput_72, keyinput_73, keyinput_74, 
        keyinput_75, keyinput_76, keyinput_77, keyinput_78, keyinput_79, 
        keyinput_80, keyinput_81, keyinput_82, keyinput_83, keyinput_84, 
        keyinput_85, keyinput_86, keyinput_87, keyinput_88, keyinput_89, 
        keyinput_90, keyinput_91, keyinput_92, keyinput_93, keyinput_94, 
        keyinput_95, keyinput_96, keyinput_97, keyinput_98, keyinput_99, 
        keyinput_100, keyinput_101, keyinput_102, keyinput_103, keyinput_104, 
        keyinput_105, keyinput_106, keyinput_107, keyinput_108, keyinput_109, 
        keyinput_110, keyinput_111, keyinput_112, keyinput_113, keyinput_114, 
        keyinput_115, keyinput_116, keyinput_117, keyinput_118, keyinput_119, 
        keyinput_120, keyinput_121, keyinput_122, keyinput_123, keyinput_124, 
        keyinput_125, keyinput_126, keyinput_127, keyinput_128, keyinput_129, 
        keyinput_130, keyinput_131, keyinput_132, keyinput_133, keyinput_134, 
        keyinput_135, keyinput_136, keyinput_137, keyinput_138, keyinput_139, 
        keyinput_140, keyinput_141, keyinput_142, keyinput_143, keyinput_144, 
        keyinput_145, keyinput_146, keyinput_147, keyinput_148, keyinput_149, 
        keyinput_150, keyinput_151, keyinput_152, keyinput_153, keyinput_154, 
        keyinput_155, keyinput_156, keyinput_157, keyinput_158, keyinput_159, 
        keyinput_160, keyinput_161, keyinput_162, keyinput_163, keyinput_164, 
        keyinput_165, keyinput_166, keyinput_167, keyinput_168, keyinput_169, 
        keyinput_170, keyinput_171, keyinput_172, keyinput_173, keyinput_174, 
        keyinput_175, keyinput_176, keyinput_177, keyinput_178, keyinput_179, 
        keyinput_180, keyinput_181, keyinput_182, keyinput_183, keyinput_184, 
        keyinput_185, keyinput_186, keyinput_187, keyinput_188, keyinput_189, 
        keyinput_190, keyinput_191, keyinput_192, keyinput_193, keyinput_194, 
        keyinput_195, keyinput_196, keyinput_197, keyinput_198, keyinput_199, 
        keyinput_200, keyinput_201, keyinput_202, keyinput_203, keyinput_204, 
        keyinput_205, keyinput_206, keyinput_207, keyinput_208, keyinput_209, 
        keyinput_210, keyinput_211, keyinput_212, keyinput_213, keyinput_214, 
        keyinput_215, keyinput_216, keyinput_217, keyinput_218, keyinput_219, 
        keyinput_220, keyinput_221, keyinput_222, keyinput_223, keyinput_224, 
        keyinput_225, keyinput_226, keyinput_227, keyinput_228, keyinput_229, 
        keyinput_230, keyinput_231, keyinput_232, keyinput_233, keyinput_234, 
        keyinput_235, keyinput_236, keyinput_237, keyinput_238, keyinput_239, 
        keyinput_240, keyinput_241, keyinput_242, keyinput_243, keyinput_244, 
        keyinput_245, keyinput_246, keyinput_247, keyinput_248, keyinput_249, 
        keyinput_250, keyinput_251, keyinput_252, keyinput_253, keyinput_254, 
        keyinput_255, P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, 
        SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, 
        SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, 
        SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_, 
        P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, 
        P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, 
        P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, 
        P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, 
        P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, 
        P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, 
        P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, 
        P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, 
        P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, 
        P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, 
        P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, 
        P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, 
        P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, 
        P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, 
        P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, 
        P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, 
        P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, 
        P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, 
        P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, 
        P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, 
        P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, 
        P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, 
        P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, 
        P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, 
        P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, 
        P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN, 
        P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN, 
        P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN, 
        P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN, 
        P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN, 
        P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN, 
        P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN, 
        P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN, 
        P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN, 
        P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN, 
        P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN, 
        P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN, 
        P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN, 
        P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN, 
        P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN, 
        P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN, 
        P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN, 
        P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN, 
        P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN, 
        P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN, 
        P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN, 
        P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN, 
        P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN, 
        P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN, 
        P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN, 
        P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN, 
        P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, 
        P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, 
        P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, 
        P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN, 
        P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN, 
        P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN, 
        P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN, 
        P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN, 
        P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN, 
        P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN, 
        P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN, 
        P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN, 
        P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN, 
        P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN, 
        P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN, 
        P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN, 
        P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN, 
        P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN, 
        P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN, 
        P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN, 
        P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN, 
        P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN, 
        P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, 
        P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN, 
        P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN, 
        P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN, 
        P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN, 
        P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN, 
        P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, ADD_1068_U4, 
        ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58, ADD_1068_U59, 
        ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63, ADD_1068_U47, 
        ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51, ADD_1068_U52, 
        ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46, U126, U123, 
        P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349, 
        P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342, 
        P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335, 
        P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328, 
        P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439, P1_U3440, P1_U3323, 
        P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316, 
        P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309, 
        P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302, 
        P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295, 
        P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462, P1_U3465, P1_U3468, 
        P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, 
        P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3509, 
        P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515, P1_U3516, 
        P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, P1_U3523, 
        P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, P1_U3530, 
        P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, P1_U3537, 
        P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, P1_U3544, 
        P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, P1_U3551, 
        P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291, P1_U3290, P1_U3289, 
        P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282, 
        P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275, 
        P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268, 
        P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, P1_U3262, 
        P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255, 
        P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248, 
        P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3554, P1_U3555, 
        P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561, P1_U3562, 
        P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, P1_U3569, 
        P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, P1_U3576, 
        P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, P1_U3583, 
        P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240, P1_U3239, P1_U3238, 
        P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231, 
        P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224, 
        P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, 
        P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, P1_U3973, 
        P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, 
        P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, 
        P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, 
        P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, 
        P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376, P2_U3377, P2_U3263, 
        P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, 
        P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, 
        P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, 
        P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, 
        P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399, P2_U3402, P2_U3405, 
        P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420, P2_U3423, P2_U3426, 
        P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441, P2_U3444, P2_U3446, 
        P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451, P2_U3452, P2_U3453, 
        P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458, P2_U3459, P2_U3460, 
        P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465, P2_U3466, P2_U3467, 
        P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472, P2_U3473, P2_U3474, 
        P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479, P2_U3480, P2_U3481, 
        P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486, P2_U3487, P2_U3488, 
        P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, 
        P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, 
        P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, 
        P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3208, 
        P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, 
        P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, 
        P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, 
        P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3491, P2_U3492, 
        P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499, 
        P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506, 
        P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, 
        P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, 
        P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180, P2_U3179, P2_U3178, 
        P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172, P2_U3171, 
        P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165, P2_U3164, 
        P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158, P2_U3157, 
        P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151, P2_U3150, P2_U3893
 );
  input keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, keyinput_5,
         keyinput_6, keyinput_7, keyinput_8, keyinput_9, keyinput_10,
         keyinput_11, keyinput_12, keyinput_13, keyinput_14, keyinput_15,
         keyinput_16, keyinput_17, keyinput_18, keyinput_19, keyinput_20,
         keyinput_21, keyinput_22, keyinput_23, keyinput_24, keyinput_25,
         keyinput_26, keyinput_27, keyinput_28, keyinput_29, keyinput_30,
         keyinput_31, keyinput_32, keyinput_33, keyinput_34, keyinput_35,
         keyinput_36, keyinput_37, keyinput_38, keyinput_39, keyinput_40,
         keyinput_41, keyinput_42, keyinput_43, keyinput_44, keyinput_45,
         keyinput_46, keyinput_47, keyinput_48, keyinput_49, keyinput_50,
         keyinput_51, keyinput_52, keyinput_53, keyinput_54, keyinput_55,
         keyinput_56, keyinput_57, keyinput_58, keyinput_59, keyinput_60,
         keyinput_61, keyinput_62, keyinput_63, keyinput_64, keyinput_65,
         keyinput_66, keyinput_67, keyinput_68, keyinput_69, keyinput_70,
         keyinput_71, keyinput_72, keyinput_73, keyinput_74, keyinput_75,
         keyinput_76, keyinput_77, keyinput_78, keyinput_79, keyinput_80,
         keyinput_81, keyinput_82, keyinput_83, keyinput_84, keyinput_85,
         keyinput_86, keyinput_87, keyinput_88, keyinput_89, keyinput_90,
         keyinput_91, keyinput_92, keyinput_93, keyinput_94, keyinput_95,
         keyinput_96, keyinput_97, keyinput_98, keyinput_99, keyinput_100,
         keyinput_101, keyinput_102, keyinput_103, keyinput_104, keyinput_105,
         keyinput_106, keyinput_107, keyinput_108, keyinput_109, keyinput_110,
         keyinput_111, keyinput_112, keyinput_113, keyinput_114, keyinput_115,
         keyinput_116, keyinput_117, keyinput_118, keyinput_119, keyinput_120,
         keyinput_121, keyinput_122, keyinput_123, keyinput_124, keyinput_125,
         keyinput_126, keyinput_127, keyinput_128, keyinput_129, keyinput_130,
         keyinput_131, keyinput_132, keyinput_133, keyinput_134, keyinput_135,
         keyinput_136, keyinput_137, keyinput_138, keyinput_139, keyinput_140,
         keyinput_141, keyinput_142, keyinput_143, keyinput_144, keyinput_145,
         keyinput_146, keyinput_147, keyinput_148, keyinput_149, keyinput_150,
         keyinput_151, keyinput_152, keyinput_153, keyinput_154, keyinput_155,
         keyinput_156, keyinput_157, keyinput_158, keyinput_159, keyinput_160,
         keyinput_161, keyinput_162, keyinput_163, keyinput_164, keyinput_165,
         keyinput_166, keyinput_167, keyinput_168, keyinput_169, keyinput_170,
         keyinput_171, keyinput_172, keyinput_173, keyinput_174, keyinput_175,
         keyinput_176, keyinput_177, keyinput_178, keyinput_179, keyinput_180,
         keyinput_181, keyinput_182, keyinput_183, keyinput_184, keyinput_185,
         keyinput_186, keyinput_187, keyinput_188, keyinput_189, keyinput_190,
         keyinput_191, keyinput_192, keyinput_193, keyinput_194, keyinput_195,
         keyinput_196, keyinput_197, keyinput_198, keyinput_199, keyinput_200,
         keyinput_201, keyinput_202, keyinput_203, keyinput_204, keyinput_205,
         keyinput_206, keyinput_207, keyinput_208, keyinput_209, keyinput_210,
         keyinput_211, keyinput_212, keyinput_213, keyinput_214, keyinput_215,
         keyinput_216, keyinput_217, keyinput_218, keyinput_219, keyinput_220,
         keyinput_221, keyinput_222, keyinput_223, keyinput_224, keyinput_225,
         keyinput_226, keyinput_227, keyinput_228, keyinput_229, keyinput_230,
         keyinput_231, keyinput_232, keyinput_233, keyinput_234, keyinput_235,
         keyinput_236, keyinput_237, keyinput_238, keyinput_239, keyinput_240,
         keyinput_241, keyinput_242, keyinput_243, keyinput_244, keyinput_245,
         keyinput_246, keyinput_247, keyinput_248, keyinput_249, keyinput_250,
         keyinput_251, keyinput_252, keyinput_253, keyinput_254, keyinput_255,
         P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN,
         P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN,
         P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN,
         P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN,
         P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN,
         P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN,
         P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN,
         P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN,
         P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN,
         P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN,
         P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN,
         P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN,
         P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN,
         P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN,
         P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN,
         P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN,
         P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN,
         P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN,
         P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN,
         P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN,
         P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN,
         P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN,
         P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN,
         P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN,
         P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN,
         P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN,
         P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN,
         P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN,
         P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN,
         P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN,
         P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN,
         P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN,
         P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN,
         P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN,
         P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN,
         P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN,
         P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN,
         P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN,
         P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN,
         P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN,
         P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN,
         P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN,
         P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN,
         P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN,
         P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN,
         P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN,
         P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN,
         P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN,
         P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN,
         P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN,
         P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN,
         P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN,
         P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN,
         P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN,
         P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN,
         P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN,
         P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN,
         P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN,
         P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN,
         P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN,
         P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN,
         P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN,
         P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN,
         P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN,
         P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN,
         P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN,
         P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN,
         P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN,
         P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN,
         P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN,
         P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN,
         P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN,
         P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN,
         P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN,
         P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN,
         P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN,
         P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN,
         P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN,
         P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN,
         P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN,
         P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN,
         P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN,
         P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN,
         P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN,
         P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN,
         P1_REG3_REG_4__SCAN_IN, P1_REG3_REG_24__SCAN_IN,
         P1_REG3_REG_17__SCAN_IN, P1_REG3_REG_5__SCAN_IN,
         P1_REG3_REG_16__SCAN_IN, P1_REG3_REG_25__SCAN_IN,
         P1_REG3_REG_12__SCAN_IN, P1_REG3_REG_21__SCAN_IN,
         P1_REG3_REG_1__SCAN_IN, P1_REG3_REG_8__SCAN_IN,
         P1_REG3_REG_28__SCAN_IN, P1_REG3_REG_19__SCAN_IN,
         P1_REG3_REG_3__SCAN_IN, P1_REG3_REG_10__SCAN_IN,
         P1_REG3_REG_23__SCAN_IN, P1_REG3_REG_14__SCAN_IN,
         P1_REG3_REG_27__SCAN_IN, P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN,
         P1_RD_REG_SCAN_IN, P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN,
         P2_IR_REG_1__SCAN_IN, P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN,
         P2_IR_REG_4__SCAN_IN, P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN,
         P2_IR_REG_7__SCAN_IN, P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN,
         P2_IR_REG_10__SCAN_IN, P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN,
         P2_IR_REG_13__SCAN_IN, P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN,
         P2_IR_REG_16__SCAN_IN, P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN,
         P2_IR_REG_19__SCAN_IN, P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN,
         P2_IR_REG_22__SCAN_IN, P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN,
         P2_IR_REG_25__SCAN_IN, P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN,
         P2_IR_REG_28__SCAN_IN, P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN,
         P2_IR_REG_31__SCAN_IN, P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN,
         P2_D_REG_2__SCAN_IN, P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN,
         P2_D_REG_5__SCAN_IN, P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN,
         P2_D_REG_8__SCAN_IN, P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN,
         P2_D_REG_11__SCAN_IN, P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN,
         P2_D_REG_14__SCAN_IN, P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN,
         P2_D_REG_17__SCAN_IN, P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN,
         P2_D_REG_20__SCAN_IN, P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN,
         P2_D_REG_23__SCAN_IN, P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN,
         P2_D_REG_26__SCAN_IN, P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN,
         P2_D_REG_29__SCAN_IN, P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN,
         P2_REG0_REG_0__SCAN_IN, P2_REG0_REG_1__SCAN_IN,
         P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN,
         P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN,
         P2_REG0_REG_6__SCAN_IN, P2_REG0_REG_7__SCAN_IN,
         P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN,
         P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN,
         P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN,
         P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN,
         P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN,
         P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN,
         P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN,
         P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN,
         P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN,
         P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN,
         P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN,
         P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN,
         P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN,
         P2_REG1_REG_2__SCAN_IN, P2_REG1_REG_3__SCAN_IN,
         P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN,
         P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN,
         P2_REG1_REG_8__SCAN_IN, P2_REG1_REG_9__SCAN_IN,
         P2_REG1_REG_10__SCAN_IN, P2_REG1_REG_11__SCAN_IN,
         P2_REG1_REG_12__SCAN_IN, P2_REG1_REG_13__SCAN_IN,
         P2_REG1_REG_14__SCAN_IN, P2_REG1_REG_15__SCAN_IN,
         P2_REG1_REG_16__SCAN_IN, P2_REG1_REG_17__SCAN_IN,
         P2_REG1_REG_18__SCAN_IN, P2_REG1_REG_19__SCAN_IN,
         P2_REG1_REG_20__SCAN_IN, P2_REG1_REG_21__SCAN_IN,
         P2_REG1_REG_22__SCAN_IN, P2_REG1_REG_23__SCAN_IN,
         P2_REG1_REG_24__SCAN_IN, P2_REG1_REG_25__SCAN_IN,
         P2_REG1_REG_26__SCAN_IN, P2_REG1_REG_27__SCAN_IN,
         P2_REG1_REG_28__SCAN_IN, P2_REG1_REG_29__SCAN_IN,
         P2_REG1_REG_30__SCAN_IN, P2_REG1_REG_31__SCAN_IN,
         P2_REG2_REG_0__SCAN_IN, P2_REG2_REG_1__SCAN_IN,
         P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN,
         P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN,
         P2_REG2_REG_6__SCAN_IN, P2_REG2_REG_7__SCAN_IN,
         P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN,
         P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN,
         P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN,
         P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN,
         P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN,
         P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN,
         P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN,
         P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN,
         P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN,
         P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN,
         P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN,
         P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN,
         P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN,
         P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN,
         P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN,
         P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN,
         P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN,
         P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN,
         P2_ADDR_REG_7__SCAN_IN, P2_ADDR_REG_6__SCAN_IN,
         P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN,
         P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN,
         P2_ADDR_REG_1__SCAN_IN, P2_ADDR_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN;
  output ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58,
         ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63,
         ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51,
         ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46,
         U126, U123, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351,
         P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344,
         P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337,
         P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330,
         P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439,
         P1_U3440, P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318,
         P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311,
         P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304,
         P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297,
         P1_U3296, P1_U3295, P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462,
         P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483,
         P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504,
         P1_U3507, P1_U3509, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291,
         P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284,
         P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277,
         P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270,
         P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264,
         P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257,
         P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250,
         P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243,
         P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240,
         P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233,
         P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226,
         P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219,
         P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086,
         P1_U3085, P1_U3973, P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291,
         P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284,
         P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277,
         P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270,
         P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376,
         P2_U3377, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258,
         P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251,
         P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244,
         P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237,
         P2_U3236, P2_U3235, P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399,
         P2_U3402, P2_U3405, P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420,
         P2_U3423, P2_U3426, P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441,
         P2_U3444, P2_U3446, P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451,
         P2_U3452, P2_U3453, P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458,
         P2_U3459, P2_U3460, P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465,
         P2_U3466, P2_U3467, P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472,
         P2_U3473, P2_U3474, P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479,
         P2_U3480, P2_U3481, P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486,
         P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231,
         P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224,
         P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217,
         P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210,
         P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203,
         P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196,
         P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189,
         P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182,
         P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497,
         P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504,
         P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511,
         P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518,
         P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180,
         P2_U3179, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173,
         P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166,
         P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159,
         P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151,
         P2_U3150, P2_U3893;
  wire   n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139,
         n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149,
         n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159,
         n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169,
         n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179,
         n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189,
         n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199,
         n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209,
         n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219,
         n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229,
         n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239,
         n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249,
         n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259,
         n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269,
         n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279,
         n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289,
         n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299,
         n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309,
         n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319,
         n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329,
         n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339,
         n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349,
         n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359,
         n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369,
         n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379,
         n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389,
         n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399,
         n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409,
         n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419,
         n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429,
         n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439,
         n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449,
         n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459,
         n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469,
         n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479,
         n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489,
         n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499,
         n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509,
         n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519,
         n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529,
         n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539,
         n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549,
         n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559,
         n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569,
         n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579,
         n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589,
         n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599,
         n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609,
         n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619,
         n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629,
         n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639,
         n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649,
         n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659,
         n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669,
         n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679,
         n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689,
         n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699,
         n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709,
         n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719,
         n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729,
         n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739,
         n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749,
         n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759,
         n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769,
         n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779,
         n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789,
         n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799,
         n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809,
         n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819,
         n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829,
         n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839,
         n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849,
         n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859,
         n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869,
         n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879,
         n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889,
         n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899,
         n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909,
         n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919,
         n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929,
         n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939,
         n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949,
         n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959,
         n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969,
         n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979,
         n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989,
         n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999,
         n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009,
         n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019,
         n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029,
         n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039,
         n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049,
         n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059,
         n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069,
         n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079,
         n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089,
         n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099,
         n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109,
         n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119,
         n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129,
         n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139,
         n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149,
         n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159,
         n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169,
         n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179,
         n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189,
         n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199,
         n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209,
         n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219,
         n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229,
         n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239,
         n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249,
         n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259,
         n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269,
         n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279,
         n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289,
         n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299,
         n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309,
         n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319,
         n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329,
         n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339,
         n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349,
         n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359,
         n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369,
         n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379,
         n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389,
         n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399,
         n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409,
         n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419,
         n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429,
         n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439,
         n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449,
         n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459,
         n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469,
         n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479,
         n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489,
         n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499,
         n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509,
         n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519,
         n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529,
         n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539,
         n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549,
         n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559,
         n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569,
         n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579,
         n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589,
         n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599,
         n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609,
         n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619,
         n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629,
         n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639,
         n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649,
         n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659,
         n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669,
         n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679,
         n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689,
         n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699,
         n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709,
         n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719,
         n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729,
         n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739,
         n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749,
         n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759,
         n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769,
         n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779,
         n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789,
         n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799,
         n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809,
         n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819,
         n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829,
         n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839,
         n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849,
         n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859,
         n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869,
         n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879,
         n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889,
         n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899,
         n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909,
         n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919,
         n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929,
         n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939,
         n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949,
         n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959,
         n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969,
         n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979,
         n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989,
         n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999,
         n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009,
         n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019,
         n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029,
         n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039,
         n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049,
         n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059,
         n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069,
         n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079,
         n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089,
         n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099,
         n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109,
         n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119,
         n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129,
         n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139,
         n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149,
         n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159,
         n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169,
         n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179,
         n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189,
         n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199,
         n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209,
         n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219,
         n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229,
         n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239,
         n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249,
         n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259,
         n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269,
         n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279,
         n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289,
         n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299,
         n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309,
         n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319,
         n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329,
         n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339,
         n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349,
         n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359,
         n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369,
         n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379,
         n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389,
         n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399,
         n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409,
         n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419,
         n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429,
         n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439,
         n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449,
         n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459,
         n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469,
         n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479,
         n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489,
         n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499,
         n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509,
         n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519,
         n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529,
         n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539,
         n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549,
         n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559,
         n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569,
         n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579,
         n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589,
         n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599,
         n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609,
         n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619,
         n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629,
         n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639,
         n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649,
         n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659,
         n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669,
         n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679,
         n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689,
         n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699,
         n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709,
         n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719,
         n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729,
         n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739,
         n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749,
         n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759,
         n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769,
         n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779,
         n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789,
         n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799,
         n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809,
         n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819,
         n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829,
         n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839,
         n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849,
         n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859,
         n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869,
         n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879,
         n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889,
         n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899,
         n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909,
         n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919,
         n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929,
         n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939,
         n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949,
         n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959,
         n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969,
         n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979,
         n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989,
         n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999,
         n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009,
         n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019,
         n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029,
         n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039,
         n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049,
         n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059,
         n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069,
         n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079,
         n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089,
         n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099,
         n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109,
         n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119,
         n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129,
         n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139,
         n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149,
         n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159,
         n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169,
         n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179,
         n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189,
         n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199,
         n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209,
         n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219,
         n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229,
         n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239,
         n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249,
         n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259,
         n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269,
         n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279,
         n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289,
         n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299,
         n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309,
         n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319,
         n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329,
         n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339,
         n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349,
         n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359,
         n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369,
         n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379,
         n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389,
         n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399,
         n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409,
         n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419,
         n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429,
         n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439,
         n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449,
         n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459,
         n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469,
         n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479,
         n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489,
         n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499,
         n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509,
         n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519,
         n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529,
         n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539,
         n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549,
         n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559,
         n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569,
         n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579,
         n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589,
         n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599,
         n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609,
         n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619,
         n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629,
         n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639,
         n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649,
         n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659,
         n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669,
         n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679,
         n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689,
         n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699,
         n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709,
         n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719,
         n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729,
         n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739,
         n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749,
         n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759,
         n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769,
         n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779,
         n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789,
         n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799,
         n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809,
         n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819,
         n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829,
         n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839,
         n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849,
         n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859,
         n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869,
         n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879,
         n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889,
         n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899,
         n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909,
         n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919,
         n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929,
         n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939,
         n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949,
         n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959,
         n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969,
         n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979,
         n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989,
         n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999,
         n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009,
         n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019,
         n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029,
         n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039,
         n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049,
         n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059,
         n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069,
         n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079,
         n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089,
         n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099,
         n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109,
         n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119,
         n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129,
         n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139,
         n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149,
         n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159,
         n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169,
         n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179,
         n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189,
         n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199,
         n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209,
         n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219,
         n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229,
         n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239,
         n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249,
         n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259,
         n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269,
         n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279,
         n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289,
         n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299,
         n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309,
         n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319,
         n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329,
         n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339,
         n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349,
         n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359,
         n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369,
         n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379,
         n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389,
         n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399,
         n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409,
         n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419,
         n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429,
         n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439,
         n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449,
         n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459,
         n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469,
         n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479,
         n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489,
         n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499,
         n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509,
         n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519,
         n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529,
         n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539,
         n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549,
         n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559,
         n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569,
         n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579,
         n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589,
         n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599,
         n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609,
         n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619,
         n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629,
         n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639,
         n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649,
         n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659,
         n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669,
         n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679,
         n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689,
         n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699,
         n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709,
         n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719,
         n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729,
         n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739,
         n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749,
         n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759,
         n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769,
         n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779,
         n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789,
         n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799,
         n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809,
         n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819,
         n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829,
         n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839,
         n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849,
         n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859,
         n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869,
         n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879,
         n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889,
         n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899,
         n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909,
         n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919,
         n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929,
         n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939,
         n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949,
         n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959,
         n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969,
         n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979,
         n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989,
         n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999,
         n10000, n10001, n10002, n10003, n10004, n10005, n10006, n10007,
         n10008, n10009, n10010, n10011, n10012, n10013, n10014, n10015,
         n10016, n10017, n10018, n10019, n10020, n10021, n10022, n10023,
         n10024, n10025, n10026, n10027, n10028, n10029, n10030, n10031,
         n10032, n10033, n10034, n10035, n10036, n10037, n10038, n10039,
         n10040, n10041, n10042, n10043, n10044, n10045, n10046, n10047,
         n10048, n10049, n10050, n10051, n10052, n10053, n10054, n10055,
         n10056, n10057, n10058, n10059, n10060, n10061, n10062, n10063,
         n10064, n10065, n10066, n10067, n10068, n10069, n10070, n10071,
         n10072, n10073, n10074, n10075, n10076, n10077, n10078, n10079,
         n10080, n10081, n10082, n10083, n10084, n10085, n10086, n10087,
         n10088, n10089, n10090, n10091, n10092, n10093, n10094, n10095,
         n10096, n10097, n10098, n10099, n10100, n10101, n10102, n10103,
         n10104, n10105, n10106, n10107, n10108, n10109, n10110, n10111,
         n10112, n10113, n10114, n10115, n10116, n10117, n10118, n10119,
         n10120, n10121, n10122, n10123, n10124, n10125, n10126, n10127,
         n10128, n10129, n10130, n10131, n10132, n10133, n10134, n10135,
         n10136, n10137, n10138, n10139, n10140, n10141, n10142, n10143,
         n10144, n10145, n10146, n10147, n10148, n10149, n10150, n10151,
         n10152, n10153, n10154, n10155, n10156, n10157, n10158, n10159,
         n10160, n10161, n10162, n10163, n10164, n10165, n10166, n10167,
         n10168, n10169, n10170, n10171, n10172, n10173, n10174, n10175,
         n10176, n10177, n10178, n10179, n10180, n10181, n10182, n10183,
         n10184, n10185, n10186, n10187, n10188, n10189, n10190, n10191,
         n10192, n10193, n10194, n10195, n10196, n10197, n10198, n10199,
         n10200, n10201, n10202, n10203, n10204, n10205, n10206, n10207,
         n10208, n10209, n10210, n10211, n10212, n10213, n10214, n10215,
         n10216, n10217, n10218, n10219, n10220, n10221, n10222, n10223,
         n10224, n10225, n10226, n10227, n10228, n10229, n10230, n10231,
         n10232, n10233, n10234, n10235, n10236, n10237, n10238, n10239,
         n10240, n10241, n10242, n10243, n10244, n10245, n10246, n10247,
         n10248, n10249, n10250, n10251, n10252, n10253, n10254, n10255,
         n10256, n10257, n10258, n10259, n10260, n10261, n10262, n10263,
         n10264, n10265, n10266, n10267, n10268, n10269, n10270, n10271,
         n10272, n10273, n10274, n10275, n10276, n10277, n10278, n10279,
         n10280, n10281, n10282, n10283, n10284, n10285, n10286, n10287,
         n10288, n10289, n10290, n10291, n10292, n10293, n10294, n10295,
         n10296, n10297, n10298, n10299, n10300, n10301, n10302, n10303,
         n10304, n10305, n10306, n10307, n10308, n10309, n10310, n10311,
         n10312, n10313, n10314, n10315, n10316, n10317, n10318, n10319,
         n10320, n10321, n10322, n10323, n10324, n10325, n10326, n10327,
         n10328, n10329, n10330, n10331, n10332, n10333, n10334, n10335,
         n10336, n10337, n10338, n10339, n10340, n10341, n10342, n10343,
         n10344, n10345, n10346, n10347, n10348, n10349, n10350, n10351,
         n10352, n10353, n10354, n10355, n10356, n10357, n10358, n10359,
         n10360, n10361, n10362, n10363, n10364, n10365, n10366, n10367,
         n10368, n10369, n10370, n10371, n10372, n10373, n10374, n10375,
         n10376, n10377, n10378, n10379, n10380, n10381, n10382, n10383,
         n10384, n10385, n10386, n10387, n10388, n10389, n10390, n10391,
         n10392, n10393, n10394, n10395, n10396, n10397, n10398, n10399,
         n10400, n10401, n10402, n10403, n10404, n10405, n10406, n10407,
         n10408, n10409, n10410, n10411, n10412, n10413, n10414, n10415,
         n10416, n10417, n10418, n10419, n10420, n10421, n10422, n10423,
         n10424, n10425, n10426, n10427, n10428, n10429, n10430, n10431,
         n10432, n10433, n10434, n10435, n10436, n10437, n10438, n10439,
         n10440, n10441, n10442, n10443, n10444, n10445, n10446, n10447,
         n10448, n10449, n10450, n10451, n10452, n10453, n10454, n10455,
         n10456, n10457, n10458, n10459, n10460, n10461, n10462, n10463,
         n10464, n10465, n10466, n10467, n10468, n10469, n10470, n10471,
         n10472, n10473, n10474, n10475, n10476, n10477, n10478, n10479,
         n10480, n10481, n10482, n10483, n10484, n10485, n10486, n10487,
         n10488, n10489, n10490, n10491, n10492, n10493, n10494, n10495,
         n10496, n10497, n10498, n10499, n10500, n10501, n10502, n10503,
         n10504, n10505, n10506, n10507, n10508, n10509, n10510, n10511,
         n10512, n10513, n10514, n10515, n10516, n10517, n10518, n10519,
         n10520, n10521, n10522, n10523, n10524, n10525, n10526, n10527,
         n10528, n10529, n10530, n10531, n10532, n10533, n10534, n10535,
         n10536, n10537, n10538, n10539, n10540, n10541, n10542, n10543,
         n10544, n10545, n10546, n10547, n10548, n10549, n10550, n10551,
         n10552, n10553, n10554, n10555, n10556, n10557, n10558, n10559,
         n10560, n10561, n10562, n10563, n10564, n10565, n10566, n10567,
         n10568, n10569, n10570, n10571, n10572, n10573, n10574, n10575,
         n10576, n10577, n10578, n10579, n10580, n10581, n10582, n10583,
         n10584, n10585, n10586, n10587, n10588, n10589, n10590, n10591,
         n10592, n10593, n10594, n10595, n10596, n10597, n10598, n10599,
         n10600, n10601, n10602, n10603, n10604, n10605, n10606, n10607,
         n10608, n10609, n10610, n10611, n10612, n10613, n10614, n10615,
         n10616, n10617, n10618, n10619, n10620, n10621, n10622, n10623,
         n10624, n10625, n10626, n10627, n10628, n10629, n10630, n10631,
         n10632, n10633, n10634, n10635, n10636, n10637, n10638, n10639,
         n10640, n10641, n10642, n10643, n10644, n10645, n10646, n10647,
         n10648, n10649, n10650, n10651, n10652, n10653, n10654, n10655,
         n10656, n10657, n10658, n10659, n10660, n10661, n10662, n10663,
         n10664, n10665, n10666, n10667, n10668, n10669, n10670, n10671,
         n10672, n10673, n10674, n10675, n10676, n10677, n10678, n10679,
         n10680, n10681, n10682, n10683, n10684, n10685, n10686, n10687,
         n10688, n10689, n10690, n10691, n10692, n10693, n10694, n10695,
         n10696, n10697, n10698, n10699, n10700, n10701, n10702, n10703,
         n10704, n10705, n10706, n10707, n10708, n10709, n10710, n10711,
         n10712, n10713, n10714, n10715, n10716, n10717, n10718, n10719,
         n10720, n10721, n10722, n10723, n10724, n10725, n10726, n10727,
         n10728, n10729, n10730, n10731, n10732, n10733, n10734, n10735,
         n10736, n10737, n10738, n10739, n10740, n10741, n10742, n10743,
         n10744, n10745, n10746, n10747, n10748, n10749, n10750, n10751,
         n10752, n10753, n10754, n10755, n10756, n10757, n10758, n10759,
         n10760, n10761, n10762, n10763, n10764, n10765, n10766, n10767,
         n10768, n10769, n10770, n10771, n10772, n10773, n10774, n10775,
         n10776, n10777, n10778, n10779, n10780, n10781, n10782, n10783,
         n10784, n10785, n10786, n10787, n10788, n10789, n10790, n10791,
         n10792, n10793, n10794, n10795, n10796, n10797, n10798, n10799,
         n10800, n10801, n10802, n10803, n10804, n10805, n10806, n10807,
         n10808, n10809, n10810, n10811, n10812, n10813, n10814, n10815,
         n10816, n10817, n10818, n10819, n10820, n10821, n10822, n10823,
         n10824, n10825, n10826, n10827, n10828, n10829, n10830, n10831,
         n10832, n10833, n10834, n10835, n10836, n10837, n10838, n10839,
         n10840, n10841, n10842, n10843, n10844, n10845, n10846, n10847,
         n10848, n10849, n10850, n10851, n10852, n10853, n10854, n10855,
         n10856, n10857, n10858, n10859, n10860, n10861, n10862, n10863,
         n10864, n10865, n10866, n10867, n10868, n10869, n10870, n10871,
         n10872, n10873, n10874, n10875, n10876, n10877, n10878, n10879,
         n10880, n10881, n10882, n10883, n10884, n10885, n10886, n10887,
         n10888, n10889, n10890, n10891, n10892, n10893, n10894, n10895,
         n10896, n10897, n10898, n10899, n10900, n10901, n10902, n10903,
         n10904, n10905, n10906, n10907, n10908, n10909, n10910, n10911,
         n10912, n10913, n10914, n10915, n10916, n10917, n10918, n10919,
         n10920, n10921, n10922, n10923, n10924, n10925, n10926, n10927,
         n10928, n10929, n10930, n10931, n10932, n10933, n10934, n10935,
         n10936, n10937, n10938, n10939, n10940, n10941, n10942, n10943,
         n10944, n10945, n10946, n10947, n10948, n10949, n10950, n10951,
         n10952, n10953, n10954, n10955, n10956, n10957, n10958, n10959,
         n10960, n10961, n10962, n10963, n10964, n10965, n10966, n10967,
         n10968, n10969, n10970, n10971, n10972, n10973, n10974, n10975,
         n10976, n10977, n10978, n10979, n10980, n10981, n10982, n10983,
         n10984, n10985, n10986, n10987, n10988, n10989, n10990, n10991,
         n10992, n10993, n10994, n10995, n10996, n10997, n10998, n10999,
         n11000, n11001, n11002, n11003, n11004, n11005, n11006, n11007,
         n11008, n11009, n11010, n11011, n11012, n11013, n11014, n11015,
         n11016, n11017, n11018, n11019, n11020, n11021, n11022, n11023,
         n11024, n11025, n11026, n11027, n11028, n11029, n11030, n11031,
         n11032, n11033, n11034, n11035, n11036, n11037, n11038, n11039,
         n11040, n11041, n11042, n11043, n11044, n11045, n11046, n11047,
         n11048, n11049, n11050, n11051, n11052, n11053, n11054, n11055,
         n11056, n11057, n11058, n11059, n11060, n11061, n11062, n11063,
         n11064, n11065, n11066, n11067, n11068, n11069, n11070, n11071,
         n11072, n11073, n11074, n11075, n11076, n11077, n11078, n11079,
         n11080, n11081, n11082, n11083, n11084, n11085, n11086, n11087,
         n11088, n11089, n11090, n11091, n11092, n11093, n11094, n11095,
         n11096, n11097, n11098, n11099, n11100, n11101, n11102, n11103,
         n11104, n11105, n11106, n11107, n11108, n11109, n11110, n11111,
         n11112, n11113, n11114, n11115, n11116, n11117, n11118, n11119,
         n11120, n11121, n11122, n11123, n11124, n11125, n11126, n11127,
         n11128, n11129, n11130, n11131, n11132, n11133, n11134, n11135,
         n11136, n11137, n11138, n11139, n11140, n11141, n11142, n11143,
         n11144, n11145, n11146, n11147, n11148, n11149, n11150, n11151,
         n11152, n11153, n11154, n11155, n11156, n11157, n11158, n11159,
         n11160, n11161, n11162, n11163, n11164, n11165, n11166, n11167,
         n11168, n11169, n11170, n11171, n11172, n11173, n11174, n11175,
         n11176, n11177, n11178;

  OR2_X1 U5194 ( .A1(n8351), .A2(n10649), .ZN(n5310) );
  OR2_X1 U5195 ( .A1(n10483), .A2(n10482), .ZN(n10486) );
  INV_X1 U5196 ( .A(n6646), .ZN(n8317) );
  INV_X1 U5197 ( .A(n8809), .ZN(n8781) );
  CLKBUF_X2 U5198 ( .A(n5755), .Z(n5598) );
  AND2_X1 U5199 ( .A1(n6455), .A2(n6454), .ZN(n6782) );
  INV_X2 U5200 ( .A(n6824), .ZN(n6520) );
  INV_X1 U5201 ( .A(n5864), .ZN(n5755) );
  NAND2_X1 U5202 ( .A1(n8094), .A2(n8093), .ZN(n8151) );
  NAND2_X1 U5203 ( .A1(n8806), .A2(n8809), .ZN(n7344) );
  INV_X1 U5204 ( .A(n5134), .ZN(n5135) );
  OR2_X1 U5205 ( .A1(n5869), .A2(n5868), .ZN(n5377) );
  INV_X1 U5206 ( .A(n5131), .ZN(n5132) );
  OR2_X1 U5207 ( .A1(n6886), .A2(n8819), .ZN(n6887) );
  NAND2_X1 U5208 ( .A1(n6474), .A2(n5755), .ZN(n6699) );
  NAND2_X1 U5209 ( .A1(n8624), .A2(n9327), .ZN(n6895) );
  NOR2_X1 U5210 ( .A1(n6886), .A2(n5432), .ZN(n9073) );
  OAI21_X1 U5211 ( .B1(n10507), .B2(n5508), .A(n5181), .ZN(n10476) );
  INV_X1 U5212 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n10692) );
  BUF_X1 U5213 ( .A(n9378), .Z(n5137) );
  AND4_X1 U5214 ( .A1(n5856), .A2(n5855), .A3(n5854), .A4(n5853), .ZN(n5130)
         );
  INV_X1 U5215 ( .A(n6729), .ZN(n5131) );
  XNOR2_X2 U5216 ( .A(n8077), .B(n8078), .ZN(n7990) );
  AOI22_X2 U5217 ( .A1(P2_REG2_REG_12__SCAN_IN), .A2(n8153), .B1(n8152), .B2(
        n8151), .ZN(n8269) );
  OAI21_X2 U5218 ( .B1(n7702), .B2(n5304), .A(n5173), .ZN(n7915) );
  XNOR2_X2 U5219 ( .A(n8257), .B(n8270), .ZN(n8145) );
  NAND2_X2 U5220 ( .A1(n6380), .A2(n8592), .ZN(n9415) );
  INV_X2 U5221 ( .A(n5131), .ZN(n5133) );
  AND2_X1 U5222 ( .A1(n9080), .A2(n10700), .ZN(n6729) );
  NAND2_X2 U5223 ( .A1(n9612), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5867) );
  OAI21_X2 U5224 ( .B1(n7394), .B2(n8509), .A(n8512), .ZN(n7474) );
  NAND2_X2 U5225 ( .A1(n7283), .A2(n8511), .ZN(n7394) );
  INV_X1 U5226 ( .A(n5956), .ZN(n5134) );
  NAND2_X1 U5227 ( .A1(n5872), .A2(n5871), .ZN(n5956) );
  AOI21_X2 U5228 ( .B1(P2_REG2_REG_16__SCAN_IN), .B2(n9336), .A(n9335), .ZN(
        n9337) );
  NOR2_X2 U5229 ( .A1(n8144), .A2(n8143), .ZN(n8257) );
  NAND2_X1 U5231 ( .A1(n5282), .A2(n5211), .ZN(n10227) );
  INV_X1 U5232 ( .A(n8806), .ZN(n8692) );
  INV_X4 U5233 ( .A(n5152), .ZN(n5136) );
  INV_X1 U5234 ( .A(n8618), .ZN(n8588) );
  CLKBUF_X2 U5235 ( .A(n7053), .Z(n8375) );
  NAND2_X1 U5236 ( .A1(n5310), .A2(n5309), .ZN(n6889) );
  AND2_X1 U5237 ( .A1(n8342), .A2(n6828), .ZN(n6829) );
  AOI21_X1 U5238 ( .B1(n5548), .B2(n5552), .A(n5546), .ZN(n5545) );
  AND2_X1 U5239 ( .A1(n5557), .A2(n5549), .ZN(n5548) );
  NAND2_X1 U5240 ( .A1(n5256), .A2(n9097), .ZN(n9110) );
  NAND2_X1 U5241 ( .A1(n10524), .A2(n10523), .ZN(n10522) );
  NAND2_X1 U5242 ( .A1(n10494), .A2(n10495), .ZN(n10493) );
  NAND2_X1 U5243 ( .A1(n5283), .A2(n5717), .ZN(n10185) );
  OAI21_X1 U5244 ( .B1(n9489), .B2(n6220), .A(n6219), .ZN(n9472) );
  NAND2_X1 U5245 ( .A1(n5574), .A2(n5214), .ZN(n5573) );
  AND3_X1 U5246 ( .A1(n5481), .A2(n5480), .A3(n5218), .ZN(n9297) );
  NAND2_X1 U5247 ( .A1(n5279), .A2(n8643), .ZN(n10091) );
  NAND2_X1 U5248 ( .A1(n10090), .A2(n10093), .ZN(n5701) );
  NAND2_X1 U5249 ( .A1(n11131), .A2(n5311), .ZN(n8065) );
  INV_X1 U5250 ( .A(n6357), .ZN(n5465) );
  OR2_X1 U5251 ( .A1(n8154), .A2(n5483), .ZN(n5480) );
  OAI21_X1 U5252 ( .B1(n8145), .B2(n5594), .A(n5593), .ZN(n9261) );
  OR2_X1 U5253 ( .A1(n11152), .A2(n11124), .ZN(n11127) );
  NAND2_X1 U5254 ( .A1(n7371), .A2(n7370), .ZN(n7493) );
  NAND2_X1 U5255 ( .A1(n7812), .A2(n6804), .ZN(n7414) );
  OR2_X1 U5256 ( .A1(n7810), .A2(n6803), .ZN(n7812) );
  NOR2_X1 U5257 ( .A1(n7749), .A2(n7748), .ZN(n7750) );
  OR2_X1 U5258 ( .A1(n7320), .A2(n5263), .ZN(n5262) );
  NAND2_X1 U5259 ( .A1(n9284), .A2(n5214), .ZN(n5572) );
  INV_X1 U5260 ( .A(n8501), .ZN(n8446) );
  NAND2_X4 U5261 ( .A1(n5265), .A2(n6898), .ZN(n6905) );
  NOR2_X1 U5262 ( .A1(n10923), .A2(n7262), .ZN(n10922) );
  INV_X2 U5263 ( .A(n6960), .ZN(n6991) );
  NAND4_X1 U5264 ( .A1(n6471), .A2(n6470), .A3(n6469), .A4(n6468), .ZN(n10297)
         );
  NAND2_X2 U5265 ( .A1(n5275), .A2(n7333), .ZN(n8809) );
  NAND4_X2 U5266 ( .A1(n6459), .A2(n6458), .A3(n6457), .A4(n6456), .ZN(n11000)
         );
  INV_X1 U5267 ( .A(n5951), .ZN(n6330) );
  INV_X1 U5268 ( .A(n7110), .ZN(n6812) );
  NAND2_X2 U5269 ( .A1(n6897), .A2(n8630), .ZN(n8618) );
  XNOR2_X1 U5270 ( .A(n6397), .B(n6396), .ZN(n8135) );
  NAND2_X1 U5271 ( .A1(n6394), .A2(n6395), .ZN(n6406) );
  XNOR2_X1 U5272 ( .A(n6339), .B(n6338), .ZN(n6896) );
  NAND2_X1 U5273 ( .A1(n6834), .A2(n6839), .ZN(n8164) );
  NAND2_X1 U5274 ( .A1(n6395), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6397) );
  INV_X2 U5275 ( .A(n9328), .ZN(n9324) );
  MUX2_X1 U5276 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6832), .S(
        P1_IR_REG_25__SCAN_IN), .Z(n6834) );
  NOR2_X1 U5277 ( .A1(n6102), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n6118) );
  XNOR2_X1 U5278 ( .A(n5377), .B(P2_IR_REG_29__SCAN_IN), .ZN(n5871) );
  NAND2_X1 U5279 ( .A1(n5618), .A2(n5617), .ZN(n6339) );
  OR2_X1 U5280 ( .A1(n6833), .A2(n10692), .ZN(n6832) );
  NAND2_X1 U5281 ( .A1(n10693), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6450) );
  NAND2_X1 U5282 ( .A1(n6474), .A2(n8306), .ZN(n6646) );
  INV_X1 U5283 ( .A(n6643), .ZN(n6644) );
  XNOR2_X1 U5284 ( .A(n5965), .B(n5964), .ZN(n7053) );
  NOR2_X1 U5285 ( .A1(n5857), .A2(n5421), .ZN(n5420) );
  NOR2_X1 U5286 ( .A1(n5624), .A2(n5622), .ZN(n6047) );
  CLKBUF_X1 U5287 ( .A(n5864), .Z(n8306) );
  INV_X1 U5288 ( .A(n6031), .ZN(n5526) );
  NAND4_X1 U5289 ( .A1(n5847), .A2(n5438), .A3(n5848), .A4(n5849), .ZN(n6031)
         );
  NAND3_X1 U5290 ( .A1(n5274), .A2(n6465), .A3(n6439), .ZN(n6513) );
  AND2_X2 U5291 ( .A1(n5944), .A2(n5439), .ZN(n5438) );
  AND2_X1 U5292 ( .A1(n9764), .A2(n9974), .ZN(n5274) );
  INV_X1 U5293 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n10013) );
  NOR2_X1 U5294 ( .A1(P1_IR_REG_21__SCAN_IN), .A2(P1_IR_REG_20__SCAN_IN), .ZN(
        n6789) );
  NOR2_X1 U5295 ( .A1(P2_IR_REG_17__SCAN_IN), .A2(P2_IR_REG_21__SCAN_IN), .ZN(
        n5853) );
  NOR2_X1 U5296 ( .A1(P2_IR_REG_18__SCAN_IN), .A2(P2_IR_REG_9__SCAN_IN), .ZN(
        n5854) );
  NOR2_X1 U5297 ( .A1(P2_IR_REG_12__SCAN_IN), .A2(P2_IR_REG_19__SCAN_IN), .ZN(
        n5855) );
  INV_X1 U5298 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n9787) );
  INV_X1 U5299 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n9995) );
  NOR2_X1 U5300 ( .A1(P2_IR_REG_3__SCAN_IN), .A2(P2_IR_REG_2__SCAN_IN), .ZN(
        n5848) );
  INV_X1 U5301 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n6206) );
  NOR2_X2 U5302 ( .A1(n10626), .A2(n10554), .ZN(n10535) );
  AOI211_X2 U5303 ( .C1(n8334), .C2(n6887), .A(n10577), .B(n9073), .ZN(n8339)
         );
  NOR2_X1 U5304 ( .A1(n8438), .A2(n5558), .ZN(n5557) );
  NOR2_X1 U5305 ( .A1(n9346), .A2(n9578), .ZN(n5558) );
  OAI21_X1 U5306 ( .B1(n6946), .B2(P2_D_REG_0__SCAN_IN), .A(n6407), .ZN(n6408)
         );
  AND2_X1 U5307 ( .A1(n6047), .A2(n6046), .ZN(n6050) );
  INV_X1 U5308 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n6046) );
  OR2_X1 U5309 ( .A1(n10450), .A2(n10462), .ZN(n9039) );
  NOR2_X1 U5310 ( .A1(n5703), .A2(n6443), .ZN(n5702) );
  NAND2_X1 U5311 ( .A1(n9781), .A2(n9780), .ZN(n5703) );
  AOI21_X1 U5312 ( .B1(n5687), .B2(n5689), .A(n5208), .ZN(n5686) );
  INV_X1 U5313 ( .A(n6149), .ZN(n5687) );
  INV_X1 U5314 ( .A(n5468), .ZN(n9361) );
  OAI21_X1 U5315 ( .B1(n9376), .B2(n5470), .A(n5469), .ZN(n5468) );
  AND2_X1 U5316 ( .A1(n9099), .A2(n9390), .ZN(n5470) );
  NAND2_X1 U5317 ( .A1(n9362), .A2(n9522), .ZN(n5469) );
  AND2_X1 U5318 ( .A1(n8593), .A2(n6379), .ZN(n5560) );
  NAND2_X1 U5319 ( .A1(n5291), .A2(n5519), .ZN(n10524) );
  AND2_X1 U5320 ( .A1(n5520), .A2(n6698), .ZN(n5519) );
  NAND2_X1 U5321 ( .A1(n8246), .A2(n5518), .ZN(n5291) );
  OR2_X1 U5322 ( .A1(n10626), .A2(n10281), .ZN(n6698) );
  INV_X1 U5323 ( .A(n6699), .ZN(n6546) );
  NAND2_X1 U5324 ( .A1(n8504), .A2(n8503), .ZN(n8514) );
  INV_X1 U5325 ( .A(n8585), .ZN(n5416) );
  OAI21_X1 U5326 ( .B1(n5387), .B2(n5386), .A(n5378), .ZN(n8580) );
  OR2_X1 U5327 ( .A1(n7317), .A2(n6899), .ZN(n8486) );
  NAND2_X1 U5328 ( .A1(n11087), .A2(n10119), .ZN(n5514) );
  AND2_X1 U5329 ( .A1(n9182), .A2(n9088), .ZN(n9093) );
  INV_X1 U5330 ( .A(n8437), .ZN(n5546) );
  OR2_X1 U5331 ( .A1(n8424), .A2(n5553), .ZN(n5552) );
  NAND2_X1 U5332 ( .A1(n8357), .A2(n8356), .ZN(n8358) );
  NOR2_X1 U5333 ( .A1(n6165), .A2(n8483), .ZN(n6372) );
  NAND2_X1 U5334 ( .A1(n7317), .A2(n6899), .ZN(n8489) );
  INV_X1 U5335 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n5849) );
  NOR2_X1 U5336 ( .A1(P2_IR_REG_4__SCAN_IN), .A2(P2_IR_REG_5__SCAN_IN), .ZN(
        n5847) );
  INV_X1 U5337 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n5439) );
  NOR2_X1 U5338 ( .A1(n8778), .A2(n5713), .ZN(n5712) );
  INV_X1 U5339 ( .A(n8765), .ZN(n5713) );
  NOR2_X1 U5340 ( .A1(n8334), .A2(n8819), .ZN(n5434) );
  NAND2_X1 U5341 ( .A1(n10444), .A2(n5139), .ZN(n5605) );
  NAND2_X1 U5342 ( .A1(n10459), .A2(n10458), .ZN(n10441) );
  NAND2_X1 U5343 ( .A1(n10486), .A2(n8980), .ZN(n10459) );
  AND2_X1 U5344 ( .A1(n9030), .A2(n10526), .ZN(n5333) );
  AOI21_X1 U5345 ( .B1(n8951), .B2(n5524), .A(n6690), .ZN(n5523) );
  OR2_X1 U5346 ( .A1(n10267), .A2(n11136), .ZN(n9015) );
  NAND2_X1 U5347 ( .A1(n11129), .A2(n6809), .ZN(n11131) );
  AOI21_X1 U5348 ( .B1(n5660), .B2(n6299), .A(n5217), .ZN(n5658) );
  INV_X1 U5349 ( .A(n5660), .ZN(n5659) );
  NOR2_X1 U5350 ( .A1(n6221), .A2(n5656), .ZN(n5655) );
  INV_X1 U5351 ( .A(n5813), .ZN(n5656) );
  INV_X1 U5352 ( .A(n5666), .ZN(n5665) );
  AOI21_X1 U5353 ( .B1(n5666), .B2(n5668), .A(n5664), .ZN(n5663) );
  INV_X1 U5354 ( .A(n6108), .ZN(n5664) );
  AOI21_X1 U5355 ( .B1(n5677), .B2(n5679), .A(n5182), .ZN(n5676) );
  INV_X1 U5356 ( .A(n6012), .ZN(n5677) );
  NAND2_X1 U5357 ( .A1(n7080), .A2(n5266), .ZN(n5265) );
  AND2_X1 U5358 ( .A1(n6895), .A2(n6896), .ZN(n5266) );
  OAI21_X1 U5359 ( .B1(n5150), .B2(n5633), .A(n5632), .ZN(n5631) );
  AND2_X1 U5360 ( .A1(n9111), .A2(n9101), .ZN(n5633) );
  NAND2_X1 U5361 ( .A1(n5150), .A2(n9101), .ZN(n5632) );
  NAND2_X1 U5362 ( .A1(n5642), .A2(n5641), .ZN(n7772) );
  AND2_X1 U5363 ( .A1(n5142), .A2(n7685), .ZN(n5641) );
  NAND2_X1 U5364 ( .A1(n6913), .A2(n7513), .ZN(n5645) );
  NAND2_X1 U5365 ( .A1(n5258), .A2(n5257), .ZN(n7384) );
  NAND2_X1 U5366 ( .A1(n5262), .A2(n6912), .ZN(n5257) );
  AOI21_X1 U5367 ( .B1(n5260), .B2(n7221), .A(n5259), .ZN(n5258) );
  AND2_X1 U5368 ( .A1(n6912), .A2(n7220), .ZN(n5260) );
  NOR2_X1 U5369 ( .A1(n5612), .A2(n9092), .ZN(n5611) );
  INV_X1 U5370 ( .A(n9152), .ZN(n5612) );
  INV_X1 U5371 ( .A(n6329), .ZN(n8428) );
  NAND2_X1 U5372 ( .A1(n6401), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5863) );
  OR2_X1 U5373 ( .A1(n7425), .A2(n5210), .ZN(n5577) );
  NOR2_X1 U5374 ( .A1(n7429), .A2(n7675), .ZN(n5583) );
  XNOR2_X1 U5375 ( .A(n7750), .B(n7761), .ZN(n7790) );
  NAND2_X1 U5376 ( .A1(n7751), .A2(n7798), .ZN(n5587) );
  NOR2_X1 U5377 ( .A1(n5168), .A2(n5647), .ZN(n5646) );
  INV_X1 U5378 ( .A(n5648), .ZN(n5647) );
  AOI21_X1 U5379 ( .B1(n9401), .B2(n6316), .A(n6315), .ZN(n9387) );
  AOI21_X1 U5380 ( .B1(n6273), .B2(n5453), .A(n5145), .ZN(n5451) );
  NAND2_X1 U5381 ( .A1(n9437), .A2(n6378), .ZN(n5561) );
  NAND2_X1 U5382 ( .A1(n5543), .A2(n5541), .ZN(n9482) );
  AOI21_X1 U5383 ( .B1(n9501), .B2(n8577), .A(n5542), .ZN(n5541) );
  NOR2_X1 U5384 ( .A1(n6372), .A2(n5531), .ZN(n5530) );
  INV_X1 U5385 ( .A(n9476), .ZN(n9495) );
  INV_X1 U5386 ( .A(n9474), .ZN(n9492) );
  INV_X1 U5387 ( .A(n5966), .ZN(n6224) );
  NAND2_X1 U5388 ( .A1(n6896), .A2(n7975), .ZN(n9565) );
  NAND2_X1 U5389 ( .A1(n6410), .A2(n6409), .ZN(n7082) );
  OR2_X1 U5390 ( .A1(n6946), .A2(P2_D_REG_1__SCAN_IN), .ZN(n6410) );
  OAI21_X1 U5391 ( .B1(n6223), .B2(P2_IR_REG_18__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n6337) );
  XNOR2_X1 U5392 ( .A(n6337), .B(P2_IR_REG_19__SCAN_IN), .ZN(n9327) );
  NAND2_X1 U5393 ( .A1(n6793), .A2(n6791), .ZN(n6842) );
  AND2_X1 U5394 ( .A1(n8684), .A2(n5718), .ZN(n5717) );
  NAND2_X1 U5395 ( .A1(n8675), .A2(n10209), .ZN(n5718) );
  INV_X1 U5396 ( .A(n6782), .ZN(n6773) );
  AOI21_X1 U5397 ( .B1(n5500), .B2(n5496), .A(n5302), .ZN(n5301) );
  INV_X1 U5398 ( .A(n5499), .ZN(n5302) );
  NAND2_X1 U5399 ( .A1(n5493), .A2(n5490), .ZN(n6879) );
  AND2_X1 U5400 ( .A1(n5498), .A2(n5491), .ZN(n5490) );
  OR2_X1 U5401 ( .A1(n10440), .A2(n5494), .ZN(n5493) );
  AND2_X1 U5402 ( .A1(n8957), .A2(n5499), .ZN(n5498) );
  NAND2_X1 U5403 ( .A1(n10440), .A2(n10442), .ZN(n5500) );
  NAND2_X1 U5404 ( .A1(n9039), .A2(n8905), .ZN(n10442) );
  AND2_X1 U5405 ( .A1(n5292), .A2(n5212), .ZN(n8246) );
  NAND2_X1 U5406 ( .A1(n8177), .A2(n8179), .ZN(n5292) );
  INV_X1 U5407 ( .A(n7915), .ZN(n6627) );
  NOR2_X1 U5408 ( .A1(n7729), .A2(n7654), .ZN(n5427) );
  OAI21_X1 U5409 ( .B1(n8928), .B2(n7723), .A(n6475), .ZN(n10994) );
  AND3_X1 U5410 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_28__SCAN_IN), .A3(
        P1_IR_REG_27__SCAN_IN), .ZN(n6464) );
  NAND2_X1 U5411 ( .A1(n6451), .A2(n5735), .ZN(n6463) );
  AND2_X1 U5412 ( .A1(n6814), .A2(n8971), .ZN(n7117) );
  NAND2_X1 U5413 ( .A1(n6750), .A2(n6749), .ZN(n10450) );
  AND2_X1 U5414 ( .A1(n9061), .A2(n6845), .ZN(n10689) );
  AND2_X1 U5415 ( .A1(n7333), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6845) );
  NAND2_X1 U5416 ( .A1(n6681), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6682) );
  OAI21_X1 U5417 ( .B1(n6150), .B2(n5688), .A(n5686), .ZN(n6186) );
  NAND2_X1 U5418 ( .A1(n6013), .A2(n6012), .ZN(n6015) );
  INV_X1 U5419 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n6439) );
  NAND2_X1 U5420 ( .A1(n5461), .A2(n9490), .ZN(n5466) );
  XOR2_X1 U5421 ( .A(n8812), .B(n8811), .Z(n8813) );
  INV_X1 U5422 ( .A(n10269), .ZN(n10244) );
  INV_X1 U5423 ( .A(n8819), .ZN(n8807) );
  NOR2_X1 U5424 ( .A1(n8853), .A2(n5223), .ZN(n5222) );
  OAI21_X1 U5425 ( .B1(n6805), .B2(n8920), .A(n5224), .ZN(n5223) );
  NAND2_X1 U5426 ( .A1(n5225), .A2(n8920), .ZN(n5224) );
  INV_X1 U5427 ( .A(n8935), .ZN(n5225) );
  NAND2_X1 U5428 ( .A1(n5364), .A2(n8588), .ZN(n5363) );
  OAI21_X1 U5429 ( .B1(n8514), .B2(n8513), .A(n5366), .ZN(n5365) );
  NAND2_X1 U5430 ( .A1(n8517), .A2(n8618), .ZN(n5362) );
  NAND2_X1 U5431 ( .A1(n5229), .A2(n5226), .ZN(n8883) );
  NOR2_X1 U5432 ( .A1(n9545), .A2(n8587), .ZN(n5419) );
  AND2_X1 U5433 ( .A1(n5383), .A2(n5382), .ZN(n8575) );
  INV_X1 U5434 ( .A(n8567), .ZN(n5382) );
  NAND2_X1 U5435 ( .A1(n8568), .A2(n8569), .ZN(n5383) );
  NAND2_X1 U5436 ( .A1(n5381), .A2(n9493), .ZN(n5380) );
  NAND2_X1 U5437 ( .A1(n5234), .A2(n8895), .ZN(n5233) );
  NAND2_X1 U5438 ( .A1(n5236), .A2(n5235), .ZN(n5234) );
  AOI21_X1 U5439 ( .B1(n5414), .B2(n5417), .A(n5413), .ZN(n5412) );
  AOI21_X1 U5440 ( .B1(n5408), .B2(n5410), .A(n5407), .ZN(n5406) );
  INV_X1 U5441 ( .A(n8594), .ZN(n5407) );
  NOR2_X1 U5442 ( .A1(n8906), .A2(n10430), .ZN(n5249) );
  NAND2_X1 U5443 ( .A1(n5248), .A2(n8907), .ZN(n5247) );
  NOR2_X1 U5444 ( .A1(n8957), .A2(n5245), .ZN(n5244) );
  INV_X1 U5445 ( .A(n8916), .ZN(n5245) );
  NOR2_X1 U5446 ( .A1(n9051), .A2(n8823), .ZN(n8919) );
  OR2_X1 U5447 ( .A1(n10603), .A2(n10496), .ZN(n8980) );
  INV_X1 U5448 ( .A(SI_9_), .ZN(n9860) );
  INV_X1 U5449 ( .A(P1_RD_REG_SCAN_IN), .ZN(n5288) );
  INV_X1 U5450 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n5290) );
  NAND2_X1 U5451 ( .A1(n5189), .A2(n5403), .ZN(n5402) );
  INV_X1 U5452 ( .A(n8619), .ZN(n5403) );
  NAND2_X1 U5453 ( .A1(n5369), .A2(n5368), .ZN(n5367) );
  INV_X1 U5454 ( .A(n8613), .ZN(n5368) );
  OAI21_X1 U5455 ( .B1(n5374), .B2(n5371), .A(n5370), .ZN(n5369) );
  OR2_X1 U5456 ( .A1(n8375), .A2(n11029), .ZN(n5476) );
  NAND2_X1 U5457 ( .A1(n8375), .A2(n11029), .ZN(n5475) );
  NAND2_X1 U5458 ( .A1(n5570), .A2(n7060), .ZN(n5569) );
  NAND2_X1 U5459 ( .A1(n5569), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n5568) );
  NAND2_X1 U5460 ( .A1(n7055), .A2(n7259), .ZN(n5571) );
  NOR2_X1 U5461 ( .A1(n6252), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n5221) );
  OR2_X1 U5462 ( .A1(n9549), .A2(n9477), .ZN(n8581) );
  INV_X1 U5463 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n9889) );
  NAND2_X1 U5464 ( .A1(n6366), .A2(n6368), .ZN(n6369) );
  NAND2_X1 U5465 ( .A1(n6165), .A2(n6370), .ZN(n8558) );
  NAND2_X1 U5466 ( .A1(n6363), .A2(n5539), .ZN(n5538) );
  INV_X1 U5467 ( .A(n8538), .ZN(n5539) );
  INV_X1 U5468 ( .A(n5538), .ZN(n5534) );
  NAND2_X1 U5469 ( .A1(n5389), .A2(n7223), .ZN(n8511) );
  OR2_X1 U5470 ( .A1(n7478), .A2(n7403), .ZN(n7396) );
  NOR2_X1 U5471 ( .A1(n6148), .A2(n5447), .ZN(n5446) );
  INV_X1 U5472 ( .A(n8560), .ZN(n5445) );
  NAND2_X1 U5473 ( .A1(n5859), .A2(n5565), .ZN(n5564) );
  INV_X1 U5474 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n5565) );
  NOR2_X1 U5475 ( .A1(n5857), .A2(P2_IR_REG_22__SCAN_IN), .ZN(n5525) );
  INV_X1 U5476 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n5964) );
  NAND3_X1 U5477 ( .A1(n5701), .A2(n10091), .A3(n5699), .ZN(n5698) );
  INV_X1 U5478 ( .A(n10165), .ZN(n5699) );
  INV_X1 U5479 ( .A(n8695), .ZN(n5715) );
  OAI21_X1 U5480 ( .B1(n5242), .B2(n5241), .A(n5238), .ZN(n8965) );
  INV_X1 U5481 ( .A(n8925), .ZN(n5241) );
  INV_X1 U5482 ( .A(n8924), .ZN(n5242) );
  INV_X1 U5483 ( .A(n5239), .ZN(n5238) );
  OR2_X1 U5484 ( .A1(n8334), .A2(n8816), .ZN(n8827) );
  NOR2_X1 U5485 ( .A1(n5497), .A2(n5155), .ZN(n5496) );
  NOR2_X1 U5486 ( .A1(n6726), .A2(n5510), .ZN(n5509) );
  INV_X1 U5487 ( .A(n6717), .ZN(n5510) );
  NAND2_X1 U5488 ( .A1(n5507), .A2(n5509), .ZN(n5506) );
  INV_X1 U5489 ( .A(n10513), .ZN(n5507) );
  AND2_X1 U5490 ( .A1(n5426), .A2(n10668), .ZN(n5425) );
  NAND2_X1 U5491 ( .A1(n9031), .A2(n9030), .ZN(n5332) );
  NOR2_X1 U5492 ( .A1(n10613), .A2(n10538), .ZN(n5426) );
  OR2_X1 U5493 ( .A1(n10568), .A2(n10626), .ZN(n10526) );
  OAI21_X1 U5494 ( .B1(n8222), .B2(n5315), .A(n5312), .ZN(n10565) );
  AOI21_X1 U5495 ( .B1(n5314), .B2(n5596), .A(n5313), .ZN(n5312) );
  INV_X1 U5496 ( .A(n5596), .ZN(n5315) );
  INV_X1 U5497 ( .A(n8889), .ZN(n5313) );
  NAND2_X1 U5498 ( .A1(n5435), .A2(n10680), .ZN(n10554) );
  INV_X1 U5499 ( .A(n6579), .ZN(n5306) );
  NAND2_X1 U5500 ( .A1(n5305), .A2(n7696), .ZN(n5303) );
  OR2_X1 U5501 ( .A1(n10101), .A2(n10170), .ZN(n8855) );
  OR2_X1 U5502 ( .A1(n11053), .A2(n10292), .ZN(n8998) );
  INV_X1 U5503 ( .A(n5325), .ZN(n5324) );
  OAI21_X1 U5504 ( .B1(n5139), .B2(n6881), .A(n8957), .ZN(n5325) );
  NAND2_X1 U5505 ( .A1(n5605), .A2(n5604), .ZN(n6882) );
  NOR2_X1 U5506 ( .A1(n8957), .A2(n6881), .ZN(n5604) );
  OR2_X1 U5507 ( .A1(n10477), .A2(n10468), .ZN(n10466) );
  NAND2_X1 U5508 ( .A1(n5328), .A2(n5326), .ZN(n10494) );
  NAND2_X1 U5509 ( .A1(n5327), .A2(n8832), .ZN(n5326) );
  INV_X1 U5510 ( .A(n5329), .ZN(n5327) );
  NOR2_X1 U5511 ( .A1(P1_IR_REG_24__SCAN_IN), .A2(n6446), .ZN(n6460) );
  INV_X1 U5512 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n6445) );
  NOR2_X1 U5513 ( .A1(P1_IR_REG_28__SCAN_IN), .A2(P1_IR_REG_27__SCAN_IN), .ZN(
        n6461) );
  AND3_X1 U5514 ( .A1(n5190), .A2(n5704), .A3(n5702), .ZN(n6831) );
  OAI21_X1 U5515 ( .B1(n6276), .B2(n6275), .A(n5831), .ZN(n6287) );
  OAI21_X1 U5516 ( .B1(n5655), .B2(n5654), .A(n6234), .ZN(n5653) );
  AND2_X1 U5517 ( .A1(n5725), .A2(n6792), .ZN(n5724) );
  OR2_X1 U5518 ( .A1(n5726), .A2(n10692), .ZN(n5725) );
  NAND2_X1 U5519 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_16__SCAN_IN), 
        .ZN(n5722) );
  INV_X1 U5520 ( .A(n6185), .ZN(n5684) );
  XNOR2_X1 U5521 ( .A(n5808), .B(n5807), .ZN(n6185) );
  INV_X1 U5522 ( .A(SI_17_), .ZN(n5807) );
  INV_X1 U5523 ( .A(n5804), .ZN(n5690) );
  NAND2_X1 U5524 ( .A1(n6644), .A2(n5193), .ZN(n6657) );
  INV_X1 U5525 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n9782) );
  INV_X1 U5526 ( .A(n5779), .ZN(n5680) );
  NAND2_X1 U5527 ( .A1(n5751), .A2(n5338), .ZN(n5337) );
  NAND2_X1 U5528 ( .A1(n5864), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n5338) );
  NAND2_X1 U5529 ( .A1(n5864), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n5741) );
  INV_X1 U5530 ( .A(n6905), .ZN(n9098) );
  INV_X1 U5531 ( .A(n8394), .ZN(n5639) );
  NAND2_X1 U5532 ( .A1(n8048), .A2(n8047), .ZN(n8112) );
  XNOR2_X1 U5533 ( .A(n6905), .B(n7074), .ZN(n6906) );
  NOR2_X1 U5534 ( .A1(n6918), .A2(n5644), .ZN(n5643) );
  INV_X1 U5535 ( .A(n5645), .ZN(n5644) );
  NAND2_X1 U5536 ( .A1(n9093), .A2(n9181), .ZN(n5613) );
  OR2_X1 U5537 ( .A1(n8618), .A2(n6870), .ZN(n7081) );
  INV_X1 U5538 ( .A(n8383), .ZN(n5636) );
  INV_X1 U5539 ( .A(n5215), .ZN(n5254) );
  AOI21_X1 U5540 ( .B1(n5732), .B2(n6896), .A(n8624), .ZN(n8473) );
  OR2_X1 U5541 ( .A1(n5959), .A2(n7016), .ZN(n5391) );
  NOR2_X1 U5542 ( .A1(n10922), .A2(n7273), .ZN(n7275) );
  NAND2_X1 U5543 ( .A1(n5577), .A2(n5575), .ZN(n5582) );
  AND2_X1 U5544 ( .A1(n5579), .A2(n5149), .ZN(n5575) );
  NAND2_X1 U5545 ( .A1(n5585), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n5584) );
  NOR2_X1 U5546 ( .A1(n7790), .A2(n6054), .ZN(n7789) );
  NAND2_X1 U5547 ( .A1(n6050), .A2(n5648), .ZN(n6205) );
  OR2_X1 U5548 ( .A1(n8273), .A2(n6120), .ZN(n5483) );
  NAND2_X1 U5549 ( .A1(n5482), .A2(n8272), .ZN(n5481) );
  INV_X1 U5550 ( .A(n5151), .ZN(n5482) );
  OR2_X1 U5551 ( .A1(n8154), .A2(n6120), .ZN(n5484) );
  AOI21_X1 U5552 ( .B1(P2_REG1_REG_14__SCAN_IN), .B2(n9269), .A(n9261), .ZN(
        n9281) );
  OAI21_X1 U5553 ( .B1(n10946), .B2(n5478), .A(n5477), .ZN(n10972) );
  NAND2_X1 U5554 ( .A1(n5479), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n5478) );
  NAND2_X1 U5555 ( .A1(n9338), .A2(n5479), .ZN(n5477) );
  INV_X1 U5556 ( .A(n10973), .ZN(n5479) );
  NOR2_X1 U5557 ( .A1(n6384), .A2(n8609), .ZN(n5556) );
  AOI21_X1 U5558 ( .B1(n8610), .B2(n5555), .A(n5184), .ZN(n5554) );
  NOR2_X1 U5559 ( .A1(n9362), .A2(n9474), .ZN(n9365) );
  NAND2_X1 U5560 ( .A1(n5471), .A2(n5162), .ZN(n9376) );
  NAND2_X1 U5561 ( .A1(n9387), .A2(n5472), .ZN(n5471) );
  OR2_X1 U5562 ( .A1(n9220), .A2(n9377), .ZN(n5472) );
  INV_X1 U5563 ( .A(n6274), .ZN(n5454) );
  INV_X1 U5564 ( .A(n9242), .ZN(n9422) );
  INV_X1 U5565 ( .A(n9433), .ZN(n5456) );
  NAND2_X1 U5566 ( .A1(n5458), .A2(n5459), .ZN(n9446) );
  AOI21_X1 U5567 ( .B1(n5138), .B2(n9483), .A(n5205), .ZN(n5459) );
  OR2_X1 U5568 ( .A1(n9502), .A2(n9501), .ZN(n9504) );
  NAND2_X1 U5569 ( .A1(n5532), .A2(n5144), .ZN(n8206) );
  OAI21_X1 U5570 ( .B1(n5972), .B2(n7282), .A(n6156), .ZN(n8477) );
  AND4_X1 U5571 ( .A1(n6074), .A2(n6073), .A3(n6072), .A4(n6071), .ZN(n8117)
         );
  NAND2_X1 U5572 ( .A1(n5540), .A2(n8456), .ZN(n7848) );
  INV_X1 U5573 ( .A(n7850), .ZN(n5540) );
  OR2_X1 U5574 ( .A1(n8618), .A2(n6930), .ZN(n9474) );
  OR2_X1 U5575 ( .A1(n6353), .A2(n5939), .ZN(n5941) );
  OR2_X1 U5576 ( .A1(n8618), .A2(n6932), .ZN(n9476) );
  INV_X1 U5577 ( .A(n6408), .ZN(n7080) );
  INV_X1 U5578 ( .A(n5972), .ZN(n8421) );
  NAND2_X1 U5579 ( .A1(n6266), .A2(n6265), .ZN(n8589) );
  INV_X1 U5580 ( .A(n9541), .ZN(n9567) );
  NAND2_X1 U5581 ( .A1(n6404), .A2(n6403), .ZN(n6946) );
  INV_X1 U5582 ( .A(n8282), .ZN(n6403) );
  NAND2_X1 U5583 ( .A1(n5858), .A2(n5473), .ZN(n5421) );
  NOR2_X1 U5584 ( .A1(n5564), .A2(P2_IR_REG_27__SCAN_IN), .ZN(n5563) );
  INV_X1 U5585 ( .A(n6348), .ZN(n9328) );
  NOR2_X1 U5586 ( .A1(P2_IR_REG_25__SCAN_IN), .A2(P2_IR_REG_24__SCAN_IN), .ZN(
        n5859) );
  NAND4_X1 U5587 ( .A1(n5526), .A2(n5525), .A3(n5562), .A4(n5473), .ZN(n6401)
         );
  INV_X1 U5588 ( .A(n5564), .ZN(n5562) );
  NAND2_X1 U5589 ( .A1(n5264), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6393) );
  INV_X1 U5590 ( .A(n6390), .ZN(n5264) );
  NAND2_X1 U5591 ( .A1(n6393), .A2(n6392), .ZN(n6395) );
  INV_X1 U5592 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n6392) );
  NAND2_X1 U5593 ( .A1(n5619), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6341) );
  INV_X1 U5594 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n6340) );
  INV_X1 U5595 ( .A(n5621), .ZN(n5620) );
  OAI21_X1 U5596 ( .B1(n6336), .B2(n5868), .A(n6340), .ZN(n5621) );
  INV_X1 U5597 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n10008) );
  NAND3_X1 U5598 ( .A1(n5278), .A2(n7111), .A3(n5276), .ZN(n5275) );
  NAND2_X1 U5599 ( .A1(n7110), .A2(n5277), .ZN(n5276) );
  OAI21_X1 U5600 ( .B1(n10104), .B2(n5281), .A(n5709), .ZN(n5280) );
  INV_X1 U5601 ( .A(n5710), .ZN(n5281) );
  INV_X1 U5602 ( .A(n6650), .ZN(n6651) );
  NAND2_X2 U5603 ( .A1(n7112), .A2(n6814), .ZN(n5152) );
  INV_X1 U5604 ( .A(n10208), .ZN(n8665) );
  NAND2_X1 U5605 ( .A1(n10185), .A2(n8691), .ZN(n10047) );
  OAI21_X1 U5606 ( .B1(n8965), .B2(n9062), .A(n6814), .ZN(n8964) );
  NAND2_X1 U5607 ( .A1(n8965), .A2(n6814), .ZN(n8974) );
  AND2_X1 U5608 ( .A1(n10416), .A2(n10271), .ZN(n9055) );
  NOR2_X1 U5609 ( .A1(n10416), .A2(n10271), .ZN(n9053) );
  INV_X1 U5610 ( .A(n7463), .ZN(n10382) );
  OR2_X1 U5611 ( .A1(n10858), .A2(n10857), .ZN(n5348) );
  AND2_X1 U5612 ( .A1(n8827), .A2(n8825), .ZN(n8961) );
  INV_X1 U5613 ( .A(n5605), .ZN(n10424) );
  NAND2_X1 U5614 ( .A1(n6745), .A2(n10484), .ZN(n6746) );
  NAND2_X1 U5615 ( .A1(n10441), .A2(n5154), .ZN(n10444) );
  AND4_X1 U5616 ( .A1(n6758), .A2(n6757), .A3(n6756), .A4(n6755), .ZN(n10462)
         );
  NAND2_X1 U5617 ( .A1(n10512), .A2(n10531), .ZN(n6717) );
  AND2_X1 U5618 ( .A1(n8901), .A2(n8977), .ZN(n10495) );
  NAND2_X1 U5619 ( .A1(n5331), .A2(n5332), .ZN(n10514) );
  NOR2_X1 U5620 ( .A1(n10513), .A2(n5330), .ZN(n5329) );
  INV_X1 U5621 ( .A(n5332), .ZN(n5330) );
  NAND2_X1 U5622 ( .A1(n10549), .A2(n5333), .ZN(n5331) );
  AND4_X1 U5623 ( .A1(n6725), .A2(n6724), .A3(n6723), .A4(n6722), .ZN(n10515)
         );
  NAND2_X1 U5624 ( .A1(n10507), .A2(n10513), .ZN(n10506) );
  AOI21_X1 U5625 ( .B1(n5523), .B2(n6678), .A(n5185), .ZN(n5521) );
  INV_X1 U5626 ( .A(n5523), .ZN(n5522) );
  OR2_X1 U5627 ( .A1(n8722), .A2(n10237), .ZN(n9021) );
  AND2_X1 U5628 ( .A1(n8887), .A2(n8889), .ZN(n8951) );
  NOR2_X1 U5629 ( .A1(n8246), .A2(n8951), .ZN(n8245) );
  OR2_X1 U5630 ( .A1(n8221), .A2(n10258), .ZN(n5731) );
  NOR2_X1 U5631 ( .A1(n8218), .A2(n10646), .ZN(n8217) );
  NAND2_X1 U5632 ( .A1(n6628), .A2(n11118), .ZN(n11123) );
  INV_X1 U5633 ( .A(n8874), .ZN(n5600) );
  OR2_X1 U5634 ( .A1(n6600), .A2(n6599), .ZN(n6606) );
  AND2_X1 U5635 ( .A1(n8872), .A2(n8874), .ZN(n8944) );
  NAND2_X1 U5636 ( .A1(n7701), .A2(n6579), .ZN(n7890) );
  NOR2_X1 U5637 ( .A1(n6562), .A2(n10167), .ZN(n6573) );
  AND4_X1 U5638 ( .A1(n6586), .A2(n6585), .A3(n6584), .A4(n6583), .ZN(n10119)
         );
  NAND2_X1 U5639 ( .A1(n5502), .A2(n5501), .ZN(n7702) );
  AOI21_X1 U5640 ( .B1(n5503), .B2(n5505), .A(n5171), .ZN(n5502) );
  NAND2_X1 U5641 ( .A1(n7702), .A2(n8940), .ZN(n7701) );
  NOR2_X2 U5642 ( .A1(n7532), .A2(n10101), .ZN(n7869) );
  INV_X1 U5643 ( .A(n5504), .ZN(n5503) );
  OAI21_X1 U5644 ( .B1(n8853), .B2(n5505), .A(n7867), .ZN(n5504) );
  INV_X1 U5645 ( .A(n6557), .ZN(n5505) );
  NAND2_X1 U5646 ( .A1(n7709), .A2(n8853), .ZN(n7708) );
  INV_X1 U5647 ( .A(n10999), .ZN(n11137) );
  AND2_X1 U5648 ( .A1(n7117), .A2(n10790), .ZN(n10999) );
  INV_X1 U5649 ( .A(n10566), .ZN(n11132) );
  NAND2_X1 U5650 ( .A1(n6760), .A2(n6759), .ZN(n10434) );
  NAND2_X1 U5651 ( .A1(n6623), .A2(n6622), .ZN(n8680) );
  NAND2_X1 U5652 ( .A1(n6841), .A2(n6859), .ZN(n10688) );
  NAND2_X1 U5653 ( .A1(n8314), .A2(n8313), .ZN(n9611) );
  XNOR2_X1 U5654 ( .A(n6452), .B(P1_IR_REG_29__SCAN_IN), .ZN(n6455) );
  NAND2_X1 U5655 ( .A1(n6302), .A2(n5839), .ZN(n5902) );
  NAND2_X1 U5656 ( .A1(n6670), .A2(n5726), .ZN(n5723) );
  NAND2_X1 U5657 ( .A1(n5651), .A2(n5816), .ZN(n6235) );
  NAND2_X1 U5658 ( .A1(n6204), .A2(n5655), .ZN(n5651) );
  NAND2_X1 U5659 ( .A1(n5284), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6680) );
  AND2_X1 U5660 ( .A1(n5286), .A2(n9791), .ZN(n5285) );
  NAND2_X1 U5661 ( .A1(n6152), .A2(n5804), .ZN(n6167) );
  NAND2_X1 U5662 ( .A1(n5320), .A2(n5318), .ZN(n6150) );
  AND2_X1 U5663 ( .A1(n5319), .A2(n5321), .ZN(n5318) );
  AND2_X1 U5664 ( .A1(n5663), .A2(n6130), .ZN(n5317) );
  AND2_X1 U5665 ( .A1(n5796), .A2(n5795), .ZN(n6108) );
  AOI21_X1 U5666 ( .B1(n6075), .B2(n5669), .A(n5667), .ZN(n5666) );
  INV_X1 U5667 ( .A(n5792), .ZN(n5667) );
  OR2_X1 U5668 ( .A1(n6076), .A2(n6075), .ZN(n5670) );
  AND2_X1 U5669 ( .A1(n5673), .A2(n5788), .ZN(n5334) );
  NAND2_X1 U5670 ( .A1(n6000), .A2(n5775), .ZN(n6013) );
  AND2_X1 U5671 ( .A1(n5779), .A2(n5778), .ZN(n6012) );
  NAND2_X1 U5672 ( .A1(n5998), .A2(n5997), .ZN(n6000) );
  INV_X1 U5673 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n5360) );
  NOR2_X2 U5674 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n6465) );
  NOR2_X1 U5675 ( .A1(n5748), .A2(n6472), .ZN(n5946) );
  NAND2_X1 U5676 ( .A1(n6138), .A2(n6137), .ZN(n9129) );
  OR2_X1 U5677 ( .A1(n8377), .A2(n5972), .ZN(n6138) );
  INV_X1 U5678 ( .A(n9125), .ZN(n9229) );
  NOR2_X1 U5679 ( .A1(n5628), .A2(n9224), .ZN(n5626) );
  AND2_X1 U5680 ( .A1(n5631), .A2(n5191), .ZN(n5628) );
  NAND2_X1 U5681 ( .A1(n5631), .A2(n5634), .ZN(n5629) );
  NAND2_X1 U5682 ( .A1(n5150), .A2(n5635), .ZN(n5634) );
  NAND2_X1 U5683 ( .A1(n5607), .A2(n5165), .ZN(n5256) );
  INV_X1 U5684 ( .A(n9244), .ZN(n9475) );
  INV_X1 U5685 ( .A(n9253), .ZN(n7936) );
  NAND2_X1 U5686 ( .A1(n7934), .A2(n7933), .ZN(n8048) );
  NAND2_X1 U5687 ( .A1(n6116), .A2(n6115), .ZN(n11103) );
  AND4_X1 U5688 ( .A1(n6284), .A2(n6283), .A3(n6282), .A4(n6281), .ZN(n9435)
         );
  AOI21_X1 U5689 ( .B1(n8412), .B2(n8411), .A(n8410), .ZN(n8414) );
  AND3_X1 U5690 ( .A1(n6929), .A2(n9553), .A3(n9609), .ZN(n9219) );
  XNOR2_X1 U5691 ( .A(n6344), .B(P2_IR_REG_22__SCAN_IN), .ZN(n8630) );
  OR2_X1 U5692 ( .A1(n7047), .A2(n9328), .ZN(n10969) );
  AND2_X1 U5693 ( .A1(P2_U3893), .A2(n6347), .ZN(n10962) );
  AND2_X1 U5694 ( .A1(n9392), .A2(n9391), .ZN(n9525) );
  OR2_X1 U5695 ( .A1(n6893), .A2(n7050), .ZN(n5440) );
  OR2_X1 U5696 ( .A1(n5972), .A2(n6949), .ZN(n5441) );
  NOR2_X1 U5697 ( .A1(n5463), .A2(n6432), .ZN(n5462) );
  INV_X1 U5698 ( .A(n5464), .ZN(n5463) );
  NAND2_X1 U5699 ( .A1(n6100), .A2(n6099), .ZN(n8203) );
  OAI21_X1 U5700 ( .B1(n10242), .B2(n5696), .A(n5694), .ZN(n5697) );
  AOI21_X1 U5701 ( .B1(n8804), .B2(n5695), .A(n8805), .ZN(n5694) );
  INV_X1 U5702 ( .A(n8804), .ZN(n5696) );
  INV_X1 U5703 ( .A(n8797), .ZN(n5695) );
  NAND2_X1 U5704 ( .A1(n6766), .A2(n6765), .ZN(n8819) );
  OR2_X1 U5705 ( .A1(n6506), .A2(n6505), .ZN(n7821) );
  AND2_X1 U5706 ( .A1(n7239), .A2(n10790), .ZN(n10261) );
  AND4_X1 U5707 ( .A1(n6764), .A2(n6763), .A3(n6762), .A4(n6761), .ZN(n10446)
         );
  NAND2_X1 U5708 ( .A1(n7127), .A2(n10580), .ZN(n10266) );
  NAND3_X1 U5709 ( .A1(n7121), .A2(n10689), .A3(n7124), .ZN(n10269) );
  NAND2_X1 U5710 ( .A1(n7449), .A2(n7450), .ZN(n10371) );
  NAND2_X1 U5711 ( .A1(n10837), .A2(n10836), .ZN(n10835) );
  NOR2_X1 U5712 ( .A1(n10851), .A2(n10850), .ZN(n10849) );
  NAND2_X1 U5713 ( .A1(n10835), .A2(n5343), .ZN(n10851) );
  OR2_X1 U5714 ( .A1(n10840), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n5343) );
  INV_X1 U5715 ( .A(n10838), .ZN(n10874) );
  NAND2_X1 U5716 ( .A1(n10881), .A2(n10854), .ZN(n5355) );
  AOI21_X1 U5717 ( .B1(n10868), .B2(P1_ADDR_REG_18__SCAN_IN), .A(n10855), .ZN(
        n5354) );
  OAI21_X1 U5718 ( .B1(n7282), .B2(n6699), .A(n6635), .ZN(n10267) );
  OR2_X1 U5719 ( .A1(n8377), .A2(n6699), .ZN(n6613) );
  NAND2_X1 U5720 ( .A1(n6598), .A2(n6597), .ZN(n8670) );
  OR2_X1 U5721 ( .A1(n7031), .A2(n6699), .ZN(n6598) );
  OR2_X1 U5722 ( .A1(n11011), .A2(n7110), .ZN(n11153) );
  OR2_X1 U5723 ( .A1(n7126), .A2(n7125), .ZN(n10580) );
  NAND2_X1 U5724 ( .A1(n5428), .A2(n5161), .ZN(n7729) );
  INV_X1 U5725 ( .A(n11014), .ZN(n11151) );
  AND2_X1 U5726 ( .A1(n8346), .A2(n8343), .ZN(n5309) );
  INV_X1 U5727 ( .A(n10434), .ZN(n10656) );
  OR2_X1 U5728 ( .A1(n6859), .A2(n6858), .ZN(n10691) );
  MUX2_X1 U5729 ( .A(n8498), .B(n8497), .S(n8588), .Z(n8499) );
  NAND2_X1 U5730 ( .A1(n8495), .A2(n8511), .ZN(n8498) );
  INV_X1 U5731 ( .A(n7831), .ZN(n8846) );
  AND2_X1 U5732 ( .A1(n8516), .A2(n8512), .ZN(n5366) );
  NAND2_X1 U5733 ( .A1(n8854), .A2(n5222), .ZN(n8859) );
  NOR4_X1 U5734 ( .A1(n8510), .A2(n8588), .A3(n8509), .A4(n8508), .ZN(n8523)
         );
  NAND2_X1 U5735 ( .A1(n5363), .A2(n5362), .ZN(n8522) );
  OAI21_X1 U5736 ( .B1(n5228), .B2(n5597), .A(n5227), .ZN(n5226) );
  NOR2_X1 U5737 ( .A1(n8984), .A2(n8920), .ZN(n5227) );
  AOI21_X1 U5738 ( .B1(n8876), .B2(n5143), .A(n6799), .ZN(n5228) );
  OAI21_X1 U5739 ( .B1(n5232), .B2(n8877), .A(n5230), .ZN(n5229) );
  NOR2_X1 U5740 ( .A1(n5597), .A2(n5231), .ZN(n5230) );
  AOI21_X1 U5741 ( .B1(n8876), .B2(n9010), .A(n8875), .ZN(n5232) );
  NAND2_X1 U5742 ( .A1(n9015), .A2(n8920), .ZN(n5231) );
  NAND2_X1 U5743 ( .A1(n5237), .A2(n8892), .ZN(n5236) );
  NAND2_X1 U5744 ( .A1(n8891), .A2(n9027), .ZN(n5237) );
  AOI21_X1 U5745 ( .B1(n8885), .B2(n5157), .A(n8896), .ZN(n5235) );
  AOI21_X1 U5746 ( .B1(n5388), .B2(n8574), .A(n8571), .ZN(n5387) );
  NAND2_X1 U5747 ( .A1(n8573), .A2(n9164), .ZN(n5388) );
  OR2_X1 U5748 ( .A1(n8576), .A2(n8588), .ZN(n5386) );
  NOR2_X1 U5749 ( .A1(n8571), .A2(n8618), .ZN(n5384) );
  OR2_X1 U5750 ( .A1(n8575), .A2(n5380), .ZN(n5379) );
  NAND2_X1 U5751 ( .A1(n8573), .A2(n8572), .ZN(n5385) );
  AOI21_X1 U5752 ( .B1(n5412), .B2(n5415), .A(n5186), .ZN(n5411) );
  AOI21_X1 U5753 ( .B1(n5233), .B2(n8900), .A(n10513), .ZN(n8903) );
  AOI21_X1 U5754 ( .B1(n5411), .B2(n5409), .A(n9424), .ZN(n5408) );
  INV_X1 U5755 ( .A(n5412), .ZN(n5409) );
  INV_X1 U5756 ( .A(n5411), .ZN(n5410) );
  INV_X1 U5757 ( .A(n5556), .ZN(n5551) );
  AOI21_X1 U5758 ( .B1(n8598), .B2(n5376), .A(n5375), .ZN(n5374) );
  OR2_X1 U5759 ( .A1(n8599), .A2(n8600), .ZN(n5376) );
  INV_X1 U5760 ( .A(n9400), .ZN(n5375) );
  NOR2_X1 U5761 ( .A1(n9380), .A2(n8607), .ZN(n5370) );
  NAND2_X1 U5762 ( .A1(n5373), .A2(n5372), .ZN(n5371) );
  INV_X1 U5763 ( .A(n8603), .ZN(n5372) );
  INV_X1 U5764 ( .A(n5554), .ZN(n5553) );
  INV_X1 U5765 ( .A(n9282), .ZN(n5574) );
  INV_X1 U5766 ( .A(n9001), .ZN(n8942) );
  OAI21_X1 U5767 ( .B1(n8926), .B2(n9053), .A(n5240), .ZN(n5239) );
  INV_X1 U5768 ( .A(n8923), .ZN(n5240) );
  AOI21_X1 U5769 ( .B1(n5246), .B2(n5244), .A(n5243), .ZN(n8917) );
  AND2_X1 U5770 ( .A1(n8915), .A2(n8920), .ZN(n5243) );
  INV_X1 U5771 ( .A(n5316), .ZN(n5314) );
  INV_X1 U5772 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n9780) );
  NOR2_X1 U5773 ( .A1(n5901), .A2(n5661), .ZN(n5660) );
  INV_X1 U5774 ( .A(n5839), .ZN(n5661) );
  INV_X1 U5775 ( .A(SI_27_), .ZN(n9825) );
  INV_X1 U5776 ( .A(SI_20_), .ZN(n9641) );
  INV_X1 U5777 ( .A(SI_16_), .ZN(n9645) );
  INV_X1 U5778 ( .A(n7385), .ZN(n5259) );
  AOI21_X1 U5779 ( .B1(n5400), .B2(n5404), .A(n5399), .ZN(n5398) );
  INV_X1 U5780 ( .A(n8623), .ZN(n5399) );
  INV_X1 U5781 ( .A(n5189), .ZN(n5404) );
  NOR2_X1 U5782 ( .A1(P2_IR_REG_15__SCAN_IN), .A2(P2_IR_REG_11__SCAN_IN), .ZN(
        n5850) );
  NOR2_X1 U5783 ( .A1(P2_IR_REG_20__SCAN_IN), .A2(P2_IR_REG_13__SCAN_IN), .ZN(
        n5851) );
  NAND2_X1 U5784 ( .A1(n8358), .A2(n7044), .ZN(n7245) );
  OR2_X1 U5785 ( .A1(n10907), .A2(n7270), .ZN(n5566) );
  NAND2_X1 U5786 ( .A1(n5566), .A2(n7272), .ZN(n7271) );
  NAND2_X1 U5787 ( .A1(n7428), .A2(n5474), .ZN(n7605) );
  OR2_X1 U5788 ( .A1(n7429), .A2(n7515), .ZN(n5474) );
  INV_X1 U5789 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n6049) );
  NAND2_X1 U5790 ( .A1(n7977), .A2(n7976), .ZN(n8091) );
  AND2_X1 U5791 ( .A1(n6049), .A2(n6077), .ZN(n5648) );
  INV_X1 U5792 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n6077) );
  OR2_X1 U5793 ( .A1(n5896), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n5889) );
  NOR2_X1 U5794 ( .A1(n6191), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n6192) );
  OR2_X1 U5795 ( .A1(n9129), .A2(n9247), .ZN(n6365) );
  AND2_X1 U5796 ( .A1(n7080), .A2(n9610), .ZN(n6865) );
  OR2_X1 U5797 ( .A1(n6946), .A2(n6421), .ZN(n6866) );
  NAND2_X1 U5798 ( .A1(n5691), .A2(n5164), .ZN(n5692) );
  NAND2_X1 U5799 ( .A1(n10106), .A2(n8765), .ZN(n10057) );
  NAND2_X1 U5800 ( .A1(n5706), .A2(n5707), .ZN(n5282) );
  AOI21_X1 U5801 ( .B1(n10135), .B2(n8718), .A(n5708), .ZN(n5707) );
  INV_X1 U5802 ( .A(n10143), .ZN(n5708) );
  NAND2_X1 U5803 ( .A1(n10656), .A2(n10446), .ZN(n5499) );
  INV_X1 U5804 ( .A(n5496), .ZN(n5494) );
  NAND2_X1 U5805 ( .A1(n5496), .A2(n5492), .ZN(n5491) );
  INV_X1 U5806 ( .A(n10442), .ZN(n5492) );
  AND2_X1 U5807 ( .A1(P1_REG3_REG_25__SCAN_IN), .A2(n6740), .ZN(n6751) );
  AND2_X1 U5808 ( .A1(n8980), .A2(n9035), .ZN(n8955) );
  AND2_X1 U5809 ( .A1(n10546), .A2(n5521), .ZN(n5518) );
  AND2_X1 U5810 ( .A1(n9030), .A2(n8897), .ZN(n10528) );
  AND2_X1 U5811 ( .A1(n8952), .A2(n9019), .ZN(n5316) );
  NOR2_X1 U5812 ( .A1(n7898), .A2(n8670), .ZN(n7883) );
  NAND2_X1 U5813 ( .A1(n9012), .A2(n8873), .ZN(n11120) );
  NAND2_X1 U5814 ( .A1(n7891), .A2(n9005), .ZN(n7876) );
  NOR2_X1 U5815 ( .A1(n10080), .A2(n10172), .ZN(n5431) );
  NOR2_X1 U5816 ( .A1(n6807), .A2(n5603), .ZN(n9001) );
  NAND2_X1 U5817 ( .A1(n6805), .A2(n7524), .ZN(n5603) );
  NAND2_X1 U5818 ( .A1(n7639), .A2(n7834), .ZN(n8935) );
  OR2_X1 U5819 ( .A1(n7839), .A2(n7639), .ZN(n7532) );
  OR2_X1 U5820 ( .A1(n11001), .A2(n11032), .ZN(n8993) );
  NAND2_X1 U5821 ( .A1(n8217), .A2(n10686), .ZN(n8251) );
  NAND2_X1 U5822 ( .A1(n6805), .A2(n8935), .ZN(n8849) );
  OR2_X1 U5823 ( .A1(n6543), .A2(n7831), .ZN(n7520) );
  XNOR2_X1 U5824 ( .A(n6321), .B(n6322), .ZN(n6319) );
  NOR2_X1 U5825 ( .A1(n6788), .A2(P1_IR_REG_17__SCAN_IN), .ZN(n5726) );
  INV_X1 U5826 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n6679) );
  INV_X1 U5827 ( .A(SI_18_), .ZN(n9845) );
  AND2_X1 U5828 ( .A1(n5193), .A2(n9999), .ZN(n5286) );
  AOI21_X1 U5829 ( .B1(n6130), .B2(n5323), .A(n5322), .ZN(n5321) );
  INV_X1 U5830 ( .A(n5800), .ZN(n5322) );
  INV_X1 U5831 ( .A(n5796), .ZN(n5323) );
  INV_X1 U5832 ( .A(SI_14_), .ZN(n9853) );
  OAI21_X1 U5833 ( .B1(n5755), .B2(n5757), .A(n5756), .ZN(n5758) );
  NAND2_X1 U5834 ( .A1(n5755), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n5756) );
  NAND2_X1 U5835 ( .A1(n5337), .A2(SI_2_), .ZN(n5754) );
  AND2_X2 U5836 ( .A1(n5251), .A2(n5250), .ZN(n5864) );
  INV_X1 U5837 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n5289) );
  INV_X1 U5838 ( .A(n9101), .ZN(n5630) );
  OR2_X1 U5839 ( .A1(n5611), .A2(n5610), .ZN(n5609) );
  NAND2_X1 U5840 ( .A1(n8392), .A2(n8391), .ZN(n9170) );
  INV_X1 U5841 ( .A(n9172), .ZN(n8392) );
  OR2_X1 U5842 ( .A1(n6082), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n6102) );
  AOI21_X1 U5843 ( .B1(n5398), .B2(n5401), .A(n8472), .ZN(n5396) );
  NAND2_X1 U5844 ( .A1(n5367), .A2(n5170), .ZN(n8614) );
  NAND2_X1 U5845 ( .A1(n5396), .A2(n5397), .ZN(n5395) );
  INV_X1 U5846 ( .A(n5398), .ZN(n5397) );
  XNOR2_X1 U5847 ( .A(n7245), .B(n7060), .ZN(n7045) );
  INV_X1 U5848 ( .A(n5568), .ZN(n5567) );
  NAND2_X1 U5849 ( .A1(n5569), .A2(n5571), .ZN(n7056) );
  AND2_X1 U5850 ( .A1(n5568), .A2(n5571), .ZN(n10909) );
  OAI21_X1 U5851 ( .B1(n5566), .B2(n7272), .A(n7271), .ZN(n10923) );
  NAND2_X1 U5852 ( .A1(n10924), .A2(n7250), .ZN(n7251) );
  NAND2_X1 U5853 ( .A1(n7251), .A2(n7252), .ZN(n7428) );
  NAND2_X1 U5854 ( .A1(n5583), .A2(n5580), .ZN(n5578) );
  XNOR2_X1 U5855 ( .A(n7605), .B(n7430), .ZN(n7431) );
  AND2_X1 U5856 ( .A1(n6050), .A2(n6049), .ZN(n6078) );
  NOR2_X1 U5857 ( .A1(n10946), .A2(n9318), .ZN(n10945) );
  NAND2_X1 U5858 ( .A1(n5886), .A2(n5885), .ZN(n9099) );
  OR2_X1 U5859 ( .A1(n6307), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n6309) );
  NAND2_X1 U5860 ( .A1(n6297), .A2(n8466), .ZN(n9401) );
  OAI21_X1 U5861 ( .B1(n9433), .B2(n5450), .A(n5449), .ZN(n6297) );
  INV_X1 U5862 ( .A(n5451), .ZN(n5450) );
  AOI21_X1 U5863 ( .B1(n5451), .B2(n5452), .A(n8597), .ZN(n5449) );
  NAND2_X1 U5864 ( .A1(n5221), .A2(n9919), .ZN(n6279) );
  OR2_X1 U5865 ( .A1(n6279), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n6290) );
  INV_X1 U5866 ( .A(n6239), .ZN(n5873) );
  INV_X1 U5867 ( .A(n5221), .ZN(n6267) );
  NAND2_X1 U5868 ( .A1(n6213), .A2(n9889), .ZN(n6239) );
  INV_X1 U5869 ( .A(n9448), .ZN(n9477) );
  INV_X1 U5870 ( .A(n6227), .ZN(n6213) );
  AOI21_X1 U5871 ( .B1(n8558), .B2(n5445), .A(n5158), .ZN(n5443) );
  OR2_X1 U5872 ( .A1(n6175), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n6191) );
  NAND2_X1 U5873 ( .A1(n8564), .A2(n8565), .ZN(n8483) );
  INV_X1 U5874 ( .A(n6372), .ZN(n5529) );
  INV_X1 U5875 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n9228) );
  NAND2_X1 U5876 ( .A1(n6369), .A2(n5740), .ZN(n8105) );
  INV_X1 U5877 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n9884) );
  AND2_X1 U5878 ( .A1(n6139), .A2(n9884), .ZN(n6157) );
  INV_X1 U5879 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n9915) );
  AND2_X1 U5880 ( .A1(n6118), .A2(n9915), .ZN(n6139) );
  INV_X1 U5881 ( .A(n8554), .ZN(n8457) );
  AND4_X1 U5882 ( .A1(n6107), .A2(n6106), .A3(n6105), .A4(n6104), .ZN(n8174)
         );
  NOR2_X1 U5883 ( .A1(n5537), .A2(n5536), .ZN(n5535) );
  NOR2_X1 U5884 ( .A1(n8456), .A2(n5538), .ZN(n5537) );
  AND2_X1 U5885 ( .A1(n8536), .A2(n8545), .ZN(n8443) );
  OR2_X1 U5886 ( .A1(n6069), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n6082) );
  INV_X1 U5887 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n6055) );
  INV_X1 U5888 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n9896) );
  AND2_X1 U5889 ( .A1(n6036), .A2(n9896), .ZN(n6056) );
  INV_X1 U5890 ( .A(n9252), .ZN(n8050) );
  AND2_X1 U5891 ( .A1(n7661), .A2(n8529), .ZN(n8521) );
  NAND2_X1 U5892 ( .A1(n7510), .A2(n8450), .ZN(n5559) );
  OR2_X1 U5893 ( .A1(n6004), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n6021) );
  NOR2_X1 U5894 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n5978) );
  OAI21_X1 U5895 ( .B1(n6899), .B2(n9259), .A(n5528), .ZN(n7315) );
  INV_X1 U5896 ( .A(n7299), .ZN(n5527) );
  OR2_X1 U5897 ( .A1(n8618), .A2(n6869), .ZN(n7091) );
  NAND2_X1 U5898 ( .A1(n7088), .A2(n7087), .ZN(n7090) );
  NAND2_X1 U5899 ( .A1(n8423), .A2(n8422), .ZN(n9346) );
  NAND2_X1 U5900 ( .A1(n7848), .A2(n6363), .ZN(n7963) );
  OR2_X1 U5901 ( .A1(n5966), .A2(n5757), .ZN(n5918) );
  XNOR2_X1 U5902 ( .A(n6429), .B(n5473), .ZN(n7011) );
  NAND2_X1 U5903 ( .A1(n5849), .A2(n5847), .ZN(n5624) );
  INV_X1 U5904 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n5623) );
  OR2_X1 U5905 ( .A1(n5926), .A2(P2_IR_REG_3__SCAN_IN), .ZN(n5928) );
  NAND2_X1 U5906 ( .A1(n5437), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5965) );
  INV_X1 U5907 ( .A(n6720), .ZN(n6721) );
  NAND2_X1 U5908 ( .A1(n6721), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n6730) );
  NAND2_X1 U5909 ( .A1(n5698), .A2(n5167), .ZN(n10072) );
  INV_X1 U5910 ( .A(n8656), .ZN(n5700) );
  AND2_X1 U5911 ( .A1(n10042), .A2(n10043), .ZN(n8804) );
  INV_X1 U5912 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n6550) );
  INV_X1 U5913 ( .A(n6739), .ZN(n6740) );
  OR2_X1 U5914 ( .A1(n10134), .A2(n10135), .ZN(n10132) );
  NAND2_X1 U5915 ( .A1(n6662), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n6673) );
  AOI21_X1 U5916 ( .B1(n5712), .B2(n10105), .A(n5176), .ZN(n5710) );
  INV_X1 U5917 ( .A(n5712), .ZN(n5711) );
  INV_X1 U5918 ( .A(n10104), .ZN(n8760) );
  NAND2_X1 U5919 ( .A1(n6685), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n6691) );
  NAND2_X1 U5920 ( .A1(n10212), .A2(n8675), .ZN(n10184) );
  INV_X1 U5921 ( .A(n6711), .ZN(n6712) );
  AND2_X1 U5922 ( .A1(n10245), .A2(n10241), .ZN(n8797) );
  NAND2_X1 U5923 ( .A1(n5716), .A2(n5714), .ZN(n8698) );
  AOI21_X1 U5924 ( .B1(n5717), .B2(n5719), .A(n5715), .ZN(n5714) );
  NAND2_X1 U5925 ( .A1(n8974), .A2(n8967), .ZN(n8968) );
  NAND2_X1 U5926 ( .A1(n8822), .A2(n10272), .ZN(n9051) );
  NAND2_X1 U5927 ( .A1(n6520), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n6476) );
  OR2_X1 U5928 ( .A1(n7163), .A2(n7162), .ZN(n5357) );
  NOR2_X1 U5929 ( .A1(n7445), .A2(n5349), .ZN(n10357) );
  AND2_X1 U5930 ( .A1(n7453), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n5349) );
  NAND2_X1 U5931 ( .A1(n10357), .A2(n10356), .ZN(n10355) );
  OR2_X1 U5932 ( .A1(n10814), .A2(n10815), .ZN(n5346) );
  AND2_X1 U5933 ( .A1(n5346), .A2(n5345), .ZN(n10373) );
  NAND2_X1 U5934 ( .A1(n10818), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n5345) );
  OR2_X1 U5935 ( .A1(n6886), .A2(n5433), .ZN(n9072) );
  NAND2_X1 U5936 ( .A1(n8822), .A2(n5434), .ZN(n5433) );
  INV_X1 U5937 ( .A(n5434), .ZN(n5432) );
  NOR2_X1 U5938 ( .A1(n10450), .A2(n10466), .ZN(n10449) );
  AND2_X1 U5939 ( .A1(n9038), .A2(n8908), .ZN(n10458) );
  AND4_X1 U5940 ( .A1(n6735), .A2(n6734), .A3(n6733), .A4(n6732), .ZN(n10496)
         );
  NOR2_X1 U5941 ( .A1(n10603), .A2(n5424), .ZN(n5423) );
  INV_X1 U5942 ( .A(n5425), .ZN(n5424) );
  INV_X1 U5943 ( .A(n5509), .ZN(n5508) );
  NAND2_X1 U5944 ( .A1(n10535), .A2(n6707), .ZN(n10536) );
  AND4_X1 U5945 ( .A1(n6695), .A2(n6694), .A3(n6693), .A4(n6692), .ZN(n10568)
         );
  AND2_X1 U5946 ( .A1(n8951), .A2(n9021), .ZN(n5596) );
  NAND2_X1 U5947 ( .A1(n8222), .A2(n5316), .ZN(n8248) );
  NAND2_X1 U5948 ( .A1(n8222), .A2(n9019), .ZN(n8178) );
  OR2_X1 U5949 ( .A1(n11127), .A2(n10267), .ZN(n8218) );
  INV_X1 U5950 ( .A(n5295), .ZN(n5294) );
  OAI21_X1 U5951 ( .B1(n6630), .B2(n5296), .A(n6642), .ZN(n5295) );
  INV_X1 U5952 ( .A(n6636), .ZN(n6637) );
  NAND2_X1 U5953 ( .A1(n6637), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n6650) );
  NAND2_X1 U5954 ( .A1(n11131), .A2(n9012), .ZN(n8063) );
  AND4_X1 U5955 ( .A1(n6656), .A2(n6655), .A3(n6654), .A4(n6653), .ZN(n10258)
         );
  NOR2_X1 U5956 ( .A1(n8948), .A2(n5597), .ZN(n5311) );
  INV_X1 U5957 ( .A(n5305), .ZN(n5304) );
  AOI21_X1 U5958 ( .B1(n5512), .B2(n5515), .A(n5169), .ZN(n5511) );
  NAND2_X1 U5959 ( .A1(n7876), .A2(n8985), .ZN(n7916) );
  NAND2_X1 U5960 ( .A1(n6581), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n6600) );
  INV_X1 U5961 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n6599) );
  NAND2_X1 U5962 ( .A1(n7869), .A2(n5429), .ZN(n7898) );
  NOR2_X1 U5963 ( .A1(n5430), .A2(n8663), .ZN(n5429) );
  INV_X1 U5964 ( .A(n5431), .ZN(n5430) );
  NAND2_X1 U5965 ( .A1(n7869), .A2(n5431), .ZN(n7897) );
  AND4_X1 U5966 ( .A1(n6578), .A2(n6577), .A3(n6576), .A4(n6575), .ZN(n8654)
         );
  AND2_X1 U5967 ( .A1(n6573), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n6581) );
  NAND2_X1 U5968 ( .A1(n9003), .A2(n5602), .ZN(n7697) );
  NAND2_X1 U5969 ( .A1(n7525), .A2(n9001), .ZN(n5602) );
  AND4_X1 U5970 ( .A1(n6567), .A2(n6566), .A3(n6565), .A4(n6564), .ZN(n10096)
         );
  OR2_X1 U5971 ( .A1(n7412), .A2(n7415), .ZN(n7829) );
  NAND2_X1 U5972 ( .A1(n7524), .A2(n8998), .ZN(n7831) );
  AND4_X1 U5973 ( .A1(n6512), .A2(n6511), .A3(n6510), .A4(n6509), .ZN(n7833)
         );
  NOR2_X1 U5974 ( .A1(n7816), .A2(n7821), .ZN(n7819) );
  NOR2_X1 U5975 ( .A1(n7128), .A2(n7729), .ZN(n10996) );
  NAND2_X1 U5976 ( .A1(n10996), .A2(n11013), .ZN(n10995) );
  INV_X1 U5977 ( .A(n10577), .ZN(n11126) );
  NAND2_X1 U5978 ( .A1(n6781), .A2(n6780), .ZN(n8334) );
  OAI21_X1 U5979 ( .B1(n10444), .B2(n6881), .A(n5324), .ZN(n6883) );
  NAND2_X1 U5980 ( .A1(n6738), .A2(n6737), .ZN(n10468) );
  OR2_X1 U5981 ( .A1(n8163), .A2(n6699), .ZN(n6738) );
  NAND2_X1 U5982 ( .A1(n6710), .A2(n6709), .ZN(n10613) );
  OR2_X1 U5983 ( .A1(n7997), .A2(n6699), .ZN(n6710) );
  OR2_X1 U5984 ( .A1(n9108), .A2(n6699), .ZN(n6701) );
  NAND2_X1 U5985 ( .A1(n6661), .A2(n6660), .ZN(n8722) );
  AND2_X1 U5986 ( .A1(n6531), .A2(n6530), .ZN(n11053) );
  NOR2_X1 U5987 ( .A1(n5278), .A2(n7107), .ZN(n10985) );
  INV_X1 U5988 ( .A(n6484), .ZN(n11013) );
  AND3_X1 U5989 ( .A1(n10689), .A2(n7119), .A3(n7130), .ZN(n7209) );
  AND2_X1 U5990 ( .A1(n7125), .A2(n7118), .ZN(n6888) );
  AND2_X1 U5991 ( .A1(n6461), .A2(n6460), .ZN(n6447) );
  INV_X1 U5992 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n10022) );
  XNOR2_X1 U5993 ( .A(n6320), .B(n6319), .ZN(n8293) );
  XNOR2_X1 U5994 ( .A(n6840), .B(P1_IR_REG_26__SCAN_IN), .ZN(n6859) );
  NAND2_X1 U5995 ( .A1(n6839), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6840) );
  NOR2_X1 U5996 ( .A1(n6835), .A2(P1_IR_REG_24__SCAN_IN), .ZN(n6833) );
  NAND2_X1 U5997 ( .A1(n6833), .A2(n10013), .ZN(n6839) );
  AND2_X1 U5998 ( .A1(n5827), .A2(n5826), .ZN(n6261) );
  OAI22_X1 U5999 ( .A1(n6204), .A2(n5650), .B1(n5652), .B2(n5818), .ZN(n6244)
         );
  NAND2_X1 U6000 ( .A1(n5816), .A2(n5657), .ZN(n5650) );
  INV_X1 U6001 ( .A(n5653), .ZN(n5652) );
  INV_X1 U6002 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n6794) );
  AND2_X1 U6003 ( .A1(n5724), .A2(n5722), .ZN(n5721) );
  INV_X1 U6004 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n9796) );
  NAND2_X1 U6005 ( .A1(n5689), .A2(n6185), .ZN(n5685) );
  INV_X1 U6006 ( .A(n5683), .ZN(n5682) );
  OAI21_X1 U6007 ( .B1(n5686), .B2(n5684), .A(n5207), .ZN(n5683) );
  NOR2_X1 U6008 ( .A1(n6443), .A2(P1_IR_REG_12__SCAN_IN), .ZN(n5705) );
  INV_X1 U6009 ( .A(n5674), .ZN(n5673) );
  OAI21_X1 U6010 ( .B1(n5676), .B2(n5675), .A(n5177), .ZN(n5674) );
  INV_X1 U6011 ( .A(n6044), .ZN(n5675) );
  NAND2_X1 U6012 ( .A1(n5336), .A2(n6000), .ZN(n5335) );
  AND2_X1 U6013 ( .A1(n5141), .A2(n5775), .ZN(n5336) );
  OR2_X1 U6014 ( .A1(n6558), .A2(P1_IR_REG_8__SCAN_IN), .ZN(n6559) );
  OAI21_X1 U6015 ( .B1(n6013), .B2(n5678), .A(n5676), .ZN(n6045) );
  OR2_X1 U6016 ( .A1(n6547), .A2(P1_IR_REG_7__SCAN_IN), .ZN(n6558) );
  NAND2_X1 U6017 ( .A1(n5987), .A2(n5770), .ZN(n5998) );
  OAI21_X1 U6018 ( .B1(SI_2_), .B2(n5337), .A(n5754), .ZN(n5968) );
  NAND2_X1 U6019 ( .A1(n5749), .A2(n5946), .ZN(n5950) );
  AND2_X1 U6020 ( .A1(n5642), .A2(n5142), .ZN(n7686) );
  NAND2_X1 U6021 ( .A1(n5255), .A2(n5635), .ZN(n9112) );
  INV_X1 U6022 ( .A(n9110), .ZN(n5255) );
  NAND2_X1 U6023 ( .A1(n6278), .A2(n6277), .ZN(n9425) );
  NAND2_X1 U6024 ( .A1(n5140), .A2(n6903), .ZN(n5615) );
  NAND2_X1 U6025 ( .A1(n7073), .A2(n5140), .ZN(n5614) );
  NAND2_X1 U6026 ( .A1(n5640), .A2(n5172), .ZN(n5638) );
  NAND2_X1 U6027 ( .A1(n6304), .A2(n6303), .ZN(n9529) );
  INV_X1 U6028 ( .A(n9255), .ZN(n7689) );
  AND4_X1 U6029 ( .A1(n5925), .A2(n5924), .A3(n5923), .A4(n5922), .ZN(n7478)
         );
  OR2_X1 U6030 ( .A1(n6353), .A2(n5919), .ZN(n5925) );
  NAND2_X1 U6031 ( .A1(n6289), .A2(n6288), .ZN(n9188) );
  AND2_X1 U6032 ( .A1(n5261), .A2(n7219), .ZN(n7387) );
  INV_X1 U6033 ( .A(n5262), .ZN(n5261) );
  NAND2_X1 U6034 ( .A1(n7219), .A2(n6910), .ZN(n7321) );
  OR2_X1 U6035 ( .A1(n6935), .A2(n6934), .ZN(n9125) );
  AOI21_X1 U6036 ( .B1(n7931), .B2(n7930), .A(n5729), .ZN(n7934) );
  INV_X1 U6037 ( .A(n9231), .ZN(n9214) );
  AOI22_X1 U6038 ( .A1(n8115), .A2(n8117), .B1(n8114), .B2(n8113), .ZN(n8194)
         );
  NAND2_X1 U6039 ( .A1(n6080), .A2(n6079), .ZN(n8122) );
  XNOR2_X1 U6040 ( .A(n6906), .B(n7289), .ZN(n7073) );
  NOR2_X1 U6041 ( .A1(n7064), .A2(n6904), .ZN(n7072) );
  NAND2_X1 U6042 ( .A1(n7384), .A2(n5645), .ZN(n6917) );
  INV_X1 U6043 ( .A(n5642), .ZN(n7683) );
  NAND2_X1 U6044 ( .A1(n5613), .A2(n5611), .ZN(n5608) );
  XNOR2_X1 U6045 ( .A(n9096), .B(n9377), .ZN(n9213) );
  NAND2_X1 U6046 ( .A1(n5904), .A2(n5903), .ZN(n9220) );
  NAND2_X1 U6047 ( .A1(n5253), .A2(n5252), .ZN(n9226) );
  AOI21_X1 U6048 ( .B1(n5254), .B2(n8380), .A(n5187), .ZN(n5252) );
  NAND2_X1 U6049 ( .A1(n9119), .A2(n8380), .ZN(n5637) );
  OR2_X1 U6050 ( .A1(n5956), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n5908) );
  NAND2_X1 U6051 ( .A1(n6329), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n5390) );
  OR2_X1 U6052 ( .A1(n5956), .A2(n7095), .ZN(n5392) );
  INV_X2 U6053 ( .A(P2_U3893), .ZN(n10977) );
  OR2_X1 U6054 ( .A1(P2_U3150), .A2(n7013), .ZN(n10938) );
  AND2_X1 U6055 ( .A1(n5581), .A2(n5582), .ZN(n7593) );
  NAND2_X1 U6056 ( .A1(n5156), .A2(n5580), .ZN(n5581) );
  INV_X1 U6057 ( .A(n5587), .ZN(n5586) );
  INV_X1 U6058 ( .A(n5591), .ZN(n8079) );
  OR2_X1 U6059 ( .A1(n7990), .A2(n6081), .ZN(n5591) );
  INV_X1 U6060 ( .A(n8080), .ZN(n5590) );
  OAI21_X1 U6061 ( .B1(n7990), .B2(n5589), .A(n5588), .ZN(n8144) );
  NAND2_X1 U6062 ( .A1(n5592), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n5589) );
  INV_X1 U6063 ( .A(n8081), .ZN(n5592) );
  NOR2_X1 U6064 ( .A1(n8145), .A2(n6117), .ZN(n8258) );
  NAND2_X1 U6065 ( .A1(n5481), .A2(n5480), .ZN(n9268) );
  NAND2_X1 U6066 ( .A1(n5595), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n5594) );
  INV_X1 U6067 ( .A(n8260), .ZN(n5595) );
  AND2_X1 U6068 ( .A1(n6187), .A2(n6172), .ZN(n9307) );
  NOR2_X1 U6069 ( .A1(n9283), .A2(n9282), .ZN(n9285) );
  INV_X1 U6070 ( .A(n10976), .ZN(n10941) );
  OAI21_X1 U6071 ( .B1(n9345), .B2(n10969), .A(n5487), .ZN(n5486) );
  INV_X1 U6072 ( .A(n9343), .ZN(n5487) );
  NOR2_X1 U6073 ( .A1(n10972), .A2(n9340), .ZN(n9341) );
  OR2_X1 U6074 ( .A1(n7047), .A2(n9324), .ZN(n10974) );
  NAND2_X1 U6075 ( .A1(n5547), .A2(n5554), .ZN(n8425) );
  OAI21_X1 U6076 ( .B1(n9367), .B2(n9471), .A(n9366), .ZN(n9516) );
  NOR2_X1 U6077 ( .A1(n9365), .A2(n9364), .ZN(n9366) );
  INV_X1 U6078 ( .A(n9099), .ZN(n9522) );
  NAND2_X1 U6079 ( .A1(n5448), .A2(n5451), .ZN(n9410) );
  NAND2_X1 U6080 ( .A1(n9433), .A2(n5453), .ZN(n5448) );
  NAND2_X1 U6081 ( .A1(n5455), .A2(n6274), .ZN(n9419) );
  NAND2_X1 U6082 ( .A1(n5456), .A2(n5457), .ZN(n5455) );
  NAND2_X1 U6083 ( .A1(n5561), .A2(n6379), .ZN(n9423) );
  NAND2_X1 U6084 ( .A1(n6250), .A2(n6249), .ZN(n9545) );
  NAND2_X1 U6085 ( .A1(n6237), .A2(n6236), .ZN(n9549) );
  NAND2_X1 U6086 ( .A1(n9473), .A2(n5138), .ZN(n9458) );
  AND2_X1 U6087 ( .A1(n9473), .A2(n6233), .ZN(n9460) );
  NAND2_X1 U6088 ( .A1(n9504), .A2(n8577), .ZN(n9484) );
  NAND2_X1 U6089 ( .A1(n6226), .A2(n6225), .ZN(n9554) );
  NAND2_X1 U6090 ( .A1(n6212), .A2(n6211), .ZN(n9508) );
  NAND2_X1 U6091 ( .A1(n5532), .A2(n5530), .ZN(n8208) );
  NAND2_X1 U6092 ( .A1(n6190), .A2(n6189), .ZN(n9178) );
  INV_X1 U6093 ( .A(n11104), .ZN(n9439) );
  OR2_X1 U6094 ( .A1(n7090), .A2(n11105), .ZN(n9441) );
  AND2_X1 U6095 ( .A1(n11111), .A2(n11110), .ZN(n9443) );
  INV_X1 U6096 ( .A(n9488), .ZN(n11111) );
  INV_X1 U6097 ( .A(n9441), .ZN(n9509) );
  NAND2_X2 U6098 ( .A1(n6874), .A2(n6873), .ZN(n9572) );
  INV_X1 U6099 ( .A(n9346), .ZN(n9575) );
  AOI21_X1 U6100 ( .B1(n9069), .B2(n8421), .A(n8420), .ZN(n9578) );
  NOR2_X1 U6101 ( .A1(n9516), .A2(n9515), .ZN(n9579) );
  AND2_X1 U6102 ( .A1(n9514), .A2(n9541), .ZN(n9515) );
  AND2_X1 U6103 ( .A1(n9525), .A2(n9524), .ZN(n9584) );
  INV_X1 U6104 ( .A(n8589), .ZN(n9600) );
  AND2_X1 U6105 ( .A1(n9560), .A2(n9559), .ZN(n9605) );
  INV_X1 U6106 ( .A(n7223), .ZN(n7468) );
  AND2_X1 U6107 ( .A1(n7011), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6947) );
  INV_X1 U6108 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n9613) );
  INV_X1 U6109 ( .A(n5871), .ZN(n8332) );
  NAND2_X1 U6110 ( .A1(n5422), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5862) );
  NAND2_X1 U6111 ( .A1(n6402), .A2(n6401), .ZN(n8282) );
  INV_X1 U6112 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n6396) );
  INV_X1 U6113 ( .A(n8630), .ZN(n7975) );
  AOI21_X1 U6114 ( .B1(n5620), .B2(n5868), .A(n5868), .ZN(n5617) );
  NAND2_X1 U6115 ( .A1(n5616), .A2(n5620), .ZN(n6343) );
  INV_X1 U6116 ( .A(n9307), .ZN(n9336) );
  INV_X1 U6117 ( .A(n8099), .ZN(n8153) );
  INV_X1 U6118 ( .A(n7757), .ZN(n7989) );
  AND2_X1 U6119 ( .A1(P2_U3151), .A2(n5598), .ZN(n9621) );
  INV_X1 U6120 ( .A(n10932), .ZN(n7272) );
  INV_X1 U6121 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n5757) );
  XNOR2_X1 U6122 ( .A(n5945), .B(n5944), .ZN(n7050) );
  OAI21_X1 U6123 ( .B1(n6842), .B2(P1_IR_REG_22__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n6843) );
  NAND2_X1 U6124 ( .A1(n6649), .A2(n6648), .ZN(n10646) );
  AND4_X1 U6125 ( .A1(n6677), .A2(n6676), .A3(n6675), .A4(n6674), .ZN(n10569)
         );
  NAND2_X1 U6126 ( .A1(n10132), .A2(n8718), .ZN(n10145) );
  AND4_X1 U6127 ( .A1(n6556), .A2(n6555), .A3(n6554), .A4(n6553), .ZN(n10170)
         );
  NAND2_X1 U6128 ( .A1(n5701), .A2(n10091), .ZN(n10164) );
  NAND2_X1 U6129 ( .A1(n10208), .A2(n8675), .ZN(n5283) );
  AND4_X1 U6130 ( .A1(n6605), .A2(n6604), .A3(n6603), .A4(n6602), .ZN(n10213)
         );
  AND4_X1 U6131 ( .A1(n6669), .A2(n6668), .A3(n6667), .A4(n6666), .ZN(n10237)
         );
  NAND2_X1 U6132 ( .A1(n7239), .A2(n10705), .ZN(n10259) );
  INV_X1 U6133 ( .A(n8654), .ZN(n10289) );
  NAND2_X1 U6134 ( .A1(n6782), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n6457) );
  XNOR2_X1 U6135 ( .A(n6818), .B(P1_IR_REG_28__SCAN_IN), .ZN(n10790) );
  AND2_X1 U6136 ( .A1(n10345), .A2(n5358), .ZN(n7163) );
  NAND2_X1 U6137 ( .A1(n10350), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n5358) );
  INV_X1 U6138 ( .A(n5357), .ZN(n7161) );
  AND2_X1 U6139 ( .A1(n5357), .A2(n5356), .ZN(n7143) );
  NAND2_X1 U6140 ( .A1(n7168), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n5356) );
  NOR2_X1 U6141 ( .A1(n7190), .A2(n7189), .ZN(n7445) );
  NOR2_X1 U6142 ( .A1(n7187), .A2(n5350), .ZN(n7190) );
  AND2_X1 U6143 ( .A1(n7192), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n5350) );
  NOR2_X1 U6144 ( .A1(n10875), .A2(n5352), .ZN(n10803) );
  AND2_X1 U6145 ( .A1(n10880), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n5352) );
  NOR2_X1 U6146 ( .A1(n10803), .A2(n10802), .ZN(n10801) );
  NOR2_X1 U6147 ( .A1(n10801), .A2(n5351), .ZN(n7449) );
  AND2_X1 U6148 ( .A1(n10806), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n5351) );
  INV_X1 U6149 ( .A(n5348), .ZN(n10856) );
  AND2_X1 U6150 ( .A1(n5348), .A2(n5347), .ZN(n10814) );
  NAND2_X1 U6151 ( .A1(n10864), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n5347) );
  INV_X1 U6152 ( .A(n5346), .ZN(n10813) );
  NAND2_X1 U6153 ( .A1(n10402), .A2(n5344), .ZN(n10837) );
  NAND2_X1 U6154 ( .A1(n10380), .A2(n10375), .ZN(n5344) );
  INV_X1 U6155 ( .A(n10870), .ZN(n10841) );
  AND2_X1 U6156 ( .A1(n6983), .A2(n7141), .ZN(n10868) );
  INV_X1 U6157 ( .A(n6825), .ZN(n6826) );
  AOI22_X1 U6158 ( .A1(n10273), .A2(n10999), .B1(n8324), .B2(n10272), .ZN(
        n6825) );
  NAND2_X1 U6159 ( .A1(n6879), .A2(n5736), .ZN(n6787) );
  OR2_X1 U6160 ( .A1(n8807), .A2(n10426), .ZN(n5736) );
  NAND2_X1 U6161 ( .A1(n5300), .A2(n5299), .ZN(n6880) );
  INV_X1 U6162 ( .A(n8957), .ZN(n5299) );
  INV_X1 U6163 ( .A(n5301), .ZN(n5300) );
  NAND2_X1 U6164 ( .A1(n10444), .A2(n8905), .ZN(n10425) );
  NOR2_X1 U6165 ( .A1(n5495), .A2(n5155), .ZN(n10431) );
  INV_X1 U6166 ( .A(n5500), .ZN(n5495) );
  OR2_X1 U6167 ( .A1(n10448), .A2(n10447), .ZN(n10592) );
  NAND2_X1 U6168 ( .A1(n10506), .A2(n6717), .ZN(n10492) );
  NAND2_X1 U6169 ( .A1(n5331), .A2(n5329), .ZN(n10517) );
  OAI21_X1 U6170 ( .B1(n8246), .B2(n5522), .A(n5521), .ZN(n10547) );
  NOR2_X1 U6171 ( .A1(n8245), .A2(n6678), .ZN(n10574) );
  NAND2_X1 U6172 ( .A1(n6672), .A2(n6671), .ZN(n10636) );
  OR2_X1 U6173 ( .A1(n7411), .A2(n6699), .ZN(n6672) );
  NAND2_X1 U6174 ( .A1(n11123), .A2(n6630), .ZN(n8069) );
  NAND2_X1 U6175 ( .A1(n5517), .A2(n5516), .ZN(n7881) );
  NAND2_X1 U6176 ( .A1(n7890), .A2(n10119), .ZN(n5516) );
  OAI21_X1 U6177 ( .B1(n7890), .B2(n10119), .A(n11087), .ZN(n5517) );
  OAI21_X1 U6178 ( .B1(n7709), .B2(n5505), .A(n5503), .ZN(n7866) );
  NAND2_X1 U6179 ( .A1(n7708), .A2(n6557), .ZN(n7868) );
  NAND2_X1 U6180 ( .A1(n5606), .A2(n6549), .ZN(n10101) );
  NAND2_X1 U6181 ( .A1(n9623), .A2(n6546), .ZN(n5606) );
  OR2_X1 U6182 ( .A1(n6495), .A2(n6494), .ZN(n7654) );
  NAND2_X1 U6183 ( .A1(n6889), .A2(n11171), .ZN(n5308) );
  NAND2_X1 U6184 ( .A1(n6697), .A2(n6696), .ZN(n10626) );
  AOI21_X1 U6185 ( .B1(n9611), .B2(n6546), .A(n5727), .ZN(n10416) );
  INV_X1 U6186 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n5341) );
  INV_X1 U6187 ( .A(n10450), .ZN(n10660) );
  INV_X1 U6188 ( .A(n10468), .ZN(n6745) );
  INV_X1 U6189 ( .A(n10626), .ZN(n10676) );
  INV_X1 U6190 ( .A(n8680), .ZN(n11116) );
  AND3_X2 U6191 ( .A1(n6888), .A2(n7209), .A3(n7206), .ZN(n11175) );
  AND2_X1 U6192 ( .A1(n10689), .A2(n10688), .ZN(n10711) );
  INV_X1 U6193 ( .A(n6455), .ZN(n10700) );
  INV_X1 U6194 ( .A(n10790), .ZN(n10705) );
  XNOR2_X1 U6195 ( .A(n6837), .B(n6836), .ZN(n8167) );
  INV_X1 U6196 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n6836) );
  NAND2_X1 U6197 ( .A1(n6151), .A2(n6152), .ZN(n7282) );
  NAND2_X1 U6198 ( .A1(n6131), .A2(n6130), .ZN(n6133) );
  OR2_X1 U6199 ( .A1(n6131), .A2(n6130), .ZN(n6132) );
  NAND2_X1 U6200 ( .A1(n6111), .A2(n5796), .ZN(n6131) );
  NAND2_X1 U6201 ( .A1(n6076), .A2(n5669), .ZN(n5662) );
  NAND2_X1 U6202 ( .A1(n5670), .A2(n5669), .ZN(n6094) );
  NAND2_X1 U6203 ( .A1(n5670), .A2(n5671), .ZN(n6093) );
  XNOR2_X1 U6204 ( .A(n6030), .B(n6029), .ZN(n9623) );
  NAND2_X1 U6205 ( .A1(n6015), .A2(n5779), .ZN(n6030) );
  NAND2_X1 U6206 ( .A1(n6014), .A2(n6015), .ZN(n6971) );
  NAND2_X1 U6207 ( .A1(n5274), .A2(n6465), .ZN(n6503) );
  NAND2_X1 U6208 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5361) );
  NAND2_X1 U6209 ( .A1(n5360), .A2(n10692), .ZN(n5359) );
  NAND2_X1 U6210 ( .A1(n5629), .A2(n9158), .ZN(n5627) );
  OAI21_X1 U6211 ( .B1(n5488), .B2(n10974), .A(n5485), .ZN(P2_U3201) );
  XNOR2_X1 U6212 ( .A(n9341), .B(n5489), .ZN(n5488) );
  AOI21_X1 U6213 ( .B1(n9344), .B2(n10962), .A(n5486), .ZN(n5485) );
  INV_X1 U6214 ( .A(n9342), .ZN(n5489) );
  INV_X1 U6215 ( .A(n6876), .ZN(n6877) );
  OAI21_X1 U6216 ( .B1(n9357), .B2(n9564), .A(n6875), .ZN(n6876) );
  NAND2_X1 U6217 ( .A1(n6435), .A2(n6436), .ZN(n6437) );
  AND2_X1 U6218 ( .A1(n10046), .A2(n5209), .ZN(n5267) );
  XNOR2_X1 U6219 ( .A(n5697), .B(n8813), .ZN(n8821) );
  OR3_X1 U6220 ( .A1(n10852), .A2(n10853), .A3(n5353), .ZN(P1_U3261) );
  NAND2_X1 U6221 ( .A1(n5355), .A2(n5354), .ZN(n5353) );
  AOI222_X1 U6222 ( .A1(n11152), .A2(n11151), .B1(n11150), .B2(n11149), .C1(
        P1_REG2_REG_14__SCAN_IN), .C2(n11011), .ZN(n11159) );
  NOR2_X1 U6223 ( .A1(n5200), .A2(n5340), .ZN(n5339) );
  NAND2_X1 U6224 ( .A1(n6889), .A2(n11175), .ZN(n5342) );
  AND2_X1 U6225 ( .A1(n9459), .A2(n6233), .ZN(n5138) );
  NAND2_X1 U6226 ( .A1(n6719), .A2(n6718), .ZN(n10068) );
  NAND4_X2 U6227 ( .A1(n5910), .A2(n5909), .A3(n5908), .A4(n5907), .ZN(n6908)
         );
  INV_X1 U6228 ( .A(n9432), .ZN(n5413) );
  NAND2_X1 U6229 ( .A1(n6572), .A2(n6571), .ZN(n10080) );
  AND2_X1 U6230 ( .A1(n5497), .A2(n8905), .ZN(n5139) );
  NAND2_X1 U6231 ( .A1(n7289), .A2(n6906), .ZN(n5140) );
  AND2_X1 U6232 ( .A1(n5613), .A2(n9091), .ZN(n9151) );
  OR2_X1 U6233 ( .A1(n10538), .A2(n10551), .ZN(n9030) );
  OR2_X1 U6234 ( .A1(n6482), .A2(n6481), .ZN(n6484) );
  INV_X1 U6235 ( .A(n6814), .ZN(n5277) );
  AND2_X1 U6236 ( .A1(n5679), .A2(n6044), .ZN(n5141) );
  NAND2_X1 U6237 ( .A1(n7682), .A2(n9255), .ZN(n5142) );
  AND4_X1 U6238 ( .A1(n6538), .A2(n6537), .A3(n6536), .A4(n6535), .ZN(n7834)
         );
  INV_X1 U6239 ( .A(n7834), .ZN(n5297) );
  AND2_X1 U6240 ( .A1(n9011), .A2(n8872), .ZN(n5143) );
  AND2_X1 U6241 ( .A1(n5530), .A2(n6374), .ZN(n5144) );
  INV_X1 U6242 ( .A(n5415), .ZN(n5414) );
  OAI21_X1 U6243 ( .B1(n5417), .B2(n5416), .A(n5418), .ZN(n5415) );
  INV_X1 U6244 ( .A(n8403), .ZN(n5640) );
  NOR2_X1 U6245 ( .A1(n11087), .A2(n10119), .ZN(n5515) );
  INV_X1 U6246 ( .A(n6678), .ZN(n5524) );
  AND2_X1 U6247 ( .A1(n10636), .A2(n10283), .ZN(n6678) );
  INV_X1 U6248 ( .A(n5401), .ZN(n5400) );
  NAND2_X1 U6249 ( .A1(n5183), .A2(n5402), .ZN(n5401) );
  NOR2_X1 U6250 ( .A1(n9425), .A2(n9243), .ZN(n5145) );
  NAND2_X1 U6251 ( .A1(n5298), .A2(n5297), .ZN(n6805) );
  OR2_X1 U6252 ( .A1(n8403), .A2(n9173), .ZN(n5146) );
  AND2_X1 U6253 ( .A1(n8521), .A2(n8518), .ZN(n5147) );
  INV_X2 U6254 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3151) );
  INV_X1 U6255 ( .A(P2_RD_REG_SCAN_IN), .ZN(n5287) );
  NAND2_X1 U6256 ( .A1(n10535), .A2(n5425), .ZN(n5148) );
  INV_X1 U6257 ( .A(n9501), .ZN(n5381) );
  INV_X1 U6258 ( .A(n6273), .ZN(n5457) );
  AND2_X1 U6259 ( .A1(n5578), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n5149) );
  INV_X1 U6260 ( .A(n5278), .ZN(n7201) );
  NAND2_X1 U6261 ( .A1(n6796), .A2(n5277), .ZN(n5278) );
  XOR2_X1 U6262 ( .A(n9368), .B(n6905), .Z(n5150) );
  INV_X1 U6263 ( .A(n6580), .ZN(n6652) );
  OR2_X1 U6264 ( .A1(n8270), .A2(n8269), .ZN(n5151) );
  INV_X1 U6265 ( .A(n9453), .ZN(n5417) );
  NOR2_X1 U6266 ( .A1(n6139), .A2(n6119), .ZN(n5153) );
  AND2_X1 U6267 ( .A1(n8319), .A2(n8318), .ZN(n8822) );
  NAND2_X1 U6268 ( .A1(n9170), .A2(n8394), .ZN(n9139) );
  OAI211_X1 U6269 ( .C1(n5966), .C2(n6942), .A(n5441), .B(n5440), .ZN(n6899)
         );
  INV_X1 U6270 ( .A(n7429), .ZN(n7426) );
  XNOR2_X1 U6271 ( .A(n9554), .B(n9494), .ZN(n9483) );
  INV_X1 U6272 ( .A(n9483), .ZN(n5542) );
  XNOR2_X1 U6273 ( .A(n6326), .B(SI_29_), .ZN(n6779) );
  NAND2_X1 U6274 ( .A1(n8486), .A2(n8489), .ZN(n5436) );
  NOR2_X1 U6275 ( .A1(n10442), .A2(n10443), .ZN(n5154) );
  AND2_X1 U6276 ( .A1(n10450), .A2(n10275), .ZN(n5155) );
  OR2_X1 U6277 ( .A1(n10434), .A2(n10446), .ZN(n9040) );
  NAND2_X1 U6278 ( .A1(n9070), .A2(n5871), .ZN(n6353) );
  NAND2_X1 U6279 ( .A1(n5723), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6793) );
  OR2_X1 U6280 ( .A1(n7425), .A2(n5583), .ZN(n5156) );
  NAND2_X1 U6281 ( .A1(n6701), .A2(n6700), .ZN(n10538) );
  NAND2_X1 U6282 ( .A1(n5608), .A2(n9095), .ZN(n9212) );
  NAND4_X1 U6283 ( .A1(n5963), .A2(n5962), .A3(n5961), .A4(n5960), .ZN(n9258)
         );
  INV_X1 U6284 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n5868) );
  AND2_X1 U6285 ( .A1(n10564), .A2(n8920), .ZN(n5157) );
  INV_X1 U6286 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n5870) );
  INV_X1 U6287 ( .A(n6908), .ZN(n5389) );
  AND2_X1 U6288 ( .A1(n8477), .A2(n9246), .ZN(n5158) );
  INV_X1 U6289 ( .A(n9386), .ZN(n5373) );
  OR2_X1 U6290 ( .A1(n11152), .A2(n10190), .ZN(n9012) );
  INV_X1 U6291 ( .A(n9012), .ZN(n5597) );
  NAND2_X1 U6292 ( .A1(n8760), .A2(n8759), .ZN(n10106) );
  AND4_X1 U6293 ( .A1(n5852), .A2(n5851), .A3(n5850), .A4(n6206), .ZN(n5159)
         );
  NAND2_X1 U6294 ( .A1(n5280), .A2(n10153), .ZN(n10124) );
  NAND2_X1 U6295 ( .A1(n9040), .A2(n9044), .ZN(n10430) );
  INV_X1 U6296 ( .A(n10430), .ZN(n5497) );
  AND2_X1 U6297 ( .A1(n5800), .A2(n5799), .ZN(n6130) );
  NAND2_X1 U6298 ( .A1(n5866), .A2(n5865), .ZN(n9105) );
  AND2_X1 U6299 ( .A1(n5466), .A2(n6357), .ZN(n5160) );
  INV_X1 U6300 ( .A(n5669), .ZN(n5668) );
  NOR2_X1 U6301 ( .A1(n6092), .A2(n5672), .ZN(n5669) );
  NAND2_X1 U6302 ( .A1(n6728), .A2(n6727), .ZN(n10603) );
  NAND2_X1 U6303 ( .A1(n6390), .A2(n5859), .ZN(n6399) );
  OR2_X1 U6304 ( .A1(n6646), .A2(n6950), .ZN(n5161) );
  OR2_X1 U6305 ( .A1(n9587), .A2(n9403), .ZN(n5162) );
  NOR2_X1 U6306 ( .A1(n10945), .A2(n9338), .ZN(n5163) );
  AND2_X1 U6307 ( .A1(n7113), .A2(n8781), .ZN(n5164) );
  AND2_X1 U6308 ( .A1(n5609), .A2(n9213), .ZN(n5165) );
  NOR2_X1 U6309 ( .A1(n9285), .A2(n9284), .ZN(n5166) );
  AND2_X1 U6310 ( .A1(n8650), .A2(n5700), .ZN(n5167) );
  NAND4_X1 U6311 ( .A1(n6209), .A2(n6208), .A3(n6207), .A4(n6206), .ZN(n5168)
         );
  AND2_X1 U6312 ( .A1(n9021), .A2(n8884), .ZN(n8952) );
  NAND2_X1 U6313 ( .A1(n6613), .A2(n6612), .ZN(n11152) );
  AND2_X1 U6314 ( .A1(n8670), .A2(n10287), .ZN(n5169) );
  OR2_X1 U6315 ( .A1(n8612), .A2(n8611), .ZN(n5170) );
  INV_X1 U6316 ( .A(n10209), .ZN(n8664) );
  INV_X1 U6317 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n5861) );
  NAND2_X1 U6318 ( .A1(n6561), .A2(n6560), .ZN(n10172) );
  NOR2_X1 U6319 ( .A1(n10172), .A2(n10290), .ZN(n5171) );
  OR2_X1 U6320 ( .A1(n8395), .A2(n5639), .ZN(n5172) );
  INV_X1 U6321 ( .A(n5672), .ZN(n5671) );
  NOR2_X1 U6322 ( .A1(n5790), .A2(SI_11_), .ZN(n5672) );
  INV_X1 U6323 ( .A(n5681), .ZN(n6201) );
  OAI21_X1 U6324 ( .B1(n6150), .B2(n5685), .A(n5682), .ZN(n5681) );
  AND2_X1 U6325 ( .A1(n5303), .A2(n5511), .ZN(n5173) );
  AND2_X1 U6326 ( .A1(n5308), .A2(n5307), .ZN(n5174) );
  NAND2_X1 U6327 ( .A1(n5335), .A2(n5673), .ZN(n5175) );
  OR2_X1 U6328 ( .A1(n8777), .A2(n8776), .ZN(n5176) );
  OR2_X1 U6329 ( .A1(n5783), .A2(SI_9_), .ZN(n5177) );
  OR2_X1 U6330 ( .A1(n10668), .A2(n10515), .ZN(n5178) );
  OR2_X1 U6331 ( .A1(n8670), .A2(n10287), .ZN(n5179) );
  INV_X1 U6332 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n5860) );
  AND3_X1 U6333 ( .A1(n9545), .A2(n9436), .A3(n8618), .ZN(n5180) );
  INV_X1 U6334 ( .A(n5679), .ZN(n5678) );
  NOR2_X1 U6335 ( .A1(n6029), .A2(n5680), .ZN(n5679) );
  INV_X1 U6336 ( .A(n5689), .ZN(n5688) );
  NOR2_X1 U6337 ( .A1(n6166), .A2(n5690), .ZN(n5689) );
  AND2_X1 U6338 ( .A1(n5178), .A2(n5506), .ZN(n5181) );
  AND2_X1 U6339 ( .A1(n5782), .A2(n5781), .ZN(n5182) );
  INV_X1 U6340 ( .A(n9459), .ZN(n9466) );
  AND2_X1 U6341 ( .A1(n8622), .A2(n8621), .ZN(n5183) );
  AND2_X1 U6342 ( .A1(n5137), .A2(n9582), .ZN(n5184) );
  NOR2_X1 U6343 ( .A1(n10680), .A2(n10550), .ZN(n5185) );
  INV_X1 U6344 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n9781) );
  OR2_X1 U6345 ( .A1(n8591), .A2(n8590), .ZN(n5186) );
  OR2_X1 U6346 ( .A1(n9225), .A2(n5636), .ZN(n5187) );
  INV_X1 U6347 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n5858) );
  INV_X1 U6348 ( .A(n7725), .ZN(n7128) );
  AND2_X1 U6349 ( .A1(n8874), .A2(n9005), .ZN(n5188) );
  AND2_X1 U6350 ( .A1(n8440), .A2(n8439), .ZN(n5189) );
  AND2_X1 U6351 ( .A1(n5734), .A2(n5733), .ZN(n5190) );
  OR2_X1 U6352 ( .A1(n5150), .A2(n5630), .ZN(n5191) );
  AND2_X1 U6353 ( .A1(n5563), .A2(n5861), .ZN(n5192) );
  AND2_X1 U6354 ( .A1(n9995), .A2(n9787), .ZN(n5193) );
  OR2_X1 U6355 ( .A1(n8985), .A2(n5600), .ZN(n5194) );
  INV_X1 U6356 ( .A(n8948), .ZN(n5296) );
  NAND2_X1 U6357 ( .A1(n9015), .A2(n8878), .ZN(n8948) );
  AND2_X1 U6358 ( .A1(n5333), .A2(n8832), .ZN(n5195) );
  AND2_X1 U6359 ( .A1(n7113), .A2(n5739), .ZN(n5196) );
  INV_X1 U6360 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n9791) );
  INV_X1 U6361 ( .A(n5513), .ZN(n5512) );
  NAND2_X1 U6362 ( .A1(n5179), .A2(n5514), .ZN(n5513) );
  INV_X1 U6363 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n9999) );
  NAND2_X1 U6364 ( .A1(n8128), .A2(n6373), .ZN(n5532) );
  INV_X1 U6365 ( .A(n9111), .ZN(n5635) );
  INV_X1 U6366 ( .A(n9254), .ZN(n7774) );
  AND2_X1 U6367 ( .A1(n10535), .A2(n5426), .ZN(n5197) );
  OAI21_X1 U6368 ( .B1(n9172), .B2(n5146), .A(n5638), .ZN(n8412) );
  INV_X1 U6369 ( .A(n5444), .ZN(n8102) );
  INV_X1 U6370 ( .A(n8542), .ZN(n5536) );
  AND2_X1 U6371 ( .A1(n5705), .A2(n5704), .ZN(n5198) );
  NAND2_X1 U6372 ( .A1(n6684), .A2(n6683), .ZN(n10579) );
  INV_X1 U6373 ( .A(n10579), .ZN(n10680) );
  NAND2_X1 U6374 ( .A1(n5460), .A2(n5542), .ZN(n9473) );
  NAND2_X1 U6375 ( .A1(n8069), .A2(n8948), .ZN(n8068) );
  NAND2_X1 U6376 ( .A1(n5637), .A2(n8383), .ZN(n9223) );
  AND2_X1 U6377 ( .A1(n8248), .A2(n5596), .ZN(n5199) );
  OR2_X1 U6378 ( .A1(n8378), .A2(n5254), .ZN(n9119) );
  NOR2_X1 U6379 ( .A1(n8807), .A2(n10685), .ZN(n5200) );
  OR2_X1 U6380 ( .A1(n9508), .A2(n9475), .ZN(n8577) );
  NOR2_X1 U6381 ( .A1(n8258), .A2(n8259), .ZN(n5201) );
  INV_X1 U6382 ( .A(n5435), .ZN(n10578) );
  NOR2_X1 U6383 ( .A1(n8251), .A2(n10636), .ZN(n5435) );
  INV_X1 U6384 ( .A(n5453), .ZN(n5452) );
  NOR2_X1 U6385 ( .A1(n6285), .A2(n5454), .ZN(n5453) );
  AND2_X1 U6386 ( .A1(n10480), .A2(n10496), .ZN(n5202) );
  AND2_X1 U6387 ( .A1(n5591), .A2(n5590), .ZN(n5203) );
  INV_X1 U6388 ( .A(n5818), .ZN(n5657) );
  OR2_X1 U6389 ( .A1(n6031), .A2(n5857), .ZN(n5204) );
  NOR2_X1 U6390 ( .A1(n9549), .A2(n9448), .ZN(n5205) );
  NAND2_X1 U6391 ( .A1(n5532), .A2(n5529), .ZN(n5206) );
  OR2_X1 U6392 ( .A1(n5808), .A2(SI_17_), .ZN(n5207) );
  AND2_X1 U6393 ( .A1(n5806), .A2(n9645), .ZN(n5208) );
  INV_X1 U6394 ( .A(n5816), .ZN(n5654) );
  OR2_X1 U6395 ( .A1(n10656), .A2(n10253), .ZN(n5209) );
  OR2_X1 U6396 ( .A1(n8387), .A2(n9232), .ZN(n8564) );
  INV_X1 U6397 ( .A(n8564), .ZN(n5531) );
  INV_X1 U6398 ( .A(n7753), .ZN(n5585) );
  OR2_X1 U6399 ( .A1(n5583), .A2(n5580), .ZN(n5210) );
  INV_X1 U6400 ( .A(n9095), .ZN(n5610) );
  AND2_X1 U6401 ( .A1(n8732), .A2(n10142), .ZN(n5211) );
  NAND2_X1 U6402 ( .A1(n8722), .A2(n10284), .ZN(n5212) );
  AND2_X1 U6403 ( .A1(n5484), .A2(n5151), .ZN(n5213) );
  NAND2_X1 U6404 ( .A1(n7384), .A2(n5643), .ZN(n5642) );
  NAND2_X1 U6405 ( .A1(n7221), .A2(n7220), .ZN(n7219) );
  INV_X1 U6406 ( .A(n9059), .ZN(n7108) );
  NAND2_X1 U6407 ( .A1(n9336), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n5214) );
  INV_X1 U6408 ( .A(n8277), .ZN(n9269) );
  XNOR2_X1 U6409 ( .A(n8112), .B(n8114), .ZN(n8115) );
  OR2_X1 U6410 ( .A1(n8237), .A2(n9248), .ZN(n5215) );
  NAND2_X1 U6411 ( .A1(n5526), .A2(n5525), .ZN(n6428) );
  NOR2_X1 U6412 ( .A1(n7789), .A2(n5586), .ZN(n5216) );
  AND2_X1 U6413 ( .A1(n9011), .A2(n11130), .ZN(n8946) );
  AND2_X1 U6414 ( .A1(n5842), .A2(n5841), .ZN(n5217) );
  OR2_X1 U6415 ( .A1(n8277), .A2(n6141), .ZN(n5218) );
  XNOR2_X1 U6416 ( .A(n5862), .B(n5861), .ZN(n6347) );
  OAI21_X1 U6417 ( .B1(n6971), .B2(n6699), .A(n6541), .ZN(n7639) );
  INV_X1 U6418 ( .A(n7639), .ZN(n5298) );
  NAND4_X1 U6419 ( .A1(n6479), .A2(n6478), .A3(n6477), .A4(n6476), .ZN(n10295)
         );
  INV_X1 U6420 ( .A(n10295), .ZN(n6483) );
  AND2_X1 U6421 ( .A1(n6346), .A2(n6345), .ZN(n9471) );
  INV_X1 U6422 ( .A(n9471), .ZN(n9490) );
  OAI22_X1 U6423 ( .A1(n7815), .A2(n6507), .B1(n11042), .B2(n7646), .ZN(n7412)
         );
  INV_X1 U6424 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n5473) );
  NOR2_X1 U6425 ( .A1(n7072), .A2(n7073), .ZN(n5219) );
  AND2_X1 U6426 ( .A1(n5567), .A2(n5571), .ZN(n5220) );
  NAND2_X1 U6427 ( .A1(n6343), .A2(n6342), .ZN(n8624) );
  INV_X1 U6428 ( .A(n9062), .ZN(n8971) );
  XNOR2_X1 U6430 ( .A(n6842), .B(P1_IR_REG_22__SCAN_IN), .ZN(n6796) );
  XNOR2_X1 U6431 ( .A(n9337), .B(n10940), .ZN(n10946) );
  XNOR2_X1 U6432 ( .A(n9310), .B(n10940), .ZN(n10949) );
  AND2_X1 U6433 ( .A1(n8625), .A2(n5395), .ZN(n5394) );
  INV_X1 U6434 ( .A(n6384), .ZN(n5555) );
  NAND2_X1 U6435 ( .A1(n5551), .A2(n5554), .ZN(n5550) );
  NAND3_X1 U6436 ( .A1(n8914), .A2(n5249), .A3(n5247), .ZN(n5246) );
  NAND3_X1 U6437 ( .A1(n8909), .A2(n10458), .A3(n8980), .ZN(n5248) );
  INV_X1 U6438 ( .A(n5864), .ZN(n5649) );
  MUX2_X1 U6439 ( .A(n5747), .B(n5953), .S(n5864), .Z(n5748) );
  NAND3_X1 U6440 ( .A1(n5287), .A2(P1_ADDR_REG_19__SCAN_IN), .A3(
        P2_ADDR_REG_19__SCAN_IN), .ZN(n5250) );
  NAND3_X1 U6441 ( .A1(n5289), .A2(n5290), .A3(n5288), .ZN(n5251) );
  NAND2_X1 U6442 ( .A1(n8378), .A2(n8380), .ZN(n5253) );
  INV_X1 U6443 ( .A(n6910), .ZN(n5263) );
  AND2_X2 U6444 ( .A1(n5420), .A2(n5526), .ZN(n6390) );
  NAND2_X1 U6445 ( .A1(n5268), .A2(n5267), .ZN(P1_U3214) );
  NAND2_X1 U6446 ( .A1(n5269), .A2(n10244), .ZN(n5268) );
  NAND2_X1 U6447 ( .A1(n5271), .A2(n5270), .ZN(n5269) );
  NAND2_X1 U6448 ( .A1(n10243), .A2(n8804), .ZN(n5270) );
  NAND2_X1 U6449 ( .A1(n5273), .A2(n5272), .ZN(n5271) );
  INV_X1 U6450 ( .A(n10042), .ZN(n5272) );
  NAND2_X1 U6451 ( .A1(n10243), .A2(n10043), .ZN(n5273) );
  NAND2_X1 U6452 ( .A1(n5698), .A2(n8650), .ZN(n8657) );
  INV_X1 U6453 ( .A(n8641), .ZN(n5279) );
  NAND2_X1 U6454 ( .A1(n8641), .A2(n8642), .ZN(n10090) );
  NAND2_X1 U6455 ( .A1(n5282), .A2(n10142), .ZN(n8735) );
  AND2_X1 U6456 ( .A1(n6644), .A2(n5286), .ZN(n6670) );
  NAND2_X1 U6457 ( .A1(n6644), .A2(n5285), .ZN(n5284) );
  NAND3_X1 U6458 ( .A1(n6628), .A2(n11118), .A3(n8948), .ZN(n5293) );
  NAND2_X1 U6459 ( .A1(n5293), .A2(n5294), .ZN(n8216) );
  NOR2_X1 U6460 ( .A1(n5513), .A2(n5306), .ZN(n5305) );
  NAND2_X1 U6461 ( .A1(n6860), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n5307) );
  NAND3_X1 U6462 ( .A1(n8946), .A2(n5599), .A3(n5194), .ZN(n11129) );
  NAND2_X1 U6463 ( .A1(n6076), .A2(n5317), .ZN(n5320) );
  OAI21_X1 U6464 ( .B1(n6076), .B2(n5665), .A(n5663), .ZN(n6111) );
  NAND3_X1 U6465 ( .A1(n5663), .A2(n5665), .A3(n6130), .ZN(n5319) );
  NAND2_X1 U6466 ( .A1(n10549), .A2(n5195), .ZN(n5328) );
  NAND2_X1 U6467 ( .A1(n5335), .A2(n5334), .ZN(n6065) );
  NAND2_X1 U6468 ( .A1(n5342), .A2(n5339), .ZN(P1_U3518) );
  NOR2_X1 U6469 ( .A1(n11175), .A2(n5341), .ZN(n5340) );
  MUX2_X1 U6470 ( .A(n10991), .B(P1_REG1_REG_1__SCAN_IN), .S(n7144), .Z(n10304) );
  NAND3_X1 U6471 ( .A1(n5365), .A2(n8515), .A3(n8518), .ZN(n5364) );
  NAND3_X1 U6472 ( .A1(n5385), .A2(n5384), .A3(n5379), .ZN(n5378) );
  OAI211_X1 U6473 ( .C1(n6893), .C2(n7259), .A(n5917), .B(n5918), .ZN(n7223)
         );
  NAND4_X2 U6474 ( .A1(n5390), .A2(n5392), .A3(n5391), .A4(n5952), .ZN(n9260)
         );
  AND2_X1 U6475 ( .A1(n9260), .A2(n7215), .ZN(n8491) );
  NAND2_X1 U6476 ( .A1(n5393), .A2(n5394), .ZN(n8626) );
  NAND2_X1 U6477 ( .A1(n8620), .A2(n5396), .ZN(n5393) );
  NAND2_X1 U6478 ( .A1(n5405), .A2(n5406), .ZN(n8595) );
  NAND2_X1 U6479 ( .A1(n8586), .A2(n5408), .ZN(n5405) );
  NOR2_X1 U6480 ( .A1(n5180), .A2(n5419), .ZN(n5418) );
  NAND3_X1 U6481 ( .A1(n5526), .A2(n5420), .A3(n5563), .ZN(n5422) );
  NAND2_X1 U6482 ( .A1(n5702), .A2(n5704), .ZN(n6643) );
  NAND4_X1 U6483 ( .A1(n5702), .A2(n5190), .A3(n6447), .A4(n5704), .ZN(n6451)
         );
  NAND2_X1 U6484 ( .A1(n10535), .A2(n5423), .ZN(n10477) );
  NAND3_X1 U6485 ( .A1(n7725), .A2(n11013), .A3(n5427), .ZN(n7816) );
  INV_X1 U6486 ( .A(n6467), .ZN(n5428) );
  NAND2_X1 U6487 ( .A1(n7883), .A2(n11116), .ZN(n11124) );
  NAND2_X1 U6488 ( .A1(n5436), .A2(n5527), .ZN(n5528) );
  INV_X1 U6489 ( .A(n5436), .ZN(n7300) );
  NAND2_X1 U6490 ( .A1(n5438), .A2(n5964), .ZN(n5926) );
  NAND2_X1 U6491 ( .A1(n5438), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n7051) );
  NAND2_X1 U6492 ( .A1(n5438), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n7042) );
  INV_X1 U6493 ( .A(n5438), .ZN(n5437) );
  NAND3_X1 U6494 ( .A1(n5438), .A2(n5848), .A3(n5623), .ZN(n5622) );
  NAND3_X1 U6495 ( .A1(n5847), .A2(n5438), .A3(n5848), .ZN(n5988) );
  NAND2_X2 U6496 ( .A1(n6893), .A2(n8306), .ZN(n5972) );
  NAND2_X2 U6497 ( .A1(n6893), .A2(n5598), .ZN(n5966) );
  NAND2_X2 U6498 ( .A1(n6348), .A2(n6347), .ZN(n6893) );
  NAND2_X1 U6499 ( .A1(n5442), .A2(n5443), .ZN(n8125) );
  NAND3_X1 U6500 ( .A1(n6129), .A2(n8558), .A3(n5446), .ZN(n5442) );
  NAND2_X1 U6501 ( .A1(n6129), .A2(n6128), .ZN(n8040) );
  AOI21_X1 U6502 ( .B1(n6129), .B2(n5446), .A(n5445), .ZN(n5444) );
  INV_X1 U6503 ( .A(n6128), .ZN(n5447) );
  INV_X1 U6504 ( .A(n9472), .ZN(n5460) );
  NAND2_X1 U6505 ( .A1(n9472), .A2(n5138), .ZN(n5458) );
  XNOR2_X1 U6506 ( .A(n6335), .B(n5467), .ZN(n5461) );
  AND2_X1 U6507 ( .A1(n5466), .A2(n5464), .ZN(n6878) );
  NAND2_X1 U6508 ( .A1(n5466), .A2(n5462), .ZN(n6434) );
  NOR2_X2 U6509 ( .A1(n6388), .A2(n5465), .ZN(n5464) );
  INV_X1 U6510 ( .A(n6385), .ZN(n5467) );
  NAND2_X1 U6511 ( .A1(n5476), .A2(n5475), .ZN(n8356) );
  INV_X1 U6512 ( .A(n5484), .ZN(n8271) );
  NAND2_X1 U6513 ( .A1(n6810), .A2(n8983), .ZN(n10549) );
  AOI211_X2 U6514 ( .C1(n10589), .C2(n11168), .A(n10588), .B(n10587), .ZN(
        n10653) );
  NAND2_X1 U6515 ( .A1(n8065), .A2(n8878), .ZN(n8223) );
  NAND2_X1 U6516 ( .A1(n8575), .A2(n8570), .ZN(n8573) );
  AOI22_X1 U6517 ( .A1(n8535), .A2(n8541), .B1(n8588), .B2(n8534), .ZN(n8544)
         );
  INV_X1 U6518 ( .A(n6513), .ZN(n5704) );
  NAND2_X1 U6519 ( .A1(n7709), .A2(n5503), .ZN(n5501) );
  INV_X1 U6520 ( .A(n10476), .ZN(n6736) );
  NAND3_X1 U6521 ( .A1(n5521), .A2(n10546), .A3(n5522), .ZN(n5520) );
  NAND3_X1 U6522 ( .A1(n8486), .A2(n8489), .A3(n7296), .ZN(n7297) );
  NAND2_X1 U6523 ( .A1(n7850), .A2(n5534), .ZN(n5533) );
  NAND2_X1 U6524 ( .A1(n5533), .A2(n5535), .ZN(n7955) );
  NAND2_X1 U6525 ( .A1(n9502), .A2(n8577), .ZN(n5543) );
  NAND2_X1 U6526 ( .A1(n9381), .A2(n5548), .ZN(n5544) );
  NAND2_X1 U6527 ( .A1(n5544), .A2(n5545), .ZN(n8474) );
  NAND2_X1 U6528 ( .A1(n9381), .A2(n5556), .ZN(n5547) );
  AOI21_X1 U6529 ( .B1(n9381), .B2(n8608), .A(n8610), .ZN(n9369) );
  OR2_X1 U6530 ( .A1(n8424), .A2(n5550), .ZN(n5549) );
  NAND2_X1 U6531 ( .A1(n5559), .A2(n5147), .ZN(n7563) );
  NAND2_X1 U6532 ( .A1(n5559), .A2(n8518), .ZN(n7565) );
  NAND2_X1 U6533 ( .A1(n5561), .A2(n5560), .ZN(n6380) );
  AND2_X2 U6534 ( .A1(n6390), .A2(n5192), .ZN(n5869) );
  INV_X1 U6535 ( .A(n7055), .ZN(n5570) );
  OAI21_X2 U6536 ( .B1(n9283), .B2(n5573), .A(n5572), .ZN(n9310) );
  NAND2_X1 U6537 ( .A1(n7425), .A2(n5580), .ZN(n5579) );
  NAND2_X1 U6538 ( .A1(n5579), .A2(n5576), .ZN(n7427) );
  AND2_X1 U6539 ( .A1(n5577), .A2(n5578), .ZN(n5576) );
  INV_X1 U6540 ( .A(n7430), .ZN(n5580) );
  INV_X1 U6541 ( .A(n5582), .ZN(n7591) );
  OAI22_X1 U6542 ( .A1(n7753), .A2(n5587), .B1(n7790), .B2(n5584), .ZN(n7988)
         );
  NAND2_X1 U6543 ( .A1(n8080), .A2(n5592), .ZN(n5588) );
  NAND2_X1 U6544 ( .A1(n8259), .A2(n5595), .ZN(n5593) );
  NAND2_X2 U6545 ( .A1(n5598), .A2(P1_U3086), .ZN(n10704) );
  MUX2_X1 U6546 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(P2_DATAO_REG_4__SCAN_IN), 
        .S(n5755), .Z(n5763) );
  MUX2_X1 U6547 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(P2_DATAO_REG_5__SCAN_IN), 
        .S(n5755), .Z(n5767) );
  MUX2_X1 U6548 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .S(n5755), .Z(n5771) );
  MUX2_X1 U6549 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(P2_DATAO_REG_8__SCAN_IN), 
        .S(n5755), .Z(n5780) );
  MUX2_X1 U6550 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .S(n5755), .Z(n5776) );
  MUX2_X1 U6551 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(P2_DATAO_REG_9__SCAN_IN), 
        .S(n5755), .Z(n5783) );
  MUX2_X1 U6552 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(P2_DATAO_REG_11__SCAN_IN), 
        .S(n5598), .Z(n5790) );
  MUX2_X1 U6553 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(P2_DATAO_REG_12__SCAN_IN), 
        .S(n5598), .Z(n5791) );
  MUX2_X1 U6554 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(P2_DATAO_REG_10__SCAN_IN), 
        .S(n5598), .Z(n5784) );
  MUX2_X1 U6555 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(P2_DATAO_REG_13__SCAN_IN), 
        .S(n5598), .Z(n5793) );
  MUX2_X1 U6556 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(P2_DATAO_REG_14__SCAN_IN), 
        .S(n5598), .Z(n5797) );
  MUX2_X1 U6557 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(P2_DATAO_REG_15__SCAN_IN), 
        .S(n5598), .Z(n5801) );
  MUX2_X1 U6558 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(P2_DATAO_REG_16__SCAN_IN), 
        .S(n5598), .Z(n5805) );
  MUX2_X1 U6559 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(P2_DATAO_REG_17__SCAN_IN), 
        .S(n5598), .Z(n5808) );
  MUX2_X1 U6560 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(P2_DATAO_REG_19__SCAN_IN), 
        .S(n5598), .Z(n5814) );
  MUX2_X1 U6561 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .S(n5598), .Z(n5809) );
  MUX2_X1 U6562 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(P2_DATAO_REG_20__SCAN_IN), 
        .S(n5598), .Z(n5817) );
  MUX2_X1 U6563 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(P2_DATAO_REG_21__SCAN_IN), 
        .S(n5598), .Z(n5819) );
  MUX2_X1 U6564 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(P2_DATAO_REG_22__SCAN_IN), 
        .S(n5598), .Z(n5824) );
  MUX2_X1 U6565 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(P2_DATAO_REG_23__SCAN_IN), 
        .S(n5598), .Z(n5828) );
  MUX2_X1 U6566 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(P2_DATAO_REG_25__SCAN_IN), 
        .S(n5598), .Z(n5835) );
  MUX2_X1 U6567 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(P2_DATAO_REG_26__SCAN_IN), 
        .S(n5598), .Z(n5840) );
  MUX2_X1 U6568 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(P2_DATAO_REG_24__SCAN_IN), 
        .S(n5598), .Z(n5833) );
  MUX2_X1 U6569 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(P2_DATAO_REG_27__SCAN_IN), 
        .S(n5598), .Z(n5843) );
  MUX2_X1 U6570 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(P2_DATAO_REG_28__SCAN_IN), 
        .S(n5598), .Z(n6321) );
  NAND2_X1 U6571 ( .A1(n7891), .A2(n5188), .ZN(n5599) );
  INV_X1 U6572 ( .A(n8946), .ZN(n5601) );
  NAND3_X1 U6573 ( .A1(n9181), .A2(n9093), .A3(n9095), .ZN(n5607) );
  OAI21_X1 U6574 ( .B1(n5615), .B2(n7064), .A(n5614), .ZN(n7221) );
  NAND2_X1 U6575 ( .A1(n6337), .A2(n6336), .ZN(n5619) );
  OR2_X1 U6576 ( .A1(n6337), .A2(n5868), .ZN(n5616) );
  NAND2_X1 U6577 ( .A1(n6337), .A2(n5620), .ZN(n5618) );
  NAND2_X1 U6578 ( .A1(n9110), .A2(n5626), .ZN(n5625) );
  OAI211_X1 U6579 ( .C1(n9110), .C2(n5627), .A(n5625), .B(n9106), .ZN(P2_U3160) );
  NAND2_X1 U6580 ( .A1(n6050), .A2(n5646), .ZN(n6223) );
  NAND2_X1 U6581 ( .A1(n5649), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n5742) );
  NAND2_X1 U6582 ( .A1(n5649), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n5751) );
  NAND2_X1 U6583 ( .A1(n6204), .A2(n5813), .ZN(n6222) );
  NAND2_X1 U6584 ( .A1(n6244), .A2(n5822), .ZN(n6248) );
  OAI21_X1 U6585 ( .B1(n6298), .B2(n5659), .A(n5658), .ZN(n5884) );
  NAND2_X1 U6586 ( .A1(n6298), .A2(n5838), .ZN(n6302) );
  NAND2_X1 U6587 ( .A1(n5884), .A2(n5883), .ZN(n5846) );
  NAND2_X1 U6588 ( .A1(n5662), .A2(n5666), .ZN(n6109) );
  NAND2_X1 U6589 ( .A1(n6150), .A2(n6149), .ZN(n6152) );
  NAND2_X1 U6590 ( .A1(n5196), .A2(n5691), .ZN(n7229) );
  NAND2_X1 U6591 ( .A1(n7344), .A2(n7128), .ZN(n5691) );
  NAND2_X1 U6592 ( .A1(n7229), .A2(n7228), .ZN(n5693) );
  NAND2_X1 U6593 ( .A1(n5693), .A2(n5692), .ZN(n7236) );
  NAND2_X1 U6594 ( .A1(n10242), .A2(n8797), .ZN(n10243) );
  NOR2_X1 U6595 ( .A1(n6513), .A2(n6443), .ZN(n6593) );
  NAND2_X1 U6596 ( .A1(n10134), .A2(n8718), .ZN(n5706) );
  OAI21_X1 U6597 ( .B1(n8760), .B2(n5711), .A(n5710), .ZN(n10152) );
  AOI21_X1 U6598 ( .B1(n5710), .B2(n5711), .A(n10155), .ZN(n5709) );
  NAND2_X1 U6599 ( .A1(n8665), .A2(n5717), .ZN(n5716) );
  INV_X1 U6600 ( .A(n8675), .ZN(n5719) );
  NAND2_X1 U6601 ( .A1(n8665), .A2(n8664), .ZN(n10212) );
  NAND2_X1 U6602 ( .A1(n6657), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5720) );
  NAND2_X1 U6603 ( .A1(n5720), .A2(n5721), .ZN(n6795) );
  NAND2_X1 U6604 ( .A1(n7313), .A2(n8446), .ZN(n7314) );
  AND2_X1 U6605 ( .A1(n10968), .A2(n10967), .ZN(n10971) );
  XNOR2_X1 U6606 ( .A(n9281), .B(n9298), .ZN(n9262) );
  NAND2_X1 U6607 ( .A1(n6449), .A2(n6448), .ZN(n10693) );
  NAND2_X1 U6608 ( .A1(n6880), .A2(n6879), .ZN(n8351) );
  NAND2_X1 U6609 ( .A1(n7783), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n7782) );
  AND2_X1 U6610 ( .A1(n11123), .A2(n11122), .ZN(n11157) );
  XNOR2_X1 U6611 ( .A(n9085), .B(n9086), .ZN(n9133) );
  OAI21_X1 U6612 ( .B1(n10966), .B2(n10971), .A(n10970), .ZN(n10983) );
  OR2_X1 U6613 ( .A1(n7101), .A2(n5972), .ZN(n6116) );
  NAND2_X2 U6614 ( .A1(n8036), .A2(n6367), .ZN(n8128) );
  INV_X1 U6615 ( .A(n6896), .ZN(n6897) );
  OAI21_X2 U6616 ( .B1(n9415), .B2(n6382), .A(n6381), .ZN(n9399) );
  INV_X1 U6617 ( .A(n6831), .ZN(n6835) );
  NAND2_X1 U6618 ( .A1(n6831), .A2(n6460), .ZN(n6816) );
  NAND2_X1 U6619 ( .A1(n5132), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n6456) );
  INV_X1 U6620 ( .A(n6451), .ZN(n6449) );
  NAND2_X1 U6621 ( .A1(n6451), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6452) );
  INV_X1 U6622 ( .A(n6670), .ZN(n6658) );
  NAND2_X1 U6623 ( .A1(n10949), .A2(n9317), .ZN(n10950) );
  NAND2_X1 U6624 ( .A1(n6815), .A2(n7111), .ZN(n10566) );
  XNOR2_X1 U6625 ( .A(n9072), .B(n10416), .ZN(n8320) );
  OAI21_X1 U6626 ( .B1(n8974), .B2(n8973), .A(n7122), .ZN(n8975) );
  XNOR2_X1 U6627 ( .A(n6793), .B(n9796), .ZN(n6813) );
  INV_X1 U6628 ( .A(n10152), .ZN(n10157) );
  NOR2_X2 U6629 ( .A1(n9260), .A2(n7215), .ZN(n7296) );
  NAND2_X1 U6630 ( .A1(n9070), .A2(n8332), .ZN(n5958) );
  INV_X1 U6631 ( .A(n9070), .ZN(n5872) );
  AND2_X1 U6632 ( .A1(n8317), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(n5727) );
  NAND2_X1 U6633 ( .A1(n10603), .A2(n10277), .ZN(n5728) );
  INV_X1 U6634 ( .A(n8462), .ZN(n6374) );
  AND2_X1 U6635 ( .A1(n7929), .A2(n7936), .ZN(n5729) );
  NOR2_X1 U6636 ( .A1(n6090), .A2(n7961), .ZN(n5730) );
  AND4_X1 U6637 ( .A1(n8471), .A2(n5189), .A3(n8470), .A4(n8623), .ZN(n5732)
         );
  AND4_X1 U6638 ( .A1(n6789), .A2(n6444), .A3(n9999), .A4(n10004), .ZN(n5733)
         );
  AND3_X1 U6639 ( .A1(n5193), .A2(n9791), .A3(n6679), .ZN(n5734) );
  OR2_X1 U6640 ( .A1(n6462), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5735) );
  OR2_X1 U6641 ( .A1(n8807), .A2(n10644), .ZN(n5737) );
  NAND2_X1 U6642 ( .A1(n7399), .A2(n7396), .ZN(n5738) );
  INV_X1 U6643 ( .A(n9493), .ZN(n9164) );
  AND4_X1 U6644 ( .A1(n6706), .A2(n6705), .A3(n6704), .A4(n6703), .ZN(n10551)
         );
  AND4_X1 U6645 ( .A1(n6641), .A2(n6640), .A3(n6639), .A4(n6638), .ZN(n11136)
         );
  AND4_X1 U6646 ( .A1(n6611), .A2(n6610), .A3(n6609), .A4(n6608), .ZN(n11138)
         );
  INV_X1 U6647 ( .A(n9105), .ZN(n9582) );
  AND4_X1 U6648 ( .A1(n6716), .A2(n6715), .A3(n6714), .A4(n6713), .ZN(n10531)
         );
  AND4_X1 U6649 ( .A1(n6619), .A2(n6618), .A3(n6617), .A4(n6616), .ZN(n10190)
         );
  INV_X1 U6650 ( .A(n10190), .ZN(n6629) );
  INV_X1 U6651 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n6405) );
  INV_X1 U6652 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n5752) );
  AND4_X1 U6653 ( .A1(n6744), .A2(n6743), .A3(n6742), .A4(n6741), .ZN(n10484)
         );
  INV_X1 U6654 ( .A(n9607), .ZN(n6436) );
  INV_X1 U6655 ( .A(n11178), .ZN(n6432) );
  OR2_X1 U6656 ( .A1(n7333), .A2(n10789), .ZN(n5739) );
  NAND2_X1 U6657 ( .A1(n7090), .A2(n11104), .ZN(n9500) );
  INV_X1 U6658 ( .A(n8521), .ZN(n7566) );
  NAND2_X2 U6659 ( .A1(n7210), .A2(n10580), .ZN(n10560) );
  INV_X2 U6660 ( .A(n10560), .ZN(n11011) );
  NAND2_X1 U6661 ( .A1(n8037), .A2(n6368), .ZN(n5740) );
  INV_X1 U6662 ( .A(n8479), .ZN(n6366) );
  INV_X1 U6663 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n10004) );
  INV_X1 U6664 ( .A(n8624), .ZN(n8472) );
  AND2_X1 U6665 ( .A1(n8775), .A2(n10060), .ZN(n8776) );
  OR2_X1 U6666 ( .A1(n7827), .A2(n8933), .ZN(n7525) );
  NAND2_X1 U6667 ( .A1(n9133), .A2(n9435), .ZN(n9181) );
  NAND2_X1 U6668 ( .A1(n8362), .A2(n8363), .ZN(n8364) );
  INV_X1 U6669 ( .A(n9390), .ZN(n9362) );
  INV_X1 U6670 ( .A(n6290), .ZN(n5875) );
  NAND2_X1 U6671 ( .A1(n9105), .A2(n5137), .ZN(n6317) );
  AOI21_X1 U6672 ( .B1(n7950), .B2(n6091), .A(n5730), .ZN(n8169) );
  INV_X1 U6673 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n6336) );
  INV_X1 U6674 ( .A(n6665), .ZN(n6662) );
  INV_X1 U6675 ( .A(n8734), .ZN(n8732) );
  INV_X1 U6676 ( .A(n10538), .ZN(n6707) );
  INV_X1 U6677 ( .A(SI_19_), .ZN(n9841) );
  INV_X1 U6678 ( .A(SI_15_), .ZN(n9846) );
  INV_X1 U6679 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n9772) );
  INV_X1 U6680 ( .A(n9173), .ZN(n8391) );
  AND2_X1 U6681 ( .A1(n6423), .A2(n6896), .ZN(n6921) );
  INV_X1 U6682 ( .A(n8364), .ZN(n8365) );
  NOR2_X1 U6683 ( .A1(n9300), .A2(n9299), .ZN(n9303) );
  NOR2_X1 U6684 ( .A1(n9363), .A2(n9476), .ZN(n9364) );
  NAND2_X1 U6685 ( .A1(n5875), .A2(n5874), .ZN(n6307) );
  INV_X1 U6686 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n9914) );
  NOR2_X1 U6687 ( .A1(n6021), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n6036) );
  INV_X1 U6688 ( .A(n10105), .ZN(n8759) );
  NOR2_X1 U6689 ( .A1(n6606), .A2(n10188), .ZN(n6614) );
  NAND2_X1 U6690 ( .A1(n6712), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n6720) );
  NAND2_X1 U6691 ( .A1(n7350), .A2(n7349), .ZN(n7353) );
  INV_X1 U6692 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n6521) );
  NOR2_X1 U6693 ( .A1(n8966), .A2(n6812), .ZN(n8963) );
  NAND2_X1 U6694 ( .A1(n10468), .A2(n10276), .ZN(n6747) );
  INV_X1 U6695 ( .A(n6730), .ZN(n6731) );
  NOR2_X1 U6696 ( .A1(n6673), .A2(n10232), .ZN(n6685) );
  INV_X1 U6697 ( .A(n8952), .ZN(n8179) );
  AND2_X1 U6698 ( .A1(n8864), .A2(n8865), .ZN(n8945) );
  OR2_X1 U6699 ( .A1(n6551), .A2(n6550), .ZN(n6562) );
  AND2_X1 U6700 ( .A1(n6812), .A2(n6813), .ZN(n7107) );
  OAI21_X1 U6701 ( .B1(n8316), .B2(n8315), .A(n8305), .ZN(n8312) );
  OR2_X1 U6702 ( .A1(P1_IR_REG_18__SCAN_IN), .A2(P1_IR_REG_19__SCAN_IN), .ZN(
        n6788) );
  INV_X1 U6703 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n9701) );
  AND2_X1 U6704 ( .A1(n9347), .A2(n5878), .ZN(n9370) );
  INV_X1 U6705 ( .A(n5959), .ZN(n6305) );
  INV_X1 U6706 ( .A(n9620), .ZN(n7758) );
  XNOR2_X1 U6707 ( .A(n8091), .B(n8078), .ZN(n7978) );
  INV_X1 U6708 ( .A(n9377), .ZN(n9403) );
  NAND2_X1 U6709 ( .A1(n6157), .A2(n9228), .ZN(n6175) );
  NAND2_X1 U6710 ( .A1(n8618), .A2(n6864), .ZN(n7083) );
  INV_X1 U6711 ( .A(n8558), .ZN(n8106) );
  INV_X1 U6712 ( .A(n9250), .ZN(n8003) );
  NAND2_X1 U6713 ( .A1(n6387), .A2(n7091), .ZN(n7968) );
  INV_X1 U6714 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n6338) );
  NAND2_X1 U6715 ( .A1(n6651), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n6665) );
  AND2_X1 U6716 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n6508) );
  NOR2_X1 U6717 ( .A1(n6691), .A2(n10178), .ZN(n6702) );
  INV_X1 U6718 ( .A(n10261), .ZN(n10236) );
  INV_X1 U6719 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n10167) );
  INV_X1 U6720 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n10188) );
  INV_X1 U6721 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n10232) );
  NAND2_X1 U6722 ( .A1(n6751), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n6770) );
  NAND2_X1 U6723 ( .A1(n10267), .A2(n10286), .ZN(n6642) );
  NAND2_X1 U6724 ( .A1(n6814), .A2(n7122), .ZN(n7111) );
  OR2_X1 U6725 ( .A1(n11011), .A2(n7533), .ZN(n11014) );
  INV_X1 U6726 ( .A(n6474), .ZN(n6529) );
  INV_X1 U6727 ( .A(n11135), .ZN(n11002) );
  INV_X1 U6728 ( .A(n7545), .ZN(n7557) );
  OR2_X1 U6729 ( .A1(n6798), .A2(n7202), .ZN(n7711) );
  AOI21_X1 U6730 ( .B1(n6287), .B2(n6286), .A(n5834), .ZN(n6298) );
  AND2_X1 U6731 ( .A1(n5804), .A2(n5803), .ZN(n6149) );
  INV_X1 U6732 ( .A(n5967), .ZN(n5969) );
  OR2_X1 U6733 ( .A1(n6935), .A2(n6931), .ZN(n9231) );
  OR2_X1 U6734 ( .A1(n5135), .A2(n9347), .ZN(n8432) );
  OR2_X1 U6735 ( .A1(n5135), .A2(n9114), .ZN(n5892) );
  OR2_X1 U6736 ( .A1(n6353), .A2(n5955), .ZN(n5963) );
  INV_X1 U6737 ( .A(n6893), .ZN(n7009) );
  INV_X1 U6738 ( .A(n10974), .ZN(n10928) );
  INV_X1 U6739 ( .A(n10969), .ZN(n10970) );
  OR2_X1 U6740 ( .A1(n9565), .A2(n6389), .ZN(n11105) );
  AND2_X1 U6741 ( .A1(n8519), .A2(n8518), .ZN(n8450) );
  AOI21_X1 U6742 ( .B1(n7082), .B2(n7083), .A(n7086), .ZN(n6874) );
  NAND2_X1 U6743 ( .A1(n7968), .A2(n8057), .ZN(n9541) );
  INV_X1 U6744 ( .A(n9565), .ZN(n9553) );
  NAND2_X1 U6745 ( .A1(n7012), .A2(n6947), .ZN(n7089) );
  NAND2_X1 U6746 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_31__SCAN_IN), .ZN(
        n5945) );
  INV_X1 U6747 ( .A(n10263), .ZN(n10250) );
  NAND2_X1 U6748 ( .A1(n6813), .A2(n7110), .ZN(n9059) );
  AND4_X1 U6749 ( .A1(n6777), .A2(n6776), .A3(n6775), .A4(n6774), .ZN(n10426)
         );
  AND4_X1 U6750 ( .A1(n6689), .A2(n6688), .A3(n6687), .A4(n6686), .ZN(n10550)
         );
  OR2_X1 U6751 ( .A1(n10796), .A2(n10310), .ZN(n10870) );
  NOR2_X1 U6752 ( .A1(n10796), .A2(n8291), .ZN(n10838) );
  INV_X1 U6753 ( .A(n8955), .ZN(n10483) );
  INV_X1 U6754 ( .A(n10563), .ZN(n10575) );
  INV_X1 U6755 ( .A(n11153), .ZN(n11018) );
  INV_X1 U6756 ( .A(n10580), .ZN(n11149) );
  INV_X1 U6757 ( .A(n11168), .ZN(n10649) );
  NAND2_X1 U6758 ( .A1(n7711), .A2(n7799), .ZN(n11168) );
  INV_X1 U6759 ( .A(n7799), .ZN(n11144) );
  OAI21_X1 U6760 ( .B1(n10688), .B2(P1_D_REG_0__SCAN_IN), .A(n10691), .ZN(
        n7206) );
  OR3_X1 U6761 ( .A1(n8135), .A2(n8282), .A3(n6406), .ZN(n7012) );
  AND2_X1 U6762 ( .A1(n6927), .A2(n6926), .ZN(n9217) );
  NAND2_X1 U6763 ( .A1(n6916), .A2(n9609), .ZN(n9224) );
  INV_X1 U6764 ( .A(n9219), .ZN(n9238) );
  INV_X1 U6765 ( .A(n9435), .ZN(n9243) );
  INV_X1 U6766 ( .A(n8174), .ZN(n9249) );
  INV_X1 U6767 ( .A(n8117), .ZN(n9251) );
  OR2_X1 U6768 ( .A1(n7010), .A2(n7009), .ZN(n10976) );
  AND2_X1 U6769 ( .A1(n9497), .A2(n9496), .ZN(n9559) );
  INV_X1 U6770 ( .A(n9443), .ZN(n9505) );
  OR3_X1 U6771 ( .A1(n9565), .A2(n7089), .A3(n6895), .ZN(n11104) );
  OR2_X1 U6772 ( .A1(n9572), .A2(n9565), .ZN(n9564) );
  INV_X1 U6773 ( .A(n9572), .ZN(n9561) );
  INV_X1 U6774 ( .A(n9220), .ZN(n9587) );
  AND2_X2 U6775 ( .A1(n6430), .A2(n9609), .ZN(n11178) );
  INV_X1 U6776 ( .A(n7089), .ZN(n9609) );
  INV_X1 U6777 ( .A(n9327), .ZN(n9334) );
  INV_X1 U6778 ( .A(n9622), .ZN(n9109) );
  XNOR2_X1 U6779 ( .A(n6843), .B(n10008), .ZN(n9061) );
  NAND2_X1 U6780 ( .A1(n7335), .A2(P1_STATE_REG_SCAN_IN), .ZN(n10263) );
  INV_X1 U6781 ( .A(n10266), .ZN(n10253) );
  AND4_X1 U6782 ( .A1(n6786), .A2(n6785), .A3(n6784), .A4(n6783), .ZN(n8816)
         );
  INV_X1 U6783 ( .A(n10550), .ZN(n10282) );
  INV_X1 U6784 ( .A(n11138), .ZN(n11115) );
  INV_X1 U6785 ( .A(n10170), .ZN(n10291) );
  INV_X1 U6786 ( .A(n10868), .ZN(n10885) );
  NAND2_X1 U6787 ( .A1(n8320), .A2(n11126), .ZN(n10419) );
  AND2_X1 U6788 ( .A1(n7896), .A2(n7895), .ZN(n11091) );
  OR2_X1 U6789 ( .A1(n11011), .A2(n7552), .ZN(n10563) );
  NAND2_X1 U6790 ( .A1(n11171), .A2(n10985), .ZN(n10644) );
  AND3_X2 U6791 ( .A1(n6888), .A2(n7209), .A3(n7120), .ZN(n11171) );
  INV_X1 U6792 ( .A(n10068), .ZN(n10668) );
  INV_X1 U6793 ( .A(n8722), .ZN(n10686) );
  INV_X1 U6794 ( .A(n11175), .ZN(n11172) );
  INV_X1 U6795 ( .A(n10711), .ZN(n10712) );
  INV_X1 U6796 ( .A(n10828), .ZN(n10385) );
  NOR2_X1 U6797 ( .A1(n7012), .A2(n6891), .ZN(P2_U3893) );
  OAI21_X1 U6798 ( .B1(n6878), .B2(n9572), .A(n6877), .ZN(P2_U3488) );
  AND2_X2 U6799 ( .A1(n9061), .A2(n6890), .ZN(P1_U3973) );
  NAND2_X1 U6800 ( .A1(n5742), .A2(n5741), .ZN(n5745) );
  INV_X1 U6801 ( .A(n5745), .ZN(n5744) );
  INV_X1 U6802 ( .A(SI_1_), .ZN(n5743) );
  NAND2_X1 U6803 ( .A1(n5744), .A2(n5743), .ZN(n5746) );
  NAND2_X1 U6804 ( .A1(n5745), .A2(SI_1_), .ZN(n5750) );
  NAND2_X1 U6805 ( .A1(n5746), .A2(n5750), .ZN(n5948) );
  INV_X1 U6806 ( .A(n5948), .ZN(n5749) );
  INV_X1 U6807 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n5747) );
  INV_X1 U6808 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n5953) );
  INV_X1 U6809 ( .A(SI_0_), .ZN(n6472) );
  NAND2_X1 U6810 ( .A1(n5950), .A2(n5750), .ZN(n5967) );
  INV_X1 U6811 ( .A(n5968), .ZN(n5753) );
  NAND2_X1 U6812 ( .A1(n5967), .A2(n5753), .ZN(n5970) );
  NAND2_X1 U6813 ( .A1(n5970), .A2(n5754), .ZN(n5914) );
  NAND2_X1 U6814 ( .A1(n5758), .A2(SI_3_), .ZN(n5762) );
  INV_X1 U6815 ( .A(n5758), .ZN(n5760) );
  INV_X1 U6816 ( .A(SI_3_), .ZN(n5759) );
  NAND2_X1 U6817 ( .A1(n5760), .A2(n5759), .ZN(n5761) );
  AND2_X1 U6818 ( .A1(n5762), .A2(n5761), .ZN(n5913) );
  NAND2_X1 U6819 ( .A1(n5914), .A2(n5913), .ZN(n5916) );
  NAND2_X1 U6820 ( .A1(n5916), .A2(n5762), .ZN(n5933) );
  NAND2_X1 U6821 ( .A1(n5763), .A2(SI_4_), .ZN(n5766) );
  INV_X1 U6822 ( .A(n5763), .ZN(n5764) );
  INV_X1 U6823 ( .A(SI_4_), .ZN(n9667) );
  NAND2_X1 U6824 ( .A1(n5764), .A2(n9667), .ZN(n5765) );
  AND2_X1 U6825 ( .A1(n5766), .A2(n5765), .ZN(n5932) );
  NAND2_X1 U6826 ( .A1(n5933), .A2(n5932), .ZN(n5935) );
  NAND2_X1 U6827 ( .A1(n5935), .A2(n5766), .ZN(n5985) );
  NAND2_X1 U6828 ( .A1(n5767), .A2(SI_5_), .ZN(n5770) );
  INV_X1 U6829 ( .A(n5767), .ZN(n5768) );
  INV_X1 U6830 ( .A(SI_5_), .ZN(n9868) );
  NAND2_X1 U6831 ( .A1(n5768), .A2(n9868), .ZN(n5769) );
  AND2_X1 U6832 ( .A1(n5770), .A2(n5769), .ZN(n5984) );
  NAND2_X1 U6833 ( .A1(n5985), .A2(n5984), .ZN(n5987) );
  NAND2_X1 U6834 ( .A1(n5771), .A2(SI_6_), .ZN(n5775) );
  INV_X1 U6835 ( .A(n5771), .ZN(n5773) );
  INV_X1 U6836 ( .A(SI_6_), .ZN(n5772) );
  NAND2_X1 U6837 ( .A1(n5773), .A2(n5772), .ZN(n5774) );
  AND2_X1 U6838 ( .A1(n5775), .A2(n5774), .ZN(n5997) );
  NAND2_X1 U6839 ( .A1(n5776), .A2(SI_7_), .ZN(n5779) );
  INV_X1 U6840 ( .A(n5776), .ZN(n5777) );
  INV_X1 U6841 ( .A(SI_7_), .ZN(n9662) );
  NAND2_X1 U6842 ( .A1(n5777), .A2(n9662), .ZN(n5778) );
  XNOR2_X1 U6843 ( .A(n5780), .B(SI_8_), .ZN(n6029) );
  INV_X1 U6844 ( .A(n5780), .ZN(n5782) );
  INV_X1 U6845 ( .A(SI_8_), .ZN(n5781) );
  XNOR2_X1 U6846 ( .A(n5783), .B(n9860), .ZN(n6044) );
  NAND2_X1 U6847 ( .A1(n5784), .A2(SI_10_), .ZN(n5789) );
  INV_X1 U6848 ( .A(n5784), .ZN(n5786) );
  INV_X1 U6849 ( .A(SI_10_), .ZN(n5785) );
  NAND2_X1 U6850 ( .A1(n5786), .A2(n5785), .ZN(n5787) );
  NAND2_X1 U6851 ( .A1(n5789), .A2(n5787), .ZN(n6063) );
  INV_X1 U6852 ( .A(n6063), .ZN(n5788) );
  NAND2_X1 U6853 ( .A1(n6065), .A2(n5789), .ZN(n6076) );
  XNOR2_X1 U6854 ( .A(n5790), .B(SI_11_), .ZN(n6075) );
  NAND2_X1 U6855 ( .A1(n5791), .A2(SI_12_), .ZN(n5792) );
  OAI21_X1 U6856 ( .B1(n5791), .B2(SI_12_), .A(n5792), .ZN(n6092) );
  NAND2_X1 U6857 ( .A1(n5793), .A2(SI_13_), .ZN(n5796) );
  INV_X1 U6858 ( .A(n5793), .ZN(n5794) );
  INV_X1 U6859 ( .A(SI_13_), .ZN(n9652) );
  NAND2_X1 U6860 ( .A1(n5794), .A2(n9652), .ZN(n5795) );
  NAND2_X1 U6861 ( .A1(n5797), .A2(SI_14_), .ZN(n5800) );
  INV_X1 U6862 ( .A(n5797), .ZN(n5798) );
  NAND2_X1 U6863 ( .A1(n5798), .A2(n9853), .ZN(n5799) );
  NAND2_X1 U6864 ( .A1(n5801), .A2(SI_15_), .ZN(n5804) );
  INV_X1 U6865 ( .A(n5801), .ZN(n5802) );
  NAND2_X1 U6866 ( .A1(n5802), .A2(n9846), .ZN(n5803) );
  XNOR2_X1 U6867 ( .A(n5805), .B(SI_16_), .ZN(n6166) );
  INV_X1 U6868 ( .A(n5805), .ZN(n5806) );
  NAND2_X1 U6869 ( .A1(n5809), .A2(SI_18_), .ZN(n5813) );
  INV_X1 U6870 ( .A(n5809), .ZN(n5810) );
  NAND2_X1 U6871 ( .A1(n5810), .A2(n9845), .ZN(n5811) );
  NAND2_X1 U6872 ( .A1(n5813), .A2(n5811), .ZN(n6202) );
  INV_X1 U6873 ( .A(n6202), .ZN(n5812) );
  NAND2_X1 U6874 ( .A1(n6201), .A2(n5812), .ZN(n6204) );
  XNOR2_X1 U6875 ( .A(n5814), .B(SI_19_), .ZN(n6221) );
  INV_X1 U6876 ( .A(n5814), .ZN(n5815) );
  NAND2_X1 U6877 ( .A1(n5815), .A2(n9841), .ZN(n5816) );
  XNOR2_X1 U6878 ( .A(n5817), .B(n9641), .ZN(n6234) );
  NOR2_X1 U6879 ( .A1(n5817), .A2(SI_20_), .ZN(n5818) );
  NAND2_X1 U6880 ( .A1(n5819), .A2(SI_21_), .ZN(n5823) );
  INV_X1 U6881 ( .A(n5819), .ZN(n5820) );
  INV_X1 U6882 ( .A(SI_21_), .ZN(n9634) );
  NAND2_X1 U6883 ( .A1(n5820), .A2(n9634), .ZN(n5821) );
  NAND2_X1 U6884 ( .A1(n5823), .A2(n5821), .ZN(n6245) );
  INV_X1 U6885 ( .A(n6245), .ZN(n5822) );
  NAND2_X1 U6886 ( .A1(n6248), .A2(n5823), .ZN(n6262) );
  NAND2_X1 U6887 ( .A1(n5824), .A2(SI_22_), .ZN(n5827) );
  INV_X1 U6888 ( .A(n5824), .ZN(n5825) );
  INV_X1 U6889 ( .A(SI_22_), .ZN(n9834) );
  NAND2_X1 U6890 ( .A1(n5825), .A2(n9834), .ZN(n5826) );
  NAND2_X1 U6891 ( .A1(n6262), .A2(n6261), .ZN(n6264) );
  NAND2_X1 U6892 ( .A1(n6264), .A2(n5827), .ZN(n6276) );
  XNOR2_X1 U6893 ( .A(n5828), .B(SI_23_), .ZN(n6275) );
  INV_X1 U6894 ( .A(n5828), .ZN(n5830) );
  INV_X1 U6895 ( .A(SI_23_), .ZN(n5829) );
  NAND2_X1 U6896 ( .A1(n5830), .A2(n5829), .ZN(n5831) );
  INV_X1 U6897 ( .A(SI_24_), .ZN(n5832) );
  XNOR2_X1 U6898 ( .A(n5833), .B(n5832), .ZN(n6286) );
  NOR2_X1 U6899 ( .A1(n5833), .A2(SI_24_), .ZN(n5834) );
  NAND2_X1 U6900 ( .A1(n5835), .A2(SI_25_), .ZN(n5839) );
  INV_X1 U6901 ( .A(n5835), .ZN(n5836) );
  INV_X1 U6902 ( .A(SI_25_), .ZN(n9830) );
  NAND2_X1 U6903 ( .A1(n5836), .A2(n9830), .ZN(n5837) );
  NAND2_X1 U6904 ( .A1(n5839), .A2(n5837), .ZN(n6299) );
  INV_X1 U6905 ( .A(n6299), .ZN(n5838) );
  XNOR2_X1 U6906 ( .A(n5840), .B(SI_26_), .ZN(n5901) );
  INV_X1 U6907 ( .A(n5840), .ZN(n5842) );
  INV_X1 U6908 ( .A(SI_26_), .ZN(n5841) );
  XNOR2_X1 U6909 ( .A(n5843), .B(n9825), .ZN(n5883) );
  INV_X1 U6910 ( .A(n5843), .ZN(n5844) );
  NAND2_X1 U6911 ( .A1(n5844), .A2(n9825), .ZN(n5845) );
  NAND2_X1 U6912 ( .A1(n5846), .A2(n5845), .ZN(n6320) );
  INV_X1 U6913 ( .A(SI_28_), .ZN(n6322) );
  NOR2_X1 U6914 ( .A1(P2_IR_REG_8__SCAN_IN), .A2(P2_IR_REG_7__SCAN_IN), .ZN(
        n5852) );
  NOR2_X1 U6915 ( .A1(P2_IR_REG_10__SCAN_IN), .A2(P2_IR_REG_14__SCAN_IN), .ZN(
        n5856) );
  NAND2_X1 U6916 ( .A1(n5159), .A2(n5130), .ZN(n5857) );
  XNOR2_X2 U6917 ( .A(n5863), .B(n5860), .ZN(n6348) );
  NAND2_X1 U6918 ( .A1(n8293), .A2(n8421), .ZN(n5866) );
  INV_X1 U6919 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n8294) );
  OR2_X1 U6920 ( .A1(n5966), .A2(n8294), .ZN(n5865) );
  NAND2_X1 U6921 ( .A1(n5869), .A2(n5870), .ZN(n9612) );
  XNOR2_X2 U6922 ( .A(n5867), .B(n9613), .ZN(n9070) );
  NAND2_X2 U6923 ( .A1(n5872), .A2(n8332), .ZN(n5959) );
  NAND2_X1 U6924 ( .A1(n6305), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n5882) );
  INV_X1 U6925 ( .A(n6353), .ZN(n6329) );
  INV_X1 U6926 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n9517) );
  OR2_X1 U6927 ( .A1(n8428), .A2(n9517), .ZN(n5881) );
  INV_X1 U6928 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n9205) );
  NAND2_X1 U6929 ( .A1(n5978), .A2(n9701), .ZN(n6004) );
  NAND2_X1 U6930 ( .A1(n6056), .A2(n6055), .ZN(n6069) );
  NAND2_X1 U6931 ( .A1(n9205), .A2(n6192), .ZN(n6227) );
  NAND2_X1 U6932 ( .A1(n5873), .A2(n9914), .ZN(n6252) );
  INV_X1 U6933 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n9919) );
  INV_X1 U6934 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n5874) );
  INV_X1 U6935 ( .A(n6309), .ZN(n5876) );
  INV_X1 U6936 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n9926) );
  NAND2_X1 U6937 ( .A1(n5876), .A2(n9926), .ZN(n5896) );
  INV_X1 U6938 ( .A(n5889), .ZN(n5877) );
  INV_X1 U6939 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n9888) );
  NAND2_X1 U6940 ( .A1(n5877), .A2(n9888), .ZN(n9347) );
  NAND2_X1 U6941 ( .A1(n5889), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n5878) );
  OR2_X1 U6942 ( .A1(n5135), .A2(n9370), .ZN(n5880) );
  INV_X2 U6943 ( .A(n5958), .ZN(n5951) );
  INV_X1 U6944 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n9580) );
  OR2_X1 U6945 ( .A1(n6330), .A2(n9580), .ZN(n5879) );
  NAND4_X1 U6946 ( .A1(n5882), .A2(n5881), .A3(n5880), .A4(n5879), .ZN(n9378)
         );
  XNOR2_X1 U6947 ( .A(n5884), .B(n5883), .ZN(n8289) );
  NAND2_X1 U6948 ( .A1(n8289), .A2(n8421), .ZN(n5886) );
  INV_X1 U6949 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n8290) );
  OR2_X1 U6950 ( .A1(n5966), .A2(n8290), .ZN(n5885) );
  NAND2_X1 U6951 ( .A1(n6329), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n5894) );
  INV_X1 U6952 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n5887) );
  OR2_X1 U6953 ( .A1(n6330), .A2(n5887), .ZN(n5893) );
  NAND2_X1 U6954 ( .A1(n5896), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n5888) );
  AND2_X1 U6955 ( .A1(n5889), .A2(n5888), .ZN(n9114) );
  INV_X1 U6956 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n5890) );
  OR2_X1 U6957 ( .A1(n5959), .A2(n5890), .ZN(n5891) );
  NAND4_X1 U6958 ( .A1(n5894), .A2(n5893), .A3(n5892), .A4(n5891), .ZN(n9390)
         );
  NAND2_X1 U6959 ( .A1(n6305), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n5900) );
  INV_X1 U6960 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n9526) );
  OR2_X1 U6961 ( .A1(n8428), .A2(n9526), .ZN(n5899) );
  NAND2_X1 U6962 ( .A1(n6309), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n5895) );
  AND2_X1 U6963 ( .A1(n5896), .A2(n5895), .ZN(n9394) );
  OR2_X1 U6964 ( .A1(n5135), .A2(n9394), .ZN(n5898) );
  INV_X1 U6965 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n9585) );
  OR2_X1 U6966 ( .A1(n6330), .A2(n9585), .ZN(n5897) );
  NAND4_X1 U6967 ( .A1(n5900), .A2(n5899), .A3(n5898), .A4(n5897), .ZN(n9377)
         );
  XNOR2_X1 U6968 ( .A(n5902), .B(n5901), .ZN(n8280) );
  NAND2_X1 U6969 ( .A1(n8280), .A2(n8421), .ZN(n5904) );
  INV_X1 U6970 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n8284) );
  OR2_X1 U6971 ( .A1(n5966), .A2(n8284), .ZN(n5903) );
  NAND2_X1 U6972 ( .A1(n5951), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n5910) );
  INV_X1 U6973 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n5905) );
  OR2_X1 U6974 ( .A1(n6353), .A2(n5905), .ZN(n5909) );
  INV_X1 U6975 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n5906) );
  OR2_X1 U6976 ( .A1(n5959), .A2(n5906), .ZN(n5907) );
  NAND2_X1 U6977 ( .A1(n5926), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5912) );
  INV_X1 U6978 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n5911) );
  XNOR2_X1 U6979 ( .A(n5912), .B(n5911), .ZN(n7259) );
  OR2_X1 U6980 ( .A1(n5914), .A2(n5913), .ZN(n5915) );
  NAND2_X1 U6981 ( .A1(n5916), .A2(n5915), .ZN(n6944) );
  OR2_X1 U6982 ( .A1(n5972), .A2(n6944), .ZN(n5917) );
  NAND2_X1 U6983 ( .A1(n6908), .A2(n7223), .ZN(n7399) );
  INV_X1 U6984 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n5919) );
  INV_X1 U6985 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n7585) );
  OR2_X1 U6986 ( .A1(n5959), .A2(n7585), .ZN(n5924) );
  AND2_X1 U6987 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n5920) );
  NOR2_X1 U6988 ( .A1(n5978), .A2(n5920), .ZN(n7322) );
  OR2_X1 U6989 ( .A1(n5956), .A2(n7322), .ZN(n5923) );
  INV_X1 U6990 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n5921) );
  OR2_X1 U6991 ( .A1(n5958), .A2(n5921), .ZN(n5922) );
  NAND2_X1 U6992 ( .A1(n5928), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5927) );
  MUX2_X1 U6993 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5927), .S(
        P2_IR_REG_4__SCAN_IN), .Z(n5931) );
  INV_X1 U6994 ( .A(n5928), .ZN(n5930) );
  INV_X1 U6995 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n5929) );
  NAND2_X1 U6996 ( .A1(n5930), .A2(n5929), .ZN(n5989) );
  NAND2_X1 U6997 ( .A1(n5931), .A2(n5989), .ZN(n7268) );
  OR2_X1 U6998 ( .A1(n5933), .A2(n5932), .ZN(n5934) );
  NAND2_X1 U6999 ( .A1(n5935), .A2(n5934), .ZN(n6953) );
  OR2_X1 U7000 ( .A1(n6953), .A2(n5972), .ZN(n5937) );
  INV_X1 U7001 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n6945) );
  OR2_X1 U7002 ( .A1(n5966), .A2(n6945), .ZN(n5936) );
  OAI211_X1 U7003 ( .C1(n6893), .C2(n7268), .A(n5937), .B(n5936), .ZN(n7587)
         );
  INV_X1 U7004 ( .A(n7587), .ZN(n7403) );
  NAND2_X1 U7005 ( .A1(n7478), .A2(n7403), .ZN(n7395) );
  INV_X1 U7006 ( .A(n7395), .ZN(n5938) );
  NAND2_X1 U7007 ( .A1(n5738), .A2(n7395), .ZN(n5977) );
  NOR2_X1 U7008 ( .A1(n6908), .A2(n7223), .ZN(n7397) );
  NOR2_X1 U7009 ( .A1(n5938), .A2(n7397), .ZN(n5975) );
  INV_X1 U7010 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n10891) );
  OR2_X1 U7011 ( .A1(n5959), .A2(n10891), .ZN(n5943) );
  INV_X1 U7012 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n10902) );
  OR2_X1 U7013 ( .A1(n5956), .A2(n10902), .ZN(n5942) );
  INV_X1 U7014 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n5939) );
  NAND2_X1 U7015 ( .A1(n5951), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n5940) );
  AND4_X2 U7016 ( .A1(n5943), .A2(n5942), .A3(n5941), .A4(n5940), .ZN(n7317)
         );
  INV_X1 U7017 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n5944) );
  INV_X1 U7018 ( .A(n5946), .ZN(n5947) );
  NAND2_X1 U7019 ( .A1(n5948), .A2(n5947), .ZN(n5949) );
  NAND2_X1 U7020 ( .A1(n5950), .A2(n5949), .ZN(n6949) );
  INV_X1 U7021 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n6942) );
  INV_X1 U7022 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n7016) );
  INV_X1 U7023 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n7095) );
  NAND2_X1 U7024 ( .A1(n5951), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n5952) );
  INV_X1 U7025 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n7048) );
  NAND2_X1 U7026 ( .A1(n8306), .A2(SI_0_), .ZN(n5954) );
  XNOR2_X1 U7027 ( .A(n5954), .B(n5953), .ZN(n10040) );
  MUX2_X1 U7028 ( .A(n7048), .B(n10040), .S(n6893), .Z(n7215) );
  INV_X1 U7029 ( .A(n7215), .ZN(n7097) );
  AND2_X1 U7030 ( .A1(n9260), .A2(n7097), .ZN(n7299) );
  INV_X1 U7031 ( .A(n7317), .ZN(n9259) );
  INV_X1 U7032 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n5955) );
  INV_X1 U7033 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n8354) );
  OR2_X1 U7034 ( .A1(n5956), .A2(n8354), .ZN(n5962) );
  INV_X1 U7035 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n5957) );
  OR2_X1 U7036 ( .A1(n5958), .A2(n5957), .ZN(n5961) );
  OR2_X1 U7037 ( .A1(n5959), .A2(n11029), .ZN(n5960) );
  OR2_X1 U7038 ( .A1(n5966), .A2(n5752), .ZN(n5974) );
  NAND2_X1 U7039 ( .A1(n5969), .A2(n5968), .ZN(n5971) );
  NAND2_X1 U7040 ( .A1(n5971), .A2(n5970), .ZN(n8374) );
  OR2_X1 U7041 ( .A1(n5972), .A2(n8374), .ZN(n5973) );
  OAI211_X1 U7042 ( .C1(n6893), .C2(n8375), .A(n5974), .B(n5973), .ZN(n7074)
         );
  INV_X1 U7043 ( .A(n7074), .ZN(n11024) );
  OR2_X2 U7044 ( .A1(n9258), .A2(n11024), .ZN(n8495) );
  NAND2_X1 U7045 ( .A1(n9258), .A2(n11024), .ZN(n8496) );
  NAND2_X2 U7046 ( .A1(n8495), .A2(n8496), .ZN(n8501) );
  NAND2_X1 U7047 ( .A1(n7315), .A2(n8501), .ZN(n7286) );
  INV_X1 U7048 ( .A(n9258), .ZN(n7289) );
  NAND2_X1 U7049 ( .A1(n7289), .A2(n11024), .ZN(n7285) );
  NAND3_X1 U7050 ( .A1(n5975), .A2(n7286), .A3(n7285), .ZN(n5976) );
  NAND2_X1 U7051 ( .A1(n5977), .A2(n5976), .ZN(n7475) );
  NAND2_X1 U7052 ( .A1(n5951), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n5983) );
  INV_X1 U7053 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n7262) );
  OR2_X1 U7054 ( .A1(n8428), .A2(n7262), .ZN(n5982) );
  OR2_X1 U7055 ( .A1(n5978), .A2(n9701), .ZN(n5979) );
  AND2_X1 U7056 ( .A1(n6004), .A2(n5979), .ZN(n7577) );
  OR2_X1 U7057 ( .A1(n5135), .A2(n7577), .ZN(n5981) );
  INV_X1 U7058 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n7576) );
  OR2_X1 U7059 ( .A1(n5959), .A2(n7576), .ZN(n5980) );
  NAND4_X1 U7060 ( .A1(n5983), .A2(n5982), .A3(n5981), .A4(n5980), .ZN(n9256)
         );
  INV_X1 U7061 ( .A(n9256), .ZN(n7513) );
  OR2_X1 U7062 ( .A1(n5985), .A2(n5984), .ZN(n5986) );
  NAND2_X1 U7063 ( .A1(n5987), .A2(n5986), .ZN(n6956) );
  OR2_X1 U7064 ( .A1(n6956), .A2(n5972), .ZN(n5993) );
  NAND2_X1 U7065 ( .A1(n5989), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5990) );
  MUX2_X1 U7066 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5990), .S(
        P2_IR_REG_5__SCAN_IN), .Z(n5991) );
  AND2_X1 U7067 ( .A1(n5988), .A2(n5991), .ZN(n10932) );
  AOI22_X1 U7068 ( .A1(n6224), .A2(P1_DATAO_REG_5__SCAN_IN), .B1(n7009), .B2(
        n10932), .ZN(n5992) );
  NAND2_X1 U7069 ( .A1(n5993), .A2(n5992), .ZN(n7579) );
  INV_X1 U7070 ( .A(n7579), .ZN(n6358) );
  NAND2_X1 U7071 ( .A1(n7513), .A2(n6358), .ZN(n5994) );
  NAND2_X1 U7072 ( .A1(n7475), .A2(n5994), .ZN(n5996) );
  NAND2_X1 U7073 ( .A1(n9256), .A2(n7579), .ZN(n5995) );
  NAND2_X1 U7074 ( .A1(n5996), .A2(n5995), .ZN(n7511) );
  OR2_X1 U7075 ( .A1(n5998), .A2(n5997), .ZN(n5999) );
  NAND2_X1 U7076 ( .A1(n6000), .A2(n5999), .ZN(n6959) );
  OR2_X1 U7077 ( .A1(n6959), .A2(n5972), .ZN(n6003) );
  NAND2_X1 U7078 ( .A1(n5988), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6001) );
  XNOR2_X1 U7079 ( .A(n6001), .B(P2_IR_REG_6__SCAN_IN), .ZN(n7429) );
  AOI22_X1 U7080 ( .A1(n6224), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n7009), .B2(
        n7429), .ZN(n6002) );
  NAND2_X1 U7081 ( .A1(n6003), .A2(n6002), .ZN(n7673) );
  NAND2_X1 U7082 ( .A1(n6329), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n6010) );
  INV_X1 U7083 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n7515) );
  OR2_X1 U7084 ( .A1(n5959), .A2(n7515), .ZN(n6009) );
  NAND2_X1 U7085 ( .A1(n6004), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n6005) );
  AND2_X1 U7086 ( .A1(n6021), .A2(n6005), .ZN(n7516) );
  OR2_X1 U7087 ( .A1(n5135), .A2(n7516), .ZN(n6008) );
  INV_X1 U7088 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n6006) );
  OR2_X1 U7089 ( .A1(n6330), .A2(n6006), .ZN(n6007) );
  NAND4_X1 U7090 ( .A1(n6010), .A2(n6009), .A3(n6008), .A4(n6007), .ZN(n9255)
         );
  AND2_X1 U7091 ( .A1(n7673), .A2(n9255), .ZN(n6011) );
  OAI22_X1 U7092 ( .A1(n7511), .A2(n6011), .B1(n9255), .B2(n7673), .ZN(n7567)
         );
  OR2_X1 U7093 ( .A1(n6013), .A2(n6012), .ZN(n6014) );
  OR2_X1 U7094 ( .A1(n6971), .A2(n5972), .ZN(n6018) );
  NAND2_X1 U7095 ( .A1(n6031), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6016) );
  XNOR2_X1 U7096 ( .A(n6016), .B(P2_IR_REG_7__SCAN_IN), .ZN(n7430) );
  AOI22_X1 U7097 ( .A1(n6224), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n7009), .B2(
        n7430), .ZN(n6017) );
  NAND2_X1 U7098 ( .A1(n6018), .A2(n6017), .ZN(n7684) );
  NAND2_X1 U7099 ( .A1(n5951), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n6026) );
  INV_X1 U7100 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n6019) );
  OR2_X1 U7101 ( .A1(n8428), .A2(n6019), .ZN(n6025) );
  INV_X1 U7102 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n6020) );
  OR2_X1 U7103 ( .A1(n5959), .A2(n6020), .ZN(n6024) );
  AND2_X1 U7104 ( .A1(n6021), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n6022) );
  NOR2_X1 U7105 ( .A1(n6036), .A2(n6022), .ZN(n7690) );
  OR2_X1 U7106 ( .A1(n5135), .A2(n7690), .ZN(n6023) );
  NAND4_X1 U7107 ( .A1(n6026), .A2(n6025), .A3(n6024), .A4(n6023), .ZN(n9254)
         );
  OR2_X1 U7108 ( .A1(n7684), .A2(n7774), .ZN(n7661) );
  NAND2_X1 U7109 ( .A1(n7684), .A2(n7774), .ZN(n8529) );
  NAND2_X1 U7110 ( .A1(n7567), .A2(n7566), .ZN(n6028) );
  OR2_X1 U7111 ( .A1(n7684), .A2(n9254), .ZN(n6027) );
  NAND2_X1 U7112 ( .A1(n6028), .A2(n6027), .ZN(n7663) );
  NAND2_X1 U7113 ( .A1(n9623), .A2(n8421), .ZN(n6034) );
  OR2_X1 U7114 ( .A1(n6047), .A2(n5868), .ZN(n6032) );
  XNOR2_X1 U7115 ( .A(n6032), .B(P2_IR_REG_8__SCAN_IN), .ZN(n9620) );
  AOI22_X1 U7116 ( .A1(n6224), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n7009), .B2(
        n9620), .ZN(n6033) );
  NAND2_X1 U7117 ( .A1(n6034), .A2(n6033), .ZN(n7946) );
  NAND2_X1 U7118 ( .A1(n6329), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n6041) );
  INV_X1 U7119 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n6035) );
  OR2_X1 U7120 ( .A1(n6330), .A2(n6035), .ZN(n6040) );
  NOR2_X1 U7121 ( .A1(n6036), .A2(n9896), .ZN(n6037) );
  OR2_X1 U7122 ( .A1(n6056), .A2(n6037), .ZN(n7667) );
  INV_X1 U7123 ( .A(n7667), .ZN(n7778) );
  OR2_X1 U7124 ( .A1(n5135), .A2(n7778), .ZN(n6039) );
  INV_X1 U7125 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n7666) );
  OR2_X1 U7126 ( .A1(n5959), .A2(n7666), .ZN(n6038) );
  NAND4_X1 U7127 ( .A1(n6041), .A2(n6040), .A3(n6039), .A4(n6038), .ZN(n9253)
         );
  NOR2_X1 U7128 ( .A1(n7946), .A2(n7936), .ZN(n8526) );
  INV_X1 U7129 ( .A(n8526), .ZN(n6360) );
  NAND2_X1 U7130 ( .A1(n7946), .A2(n7936), .ZN(n8528) );
  NAND2_X1 U7131 ( .A1(n6360), .A2(n8528), .ZN(n8453) );
  NAND2_X1 U7132 ( .A1(n7663), .A2(n8453), .ZN(n6043) );
  OR2_X1 U7133 ( .A1(n7946), .A2(n9253), .ZN(n6042) );
  NAND2_X1 U7134 ( .A1(n6043), .A2(n6042), .ZN(n7852) );
  XNOR2_X1 U7135 ( .A(n6045), .B(n6044), .ZN(n6984) );
  NAND2_X1 U7136 ( .A1(n6984), .A2(n8421), .ZN(n6053) );
  NOR2_X1 U7137 ( .A1(n6050), .A2(n5868), .ZN(n6048) );
  MUX2_X1 U7138 ( .A(n5868), .B(n6048), .S(P2_IR_REG_9__SCAN_IN), .Z(n6051) );
  NOR2_X1 U7139 ( .A1(n6051), .A2(n6078), .ZN(n7761) );
  AOI22_X1 U7140 ( .A1(n6224), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n7009), .B2(
        n7761), .ZN(n6052) );
  NAND2_X1 U7141 ( .A1(n6053), .A2(n6052), .ZN(n7932) );
  NAND2_X1 U7142 ( .A1(n5951), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n6062) );
  INV_X1 U7143 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n6054) );
  OR2_X1 U7144 ( .A1(n8428), .A2(n6054), .ZN(n6061) );
  OR2_X1 U7145 ( .A1(n6056), .A2(n6055), .ZN(n6057) );
  AND2_X1 U7146 ( .A1(n6069), .A2(n6057), .ZN(n7937) );
  OR2_X1 U7147 ( .A1(n5135), .A2(n7937), .ZN(n6060) );
  INV_X1 U7148 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n6058) );
  OR2_X1 U7149 ( .A1(n5959), .A2(n6058), .ZN(n6059) );
  NAND4_X1 U7150 ( .A1(n6062), .A2(n6061), .A3(n6060), .A4(n6059), .ZN(n9252)
         );
  NOR2_X1 U7151 ( .A1(n7932), .A2(n8050), .ZN(n8539) );
  INV_X1 U7152 ( .A(n8539), .ZN(n6363) );
  NAND2_X1 U7153 ( .A1(n7932), .A2(n8050), .ZN(n8532) );
  NAND2_X1 U7154 ( .A1(n6363), .A2(n8532), .ZN(n7851) );
  NAND2_X1 U7155 ( .A1(n7852), .A2(n7851), .ZN(n7950) );
  OR2_X1 U7156 ( .A1(n7932), .A2(n9252), .ZN(n7949) );
  NAND2_X1 U7157 ( .A1(n5175), .A2(n6063), .ZN(n6064) );
  NAND2_X1 U7158 ( .A1(n6065), .A2(n6064), .ZN(n6990) );
  OR2_X1 U7159 ( .A1(n6990), .A2(n5972), .ZN(n6068) );
  OR2_X1 U7160 ( .A1(n6078), .A2(n5868), .ZN(n6066) );
  XNOR2_X1 U7161 ( .A(n6066), .B(P2_IR_REG_10__SCAN_IN), .ZN(n7757) );
  AOI22_X1 U7162 ( .A1(n6224), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n7009), .B2(
        n7757), .ZN(n6067) );
  NAND2_X1 U7163 ( .A1(n6068), .A2(n6067), .ZN(n8061) );
  NAND2_X1 U7164 ( .A1(n5951), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n6074) );
  INV_X1 U7165 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n7743) );
  OR2_X1 U7166 ( .A1(n5959), .A2(n7743), .ZN(n6073) );
  INV_X1 U7167 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n7742) );
  OR2_X1 U7168 ( .A1(n8428), .A2(n7742), .ZN(n6072) );
  NAND2_X1 U7169 ( .A1(n6069), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n6070) );
  AND2_X1 U7170 ( .A1(n6082), .A2(n6070), .ZN(n8053) );
  OR2_X1 U7171 ( .A1(n5135), .A2(n8053), .ZN(n6071) );
  OR2_X1 U7172 ( .A1(n8061), .A2(n9251), .ZN(n7962) );
  XNOR2_X1 U7173 ( .A(n6076), .B(n6075), .ZN(n6587) );
  NAND2_X1 U7174 ( .A1(n6587), .A2(n8421), .ZN(n6080) );
  NAND2_X1 U7175 ( .A1(n6205), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6097) );
  XNOR2_X1 U7176 ( .A(n6097), .B(P2_IR_REG_11__SCAN_IN), .ZN(n8078) );
  AOI22_X1 U7177 ( .A1(n6224), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n7009), .B2(
        n8078), .ZN(n6079) );
  NAND2_X1 U7178 ( .A1(n5951), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n6087) );
  INV_X1 U7179 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n7956) );
  OR2_X1 U7180 ( .A1(n5959), .A2(n7956), .ZN(n6086) );
  INV_X1 U7181 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n6081) );
  OR2_X1 U7182 ( .A1(n8428), .A2(n6081), .ZN(n6085) );
  NAND2_X1 U7183 ( .A1(n6082), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n6083) );
  AND2_X1 U7184 ( .A1(n6102), .A2(n6083), .ZN(n8120) );
  OR2_X1 U7185 ( .A1(n5135), .A2(n8120), .ZN(n6084) );
  NAND4_X1 U7186 ( .A1(n6087), .A2(n6086), .A3(n6085), .A4(n6084), .ZN(n9250)
         );
  OR2_X1 U7187 ( .A1(n8122), .A2(n9250), .ZN(n6088) );
  AND2_X1 U7188 ( .A1(n7962), .A2(n6088), .ZN(n6089) );
  AND2_X1 U7189 ( .A1(n7949), .A2(n6089), .ZN(n6091) );
  INV_X1 U7190 ( .A(n6089), .ZN(n6090) );
  NAND2_X1 U7191 ( .A1(n8061), .A2(n9251), .ZN(n7961) );
  NAND2_X1 U7192 ( .A1(n8122), .A2(n9250), .ZN(n8000) );
  NAND2_X1 U7193 ( .A1(n6093), .A2(n6092), .ZN(n6095) );
  NAND2_X1 U7194 ( .A1(n6095), .A2(n6094), .ZN(n7031) );
  OR2_X1 U7195 ( .A1(n7031), .A2(n5972), .ZN(n6100) );
  INV_X1 U7196 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n6096) );
  NAND2_X1 U7197 ( .A1(n6097), .A2(n6096), .ZN(n6098) );
  NAND2_X1 U7198 ( .A1(n6098), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6113) );
  XNOR2_X1 U7199 ( .A(n6113), .B(P2_IR_REG_12__SCAN_IN), .ZN(n8099) );
  AOI22_X1 U7200 ( .A1(n6224), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n7009), .B2(
        n8099), .ZN(n6099) );
  NAND2_X1 U7201 ( .A1(n5951), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n6107) );
  INV_X1 U7202 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n6101) );
  OR2_X1 U7203 ( .A1(n8428), .A2(n6101), .ZN(n6106) );
  AND2_X1 U7204 ( .A1(n6102), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n6103) );
  NOR2_X1 U7205 ( .A1(n6118), .A2(n6103), .ZN(n8201) );
  OR2_X1 U7206 ( .A1(n5135), .A2(n8201), .ZN(n6105) );
  INV_X1 U7207 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n8004) );
  OR2_X1 U7208 ( .A1(n5959), .A2(n8004), .ZN(n6104) );
  NAND2_X1 U7209 ( .A1(n8203), .A2(n9249), .ZN(n8196) );
  AND2_X1 U7210 ( .A1(n8000), .A2(n8196), .ZN(n8168) );
  OR2_X1 U7211 ( .A1(n6109), .A2(n6108), .ZN(n6110) );
  NAND2_X1 U7212 ( .A1(n6111), .A2(n6110), .ZN(n7101) );
  INV_X1 U7213 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n6112) );
  NAND2_X1 U7214 ( .A1(n6113), .A2(n6112), .ZN(n6114) );
  NAND2_X1 U7215 ( .A1(n6114), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6135) );
  XNOR2_X1 U7216 ( .A(n6135), .B(P2_IR_REG_13__SCAN_IN), .ZN(n8270) );
  AOI22_X1 U7217 ( .A1(n6224), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n7009), .B2(
        n8270), .ZN(n6115) );
  NAND2_X1 U7218 ( .A1(n5951), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n6124) );
  INV_X1 U7219 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n6117) );
  OR2_X1 U7220 ( .A1(n8428), .A2(n6117), .ZN(n6123) );
  NOR2_X1 U7221 ( .A1(n6118), .A2(n9915), .ZN(n6119) );
  OR2_X1 U7222 ( .A1(n5135), .A2(n5153), .ZN(n6122) );
  INV_X1 U7223 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n6120) );
  OR2_X1 U7224 ( .A1(n5959), .A2(n6120), .ZN(n6121) );
  NAND4_X1 U7225 ( .A1(n6124), .A2(n6123), .A3(n6122), .A4(n6121), .ZN(n9248)
         );
  NAND2_X1 U7226 ( .A1(n11103), .A2(n9248), .ZN(n6125) );
  AND2_X1 U7227 ( .A1(n8168), .A2(n6125), .ZN(n6127) );
  OR2_X1 U7228 ( .A1(n8203), .A2(n9249), .ZN(n8195) );
  INV_X1 U7229 ( .A(n8195), .ZN(n8170) );
  AND2_X1 U7230 ( .A1(n6125), .A2(n8170), .ZN(n6126) );
  AOI21_X1 U7231 ( .B1(n8169), .B2(n6127), .A(n6126), .ZN(n6129) );
  OR2_X1 U7232 ( .A1(n11103), .A2(n9248), .ZN(n6128) );
  NAND2_X1 U7233 ( .A1(n6133), .A2(n6132), .ZN(n8377) );
  INV_X1 U7234 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n6134) );
  NAND2_X1 U7235 ( .A1(n6135), .A2(n6134), .ZN(n6136) );
  NAND2_X1 U7236 ( .A1(n6136), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6154) );
  XNOR2_X1 U7237 ( .A(n6154), .B(P2_IR_REG_14__SCAN_IN), .ZN(n8277) );
  AOI22_X1 U7238 ( .A1(n8277), .A2(n7009), .B1(n6224), .B2(
        P1_DATAO_REG_14__SCAN_IN), .ZN(n6137) );
  NOR2_X1 U7239 ( .A1(n6139), .A2(n9884), .ZN(n6140) );
  OR2_X1 U7240 ( .A1(n6157), .A2(n6140), .ZN(n9128) );
  NAND2_X1 U7241 ( .A1(n5134), .A2(n9128), .ZN(n6147) );
  INV_X1 U7242 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n6141) );
  OR2_X1 U7243 ( .A1(n5959), .A2(n6141), .ZN(n6146) );
  INV_X1 U7244 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n6142) );
  OR2_X1 U7245 ( .A1(n8428), .A2(n6142), .ZN(n6145) );
  INV_X1 U7246 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n6143) );
  OR2_X1 U7247 ( .A1(n6330), .A2(n6143), .ZN(n6144) );
  NAND4_X1 U7248 ( .A1(n6147), .A2(n6146), .A3(n6145), .A4(n6144), .ZN(n9247)
         );
  INV_X1 U7249 ( .A(n6365), .ZN(n6148) );
  NAND2_X1 U7250 ( .A1(n9129), .A2(n9247), .ZN(n8560) );
  OR2_X1 U7251 ( .A1(n6150), .A2(n6149), .ZN(n6151) );
  INV_X1 U7252 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n6153) );
  NAND2_X1 U7253 ( .A1(n6154), .A2(n6153), .ZN(n6155) );
  NAND2_X1 U7254 ( .A1(n6155), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6169) );
  XNOR2_X1 U7255 ( .A(n6169), .B(P2_IR_REG_15__SCAN_IN), .ZN(n9298) );
  AOI22_X1 U7256 ( .A1(n9298), .A2(n7009), .B1(n6224), .B2(
        P1_DATAO_REG_15__SCAN_IN), .ZN(n6156) );
  OR2_X1 U7257 ( .A1(n6157), .A2(n9228), .ZN(n6158) );
  NAND2_X1 U7258 ( .A1(n6175), .A2(n6158), .ZN(n9235) );
  NAND2_X1 U7259 ( .A1(n5134), .A2(n9235), .ZN(n6164) );
  INV_X1 U7260 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n8108) );
  OR2_X1 U7261 ( .A1(n5959), .A2(n8108), .ZN(n6163) );
  INV_X1 U7262 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n6159) );
  OR2_X1 U7263 ( .A1(n8428), .A2(n6159), .ZN(n6162) );
  INV_X1 U7264 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n6160) );
  OR2_X1 U7265 ( .A1(n6330), .A2(n6160), .ZN(n6161) );
  NAND4_X1 U7266 ( .A1(n6164), .A2(n6163), .A3(n6162), .A4(n6161), .ZN(n9246)
         );
  INV_X1 U7267 ( .A(n9246), .ZN(n8478) );
  NOR2_X1 U7268 ( .A1(n8477), .A2(n8478), .ZN(n8481) );
  INV_X1 U7269 ( .A(n8481), .ZN(n6165) );
  AND2_X1 U7270 ( .A1(n8477), .A2(n8478), .ZN(n8480) );
  INV_X1 U7271 ( .A(n8480), .ZN(n6370) );
  XNOR2_X1 U7272 ( .A(n6167), .B(n6166), .ZN(n7329) );
  NAND2_X1 U7273 ( .A1(n7329), .A2(n8421), .ZN(n6174) );
  INV_X1 U7274 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n6168) );
  NAND2_X1 U7275 ( .A1(n6169), .A2(n6168), .ZN(n6170) );
  NAND2_X1 U7276 ( .A1(n6170), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6171) );
  NAND2_X1 U7277 ( .A1(n6171), .A2(n6206), .ZN(n6187) );
  OR2_X1 U7278 ( .A1(n6171), .A2(n6206), .ZN(n6172) );
  AOI22_X1 U7279 ( .A1(n9307), .A2(n7009), .B1(n6224), .B2(
        P1_DATAO_REG_16__SCAN_IN), .ZN(n6173) );
  NAND2_X1 U7280 ( .A1(n6174), .A2(n6173), .ZN(n8387) );
  NAND2_X1 U7281 ( .A1(n6175), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n6176) );
  NAND2_X1 U7282 ( .A1(n6191), .A2(n6176), .ZN(n9166) );
  NAND2_X1 U7283 ( .A1(n5134), .A2(n9166), .ZN(n6182) );
  INV_X1 U7284 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n9301) );
  OR2_X1 U7285 ( .A1(n5959), .A2(n9301), .ZN(n6181) );
  INV_X1 U7286 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n6177) );
  OR2_X1 U7287 ( .A1(n8428), .A2(n6177), .ZN(n6180) );
  INV_X1 U7288 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n6178) );
  OR2_X1 U7289 ( .A1(n6330), .A2(n6178), .ZN(n6179) );
  NAND4_X1 U7290 ( .A1(n6182), .A2(n6181), .A3(n6180), .A4(n6179), .ZN(n9245)
         );
  INV_X1 U7291 ( .A(n9245), .ZN(n9232) );
  NAND2_X1 U7292 ( .A1(n8387), .A2(n9232), .ZN(n8565) );
  NAND2_X1 U7293 ( .A1(n8125), .A2(n8483), .ZN(n6184) );
  NAND2_X1 U7294 ( .A1(n8387), .A2(n9245), .ZN(n6183) );
  NAND2_X1 U7295 ( .A1(n6184), .A2(n6183), .ZN(n8209) );
  XNOR2_X1 U7296 ( .A(n6186), .B(n6185), .ZN(n7406) );
  NAND2_X1 U7297 ( .A1(n7406), .A2(n8421), .ZN(n6190) );
  NAND2_X1 U7298 ( .A1(n6187), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6188) );
  XNOR2_X1 U7299 ( .A(n6188), .B(P2_IR_REG_17__SCAN_IN), .ZN(n10940) );
  AOI22_X1 U7300 ( .A1(n10940), .A2(n7009), .B1(n6224), .B2(
        P1_DATAO_REG_17__SCAN_IN), .ZN(n6189) );
  NAND2_X1 U7301 ( .A1(n6191), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n6193) );
  INV_X1 U7302 ( .A(n6192), .ZN(n6214) );
  NAND2_X1 U7303 ( .A1(n6193), .A2(n6214), .ZN(n9174) );
  NAND2_X1 U7304 ( .A1(n5134), .A2(n9174), .ZN(n6198) );
  INV_X1 U7305 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n9318) );
  OR2_X1 U7306 ( .A1(n5959), .A2(n9318), .ZN(n6197) );
  INV_X1 U7307 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n9317) );
  OR2_X1 U7308 ( .A1(n8428), .A2(n9317), .ZN(n6196) );
  INV_X1 U7309 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n6194) );
  OR2_X1 U7310 ( .A1(n6330), .A2(n6194), .ZN(n6195) );
  NAND4_X1 U7311 ( .A1(n6198), .A2(n6197), .A3(n6196), .A4(n6195), .ZN(n9493)
         );
  XNOR2_X1 U7312 ( .A(n9178), .B(n9164), .ZN(n8462) );
  NAND2_X1 U7313 ( .A1(n8209), .A2(n8462), .ZN(n6200) );
  NAND2_X1 U7314 ( .A1(n9178), .A2(n9493), .ZN(n6199) );
  NAND2_X1 U7315 ( .A1(n6200), .A2(n6199), .ZN(n9489) );
  NAND2_X1 U7316 ( .A1(n5681), .A2(n6202), .ZN(n6203) );
  NAND2_X1 U7317 ( .A1(n6204), .A2(n6203), .ZN(n7411) );
  OR2_X1 U7318 ( .A1(n7411), .A2(n5972), .ZN(n6212) );
  NOR2_X1 U7319 ( .A1(P2_IR_REG_13__SCAN_IN), .A2(P2_IR_REG_15__SCAN_IN), .ZN(
        n6209) );
  NOR2_X1 U7320 ( .A1(P2_IR_REG_11__SCAN_IN), .A2(P2_IR_REG_14__SCAN_IN), .ZN(
        n6208) );
  NOR2_X1 U7321 ( .A1(P2_IR_REG_12__SCAN_IN), .A2(P2_IR_REG_17__SCAN_IN), .ZN(
        n6207) );
  NAND2_X1 U7322 ( .A1(n6223), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6210) );
  XNOR2_X1 U7323 ( .A(n6210), .B(P2_IR_REG_18__SCAN_IN), .ZN(n10979) );
  AOI22_X1 U7324 ( .A1(n6224), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n7009), .B2(
        n10979), .ZN(n6211) );
  NAND2_X1 U7325 ( .A1(n6305), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n6218) );
  INV_X1 U7326 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n9562) );
  OR2_X1 U7327 ( .A1(n8428), .A2(n9562), .ZN(n6217) );
  AOI21_X1 U7328 ( .B1(P2_REG3_REG_18__SCAN_IN), .B2(n6214), .A(n6213), .ZN(
        n9498) );
  OR2_X1 U7329 ( .A1(n5135), .A2(n9498), .ZN(n6216) );
  INV_X1 U7330 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n9604) );
  OR2_X1 U7331 ( .A1(n6330), .A2(n9604), .ZN(n6215) );
  NAND4_X1 U7332 ( .A1(n6218), .A2(n6217), .A3(n6216), .A4(n6215), .ZN(n9244)
         );
  AND2_X1 U7333 ( .A1(n9508), .A2(n9244), .ZN(n6220) );
  OR2_X1 U7334 ( .A1(n9508), .A2(n9244), .ZN(n6219) );
  XNOR2_X1 U7335 ( .A(n6222), .B(n6221), .ZN(n7657) );
  NAND2_X1 U7336 ( .A1(n7657), .A2(n8421), .ZN(n6226) );
  AOI22_X1 U7337 ( .A1(n6224), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n9327), .B2(
        n7009), .ZN(n6225) );
  NAND2_X1 U7338 ( .A1(n5951), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n6232) );
  INV_X1 U7339 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n9314) );
  OR2_X1 U7340 ( .A1(n8428), .A2(n9314), .ZN(n6231) );
  NAND2_X1 U7341 ( .A1(P2_REG3_REG_19__SCAN_IN), .A2(n6227), .ZN(n6228) );
  AND2_X1 U7342 ( .A1(n6239), .A2(n6228), .ZN(n9480) );
  OR2_X1 U7343 ( .A1(n5135), .A2(n9480), .ZN(n6230) );
  INV_X1 U7344 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n9481) );
  OR2_X1 U7345 ( .A1(n5959), .A2(n9481), .ZN(n6229) );
  NAND4_X1 U7346 ( .A1(n6232), .A2(n6231), .A3(n6230), .A4(n6229), .ZN(n9494)
         );
  NAND2_X1 U7347 ( .A1(n9554), .A2(n9494), .ZN(n6233) );
  XNOR2_X1 U7348 ( .A(n6235), .B(n6234), .ZN(n7905) );
  NAND2_X1 U7349 ( .A1(n7905), .A2(n8421), .ZN(n6237) );
  INV_X1 U7350 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n7906) );
  OR2_X1 U7351 ( .A1(n5966), .A2(n7906), .ZN(n6236) );
  NAND2_X1 U7352 ( .A1(n6329), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n6243) );
  INV_X1 U7353 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n6238) );
  OR2_X1 U7354 ( .A1(n6330), .A2(n6238), .ZN(n6242) );
  XNOR2_X1 U7355 ( .A(n6239), .B(n9914), .ZN(n9463) );
  OR2_X1 U7356 ( .A1(n5135), .A2(n9463), .ZN(n6241) );
  INV_X1 U7357 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n9464) );
  OR2_X1 U7358 ( .A1(n5959), .A2(n9464), .ZN(n6240) );
  NAND4_X1 U7359 ( .A1(n6243), .A2(n6242), .A3(n6241), .A4(n6240), .ZN(n9448)
         );
  NAND2_X1 U7360 ( .A1(n9549), .A2(n9477), .ZN(n8582) );
  NAND2_X1 U7361 ( .A1(n8581), .A2(n8582), .ZN(n9459) );
  INV_X1 U7362 ( .A(n6244), .ZN(n6246) );
  NAND2_X1 U7363 ( .A1(n6246), .A2(n6245), .ZN(n6247) );
  NAND2_X1 U7364 ( .A1(n6248), .A2(n6247), .ZN(n9108) );
  OR2_X1 U7365 ( .A1(n9108), .A2(n5972), .ZN(n6250) );
  INV_X1 U7366 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n9107) );
  OR2_X1 U7367 ( .A1(n5966), .A2(n9107), .ZN(n6249) );
  NAND2_X1 U7368 ( .A1(n6305), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n6258) );
  INV_X1 U7369 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n6251) );
  OR2_X1 U7370 ( .A1(n8428), .A2(n6251), .ZN(n6257) );
  NAND2_X1 U7371 ( .A1(n6252), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n6253) );
  AND2_X1 U7372 ( .A1(n6267), .A2(n6253), .ZN(n9450) );
  OR2_X1 U7373 ( .A1(n5135), .A2(n9450), .ZN(n6256) );
  INV_X1 U7374 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n6254) );
  OR2_X1 U7375 ( .A1(n6330), .A2(n6254), .ZN(n6255) );
  NAND4_X1 U7376 ( .A1(n6258), .A2(n6257), .A3(n6256), .A4(n6255), .ZN(n9461)
         );
  XNOR2_X1 U7377 ( .A(n9545), .B(n9461), .ZN(n9453) );
  NAND2_X1 U7378 ( .A1(n9446), .A2(n5417), .ZN(n6260) );
  OR2_X1 U7379 ( .A1(n9545), .A2(n9461), .ZN(n6259) );
  NAND2_X1 U7380 ( .A1(n6260), .A2(n6259), .ZN(n9433) );
  OR2_X1 U7381 ( .A1(n6262), .A2(n6261), .ZN(n6263) );
  NAND2_X1 U7382 ( .A1(n6264), .A2(n6263), .ZN(n7997) );
  OR2_X1 U7383 ( .A1(n7997), .A2(n5972), .ZN(n6266) );
  INV_X1 U7384 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n7974) );
  OR2_X1 U7385 ( .A1(n5966), .A2(n7974), .ZN(n6265) );
  NAND2_X1 U7386 ( .A1(n6305), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n6272) );
  INV_X1 U7387 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n9543) );
  OR2_X1 U7388 ( .A1(n8428), .A2(n9543), .ZN(n6271) );
  NAND2_X1 U7389 ( .A1(n6267), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n6268) );
  AND2_X1 U7390 ( .A1(n6279), .A2(n6268), .ZN(n8415) );
  OR2_X1 U7391 ( .A1(n5135), .A2(n8415), .ZN(n6270) );
  INV_X1 U7392 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n9598) );
  OR2_X1 U7393 ( .A1(n6330), .A2(n9598), .ZN(n6269) );
  NAND4_X1 U7394 ( .A1(n6272), .A2(n6271), .A3(n6270), .A4(n6269), .ZN(n9447)
         );
  NOR2_X1 U7395 ( .A1(n8589), .A2(n9447), .ZN(n6273) );
  NAND2_X1 U7396 ( .A1(n8589), .A2(n9447), .ZN(n6274) );
  XNOR2_X1 U7397 ( .A(n6276), .B(n6275), .ZN(n8032) );
  NAND2_X1 U7398 ( .A1(n8032), .A2(n8421), .ZN(n6278) );
  INV_X1 U7399 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n8035) );
  OR2_X1 U7400 ( .A1(n5966), .A2(n8035), .ZN(n6277) );
  NAND2_X1 U7401 ( .A1(n6329), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n6284) );
  INV_X1 U7402 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n9427) );
  OR2_X1 U7403 ( .A1(n5959), .A2(n9427), .ZN(n6283) );
  NAND2_X1 U7404 ( .A1(n6279), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n6280) );
  AND2_X1 U7405 ( .A1(n6290), .A2(n6280), .ZN(n9426) );
  OR2_X1 U7406 ( .A1(n5135), .A2(n9426), .ZN(n6282) );
  INV_X1 U7407 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n9594) );
  OR2_X1 U7408 ( .A1(n6330), .A2(n9594), .ZN(n6281) );
  AND2_X1 U7409 ( .A1(n9425), .A2(n9243), .ZN(n6285) );
  XNOR2_X1 U7410 ( .A(n6287), .B(n6286), .ZN(n8140) );
  NAND2_X1 U7411 ( .A1(n8140), .A2(n8421), .ZN(n6289) );
  INV_X1 U7412 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n8141) );
  OR2_X1 U7413 ( .A1(n5966), .A2(n8141), .ZN(n6288) );
  NAND2_X1 U7414 ( .A1(n6329), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n6296) );
  INV_X1 U7415 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n9590) );
  OR2_X1 U7416 ( .A1(n6330), .A2(n9590), .ZN(n6295) );
  NAND2_X1 U7417 ( .A1(n6290), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n6291) );
  AND2_X1 U7418 ( .A1(n6307), .A2(n6291), .ZN(n9413) );
  OR2_X1 U7419 ( .A1(n5135), .A2(n9413), .ZN(n6294) );
  INV_X1 U7420 ( .A(P2_REG2_REG_24__SCAN_IN), .ZN(n6292) );
  OR2_X1 U7421 ( .A1(n5959), .A2(n6292), .ZN(n6293) );
  NAND4_X1 U7422 ( .A1(n6296), .A2(n6295), .A3(n6294), .A4(n6293), .ZN(n9242)
         );
  AND2_X1 U7423 ( .A1(n9188), .A2(n9242), .ZN(n8597) );
  INV_X1 U7424 ( .A(n8597), .ZN(n8465) );
  NOR2_X1 U7425 ( .A1(n9188), .A2(n9242), .ZN(n8600) );
  INV_X1 U7426 ( .A(n8600), .ZN(n8466) );
  INV_X1 U7427 ( .A(n6298), .ZN(n6300) );
  NAND2_X1 U7428 ( .A1(n6300), .A2(n6299), .ZN(n6301) );
  NAND2_X1 U7429 ( .A1(n6302), .A2(n6301), .ZN(n8163) );
  OR2_X1 U7430 ( .A1(n8163), .A2(n5972), .ZN(n6304) );
  INV_X1 U7431 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n8134) );
  OR2_X1 U7432 ( .A1(n5966), .A2(n8134), .ZN(n6303) );
  NAND2_X1 U7433 ( .A1(n6305), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n6314) );
  INV_X1 U7434 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n6306) );
  OR2_X1 U7435 ( .A1(n8428), .A2(n6306), .ZN(n6313) );
  NAND2_X1 U7436 ( .A1(n6307), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n6308) );
  AND2_X1 U7437 ( .A1(n6309), .A2(n6308), .ZN(n9406) );
  OR2_X1 U7438 ( .A1(n5135), .A2(n9406), .ZN(n6312) );
  INV_X1 U7439 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n6310) );
  OR2_X1 U7440 ( .A1(n6330), .A2(n6310), .ZN(n6311) );
  NAND4_X1 U7441 ( .A1(n6314), .A2(n6313), .A3(n6312), .A4(n6311), .ZN(n9389)
         );
  NAND2_X1 U7442 ( .A1(n9529), .A2(n9389), .ZN(n6316) );
  NOR2_X1 U7443 ( .A1(n9529), .A2(n9389), .ZN(n6315) );
  OAI21_X1 U7444 ( .B1(n9105), .B2(n5137), .A(n9361), .ZN(n6318) );
  INV_X1 U7445 ( .A(n5137), .ZN(n8475) );
  NAND2_X1 U7446 ( .A1(n6318), .A2(n6317), .ZN(n6335) );
  NAND2_X1 U7447 ( .A1(n6320), .A2(n6319), .ZN(n6325) );
  INV_X1 U7448 ( .A(n6321), .ZN(n6323) );
  NAND2_X1 U7449 ( .A1(n6323), .A2(n6322), .ZN(n6324) );
  NAND2_X1 U7450 ( .A1(n6325), .A2(n6324), .ZN(n8296) );
  MUX2_X1 U7451 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(P1_DATAO_REG_29__SCAN_IN), 
        .S(n8306), .Z(n8297) );
  XNOR2_X1 U7452 ( .A(n8296), .B(n8297), .ZN(n8295) );
  INV_X1 U7453 ( .A(n8295), .ZN(n6326) );
  NAND2_X1 U7454 ( .A1(n6779), .A2(n8421), .ZN(n6328) );
  INV_X1 U7455 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n8331) );
  OR2_X1 U7456 ( .A1(n5966), .A2(n8331), .ZN(n6327) );
  NAND2_X1 U7457 ( .A1(n6328), .A2(n6327), .ZN(n6435) );
  NAND2_X1 U7458 ( .A1(n6329), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n6334) );
  INV_X1 U7459 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n6431) );
  OR2_X1 U7460 ( .A1(n6330), .A2(n6431), .ZN(n6333) );
  INV_X1 U7461 ( .A(P2_REG2_REG_29__SCAN_IN), .ZN(n6331) );
  OR2_X1 U7462 ( .A1(n5959), .A2(n6331), .ZN(n6332) );
  NAND4_X1 U7463 ( .A1(n8432), .A2(n6334), .A3(n6333), .A4(n6332), .ZN(n9241)
         );
  INV_X1 U7464 ( .A(n9241), .ZN(n9363) );
  OR2_X1 U7465 ( .A1(n6435), .A2(n9363), .ZN(n8439) );
  NAND2_X1 U7466 ( .A1(n6435), .A2(n9363), .ZN(n8619) );
  NAND2_X1 U7467 ( .A1(n8439), .A2(n8619), .ZN(n6385) );
  OR2_X1 U7468 ( .A1(n6341), .A2(n6340), .ZN(n6342) );
  OR2_X1 U7469 ( .A1(n6896), .A2(n8624), .ZN(n6346) );
  NAND2_X1 U7470 ( .A1(n5204), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6344) );
  NAND2_X1 U7471 ( .A1(n9327), .A2(n8630), .ZN(n6345) );
  INV_X1 U7472 ( .A(n6347), .ZN(n8627) );
  NAND2_X1 U7473 ( .A1(n8627), .A2(n9328), .ZN(n6349) );
  AND2_X1 U7474 ( .A1(n6893), .A2(n6349), .ZN(n6932) );
  AND2_X1 U7475 ( .A1(n6893), .A2(P2_B_REG_SCAN_IN), .ZN(n6350) );
  NOR2_X1 U7476 ( .A1(n9476), .A2(n6350), .ZN(n9350) );
  NAND2_X1 U7477 ( .A1(n5951), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n6356) );
  INV_X1 U7478 ( .A(P2_REG2_REG_30__SCAN_IN), .ZN(n6351) );
  OR2_X1 U7479 ( .A1(n5959), .A2(n6351), .ZN(n6355) );
  INV_X1 U7480 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n6352) );
  OR2_X1 U7481 ( .A1(n6353), .A2(n6352), .ZN(n6354) );
  NAND4_X1 U7482 ( .A1(n8432), .A2(n6356), .A3(n6355), .A4(n6354), .ZN(n9240)
         );
  INV_X1 U7483 ( .A(n6932), .ZN(n6930) );
  AOI22_X1 U7484 ( .A1(n9350), .A2(n9240), .B1(n9492), .B2(n5137), .ZN(n6357)
         );
  NAND2_X1 U7485 ( .A1(n6908), .A2(n7468), .ZN(n8505) );
  NAND2_X1 U7486 ( .A1(n8511), .A2(n8505), .ZN(n8444) );
  INV_X1 U7487 ( .A(n8444), .ZN(n7287) );
  NAND2_X1 U7488 ( .A1(n7297), .A2(n8489), .ZN(n7313) );
  NAND2_X1 U7489 ( .A1(n7314), .A2(n8495), .ZN(n7284) );
  NAND2_X1 U7490 ( .A1(n7287), .A2(n7284), .ZN(n7283) );
  NAND2_X1 U7491 ( .A1(n7478), .A2(n7587), .ZN(n8503) );
  INV_X1 U7492 ( .A(n8503), .ZN(n8509) );
  NOR2_X1 U7493 ( .A1(n7478), .A2(n7587), .ZN(n8506) );
  INV_X1 U7494 ( .A(n8506), .ZN(n8512) );
  NAND2_X1 U7495 ( .A1(n9256), .A2(n6358), .ZN(n8516) );
  INV_X1 U7496 ( .A(n8516), .ZN(n6359) );
  NOR2_X1 U7497 ( .A1(n9256), .A2(n6358), .ZN(n8508) );
  INV_X1 U7498 ( .A(n8508), .ZN(n8515) );
  OAI21_X2 U7499 ( .B1(n7474), .B2(n6359), .A(n8515), .ZN(n7510) );
  OR2_X1 U7500 ( .A1(n7689), .A2(n7673), .ZN(n8519) );
  NAND2_X1 U7501 ( .A1(n7689), .A2(n7673), .ZN(n8518) );
  NAND2_X1 U7502 ( .A1(n6360), .A2(n7661), .ZN(n8540) );
  INV_X1 U7503 ( .A(n8540), .ZN(n6361) );
  NAND2_X1 U7504 ( .A1(n7563), .A2(n6361), .ZN(n6362) );
  NAND2_X1 U7505 ( .A1(n6362), .A2(n8528), .ZN(n7850) );
  NOR2_X1 U7506 ( .A1(n8061), .A2(n8117), .ZN(n8538) );
  NAND2_X1 U7507 ( .A1(n8061), .A2(n8117), .ZN(n8542) );
  NOR2_X1 U7508 ( .A1(n8122), .A2(n8003), .ZN(n8546) );
  INV_X1 U7509 ( .A(n8546), .ZN(n8536) );
  NAND2_X1 U7510 ( .A1(n8122), .A2(n8003), .ZN(n8545) );
  NAND2_X1 U7511 ( .A1(n7955), .A2(n8443), .ZN(n7954) );
  NAND2_X1 U7512 ( .A1(n7954), .A2(n8545), .ZN(n7999) );
  OR2_X1 U7513 ( .A1(n8203), .A2(n8174), .ZN(n8550) );
  NAND2_X1 U7514 ( .A1(n7999), .A2(n8550), .ZN(n6364) );
  NAND2_X1 U7515 ( .A1(n8203), .A2(n8174), .ZN(n8551) );
  NAND2_X1 U7516 ( .A1(n6364), .A2(n8551), .ZN(n8036) );
  XNOR2_X1 U7517 ( .A(n11103), .B(n9248), .ZN(n8553) );
  NAND2_X1 U7518 ( .A1(n6365), .A2(n8560), .ZN(n8479) );
  INV_X1 U7519 ( .A(n9247), .ZN(n8381) );
  NAND2_X1 U7520 ( .A1(n9129), .A2(n8381), .ZN(n6368) );
  AND2_X1 U7521 ( .A1(n8553), .A2(n6369), .ZN(n6367) );
  INV_X1 U7522 ( .A(n9248), .ZN(n9126) );
  AND2_X1 U7523 ( .A1(n11103), .A2(n9126), .ZN(n8557) );
  INV_X1 U7524 ( .A(n8557), .ZN(n8037) );
  AND2_X1 U7525 ( .A1(n8105), .A2(n6370), .ZN(n8127) );
  INV_X1 U7526 ( .A(n8483), .ZN(n6371) );
  AND2_X1 U7527 ( .A1(n8127), .A2(n6371), .ZN(n6373) );
  NAND2_X1 U7528 ( .A1(n9178), .A2(n9164), .ZN(n6375) );
  NAND2_X1 U7529 ( .A1(n8206), .A2(n6375), .ZN(n9502) );
  NAND2_X1 U7530 ( .A1(n9508), .A2(n9475), .ZN(n8574) );
  NAND2_X1 U7531 ( .A1(n8577), .A2(n8574), .ZN(n9501) );
  INV_X1 U7532 ( .A(n9494), .ZN(n9207) );
  OR2_X1 U7533 ( .A1(n9554), .A2(n9207), .ZN(n6376) );
  NAND2_X1 U7534 ( .A1(n9482), .A2(n6376), .ZN(n9467) );
  NAND2_X1 U7535 ( .A1(n9467), .A2(n9466), .ZN(n9465) );
  NAND2_X1 U7536 ( .A1(n9465), .A2(n8581), .ZN(n9454) );
  NAND2_X1 U7537 ( .A1(n9454), .A2(n9453), .ZN(n9452) );
  INV_X1 U7538 ( .A(n9461), .ZN(n9436) );
  OR2_X1 U7539 ( .A1(n9545), .A2(n9436), .ZN(n6377) );
  NAND2_X1 U7540 ( .A1(n9452), .A2(n6377), .ZN(n9437) );
  INV_X1 U7541 ( .A(n9447), .ZN(n9421) );
  NAND2_X1 U7542 ( .A1(n8589), .A2(n9421), .ZN(n6378) );
  OR2_X1 U7543 ( .A1(n8589), .A2(n9421), .ZN(n6379) );
  OR2_X1 U7544 ( .A1(n9425), .A2(n9435), .ZN(n8593) );
  NAND2_X1 U7545 ( .A1(n9425), .A2(n9435), .ZN(n8592) );
  AND2_X1 U7546 ( .A1(n9188), .A2(n9422), .ZN(n6382) );
  OR2_X1 U7547 ( .A1(n9188), .A2(n9422), .ZN(n6381) );
  INV_X1 U7548 ( .A(n9389), .ZN(n9412) );
  NOR2_X1 U7549 ( .A1(n9529), .A2(n9412), .ZN(n8602) );
  AND2_X1 U7550 ( .A1(n9529), .A2(n9412), .ZN(n8601) );
  INV_X1 U7551 ( .A(n8601), .ZN(n6383) );
  OAI21_X2 U7552 ( .B1(n9399), .B2(n8602), .A(n6383), .ZN(n9393) );
  OR2_X1 U7553 ( .A1(n9220), .A2(n9403), .ZN(n8604) );
  NAND2_X1 U7554 ( .A1(n9220), .A2(n9403), .ZN(n8442) );
  INV_X1 U7555 ( .A(n8442), .ZN(n8606) );
  AOI21_X2 U7556 ( .B1(n9393), .B2(n8604), .A(n8606), .ZN(n9381) );
  NAND2_X1 U7557 ( .A1(n9099), .A2(n9362), .ZN(n8608) );
  OR2_X1 U7558 ( .A1(n9099), .A2(n9362), .ZN(n8441) );
  INV_X1 U7559 ( .A(n8441), .ZN(n8610) );
  NOR2_X1 U7560 ( .A1(n9582), .A2(n5137), .ZN(n6384) );
  XNOR2_X1 U7561 ( .A(n8425), .B(n6385), .ZN(n9354) );
  NAND2_X1 U7562 ( .A1(n8624), .A2(n9334), .ZN(n6869) );
  OR2_X1 U7563 ( .A1(n9327), .A2(n7975), .ZN(n6863) );
  NAND2_X1 U7564 ( .A1(n6869), .A2(n6863), .ZN(n6386) );
  AND2_X1 U7565 ( .A1(n9565), .A2(n6386), .ZN(n6387) );
  OR2_X1 U7566 ( .A1(n6895), .A2(n8630), .ZN(n8057) );
  AND2_X2 U7567 ( .A1(n9354), .A2(n9541), .ZN(n6388) );
  NAND3_X1 U7568 ( .A1(n8472), .A2(n8630), .A3(n9327), .ZN(n6422) );
  NAND3_X1 U7569 ( .A1(n8618), .A2(n9565), .A3(n6422), .ZN(n6915) );
  INV_X1 U7570 ( .A(n6895), .ZN(n6389) );
  NAND2_X1 U7571 ( .A1(n6915), .A2(n11105), .ZN(n6919) );
  INV_X1 U7572 ( .A(n6393), .ZN(n6391) );
  NAND2_X1 U7573 ( .A1(n6391), .A2(P2_IR_REG_24__SCAN_IN), .ZN(n6394) );
  XNOR2_X1 U7574 ( .A(n6406), .B(P2_B_REG_SCAN_IN), .ZN(n6398) );
  NAND2_X1 U7575 ( .A1(n6398), .A2(n8135), .ZN(n6404) );
  NAND2_X1 U7576 ( .A1(n6399), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6400) );
  MUX2_X1 U7577 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6400), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n6402) );
  NAND2_X1 U7578 ( .A1(n8282), .A2(n6406), .ZN(n6407) );
  NAND2_X1 U7579 ( .A1(n8282), .A2(n8135), .ZN(n6409) );
  NOR2_X1 U7580 ( .A1(P2_D_REG_31__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .ZN(
        n6414) );
  NOR4_X1 U7581 ( .A1(P2_D_REG_4__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .A3(
        P2_D_REG_29__SCAN_IN), .A4(P2_D_REG_28__SCAN_IN), .ZN(n6413) );
  NOR4_X1 U7582 ( .A1(P2_D_REG_23__SCAN_IN), .A2(P2_D_REG_22__SCAN_IN), .A3(
        P2_D_REG_21__SCAN_IN), .A4(P2_D_REG_20__SCAN_IN), .ZN(n6412) );
  NOR4_X1 U7583 ( .A1(P2_D_REG_27__SCAN_IN), .A2(P2_D_REG_26__SCAN_IN), .A3(
        P2_D_REG_25__SCAN_IN), .A4(P2_D_REG_24__SCAN_IN), .ZN(n6411) );
  NAND4_X1 U7584 ( .A1(n6414), .A2(n6413), .A3(n6412), .A4(n6411), .ZN(n6420)
         );
  NOR4_X1 U7585 ( .A1(P2_D_REG_15__SCAN_IN), .A2(P2_D_REG_14__SCAN_IN), .A3(
        P2_D_REG_13__SCAN_IN), .A4(P2_D_REG_12__SCAN_IN), .ZN(n6418) );
  NOR4_X1 U7586 ( .A1(P2_D_REG_17__SCAN_IN), .A2(P2_D_REG_19__SCAN_IN), .A3(
        P2_D_REG_18__SCAN_IN), .A4(P2_D_REG_16__SCAN_IN), .ZN(n6417) );
  NOR4_X1 U7587 ( .A1(P2_D_REG_7__SCAN_IN), .A2(P2_D_REG_6__SCAN_IN), .A3(
        P2_D_REG_5__SCAN_IN), .A4(P2_D_REG_2__SCAN_IN), .ZN(n6416) );
  NOR4_X1 U7588 ( .A1(P2_D_REG_11__SCAN_IN), .A2(P2_D_REG_10__SCAN_IN), .A3(
        P2_D_REG_9__SCAN_IN), .A4(P2_D_REG_8__SCAN_IN), .ZN(n6415) );
  NAND4_X1 U7589 ( .A1(n6418), .A2(n6417), .A3(n6416), .A4(n6415), .ZN(n6419)
         );
  NOR2_X1 U7590 ( .A1(n6420), .A2(n6419), .ZN(n6421) );
  AND3_X1 U7591 ( .A1(n6408), .A2(n7082), .A3(n6866), .ZN(n6933) );
  NAND2_X1 U7592 ( .A1(n6919), .A2(n6933), .ZN(n6427) );
  INV_X1 U7593 ( .A(n6422), .ZN(n6423) );
  INV_X1 U7594 ( .A(n6921), .ZN(n6914) );
  NAND2_X1 U7595 ( .A1(n6914), .A2(n7091), .ZN(n6425) );
  INV_X1 U7596 ( .A(n7082), .ZN(n9610) );
  NAND2_X1 U7597 ( .A1(n6865), .A2(n6866), .ZN(n6928) );
  INV_X1 U7598 ( .A(n6928), .ZN(n6424) );
  NAND2_X1 U7599 ( .A1(n6425), .A2(n6424), .ZN(n6426) );
  NAND2_X1 U7600 ( .A1(n6427), .A2(n6426), .ZN(n6430) );
  NAND2_X1 U7601 ( .A1(n6428), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6429) );
  NAND2_X1 U7602 ( .A1(n6432), .A2(n6431), .ZN(n6433) );
  NAND2_X1 U7603 ( .A1(n6434), .A2(n6433), .ZN(n6438) );
  INV_X1 U7604 ( .A(n6435), .ZN(n9357) );
  NAND2_X1 U7605 ( .A1(n11178), .A2(n9553), .ZN(n9607) );
  NAND2_X1 U7606 ( .A1(n6438), .A2(n6437), .ZN(P2_U3456) );
  NOR2_X1 U7607 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_8__SCAN_IN), .ZN(
        n6442) );
  NOR2_X1 U7608 ( .A1(P1_IR_REG_6__SCAN_IN), .A2(P1_IR_REG_7__SCAN_IN), .ZN(
        n6441) );
  NOR2_X1 U7609 ( .A1(P1_IR_REG_5__SCAN_IN), .A2(P1_IR_REG_10__SCAN_IN), .ZN(
        n6440) );
  NAND4_X1 U7610 ( .A1(n6442), .A2(n6441), .A3(n6440), .A4(n9782), .ZN(n6443)
         );
  NOR2_X1 U7611 ( .A1(P1_IR_REG_23__SCAN_IN), .A2(P1_IR_REG_22__SCAN_IN), .ZN(
        n6444) );
  NAND2_X1 U7612 ( .A1(n6445), .A2(n10013), .ZN(n6446) );
  INV_X1 U7613 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n6448) );
  XNOR2_X2 U7614 ( .A(n6450), .B(n10022), .ZN(n9080) );
  INV_X1 U7615 ( .A(n9080), .ZN(n6454) );
  NAND2_X1 U7616 ( .A1(n6454), .A2(n10700), .ZN(n6824) );
  INV_X1 U7617 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n6453) );
  OR2_X1 U7618 ( .A1(n6824), .A2(n6453), .ZN(n6459) );
  AND2_X2 U7619 ( .A1(n9080), .A2(n6455), .ZN(n6580) );
  NAND2_X1 U7620 ( .A1(n6580), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n6458) );
  INV_X1 U7621 ( .A(n6461), .ZN(n6462) );
  AOI21_X4 U7622 ( .B1(n6464), .B2(n6816), .A(n6463), .ZN(n6474) );
  INV_X1 U7623 ( .A(n6465), .ZN(n6466) );
  OAI22_X1 U7624 ( .A1(n6699), .A2(n6949), .B1(n6474), .B2(n7144), .ZN(n6467)
         );
  INV_X1 U7625 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n6950) );
  XNOR2_X2 U7626 ( .A(n11000), .B(n7729), .ZN(n8928) );
  NAND2_X1 U7627 ( .A1(n6520), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n6471) );
  NAND2_X1 U7628 ( .A1(n6580), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n6470) );
  NAND2_X1 U7629 ( .A1(n6782), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n6469) );
  NAND2_X1 U7630 ( .A1(n5133), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n6468) );
  NOR2_X1 U7631 ( .A1(n8306), .A2(n6472), .ZN(n6473) );
  XNOR2_X1 U7632 ( .A(n6473), .B(P2_DATAO_REG_0__SCAN_IN), .ZN(n10706) );
  INV_X1 U7633 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n10793) );
  MUX2_X1 U7634 ( .A(n10706), .B(n10793), .S(n6529), .Z(n7725) );
  AND2_X1 U7635 ( .A1(n10297), .A2(n7128), .ZN(n7723) );
  OR2_X1 U7636 ( .A1(n11000), .A2(n7729), .ZN(n6475) );
  NAND2_X1 U7637 ( .A1(n6580), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n6479) );
  NAND2_X1 U7638 ( .A1(n6782), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n6478) );
  NAND2_X1 U7639 ( .A1(n6729), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n6477) );
  NOR2_X1 U7640 ( .A1(n6699), .A2(n8374), .ZN(n6482) );
  INV_X1 U7641 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n6951) );
  OR2_X1 U7642 ( .A1(n6465), .A2(n10692), .ZN(n6480) );
  INV_X1 U7643 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n9764) );
  NAND2_X1 U7644 ( .A1(n6480), .A2(n9764), .ZN(n6492) );
  OAI21_X1 U7645 ( .B1(n6480), .B2(n9764), .A(n6492), .ZN(n7146) );
  OAI22_X1 U7646 ( .A1(n6646), .A2(n6951), .B1(n6474), .B2(n7146), .ZN(n6481)
         );
  NAND2_X1 U7647 ( .A1(n10295), .A2(n11013), .ZN(n8836) );
  NAND2_X1 U7648 ( .A1(n6483), .A2(n6484), .ZN(n8988) );
  NAND2_X2 U7649 ( .A1(n8836), .A2(n8988), .ZN(n10997) );
  NAND2_X1 U7650 ( .A1(n10994), .A2(n10997), .ZN(n6486) );
  OR2_X1 U7651 ( .A1(n10295), .A2(n6484), .ZN(n6485) );
  NAND2_X1 U7652 ( .A1(n6486), .A2(n6485), .ZN(n7642) );
  NAND2_X1 U7653 ( .A1(n6520), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n6491) );
  NAND2_X1 U7654 ( .A1(n6580), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n6490) );
  INV_X1 U7655 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n6487) );
  NAND2_X1 U7656 ( .A1(n6782), .A2(n6487), .ZN(n6489) );
  NAND2_X1 U7657 ( .A1(n5133), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n6488) );
  NAND4_X1 U7658 ( .A1(n6491), .A2(n6490), .A3(n6489), .A4(n6488), .ZN(n11001)
         );
  INV_X1 U7659 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n6943) );
  NAND2_X1 U7660 ( .A1(n6492), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6493) );
  INV_X1 U7661 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n9974) );
  XNOR2_X1 U7662 ( .A(n6493), .B(n9974), .ZN(n7148) );
  OAI22_X1 U7663 ( .A1(n6646), .A2(n6943), .B1(n6474), .B2(n7148), .ZN(n6495)
         );
  NOR2_X1 U7664 ( .A1(n6699), .A2(n6944), .ZN(n6494) );
  INV_X1 U7665 ( .A(n7654), .ZN(n11032) );
  NAND2_X1 U7666 ( .A1(n11001), .A2(n11032), .ZN(n8837) );
  NAND2_X1 U7667 ( .A1(n8993), .A2(n8837), .ZN(n8934) );
  NAND2_X1 U7668 ( .A1(n7642), .A2(n8934), .ZN(n6497) );
  OR2_X1 U7669 ( .A1(n11001), .A2(n7654), .ZN(n6496) );
  NAND2_X1 U7670 ( .A1(n6497), .A2(n6496), .ZN(n7815) );
  NAND2_X1 U7671 ( .A1(n6580), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n6502) );
  NAND2_X1 U7672 ( .A1(n5133), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n6501) );
  NOR2_X1 U7673 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n6498) );
  NOR2_X1 U7674 ( .A1(n6508), .A2(n6498), .ZN(n7820) );
  NAND2_X1 U7675 ( .A1(n6782), .A2(n7820), .ZN(n6500) );
  NAND2_X1 U7676 ( .A1(n6520), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n6499) );
  NAND4_X1 U7677 ( .A1(n6502), .A2(n6501), .A3(n6500), .A4(n6499), .ZN(n10294)
         );
  INV_X1 U7678 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n6952) );
  NAND2_X1 U7679 ( .A1(n6503), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6504) );
  XNOR2_X1 U7680 ( .A(n6504), .B(n6439), .ZN(n7150) );
  OAI22_X1 U7681 ( .A1(n6646), .A2(n6952), .B1(n6474), .B2(n7150), .ZN(n6506)
         );
  NOR2_X1 U7682 ( .A1(n6953), .A2(n6699), .ZN(n6505) );
  NOR2_X1 U7683 ( .A1(n10294), .A2(n7821), .ZN(n6507) );
  INV_X1 U7684 ( .A(n7821), .ZN(n11042) );
  INV_X1 U7685 ( .A(n10294), .ZN(n7646) );
  NAND2_X1 U7686 ( .A1(n6520), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n6512) );
  NAND2_X1 U7687 ( .A1(n6580), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n6511) );
  NAND2_X1 U7688 ( .A1(n5132), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n6510) );
  NAND2_X1 U7689 ( .A1(n6508), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n6522) );
  OAI21_X1 U7690 ( .B1(n6508), .B2(P1_REG3_REG_5__SCAN_IN), .A(n6522), .ZN(
        n7556) );
  OR2_X1 U7691 ( .A1(n6773), .A2(n7556), .ZN(n6509) );
  OR2_X1 U7692 ( .A1(n6956), .A2(n6699), .ZN(n6519) );
  INV_X1 U7693 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n6955) );
  NOR2_X1 U7694 ( .A1(n6513), .A2(P1_IR_REG_5__SCAN_IN), .ZN(n6539) );
  INV_X1 U7695 ( .A(n6539), .ZN(n6516) );
  NAND2_X1 U7696 ( .A1(n6513), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6514) );
  MUX2_X1 U7697 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6514), .S(
        P1_IR_REG_5__SCAN_IN), .Z(n6515) );
  NAND2_X1 U7698 ( .A1(n6516), .A2(n6515), .ZN(n7152) );
  OAI22_X1 U7699 ( .A1(n6646), .A2(n6955), .B1(n6474), .B2(n7152), .ZN(n6517)
         );
  INV_X1 U7700 ( .A(n6517), .ZN(n6518) );
  NAND2_X1 U7701 ( .A1(n6519), .A2(n6518), .ZN(n7545) );
  NAND2_X1 U7702 ( .A1(n7833), .A2(n7545), .ZN(n8843) );
  INV_X1 U7703 ( .A(n7833), .ZN(n10293) );
  NAND2_X1 U7704 ( .A1(n10293), .A2(n7557), .ZN(n8995) );
  NAND2_X1 U7705 ( .A1(n8843), .A2(n8995), .ZN(n8932) );
  INV_X1 U7706 ( .A(n8932), .ZN(n7415) );
  NAND2_X1 U7707 ( .A1(n7833), .A2(n7557), .ZN(n7828) );
  NAND2_X1 U7708 ( .A1(n6580), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n6527) );
  NAND2_X1 U7709 ( .A1(n6520), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n6526) );
  NOR2_X1 U7710 ( .A1(n6522), .A2(n6521), .ZN(n6533) );
  AND2_X1 U7711 ( .A1(n6522), .A2(n6521), .ZN(n6523) );
  NOR2_X1 U7712 ( .A1(n6533), .A2(n6523), .ZN(n7841) );
  NAND2_X1 U7713 ( .A1(n6782), .A2(n7841), .ZN(n6525) );
  NAND2_X1 U7714 ( .A1(n5133), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n6524) );
  NAND4_X1 U7715 ( .A1(n6527), .A2(n6526), .A3(n6525), .A4(n6524), .ZN(n10292)
         );
  INV_X1 U7716 ( .A(n10292), .ZN(n7528) );
  OR2_X1 U7717 ( .A1(n6959), .A2(n6699), .ZN(n6531) );
  OR2_X1 U7718 ( .A1(n6539), .A2(n10692), .ZN(n6528) );
  XNOR2_X1 U7719 ( .A(n6528), .B(P1_IR_REG_6__SCAN_IN), .ZN(n7178) );
  AOI22_X1 U7720 ( .A1(n8317), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n7178), .B2(
        n6529), .ZN(n6530) );
  NAND2_X1 U7721 ( .A1(n7528), .A2(n11053), .ZN(n6542) );
  AND2_X1 U7722 ( .A1(n7828), .A2(n6542), .ZN(n6532) );
  NAND2_X1 U7723 ( .A1(n7829), .A2(n6532), .ZN(n7521) );
  NAND2_X1 U7724 ( .A1(n6580), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n6538) );
  NAND2_X1 U7725 ( .A1(n6520), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n6537) );
  NAND2_X1 U7726 ( .A1(n5132), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n6536) );
  NAND2_X1 U7727 ( .A1(n6533), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n6551) );
  OR2_X1 U7728 ( .A1(n6533), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n6534) );
  NAND2_X1 U7729 ( .A1(n6551), .A2(n6534), .ZN(n7637) );
  OR2_X1 U7730 ( .A1(n6773), .A2(n7637), .ZN(n6535) );
  NAND2_X1 U7731 ( .A1(n6539), .A2(n9772), .ZN(n6547) );
  NAND2_X1 U7732 ( .A1(n6547), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6540) );
  XNOR2_X1 U7733 ( .A(n6540), .B(P1_IR_REG_7__SCAN_IN), .ZN(n7192) );
  AOI22_X1 U7734 ( .A1(n8317), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n7192), .B2(
        n6529), .ZN(n6541) );
  INV_X1 U7735 ( .A(n6542), .ZN(n6543) );
  NAND2_X1 U7736 ( .A1(n11053), .A2(n10292), .ZN(n7524) );
  AND2_X1 U7737 ( .A1(n8849), .A2(n7520), .ZN(n6544) );
  NAND2_X1 U7738 ( .A1(n7521), .A2(n6544), .ZN(n7522) );
  OR2_X1 U7739 ( .A1(n5297), .A2(n7639), .ZN(n6545) );
  NAND2_X1 U7740 ( .A1(n7522), .A2(n6545), .ZN(n7709) );
  NAND2_X1 U7741 ( .A1(n6558), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6548) );
  XNOR2_X1 U7742 ( .A(n6548), .B(P1_IR_REG_8__SCAN_IN), .ZN(n7453) );
  AOI22_X1 U7743 ( .A1(n8317), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n7453), .B2(
        n6529), .ZN(n6549) );
  NAND2_X1 U7744 ( .A1(n6520), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n6556) );
  NAND2_X1 U7745 ( .A1(n6580), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n6555) );
  NAND2_X1 U7746 ( .A1(n5133), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n6554) );
  NAND2_X1 U7747 ( .A1(n6551), .A2(n6550), .ZN(n6552) );
  NAND2_X1 U7748 ( .A1(n6562), .A2(n6552), .ZN(n10099) );
  OR2_X1 U7749 ( .A1(n6773), .A2(n10099), .ZN(n6553) );
  NAND2_X1 U7750 ( .A1(n10101), .A2(n10170), .ZN(n8936) );
  NAND2_X1 U7751 ( .A1(n8855), .A2(n8936), .ZN(n8853) );
  OR2_X1 U7752 ( .A1(n10101), .A2(n10291), .ZN(n6557) );
  NAND2_X1 U7753 ( .A1(n6984), .A2(n6546), .ZN(n6561) );
  NAND2_X1 U7754 ( .A1(n6559), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6568) );
  XNOR2_X1 U7755 ( .A(n6568), .B(P1_IR_REG_9__SCAN_IN), .ZN(n10364) );
  AOI22_X1 U7756 ( .A1(n8317), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n10364), .B2(
        n6529), .ZN(n6560) );
  NAND2_X1 U7757 ( .A1(n6580), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n6567) );
  NAND2_X1 U7758 ( .A1(n5133), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n6566) );
  AND2_X1 U7759 ( .A1(n6562), .A2(n10167), .ZN(n6563) );
  NOR2_X1 U7760 ( .A1(n6573), .A2(n6563), .ZN(n10166) );
  NAND2_X1 U7761 ( .A1(n6782), .A2(n10166), .ZN(n6565) );
  NAND2_X1 U7762 ( .A1(n6520), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n6564) );
  OR2_X1 U7763 ( .A1(n10172), .A2(n10096), .ZN(n8860) );
  NAND2_X1 U7764 ( .A1(n10172), .A2(n10096), .ZN(n8927) );
  NAND2_X1 U7765 ( .A1(n8860), .A2(n8927), .ZN(n7867) );
  INV_X1 U7766 ( .A(n10096), .ZN(n10290) );
  OR2_X1 U7767 ( .A1(n6990), .A2(n6699), .ZN(n6572) );
  INV_X1 U7768 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n6989) );
  INV_X1 U7769 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n9986) );
  NAND2_X1 U7770 ( .A1(n6568), .A2(n9986), .ZN(n6569) );
  NAND2_X1 U7771 ( .A1(n6569), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6588) );
  XNOR2_X1 U7772 ( .A(n6588), .B(P1_IR_REG_10__SCAN_IN), .ZN(n10880) );
  INV_X1 U7773 ( .A(n10880), .ZN(n7456) );
  OAI22_X1 U7774 ( .A1(n6646), .A2(n6989), .B1(n6474), .B2(n7456), .ZN(n6570)
         );
  INV_X1 U7775 ( .A(n6570), .ZN(n6571) );
  NAND2_X1 U7776 ( .A1(n6520), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n6578) );
  NAND2_X1 U7777 ( .A1(n6580), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n6577) );
  NAND2_X1 U7778 ( .A1(n5132), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n6576) );
  NOR2_X1 U7779 ( .A1(n6573), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n6574) );
  OR2_X1 U7780 ( .A1(n6581), .A2(n6574), .ZN(n10078) );
  OR2_X1 U7781 ( .A1(n6773), .A2(n10078), .ZN(n6575) );
  OR2_X1 U7782 ( .A1(n10080), .A2(n8654), .ZN(n8867) );
  NAND2_X1 U7783 ( .A1(n10080), .A2(n8654), .ZN(n8862) );
  NAND2_X1 U7784 ( .A1(n8867), .A2(n8862), .ZN(n8940) );
  OR2_X1 U7785 ( .A1(n10080), .A2(n10289), .ZN(n6579) );
  NAND2_X1 U7786 ( .A1(n6580), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n6586) );
  NAND2_X1 U7787 ( .A1(n6520), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n6585) );
  NAND2_X1 U7788 ( .A1(n5133), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n6584) );
  OR2_X1 U7789 ( .A1(n6581), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n6582) );
  NAND2_X1 U7790 ( .A1(n6600), .A2(n6582), .ZN(n10214) );
  OR2_X1 U7791 ( .A1(n6773), .A2(n10214), .ZN(n6583) );
  NAND2_X1 U7792 ( .A1(n6587), .A2(n6546), .ZN(n6592) );
  INV_X1 U7793 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n9987) );
  NAND2_X1 U7794 ( .A1(n6588), .A2(n9987), .ZN(n6589) );
  NAND2_X1 U7795 ( .A1(n6589), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6590) );
  XNOR2_X1 U7796 ( .A(n6590), .B(P1_IR_REG_11__SCAN_IN), .ZN(n10806) );
  AOI22_X1 U7797 ( .A1(n8317), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n10806), 
        .B2(n6529), .ZN(n6591) );
  NAND2_X1 U7798 ( .A1(n6592), .A2(n6591), .ZN(n8663) );
  INV_X1 U7799 ( .A(n8663), .ZN(n11087) );
  INV_X1 U7800 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n7030) );
  NOR2_X1 U7801 ( .A1(n6593), .A2(n10692), .ZN(n6594) );
  MUX2_X1 U7802 ( .A(n10692), .B(n6594), .S(P1_IR_REG_12__SCAN_IN), .Z(n6595)
         );
  OR2_X1 U7803 ( .A1(n6595), .A2(n5198), .ZN(n7463) );
  OAI22_X1 U7804 ( .A1(n6646), .A2(n7030), .B1(n6474), .B2(n7463), .ZN(n6596)
         );
  INV_X1 U7805 ( .A(n6596), .ZN(n6597) );
  NAND2_X1 U7806 ( .A1(n6580), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n6605) );
  NAND2_X1 U7807 ( .A1(n5133), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n6604) );
  NAND2_X1 U7808 ( .A1(n6520), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n6603) );
  NAND2_X1 U7809 ( .A1(n6600), .A2(n6599), .ZN(n6601) );
  NAND2_X1 U7810 ( .A1(n6606), .A2(n6601), .ZN(n10116) );
  OR2_X1 U7811 ( .A1(n6773), .A2(n10116), .ZN(n6602) );
  INV_X1 U7812 ( .A(n10213), .ZN(n10287) );
  NAND2_X1 U7813 ( .A1(n6520), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n6611) );
  NAND2_X1 U7814 ( .A1(n6580), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n6610) );
  NAND2_X1 U7815 ( .A1(n5132), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n6609) );
  AND2_X1 U7816 ( .A1(n6606), .A2(n10188), .ZN(n6607) );
  OR2_X1 U7817 ( .A1(n6614), .A2(n6607), .ZN(n7922) );
  OR2_X1 U7818 ( .A1(n6773), .A2(n7922), .ZN(n6608) );
  NAND2_X1 U7819 ( .A1(n6643), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6631) );
  XNOR2_X1 U7820 ( .A(n6631), .B(P1_IR_REG_14__SCAN_IN), .ZN(n10818) );
  AOI22_X1 U7821 ( .A1(n8317), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n10818), 
        .B2(n6529), .ZN(n6612) );
  NAND2_X1 U7822 ( .A1(n6580), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n6619) );
  NAND2_X1 U7823 ( .A1(n6520), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n6618) );
  NAND2_X1 U7824 ( .A1(n5133), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n6617) );
  OR2_X1 U7825 ( .A1(n6614), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n6615) );
  NAND2_X1 U7826 ( .A1(n6614), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n6636) );
  NAND2_X1 U7827 ( .A1(n6615), .A2(n6636), .ZN(n11148) );
  OR2_X1 U7828 ( .A1(n6773), .A2(n11148), .ZN(n6616) );
  AND2_X1 U7829 ( .A1(n11152), .A2(n10190), .ZN(n8877) );
  INV_X1 U7830 ( .A(n8877), .ZN(n8873) );
  AND2_X1 U7831 ( .A1(n11115), .A2(n11120), .ZN(n6620) );
  NAND2_X1 U7832 ( .A1(n7915), .A2(n6620), .ZN(n6626) );
  INV_X1 U7833 ( .A(n11120), .ZN(n6624) );
  OR2_X1 U7834 ( .A1(n7101), .A2(n6699), .ZN(n6623) );
  OR2_X1 U7835 ( .A1(n5198), .A2(n10692), .ZN(n6621) );
  XNOR2_X1 U7836 ( .A(n6621), .B(P1_IR_REG_13__SCAN_IN), .ZN(n10864) );
  AOI22_X1 U7837 ( .A1(n8317), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n10864), 
        .B2(n6529), .ZN(n6622) );
  OR2_X1 U7838 ( .A1(n6624), .A2(n11116), .ZN(n6625) );
  NAND2_X1 U7839 ( .A1(n6626), .A2(n6625), .ZN(n6628) );
  NAND2_X1 U7840 ( .A1(n6627), .A2(n11138), .ZN(n11118) );
  INV_X1 U7841 ( .A(n11152), .ZN(n11128) );
  NAND2_X1 U7842 ( .A1(n11152), .A2(n6629), .ZN(n6630) );
  INV_X1 U7843 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n7281) );
  NAND2_X1 U7844 ( .A1(n6631), .A2(n9995), .ZN(n6632) );
  NAND2_X1 U7845 ( .A1(n6632), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6633) );
  XNOR2_X1 U7846 ( .A(n6633), .B(P1_IR_REG_15__SCAN_IN), .ZN(n10828) );
  OAI22_X1 U7847 ( .A1(n6646), .A2(n7281), .B1(n6474), .B2(n10385), .ZN(n6634)
         );
  INV_X1 U7848 ( .A(n6634), .ZN(n6635) );
  NAND2_X1 U7849 ( .A1(n6520), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n6641) );
  NAND2_X1 U7850 ( .A1(n6580), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n6640) );
  NAND2_X1 U7851 ( .A1(n5133), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n6639) );
  OAI21_X1 U7852 ( .B1(n6637), .B2(P1_REG3_REG_15__SCAN_IN), .A(n6650), .ZN(
        n10264) );
  OR2_X1 U7853 ( .A1(n6773), .A2(n10264), .ZN(n6638) );
  NAND2_X1 U7854 ( .A1(n10267), .A2(n11136), .ZN(n8878) );
  INV_X1 U7855 ( .A(n10267), .ZN(n11166) );
  NAND2_X1 U7856 ( .A1(n7329), .A2(n6546), .ZN(n6649) );
  INV_X1 U7857 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n7330) );
  NAND2_X1 U7858 ( .A1(n6657), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6645) );
  XNOR2_X1 U7859 ( .A(n6645), .B(P1_IR_REG_16__SCAN_IN), .ZN(n10403) );
  INV_X1 U7860 ( .A(n10403), .ZN(n10380) );
  OAI22_X1 U7861 ( .A1(n6646), .A2(n7330), .B1(n6474), .B2(n10380), .ZN(n6647)
         );
  INV_X1 U7862 ( .A(n6647), .ZN(n6648) );
  NAND2_X1 U7863 ( .A1(n6520), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n6656) );
  OAI21_X1 U7864 ( .B1(n6651), .B2(P1_REG3_REG_16__SCAN_IN), .A(n6665), .ZN(
        n10138) );
  INV_X1 U7865 ( .A(n10138), .ZN(n8219) );
  NAND2_X1 U7866 ( .A1(n6782), .A2(n8219), .ZN(n6655) );
  NAND2_X1 U7867 ( .A1(n5133), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n6654) );
  INV_X1 U7868 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n10375) );
  OR2_X1 U7869 ( .A1(n6652), .A2(n10375), .ZN(n6653) );
  OR2_X1 U7870 ( .A1(n10646), .A2(n10258), .ZN(n9020) );
  NAND2_X1 U7871 ( .A1(n10646), .A2(n10258), .ZN(n9019) );
  NAND2_X1 U7872 ( .A1(n9020), .A2(n9019), .ZN(n8949) );
  NAND2_X1 U7873 ( .A1(n8216), .A2(n8949), .ZN(n8215) );
  INV_X1 U7874 ( .A(n10646), .ZN(n8221) );
  NAND2_X1 U7875 ( .A1(n8215), .A2(n5731), .ZN(n8177) );
  NAND2_X1 U7876 ( .A1(n7406), .A2(n6546), .ZN(n6661) );
  NAND2_X1 U7877 ( .A1(n6658), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6659) );
  XNOR2_X1 U7878 ( .A(n6659), .B(P1_IR_REG_17__SCAN_IN), .ZN(n10840) );
  AOI22_X1 U7879 ( .A1(n8317), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n10840), 
        .B2(n6529), .ZN(n6660) );
  NAND2_X1 U7880 ( .A1(n6520), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n6669) );
  NAND2_X1 U7881 ( .A1(n6580), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n6668) );
  INV_X1 U7882 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n6664) );
  INV_X1 U7883 ( .A(n6673), .ZN(n6663) );
  AOI21_X1 U7884 ( .B1(n6665), .B2(n6664), .A(n6663), .ZN(n10149) );
  NAND2_X1 U7885 ( .A1(n6782), .A2(n10149), .ZN(n6667) );
  NAND2_X1 U7886 ( .A1(n5132), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n6666) );
  NAND2_X1 U7887 ( .A1(n8722), .A2(n10237), .ZN(n8884) );
  INV_X1 U7888 ( .A(n10237), .ZN(n10284) );
  XNOR2_X1 U7889 ( .A(n6680), .B(P1_IR_REG_18__SCAN_IN), .ZN(n10854) );
  AOI22_X1 U7890 ( .A1(n8317), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n10854), 
        .B2(n6529), .ZN(n6671) );
  NAND2_X1 U7891 ( .A1(n6580), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n6677) );
  NAND2_X1 U7892 ( .A1(n5133), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n6676) );
  AOI21_X1 U7893 ( .B1(n10232), .B2(n6673), .A(n6685), .ZN(n10231) );
  NAND2_X1 U7894 ( .A1(n6782), .A2(n10231), .ZN(n6675) );
  NAND2_X1 U7895 ( .A1(n6520), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n6674) );
  OR2_X1 U7896 ( .A1(n10636), .A2(n10569), .ZN(n8887) );
  NAND2_X1 U7897 ( .A1(n10636), .A2(n10569), .ZN(n8889) );
  INV_X1 U7898 ( .A(n10569), .ZN(n10283) );
  NAND2_X1 U7899 ( .A1(n7657), .A2(n6546), .ZN(n6684) );
  NAND2_X1 U7900 ( .A1(n6680), .A2(n6679), .ZN(n6681) );
  XNOR2_X2 U7901 ( .A(n6682), .B(P1_IR_REG_19__SCAN_IN), .ZN(n7110) );
  AOI22_X1 U7902 ( .A1(n8317), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n7110), .B2(
        n6529), .ZN(n6683) );
  NAND2_X1 U7903 ( .A1(n6580), .A2(P1_REG1_REG_19__SCAN_IN), .ZN(n6689) );
  NAND2_X1 U7904 ( .A1(n6520), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n6688) );
  NAND2_X1 U7905 ( .A1(n5132), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n6687) );
  OAI21_X1 U7906 ( .B1(P1_REG3_REG_19__SCAN_IN), .B2(n6685), .A(n6691), .ZN(
        n10581) );
  OR2_X1 U7907 ( .A1(n6773), .A2(n10581), .ZN(n6686) );
  NOR2_X1 U7908 ( .A1(n10579), .A2(n10282), .ZN(n6690) );
  NAND2_X1 U7909 ( .A1(n6580), .A2(P1_REG1_REG_20__SCAN_IN), .ZN(n6695) );
  NAND2_X1 U7910 ( .A1(n5132), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n6694) );
  INV_X1 U7911 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n10178) );
  AOI21_X1 U7912 ( .B1(n10178), .B2(n6691), .A(n6702), .ZN(n10556) );
  NAND2_X1 U7913 ( .A1(n6782), .A2(n10556), .ZN(n6693) );
  NAND2_X1 U7914 ( .A1(n6520), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n6692) );
  NAND2_X1 U7915 ( .A1(n7905), .A2(n6546), .ZN(n6697) );
  NAND2_X1 U7916 ( .A1(n8317), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n6696) );
  NAND2_X1 U7917 ( .A1(n10626), .A2(n10568), .ZN(n10525) );
  NAND2_X1 U7918 ( .A1(n10526), .A2(n10525), .ZN(n10546) );
  INV_X1 U7919 ( .A(n10546), .ZN(n10548) );
  INV_X1 U7920 ( .A(n10568), .ZN(n10281) );
  NAND2_X1 U7921 ( .A1(n8317), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n6700) );
  NAND2_X1 U7922 ( .A1(n6520), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n6706) );
  NAND2_X1 U7923 ( .A1(n6580), .A2(P1_REG1_REG_21__SCAN_IN), .ZN(n6705) );
  NAND2_X1 U7924 ( .A1(n5133), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n6704) );
  NAND2_X1 U7925 ( .A1(n6702), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n6711) );
  OAI21_X1 U7926 ( .B1(P1_REG3_REG_21__SCAN_IN), .B2(n6702), .A(n6711), .ZN(
        n10539) );
  OR2_X1 U7927 ( .A1(n6773), .A2(n10539), .ZN(n6703) );
  NAND2_X1 U7928 ( .A1(n10538), .A2(n10551), .ZN(n8897) );
  INV_X1 U7929 ( .A(n10528), .ZN(n10523) );
  INV_X1 U7930 ( .A(n10551), .ZN(n10280) );
  NAND2_X1 U7931 ( .A1(n6707), .A2(n10551), .ZN(n6708) );
  NAND2_X1 U7932 ( .A1(n10522), .A2(n6708), .ZN(n10507) );
  NAND2_X1 U7933 ( .A1(n8317), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n6709) );
  NAND2_X1 U7934 ( .A1(n6580), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n6716) );
  NAND2_X1 U7935 ( .A1(n6520), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n6715) );
  NAND2_X1 U7936 ( .A1(n5133), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n6714) );
  OAI21_X1 U7937 ( .B1(P1_REG3_REG_22__SCAN_IN), .B2(n6712), .A(n6720), .ZN(
        n10509) );
  OR2_X1 U7938 ( .A1(n6773), .A2(n10509), .ZN(n6713) );
  OR2_X1 U7939 ( .A1(n10613), .A2(n10531), .ZN(n8832) );
  NAND2_X1 U7940 ( .A1(n10613), .A2(n10531), .ZN(n8831) );
  NAND2_X1 U7941 ( .A1(n8832), .A2(n8831), .ZN(n10513) );
  INV_X1 U7942 ( .A(n10531), .ZN(n10279) );
  NAND2_X1 U7943 ( .A1(n8032), .A2(n6546), .ZN(n6719) );
  NAND2_X1 U7944 ( .A1(n8317), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n6718) );
  NAND2_X1 U7945 ( .A1(n6580), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n6725) );
  NAND2_X1 U7946 ( .A1(n5133), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n6724) );
  NAND2_X1 U7947 ( .A1(n6520), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n6723) );
  OAI21_X1 U7948 ( .B1(P1_REG3_REG_23__SCAN_IN), .B2(n6721), .A(n6730), .ZN(
        n10499) );
  OR2_X1 U7949 ( .A1(n6773), .A2(n10499), .ZN(n6722) );
  INV_X1 U7950 ( .A(n10515), .ZN(n10278) );
  NOR2_X1 U7951 ( .A1(n10068), .A2(n10278), .ZN(n6726) );
  NAND2_X1 U7952 ( .A1(n8140), .A2(n6546), .ZN(n6728) );
  NAND2_X1 U7953 ( .A1(n8317), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n6727) );
  NAND2_X1 U7954 ( .A1(n6580), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n6735) );
  NAND2_X1 U7955 ( .A1(n5133), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n6734) );
  NAND2_X1 U7956 ( .A1(n6520), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n6733) );
  NAND2_X1 U7957 ( .A1(n6731), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n6739) );
  OAI21_X1 U7958 ( .B1(P1_REG3_REG_24__SCAN_IN), .B2(n6731), .A(n6739), .ZN(
        n10488) );
  OR2_X1 U7959 ( .A1(n6773), .A2(n10488), .ZN(n6732) );
  INV_X1 U7960 ( .A(n10496), .ZN(n10277) );
  INV_X1 U7961 ( .A(n10603), .ZN(n10480) );
  AOI21_X1 U7962 ( .B1(n6736), .B2(n5728), .A(n5202), .ZN(n10457) );
  NAND2_X1 U7963 ( .A1(n8317), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n6737) );
  NAND2_X1 U7964 ( .A1(n6520), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n6744) );
  NAND2_X1 U7965 ( .A1(n6580), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n6743) );
  NAND2_X1 U7966 ( .A1(n5132), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n6742) );
  INV_X1 U7967 ( .A(n6751), .ZN(n6753) );
  OAI21_X1 U7968 ( .B1(P1_REG3_REG_25__SCAN_IN), .B2(n6740), .A(n6753), .ZN(
        n10469) );
  OR2_X1 U7969 ( .A1(n6773), .A2(n10469), .ZN(n6741) );
  INV_X1 U7970 ( .A(n10484), .ZN(n10276) );
  NAND2_X1 U7971 ( .A1(n10457), .A2(n6746), .ZN(n6748) );
  NAND2_X1 U7972 ( .A1(n6748), .A2(n6747), .ZN(n10440) );
  NAND2_X1 U7973 ( .A1(n8280), .A2(n6546), .ZN(n6750) );
  NAND2_X1 U7974 ( .A1(n8317), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n6749) );
  NAND2_X1 U7975 ( .A1(n6520), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n6758) );
  NAND2_X1 U7976 ( .A1(n6580), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n6757) );
  NAND2_X1 U7977 ( .A1(n5133), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n6756) );
  INV_X1 U7978 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n6752) );
  NAND2_X1 U7979 ( .A1(n6753), .A2(n6752), .ZN(n6754) );
  NAND2_X1 U7980 ( .A1(n6770), .A2(n6754), .ZN(n10247) );
  OR2_X1 U7981 ( .A1(n6773), .A2(n10247), .ZN(n6755) );
  NAND2_X1 U7982 ( .A1(n10450), .A2(n10462), .ZN(n8905) );
  INV_X1 U7983 ( .A(n10462), .ZN(n10275) );
  NAND2_X1 U7984 ( .A1(n8289), .A2(n6546), .ZN(n6760) );
  NAND2_X1 U7985 ( .A1(n8317), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n6759) );
  NAND2_X1 U7986 ( .A1(n6520), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n6764) );
  NAND2_X1 U7987 ( .A1(n6580), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n6763) );
  XNOR2_X1 U7988 ( .A(n6770), .B(P1_REG3_REG_27__SCAN_IN), .ZN(n10429) );
  NAND2_X1 U7989 ( .A1(n6782), .A2(n10429), .ZN(n6762) );
  NAND2_X1 U7990 ( .A1(n5133), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n6761) );
  NAND2_X1 U7991 ( .A1(n10434), .A2(n10446), .ZN(n9044) );
  NAND2_X1 U7992 ( .A1(n8293), .A2(n6546), .ZN(n6766) );
  NAND2_X1 U7993 ( .A1(n8317), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n6765) );
  NAND2_X1 U7994 ( .A1(n6520), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n6777) );
  NAND2_X1 U7995 ( .A1(n6580), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n6776) );
  NAND2_X1 U7996 ( .A1(n5132), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n6775) );
  INV_X1 U7997 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n6768) );
  INV_X1 U7998 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n6767) );
  OAI21_X1 U7999 ( .B1(n6770), .B2(n6768), .A(n6767), .ZN(n6772) );
  NAND2_X1 U8000 ( .A1(P1_REG3_REG_28__SCAN_IN), .A2(P1_REG3_REG_27__SCAN_IN), 
        .ZN(n6769) );
  NOR2_X1 U8001 ( .A1(n6770), .A2(n6769), .ZN(n8335) );
  INV_X1 U8002 ( .A(n8335), .ZN(n6771) );
  NAND2_X1 U8003 ( .A1(n6772), .A2(n6771), .ZN(n8814) );
  OR2_X1 U8004 ( .A1(n6773), .A2(n8814), .ZN(n6774) );
  NOR2_X1 U8005 ( .A1(n8819), .A2(n10426), .ZN(n8828) );
  INV_X1 U8006 ( .A(n8828), .ZN(n6778) );
  NAND2_X1 U8007 ( .A1(n8819), .A2(n10426), .ZN(n9045) );
  NAND2_X1 U8008 ( .A1(n6778), .A2(n9045), .ZN(n8957) );
  NAND2_X1 U8009 ( .A1(n6779), .A2(n6546), .ZN(n6781) );
  NAND2_X1 U8010 ( .A1(n8317), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n6780) );
  NAND2_X1 U8011 ( .A1(n6520), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n6786) );
  NAND2_X1 U8012 ( .A1(n6580), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n6785) );
  NAND2_X1 U8013 ( .A1(n6782), .A2(n8335), .ZN(n6784) );
  NAND2_X1 U8014 ( .A1(n5133), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n6783) );
  NAND2_X1 U8015 ( .A1(n8334), .A2(n8816), .ZN(n8825) );
  XNOR2_X1 U8016 ( .A(n6787), .B(n8961), .ZN(n8333) );
  INV_X1 U8017 ( .A(n6789), .ZN(n6790) );
  NAND2_X1 U8018 ( .A1(n6790), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6791) );
  NOR2_X1 U8019 ( .A1(n9062), .A2(n7110), .ZN(n6797) );
  OR2_X1 U8020 ( .A1(n10692), .A2(n9796), .ZN(n6792) );
  XNOR2_X2 U8021 ( .A(n6795), .B(n6794), .ZN(n6814) );
  OAI21_X1 U8022 ( .B1(n6797), .B2(n7107), .A(n5278), .ZN(n6798) );
  AND2_X1 U8023 ( .A1(n7117), .A2(n7107), .ZN(n7202) );
  OR2_X1 U8024 ( .A1(n8971), .A2(n9059), .ZN(n7799) );
  NAND2_X1 U8025 ( .A1(n8333), .A2(n11168), .ZN(n6830) );
  NAND2_X1 U8026 ( .A1(n10603), .A2(n10496), .ZN(n9035) );
  NAND2_X1 U8027 ( .A1(n8897), .A2(n10525), .ZN(n9031) );
  NAND2_X1 U8028 ( .A1(n8680), .A2(n11138), .ZN(n11130) );
  INV_X1 U8029 ( .A(n11130), .ZN(n6799) );
  NOR2_X1 U8030 ( .A1(n11120), .A2(n6799), .ZN(n6809) );
  NOR2_X1 U8031 ( .A1(n10297), .A2(n7725), .ZN(n7025) );
  NAND2_X1 U8032 ( .A1(n8928), .A2(n7025), .ZN(n6801) );
  INV_X1 U8033 ( .A(n7729), .ZN(n10987) );
  OR2_X1 U8034 ( .A1(n11000), .A2(n10987), .ZN(n6800) );
  NAND2_X1 U8035 ( .A1(n6801), .A2(n6800), .ZN(n10998) );
  INV_X1 U8036 ( .A(n10997), .ZN(n6802) );
  NAND2_X1 U8037 ( .A1(n10998), .A2(n6802), .ZN(n8833) );
  NAND2_X1 U8038 ( .A1(n8833), .A2(n8988), .ZN(n7644) );
  INV_X1 U8039 ( .A(n8934), .ZN(n7645) );
  NAND2_X1 U8040 ( .A1(n7644), .A2(n7645), .ZN(n7643) );
  NAND2_X1 U8041 ( .A1(n7643), .A2(n8993), .ZN(n7810) );
  OR2_X1 U8042 ( .A1(n10294), .A2(n11042), .ZN(n8842) );
  INV_X1 U8043 ( .A(n8842), .ZN(n6803) );
  AND2_X1 U8044 ( .A1(n10294), .A2(n11042), .ZN(n8992) );
  NOR2_X1 U8045 ( .A1(n8932), .A2(n8992), .ZN(n6804) );
  NAND2_X1 U8046 ( .A1(n7414), .A2(n8843), .ZN(n7827) );
  INV_X1 U8047 ( .A(n8998), .ZN(n8933) );
  NAND2_X1 U8048 ( .A1(n8860), .A2(n8855), .ZN(n6807) );
  INV_X1 U8049 ( .A(n7524), .ZN(n8848) );
  AND2_X1 U8050 ( .A1(n8936), .A2(n8935), .ZN(n6806) );
  OR2_X1 U8051 ( .A1(n6807), .A2(n6806), .ZN(n6808) );
  AND2_X1 U8052 ( .A1(n6808), .A2(n8927), .ZN(n9003) );
  INV_X1 U8053 ( .A(n8940), .ZN(n7696) );
  NAND2_X2 U8054 ( .A1(n7697), .A2(n7696), .ZN(n7891) );
  NAND2_X1 U8055 ( .A1(n8663), .A2(n10119), .ZN(n8865) );
  AND2_X1 U8056 ( .A1(n8865), .A2(n8862), .ZN(n9005) );
  OR2_X1 U8057 ( .A1(n8670), .A2(n10213), .ZN(n8872) );
  OR2_X1 U8058 ( .A1(n8663), .A2(n10119), .ZN(n8864) );
  AND2_X1 U8059 ( .A1(n8872), .A2(n8864), .ZN(n8985) );
  NAND2_X1 U8060 ( .A1(n8670), .A2(n10213), .ZN(n8874) );
  AND2_X1 U8061 ( .A1(n11116), .A2(n11115), .ZN(n8875) );
  INV_X1 U8062 ( .A(n8875), .ZN(n9011) );
  INV_X1 U8063 ( .A(n8949), .ZN(n8224) );
  NAND2_X1 U8064 ( .A1(n8223), .A2(n8224), .ZN(n8222) );
  XNOR2_X1 U8065 ( .A(n10579), .B(n10282), .ZN(n10564) );
  NAND2_X1 U8066 ( .A1(n10565), .A2(n10564), .ZN(n6810) );
  NAND2_X1 U8067 ( .A1(n10579), .A2(n10550), .ZN(n8983) );
  OR2_X1 U8068 ( .A1(n10068), .A2(n10515), .ZN(n8901) );
  NAND2_X1 U8069 ( .A1(n10068), .A2(n10515), .ZN(n8977) );
  NAND2_X1 U8070 ( .A1(n10493), .A2(n8977), .ZN(n10482) );
  OR2_X1 U8071 ( .A1(n10468), .A2(n10484), .ZN(n9038) );
  NAND2_X1 U8072 ( .A1(n10468), .A2(n10484), .ZN(n8908) );
  INV_X1 U8073 ( .A(n9038), .ZN(n10443) );
  INV_X1 U8074 ( .A(n9040), .ZN(n6881) );
  NAND2_X1 U8075 ( .A1(n6882), .A2(n9045), .ZN(n6811) );
  XNOR2_X1 U8076 ( .A(n6811), .B(n8961), .ZN(n6827) );
  OR2_X1 U8077 ( .A1(n6812), .A2(n9062), .ZN(n6815) );
  INV_X1 U8078 ( .A(n6813), .ZN(n7122) );
  INV_X1 U8079 ( .A(n10426), .ZN(n10273) );
  NAND2_X1 U8080 ( .A1(n6816), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6819) );
  INV_X1 U8081 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n10018) );
  NAND2_X1 U8082 ( .A1(n6819), .A2(n10018), .ZN(n6817) );
  NAND2_X1 U8083 ( .A1(n6817), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6818) );
  NAND2_X2 U8084 ( .A1(n7117), .A2(n10705), .ZN(n11135) );
  XNOR2_X1 U8085 ( .A(n6819), .B(P1_IR_REG_27__SCAN_IN), .ZN(n8291) );
  AND2_X1 U8086 ( .A1(n8291), .A2(P1_B_REG_SCAN_IN), .ZN(n6820) );
  NOR2_X1 U8087 ( .A1(n11135), .A2(n6820), .ZN(n8324) );
  INV_X1 U8088 ( .A(P1_REG2_REG_30__SCAN_IN), .ZN(n6823) );
  NAND2_X1 U8089 ( .A1(n6580), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n6822) );
  NAND2_X1 U8090 ( .A1(n5133), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n6821) );
  OAI211_X1 U8091 ( .C1(n6824), .C2(n6823), .A(n6822), .B(n6821), .ZN(n10272)
         );
  AOI21_X2 U8092 ( .B1(n6827), .B2(n10566), .A(n6826), .ZN(n8342) );
  AND2_X1 U8093 ( .A1(n7819), .A2(n7557), .ZN(n7840) );
  NAND2_X1 U8094 ( .A1(n7840), .A2(n11053), .ZN(n7839) );
  INV_X1 U8095 ( .A(n10080), .ZN(n11077) );
  INV_X1 U8096 ( .A(n10172), .ZN(n11069) );
  NAND2_X1 U8097 ( .A1(n10656), .A2(n10449), .ZN(n6886) );
  NAND2_X1 U8098 ( .A1(n7201), .A2(n6813), .ZN(n10577) );
  AOI21_X1 U8099 ( .B1(n10985), .B2(n8334), .A(n8339), .ZN(n6828) );
  NAND2_X1 U8100 ( .A1(n6830), .A2(n6829), .ZN(n10652) );
  NAND2_X1 U8101 ( .A1(n7201), .A2(n7108), .ZN(n7125) );
  NAND2_X1 U8102 ( .A1(n8164), .A2(P1_B_REG_SCAN_IN), .ZN(n6838) );
  NAND2_X1 U8103 ( .A1(n6835), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6837) );
  MUX2_X1 U8104 ( .A(P1_B_REG_SCAN_IN), .B(n6838), .S(n8167), .Z(n6841) );
  INV_X1 U8105 ( .A(n6859), .ZN(n8281) );
  NAND2_X1 U8106 ( .A1(n8281), .A2(n8164), .ZN(n10690) );
  OAI21_X1 U8107 ( .B1(n10688), .B2(P1_D_REG_1__SCAN_IN), .A(n10690), .ZN(
        n7118) );
  NOR2_X1 U8108 ( .A1(n8164), .A2(n8167), .ZN(n6844) );
  NAND2_X2 U8109 ( .A1(n6844), .A2(n6859), .ZN(n7333) );
  NOR4_X1 U8110 ( .A1(P1_D_REG_18__SCAN_IN), .A2(P1_D_REG_17__SCAN_IN), .A3(
        P1_D_REG_16__SCAN_IN), .A4(P1_D_REG_15__SCAN_IN), .ZN(n6849) );
  NOR4_X1 U8111 ( .A1(P1_D_REG_20__SCAN_IN), .A2(P1_D_REG_22__SCAN_IN), .A3(
        P1_D_REG_21__SCAN_IN), .A4(P1_D_REG_19__SCAN_IN), .ZN(n6848) );
  NOR4_X1 U8112 ( .A1(P1_D_REG_10__SCAN_IN), .A2(P1_D_REG_9__SCAN_IN), .A3(
        P1_D_REG_8__SCAN_IN), .A4(P1_D_REG_5__SCAN_IN), .ZN(n6847) );
  NOR4_X1 U8113 ( .A1(P1_D_REG_14__SCAN_IN), .A2(P1_D_REG_13__SCAN_IN), .A3(
        P1_D_REG_12__SCAN_IN), .A4(P1_D_REG_11__SCAN_IN), .ZN(n6846) );
  NAND4_X1 U8114 ( .A1(n6849), .A2(n6848), .A3(n6847), .A4(n6846), .ZN(n6856)
         );
  NOR2_X1 U8115 ( .A1(P1_D_REG_3__SCAN_IN), .A2(P1_D_REG_2__SCAN_IN), .ZN(
        n6853) );
  NOR4_X1 U8116 ( .A1(P1_D_REG_7__SCAN_IN), .A2(P1_D_REG_6__SCAN_IN), .A3(
        P1_D_REG_4__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n6852) );
  NOR4_X1 U8117 ( .A1(P1_D_REG_26__SCAN_IN), .A2(P1_D_REG_25__SCAN_IN), .A3(
        P1_D_REG_24__SCAN_IN), .A4(P1_D_REG_23__SCAN_IN), .ZN(n6851) );
  NOR4_X1 U8118 ( .A1(P1_D_REG_30__SCAN_IN), .A2(P1_D_REG_29__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_27__SCAN_IN), .ZN(n6850) );
  NAND4_X1 U8119 ( .A1(n6853), .A2(n6852), .A3(n6851), .A4(n6850), .ZN(n6855)
         );
  INV_X1 U8120 ( .A(n10688), .ZN(n6854) );
  OAI21_X1 U8121 ( .B1(n6856), .B2(n6855), .A(n6854), .ZN(n7119) );
  INV_X1 U8122 ( .A(n7107), .ZN(n6857) );
  NAND2_X1 U8123 ( .A1(n6857), .A2(n7117), .ZN(n7130) );
  INV_X1 U8124 ( .A(n8167), .ZN(n6858) );
  INV_X1 U8125 ( .A(n7206), .ZN(n7120) );
  NAND2_X1 U8126 ( .A1(n10652), .A2(n11171), .ZN(n6862) );
  INV_X1 U8127 ( .A(n11171), .ZN(n6860) );
  NAND2_X1 U8128 ( .A1(n6860), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n6861) );
  NAND2_X1 U8129 ( .A1(n6862), .A2(n6861), .ZN(P1_U3551) );
  OR2_X1 U8130 ( .A1(n8624), .A2(n6863), .ZN(n6864) );
  INV_X1 U8131 ( .A(n6865), .ZN(n6868) );
  AND2_X1 U8132 ( .A1(n9609), .A2(n6866), .ZN(n6867) );
  NAND2_X1 U8133 ( .A1(n6868), .A2(n6867), .ZN(n7086) );
  INV_X1 U8134 ( .A(n6869), .ZN(n6870) );
  NAND2_X1 U8135 ( .A1(n7081), .A2(n7083), .ZN(n6872) );
  OAI21_X1 U8136 ( .B1(n6897), .B2(n8057), .A(n7080), .ZN(n6871) );
  NAND2_X1 U8137 ( .A1(n6872), .A2(n6871), .ZN(n6873) );
  NAND2_X1 U8138 ( .A1(n9572), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n6875) );
  NAND2_X1 U8139 ( .A1(n6883), .A2(n6882), .ZN(n6885) );
  OAI22_X1 U8140 ( .A1(n10446), .A2(n11137), .B1(n8816), .B2(n11135), .ZN(
        n6884) );
  AOI21_X1 U8141 ( .B1(n6885), .B2(n10566), .A(n6884), .ZN(n8346) );
  INV_X1 U8142 ( .A(n6886), .ZN(n10432) );
  OAI211_X1 U8143 ( .C1(n8807), .C2(n10432), .A(n11126), .B(n6887), .ZN(n8343)
         );
  NAND2_X1 U8144 ( .A1(n5174), .A2(n5737), .ZN(P1_U3550) );
  NAND2_X1 U8145 ( .A1(n11175), .A2(n10985), .ZN(n10685) );
  INV_X2 U8146 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  NOR2_X1 U8147 ( .A1(n7333), .A2(P1_U3086), .ZN(n6890) );
  INV_X1 U8148 ( .A(n6947), .ZN(n6891) );
  NAND2_X1 U8149 ( .A1(n8618), .A2(n7012), .ZN(n6892) );
  NAND2_X1 U8150 ( .A1(n6892), .A2(n7011), .ZN(n7008) );
  NAND2_X1 U8151 ( .A1(n7008), .A2(n6893), .ZN(n6894) );
  NAND2_X1 U8152 ( .A1(n6894), .A2(P2_STATE_REG_SCAN_IN), .ZN(P2_U3150) );
  NAND2_X1 U8153 ( .A1(n6897), .A2(n8624), .ZN(n6898) );
  XNOR2_X1 U8154 ( .A(n7673), .B(n6905), .ZN(n7681) );
  XOR2_X1 U8155 ( .A(n9255), .B(n7681), .Z(n6918) );
  XNOR2_X1 U8156 ( .A(n7579), .B(n6905), .ZN(n6913) );
  XNOR2_X1 U8157 ( .A(n6905), .B(n6899), .ZN(n6900) );
  NAND2_X1 U8158 ( .A1(n6900), .A2(n7317), .ZN(n6903) );
  INV_X1 U8159 ( .A(n6900), .ZN(n6901) );
  NAND2_X1 U8160 ( .A1(n6901), .A2(n9259), .ZN(n6902) );
  NAND2_X1 U8161 ( .A1(n6903), .A2(n6902), .ZN(n7066) );
  AOI21_X1 U8162 ( .B1(n9098), .B2(n7215), .A(n7296), .ZN(n7065) );
  NOR2_X1 U8163 ( .A1(n7066), .A2(n7065), .ZN(n7064) );
  INV_X1 U8164 ( .A(n6903), .ZN(n6904) );
  XNOR2_X1 U8165 ( .A(n6905), .B(n7223), .ZN(n6907) );
  XNOR2_X1 U8166 ( .A(n6907), .B(n6908), .ZN(n7220) );
  INV_X1 U8167 ( .A(n6907), .ZN(n6909) );
  NAND2_X1 U8168 ( .A1(n6909), .A2(n6908), .ZN(n6910) );
  XNOR2_X1 U8169 ( .A(n6905), .B(n7587), .ZN(n6911) );
  NAND2_X1 U8170 ( .A1(n6911), .A2(n7478), .ZN(n6912) );
  OAI21_X1 U8171 ( .B1(n6911), .B2(n7478), .A(n6912), .ZN(n7320) );
  INV_X1 U8172 ( .A(n6912), .ZN(n7386) );
  XNOR2_X1 U8173 ( .A(n6913), .B(n9256), .ZN(n7385) );
  INV_X1 U8174 ( .A(n6933), .ZN(n6925) );
  OAI22_X1 U8175 ( .A1(n6915), .A2(n6928), .B1(n6925), .B2(n6914), .ZN(n6916)
         );
  AOI211_X1 U8176 ( .C1(n6918), .C2(n6917), .A(n9224), .B(n7683), .ZN(n6941)
         );
  NAND2_X1 U8177 ( .A1(n6919), .A2(n6928), .ZN(n6923) );
  NAND2_X1 U8178 ( .A1(n7012), .A2(n7011), .ZN(n6920) );
  AOI21_X1 U8179 ( .B1(n6921), .B2(n6925), .A(n6920), .ZN(n6922) );
  NAND3_X1 U8180 ( .A1(n6923), .A2(n6922), .A3(n7081), .ZN(n6924) );
  NAND2_X1 U8181 ( .A1(n6924), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6927) );
  OR2_X1 U8182 ( .A1(n7091), .A2(n7089), .ZN(n6935) );
  INV_X1 U8183 ( .A(n6935), .ZN(n8628) );
  NAND2_X1 U8184 ( .A1(n8628), .A2(n6925), .ZN(n6926) );
  NOR2_X1 U8185 ( .A1(n9217), .A2(n7516), .ZN(n6940) );
  NAND2_X1 U8186 ( .A1(n6928), .A2(n6895), .ZN(n6929) );
  AND2_X1 U8187 ( .A1(n7673), .A2(n9219), .ZN(n6939) );
  NAND2_X1 U8188 ( .A1(n6933), .A2(n6930), .ZN(n6931) );
  NAND2_X1 U8189 ( .A1(n6933), .A2(n6932), .ZN(n6934) );
  NAND2_X1 U8190 ( .A1(n9229), .A2(n9256), .ZN(n6937) );
  INV_X1 U8191 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n6936) );
  OR2_X1 U8192 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6936), .ZN(n7254) );
  OAI211_X1 U8193 ( .C1(n7774), .C2(n9231), .A(n6937), .B(n7254), .ZN(n6938)
         );
  OR4_X1 U8194 ( .A1(n6941), .A2(n6940), .A3(n6939), .A4(n6938), .ZN(P2_U3179)
         );
  INV_X2 U8195 ( .A(n9621), .ZN(n9614) );
  NAND2_X1 U8196 ( .A1(n8306), .A2(P2_U3151), .ZN(n9619) );
  OAI222_X1 U8197 ( .A1(n9614), .A2(n6942), .B1(n7050), .B2(P2_U3151), .C1(
        n9619), .C2(n6949), .ZN(P2_U3294) );
  NAND2_X1 U8198 ( .A1(n8306), .A2(P1_U3086), .ZN(n10701) );
  OAI222_X1 U8199 ( .A1(P1_U3086), .A2(n7148), .B1(n10704), .B2(n6944), .C1(
        n6943), .C2(n10701), .ZN(P1_U3352) );
  OAI222_X1 U8200 ( .A1(n9614), .A2(n5757), .B1(n7259), .B2(P2_U3151), .C1(
        n9619), .C2(n6944), .ZN(P2_U3292) );
  INV_X1 U8201 ( .A(n9619), .ZN(n9622) );
  OAI222_X1 U8202 ( .A1(n9109), .A2(n6953), .B1(n7268), .B2(P2_U3151), .C1(
        n6945), .C2(n9614), .ZN(P2_U3291) );
  NAND2_X1 U8203 ( .A1(n9609), .A2(n6946), .ZN(n6960) );
  AND2_X1 U8204 ( .A1(n6947), .A2(n6406), .ZN(n6948) );
  AOI22_X1 U8205 ( .A1(n6960), .A2(n6405), .B1(n6948), .B2(n8282), .ZN(
        P2_U3376) );
  OAI222_X1 U8206 ( .A1(n10701), .A2(n6950), .B1(n10704), .B2(n6949), .C1(
        P1_U3086), .C2(n7144), .ZN(P1_U3354) );
  OAI222_X1 U8207 ( .A1(P1_U3086), .A2(n7146), .B1(n10704), .B2(n8374), .C1(
        n6951), .C2(n10701), .ZN(P1_U3353) );
  OAI222_X1 U8208 ( .A1(P1_U3086), .A2(n7150), .B1(n10704), .B2(n6953), .C1(
        n6952), .C2(n10701), .ZN(P1_U3351) );
  INV_X1 U8209 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n6954) );
  OAI222_X1 U8210 ( .A1(n9109), .A2(n6956), .B1(n7272), .B2(P2_U3151), .C1(
        n6954), .C2(n9614), .ZN(P2_U3290) );
  OAI222_X1 U8211 ( .A1(P1_U3086), .A2(n7152), .B1(n10704), .B2(n6956), .C1(
        n6955), .C2(n10701), .ZN(P1_U3350) );
  INV_X1 U8212 ( .A(n10701), .ZN(n10695) );
  AOI22_X1 U8213 ( .A1(n7178), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_6__SCAN_IN), .B2(n10695), .ZN(n6957) );
  OAI21_X1 U8214 ( .B1(n6959), .B2(n10704), .A(n6957), .ZN(P1_U3349) );
  INV_X1 U8215 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n6958) );
  OAI222_X1 U8216 ( .A1(n9109), .A2(n6959), .B1(n7426), .B2(P2_U3151), .C1(
        n6958), .C2(n9614), .ZN(P2_U3289) );
  INV_X1 U8217 ( .A(P2_D_REG_24__SCAN_IN), .ZN(n6961) );
  NOR2_X1 U8218 ( .A1(n6991), .A2(n6961), .ZN(P2_U3241) );
  INV_X1 U8219 ( .A(P2_D_REG_25__SCAN_IN), .ZN(n6962) );
  NOR2_X1 U8220 ( .A1(n6991), .A2(n6962), .ZN(P2_U3240) );
  INV_X1 U8221 ( .A(P2_D_REG_30__SCAN_IN), .ZN(n6963) );
  NOR2_X1 U8222 ( .A1(n6991), .A2(n6963), .ZN(P2_U3235) );
  INV_X1 U8223 ( .A(P2_D_REG_23__SCAN_IN), .ZN(n6964) );
  NOR2_X1 U8224 ( .A1(n6991), .A2(n6964), .ZN(P2_U3242) );
  INV_X1 U8225 ( .A(P2_D_REG_29__SCAN_IN), .ZN(n6965) );
  NOR2_X1 U8226 ( .A1(n6991), .A2(n6965), .ZN(P2_U3236) );
  INV_X1 U8227 ( .A(P2_D_REG_28__SCAN_IN), .ZN(n6966) );
  NOR2_X1 U8228 ( .A1(n6991), .A2(n6966), .ZN(P2_U3237) );
  INV_X1 U8229 ( .A(P2_D_REG_27__SCAN_IN), .ZN(n6967) );
  NOR2_X1 U8230 ( .A1(n6991), .A2(n6967), .ZN(P2_U3238) );
  INV_X1 U8231 ( .A(P2_D_REG_31__SCAN_IN), .ZN(n6968) );
  NOR2_X1 U8232 ( .A1(n6991), .A2(n6968), .ZN(P2_U3234) );
  INV_X1 U8233 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n6969) );
  OAI222_X1 U8234 ( .A1(n9109), .A2(n6971), .B1(n5580), .B2(P2_U3151), .C1(
        n6969), .C2(n9614), .ZN(P2_U3288) );
  INV_X1 U8235 ( .A(n7192), .ZN(n7183) );
  INV_X1 U8236 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n6970) );
  OAI222_X1 U8237 ( .A1(P1_U3086), .A2(n7183), .B1(n10704), .B2(n6971), .C1(
        n6970), .C2(n10701), .ZN(P1_U3348) );
  INV_X1 U8238 ( .A(n9623), .ZN(n6973) );
  AOI22_X1 U8239 ( .A1(n7453), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(n10695), .ZN(n6972) );
  OAI21_X1 U8240 ( .B1(n6973), .B2(n10704), .A(n6972), .ZN(P1_U3347) );
  INV_X1 U8241 ( .A(P2_D_REG_6__SCAN_IN), .ZN(n6974) );
  NOR2_X1 U8242 ( .A1(n6991), .A2(n6974), .ZN(P2_U3259) );
  INV_X1 U8243 ( .A(P2_D_REG_26__SCAN_IN), .ZN(n6975) );
  NOR2_X1 U8244 ( .A1(n6991), .A2(n6975), .ZN(P2_U3239) );
  INV_X1 U8245 ( .A(P2_D_REG_7__SCAN_IN), .ZN(n6976) );
  NOR2_X1 U8246 ( .A1(n6991), .A2(n6976), .ZN(P2_U3258) );
  INV_X1 U8247 ( .A(P2_D_REG_2__SCAN_IN), .ZN(n6977) );
  NOR2_X1 U8248 ( .A1(n6991), .A2(n6977), .ZN(P2_U3263) );
  INV_X1 U8249 ( .A(P2_D_REG_4__SCAN_IN), .ZN(n6978) );
  NOR2_X1 U8250 ( .A1(n6991), .A2(n6978), .ZN(P2_U3261) );
  INV_X1 U8251 ( .A(P2_D_REG_3__SCAN_IN), .ZN(n6979) );
  NOR2_X1 U8252 ( .A1(n6991), .A2(n6979), .ZN(P2_U3262) );
  INV_X1 U8253 ( .A(P2_D_REG_5__SCAN_IN), .ZN(n6980) );
  NOR2_X1 U8254 ( .A1(n6991), .A2(n6980), .ZN(P2_U3260) );
  INV_X1 U8255 ( .A(n7333), .ZN(n7106) );
  NAND2_X1 U8256 ( .A1(n9061), .A2(n7106), .ZN(n6981) );
  NAND2_X1 U8257 ( .A1(n6981), .A2(P1_STATE_REG_SCAN_IN), .ZN(n7140) );
  INV_X1 U8258 ( .A(n7140), .ZN(n6983) );
  NAND2_X1 U8259 ( .A1(n7117), .A2(n9061), .ZN(n6982) );
  NAND2_X1 U8260 ( .A1(n6982), .A2(n6474), .ZN(n7141) );
  NOR2_X1 U8261 ( .A1(n10868), .A2(P1_U3973), .ZN(P1_U3085) );
  INV_X1 U8262 ( .A(n6984), .ZN(n6988) );
  AOI22_X1 U8263 ( .A1(n10364), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_9__SCAN_IN), .B2(n10695), .ZN(n6985) );
  OAI21_X1 U8264 ( .B1(n6988), .B2(n10704), .A(n6985), .ZN(P1_U3346) );
  INV_X1 U8265 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n6986) );
  OAI222_X1 U8266 ( .A1(n9109), .A2(n6990), .B1(n7989), .B2(P2_U3151), .C1(
        n6986), .C2(n9614), .ZN(P2_U3285) );
  INV_X1 U8267 ( .A(n7761), .ZN(n7798) );
  INV_X1 U8268 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n6987) );
  OAI222_X1 U8269 ( .A1(n9109), .A2(n6988), .B1(n7798), .B2(P2_U3151), .C1(
        n6987), .C2(n9614), .ZN(P2_U3286) );
  OAI222_X1 U8270 ( .A1(P1_U3086), .A2(n7456), .B1(n10704), .B2(n6990), .C1(
        n6989), .C2(n10701), .ZN(P1_U3345) );
  INV_X1 U8271 ( .A(P2_D_REG_21__SCAN_IN), .ZN(n6992) );
  NOR2_X1 U8272 ( .A1(n6991), .A2(n6992), .ZN(P2_U3244) );
  INV_X1 U8273 ( .A(P2_D_REG_17__SCAN_IN), .ZN(n6993) );
  NOR2_X1 U8274 ( .A1(n6991), .A2(n6993), .ZN(P2_U3248) );
  INV_X1 U8275 ( .A(P2_D_REG_22__SCAN_IN), .ZN(n6994) );
  NOR2_X1 U8276 ( .A1(n6991), .A2(n6994), .ZN(P2_U3243) );
  INV_X1 U8277 ( .A(P2_D_REG_20__SCAN_IN), .ZN(n6995) );
  NOR2_X1 U8278 ( .A1(n6991), .A2(n6995), .ZN(P2_U3245) );
  INV_X1 U8279 ( .A(P2_D_REG_11__SCAN_IN), .ZN(n6996) );
  NOR2_X1 U8280 ( .A1(n6991), .A2(n6996), .ZN(P2_U3254) );
  INV_X1 U8281 ( .A(P2_D_REG_10__SCAN_IN), .ZN(n6997) );
  NOR2_X1 U8282 ( .A1(n6991), .A2(n6997), .ZN(P2_U3255) );
  INV_X1 U8283 ( .A(P2_D_REG_9__SCAN_IN), .ZN(n6998) );
  NOR2_X1 U8284 ( .A1(n6991), .A2(n6998), .ZN(P2_U3256) );
  INV_X1 U8285 ( .A(P2_D_REG_8__SCAN_IN), .ZN(n6999) );
  NOR2_X1 U8286 ( .A1(n6991), .A2(n6999), .ZN(P2_U3257) );
  INV_X1 U8287 ( .A(P2_D_REG_19__SCAN_IN), .ZN(n7000) );
  NOR2_X1 U8288 ( .A1(n6991), .A2(n7000), .ZN(P2_U3246) );
  INV_X1 U8289 ( .A(P2_D_REG_16__SCAN_IN), .ZN(n7001) );
  NOR2_X1 U8290 ( .A1(n6991), .A2(n7001), .ZN(P2_U3249) );
  INV_X1 U8291 ( .A(P2_D_REG_15__SCAN_IN), .ZN(n7002) );
  NOR2_X1 U8292 ( .A1(n6991), .A2(n7002), .ZN(P2_U3250) );
  INV_X1 U8293 ( .A(P2_D_REG_14__SCAN_IN), .ZN(n7003) );
  NOR2_X1 U8294 ( .A1(n6991), .A2(n7003), .ZN(P2_U3251) );
  INV_X1 U8295 ( .A(P2_D_REG_13__SCAN_IN), .ZN(n7004) );
  NOR2_X1 U8296 ( .A1(n6991), .A2(n7004), .ZN(P2_U3252) );
  INV_X1 U8297 ( .A(P2_D_REG_18__SCAN_IN), .ZN(n7005) );
  NOR2_X1 U8298 ( .A1(n6991), .A2(n7005), .ZN(P2_U3247) );
  INV_X1 U8299 ( .A(P2_D_REG_12__SCAN_IN), .ZN(n7006) );
  NOR2_X1 U8300 ( .A1(n6991), .A2(n7006), .ZN(P2_U3253) );
  INV_X1 U8301 ( .A(n6587), .ZN(n7023) );
  AOI22_X1 U8302 ( .A1(n10806), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_11__SCAN_IN), .B2(n10695), .ZN(n7007) );
  OAI21_X1 U8303 ( .B1(n7023), .B2(n10704), .A(n7007), .ZN(P1_U3344) );
  NAND2_X1 U8304 ( .A1(n7008), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7014) );
  MUX2_X1 U8305 ( .A(n10977), .B(n7014), .S(n6347), .Z(n7010) );
  INV_X1 U8306 ( .A(n7011), .ZN(n8033) );
  NOR2_X1 U8307 ( .A1(n7012), .A2(n8033), .ZN(n7013) );
  INV_X1 U8308 ( .A(n10938), .ZN(n10965) );
  NOR2_X1 U8309 ( .A1(n7095), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7021) );
  OR2_X1 U8310 ( .A1(n7014), .A2(n6347), .ZN(n7047) );
  INV_X1 U8311 ( .A(n10962), .ZN(n10915) );
  INV_X1 U8312 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n7015) );
  MUX2_X1 U8313 ( .A(n7016), .B(n7015), .S(n6348), .Z(n7017) );
  NAND2_X1 U8314 ( .A1(n7017), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n10898) );
  MUX2_X1 U8315 ( .A(P2_REG2_REG_0__SCAN_IN), .B(P2_REG1_REG_0__SCAN_IN), .S(
        n9324), .Z(n7018) );
  NAND2_X1 U8316 ( .A1(n7018), .A2(n7048), .ZN(n7019) );
  AOI22_X1 U8317 ( .A1(n7047), .A2(n10915), .B1(n10898), .B2(n7019), .ZN(n7020) );
  AOI211_X1 U8318 ( .C1(P2_ADDR_REG_0__SCAN_IN), .C2(n10965), .A(n7021), .B(
        n7020), .ZN(n7022) );
  OAI21_X1 U8319 ( .B1(n7048), .B2(n10976), .A(n7022), .ZN(P2_U3182) );
  INV_X1 U8320 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n7024) );
  INV_X1 U8321 ( .A(n8078), .ZN(n8092) );
  OAI222_X1 U8322 ( .A1(n9614), .A2(n7024), .B1(n9619), .B2(n7023), .C1(
        P2_U3151), .C2(n8092), .ZN(P2_U3284) );
  INV_X1 U8323 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n7028) );
  INV_X1 U8324 ( .A(n7025), .ZN(n7730) );
  NAND2_X1 U8325 ( .A1(n10297), .A2(n7725), .ZN(n8987) );
  NAND2_X1 U8326 ( .A1(n7730), .A2(n8987), .ZN(n8929) );
  OAI21_X1 U8327 ( .B1(n11168), .B2(n10566), .A(n8929), .ZN(n7026) );
  NAND2_X1 U8328 ( .A1(n11000), .A2(n11002), .ZN(n7200) );
  OAI211_X1 U8329 ( .C1(n5278), .C2(n7725), .A(n7026), .B(n7200), .ZN(n10651)
         );
  NAND2_X1 U8330 ( .A1(n10651), .A2(n11175), .ZN(n7027) );
  OAI21_X1 U8331 ( .B1(n11175), .B2(n7028), .A(n7027), .ZN(P1_U3453) );
  INV_X1 U8332 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n7029) );
  OAI222_X1 U8333 ( .A1(n9109), .A2(n7031), .B1(n8153), .B2(P2_U3151), .C1(
        n7029), .C2(n9614), .ZN(P2_U3283) );
  OAI222_X1 U8334 ( .A1(P1_U3086), .A2(n7463), .B1(n10704), .B2(n7031), .C1(
        n7030), .C2(n10701), .ZN(P1_U3343) );
  OR2_X1 U8335 ( .A1(n8491), .A2(n7296), .ZN(n7093) );
  INV_X1 U8336 ( .A(n7093), .ZN(n8447) );
  NAND2_X1 U8337 ( .A1(n9217), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7077) );
  NAND2_X1 U8338 ( .A1(n7077), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n7033) );
  AOI22_X1 U8339 ( .A1(n9214), .A2(n9259), .B1(n9219), .B2(n7097), .ZN(n7032)
         );
  OAI211_X1 U8340 ( .C1(n8447), .C2(n9224), .A(n7033), .B(n7032), .ZN(P2_U3172) );
  MUX2_X1 U8341 ( .A(P2_REG2_REG_1__SCAN_IN), .B(P2_REG1_REG_1__SCAN_IN), .S(
        n6348), .Z(n7034) );
  INV_X1 U8342 ( .A(n7050), .ZN(n10896) );
  XNOR2_X1 U8343 ( .A(n7034), .B(n10896), .ZN(n10897) );
  AOI22_X1 U8344 ( .A1(n10897), .A2(n10898), .B1(n7034), .B2(n7050), .ZN(n8352) );
  MUX2_X1 U8345 ( .A(P2_REG2_REG_2__SCAN_IN), .B(P2_REG1_REG_2__SCAN_IN), .S(
        n6348), .Z(n7035) );
  XNOR2_X1 U8346 ( .A(n7035), .B(n8375), .ZN(n8353) );
  INV_X1 U8347 ( .A(n8375), .ZN(n7037) );
  INV_X1 U8348 ( .A(n7035), .ZN(n7036) );
  OAI22_X1 U8349 ( .A1(n8352), .A2(n8353), .B1(n7037), .B2(n7036), .ZN(n7039)
         );
  MUX2_X1 U8350 ( .A(P2_REG2_REG_3__SCAN_IN), .B(P2_REG1_REG_3__SCAN_IN), .S(
        n9324), .Z(n7260) );
  XNOR2_X1 U8351 ( .A(n7260), .B(n7259), .ZN(n7038) );
  NOR2_X1 U8352 ( .A1(n7038), .A2(n7039), .ZN(n7257) );
  AOI21_X1 U8353 ( .B1(n7039), .B2(n7038), .A(n7257), .ZN(n7063) );
  INV_X1 U8354 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n7040) );
  NOR2_X1 U8355 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7040), .ZN(n7222) );
  AND2_X1 U8356 ( .A1(P2_REG2_REG_0__SCAN_IN), .A2(n7048), .ZN(n7041) );
  OAI21_X1 U8357 ( .B1(n7050), .B2(n7041), .A(n7042), .ZN(n10890) );
  NOR2_X1 U8358 ( .A1(n10890), .A2(n10891), .ZN(n10889) );
  INV_X1 U8359 ( .A(n7042), .ZN(n7043) );
  OR2_X1 U8360 ( .A1(n10889), .A2(n7043), .ZN(n8357) );
  NAND2_X1 U8361 ( .A1(n8375), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n7044) );
  INV_X1 U8362 ( .A(n7259), .ZN(n7060) );
  NAND2_X1 U8363 ( .A1(P2_REG2_REG_3__SCAN_IN), .A2(n7045), .ZN(n7246) );
  OAI21_X1 U8364 ( .B1(n7045), .B2(P2_REG2_REG_3__SCAN_IN), .A(n7246), .ZN(
        n7046) );
  INV_X1 U8365 ( .A(n7046), .ZN(n7058) );
  AND2_X1 U8366 ( .A1(n7048), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n7049) );
  OAI21_X1 U8367 ( .B1(n7050), .B2(n7049), .A(n7051), .ZN(n10887) );
  NOR2_X1 U8368 ( .A1(n10887), .A2(n5939), .ZN(n10886) );
  INV_X1 U8369 ( .A(n7051), .ZN(n7052) );
  OR2_X1 U8370 ( .A1(n10886), .A2(n7052), .ZN(n8362) );
  MUX2_X1 U8371 ( .A(P2_REG1_REG_2__SCAN_IN), .B(n5955), .S(n7053), .Z(n8363)
         );
  NAND2_X1 U8372 ( .A1(n8375), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n7054) );
  NAND2_X1 U8373 ( .A1(n8364), .A2(n7054), .ZN(n7055) );
  AOI21_X1 U8374 ( .B1(n7056), .B2(n5905), .A(n5220), .ZN(n7057) );
  OAI22_X1 U8375 ( .A1(n7058), .A2(n10974), .B1(n10969), .B2(n7057), .ZN(n7059) );
  AOI211_X1 U8376 ( .C1(n10965), .C2(P2_ADDR_REG_3__SCAN_IN), .A(n7222), .B(
        n7059), .ZN(n7062) );
  NAND2_X1 U8377 ( .A1(n10941), .A2(n7060), .ZN(n7061) );
  OAI211_X1 U8378 ( .C1(n7063), .C2(n10915), .A(n7062), .B(n7061), .ZN(
        P2_U3185) );
  AOI21_X1 U8379 ( .B1(n7066), .B2(n7065), .A(n7064), .ZN(n7070) );
  AOI22_X1 U8380 ( .A1(n9229), .A2(n9260), .B1(n9219), .B2(n6899), .ZN(n7067)
         );
  OAI21_X1 U8381 ( .B1(n7289), .B2(n9231), .A(n7067), .ZN(n7068) );
  AOI21_X1 U8382 ( .B1(P2_REG3_REG_1__SCAN_IN), .B2(n7077), .A(n7068), .ZN(
        n7069) );
  OAI21_X1 U8383 ( .B1(n7070), .B2(n9224), .A(n7069), .ZN(P2_U3162) );
  AOI22_X1 U8384 ( .A1(n10864), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n10695), .ZN(n7071) );
  OAI21_X1 U8385 ( .B1(n7101), .B2(n10704), .A(n7071), .ZN(P1_U3342) );
  AOI21_X1 U8386 ( .B1(n7073), .B2(n7072), .A(n5219), .ZN(n7079) );
  AOI22_X1 U8387 ( .A1(n9229), .A2(n9259), .B1(n9219), .B2(n7074), .ZN(n7075)
         );
  OAI21_X1 U8388 ( .B1(n5389), .B2(n9231), .A(n7075), .ZN(n7076) );
  AOI21_X1 U8389 ( .B1(P2_REG3_REG_2__SCAN_IN), .B2(n7077), .A(n7076), .ZN(
        n7078) );
  OAI21_X1 U8390 ( .B1(n7079), .B2(n9224), .A(n7078), .ZN(P2_U3177) );
  NAND3_X1 U8391 ( .A1(n7081), .A2(n7083), .A3(n7080), .ZN(n7085) );
  OR2_X1 U8392 ( .A1(n7083), .A2(n7082), .ZN(n7084) );
  NAND2_X1 U8393 ( .A1(n7085), .A2(n7084), .ZN(n7088) );
  INV_X1 U8394 ( .A(n7086), .ZN(n7087) );
  INV_X1 U8395 ( .A(n7090), .ZN(n7092) );
  NAND4_X1 U8396 ( .A1(n7093), .A2(n7092), .A3(n7091), .A4(n9565), .ZN(n7094)
         );
  OAI21_X1 U8397 ( .B1(n11104), .B2(n7095), .A(n7094), .ZN(n7096) );
  AOI21_X1 U8398 ( .B1(n7097), .B2(n9509), .A(n7096), .ZN(n7099) );
  NOR2_X1 U8399 ( .A1(n7317), .A2(n9476), .ZN(n7102) );
  NAND2_X1 U8400 ( .A1(n7102), .A2(n9500), .ZN(n7098) );
  OAI211_X1 U8401 ( .C1(n7016), .C2(n9500), .A(n7099), .B(n7098), .ZN(P2_U3233) );
  INV_X1 U8402 ( .A(n8270), .ZN(n8263) );
  INV_X1 U8403 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n7100) );
  OAI222_X1 U8404 ( .A1(n9109), .A2(n7101), .B1(n8263), .B2(P2_U3151), .C1(
        n7100), .C2(n9614), .ZN(P2_U3282) );
  INV_X1 U8405 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n7104) );
  AOI21_X1 U8406 ( .B1(n9567), .B2(n9471), .A(n8447), .ZN(n7103) );
  NOR2_X1 U8407 ( .A1(n7103), .A2(n7102), .ZN(n7218) );
  MUX2_X1 U8408 ( .A(n7104), .B(n7218), .S(n11178), .Z(n7105) );
  OAI21_X1 U8409 ( .B1(n7215), .B2(n9607), .A(n7105), .ZN(P2_U3390) );
  AOI21_X1 U8410 ( .B1(n7107), .B2(n9062), .A(n7106), .ZN(n7109) );
  NAND2_X1 U8411 ( .A1(n7108), .A2(n6814), .ZN(n7551) );
  NAND2_X2 U8412 ( .A1(n7109), .A2(n7551), .ZN(n8806) );
  AND2_X1 U8413 ( .A1(n7333), .A2(n6813), .ZN(n7112) );
  NAND2_X1 U8414 ( .A1(n10297), .A2(n5136), .ZN(n7113) );
  INV_X1 U8415 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n10789) );
  NAND2_X1 U8416 ( .A1(n10297), .A2(n8692), .ZN(n7116) );
  OAI22_X1 U8417 ( .A1(n7725), .A2(n5152), .B1(n7333), .B2(n10793), .ZN(n7114)
         );
  INV_X1 U8418 ( .A(n7114), .ZN(n7115) );
  NAND2_X1 U8419 ( .A1(n7116), .A2(n7115), .ZN(n7228) );
  XNOR2_X1 U8420 ( .A(n7229), .B(n7228), .ZN(n10309) );
  OR2_X1 U8421 ( .A1(n10985), .A2(n7117), .ZN(n7129) );
  INV_X1 U8422 ( .A(n7129), .ZN(n7121) );
  INV_X1 U8423 ( .A(n7118), .ZN(n7207) );
  NAND3_X1 U8424 ( .A1(n7120), .A2(n7207), .A3(n7119), .ZN(n7132) );
  INV_X1 U8425 ( .A(n7132), .ZN(n7124) );
  NAND2_X1 U8426 ( .A1(n7202), .A2(n10689), .ZN(n9065) );
  NOR2_X1 U8427 ( .A1(n7132), .A2(n9065), .ZN(n7239) );
  INV_X1 U8428 ( .A(n10259), .ZN(n10233) );
  INV_X1 U8429 ( .A(n10689), .ZN(n7126) );
  NAND2_X1 U8430 ( .A1(n7201), .A2(n7122), .ZN(n7533) );
  NOR2_X1 U8431 ( .A1(n7126), .A2(n7533), .ZN(n7123) );
  NAND2_X1 U8432 ( .A1(n7124), .A2(n7123), .ZN(n7127) );
  AOI22_X1 U8433 ( .A1(n10233), .A2(n11000), .B1(n7128), .B2(n10266), .ZN(
        n7135) );
  NAND3_X1 U8434 ( .A1(n7129), .A2(n9065), .A3(n7533), .ZN(n7133) );
  INV_X1 U8435 ( .A(n7130), .ZN(n7131) );
  AOI21_X1 U8436 ( .B1(n7133), .B2(n7132), .A(n7131), .ZN(n7334) );
  NAND2_X1 U8437 ( .A1(n7334), .A2(n10689), .ZN(n10223) );
  NAND2_X1 U8438 ( .A1(n10223), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n7134) );
  OAI211_X1 U8439 ( .C1(n10309), .C2(n10269), .A(n7135), .B(n7134), .ZN(
        P1_U3232) );
  INV_X1 U8440 ( .A(n7152), .ZN(n7168) );
  INV_X1 U8441 ( .A(n7150), .ZN(n10350) );
  INV_X1 U8442 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n10991) );
  AND2_X1 U8443 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(
        n10303) );
  NAND2_X1 U8444 ( .A1(n10304), .A2(n10303), .ZN(n10302) );
  INV_X1 U8445 ( .A(n7144), .ZN(n10301) );
  NAND2_X1 U8446 ( .A1(n10301), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n7136) );
  NAND2_X1 U8447 ( .A1(n10302), .A2(n7136), .ZN(n10320) );
  XNOR2_X1 U8448 ( .A(n7146), .B(P1_REG1_REG_2__SCAN_IN), .ZN(n10321) );
  NAND2_X1 U8449 ( .A1(n10320), .A2(n10321), .ZN(n10319) );
  INV_X1 U8450 ( .A(n7146), .ZN(n10324) );
  NAND2_X1 U8451 ( .A1(n10324), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n7137) );
  NAND2_X1 U8452 ( .A1(n10319), .A2(n7137), .ZN(n10336) );
  XNOR2_X1 U8453 ( .A(n7148), .B(P1_REG1_REG_3__SCAN_IN), .ZN(n10337) );
  NAND2_X1 U8454 ( .A1(n10336), .A2(n10337), .ZN(n10335) );
  INV_X1 U8455 ( .A(n7148), .ZN(n10331) );
  NAND2_X1 U8456 ( .A1(n10331), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n7138) );
  NAND2_X1 U8457 ( .A1(n10335), .A2(n7138), .ZN(n10346) );
  XNOR2_X1 U8458 ( .A(n7150), .B(P1_REG1_REG_4__SCAN_IN), .ZN(n10347) );
  NAND2_X1 U8459 ( .A1(n10346), .A2(n10347), .ZN(n10345) );
  INV_X1 U8460 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n7139) );
  MUX2_X1 U8461 ( .A(P1_REG1_REG_5__SCAN_IN), .B(n7139), .S(n7152), .Z(n7162)
         );
  XNOR2_X1 U8462 ( .A(n7178), .B(P1_REG1_REG_6__SCAN_IN), .ZN(n7142) );
  NOR2_X1 U8463 ( .A1(n7143), .A2(n7142), .ZN(n7174) );
  OR2_X1 U8464 ( .A1(n7141), .A2(n7140), .ZN(n10796) );
  AOI211_X1 U8465 ( .C1(n7143), .C2(n7142), .A(n7174), .B(n10874), .ZN(n7160)
         );
  INV_X1 U8466 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n7151) );
  MUX2_X1 U8467 ( .A(n6453), .B(P1_REG2_REG_1__SCAN_IN), .S(n7144), .Z(n10300)
         );
  NAND2_X1 U8468 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n10311) );
  INV_X1 U8469 ( .A(n10311), .ZN(n10299) );
  NAND2_X1 U8470 ( .A1(n10300), .A2(n10299), .ZN(n10298) );
  NAND2_X1 U8471 ( .A1(n10301), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n7145) );
  NAND2_X1 U8472 ( .A1(n10298), .A2(n7145), .ZN(n10317) );
  XNOR2_X1 U8473 ( .A(n7146), .B(P1_REG2_REG_2__SCAN_IN), .ZN(n10318) );
  NAND2_X1 U8474 ( .A1(n10317), .A2(n10318), .ZN(n10316) );
  NAND2_X1 U8475 ( .A1(n10324), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n7147) );
  NAND2_X1 U8476 ( .A1(n10316), .A2(n7147), .ZN(n10333) );
  XNOR2_X1 U8477 ( .A(n7148), .B(P1_REG2_REG_3__SCAN_IN), .ZN(n10334) );
  NAND2_X1 U8478 ( .A1(n10333), .A2(n10334), .ZN(n10332) );
  NAND2_X1 U8479 ( .A1(n10331), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n7149) );
  NAND2_X1 U8480 ( .A1(n10332), .A2(n7149), .ZN(n10343) );
  XNOR2_X1 U8481 ( .A(n7150), .B(P1_REG2_REG_4__SCAN_IN), .ZN(n10344) );
  NAND2_X1 U8482 ( .A1(n10343), .A2(n10344), .ZN(n10342) );
  OAI21_X1 U8483 ( .B1(n7151), .B2(n7150), .A(n10342), .ZN(n7165) );
  INV_X1 U8484 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n7153) );
  MUX2_X1 U8485 ( .A(n7153), .B(P1_REG2_REG_5__SCAN_IN), .S(n7152), .Z(n7164)
         );
  AND2_X1 U8486 ( .A1(n7165), .A2(n7164), .ZN(n7167) );
  AOI21_X1 U8487 ( .B1(n7168), .B2(P1_REG2_REG_5__SCAN_IN), .A(n7167), .ZN(
        n7155) );
  XNOR2_X1 U8488 ( .A(n7178), .B(P1_REG2_REG_6__SCAN_IN), .ZN(n7154) );
  NOR2_X1 U8489 ( .A1(n7155), .A2(n7154), .ZN(n7177) );
  NAND2_X1 U8490 ( .A1(n10790), .A2(n8291), .ZN(n10310) );
  AOI211_X1 U8491 ( .C1(n7155), .C2(n7154), .A(n7177), .B(n10870), .ZN(n7159)
         );
  INV_X1 U8492 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n7157) );
  NOR2_X2 U8493 ( .A1(n10796), .A2(n10790), .ZN(n10881) );
  NAND2_X1 U8494 ( .A1(n10881), .A2(n7178), .ZN(n7156) );
  NAND2_X1 U8495 ( .A1(P1_U3086), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n7504) );
  OAI211_X1 U8496 ( .C1(n10885), .C2(n7157), .A(n7156), .B(n7504), .ZN(n7158)
         );
  OR3_X1 U8497 ( .A1(n7160), .A2(n7159), .A3(n7158), .ZN(P1_U3249) );
  AOI211_X1 U8498 ( .C1(n7163), .C2(n7162), .A(n7161), .B(n10874), .ZN(n7173)
         );
  NOR2_X1 U8499 ( .A1(n7165), .A2(n7164), .ZN(n7166) );
  NOR3_X1 U8500 ( .A1(n10870), .A2(n7167), .A3(n7166), .ZN(n7172) );
  INV_X1 U8501 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n7170) );
  NAND2_X1 U8502 ( .A1(n10881), .A2(n7168), .ZN(n7169) );
  NAND2_X1 U8503 ( .A1(P1_U3086), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n7543) );
  OAI211_X1 U8504 ( .C1(n10885), .C2(n7170), .A(n7169), .B(n7543), .ZN(n7171)
         );
  OR3_X1 U8505 ( .A1(n7173), .A2(n7172), .A3(n7171), .ZN(P1_U3248) );
  AOI21_X1 U8506 ( .B1(n7178), .B2(P1_REG1_REG_6__SCAN_IN), .A(n7174), .ZN(
        n7176) );
  XNOR2_X1 U8507 ( .A(n7192), .B(P1_REG1_REG_7__SCAN_IN), .ZN(n7175) );
  NOR2_X1 U8508 ( .A1(n7176), .A2(n7175), .ZN(n7187) );
  AOI211_X1 U8509 ( .C1(n7176), .C2(n7175), .A(n10874), .B(n7187), .ZN(n7186)
         );
  AOI21_X1 U8510 ( .B1(n7178), .B2(P1_REG2_REG_6__SCAN_IN), .A(n7177), .ZN(
        n7180) );
  XNOR2_X1 U8511 ( .A(n7192), .B(P1_REG2_REG_7__SCAN_IN), .ZN(n7179) );
  NOR2_X1 U8512 ( .A1(n7180), .A2(n7179), .ZN(n7191) );
  AOI211_X1 U8513 ( .C1(n7180), .C2(n7179), .A(n10870), .B(n7191), .ZN(n7185)
         );
  INV_X1 U8514 ( .A(n10881), .ZN(n10414) );
  INV_X1 U8515 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n7181) );
  NOR2_X1 U8516 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7181), .ZN(n7634) );
  AOI21_X1 U8517 ( .B1(n10868), .B2(P1_ADDR_REG_7__SCAN_IN), .A(n7634), .ZN(
        n7182) );
  OAI21_X1 U8518 ( .B1(n10414), .B2(n7183), .A(n7182), .ZN(n7184) );
  OR3_X1 U8519 ( .A1(n7186), .A2(n7185), .A3(n7184), .ZN(P1_U3250) );
  INV_X1 U8520 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n7188) );
  MUX2_X1 U8521 ( .A(n7188), .B(P1_REG1_REG_8__SCAN_IN), .S(n7453), .Z(n7189)
         );
  AOI211_X1 U8522 ( .C1(n7190), .C2(n7189), .A(n10874), .B(n7445), .ZN(n7199)
         );
  AOI21_X1 U8523 ( .B1(n7192), .B2(P1_REG2_REG_7__SCAN_IN), .A(n7191), .ZN(
        n7194) );
  XNOR2_X1 U8524 ( .A(n7453), .B(P1_REG2_REG_8__SCAN_IN), .ZN(n7193) );
  NOR2_X1 U8525 ( .A1(n7194), .A2(n7193), .ZN(n7452) );
  AOI211_X1 U8526 ( .C1(n7194), .C2(n7193), .A(n10870), .B(n7452), .ZN(n7198)
         );
  INV_X1 U8527 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n7196) );
  NAND2_X1 U8528 ( .A1(n10881), .A2(n7453), .ZN(n7195) );
  NAND2_X1 U8529 ( .A1(P1_U3086), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n10094) );
  OAI211_X1 U8530 ( .C1(n10885), .C2(n7196), .A(n7195), .B(n10094), .ZN(n7197)
         );
  OR3_X1 U8531 ( .A1(n7199), .A2(n7198), .A3(n7197), .ZN(P1_U3251) );
  INV_X1 U8532 ( .A(n7200), .ZN(n7205) );
  INV_X1 U8533 ( .A(n8929), .ZN(n7203) );
  NOR3_X1 U8534 ( .A1(n7203), .A2(n7202), .A3(n7201), .ZN(n7204) );
  AOI211_X1 U8535 ( .C1(n11149), .C2(P1_REG3_REG_0__SCAN_IN), .A(n7205), .B(
        n7204), .ZN(n7213) );
  AND2_X1 U8536 ( .A1(n7207), .A2(n7206), .ZN(n7208) );
  NAND2_X1 U8537 ( .A1(n7209), .A2(n7208), .ZN(n7210) );
  NOR4_X1 U8538 ( .A1(n7210), .A2(n7108), .A3(n5278), .A4(n7725), .ZN(n7211)
         );
  AOI21_X1 U8539 ( .B1(n11011), .B2(P1_REG2_REG_0__SCAN_IN), .A(n7211), .ZN(
        n7212) );
  OAI21_X1 U8540 ( .B1(n7213), .B2(n11011), .A(n7212), .ZN(P1_U3293) );
  INV_X1 U8541 ( .A(P1_U3973), .ZN(n10296) );
  NAND2_X1 U8542 ( .A1(n10296), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n7214) );
  OAI21_X1 U8543 ( .B1(n8816), .B2(n10296), .A(n7214), .ZN(P1_U3583) );
  OAI22_X1 U8544 ( .A1(n7215), .A2(n9564), .B1(n9561), .B2(n7015), .ZN(n7216)
         );
  INV_X1 U8545 ( .A(n7216), .ZN(n7217) );
  OAI21_X1 U8546 ( .B1(n7218), .B2(n9572), .A(n7217), .ZN(P2_U3459) );
  INV_X1 U8547 ( .A(n9224), .ZN(n9158) );
  OAI211_X1 U8548 ( .C1(n7221), .C2(n7220), .A(n7219), .B(n9158), .ZN(n7227)
         );
  INV_X1 U8549 ( .A(n7478), .ZN(n9257) );
  AOI21_X1 U8550 ( .B1(n9219), .B2(n7223), .A(n7222), .ZN(n7224) );
  OAI21_X1 U8551 ( .B1(n9125), .B2(n7289), .A(n7224), .ZN(n7225) );
  AOI21_X1 U8552 ( .B1(n9214), .B2(n9257), .A(n7225), .ZN(n7226) );
  OAI211_X1 U8553 ( .C1(P2_REG3_REG_3__SCAN_IN), .C2(n9217), .A(n7227), .B(
        n7226), .ZN(P2_U3158) );
  INV_X1 U8554 ( .A(n7236), .ZN(n7234) );
  NAND2_X1 U8555 ( .A1(n7344), .A2(n7729), .ZN(n7231) );
  NAND2_X1 U8556 ( .A1(n11000), .A2(n5136), .ZN(n7230) );
  NAND2_X1 U8557 ( .A1(n7231), .A2(n7230), .ZN(n7232) );
  XNOR2_X1 U8558 ( .A(n7232), .B(n8809), .ZN(n7235) );
  INV_X1 U8559 ( .A(n7235), .ZN(n7233) );
  NAND2_X1 U8560 ( .A1(n7234), .A2(n7233), .ZN(n7342) );
  NAND2_X1 U8561 ( .A1(n7236), .A2(n7235), .ZN(n7341) );
  NAND2_X1 U8562 ( .A1(n7342), .A2(n7341), .ZN(n7238) );
  AND2_X1 U8563 ( .A1(n7729), .A2(n5136), .ZN(n7237) );
  AOI21_X1 U8564 ( .B1(n11000), .B2(n8692), .A(n7237), .ZN(n7340) );
  XNOR2_X1 U8565 ( .A(n7238), .B(n7340), .ZN(n7242) );
  AOI22_X1 U8566 ( .A1(n10233), .A2(n10295), .B1(n7729), .B2(n10266), .ZN(
        n7241) );
  AOI22_X1 U8567 ( .A1(n10223), .A2(P1_REG3_REG_1__SCAN_IN), .B1(n10261), .B2(
        n10297), .ZN(n7240) );
  OAI211_X1 U8568 ( .C1(n7242), .C2(n10269), .A(n7241), .B(n7240), .ZN(
        P1_U3222) );
  INV_X1 U8569 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n7243) );
  OAI222_X1 U8570 ( .A1(n9109), .A2(n8377), .B1(n9269), .B2(P2_U3151), .C1(
        n7243), .C2(n9614), .ZN(P2_U3281) );
  INV_X1 U8571 ( .A(n9298), .ZN(n9286) );
  INV_X1 U8572 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n7244) );
  OAI222_X1 U8573 ( .A1(n9109), .A2(n7282), .B1(n9286), .B2(P2_U3151), .C1(
        n7244), .C2(n9614), .ZN(P2_U3280) );
  INV_X1 U8574 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n7256) );
  AOI22_X1 U8575 ( .A1(n7429), .A2(n7515), .B1(P2_REG2_REG_6__SCAN_IN), .B2(
        n7426), .ZN(n7252) );
  NAND2_X1 U8576 ( .A1(P2_REG2_REG_4__SCAN_IN), .A2(n7268), .ZN(n7248) );
  INV_X1 U8577 ( .A(n7268), .ZN(n10913) );
  AOI22_X1 U8578 ( .A1(n10913), .A2(n7585), .B1(P2_REG2_REG_4__SCAN_IN), .B2(
        n7268), .ZN(n10905) );
  NAND2_X1 U8579 ( .A1(n7245), .A2(n7259), .ZN(n7247) );
  NAND2_X1 U8580 ( .A1(n7247), .A2(n7246), .ZN(n10904) );
  NAND2_X1 U8581 ( .A1(n10905), .A2(n10904), .ZN(n10903) );
  NAND2_X1 U8582 ( .A1(n7248), .A2(n10903), .ZN(n7249) );
  NAND2_X1 U8583 ( .A1(n7249), .A2(n7272), .ZN(n7250) );
  XNOR2_X1 U8584 ( .A(n7249), .B(n10932), .ZN(n10925) );
  NAND2_X1 U8585 ( .A1(P2_REG2_REG_5__SCAN_IN), .A2(n10925), .ZN(n10924) );
  OAI21_X1 U8586 ( .B1(n7252), .B2(n7251), .A(n7428), .ZN(n7253) );
  NAND2_X1 U8587 ( .A1(n10928), .A2(n7253), .ZN(n7255) );
  OAI211_X1 U8588 ( .C1(n7256), .C2(n10938), .A(n7255), .B(n7254), .ZN(n7279)
         );
  MUX2_X1 U8589 ( .A(P2_REG2_REG_4__SCAN_IN), .B(P2_REG1_REG_4__SCAN_IN), .S(
        n9324), .Z(n7261) );
  XNOR2_X1 U8590 ( .A(n7261), .B(n7268), .ZN(n10917) );
  INV_X1 U8591 ( .A(n7257), .ZN(n7258) );
  OAI21_X1 U8592 ( .B1(n7260), .B2(n7259), .A(n7258), .ZN(n10916) );
  NOR2_X1 U8593 ( .A1(n10917), .A2(n10916), .ZN(n10914) );
  AOI21_X1 U8594 ( .B1(n7261), .B2(n7268), .A(n10914), .ZN(n10933) );
  MUX2_X1 U8595 ( .A(n7576), .B(n7262), .S(n9324), .Z(n7263) );
  XNOR2_X1 U8596 ( .A(n7263), .B(n10932), .ZN(n10934) );
  OAI22_X1 U8597 ( .A1(n10933), .A2(n10934), .B1(n10932), .B2(n7263), .ZN(
        n7267) );
  MUX2_X1 U8598 ( .A(P2_REG2_REG_6__SCAN_IN), .B(P2_REG1_REG_6__SCAN_IN), .S(
        n9324), .Z(n7264) );
  NOR2_X1 U8599 ( .A1(n7264), .A2(n7426), .ZN(n7435) );
  AOI21_X1 U8600 ( .B1(n7264), .B2(n7426), .A(n7435), .ZN(n7265) );
  INV_X1 U8601 ( .A(n7265), .ZN(n7266) );
  NOR2_X1 U8602 ( .A1(n7267), .A2(n7266), .ZN(n7434) );
  AOI21_X1 U8603 ( .B1(n7267), .B2(n7266), .A(n7434), .ZN(n7277) );
  NAND2_X1 U8604 ( .A1(P2_REG1_REG_4__SCAN_IN), .A2(n7268), .ZN(n7269) );
  OAI21_X1 U8605 ( .B1(P2_REG1_REG_4__SCAN_IN), .B2(n7268), .A(n7269), .ZN(
        n10908) );
  NOR2_X1 U8606 ( .A1(n10909), .A2(n10908), .ZN(n10907) );
  INV_X1 U8607 ( .A(n7269), .ZN(n7270) );
  INV_X1 U8608 ( .A(n7271), .ZN(n7273) );
  INV_X1 U8609 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n7675) );
  AOI22_X1 U8610 ( .A1(n7429), .A2(P2_REG1_REG_6__SCAN_IN), .B1(n7675), .B2(
        n7426), .ZN(n7274) );
  NOR2_X1 U8611 ( .A1(n7275), .A2(n7274), .ZN(n7425) );
  AOI21_X1 U8612 ( .B1(n7275), .B2(n7274), .A(n7425), .ZN(n7276) );
  OAI22_X1 U8613 ( .A1(n7277), .A2(n10915), .B1(n7276), .B2(n10969), .ZN(n7278) );
  AOI211_X1 U8614 ( .C1(n7429), .C2(n10941), .A(n7279), .B(n7278), .ZN(n7280)
         );
  INV_X1 U8615 ( .A(n7280), .ZN(P2_U3188) );
  OAI222_X1 U8616 ( .A1(P1_U3086), .A2(n10385), .B1(n10704), .B2(n7282), .C1(
        n7281), .C2(n10701), .ZN(P1_U3340) );
  OAI21_X1 U8617 ( .B1(n7284), .B2(n7287), .A(n7283), .ZN(n7472) );
  NAND2_X1 U8618 ( .A1(n7286), .A2(n7285), .ZN(n7398) );
  XNOR2_X1 U8619 ( .A(n7287), .B(n7398), .ZN(n7288) );
  OAI222_X1 U8620 ( .A1(n9476), .A2(n7478), .B1(n9474), .B2(n7289), .C1(n9471), 
        .C2(n7288), .ZN(n7469) );
  AOI21_X1 U8621 ( .B1(n9541), .B2(n7472), .A(n7469), .ZN(n7295) );
  INV_X1 U8622 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n7290) );
  OAI22_X1 U8623 ( .A1(n9607), .A2(n7468), .B1(n11178), .B2(n7290), .ZN(n7291)
         );
  INV_X1 U8624 ( .A(n7291), .ZN(n7292) );
  OAI21_X1 U8625 ( .B1(n7295), .B2(n6432), .A(n7292), .ZN(P2_U3399) );
  OAI22_X1 U8626 ( .A1(n7468), .A2(n9564), .B1(n9561), .B2(n5905), .ZN(n7293)
         );
  INV_X1 U8627 ( .A(n7293), .ZN(n7294) );
  OAI21_X1 U8628 ( .B1(n7295), .B2(n9572), .A(n7294), .ZN(P2_U3462) );
  INV_X1 U8629 ( .A(n8057), .ZN(n7305) );
  INV_X1 U8630 ( .A(n7296), .ZN(n8490) );
  INV_X1 U8631 ( .A(n7297), .ZN(n7298) );
  AOI21_X1 U8632 ( .B1(n8490), .B2(n5436), .A(n7298), .ZN(n7304) );
  INV_X1 U8633 ( .A(n7304), .ZN(n7380) );
  AOI22_X1 U8634 ( .A1(n9492), .A2(n9260), .B1(n9258), .B2(n9495), .ZN(n7303)
         );
  XNOR2_X1 U8635 ( .A(n7300), .B(n7299), .ZN(n7301) );
  NAND2_X1 U8636 ( .A1(n7301), .A2(n9490), .ZN(n7302) );
  OAI211_X1 U8637 ( .C1(n7304), .C2(n7968), .A(n7303), .B(n7302), .ZN(n7379)
         );
  AOI21_X1 U8638 ( .B1(n7305), .B2(n7380), .A(n7379), .ZN(n7312) );
  INV_X1 U8639 ( .A(n6899), .ZN(n7309) );
  INV_X1 U8640 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n7306) );
  OAI22_X1 U8641 ( .A1(n9607), .A2(n7309), .B1(n11178), .B2(n7306), .ZN(n7307)
         );
  INV_X1 U8642 ( .A(n7307), .ZN(n7308) );
  OAI21_X1 U8643 ( .B1(n7312), .B2(n6432), .A(n7308), .ZN(P2_U3393) );
  OAI22_X1 U8644 ( .A1(n7309), .A2(n9564), .B1(n9561), .B2(n5939), .ZN(n7310)
         );
  INV_X1 U8645 ( .A(n7310), .ZN(n7311) );
  OAI21_X1 U8646 ( .B1(n7312), .B2(n9572), .A(n7311), .ZN(P2_U3460) );
  OAI21_X1 U8647 ( .B1(n7313), .B2(n8446), .A(n7314), .ZN(n11027) );
  NOR2_X1 U8648 ( .A1(n11024), .A2(n9565), .ZN(n7318) );
  XNOR2_X1 U8649 ( .A(n7315), .B(n8446), .ZN(n7316) );
  OAI222_X1 U8650 ( .A1(n9476), .A2(n5389), .B1(n9474), .B2(n7317), .C1(n9471), 
        .C2(n7316), .ZN(n11025) );
  AOI211_X1 U8651 ( .C1(n9541), .C2(n11027), .A(n7318), .B(n11025), .ZN(n11023) );
  OR2_X1 U8652 ( .A1(n11023), .A2(n9572), .ZN(n7319) );
  OAI21_X1 U8653 ( .B1(n9561), .B2(n5955), .A(n7319), .ZN(P2_U3461) );
  AOI21_X1 U8654 ( .B1(n7321), .B2(n7320), .A(n7387), .ZN(n7328) );
  INV_X1 U8655 ( .A(n7322), .ZN(n7586) );
  INV_X1 U8656 ( .A(n9217), .ZN(n9234) );
  INV_X1 U8657 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n7323) );
  NOR2_X1 U8658 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7323), .ZN(n10912) );
  NOR2_X1 U8659 ( .A1(n9125), .A2(n5389), .ZN(n7324) );
  AOI211_X1 U8660 ( .C1(n9219), .C2(n7587), .A(n10912), .B(n7324), .ZN(n7325)
         );
  OAI21_X1 U8661 ( .B1(n7513), .B2(n9231), .A(n7325), .ZN(n7326) );
  AOI21_X1 U8662 ( .B1(n7586), .B2(n9234), .A(n7326), .ZN(n7327) );
  OAI21_X1 U8663 ( .B1(n7328), .B2(n9224), .A(n7327), .ZN(P2_U3170) );
  INV_X1 U8664 ( .A(n7329), .ZN(n7331) );
  OAI222_X1 U8665 ( .A1(n10380), .A2(P1_U3086), .B1(n10704), .B2(n7331), .C1(
        n7330), .C2(n10701), .ZN(P1_U3339) );
  INV_X1 U8666 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n7332) );
  OAI222_X1 U8667 ( .A1(n9614), .A2(n7332), .B1(n9619), .B2(n7331), .C1(
        P2_U3151), .C2(n9336), .ZN(P2_U3279) );
  NAND3_X1 U8668 ( .A1(n7334), .A2(n9061), .A3(n7333), .ZN(n7335) );
  INV_X1 U8669 ( .A(n7344), .ZN(n7484) );
  NAND2_X1 U8670 ( .A1(n7344), .A2(n7654), .ZN(n7337) );
  NAND2_X1 U8671 ( .A1(n11001), .A2(n5136), .ZN(n7336) );
  NAND2_X1 U8672 ( .A1(n7337), .A2(n7336), .ZN(n7338) );
  XNOR2_X1 U8673 ( .A(n7338), .B(n8809), .ZN(n7362) );
  AND2_X1 U8674 ( .A1(n7654), .A2(n5136), .ZN(n7339) );
  AOI21_X1 U8675 ( .B1(n11001), .B2(n8692), .A(n7339), .ZN(n7363) );
  XNOR2_X1 U8676 ( .A(n7362), .B(n7363), .ZN(n7356) );
  NAND2_X1 U8677 ( .A1(n7341), .A2(n7340), .ZN(n7343) );
  NAND2_X1 U8678 ( .A1(n7343), .A2(n7342), .ZN(n10220) );
  NAND2_X1 U8679 ( .A1(n7344), .A2(n6484), .ZN(n7346) );
  NAND2_X1 U8680 ( .A1(n10295), .A2(n5136), .ZN(n7345) );
  NAND2_X1 U8681 ( .A1(n7346), .A2(n7345), .ZN(n7347) );
  XNOR2_X1 U8682 ( .A(n7347), .B(n8781), .ZN(n7352) );
  INV_X1 U8683 ( .A(n7352), .ZN(n7350) );
  AND2_X1 U8684 ( .A1(n6484), .A2(n5136), .ZN(n7348) );
  AOI21_X1 U8685 ( .B1(n10295), .B2(n8692), .A(n7348), .ZN(n7351) );
  INV_X1 U8686 ( .A(n7351), .ZN(n7349) );
  NAND2_X1 U8687 ( .A1(n7352), .A2(n7351), .ZN(n7354) );
  AND2_X1 U8688 ( .A1(n7353), .A2(n7354), .ZN(n10221) );
  NAND2_X1 U8689 ( .A1(n10220), .A2(n10221), .ZN(n10219) );
  NAND2_X1 U8690 ( .A1(n10219), .A2(n7354), .ZN(n7355) );
  NAND2_X1 U8691 ( .A1(n7355), .A2(n7356), .ZN(n7371) );
  OAI21_X1 U8692 ( .B1(n7356), .B2(n7355), .A(n7371), .ZN(n7357) );
  NAND2_X1 U8693 ( .A1(n7357), .A2(n10244), .ZN(n7361) );
  NAND2_X1 U8694 ( .A1(P1_U3086), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n10328) );
  INV_X1 U8695 ( .A(n10328), .ZN(n7359) );
  OAI22_X1 U8696 ( .A1(n10236), .A2(n6483), .B1(n7646), .B2(n10259), .ZN(n7358) );
  AOI211_X1 U8697 ( .C1(n7654), .C2(n10266), .A(n7359), .B(n7358), .ZN(n7360)
         );
  OAI211_X1 U8698 ( .C1(P1_REG3_REG_3__SCAN_IN), .C2(n10263), .A(n7361), .B(
        n7360), .ZN(P1_U3218) );
  INV_X1 U8699 ( .A(n7820), .ZN(n7378) );
  INV_X1 U8700 ( .A(n7362), .ZN(n7364) );
  NAND2_X1 U8701 ( .A1(n7364), .A2(n7363), .ZN(n7369) );
  AND2_X1 U8702 ( .A1(n7371), .A2(n7369), .ZN(n7373) );
  NAND2_X1 U8703 ( .A1(n7344), .A2(n7821), .ZN(n7366) );
  NAND2_X1 U8704 ( .A1(n10294), .A2(n5136), .ZN(n7365) );
  NAND2_X1 U8705 ( .A1(n7366), .A2(n7365), .ZN(n7367) );
  XNOR2_X1 U8706 ( .A(n7367), .B(n8809), .ZN(n7483) );
  AND2_X1 U8707 ( .A1(n7821), .A2(n5136), .ZN(n7368) );
  AOI21_X1 U8708 ( .B1(n10294), .B2(n8692), .A(n7368), .ZN(n7481) );
  XNOR2_X1 U8709 ( .A(n7483), .B(n7481), .ZN(n7372) );
  AND2_X1 U8710 ( .A1(n7372), .A2(n7369), .ZN(n7370) );
  OAI211_X1 U8711 ( .C1(n7373), .C2(n7372), .A(n10244), .B(n7493), .ZN(n7377)
         );
  AND2_X1 U8712 ( .A1(P1_U3086), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n10341) );
  INV_X1 U8713 ( .A(n11001), .ZN(n7374) );
  OAI22_X1 U8714 ( .A1(n10236), .A2(n7374), .B1(n7833), .B2(n10259), .ZN(n7375) );
  AOI211_X1 U8715 ( .C1(n7821), .C2(n10266), .A(n10341), .B(n7375), .ZN(n7376)
         );
  OAI211_X1 U8716 ( .C1(n10263), .C2(n7378), .A(n7377), .B(n7376), .ZN(
        P1_U3230) );
  OR2_X1 U8717 ( .A1(n6896), .A2(n6895), .ZN(n7467) );
  INV_X1 U8718 ( .A(n7467), .ZN(n7970) );
  AOI21_X1 U8719 ( .B1(n7970), .B2(n7380), .A(n7379), .ZN(n7381) );
  INV_X2 U8720 ( .A(n9500), .ZN(n9488) );
  MUX2_X1 U8721 ( .A(n10891), .B(n7381), .S(n11111), .Z(n7383) );
  NAND2_X1 U8722 ( .A1(n9509), .A2(n6899), .ZN(n7382) );
  OAI211_X1 U8723 ( .C1(n11104), .C2(n10902), .A(n7383), .B(n7382), .ZN(
        P2_U3232) );
  INV_X1 U8724 ( .A(n7384), .ZN(n7389) );
  NOR3_X1 U8725 ( .A1(n7387), .A2(n7386), .A3(n7385), .ZN(n7388) );
  OAI21_X1 U8726 ( .B1(n7389), .B2(n7388), .A(n9158), .ZN(n7392) );
  NOR2_X1 U8727 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9701), .ZN(n10926) );
  OAI22_X1 U8728 ( .A1(n7478), .A2(n9125), .B1(n9231), .B2(n7689), .ZN(n7390)
         );
  AOI211_X1 U8729 ( .C1(n9219), .C2(n7579), .A(n10926), .B(n7390), .ZN(n7391)
         );
  OAI211_X1 U8730 ( .C1(n7577), .C2(n9217), .A(n7392), .B(n7391), .ZN(P2_U3167) );
  AOI22_X1 U8731 ( .A1(n10854), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n10695), .ZN(n7393) );
  OAI21_X1 U8732 ( .B1(n7411), .B2(n10704), .A(n7393), .ZN(P1_U3337) );
  NAND2_X1 U8733 ( .A1(n7396), .A2(n7395), .ZN(n8445) );
  XNOR2_X1 U8734 ( .A(n7394), .B(n8445), .ZN(n7583) );
  OR2_X1 U8735 ( .A1(n7398), .A2(n7397), .ZN(n7400) );
  NAND2_X1 U8736 ( .A1(n7400), .A2(n7399), .ZN(n7401) );
  XNOR2_X1 U8737 ( .A(n7401), .B(n8445), .ZN(n7402) );
  AOI222_X1 U8738 ( .A1(n9490), .A2(n7402), .B1(n9256), .B2(n9495), .C1(n6908), 
        .C2(n9492), .ZN(n7584) );
  OAI21_X1 U8739 ( .B1(n7403), .B2(n9565), .A(n7584), .ZN(n7404) );
  AOI21_X1 U8740 ( .B1(n9541), .B2(n7583), .A(n7404), .ZN(n11039) );
  OR2_X1 U8741 ( .A1(n9561), .A2(n5919), .ZN(n7405) );
  OAI21_X1 U8742 ( .B1(n11039), .B2(n9572), .A(n7405), .ZN(P2_U3463) );
  INV_X1 U8743 ( .A(n7406), .ZN(n7409) );
  AOI22_X1 U8744 ( .A1(n10840), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n10695), .ZN(n7407) );
  OAI21_X1 U8745 ( .B1(n7409), .B2(n10704), .A(n7407), .ZN(P1_U3338) );
  AOI22_X1 U8746 ( .A1(n10940), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_17__SCAN_IN), .B2(n9621), .ZN(n7408) );
  OAI21_X1 U8747 ( .B1(n7409), .B2(n9619), .A(n7408), .ZN(P2_U3278) );
  INV_X1 U8748 ( .A(n10979), .ZN(n10961) );
  INV_X1 U8749 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n7410) );
  OAI222_X1 U8750 ( .A1(n9109), .A2(n7411), .B1(n10961), .B2(P2_U3151), .C1(
        n7410), .C2(n9614), .ZN(P2_U3277) );
  XNOR2_X1 U8751 ( .A(n7412), .B(n7415), .ZN(n7553) );
  OAI21_X1 U8752 ( .B1(n7819), .B2(n7557), .A(n11126), .ZN(n7413) );
  NOR2_X1 U8753 ( .A1(n7413), .A2(n7840), .ZN(n7559) );
  INV_X1 U8754 ( .A(n7414), .ZN(n7417) );
  INV_X1 U8755 ( .A(n8992), .ZN(n8834) );
  AOI21_X1 U8756 ( .B1(n7812), .B2(n8834), .A(n7415), .ZN(n7416) );
  NOR2_X1 U8757 ( .A1(n7417), .A2(n7416), .ZN(n7418) );
  OAI222_X1 U8758 ( .A1(n11137), .A2(n7646), .B1(n11135), .B2(n7528), .C1(
        n11132), .C2(n7418), .ZN(n7554) );
  AOI211_X1 U8759 ( .C1(n7553), .C2(n11168), .A(n7559), .B(n7554), .ZN(n7424)
         );
  OAI22_X1 U8760 ( .A1(n10644), .A2(n7557), .B1(n11171), .B2(n7139), .ZN(n7419) );
  INV_X1 U8761 ( .A(n7419), .ZN(n7420) );
  OAI21_X1 U8762 ( .B1(n7424), .B2(n6860), .A(n7420), .ZN(P1_U3527) );
  INV_X1 U8763 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n7421) );
  OAI22_X1 U8764 ( .A1(n10685), .A2(n7557), .B1(n11175), .B2(n7421), .ZN(n7422) );
  INV_X1 U8765 ( .A(n7422), .ZN(n7423) );
  OAI21_X1 U8766 ( .B1(n7424), .B2(n11172), .A(n7423), .ZN(P1_U3468) );
  AOI21_X1 U8767 ( .B1(n7427), .B2(n6019), .A(n7591), .ZN(n7444) );
  NAND2_X1 U8768 ( .A1(P2_REG2_REG_7__SCAN_IN), .A2(n7431), .ZN(n7606) );
  OAI21_X1 U8769 ( .B1(n7431), .B2(P2_REG2_REG_7__SCAN_IN), .A(n7606), .ZN(
        n7442) );
  MUX2_X1 U8770 ( .A(P2_REG2_REG_7__SCAN_IN), .B(P2_REG1_REG_7__SCAN_IN), .S(
        n9324), .Z(n7432) );
  NOR2_X1 U8771 ( .A1(n7432), .A2(n5580), .ZN(n7598) );
  AOI21_X1 U8772 ( .B1(n7432), .B2(n5580), .A(n7598), .ZN(n7433) );
  INV_X1 U8773 ( .A(n7433), .ZN(n7437) );
  NOR2_X1 U8774 ( .A1(n7435), .A2(n7434), .ZN(n7436) );
  NOR2_X1 U8775 ( .A1(n7436), .A2(n7437), .ZN(n7597) );
  AOI21_X1 U8776 ( .B1(n7437), .B2(n7436), .A(n7597), .ZN(n7438) );
  NAND2_X1 U8777 ( .A1(P2_U3151), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n7688) );
  OAI21_X1 U8778 ( .B1(n7438), .B2(n10915), .A(n7688), .ZN(n7439) );
  AOI21_X1 U8779 ( .B1(n10965), .B2(P2_ADDR_REG_7__SCAN_IN), .A(n7439), .ZN(
        n7440) );
  OAI21_X1 U8780 ( .B1(n5580), .B2(n10976), .A(n7440), .ZN(n7441) );
  AOI21_X1 U8781 ( .B1(n10928), .B2(n7442), .A(n7441), .ZN(n7443) );
  OAI21_X1 U8782 ( .B1(n7444), .B2(n10969), .A(n7443), .ZN(P2_U3189) );
  INV_X1 U8783 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n11099) );
  AOI22_X1 U8784 ( .A1(P1_REG1_REG_12__SCAN_IN), .A2(n10382), .B1(n7463), .B2(
        n11099), .ZN(n7450) );
  INV_X1 U8785 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n7446) );
  MUX2_X1 U8786 ( .A(P1_REG1_REG_9__SCAN_IN), .B(n7446), .S(n10364), .Z(n10356) );
  OAI21_X1 U8787 ( .B1(n10364), .B2(P1_REG1_REG_9__SCAN_IN), .A(n10355), .ZN(
        n10877) );
  INV_X1 U8788 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n7447) );
  MUX2_X1 U8789 ( .A(n7447), .B(P1_REG1_REG_10__SCAN_IN), .S(n10880), .Z(
        n10876) );
  NOR2_X1 U8790 ( .A1(n10877), .A2(n10876), .ZN(n10875) );
  INV_X1 U8791 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n7448) );
  MUX2_X1 U8792 ( .A(n7448), .B(P1_REG1_REG_11__SCAN_IN), .S(n10806), .Z(
        n10802) );
  OAI21_X1 U8793 ( .B1(n7450), .B2(n7449), .A(n10371), .ZN(n7465) );
  NOR2_X1 U8794 ( .A1(P1_REG2_REG_12__SCAN_IN), .A2(n10382), .ZN(n7451) );
  AOI21_X1 U8795 ( .B1(n10382), .B2(P1_REG2_REG_12__SCAN_IN), .A(n7451), .ZN(
        n7459) );
  AOI21_X1 U8796 ( .B1(n7453), .B2(P1_REG2_REG_8__SCAN_IN), .A(n7452), .ZN(
        n10361) );
  NOR2_X1 U8797 ( .A1(n10364), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n7454) );
  AOI21_X1 U8798 ( .B1(n10364), .B2(P1_REG2_REG_9__SCAN_IN), .A(n7454), .ZN(
        n10362) );
  NAND2_X1 U8799 ( .A1(n10361), .A2(n10362), .ZN(n10360) );
  OAI21_X1 U8800 ( .B1(n10364), .B2(P1_REG2_REG_9__SCAN_IN), .A(n10360), .ZN(
        n10873) );
  INV_X1 U8801 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n7455) );
  AOI22_X1 U8802 ( .A1(P1_REG2_REG_10__SCAN_IN), .A2(n7456), .B1(n10880), .B2(
        n7455), .ZN(n10872) );
  NOR2_X1 U8803 ( .A1(n10873), .A2(n10872), .ZN(n10871) );
  AOI21_X1 U8804 ( .B1(n10880), .B2(P1_REG2_REG_10__SCAN_IN), .A(n10871), .ZN(
        n10800) );
  NAND2_X1 U8805 ( .A1(n10806), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n7457) );
  OAI21_X1 U8806 ( .B1(n10806), .B2(P1_REG2_REG_11__SCAN_IN), .A(n7457), .ZN(
        n10799) );
  NOR2_X1 U8807 ( .A1(n10800), .A2(n10799), .ZN(n10798) );
  AOI21_X1 U8808 ( .B1(P1_REG2_REG_11__SCAN_IN), .B2(n10806), .A(n10798), .ZN(
        n7458) );
  NAND2_X1 U8809 ( .A1(n7459), .A2(n7458), .ZN(n10381) );
  OAI21_X1 U8810 ( .B1(n7459), .B2(n7458), .A(n10381), .ZN(n7460) );
  NAND2_X1 U8811 ( .A1(n7460), .A2(n10841), .ZN(n7462) );
  AND2_X1 U8812 ( .A1(P1_U3086), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n10117) );
  AOI21_X1 U8813 ( .B1(n10868), .B2(P1_ADDR_REG_12__SCAN_IN), .A(n10117), .ZN(
        n7461) );
  OAI211_X1 U8814 ( .C1(n10414), .C2(n7463), .A(n7462), .B(n7461), .ZN(n7464)
         );
  AOI21_X1 U8815 ( .B1(n10838), .B2(n7465), .A(n7464), .ZN(n7466) );
  INV_X1 U8816 ( .A(n7466), .ZN(P1_U3255) );
  NAND2_X1 U8817 ( .A1(n7968), .A2(n7467), .ZN(n11110) );
  OAI22_X1 U8818 ( .A1(n9441), .A2(n7468), .B1(P2_REG3_REG_3__SCAN_IN), .B2(
        n11104), .ZN(n7471) );
  MUX2_X1 U8819 ( .A(P2_REG2_REG_3__SCAN_IN), .B(n7469), .S(n11111), .Z(n7470)
         );
  AOI211_X1 U8820 ( .C1(n9443), .C2(n7472), .A(n7471), .B(n7470), .ZN(n7473)
         );
  INV_X1 U8821 ( .A(n7473), .ZN(P2_U3230) );
  NAND2_X1 U8822 ( .A1(n8515), .A2(n8516), .ZN(n7476) );
  INV_X1 U8823 ( .A(n7476), .ZN(n8449) );
  XNOR2_X1 U8824 ( .A(n7474), .B(n8449), .ZN(n7582) );
  NOR2_X1 U8825 ( .A1(n7582), .A2(n9567), .ZN(n7479) );
  XNOR2_X1 U8826 ( .A(n7475), .B(n7476), .ZN(n7477) );
  OAI222_X1 U8827 ( .A1(n9476), .A2(n7689), .B1(n9474), .B2(n7478), .C1(n7477), 
        .C2(n9471), .ZN(n7574) );
  AOI211_X1 U8828 ( .C1(n9553), .C2(n7579), .A(n7479), .B(n7574), .ZN(n11050)
         );
  OR2_X1 U8829 ( .A1(n11050), .A2(n9572), .ZN(n7480) );
  OAI21_X1 U8830 ( .B1(n9561), .B2(n7262), .A(n7480), .ZN(P2_U3464) );
  INV_X1 U8831 ( .A(n7481), .ZN(n7482) );
  NAND2_X1 U8832 ( .A1(n7483), .A2(n7482), .ZN(n7490) );
  NAND2_X1 U8833 ( .A1(n7493), .A2(n7490), .ZN(n7487) );
  INV_X2 U8834 ( .A(n7484), .ZN(n8808) );
  NAND2_X1 U8835 ( .A1(n8808), .A2(n7545), .ZN(n7485) );
  OAI21_X1 U8836 ( .B1(n7833), .B2(n5152), .A(n7485), .ZN(n7486) );
  XNOR2_X1 U8837 ( .A(n7486), .B(n8809), .ZN(n7489) );
  NAND2_X1 U8838 ( .A1(n7487), .A2(n7489), .ZN(n7540) );
  OAI22_X1 U8839 ( .A1(n7833), .A2(n8806), .B1(n7557), .B2(n5152), .ZN(n7541)
         );
  INV_X1 U8840 ( .A(n7541), .ZN(n7488) );
  NAND2_X1 U8841 ( .A1(n7540), .A2(n7488), .ZN(n7617) );
  INV_X1 U8842 ( .A(n7489), .ZN(n7491) );
  AND2_X1 U8843 ( .A1(n7491), .A2(n7490), .ZN(n7492) );
  NAND2_X1 U8844 ( .A1(n7493), .A2(n7492), .ZN(n7615) );
  NAND2_X1 U8845 ( .A1(n7617), .A2(n7615), .ZN(n7503) );
  NAND2_X1 U8846 ( .A1(n10292), .A2(n5136), .ZN(n7494) );
  OAI21_X1 U8847 ( .B1(n7484), .B2(n11053), .A(n7494), .ZN(n7495) );
  XNOR2_X1 U8848 ( .A(n7495), .B(n8781), .ZN(n7499) );
  OR2_X1 U8849 ( .A1(n11053), .A2(n5152), .ZN(n7497) );
  NAND2_X1 U8850 ( .A1(n10292), .A2(n8692), .ZN(n7496) );
  NAND2_X1 U8851 ( .A1(n7497), .A2(n7496), .ZN(n7500) );
  INV_X1 U8852 ( .A(n7500), .ZN(n7498) );
  NAND2_X1 U8853 ( .A1(n7499), .A2(n7498), .ZN(n7614) );
  INV_X1 U8854 ( .A(n7499), .ZN(n7501) );
  NAND2_X1 U8855 ( .A1(n7501), .A2(n7500), .ZN(n7628) );
  NAND2_X1 U8856 ( .A1(n7614), .A2(n7628), .ZN(n7502) );
  XNOR2_X1 U8857 ( .A(n7503), .B(n7502), .ZN(n7509) );
  INV_X1 U8858 ( .A(n11053), .ZN(n7842) );
  INV_X1 U8859 ( .A(n7504), .ZN(n7506) );
  OAI22_X1 U8860 ( .A1(n10236), .A2(n7833), .B1(n7834), .B2(n10259), .ZN(n7505) );
  AOI211_X1 U8861 ( .C1(n7842), .C2(n10266), .A(n7506), .B(n7505), .ZN(n7508)
         );
  NAND2_X1 U8862 ( .A1(n10250), .A2(n7841), .ZN(n7507) );
  OAI211_X1 U8863 ( .C1(n7509), .C2(n10269), .A(n7508), .B(n7507), .ZN(
        P1_U3239) );
  XOR2_X1 U8864 ( .A(n7510), .B(n8450), .Z(n7670) );
  XOR2_X1 U8865 ( .A(n8450), .B(n7511), .Z(n7512) );
  OAI222_X1 U8866 ( .A1(n9476), .A2(n7774), .B1(n9474), .B2(n7513), .C1(n7512), 
        .C2(n9471), .ZN(n7671) );
  INV_X1 U8867 ( .A(n7671), .ZN(n7514) );
  MUX2_X1 U8868 ( .A(n7515), .B(n7514), .S(n11111), .Z(n7519) );
  INV_X1 U8869 ( .A(n7516), .ZN(n7517) );
  AOI22_X1 U8870 ( .A1(n9509), .A2(n7673), .B1(n9439), .B2(n7517), .ZN(n7518)
         );
  OAI211_X1 U8871 ( .C1(n9505), .C2(n7670), .A(n7519), .B(n7518), .ZN(P2_U3227) );
  AND2_X1 U8872 ( .A1(n7521), .A2(n7520), .ZN(n7523) );
  OAI21_X1 U8873 ( .B1(n7523), .B2(n8849), .A(n7522), .ZN(n7802) );
  INV_X1 U8874 ( .A(n7802), .ZN(n7539) );
  OR2_X1 U8875 ( .A1(n11011), .A2(n7551), .ZN(n7838) );
  INV_X1 U8876 ( .A(n8849), .ZN(n7527) );
  AND2_X1 U8877 ( .A1(n7525), .A2(n7524), .ZN(n7526) );
  NAND2_X1 U8878 ( .A1(n7526), .A2(n7527), .ZN(n7860) );
  OAI21_X1 U8879 ( .B1(n7527), .B2(n7526), .A(n7860), .ZN(n7530) );
  OAI22_X1 U8880 ( .A1(n7528), .A2(n11137), .B1(n10170), .B2(n11135), .ZN(
        n7529) );
  AOI21_X1 U8881 ( .B1(n7530), .B2(n10566), .A(n7529), .ZN(n7531) );
  OAI21_X1 U8882 ( .B1(n7539), .B2(n7711), .A(n7531), .ZN(n7800) );
  NAND2_X1 U8883 ( .A1(n7800), .A2(n10560), .ZN(n7538) );
  INV_X1 U8884 ( .A(n7532), .ZN(n7717) );
  AOI211_X1 U8885 ( .C1(n7639), .C2(n7839), .A(n10577), .B(n7717), .ZN(n7801)
         );
  INV_X1 U8886 ( .A(n7637), .ZN(n7534) );
  AOI22_X1 U8887 ( .A1(n11011), .A2(P1_REG2_REG_7__SCAN_IN), .B1(n7534), .B2(
        n11149), .ZN(n7535) );
  OAI21_X1 U8888 ( .B1(n11014), .B2(n5298), .A(n7535), .ZN(n7536) );
  AOI21_X1 U8889 ( .B1(n7801), .B2(n11018), .A(n7536), .ZN(n7537) );
  OAI211_X1 U8890 ( .C1(n7539), .C2(n7838), .A(n7538), .B(n7537), .ZN(P1_U3286) );
  NAND2_X1 U8891 ( .A1(n7615), .A2(n7540), .ZN(n7542) );
  XNOR2_X1 U8892 ( .A(n7542), .B(n7541), .ZN(n7549) );
  AOI22_X1 U8893 ( .A1(n10233), .A2(n10292), .B1(n10261), .B2(n10294), .ZN(
        n7547) );
  INV_X1 U8894 ( .A(n7543), .ZN(n7544) );
  AOI21_X1 U8895 ( .B1(n10266), .B2(n7545), .A(n7544), .ZN(n7546) );
  OAI211_X1 U8896 ( .C1(n10263), .C2(n7556), .A(n7547), .B(n7546), .ZN(n7548)
         );
  AOI21_X1 U8897 ( .B1(n7549), .B2(n10244), .A(n7548), .ZN(n7550) );
  INV_X1 U8898 ( .A(n7550), .ZN(P1_U3227) );
  AND2_X1 U8899 ( .A1(n7711), .A2(n7551), .ZN(n7552) );
  INV_X1 U8900 ( .A(n7553), .ZN(n7562) );
  INV_X1 U8901 ( .A(n7554), .ZN(n7555) );
  MUX2_X1 U8902 ( .A(n7153), .B(n7555), .S(n10560), .Z(n7561) );
  OAI22_X1 U8903 ( .A1(n11014), .A2(n7557), .B1(n7556), .B2(n10580), .ZN(n7558) );
  AOI21_X1 U8904 ( .B1(n7559), .B2(n11018), .A(n7558), .ZN(n7560) );
  OAI211_X1 U8905 ( .C1(n10563), .C2(n7562), .A(n7561), .B(n7560), .ZN(
        P1_U3288) );
  INV_X1 U8906 ( .A(n7563), .ZN(n7564) );
  AOI21_X1 U8907 ( .B1(n7566), .B2(n7565), .A(n7564), .ZN(n7679) );
  XNOR2_X1 U8908 ( .A(n7567), .B(n8521), .ZN(n7568) );
  OAI222_X1 U8909 ( .A1(n9476), .A2(n7936), .B1(n9474), .B2(n7689), .C1(n9471), 
        .C2(n7568), .ZN(n7676) );
  AOI21_X1 U8910 ( .B1(n7679), .B2(n9541), .A(n7676), .ZN(n7573) );
  INV_X1 U8911 ( .A(n9564), .ZN(n8024) );
  AOI22_X1 U8912 ( .A1(n8024), .A2(n7684), .B1(n9572), .B2(
        P2_REG1_REG_7__SCAN_IN), .ZN(n7569) );
  OAI21_X1 U8913 ( .B1(n7573), .B2(n9572), .A(n7569), .ZN(P2_U3466) );
  INV_X1 U8914 ( .A(n7684), .ZN(n7695) );
  INV_X1 U8915 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n7570) );
  OAI22_X1 U8916 ( .A1(n9607), .A2(n7695), .B1(n11178), .B2(n7570), .ZN(n7571)
         );
  INV_X1 U8917 ( .A(n7571), .ZN(n7572) );
  OAI21_X1 U8918 ( .B1(n7573), .B2(n6432), .A(n7572), .ZN(P2_U3411) );
  INV_X1 U8919 ( .A(n7574), .ZN(n7575) );
  MUX2_X1 U8920 ( .A(n7576), .B(n7575), .S(n11111), .Z(n7581) );
  INV_X1 U8921 ( .A(n7577), .ZN(n7578) );
  AOI22_X1 U8922 ( .A1(n9509), .A2(n7579), .B1(n9439), .B2(n7578), .ZN(n7580)
         );
  OAI211_X1 U8923 ( .C1(n7582), .C2(n9505), .A(n7581), .B(n7580), .ZN(P2_U3228) );
  INV_X1 U8924 ( .A(n7583), .ZN(n7590) );
  MUX2_X1 U8925 ( .A(n7585), .B(n7584), .S(n11111), .Z(n7589) );
  AOI22_X1 U8926 ( .A1(n9509), .A2(n7587), .B1(n9439), .B2(n7586), .ZN(n7588)
         );
  OAI211_X1 U8927 ( .C1(n7590), .C2(n9505), .A(n7589), .B(n7588), .ZN(P2_U3229) );
  NAND2_X1 U8928 ( .A1(P2_REG1_REG_8__SCAN_IN), .A2(n7758), .ZN(n7747) );
  OAI21_X1 U8929 ( .B1(n7758), .B2(P2_REG1_REG_8__SCAN_IN), .A(n7747), .ZN(
        n7592) );
  NOR2_X1 U8930 ( .A1(n7593), .A2(n7592), .ZN(n7749) );
  AOI21_X1 U8931 ( .B1(n7593), .B2(n7592), .A(n7749), .ZN(n7613) );
  INV_X1 U8932 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n7594) );
  NOR2_X1 U8933 ( .A1(n10938), .A2(n7594), .ZN(n7604) );
  MUX2_X1 U8934 ( .A(P2_REG2_REG_8__SCAN_IN), .B(P2_REG1_REG_8__SCAN_IN), .S(
        n9324), .Z(n7595) );
  NOR2_X1 U8935 ( .A1(n7595), .A2(n7758), .ZN(n7738) );
  AOI21_X1 U8936 ( .B1(n7595), .B2(n7758), .A(n7738), .ZN(n7596) );
  INV_X1 U8937 ( .A(n7596), .ZN(n7600) );
  NOR2_X1 U8938 ( .A1(n7598), .A2(n7597), .ZN(n7599) );
  NOR2_X1 U8939 ( .A1(n7599), .A2(n7600), .ZN(n7737) );
  AOI21_X1 U8940 ( .B1(n7600), .B2(n7599), .A(n7737), .ZN(n7602) );
  NOR2_X1 U8941 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9896), .ZN(n7776) );
  INV_X1 U8942 ( .A(n7776), .ZN(n7601) );
  OAI21_X1 U8943 ( .B1(n7602), .B2(n10915), .A(n7601), .ZN(n7603) );
  AOI211_X1 U8944 ( .C1(n10941), .C2(n9620), .A(n7604), .B(n7603), .ZN(n7612)
         );
  AOI22_X1 U8945 ( .A1(n9620), .A2(n7666), .B1(P2_REG2_REG_8__SCAN_IN), .B2(
        n7758), .ZN(n7609) );
  NAND2_X1 U8946 ( .A1(n7605), .A2(n5580), .ZN(n7607) );
  NAND2_X1 U8947 ( .A1(n7607), .A2(n7606), .ZN(n7608) );
  NAND2_X1 U8948 ( .A1(n7609), .A2(n7608), .ZN(n7759) );
  OAI21_X1 U8949 ( .B1(n7609), .B2(n7608), .A(n7759), .ZN(n7610) );
  NAND2_X1 U8950 ( .A1(n7610), .A2(n10928), .ZN(n7611) );
  OAI211_X1 U8951 ( .C1(n7613), .C2(n10969), .A(n7612), .B(n7611), .ZN(
        P2_U3190) );
  AND2_X1 U8952 ( .A1(n7615), .A2(n7614), .ZN(n7616) );
  NAND2_X1 U8953 ( .A1(n7617), .A2(n7616), .ZN(n7630) );
  NAND2_X1 U8954 ( .A1(n7630), .A2(n7628), .ZN(n7633) );
  NAND2_X1 U8955 ( .A1(n7639), .A2(n8808), .ZN(n7618) );
  OAI21_X1 U8956 ( .B1(n7834), .B2(n5152), .A(n7618), .ZN(n7619) );
  XNOR2_X1 U8957 ( .A(n7619), .B(n8781), .ZN(n7622) );
  NAND2_X1 U8958 ( .A1(n5297), .A2(n8692), .ZN(n7621) );
  NAND2_X1 U8959 ( .A1(n7639), .A2(n5136), .ZN(n7620) );
  AND2_X1 U8960 ( .A1(n7621), .A2(n7620), .ZN(n7623) );
  NAND2_X1 U8961 ( .A1(n7622), .A2(n7623), .ZN(n8634) );
  INV_X1 U8962 ( .A(n7622), .ZN(n7625) );
  INV_X1 U8963 ( .A(n7623), .ZN(n7624) );
  NAND2_X1 U8964 ( .A1(n7625), .A2(n7624), .ZN(n7626) );
  NAND2_X1 U8965 ( .A1(n8634), .A2(n7626), .ZN(n7632) );
  INV_X1 U8966 ( .A(n7632), .ZN(n7627) );
  AND2_X1 U8967 ( .A1(n7628), .A2(n7627), .ZN(n7629) );
  NAND2_X1 U8968 ( .A1(n7630), .A2(n7629), .ZN(n8635) );
  INV_X1 U8969 ( .A(n8635), .ZN(n7631) );
  AOI21_X1 U8970 ( .B1(n7633), .B2(n7632), .A(n7631), .ZN(n7641) );
  AOI21_X1 U8971 ( .B1(n10233), .B2(n10291), .A(n7634), .ZN(n7636) );
  NAND2_X1 U8972 ( .A1(n10261), .A2(n10292), .ZN(n7635) );
  OAI211_X1 U8973 ( .C1(n10263), .C2(n7637), .A(n7636), .B(n7635), .ZN(n7638)
         );
  AOI21_X1 U8974 ( .B1(n7639), .B2(n10266), .A(n7638), .ZN(n7640) );
  OAI21_X1 U8975 ( .B1(n7641), .B2(n10269), .A(n7640), .ZN(P1_U3213) );
  XNOR2_X1 U8976 ( .A(n7642), .B(n7645), .ZN(n11030) );
  OAI21_X1 U8977 ( .B1(n7645), .B2(n7644), .A(n7643), .ZN(n7648) );
  OAI22_X1 U8978 ( .A1(n7646), .A2(n11135), .B1(n6483), .B2(n11137), .ZN(n7647) );
  AOI21_X1 U8979 ( .B1(n7648), .B2(n10566), .A(n7647), .ZN(n7649) );
  OAI21_X1 U8980 ( .B1(n11030), .B2(n7711), .A(n7649), .ZN(n11033) );
  NAND2_X1 U8981 ( .A1(n11033), .A2(n10560), .ZN(n7656) );
  INV_X1 U8982 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n7650) );
  OAI22_X1 U8983 ( .A1(n10560), .A2(n7650), .B1(P1_REG3_REG_3__SCAN_IN), .B2(
        n10580), .ZN(n7653) );
  INV_X1 U8984 ( .A(n10995), .ZN(n7651) );
  OAI211_X1 U8985 ( .C1(n7651), .C2(n11032), .A(n11126), .B(n7816), .ZN(n11031) );
  NOR2_X1 U8986 ( .A1(n11031), .A2(n11153), .ZN(n7652) );
  AOI211_X1 U8987 ( .C1(n11151), .C2(n7654), .A(n7653), .B(n7652), .ZN(n7655)
         );
  OAI211_X1 U8988 ( .C1(n11030), .C2(n7838), .A(n7656), .B(n7655), .ZN(
        P1_U3290) );
  INV_X1 U8989 ( .A(n7657), .ZN(n7659) );
  INV_X1 U8990 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n7658) );
  OAI222_X1 U8991 ( .A1(n6812), .A2(P1_U3086), .B1(n10704), .B2(n7659), .C1(
        n7658), .C2(n10701), .ZN(P1_U3336) );
  INV_X1 U8992 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n7660) );
  OAI222_X1 U8993 ( .A1(n9614), .A2(n7660), .B1(n9619), .B2(n7659), .C1(
        P2_U3151), .C2(n9334), .ZN(P2_U3276) );
  NAND2_X1 U8994 ( .A1(n7563), .A2(n7661), .ZN(n7662) );
  XOR2_X1 U8995 ( .A(n8453), .B(n7662), .Z(n7943) );
  XOR2_X1 U8996 ( .A(n7663), .B(n8453), .Z(n7664) );
  OAI222_X1 U8997 ( .A1(n9476), .A2(n8050), .B1(n9474), .B2(n7774), .C1(n9471), 
        .C2(n7664), .ZN(n7944) );
  INV_X1 U8998 ( .A(n7944), .ZN(n7665) );
  MUX2_X1 U8999 ( .A(n7666), .B(n7665), .S(n11111), .Z(n7669) );
  AOI22_X1 U9000 ( .A1(n7946), .A2(n9509), .B1(n9439), .B2(n7667), .ZN(n7668)
         );
  OAI211_X1 U9001 ( .C1(n7943), .C2(n9505), .A(n7669), .B(n7668), .ZN(P2_U3225) );
  NOR2_X1 U9002 ( .A1(n7670), .A2(n9567), .ZN(n7672) );
  AOI211_X1 U9003 ( .C1(n9553), .C2(n7673), .A(n7672), .B(n7671), .ZN(n11051)
         );
  OR2_X1 U9004 ( .A1(n11051), .A2(n9572), .ZN(n7674) );
  OAI21_X1 U9005 ( .B1(n9561), .B2(n7675), .A(n7674), .ZN(P2_U3465) );
  OAI22_X1 U9006 ( .A1(n7695), .A2(n9441), .B1(n7690), .B2(n11104), .ZN(n7678)
         );
  MUX2_X1 U9007 ( .A(P2_REG2_REG_7__SCAN_IN), .B(n7676), .S(n11111), .Z(n7677)
         );
  AOI211_X1 U9008 ( .C1(n9443), .C2(n7679), .A(n7678), .B(n7677), .ZN(n7680)
         );
  INV_X1 U9009 ( .A(n7680), .ZN(P2_U3226) );
  INV_X1 U9010 ( .A(n7681), .ZN(n7682) );
  XNOR2_X1 U9011 ( .A(n7684), .B(n6905), .ZN(n7770) );
  XNOR2_X1 U9012 ( .A(n7770), .B(n9254), .ZN(n7685) );
  OAI21_X1 U9013 ( .B1(n7686), .B2(n7685), .A(n7772), .ZN(n7687) );
  NAND2_X1 U9014 ( .A1(n7687), .A2(n9158), .ZN(n7694) );
  OAI21_X1 U9015 ( .B1(n9125), .B2(n7689), .A(n7688), .ZN(n7692) );
  NOR2_X1 U9016 ( .A1(n9217), .A2(n7690), .ZN(n7691) );
  AOI211_X1 U9017 ( .C1(n9214), .C2(n9253), .A(n7692), .B(n7691), .ZN(n7693)
         );
  OAI211_X1 U9018 ( .C1(n7695), .C2(n9238), .A(n7694), .B(n7693), .ZN(P2_U3153) );
  OR2_X1 U9019 ( .A1(n7697), .A2(n7696), .ZN(n7698) );
  NAND2_X1 U9020 ( .A1(n7891), .A2(n7698), .ZN(n7700) );
  OAI22_X1 U9021 ( .A1(n10096), .A2(n11137), .B1(n10119), .B2(n11135), .ZN(
        n7699) );
  AOI21_X1 U9022 ( .B1(n7700), .B2(n10566), .A(n7699), .ZN(n11076) );
  OAI21_X1 U9023 ( .B1(n7702), .B2(n8940), .A(n7701), .ZN(n11079) );
  NAND2_X1 U9024 ( .A1(n11079), .A2(n10575), .ZN(n7707) );
  OAI22_X1 U9025 ( .A1(n10560), .A2(n7455), .B1(n10078), .B2(n10580), .ZN(
        n7705) );
  INV_X1 U9026 ( .A(n7869), .ZN(n7716) );
  OAI21_X1 U9027 ( .B1(n7716), .B2(n10172), .A(n10080), .ZN(n7703) );
  NAND3_X1 U9028 ( .A1(n7703), .A2(n11126), .A3(n7897), .ZN(n11075) );
  NOR2_X1 U9029 ( .A1(n11075), .A2(n11153), .ZN(n7704) );
  AOI211_X1 U9030 ( .C1(n11151), .C2(n10080), .A(n7705), .B(n7704), .ZN(n7706)
         );
  OAI211_X1 U9031 ( .C1(n11011), .C2(n11076), .A(n7707), .B(n7706), .ZN(
        P1_U3283) );
  OAI21_X1 U9032 ( .B1(n7709), .B2(n8853), .A(n7708), .ZN(n11064) );
  INV_X1 U9033 ( .A(n11064), .ZN(n7722) );
  NAND2_X1 U9034 ( .A1(n7860), .A2(n8935), .ZN(n7710) );
  XNOR2_X1 U9035 ( .A(n7710), .B(n8853), .ZN(n7714) );
  INV_X1 U9036 ( .A(n7711), .ZN(n11141) );
  OAI22_X1 U9037 ( .A1(n10096), .A2(n11135), .B1(n7834), .B2(n11137), .ZN(
        n7712) );
  AOI21_X1 U9038 ( .B1(n11064), .B2(n11141), .A(n7712), .ZN(n7713) );
  OAI21_X1 U9039 ( .B1(n11132), .B2(n7714), .A(n7713), .ZN(n11062) );
  NAND2_X1 U9040 ( .A1(n11062), .A2(n10560), .ZN(n7721) );
  INV_X1 U9041 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n7715) );
  OAI22_X1 U9042 ( .A1(n10560), .A2(n7715), .B1(n10099), .B2(n10580), .ZN(
        n7719) );
  INV_X1 U9043 ( .A(n10101), .ZN(n11061) );
  OAI211_X1 U9044 ( .C1(n11061), .C2(n7717), .A(n7716), .B(n11126), .ZN(n11060) );
  NOR2_X1 U9045 ( .A1(n11060), .A2(n11153), .ZN(n7718) );
  AOI211_X1 U9046 ( .C1(n11151), .C2(n10101), .A(n7719), .B(n7718), .ZN(n7720)
         );
  OAI211_X1 U9047 ( .C1(n7722), .C2(n7838), .A(n7721), .B(n7720), .ZN(P1_U3285) );
  XNOR2_X1 U9048 ( .A(n8928), .B(n7723), .ZN(n10990) );
  INV_X1 U9049 ( .A(n10990), .ZN(n7736) );
  INV_X1 U9050 ( .A(n10996), .ZN(n7724) );
  OAI211_X1 U9051 ( .C1(n10987), .C2(n7725), .A(n7724), .B(n11126), .ZN(n10986) );
  NOR2_X1 U9052 ( .A1(n11153), .A2(n10986), .ZN(n7728) );
  INV_X1 U9053 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n7726) );
  OAI22_X1 U9054 ( .A1(n10560), .A2(n6453), .B1(n7726), .B2(n10580), .ZN(n7727) );
  AOI211_X1 U9055 ( .C1(n11151), .C2(n7729), .A(n7728), .B(n7727), .ZN(n7735)
         );
  XNOR2_X1 U9056 ( .A(n7730), .B(n8928), .ZN(n7733) );
  NAND2_X1 U9057 ( .A1(n10990), .A2(n11141), .ZN(n7732) );
  AOI22_X1 U9058 ( .A1(n10999), .A2(n10297), .B1(n10295), .B2(n11002), .ZN(
        n7731) );
  OAI211_X1 U9059 ( .C1(n7733), .C2(n11132), .A(n7732), .B(n7731), .ZN(n10988)
         );
  NAND2_X1 U9060 ( .A1(n10988), .A2(n10560), .ZN(n7734) );
  OAI211_X1 U9061 ( .C1(n7736), .C2(n7838), .A(n7735), .B(n7734), .ZN(P1_U3292) );
  MUX2_X1 U9062 ( .A(P2_REG2_REG_9__SCAN_IN), .B(P2_REG1_REG_9__SCAN_IN), .S(
        n9324), .Z(n7739) );
  NOR2_X1 U9063 ( .A1(n7739), .A2(n7798), .ZN(n7741) );
  NOR2_X1 U9064 ( .A1(n7738), .A2(n7737), .ZN(n7786) );
  AOI21_X1 U9065 ( .B1(n7739), .B2(n7798), .A(n7741), .ZN(n7740) );
  INV_X1 U9066 ( .A(n7740), .ZN(n7787) );
  NOR2_X1 U9067 ( .A1(n7786), .A2(n7787), .ZN(n7785) );
  NOR2_X1 U9068 ( .A1(n7741), .A2(n7785), .ZN(n7982) );
  MUX2_X1 U9069 ( .A(n7743), .B(n7742), .S(n9324), .Z(n7744) );
  AND2_X1 U9070 ( .A1(n7744), .A2(n7757), .ZN(n7980) );
  NOR2_X1 U9071 ( .A1(n7744), .A2(n7757), .ZN(n7983) );
  NOR2_X1 U9072 ( .A1(n7980), .A2(n7983), .ZN(n7745) );
  XNOR2_X1 U9073 ( .A(n7982), .B(n7745), .ZN(n7769) );
  INV_X1 U9074 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n7746) );
  NAND2_X1 U9075 ( .A1(P2_U3151), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n8049) );
  OAI21_X1 U9076 ( .B1(n10938), .B2(n7746), .A(n8049), .ZN(n7756) );
  INV_X1 U9077 ( .A(n7747), .ZN(n7748) );
  INV_X1 U9078 ( .A(n7750), .ZN(n7751) );
  NAND2_X1 U9079 ( .A1(P2_REG1_REG_10__SCAN_IN), .A2(n7989), .ZN(n7752) );
  OAI21_X1 U9080 ( .B1(n7989), .B2(P2_REG1_REG_10__SCAN_IN), .A(n7752), .ZN(
        n7753) );
  AOI21_X1 U9081 ( .B1(n5216), .B2(n7753), .A(n7988), .ZN(n7754) );
  NOR2_X1 U9082 ( .A1(n10969), .A2(n7754), .ZN(n7755) );
  AOI211_X1 U9083 ( .C1(n10941), .C2(n7757), .A(n7756), .B(n7755), .ZN(n7768)
         );
  AOI22_X1 U9084 ( .A1(n7757), .A2(n7743), .B1(P2_REG2_REG_10__SCAN_IN), .B2(
        n7989), .ZN(n7765) );
  NAND2_X1 U9085 ( .A1(P2_REG2_REG_8__SCAN_IN), .A2(n7758), .ZN(n7760) );
  NAND2_X1 U9086 ( .A1(n7760), .A2(n7759), .ZN(n7762) );
  NAND2_X1 U9087 ( .A1(n7762), .A2(n7798), .ZN(n7763) );
  XNOR2_X1 U9088 ( .A(n7762), .B(n7761), .ZN(n7783) );
  NAND2_X1 U9089 ( .A1(n7763), .A2(n7782), .ZN(n7764) );
  NAND2_X1 U9090 ( .A1(n7765), .A2(n7764), .ZN(n7977) );
  OAI21_X1 U9091 ( .B1(n7765), .B2(n7764), .A(n7977), .ZN(n7766) );
  NAND2_X1 U9092 ( .A1(n7766), .A2(n10928), .ZN(n7767) );
  OAI211_X1 U9093 ( .C1(n7769), .C2(n10915), .A(n7768), .B(n7767), .ZN(
        P2_U3192) );
  NAND2_X1 U9094 ( .A1(n7770), .A2(n7774), .ZN(n7771) );
  NAND2_X1 U9095 ( .A1(n7772), .A2(n7771), .ZN(n7931) );
  XNOR2_X1 U9096 ( .A(n7946), .B(n9098), .ZN(n7928) );
  XNOR2_X1 U9097 ( .A(n7928), .B(n9253), .ZN(n7773) );
  XNOR2_X1 U9098 ( .A(n7931), .B(n7773), .ZN(n7781) );
  NOR2_X1 U9099 ( .A1(n9125), .A2(n7774), .ZN(n7775) );
  AOI211_X1 U9100 ( .C1(n9214), .C2(n9252), .A(n7776), .B(n7775), .ZN(n7777)
         );
  OAI21_X1 U9101 ( .B1(n7778), .B2(n9217), .A(n7777), .ZN(n7779) );
  AOI21_X1 U9102 ( .B1(n9219), .B2(n7946), .A(n7779), .ZN(n7780) );
  OAI21_X1 U9103 ( .B1(n7781), .B2(n9224), .A(n7780), .ZN(P2_U3161) );
  OAI21_X1 U9104 ( .B1(n7783), .B2(P2_REG2_REG_9__SCAN_IN), .A(n7782), .ZN(
        n7784) );
  NAND2_X1 U9105 ( .A1(n7784), .A2(n10928), .ZN(n7797) );
  AOI21_X1 U9106 ( .B1(n7787), .B2(n7786), .A(n7785), .ZN(n7788) );
  NAND2_X1 U9107 ( .A1(P2_U3151), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n7935) );
  OAI21_X1 U9108 ( .B1(n7788), .B2(n10915), .A(n7935), .ZN(n7795) );
  AOI21_X1 U9109 ( .B1(n6054), .B2(n7790), .A(n7789), .ZN(n7791) );
  NOR2_X1 U9110 ( .A1(n10969), .A2(n7791), .ZN(n7794) );
  INV_X1 U9111 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n7792) );
  NOR2_X1 U9112 ( .A1(n10938), .A2(n7792), .ZN(n7793) );
  NOR3_X1 U9113 ( .A1(n7795), .A2(n7794), .A3(n7793), .ZN(n7796) );
  OAI211_X1 U9114 ( .C1(n10976), .C2(n7798), .A(n7797), .B(n7796), .ZN(
        P2_U3191) );
  AOI211_X1 U9115 ( .C1(n11144), .C2(n7802), .A(n7801), .B(n7800), .ZN(n7809)
         );
  INV_X1 U9116 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n7803) );
  OAI22_X1 U9117 ( .A1(n10685), .A2(n5298), .B1(n11175), .B2(n7803), .ZN(n7804) );
  INV_X1 U9118 ( .A(n7804), .ZN(n7805) );
  OAI21_X1 U9119 ( .B1(n7809), .B2(n11172), .A(n7805), .ZN(P1_U3474) );
  INV_X1 U9120 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n7806) );
  OAI22_X1 U9121 ( .A1(n10644), .A2(n5298), .B1(n11171), .B2(n7806), .ZN(n7807) );
  INV_X1 U9122 ( .A(n7807), .ZN(n7808) );
  OAI21_X1 U9123 ( .B1(n7809), .B2(n6860), .A(n7808), .ZN(P1_U3529) );
  NAND2_X1 U9124 ( .A1(n8842), .A2(n8834), .ZN(n8931) );
  AOI21_X1 U9125 ( .B1(n7810), .B2(n8931), .A(n11132), .ZN(n7811) );
  OAI21_X1 U9126 ( .B1(n7812), .B2(n8992), .A(n7811), .ZN(n7814) );
  AOI22_X1 U9127 ( .A1(n10293), .A2(n11002), .B1(n10999), .B2(n11001), .ZN(
        n7813) );
  NAND2_X1 U9128 ( .A1(n7814), .A2(n7813), .ZN(n11044) );
  INV_X1 U9129 ( .A(n11044), .ZN(n7826) );
  XNOR2_X1 U9130 ( .A(n7815), .B(n8931), .ZN(n11040) );
  NAND2_X1 U9131 ( .A1(n7816), .A2(n7821), .ZN(n7817) );
  NAND2_X1 U9132 ( .A1(n7817), .A2(n11126), .ZN(n7818) );
  OR2_X1 U9133 ( .A1(n7819), .A2(n7818), .ZN(n11041) );
  AOI22_X1 U9134 ( .A1(n11011), .A2(P1_REG2_REG_4__SCAN_IN), .B1(n7820), .B2(
        n11149), .ZN(n7823) );
  NAND2_X1 U9135 ( .A1(n11151), .A2(n7821), .ZN(n7822) );
  OAI211_X1 U9136 ( .C1(n11041), .C2(n11153), .A(n7823), .B(n7822), .ZN(n7824)
         );
  AOI21_X1 U9137 ( .B1(n11040), .B2(n10575), .A(n7824), .ZN(n7825) );
  OAI21_X1 U9138 ( .B1(n7826), .B2(n11011), .A(n7825), .ZN(P1_U3289) );
  XNOR2_X1 U9139 ( .A(n7827), .B(n7831), .ZN(n7837) );
  NAND2_X1 U9140 ( .A1(n7829), .A2(n7828), .ZN(n7832) );
  NAND2_X1 U9141 ( .A1(n7832), .A2(n7831), .ZN(n7830) );
  OAI21_X1 U9142 ( .B1(n7832), .B2(n7831), .A(n7830), .ZN(n11056) );
  OAI22_X1 U9143 ( .A1(n7834), .A2(n11135), .B1(n7833), .B2(n11137), .ZN(n7835) );
  AOI21_X1 U9144 ( .B1(n11056), .B2(n11141), .A(n7835), .ZN(n7836) );
  OAI21_X1 U9145 ( .B1(n11132), .B2(n7837), .A(n7836), .ZN(n11054) );
  INV_X1 U9146 ( .A(n11054), .ZN(n7847) );
  INV_X1 U9147 ( .A(n7838), .ZN(n11156) );
  OAI211_X1 U9148 ( .C1(n7840), .C2(n11053), .A(n11126), .B(n7839), .ZN(n11052) );
  AOI22_X1 U9149 ( .A1(n11011), .A2(P1_REG2_REG_6__SCAN_IN), .B1(n7841), .B2(
        n11149), .ZN(n7844) );
  NAND2_X1 U9150 ( .A1(n11151), .A2(n7842), .ZN(n7843) );
  OAI211_X1 U9151 ( .C1(n11052), .C2(n11153), .A(n7844), .B(n7843), .ZN(n7845)
         );
  AOI21_X1 U9152 ( .B1(n11056), .B2(n11156), .A(n7845), .ZN(n7846) );
  OAI21_X1 U9153 ( .B1(n7847), .B2(n11011), .A(n7846), .ZN(P1_U3287) );
  INV_X1 U9154 ( .A(n7848), .ZN(n7849) );
  AOI21_X1 U9155 ( .B1(n7851), .B2(n7850), .A(n7849), .ZN(n7913) );
  INV_X1 U9156 ( .A(n7851), .ZN(n8456) );
  XNOR2_X1 U9157 ( .A(n7852), .B(n8456), .ZN(n7853) );
  OAI222_X1 U9158 ( .A1(n9476), .A2(n8117), .B1(n9474), .B2(n7936), .C1(n9471), 
        .C2(n7853), .ZN(n7910) );
  AOI21_X1 U9159 ( .B1(n7913), .B2(n9541), .A(n7910), .ZN(n7858) );
  INV_X1 U9160 ( .A(n7932), .ZN(n7942) );
  INV_X1 U9161 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n7854) );
  OAI22_X1 U9162 ( .A1(n7942), .A2(n9607), .B1(n11178), .B2(n7854), .ZN(n7855)
         );
  INV_X1 U9163 ( .A(n7855), .ZN(n7856) );
  OAI21_X1 U9164 ( .B1(n7858), .B2(n6432), .A(n7856), .ZN(P2_U3417) );
  AOI22_X1 U9165 ( .A1(n7932), .A2(n8024), .B1(n9572), .B2(
        P2_REG1_REG_9__SCAN_IN), .ZN(n7857) );
  OAI21_X1 U9166 ( .B1(n7858), .B2(n9572), .A(n7857), .ZN(P2_U3468) );
  INV_X1 U9167 ( .A(n8853), .ZN(n7859) );
  NAND3_X1 U9168 ( .A1(n7860), .A2(n7859), .A3(n8935), .ZN(n7861) );
  NAND2_X1 U9169 ( .A1(n7861), .A2(n8855), .ZN(n7862) );
  XNOR2_X1 U9170 ( .A(n7862), .B(n7867), .ZN(n7863) );
  NAND2_X1 U9171 ( .A1(n7863), .A2(n10566), .ZN(n7865) );
  NAND2_X1 U9172 ( .A1(n10291), .A2(n10999), .ZN(n7864) );
  NAND2_X1 U9173 ( .A1(n7865), .A2(n7864), .ZN(n11070) );
  INV_X1 U9174 ( .A(n11070), .ZN(n7875) );
  OAI21_X1 U9175 ( .B1(n7868), .B2(n7867), .A(n7866), .ZN(n11072) );
  XNOR2_X1 U9176 ( .A(n7869), .B(n10172), .ZN(n7870) );
  AOI22_X1 U9177 ( .A1(n7870), .A2(n11126), .B1(n11002), .B2(n10289), .ZN(
        n11068) );
  AOI22_X1 U9178 ( .A1(n11011), .A2(P1_REG2_REG_9__SCAN_IN), .B1(n10166), .B2(
        n11149), .ZN(n7872) );
  NAND2_X1 U9179 ( .A1(n10172), .A2(n11151), .ZN(n7871) );
  OAI211_X1 U9180 ( .C1(n11068), .C2(n11153), .A(n7872), .B(n7871), .ZN(n7873)
         );
  AOI21_X1 U9181 ( .B1(n11072), .B2(n10575), .A(n7873), .ZN(n7874) );
  OAI21_X1 U9182 ( .B1(n7875), .B2(n11011), .A(n7874), .ZN(P1_U3284) );
  NAND2_X1 U9183 ( .A1(n7876), .A2(n8864), .ZN(n7878) );
  INV_X1 U9184 ( .A(n8944), .ZN(n7877) );
  XNOR2_X1 U9185 ( .A(n7878), .B(n7877), .ZN(n7880) );
  OAI22_X1 U9186 ( .A1(n10119), .A2(n11137), .B1(n11138), .B2(n11135), .ZN(
        n7879) );
  AOI21_X1 U9187 ( .B1(n7880), .B2(n10566), .A(n7879), .ZN(n11095) );
  XOR2_X1 U9188 ( .A(n7881), .B(n8944), .Z(n11098) );
  NAND2_X1 U9189 ( .A1(n11098), .A2(n10575), .ZN(n7888) );
  INV_X1 U9190 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n7882) );
  OAI22_X1 U9191 ( .A1(n10560), .A2(n7882), .B1(n10116), .B2(n10580), .ZN(
        n7886) );
  INV_X1 U9192 ( .A(n8670), .ZN(n11096) );
  INV_X1 U9193 ( .A(n7898), .ZN(n7884) );
  INV_X1 U9194 ( .A(n7883), .ZN(n7921) );
  OAI211_X1 U9195 ( .C1(n11096), .C2(n7884), .A(n7921), .B(n11126), .ZN(n11094) );
  NOR2_X1 U9196 ( .A1(n11094), .A2(n11153), .ZN(n7885) );
  AOI211_X1 U9197 ( .C1(n11151), .C2(n8670), .A(n7886), .B(n7885), .ZN(n7887)
         );
  OAI211_X1 U9198 ( .C1(n11011), .C2(n11095), .A(n7888), .B(n7887), .ZN(
        P1_U3281) );
  INV_X1 U9199 ( .A(n8945), .ZN(n7889) );
  XNOR2_X1 U9200 ( .A(n7890), .B(n7889), .ZN(n11089) );
  NAND2_X1 U9201 ( .A1(n11089), .A2(n11141), .ZN(n7896) );
  NAND2_X1 U9202 ( .A1(n7891), .A2(n8862), .ZN(n7892) );
  XNOR2_X1 U9203 ( .A(n7892), .B(n8945), .ZN(n7894) );
  OAI22_X1 U9204 ( .A1(n8654), .A2(n11137), .B1(n10213), .B2(n11135), .ZN(
        n7893) );
  AOI21_X1 U9205 ( .B1(n7894), .B2(n10566), .A(n7893), .ZN(n7895) );
  AOI21_X1 U9206 ( .B1(n7897), .B2(n8663), .A(n10577), .ZN(n7899) );
  NAND2_X1 U9207 ( .A1(n7899), .A2(n7898), .ZN(n11086) );
  INV_X1 U9208 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n7900) );
  OAI22_X1 U9209 ( .A1(n10560), .A2(n7900), .B1(n10214), .B2(n10580), .ZN(
        n7901) );
  AOI21_X1 U9210 ( .B1(n8663), .B2(n11151), .A(n7901), .ZN(n7902) );
  OAI21_X1 U9211 ( .B1(n11086), .B2(n11153), .A(n7902), .ZN(n7903) );
  AOI21_X1 U9212 ( .B1(n11089), .B2(n11156), .A(n7903), .ZN(n7904) );
  OAI21_X1 U9213 ( .B1(n11091), .B2(n11011), .A(n7904), .ZN(P1_U3282) );
  INV_X1 U9214 ( .A(n7905), .ZN(n7909) );
  OAI222_X1 U9215 ( .A1(n9109), .A2(n7909), .B1(n8624), .B2(P2_U3151), .C1(
        n7906), .C2(n9614), .ZN(P2_U3275) );
  INV_X1 U9216 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n7907) );
  OAI222_X1 U9217 ( .A1(P1_U3086), .A2(n5277), .B1(n10704), .B2(n9108), .C1(
        n7907), .C2(n10701), .ZN(P1_U3334) );
  INV_X1 U9218 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n7908) );
  OAI222_X1 U9219 ( .A1(P1_U3086), .A2(n6813), .B1(n10704), .B2(n7909), .C1(
        n7908), .C2(n10701), .ZN(P1_U3335) );
  OAI22_X1 U9220 ( .A1(n7942), .A2(n9441), .B1(n7937), .B2(n11104), .ZN(n7912)
         );
  MUX2_X1 U9221 ( .A(P2_REG2_REG_9__SCAN_IN), .B(n7910), .S(n11111), .Z(n7911)
         );
  AOI211_X1 U9222 ( .C1(n9443), .C2(n7913), .A(n7912), .B(n7911), .ZN(n7914)
         );
  INV_X1 U9223 ( .A(n7914), .ZN(P2_U3224) );
  XNOR2_X1 U9224 ( .A(n7915), .B(n8946), .ZN(n8016) );
  INV_X1 U9225 ( .A(n8016), .ZN(n7927) );
  NAND3_X1 U9226 ( .A1(n5601), .A2(n7916), .A3(n8874), .ZN(n7917) );
  AOI21_X1 U9227 ( .B1(n11129), .B2(n7917), .A(n11132), .ZN(n7919) );
  OAI22_X1 U9228 ( .A1(n10213), .A2(n11137), .B1(n10190), .B2(n11135), .ZN(
        n7918) );
  OR2_X1 U9229 ( .A1(n7919), .A2(n7918), .ZN(n8014) );
  INV_X1 U9230 ( .A(n11124), .ZN(n7920) );
  AOI211_X1 U9231 ( .C1(n8680), .C2(n7921), .A(n10577), .B(n7920), .ZN(n8015)
         );
  NAND2_X1 U9232 ( .A1(n8015), .A2(n11018), .ZN(n7924) );
  INV_X1 U9233 ( .A(n7922), .ZN(n10192) );
  AOI22_X1 U9234 ( .A1(n11011), .A2(P1_REG2_REG_13__SCAN_IN), .B1(n10192), 
        .B2(n11149), .ZN(n7923) );
  OAI211_X1 U9235 ( .C1(n11116), .C2(n11014), .A(n7924), .B(n7923), .ZN(n7925)
         );
  AOI21_X1 U9236 ( .B1(n10560), .B2(n8014), .A(n7925), .ZN(n7926) );
  OAI21_X1 U9237 ( .B1(n7927), .B2(n10563), .A(n7926), .ZN(P1_U3280) );
  NAND2_X1 U9238 ( .A1(n7928), .A2(n9253), .ZN(n7930) );
  INV_X1 U9239 ( .A(n7928), .ZN(n7929) );
  XNOR2_X1 U9240 ( .A(n7932), .B(n6905), .ZN(n8046) );
  XNOR2_X1 U9241 ( .A(n8046), .B(n9252), .ZN(n7933) );
  OAI211_X1 U9242 ( .C1(n7934), .C2(n7933), .A(n8048), .B(n9158), .ZN(n7941)
         );
  OAI21_X1 U9243 ( .B1(n9125), .B2(n7936), .A(n7935), .ZN(n7939) );
  NOR2_X1 U9244 ( .A1(n9217), .A2(n7937), .ZN(n7938) );
  AOI211_X1 U9245 ( .C1(n9214), .C2(n9251), .A(n7939), .B(n7938), .ZN(n7940)
         );
  OAI211_X1 U9246 ( .C1(n7942), .C2(n9238), .A(n7941), .B(n7940), .ZN(P2_U3171) );
  INV_X1 U9247 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n7948) );
  NOR2_X1 U9248 ( .A1(n7943), .A2(n9567), .ZN(n7945) );
  AOI211_X1 U9249 ( .C1(n9553), .C2(n7946), .A(n7945), .B(n7944), .ZN(n11067)
         );
  OR2_X1 U9250 ( .A1(n11067), .A2(n9572), .ZN(n7947) );
  OAI21_X1 U9251 ( .B1(n9561), .B2(n7948), .A(n7947), .ZN(P2_U3467) );
  NAND2_X1 U9252 ( .A1(n7950), .A2(n7949), .ZN(n7964) );
  NAND2_X1 U9253 ( .A1(n7964), .A2(n7961), .ZN(n7951) );
  NAND2_X1 U9254 ( .A1(n7951), .A2(n7962), .ZN(n7952) );
  XNOR2_X1 U9255 ( .A(n7952), .B(n8443), .ZN(n7953) );
  OAI222_X1 U9256 ( .A1(n9476), .A2(n8174), .B1(n9474), .B2(n8117), .C1(n9471), 
        .C2(n7953), .ZN(n8010) );
  INV_X1 U9257 ( .A(n8010), .ZN(n7960) );
  OAI21_X1 U9258 ( .B1(n7955), .B2(n8443), .A(n7954), .ZN(n8012) );
  INV_X1 U9259 ( .A(n8122), .ZN(n8009) );
  NOR2_X1 U9260 ( .A1(n8009), .A2(n9441), .ZN(n7958) );
  OAI22_X1 U9261 ( .A1(n11111), .A2(n7956), .B1(n8120), .B2(n11104), .ZN(n7957) );
  AOI211_X1 U9262 ( .C1(n8012), .C2(n9443), .A(n7958), .B(n7957), .ZN(n7959)
         );
  OAI21_X1 U9263 ( .B1(n7960), .B2(n9488), .A(n7959), .ZN(P2_U3222) );
  NAND2_X1 U9264 ( .A1(n7962), .A2(n7961), .ZN(n8454) );
  XNOR2_X1 U9265 ( .A(n7963), .B(n8454), .ZN(n8058) );
  INV_X1 U9266 ( .A(n8058), .ZN(n7969) );
  XOR2_X1 U9267 ( .A(n8454), .B(n7964), .Z(n7966) );
  OAI22_X1 U9268 ( .A1(n8050), .A2(n9474), .B1(n8003), .B2(n9476), .ZN(n7965)
         );
  AOI21_X1 U9269 ( .B1(n7966), .B2(n9490), .A(n7965), .ZN(n7967) );
  OAI21_X1 U9270 ( .B1(n7968), .B2(n8058), .A(n7967), .ZN(n8059) );
  AOI21_X1 U9271 ( .B1(n7970), .B2(n7969), .A(n8059), .ZN(n7973) );
  OAI22_X1 U9272 ( .A1(n9500), .A2(n7743), .B1(n8053), .B2(n11104), .ZN(n7971)
         );
  AOI21_X1 U9273 ( .B1(n8061), .B2(n9509), .A(n7971), .ZN(n7972) );
  OAI21_X1 U9274 ( .B1(n7973), .B2(n9488), .A(n7972), .ZN(P2_U3223) );
  OAI222_X1 U9275 ( .A1(n9109), .A2(n7997), .B1(n7975), .B2(P2_U3151), .C1(
        n7974), .C2(n9614), .ZN(P2_U3273) );
  NAND2_X1 U9276 ( .A1(P2_REG2_REG_10__SCAN_IN), .A2(n7989), .ZN(n7976) );
  NAND2_X1 U9277 ( .A1(P2_REG2_REG_11__SCAN_IN), .A2(n7978), .ZN(n8093) );
  OAI21_X1 U9278 ( .B1(P2_REG2_REG_11__SCAN_IN), .B2(n7978), .A(n8093), .ZN(
        n7979) );
  INV_X1 U9279 ( .A(n7979), .ZN(n7996) );
  INV_X1 U9280 ( .A(n7980), .ZN(n7981) );
  OAI21_X1 U9281 ( .B1(n7983), .B2(n7982), .A(n7981), .ZN(n7985) );
  MUX2_X1 U9282 ( .A(P2_REG2_REG_11__SCAN_IN), .B(P2_REG1_REG_11__SCAN_IN), 
        .S(n9324), .Z(n8082) );
  XNOR2_X1 U9283 ( .A(n8082), .B(n8078), .ZN(n7984) );
  NAND2_X1 U9284 ( .A1(n7984), .A2(n7985), .ZN(n8083) );
  OAI21_X1 U9285 ( .B1(n7985), .B2(n7984), .A(n8083), .ZN(n7986) );
  NAND2_X1 U9286 ( .A1(n7986), .A2(n10962), .ZN(n7995) );
  INV_X1 U9287 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n7987) );
  NAND2_X1 U9288 ( .A1(P2_U3151), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n8116) );
  OAI21_X1 U9289 ( .B1(n10938), .B2(n7987), .A(n8116), .ZN(n7993) );
  AOI21_X2 U9290 ( .B1(P2_REG1_REG_10__SCAN_IN), .B2(n7989), .A(n7988), .ZN(
        n8077) );
  AOI21_X1 U9291 ( .B1(n7990), .B2(n6081), .A(n8079), .ZN(n7991) );
  NOR2_X1 U9292 ( .A1(n10969), .A2(n7991), .ZN(n7992) );
  AOI211_X1 U9293 ( .C1(n10941), .C2(n8078), .A(n7993), .B(n7992), .ZN(n7994)
         );
  OAI211_X1 U9294 ( .C1(n10974), .C2(n7996), .A(n7995), .B(n7994), .ZN(
        P2_U3193) );
  INV_X1 U9295 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n7998) );
  OAI222_X1 U9296 ( .A1(n10701), .A2(n7998), .B1(P1_U3086), .B2(n9062), .C1(
        n7997), .C2(n10704), .ZN(P1_U3333) );
  AND2_X1 U9297 ( .A1(n8195), .A2(n8196), .ZN(n8554) );
  XNOR2_X1 U9298 ( .A(n7999), .B(n8457), .ZN(n8022) );
  INV_X1 U9299 ( .A(n8022), .ZN(n8008) );
  AND2_X1 U9300 ( .A1(n8169), .A2(n8000), .ZN(n8001) );
  XNOR2_X1 U9301 ( .A(n8001), .B(n8457), .ZN(n8002) );
  OAI222_X1 U9302 ( .A1(n9474), .A2(n8003), .B1(n9476), .B2(n9126), .C1(n8002), 
        .C2(n9471), .ZN(n8021) );
  NAND2_X1 U9303 ( .A1(n8021), .A2(n9500), .ZN(n8007) );
  OAI22_X1 U9304 ( .A1(n9500), .A2(n8004), .B1(n8201), .B2(n11104), .ZN(n8005)
         );
  AOI21_X1 U9305 ( .B1(n8203), .B2(n9509), .A(n8005), .ZN(n8006) );
  OAI211_X1 U9306 ( .C1(n8008), .C2(n9505), .A(n8007), .B(n8006), .ZN(P2_U3221) );
  NOR2_X1 U9307 ( .A1(n8009), .A2(n9565), .ZN(n8011) );
  AOI211_X1 U9308 ( .C1(n9541), .C2(n8012), .A(n8011), .B(n8010), .ZN(n11085)
         );
  OR2_X1 U9309 ( .A1(n11085), .A2(n9572), .ZN(n8013) );
  OAI21_X1 U9310 ( .B1(n9561), .B2(n6081), .A(n8013), .ZN(P2_U3470) );
  INV_X1 U9311 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n8017) );
  AOI211_X1 U9312 ( .C1(n8016), .C2(n11168), .A(n8015), .B(n8014), .ZN(n8019)
         );
  MUX2_X1 U9313 ( .A(n8017), .B(n8019), .S(n11175), .Z(n8018) );
  OAI21_X1 U9314 ( .B1(n11116), .B2(n10685), .A(n8018), .ZN(P1_U3492) );
  INV_X1 U9315 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n10370) );
  MUX2_X1 U9316 ( .A(n10370), .B(n8019), .S(n11171), .Z(n8020) );
  OAI21_X1 U9317 ( .B1(n11116), .B2(n10644), .A(n8020), .ZN(P1_U3535) );
  AOI21_X1 U9318 ( .B1(n9541), .B2(n8022), .A(n8021), .ZN(n8029) );
  NOR2_X1 U9319 ( .A1(n9561), .A2(n6101), .ZN(n8023) );
  AOI21_X1 U9320 ( .B1(n8203), .B2(n8024), .A(n8023), .ZN(n8025) );
  OAI21_X1 U9321 ( .B1(n8029), .B2(n9572), .A(n8025), .ZN(P2_U3471) );
  INV_X1 U9322 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n8026) );
  NOR2_X1 U9323 ( .A1(n11178), .A2(n8026), .ZN(n8027) );
  AOI21_X1 U9324 ( .B1(n8203), .B2(n6436), .A(n8027), .ZN(n8028) );
  OAI21_X1 U9325 ( .B1(n8029), .B2(n6432), .A(n8028), .ZN(P2_U3426) );
  INV_X1 U9326 ( .A(n8032), .ZN(n8031) );
  NOR2_X1 U9327 ( .A1(n9061), .A2(P1_U3086), .ZN(n9057) );
  AOI21_X1 U9328 ( .B1(P2_DATAO_REG_23__SCAN_IN), .B2(n10695), .A(n9057), .ZN(
        n8030) );
  OAI21_X1 U9329 ( .B1(n8031), .B2(n10704), .A(n8030), .ZN(P1_U3332) );
  NAND2_X1 U9330 ( .A1(n8032), .A2(n9622), .ZN(n8034) );
  NAND2_X1 U9331 ( .A1(n8033), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8632) );
  OAI211_X1 U9332 ( .C1(n8035), .C2(n9614), .A(n8034), .B(n8632), .ZN(P2_U3272) );
  NAND2_X1 U9333 ( .A1(n8036), .A2(n8553), .ZN(n8038) );
  NAND2_X1 U9334 ( .A1(n8038), .A2(n8037), .ZN(n8039) );
  XNOR2_X1 U9335 ( .A(n8039), .B(n6366), .ZN(n8285) );
  XNOR2_X1 U9336 ( .A(n8040), .B(n8479), .ZN(n8041) );
  OAI222_X1 U9337 ( .A1(n9474), .A2(n9126), .B1(n9476), .B2(n8478), .C1(n8041), 
        .C2(n9471), .ZN(n8286) );
  INV_X1 U9338 ( .A(n9129), .ZN(n8042) );
  NOR2_X1 U9339 ( .A1(n8042), .A2(n11105), .ZN(n8043) );
  OAI21_X1 U9340 ( .B1(n8286), .B2(n8043), .A(n9500), .ZN(n8045) );
  AOI22_X1 U9341 ( .A1(n9488), .A2(P2_REG2_REG_14__SCAN_IN), .B1(n9439), .B2(
        n9128), .ZN(n8044) );
  OAI211_X1 U9342 ( .C1(n8285), .C2(n9505), .A(n8045), .B(n8044), .ZN(P2_U3219) );
  OR2_X1 U9343 ( .A1(n8046), .A2(n8050), .ZN(n8047) );
  XNOR2_X1 U9344 ( .A(n8061), .B(n6905), .ZN(n8114) );
  XNOR2_X1 U9345 ( .A(n8115), .B(n9251), .ZN(n8056) );
  OAI21_X1 U9346 ( .B1(n9125), .B2(n8050), .A(n8049), .ZN(n8051) );
  AOI21_X1 U9347 ( .B1(n9214), .B2(n9250), .A(n8051), .ZN(n8052) );
  OAI21_X1 U9348 ( .B1(n8053), .B2(n9217), .A(n8052), .ZN(n8054) );
  AOI21_X1 U9349 ( .B1(n8061), .B2(n9219), .A(n8054), .ZN(n8055) );
  OAI21_X1 U9350 ( .B1(n8056), .B2(n9224), .A(n8055), .ZN(P2_U3157) );
  NOR2_X1 U9351 ( .A1(n8058), .A2(n8057), .ZN(n8060) );
  AOI211_X1 U9352 ( .C1(n9553), .C2(n8061), .A(n8060), .B(n8059), .ZN(n11083)
         );
  OR2_X1 U9353 ( .A1(n11083), .A2(n9572), .ZN(n8062) );
  OAI21_X1 U9354 ( .B1(n9561), .B2(n7742), .A(n8062), .ZN(P2_U3469) );
  NAND2_X1 U9355 ( .A1(n8063), .A2(n8948), .ZN(n8064) );
  NAND2_X1 U9356 ( .A1(n8065), .A2(n8064), .ZN(n8067) );
  OAI22_X1 U9357 ( .A1(n10190), .A2(n11137), .B1(n10258), .B2(n11135), .ZN(
        n8066) );
  AOI21_X1 U9358 ( .B1(n8067), .B2(n10566), .A(n8066), .ZN(n11164) );
  OAI21_X1 U9359 ( .B1(n8069), .B2(n8948), .A(n8068), .ZN(n8070) );
  INV_X1 U9360 ( .A(n8070), .ZN(n11169) );
  NAND2_X1 U9361 ( .A1(n11169), .A2(n10575), .ZN(n8076) );
  INV_X1 U9362 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n8071) );
  OAI22_X1 U9363 ( .A1(n10560), .A2(n8071), .B1(n10264), .B2(n10580), .ZN(
        n8074) );
  INV_X1 U9364 ( .A(n11127), .ZN(n8072) );
  OAI211_X1 U9365 ( .C1(n11166), .C2(n8072), .A(n11126), .B(n8218), .ZN(n11163) );
  NOR2_X1 U9366 ( .A1(n11163), .A2(n11153), .ZN(n8073) );
  AOI211_X1 U9367 ( .C1(n11151), .C2(n10267), .A(n8074), .B(n8073), .ZN(n8075)
         );
  OAI211_X1 U9368 ( .C1(n11011), .C2(n11164), .A(n8076), .B(n8075), .ZN(
        P1_U3278) );
  NOR2_X1 U9369 ( .A1(n8078), .A2(n8077), .ZN(n8080) );
  NAND2_X1 U9370 ( .A1(P2_REG1_REG_12__SCAN_IN), .A2(n8153), .ZN(n8142) );
  OAI21_X1 U9371 ( .B1(P2_REG1_REG_12__SCAN_IN), .B2(n8153), .A(n8142), .ZN(
        n8081) );
  AOI21_X1 U9372 ( .B1(n5203), .B2(n8081), .A(n8144), .ZN(n8101) );
  INV_X1 U9373 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n8090) );
  MUX2_X1 U9374 ( .A(P2_REG2_REG_12__SCAN_IN), .B(P2_REG1_REG_12__SCAN_IN), 
        .S(n9324), .Z(n8146) );
  XNOR2_X1 U9375 ( .A(n8146), .B(n8099), .ZN(n8086) );
  OR2_X1 U9376 ( .A1(n8082), .A2(n8092), .ZN(n8084) );
  NAND2_X1 U9377 ( .A1(n8084), .A2(n8083), .ZN(n8085) );
  NAND2_X1 U9378 ( .A1(n8086), .A2(n8085), .ZN(n8147) );
  OAI21_X1 U9379 ( .B1(n8086), .B2(n8085), .A(n8147), .ZN(n8088) );
  INV_X1 U9380 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n8087) );
  NOR2_X1 U9381 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8087), .ZN(n8199) );
  AOI21_X1 U9382 ( .B1(n8088), .B2(n10962), .A(n8199), .ZN(n8089) );
  OAI21_X1 U9383 ( .B1(n10938), .B2(n8090), .A(n8089), .ZN(n8098) );
  NAND2_X1 U9384 ( .A1(n8092), .A2(n8091), .ZN(n8094) );
  NAND2_X1 U9385 ( .A1(n8099), .A2(n8004), .ZN(n8152) );
  OAI21_X1 U9386 ( .B1(n8099), .B2(n8004), .A(n8152), .ZN(n8095) );
  XNOR2_X1 U9387 ( .A(n8151), .B(n8095), .ZN(n8096) );
  NOR2_X1 U9388 ( .A1(n8096), .A2(n10974), .ZN(n8097) );
  AOI211_X1 U9389 ( .C1(n10941), .C2(n8099), .A(n8098), .B(n8097), .ZN(n8100)
         );
  OAI21_X1 U9390 ( .B1(n8101), .B2(n10969), .A(n8100), .ZN(P2_U3194) );
  XNOR2_X1 U9391 ( .A(n8102), .B(n8106), .ZN(n8103) );
  AOI222_X1 U9392 ( .A1(n9490), .A2(n8103), .B1(n9247), .B2(n9492), .C1(n9245), 
        .C2(n9495), .ZN(n8136) );
  INV_X1 U9393 ( .A(n8136), .ZN(n8104) );
  AOI21_X1 U9394 ( .B1(n9439), .B2(n9235), .A(n8104), .ZN(n8111) );
  NAND2_X1 U9395 ( .A1(n8128), .A2(n8105), .ZN(n8107) );
  XNOR2_X1 U9396 ( .A(n8107), .B(n8106), .ZN(n8138) );
  INV_X1 U9397 ( .A(n8477), .ZN(n9239) );
  OAI22_X1 U9398 ( .A1(n9239), .A2(n9441), .B1(n9500), .B2(n8108), .ZN(n8109)
         );
  AOI21_X1 U9399 ( .B1(n8138), .B2(n9443), .A(n8109), .ZN(n8110) );
  OAI21_X1 U9400 ( .B1(n8111), .B2(n9488), .A(n8110), .ZN(P2_U3218) );
  INV_X1 U9401 ( .A(n8112), .ZN(n8113) );
  XNOR2_X1 U9402 ( .A(n8122), .B(n6905), .ZN(n8191) );
  XOR2_X1 U9403 ( .A(n9250), .B(n8191), .Z(n8193) );
  XOR2_X1 U9404 ( .A(n8194), .B(n8193), .Z(n8124) );
  OAI21_X1 U9405 ( .B1(n9125), .B2(n8117), .A(n8116), .ZN(n8118) );
  AOI21_X1 U9406 ( .B1(n9214), .B2(n9249), .A(n8118), .ZN(n8119) );
  OAI21_X1 U9407 ( .B1(n8120), .B2(n9217), .A(n8119), .ZN(n8121) );
  AOI21_X1 U9408 ( .B1(n8122), .B2(n9219), .A(n8121), .ZN(n8123) );
  OAI21_X1 U9409 ( .B1(n8124), .B2(n9224), .A(n8123), .ZN(P2_U3176) );
  XNOR2_X1 U9410 ( .A(n8125), .B(n8483), .ZN(n8126) );
  OAI222_X1 U9411 ( .A1(n9474), .A2(n8478), .B1(n9476), .B2(n9164), .C1(n8126), 
        .C2(n9471), .ZN(n8229) );
  AOI21_X1 U9412 ( .B1(n9439), .B2(n9166), .A(n8229), .ZN(n8133) );
  NAND2_X1 U9413 ( .A1(n8128), .A2(n8127), .ZN(n8129) );
  AND2_X1 U9414 ( .A1(n8129), .A2(n6165), .ZN(n8130) );
  AOI21_X1 U9415 ( .B1(n8483), .B2(n8130), .A(n5206), .ZN(n8231) );
  INV_X1 U9416 ( .A(n8387), .ZN(n9169) );
  OAI22_X1 U9417 ( .A1(n9169), .A2(n9441), .B1(n9301), .B2(n9500), .ZN(n8131)
         );
  AOI21_X1 U9418 ( .B1(n8231), .B2(n9443), .A(n8131), .ZN(n8132) );
  OAI21_X1 U9419 ( .B1(n8133), .B2(n9488), .A(n8132), .ZN(P2_U3217) );
  OAI222_X1 U9420 ( .A1(n9619), .A2(n8163), .B1(P2_U3151), .B2(n8135), .C1(
        n8134), .C2(n9614), .ZN(P2_U3270) );
  OAI21_X1 U9421 ( .B1(n9239), .B2(n9565), .A(n8136), .ZN(n8137) );
  AOI21_X1 U9422 ( .B1(n8138), .B2(n9541), .A(n8137), .ZN(n11162) );
  NAND2_X1 U9423 ( .A1(n9572), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n8139) );
  OAI21_X1 U9424 ( .B1(n11162), .B2(n9572), .A(n8139), .ZN(P2_U3474) );
  INV_X1 U9425 ( .A(n8140), .ZN(n8166) );
  OAI222_X1 U9426 ( .A1(n9619), .A2(n8166), .B1(P2_U3151), .B2(n6406), .C1(
        n8141), .C2(n9614), .ZN(P2_U3271) );
  INV_X1 U9427 ( .A(n8142), .ZN(n8143) );
  AOI21_X1 U9428 ( .B1(n6117), .B2(n8145), .A(n8258), .ZN(n8161) );
  MUX2_X1 U9429 ( .A(P2_REG2_REG_13__SCAN_IN), .B(P2_REG1_REG_13__SCAN_IN), 
        .S(n9324), .Z(n8262) );
  XNOR2_X1 U9430 ( .A(n8262), .B(n8270), .ZN(n8150) );
  OR2_X1 U9431 ( .A1(n8146), .A2(n8153), .ZN(n8148) );
  NAND2_X1 U9432 ( .A1(n8148), .A2(n8147), .ZN(n8149) );
  NAND2_X1 U9433 ( .A1(n8150), .A2(n8149), .ZN(n8261) );
  OAI21_X1 U9434 ( .B1(n8150), .B2(n8149), .A(n8261), .ZN(n8158) );
  NOR2_X1 U9435 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9915), .ZN(n8240) );
  XNOR2_X1 U9436 ( .A(n8270), .B(n8269), .ZN(n8154) );
  AOI21_X1 U9437 ( .B1(n8154), .B2(n6120), .A(n8271), .ZN(n8156) );
  INV_X1 U9438 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n8155) );
  OAI22_X1 U9439 ( .A1(n10974), .A2(n8156), .B1(n10938), .B2(n8155), .ZN(n8157) );
  AOI211_X1 U9440 ( .C1(n10962), .C2(n8158), .A(n8240), .B(n8157), .ZN(n8160)
         );
  NAND2_X1 U9441 ( .A1(n10941), .A2(n8270), .ZN(n8159) );
  OAI211_X1 U9442 ( .C1(n8161), .C2(n10969), .A(n8160), .B(n8159), .ZN(
        P2_U3195) );
  INV_X1 U9443 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n8162) );
  OAI222_X1 U9444 ( .A1(P1_U3086), .A2(n8164), .B1(n10704), .B2(n8163), .C1(
        n8162), .C2(n10701), .ZN(P1_U3330) );
  INV_X1 U9445 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n8165) );
  OAI222_X1 U9446 ( .A1(P1_U3086), .A2(n8167), .B1(n10704), .B2(n8166), .C1(
        n8165), .C2(n10701), .ZN(P1_U3331) );
  INV_X1 U9447 ( .A(n8553), .ZN(n8460) );
  XNOR2_X1 U9448 ( .A(n8036), .B(n8460), .ZN(n11102) );
  NOR2_X1 U9449 ( .A1(n11102), .A2(n9567), .ZN(n8175) );
  AND2_X1 U9450 ( .A1(n8169), .A2(n8168), .ZN(n8171) );
  NOR2_X1 U9451 ( .A1(n8171), .A2(n8170), .ZN(n8172) );
  XNOR2_X1 U9452 ( .A(n8172), .B(n8460), .ZN(n8173) );
  OAI222_X1 U9453 ( .A1(n9474), .A2(n8174), .B1(n9476), .B2(n8381), .C1(n9471), 
        .C2(n8173), .ZN(n11107) );
  AOI211_X1 U9454 ( .C1(n9553), .C2(n11103), .A(n8175), .B(n11107), .ZN(n11114) );
  NAND2_X1 U9455 ( .A1(n9572), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n8176) );
  OAI21_X1 U9456 ( .B1(n11114), .B2(n9572), .A(n8176), .ZN(P2_U3472) );
  XNOR2_X1 U9457 ( .A(n8177), .B(n8952), .ZN(n10641) );
  INV_X1 U9458 ( .A(n10641), .ZN(n8190) );
  NAND2_X1 U9459 ( .A1(n8179), .A2(n8178), .ZN(n8180) );
  NAND3_X1 U9460 ( .A1(n8248), .A2(n10566), .A3(n8180), .ZN(n8183) );
  OAI22_X1 U9461 ( .A1(n10569), .A2(n11135), .B1(n10258), .B2(n11137), .ZN(
        n8181) );
  INV_X1 U9462 ( .A(n8181), .ZN(n8182) );
  NAND2_X1 U9463 ( .A1(n8183), .A2(n8182), .ZN(n10639) );
  INV_X1 U9464 ( .A(n8217), .ZN(n8185) );
  INV_X1 U9465 ( .A(n8251), .ZN(n8184) );
  AOI211_X1 U9466 ( .C1(n8722), .C2(n8185), .A(n10577), .B(n8184), .ZN(n10640)
         );
  NAND2_X1 U9467 ( .A1(n10640), .A2(n11018), .ZN(n8187) );
  AOI22_X1 U9468 ( .A1(n11011), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n10149), 
        .B2(n11149), .ZN(n8186) );
  OAI211_X1 U9469 ( .C1(n10686), .C2(n11014), .A(n8187), .B(n8186), .ZN(n8188)
         );
  AOI21_X1 U9470 ( .B1(n10560), .B2(n10639), .A(n8188), .ZN(n8189) );
  OAI21_X1 U9471 ( .B1(n8190), .B2(n10563), .A(n8189), .ZN(P1_U3276) );
  INV_X1 U9472 ( .A(n8191), .ZN(n8192) );
  OAI22_X1 U9473 ( .A1(n8194), .A2(n8193), .B1(n8192), .B2(n9250), .ZN(n8234)
         );
  MUX2_X1 U9474 ( .A(n8195), .B(n8551), .S(n6905), .Z(n8235) );
  MUX2_X1 U9475 ( .A(n8196), .B(n8550), .S(n6905), .Z(n8233) );
  NAND2_X1 U9476 ( .A1(n8235), .A2(n8233), .ZN(n8197) );
  XNOR2_X1 U9477 ( .A(n8234), .B(n8197), .ZN(n8205) );
  NOR2_X1 U9478 ( .A1(n9231), .A2(n9126), .ZN(n8198) );
  AOI211_X1 U9479 ( .C1(n9229), .C2(n9250), .A(n8199), .B(n8198), .ZN(n8200)
         );
  OAI21_X1 U9480 ( .B1(n8201), .B2(n9217), .A(n8200), .ZN(n8202) );
  AOI21_X1 U9481 ( .B1(n8203), .B2(n9219), .A(n8202), .ZN(n8204) );
  OAI21_X1 U9482 ( .B1(n8205), .B2(n9224), .A(n8204), .ZN(P2_U3164) );
  INV_X1 U9483 ( .A(n8206), .ZN(n8207) );
  AOI21_X1 U9484 ( .B1(n8462), .B2(n8208), .A(n8207), .ZN(n9568) );
  XNOR2_X1 U9485 ( .A(n8209), .B(n8462), .ZN(n8210) );
  OAI222_X1 U9486 ( .A1(n9474), .A2(n9232), .B1(n9476), .B2(n9475), .C1(n9471), 
        .C2(n8210), .ZN(n9569) );
  NAND2_X1 U9487 ( .A1(n9569), .A2(n9500), .ZN(n8214) );
  INV_X1 U9488 ( .A(n9174), .ZN(n8211) );
  OAI22_X1 U9489 ( .A1(n9500), .A2(n9318), .B1(n8211), .B2(n11104), .ZN(n8212)
         );
  AOI21_X1 U9490 ( .B1(n9178), .B2(n9509), .A(n8212), .ZN(n8213) );
  OAI211_X1 U9491 ( .C1(n9568), .C2(n9505), .A(n8214), .B(n8213), .ZN(P2_U3216) );
  OAI21_X1 U9492 ( .B1(n8216), .B2(n8949), .A(n8215), .ZN(n10650) );
  AOI211_X1 U9493 ( .C1(n10646), .C2(n8218), .A(n10577), .B(n8217), .ZN(n10645) );
  AOI22_X1 U9494 ( .A1(n11011), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n11149), 
        .B2(n8219), .ZN(n8220) );
  OAI21_X1 U9495 ( .B1(n8221), .B2(n11014), .A(n8220), .ZN(n8227) );
  OAI21_X1 U9496 ( .B1(n8224), .B2(n8223), .A(n8222), .ZN(n8225) );
  INV_X1 U9497 ( .A(n11136), .ZN(n10286) );
  AOI222_X1 U9498 ( .A1(n10566), .A2(n8225), .B1(n10286), .B2(n10999), .C1(
        n10284), .C2(n11002), .ZN(n10648) );
  NOR2_X1 U9499 ( .A1(n10648), .A2(n11011), .ZN(n8226) );
  AOI211_X1 U9500 ( .C1(n10645), .C2(n11018), .A(n8227), .B(n8226), .ZN(n8228)
         );
  OAI21_X1 U9501 ( .B1(n10650), .B2(n10563), .A(n8228), .ZN(P1_U3277) );
  NOR2_X1 U9502 ( .A1(n9169), .A2(n9565), .ZN(n8230) );
  AOI211_X1 U9503 ( .C1(n8231), .C2(n9541), .A(n8230), .B(n8229), .ZN(n11176)
         );
  OR2_X1 U9504 ( .A1(n11176), .A2(n9572), .ZN(n8232) );
  OAI21_X1 U9505 ( .B1(n9561), .B2(n6177), .A(n8232), .ZN(P2_U3475) );
  NAND2_X1 U9506 ( .A1(n8234), .A2(n8233), .ZN(n8236) );
  NAND2_X1 U9507 ( .A1(n8236), .A2(n8235), .ZN(n8378) );
  XNOR2_X1 U9508 ( .A(n11103), .B(n9098), .ZN(n8237) );
  NAND2_X1 U9509 ( .A1(n8237), .A2(n9248), .ZN(n9120) );
  NAND2_X1 U9510 ( .A1(n5215), .A2(n9120), .ZN(n8238) );
  XNOR2_X1 U9511 ( .A(n8378), .B(n8238), .ZN(n8244) );
  NOR2_X1 U9512 ( .A1(n9231), .A2(n8381), .ZN(n8239) );
  AOI211_X1 U9513 ( .C1(n9229), .C2(n9249), .A(n8240), .B(n8239), .ZN(n8241)
         );
  OAI21_X1 U9514 ( .B1(n5153), .B2(n9217), .A(n8241), .ZN(n8242) );
  AOI21_X1 U9515 ( .B1(n11103), .B2(n9219), .A(n8242), .ZN(n8243) );
  OAI21_X1 U9516 ( .B1(n8244), .B2(n9224), .A(n8243), .ZN(P2_U3174) );
  AOI21_X1 U9517 ( .B1(n8246), .B2(n8951), .A(n8245), .ZN(n8247) );
  INV_X1 U9518 ( .A(n8247), .ZN(n10638) );
  AOI21_X1 U9519 ( .B1(n9021), .B2(n8248), .A(n8951), .ZN(n8249) );
  NOR2_X1 U9520 ( .A1(n5199), .A2(n8249), .ZN(n8250) );
  OAI222_X1 U9521 ( .A1(n11135), .A2(n10550), .B1(n11137), .B2(n10237), .C1(
        n11132), .C2(n8250), .ZN(n10634) );
  INV_X1 U9522 ( .A(n10636), .ZN(n8254) );
  AOI211_X1 U9523 ( .C1(n10636), .C2(n8251), .A(n10577), .B(n5435), .ZN(n10635) );
  NAND2_X1 U9524 ( .A1(n10635), .A2(n11018), .ZN(n8253) );
  AOI22_X1 U9525 ( .A1(n11011), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n10231), 
        .B2(n11149), .ZN(n8252) );
  OAI211_X1 U9526 ( .C1(n8254), .C2(n11014), .A(n8253), .B(n8252), .ZN(n8255)
         );
  AOI21_X1 U9527 ( .B1(n10634), .B2(n10560), .A(n8255), .ZN(n8256) );
  OAI21_X1 U9528 ( .B1(n10638), .B2(n10563), .A(n8256), .ZN(P1_U3275) );
  NOR2_X1 U9529 ( .A1(n8270), .A2(n8257), .ZN(n8259) );
  AOI22_X1 U9530 ( .A1(n8277), .A2(P2_REG1_REG_14__SCAN_IN), .B1(n6142), .B2(
        n9269), .ZN(n8260) );
  AOI21_X1 U9531 ( .B1(n5201), .B2(n8260), .A(n9261), .ZN(n8279) );
  INV_X1 U9532 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n8268) );
  OAI21_X1 U9533 ( .B1(n8263), .B2(n8262), .A(n8261), .ZN(n8265) );
  MUX2_X1 U9534 ( .A(P2_REG2_REG_14__SCAN_IN), .B(P2_REG1_REG_14__SCAN_IN), 
        .S(n9324), .Z(n9263) );
  XNOR2_X1 U9535 ( .A(n8277), .B(n9263), .ZN(n8264) );
  NAND2_X1 U9536 ( .A1(n8264), .A2(n8265), .ZN(n9264) );
  OAI21_X1 U9537 ( .B1(n8265), .B2(n8264), .A(n9264), .ZN(n8266) );
  NAND2_X1 U9538 ( .A1(n8266), .A2(n10962), .ZN(n8267) );
  NAND2_X1 U9539 ( .A1(P2_U3151), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n9123) );
  OAI211_X1 U9540 ( .C1(n10938), .C2(n8268), .A(n8267), .B(n9123), .ZN(n8276)
         );
  MUX2_X1 U9541 ( .A(n6141), .B(P2_REG2_REG_14__SCAN_IN), .S(n8277), .Z(n8272)
         );
  INV_X1 U9542 ( .A(n8272), .ZN(n8273) );
  AOI21_X1 U9543 ( .B1(n5213), .B2(n8273), .A(n9268), .ZN(n8274) );
  NOR2_X1 U9544 ( .A1(n8274), .A2(n10974), .ZN(n8275) );
  AOI211_X1 U9545 ( .C1(n10941), .C2(n8277), .A(n8276), .B(n8275), .ZN(n8278)
         );
  OAI21_X1 U9546 ( .B1(n8279), .B2(n10969), .A(n8278), .ZN(P2_U3196) );
  INV_X1 U9547 ( .A(n8280), .ZN(n8283) );
  INV_X1 U9548 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n9732) );
  OAI222_X1 U9549 ( .A1(n8281), .A2(P1_U3086), .B1(n10704), .B2(n8283), .C1(
        n9732), .C2(n10701), .ZN(P1_U3329) );
  OAI222_X1 U9550 ( .A1(n9614), .A2(n8284), .B1(n9619), .B2(n8283), .C1(n8282), 
        .C2(P2_U3151), .ZN(P2_U3269) );
  NOR2_X1 U9551 ( .A1(n8285), .A2(n9567), .ZN(n8287) );
  AOI211_X1 U9552 ( .C1(n9553), .C2(n9129), .A(n8287), .B(n8286), .ZN(n11161)
         );
  OR2_X1 U9553 ( .A1(n11161), .A2(n9572), .ZN(n8288) );
  OAI21_X1 U9554 ( .B1(n9561), .B2(n6142), .A(n8288), .ZN(P2_U3473) );
  INV_X1 U9555 ( .A(n8289), .ZN(n8292) );
  OAI222_X1 U9556 ( .A1(n9619), .A2(n8292), .B1(n9324), .B2(P2_U3151), .C1(
        n8290), .C2(n9614), .ZN(P2_U3268) );
  INV_X1 U9557 ( .A(n8291), .ZN(n10792) );
  INV_X1 U9558 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n9942) );
  OAI222_X1 U9559 ( .A1(P1_U3086), .A2(n10792), .B1(n10704), .B2(n8292), .C1(
        n9942), .C2(n10701), .ZN(P1_U3328) );
  INV_X1 U9560 ( .A(n8293), .ZN(n10703) );
  OAI222_X1 U9561 ( .A1(n9619), .A2(n10703), .B1(n6347), .B2(P2_U3151), .C1(
        n8294), .C2(n9614), .ZN(P2_U3267) );
  NAND2_X1 U9562 ( .A1(n8295), .A2(SI_29_), .ZN(n8300) );
  INV_X1 U9563 ( .A(n8296), .ZN(n8298) );
  NAND2_X1 U9564 ( .A1(n8298), .A2(n8297), .ZN(n8299) );
  NAND2_X1 U9565 ( .A1(n8300), .A2(n8299), .ZN(n8316) );
  INV_X1 U9566 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n9933) );
  INV_X1 U9567 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n9071) );
  MUX2_X1 U9568 ( .A(n9933), .B(n9071), .S(n8306), .Z(n8302) );
  INV_X1 U9569 ( .A(SI_30_), .ZN(n8301) );
  NAND2_X1 U9570 ( .A1(n8302), .A2(n8301), .ZN(n8305) );
  INV_X1 U9571 ( .A(n8302), .ZN(n8303) );
  NAND2_X1 U9572 ( .A1(n8303), .A2(SI_30_), .ZN(n8304) );
  NAND2_X1 U9573 ( .A1(n8305), .A2(n8304), .ZN(n8315) );
  INV_X1 U9574 ( .A(n8312), .ZN(n8310) );
  MUX2_X1 U9575 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n8306), .Z(n8308) );
  INV_X1 U9576 ( .A(SI_31_), .ZN(n8307) );
  XNOR2_X1 U9577 ( .A(n8308), .B(n8307), .ZN(n8311) );
  INV_X1 U9578 ( .A(n8311), .ZN(n8309) );
  NAND2_X1 U9579 ( .A1(n8310), .A2(n8309), .ZN(n8314) );
  NAND2_X1 U9580 ( .A1(n8312), .A2(n8311), .ZN(n8313) );
  INV_X1 U9581 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n8326) );
  XNOR2_X1 U9582 ( .A(n8316), .B(n8315), .ZN(n9069) );
  NAND2_X1 U9583 ( .A1(n9069), .A2(n6546), .ZN(n8319) );
  NAND2_X1 U9584 ( .A1(n8317), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n8318) );
  NAND2_X1 U9585 ( .A1(n6580), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n8323) );
  NAND2_X1 U9586 ( .A1(n6520), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n8322) );
  NAND2_X1 U9587 ( .A1(n5132), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n8321) );
  AND3_X1 U9588 ( .A1(n8323), .A2(n8322), .A3(n8321), .ZN(n8823) );
  INV_X1 U9589 ( .A(n8324), .ZN(n8325) );
  OR2_X1 U9590 ( .A1(n8823), .A2(n8325), .ZN(n10415) );
  AND2_X1 U9591 ( .A1(n10419), .A2(n10415), .ZN(n8328) );
  MUX2_X1 U9592 ( .A(n8326), .B(n8328), .S(n11171), .Z(n8327) );
  OAI21_X1 U9593 ( .B1(n10416), .B2(n10644), .A(n8327), .ZN(P1_U3553) );
  INV_X1 U9594 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n8329) );
  MUX2_X1 U9595 ( .A(n8329), .B(n8328), .S(n11175), .Z(n8330) );
  OAI21_X1 U9596 ( .B1(n10416), .B2(n10685), .A(n8330), .ZN(P1_U3521) );
  INV_X1 U9597 ( .A(n6779), .ZN(n10699) );
  OAI222_X1 U9598 ( .A1(n9619), .A2(n10699), .B1(n8332), .B2(P2_U3151), .C1(
        n8331), .C2(n9614), .ZN(P2_U3266) );
  NAND2_X1 U9599 ( .A1(n8333), .A2(n10575), .ZN(n8341) );
  INV_X1 U9600 ( .A(n8334), .ZN(n8337) );
  AOI22_X1 U9601 ( .A1(n11011), .A2(P1_REG2_REG_29__SCAN_IN), .B1(n8335), .B2(
        n11149), .ZN(n8336) );
  OAI21_X1 U9602 ( .B1(n8337), .B2(n11014), .A(n8336), .ZN(n8338) );
  AOI21_X1 U9603 ( .B1(n8339), .B2(n11018), .A(n8338), .ZN(n8340) );
  OAI211_X1 U9604 ( .C1(n8342), .C2(n11011), .A(n8341), .B(n8340), .ZN(
        P1_U3356) );
  INV_X1 U9605 ( .A(n8343), .ZN(n8349) );
  INV_X1 U9606 ( .A(n8814), .ZN(n8344) );
  AOI22_X1 U9607 ( .A1(n11011), .A2(P1_REG2_REG_28__SCAN_IN), .B1(n8344), .B2(
        n11149), .ZN(n8345) );
  OAI21_X1 U9608 ( .B1(n8807), .B2(n11014), .A(n8345), .ZN(n8348) );
  NOR2_X1 U9609 ( .A1(n8346), .A2(n11011), .ZN(n8347) );
  AOI211_X1 U9610 ( .C1(n11018), .C2(n8349), .A(n8348), .B(n8347), .ZN(n8350)
         );
  OAI21_X1 U9611 ( .B1(n8351), .B2(n10563), .A(n8350), .ZN(P1_U3265) );
  XOR2_X1 U9612 ( .A(n8353), .B(n8352), .Z(n8372) );
  INV_X1 U9613 ( .A(P2_ADDR_REG_2__SCAN_IN), .ZN(n8355) );
  OAI22_X1 U9614 ( .A1(n10938), .A2(n8355), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8354), .ZN(n8371) );
  INV_X1 U9615 ( .A(n8356), .ZN(n8361) );
  INV_X1 U9616 ( .A(n8357), .ZN(n8360) );
  INV_X1 U9617 ( .A(n8358), .ZN(n8359) );
  AOI21_X1 U9618 ( .B1(n8361), .B2(n8360), .A(n8359), .ZN(n8369) );
  INV_X1 U9619 ( .A(n8362), .ZN(n8367) );
  INV_X1 U9620 ( .A(n8363), .ZN(n8366) );
  AOI21_X1 U9621 ( .B1(n8367), .B2(n8366), .A(n8365), .ZN(n8368) );
  OAI22_X1 U9622 ( .A1(n8369), .A2(n10974), .B1(n10969), .B2(n8368), .ZN(n8370) );
  AOI211_X1 U9623 ( .C1(n10962), .C2(n8372), .A(n8371), .B(n8370), .ZN(n8373)
         );
  OAI21_X1 U9624 ( .B1(n8375), .B2(n10976), .A(n8373), .ZN(P2_U3184) );
  OAI222_X1 U9625 ( .A1(n9614), .A2(n5752), .B1(n8375), .B2(P2_U3151), .C1(
        n9619), .C2(n8374), .ZN(P2_U3293) );
  AOI22_X1 U9626 ( .A1(n10818), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_14__SCAN_IN), .B2(n10695), .ZN(n8376) );
  OAI21_X1 U9627 ( .B1(n8377), .B2(n10704), .A(n8376), .ZN(P1_U3341) );
  XNOR2_X1 U9628 ( .A(n9545), .B(n6905), .ZN(n8409) );
  XNOR2_X1 U9629 ( .A(n8409), .B(n9461), .ZN(n8411) );
  XNOR2_X1 U9630 ( .A(n9129), .B(n6905), .ZN(n8382) );
  XOR2_X1 U9631 ( .A(n9247), .B(n8382), .Z(n9122) );
  INV_X1 U9632 ( .A(n9122), .ZN(n8379) );
  AND2_X1 U9633 ( .A1(n8379), .A2(n9120), .ZN(n8380) );
  NAND2_X1 U9634 ( .A1(n8382), .A2(n8381), .ZN(n8383) );
  XNOR2_X1 U9635 ( .A(n8477), .B(n6905), .ZN(n8384) );
  XOR2_X1 U9636 ( .A(n9246), .B(n8384), .Z(n9225) );
  INV_X1 U9637 ( .A(n8384), .ZN(n8385) );
  NAND2_X1 U9638 ( .A1(n8385), .A2(n9246), .ZN(n8386) );
  NAND2_X1 U9639 ( .A1(n9226), .A2(n8386), .ZN(n9161) );
  XNOR2_X1 U9640 ( .A(n8387), .B(n6905), .ZN(n8388) );
  XNOR2_X1 U9641 ( .A(n8388), .B(n9245), .ZN(n9160) );
  NAND2_X1 U9642 ( .A1(n9161), .A2(n9160), .ZN(n9159) );
  INV_X1 U9643 ( .A(n8388), .ZN(n8389) );
  NAND2_X1 U9644 ( .A1(n8389), .A2(n9245), .ZN(n8390) );
  NAND2_X1 U9645 ( .A1(n9159), .A2(n8390), .ZN(n9172) );
  XNOR2_X1 U9646 ( .A(n9178), .B(n6905), .ZN(n8393) );
  XOR2_X1 U9647 ( .A(n9493), .B(n8393), .Z(n9173) );
  NAND2_X1 U9648 ( .A1(n8393), .A2(n9164), .ZN(n8394) );
  XNOR2_X1 U9649 ( .A(n9508), .B(n6905), .ZN(n8397) );
  XOR2_X1 U9650 ( .A(n9244), .B(n8397), .Z(n9202) );
  XNOR2_X1 U9651 ( .A(n9483), .B(n6905), .ZN(n9144) );
  INV_X1 U9652 ( .A(n9144), .ZN(n8399) );
  OR2_X1 U9653 ( .A1(n9202), .A2(n8399), .ZN(n9141) );
  XNOR2_X1 U9654 ( .A(n9549), .B(n6905), .ZN(n8396) );
  AND2_X1 U9655 ( .A1(n8396), .A2(n9477), .ZN(n8402) );
  OR2_X1 U9656 ( .A1(n9141), .A2(n8402), .ZN(n8395) );
  XOR2_X1 U9657 ( .A(n9448), .B(n8396), .Z(n9196) );
  INV_X1 U9658 ( .A(n9196), .ZN(n8401) );
  NAND2_X1 U9659 ( .A1(n8399), .A2(n9494), .ZN(n8400) );
  INV_X1 U9660 ( .A(n8397), .ZN(n8398) );
  NAND2_X1 U9661 ( .A1(n8398), .A2(n9244), .ZN(n9140) );
  OR2_X1 U9662 ( .A1(n8399), .A2(n9140), .ZN(n9142) );
  AND2_X1 U9663 ( .A1(n8400), .A2(n9142), .ZN(n9191) );
  AND2_X1 U9664 ( .A1(n8401), .A2(n9191), .ZN(n9192) );
  NOR2_X1 U9665 ( .A1(n8402), .A2(n9192), .ZN(n8403) );
  XOR2_X1 U9666 ( .A(n8411), .B(n8412), .Z(n8408) );
  AOI22_X1 U9667 ( .A1(n9214), .A2(n9447), .B1(P2_REG3_REG_21__SCAN_IN), .B2(
        P2_U3151), .ZN(n8405) );
  NAND2_X1 U9668 ( .A1(n9229), .A2(n9448), .ZN(n8404) );
  OAI211_X1 U9669 ( .C1(n9217), .C2(n9450), .A(n8405), .B(n8404), .ZN(n8406)
         );
  AOI21_X1 U9670 ( .B1(n9545), .B2(n9219), .A(n8406), .ZN(n8407) );
  OAI21_X1 U9671 ( .B1(n8408), .B2(n9224), .A(n8407), .ZN(P2_U3163) );
  AND2_X1 U9672 ( .A1(n8409), .A2(n9436), .ZN(n8410) );
  XNOR2_X1 U9673 ( .A(n8589), .B(n6905), .ZN(n9081) );
  XNOR2_X1 U9674 ( .A(n9081), .B(n9447), .ZN(n8413) );
  NAND2_X1 U9675 ( .A1(n8414), .A2(n8413), .ZN(n9084) );
  OAI211_X1 U9676 ( .C1(n8414), .C2(n8413), .A(n9084), .B(n9158), .ZN(n8419)
         );
  INV_X1 U9677 ( .A(n8415), .ZN(n9438) );
  AOI22_X1 U9678 ( .A1(n9229), .A2(n9461), .B1(P2_REG3_REG_22__SCAN_IN), .B2(
        P2_U3151), .ZN(n8416) );
  OAI21_X1 U9679 ( .B1(n9435), .B2(n9231), .A(n8416), .ZN(n8417) );
  AOI21_X1 U9680 ( .B1(n9438), .B2(n9234), .A(n8417), .ZN(n8418) );
  OAI211_X1 U9681 ( .C1(n9600), .C2(n9238), .A(n8419), .B(n8418), .ZN(P2_U3175) );
  INV_X1 U9682 ( .A(n8439), .ZN(n8424) );
  NOR2_X1 U9683 ( .A1(n5966), .A2(n9071), .ZN(n8420) );
  NAND2_X1 U9684 ( .A1(n9611), .A2(n8421), .ZN(n8423) );
  INV_X1 U9685 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n9615) );
  OR2_X1 U9686 ( .A1(n5966), .A2(n9615), .ZN(n8422) );
  NAND2_X1 U9687 ( .A1(n5951), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n8431) );
  INV_X1 U9688 ( .A(P2_REG2_REG_31__SCAN_IN), .ZN(n8426) );
  OR2_X1 U9689 ( .A1(n5959), .A2(n8426), .ZN(n8430) );
  INV_X1 U9690 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n8427) );
  OR2_X1 U9691 ( .A1(n8428), .A2(n8427), .ZN(n8429) );
  NAND4_X1 U9692 ( .A1(n8432), .A2(n8431), .A3(n8430), .A4(n8429), .ZN(n9349)
         );
  INV_X1 U9693 ( .A(n9349), .ZN(n8469) );
  OR2_X1 U9694 ( .A1(n9346), .A2(n8469), .ZN(n8622) );
  INV_X1 U9695 ( .A(n9578), .ZN(n8434) );
  INV_X1 U9696 ( .A(n9240), .ZN(n8433) );
  NAND2_X1 U9697 ( .A1(n8434), .A2(n8433), .ZN(n8621) );
  AND2_X1 U9698 ( .A1(n8621), .A2(n8619), .ZN(n8435) );
  NAND2_X1 U9699 ( .A1(n8622), .A2(n8435), .ZN(n8438) );
  NAND2_X1 U9700 ( .A1(n9578), .A2(n9240), .ZN(n8440) );
  INV_X1 U9701 ( .A(n8440), .ZN(n8436) );
  OAI21_X1 U9702 ( .B1(n8436), .B2(n8469), .A(n9346), .ZN(n8437) );
  INV_X1 U9703 ( .A(n8438), .ZN(n8471) );
  XNOR2_X1 U9704 ( .A(n9105), .B(n5137), .ZN(n9368) );
  INV_X1 U9705 ( .A(n9368), .ZN(n9360) );
  NAND2_X1 U9706 ( .A1(n8441), .A2(n8608), .ZN(n9380) );
  NAND2_X1 U9707 ( .A1(n8604), .A2(n8442), .ZN(n9386) );
  XNOR2_X1 U9708 ( .A(n9529), .B(n9389), .ZN(n9400) );
  NAND2_X1 U9709 ( .A1(n8593), .A2(n8592), .ZN(n9424) );
  XNOR2_X1 U9710 ( .A(n8589), .B(n9447), .ZN(n9432) );
  INV_X1 U9711 ( .A(n8443), .ZN(n8459) );
  NOR2_X1 U9712 ( .A1(n5436), .A2(n8444), .ZN(n8448) );
  AND4_X1 U9713 ( .A1(n8448), .A2(n8447), .A3(n8446), .A4(n8445), .ZN(n8451)
         );
  NAND4_X1 U9714 ( .A1(n8451), .A2(n8521), .A3(n8450), .A4(n8449), .ZN(n8452)
         );
  NOR2_X1 U9715 ( .A1(n8453), .A2(n8452), .ZN(n8455) );
  NAND4_X1 U9716 ( .A1(n8457), .A2(n8456), .A3(n8455), .A4(n8454), .ZN(n8458)
         );
  OR4_X1 U9717 ( .A1(n6366), .A2(n8460), .A3(n8459), .A4(n8458), .ZN(n8461) );
  NOR4_X1 U9718 ( .A1(n8461), .A2(n8558), .A3(n8483), .A4(n9501), .ZN(n8463)
         );
  NAND4_X1 U9719 ( .A1(n9466), .A2(n8463), .A3(n9483), .A4(n6374), .ZN(n8464)
         );
  NOR4_X1 U9720 ( .A1(n9424), .A2(n5413), .A3(n5417), .A4(n8464), .ZN(n8467)
         );
  NAND2_X1 U9721 ( .A1(n8466), .A2(n8465), .ZN(n9416) );
  NAND3_X1 U9722 ( .A1(n9400), .A2(n8467), .A3(n9416), .ZN(n8468) );
  NOR4_X1 U9723 ( .A1(n9360), .A2(n9380), .A3(n9386), .A4(n8468), .ZN(n8470)
         );
  NAND2_X1 U9724 ( .A1(n9346), .A2(n8469), .ZN(n8623) );
  OAI21_X1 U9725 ( .B1(n8474), .B2(n6896), .A(n8473), .ZN(n8625) );
  MUX2_X1 U9726 ( .A(n5137), .B(n9105), .S(n8618), .Z(n8611) );
  INV_X1 U9727 ( .A(n8611), .ZN(n8616) );
  MUX2_X1 U9728 ( .A(n9582), .B(n8475), .S(n8618), .Z(n8612) );
  INV_X1 U9729 ( .A(n8612), .ZN(n8615) );
  INV_X1 U9730 ( .A(n9188), .ZN(n9592) );
  MUX2_X1 U9731 ( .A(n9592), .B(n9422), .S(n8618), .Z(n8596) );
  INV_X1 U9732 ( .A(n8596), .ZN(n8599) );
  NAND2_X1 U9733 ( .A1(n9461), .A2(n8588), .ZN(n8587) );
  INV_X1 U9734 ( .A(n8574), .ZN(n8476) );
  NOR2_X1 U9735 ( .A1(n8476), .A2(n9178), .ZN(n8572) );
  OAI21_X1 U9736 ( .B1(n8618), .B2(n9246), .A(n8477), .ZN(n8485) );
  OAI21_X1 U9737 ( .B1(n8588), .B2(n8478), .A(n9239), .ZN(n8484) );
  MUX2_X1 U9738 ( .A(n9247), .B(n9129), .S(n8618), .Z(n8561) );
  NOR4_X1 U9739 ( .A1(n8481), .A2(n8480), .A3(n8561), .A4(n8479), .ZN(n8482)
         );
  AOI211_X1 U9740 ( .C1(n8485), .C2(n8484), .A(n8483), .B(n8482), .ZN(n8569)
         );
  INV_X1 U9741 ( .A(n8491), .ZN(n8487) );
  NAND2_X1 U9742 ( .A1(n8486), .A2(n8487), .ZN(n8488) );
  NAND2_X1 U9743 ( .A1(n8488), .A2(n8489), .ZN(n8494) );
  OAI211_X1 U9744 ( .C1(n8491), .C2(n6896), .A(n8490), .B(n8489), .ZN(n8492)
         );
  NAND2_X1 U9745 ( .A1(n8492), .A2(n8486), .ZN(n8493) );
  MUX2_X1 U9746 ( .A(n8494), .B(n8493), .S(n8618), .Z(n8502) );
  NAND2_X1 U9747 ( .A1(n8505), .A2(n8496), .ZN(n8497) );
  INV_X1 U9748 ( .A(n8499), .ZN(n8500) );
  OAI21_X1 U9749 ( .B1(n8502), .B2(n8501), .A(n8500), .ZN(n8504) );
  INV_X1 U9750 ( .A(n8505), .ZN(n8507) );
  NOR3_X1 U9751 ( .A1(n8514), .A2(n8507), .A3(n8506), .ZN(n8510) );
  INV_X1 U9752 ( .A(n8511), .ZN(n8513) );
  NAND2_X1 U9753 ( .A1(n8519), .A2(n8516), .ZN(n8517) );
  MUX2_X1 U9754 ( .A(n8519), .B(n8518), .S(n8618), .Z(n8520) );
  OAI211_X1 U9755 ( .C1(n8523), .C2(n8522), .A(n8521), .B(n8520), .ZN(n8524)
         );
  INV_X1 U9756 ( .A(n8524), .ZN(n8535) );
  NAND2_X1 U9757 ( .A1(n8532), .A2(n8528), .ZN(n8525) );
  MUX2_X1 U9758 ( .A(n8526), .B(n8525), .S(n8618), .Z(n8527) );
  NOR2_X1 U9759 ( .A1(n8527), .A2(n8539), .ZN(n8541) );
  INV_X1 U9760 ( .A(n8528), .ZN(n8531) );
  INV_X1 U9761 ( .A(n8529), .ZN(n8530) );
  OAI21_X1 U9762 ( .B1(n8531), .B2(n8530), .A(n8541), .ZN(n8533) );
  NAND3_X1 U9763 ( .A1(n8533), .A2(n8542), .A3(n8532), .ZN(n8534) );
  OAI21_X1 U9764 ( .B1(n8544), .B2(n8538), .A(n8545), .ZN(n8537) );
  NAND2_X1 U9765 ( .A1(n8537), .A2(n8536), .ZN(n8549) );
  AOI211_X1 U9766 ( .C1(n8541), .C2(n8540), .A(n8539), .B(n8538), .ZN(n8543)
         );
  AOI21_X1 U9767 ( .B1(n8544), .B2(n8543), .A(n5536), .ZN(n8547) );
  OAI21_X1 U9768 ( .B1(n8547), .B2(n8546), .A(n8545), .ZN(n8548) );
  MUX2_X1 U9769 ( .A(n8549), .B(n8548), .S(n8618), .Z(n8555) );
  MUX2_X1 U9770 ( .A(n8551), .B(n8550), .S(n8618), .Z(n8552) );
  OAI211_X1 U9771 ( .C1(n8555), .C2(n8554), .A(n8553), .B(n8552), .ZN(n8563)
         );
  NOR2_X1 U9772 ( .A1(n11103), .A2(n9126), .ZN(n8556) );
  MUX2_X1 U9773 ( .A(n8557), .B(n8556), .S(n8588), .Z(n8559) );
  AOI211_X1 U9774 ( .C1(n8561), .C2(n8560), .A(n8559), .B(n8558), .ZN(n8562)
         );
  NAND2_X1 U9775 ( .A1(n8563), .A2(n8562), .ZN(n8568) );
  INV_X1 U9776 ( .A(n8565), .ZN(n8566) );
  MUX2_X1 U9777 ( .A(n5531), .B(n8566), .S(n8618), .Z(n8567) );
  INV_X1 U9778 ( .A(n9178), .ZN(n9566) );
  MUX2_X1 U9779 ( .A(n9164), .B(n9566), .S(n8618), .Z(n8570) );
  INV_X1 U9780 ( .A(n8577), .ZN(n8571) );
  NOR3_X1 U9781 ( .A1(n8575), .A2(n9566), .A3(n9501), .ZN(n8576) );
  MUX2_X1 U9782 ( .A(n8588), .B(n9494), .S(n9554), .Z(n8578) );
  AOI21_X1 U9783 ( .B1(n9207), .B2(n8618), .A(n8578), .ZN(n8579) );
  AOI211_X1 U9784 ( .C1(n8580), .C2(n9483), .A(n8579), .B(n9459), .ZN(n8586)
         );
  INV_X1 U9785 ( .A(n8581), .ZN(n8584) );
  INV_X1 U9786 ( .A(n8582), .ZN(n8583) );
  MUX2_X1 U9787 ( .A(n8584), .B(n8583), .S(n8618), .Z(n8585) );
  NOR3_X1 U9788 ( .A1(n9600), .A2(n8588), .A3(n9447), .ZN(n8591) );
  NOR3_X1 U9789 ( .A1(n8589), .A2(n9421), .A3(n8618), .ZN(n8590) );
  MUX2_X1 U9790 ( .A(n8593), .B(n8592), .S(n8618), .Z(n8594) );
  OAI21_X1 U9791 ( .B1(n8597), .B2(n8596), .A(n8595), .ZN(n8598) );
  MUX2_X1 U9792 ( .A(n8602), .B(n8601), .S(n8618), .Z(n8603) );
  INV_X1 U9793 ( .A(n8604), .ZN(n8605) );
  MUX2_X1 U9794 ( .A(n8606), .B(n8605), .S(n8618), .Z(n8607) );
  INV_X1 U9795 ( .A(n8608), .ZN(n8609) );
  MUX2_X1 U9796 ( .A(n8610), .B(n8609), .S(n8618), .Z(n8613) );
  OAI21_X1 U9797 ( .B1(n8616), .B2(n8615), .A(n8614), .ZN(n8617) );
  XOR2_X1 U9798 ( .A(n8618), .B(n8617), .Z(n8620) );
  XNOR2_X1 U9799 ( .A(n8626), .B(n9334), .ZN(n8633) );
  NAND3_X1 U9800 ( .A1(n8628), .A2(n8627), .A3(n9324), .ZN(n8629) );
  OAI211_X1 U9801 ( .C1(n8630), .C2(n8632), .A(n8629), .B(P2_B_REG_SCAN_IN), 
        .ZN(n8631) );
  OAI21_X1 U9802 ( .B1(n8633), .B2(n8632), .A(n8631), .ZN(P2_U3296) );
  NAND2_X1 U9803 ( .A1(n8635), .A2(n8634), .ZN(n8641) );
  NAND2_X1 U9804 ( .A1(n10101), .A2(n8808), .ZN(n8637) );
  NAND2_X1 U9805 ( .A1(n10291), .A2(n5136), .ZN(n8636) );
  NAND2_X1 U9806 ( .A1(n8637), .A2(n8636), .ZN(n8638) );
  XNOR2_X1 U9807 ( .A(n8638), .B(n8781), .ZN(n8642) );
  NAND2_X1 U9808 ( .A1(n10101), .A2(n5136), .ZN(n8640) );
  NAND2_X1 U9809 ( .A1(n10291), .A2(n8692), .ZN(n8639) );
  NAND2_X1 U9810 ( .A1(n8640), .A2(n8639), .ZN(n10093) );
  INV_X1 U9811 ( .A(n8642), .ZN(n8643) );
  NAND2_X1 U9812 ( .A1(n10172), .A2(n8808), .ZN(n8645) );
  OR2_X1 U9813 ( .A1(n10096), .A2(n5152), .ZN(n8644) );
  NAND2_X1 U9814 ( .A1(n8645), .A2(n8644), .ZN(n8646) );
  XNOR2_X1 U9815 ( .A(n8646), .B(n8781), .ZN(n8649) );
  NOR2_X1 U9816 ( .A1(n10096), .A2(n8806), .ZN(n8647) );
  AOI21_X1 U9817 ( .B1(n10172), .B2(n5136), .A(n8647), .ZN(n8648) );
  XNOR2_X1 U9818 ( .A(n8649), .B(n8648), .ZN(n10165) );
  NAND2_X1 U9819 ( .A1(n8649), .A2(n8648), .ZN(n8650) );
  NAND2_X1 U9820 ( .A1(n10080), .A2(n8808), .ZN(n8652) );
  NAND2_X1 U9821 ( .A1(n10289), .A2(n5136), .ZN(n8651) );
  NAND2_X1 U9822 ( .A1(n8652), .A2(n8651), .ZN(n8653) );
  XNOR2_X1 U9823 ( .A(n8653), .B(n8781), .ZN(n8656) );
  NOR2_X1 U9824 ( .A1(n8654), .A2(n8806), .ZN(n8655) );
  AOI21_X1 U9825 ( .B1(n10080), .B2(n5136), .A(n8655), .ZN(n10073) );
  NAND2_X1 U9826 ( .A1(n10072), .A2(n10073), .ZN(n8658) );
  NAND2_X1 U9827 ( .A1(n8657), .A2(n8656), .ZN(n10071) );
  NAND2_X1 U9828 ( .A1(n8658), .A2(n10071), .ZN(n10208) );
  NAND2_X1 U9829 ( .A1(n8663), .A2(n8808), .ZN(n8660) );
  INV_X1 U9830 ( .A(n10119), .ZN(n10288) );
  NAND2_X1 U9831 ( .A1(n10288), .A2(n5136), .ZN(n8659) );
  NAND2_X1 U9832 ( .A1(n8660), .A2(n8659), .ZN(n8661) );
  XNOR2_X1 U9833 ( .A(n8661), .B(n8781), .ZN(n8671) );
  NOR2_X1 U9834 ( .A1(n10119), .A2(n8806), .ZN(n8662) );
  AOI21_X1 U9835 ( .B1(n8663), .B2(n5136), .A(n8662), .ZN(n8672) );
  AND2_X1 U9836 ( .A1(n8671), .A2(n8672), .ZN(n10209) );
  NAND2_X1 U9837 ( .A1(n8670), .A2(n8808), .ZN(n8667) );
  NAND2_X1 U9838 ( .A1(n10287), .A2(n5136), .ZN(n8666) );
  NAND2_X1 U9839 ( .A1(n8667), .A2(n8666), .ZN(n8668) );
  XNOR2_X1 U9840 ( .A(n8668), .B(n8809), .ZN(n8681) );
  NOR2_X1 U9841 ( .A1(n10213), .A2(n8806), .ZN(n8669) );
  AOI21_X1 U9842 ( .B1(n8670), .B2(n5136), .A(n8669), .ZN(n8682) );
  XNOR2_X1 U9843 ( .A(n8681), .B(n8682), .ZN(n10113) );
  INV_X1 U9844 ( .A(n8671), .ZN(n8674) );
  INV_X1 U9845 ( .A(n8672), .ZN(n8673) );
  NAND2_X1 U9846 ( .A1(n8674), .A2(n8673), .ZN(n10207) );
  AND2_X1 U9847 ( .A1(n10113), .A2(n10207), .ZN(n8675) );
  NAND2_X1 U9848 ( .A1(n8680), .A2(n8808), .ZN(n8677) );
  NAND2_X1 U9849 ( .A1(n11115), .A2(n5136), .ZN(n8676) );
  NAND2_X1 U9850 ( .A1(n8677), .A2(n8676), .ZN(n8678) );
  XNOR2_X1 U9851 ( .A(n8678), .B(n8809), .ZN(n8690) );
  NOR2_X1 U9852 ( .A1(n11138), .A2(n8806), .ZN(n8679) );
  AOI21_X1 U9853 ( .B1(n8680), .B2(n5136), .A(n8679), .ZN(n8688) );
  XNOR2_X1 U9854 ( .A(n8690), .B(n8688), .ZN(n10186) );
  INV_X1 U9855 ( .A(n8681), .ZN(n8683) );
  NAND2_X1 U9856 ( .A1(n8683), .A2(n8682), .ZN(n10183) );
  AND2_X1 U9857 ( .A1(n10186), .A2(n10183), .ZN(n8684) );
  NAND2_X1 U9858 ( .A1(n11152), .A2(n8808), .ZN(n8686) );
  NAND2_X1 U9859 ( .A1(n6629), .A2(n5136), .ZN(n8685) );
  NAND2_X1 U9860 ( .A1(n8686), .A2(n8685), .ZN(n8687) );
  XNOR2_X1 U9861 ( .A(n8687), .B(n8781), .ZN(n8696) );
  INV_X1 U9862 ( .A(n8688), .ZN(n8689) );
  NAND2_X1 U9863 ( .A1(n8690), .A2(n8689), .ZN(n8695) );
  AND2_X1 U9864 ( .A1(n8696), .A2(n8695), .ZN(n8691) );
  NAND2_X1 U9865 ( .A1(n11152), .A2(n5136), .ZN(n8694) );
  NAND2_X1 U9866 ( .A1(n6629), .A2(n8692), .ZN(n8693) );
  NAND2_X1 U9867 ( .A1(n8694), .A2(n8693), .ZN(n10050) );
  NAND2_X1 U9868 ( .A1(n10047), .A2(n10050), .ZN(n8699) );
  INV_X1 U9869 ( .A(n8696), .ZN(n8697) );
  NAND2_X1 U9870 ( .A1(n8698), .A2(n8697), .ZN(n10048) );
  NAND2_X1 U9871 ( .A1(n8699), .A2(n10048), .ZN(n10257) );
  NAND2_X1 U9872 ( .A1(n10267), .A2(n8808), .ZN(n8701) );
  NAND2_X1 U9873 ( .A1(n10286), .A2(n5136), .ZN(n8700) );
  NAND2_X1 U9874 ( .A1(n8701), .A2(n8700), .ZN(n8702) );
  XNOR2_X1 U9875 ( .A(n8702), .B(n8781), .ZN(n10255) );
  NOR2_X1 U9876 ( .A1(n11136), .A2(n8806), .ZN(n8703) );
  AOI21_X1 U9877 ( .B1(n10267), .B2(n5136), .A(n8703), .ZN(n8705) );
  NAND2_X1 U9878 ( .A1(n10255), .A2(n8705), .ZN(n8704) );
  NAND2_X1 U9879 ( .A1(n10257), .A2(n8704), .ZN(n8708) );
  INV_X1 U9880 ( .A(n10255), .ZN(n8706) );
  INV_X1 U9881 ( .A(n8705), .ZN(n10254) );
  NAND2_X1 U9882 ( .A1(n8706), .A2(n10254), .ZN(n8707) );
  NAND2_X1 U9883 ( .A1(n8708), .A2(n8707), .ZN(n10134) );
  NAND2_X1 U9884 ( .A1(n10646), .A2(n8808), .ZN(n8710) );
  INV_X1 U9885 ( .A(n10258), .ZN(n10285) );
  NAND2_X1 U9886 ( .A1(n10285), .A2(n5136), .ZN(n8709) );
  NAND2_X1 U9887 ( .A1(n8710), .A2(n8709), .ZN(n8711) );
  XNOR2_X1 U9888 ( .A(n8711), .B(n8781), .ZN(n8713) );
  NOR2_X1 U9889 ( .A1(n10258), .A2(n8806), .ZN(n8712) );
  AOI21_X1 U9890 ( .B1(n10646), .B2(n5136), .A(n8712), .ZN(n8714) );
  NAND2_X1 U9891 ( .A1(n8713), .A2(n8714), .ZN(n8718) );
  INV_X1 U9892 ( .A(n8713), .ZN(n8716) );
  INV_X1 U9893 ( .A(n8714), .ZN(n8715) );
  NAND2_X1 U9894 ( .A1(n8716), .A2(n8715), .ZN(n8717) );
  NAND2_X1 U9895 ( .A1(n8718), .A2(n8717), .ZN(n10135) );
  NAND2_X1 U9896 ( .A1(n8722), .A2(n8808), .ZN(n8720) );
  OR2_X1 U9897 ( .A1(n10237), .A2(n5152), .ZN(n8719) );
  NAND2_X1 U9898 ( .A1(n8720), .A2(n8719), .ZN(n8721) );
  XNOR2_X1 U9899 ( .A(n8721), .B(n8809), .ZN(n8725) );
  NAND2_X1 U9900 ( .A1(n8722), .A2(n5136), .ZN(n8724) );
  OR2_X1 U9901 ( .A1(n10237), .A2(n8806), .ZN(n8723) );
  NAND2_X1 U9902 ( .A1(n8724), .A2(n8723), .ZN(n8726) );
  NAND2_X1 U9903 ( .A1(n8725), .A2(n8726), .ZN(n10143) );
  INV_X1 U9904 ( .A(n8725), .ZN(n8728) );
  INV_X1 U9905 ( .A(n8726), .ZN(n8727) );
  NAND2_X1 U9906 ( .A1(n8728), .A2(n8727), .ZN(n10142) );
  NAND2_X1 U9907 ( .A1(n10636), .A2(n8808), .ZN(n8730) );
  OR2_X1 U9908 ( .A1(n10569), .A2(n5152), .ZN(n8729) );
  NAND2_X1 U9909 ( .A1(n8730), .A2(n8729), .ZN(n8731) );
  XNOR2_X1 U9910 ( .A(n8731), .B(n8781), .ZN(n8734) );
  NOR2_X1 U9911 ( .A1(n10569), .A2(n8806), .ZN(n8733) );
  AOI21_X1 U9912 ( .B1(n10636), .B2(n5136), .A(n8733), .ZN(n10229) );
  NAND2_X1 U9913 ( .A1(n10227), .A2(n10229), .ZN(n8736) );
  NAND2_X1 U9914 ( .A1(n8735), .A2(n8734), .ZN(n10228) );
  NAND2_X1 U9915 ( .A1(n8736), .A2(n10228), .ZN(n10084) );
  NAND2_X1 U9916 ( .A1(n10579), .A2(n8808), .ZN(n8738) );
  NAND2_X1 U9917 ( .A1(n10282), .A2(n5136), .ZN(n8737) );
  NAND2_X1 U9918 ( .A1(n8738), .A2(n8737), .ZN(n8739) );
  XNOR2_X1 U9919 ( .A(n8739), .B(n8809), .ZN(n8741) );
  NOR2_X1 U9920 ( .A1(n10550), .A2(n8806), .ZN(n8740) );
  AOI21_X1 U9921 ( .B1(n10579), .B2(n5136), .A(n8740), .ZN(n8742) );
  XNOR2_X1 U9922 ( .A(n8741), .B(n8742), .ZN(n10083) );
  NAND2_X1 U9923 ( .A1(n10084), .A2(n10083), .ZN(n8745) );
  INV_X1 U9924 ( .A(n8741), .ZN(n8743) );
  NAND2_X1 U9925 ( .A1(n8743), .A2(n8742), .ZN(n8744) );
  NAND2_X1 U9926 ( .A1(n8745), .A2(n8744), .ZN(n10175) );
  NAND2_X1 U9927 ( .A1(n10626), .A2(n8808), .ZN(n8747) );
  OR2_X1 U9928 ( .A1(n10568), .A2(n5152), .ZN(n8746) );
  NAND2_X1 U9929 ( .A1(n8747), .A2(n8746), .ZN(n8748) );
  XNOR2_X1 U9930 ( .A(n8748), .B(n8809), .ZN(n8750) );
  NOR2_X1 U9931 ( .A1(n10568), .A2(n8806), .ZN(n8749) );
  AOI21_X1 U9932 ( .B1(n10626), .B2(n5136), .A(n8749), .ZN(n8751) );
  XNOR2_X1 U9933 ( .A(n8750), .B(n8751), .ZN(n10176) );
  NAND2_X1 U9934 ( .A1(n10175), .A2(n10176), .ZN(n8754) );
  INV_X1 U9935 ( .A(n8750), .ZN(n8752) );
  NAND2_X1 U9936 ( .A1(n8752), .A2(n8751), .ZN(n8753) );
  NAND2_X1 U9937 ( .A1(n8754), .A2(n8753), .ZN(n10104) );
  NAND2_X1 U9938 ( .A1(n10538), .A2(n8808), .ZN(n8756) );
  NAND2_X1 U9939 ( .A1(n10280), .A2(n5136), .ZN(n8755) );
  NAND2_X1 U9940 ( .A1(n8756), .A2(n8755), .ZN(n8757) );
  XNOR2_X1 U9941 ( .A(n8757), .B(n8781), .ZN(n8761) );
  NOR2_X1 U9942 ( .A1(n10551), .A2(n8806), .ZN(n8758) );
  AOI21_X1 U9943 ( .B1(n10538), .B2(n5136), .A(n8758), .ZN(n8762) );
  XNOR2_X1 U9944 ( .A(n8761), .B(n8762), .ZN(n10105) );
  INV_X1 U9945 ( .A(n8761), .ZN(n8764) );
  INV_X1 U9946 ( .A(n8762), .ZN(n8763) );
  NAND2_X1 U9947 ( .A1(n8764), .A2(n8763), .ZN(n8765) );
  AOI22_X1 U9948 ( .A1(n10068), .A2(n8808), .B1(n5136), .B2(n10278), .ZN(n8766) );
  XNOR2_X1 U9949 ( .A(n8766), .B(n8809), .ZN(n10061) );
  NOR2_X1 U9950 ( .A1(n10515), .A2(n8806), .ZN(n8767) );
  AOI21_X1 U9951 ( .B1(n10068), .B2(n5136), .A(n8767), .ZN(n10060) );
  NOR2_X1 U9952 ( .A1(n10531), .A2(n8806), .ZN(n8768) );
  AOI21_X1 U9953 ( .B1(n10613), .B2(n5136), .A(n8768), .ZN(n10197) );
  NAND2_X1 U9954 ( .A1(n10613), .A2(n8808), .ZN(n8770) );
  NAND2_X1 U9955 ( .A1(n10279), .A2(n5136), .ZN(n8769) );
  NAND2_X1 U9956 ( .A1(n8770), .A2(n8769), .ZN(n8771) );
  XNOR2_X1 U9957 ( .A(n8771), .B(n8781), .ZN(n10058) );
  OAI22_X1 U9958 ( .A1(n10061), .A2(n10060), .B1(n10197), .B2(n10058), .ZN(
        n8778) );
  INV_X1 U9959 ( .A(n10060), .ZN(n8773) );
  NAND2_X1 U9960 ( .A1(n10058), .A2(n10197), .ZN(n8774) );
  INV_X1 U9961 ( .A(n10061), .ZN(n8772) );
  AOI21_X1 U9962 ( .B1(n8773), .B2(n8774), .A(n8772), .ZN(n8777) );
  INV_X1 U9963 ( .A(n8774), .ZN(n8775) );
  NAND2_X1 U9964 ( .A1(n10603), .A2(n8808), .ZN(n8780) );
  NAND2_X1 U9965 ( .A1(n10277), .A2(n5136), .ZN(n8779) );
  NAND2_X1 U9966 ( .A1(n8780), .A2(n8779), .ZN(n8782) );
  XNOR2_X1 U9967 ( .A(n8782), .B(n8781), .ZN(n8785) );
  NOR2_X1 U9968 ( .A1(n10496), .A2(n8806), .ZN(n8783) );
  AOI21_X1 U9969 ( .B1(n10603), .B2(n5136), .A(n8783), .ZN(n8784) );
  NOR2_X1 U9970 ( .A1(n8785), .A2(n8784), .ZN(n10155) );
  NAND2_X1 U9971 ( .A1(n8785), .A2(n8784), .ZN(n10153) );
  OAI22_X1 U9972 ( .A1(n6745), .A2(n5152), .B1(n10484), .B2(n8806), .ZN(n8794)
         );
  NAND2_X1 U9973 ( .A1(n10468), .A2(n8808), .ZN(n8787) );
  NAND2_X1 U9974 ( .A1(n10276), .A2(n5136), .ZN(n8786) );
  NAND2_X1 U9975 ( .A1(n8787), .A2(n8786), .ZN(n8788) );
  XNOR2_X1 U9976 ( .A(n8788), .B(n8809), .ZN(n8793) );
  XOR2_X1 U9977 ( .A(n8794), .B(n8793), .Z(n10125) );
  NAND2_X1 U9978 ( .A1(n10124), .A2(n10125), .ZN(n10242) );
  NAND2_X1 U9979 ( .A1(n10450), .A2(n8808), .ZN(n8790) );
  NAND2_X1 U9980 ( .A1(n10275), .A2(n5136), .ZN(n8789) );
  NAND2_X1 U9981 ( .A1(n8790), .A2(n8789), .ZN(n8791) );
  XNOR2_X1 U9982 ( .A(n8791), .B(n8809), .ZN(n8803) );
  NOR2_X1 U9983 ( .A1(n10462), .A2(n8806), .ZN(n8792) );
  AOI21_X1 U9984 ( .B1(n10450), .B2(n5136), .A(n8792), .ZN(n8801) );
  XNOR2_X1 U9985 ( .A(n8803), .B(n8801), .ZN(n10245) );
  INV_X1 U9986 ( .A(n8793), .ZN(n8796) );
  INV_X1 U9987 ( .A(n8794), .ZN(n8795) );
  NAND2_X1 U9988 ( .A1(n8796), .A2(n8795), .ZN(n10241) );
  OAI22_X1 U9989 ( .A1(n10656), .A2(n7484), .B1(n10446), .B2(n5152), .ZN(n8798) );
  XNOR2_X1 U9990 ( .A(n8798), .B(n8809), .ZN(n8800) );
  OAI22_X1 U9991 ( .A1(n10656), .A2(n5152), .B1(n10446), .B2(n8806), .ZN(n8799) );
  NOR2_X1 U9992 ( .A1(n8800), .A2(n8799), .ZN(n8805) );
  AOI21_X1 U9993 ( .B1(n8800), .B2(n8799), .A(n8805), .ZN(n10042) );
  INV_X1 U9994 ( .A(n8801), .ZN(n8802) );
  NAND2_X1 U9995 ( .A1(n8803), .A2(n8802), .ZN(n10043) );
  OAI22_X1 U9996 ( .A1(n8807), .A2(n5152), .B1(n10426), .B2(n8806), .ZN(n8812)
         );
  AOI22_X1 U9997 ( .A1(n8819), .A2(n8808), .B1(n5136), .B2(n10273), .ZN(n8810)
         );
  XNOR2_X1 U9998 ( .A(n8810), .B(n8809), .ZN(n8811) );
  NOR2_X1 U9999 ( .A1(n10263), .A2(n8814), .ZN(n8818) );
  INV_X1 U10000 ( .A(n10446), .ZN(n10274) );
  AOI22_X1 U10001 ( .A1(n10261), .A2(n10274), .B1(P1_REG3_REG_28__SCAN_IN), 
        .B2(P1_U3086), .ZN(n8815) );
  OAI21_X1 U10002 ( .B1(n8816), .B2(n10259), .A(n8815), .ZN(n8817) );
  AOI211_X1 U10003 ( .C1(n8819), .C2(n10266), .A(n8818), .B(n8817), .ZN(n8820)
         );
  OAI21_X1 U10004 ( .B1(n8821), .B2(n10269), .A(n8820), .ZN(P1_U3220) );
  INV_X1 U10005 ( .A(n8823), .ZN(n10271) );
  AOI21_X1 U10006 ( .B1(n10272), .B2(n10271), .A(n8822), .ZN(n8826) );
  NAND2_X1 U10007 ( .A1(n9062), .A2(n7110), .ZN(n8920) );
  NAND2_X1 U10008 ( .A1(n8827), .A2(n8920), .ZN(n8830) );
  NOR3_X1 U10009 ( .A1(n8919), .A2(n8825), .A3(n8830), .ZN(n8824) );
  AOI211_X1 U10010 ( .C1(n8826), .C2(n8920), .A(n9055), .B(n8824), .ZN(n8926)
         );
  INV_X1 U10011 ( .A(n8825), .ZN(n9048) );
  OAI33_X1 U10012 ( .A1(n8830), .A2(n8919), .A3(n9053), .B1(n8920), .B2(n9048), 
        .B3(n8826), .ZN(n8925) );
  INV_X1 U10013 ( .A(n8827), .ZN(n8829) );
  NOR2_X1 U10014 ( .A1(n8829), .A2(n8828), .ZN(n9050) );
  INV_X1 U10015 ( .A(n8830), .ZN(n8918) );
  NAND2_X1 U10016 ( .A1(n8905), .A2(n8908), .ZN(n9041) );
  NOR2_X1 U10017 ( .A1(n9041), .A2(n8920), .ZN(n8907) );
  NAND2_X1 U10018 ( .A1(n8977), .A2(n8831), .ZN(n8982) );
  NAND2_X1 U10019 ( .A1(n8901), .A2(n8832), .ZN(n8978) );
  INV_X1 U10020 ( .A(n8920), .ZN(n8892) );
  MUX2_X1 U10021 ( .A(n8982), .B(n8978), .S(n8892), .Z(n8904) );
  AOI21_X1 U10022 ( .B1(n10525), .B2(n8983), .A(n8892), .ZN(n8896) );
  NAND3_X1 U10023 ( .A1(n8833), .A2(n8988), .A3(n8993), .ZN(n8835) );
  NAND3_X1 U10024 ( .A1(n8835), .A2(n8837), .A3(n8834), .ZN(n8841) );
  AND2_X1 U10025 ( .A1(n8837), .A2(n8836), .ZN(n8990) );
  OAI21_X1 U10026 ( .B1(n10998), .B2(n10997), .A(n8990), .ZN(n8839) );
  AND2_X1 U10027 ( .A1(n8993), .A2(n8842), .ZN(n8838) );
  AOI21_X1 U10028 ( .B1(n8839), .B2(n8838), .A(n8992), .ZN(n8840) );
  MUX2_X1 U10029 ( .A(n8841), .B(n8840), .S(n8892), .Z(n8847) );
  NAND2_X1 U10030 ( .A1(n8843), .A2(n8842), .ZN(n8996) );
  NAND2_X1 U10031 ( .A1(n8996), .A2(n8995), .ZN(n8844) );
  MUX2_X1 U10032 ( .A(n8995), .B(n8844), .S(n8920), .Z(n8845) );
  OAI211_X1 U10033 ( .C1(n8847), .C2(n8932), .A(n8846), .B(n8845), .ZN(n8852)
         );
  MUX2_X1 U10034 ( .A(n8933), .B(n8848), .S(n8920), .Z(n8850) );
  NOR2_X1 U10035 ( .A1(n8850), .A2(n8849), .ZN(n8851) );
  NAND2_X1 U10036 ( .A1(n8852), .A2(n8851), .ZN(n8854) );
  AND2_X1 U10037 ( .A1(n8927), .A2(n8936), .ZN(n8857) );
  AND2_X1 U10038 ( .A1(n8867), .A2(n8855), .ZN(n8856) );
  MUX2_X1 U10039 ( .A(n8857), .B(n8856), .S(n8920), .Z(n8858) );
  NAND4_X1 U10040 ( .A1(n8859), .A2(n8858), .A3(n8862), .A4(n8860), .ZN(n8868)
         );
  INV_X1 U10041 ( .A(n8860), .ZN(n8861) );
  NAND2_X1 U10042 ( .A1(n8862), .A2(n8861), .ZN(n8863) );
  NAND4_X1 U10043 ( .A1(n8868), .A2(n8864), .A3(n8867), .A4(n8863), .ZN(n8866)
         );
  NAND3_X1 U10044 ( .A1(n8866), .A2(n8865), .A3(n8874), .ZN(n8871) );
  INV_X1 U10045 ( .A(n8867), .ZN(n9002) );
  OAI211_X1 U10046 ( .C1(n9002), .C2(n8927), .A(n8868), .B(n9005), .ZN(n8869)
         );
  NAND2_X1 U10047 ( .A1(n8869), .A2(n8985), .ZN(n8870) );
  MUX2_X1 U10048 ( .A(n8871), .B(n8870), .S(n8920), .Z(n8876) );
  NAND2_X1 U10049 ( .A1(n8878), .A2(n8873), .ZN(n8984) );
  AND2_X1 U10050 ( .A1(n11130), .A2(n8874), .ZN(n9010) );
  NAND2_X1 U10051 ( .A1(n9019), .A2(n8878), .ZN(n8880) );
  NAND2_X1 U10052 ( .A1(n9020), .A2(n9015), .ZN(n8879) );
  MUX2_X1 U10053 ( .A(n8880), .B(n8879), .S(n8892), .Z(n8882) );
  MUX2_X1 U10054 ( .A(n9019), .B(n9020), .S(n8920), .Z(n8881) );
  OAI211_X1 U10055 ( .C1(n8883), .C2(n8882), .A(n8952), .B(n8881), .ZN(n8888)
         );
  AND2_X1 U10056 ( .A1(n8889), .A2(n8884), .ZN(n9026) );
  INV_X1 U10057 ( .A(n8887), .ZN(n9024) );
  AOI21_X1 U10058 ( .B1(n8888), .B2(n9026), .A(n9024), .ZN(n8885) );
  OR2_X1 U10059 ( .A1(n10579), .A2(n10550), .ZN(n8886) );
  AND2_X1 U10060 ( .A1(n10526), .A2(n8886), .ZN(n9027) );
  NAND3_X1 U10061 ( .A1(n8888), .A2(n8887), .A3(n9021), .ZN(n8890) );
  NAND3_X1 U10062 ( .A1(n8890), .A2(n8983), .A3(n8889), .ZN(n8891) );
  NAND2_X1 U10063 ( .A1(n9030), .A2(n8892), .ZN(n8899) );
  NAND2_X1 U10064 ( .A1(n9030), .A2(n10526), .ZN(n8894) );
  OAI21_X1 U10065 ( .B1(n10525), .B2(n8920), .A(n8897), .ZN(n8893) );
  AOI21_X1 U10066 ( .B1(n8899), .B2(n8894), .A(n8893), .ZN(n8895) );
  NAND2_X1 U10067 ( .A1(n8897), .A2(n8920), .ZN(n8898) );
  NAND2_X1 U10068 ( .A1(n8899), .A2(n8898), .ZN(n8900) );
  MUX2_X1 U10069 ( .A(n8977), .B(n8901), .S(n8920), .Z(n8902) );
  OAI211_X1 U10070 ( .C1(n8904), .C2(n8903), .A(n8955), .B(n8902), .ZN(n8909)
         );
  NAND2_X1 U10071 ( .A1(n9039), .A2(n8920), .ZN(n8910) );
  OAI22_X1 U10072 ( .A1(n8910), .A2(n8905), .B1(n8920), .B2(n9039), .ZN(n8906)
         );
  INV_X1 U10073 ( .A(n8908), .ZN(n8913) );
  AOI21_X1 U10074 ( .B1(n8909), .B2(n9035), .A(n10443), .ZN(n8912) );
  INV_X1 U10075 ( .A(n8910), .ZN(n8911) );
  OAI21_X1 U10076 ( .B1(n8913), .B2(n8912), .A(n8911), .ZN(n8914) );
  MUX2_X1 U10077 ( .A(n9044), .B(n9040), .S(n8920), .Z(n8916) );
  INV_X1 U10078 ( .A(n9045), .ZN(n8915) );
  OAI21_X1 U10079 ( .B1(n9050), .B2(n8918), .A(n8917), .ZN(n8924) );
  INV_X1 U10080 ( .A(n8919), .ZN(n8922) );
  INV_X1 U10081 ( .A(n9053), .ZN(n8921) );
  AOI21_X1 U10082 ( .B1(n8922), .B2(n8921), .A(n8920), .ZN(n8923) );
  INV_X1 U10083 ( .A(n10564), .ZN(n10573) );
  INV_X1 U10084 ( .A(n8927), .ZN(n8941) );
  INV_X1 U10085 ( .A(n8928), .ZN(n8930) );
  NOR4_X1 U10086 ( .A1(n10997), .A2(n6814), .A3(n8930), .A4(n8929), .ZN(n8938)
         );
  NOR4_X1 U10087 ( .A1(n8934), .A2(n8933), .A3(n8932), .A4(n8931), .ZN(n8937)
         );
  NAND4_X1 U10088 ( .A1(n8938), .A2(n8937), .A3(n8936), .A4(n8935), .ZN(n8939)
         );
  NOR4_X1 U10089 ( .A1(n8942), .A2(n8941), .A3(n8940), .A4(n8939), .ZN(n8943)
         );
  NAND4_X1 U10090 ( .A1(n8946), .A2(n8945), .A3(n8944), .A4(n8943), .ZN(n8947)
         );
  NOR4_X1 U10091 ( .A1(n8949), .A2(n8948), .A3(n8947), .A4(n11120), .ZN(n8950)
         );
  NAND4_X1 U10092 ( .A1(n10528), .A2(n8952), .A3(n8951), .A4(n8950), .ZN(n8953) );
  NOR4_X1 U10093 ( .A1(n10513), .A2(n10573), .A3(n10546), .A4(n8953), .ZN(
        n8954) );
  NAND4_X1 U10094 ( .A1(n10458), .A2(n8955), .A3(n10495), .A4(n8954), .ZN(
        n8956) );
  NOR4_X1 U10095 ( .A1(n8957), .A2(n10430), .A3(n10442), .A4(n8956), .ZN(n8960) );
  INV_X1 U10096 ( .A(n8822), .ZN(n8959) );
  INV_X1 U10097 ( .A(n10272), .ZN(n8958) );
  NAND2_X1 U10098 ( .A1(n8959), .A2(n8958), .ZN(n9046) );
  NAND4_X1 U10099 ( .A1(n9051), .A2(n8961), .A3(n8960), .A4(n9046), .ZN(n8962)
         );
  NOR3_X1 U10100 ( .A1(n9053), .A2(n9055), .A3(n8962), .ZN(n8966) );
  NAND2_X1 U10101 ( .A1(n8964), .A2(n8963), .ZN(n8970) );
  INV_X1 U10102 ( .A(n8966), .ZN(n8967) );
  NAND2_X1 U10103 ( .A1(n8968), .A2(n6812), .ZN(n8969) );
  NAND2_X1 U10104 ( .A1(n8970), .A2(n8969), .ZN(n8976) );
  INV_X1 U10105 ( .A(n9055), .ZN(n8972) );
  NAND2_X1 U10106 ( .A1(n8972), .A2(n6796), .ZN(n8973) );
  NOR2_X1 U10107 ( .A1(n8976), .A2(n8975), .ZN(n9068) );
  NAND2_X1 U10108 ( .A1(n8978), .A2(n8977), .ZN(n8979) );
  NAND2_X1 U10109 ( .A1(n8980), .A2(n8979), .ZN(n8981) );
  NAND2_X1 U10110 ( .A1(n8981), .A2(n9035), .ZN(n9037) );
  INV_X1 U10111 ( .A(n8982), .ZN(n9034) );
  INV_X1 U10112 ( .A(n8983), .ZN(n9029) );
  INV_X1 U10113 ( .A(n8984), .ZN(n9018) );
  INV_X1 U10114 ( .A(n8985), .ZN(n9009) );
  NAND2_X1 U10115 ( .A1(n11000), .A2(n10987), .ZN(n8986) );
  NAND3_X1 U10116 ( .A1(n8987), .A2(n6814), .A3(n8986), .ZN(n8989) );
  NAND2_X1 U10117 ( .A1(n8989), .A2(n8988), .ZN(n8991) );
  OAI21_X1 U10118 ( .B1(n10998), .B2(n8991), .A(n8990), .ZN(n8994) );
  AOI21_X1 U10119 ( .B1(n8994), .B2(n8993), .A(n8992), .ZN(n8997) );
  OAI21_X1 U10120 ( .B1(n8997), .B2(n8996), .A(n8995), .ZN(n8999) );
  NAND2_X1 U10121 ( .A1(n8999), .A2(n8998), .ZN(n9000) );
  NAND2_X1 U10122 ( .A1(n9001), .A2(n9000), .ZN(n9004) );
  AOI21_X1 U10123 ( .B1(n9004), .B2(n9003), .A(n9002), .ZN(n9007) );
  INV_X1 U10124 ( .A(n9005), .ZN(n9006) );
  NOR2_X1 U10125 ( .A1(n9007), .A2(n9006), .ZN(n9008) );
  NOR2_X1 U10126 ( .A1(n9009), .A2(n9008), .ZN(n9014) );
  INV_X1 U10127 ( .A(n9010), .ZN(n9013) );
  OAI211_X1 U10128 ( .C1(n9014), .C2(n9013), .A(n9012), .B(n9011), .ZN(n9017)
         );
  INV_X1 U10129 ( .A(n9015), .ZN(n9016) );
  AOI21_X1 U10130 ( .B1(n9018), .B2(n9017), .A(n9016), .ZN(n9023) );
  INV_X1 U10131 ( .A(n9019), .ZN(n9022) );
  OAI211_X1 U10132 ( .C1(n9023), .C2(n9022), .A(n9021), .B(n9020), .ZN(n9025)
         );
  AOI21_X1 U10133 ( .B1(n9026), .B2(n9025), .A(n9024), .ZN(n9028) );
  OAI211_X1 U10134 ( .C1(n9029), .C2(n9028), .A(n9030), .B(n9027), .ZN(n9033)
         );
  NAND2_X1 U10135 ( .A1(n9031), .A2(n9030), .ZN(n9032) );
  NAND4_X1 U10136 ( .A1(n9035), .A2(n9034), .A3(n9033), .A4(n9032), .ZN(n9036)
         );
  AND3_X1 U10137 ( .A1(n9038), .A2(n9037), .A3(n9036), .ZN(n9042) );
  OAI211_X1 U10138 ( .C1(n9042), .C2(n9041), .A(n9040), .B(n9039), .ZN(n9043)
         );
  NAND3_X1 U10139 ( .A1(n9045), .A2(n9044), .A3(n9043), .ZN(n9049) );
  INV_X1 U10140 ( .A(n9046), .ZN(n9047) );
  AOI211_X1 U10141 ( .C1(n9050), .C2(n9049), .A(n9048), .B(n9047), .ZN(n9054)
         );
  INV_X1 U10142 ( .A(n9051), .ZN(n9052) );
  NOR3_X1 U10143 ( .A1(n9054), .A2(n9053), .A3(n9052), .ZN(n9056) );
  NOR2_X1 U10144 ( .A1(n9056), .A2(n9055), .ZN(n9060) );
  NAND2_X1 U10145 ( .A1(n9060), .A2(n7107), .ZN(n9058) );
  OAI211_X1 U10146 ( .C1(n9060), .C2(n9059), .A(n9058), .B(n9057), .ZN(n9067)
         );
  INV_X1 U10147 ( .A(n9061), .ZN(n9063) );
  NAND3_X1 U10148 ( .A1(n9063), .A2(P1_STATE_REG_SCAN_IN), .A3(n9062), .ZN(
        n9064) );
  OAI211_X1 U10149 ( .C1(n9065), .C2(n10310), .A(P1_B_REG_SCAN_IN), .B(n9064), 
        .ZN(n9066) );
  OAI21_X1 U10150 ( .B1(n9068), .B2(n9067), .A(n9066), .ZN(P1_U3242) );
  INV_X1 U10151 ( .A(n9069), .ZN(n9079) );
  OAI222_X1 U10152 ( .A1(n9614), .A2(n9071), .B1(n9619), .B2(n9079), .C1(
        P2_U3151), .C2(n9070), .ZN(P2_U3265) );
  INV_X1 U10153 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n9074) );
  OAI211_X1 U10154 ( .C1(n9073), .C2(n8822), .A(n11126), .B(n9072), .ZN(n10423) );
  AND2_X1 U10155 ( .A1(n10423), .A2(n10415), .ZN(n9076) );
  MUX2_X1 U10156 ( .A(n9074), .B(n9076), .S(n11175), .Z(n9075) );
  OAI21_X1 U10157 ( .B1(n8822), .B2(n10685), .A(n9075), .ZN(P1_U3520) );
  INV_X1 U10158 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n9077) );
  MUX2_X1 U10159 ( .A(n9077), .B(n9076), .S(n11171), .Z(n9078) );
  OAI21_X1 U10160 ( .B1(n8822), .B2(n10644), .A(n9078), .ZN(P1_U3552) );
  OAI222_X1 U10161 ( .A1(n9080), .A2(P1_U3086), .B1(n10704), .B2(n9079), .C1(
        n9933), .C2(n10701), .ZN(P1_U3325) );
  INV_X1 U10162 ( .A(n9081), .ZN(n9082) );
  NAND2_X1 U10163 ( .A1(n9082), .A2(n9447), .ZN(n9083) );
  NAND2_X1 U10164 ( .A1(n9084), .A2(n9083), .ZN(n9085) );
  XNOR2_X1 U10165 ( .A(n9425), .B(n6905), .ZN(n9086) );
  INV_X1 U10166 ( .A(n9085), .ZN(n9087) );
  NAND2_X1 U10167 ( .A1(n9087), .A2(n9086), .ZN(n9182) );
  XNOR2_X1 U10168 ( .A(n9188), .B(n6905), .ZN(n9089) );
  NAND2_X1 U10169 ( .A1(n9089), .A2(n9422), .ZN(n9088) );
  INV_X1 U10170 ( .A(n9088), .ZN(n9090) );
  XNOR2_X1 U10171 ( .A(n9089), .B(n9242), .ZN(n9184) );
  OR2_X1 U10172 ( .A1(n9090), .A2(n9184), .ZN(n9091) );
  INV_X1 U10173 ( .A(n9091), .ZN(n9092) );
  XNOR2_X1 U10174 ( .A(n9529), .B(n6905), .ZN(n9094) );
  XNOR2_X1 U10175 ( .A(n9094), .B(n9389), .ZN(n9152) );
  NAND2_X1 U10176 ( .A1(n9094), .A2(n9412), .ZN(n9095) );
  XNOR2_X1 U10177 ( .A(n9220), .B(n6905), .ZN(n9096) );
  NAND2_X1 U10178 ( .A1(n9096), .A2(n9403), .ZN(n9097) );
  XNOR2_X1 U10179 ( .A(n9099), .B(n9098), .ZN(n9100) );
  NAND2_X1 U10180 ( .A1(n9100), .A2(n9390), .ZN(n9101) );
  OAI21_X1 U10181 ( .B1(n9100), .B2(n9390), .A(n9101), .ZN(n9111) );
  AOI22_X1 U10182 ( .A1(n9229), .A2(n9390), .B1(P2_REG3_REG_28__SCAN_IN), .B2(
        P2_U3151), .ZN(n9103) );
  NAND2_X1 U10183 ( .A1(n9214), .A2(n9241), .ZN(n9102) );
  OAI211_X1 U10184 ( .C1(n9217), .C2(n9370), .A(n9103), .B(n9102), .ZN(n9104)
         );
  AOI21_X1 U10185 ( .B1(n9105), .B2(n9219), .A(n9104), .ZN(n9106) );
  OAI222_X1 U10186 ( .A1(n9109), .A2(n9108), .B1(n6896), .B2(P2_U3151), .C1(
        n9107), .C2(n9614), .ZN(P2_U3274) );
  AOI21_X1 U10187 ( .B1(n9110), .B2(n9111), .A(n9224), .ZN(n9113) );
  NAND2_X1 U10188 ( .A1(n9113), .A2(n9112), .ZN(n9118) );
  INV_X1 U10189 ( .A(n9114), .ZN(n9382) );
  AOI22_X1 U10190 ( .A1(n9214), .A2(n5137), .B1(P2_REG3_REG_27__SCAN_IN), .B2(
        P2_U3151), .ZN(n9115) );
  OAI21_X1 U10191 ( .B1(n9403), .B2(n9125), .A(n9115), .ZN(n9116) );
  AOI21_X1 U10192 ( .B1(n9382), .B2(n9234), .A(n9116), .ZN(n9117) );
  OAI211_X1 U10193 ( .C1(n9522), .C2(n9238), .A(n9118), .B(n9117), .ZN(
        P2_U3154) );
  NAND2_X1 U10194 ( .A1(n9119), .A2(n9120), .ZN(n9121) );
  XOR2_X1 U10195 ( .A(n9122), .B(n9121), .Z(n9132) );
  NAND2_X1 U10196 ( .A1(n9214), .A2(n9246), .ZN(n9124) );
  OAI211_X1 U10197 ( .C1(n9126), .C2(n9125), .A(n9124), .B(n9123), .ZN(n9127)
         );
  AOI21_X1 U10198 ( .B1(n9234), .B2(n9128), .A(n9127), .ZN(n9131) );
  NAND2_X1 U10199 ( .A1(n9129), .A2(n9219), .ZN(n9130) );
  OAI211_X1 U10200 ( .C1(n9132), .C2(n9224), .A(n9131), .B(n9130), .ZN(
        P2_U3155) );
  XNOR2_X1 U10201 ( .A(n9133), .B(n9243), .ZN(n9138) );
  AOI22_X1 U10202 ( .A1(n9214), .A2(n9242), .B1(P2_REG3_REG_23__SCAN_IN), .B2(
        P2_U3151), .ZN(n9135) );
  NAND2_X1 U10203 ( .A1(n9229), .A2(n9447), .ZN(n9134) );
  OAI211_X1 U10204 ( .C1(n9217), .C2(n9426), .A(n9135), .B(n9134), .ZN(n9136)
         );
  AOI21_X1 U10205 ( .B1(n9425), .B2(n9219), .A(n9136), .ZN(n9137) );
  OAI21_X1 U10206 ( .B1(n9138), .B2(n9224), .A(n9137), .ZN(P2_U3156) );
  INV_X1 U10207 ( .A(n9554), .ZN(n9150) );
  OR2_X1 U10208 ( .A1(n9139), .A2(n9202), .ZN(n9203) );
  NAND2_X1 U10209 ( .A1(n9203), .A2(n9140), .ZN(n9145) );
  OR2_X1 U10210 ( .A1(n9139), .A2(n9141), .ZN(n9193) );
  AND2_X1 U10211 ( .A1(n9193), .A2(n9142), .ZN(n9143) );
  OAI211_X1 U10212 ( .C1(n9145), .C2(n9144), .A(n9143), .B(n9158), .ZN(n9149)
         );
  NAND2_X1 U10213 ( .A1(P2_U3151), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n9332) );
  OAI21_X1 U10214 ( .B1(n9231), .B2(n9477), .A(n9332), .ZN(n9147) );
  NOR2_X1 U10215 ( .A1(n9217), .A2(n9480), .ZN(n9146) );
  AOI211_X1 U10216 ( .C1(n9229), .C2(n9244), .A(n9147), .B(n9146), .ZN(n9148)
         );
  OAI211_X1 U10217 ( .C1(n9150), .C2(n9238), .A(n9149), .B(n9148), .ZN(
        P2_U3159) );
  XOR2_X1 U10218 ( .A(n9152), .B(n9151), .Z(n9157) );
  AOI22_X1 U10219 ( .A1(n9214), .A2(n9377), .B1(P2_REG3_REG_25__SCAN_IN), .B2(
        P2_U3151), .ZN(n9154) );
  NAND2_X1 U10220 ( .A1(n9229), .A2(n9242), .ZN(n9153) );
  OAI211_X1 U10221 ( .C1(n9217), .C2(n9406), .A(n9154), .B(n9153), .ZN(n9155)
         );
  AOI21_X1 U10222 ( .B1(n9529), .B2(n9219), .A(n9155), .ZN(n9156) );
  OAI21_X1 U10223 ( .B1(n9157), .B2(n9224), .A(n9156), .ZN(P2_U3165) );
  OAI211_X1 U10224 ( .C1(n9161), .C2(n9160), .A(n9159), .B(n9158), .ZN(n9168)
         );
  INV_X1 U10225 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n9162) );
  NOR2_X1 U10226 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9162), .ZN(n9293) );
  AOI21_X1 U10227 ( .B1(n9229), .B2(n9246), .A(n9293), .ZN(n9163) );
  OAI21_X1 U10228 ( .B1(n9164), .B2(n9231), .A(n9163), .ZN(n9165) );
  AOI21_X1 U10229 ( .B1(n9166), .B2(n9234), .A(n9165), .ZN(n9167) );
  OAI211_X1 U10230 ( .C1(n9169), .C2(n9238), .A(n9168), .B(n9167), .ZN(
        P2_U3166) );
  INV_X1 U10231 ( .A(n9170), .ZN(n9171) );
  AOI21_X1 U10232 ( .B1(n9173), .B2(n9172), .A(n9171), .ZN(n9180) );
  NAND2_X1 U10233 ( .A1(n9234), .A2(n9174), .ZN(n9176) );
  AOI22_X1 U10234 ( .A1(n9229), .A2(n9245), .B1(P2_REG3_REG_17__SCAN_IN), .B2(
        P2_U3151), .ZN(n9175) );
  OAI211_X1 U10235 ( .C1(n9475), .C2(n9231), .A(n9176), .B(n9175), .ZN(n9177)
         );
  AOI21_X1 U10236 ( .B1(n9178), .B2(n9219), .A(n9177), .ZN(n9179) );
  OAI21_X1 U10237 ( .B1(n9180), .B2(n9224), .A(n9179), .ZN(P2_U3168) );
  NAND2_X1 U10238 ( .A1(n9181), .A2(n9182), .ZN(n9183) );
  XOR2_X1 U10239 ( .A(n9184), .B(n9183), .Z(n9190) );
  AOI22_X1 U10240 ( .A1(n9214), .A2(n9389), .B1(P2_REG3_REG_24__SCAN_IN), .B2(
        P2_U3151), .ZN(n9186) );
  NAND2_X1 U10241 ( .A1(n9229), .A2(n9243), .ZN(n9185) );
  OAI211_X1 U10242 ( .C1(n9217), .C2(n9413), .A(n9186), .B(n9185), .ZN(n9187)
         );
  AOI21_X1 U10243 ( .B1(n9188), .B2(n9219), .A(n9187), .ZN(n9189) );
  OAI21_X1 U10244 ( .B1(n9190), .B2(n9224), .A(n9189), .ZN(P2_U3169) );
  NAND2_X1 U10245 ( .A1(n9193), .A2(n9191), .ZN(n9195) );
  AND2_X1 U10246 ( .A1(n9193), .A2(n9192), .ZN(n9194) );
  AOI21_X1 U10247 ( .B1(n9196), .B2(n9195), .A(n9194), .ZN(n9201) );
  OAI22_X1 U10248 ( .A1(n9231), .A2(n9436), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9914), .ZN(n9197) );
  AOI21_X1 U10249 ( .B1(n9229), .B2(n9494), .A(n9197), .ZN(n9198) );
  OAI21_X1 U10250 ( .B1(n9217), .B2(n9463), .A(n9198), .ZN(n9199) );
  AOI21_X1 U10251 ( .B1(n9549), .B2(n9219), .A(n9199), .ZN(n9200) );
  OAI21_X1 U10252 ( .B1(n9201), .B2(n9224), .A(n9200), .ZN(P2_U3173) );
  INV_X1 U10253 ( .A(n9508), .ZN(n9608) );
  AOI21_X1 U10254 ( .B1(n9139), .B2(n9202), .A(n9224), .ZN(n9204) );
  NAND2_X1 U10255 ( .A1(n9204), .A2(n9203), .ZN(n9211) );
  INV_X1 U10256 ( .A(n9498), .ZN(n9209) );
  NOR2_X1 U10257 ( .A1(n9205), .A2(P2_STATE_REG_SCAN_IN), .ZN(n10964) );
  AOI21_X1 U10258 ( .B1(n9229), .B2(n9493), .A(n10964), .ZN(n9206) );
  OAI21_X1 U10259 ( .B1(n9207), .B2(n9231), .A(n9206), .ZN(n9208) );
  AOI21_X1 U10260 ( .B1(n9209), .B2(n9234), .A(n9208), .ZN(n9210) );
  OAI211_X1 U10261 ( .C1(n9608), .C2(n9238), .A(n9211), .B(n9210), .ZN(
        P2_U3178) );
  XOR2_X1 U10262 ( .A(n9213), .B(n9212), .Z(n9222) );
  AOI22_X1 U10263 ( .A1(n9229), .A2(n9389), .B1(P2_REG3_REG_26__SCAN_IN), .B2(
        P2_U3151), .ZN(n9216) );
  NAND2_X1 U10264 ( .A1(n9214), .A2(n9390), .ZN(n9215) );
  OAI211_X1 U10265 ( .C1(n9217), .C2(n9394), .A(n9216), .B(n9215), .ZN(n9218)
         );
  AOI21_X1 U10266 ( .B1(n9220), .B2(n9219), .A(n9218), .ZN(n9221) );
  OAI21_X1 U10267 ( .B1(n9222), .B2(n9224), .A(n9221), .ZN(P2_U3180) );
  AOI21_X1 U10268 ( .B1(n9223), .B2(n9225), .A(n9224), .ZN(n9227) );
  NAND2_X1 U10269 ( .A1(n9227), .A2(n9226), .ZN(n9237) );
  NOR2_X1 U10270 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9228), .ZN(n9271) );
  AOI21_X1 U10271 ( .B1(n9229), .B2(n9247), .A(n9271), .ZN(n9230) );
  OAI21_X1 U10272 ( .B1(n9232), .B2(n9231), .A(n9230), .ZN(n9233) );
  AOI21_X1 U10273 ( .B1(n9235), .B2(n9234), .A(n9233), .ZN(n9236) );
  OAI211_X1 U10274 ( .C1(n9239), .C2(n9238), .A(n9237), .B(n9236), .ZN(
        P2_U3181) );
  MUX2_X1 U10275 ( .A(n9349), .B(P2_DATAO_REG_31__SCAN_IN), .S(n10977), .Z(
        P2_U3522) );
  MUX2_X1 U10276 ( .A(n9240), .B(P2_DATAO_REG_30__SCAN_IN), .S(n10977), .Z(
        P2_U3521) );
  MUX2_X1 U10277 ( .A(n9241), .B(P2_DATAO_REG_29__SCAN_IN), .S(n10977), .Z(
        P2_U3520) );
  MUX2_X1 U10278 ( .A(n5137), .B(P2_DATAO_REG_28__SCAN_IN), .S(n10977), .Z(
        P2_U3519) );
  MUX2_X1 U10279 ( .A(n9390), .B(P2_DATAO_REG_27__SCAN_IN), .S(n10977), .Z(
        P2_U3518) );
  MUX2_X1 U10280 ( .A(n9377), .B(P2_DATAO_REG_26__SCAN_IN), .S(n10977), .Z(
        P2_U3517) );
  MUX2_X1 U10281 ( .A(n9389), .B(P2_DATAO_REG_25__SCAN_IN), .S(n10977), .Z(
        P2_U3516) );
  MUX2_X1 U10282 ( .A(n9242), .B(P2_DATAO_REG_24__SCAN_IN), .S(n10977), .Z(
        P2_U3515) );
  MUX2_X1 U10283 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(n9243), .S(P2_U3893), .Z(
        P2_U3514) );
  MUX2_X1 U10284 ( .A(n9447), .B(P2_DATAO_REG_22__SCAN_IN), .S(n10977), .Z(
        P2_U3513) );
  MUX2_X1 U10285 ( .A(n9461), .B(P2_DATAO_REG_21__SCAN_IN), .S(n10977), .Z(
        P2_U3512) );
  MUX2_X1 U10286 ( .A(n9448), .B(P2_DATAO_REG_20__SCAN_IN), .S(n10977), .Z(
        P2_U3511) );
  MUX2_X1 U10287 ( .A(n9494), .B(P2_DATAO_REG_19__SCAN_IN), .S(n10977), .Z(
        P2_U3510) );
  MUX2_X1 U10288 ( .A(n9244), .B(P2_DATAO_REG_18__SCAN_IN), .S(n10977), .Z(
        P2_U3509) );
  MUX2_X1 U10289 ( .A(n9493), .B(P2_DATAO_REG_17__SCAN_IN), .S(n10977), .Z(
        P2_U3508) );
  MUX2_X1 U10290 ( .A(n9245), .B(P2_DATAO_REG_16__SCAN_IN), .S(n10977), .Z(
        P2_U3507) );
  MUX2_X1 U10291 ( .A(n9246), .B(P2_DATAO_REG_15__SCAN_IN), .S(n10977), .Z(
        P2_U3506) );
  MUX2_X1 U10292 ( .A(n9247), .B(P2_DATAO_REG_14__SCAN_IN), .S(n10977), .Z(
        P2_U3505) );
  MUX2_X1 U10293 ( .A(n9248), .B(P2_DATAO_REG_13__SCAN_IN), .S(n10977), .Z(
        P2_U3504) );
  MUX2_X1 U10294 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(n9249), .S(P2_U3893), .Z(
        P2_U3503) );
  MUX2_X1 U10295 ( .A(n9250), .B(P2_DATAO_REG_11__SCAN_IN), .S(n10977), .Z(
        P2_U3502) );
  MUX2_X1 U10296 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(n9251), .S(P2_U3893), .Z(
        P2_U3501) );
  MUX2_X1 U10297 ( .A(n9252), .B(P2_DATAO_REG_9__SCAN_IN), .S(n10977), .Z(
        P2_U3500) );
  MUX2_X1 U10298 ( .A(n9253), .B(P2_DATAO_REG_8__SCAN_IN), .S(n10977), .Z(
        P2_U3499) );
  MUX2_X1 U10299 ( .A(n9254), .B(P2_DATAO_REG_7__SCAN_IN), .S(n10977), .Z(
        P2_U3498) );
  MUX2_X1 U10300 ( .A(n9255), .B(P2_DATAO_REG_6__SCAN_IN), .S(n10977), .Z(
        P2_U3497) );
  MUX2_X1 U10301 ( .A(n9256), .B(P2_DATAO_REG_5__SCAN_IN), .S(n10977), .Z(
        P2_U3496) );
  MUX2_X1 U10302 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(n9257), .S(P2_U3893), .Z(
        P2_U3495) );
  MUX2_X1 U10303 ( .A(n6908), .B(P2_DATAO_REG_3__SCAN_IN), .S(n10977), .Z(
        P2_U3494) );
  MUX2_X1 U10304 ( .A(n9258), .B(P2_DATAO_REG_2__SCAN_IN), .S(n10977), .Z(
        P2_U3493) );
  MUX2_X1 U10305 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(n9259), .S(P2_U3893), .Z(
        P2_U3492) );
  MUX2_X1 U10306 ( .A(n9260), .B(P2_DATAO_REG_0__SCAN_IN), .S(n10977), .Z(
        P2_U3491) );
  NOR2_X2 U10307 ( .A1(n9262), .A2(n6159), .ZN(n9283) );
  AOI21_X1 U10308 ( .B1(n6159), .B2(n9262), .A(n9283), .ZN(n9280) );
  MUX2_X1 U10309 ( .A(P2_REG2_REG_15__SCAN_IN), .B(P2_REG1_REG_15__SCAN_IN), 
        .S(n9324), .Z(n9287) );
  XNOR2_X1 U10310 ( .A(n9298), .B(n9287), .ZN(n9267) );
  OR2_X1 U10311 ( .A1(n9263), .A2(n9269), .ZN(n9265) );
  NAND2_X1 U10312 ( .A1(n9265), .A2(n9264), .ZN(n9266) );
  NAND2_X1 U10313 ( .A1(n9267), .A2(n9266), .ZN(n9288) );
  OAI21_X1 U10314 ( .B1(n9267), .B2(n9266), .A(n9288), .ZN(n9278) );
  XNOR2_X1 U10315 ( .A(n9298), .B(n9297), .ZN(n9270) );
  NOR2_X1 U10316 ( .A1(n8108), .A2(n9270), .ZN(n9299) );
  AOI21_X1 U10317 ( .B1(n9270), .B2(n8108), .A(n9299), .ZN(n9275) );
  INV_X1 U10318 ( .A(n9271), .ZN(n9274) );
  INV_X1 U10319 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n9272) );
  OR2_X1 U10320 ( .A1(n10938), .A2(n9272), .ZN(n9273) );
  OAI211_X1 U10321 ( .C1(n10974), .C2(n9275), .A(n9274), .B(n9273), .ZN(n9277)
         );
  NOR2_X1 U10322 ( .A1(n10976), .A2(n9286), .ZN(n9276) );
  AOI211_X1 U10323 ( .C1(n10962), .C2(n9278), .A(n9277), .B(n9276), .ZN(n9279)
         );
  OAI21_X1 U10324 ( .B1(n9280), .B2(n10969), .A(n9279), .ZN(P2_U3197) );
  NOR2_X1 U10325 ( .A1(n9298), .A2(n9281), .ZN(n9282) );
  AOI22_X1 U10326 ( .A1(n9307), .A2(P2_REG1_REG_16__SCAN_IN), .B1(n6177), .B2(
        n9336), .ZN(n9284) );
  AOI21_X1 U10327 ( .B1(n9285), .B2(n9284), .A(n5166), .ZN(n9309) );
  INV_X1 U10328 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n9296) );
  MUX2_X1 U10329 ( .A(P2_REG2_REG_16__SCAN_IN), .B(P2_REG1_REG_16__SCAN_IN), 
        .S(n9324), .Z(n9319) );
  XNOR2_X1 U10330 ( .A(n9307), .B(n9319), .ZN(n9291) );
  OR2_X1 U10331 ( .A1(n9287), .A2(n9286), .ZN(n9289) );
  NAND2_X1 U10332 ( .A1(n9289), .A2(n9288), .ZN(n9290) );
  NAND2_X1 U10333 ( .A1(n9291), .A2(n9290), .ZN(n9320) );
  OAI21_X1 U10334 ( .B1(n9291), .B2(n9290), .A(n9320), .ZN(n9292) );
  NAND2_X1 U10335 ( .A1(n9292), .A2(n10962), .ZN(n9295) );
  INV_X1 U10336 ( .A(n9293), .ZN(n9294) );
  OAI211_X1 U10337 ( .C1(n9296), .C2(n10938), .A(n9295), .B(n9294), .ZN(n9306)
         );
  NOR2_X1 U10338 ( .A1(n9298), .A2(n9297), .ZN(n9300) );
  MUX2_X1 U10339 ( .A(P2_REG2_REG_16__SCAN_IN), .B(n9301), .S(n9307), .Z(n9302) );
  NOR2_X1 U10340 ( .A1(n9303), .A2(n9302), .ZN(n9335) );
  AOI21_X1 U10341 ( .B1(n9303), .B2(n9302), .A(n9335), .ZN(n9304) );
  NOR2_X1 U10342 ( .A1(n9304), .A2(n10974), .ZN(n9305) );
  AOI211_X1 U10343 ( .C1(n10941), .C2(n9307), .A(n9306), .B(n9305), .ZN(n9308)
         );
  OAI21_X1 U10344 ( .B1(n9309), .B2(n10969), .A(n9308), .ZN(P2_U3198) );
  NOR2_X1 U10345 ( .A1(n10940), .A2(n9310), .ZN(n9311) );
  NOR2_X1 U10346 ( .A1(n9317), .A2(n10949), .ZN(n10948) );
  NOR2_X1 U10347 ( .A1(n9311), .A2(n10948), .ZN(n10968) );
  NAND2_X1 U10348 ( .A1(n10961), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n9312) );
  OAI21_X1 U10349 ( .B1(n10961), .B2(P2_REG1_REG_18__SCAN_IN), .A(n9312), .ZN(
        n10967) );
  NOR2_X1 U10350 ( .A1(n10968), .A2(n10967), .ZN(n10966) );
  INV_X1 U10351 ( .A(n9312), .ZN(n9313) );
  NOR2_X1 U10352 ( .A1(n10966), .A2(n9313), .ZN(n9316) );
  XNOR2_X1 U10353 ( .A(n9327), .B(n9314), .ZN(n9329) );
  INV_X1 U10354 ( .A(n9329), .ZN(n9315) );
  XNOR2_X1 U10355 ( .A(n9316), .B(n9315), .ZN(n9345) );
  MUX2_X1 U10356 ( .A(n9318), .B(n9317), .S(n9324), .Z(n9323) );
  XOR2_X1 U10357 ( .A(n9323), .B(n10940), .Z(n10944) );
  OR2_X1 U10358 ( .A1(n9319), .A2(n9336), .ZN(n9321) );
  NAND2_X1 U10359 ( .A1(n9321), .A2(n9320), .ZN(n10943) );
  NAND2_X1 U10360 ( .A1(n10944), .A2(n10943), .ZN(n10942) );
  INV_X1 U10361 ( .A(n10942), .ZN(n9322) );
  AOI21_X1 U10362 ( .B1(n10940), .B2(n9323), .A(n9322), .ZN(n9326) );
  MUX2_X1 U10363 ( .A(P2_REG2_REG_18__SCAN_IN), .B(P2_REG1_REG_18__SCAN_IN), 
        .S(n9324), .Z(n9325) );
  NOR2_X1 U10364 ( .A1(n9326), .A2(n9325), .ZN(n10958) );
  NAND2_X1 U10365 ( .A1(n9326), .A2(n9325), .ZN(n10959) );
  OAI21_X1 U10366 ( .B1(n10958), .B2(n10979), .A(n10959), .ZN(n9331) );
  MUX2_X1 U10367 ( .A(P2_REG2_REG_19__SCAN_IN), .B(n9481), .S(n9327), .Z(n9342) );
  MUX2_X1 U10368 ( .A(n9329), .B(n9342), .S(n9328), .Z(n9330) );
  XNOR2_X1 U10369 ( .A(n9331), .B(n9330), .ZN(n9344) );
  NAND2_X1 U10370 ( .A1(n10965), .A2(P2_ADDR_REG_19__SCAN_IN), .ZN(n9333) );
  OAI211_X1 U10371 ( .C1(n10976), .C2(n9334), .A(n9333), .B(n9332), .ZN(n9343)
         );
  NOR2_X1 U10372 ( .A1(n10940), .A2(n9337), .ZN(n9338) );
  NAND2_X1 U10373 ( .A1(n10961), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n9339) );
  OAI21_X1 U10374 ( .B1(n10961), .B2(P2_REG2_REG_18__SCAN_IN), .A(n9339), .ZN(
        n10973) );
  INV_X1 U10375 ( .A(n9339), .ZN(n9340) );
  INV_X1 U10376 ( .A(n9347), .ZN(n9348) );
  NAND2_X1 U10377 ( .A1(n9439), .A2(n9348), .ZN(n9356) );
  NAND2_X1 U10378 ( .A1(n9350), .A2(n9349), .ZN(n9573) );
  NAND3_X1 U10379 ( .A1(n9356), .A2(n11111), .A3(n9573), .ZN(n9352) );
  OAI21_X1 U10380 ( .B1(n9500), .B2(P2_REG2_REG_31__SCAN_IN), .A(n9352), .ZN(
        n9351) );
  OAI21_X1 U10381 ( .B1(n9575), .B2(n9441), .A(n9351), .ZN(P2_U3202) );
  OAI21_X1 U10382 ( .B1(n11111), .B2(P2_REG2_REG_30__SCAN_IN), .A(n9352), .ZN(
        n9353) );
  OAI21_X1 U10383 ( .B1(n9578), .B2(n9441), .A(n9353), .ZN(P2_U3203) );
  NAND2_X1 U10384 ( .A1(n9488), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n9355) );
  OAI211_X1 U10385 ( .C1(n9357), .C2(n9441), .A(n9356), .B(n9355), .ZN(n9358)
         );
  AOI21_X1 U10386 ( .B1(n9354), .B2(n9443), .A(n9358), .ZN(n9359) );
  OAI21_X1 U10387 ( .B1(n5160), .B2(n9488), .A(n9359), .ZN(P2_U3204) );
  XNOR2_X1 U10388 ( .A(n9361), .B(n9360), .ZN(n9367) );
  INV_X1 U10389 ( .A(n9516), .ZN(n9375) );
  XNOR2_X1 U10390 ( .A(n9369), .B(n9368), .ZN(n9514) );
  INV_X1 U10391 ( .A(n9370), .ZN(n9371) );
  AOI22_X1 U10392 ( .A1(n9488), .A2(P2_REG2_REG_28__SCAN_IN), .B1(n9439), .B2(
        n9371), .ZN(n9372) );
  OAI21_X1 U10393 ( .B1(n9582), .B2(n9441), .A(n9372), .ZN(n9373) );
  AOI21_X1 U10394 ( .B1(n9514), .B2(n9443), .A(n9373), .ZN(n9374) );
  OAI21_X1 U10395 ( .B1(n9375), .B2(n9488), .A(n9374), .ZN(P2_U3205) );
  XOR2_X1 U10396 ( .A(n9380), .B(n9376), .Z(n9379) );
  AOI222_X1 U10397 ( .A1(n9490), .A2(n9379), .B1(n5137), .B2(n9495), .C1(n9377), .C2(n9492), .ZN(n9521) );
  XNOR2_X1 U10398 ( .A(n9381), .B(n9380), .ZN(n9519) );
  AOI22_X1 U10399 ( .A1(n9488), .A2(P2_REG2_REG_27__SCAN_IN), .B1(n9439), .B2(
        n9382), .ZN(n9383) );
  OAI21_X1 U10400 ( .B1(n9522), .B2(n9441), .A(n9383), .ZN(n9384) );
  AOI21_X1 U10401 ( .B1(n9519), .B2(n9443), .A(n9384), .ZN(n9385) );
  OAI21_X1 U10402 ( .B1(n9521), .B2(n9488), .A(n9385), .ZN(P2_U3206) );
  XNOR2_X1 U10403 ( .A(n9387), .B(n5373), .ZN(n9388) );
  NAND2_X1 U10404 ( .A1(n9388), .A2(n9490), .ZN(n9392) );
  AOI22_X1 U10405 ( .A1(n9495), .A2(n9390), .B1(n9389), .B2(n9492), .ZN(n9391)
         );
  XNOR2_X1 U10406 ( .A(n9393), .B(n5373), .ZN(n9523) );
  INV_X1 U10407 ( .A(n9394), .ZN(n9395) );
  AOI22_X1 U10408 ( .A1(n9488), .A2(P2_REG2_REG_26__SCAN_IN), .B1(n9439), .B2(
        n9395), .ZN(n9396) );
  OAI21_X1 U10409 ( .B1(n9587), .B2(n9441), .A(n9396), .ZN(n9397) );
  AOI21_X1 U10410 ( .B1(n9523), .B2(n9443), .A(n9397), .ZN(n9398) );
  OAI21_X1 U10411 ( .B1(n9525), .B2(n9488), .A(n9398), .ZN(P2_U3207) );
  XNOR2_X1 U10412 ( .A(n9399), .B(n9400), .ZN(n9531) );
  XNOR2_X1 U10413 ( .A(n9401), .B(n9400), .ZN(n9402) );
  OAI222_X1 U10414 ( .A1(n9474), .A2(n9422), .B1(n9476), .B2(n9403), .C1(n9402), .C2(n9471), .ZN(n9528) );
  INV_X1 U10415 ( .A(n9529), .ZN(n9404) );
  NOR2_X1 U10416 ( .A1(n9404), .A2(n11105), .ZN(n9405) );
  OAI21_X1 U10417 ( .B1(n9528), .B2(n9405), .A(n9500), .ZN(n9409) );
  INV_X1 U10418 ( .A(n9406), .ZN(n9407) );
  AOI22_X1 U10419 ( .A1(n9488), .A2(P2_REG2_REG_25__SCAN_IN), .B1(n9439), .B2(
        n9407), .ZN(n9408) );
  OAI211_X1 U10420 ( .C1(n9531), .C2(n9505), .A(n9409), .B(n9408), .ZN(
        P2_U3208) );
  XNOR2_X1 U10421 ( .A(n9410), .B(n9416), .ZN(n9411) );
  OAI222_X1 U10422 ( .A1(n9474), .A2(n9435), .B1(n9476), .B2(n9412), .C1(n9411), .C2(n9471), .ZN(n9532) );
  OAI22_X1 U10423 ( .A1(n9592), .A2(n11105), .B1(n9413), .B2(n11104), .ZN(
        n9414) );
  OAI21_X1 U10424 ( .B1(n9532), .B2(n9414), .A(n9500), .ZN(n9418) );
  XNOR2_X1 U10425 ( .A(n9415), .B(n9416), .ZN(n9533) );
  AOI22_X1 U10426 ( .A1(n9533), .A2(n9443), .B1(P2_REG2_REG_24__SCAN_IN), .B2(
        n9488), .ZN(n9417) );
  NAND2_X1 U10427 ( .A1(n9418), .A2(n9417), .ZN(P2_U3209) );
  XNOR2_X1 U10428 ( .A(n9419), .B(n9424), .ZN(n9420) );
  OAI222_X1 U10429 ( .A1(n9476), .A2(n9422), .B1(n9474), .B2(n9421), .C1(n9420), .C2(n9471), .ZN(n9536) );
  INV_X1 U10430 ( .A(n9536), .ZN(n9431) );
  XNOR2_X1 U10431 ( .A(n9423), .B(n9424), .ZN(n9537) );
  INV_X1 U10432 ( .A(n9425), .ZN(n9596) );
  NOR2_X1 U10433 ( .A1(n9596), .A2(n9441), .ZN(n9429) );
  OAI22_X1 U10434 ( .A1(n9500), .A2(n9427), .B1(n9426), .B2(n11104), .ZN(n9428) );
  AOI211_X1 U10435 ( .C1(n9537), .C2(n9443), .A(n9429), .B(n9428), .ZN(n9430)
         );
  OAI21_X1 U10436 ( .B1(n9431), .B2(n9488), .A(n9430), .ZN(P2_U3210) );
  XNOR2_X1 U10437 ( .A(n9433), .B(n9432), .ZN(n9434) );
  OAI222_X1 U10438 ( .A1(n9474), .A2(n9436), .B1(n9476), .B2(n9435), .C1(n9434), .C2(n9471), .ZN(n9540) );
  INV_X1 U10439 ( .A(n9540), .ZN(n9445) );
  XNOR2_X1 U10440 ( .A(n9437), .B(n5413), .ZN(n9542) );
  AOI22_X1 U10441 ( .A1(n9488), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n9439), .B2(
        n9438), .ZN(n9440) );
  OAI21_X1 U10442 ( .B1(n9600), .B2(n9441), .A(n9440), .ZN(n9442) );
  AOI21_X1 U10443 ( .B1(n9542), .B2(n9443), .A(n9442), .ZN(n9444) );
  OAI21_X1 U10444 ( .B1(n9445), .B2(n9488), .A(n9444), .ZN(P2_U3211) );
  XNOR2_X1 U10445 ( .A(n9446), .B(n5417), .ZN(n9449) );
  AOI222_X1 U10446 ( .A1(n9490), .A2(n9449), .B1(n9448), .B2(n9492), .C1(n9447), .C2(n9495), .ZN(n9547) );
  INV_X1 U10447 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n9451) );
  OAI22_X1 U10448 ( .A1(n9500), .A2(n9451), .B1(n9450), .B2(n11104), .ZN(n9456) );
  OAI21_X1 U10449 ( .B1(n9454), .B2(n9453), .A(n9452), .ZN(n9548) );
  NOR2_X1 U10450 ( .A1(n9548), .A2(n9505), .ZN(n9455) );
  AOI211_X1 U10451 ( .C1(n9509), .C2(n9545), .A(n9456), .B(n9455), .ZN(n9457)
         );
  OAI21_X1 U10452 ( .B1(n9488), .B2(n9547), .A(n9457), .ZN(P2_U3212) );
  OAI21_X1 U10453 ( .B1(n9460), .B2(n9459), .A(n9458), .ZN(n9462) );
  AOI222_X1 U10454 ( .A1(n9490), .A2(n9462), .B1(n9494), .B2(n9492), .C1(n9461), .C2(n9495), .ZN(n9551) );
  OAI22_X1 U10455 ( .A1(n9500), .A2(n9464), .B1(n9463), .B2(n11104), .ZN(n9469) );
  OAI21_X1 U10456 ( .B1(n9467), .B2(n9466), .A(n9465), .ZN(n9552) );
  NOR2_X1 U10457 ( .A1(n9552), .A2(n9505), .ZN(n9468) );
  AOI211_X1 U10458 ( .C1(n9509), .C2(n9549), .A(n9469), .B(n9468), .ZN(n9470)
         );
  OAI21_X1 U10459 ( .B1(n9488), .B2(n9551), .A(n9470), .ZN(P2_U3213) );
  AOI21_X1 U10460 ( .B1(n9472), .B2(n9483), .A(n9471), .ZN(n9479) );
  OAI22_X1 U10461 ( .A1(n9477), .A2(n9476), .B1(n9475), .B2(n9474), .ZN(n9478)
         );
  AOI21_X1 U10462 ( .B1(n9479), .B2(n9473), .A(n9478), .ZN(n9556) );
  OAI22_X1 U10463 ( .A1(n9500), .A2(n9481), .B1(n9480), .B2(n11104), .ZN(n9486) );
  OAI21_X1 U10464 ( .B1(n9484), .B2(n9483), .A(n9482), .ZN(n9557) );
  NOR2_X1 U10465 ( .A1(n9557), .A2(n9505), .ZN(n9485) );
  AOI211_X1 U10466 ( .C1(n9509), .C2(n9554), .A(n9486), .B(n9485), .ZN(n9487)
         );
  OAI21_X1 U10467 ( .B1(n9488), .B2(n9556), .A(n9487), .ZN(P2_U3214) );
  XNOR2_X1 U10468 ( .A(n9489), .B(n5381), .ZN(n9491) );
  NAND2_X1 U10469 ( .A1(n9491), .A2(n9490), .ZN(n9497) );
  AOI22_X1 U10470 ( .A1(n9495), .A2(n9494), .B1(n9493), .B2(n9492), .ZN(n9496)
         );
  INV_X1 U10471 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n9499) );
  OAI22_X1 U10472 ( .A1(n9500), .A2(n9499), .B1(n9498), .B2(n11104), .ZN(n9507) );
  NAND2_X1 U10473 ( .A1(n9502), .A2(n9501), .ZN(n9503) );
  NAND2_X1 U10474 ( .A1(n9504), .A2(n9503), .ZN(n9558) );
  NOR2_X1 U10475 ( .A1(n9558), .A2(n9505), .ZN(n9506) );
  AOI211_X1 U10476 ( .C1(n9509), .C2(n9508), .A(n9507), .B(n9506), .ZN(n9510)
         );
  OAI21_X1 U10477 ( .B1(n9488), .B2(n9559), .A(n9510), .ZN(P2_U3215) );
  NOR2_X1 U10478 ( .A1(n9573), .A2(n9572), .ZN(n9512) );
  AOI21_X1 U10479 ( .B1(P2_REG1_REG_31__SCAN_IN), .B2(n9572), .A(n9512), .ZN(
        n9511) );
  OAI21_X1 U10480 ( .B1(n9575), .B2(n9564), .A(n9511), .ZN(P2_U3490) );
  AOI21_X1 U10481 ( .B1(P2_REG1_REG_30__SCAN_IN), .B2(n9572), .A(n9512), .ZN(
        n9513) );
  OAI21_X1 U10482 ( .B1(n9578), .B2(n9564), .A(n9513), .ZN(P2_U3489) );
  MUX2_X1 U10483 ( .A(n9579), .B(n9517), .S(n9572), .Z(n9518) );
  OAI21_X1 U10484 ( .B1(n9582), .B2(n9564), .A(n9518), .ZN(P2_U3487) );
  NAND2_X1 U10485 ( .A1(n9519), .A2(n9541), .ZN(n9520) );
  OAI211_X1 U10486 ( .C1(n9522), .C2(n9565), .A(n9521), .B(n9520), .ZN(n9583)
         );
  MUX2_X1 U10487 ( .A(n9583), .B(P2_REG1_REG_27__SCAN_IN), .S(n9572), .Z(
        P2_U3486) );
  NAND2_X1 U10488 ( .A1(n9523), .A2(n9541), .ZN(n9524) );
  MUX2_X1 U10489 ( .A(n9526), .B(n9584), .S(n9561), .Z(n9527) );
  OAI21_X1 U10490 ( .B1(n9587), .B2(n9564), .A(n9527), .ZN(P2_U3485) );
  AOI21_X1 U10491 ( .B1(n9553), .B2(n9529), .A(n9528), .ZN(n9530) );
  OAI21_X1 U10492 ( .B1(n9567), .B2(n9531), .A(n9530), .ZN(n9588) );
  MUX2_X1 U10493 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n9588), .S(n9561), .Z(
        P2_U3484) );
  INV_X1 U10494 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n9534) );
  AOI21_X1 U10495 ( .B1(n9541), .B2(n9533), .A(n9532), .ZN(n9589) );
  MUX2_X1 U10496 ( .A(n9534), .B(n9589), .S(n9561), .Z(n9535) );
  OAI21_X1 U10497 ( .B1(n9592), .B2(n9564), .A(n9535), .ZN(P2_U3483) );
  INV_X1 U10498 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n9538) );
  AOI21_X1 U10499 ( .B1(n9541), .B2(n9537), .A(n9536), .ZN(n9593) );
  MUX2_X1 U10500 ( .A(n9538), .B(n9593), .S(n9561), .Z(n9539) );
  OAI21_X1 U10501 ( .B1(n9596), .B2(n9564), .A(n9539), .ZN(P2_U3482) );
  AOI21_X1 U10502 ( .B1(n9542), .B2(n9541), .A(n9540), .ZN(n9597) );
  MUX2_X1 U10503 ( .A(n9543), .B(n9597), .S(n9561), .Z(n9544) );
  OAI21_X1 U10504 ( .B1(n9600), .B2(n9564), .A(n9544), .ZN(P2_U3481) );
  NAND2_X1 U10505 ( .A1(n9545), .A2(n9553), .ZN(n9546) );
  OAI211_X1 U10506 ( .C1(n9567), .C2(n9548), .A(n9547), .B(n9546), .ZN(n9601)
         );
  MUX2_X1 U10507 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n9601), .S(n9561), .Z(
        P2_U3480) );
  NAND2_X1 U10508 ( .A1(n9549), .A2(n9553), .ZN(n9550) );
  OAI211_X1 U10509 ( .C1(n9567), .C2(n9552), .A(n9551), .B(n9550), .ZN(n9602)
         );
  MUX2_X1 U10510 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n9602), .S(n9561), .Z(
        P2_U3479) );
  NAND2_X1 U10511 ( .A1(n9554), .A2(n9553), .ZN(n9555) );
  OAI211_X1 U10512 ( .C1(n9557), .C2(n9567), .A(n9556), .B(n9555), .ZN(n9603)
         );
  MUX2_X1 U10513 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n9603), .S(n9561), .Z(
        P2_U3478) );
  OR2_X1 U10514 ( .A1(n9558), .A2(n9567), .ZN(n9560) );
  MUX2_X1 U10515 ( .A(n9562), .B(n9605), .S(n9561), .Z(n9563) );
  OAI21_X1 U10516 ( .B1(n9608), .B2(n9564), .A(n9563), .ZN(P2_U3477) );
  OAI22_X1 U10517 ( .A1(n9568), .A2(n9567), .B1(n9566), .B2(n9565), .ZN(n9570)
         );
  NOR2_X1 U10518 ( .A1(n9570), .A2(n9569), .ZN(n11177) );
  NAND2_X1 U10519 ( .A1(n9572), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n9571) );
  OAI21_X1 U10520 ( .B1(n11177), .B2(n9572), .A(n9571), .ZN(P2_U3476) );
  NOR2_X1 U10521 ( .A1(n6432), .A2(n9573), .ZN(n9576) );
  AOI21_X1 U10522 ( .B1(n6432), .B2(P2_REG0_REG_31__SCAN_IN), .A(n9576), .ZN(
        n9574) );
  OAI21_X1 U10523 ( .B1(n9575), .B2(n9607), .A(n9574), .ZN(P2_U3458) );
  AOI21_X1 U10524 ( .B1(n6432), .B2(P2_REG0_REG_30__SCAN_IN), .A(n9576), .ZN(
        n9577) );
  OAI21_X1 U10525 ( .B1(n9578), .B2(n9607), .A(n9577), .ZN(P2_U3457) );
  MUX2_X1 U10526 ( .A(n9580), .B(n9579), .S(n11178), .Z(n9581) );
  OAI21_X1 U10527 ( .B1(n9582), .B2(n9607), .A(n9581), .ZN(P2_U3455) );
  MUX2_X1 U10528 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n9583), .S(n11178), .Z(
        P2_U3454) );
  MUX2_X1 U10529 ( .A(n9585), .B(n9584), .S(n11178), .Z(n9586) );
  OAI21_X1 U10530 ( .B1(n9587), .B2(n9607), .A(n9586), .ZN(P2_U3453) );
  MUX2_X1 U10531 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n9588), .S(n11178), .Z(
        P2_U3452) );
  MUX2_X1 U10532 ( .A(n9590), .B(n9589), .S(n11178), .Z(n9591) );
  OAI21_X1 U10533 ( .B1(n9592), .B2(n9607), .A(n9591), .ZN(P2_U3451) );
  MUX2_X1 U10534 ( .A(n9594), .B(n9593), .S(n11178), .Z(n9595) );
  OAI21_X1 U10535 ( .B1(n9596), .B2(n9607), .A(n9595), .ZN(P2_U3450) );
  MUX2_X1 U10536 ( .A(n9598), .B(n9597), .S(n11178), .Z(n9599) );
  OAI21_X1 U10537 ( .B1(n9600), .B2(n9607), .A(n9599), .ZN(P2_U3449) );
  MUX2_X1 U10538 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n9601), .S(n11178), .Z(
        P2_U3448) );
  MUX2_X1 U10539 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n9602), .S(n11178), .Z(
        P2_U3447) );
  MUX2_X1 U10540 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n9603), .S(n11178), .Z(
        P2_U3446) );
  MUX2_X1 U10541 ( .A(n9605), .B(n9604), .S(n6432), .Z(n9606) );
  OAI21_X1 U10542 ( .B1(n9608), .B2(n9607), .A(n9606), .ZN(P2_U3444) );
  MUX2_X1 U10543 ( .A(P2_D_REG_1__SCAN_IN), .B(n9610), .S(n9609), .Z(P2_U3377)
         );
  INV_X1 U10544 ( .A(n9611), .ZN(n10697) );
  NAND3_X1 U10545 ( .A1(n9613), .A2(P2_STATE_REG_SCAN_IN), .A3(
        P2_IR_REG_31__SCAN_IN), .ZN(n9616) );
  OAI22_X1 U10546 ( .A1(n9612), .A2(n9616), .B1(n9615), .B2(n9614), .ZN(n9617)
         );
  INV_X1 U10547 ( .A(n9617), .ZN(n9618) );
  OAI21_X1 U10548 ( .B1(n10697), .B2(n9619), .A(n9618), .ZN(P2_U3264) );
  AOI222_X1 U10549 ( .A1(n9623), .A2(n9622), .B1(P1_DATAO_REG_8__SCAN_IN), 
        .B2(n9621), .C1(P2_STATE_REG_SCAN_IN), .C2(n9620), .ZN(n10039) );
  XNOR2_X1 U10550 ( .A(SI_31_), .B(keyinput_129), .ZN(n9626) );
  XNOR2_X1 U10551 ( .A(P2_WR_REG_SCAN_IN), .B(keyinput_128), .ZN(n9625) );
  XNOR2_X1 U10552 ( .A(SI_30_), .B(keyinput_130), .ZN(n9624) );
  OAI21_X1 U10553 ( .B1(n9626), .B2(n9625), .A(n9624), .ZN(n9630) );
  XNOR2_X1 U10554 ( .A(SI_29_), .B(keyinput_131), .ZN(n9629) );
  XNOR2_X1 U10555 ( .A(SI_28_), .B(keyinput_132), .ZN(n9628) );
  XNOR2_X1 U10556 ( .A(n9825), .B(keyinput_133), .ZN(n9627) );
  AOI211_X1 U10557 ( .C1(n9630), .C2(n9629), .A(n9628), .B(n9627), .ZN(n9633)
         );
  XNOR2_X1 U10558 ( .A(SI_26_), .B(keyinput_134), .ZN(n9632) );
  XNOR2_X1 U10559 ( .A(n9830), .B(keyinput_135), .ZN(n9631) );
  OAI21_X1 U10560 ( .B1(n9633), .B2(n9632), .A(n9631), .ZN(n9640) );
  XNOR2_X1 U10561 ( .A(SI_24_), .B(keyinput_136), .ZN(n9639) );
  XNOR2_X1 U10562 ( .A(n9634), .B(keyinput_139), .ZN(n9637) );
  XNOR2_X1 U10563 ( .A(SI_23_), .B(keyinput_137), .ZN(n9636) );
  XNOR2_X1 U10564 ( .A(SI_22_), .B(keyinput_138), .ZN(n9635) );
  NAND3_X1 U10565 ( .A1(n9637), .A2(n9636), .A3(n9635), .ZN(n9638) );
  AOI21_X1 U10566 ( .B1(n9640), .B2(n9639), .A(n9638), .ZN(n9644) );
  XNOR2_X1 U10567 ( .A(n9641), .B(keyinput_140), .ZN(n9643) );
  XNOR2_X1 U10568 ( .A(n9841), .B(keyinput_141), .ZN(n9642) );
  NOR3_X1 U10569 ( .A1(n9644), .A2(n9643), .A3(n9642), .ZN(n9651) );
  XNOR2_X1 U10570 ( .A(n9845), .B(keyinput_142), .ZN(n9650) );
  XNOR2_X1 U10571 ( .A(n9645), .B(keyinput_144), .ZN(n9648) );
  XNOR2_X1 U10572 ( .A(SI_15_), .B(keyinput_145), .ZN(n9647) );
  XNOR2_X1 U10573 ( .A(SI_17_), .B(keyinput_143), .ZN(n9646) );
  NOR3_X1 U10574 ( .A1(n9648), .A2(n9647), .A3(n9646), .ZN(n9649) );
  OAI21_X1 U10575 ( .B1(n9651), .B2(n9650), .A(n9649), .ZN(n9658) );
  XNOR2_X1 U10576 ( .A(n9853), .B(keyinput_146), .ZN(n9657) );
  XOR2_X1 U10577 ( .A(SI_11_), .B(keyinput_149), .Z(n9655) );
  XNOR2_X1 U10578 ( .A(n9652), .B(keyinput_147), .ZN(n9654) );
  XNOR2_X1 U10579 ( .A(SI_12_), .B(keyinput_148), .ZN(n9653) );
  NAND3_X1 U10580 ( .A1(n9655), .A2(n9654), .A3(n9653), .ZN(n9656) );
  AOI21_X1 U10581 ( .B1(n9658), .B2(n9657), .A(n9656), .ZN(n9661) );
  XNOR2_X1 U10582 ( .A(n9860), .B(keyinput_151), .ZN(n9660) );
  XNOR2_X1 U10583 ( .A(SI_10_), .B(keyinput_150), .ZN(n9659) );
  NOR3_X1 U10584 ( .A1(n9661), .A2(n9660), .A3(n9659), .ZN(n9666) );
  XNOR2_X1 U10585 ( .A(SI_8_), .B(keyinput_152), .ZN(n9665) );
  XNOR2_X1 U10586 ( .A(n9662), .B(keyinput_153), .ZN(n9664) );
  XNOR2_X1 U10587 ( .A(SI_6_), .B(keyinput_154), .ZN(n9663) );
  OAI211_X1 U10588 ( .C1(n9666), .C2(n9665), .A(n9664), .B(n9663), .ZN(n9670)
         );
  XNOR2_X1 U10589 ( .A(n9868), .B(keyinput_155), .ZN(n9669) );
  XNOR2_X1 U10590 ( .A(n9667), .B(keyinput_156), .ZN(n9668) );
  AOI21_X1 U10591 ( .B1(n9670), .B2(n9669), .A(n9668), .ZN(n9673) );
  XNOR2_X1 U10592 ( .A(SI_3_), .B(keyinput_157), .ZN(n9672) );
  XNOR2_X1 U10593 ( .A(SI_2_), .B(keyinput_158), .ZN(n9671) );
  NOR3_X1 U10594 ( .A1(n9673), .A2(n9672), .A3(n9671), .ZN(n9676) );
  XNOR2_X1 U10595 ( .A(SI_1_), .B(keyinput_159), .ZN(n9675) );
  XNOR2_X1 U10596 ( .A(SI_0_), .B(keyinput_160), .ZN(n9674) );
  NOR3_X1 U10597 ( .A1(n9676), .A2(n9675), .A3(n9674), .ZN(n9679) );
  XNOR2_X1 U10598 ( .A(n5287), .B(keyinput_161), .ZN(n9678) );
  XNOR2_X1 U10599 ( .A(P2_STATE_REG_SCAN_IN), .B(keyinput_162), .ZN(n9677) );
  OAI21_X1 U10600 ( .B1(n9679), .B2(n9678), .A(n9677), .ZN(n9682) );
  XOR2_X1 U10601 ( .A(P2_REG3_REG_27__SCAN_IN), .B(keyinput_164), .Z(n9681) );
  XNOR2_X1 U10602 ( .A(P2_REG3_REG_7__SCAN_IN), .B(keyinput_163), .ZN(n9680)
         );
  NAND3_X1 U10603 ( .A1(n9682), .A2(n9681), .A3(n9680), .ZN(n9685) );
  XNOR2_X1 U10604 ( .A(P2_REG3_REG_14__SCAN_IN), .B(keyinput_165), .ZN(n9684)
         );
  XNOR2_X1 U10605 ( .A(P2_REG3_REG_23__SCAN_IN), .B(keyinput_166), .ZN(n9683)
         );
  AOI21_X1 U10606 ( .B1(n9685), .B2(n9684), .A(n9683), .ZN(n9691) );
  XNOR2_X1 U10607 ( .A(P2_REG3_REG_10__SCAN_IN), .B(keyinput_167), .ZN(n9690)
         );
  XNOR2_X1 U10608 ( .A(n9889), .B(keyinput_169), .ZN(n9688) );
  XNOR2_X1 U10609 ( .A(P2_REG3_REG_3__SCAN_IN), .B(keyinput_168), .ZN(n9687)
         );
  XNOR2_X1 U10610 ( .A(P2_REG3_REG_28__SCAN_IN), .B(keyinput_170), .ZN(n9686)
         );
  NOR3_X1 U10611 ( .A1(n9688), .A2(n9687), .A3(n9686), .ZN(n9689) );
  OAI21_X1 U10612 ( .B1(n9691), .B2(n9690), .A(n9689), .ZN(n9694) );
  XNOR2_X1 U10613 ( .A(n9896), .B(keyinput_171), .ZN(n9693) );
  XNOR2_X1 U10614 ( .A(P2_REG3_REG_1__SCAN_IN), .B(keyinput_172), .ZN(n9692)
         );
  NAND3_X1 U10615 ( .A1(n9694), .A2(n9693), .A3(n9692), .ZN(n9697) );
  XNOR2_X1 U10616 ( .A(P2_REG3_REG_21__SCAN_IN), .B(keyinput_173), .ZN(n9696)
         );
  XNOR2_X1 U10617 ( .A(P2_REG3_REG_12__SCAN_IN), .B(keyinput_174), .ZN(n9695)
         );
  AOI21_X1 U10618 ( .B1(n9697), .B2(n9696), .A(n9695), .ZN(n9700) );
  XOR2_X1 U10619 ( .A(P2_REG3_REG_16__SCAN_IN), .B(keyinput_176), .Z(n9699) );
  XNOR2_X1 U10620 ( .A(P2_REG3_REG_25__SCAN_IN), .B(keyinput_175), .ZN(n9698)
         );
  NOR3_X1 U10621 ( .A1(n9700), .A2(n9699), .A3(n9698), .ZN(n9709) );
  XNOR2_X1 U10622 ( .A(n9701), .B(keyinput_177), .ZN(n9708) );
  XNOR2_X1 U10623 ( .A(P2_REG3_REG_9__SCAN_IN), .B(keyinput_181), .ZN(n9707)
         );
  XNOR2_X1 U10624 ( .A(P2_REG3_REG_17__SCAN_IN), .B(keyinput_178), .ZN(n9705)
         );
  XNOR2_X1 U10625 ( .A(P2_REG3_REG_4__SCAN_IN), .B(keyinput_180), .ZN(n9704)
         );
  XNOR2_X1 U10626 ( .A(P2_REG3_REG_24__SCAN_IN), .B(keyinput_179), .ZN(n9703)
         );
  XNOR2_X1 U10627 ( .A(P2_REG3_REG_0__SCAN_IN), .B(keyinput_182), .ZN(n9702)
         );
  NAND4_X1 U10628 ( .A1(n9705), .A2(n9704), .A3(n9703), .A4(n9702), .ZN(n9706)
         );
  NOR4_X1 U10629 ( .A1(n9709), .A2(n9708), .A3(n9707), .A4(n9706), .ZN(n9712)
         );
  XNOR2_X1 U10630 ( .A(n9914), .B(keyinput_183), .ZN(n9711) );
  XNOR2_X1 U10631 ( .A(P2_REG3_REG_13__SCAN_IN), .B(keyinput_184), .ZN(n9710)
         );
  OAI21_X1 U10632 ( .B1(n9712), .B2(n9711), .A(n9710), .ZN(n9717) );
  XOR2_X1 U10633 ( .A(P2_REG3_REG_2__SCAN_IN), .B(keyinput_187), .Z(n9716) );
  OAI22_X1 U10634 ( .A1(P2_REG3_REG_22__SCAN_IN), .A2(keyinput_185), .B1(
        P2_REG3_REG_11__SCAN_IN), .B2(keyinput_186), .ZN(n9713) );
  AOI21_X1 U10635 ( .B1(P2_REG3_REG_22__SCAN_IN), .B2(keyinput_185), .A(n9713), 
        .ZN(n9715) );
  NAND2_X1 U10636 ( .A1(P2_REG3_REG_11__SCAN_IN), .A2(keyinput_186), .ZN(n9714) );
  NAND4_X1 U10637 ( .A1(n9717), .A2(n9716), .A3(n9715), .A4(n9714), .ZN(n9723)
         );
  XNOR2_X1 U10638 ( .A(P2_REG3_REG_6__SCAN_IN), .B(keyinput_189), .ZN(n9720)
         );
  XNOR2_X1 U10639 ( .A(P2_REG3_REG_26__SCAN_IN), .B(keyinput_190), .ZN(n9719)
         );
  XNOR2_X1 U10640 ( .A(P2_REG3_REG_18__SCAN_IN), .B(keyinput_188), .ZN(n9718)
         );
  NOR3_X1 U10641 ( .A1(n9720), .A2(n9719), .A3(n9718), .ZN(n9722) );
  XNOR2_X1 U10642 ( .A(P2_REG3_REG_15__SCAN_IN), .B(keyinput_191), .ZN(n9721)
         );
  AOI21_X1 U10643 ( .B1(n9723), .B2(n9722), .A(n9721), .ZN(n9727) );
  XNOR2_X1 U10644 ( .A(P2_B_REG_SCAN_IN), .B(keyinput_192), .ZN(n9726) );
  XNOR2_X1 U10645 ( .A(n9933), .B(keyinput_194), .ZN(n9725) );
  XNOR2_X1 U10646 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(keyinput_193), .ZN(n9724)
         );
  OAI211_X1 U10647 ( .C1(n9727), .C2(n9726), .A(n9725), .B(n9724), .ZN(n9730)
         );
  XNOR2_X1 U10648 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(keyinput_195), .ZN(n9729)
         );
  XNOR2_X1 U10649 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(keyinput_196), .ZN(n9728)
         );
  NAND3_X1 U10650 ( .A1(n9730), .A2(n9729), .A3(n9728), .ZN(n9736) );
  OAI22_X1 U10651 ( .A1(n9942), .A2(keyinput_197), .B1(n9732), .B2(
        keyinput_198), .ZN(n9731) );
  AOI21_X1 U10652 ( .B1(n9942), .B2(keyinput_197), .A(n9731), .ZN(n9735) );
  XNOR2_X1 U10653 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(keyinput_199), .ZN(n9734)
         );
  NAND2_X1 U10654 ( .A1(n9732), .A2(keyinput_198), .ZN(n9733) );
  NAND4_X1 U10655 ( .A1(n9736), .A2(n9735), .A3(n9734), .A4(n9733), .ZN(n9740)
         );
  XNOR2_X1 U10656 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(keyinput_200), .ZN(n9739)
         );
  XOR2_X1 U10657 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(keyinput_201), .Z(n9738)
         );
  XNOR2_X1 U10658 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(keyinput_202), .ZN(n9737)
         );
  AOI211_X1 U10659 ( .C1(n9740), .C2(n9739), .A(n9738), .B(n9737), .ZN(n9743)
         );
  XOR2_X1 U10660 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(keyinput_203), .Z(n9742)
         );
  XOR2_X1 U10661 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(keyinput_204), .Z(n9741)
         );
  OAI21_X1 U10662 ( .B1(n9743), .B2(n9742), .A(n9741), .ZN(n9749) );
  XOR2_X1 U10663 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(keyinput_206), .Z(n9745)
         );
  XNOR2_X1 U10664 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(keyinput_205), .ZN(n9744)
         );
  NOR2_X1 U10665 ( .A1(n9745), .A2(n9744), .ZN(n9748) );
  XOR2_X1 U10666 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(keyinput_207), .Z(n9747)
         );
  XNOR2_X1 U10667 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(keyinput_208), .ZN(n9746)
         );
  AOI211_X1 U10668 ( .C1(n9749), .C2(n9748), .A(n9747), .B(n9746), .ZN(n9752)
         );
  XNOR2_X1 U10669 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(keyinput_209), .ZN(n9751)
         );
  XOR2_X1 U10670 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(keyinput_210), .Z(n9750)
         );
  OAI21_X1 U10671 ( .B1(n9752), .B2(n9751), .A(n9750), .ZN(n9756) );
  XOR2_X1 U10672 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(keyinput_211), .Z(n9755)
         );
  XNOR2_X1 U10673 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(keyinput_213), .ZN(n9754)
         );
  XNOR2_X1 U10674 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(keyinput_212), .ZN(n9753)
         );
  AOI211_X1 U10675 ( .C1(n9756), .C2(n9755), .A(n9754), .B(n9753), .ZN(n9759)
         );
  XOR2_X1 U10676 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(keyinput_214), .Z(n9758)
         );
  XOR2_X1 U10677 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(keyinput_215), .Z(n9757) );
  NOR3_X1 U10678 ( .A1(n9759), .A2(n9758), .A3(n9757), .ZN(n9768) );
  XOR2_X1 U10679 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(keyinput_216), .Z(n9763) );
  XNOR2_X1 U10680 ( .A(P1_IR_REG_0__SCAN_IN), .B(keyinput_218), .ZN(n9762) );
  XNOR2_X1 U10681 ( .A(P1_IR_REG_1__SCAN_IN), .B(keyinput_219), .ZN(n9761) );
  XNOR2_X1 U10682 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(keyinput_217), .ZN(n9760)
         );
  NAND4_X1 U10683 ( .A1(n9763), .A2(n9762), .A3(n9761), .A4(n9760), .ZN(n9767)
         );
  XNOR2_X1 U10684 ( .A(n9764), .B(keyinput_220), .ZN(n9766) );
  XNOR2_X1 U10685 ( .A(n9974), .B(keyinput_221), .ZN(n9765) );
  OAI211_X1 U10686 ( .C1(n9768), .C2(n9767), .A(n9766), .B(n9765), .ZN(n9771)
         );
  XNOR2_X1 U10687 ( .A(P1_IR_REG_4__SCAN_IN), .B(keyinput_222), .ZN(n9770) );
  XNOR2_X1 U10688 ( .A(P1_IR_REG_5__SCAN_IN), .B(keyinput_223), .ZN(n9769) );
  AOI21_X1 U10689 ( .B1(n9771), .B2(n9770), .A(n9769), .ZN(n9776) );
  XOR2_X1 U10690 ( .A(P1_IR_REG_7__SCAN_IN), .B(keyinput_225), .Z(n9775) );
  XNOR2_X1 U10691 ( .A(n9772), .B(keyinput_224), .ZN(n9774) );
  XNOR2_X1 U10692 ( .A(P1_IR_REG_8__SCAN_IN), .B(keyinput_226), .ZN(n9773) );
  NOR4_X1 U10693 ( .A1(n9776), .A2(n9775), .A3(n9774), .A4(n9773), .ZN(n9779)
         );
  XNOR2_X1 U10694 ( .A(n9986), .B(keyinput_227), .ZN(n9778) );
  XNOR2_X1 U10695 ( .A(P1_IR_REG_10__SCAN_IN), .B(keyinput_228), .ZN(n9777) );
  OAI21_X1 U10696 ( .B1(n9779), .B2(n9778), .A(n9777), .ZN(n9786) );
  XNOR2_X1 U10697 ( .A(n9780), .B(keyinput_231), .ZN(n9785) );
  XNOR2_X1 U10698 ( .A(n9781), .B(keyinput_230), .ZN(n9784) );
  XNOR2_X1 U10699 ( .A(n9782), .B(keyinput_229), .ZN(n9783) );
  NAND4_X1 U10700 ( .A1(n9786), .A2(n9785), .A3(n9784), .A4(n9783), .ZN(n9790)
         );
  XNOR2_X1 U10701 ( .A(P1_IR_REG_14__SCAN_IN), .B(keyinput_232), .ZN(n9789) );
  XNOR2_X1 U10702 ( .A(n9787), .B(keyinput_233), .ZN(n9788) );
  AOI21_X1 U10703 ( .B1(n9790), .B2(n9789), .A(n9788), .ZN(n9795) );
  XNOR2_X1 U10704 ( .A(P1_IR_REG_16__SCAN_IN), .B(keyinput_234), .ZN(n9794) );
  XNOR2_X1 U10705 ( .A(n9791), .B(keyinput_235), .ZN(n9793) );
  XNOR2_X1 U10706 ( .A(P1_IR_REG_18__SCAN_IN), .B(keyinput_236), .ZN(n9792) );
  OAI211_X1 U10707 ( .C1(n9795), .C2(n9794), .A(n9793), .B(n9792), .ZN(n9799)
         );
  XNOR2_X1 U10708 ( .A(n9796), .B(keyinput_238), .ZN(n9798) );
  XNOR2_X1 U10709 ( .A(P1_IR_REG_19__SCAN_IN), .B(keyinput_237), .ZN(n9797) );
  NAND3_X1 U10710 ( .A1(n9799), .A2(n9798), .A3(n9797), .ZN(n9803) );
  XNOR2_X1 U10711 ( .A(P1_IR_REG_21__SCAN_IN), .B(keyinput_239), .ZN(n9802) );
  XNOR2_X1 U10712 ( .A(n10008), .B(keyinput_241), .ZN(n9801) );
  XNOR2_X1 U10713 ( .A(P1_IR_REG_22__SCAN_IN), .B(keyinput_240), .ZN(n9800) );
  AOI211_X1 U10714 ( .C1(n9803), .C2(n9802), .A(n9801), .B(n9800), .ZN(n9807)
         );
  XNOR2_X1 U10715 ( .A(P1_IR_REG_26__SCAN_IN), .B(keyinput_244), .ZN(n9806) );
  XNOR2_X1 U10716 ( .A(P1_IR_REG_24__SCAN_IN), .B(keyinput_242), .ZN(n9805) );
  XNOR2_X1 U10717 ( .A(P1_IR_REG_25__SCAN_IN), .B(keyinput_243), .ZN(n9804) );
  NOR4_X1 U10718 ( .A1(n9807), .A2(n9806), .A3(n9805), .A4(n9804), .ZN(n9810)
         );
  XNOR2_X1 U10719 ( .A(n10018), .B(keyinput_245), .ZN(n9809) );
  XOR2_X1 U10720 ( .A(P1_IR_REG_28__SCAN_IN), .B(keyinput_246), .Z(n9808) );
  OAI21_X1 U10721 ( .B1(n9810), .B2(n9809), .A(n9808), .ZN(n9814) );
  XOR2_X1 U10722 ( .A(P1_IR_REG_29__SCAN_IN), .B(keyinput_247), .Z(n9813) );
  XNOR2_X1 U10723 ( .A(P1_IR_REG_30__SCAN_IN), .B(keyinput_248), .ZN(n9812) );
  XNOR2_X1 U10724 ( .A(P1_IR_REG_31__SCAN_IN), .B(keyinput_249), .ZN(n9811) );
  AOI211_X1 U10725 ( .C1(n9814), .C2(n9813), .A(n9812), .B(n9811), .ZN(n9817)
         );
  XNOR2_X1 U10726 ( .A(P1_D_REG_0__SCAN_IN), .B(keyinput_250), .ZN(n9816) );
  XOR2_X1 U10727 ( .A(P1_D_REG_1__SCAN_IN), .B(keyinput_251), .Z(n9815) );
  OAI21_X1 U10728 ( .B1(n9817), .B2(n9816), .A(n9815), .ZN(n9821) );
  XNOR2_X1 U10729 ( .A(P1_D_REG_2__SCAN_IN), .B(keyinput_252), .ZN(n9820) );
  INV_X1 U10730 ( .A(P1_D_REG_4__SCAN_IN), .ZN(n10710) );
  XNOR2_X1 U10731 ( .A(n10710), .B(keyinput_254), .ZN(n9819) );
  INV_X1 U10732 ( .A(P1_D_REG_3__SCAN_IN), .ZN(n10709) );
  XNOR2_X1 U10733 ( .A(n10709), .B(keyinput_253), .ZN(n9818) );
  AOI211_X1 U10734 ( .C1(n9821), .C2(n9820), .A(n9819), .B(n9818), .ZN(n10037)
         );
  XNOR2_X1 U10735 ( .A(P1_D_REG_5__SCAN_IN), .B(keyinput_255), .ZN(n10036) );
  XOR2_X1 U10736 ( .A(P1_D_REG_5__SCAN_IN), .B(keyinput_127), .Z(n10035) );
  XNOR2_X1 U10737 ( .A(P2_WR_REG_SCAN_IN), .B(keyinput_0), .ZN(n9824) );
  XNOR2_X1 U10738 ( .A(SI_31_), .B(keyinput_1), .ZN(n9823) );
  XNOR2_X1 U10739 ( .A(SI_30_), .B(keyinput_2), .ZN(n9822) );
  OAI21_X1 U10740 ( .B1(n9824), .B2(n9823), .A(n9822), .ZN(n9829) );
  XNOR2_X1 U10741 ( .A(SI_29_), .B(keyinput_3), .ZN(n9828) );
  XNOR2_X1 U10742 ( .A(SI_28_), .B(keyinput_4), .ZN(n9827) );
  XNOR2_X1 U10743 ( .A(n9825), .B(keyinput_5), .ZN(n9826) );
  AOI211_X1 U10744 ( .C1(n9829), .C2(n9828), .A(n9827), .B(n9826), .ZN(n9833)
         );
  XNOR2_X1 U10745 ( .A(SI_26_), .B(keyinput_6), .ZN(n9832) );
  XNOR2_X1 U10746 ( .A(n9830), .B(keyinput_7), .ZN(n9831) );
  OAI21_X1 U10747 ( .B1(n9833), .B2(n9832), .A(n9831), .ZN(n9840) );
  XNOR2_X1 U10748 ( .A(SI_24_), .B(keyinput_8), .ZN(n9839) );
  XNOR2_X1 U10749 ( .A(n9834), .B(keyinput_10), .ZN(n9837) );
  XNOR2_X1 U10750 ( .A(SI_21_), .B(keyinput_11), .ZN(n9836) );
  XNOR2_X1 U10751 ( .A(SI_23_), .B(keyinput_9), .ZN(n9835) );
  NAND3_X1 U10752 ( .A1(n9837), .A2(n9836), .A3(n9835), .ZN(n9838) );
  AOI21_X1 U10753 ( .B1(n9840), .B2(n9839), .A(n9838), .ZN(n9844) );
  XNOR2_X1 U10754 ( .A(n9841), .B(keyinput_13), .ZN(n9843) );
  XNOR2_X1 U10755 ( .A(SI_20_), .B(keyinput_12), .ZN(n9842) );
  NOR3_X1 U10756 ( .A1(n9844), .A2(n9843), .A3(n9842), .ZN(n9852) );
  XNOR2_X1 U10757 ( .A(n9845), .B(keyinput_14), .ZN(n9851) );
  XNOR2_X1 U10758 ( .A(n9846), .B(keyinput_17), .ZN(n9849) );
  XNOR2_X1 U10759 ( .A(SI_17_), .B(keyinput_15), .ZN(n9848) );
  XNOR2_X1 U10760 ( .A(SI_16_), .B(keyinput_16), .ZN(n9847) );
  NOR3_X1 U10761 ( .A1(n9849), .A2(n9848), .A3(n9847), .ZN(n9850) );
  OAI21_X1 U10762 ( .B1(n9852), .B2(n9851), .A(n9850), .ZN(n9859) );
  XNOR2_X1 U10763 ( .A(n9853), .B(keyinput_18), .ZN(n9858) );
  XOR2_X1 U10764 ( .A(SI_12_), .B(keyinput_20), .Z(n9856) );
  XNOR2_X1 U10765 ( .A(SI_11_), .B(keyinput_21), .ZN(n9855) );
  XNOR2_X1 U10766 ( .A(SI_13_), .B(keyinput_19), .ZN(n9854) );
  NAND3_X1 U10767 ( .A1(n9856), .A2(n9855), .A3(n9854), .ZN(n9857) );
  AOI21_X1 U10768 ( .B1(n9859), .B2(n9858), .A(n9857), .ZN(n9863) );
  XNOR2_X1 U10769 ( .A(n9860), .B(keyinput_23), .ZN(n9862) );
  XNOR2_X1 U10770 ( .A(SI_10_), .B(keyinput_22), .ZN(n9861) );
  NOR3_X1 U10771 ( .A1(n9863), .A2(n9862), .A3(n9861), .ZN(n9867) );
  XNOR2_X1 U10772 ( .A(SI_8_), .B(keyinput_24), .ZN(n9866) );
  XNOR2_X1 U10773 ( .A(SI_6_), .B(keyinput_26), .ZN(n9865) );
  XNOR2_X1 U10774 ( .A(SI_7_), .B(keyinput_25), .ZN(n9864) );
  OAI211_X1 U10775 ( .C1(n9867), .C2(n9866), .A(n9865), .B(n9864), .ZN(n9871)
         );
  XNOR2_X1 U10776 ( .A(n9868), .B(keyinput_27), .ZN(n9870) );
  XNOR2_X1 U10777 ( .A(SI_4_), .B(keyinput_28), .ZN(n9869) );
  AOI21_X1 U10778 ( .B1(n9871), .B2(n9870), .A(n9869), .ZN(n9874) );
  XOR2_X1 U10779 ( .A(SI_2_), .B(keyinput_30), .Z(n9873) );
  XNOR2_X1 U10780 ( .A(SI_3_), .B(keyinput_29), .ZN(n9872) );
  NOR3_X1 U10781 ( .A1(n9874), .A2(n9873), .A3(n9872), .ZN(n9877) );
  XOR2_X1 U10782 ( .A(SI_0_), .B(keyinput_32), .Z(n9876) );
  XNOR2_X1 U10783 ( .A(SI_1_), .B(keyinput_31), .ZN(n9875) );
  NOR3_X1 U10784 ( .A1(n9877), .A2(n9876), .A3(n9875), .ZN(n9880) );
  XNOR2_X1 U10785 ( .A(P2_RD_REG_SCAN_IN), .B(keyinput_33), .ZN(n9879) );
  XNOR2_X1 U10786 ( .A(P2_U3151), .B(keyinput_34), .ZN(n9878) );
  OAI21_X1 U10787 ( .B1(n9880), .B2(n9879), .A(n9878), .ZN(n9883) );
  XOR2_X1 U10788 ( .A(P2_REG3_REG_27__SCAN_IN), .B(keyinput_36), .Z(n9882) );
  XNOR2_X1 U10789 ( .A(P2_REG3_REG_7__SCAN_IN), .B(keyinput_35), .ZN(n9881) );
  NAND3_X1 U10790 ( .A1(n9883), .A2(n9882), .A3(n9881), .ZN(n9887) );
  XNOR2_X1 U10791 ( .A(n9884), .B(keyinput_37), .ZN(n9886) );
  XNOR2_X1 U10792 ( .A(P2_REG3_REG_23__SCAN_IN), .B(keyinput_38), .ZN(n9885)
         );
  AOI21_X1 U10793 ( .B1(n9887), .B2(n9886), .A(n9885), .ZN(n9895) );
  XOR2_X1 U10794 ( .A(P2_REG3_REG_10__SCAN_IN), .B(keyinput_39), .Z(n9894) );
  XOR2_X1 U10795 ( .A(P2_REG3_REG_3__SCAN_IN), .B(keyinput_40), .Z(n9892) );
  XNOR2_X1 U10796 ( .A(n9888), .B(keyinput_42), .ZN(n9891) );
  XNOR2_X1 U10797 ( .A(n9889), .B(keyinput_41), .ZN(n9890) );
  NOR3_X1 U10798 ( .A1(n9892), .A2(n9891), .A3(n9890), .ZN(n9893) );
  OAI21_X1 U10799 ( .B1(n9895), .B2(n9894), .A(n9893), .ZN(n9899) );
  XOR2_X1 U10800 ( .A(P2_REG3_REG_1__SCAN_IN), .B(keyinput_44), .Z(n9898) );
  XNOR2_X1 U10801 ( .A(n9896), .B(keyinput_43), .ZN(n9897) );
  NAND3_X1 U10802 ( .A1(n9899), .A2(n9898), .A3(n9897), .ZN(n9902) );
  XOR2_X1 U10803 ( .A(P2_REG3_REG_21__SCAN_IN), .B(keyinput_45), .Z(n9901) );
  XOR2_X1 U10804 ( .A(P2_REG3_REG_12__SCAN_IN), .B(keyinput_46), .Z(n9900) );
  AOI21_X1 U10805 ( .B1(n9902), .B2(n9901), .A(n9900), .ZN(n9905) );
  XOR2_X1 U10806 ( .A(P2_REG3_REG_16__SCAN_IN), .B(keyinput_48), .Z(n9904) );
  XNOR2_X1 U10807 ( .A(P2_REG3_REG_25__SCAN_IN), .B(keyinput_47), .ZN(n9903)
         );
  NOR3_X1 U10808 ( .A1(n9905), .A2(n9904), .A3(n9903), .ZN(n9913) );
  XNOR2_X1 U10809 ( .A(P2_REG3_REG_9__SCAN_IN), .B(keyinput_53), .ZN(n9912) );
  XNOR2_X1 U10810 ( .A(P2_REG3_REG_24__SCAN_IN), .B(keyinput_51), .ZN(n9911)
         );
  XNOR2_X1 U10811 ( .A(P2_REG3_REG_5__SCAN_IN), .B(keyinput_49), .ZN(n9909) );
  XNOR2_X1 U10812 ( .A(P2_REG3_REG_4__SCAN_IN), .B(keyinput_52), .ZN(n9908) );
  XNOR2_X1 U10813 ( .A(P2_REG3_REG_17__SCAN_IN), .B(keyinput_50), .ZN(n9907)
         );
  XNOR2_X1 U10814 ( .A(P2_REG3_REG_0__SCAN_IN), .B(keyinput_54), .ZN(n9906) );
  NAND4_X1 U10815 ( .A1(n9909), .A2(n9908), .A3(n9907), .A4(n9906), .ZN(n9910)
         );
  NOR4_X1 U10816 ( .A1(n9913), .A2(n9912), .A3(n9911), .A4(n9910), .ZN(n9918)
         );
  XNOR2_X1 U10817 ( .A(n9914), .B(keyinput_55), .ZN(n9917) );
  XNOR2_X1 U10818 ( .A(n9915), .B(keyinput_56), .ZN(n9916) );
  OAI21_X1 U10819 ( .B1(n9918), .B2(n9917), .A(n9916), .ZN(n9925) );
  XNOR2_X1 U10820 ( .A(n9919), .B(keyinput_57), .ZN(n9924) );
  INV_X1 U10821 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n9921) );
  OAI22_X1 U10822 ( .A1(n9921), .A2(keyinput_58), .B1(keyinput_59), .B2(
        P2_REG3_REG_2__SCAN_IN), .ZN(n9920) );
  AOI21_X1 U10823 ( .B1(n9921), .B2(keyinput_58), .A(n9920), .ZN(n9923) );
  NAND2_X1 U10824 ( .A1(P2_REG3_REG_2__SCAN_IN), .A2(keyinput_59), .ZN(n9922)
         );
  NAND4_X1 U10825 ( .A1(n9925), .A2(n9924), .A3(n9923), .A4(n9922), .ZN(n9932)
         );
  XOR2_X1 U10826 ( .A(P2_REG3_REG_6__SCAN_IN), .B(keyinput_61), .Z(n9929) );
  XNOR2_X1 U10827 ( .A(n9926), .B(keyinput_62), .ZN(n9928) );
  XNOR2_X1 U10828 ( .A(P2_REG3_REG_18__SCAN_IN), .B(keyinput_60), .ZN(n9927)
         );
  NOR3_X1 U10829 ( .A1(n9929), .A2(n9928), .A3(n9927), .ZN(n9931) );
  XNOR2_X1 U10830 ( .A(P2_REG3_REG_15__SCAN_IN), .B(keyinput_63), .ZN(n9930)
         );
  AOI21_X1 U10831 ( .B1(n9932), .B2(n9931), .A(n9930), .ZN(n9937) );
  XOR2_X1 U10832 ( .A(P2_B_REG_SCAN_IN), .B(keyinput_64), .Z(n9936) );
  XNOR2_X1 U10833 ( .A(n9933), .B(keyinput_66), .ZN(n9935) );
  XNOR2_X1 U10834 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(keyinput_65), .ZN(n9934)
         );
  OAI211_X1 U10835 ( .C1(n9937), .C2(n9936), .A(n9935), .B(n9934), .ZN(n9940)
         );
  XNOR2_X1 U10836 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(keyinput_67), .ZN(n9939)
         );
  XNOR2_X1 U10837 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(keyinput_68), .ZN(n9938)
         );
  NAND3_X1 U10838 ( .A1(n9940), .A2(n9939), .A3(n9938), .ZN(n9946) );
  OAI22_X1 U10839 ( .A1(n9942), .A2(keyinput_69), .B1(P2_DATAO_REG_26__SCAN_IN), .B2(keyinput_70), .ZN(n9941) );
  AOI21_X1 U10840 ( .B1(n9942), .B2(keyinput_69), .A(n9941), .ZN(n9945) );
  XNOR2_X1 U10841 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(keyinput_71), .ZN(n9944)
         );
  NAND2_X1 U10842 ( .A1(P2_DATAO_REG_26__SCAN_IN), .A2(keyinput_70), .ZN(n9943) );
  NAND4_X1 U10843 ( .A1(n9946), .A2(n9945), .A3(n9944), .A4(n9943), .ZN(n9950)
         );
  XOR2_X1 U10844 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(keyinput_72), .Z(n9949) );
  XOR2_X1 U10845 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(keyinput_74), .Z(n9948) );
  XNOR2_X1 U10846 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(keyinput_73), .ZN(n9947)
         );
  AOI211_X1 U10847 ( .C1(n9950), .C2(n9949), .A(n9948), .B(n9947), .ZN(n9953)
         );
  XOR2_X1 U10848 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(keyinput_75), .Z(n9952) );
  XNOR2_X1 U10849 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(keyinput_76), .ZN(n9951)
         );
  OAI21_X1 U10850 ( .B1(n9953), .B2(n9952), .A(n9951), .ZN(n9956) );
  XNOR2_X1 U10851 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(keyinput_77), .ZN(n9955)
         );
  XNOR2_X1 U10852 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(keyinput_78), .ZN(n9954)
         );
  NAND3_X1 U10853 ( .A1(n9956), .A2(n9955), .A3(n9954), .ZN(n9959) );
  XNOR2_X1 U10854 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(keyinput_79), .ZN(n9958)
         );
  XNOR2_X1 U10855 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(keyinput_80), .ZN(n9957)
         );
  NAND3_X1 U10856 ( .A1(n9959), .A2(n9958), .A3(n9957), .ZN(n9962) );
  XOR2_X1 U10857 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(keyinput_81), .Z(n9961) );
  XNOR2_X1 U10858 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(keyinput_82), .ZN(n9960)
         );
  AOI21_X1 U10859 ( .B1(n9962), .B2(n9961), .A(n9960), .ZN(n9966) );
  XNOR2_X1 U10860 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(keyinput_83), .ZN(n9965)
         );
  XNOR2_X1 U10861 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(keyinput_85), .ZN(n9964)
         );
  XNOR2_X1 U10862 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(keyinput_84), .ZN(n9963)
         );
  OAI211_X1 U10863 ( .C1(n9966), .C2(n9965), .A(n9964), .B(n9963), .ZN(n9969)
         );
  XOR2_X1 U10864 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(keyinput_87), .Z(n9968) );
  XNOR2_X1 U10865 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(keyinput_86), .ZN(n9967)
         );
  NAND3_X1 U10866 ( .A1(n9969), .A2(n9968), .A3(n9967), .ZN(n9978) );
  XOR2_X1 U10867 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(keyinput_89), .Z(n9973) );
  XNOR2_X1 U10868 ( .A(P1_IR_REG_1__SCAN_IN), .B(keyinput_91), .ZN(n9972) );
  XNOR2_X1 U10869 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(keyinput_88), .ZN(n9971)
         );
  XNOR2_X1 U10870 ( .A(P1_IR_REG_0__SCAN_IN), .B(keyinput_90), .ZN(n9970) );
  NOR4_X1 U10871 ( .A1(n9973), .A2(n9972), .A3(n9971), .A4(n9970), .ZN(n9977)
         );
  XNOR2_X1 U10872 ( .A(n9974), .B(keyinput_93), .ZN(n9976) );
  XNOR2_X1 U10873 ( .A(P1_IR_REG_2__SCAN_IN), .B(keyinput_92), .ZN(n9975) );
  AOI211_X1 U10874 ( .C1(n9978), .C2(n9977), .A(n9976), .B(n9975), .ZN(n9981)
         );
  XNOR2_X1 U10875 ( .A(n6439), .B(keyinput_94), .ZN(n9980) );
  XNOR2_X1 U10876 ( .A(P1_IR_REG_5__SCAN_IN), .B(keyinput_95), .ZN(n9979) );
  OAI21_X1 U10877 ( .B1(n9981), .B2(n9980), .A(n9979), .ZN(n9985) );
  XOR2_X1 U10878 ( .A(P1_IR_REG_7__SCAN_IN), .B(keyinput_97), .Z(n9984) );
  XNOR2_X1 U10879 ( .A(P1_IR_REG_8__SCAN_IN), .B(keyinput_98), .ZN(n9983) );
  XNOR2_X1 U10880 ( .A(P1_IR_REG_6__SCAN_IN), .B(keyinput_96), .ZN(n9982) );
  NAND4_X1 U10881 ( .A1(n9985), .A2(n9984), .A3(n9983), .A4(n9982), .ZN(n9990)
         );
  XNOR2_X1 U10882 ( .A(n9986), .B(keyinput_99), .ZN(n9989) );
  XNOR2_X1 U10883 ( .A(n9987), .B(keyinput_100), .ZN(n9988) );
  AOI21_X1 U10884 ( .B1(n9990), .B2(n9989), .A(n9988), .ZN(n9994) );
  XNOR2_X1 U10885 ( .A(P1_IR_REG_11__SCAN_IN), .B(keyinput_101), .ZN(n9993) );
  XNOR2_X1 U10886 ( .A(P1_IR_REG_13__SCAN_IN), .B(keyinput_103), .ZN(n9992) );
  XNOR2_X1 U10887 ( .A(P1_IR_REG_12__SCAN_IN), .B(keyinput_102), .ZN(n9991) );
  NOR4_X1 U10888 ( .A1(n9994), .A2(n9993), .A3(n9992), .A4(n9991), .ZN(n9998)
         );
  XNOR2_X1 U10889 ( .A(n9995), .B(keyinput_104), .ZN(n9997) );
  XNOR2_X1 U10890 ( .A(P1_IR_REG_15__SCAN_IN), .B(keyinput_105), .ZN(n9996) );
  OAI21_X1 U10891 ( .B1(n9998), .B2(n9997), .A(n9996), .ZN(n10003) );
  XNOR2_X1 U10892 ( .A(n9999), .B(keyinput_106), .ZN(n10002) );
  XNOR2_X1 U10893 ( .A(P1_IR_REG_18__SCAN_IN), .B(keyinput_108), .ZN(n10001)
         );
  XNOR2_X1 U10894 ( .A(P1_IR_REG_17__SCAN_IN), .B(keyinput_107), .ZN(n10000)
         );
  AOI211_X1 U10895 ( .C1(n10003), .C2(n10002), .A(n10001), .B(n10000), .ZN(
        n10007) );
  XNOR2_X1 U10896 ( .A(n10004), .B(keyinput_109), .ZN(n10006) );
  XNOR2_X1 U10897 ( .A(P1_IR_REG_20__SCAN_IN), .B(keyinput_110), .ZN(n10005)
         );
  NOR3_X1 U10898 ( .A1(n10007), .A2(n10006), .A3(n10005), .ZN(n10012) );
  XNOR2_X1 U10899 ( .A(P1_IR_REG_21__SCAN_IN), .B(keyinput_111), .ZN(n10011)
         );
  XNOR2_X1 U10900 ( .A(n10008), .B(keyinput_113), .ZN(n10010) );
  XNOR2_X1 U10901 ( .A(P1_IR_REG_22__SCAN_IN), .B(keyinput_112), .ZN(n10009)
         );
  OAI211_X1 U10902 ( .C1(n10012), .C2(n10011), .A(n10010), .B(n10009), .ZN(
        n10017) );
  XNOR2_X1 U10903 ( .A(n10013), .B(keyinput_115), .ZN(n10016) );
  XNOR2_X1 U10904 ( .A(P1_IR_REG_24__SCAN_IN), .B(keyinput_114), .ZN(n10015)
         );
  XNOR2_X1 U10905 ( .A(P1_IR_REG_26__SCAN_IN), .B(keyinput_116), .ZN(n10014)
         );
  NAND4_X1 U10906 ( .A1(n10017), .A2(n10016), .A3(n10015), .A4(n10014), .ZN(
        n10021) );
  XNOR2_X1 U10907 ( .A(n10018), .B(keyinput_117), .ZN(n10020) );
  XOR2_X1 U10908 ( .A(P1_IR_REG_28__SCAN_IN), .B(keyinput_118), .Z(n10019) );
  AOI21_X1 U10909 ( .B1(n10021), .B2(n10020), .A(n10019), .ZN(n10026) );
  XOR2_X1 U10910 ( .A(P1_IR_REG_29__SCAN_IN), .B(keyinput_119), .Z(n10025) );
  XOR2_X1 U10911 ( .A(P1_IR_REG_31__SCAN_IN), .B(keyinput_121), .Z(n10024) );
  XNOR2_X1 U10912 ( .A(n10022), .B(keyinput_120), .ZN(n10023) );
  OAI211_X1 U10913 ( .C1(n10026), .C2(n10025), .A(n10024), .B(n10023), .ZN(
        n10029) );
  XNOR2_X1 U10914 ( .A(P1_D_REG_0__SCAN_IN), .B(keyinput_122), .ZN(n10028) );
  XNOR2_X1 U10915 ( .A(P1_D_REG_1__SCAN_IN), .B(keyinput_123), .ZN(n10027) );
  AOI21_X1 U10916 ( .B1(n10029), .B2(n10028), .A(n10027), .ZN(n10033) );
  INV_X1 U10917 ( .A(P1_D_REG_2__SCAN_IN), .ZN(n10708) );
  XNOR2_X1 U10918 ( .A(n10708), .B(keyinput_124), .ZN(n10032) );
  XNOR2_X1 U10919 ( .A(n10710), .B(keyinput_126), .ZN(n10031) );
  XNOR2_X1 U10920 ( .A(P1_D_REG_3__SCAN_IN), .B(keyinput_125), .ZN(n10030) );
  OAI211_X1 U10921 ( .C1(n10033), .C2(n10032), .A(n10031), .B(n10030), .ZN(
        n10034) );
  OAI211_X1 U10922 ( .C1(n10037), .C2(n10036), .A(n10035), .B(n10034), .ZN(
        n10038) );
  XOR2_X1 U10923 ( .A(n10039), .B(n10038), .Z(P2_U3287) );
  INV_X1 U10924 ( .A(n10040), .ZN(n10041) );
  MUX2_X1 U10925 ( .A(n10041), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3295) );
  AOI22_X1 U10926 ( .A1(n10261), .A2(n10275), .B1(P1_REG3_REG_27__SCAN_IN), 
        .B2(P1_U3086), .ZN(n10044) );
  OAI21_X1 U10927 ( .B1(n10426), .B2(n10259), .A(n10044), .ZN(n10045) );
  AOI21_X1 U10928 ( .B1(n10429), .B2(n10250), .A(n10045), .ZN(n10046) );
  NAND2_X1 U10929 ( .A1(n10048), .A2(n10047), .ZN(n10049) );
  XOR2_X1 U10930 ( .A(n10050), .B(n10049), .Z(n10055) );
  NAND2_X1 U10931 ( .A1(P1_REG3_REG_14__SCAN_IN), .A2(P1_U3086), .ZN(n10819)
         );
  OAI21_X1 U10932 ( .B1(n10259), .B2(n11136), .A(n10819), .ZN(n10051) );
  AOI21_X1 U10933 ( .B1(n10261), .B2(n11115), .A(n10051), .ZN(n10052) );
  OAI21_X1 U10934 ( .B1(n11148), .B2(n10263), .A(n10052), .ZN(n10053) );
  AOI21_X1 U10935 ( .B1(n11152), .B2(n10266), .A(n10053), .ZN(n10054) );
  OAI21_X1 U10936 ( .B1(n10055), .B2(n10269), .A(n10054), .ZN(P1_U3215) );
  INV_X1 U10937 ( .A(n10058), .ZN(n10056) );
  NAND2_X1 U10938 ( .A1(n10057), .A2(n10056), .ZN(n10198) );
  NAND2_X1 U10939 ( .A1(n10198), .A2(n10197), .ZN(n10195) );
  INV_X1 U10940 ( .A(n10057), .ZN(n10059) );
  NAND2_X1 U10941 ( .A1(n10059), .A2(n10058), .ZN(n10199) );
  NAND2_X1 U10942 ( .A1(n10195), .A2(n10199), .ZN(n10063) );
  XNOR2_X1 U10943 ( .A(n10061), .B(n10060), .ZN(n10062) );
  XNOR2_X1 U10944 ( .A(n10063), .B(n10062), .ZN(n10070) );
  INV_X1 U10945 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n10064) );
  OAI22_X1 U10946 ( .A1(n10259), .A2(n10496), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n10064), .ZN(n10065) );
  AOI21_X1 U10947 ( .B1(n10261), .B2(n10279), .A(n10065), .ZN(n10066) );
  OAI21_X1 U10948 ( .B1(n10499), .B2(n10263), .A(n10066), .ZN(n10067) );
  AOI21_X1 U10949 ( .B1(n10068), .B2(n10266), .A(n10067), .ZN(n10069) );
  OAI21_X1 U10950 ( .B1(n10070), .B2(n10269), .A(n10069), .ZN(P1_U3216) );
  NAND2_X1 U10951 ( .A1(n10072), .A2(n10071), .ZN(n10074) );
  XNOR2_X1 U10952 ( .A(n10074), .B(n10073), .ZN(n10082) );
  NAND2_X1 U10953 ( .A1(P1_U3086), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n10882)
         );
  INV_X1 U10954 ( .A(n10882), .ZN(n10076) );
  NOR2_X1 U10955 ( .A1(n10259), .A2(n10119), .ZN(n10075) );
  AOI211_X1 U10956 ( .C1(n10261), .C2(n10290), .A(n10076), .B(n10075), .ZN(
        n10077) );
  OAI21_X1 U10957 ( .B1(n10078), .B2(n10263), .A(n10077), .ZN(n10079) );
  AOI21_X1 U10958 ( .B1(n10080), .B2(n10266), .A(n10079), .ZN(n10081) );
  OAI21_X1 U10959 ( .B1(n10082), .B2(n10269), .A(n10081), .ZN(P1_U3217) );
  XOR2_X1 U10960 ( .A(n10084), .B(n10083), .Z(n10089) );
  NAND2_X1 U10961 ( .A1(P1_U3086), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n10410)
         );
  OAI21_X1 U10962 ( .B1(n10259), .B2(n10568), .A(n10410), .ZN(n10085) );
  AOI21_X1 U10963 ( .B1(n10261), .B2(n10283), .A(n10085), .ZN(n10086) );
  OAI21_X1 U10964 ( .B1(n10581), .B2(n10263), .A(n10086), .ZN(n10087) );
  AOI21_X1 U10965 ( .B1(n10579), .B2(n10266), .A(n10087), .ZN(n10088) );
  OAI21_X1 U10966 ( .B1(n10089), .B2(n10269), .A(n10088), .ZN(P1_U3219) );
  NAND2_X1 U10967 ( .A1(n10091), .A2(n10090), .ZN(n10092) );
  XOR2_X1 U10968 ( .A(n10093), .B(n10092), .Z(n10103) );
  INV_X1 U10969 ( .A(n10094), .ZN(n10095) );
  AOI21_X1 U10970 ( .B1(n10261), .B2(n5297), .A(n10095), .ZN(n10098) );
  OR2_X1 U10971 ( .A1(n10259), .A2(n10096), .ZN(n10097) );
  OAI211_X1 U10972 ( .C1(n10263), .C2(n10099), .A(n10098), .B(n10097), .ZN(
        n10100) );
  AOI21_X1 U10973 ( .B1(n10101), .B2(n10266), .A(n10100), .ZN(n10102) );
  OAI21_X1 U10974 ( .B1(n10103), .B2(n10269), .A(n10102), .ZN(P1_U3221) );
  AOI21_X1 U10975 ( .B1(n10104), .B2(n10105), .A(n10269), .ZN(n10107) );
  NAND2_X1 U10976 ( .A1(n10107), .A2(n10106), .ZN(n10112) );
  INV_X1 U10977 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n10108) );
  OAI22_X1 U10978 ( .A1(n10259), .A2(n10531), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n10108), .ZN(n10110) );
  NOR2_X1 U10979 ( .A1(n10263), .A2(n10539), .ZN(n10109) );
  AOI211_X1 U10980 ( .C1(n10261), .C2(n10281), .A(n10110), .B(n10109), .ZN(
        n10111) );
  OAI211_X1 U10981 ( .C1(n6707), .C2(n10253), .A(n10112), .B(n10111), .ZN(
        P1_U3223) );
  INV_X1 U10982 ( .A(n10184), .ZN(n10115) );
  AOI21_X1 U10983 ( .B1(n10212), .B2(n10207), .A(n10113), .ZN(n10114) );
  OAI21_X1 U10984 ( .B1(n10115), .B2(n10114), .A(n10244), .ZN(n10123) );
  INV_X1 U10985 ( .A(n10116), .ZN(n10121) );
  AOI21_X1 U10986 ( .B1(n10233), .B2(n11115), .A(n10117), .ZN(n10118) );
  OAI21_X1 U10987 ( .B1(n10119), .B2(n10236), .A(n10118), .ZN(n10120) );
  AOI21_X1 U10988 ( .B1(n10121), .B2(n10250), .A(n10120), .ZN(n10122) );
  OAI211_X1 U10989 ( .C1(n11096), .C2(n10253), .A(n10123), .B(n10122), .ZN(
        P1_U3224) );
  OAI21_X1 U10990 ( .B1(n10125), .B2(n10124), .A(n10242), .ZN(n10126) );
  NAND2_X1 U10991 ( .A1(n10126), .A2(n10244), .ZN(n10131) );
  INV_X1 U10992 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n10127) );
  OAI22_X1 U10993 ( .A1(n10259), .A2(n10462), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n10127), .ZN(n10129) );
  NOR2_X1 U10994 ( .A1(n10263), .A2(n10469), .ZN(n10128) );
  AOI211_X1 U10995 ( .C1(n10261), .C2(n10277), .A(n10129), .B(n10128), .ZN(
        n10130) );
  OAI211_X1 U10996 ( .C1(n6745), .C2(n10253), .A(n10131), .B(n10130), .ZN(
        P1_U3225) );
  INV_X1 U10997 ( .A(n10132), .ZN(n10133) );
  AOI21_X1 U10998 ( .B1(n10135), .B2(n10134), .A(n10133), .ZN(n10141) );
  AND2_X1 U10999 ( .A1(P1_U3086), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n10378) );
  NOR2_X1 U11000 ( .A1(n10259), .A2(n10237), .ZN(n10136) );
  AOI211_X1 U11001 ( .C1(n10261), .C2(n10286), .A(n10378), .B(n10136), .ZN(
        n10137) );
  OAI21_X1 U11002 ( .B1(n10138), .B2(n10263), .A(n10137), .ZN(n10139) );
  AOI21_X1 U11003 ( .B1(n10646), .B2(n10266), .A(n10139), .ZN(n10140) );
  OAI21_X1 U11004 ( .B1(n10141), .B2(n10269), .A(n10140), .ZN(P1_U3226) );
  NAND2_X1 U11005 ( .A1(n10143), .A2(n10142), .ZN(n10144) );
  XNOR2_X1 U11006 ( .A(n10145), .B(n10144), .ZN(n10151) );
  NAND2_X1 U11007 ( .A1(n10261), .A2(n10285), .ZN(n10146) );
  NAND2_X1 U11008 ( .A1(P1_REG3_REG_17__SCAN_IN), .A2(P1_U3086), .ZN(n10843)
         );
  OAI211_X1 U11009 ( .C1(n10569), .C2(n10259), .A(n10146), .B(n10843), .ZN(
        n10148) );
  NOR2_X1 U11010 ( .A1(n10686), .A2(n10253), .ZN(n10147) );
  AOI211_X1 U11011 ( .C1(n10250), .C2(n10149), .A(n10148), .B(n10147), .ZN(
        n10150) );
  OAI21_X1 U11012 ( .B1(n10151), .B2(n10269), .A(n10150), .ZN(P1_U3228) );
  INV_X1 U11013 ( .A(n10153), .ZN(n10154) );
  NOR2_X1 U11014 ( .A1(n10155), .A2(n10154), .ZN(n10156) );
  XNOR2_X1 U11015 ( .A(n10157), .B(n10156), .ZN(n10163) );
  INV_X1 U11016 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n10158) );
  OAI22_X1 U11017 ( .A1(n10259), .A2(n10484), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n10158), .ZN(n10159) );
  AOI21_X1 U11018 ( .B1(n10261), .B2(n10278), .A(n10159), .ZN(n10160) );
  OAI21_X1 U11019 ( .B1(n10488), .B2(n10263), .A(n10160), .ZN(n10161) );
  AOI21_X1 U11020 ( .B1(n10603), .B2(n10266), .A(n10161), .ZN(n10162) );
  OAI21_X1 U11021 ( .B1(n10163), .B2(n10269), .A(n10162), .ZN(P1_U3229) );
  XOR2_X1 U11022 ( .A(n10165), .B(n10164), .Z(n10174) );
  NAND2_X1 U11023 ( .A1(n10250), .A2(n10166), .ZN(n10169) );
  NOR2_X1 U11024 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n10167), .ZN(n10359) );
  AOI21_X1 U11025 ( .B1(n10233), .B2(n10289), .A(n10359), .ZN(n10168) );
  OAI211_X1 U11026 ( .C1(n10170), .C2(n10236), .A(n10169), .B(n10168), .ZN(
        n10171) );
  AOI21_X1 U11027 ( .B1(n10172), .B2(n10266), .A(n10171), .ZN(n10173) );
  OAI21_X1 U11028 ( .B1(n10174), .B2(n10269), .A(n10173), .ZN(P1_U3231) );
  XNOR2_X1 U11029 ( .A(n10175), .B(n10176), .ZN(n10177) );
  NAND2_X1 U11030 ( .A1(n10177), .A2(n10244), .ZN(n10182) );
  OAI22_X1 U11031 ( .A1(n10259), .A2(n10551), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n10178), .ZN(n10180) );
  NOR2_X1 U11032 ( .A1(n10236), .A2(n10550), .ZN(n10179) );
  AOI211_X1 U11033 ( .C1(n10250), .C2(n10556), .A(n10180), .B(n10179), .ZN(
        n10181) );
  OAI211_X1 U11034 ( .C1(n10676), .C2(n10253), .A(n10182), .B(n10181), .ZN(
        P1_U3233) );
  AND2_X1 U11035 ( .A1(n10184), .A2(n10183), .ZN(n10187) );
  OAI211_X1 U11036 ( .C1(n10187), .C2(n10186), .A(n10244), .B(n10185), .ZN(
        n10194) );
  NOR2_X1 U11037 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n10188), .ZN(n10866) );
  AOI21_X1 U11038 ( .B1(n10261), .B2(n10287), .A(n10866), .ZN(n10189) );
  OAI21_X1 U11039 ( .B1(n10190), .B2(n10259), .A(n10189), .ZN(n10191) );
  AOI21_X1 U11040 ( .B1(n10192), .B2(n10250), .A(n10191), .ZN(n10193) );
  OAI211_X1 U11041 ( .C1(n11116), .C2(n10253), .A(n10194), .B(n10193), .ZN(
        P1_U3234) );
  INV_X1 U11042 ( .A(n10613), .ZN(n10512) );
  INV_X1 U11043 ( .A(n10199), .ZN(n10196) );
  NOR2_X1 U11044 ( .A1(n10196), .A2(n10195), .ZN(n10201) );
  AOI21_X1 U11045 ( .B1(n10199), .B2(n10198), .A(n10197), .ZN(n10200) );
  OAI21_X1 U11046 ( .B1(n10201), .B2(n10200), .A(n10244), .ZN(n10206) );
  INV_X1 U11047 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n10202) );
  OAI22_X1 U11048 ( .A1(n10259), .A2(n10515), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n10202), .ZN(n10204) );
  NOR2_X1 U11049 ( .A1(n10263), .A2(n10509), .ZN(n10203) );
  AOI211_X1 U11050 ( .C1(n10261), .C2(n10280), .A(n10204), .B(n10203), .ZN(
        n10205) );
  OAI211_X1 U11051 ( .C1(n10512), .C2(n10253), .A(n10206), .B(n10205), .ZN(
        P1_U3235) );
  INV_X1 U11052 ( .A(n10207), .ZN(n10211) );
  OAI21_X1 U11053 ( .B1(n10209), .B2(n10211), .A(n10208), .ZN(n10210) );
  OAI211_X1 U11054 ( .C1(n10212), .C2(n10211), .A(n10244), .B(n10210), .ZN(
        n10218) );
  NAND2_X1 U11055 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_U3086), .ZN(n10807)
         );
  OAI21_X1 U11056 ( .B1(n10259), .B2(n10213), .A(n10807), .ZN(n10216) );
  NOR2_X1 U11057 ( .A1(n10263), .A2(n10214), .ZN(n10215) );
  AOI211_X1 U11058 ( .C1(n10261), .C2(n10289), .A(n10216), .B(n10215), .ZN(
        n10217) );
  OAI211_X1 U11059 ( .C1(n11087), .C2(n10253), .A(n10218), .B(n10217), .ZN(
        P1_U3236) );
  OAI21_X1 U11060 ( .B1(n10221), .B2(n10220), .A(n10219), .ZN(n10222) );
  NAND2_X1 U11061 ( .A1(n10222), .A2(n10244), .ZN(n10226) );
  AOI22_X1 U11062 ( .A1(n10233), .A2(n11001), .B1(n6484), .B2(n10266), .ZN(
        n10225) );
  AOI22_X1 U11063 ( .A1(n10223), .A2(P1_REG3_REG_2__SCAN_IN), .B1(n10261), 
        .B2(n11000), .ZN(n10224) );
  NAND3_X1 U11064 ( .A1(n10226), .A2(n10225), .A3(n10224), .ZN(P1_U3237) );
  NAND2_X1 U11065 ( .A1(n10227), .A2(n10228), .ZN(n10230) );
  XNOR2_X1 U11066 ( .A(n10230), .B(n10229), .ZN(n10240) );
  NAND2_X1 U11067 ( .A1(n10250), .A2(n10231), .ZN(n10235) );
  NOR2_X1 U11068 ( .A1(n10232), .A2(P1_STATE_REG_SCAN_IN), .ZN(n10855) );
  AOI21_X1 U11069 ( .B1(n10233), .B2(n10282), .A(n10855), .ZN(n10234) );
  OAI211_X1 U11070 ( .C1(n10237), .C2(n10236), .A(n10235), .B(n10234), .ZN(
        n10238) );
  AOI21_X1 U11071 ( .B1(n10636), .B2(n10266), .A(n10238), .ZN(n10239) );
  OAI21_X1 U11072 ( .B1(n10240), .B2(n10269), .A(n10239), .ZN(P1_U3238) );
  AND2_X1 U11073 ( .A1(n10242), .A2(n10241), .ZN(n10246) );
  OAI211_X1 U11074 ( .C1(n10246), .C2(n10245), .A(n10244), .B(n10243), .ZN(
        n10252) );
  INV_X1 U11075 ( .A(n10247), .ZN(n10451) );
  AOI22_X1 U11076 ( .A1(n10261), .A2(n10276), .B1(P1_REG3_REG_26__SCAN_IN), 
        .B2(P1_U3086), .ZN(n10248) );
  OAI21_X1 U11077 ( .B1(n10446), .B2(n10259), .A(n10248), .ZN(n10249) );
  AOI21_X1 U11078 ( .B1(n10451), .B2(n10250), .A(n10249), .ZN(n10251) );
  OAI211_X1 U11079 ( .C1(n10660), .C2(n10253), .A(n10252), .B(n10251), .ZN(
        P1_U3240) );
  XNOR2_X1 U11080 ( .A(n10255), .B(n10254), .ZN(n10256) );
  XNOR2_X1 U11081 ( .A(n10257), .B(n10256), .ZN(n10270) );
  NAND2_X1 U11082 ( .A1(P1_REG3_REG_15__SCAN_IN), .A2(P1_U3086), .ZN(n10829)
         );
  OAI21_X1 U11083 ( .B1(n10259), .B2(n10258), .A(n10829), .ZN(n10260) );
  AOI21_X1 U11084 ( .B1(n10261), .B2(n6629), .A(n10260), .ZN(n10262) );
  OAI21_X1 U11085 ( .B1(n10264), .B2(n10263), .A(n10262), .ZN(n10265) );
  AOI21_X1 U11086 ( .B1(n10267), .B2(n10266), .A(n10265), .ZN(n10268) );
  OAI21_X1 U11087 ( .B1(n10270), .B2(n10269), .A(n10268), .ZN(P1_U3241) );
  MUX2_X1 U11088 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(n10271), .S(P1_U3973), .Z(
        P1_U3585) );
  MUX2_X1 U11089 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n10272), .S(P1_U3973), .Z(
        P1_U3584) );
  MUX2_X1 U11090 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n10273), .S(P1_U3973), .Z(
        P1_U3582) );
  MUX2_X1 U11091 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n10274), .S(P1_U3973), .Z(
        P1_U3581) );
  MUX2_X1 U11092 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n10275), .S(P1_U3973), .Z(
        P1_U3580) );
  MUX2_X1 U11093 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n10276), .S(P1_U3973), .Z(
        P1_U3579) );
  MUX2_X1 U11094 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n10277), .S(P1_U3973), .Z(
        P1_U3578) );
  MUX2_X1 U11095 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n10278), .S(P1_U3973), .Z(
        P1_U3577) );
  MUX2_X1 U11096 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n10279), .S(P1_U3973), .Z(
        P1_U3576) );
  MUX2_X1 U11097 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n10280), .S(P1_U3973), .Z(
        P1_U3575) );
  MUX2_X1 U11098 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n10281), .S(P1_U3973), .Z(
        P1_U3574) );
  MUX2_X1 U11099 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n10282), .S(P1_U3973), .Z(
        P1_U3573) );
  MUX2_X1 U11100 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n10283), .S(P1_U3973), .Z(
        P1_U3572) );
  MUX2_X1 U11101 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n10284), .S(P1_U3973), .Z(
        P1_U3571) );
  MUX2_X1 U11102 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n10285), .S(P1_U3973), .Z(
        P1_U3570) );
  MUX2_X1 U11103 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n10286), .S(P1_U3973), .Z(
        P1_U3569) );
  MUX2_X1 U11104 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n6629), .S(P1_U3973), .Z(
        P1_U3568) );
  MUX2_X1 U11105 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n11115), .S(P1_U3973), .Z(
        P1_U3567) );
  MUX2_X1 U11106 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n10287), .S(P1_U3973), .Z(
        P1_U3566) );
  MUX2_X1 U11107 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n10288), .S(P1_U3973), .Z(
        P1_U3565) );
  MUX2_X1 U11108 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n10289), .S(P1_U3973), .Z(
        P1_U3564) );
  MUX2_X1 U11109 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n10290), .S(P1_U3973), .Z(
        P1_U3563) );
  MUX2_X1 U11110 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n10291), .S(P1_U3973), .Z(
        P1_U3562) );
  MUX2_X1 U11111 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n5297), .S(P1_U3973), .Z(
        P1_U3561) );
  MUX2_X1 U11112 ( .A(n10292), .B(P1_DATAO_REG_6__SCAN_IN), .S(n10296), .Z(
        P1_U3560) );
  MUX2_X1 U11113 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n10293), .S(P1_U3973), .Z(
        P1_U3559) );
  MUX2_X1 U11114 ( .A(n10294), .B(P1_DATAO_REG_4__SCAN_IN), .S(n10296), .Z(
        P1_U3558) );
  MUX2_X1 U11115 ( .A(n11001), .B(P1_DATAO_REG_3__SCAN_IN), .S(n10296), .Z(
        P1_U3557) );
  MUX2_X1 U11116 ( .A(n10295), .B(P1_DATAO_REG_2__SCAN_IN), .S(n10296), .Z(
        P1_U3556) );
  MUX2_X1 U11117 ( .A(n11000), .B(P1_DATAO_REG_1__SCAN_IN), .S(n10296), .Z(
        P1_U3555) );
  MUX2_X1 U11118 ( .A(n10297), .B(P1_DATAO_REG_0__SCAN_IN), .S(n10296), .Z(
        P1_U3554) );
  OAI211_X1 U11119 ( .C1(n10300), .C2(n10299), .A(n10841), .B(n10298), .ZN(
        n10308) );
  AOI22_X1 U11120 ( .A1(n10868), .A2(P1_ADDR_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(P1_U3086), .ZN(n10307) );
  NAND2_X1 U11121 ( .A1(n10881), .A2(n10301), .ZN(n10306) );
  OAI211_X1 U11122 ( .C1(n10304), .C2(n10303), .A(n10838), .B(n10302), .ZN(
        n10305) );
  NAND4_X1 U11123 ( .A1(n10308), .A2(n10307), .A3(n10306), .A4(n10305), .ZN(
        P1_U3244) );
  NAND3_X1 U11124 ( .A1(n10309), .A2(n10790), .A3(n10792), .ZN(n10315) );
  INV_X1 U11125 ( .A(n10310), .ZN(n10313) );
  OAI21_X1 U11126 ( .B1(P1_IR_REG_0__SCAN_IN), .B2(P1_REG2_REG_0__SCAN_IN), 
        .A(n10311), .ZN(n10312) );
  AOI22_X1 U11127 ( .A1(n10313), .A2(n10312), .B1(n10705), .B2(n10793), .ZN(
        n10314) );
  NAND3_X1 U11128 ( .A1(n10315), .A2(P1_U3973), .A3(n10314), .ZN(n10354) );
  AOI22_X1 U11129 ( .A1(n10868), .A2(P1_ADDR_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(P1_U3086), .ZN(n10327) );
  OAI211_X1 U11130 ( .C1(n10318), .C2(n10317), .A(n10841), .B(n10316), .ZN(
        n10323) );
  OAI211_X1 U11131 ( .C1(n10321), .C2(n10320), .A(n10838), .B(n10319), .ZN(
        n10322) );
  AND2_X1 U11132 ( .A1(n10323), .A2(n10322), .ZN(n10326) );
  NAND2_X1 U11133 ( .A1(n10881), .A2(n10324), .ZN(n10325) );
  NAND4_X1 U11134 ( .A1(n10354), .A2(n10327), .A3(n10326), .A4(n10325), .ZN(
        P1_U3245) );
  INV_X1 U11135 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n10329) );
  OAI21_X1 U11136 ( .B1(n10885), .B2(n10329), .A(n10328), .ZN(n10330) );
  AOI21_X1 U11137 ( .B1(n10331), .B2(n10881), .A(n10330), .ZN(n10340) );
  OAI211_X1 U11138 ( .C1(n10334), .C2(n10333), .A(n10841), .B(n10332), .ZN(
        n10339) );
  OAI211_X1 U11139 ( .C1(n10337), .C2(n10336), .A(n10838), .B(n10335), .ZN(
        n10338) );
  NAND3_X1 U11140 ( .A1(n10340), .A2(n10339), .A3(n10338), .ZN(P1_U3246) );
  AOI21_X1 U11141 ( .B1(n10868), .B2(P1_ADDR_REG_4__SCAN_IN), .A(n10341), .ZN(
        n10353) );
  OAI211_X1 U11142 ( .C1(n10344), .C2(n10343), .A(n10841), .B(n10342), .ZN(
        n10349) );
  OAI211_X1 U11143 ( .C1(n10347), .C2(n10346), .A(n10838), .B(n10345), .ZN(
        n10348) );
  AND2_X1 U11144 ( .A1(n10349), .A2(n10348), .ZN(n10352) );
  NAND2_X1 U11145 ( .A1(n10881), .A2(n10350), .ZN(n10351) );
  NAND4_X1 U11146 ( .A1(n10354), .A2(n10353), .A3(n10352), .A4(n10351), .ZN(
        P1_U3247) );
  OAI21_X1 U11147 ( .B1(n10357), .B2(n10356), .A(n10355), .ZN(n10358) );
  NAND2_X1 U11148 ( .A1(n10358), .A2(n10838), .ZN(n10368) );
  AOI21_X1 U11149 ( .B1(n10868), .B2(P1_ADDR_REG_9__SCAN_IN), .A(n10359), .ZN(
        n10367) );
  OAI21_X1 U11150 ( .B1(n10362), .B2(n10361), .A(n10360), .ZN(n10363) );
  NAND2_X1 U11151 ( .A1(n10363), .A2(n10841), .ZN(n10366) );
  NAND2_X1 U11152 ( .A1(n10881), .A2(n10364), .ZN(n10365) );
  NAND4_X1 U11153 ( .A1(n10368), .A2(n10367), .A3(n10366), .A4(n10365), .ZN(
        P1_U3252) );
  NOR2_X1 U11154 ( .A1(n10864), .A2(n10370), .ZN(n10369) );
  AOI21_X1 U11155 ( .B1(n10370), .B2(n10864), .A(n10369), .ZN(n10857) );
  OAI21_X1 U11156 ( .B1(P1_REG1_REG_12__SCAN_IN), .B2(n10382), .A(n10371), 
        .ZN(n10858) );
  INV_X1 U11157 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n11145) );
  NOR2_X1 U11158 ( .A1(n10818), .A2(n11145), .ZN(n10372) );
  AOI21_X1 U11159 ( .B1(n10818), .B2(n11145), .A(n10372), .ZN(n10815) );
  NOR2_X1 U11160 ( .A1(n10373), .A2(n10385), .ZN(n10374) );
  INV_X1 U11161 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n11170) );
  XNOR2_X1 U11162 ( .A(n10385), .B(n10373), .ZN(n10823) );
  NOR2_X1 U11163 ( .A1(n11170), .A2(n10823), .ZN(n10822) );
  NOR2_X1 U11164 ( .A1(n10374), .A2(n10822), .ZN(n10377) );
  AOI22_X1 U11165 ( .A1(n10403), .A2(P1_REG1_REG_16__SCAN_IN), .B1(n10375), 
        .B2(n10380), .ZN(n10376) );
  NAND2_X1 U11166 ( .A1(n10376), .A2(n10377), .ZN(n10402) );
  OAI21_X1 U11167 ( .B1(n10377), .B2(n10376), .A(n10402), .ZN(n10393) );
  AOI21_X1 U11168 ( .B1(n10868), .B2(P1_ADDR_REG_16__SCAN_IN), .A(n10378), 
        .ZN(n10379) );
  OAI21_X1 U11169 ( .B1(n10414), .B2(n10380), .A(n10379), .ZN(n10392) );
  OAI21_X1 U11170 ( .B1(P1_REG2_REG_12__SCAN_IN), .B2(n10382), .A(n10381), 
        .ZN(n10861) );
  NAND2_X1 U11171 ( .A1(n10864), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n10383) );
  OAI21_X1 U11172 ( .B1(n10864), .B2(P1_REG2_REG_13__SCAN_IN), .A(n10383), 
        .ZN(n10860) );
  NOR2_X1 U11173 ( .A1(n10861), .A2(n10860), .ZN(n10859) );
  AOI21_X1 U11174 ( .B1(P1_REG2_REG_13__SCAN_IN), .B2(n10864), .A(n10859), 
        .ZN(n10812) );
  NAND2_X1 U11175 ( .A1(n10818), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n10384) );
  OAI21_X1 U11176 ( .B1(n10818), .B2(P1_REG2_REG_14__SCAN_IN), .A(n10384), 
        .ZN(n10811) );
  NOR2_X1 U11177 ( .A1(n10812), .A2(n10811), .ZN(n10810) );
  AOI21_X1 U11178 ( .B1(P1_REG2_REG_14__SCAN_IN), .B2(n10818), .A(n10810), 
        .ZN(n10386) );
  NOR2_X1 U11179 ( .A1(n10386), .A2(n10385), .ZN(n10387) );
  XOR2_X1 U11180 ( .A(n10828), .B(n10386), .Z(n10825) );
  NOR2_X1 U11181 ( .A1(n8071), .A2(n10825), .ZN(n10824) );
  NOR2_X1 U11182 ( .A1(n10387), .A2(n10824), .ZN(n10390) );
  NAND2_X1 U11183 ( .A1(n10403), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n10388) );
  OAI21_X1 U11184 ( .B1(n10403), .B2(P1_REG2_REG_16__SCAN_IN), .A(n10388), 
        .ZN(n10389) );
  NOR2_X1 U11185 ( .A1(n10390), .A2(n10389), .ZN(n10396) );
  AOI211_X1 U11186 ( .C1(n10390), .C2(n10389), .A(n10396), .B(n10870), .ZN(
        n10391) );
  AOI211_X1 U11187 ( .C1(n10838), .C2(n10393), .A(n10392), .B(n10391), .ZN(
        n10394) );
  INV_X1 U11188 ( .A(n10394), .ZN(P1_U3259) );
  NAND2_X1 U11189 ( .A1(n10854), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n10397) );
  OAI21_X1 U11190 ( .B1(n10854), .B2(P1_REG2_REG_18__SCAN_IN), .A(n10397), 
        .ZN(n10847) );
  NOR2_X1 U11191 ( .A1(n10840), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n10395) );
  AOI21_X1 U11192 ( .B1(P1_REG2_REG_17__SCAN_IN), .B2(n10840), .A(n10395), 
        .ZN(n10833) );
  AOI21_X1 U11193 ( .B1(P1_REG2_REG_16__SCAN_IN), .B2(n10403), .A(n10396), 
        .ZN(n10834) );
  NAND2_X1 U11194 ( .A1(n10833), .A2(n10834), .ZN(n10832) );
  OAI21_X1 U11195 ( .B1(n10840), .B2(P1_REG2_REG_17__SCAN_IN), .A(n10832), 
        .ZN(n10848) );
  NOR2_X1 U11196 ( .A1(n10847), .A2(n10848), .ZN(n10846) );
  INV_X1 U11197 ( .A(n10846), .ZN(n10398) );
  NAND2_X1 U11198 ( .A1(n10398), .A2(n10397), .ZN(n10401) );
  INV_X1 U11199 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n10399) );
  MUX2_X1 U11200 ( .A(n10399), .B(P1_REG2_REG_19__SCAN_IN), .S(n7110), .Z(
        n10400) );
  XNOR2_X1 U11201 ( .A(n10401), .B(n10400), .ZN(n10409) );
  NAND2_X1 U11202 ( .A1(n10854), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n10404) );
  OAI21_X1 U11203 ( .B1(n10854), .B2(P1_REG1_REG_18__SCAN_IN), .A(n10404), 
        .ZN(n10850) );
  INV_X1 U11204 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n10642) );
  XNOR2_X1 U11205 ( .A(n10840), .B(n10642), .ZN(n10836) );
  INV_X1 U11206 ( .A(n10404), .ZN(n10405) );
  NOR2_X1 U11207 ( .A1(n10849), .A2(n10405), .ZN(n10407) );
  INV_X1 U11208 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n10632) );
  XNOR2_X1 U11209 ( .A(n7110), .B(n10632), .ZN(n10406) );
  XNOR2_X1 U11210 ( .A(n10407), .B(n10406), .ZN(n10408) );
  AOI22_X1 U11211 ( .A1(n10841), .A2(n10409), .B1(n10838), .B2(n10408), .ZN(
        n10413) );
  INV_X1 U11212 ( .A(n10410), .ZN(n10411) );
  AOI21_X1 U11213 ( .B1(n10868), .B2(P1_ADDR_REG_19__SCAN_IN), .A(n10411), 
        .ZN(n10412) );
  OAI211_X1 U11214 ( .C1(n6812), .C2(n10414), .A(n10413), .B(n10412), .ZN(
        P1_U3262) );
  NOR2_X1 U11215 ( .A1(n11011), .A2(n10415), .ZN(n10421) );
  NOR2_X1 U11216 ( .A1(n10416), .A2(n11014), .ZN(n10417) );
  AOI211_X1 U11217 ( .C1(n11011), .C2(P1_REG2_REG_31__SCAN_IN), .A(n10421), 
        .B(n10417), .ZN(n10418) );
  OAI21_X1 U11218 ( .B1(n10419), .B2(n11153), .A(n10418), .ZN(P1_U3263) );
  NOR2_X1 U11219 ( .A1(n8822), .A2(n11014), .ZN(n10420) );
  AOI211_X1 U11220 ( .C1(n11011), .C2(P1_REG2_REG_30__SCAN_IN), .A(n10421), 
        .B(n10420), .ZN(n10422) );
  OAI21_X1 U11221 ( .B1(n11153), .B2(n10423), .A(n10422), .ZN(P1_U3264) );
  AOI211_X1 U11222 ( .C1(n10430), .C2(n10425), .A(n11132), .B(n10424), .ZN(
        n10428) );
  OAI22_X1 U11223 ( .A1(n10462), .A2(n11137), .B1(n10426), .B2(n11135), .ZN(
        n10427) );
  OR2_X1 U11224 ( .A1(n10428), .A2(n10427), .ZN(n10587) );
  AOI21_X1 U11225 ( .B1(n10429), .B2(n11149), .A(n10587), .ZN(n10439) );
  XNOR2_X1 U11226 ( .A(n10431), .B(n10430), .ZN(n10589) );
  NAND2_X1 U11227 ( .A1(n10589), .A2(n10575), .ZN(n10438) );
  INV_X1 U11228 ( .A(n10449), .ZN(n10433) );
  AOI211_X1 U11229 ( .C1(n10434), .C2(n10433), .A(n10577), .B(n10432), .ZN(
        n10588) );
  INV_X1 U11230 ( .A(P1_REG2_REG_27__SCAN_IN), .ZN(n10435) );
  OAI22_X1 U11231 ( .A1(n10656), .A2(n11014), .B1(n10435), .B2(n10560), .ZN(
        n10436) );
  AOI21_X1 U11232 ( .B1(n10588), .B2(n11018), .A(n10436), .ZN(n10437) );
  OAI211_X1 U11233 ( .C1(n11011), .C2(n10439), .A(n10438), .B(n10437), .ZN(
        P1_U3266) );
  XOR2_X1 U11234 ( .A(n10442), .B(n10440), .Z(n10594) );
  INV_X1 U11235 ( .A(n10594), .ZN(n10456) );
  INV_X1 U11236 ( .A(n10441), .ZN(n10461) );
  OAI21_X1 U11237 ( .B1(n10461), .B2(n10443), .A(n10442), .ZN(n10445) );
  AOI21_X1 U11238 ( .B1(n10445), .B2(n10444), .A(n11132), .ZN(n10448) );
  OAI22_X1 U11239 ( .A1(n10446), .A2(n11135), .B1(n10484), .B2(n11137), .ZN(
        n10447) );
  AOI211_X1 U11240 ( .C1(n10450), .C2(n10466), .A(n10577), .B(n10449), .ZN(
        n10593) );
  NAND2_X1 U11241 ( .A1(n10593), .A2(n11018), .ZN(n10453) );
  AOI22_X1 U11242 ( .A1(n11011), .A2(P1_REG2_REG_26__SCAN_IN), .B1(n10451), 
        .B2(n11149), .ZN(n10452) );
  OAI211_X1 U11243 ( .C1(n10660), .C2(n11014), .A(n10453), .B(n10452), .ZN(
        n10454) );
  AOI21_X1 U11244 ( .B1(n10560), .B2(n10592), .A(n10454), .ZN(n10455) );
  OAI21_X1 U11245 ( .B1(n10456), .B2(n10563), .A(n10455), .ZN(P1_U3267) );
  XNOR2_X1 U11246 ( .A(n10457), .B(n10458), .ZN(n10599) );
  INV_X1 U11247 ( .A(n10599), .ZN(n10475) );
  OAI21_X1 U11248 ( .B1(n10459), .B2(n10458), .A(n10566), .ZN(n10460) );
  OR2_X1 U11249 ( .A1(n10461), .A2(n10460), .ZN(n10465) );
  OAI22_X1 U11250 ( .A1(n10496), .A2(n11137), .B1(n10462), .B2(n11135), .ZN(
        n10463) );
  INV_X1 U11251 ( .A(n10463), .ZN(n10464) );
  NAND2_X1 U11252 ( .A1(n10465), .A2(n10464), .ZN(n10597) );
  INV_X1 U11253 ( .A(n10466), .ZN(n10467) );
  AOI211_X1 U11254 ( .C1(n10468), .C2(n10477), .A(n10577), .B(n10467), .ZN(
        n10598) );
  NAND2_X1 U11255 ( .A1(n10598), .A2(n11018), .ZN(n10472) );
  INV_X1 U11256 ( .A(n10469), .ZN(n10470) );
  AOI22_X1 U11257 ( .A1(n11011), .A2(P1_REG2_REG_25__SCAN_IN), .B1(n10470), 
        .B2(n11149), .ZN(n10471) );
  OAI211_X1 U11258 ( .C1(n6745), .C2(n11014), .A(n10472), .B(n10471), .ZN(
        n10473) );
  AOI21_X1 U11259 ( .B1(n10560), .B2(n10597), .A(n10473), .ZN(n10474) );
  OAI21_X1 U11260 ( .B1(n10475), .B2(n10563), .A(n10474), .ZN(P1_U3268) );
  XNOR2_X1 U11261 ( .A(n10476), .B(n10483), .ZN(n10606) );
  INV_X1 U11262 ( .A(n10477), .ZN(n10478) );
  AOI211_X1 U11263 ( .C1(n10603), .C2(n5148), .A(n10577), .B(n10478), .ZN(
        n10602) );
  INV_X1 U11264 ( .A(P1_REG2_REG_24__SCAN_IN), .ZN(n10479) );
  OAI22_X1 U11265 ( .A1(n10480), .A2(n11014), .B1(n10479), .B2(n10560), .ZN(
        n10481) );
  AOI21_X1 U11266 ( .B1(n10602), .B2(n11018), .A(n10481), .ZN(n10491) );
  AOI21_X1 U11267 ( .B1(n10483), .B2(n10482), .A(n11132), .ZN(n10487) );
  OAI22_X1 U11268 ( .A1(n10515), .A2(n11137), .B1(n10484), .B2(n11135), .ZN(
        n10485) );
  AOI21_X1 U11269 ( .B1(n10487), .B2(n10486), .A(n10485), .ZN(n10605) );
  OAI21_X1 U11270 ( .B1(n10488), .B2(n10580), .A(n10605), .ZN(n10489) );
  NAND2_X1 U11271 ( .A1(n10489), .A2(n10560), .ZN(n10490) );
  OAI211_X1 U11272 ( .C1(n10606), .C2(n10563), .A(n10491), .B(n10490), .ZN(
        P1_U3269) );
  XNOR2_X1 U11273 ( .A(n10492), .B(n10495), .ZN(n10609) );
  OAI21_X1 U11274 ( .B1(n10495), .B2(n10494), .A(n10493), .ZN(n10498) );
  OAI22_X1 U11275 ( .A1(n10531), .A2(n11137), .B1(n10496), .B2(n11135), .ZN(
        n10497) );
  AOI21_X1 U11276 ( .B1(n10498), .B2(n10566), .A(n10497), .ZN(n10608) );
  INV_X1 U11277 ( .A(n10608), .ZN(n10504) );
  OAI211_X1 U11278 ( .C1(n10668), .C2(n5197), .A(n11126), .B(n5148), .ZN(
        n10607) );
  NOR2_X1 U11279 ( .A1(n10607), .A2(n11153), .ZN(n10503) );
  INV_X1 U11280 ( .A(n10499), .ZN(n10500) );
  AOI22_X1 U11281 ( .A1(n11011), .A2(P1_REG2_REG_23__SCAN_IN), .B1(n10500), 
        .B2(n11149), .ZN(n10501) );
  OAI21_X1 U11282 ( .B1(n10668), .B2(n11014), .A(n10501), .ZN(n10502) );
  AOI211_X1 U11283 ( .C1(n10504), .C2(n10560), .A(n10503), .B(n10502), .ZN(
        n10505) );
  OAI21_X1 U11284 ( .B1(n10609), .B2(n10563), .A(n10505), .ZN(P1_U3270) );
  OAI21_X1 U11285 ( .B1(n10507), .B2(n10513), .A(n10506), .ZN(n10508) );
  INV_X1 U11286 ( .A(n10508), .ZN(n10616) );
  AOI211_X1 U11287 ( .C1(n10613), .C2(n10536), .A(n10577), .B(n5197), .ZN(
        n10612) );
  INV_X1 U11288 ( .A(n10509), .ZN(n10510) );
  AOI22_X1 U11289 ( .A1(n11011), .A2(P1_REG2_REG_22__SCAN_IN), .B1(n10510), 
        .B2(n11149), .ZN(n10511) );
  OAI21_X1 U11290 ( .B1(n10512), .B2(n11014), .A(n10511), .ZN(n10520) );
  AOI21_X1 U11291 ( .B1(n10514), .B2(n10513), .A(n11132), .ZN(n10518) );
  OAI22_X1 U11292 ( .A1(n10551), .A2(n11137), .B1(n10515), .B2(n11135), .ZN(
        n10516) );
  AOI21_X1 U11293 ( .B1(n10518), .B2(n10517), .A(n10516), .ZN(n10615) );
  NOR2_X1 U11294 ( .A1(n10615), .A2(n11011), .ZN(n10519) );
  AOI211_X1 U11295 ( .C1(n10612), .C2(n11018), .A(n10520), .B(n10519), .ZN(
        n10521) );
  OAI21_X1 U11296 ( .B1(n10616), .B2(n10563), .A(n10521), .ZN(P1_U3271) );
  OAI21_X1 U11297 ( .B1(n10524), .B2(n10523), .A(n10522), .ZN(n10619) );
  INV_X1 U11298 ( .A(n10619), .ZN(n10545) );
  INV_X1 U11299 ( .A(n10525), .ZN(n10527) );
  OAI21_X1 U11300 ( .B1(n10549), .B2(n10527), .A(n10526), .ZN(n10529) );
  XNOR2_X1 U11301 ( .A(n10529), .B(n10528), .ZN(n10530) );
  OR2_X1 U11302 ( .A1(n10530), .A2(n11132), .ZN(n10534) );
  OAI22_X1 U11303 ( .A1(n10568), .A2(n11137), .B1(n10531), .B2(n11135), .ZN(
        n10532) );
  INV_X1 U11304 ( .A(n10532), .ZN(n10533) );
  NAND2_X1 U11305 ( .A1(n10534), .A2(n10533), .ZN(n10617) );
  INV_X1 U11306 ( .A(n10535), .ZN(n10555) );
  INV_X1 U11307 ( .A(n10536), .ZN(n10537) );
  AOI211_X1 U11308 ( .C1(n10538), .C2(n10555), .A(n10577), .B(n10537), .ZN(
        n10618) );
  NAND2_X1 U11309 ( .A1(n10618), .A2(n11018), .ZN(n10542) );
  INV_X1 U11310 ( .A(n10539), .ZN(n10540) );
  AOI22_X1 U11311 ( .A1(n11011), .A2(P1_REG2_REG_21__SCAN_IN), .B1(n10540), 
        .B2(n11149), .ZN(n10541) );
  OAI211_X1 U11312 ( .C1(n6707), .C2(n11014), .A(n10542), .B(n10541), .ZN(
        n10543) );
  AOI21_X1 U11313 ( .B1(n10560), .B2(n10617), .A(n10543), .ZN(n10544) );
  OAI21_X1 U11314 ( .B1(n10545), .B2(n10563), .A(n10544), .ZN(P1_U3272) );
  XNOR2_X1 U11315 ( .A(n10547), .B(n10546), .ZN(n10624) );
  XNOR2_X1 U11316 ( .A(n10549), .B(n10548), .ZN(n10553) );
  OAI22_X1 U11317 ( .A1(n10551), .A2(n11135), .B1(n10550), .B2(n11137), .ZN(
        n10552) );
  AOI21_X1 U11318 ( .B1(n10553), .B2(n10566), .A(n10552), .ZN(n10623) );
  INV_X1 U11319 ( .A(n10623), .ZN(n10561) );
  INV_X1 U11320 ( .A(n10554), .ZN(n10576) );
  OAI211_X1 U11321 ( .C1(n10676), .C2(n10576), .A(n10555), .B(n11126), .ZN(
        n10622) );
  NOR2_X1 U11322 ( .A1(n10622), .A2(n11153), .ZN(n10559) );
  AOI22_X1 U11323 ( .A1(n11011), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n10556), 
        .B2(n11149), .ZN(n10557) );
  OAI21_X1 U11324 ( .B1(n10676), .B2(n11014), .A(n10557), .ZN(n10558) );
  AOI211_X1 U11325 ( .C1(n10561), .C2(n10560), .A(n10559), .B(n10558), .ZN(
        n10562) );
  OAI21_X1 U11326 ( .B1(n10624), .B2(n10563), .A(n10562), .ZN(P1_U3273) );
  XNOR2_X1 U11327 ( .A(n10565), .B(n10564), .ZN(n10567) );
  NAND2_X1 U11328 ( .A1(n10567), .A2(n10566), .ZN(n10572) );
  OAI22_X1 U11329 ( .A1(n10569), .A2(n11137), .B1(n10568), .B2(n11135), .ZN(
        n10570) );
  INV_X1 U11330 ( .A(n10570), .ZN(n10571) );
  NAND2_X1 U11331 ( .A1(n10572), .A2(n10571), .ZN(n10629) );
  INV_X1 U11332 ( .A(n10629), .ZN(n10586) );
  XNOR2_X1 U11333 ( .A(n10574), .B(n10573), .ZN(n10631) );
  NAND2_X1 U11334 ( .A1(n10631), .A2(n10575), .ZN(n10585) );
  AOI211_X1 U11335 ( .C1(n10579), .C2(n10578), .A(n10577), .B(n10576), .ZN(
        n10630) );
  NOR2_X1 U11336 ( .A1(n10680), .A2(n11014), .ZN(n10583) );
  OAI22_X1 U11337 ( .A1(n10560), .A2(n10399), .B1(n10581), .B2(n10580), .ZN(
        n10582) );
  AOI211_X1 U11338 ( .C1(n10630), .C2(n11018), .A(n10583), .B(n10582), .ZN(
        n10584) );
  OAI211_X1 U11339 ( .C1(n11011), .C2(n10586), .A(n10585), .B(n10584), .ZN(
        P1_U3274) );
  INV_X1 U11340 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n10590) );
  MUX2_X1 U11341 ( .A(n10590), .B(n10653), .S(n11171), .Z(n10591) );
  OAI21_X1 U11342 ( .B1(n10656), .B2(n10644), .A(n10591), .ZN(P1_U3549) );
  INV_X1 U11343 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n10595) );
  AOI211_X1 U11344 ( .C1(n10594), .C2(n11168), .A(n10593), .B(n10592), .ZN(
        n10657) );
  MUX2_X1 U11345 ( .A(n10595), .B(n10657), .S(n11171), .Z(n10596) );
  OAI21_X1 U11346 ( .B1(n10660), .B2(n10644), .A(n10596), .ZN(P1_U3548) );
  INV_X1 U11347 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n10600) );
  AOI211_X1 U11348 ( .C1(n10599), .C2(n11168), .A(n10598), .B(n10597), .ZN(
        n10661) );
  MUX2_X1 U11349 ( .A(n10600), .B(n10661), .S(n11171), .Z(n10601) );
  OAI21_X1 U11350 ( .B1(n6745), .B2(n10644), .A(n10601), .ZN(P1_U3547) );
  AOI21_X1 U11351 ( .B1(n10985), .B2(n10603), .A(n10602), .ZN(n10604) );
  OAI211_X1 U11352 ( .C1(n10606), .C2(n10649), .A(n10605), .B(n10604), .ZN(
        n10664) );
  MUX2_X1 U11353 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n10664), .S(n11171), .Z(
        P1_U3546) );
  OAI211_X1 U11354 ( .C1(n10609), .C2(n10649), .A(n10608), .B(n10607), .ZN(
        n10665) );
  MUX2_X1 U11355 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n10665), .S(n11171), .Z(
        n10610) );
  INV_X1 U11356 ( .A(n10610), .ZN(n10611) );
  OAI21_X1 U11357 ( .B1(n10668), .B2(n10644), .A(n10611), .ZN(P1_U3545) );
  AOI21_X1 U11358 ( .B1(n10985), .B2(n10613), .A(n10612), .ZN(n10614) );
  OAI211_X1 U11359 ( .C1(n10616), .C2(n10649), .A(n10615), .B(n10614), .ZN(
        n10669) );
  MUX2_X1 U11360 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n10669), .S(n11171), .Z(
        P1_U3544) );
  INV_X1 U11361 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n10620) );
  AOI211_X1 U11362 ( .C1(n10619), .C2(n11168), .A(n10618), .B(n10617), .ZN(
        n10670) );
  MUX2_X1 U11363 ( .A(n10620), .B(n10670), .S(n11171), .Z(n10621) );
  OAI21_X1 U11364 ( .B1(n6707), .B2(n10644), .A(n10621), .ZN(P1_U3543) );
  INV_X1 U11365 ( .A(n10644), .ZN(n10627) );
  OAI211_X1 U11366 ( .C1(n10624), .C2(n10649), .A(n10623), .B(n10622), .ZN(
        n10673) );
  MUX2_X1 U11367 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n10673), .S(n11171), .Z(
        n10625) );
  AOI21_X1 U11368 ( .B1(n10627), .B2(n10626), .A(n10625), .ZN(n10628) );
  INV_X1 U11369 ( .A(n10628), .ZN(P1_U3542) );
  AOI211_X1 U11370 ( .C1(n10631), .C2(n11168), .A(n10630), .B(n10629), .ZN(
        n10677) );
  MUX2_X1 U11371 ( .A(n10632), .B(n10677), .S(n11171), .Z(n10633) );
  OAI21_X1 U11372 ( .B1(n10680), .B2(n10644), .A(n10633), .ZN(P1_U3541) );
  AOI211_X1 U11373 ( .C1(n10985), .C2(n10636), .A(n10635), .B(n10634), .ZN(
        n10637) );
  OAI21_X1 U11374 ( .B1(n10638), .B2(n10649), .A(n10637), .ZN(n10681) );
  MUX2_X1 U11375 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n10681), .S(n11171), .Z(
        P1_U3540) );
  AOI211_X1 U11376 ( .C1(n10641), .C2(n11168), .A(n10640), .B(n10639), .ZN(
        n10682) );
  MUX2_X1 U11377 ( .A(n10642), .B(n10682), .S(n11171), .Z(n10643) );
  OAI21_X1 U11378 ( .B1(n10686), .B2(n10644), .A(n10643), .ZN(P1_U3539) );
  AOI21_X1 U11379 ( .B1(n10985), .B2(n10646), .A(n10645), .ZN(n10647) );
  OAI211_X1 U11380 ( .C1(n10650), .C2(n10649), .A(n10648), .B(n10647), .ZN(
        n10687) );
  MUX2_X1 U11381 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n10687), .S(n11171), .Z(
        P1_U3538) );
  MUX2_X1 U11382 ( .A(n10651), .B(P1_REG1_REG_0__SCAN_IN), .S(n6860), .Z(
        P1_U3522) );
  MUX2_X1 U11383 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n10652), .S(n11175), .Z(
        P1_U3519) );
  INV_X1 U11384 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n10654) );
  MUX2_X1 U11385 ( .A(n10654), .B(n10653), .S(n11175), .Z(n10655) );
  OAI21_X1 U11386 ( .B1(n10656), .B2(n10685), .A(n10655), .ZN(P1_U3517) );
  INV_X1 U11387 ( .A(P1_REG0_REG_26__SCAN_IN), .ZN(n10658) );
  MUX2_X1 U11388 ( .A(n10658), .B(n10657), .S(n11175), .Z(n10659) );
  OAI21_X1 U11389 ( .B1(n10660), .B2(n10685), .A(n10659), .ZN(P1_U3516) );
  INV_X1 U11390 ( .A(P1_REG0_REG_25__SCAN_IN), .ZN(n10662) );
  MUX2_X1 U11391 ( .A(n10662), .B(n10661), .S(n11175), .Z(n10663) );
  OAI21_X1 U11392 ( .B1(n6745), .B2(n10685), .A(n10663), .ZN(P1_U3515) );
  MUX2_X1 U11393 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n10664), .S(n11175), .Z(
        P1_U3514) );
  MUX2_X1 U11394 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n10665), .S(n11175), .Z(
        n10666) );
  INV_X1 U11395 ( .A(n10666), .ZN(n10667) );
  OAI21_X1 U11396 ( .B1(n10668), .B2(n10685), .A(n10667), .ZN(P1_U3513) );
  MUX2_X1 U11397 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n10669), .S(n11175), .Z(
        P1_U3512) );
  INV_X1 U11398 ( .A(P1_REG0_REG_21__SCAN_IN), .ZN(n10671) );
  MUX2_X1 U11399 ( .A(n10671), .B(n10670), .S(n11175), .Z(n10672) );
  OAI21_X1 U11400 ( .B1(n6707), .B2(n10685), .A(n10672), .ZN(P1_U3511) );
  MUX2_X1 U11401 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n10673), .S(n11175), .Z(
        n10674) );
  INV_X1 U11402 ( .A(n10674), .ZN(n10675) );
  OAI21_X1 U11403 ( .B1(n10676), .B2(n10685), .A(n10675), .ZN(P1_U3510) );
  INV_X1 U11404 ( .A(P1_REG0_REG_19__SCAN_IN), .ZN(n10678) );
  MUX2_X1 U11405 ( .A(n10678), .B(n10677), .S(n11175), .Z(n10679) );
  OAI21_X1 U11406 ( .B1(n10680), .B2(n10685), .A(n10679), .ZN(P1_U3509) );
  MUX2_X1 U11407 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n10681), .S(n11175), .Z(
        P1_U3507) );
  INV_X1 U11408 ( .A(P1_REG0_REG_17__SCAN_IN), .ZN(n10683) );
  MUX2_X1 U11409 ( .A(n10683), .B(n10682), .S(n11175), .Z(n10684) );
  OAI21_X1 U11410 ( .B1(n10686), .B2(n10685), .A(n10684), .ZN(P1_U3504) );
  MUX2_X1 U11411 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n10687), .S(n11175), .Z(
        P1_U3501) );
  MUX2_X1 U11412 ( .A(P1_D_REG_1__SCAN_IN), .B(n10690), .S(n10711), .Z(
        P1_U3440) );
  MUX2_X1 U11413 ( .A(P1_D_REG_0__SCAN_IN), .B(n10691), .S(n10711), .Z(
        P1_U3439) );
  NOR4_X1 U11414 ( .A1(n10693), .A2(P1_IR_REG_30__SCAN_IN), .A3(P1_U3086), 
        .A4(n10692), .ZN(n10694) );
  AOI21_X1 U11415 ( .B1(P2_DATAO_REG_31__SCAN_IN), .B2(n10695), .A(n10694), 
        .ZN(n10696) );
  OAI21_X1 U11416 ( .B1(n10697), .B2(n10704), .A(n10696), .ZN(P1_U3324) );
  INV_X1 U11417 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n10698) );
  OAI222_X1 U11418 ( .A1(P1_U3086), .A2(n10700), .B1(n10704), .B2(n10699), 
        .C1(n10698), .C2(n10701), .ZN(P1_U3326) );
  INV_X1 U11419 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n10702) );
  OAI222_X1 U11420 ( .A1(P1_U3086), .A2(n10705), .B1(n10704), .B2(n10703), 
        .C1(n10702), .C2(n10701), .ZN(P1_U3327) );
  INV_X1 U11421 ( .A(n10706), .ZN(n10707) );
  MUX2_X1 U11422 ( .A(n10707), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  NOR2_X1 U11423 ( .A1(n10711), .A2(n10708), .ZN(P1_U3323) );
  NOR2_X1 U11424 ( .A1(n10711), .A2(n10709), .ZN(P1_U3322) );
  NOR2_X1 U11425 ( .A1(n10711), .A2(n10710), .ZN(P1_U3321) );
  AND2_X1 U11426 ( .A1(n10712), .A2(P1_D_REG_5__SCAN_IN), .ZN(P1_U3320) );
  AND2_X1 U11427 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n10712), .ZN(P1_U3319) );
  AND2_X1 U11428 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n10712), .ZN(P1_U3318) );
  AND2_X1 U11429 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n10712), .ZN(P1_U3317) );
  AND2_X1 U11430 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n10712), .ZN(P1_U3316) );
  AND2_X1 U11431 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n10712), .ZN(P1_U3315) );
  AND2_X1 U11432 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n10712), .ZN(P1_U3314) );
  AND2_X1 U11433 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n10712), .ZN(P1_U3313) );
  AND2_X1 U11434 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n10712), .ZN(P1_U3312) );
  AND2_X1 U11435 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n10712), .ZN(P1_U3311) );
  AND2_X1 U11436 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n10712), .ZN(P1_U3310) );
  AND2_X1 U11437 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n10712), .ZN(P1_U3309) );
  AND2_X1 U11438 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n10712), .ZN(P1_U3308) );
  AND2_X1 U11439 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n10712), .ZN(P1_U3307) );
  AND2_X1 U11440 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n10712), .ZN(P1_U3306) );
  AND2_X1 U11441 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n10712), .ZN(P1_U3305) );
  AND2_X1 U11442 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n10712), .ZN(P1_U3304) );
  AND2_X1 U11443 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n10712), .ZN(P1_U3303) );
  AND2_X1 U11444 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n10712), .ZN(P1_U3302) );
  AND2_X1 U11445 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n10712), .ZN(P1_U3301) );
  AND2_X1 U11446 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n10712), .ZN(P1_U3300) );
  AND2_X1 U11447 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n10712), .ZN(P1_U3299) );
  AND2_X1 U11448 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n10712), .ZN(P1_U3298) );
  AND2_X1 U11449 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n10712), .ZN(P1_U3297) );
  AND2_X1 U11450 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n10712), .ZN(P1_U3296) );
  AND2_X1 U11451 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n10712), .ZN(P1_U3295) );
  AND2_X1 U11452 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n10712), .ZN(P1_U3294) );
  NAND2_X1 U11453 ( .A1(P2_ADDR_REG_0__SCAN_IN), .A2(P1_ADDR_REG_0__SCAN_IN), 
        .ZN(n10716) );
  OAI21_X1 U11454 ( .B1(P2_ADDR_REG_0__SCAN_IN), .B2(P1_ADDR_REG_0__SCAN_IN), 
        .A(n10716), .ZN(n10713) );
  INV_X1 U11455 ( .A(n10713), .ZN(ADD_1068_U46) );
  INV_X1 U11456 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n10714) );
  NAND2_X1 U11457 ( .A1(n10714), .A2(n10716), .ZN(n10717) );
  OAI21_X1 U11458 ( .B1(n10714), .B2(n10716), .A(n10717), .ZN(n10715) );
  INV_X1 U11459 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n10892) );
  XOR2_X1 U11460 ( .A(n10715), .B(n10892), .Z(ADD_1068_U5) );
  INV_X1 U11461 ( .A(n10716), .ZN(n10718) );
  AOI22_X1 U11462 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(n10718), .B1(
        P2_ADDR_REG_1__SCAN_IN), .B2(n10717), .ZN(n10721) );
  NAND2_X1 U11463 ( .A1(P1_ADDR_REG_2__SCAN_IN), .A2(P2_ADDR_REG_2__SCAN_IN), 
        .ZN(n10719) );
  OAI21_X1 U11464 ( .B1(P1_ADDR_REG_2__SCAN_IN), .B2(P2_ADDR_REG_2__SCAN_IN), 
        .A(n10719), .ZN(n10720) );
  NOR2_X1 U11465 ( .A1(n10721), .A2(n10720), .ZN(n10722) );
  AOI21_X1 U11466 ( .B1(n10721), .B2(n10720), .A(n10722), .ZN(ADD_1068_U54) );
  AOI21_X1 U11467 ( .B1(P2_ADDR_REG_2__SCAN_IN), .B2(P1_ADDR_REG_2__SCAN_IN), 
        .A(n10722), .ZN(n10725) );
  NAND2_X1 U11468 ( .A1(P2_ADDR_REG_3__SCAN_IN), .A2(P1_ADDR_REG_3__SCAN_IN), 
        .ZN(n10723) );
  OAI21_X1 U11469 ( .B1(P2_ADDR_REG_3__SCAN_IN), .B2(P1_ADDR_REG_3__SCAN_IN), 
        .A(n10723), .ZN(n10724) );
  NOR2_X1 U11470 ( .A1(n10725), .A2(n10724), .ZN(n10726) );
  AOI21_X1 U11471 ( .B1(n10725), .B2(n10724), .A(n10726), .ZN(ADD_1068_U53) );
  AOI21_X1 U11472 ( .B1(P1_ADDR_REG_3__SCAN_IN), .B2(P2_ADDR_REG_3__SCAN_IN), 
        .A(n10726), .ZN(n10729) );
  NOR2_X1 U11473 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n10727) );
  AOI21_X1 U11474 ( .B1(P2_ADDR_REG_4__SCAN_IN), .B2(P1_ADDR_REG_4__SCAN_IN), 
        .A(n10727), .ZN(n10728) );
  NAND2_X1 U11475 ( .A1(n10729), .A2(n10728), .ZN(n10731) );
  OAI21_X1 U11476 ( .B1(n10729), .B2(n10728), .A(n10731), .ZN(ADD_1068_U52) );
  NOR2_X1 U11477 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(P1_ADDR_REG_5__SCAN_IN), 
        .ZN(n10730) );
  AOI21_X1 U11478 ( .B1(P1_ADDR_REG_5__SCAN_IN), .B2(P2_ADDR_REG_5__SCAN_IN), 
        .A(n10730), .ZN(n10733) );
  OAI21_X1 U11479 ( .B1(P1_ADDR_REG_4__SCAN_IN), .B2(P2_ADDR_REG_4__SCAN_IN), 
        .A(n10731), .ZN(n10732) );
  NAND2_X1 U11480 ( .A1(n10733), .A2(n10732), .ZN(n10735) );
  OAI21_X1 U11481 ( .B1(n10733), .B2(n10732), .A(n10735), .ZN(ADD_1068_U51) );
  NOR2_X1 U11482 ( .A1(P2_ADDR_REG_6__SCAN_IN), .A2(P1_ADDR_REG_6__SCAN_IN), 
        .ZN(n10734) );
  AOI21_X1 U11483 ( .B1(P1_ADDR_REG_6__SCAN_IN), .B2(P2_ADDR_REG_6__SCAN_IN), 
        .A(n10734), .ZN(n10737) );
  OAI21_X1 U11484 ( .B1(P2_ADDR_REG_5__SCAN_IN), .B2(P1_ADDR_REG_5__SCAN_IN), 
        .A(n10735), .ZN(n10736) );
  NAND2_X1 U11485 ( .A1(n10737), .A2(n10736), .ZN(n10739) );
  OAI21_X1 U11486 ( .B1(n10737), .B2(n10736), .A(n10739), .ZN(ADD_1068_U50) );
  NOR2_X1 U11487 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(P1_ADDR_REG_7__SCAN_IN), 
        .ZN(n10738) );
  AOI21_X1 U11488 ( .B1(P1_ADDR_REG_7__SCAN_IN), .B2(P2_ADDR_REG_7__SCAN_IN), 
        .A(n10738), .ZN(n10741) );
  OAI21_X1 U11489 ( .B1(P2_ADDR_REG_6__SCAN_IN), .B2(P1_ADDR_REG_6__SCAN_IN), 
        .A(n10739), .ZN(n10740) );
  NAND2_X1 U11490 ( .A1(n10741), .A2(n10740), .ZN(n10743) );
  OAI21_X1 U11491 ( .B1(n10741), .B2(n10740), .A(n10743), .ZN(ADD_1068_U49) );
  NOR2_X1 U11492 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(P1_ADDR_REG_8__SCAN_IN), 
        .ZN(n10742) );
  AOI21_X1 U11493 ( .B1(P1_ADDR_REG_8__SCAN_IN), .B2(P2_ADDR_REG_8__SCAN_IN), 
        .A(n10742), .ZN(n10745) );
  OAI21_X1 U11494 ( .B1(P2_ADDR_REG_7__SCAN_IN), .B2(P1_ADDR_REG_7__SCAN_IN), 
        .A(n10743), .ZN(n10744) );
  NAND2_X1 U11495 ( .A1(n10745), .A2(n10744), .ZN(n10747) );
  OAI21_X1 U11496 ( .B1(n10745), .B2(n10744), .A(n10747), .ZN(ADD_1068_U48) );
  NOR2_X1 U11497 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(P1_ADDR_REG_9__SCAN_IN), 
        .ZN(n10746) );
  AOI21_X1 U11498 ( .B1(P1_ADDR_REG_9__SCAN_IN), .B2(P2_ADDR_REG_9__SCAN_IN), 
        .A(n10746), .ZN(n10749) );
  OAI21_X1 U11499 ( .B1(P2_ADDR_REG_8__SCAN_IN), .B2(P1_ADDR_REG_8__SCAN_IN), 
        .A(n10747), .ZN(n10748) );
  NAND2_X1 U11500 ( .A1(n10749), .A2(n10748), .ZN(n10751) );
  OAI21_X1 U11501 ( .B1(n10749), .B2(n10748), .A(n10751), .ZN(ADD_1068_U47) );
  NOR2_X1 U11502 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(P1_ADDR_REG_10__SCAN_IN), 
        .ZN(n10750) );
  AOI21_X1 U11503 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(P2_ADDR_REG_10__SCAN_IN), 
        .A(n10750), .ZN(n10753) );
  OAI21_X1 U11504 ( .B1(P2_ADDR_REG_9__SCAN_IN), .B2(P1_ADDR_REG_9__SCAN_IN), 
        .A(n10751), .ZN(n10752) );
  NAND2_X1 U11505 ( .A1(n10753), .A2(n10752), .ZN(n10755) );
  OAI21_X1 U11506 ( .B1(n10753), .B2(n10752), .A(n10755), .ZN(ADD_1068_U63) );
  NOR2_X1 U11507 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(P1_ADDR_REG_11__SCAN_IN), 
        .ZN(n10754) );
  AOI21_X1 U11508 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(P2_ADDR_REG_11__SCAN_IN), 
        .A(n10754), .ZN(n10757) );
  OAI21_X1 U11509 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(P1_ADDR_REG_10__SCAN_IN), 
        .A(n10755), .ZN(n10756) );
  NAND2_X1 U11510 ( .A1(n10757), .A2(n10756), .ZN(n10759) );
  OAI21_X1 U11511 ( .B1(n10757), .B2(n10756), .A(n10759), .ZN(ADD_1068_U62) );
  NOR2_X1 U11512 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n10758) );
  AOI21_X1 U11513 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(P2_ADDR_REG_12__SCAN_IN), 
        .A(n10758), .ZN(n10761) );
  OAI21_X1 U11514 ( .B1(P2_ADDR_REG_11__SCAN_IN), .B2(P1_ADDR_REG_11__SCAN_IN), 
        .A(n10759), .ZN(n10760) );
  NAND2_X1 U11515 ( .A1(n10761), .A2(n10760), .ZN(n10763) );
  OAI21_X1 U11516 ( .B1(n10761), .B2(n10760), .A(n10763), .ZN(ADD_1068_U61) );
  NOR2_X1 U11517 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n10762) );
  AOI21_X1 U11518 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(P2_ADDR_REG_13__SCAN_IN), 
        .A(n10762), .ZN(n10765) );
  OAI21_X1 U11519 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(P1_ADDR_REG_12__SCAN_IN), 
        .A(n10763), .ZN(n10764) );
  NAND2_X1 U11520 ( .A1(n10765), .A2(n10764), .ZN(n10767) );
  OAI21_X1 U11521 ( .B1(n10765), .B2(n10764), .A(n10767), .ZN(ADD_1068_U60) );
  NOR2_X1 U11522 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n10766) );
  AOI21_X1 U11523 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(P2_ADDR_REG_14__SCAN_IN), 
        .A(n10766), .ZN(n10769) );
  OAI21_X1 U11524 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(P1_ADDR_REG_13__SCAN_IN), 
        .A(n10767), .ZN(n10768) );
  NAND2_X1 U11525 ( .A1(n10769), .A2(n10768), .ZN(n10771) );
  OAI21_X1 U11526 ( .B1(n10769), .B2(n10768), .A(n10771), .ZN(ADD_1068_U59) );
  NOR2_X1 U11527 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n10770) );
  AOI21_X1 U11528 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(P2_ADDR_REG_15__SCAN_IN), 
        .A(n10770), .ZN(n10773) );
  OAI21_X1 U11529 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(P1_ADDR_REG_14__SCAN_IN), 
        .A(n10771), .ZN(n10772) );
  NAND2_X1 U11530 ( .A1(n10773), .A2(n10772), .ZN(n10775) );
  OAI21_X1 U11531 ( .B1(n10773), .B2(n10772), .A(n10775), .ZN(ADD_1068_U58) );
  NOR2_X1 U11532 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n10774) );
  AOI21_X1 U11533 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(P2_ADDR_REG_16__SCAN_IN), 
        .A(n10774), .ZN(n10777) );
  OAI21_X1 U11534 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(P1_ADDR_REG_15__SCAN_IN), 
        .A(n10775), .ZN(n10776) );
  NAND2_X1 U11535 ( .A1(n10777), .A2(n10776), .ZN(n10779) );
  OAI21_X1 U11536 ( .B1(n10777), .B2(n10776), .A(n10779), .ZN(ADD_1068_U57) );
  NOR2_X1 U11537 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n10778) );
  AOI21_X1 U11538 ( .B1(P1_ADDR_REG_17__SCAN_IN), .B2(P2_ADDR_REG_17__SCAN_IN), 
        .A(n10778), .ZN(n10781) );
  OAI21_X1 U11539 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(P1_ADDR_REG_16__SCAN_IN), 
        .A(n10779), .ZN(n10780) );
  NAND2_X1 U11540 ( .A1(n10781), .A2(n10780), .ZN(n10783) );
  OAI21_X1 U11541 ( .B1(n10781), .B2(n10780), .A(n10783), .ZN(ADD_1068_U56) );
  NOR2_X1 U11542 ( .A1(P2_ADDR_REG_18__SCAN_IN), .A2(P1_ADDR_REG_18__SCAN_IN), 
        .ZN(n10782) );
  AOI21_X1 U11543 ( .B1(P1_ADDR_REG_18__SCAN_IN), .B2(P2_ADDR_REG_18__SCAN_IN), 
        .A(n10782), .ZN(n10785) );
  OAI21_X1 U11544 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(P1_ADDR_REG_17__SCAN_IN), 
        .A(n10783), .ZN(n10784) );
  NAND2_X1 U11545 ( .A1(n10785), .A2(n10784), .ZN(n10786) );
  OAI21_X1 U11546 ( .B1(n10785), .B2(n10784), .A(n10786), .ZN(ADD_1068_U55) );
  OAI21_X1 U11547 ( .B1(P2_ADDR_REG_18__SCAN_IN), .B2(P1_ADDR_REG_18__SCAN_IN), 
        .A(n10786), .ZN(n10788) );
  XOR2_X1 U11548 ( .A(P1_ADDR_REG_19__SCAN_IN), .B(P2_ADDR_REG_19__SCAN_IN), 
        .Z(n10787) );
  XNOR2_X1 U11549 ( .A(n10788), .B(n10787), .ZN(ADD_1068_U4) );
  NAND2_X1 U11550 ( .A1(n10792), .A2(n10789), .ZN(n10791) );
  OAI211_X1 U11551 ( .C1(n10792), .C2(P1_REG2_REG_0__SCAN_IN), .A(n10791), .B(
        n10790), .ZN(n10794) );
  XNOR2_X1 U11552 ( .A(n10794), .B(n10793), .ZN(n10797) );
  AOI22_X1 U11553 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(n10868), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(P1_U3086), .ZN(n10795) );
  OAI21_X1 U11554 ( .B1(n10797), .B2(n10796), .A(n10795), .ZN(P1_U3243) );
  INV_X1 U11555 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n10809) );
  AOI211_X1 U11556 ( .C1(n10800), .C2(n10799), .A(n10798), .B(n10870), .ZN(
        n10805) );
  AOI211_X1 U11557 ( .C1(n10803), .C2(n10802), .A(n10801), .B(n10874), .ZN(
        n10804) );
  AOI211_X1 U11558 ( .C1(n10881), .C2(n10806), .A(n10805), .B(n10804), .ZN(
        n10808) );
  OAI211_X1 U11559 ( .C1(n10885), .C2(n10809), .A(n10808), .B(n10807), .ZN(
        P1_U3254) );
  INV_X1 U11560 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n10821) );
  AOI211_X1 U11561 ( .C1(n10812), .C2(n10811), .A(n10810), .B(n10870), .ZN(
        n10817) );
  AOI211_X1 U11562 ( .C1(n10815), .C2(n10814), .A(n10813), .B(n10874), .ZN(
        n10816) );
  AOI211_X1 U11563 ( .C1(n10881), .C2(n10818), .A(n10817), .B(n10816), .ZN(
        n10820) );
  OAI211_X1 U11564 ( .C1(n10885), .C2(n10821), .A(n10820), .B(n10819), .ZN(
        P1_U3257) );
  INV_X1 U11565 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n10831) );
  AOI211_X1 U11566 ( .C1(n10823), .C2(n11170), .A(n10822), .B(n10874), .ZN(
        n10827) );
  AOI211_X1 U11567 ( .C1(n10825), .C2(n8071), .A(n10824), .B(n10870), .ZN(
        n10826) );
  AOI211_X1 U11568 ( .C1(n10881), .C2(n10828), .A(n10827), .B(n10826), .ZN(
        n10830) );
  OAI211_X1 U11569 ( .C1(n10885), .C2(n10831), .A(n10830), .B(n10829), .ZN(
        P1_U3258) );
  INV_X1 U11570 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n10845) );
  OAI21_X1 U11571 ( .B1(n10834), .B2(n10833), .A(n10832), .ZN(n10842) );
  OAI21_X1 U11572 ( .B1(n10837), .B2(n10836), .A(n10835), .ZN(n10839) );
  AOI222_X1 U11573 ( .A1(n10842), .A2(n10841), .B1(n10840), .B2(n10881), .C1(
        n10839), .C2(n10838), .ZN(n10844) );
  OAI211_X1 U11574 ( .C1(n10885), .C2(n10845), .A(n10844), .B(n10843), .ZN(
        P1_U3260) );
  AOI211_X1 U11575 ( .C1(n10848), .C2(n10847), .A(n10846), .B(n10870), .ZN(
        n10853) );
  AOI211_X1 U11576 ( .C1(n10851), .C2(n10850), .A(n10849), .B(n10874), .ZN(
        n10852) );
  AOI211_X1 U11577 ( .C1(n10858), .C2(n10857), .A(n10856), .B(n10874), .ZN(
        n10863) );
  AOI211_X1 U11578 ( .C1(n10861), .C2(n10860), .A(n10859), .B(n10870), .ZN(
        n10862) );
  AOI211_X1 U11579 ( .C1(n10881), .C2(n10864), .A(n10863), .B(n10862), .ZN(
        n10865) );
  INV_X1 U11580 ( .A(n10865), .ZN(n10867) );
  AOI211_X1 U11581 ( .C1(n10868), .C2(P1_ADDR_REG_13__SCAN_IN), .A(n10867), 
        .B(n10866), .ZN(n10869) );
  INV_X1 U11582 ( .A(n10869), .ZN(P1_U3256) );
  INV_X1 U11583 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n10884) );
  AOI211_X1 U11584 ( .C1(n10873), .C2(n10872), .A(n10871), .B(n10870), .ZN(
        n10879) );
  AOI211_X1 U11585 ( .C1(n10877), .C2(n10876), .A(n10875), .B(n10874), .ZN(
        n10878) );
  AOI211_X1 U11586 ( .C1(n10881), .C2(n10880), .A(n10879), .B(n10878), .ZN(
        n10883) );
  OAI211_X1 U11587 ( .C1(n10885), .C2(n10884), .A(n10883), .B(n10882), .ZN(
        P1_U3253) );
  AOI21_X1 U11588 ( .B1(n5939), .B2(n10887), .A(n10886), .ZN(n10888) );
  NOR2_X1 U11589 ( .A1(n10969), .A2(n10888), .ZN(n10895) );
  AOI21_X1 U11590 ( .B1(n10891), .B2(n10890), .A(n10889), .ZN(n10893) );
  OAI22_X1 U11591 ( .A1(n10974), .A2(n10893), .B1(n10938), .B2(n10892), .ZN(
        n10894) );
  AOI211_X1 U11592 ( .C1(n10941), .C2(n10896), .A(n10895), .B(n10894), .ZN(
        n10901) );
  XOR2_X1 U11593 ( .A(n10898), .B(n10897), .Z(n10899) );
  NAND2_X1 U11594 ( .A1(n10899), .A2(n10962), .ZN(n10900) );
  OAI211_X1 U11595 ( .C1(P2_STATE_REG_SCAN_IN), .C2(n10902), .A(n10901), .B(
        n10900), .ZN(P2_U3183) );
  OAI21_X1 U11596 ( .B1(n10905), .B2(n10904), .A(n10903), .ZN(n10906) );
  AOI22_X1 U11597 ( .A1(n10928), .A2(n10906), .B1(n10965), .B2(
        P2_ADDR_REG_4__SCAN_IN), .ZN(n10921) );
  AOI21_X1 U11598 ( .B1(n10909), .B2(n10908), .A(n10907), .ZN(n10910) );
  NOR2_X1 U11599 ( .A1(n10969), .A2(n10910), .ZN(n10911) );
  AOI211_X1 U11600 ( .C1(n10941), .C2(n10913), .A(n10912), .B(n10911), .ZN(
        n10920) );
  AOI211_X1 U11601 ( .C1(n10917), .C2(n10916), .A(n10915), .B(n10914), .ZN(
        n10918) );
  INV_X1 U11602 ( .A(n10918), .ZN(n10919) );
  NAND3_X1 U11603 ( .A1(n10921), .A2(n10920), .A3(n10919), .ZN(P2_U3186) );
  INV_X1 U11604 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n10939) );
  AOI21_X1 U11605 ( .B1(n10923), .B2(n7262), .A(n10922), .ZN(n10930) );
  OAI21_X1 U11606 ( .B1(n10925), .B2(P2_REG2_REG_5__SCAN_IN), .A(n10924), .ZN(
        n10927) );
  AOI21_X1 U11607 ( .B1(n10928), .B2(n10927), .A(n10926), .ZN(n10929) );
  OAI21_X1 U11608 ( .B1(n10930), .B2(n10969), .A(n10929), .ZN(n10931) );
  AOI21_X1 U11609 ( .B1(n10932), .B2(n10941), .A(n10931), .ZN(n10937) );
  XOR2_X1 U11610 ( .A(n10934), .B(n10933), .Z(n10935) );
  NAND2_X1 U11611 ( .A1(n10935), .A2(n10962), .ZN(n10936) );
  OAI211_X1 U11612 ( .C1(n10939), .C2(n10938), .A(n10937), .B(n10936), .ZN(
        P2_U3187) );
  INV_X1 U11613 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n10957) );
  AOI22_X1 U11614 ( .A1(n10941), .A2(n10940), .B1(n10965), .B2(
        P2_ADDR_REG_17__SCAN_IN), .ZN(n10956) );
  OAI21_X1 U11615 ( .B1(n10944), .B2(n10943), .A(n10942), .ZN(n10954) );
  AOI21_X1 U11616 ( .B1(n9318), .B2(n10946), .A(n10945), .ZN(n10947) );
  NOR2_X1 U11617 ( .A1(n10947), .A2(n10974), .ZN(n10953) );
  INV_X1 U11618 ( .A(n10948), .ZN(n10951) );
  AOI21_X1 U11619 ( .B1(n10951), .B2(n10950), .A(n10969), .ZN(n10952) );
  AOI211_X1 U11620 ( .C1(n10962), .C2(n10954), .A(n10953), .B(n10952), .ZN(
        n10955) );
  OAI211_X1 U11621 ( .C1(P2_STATE_REG_SCAN_IN), .C2(n10957), .A(n10956), .B(
        n10955), .ZN(P2_U3199) );
  INV_X1 U11622 ( .A(n10958), .ZN(n10960) );
  NAND2_X1 U11623 ( .A1(n10960), .A2(n10959), .ZN(n10978) );
  AND3_X1 U11624 ( .A1(n10978), .A2(n10962), .A3(n10961), .ZN(n10963) );
  AOI211_X1 U11625 ( .C1(n10965), .C2(P2_ADDR_REG_18__SCAN_IN), .A(n10964), 
        .B(n10963), .ZN(n10984) );
  AOI21_X1 U11626 ( .B1(n5163), .B2(n10973), .A(n10972), .ZN(n10975) );
  OR2_X1 U11627 ( .A1(n10975), .A2(n10974), .ZN(n10982) );
  OAI21_X1 U11628 ( .B1(n10978), .B2(n10977), .A(n10976), .ZN(n10980) );
  NAND2_X1 U11629 ( .A1(n10980), .A2(n10979), .ZN(n10981) );
  NAND4_X1 U11630 ( .A1(n10984), .A2(n10983), .A3(n10982), .A4(n10981), .ZN(
        P2_U3200) );
  XNOR2_X1 U11631 ( .A(P2_RD_REG_SCAN_IN), .B(P1_RD_REG_SCAN_IN), .ZN(U126) );
  INV_X1 U11632 ( .A(n10985), .ZN(n11165) );
  OAI21_X1 U11633 ( .B1(n10987), .B2(n11165), .A(n10986), .ZN(n10989) );
  AOI211_X1 U11634 ( .C1(n11144), .C2(n10990), .A(n10989), .B(n10988), .ZN(
        n10993) );
  AOI22_X1 U11635 ( .A1(n11171), .A2(n10993), .B1(n10991), .B2(n6860), .ZN(
        P1_U3523) );
  INV_X1 U11636 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n10992) );
  AOI22_X1 U11637 ( .A1(n11175), .A2(n10993), .B1(n10992), .B2(n11172), .ZN(
        P1_U3456) );
  XNOR2_X1 U11638 ( .A(n10994), .B(n10997), .ZN(n11019) );
  OAI211_X1 U11639 ( .C1(n10996), .C2(n11013), .A(n10995), .B(n11126), .ZN(
        n11016) );
  OAI21_X1 U11640 ( .B1(n11013), .B2(n11165), .A(n11016), .ZN(n11007) );
  XNOR2_X1 U11641 ( .A(n10998), .B(n10997), .ZN(n11004) );
  AOI22_X1 U11642 ( .A1(n11002), .A2(n11001), .B1(n11000), .B2(n10999), .ZN(
        n11003) );
  OAI21_X1 U11643 ( .B1(n11004), .B2(n11132), .A(n11003), .ZN(n11005) );
  AOI21_X1 U11644 ( .B1(n11141), .B2(n11019), .A(n11005), .ZN(n11022) );
  INV_X1 U11645 ( .A(n11022), .ZN(n11006) );
  AOI211_X1 U11646 ( .C1(n11144), .C2(n11019), .A(n11007), .B(n11006), .ZN(
        n11010) );
  INV_X1 U11647 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n11008) );
  AOI22_X1 U11648 ( .A1(n11171), .A2(n11010), .B1(n11008), .B2(n6860), .ZN(
        P1_U3524) );
  INV_X1 U11649 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n11009) );
  AOI22_X1 U11650 ( .A1(n11175), .A2(n11010), .B1(n11009), .B2(n11172), .ZN(
        P1_U3459) );
  AOI22_X1 U11651 ( .A1(n11011), .A2(P1_REG2_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(n11149), .ZN(n11012) );
  OAI21_X1 U11652 ( .B1(n11014), .B2(n11013), .A(n11012), .ZN(n11015) );
  INV_X1 U11653 ( .A(n11015), .ZN(n11021) );
  INV_X1 U11654 ( .A(n11016), .ZN(n11017) );
  AOI22_X1 U11655 ( .A1(n11019), .A2(n11156), .B1(n11018), .B2(n11017), .ZN(
        n11020) );
  OAI211_X1 U11656 ( .C1(n11011), .C2(n11022), .A(n11021), .B(n11020), .ZN(
        P1_U3291) );
  AOI22_X1 U11657 ( .A1(n11178), .A2(n11023), .B1(n5957), .B2(n6432), .ZN(
        P2_U3396) );
  INV_X1 U11658 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n11029) );
  OAI22_X1 U11659 ( .A1(n11024), .A2(n11105), .B1(n11104), .B2(n8354), .ZN(
        n11026) );
  AOI211_X1 U11660 ( .C1(n11110), .C2(n11027), .A(n11026), .B(n11025), .ZN(
        n11028) );
  AOI22_X1 U11661 ( .A1(n9488), .A2(n11029), .B1(n11028), .B2(n11111), .ZN(
        P2_U3231) );
  INV_X1 U11662 ( .A(n11030), .ZN(n11035) );
  OAI21_X1 U11663 ( .B1(n11032), .B2(n11165), .A(n11031), .ZN(n11034) );
  AOI211_X1 U11664 ( .C1(n11144), .C2(n11035), .A(n11034), .B(n11033), .ZN(
        n11038) );
  INV_X1 U11665 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n11036) );
  AOI22_X1 U11666 ( .A1(n11171), .A2(n11038), .B1(n11036), .B2(n6860), .ZN(
        P1_U3525) );
  INV_X1 U11667 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n11037) );
  AOI22_X1 U11668 ( .A1(n11175), .A2(n11038), .B1(n11037), .B2(n11172), .ZN(
        P1_U3462) );
  AOI22_X1 U11669 ( .A1(n11178), .A2(n11039), .B1(n5921), .B2(n6432), .ZN(
        P2_U3402) );
  AND2_X1 U11670 ( .A1(n11040), .A2(n11168), .ZN(n11045) );
  OAI21_X1 U11671 ( .B1(n11042), .B2(n11165), .A(n11041), .ZN(n11043) );
  NOR3_X1 U11672 ( .A1(n11045), .A2(n11044), .A3(n11043), .ZN(n11048) );
  INV_X1 U11673 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n11046) );
  AOI22_X1 U11674 ( .A1(n11171), .A2(n11048), .B1(n11046), .B2(n6860), .ZN(
        P1_U3526) );
  INV_X1 U11675 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n11047) );
  AOI22_X1 U11676 ( .A1(n11175), .A2(n11048), .B1(n11047), .B2(n11172), .ZN(
        P1_U3465) );
  INV_X1 U11677 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n11049) );
  AOI22_X1 U11678 ( .A1(n11178), .A2(n11050), .B1(n11049), .B2(n6432), .ZN(
        P2_U3405) );
  AOI22_X1 U11679 ( .A1(n11178), .A2(n11051), .B1(n6006), .B2(n6432), .ZN(
        P2_U3408) );
  OAI21_X1 U11680 ( .B1(n11053), .B2(n11165), .A(n11052), .ZN(n11055) );
  AOI211_X1 U11681 ( .C1(n11144), .C2(n11056), .A(n11055), .B(n11054), .ZN(
        n11059) );
  INV_X1 U11682 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n11057) );
  AOI22_X1 U11683 ( .A1(n11171), .A2(n11059), .B1(n11057), .B2(n6860), .ZN(
        P1_U3528) );
  INV_X1 U11684 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n11058) );
  AOI22_X1 U11685 ( .A1(n11175), .A2(n11059), .B1(n11058), .B2(n11172), .ZN(
        P1_U3471) );
  OAI21_X1 U11686 ( .B1(n11061), .B2(n11165), .A(n11060), .ZN(n11063) );
  AOI211_X1 U11687 ( .C1(n11144), .C2(n11064), .A(n11063), .B(n11062), .ZN(
        n11066) );
  AOI22_X1 U11688 ( .A1(n11171), .A2(n11066), .B1(n7188), .B2(n6860), .ZN(
        P1_U3530) );
  INV_X1 U11689 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n11065) );
  AOI22_X1 U11690 ( .A1(n11175), .A2(n11066), .B1(n11065), .B2(n11172), .ZN(
        P1_U3477) );
  AOI22_X1 U11691 ( .A1(n11178), .A2(n11067), .B1(n6035), .B2(n6432), .ZN(
        P2_U3414) );
  OAI21_X1 U11692 ( .B1(n11069), .B2(n11165), .A(n11068), .ZN(n11071) );
  AOI211_X1 U11693 ( .C1(n11168), .C2(n11072), .A(n11071), .B(n11070), .ZN(
        n11074) );
  AOI22_X1 U11694 ( .A1(n11171), .A2(n11074), .B1(n7446), .B2(n6860), .ZN(
        P1_U3531) );
  INV_X1 U11695 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n11073) );
  AOI22_X1 U11696 ( .A1(n11175), .A2(n11074), .B1(n11073), .B2(n11172), .ZN(
        P1_U3480) );
  OAI211_X1 U11697 ( .C1(n11077), .C2(n11165), .A(n11076), .B(n11075), .ZN(
        n11078) );
  AOI21_X1 U11698 ( .B1(n11079), .B2(n11168), .A(n11078), .ZN(n11081) );
  AOI22_X1 U11699 ( .A1(n11171), .A2(n11081), .B1(n7447), .B2(n6860), .ZN(
        P1_U3532) );
  INV_X1 U11700 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n11080) );
  AOI22_X1 U11701 ( .A1(n11175), .A2(n11081), .B1(n11080), .B2(n11172), .ZN(
        P1_U3483) );
  INV_X1 U11702 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n11082) );
  AOI22_X1 U11703 ( .A1(n11178), .A2(n11083), .B1(n11082), .B2(n6432), .ZN(
        P2_U3420) );
  INV_X1 U11704 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n11084) );
  AOI22_X1 U11705 ( .A1(n11178), .A2(n11085), .B1(n11084), .B2(n6432), .ZN(
        P2_U3423) );
  OAI21_X1 U11706 ( .B1(n11087), .B2(n11165), .A(n11086), .ZN(n11088) );
  AOI21_X1 U11707 ( .B1(n11089), .B2(n11144), .A(n11088), .ZN(n11090) );
  AND2_X1 U11708 ( .A1(n11091), .A2(n11090), .ZN(n11093) );
  AOI22_X1 U11709 ( .A1(n11171), .A2(n11093), .B1(n7448), .B2(n6860), .ZN(
        P1_U3533) );
  INV_X1 U11710 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n11092) );
  AOI22_X1 U11711 ( .A1(n11175), .A2(n11093), .B1(n11092), .B2(n11172), .ZN(
        P1_U3486) );
  OAI211_X1 U11712 ( .C1(n11096), .C2(n11165), .A(n11095), .B(n11094), .ZN(
        n11097) );
  AOI21_X1 U11713 ( .B1(n11098), .B2(n11168), .A(n11097), .ZN(n11101) );
  AOI22_X1 U11714 ( .A1(n11171), .A2(n11101), .B1(n11099), .B2(n6860), .ZN(
        P1_U3534) );
  INV_X1 U11715 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n11100) );
  AOI22_X1 U11716 ( .A1(n11175), .A2(n11101), .B1(n11100), .B2(n11172), .ZN(
        P1_U3489) );
  INV_X1 U11717 ( .A(n11102), .ZN(n11109) );
  INV_X1 U11718 ( .A(n11103), .ZN(n11106) );
  OAI22_X1 U11719 ( .A1(n11106), .A2(n11105), .B1(n5153), .B2(n11104), .ZN(
        n11108) );
  AOI211_X1 U11720 ( .C1(n11110), .C2(n11109), .A(n11108), .B(n11107), .ZN(
        n11112) );
  AOI22_X1 U11721 ( .A1(n9488), .A2(n6120), .B1(n11112), .B2(n11111), .ZN(
        P2_U3220) );
  INV_X1 U11722 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n11113) );
  AOI22_X1 U11723 ( .A1(n11178), .A2(n11114), .B1(n11113), .B2(n6432), .ZN(
        P2_U3429) );
  NAND2_X1 U11724 ( .A1(n7915), .A2(n11115), .ZN(n11117) );
  NAND2_X1 U11725 ( .A1(n11117), .A2(n11116), .ZN(n11119) );
  NAND2_X1 U11726 ( .A1(n11119), .A2(n11118), .ZN(n11121) );
  NAND2_X1 U11727 ( .A1(n11121), .A2(n6624), .ZN(n11122) );
  NAND2_X1 U11728 ( .A1(n11124), .A2(n11152), .ZN(n11125) );
  NAND3_X1 U11729 ( .A1(n11127), .A2(n11126), .A3(n11125), .ZN(n11154) );
  OAI21_X1 U11730 ( .B1(n11128), .B2(n11165), .A(n11154), .ZN(n11143) );
  AOI21_X1 U11731 ( .B1(n11130), .B2(n11129), .A(n6624), .ZN(n11134) );
  INV_X1 U11732 ( .A(n11131), .ZN(n11133) );
  NOR3_X1 U11733 ( .A1(n11134), .A2(n11133), .A3(n11132), .ZN(n11140) );
  OAI22_X1 U11734 ( .A1(n11138), .A2(n11137), .B1(n11136), .B2(n11135), .ZN(
        n11139) );
  AOI211_X1 U11735 ( .C1(n11157), .C2(n11141), .A(n11140), .B(n11139), .ZN(
        n11160) );
  INV_X1 U11736 ( .A(n11160), .ZN(n11142) );
  AOI211_X1 U11737 ( .C1(n11144), .C2(n11157), .A(n11143), .B(n11142), .ZN(
        n11147) );
  AOI22_X1 U11738 ( .A1(n11171), .A2(n11147), .B1(n11145), .B2(n6860), .ZN(
        P1_U3536) );
  INV_X1 U11739 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n11146) );
  AOI22_X1 U11740 ( .A1(n11175), .A2(n11147), .B1(n11146), .B2(n11172), .ZN(
        P1_U3495) );
  INV_X1 U11741 ( .A(n11148), .ZN(n11150) );
  NOR2_X1 U11742 ( .A1(n11154), .A2(n11153), .ZN(n11155) );
  AOI21_X1 U11743 ( .B1(n11157), .B2(n11156), .A(n11155), .ZN(n11158) );
  OAI211_X1 U11744 ( .C1(n11011), .C2(n11160), .A(n11159), .B(n11158), .ZN(
        P1_U3279) );
  AOI22_X1 U11745 ( .A1(n11178), .A2(n11161), .B1(n6143), .B2(n6432), .ZN(
        P2_U3432) );
  AOI22_X1 U11746 ( .A1(n11178), .A2(n11162), .B1(n6160), .B2(n6432), .ZN(
        P2_U3435) );
  OAI211_X1 U11747 ( .C1(n11166), .C2(n11165), .A(n11164), .B(n11163), .ZN(
        n11167) );
  AOI21_X1 U11748 ( .B1(n11169), .B2(n11168), .A(n11167), .ZN(n11174) );
  AOI22_X1 U11749 ( .A1(n11171), .A2(n11174), .B1(n11170), .B2(n6860), .ZN(
        P1_U3537) );
  INV_X1 U11750 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n11173) );
  AOI22_X1 U11751 ( .A1(n11175), .A2(n11174), .B1(n11173), .B2(n11172), .ZN(
        P1_U3498) );
  AOI22_X1 U11752 ( .A1(n11178), .A2(n11176), .B1(n6178), .B2(n6432), .ZN(
        P2_U3438) );
  AOI22_X1 U11753 ( .A1(n11178), .A2(n11177), .B1(n6194), .B2(n6432), .ZN(
        P2_U3441) );
  XNOR2_X1 U11754 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  CLKBUF_X1 U5230 ( .A(n6796), .Z(n9062) );
  OAI211_X1 U6429 ( .C1(n5361), .C2(n10692), .A(n6466), .B(n5359), .ZN(n7144)
         );
endmodule

