

module b22_C_2inp_gates_syn ( P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN, 
        P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN, 
        P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN, 
        P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN, 
        P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN, 
        P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN, 
        P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN, 
        P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN, 
        P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN, 
        P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN, P3_REG3_REG_0__SCAN_IN, 
        P3_REG3_REG_20__SCAN_IN, P3_REG3_REG_13__SCAN_IN, 
        P3_REG3_REG_22__SCAN_IN, P3_REG3_REG_11__SCAN_IN, 
        P3_REG3_REG_2__SCAN_IN, P3_REG3_REG_18__SCAN_IN, 
        P3_REG3_REG_6__SCAN_IN, P3_REG3_REG_26__SCAN_IN, 
        P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_ADDR_REG_0__SCAN_IN, 
        P3_ADDR_REG_1__SCAN_IN, P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN, 
        P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN, P3_ADDR_REG_6__SCAN_IN, 
        P3_ADDR_REG_7__SCAN_IN, P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, 
        P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, 
        P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, 
        P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, 
        P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, 
        P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, 
        P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, 
        P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, 
        P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, 
        P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, 
        P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, 
        P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, 
        P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, 
        P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, 
        P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, 
        P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, 
        P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, 
        P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, 
        P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, 
        P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, 
        P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, 
        P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, 
        P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, 
        P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, 
        P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, 
        P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, 
        P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN, 
        P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN, 
        P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN, 
        P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN, 
        P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN, 
        P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN, 
        P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN, 
        P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN, 
        P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN, 
        P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN, 
        P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN, 
        P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN, 
        P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN, 
        P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN, 
        P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN, 
        P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN, 
        P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN, 
        P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_4__SCAN_IN, 
        P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_17__SCAN_IN, 
        P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_16__SCAN_IN, 
        P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_12__SCAN_IN, 
        P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_1__SCAN_IN, 
        P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_28__SCAN_IN, 
        P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_3__SCAN_IN, 
        P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_23__SCAN_IN, 
        P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_27__SCAN_IN, 
        P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN, P2_RD_REG_SCAN_IN, 
        P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN, P3_IR_REG_1__SCAN_IN, 
        P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN, P3_IR_REG_4__SCAN_IN, 
        P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN, P3_IR_REG_7__SCAN_IN, 
        P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN, P3_IR_REG_10__SCAN_IN, 
        P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN, P3_IR_REG_13__SCAN_IN, 
        P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN, P3_IR_REG_16__SCAN_IN, 
        P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN, P3_IR_REG_19__SCAN_IN, 
        P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN, P3_IR_REG_22__SCAN_IN, 
        P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN, P3_IR_REG_25__SCAN_IN, 
        P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN, P3_IR_REG_28__SCAN_IN, 
        P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN, P3_IR_REG_31__SCAN_IN, 
        P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN, P3_D_REG_2__SCAN_IN, 
        P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN, P3_D_REG_5__SCAN_IN, 
        P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN, P3_D_REG_8__SCAN_IN, 
        P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN, P3_D_REG_11__SCAN_IN, 
        P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN, P3_D_REG_14__SCAN_IN, 
        P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN, P3_D_REG_17__SCAN_IN, 
        P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN, P3_D_REG_20__SCAN_IN, 
        P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN, P3_D_REG_23__SCAN_IN, 
        P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN, P3_D_REG_26__SCAN_IN, 
        P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN, P3_D_REG_29__SCAN_IN, 
        P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN, P3_REG0_REG_0__SCAN_IN, 
        P3_REG0_REG_1__SCAN_IN, P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN, 
        P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN, P3_REG0_REG_6__SCAN_IN, 
        P3_REG0_REG_7__SCAN_IN, P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN, 
        P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN, 
        P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN, 
        P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN, 
        P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN, 
        P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN, 
        P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN, 
        P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN, 
        P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN, 
        P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN, 
        P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN, 
        P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN, 
        P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN, P3_REG1_REG_2__SCAN_IN, 
        P3_REG1_REG_3__SCAN_IN, P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN, 
        P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN, P3_REG1_REG_8__SCAN_IN, 
        P3_REG1_REG_9__SCAN_IN, P3_REG1_REG_10__SCAN_IN, 
        P3_REG1_REG_11__SCAN_IN, P3_REG1_REG_12__SCAN_IN, 
        P3_REG1_REG_13__SCAN_IN, P3_REG1_REG_14__SCAN_IN, 
        P3_REG1_REG_15__SCAN_IN, P3_REG1_REG_16__SCAN_IN, 
        P3_REG1_REG_17__SCAN_IN, P3_REG1_REG_18__SCAN_IN, 
        P3_REG1_REG_19__SCAN_IN, P3_REG1_REG_20__SCAN_IN, 
        P3_REG1_REG_21__SCAN_IN, P3_REG1_REG_22__SCAN_IN, 
        P3_REG1_REG_23__SCAN_IN, P3_REG1_REG_24__SCAN_IN, 
        P3_REG1_REG_25__SCAN_IN, P3_REG1_REG_26__SCAN_IN, 
        P3_REG1_REG_27__SCAN_IN, P3_REG1_REG_28__SCAN_IN, 
        P3_REG1_REG_29__SCAN_IN, P3_REG1_REG_30__SCAN_IN, 
        P3_REG1_REG_31__SCAN_IN, P3_REG2_REG_0__SCAN_IN, 
        P3_REG2_REG_1__SCAN_IN, P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN, 
        P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN, P3_REG2_REG_6__SCAN_IN, 
        P3_REG2_REG_7__SCAN_IN, P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN, 
        P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN, 
        P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN, 
        P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN, 
        P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN, 
        P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN, 
        P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN, 
        P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN, 
        P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN, 
        P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN, 
        P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN, 
        P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN, 
        P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN, 
        P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN, 
        P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN, 
        P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN, 
        P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, SUB_1596_U4, 
        SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65, SUB_1596_U66, 
        SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70, SUB_1596_U54, 
        SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58, SUB_1596_U59, 
        SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53, U29, U28, 
        P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349, 
        P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342, 
        P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335, 
        P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328, 
        P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446, P1_U3323, 
        P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316, 
        P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309, 
        P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302, 
        P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295, 
        P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471, P1_U3474, 
        P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492, P1_U3495, 
        P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513, P1_U3515, 
        P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, 
        P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, 
        P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, 
        P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, 
        P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, 
        P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556, P1_U3557, 
        P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290, P1_U3289, 
        P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282, 
        P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275, 
        P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268, 
        P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, P1_U3262, 
        P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255, 
        P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248, 
        P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560, P1_U3561, 
        P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, 
        P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, 
        P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, 
        P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588, P1_U3589, 
        P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239, P1_U3238, 
        P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231, 
        P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224, 
        P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, 
        P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, P1_U4016, 
        P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321, 
        P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314, 
        P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307, 
        P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300, 
        P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417, P2_U3295, 
        P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, 
        P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, 
        P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, 
        P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, 
        P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442, P2_U3445, 
        P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463, P2_U3466, 
        P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484, P2_U3486, 
        P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492, P2_U3493, 
        P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499, P2_U3500, 
        P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506, P2_U3507, 
        P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, P2_U3514, 
        P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, P2_U3521, 
        P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527, P2_U3528, 
        P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, 
        P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, 
        P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, 
        P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241, P2_U3240, 
        P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, 
        P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, 
        P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, 
        P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531, P2_U3532, 
        P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, 
        P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, 
        P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552, P2_U3553, 
        P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559, P2_U3560, 
        P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211, P2_U3210, 
        P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, 
        P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, 
        P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, 
        P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087, P2_U3947, 
        P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290, P3_U3289, 
        P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283, P3_U3282, 
        P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276, P3_U3275, 
        P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269, P3_U3268, 
        P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377, P3_U3263, 
        P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257, P3_U3256, 
        P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250, P3_U3249, 
        P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243, P3_U3242, 
        P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236, P3_U3235, 
        P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402, P3_U3405, 
        P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423, P3_U3426, 
        P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444, P3_U3446, 
        P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452, P3_U3453, 
        P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459, P3_U3460, 
        P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466, P3_U3467, 
        P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473, P3_U3474, 
        P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480, P3_U3481, 
        P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487, P3_U3488, 
        P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230, P3_U3229, 
        P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223, P3_U3222, 
        P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216, P3_U3215, 
        P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209, P3_U3208, 
        P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202, P3_U3201, 
        P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195, P3_U3194, 
        P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188, P3_U3187, 
        P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491, P3_U3492, 
        P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498, P3_U3499, 
        P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505, P3_U3506, 
        P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512, P3_U3513, 
        P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519, P3_U3520, 
        P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179, P3_U3178, 
        P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172, P3_U3171, 
        P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165, P3_U3164, 
        P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158, P3_U3157, 
        P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150, P3_U3897, 
        keyinput127, keyinput126, keyinput125, keyinput124, keyinput123, 
        keyinput122, keyinput121, keyinput120, keyinput119, keyinput118, 
        keyinput117, keyinput116, keyinput115, keyinput114, keyinput113, 
        keyinput112, keyinput111, keyinput110, keyinput109, keyinput108, 
        keyinput107, keyinput106, keyinput105, keyinput104, keyinput103, 
        keyinput102, keyinput101, keyinput100, keyinput99, keyinput98, 
        keyinput97, keyinput96, keyinput95, keyinput94, keyinput93, keyinput92, 
        keyinput91, keyinput90, keyinput89, keyinput88, keyinput87, keyinput86, 
        keyinput85, keyinput84, keyinput83, keyinput82, keyinput81, keyinput80, 
        keyinput79, keyinput78, keyinput77, keyinput76, keyinput75, keyinput74, 
        keyinput73, keyinput72, keyinput71, keyinput70, keyinput69, keyinput68, 
        keyinput67, keyinput66, keyinput65, keyinput64, keyinput63, keyinput62, 
        keyinput61, keyinput60, keyinput59, keyinput58, keyinput57, keyinput56, 
        keyinput55, keyinput54, keyinput53, keyinput52, keyinput51, keyinput50, 
        keyinput49, keyinput48, keyinput47, keyinput46, keyinput45, keyinput44, 
        keyinput43, keyinput42, keyinput41, keyinput40, keyinput39, keyinput38, 
        keyinput37, keyinput36, keyinput35, keyinput34, keyinput33, keyinput32, 
        keyinput31, keyinput30, keyinput29, keyinput28, keyinput27, keyinput26, 
        keyinput25, keyinput24, keyinput23, keyinput22, keyinput21, keyinput20, 
        keyinput19, keyinput18, keyinput17, keyinput16, keyinput15, keyinput14, 
        keyinput13, keyinput12, keyinput11, keyinput10, keyinput9, keyinput8, 
        keyinput7, keyinput6, keyinput5, keyinput4, keyinput3, keyinput2, 
        keyinput1, keyinput0 );
  input P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN,
         P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN,
         P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN,
         P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN,
         P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN,
         P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN,
         P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN,
         P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN,
         P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN,
         P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN,
         P3_REG3_REG_0__SCAN_IN, P3_REG3_REG_20__SCAN_IN,
         P3_REG3_REG_13__SCAN_IN, P3_REG3_REG_22__SCAN_IN,
         P3_REG3_REG_11__SCAN_IN, P3_REG3_REG_2__SCAN_IN,
         P3_REG3_REG_18__SCAN_IN, P3_REG3_REG_6__SCAN_IN,
         P3_REG3_REG_26__SCAN_IN, P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN,
         P3_DATAO_REG_31__SCAN_IN, P3_DATAO_REG_30__SCAN_IN,
         P3_DATAO_REG_29__SCAN_IN, P3_DATAO_REG_28__SCAN_IN,
         P3_DATAO_REG_27__SCAN_IN, P3_DATAO_REG_26__SCAN_IN,
         P3_DATAO_REG_25__SCAN_IN, P3_DATAO_REG_24__SCAN_IN,
         P3_DATAO_REG_23__SCAN_IN, P3_DATAO_REG_22__SCAN_IN,
         P3_DATAO_REG_21__SCAN_IN, P3_DATAO_REG_20__SCAN_IN,
         P3_DATAO_REG_19__SCAN_IN, P3_DATAO_REG_18__SCAN_IN,
         P3_DATAO_REG_17__SCAN_IN, P3_DATAO_REG_16__SCAN_IN,
         P3_DATAO_REG_15__SCAN_IN, P3_DATAO_REG_14__SCAN_IN,
         P3_DATAO_REG_13__SCAN_IN, P3_DATAO_REG_12__SCAN_IN,
         P3_DATAO_REG_11__SCAN_IN, P3_DATAO_REG_10__SCAN_IN,
         P3_DATAO_REG_9__SCAN_IN, P3_DATAO_REG_8__SCAN_IN,
         P3_DATAO_REG_7__SCAN_IN, P3_DATAO_REG_6__SCAN_IN,
         P3_DATAO_REG_5__SCAN_IN, P3_DATAO_REG_4__SCAN_IN,
         P3_DATAO_REG_3__SCAN_IN, P3_DATAO_REG_2__SCAN_IN,
         P3_DATAO_REG_1__SCAN_IN, P3_DATAO_REG_0__SCAN_IN,
         P3_ADDR_REG_0__SCAN_IN, P3_ADDR_REG_1__SCAN_IN,
         P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN,
         P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN,
         P3_ADDR_REG_6__SCAN_IN, P3_ADDR_REG_7__SCAN_IN,
         P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, P1_IR_REG_0__SCAN_IN,
         P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN,
         P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN,
         P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN,
         P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN,
         P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN,
         P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN,
         P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN,
         P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN,
         P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN,
         P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN,
         P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN,
         P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN,
         P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN,
         P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN,
         P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN,
         P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN,
         P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN,
         P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN,
         P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN,
         P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN,
         P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN,
         P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN,
         P2_RD_REG_SCAN_IN, P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN,
         P3_IR_REG_1__SCAN_IN, P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN,
         P3_IR_REG_4__SCAN_IN, P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN,
         P3_IR_REG_7__SCAN_IN, P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN,
         P3_IR_REG_10__SCAN_IN, P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN,
         P3_IR_REG_13__SCAN_IN, P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN,
         P3_IR_REG_16__SCAN_IN, P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN,
         P3_IR_REG_19__SCAN_IN, P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN,
         P3_IR_REG_22__SCAN_IN, P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN,
         P3_IR_REG_25__SCAN_IN, P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN,
         P3_IR_REG_28__SCAN_IN, P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN,
         P3_IR_REG_31__SCAN_IN, P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN,
         P3_D_REG_2__SCAN_IN, P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN,
         P3_D_REG_5__SCAN_IN, P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN,
         P3_D_REG_8__SCAN_IN, P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN,
         P3_D_REG_11__SCAN_IN, P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN,
         P3_D_REG_14__SCAN_IN, P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN,
         P3_D_REG_17__SCAN_IN, P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN,
         P3_D_REG_20__SCAN_IN, P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN,
         P3_D_REG_23__SCAN_IN, P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN,
         P3_D_REG_26__SCAN_IN, P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN,
         P3_D_REG_29__SCAN_IN, P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN,
         P3_REG0_REG_0__SCAN_IN, P3_REG0_REG_1__SCAN_IN,
         P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN,
         P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN,
         P3_REG0_REG_6__SCAN_IN, P3_REG0_REG_7__SCAN_IN,
         P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN,
         P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN,
         P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN,
         P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN,
         P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN,
         P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN,
         P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN,
         P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN,
         P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN,
         P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN,
         P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN,
         P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN,
         P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN,
         P3_REG1_REG_2__SCAN_IN, P3_REG1_REG_3__SCAN_IN,
         P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN,
         P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN,
         P3_REG1_REG_8__SCAN_IN, P3_REG1_REG_9__SCAN_IN,
         P3_REG1_REG_10__SCAN_IN, P3_REG1_REG_11__SCAN_IN,
         P3_REG1_REG_12__SCAN_IN, P3_REG1_REG_13__SCAN_IN,
         P3_REG1_REG_14__SCAN_IN, P3_REG1_REG_15__SCAN_IN,
         P3_REG1_REG_16__SCAN_IN, P3_REG1_REG_17__SCAN_IN,
         P3_REG1_REG_18__SCAN_IN, P3_REG1_REG_19__SCAN_IN,
         P3_REG1_REG_20__SCAN_IN, P3_REG1_REG_21__SCAN_IN,
         P3_REG1_REG_22__SCAN_IN, P3_REG1_REG_23__SCAN_IN,
         P3_REG1_REG_24__SCAN_IN, P3_REG1_REG_25__SCAN_IN,
         P3_REG1_REG_26__SCAN_IN, P3_REG1_REG_27__SCAN_IN,
         P3_REG1_REG_28__SCAN_IN, P3_REG1_REG_29__SCAN_IN,
         P3_REG1_REG_30__SCAN_IN, P3_REG1_REG_31__SCAN_IN,
         P3_REG2_REG_0__SCAN_IN, P3_REG2_REG_1__SCAN_IN,
         P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN,
         P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN,
         P3_REG2_REG_6__SCAN_IN, P3_REG2_REG_7__SCAN_IN,
         P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN,
         P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN,
         P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN,
         P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN,
         P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN,
         P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN,
         P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN,
         P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN,
         P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN,
         P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN,
         P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN,
         P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN,
         P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN,
         P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN,
         P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN,
         P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN,
         P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, keyinput127,
         keyinput126, keyinput125, keyinput124, keyinput123, keyinput122,
         keyinput121, keyinput120, keyinput119, keyinput118, keyinput117,
         keyinput116, keyinput115, keyinput114, keyinput113, keyinput112,
         keyinput111, keyinput110, keyinput109, keyinput108, keyinput107,
         keyinput106, keyinput105, keyinput104, keyinput103, keyinput102,
         keyinput101, keyinput100, keyinput99, keyinput98, keyinput97,
         keyinput96, keyinput95, keyinput94, keyinput93, keyinput92,
         keyinput91, keyinput90, keyinput89, keyinput88, keyinput87,
         keyinput86, keyinput85, keyinput84, keyinput83, keyinput82,
         keyinput81, keyinput80, keyinput79, keyinput78, keyinput77,
         keyinput76, keyinput75, keyinput74, keyinput73, keyinput72,
         keyinput71, keyinput70, keyinput69, keyinput68, keyinput67,
         keyinput66, keyinput65, keyinput64, keyinput63, keyinput62,
         keyinput61, keyinput60, keyinput59, keyinput58, keyinput57,
         keyinput56, keyinput55, keyinput54, keyinput53, keyinput52,
         keyinput51, keyinput50, keyinput49, keyinput48, keyinput47,
         keyinput46, keyinput45, keyinput44, keyinput43, keyinput42,
         keyinput41, keyinput40, keyinput39, keyinput38, keyinput37,
         keyinput36, keyinput35, keyinput34, keyinput33, keyinput32,
         keyinput31, keyinput30, keyinput29, keyinput28, keyinput27,
         keyinput26, keyinput25, keyinput24, keyinput23, keyinput22,
         keyinput21, keyinput20, keyinput19, keyinput18, keyinput17,
         keyinput16, keyinput15, keyinput14, keyinput13, keyinput12,
         keyinput11, keyinput10, keyinput9, keyinput8, keyinput7, keyinput6,
         keyinput5, keyinput4, keyinput3, keyinput2, keyinput1, keyinput0;
  output SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65,
         SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70,
         SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58,
         SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53,
         U29, U28, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350,
         P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343,
         P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336,
         P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329,
         P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446,
         P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317,
         P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310,
         P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303,
         P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296,
         P1_U3295, P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471,
         P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492,
         P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556,
         P1_U3557, P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290,
         P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283,
         P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276,
         P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269,
         P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263,
         P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256,
         P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249,
         P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588,
         P1_U3589, P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239,
         P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232,
         P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085,
         P1_U4016, P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322,
         P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315,
         P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308,
         P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301,
         P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417,
         P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289,
         P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282,
         P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275,
         P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268,
         P2_U3267, P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442,
         P2_U3445, P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463,
         P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484,
         P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492,
         P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499,
         P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506,
         P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513,
         P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520,
         P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527,
         P2_U3528, P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262,
         P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255,
         P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248,
         P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241,
         P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234,
         P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227,
         P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220,
         P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531,
         P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538,
         P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545,
         P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552,
         P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559,
         P2_U3560, P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204,
         P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197,
         P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190,
         P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087,
         P2_U3947, P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290,
         P3_U3289, P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283,
         P3_U3282, P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276,
         P3_U3275, P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269,
         P3_U3268, P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377,
         P3_U3263, P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257,
         P3_U3256, P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250,
         P3_U3249, P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243,
         P3_U3242, P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236,
         P3_U3235, P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402,
         P3_U3405, P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423,
         P3_U3426, P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444,
         P3_U3446, P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452,
         P3_U3453, P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459,
         P3_U3460, P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466,
         P3_U3467, P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473,
         P3_U3474, P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480,
         P3_U3481, P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487,
         P3_U3488, P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230,
         P3_U3229, P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223,
         P3_U3222, P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216,
         P3_U3215, P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209,
         P3_U3208, P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202,
         P3_U3201, P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195,
         P3_U3194, P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188,
         P3_U3187, P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491,
         P3_U3492, P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498,
         P3_U3499, P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505,
         P3_U3506, P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512,
         P3_U3513, P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519,
         P3_U3520, P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179,
         P3_U3178, P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172,
         P3_U3171, P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165,
         P3_U3164, P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158,
         P3_U3157, P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150,
         P3_U3897;
  wire   n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531,
         n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541,
         n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551,
         n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561,
         n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571,
         n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581,
         n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591,
         n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601,
         n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611,
         n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621,
         n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631,
         n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641,
         n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651,
         n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661,
         n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671,
         n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681,
         n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691,
         n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701,
         n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711,
         n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721,
         n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731,
         n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741,
         n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751,
         n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761,
         n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771,
         n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781,
         n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791,
         n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801,
         n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811,
         n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821,
         n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831,
         n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841,
         n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851,
         n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861,
         n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871,
         n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881,
         n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891,
         n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901,
         n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911,
         n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921,
         n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931,
         n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941,
         n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951,
         n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961,
         n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971,
         n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981,
         n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991,
         n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001,
         n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011,
         n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021,
         n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031,
         n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041,
         n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051,
         n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061,
         n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071,
         n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081,
         n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091,
         n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101,
         n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111,
         n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121,
         n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131,
         n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141,
         n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151,
         n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161,
         n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171,
         n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181,
         n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191,
         n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201,
         n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211,
         n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221,
         n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231,
         n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241,
         n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251,
         n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261,
         n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271,
         n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281,
         n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291,
         n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301,
         n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311,
         n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321,
         n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331,
         n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341,
         n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351,
         n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361,
         n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371,
         n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381,
         n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391,
         n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401,
         n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411,
         n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421,
         n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431,
         n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443,
         n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453,
         n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463,
         n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473,
         n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483,
         n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493,
         n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503,
         n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513,
         n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523,
         n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533,
         n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543,
         n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553,
         n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563,
         n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573,
         n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583,
         n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593,
         n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603,
         n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613,
         n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623,
         n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633,
         n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643,
         n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653,
         n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663,
         n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673,
         n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683,
         n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693,
         n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703,
         n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713,
         n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723,
         n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733,
         n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743,
         n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753,
         n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763,
         n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773,
         n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783,
         n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793,
         n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803,
         n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813,
         n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823,
         n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833,
         n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843,
         n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853,
         n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863,
         n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873,
         n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883,
         n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893,
         n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903,
         n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913,
         n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923,
         n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933,
         n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943,
         n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953,
         n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963,
         n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973,
         n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983,
         n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993,
         n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003,
         n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013,
         n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023,
         n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033,
         n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043,
         n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053,
         n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063,
         n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073,
         n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083,
         n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093,
         n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103,
         n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113,
         n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123,
         n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133,
         n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143,
         n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153,
         n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163,
         n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173,
         n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183,
         n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193,
         n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203,
         n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213,
         n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223,
         n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233,
         n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243,
         n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253,
         n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263,
         n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273,
         n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283,
         n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293,
         n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303,
         n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313,
         n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323,
         n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333,
         n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343,
         n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353,
         n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363,
         n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373,
         n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383,
         n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393,
         n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403,
         n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413,
         n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423,
         n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433,
         n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443,
         n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453,
         n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463,
         n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473,
         n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483,
         n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493,
         n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503,
         n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513,
         n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523,
         n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533,
         n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543,
         n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553,
         n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563,
         n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573,
         n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583,
         n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593,
         n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603,
         n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613,
         n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623,
         n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633,
         n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643,
         n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653,
         n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663,
         n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673,
         n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683,
         n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693,
         n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703,
         n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713,
         n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723,
         n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733,
         n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743,
         n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753,
         n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763,
         n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773,
         n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783,
         n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793,
         n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803,
         n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813,
         n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823,
         n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833,
         n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843,
         n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853,
         n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863,
         n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873,
         n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883,
         n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893,
         n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903,
         n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913,
         n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923,
         n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933,
         n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943,
         n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953,
         n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963,
         n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973,
         n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983,
         n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993,
         n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003,
         n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013,
         n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023,
         n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033,
         n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043,
         n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053,
         n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063,
         n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073,
         n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083,
         n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093,
         n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103,
         n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113,
         n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123,
         n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133,
         n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143,
         n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153,
         n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163,
         n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173,
         n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183,
         n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193,
         n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203,
         n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213,
         n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223,
         n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233,
         n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243,
         n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253,
         n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263,
         n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273,
         n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283,
         n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293,
         n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303,
         n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313,
         n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323,
         n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333,
         n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343,
         n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353,
         n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363,
         n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373,
         n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383,
         n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393,
         n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403,
         n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413,
         n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423,
         n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433,
         n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443,
         n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453,
         n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463,
         n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473,
         n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483,
         n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493,
         n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503,
         n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513,
         n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523,
         n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533,
         n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543,
         n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553,
         n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563,
         n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573,
         n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583,
         n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593,
         n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603,
         n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613,
         n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623,
         n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633,
         n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643,
         n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653,
         n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663,
         n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673,
         n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683,
         n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693,
         n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703,
         n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713,
         n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723,
         n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733,
         n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743,
         n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753,
         n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763,
         n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773,
         n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783,
         n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793,
         n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803,
         n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813,
         n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823,
         n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833,
         n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843,
         n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853,
         n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863,
         n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873,
         n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883,
         n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893,
         n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903,
         n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913,
         n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923,
         n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933,
         n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943,
         n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953,
         n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963,
         n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973,
         n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983,
         n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993,
         n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001, n10002,
         n10003, n10004, n10005, n10006, n10007, n10008, n10009, n10010,
         n10011, n10012, n10013, n10014, n10015, n10016, n10017, n10018,
         n10019, n10020, n10021, n10022, n10023, n10024, n10025, n10026,
         n10027, n10028, n10029, n10030, n10031, n10032, n10033, n10034,
         n10035, n10036, n10037, n10038, n10039, n10040, n10041, n10042,
         n10043, n10044, n10045, n10046, n10047, n10048, n10049, n10050,
         n10051, n10052, n10053, n10054, n10055, n10056, n10057, n10058,
         n10059, n10060, n10061, n10062, n10063, n10064, n10065, n10066,
         n10067, n10068, n10069, n10070, n10071, n10072, n10073, n10074,
         n10075, n10076, n10077, n10078, n10079, n10080, n10081, n10082,
         n10083, n10084, n10085, n10086, n10087, n10088, n10089, n10090,
         n10091, n10092, n10093, n10094, n10095, n10096, n10097, n10098,
         n10099, n10100, n10101, n10102, n10103, n10104, n10105, n10106,
         n10107, n10108, n10109, n10110, n10111, n10112, n10113, n10114,
         n10115, n10116, n10117, n10118, n10119, n10120, n10121, n10122,
         n10123, n10124, n10125, n10126, n10127, n10128, n10129, n10130,
         n10131, n10132, n10133, n10134, n10135, n10136, n10137, n10138,
         n10139, n10140, n10141, n10142, n10143, n10144, n10145, n10146,
         n10147, n10148, n10149, n10150, n10151, n10152, n10153, n10154,
         n10155, n10156, n10157, n10158, n10159, n10160, n10161, n10162,
         n10163, n10164, n10165, n10166, n10167, n10168, n10169, n10170,
         n10171, n10172, n10173, n10174, n10175, n10176, n10177, n10178,
         n10179, n10180, n10181, n10182, n10183, n10184, n10185, n10186,
         n10187, n10188, n10189, n10190, n10191, n10192, n10193, n10194,
         n10195, n10196, n10197, n10198, n10199, n10200, n10201, n10202,
         n10203, n10204, n10205, n10206, n10207, n10208, n10209, n10210,
         n10211, n10212, n10213, n10214, n10215, n10216, n10217, n10218,
         n10219, n10220, n10221, n10222, n10223, n10224, n10225, n10226,
         n10227, n10228, n10229, n10230, n10231, n10232, n10233, n10234,
         n10235, n10236, n10237, n10238, n10239, n10240, n10241, n10242,
         n10243, n10244, n10245, n10246, n10247, n10248, n10249, n10250,
         n10251, n10252, n10253, n10254, n10255, n10256, n10257, n10258,
         n10259, n10260, n10261, n10262, n10263, n10264, n10265, n10266,
         n10267, n10268, n10269, n10270, n10271, n10272, n10273, n10274,
         n10275, n10276, n10277, n10278, n10279, n10280, n10281, n10282,
         n10283, n10284, n10285, n10286, n10287, n10288, n10289, n10290,
         n10291, n10292, n10293, n10294, n10295, n10296, n10297, n10298,
         n10299, n10300, n10301, n10302, n10303, n10304, n10305, n10306,
         n10307, n10308, n10309, n10310, n10311, n10312, n10313, n10314,
         n10315, n10316, n10317, n10318, n10319, n10320, n10321, n10322,
         n10323, n10324, n10325, n10326, n10327, n10328, n10329, n10330,
         n10331, n10332, n10333, n10334, n10335, n10336, n10337, n10338,
         n10339, n10340, n10341, n10342, n10343, n10344, n10345, n10346,
         n10347, n10348, n10349, n10350, n10351, n10352, n10353, n10354,
         n10355, n10356, n10357, n10358, n10359, n10360, n10361, n10362,
         n10363, n10364, n10365, n10366, n10367, n10368, n10369, n10370,
         n10371, n10372, n10373, n10374, n10375, n10376, n10377, n10378,
         n10379, n10380, n10381, n10382, n10383, n10384, n10385, n10386,
         n10387, n10388, n10389, n10390, n10391, n10392, n10393, n10394,
         n10395, n10396, n10397, n10398, n10399, n10400, n10401, n10402,
         n10403, n10404, n10405, n10406, n10407, n10408, n10409, n10410,
         n10411, n10412, n10413, n10414, n10415, n10416, n10417, n10418,
         n10419, n10420, n10421, n10422, n10423, n10424, n10425, n10426,
         n10427, n10428, n10429, n10430, n10431, n10432, n10433, n10434,
         n10435, n10436, n10437, n10438, n10439, n10440, n10441, n10442,
         n10443, n10444, n10445, n10446, n10447, n10448, n10449, n10450,
         n10451, n10452, n10453, n10454, n10455, n10456, n10457, n10458,
         n10459, n10460, n10461, n10462, n10463, n10464, n10465, n10466,
         n10467, n10468, n10469, n10470, n10471, n10472, n10473, n10474,
         n10475, n10476, n10477, n10478, n10479, n10480, n10481, n10482,
         n10483, n10484, n10485, n10486, n10487, n10488, n10489, n10490,
         n10491, n10492, n10493, n10494, n10495, n10496, n10497, n10498,
         n10499, n10500, n10501, n10502, n10503, n10504, n10505, n10506,
         n10507, n10508, n10509, n10510, n10511, n10512, n10513, n10514,
         n10515, n10516, n10517, n10518, n10519, n10520, n10521, n10522,
         n10523, n10524, n10525, n10526, n10527, n10528, n10529, n10530,
         n10531, n10532, n10533, n10534, n10535, n10536, n10537, n10538,
         n10539, n10540, n10541, n10542, n10543, n10544, n10545, n10546,
         n10547, n10548, n10549, n10550, n10551, n10552, n10553, n10554,
         n10555, n10556, n10557, n10558, n10559, n10560, n10561, n10562,
         n10563, n10564, n10565, n10566, n10567, n10568, n10569, n10570,
         n10571, n10572, n10573, n10574, n10575, n10576, n10577, n10578,
         n10579, n10580, n10581, n10582, n10583, n10584, n10585, n10586,
         n10587, n10588, n10589, n10590, n10591, n10592, n10593, n10594,
         n10595, n10596, n10597, n10598, n10599, n10600, n10601, n10602,
         n10603, n10604, n10605, n10606, n10607, n10608, n10609, n10610,
         n10611, n10612, n10613, n10614, n10615, n10616, n10617, n10618,
         n10619, n10620, n10621, n10622, n10623, n10624, n10625, n10626,
         n10627, n10628, n10629, n10630, n10631, n10632, n10633, n10634,
         n10635, n10636, n10637, n10638, n10639, n10640, n10641, n10642,
         n10643, n10644, n10645, n10646, n10647, n10648, n10649, n10650,
         n10651, n10652, n10653, n10654, n10655, n10656, n10657, n10658,
         n10659, n10660, n10661, n10662, n10663, n10664, n10665, n10666,
         n10667, n10668, n10669, n10670, n10671, n10672, n10673, n10674,
         n10675, n10676, n10677, n10678, n10679, n10680, n10681, n10682,
         n10683, n10684, n10685, n10686, n10687, n10688, n10689, n10690,
         n10691, n10692, n10693, n10694, n10695, n10696, n10697, n10698,
         n10699, n10700, n10701, n10702, n10703, n10704, n10705, n10706,
         n10707, n10708, n10709, n10710, n10711, n10712, n10713, n10714,
         n10715, n10716, n10717, n10718, n10719, n10720, n10721, n10722,
         n10723, n10724, n10725, n10726, n10727, n10728, n10729, n10730,
         n10731, n10732, n10733, n10734, n10735, n10736, n10737, n10738,
         n10739, n10740, n10741, n10742, n10743, n10744, n10745, n10746,
         n10747, n10748, n10749, n10750, n10751, n10752, n10753, n10754,
         n10755, n10756, n10757, n10758, n10759, n10760, n10761, n10762,
         n10763, n10764, n10765, n10766, n10767, n10768, n10769, n10770,
         n10771, n10772, n10773, n10774, n10775, n10776, n10777, n10778,
         n10779, n10780, n10781, n10782, n10783, n10784, n10785, n10786,
         n10787, n10788, n10789, n10790, n10791, n10792, n10793, n10794,
         n10795, n10796, n10797, n10798, n10799, n10800, n10801, n10802,
         n10803, n10804, n10805, n10806, n10807, n10808, n10809, n10810,
         n10811, n10812, n10813, n10814, n10815, n10816, n10817, n10818,
         n10819, n10820, n10821, n10822, n10823, n10824, n10825, n10826,
         n10827, n10828, n10829, n10830, n10831, n10832, n10833, n10834,
         n10835, n10836, n10837, n10838, n10839, n10840, n10841, n10842,
         n10843, n10844, n10845, n10846, n10847, n10848, n10849, n10850,
         n10851, n10852, n10853, n10854, n10855, n10856, n10857, n10858,
         n10859, n10860, n10861, n10862, n10863, n10864, n10865, n10866,
         n10867, n10868, n10869, n10870, n10871, n10872, n10873, n10874,
         n10875, n10876, n10877, n10878, n10879, n10880, n10881, n10882,
         n10883, n10884, n10885, n10886, n10887, n10888, n10889, n10890,
         n10891, n10892, n10893, n10894, n10895, n10896, n10897, n10898,
         n10899, n10900, n10901, n10902, n10903, n10904, n10905, n10906,
         n10907, n10908, n10909, n10910, n10911, n10912, n10913, n10914,
         n10915, n10916, n10917, n10918, n10919, n10920, n10921, n10922,
         n10923, n10924, n10925, n10926, n10927, n10928, n10929, n10930,
         n10931, n10932, n10933, n10934, n10935, n10936, n10937, n10938,
         n10939, n10940, n10941, n10942, n10943, n10944, n10945, n10946,
         n10947, n10948, n10949, n10950, n10951, n10952, n10953, n10954,
         n10955, n10956, n10957, n10958, n10959, n10960, n10961, n10962,
         n10963, n10964, n10965, n10966, n10967, n10968, n10969, n10970,
         n10971, n10972, n10973, n10974, n10975, n10976, n10977, n10978,
         n10979, n10980, n10981, n10982, n10983, n10984, n10985, n10986,
         n10987, n10988, n10989, n10990, n10991, n10992, n10993, n10994,
         n10995, n10996, n10997, n10998, n10999, n11000, n11001, n11002,
         n11003, n11004, n11005, n11006, n11007, n11008, n11009, n11010,
         n11011, n11012, n11013, n11014, n11015, n11016, n11017, n11018,
         n11019, n11020, n11021, n11022, n11023, n11024, n11025, n11026,
         n11027, n11028, n11029, n11030, n11031, n11032, n11033, n11034,
         n11035, n11036, n11037, n11038, n11039, n11040, n11041, n11042,
         n11043, n11044, n11045, n11046, n11047, n11048, n11049, n11050,
         n11051, n11052, n11053, n11054, n11055, n11056, n11057, n11058,
         n11059, n11060, n11061, n11062, n11063, n11064, n11065, n11066,
         n11067, n11068, n11069, n11070, n11071, n11072, n11073, n11074,
         n11075, n11076, n11077, n11078, n11079, n11080, n11081, n11082,
         n11083, n11084, n11085, n11086, n11087, n11088, n11089, n11090,
         n11091, n11092, n11093, n11094, n11095, n11096, n11097, n11098,
         n11099, n11100, n11101, n11102, n11103, n11104, n11105, n11106,
         n11107, n11108, n11109, n11110, n11111, n11112, n11113, n11114,
         n11115, n11116, n11117, n11118, n11119, n11120, n11121, n11122,
         n11123, n11124, n11125, n11126, n11127, n11128, n11129, n11130,
         n11131, n11132, n11133, n11134, n11135, n11136, n11137, n11138,
         n11139, n11140, n11141, n11142, n11143, n11144, n11145, n11146,
         n11147, n11148, n11149, n11150, n11151, n11152, n11153, n11154,
         n11155, n11156, n11157, n11158, n11159, n11160, n11161, n11162,
         n11163, n11164, n11165, n11166, n11167, n11168, n11169, n11170,
         n11171, n11172, n11173, n11174, n11175, n11176, n11177, n11178,
         n11179, n11180, n11181, n11182, n11183, n11184, n11185, n11186,
         n11187, n11188, n11189, n11190, n11191, n11192, n11193, n11194,
         n11195, n11196, n11197, n11198, n11199, n11200, n11201, n11202,
         n11203, n11204, n11205, n11206, n11207, n11208, n11209, n11210,
         n11211, n11212, n11213, n11214, n11215, n11216, n11217, n11218,
         n11219, n11220, n11221, n11222, n11223, n11224, n11225, n11226,
         n11227, n11228, n11229, n11230, n11231, n11232, n11233, n11234,
         n11235, n11236, n11237, n11238, n11239, n11240, n11241, n11242,
         n11243, n11244, n11245, n11246, n11247, n11248, n11249, n11250,
         n11251, n11252, n11253, n11254, n11255, n11256, n11257, n11258,
         n11259, n11260, n11261, n11262, n11263, n11264, n11265, n11266,
         n11267, n11268, n11269, n11270, n11271, n11272, n11273, n11274,
         n11275, n11276, n11277, n11278, n11279, n11280, n11281, n11282,
         n11283, n11284, n11285, n11286, n11287, n11288, n11289, n11290,
         n11291, n11292, n11293, n11294, n11295, n11296, n11297, n11298,
         n11299, n11300, n11301, n11302, n11303, n11304, n11305, n11306,
         n11307, n11308, n11309, n11310, n11311, n11312, n11313, n11314,
         n11315, n11316, n11317, n11318, n11319, n11320, n11321, n11322,
         n11323, n11324, n11325, n11326, n11327, n11328, n11329, n11330,
         n11331, n11332, n11333, n11334, n11335, n11336, n11337, n11338,
         n11339, n11340, n11341, n11342, n11343, n11344, n11345, n11346,
         n11347, n11348, n11349, n11350, n11351, n11352, n11353, n11354,
         n11355, n11356, n11357, n11358, n11359, n11360, n11361, n11362,
         n11363, n11364, n11365, n11366, n11367, n11368, n11369, n11370,
         n11371, n11372, n11373, n11374, n11375, n11376, n11377, n11378,
         n11379, n11380, n11381, n11382, n11383, n11384, n11385, n11386,
         n11387, n11388, n11389, n11390, n11391, n11392, n11393, n11394,
         n11395, n11396, n11397, n11398, n11399, n11400, n11401, n11402,
         n11403, n11404, n11405, n11406, n11407, n11408, n11409, n11410,
         n11411, n11412, n11413, n11414, n11415, n11416, n11417, n11418,
         n11419, n11420, n11421, n11422, n11423, n11424, n11425, n11426,
         n11427, n11428, n11429, n11430, n11431, n11432, n11433, n11434,
         n11435, n11436, n11437, n11438, n11439, n11440, n11441, n11442,
         n11443, n11444, n11445, n11446, n11447, n11448, n11449, n11450,
         n11451, n11452, n11453, n11454, n11455, n11456, n11457, n11458,
         n11459, n11460, n11461, n11462, n11463, n11464, n11465, n11466,
         n11467, n11468, n11469, n11470, n11471, n11472, n11473, n11474,
         n11475, n11476, n11477, n11478, n11479, n11480, n11481, n11482,
         n11483, n11484, n11485, n11486, n11487, n11488, n11489, n11490,
         n11491, n11492, n11493, n11494, n11495, n11496, n11497, n11498,
         n11499, n11500, n11501, n11502, n11503, n11504, n11505, n11506,
         n11507, n11508, n11509, n11510, n11511, n11512, n11513, n11514,
         n11515, n11516, n11517, n11518, n11519, n11520, n11521, n11522,
         n11523, n11524, n11525, n11526, n11527, n11528, n11529, n11530,
         n11531, n11532, n11533, n11534, n11535, n11536, n11537, n11538,
         n11539, n11540, n11541, n11542, n11543, n11544, n11545, n11546,
         n11547, n11548, n11549, n11550, n11551, n11552, n11553, n11554,
         n11555, n11556, n11557, n11558, n11559, n11560, n11561, n11562,
         n11563, n11564, n11565, n11566, n11567, n11568, n11569, n11570,
         n11571, n11572, n11573, n11574, n11575, n11576, n11577, n11578,
         n11579, n11580, n11581, n11582, n11583, n11584, n11585, n11586,
         n11587, n11588, n11589, n11590, n11591, n11592, n11593, n11594,
         n11595, n11596, n11597, n11598, n11599, n11600, n11601, n11602,
         n11603, n11604, n11605, n11606, n11607, n11608, n11609, n11610,
         n11611, n11612, n11613, n11614, n11615, n11616, n11617, n11618,
         n11619, n11620, n11621, n11622, n11623, n11624, n11625, n11626,
         n11627, n11628, n11629, n11630, n11631, n11632, n11633, n11634,
         n11635, n11636, n11637, n11638, n11639, n11640, n11641, n11642,
         n11643, n11644, n11645, n11646, n11647, n11648, n11649, n11650,
         n11651, n11652, n11653, n11654, n11655, n11656, n11657, n11658,
         n11659, n11660, n11661, n11662, n11663, n11664, n11665, n11666,
         n11667, n11668, n11669, n11670, n11671, n11672, n11673, n11674,
         n11675, n11676, n11677, n11678, n11679, n11680, n11681, n11682,
         n11683, n11684, n11685, n11686, n11687, n11688, n11689, n11690,
         n11691, n11692, n11693, n11694, n11695, n11696, n11697, n11698,
         n11699, n11700, n11701, n11702, n11703, n11704, n11705, n11706,
         n11707, n11708, n11709, n11710, n11711, n11712, n11713, n11714,
         n11715, n11716, n11717, n11718, n11719, n11720, n11721, n11722,
         n11723, n11724, n11725, n11726, n11727, n11728, n11729, n11730,
         n11731, n11732, n11733, n11734, n11735, n11736, n11737, n11738,
         n11739, n11740, n11741, n11742, n11743, n11744, n11745, n11746,
         n11747, n11748, n11749, n11750, n11751, n11752, n11753, n11754,
         n11755, n11756, n11757, n11758, n11759, n11760, n11761, n11762,
         n11763, n11764, n11765, n11766, n11767, n11768, n11769, n11770,
         n11771, n11772, n11773, n11774, n11775, n11776, n11777, n11778,
         n11779, n11780, n11781, n11782, n11783, n11784, n11785, n11786,
         n11787, n11788, n11789, n11790, n11791, n11792, n11793, n11794,
         n11795, n11796, n11797, n11798, n11799, n11800, n11801, n11802,
         n11803, n11804, n11805, n11806, n11807, n11808, n11809, n11810,
         n11811, n11812, n11813, n11814, n11815, n11816, n11817, n11818,
         n11819, n11820, n11821, n11822, n11823, n11824, n11825, n11826,
         n11827, n11828, n11829, n11830, n11831, n11832, n11833, n11834,
         n11835, n11836, n11837, n11838, n11839, n11840, n11841, n11842,
         n11843, n11844, n11845, n11846, n11847, n11848, n11849, n11850,
         n11851, n11852, n11853, n11854, n11855, n11856, n11857, n11858,
         n11859, n11860, n11861, n11862, n11863, n11864, n11865, n11866,
         n11867, n11868, n11869, n11870, n11871, n11872, n11873, n11874,
         n11875, n11876, n11877, n11878, n11879, n11880, n11881, n11882,
         n11883, n11884, n11885, n11886, n11887, n11888, n11889, n11890,
         n11891, n11892, n11893, n11894, n11895, n11896, n11897, n11898,
         n11899, n11900, n11901, n11902, n11903, n11904, n11905, n11906,
         n11907, n11908, n11909, n11910, n11911, n11912, n11913, n11914,
         n11915, n11916, n11917, n11918, n11919, n11920, n11921, n11922,
         n11923, n11924, n11925, n11926, n11927, n11928, n11929, n11930,
         n11931, n11932, n11933, n11934, n11935, n11936, n11937, n11938,
         n11939, n11940, n11941, n11942, n11943, n11944, n11945, n11946,
         n11947, n11948, n11949, n11950, n11951, n11952, n11953, n11954,
         n11955, n11956, n11957, n11958, n11959, n11960, n11961, n11962,
         n11963, n11964, n11965, n11966, n11967, n11968, n11969, n11970,
         n11971, n11972, n11973, n11974, n11975, n11976, n11977, n11978,
         n11979, n11980, n11981, n11982, n11983, n11984, n11985, n11986,
         n11987, n11988, n11989, n11990, n11991, n11992, n11993, n11994,
         n11995, n11996, n11997, n11998, n11999, n12000, n12001, n12002,
         n12003, n12004, n12005, n12006, n12007, n12008, n12009, n12010,
         n12011, n12012, n12013, n12014, n12015, n12016, n12017, n12018,
         n12019, n12020, n12021, n12022, n12023, n12024, n12025, n12026,
         n12027, n12028, n12029, n12030, n12031, n12032, n12033, n12034,
         n12035, n12036, n12037, n12038, n12039, n12040, n12041, n12042,
         n12043, n12044, n12045, n12046, n12047, n12048, n12049, n12050,
         n12051, n12052, n12053, n12054, n12055, n12056, n12057, n12058,
         n12059, n12060, n12061, n12062, n12063, n12064, n12065, n12066,
         n12067, n12068, n12069, n12070, n12071, n12072, n12073, n12074,
         n12075, n12076, n12077, n12078, n12079, n12080, n12081, n12082,
         n12083, n12084, n12085, n12086, n12087, n12088, n12089, n12090,
         n12091, n12092, n12093, n12094, n12095, n12096, n12097, n12098,
         n12099, n12100, n12101, n12102, n12103, n12104, n12105, n12106,
         n12107, n12108, n12109, n12110, n12111, n12112, n12113, n12114,
         n12115, n12116, n12117, n12118, n12119, n12120, n12121, n12122,
         n12123, n12124, n12125, n12126, n12127, n12128, n12129, n12130,
         n12131, n12132, n12133, n12134, n12135, n12136, n12137, n12138,
         n12139, n12140, n12141, n12142, n12143, n12144, n12145, n12146,
         n12147, n12148, n12149, n12150, n12151, n12152, n12153, n12154,
         n12155, n12156, n12157, n12158, n12159, n12160, n12161, n12162,
         n12163, n12164, n12165, n12166, n12167, n12168, n12169, n12170,
         n12171, n12172, n12173, n12174, n12175, n12176, n12177, n12178,
         n12179, n12180, n12181, n12182, n12183, n12184, n12185, n12186,
         n12187, n12188, n12189, n12190, n12191, n12192, n12193, n12194,
         n12195, n12196, n12197, n12198, n12199, n12200, n12201, n12202,
         n12203, n12204, n12205, n12206, n12207, n12208, n12209, n12210,
         n12211, n12212, n12213, n12214, n12215, n12216, n12217, n12218,
         n12219, n12220, n12221, n12222, n12223, n12224, n12225, n12226,
         n12227, n12228, n12229, n12230, n12231, n12232, n12233, n12234,
         n12235, n12236, n12237, n12238, n12239, n12240, n12241, n12242,
         n12243, n12244, n12245, n12246, n12247, n12248, n12249, n12250,
         n12251, n12252, n12253, n12254, n12255, n12256, n12257, n12258,
         n12259, n12260, n12261, n12262, n12263, n12264, n12265, n12266,
         n12267, n12268, n12269, n12270, n12271, n12272, n12273, n12274,
         n12275, n12276, n12277, n12278, n12279, n12280, n12281, n12282,
         n12283, n12284, n12285, n12286, n12287, n12288, n12289, n12290,
         n12291, n12292, n12293, n12294, n12295, n12296, n12297, n12298,
         n12299, n12300, n12301, n12302, n12303, n12304, n12305, n12306,
         n12307, n12308, n12309, n12310, n12311, n12312, n12313, n12314,
         n12315, n12316, n12317, n12318, n12319, n12320, n12321, n12323,
         n12324, n12325, n12326, n12327, n12328, n12329, n12330, n12331,
         n12332, n12333, n12334, n12335, n12336, n12337, n12338, n12339,
         n12340, n12341, n12342, n12343, n12344, n12345, n12346, n12347,
         n12348, n12349, n12350, n12351, n12352, n12353, n12354, n12355,
         n12356, n12357, n12358, n12359, n12360, n12361, n12362, n12363,
         n12364, n12365, n12366, n12367, n12368, n12369, n12370, n12371,
         n12372, n12373, n12374, n12375, n12376, n12377, n12378, n12379,
         n12380, n12381, n12382, n12383, n12384, n12385, n12386, n12387,
         n12388, n12389, n12390, n12391, n12392, n12393, n12394, n12395,
         n12396, n12397, n12398, n12399, n12400, n12401, n12402, n12403,
         n12404, n12405, n12406, n12407, n12408, n12409, n12410, n12411,
         n12412, n12413, n12414, n12415, n12416, n12417, n12418, n12419,
         n12420, n12421, n12422, n12423, n12424, n12425, n12426, n12427,
         n12428, n12429, n12430, n12431, n12432, n12433, n12434, n12435,
         n12436, n12437, n12438, n12439, n12440, n12441, n12442, n12443,
         n12444, n12445, n12446, n12447, n12448, n12449, n12450, n12451,
         n12452, n12453, n12454, n12455, n12456, n12457, n12458, n12459,
         n12460, n12461, n12462, n12463, n12464, n12465, n12466, n12467,
         n12468, n12469, n12470, n12471, n12472, n12473, n12474, n12475,
         n12476, n12477, n12478, n12479, n12480, n12481, n12482, n12483,
         n12484, n12485, n12486, n12487, n12488, n12489, n12490, n12491,
         n12492, n12493, n12494, n12495, n12496, n12497, n12498, n12499,
         n12500, n12501, n12502, n12503, n12504, n12505, n12506, n12507,
         n12508, n12509, n12510, n12511, n12512, n12513, n12514, n12515,
         n12516, n12517, n12518, n12519, n12520, n12521, n12522, n12523,
         n12524, n12525, n12526, n12527, n12528, n12529, n12530, n12531,
         n12532, n12533, n12534, n12535, n12536, n12537, n12538, n12539,
         n12540, n12541, n12542, n12543, n12544, n12545, n12546, n12547,
         n12548, n12549, n12550, n12551, n12552, n12553, n12554, n12555,
         n12556, n12557, n12558, n12559, n12560, n12561, n12562, n12563,
         n12564, n12565, n12566, n12567, n12568, n12569, n12570, n12571,
         n12572, n12573, n12574, n12575, n12576, n12577, n12578, n12579,
         n12580, n12581, n12582, n12583, n12584, n12585, n12586, n12587,
         n12588, n12589, n12590, n12591, n12592, n12593, n12594, n12595,
         n12596, n12597, n12598, n12599, n12600, n12601, n12602, n12603,
         n12604, n12605, n12606, n12607, n12608, n12609, n12610, n12611,
         n12612, n12613, n12614, n12615, n12616, n12617, n12618, n12619,
         n12620, n12621, n12622, n12623, n12624, n12625, n12626, n12627,
         n12628, n12629, n12630, n12631, n12632, n12633, n12634, n12635,
         n12636, n12637, n12638, n12639, n12640, n12641, n12642, n12643,
         n12644, n12645, n12646, n12647, n12648, n12649, n12650, n12651,
         n12652, n12653, n12654, n12655, n12656, n12657, n12658, n12659,
         n12660, n12661, n12662, n12663, n12664, n12665, n12666, n12667,
         n12668, n12669, n12670, n12671, n12672, n12673, n12674, n12675,
         n12676, n12677, n12678, n12679, n12680, n12681, n12682, n12683,
         n12684, n12685, n12686, n12687, n12688, n12689, n12690, n12691,
         n12692, n12693, n12694, n12695, n12696, n12697, n12698, n12699,
         n12700, n12701, n12702, n12703, n12704, n12705, n12706, n12707,
         n12708, n12709, n12710, n12711, n12712, n12713, n12714, n12715,
         n12716, n12717, n12718, n12719, n12720, n12721, n12722, n12723,
         n12724, n12725, n12726, n12727, n12728, n12729, n12730, n12731,
         n12732, n12733, n12734, n12735, n12736, n12737, n12738, n12739,
         n12740, n12741, n12742, n12743, n12744, n12745, n12746, n12747,
         n12748, n12749, n12750, n12751, n12752, n12753, n12754, n12755,
         n12756, n12757, n12758, n12759, n12760, n12761, n12762, n12763,
         n12764, n12765, n12766, n12767, n12768, n12769, n12770, n12771,
         n12772, n12773, n12774, n12775, n12776, n12777, n12778, n12779,
         n12780, n12781, n12782, n12783, n12784, n12785, n12786, n12787,
         n12788, n12789, n12790, n12791, n12792, n12793, n12794, n12795,
         n12796, n12797, n12798, n12799, n12800, n12801, n12802, n12803,
         n12804, n12805, n12806, n12807, n12808, n12809, n12810, n12811,
         n12812, n12813, n12814, n12815, n12816, n12817, n12818, n12819,
         n12820, n12821, n12822, n12823, n12824, n12825, n12826, n12827,
         n12828, n12829, n12830, n12831, n12832, n12833, n12834, n12835,
         n12836, n12837, n12838, n12839, n12840, n12841, n12842, n12843,
         n12844, n12845, n12846, n12847, n12848, n12849, n12850, n12851,
         n12852, n12853, n12854, n12855, n12856, n12857, n12858, n12859,
         n12860, n12861, n12862, n12863, n12864, n12865, n12866, n12867,
         n12868, n12869, n12870, n12871, n12872, n12873, n12874, n12875,
         n12876, n12877, n12878, n12879, n12880, n12881, n12882, n12883,
         n12884, n12885, n12886, n12887, n12888, n12889, n12890, n12891,
         n12892, n12893, n12894, n12895, n12896, n12897, n12898, n12899,
         n12900, n12901, n12902, n12903, n12904, n12905, n12906, n12907,
         n12908, n12909, n12910, n12911, n12912, n12913, n12914, n12915,
         n12916, n12917, n12918, n12919, n12920, n12921, n12922, n12923,
         n12924, n12925, n12926, n12927, n12928, n12929, n12930, n12931,
         n12932, n12933, n12934, n12935, n12936, n12937, n12938, n12939,
         n12940, n12941, n12942, n12943, n12944, n12945, n12946, n12947,
         n12948, n12949, n12950, n12951, n12952, n12953, n12954, n12955,
         n12956, n12957, n12958, n12959, n12960, n12961, n12962, n12963,
         n12964, n12965, n12966, n12967, n12968, n12969, n12970, n12971,
         n12972, n12973, n12974, n12975, n12976, n12977, n12978, n12979,
         n12980, n12981, n12982, n12983, n12984, n12985, n12986, n12987,
         n12988, n12989, n12990, n12991, n12992, n12993, n12994, n12995,
         n12996, n12997, n12998, n12999, n13000, n13001, n13002, n13003,
         n13004, n13005, n13006, n13007, n13008, n13009, n13010, n13011,
         n13012, n13013, n13014, n13015, n13016, n13017, n13018, n13019,
         n13020, n13021, n13022, n13023, n13024, n13025, n13026, n13027,
         n13028, n13029, n13030, n13031, n13032, n13033, n13034, n13035,
         n13036, n13037, n13038, n13039, n13040, n13041, n13042, n13043,
         n13044, n13045, n13046, n13047, n13048, n13049, n13050, n13051,
         n13052, n13053, n13054, n13055, n13056, n13057, n13058, n13059,
         n13060, n13061, n13062, n13063, n13064, n13065, n13066, n13067,
         n13068, n13069, n13070, n13071, n13072, n13073, n13074, n13075,
         n13076, n13077, n13078, n13079, n13080, n13081, n13082, n13083,
         n13084, n13085, n13086, n13087, n13088, n13089, n13090, n13091,
         n13092, n13093, n13094, n13095, n13096, n13097, n13098, n13099,
         n13100, n13101, n13102, n13103, n13104, n13105, n13106, n13107,
         n13108, n13109, n13110, n13111, n13112, n13113, n13114, n13115,
         n13116, n13117, n13118, n13119, n13120, n13121, n13122, n13123,
         n13124, n13125, n13126, n13127, n13128, n13129, n13130, n13131,
         n13132, n13133, n13134, n13135, n13136, n13137, n13138, n13139,
         n13140, n13141, n13142, n13143, n13144, n13145, n13146, n13147,
         n13148, n13149, n13150, n13151, n13152, n13153, n13154, n13155,
         n13156, n13157, n13158, n13159, n13160, n13161, n13162, n13163,
         n13164, n13165, n13166, n13167, n13168, n13169, n13170, n13171,
         n13172, n13173, n13174, n13175, n13176, n13177, n13178, n13179,
         n13180, n13181, n13182, n13183, n13184, n13185, n13186, n13187,
         n13188, n13189, n13190, n13191, n13192, n13193, n13194, n13195,
         n13196, n13197, n13198, n13199, n13200, n13201, n13202, n13203,
         n13204, n13205, n13206, n13207, n13208, n13209, n13210, n13211,
         n13212, n13213, n13214, n13215, n13216, n13217, n13218, n13219,
         n13220, n13221, n13222, n13223, n13224, n13225, n13226, n13227,
         n13228, n13229, n13230, n13231, n13232, n13233, n13234, n13235,
         n13236, n13237, n13238, n13239, n13240, n13241, n13242, n13243,
         n13244, n13245, n13246, n13247, n13248, n13249, n13250, n13251,
         n13252, n13253, n13254, n13255, n13256, n13257, n13258, n13259,
         n13260, n13261, n13262, n13263, n13264, n13265, n13266, n13267,
         n13268, n13269, n13270, n13271, n13272, n13273, n13274, n13275,
         n13276, n13277, n13278, n13279, n13280, n13281, n13282, n13283,
         n13284, n13285, n13286, n13287, n13288, n13289, n13290, n13291,
         n13292, n13293, n13294, n13295, n13296, n13297, n13298, n13299,
         n13300, n13301, n13302, n13303, n13304, n13305, n13306, n13307,
         n13308, n13309, n13310, n13311, n13312, n13313, n13314, n13315,
         n13316, n13317, n13318, n13319, n13320, n13321, n13322, n13323,
         n13324, n13325, n13326, n13327, n13328, n13329, n13330, n13331,
         n13332, n13333, n13334, n13335, n13336, n13337, n13338, n13339,
         n13340, n13341, n13342, n13343, n13344, n13345, n13346, n13347,
         n13348, n13349, n13350, n13351, n13352, n13353, n13354, n13355,
         n13356, n13357, n13358, n13359, n13360, n13361, n13362, n13363,
         n13364, n13365, n13366, n13367, n13368, n13369, n13370, n13371,
         n13372, n13373, n13374, n13375, n13376, n13377, n13378, n13379,
         n13380, n13381, n13382, n13383, n13384, n13385, n13386, n13387,
         n13388, n13389, n13390, n13391, n13392, n13393, n13394, n13395,
         n13396, n13397, n13398, n13399, n13400, n13401, n13402, n13403,
         n13404, n13405, n13406, n13407, n13408, n13409, n13410, n13411,
         n13412, n13413, n13414, n13415, n13416, n13417, n13418, n13419,
         n13420, n13421, n13422, n13423, n13424, n13425, n13426, n13427,
         n13428, n13429, n13430, n13431, n13432, n13433, n13434, n13435,
         n13436, n13437, n13438, n13439, n13440, n13441, n13442, n13443,
         n13444, n13445, n13446, n13447, n13448, n13449, n13450, n13451,
         n13452, n13453, n13454, n13455, n13456, n13457, n13458, n13459,
         n13460, n13461, n13462, n13463, n13464, n13465, n13466, n13467,
         n13468, n13469, n13470, n13471, n13472, n13473, n13474, n13475,
         n13476, n13477, n13478, n13479, n13480, n13481, n13482, n13483,
         n13484, n13485, n13486, n13487, n13488, n13489, n13490, n13491,
         n13492, n13493, n13494, n13495, n13496, n13497, n13498, n13499,
         n13500, n13501, n13502, n13503, n13504, n13505, n13506, n13507,
         n13508, n13509, n13510, n13511, n13512, n13513, n13514, n13515,
         n13516, n13517, n13518, n13519, n13520, n13521, n13522, n13523,
         n13524, n13525, n13526, n13527, n13528, n13529, n13530, n13531,
         n13532, n13533, n13534, n13535, n13536, n13537, n13538, n13539,
         n13540, n13541, n13542, n13543, n13544, n13545, n13546, n13547,
         n13548, n13549, n13550, n13551, n13552, n13553, n13554, n13555,
         n13556, n13557, n13558, n13559, n13560, n13561, n13562, n13563,
         n13564, n13565, n13566, n13567, n13568, n13569, n13570, n13571,
         n13572, n13573, n13574, n13575, n13576, n13577, n13578, n13579,
         n13580, n13581, n13582, n13583, n13584, n13585, n13586, n13587,
         n13588, n13589, n13590, n13591, n13592, n13593, n13594, n13595,
         n13596, n13597, n13598, n13599, n13600, n13601, n13602, n13603,
         n13604, n13605, n13606, n13607, n13608, n13609, n13610, n13611,
         n13612, n13613, n13614, n13615, n13616, n13617, n13618, n13619,
         n13620, n13621, n13622, n13623, n13624, n13625, n13626, n13627,
         n13628, n13629, n13630, n13631, n13632, n13633, n13634, n13635,
         n13636, n13637, n13638, n13639, n13640, n13641, n13642, n13643,
         n13644, n13645, n13646, n13647, n13648, n13649, n13650, n13651,
         n13652, n13653, n13654, n13655, n13656, n13657, n13658, n13659,
         n13660, n13661, n13662, n13663, n13664, n13665, n13666, n13667,
         n13668, n13669, n13670, n13671, n13672, n13673, n13674, n13675,
         n13676, n13677, n13678, n13679, n13680, n13681, n13682, n13683,
         n13684, n13685, n13686, n13687, n13688, n13689, n13690, n13691,
         n13692, n13693, n13694, n13695, n13696, n13697, n13698, n13699,
         n13700, n13701, n13702, n13703, n13704, n13705, n13706, n13707,
         n13708, n13709, n13710, n13711, n13712, n13713, n13714, n13715,
         n13716, n13717, n13718, n13719, n13720, n13721, n13722, n13723,
         n13724, n13725, n13726, n13727, n13728, n13729, n13730, n13731,
         n13732, n13733, n13734, n13735, n13736, n13737, n13738, n13739,
         n13740, n13741, n13742, n13743, n13744, n13745, n13746, n13747,
         n13748, n13749, n13750, n13751, n13752, n13753, n13754, n13755,
         n13756, n13757, n13758, n13759, n13760, n13761, n13762, n13763,
         n13764, n13765, n13766, n13767, n13768, n13769, n13770, n13771,
         n13772, n13773, n13774, n13775, n13776, n13777, n13778, n13779,
         n13780, n13781, n13782, n13783, n13784, n13785, n13786, n13787,
         n13788, n13789, n13790, n13791, n13792, n13793, n13794, n13795,
         n13796, n13797, n13798, n13799, n13800, n13801, n13802, n13803,
         n13804, n13805, n13806, n13807, n13808, n13809, n13810, n13811,
         n13812, n13813, n13814, n13815, n13816, n13817, n13818, n13819,
         n13820, n13821, n13822, n13823, n13824, n13825, n13826, n13827,
         n13828, n13829, n13830, n13831, n13832, n13833, n13834, n13835,
         n13836, n13837, n13838, n13839, n13840, n13841, n13842, n13843,
         n13844, n13845, n13846, n13847, n13848, n13849, n13850, n13851,
         n13852, n13853, n13854, n13855, n13856, n13857, n13858, n13859,
         n13860, n13861, n13862, n13863, n13864, n13865, n13866, n13867,
         n13868, n13869, n13870, n13871, n13872, n13873, n13874, n13875,
         n13876, n13877, n13878, n13879, n13880, n13881, n13882, n13883,
         n13884, n13885, n13886, n13887, n13888, n13889, n13890, n13891,
         n13892, n13893, n13894, n13895, n13896, n13897, n13898, n13899,
         n13900, n13901, n13902, n13903, n13904, n13905, n13906, n13907,
         n13908, n13909, n13910, n13911, n13912, n13913, n13914, n13915,
         n13916, n13917, n13918, n13919, n13920, n13921, n13922, n13923,
         n13924, n13925, n13926, n13927, n13928, n13929, n13930, n13931,
         n13932, n13933, n13934, n13935, n13936, n13937, n13938, n13939,
         n13940, n13941, n13942, n13943, n13944, n13945, n13946, n13947,
         n13948, n13949, n13950, n13951, n13952, n13953, n13954, n13955,
         n13956, n13957, n13958, n13959, n13960, n13961, n13962, n13963,
         n13964, n13965, n13966, n13967, n13968, n13969, n13970, n13971,
         n13972, n13973, n13974, n13975, n13976, n13977, n13978, n13979,
         n13980, n13981, n13982, n13983, n13984, n13985, n13986, n13987,
         n13988, n13989, n13990, n13991, n13992, n13993, n13994, n13995,
         n13996, n13997, n13998, n13999, n14000, n14001, n14002, n14003,
         n14004, n14005, n14006, n14007, n14008, n14009, n14010, n14011,
         n14012, n14013, n14014, n14015, n14016, n14017, n14018, n14019,
         n14020, n14021, n14022, n14023, n14024, n14025, n14026, n14027,
         n14028, n14029, n14030, n14031, n14032, n14033, n14034, n14035,
         n14036, n14037, n14038, n14039, n14040, n14041, n14042, n14043,
         n14044, n14045, n14046, n14047, n14048, n14049, n14050, n14051,
         n14052, n14053, n14054, n14055, n14056, n14057, n14058, n14059,
         n14060, n14061, n14062, n14063, n14064, n14065, n14066, n14067,
         n14068, n14069, n14070, n14071, n14072, n14073, n14074, n14075,
         n14076, n14077, n14078, n14079, n14080, n14081, n14082, n14083,
         n14084, n14085, n14086, n14087, n14088, n14089, n14090, n14091,
         n14092, n14093, n14094, n14095, n14096, n14097, n14098, n14099,
         n14100, n14101, n14102, n14103, n14104, n14105, n14106, n14107,
         n14108, n14109, n14110, n14111, n14112, n14113, n14114, n14115,
         n14116, n14117, n14118, n14119, n14120, n14121, n14122, n14123,
         n14124, n14125, n14126, n14127, n14128, n14129, n14130, n14131,
         n14132, n14133, n14134, n14135, n14136, n14137, n14138, n14139,
         n14140, n14141, n14142, n14143, n14144, n14145, n14146, n14147,
         n14148, n14149, n14150, n14151, n14152, n14153, n14154, n14155,
         n14156, n14157, n14158, n14159, n14160, n14161, n14162, n14163,
         n14164, n14165, n14166, n14167, n14168, n14169, n14170, n14171,
         n14172, n14173, n14174, n14175, n14176, n14177, n14178, n14179,
         n14180, n14181, n14182, n14183, n14184, n14185, n14186, n14187,
         n14188, n14189, n14190, n14191, n14192, n14193, n14194, n14195,
         n14196, n14197, n14198, n14199, n14200, n14201, n14202, n14203,
         n14204, n14205, n14206, n14207, n14208, n14209, n14210, n14211,
         n14212, n14213, n14214, n14215, n14216, n14217, n14218, n14219,
         n14220, n14221, n14222, n14223, n14224, n14225, n14226, n14227,
         n14228, n14229, n14230, n14231, n14232, n14233, n14234, n14235,
         n14236, n14237, n14238, n14239, n14240, n14241, n14242, n14243,
         n14244, n14245, n14246, n14247, n14248, n14249, n14250, n14251,
         n14252, n14253, n14254, n14255, n14256, n14257, n14258, n14259,
         n14260, n14261, n14262, n14263, n14264, n14265, n14266, n14267,
         n14268, n14269, n14270, n14271, n14272, n14273, n14274, n14275,
         n14276, n14277, n14278, n14279, n14280, n14281, n14282, n14283,
         n14284, n14285, n14286, n14287, n14288, n14289, n14290, n14291,
         n14292, n14293, n14294, n14295, n14296, n14297, n14298, n14299,
         n14300, n14301, n14302, n14303, n14304, n14305, n14306, n14307,
         n14308, n14309, n14310, n14311, n14312, n14313, n14314, n14315,
         n14316, n14317, n14318, n14319, n14320, n14321, n14322, n14323,
         n14324, n14325, n14326, n14327, n14328, n14329, n14330, n14331,
         n14332, n14333, n14334, n14335, n14336, n14337, n14338, n14339,
         n14340, n14341, n14342, n14343, n14344, n14345, n14346, n14347,
         n14348, n14349, n14350, n14351, n14352, n14353, n14354, n14355,
         n14356, n14357, n14358, n14359, n14360, n14361, n14362, n14363,
         n14364, n14365, n14366, n14367, n14368, n14369, n14370, n14371,
         n14372, n14373, n14374, n14375, n14376, n14377, n14378, n14379,
         n14380, n14381, n14382, n14383, n14384, n14385, n14386, n14387,
         n14388, n14389, n14390, n14391, n14392, n14393, n14394, n14395,
         n14396, n14397, n14398, n14399, n14400, n14401, n14402, n14403,
         n14404, n14405, n14406, n14407, n14408, n14409, n14410, n14411,
         n14412, n14413, n14414, n14415, n14416, n14417, n14418, n14419,
         n14420, n14421, n14422, n14423, n14424, n14425, n14426, n14427,
         n14428, n14429, n14430, n14431, n14432, n14433, n14434, n14435,
         n14436, n14437, n14438, n14439, n14440, n14441, n14442, n14443,
         n14444, n14445, n14446, n14447, n14448, n14449, n14450, n14451,
         n14452, n14453, n14454, n14455, n14456, n14457, n14458, n14459,
         n14460, n14461, n14462, n14463, n14464, n14465, n14466, n14467,
         n14468, n14469, n14470, n14471, n14472, n14473, n14474, n14475,
         n14476, n14477, n14478, n14479, n14480, n14481, n14482, n14483,
         n14484, n14485, n14486, n14487, n14488, n14489, n14490, n14491,
         n14492, n14493, n14494, n14495, n14496, n14497, n14498, n14499,
         n14500, n14501, n14502, n14503, n14504, n14505, n14506, n14507,
         n14508, n14509, n14510, n14511, n14512, n14513, n14514, n14515,
         n14516, n14517, n14518, n14519, n14520, n14521, n14522, n14523,
         n14524, n14525, n14526, n14527, n14528, n14529, n14530, n14531,
         n14532, n14533, n14534, n14535, n14536, n14537, n14538, n14539,
         n14540, n14541, n14542, n14543, n14544, n14545, n14546, n14547,
         n14548, n14549, n14550, n14551, n14552, n14553, n14554, n14555,
         n14556, n14557, n14558, n14559, n14560, n14561, n14562, n14563,
         n14564, n14565, n14566, n14567, n14568, n14569, n14570, n14571,
         n14572, n14573, n14574, n14575, n14576, n14577, n14578, n14579,
         n14580, n14581, n14582, n14583, n14584, n14585, n14586, n14587,
         n14588, n14589, n14590, n14591, n14592, n14593, n14594, n14595,
         n14596, n14597, n14598, n14599, n14600, n14601, n14602, n14603,
         n14604, n14605, n14606, n14607, n14608, n14609, n14610, n14611,
         n14612, n14613, n14614, n14615, n14616, n14617, n14618, n14619,
         n14620, n14621, n14622, n14623, n14624, n14625, n14626, n14627,
         n14628, n14629, n14630, n14631, n14632, n14633, n14634, n14635,
         n14636, n14637, n14638, n14639, n14640, n14641, n14642, n14643,
         n14644, n14645, n14646, n14647, n14648, n14649, n14650, n14651,
         n14652, n14653, n14654, n14655, n14656, n14657, n14658, n14659,
         n14660, n14661, n14662, n14663, n14664, n14665, n14666, n14667,
         n14668, n14669, n14670, n14671, n14672, n14673, n14674, n14675,
         n14676, n14677, n14678, n14679, n14680, n14681, n14682, n14683,
         n14684, n14685, n14686, n14687, n14688, n14689, n14690, n14691,
         n14692, n14693, n14694, n14695, n14696, n14697, n14698, n14699,
         n14700, n14701, n14702, n14703, n14704, n14705, n14706, n14707,
         n14708, n14709, n14710, n14711, n14712, n14713, n14714, n14715,
         n14716, n14717, n14718, n14719, n14720, n14721, n14722, n14723,
         n14724, n14725, n14726, n14727, n14728, n14729, n14730, n14731,
         n14732, n14733, n14734, n14735, n14736, n14737, n14738, n14739,
         n14740, n14741, n14742, n14743, n14744, n14745, n14746, n14747,
         n14748, n14749, n14750, n14751, n14752, n14753, n14754, n14755,
         n14756, n14757, n14758, n14759, n14760, n14761, n14762, n14763,
         n14764, n14765, n14766, n14767, n14768, n14769, n14770, n14771,
         n14772, n14773, n14774, n14775, n14776, n14777, n14778, n14779,
         n14780, n14781, n14782, n14783, n14784, n14785, n14786, n14787,
         n14788, n14789, n14790, n14791, n14792, n14793, n14794, n14795,
         n14796, n14797, n14798, n14799, n14800, n14801, n14802, n14803,
         n14804, n14805, n14806, n14807, n14808, n14809, n14810, n14811,
         n14812, n14813, n14814, n14815, n14816, n14817, n14818, n14819,
         n14820, n14821, n14822, n14823, n14824, n14825, n14826, n14827,
         n14828, n14829, n14830, n14831, n14832, n14833, n14834, n14835,
         n14836, n14837, n14838, n14839, n14840, n14841, n14842, n14843,
         n14844, n14845, n14846, n14847, n14848, n14849, n14850, n14851,
         n14852, n14853, n14854, n14855, n14856, n14857, n14858, n14859,
         n14860, n14861, n14862, n14863, n14864, n14865, n14866, n14867,
         n14868, n14869, n14870, n14871, n14872, n14873, n14874, n14875,
         n14876, n14877, n14878, n14879, n14880, n14881, n14882, n14883,
         n14884, n14885, n14886, n14887, n14888, n14889, n14890, n14891,
         n14892, n14893, n14894, n14895, n14896, n14897, n14898, n14899,
         n14900, n14901, n14902, n14903, n14904, n14905, n14906, n14907,
         n14908, n14909, n14910, n14911, n14912, n14913, n14914, n14915,
         n14916, n14917, n14918, n14919, n14920, n14921, n14922, n14923,
         n14924, n14925, n14926, n14927, n14928, n14929, n14930, n14931,
         n14932, n14933, n14934, n14935, n14936, n14937, n14938, n14939,
         n14940, n14941, n14942, n14943, n14944, n14945, n14946, n14947,
         n14948, n14949, n14950, n14951, n14952, n14953, n14954, n14955,
         n14956, n14957, n14958, n14959, n14960, n14961, n14962, n14963,
         n14964, n14965, n14966, n14967, n14968, n14969, n14970, n14971,
         n14972, n14973, n14974, n14975, n14976, n14977, n14978, n14979,
         n14980, n14981, n14982, n14983, n14984, n14985, n14986, n14987,
         n14988, n14989, n14990, n14991, n14992, n14993, n14994, n14995,
         n14996, n14997, n14998, n14999, n15000, n15001, n15002, n15003,
         n15004, n15005, n15006, n15007, n15008, n15009, n15010, n15011,
         n15012, n15013, n15014, n15015, n15016, n15017, n15018, n15019,
         n15020, n15021, n15022, n15023, n15024, n15025, n15026, n15027,
         n15028, n15029, n15030, n15031, n15032, n15033, n15034, n15035,
         n15036, n15037, n15038, n15039, n15040, n15041, n15042, n15043,
         n15044, n15045, n15046, n15047, n15048, n15049, n15050, n15051,
         n15052, n15053, n15054, n15055, n15056, n15057, n15058, n15059,
         n15060, n15061, n15062, n15063, n15064, n15065, n15066, n15067,
         n15068, n15069, n15070, n15071, n15072, n15073, n15074, n15075,
         n15076, n15077, n15078, n15079, n15080, n15081, n15082, n15083,
         n15084, n15085, n15086, n15087, n15088, n15089, n15090, n15091,
         n15092, n15093, n15094, n15095, n15096, n15097, n15098, n15099,
         n15100, n15101, n15102, n15103, n15104, n15105, n15106, n15107,
         n15108, n15109, n15110, n15111, n15112, n15113, n15114, n15115,
         n15116, n15117, n15118, n15119, n15120, n15121, n15122, n15123,
         n15124, n15125, n15126, n15127, n15128, n15129, n15130, n15131,
         n15132, n15133, n15134, n15135, n15136, n15137, n15138, n15139,
         n15140, n15141, n15142, n15143, n15144, n15145, n15146, n15147,
         n15148, n15149, n15150, n15151, n15152, n15153, n15154, n15155,
         n15156, n15157, n15158, n15159, n15160, n15161, n15162, n15163,
         n15164, n15165, n15166, n15167, n15168, n15169, n15170, n15171,
         n15172, n15173, n15174, n15175, n15176, n15177, n15178, n15179,
         n15180, n15181, n15182, n15183, n15184, n15185, n15186, n15187,
         n15188, n15189, n15190, n15191, n15192, n15193, n15194, n15195,
         n15196, n15197, n15198, n15199, n15200, n15201, n15202, n15203,
         n15204, n15205, n15206, n15207, n15208, n15209, n15210, n15211,
         n15212, n15213, n15214, n15215, n15216, n15217, n15218, n15219,
         n15220, n15221, n15222, n15223, n15224, n15225, n15226, n15227,
         n15228, n15229, n15230, n15231, n15232, n15233, n15234, n15235,
         n15236, n15237, n15238, n15239, n15240, n15241, n15242, n15243,
         n15244, n15245, n15246, n15247, n15248, n15249, n15250, n15251,
         n15252, n15253, n15254, n15255, n15256, n15257, n15258, n15259,
         n15260, n15261, n15262, n15263, n15264, n15265, n15266, n15267,
         n15268, n15269, n15270, n15271, n15272, n15273, n15274, n15275,
         n15276, n15277, n15278, n15279, n15280, n15281, n15282, n15283,
         n15284, n15285, n15286, n15287, n15288, n15289, n15290, n15291,
         n15292, n15293, n15294, n15295, n15296, n15297, n15298, n15299,
         n15300, n15301, n15302, n15303, n15304, n15305, n15306, n15307,
         n15308, n15309, n15310, n15311, n15312, n15313, n15314, n15315,
         n15316, n15317, n15318, n15319, n15320, n15321, n15322, n15323,
         n15324, n15325, n15326, n15327, n15328, n15329, n15330, n15331,
         n15332, n15333, n15334, n15335, n15336, n15337, n15338, n15339,
         n15340, n15341, n15342, n15343, n15344, n15345, n15346, n15347,
         n15348, n15349, n15350, n15351, n15352, n15353, n15354, n15355,
         n15356, n15357, n15358, n15359, n15360, n15361, n15362, n15363,
         n15364, n15365, n15366, n15367, n15368, n15369, n15370, n15371,
         n15372, n15373, n15374, n15375, n15376, n15377, n15378, n15379,
         n15380, n15381, n15382, n15383, n15384, n15385, n15386, n15387,
         n15388, n15389, n15390, n15391, n15392, n15393, n15394, n15395,
         n15396, n15397, n15398, n15399, n15400, n15401, n15402, n15403,
         n15404, n15405, n15406, n15407, n15408, n15409, n15410, n15411,
         n15412, n15413, n15414, n15415, n15416, n15417, n15418, n15419,
         n15420, n15421, n15422;

  NAND2_X1 U7270 ( .A1(n8139), .A2(n8138), .ZN(n13272) );
  NAND2_X1 U7271 ( .A1(n11802), .A2(n11810), .ZN(n12531) );
  NOR2_X1 U7272 ( .A1(n11563), .A2(P3_REG3_REG_27__SCAN_IN), .ZN(n11562) );
  AND2_X1 U7273 ( .A1(n10578), .A2(n10579), .ZN(n11060) );
  INV_X1 U7274 ( .A(n12191), .ZN(n9534) );
  INV_X2 U7275 ( .A(n9445), .ZN(n9550) );
  INV_X2 U7276 ( .A(n11815), .ZN(n11811) );
  BUF_X2 U7277 ( .A(n11686), .Z(n6527) );
  CLKBUF_X2 U7278 ( .A(n10193), .Z(n11662) );
  AND4_X1 U7279 ( .A1(n9974), .A2(n9973), .A3(n9972), .A4(n9971), .ZN(n15030)
         );
  BUF_X1 U7280 ( .A(n9726), .Z(n10530) );
  INV_X1 U7281 ( .A(n12023), .ZN(n12137) );
  CLKBUF_X2 U7282 ( .A(n7607), .Z(n8156) );
  NAND4_X2 U7283 ( .A1(n8374), .A2(n8375), .A3(n8373), .A4(n8372), .ZN(n13772)
         );
  OR2_X2 U7284 ( .A1(n8092), .A2(n12230), .ZN(n11924) );
  NAND2_X1 U7285 ( .A1(n8053), .A2(P2_IR_REG_21__SCAN_IN), .ZN(n8056) );
  NAND2_X1 U7286 ( .A1(n8320), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8322) );
  INV_X4 U7287 ( .A(n14543), .ZN(n6531) );
  BUF_X1 U7288 ( .A(n11977), .Z(n6532) );
  INV_X2 U7289 ( .A(n12149), .ZN(n12157) );
  AOI21_X1 U7290 ( .B1(n7642), .B2(n7496), .A(n7663), .ZN(n7249) );
  AND2_X1 U7291 ( .A1(n13004), .A2(n12884), .ZN(n7130) );
  NAND2_X1 U7292 ( .A1(n8094), .A2(n11924), .ZN(n9444) );
  INV_X2 U7293 ( .A(n8788), .ZN(n8770) );
  INV_X2 U7294 ( .A(n10525), .ZN(n10531) );
  AND2_X1 U7295 ( .A1(n9683), .A2(n9682), .ZN(n9701) );
  XNOR2_X1 U7296 ( .A(n13050), .B(n11946), .ZN(n12191) );
  INV_X1 U7297 ( .A(n13637), .ZN(n13591) );
  OR2_X1 U7298 ( .A1(n12807), .A2(n12331), .ZN(n11613) );
  INV_X2 U7299 ( .A(n10530), .ZN(n11492) );
  INV_X1 U7300 ( .A(P3_IR_REG_31__SCAN_IN), .ZN(n9718) );
  NAND2_X1 U7301 ( .A1(n10243), .A2(n10244), .ZN(n10329) );
  INV_X1 U7302 ( .A(n8156), .ZN(n8195) );
  INV_X1 U7303 ( .A(n9550), .ZN(n12940) );
  INV_X1 U7304 ( .A(n8781), .ZN(n8776) );
  NAND2_X1 U7305 ( .A1(n8325), .A2(n8324), .ZN(n8399) );
  AND3_X1 U7306 ( .A1(n9756), .A2(n6548), .A3(n6966), .ZN(n14519) );
  OR2_X1 U7307 ( .A1(n9248), .A2(n9242), .ZN(n14572) );
  OAI21_X1 U7308 ( .B1(n7494), .B2(SI_4_), .A(n7496), .ZN(n7642) );
  OAI211_X1 U7309 ( .C1(n10530), .C2(n9999), .A(n9803), .B(n9802), .ZN(n15048)
         );
  OAI21_X1 U7310 ( .B1(n12295), .B2(n12296), .A(n6551), .ZN(n12279) );
  XNOR2_X1 U7311 ( .A(n11880), .B(n11878), .ZN(n12310) );
  XNOR2_X1 U7312 ( .A(n12372), .B(n12383), .ZN(n11125) );
  INV_X1 U7313 ( .A(n10001), .ZN(n11664) );
  AOI21_X1 U7314 ( .B1(n12588), .B2(n11792), .A(n11525), .ZN(n12573) );
  NAND2_X1 U7315 ( .A1(n6876), .A2(n6875), .ZN(n9379) );
  NAND2_X1 U7316 ( .A1(n7755), .A2(n7754), .ZN(n14811) );
  NOR2_X1 U7317 ( .A1(n11378), .A2(n11379), .ZN(n11461) );
  AOI21_X1 U7318 ( .B1(n8166), .B2(n13335), .A(n8165), .ZN(n13353) );
  NAND2_X1 U7319 ( .A1(n7842), .A2(n7841), .ZN(n12050) );
  AND2_X1 U7320 ( .A1(n8392), .A2(n8391), .ZN(n14599) );
  BUF_X1 U7321 ( .A(n8376), .Z(n9059) );
  AND2_X1 U7322 ( .A1(n14270), .A2(n9059), .ZN(n14186) );
  NAND2_X1 U7323 ( .A1(n8733), .A2(n8732), .ZN(n14162) );
  CLKBUF_X3 U7324 ( .A(n8399), .Z(n8752) );
  NAND2_X1 U7325 ( .A1(n8503), .A2(n8502), .ZN(n14635) );
  NAND2_X1 U7326 ( .A1(n8468), .A2(n8467), .ZN(n10600) );
  INV_X1 U7327 ( .A(n9854), .ZN(n14608) );
  NAND2_X1 U7328 ( .A1(n7302), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8334) );
  INV_X1 U7329 ( .A(n8153), .ZN(n11925) );
  XNOR2_X1 U7330 ( .A(n9706), .B(n9705), .ZN(n11686) );
  CLKBUF_X3 U7331 ( .A(n13412), .Z(n6523) );
  BUF_X1 U7332 ( .A(n9444), .Z(n12942) );
  NAND4_X2 U7333 ( .A1(n7629), .A2(n7628), .A3(n7627), .A4(n7626), .ZN(n13049)
         );
  NAND2_X2 U7334 ( .A1(n7700), .A2(n7699), .ZN(n7698) );
  INV_X1 U7335 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n6522) );
  NAND2_X2 U7336 ( .A1(n10469), .A2(n7731), .ZN(n10486) );
  NAND2_X2 U7337 ( .A1(n7099), .A2(n7097), .ZN(n10469) );
  NAND2_X2 U7338 ( .A1(n6956), .A2(n11600), .ZN(n12690) );
  XNOR2_X2 U7339 ( .A(n6741), .B(n12422), .ZN(n12397) );
  OR2_X2 U7340 ( .A1(n12396), .A2(n6742), .ZN(n6741) );
  NOR2_X2 U7341 ( .A1(n11533), .A2(P3_REG3_REG_24__SCAN_IN), .ZN(n11544) );
  NAND2_X2 U7342 ( .A1(n9726), .A2(n7499), .ZN(n10001) );
  NAND2_X2 U7343 ( .A1(n11720), .A2(n11717), .ZN(n10752) );
  INV_X2 U7344 ( .A(P3_ADDR_REG_19__SCAN_IN), .ZN(n8302) );
  NOR2_X4 U7345 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n8365) );
  NAND2_X2 U7346 ( .A1(n9640), .A2(n9639), .ZN(n12592) );
  NAND2_X2 U7347 ( .A1(n10552), .A2(n10551), .ZN(n11066) );
  INV_X2 U7348 ( .A(n11649), .ZN(n9387) );
  BUF_X2 U7349 ( .A(n9381), .Z(n9386) );
  NAND2_X1 U7350 ( .A1(n7889), .A2(n7888), .ZN(n13412) );
  NAND3_X4 U7351 ( .A1(n7091), .A2(n7581), .A3(n7582), .ZN(n13051) );
  OR2_X4 U7352 ( .A1(n11921), .A2(n12230), .ZN(n12180) );
  NAND2_X2 U7353 ( .A1(n7595), .A2(n7594), .ZN(n11932) );
  XNOR2_X2 U7354 ( .A(n7906), .B(P2_IR_REG_19__SCAN_IN), .ZN(n11921) );
  INV_X1 U7356 ( .A(n12023), .ZN(n6525) );
  INV_X1 U7357 ( .A(n12023), .ZN(n6526) );
  INV_X2 U7358 ( .A(n7499), .ZN(n9729) );
  INV_X4 U7359 ( .A(n7488), .ZN(n7499) );
  BUF_X4 U7360 ( .A(n12942), .Z(n6528) );
  XNOR2_X2 U7361 ( .A(n7465), .B(n7461), .ZN(n7470) );
  AOI21_X2 U7362 ( .B1(n11476), .B2(n11475), .A(n7440), .ZN(n14980) );
  OR2_X2 U7363 ( .A1(n9003), .A2(n9718), .ZN(n9004) );
  NOR3_X2 U7364 ( .A1(n12519), .A2(n12518), .A3(n15027), .ZN(n12523) );
  NAND2_X2 U7365 ( .A1(n7825), .A2(n7824), .ZN(n14356) );
  CLKBUF_X1 U7366 ( .A(n9740), .Z(n6529) );
  XNOR2_X2 U7368 ( .A(n8104), .B(n11965), .ZN(n12194) );
  INV_X1 U7369 ( .A(n13049), .ZN(n8104) );
  XNOR2_X2 U7370 ( .A(n9720), .B(n9719), .ZN(n12242) );
  AOI21_X2 U7371 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(n8289), .A(n14438), .ZN(
        n14301) );
  AOI21_X1 U7372 ( .B1(n7386), .B2(n7385), .A(n7383), .ZN(n11671) );
  XNOR2_X1 U7373 ( .A(n11619), .B(n11618), .ZN(n11624) );
  AOI21_X1 U7374 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(n8284), .A(n14434), .ZN(
        n14440) );
  INV_X1 U7375 ( .A(n12021), .ZN(n10782) );
  NAND2_X1 U7376 ( .A1(n7722), .A2(n7721), .ZN(n14795) );
  AND2_X1 U7377 ( .A1(n8423), .A2(n8422), .ZN(n14615) );
  INV_X1 U7379 ( .A(n6528), .ZN(n12915) );
  NAND2_X2 U7380 ( .A1(n10098), .A2(n12349), .ZN(n11685) );
  CLKBUF_X1 U7381 ( .A(n8094), .Z(n6538) );
  INV_X1 U7382 ( .A(n8944), .ZN(n13770) );
  AND4_X1 U7383 ( .A1(n8416), .A2(n8415), .A3(n8414), .A4(n8413), .ZN(n9866)
         );
  NAND2_X1 U7384 ( .A1(n7487), .A2(n7489), .ZN(n7237) );
  NAND2_X1 U7385 ( .A1(n9726), .A2(n9727), .ZN(n10193) );
  AND2_X1 U7386 ( .A1(n7784), .A2(n7782), .ZN(n7522) );
  NAND2_X2 U7387 ( .A1(n12242), .A2(n12463), .ZN(n9726) );
  INV_X1 U7388 ( .A(n7592), .ZN(n8037) );
  CLKBUF_X2 U7389 ( .A(n8041), .Z(n7995) );
  INV_X1 U7390 ( .A(n8199), .ZN(n7605) );
  OAI21_X1 U7391 ( .B1(n8852), .B2(P1_IR_REG_25__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n8853) );
  OAI21_X1 U7392 ( .B1(n7905), .B2(P2_IR_REG_18__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n7906) );
  NAND2_X2 U7393 ( .A1(n9727), .A2(P1_U3086), .ZN(n14266) );
  NAND2_X1 U7394 ( .A1(n9727), .A2(P3_U3151), .ZN(n11338) );
  INV_X1 U7395 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n13473) );
  NOR2_X1 U7396 ( .A1(n6976), .A2(n6793), .ZN(n6792) );
  NAND2_X1 U7397 ( .A1(n14155), .A2(n14154), .ZN(n14240) );
  AND2_X1 U7398 ( .A1(n7340), .A2(n7339), .ZN(n11822) );
  NAND2_X1 U7399 ( .A1(n13732), .A2(n13733), .ZN(n13731) );
  NAND2_X1 U7400 ( .A1(n13966), .A2(n6740), .ZN(n13965) );
  NAND2_X1 U7401 ( .A1(n13182), .A2(n13181), .ZN(n13180) );
  NAND2_X1 U7402 ( .A1(n6645), .A2(n7384), .ZN(n7383) );
  AOI21_X1 U7403 ( .B1(n11624), .B2(n15046), .A(n11623), .ZN(n11915) );
  AOI21_X1 U7404 ( .B1(n6959), .B2(n15046), .A(n6957), .ZN(n12737) );
  NAND2_X1 U7405 ( .A1(n13651), .A2(n13650), .ZN(n13716) );
  AND2_X1 U7406 ( .A1(n8804), .A2(n8832), .ZN(n8828) );
  AND2_X1 U7407 ( .A1(n7084), .A2(n6661), .ZN(n8002) );
  AND2_X1 U7408 ( .A1(n7387), .A2(n11814), .ZN(n11670) );
  NAND2_X1 U7409 ( .A1(n6878), .A2(n6882), .ZN(n12528) );
  NAND2_X1 U7410 ( .A1(n6850), .A2(n6552), .ZN(n6755) );
  AOI21_X1 U7411 ( .B1(n7290), .B2(n7289), .A(n6544), .ZN(n7288) );
  AND2_X1 U7412 ( .A1(n6722), .A2(n12540), .ZN(n6721) );
  NAND2_X1 U7413 ( .A1(n12954), .A2(n12897), .ZN(n12899) );
  OR2_X1 U7414 ( .A1(n11798), .A2(n11797), .ZN(n6722) );
  NAND2_X1 U7415 ( .A1(n8189), .A2(n8185), .ZN(n11907) );
  NAND2_X1 U7416 ( .A1(n13912), .A2(n8809), .ZN(n13936) );
  NOR2_X1 U7417 ( .A1(n14301), .A2(n14300), .ZN(n14299) );
  AND2_X1 U7418 ( .A1(n11799), .A2(n11615), .ZN(n12540) );
  NAND2_X2 U7419 ( .A1(n8758), .A2(n8757), .ZN(n14143) );
  XNOR2_X1 U7420 ( .A(n8014), .B(n8006), .ZN(n13483) );
  NOR2_X1 U7421 ( .A1(n7107), .A2(n7106), .ZN(n7105) );
  NAND2_X1 U7422 ( .A1(n6873), .A2(n6951), .ZN(n12602) );
  NAND2_X1 U7423 ( .A1(n7990), .A2(n7989), .ZN(n13375) );
  AND2_X1 U7424 ( .A1(n7102), .A2(n7917), .ZN(n7101) );
  NAND2_X1 U7425 ( .A1(n7978), .A2(n7977), .ZN(n13233) );
  OR2_X1 U7426 ( .A1(n12397), .A2(n7033), .ZN(n7031) );
  OR2_X1 U7427 ( .A1(n6607), .A2(n7104), .ZN(n7102) );
  NAND2_X1 U7428 ( .A1(n7564), .A2(n7563), .ZN(n7988) );
  NAND2_X1 U7429 ( .A1(n7242), .A2(n7240), .ZN(n7976) );
  NAND2_X2 U7430 ( .A1(n6715), .A2(n7909), .ZN(n13406) );
  OAI21_X1 U7431 ( .B1(n7557), .B2(n6694), .A(n7560), .ZN(n7241) );
  NAND2_X1 U7432 ( .A1(n8669), .A2(n8668), .ZN(n14190) );
  XNOR2_X1 U7433 ( .A(n7556), .B(SI_22_), .ZN(n7948) );
  NAND2_X1 U7434 ( .A1(n7881), .A2(n7880), .ZN(n12065) );
  NAND2_X1 U7435 ( .A1(n10242), .A2(n10241), .ZN(n10243) );
  OR2_X1 U7436 ( .A1(n7535), .A2(n7256), .ZN(n7254) );
  NAND2_X1 U7437 ( .A1(n7535), .A2(n7259), .ZN(n7258) );
  NAND2_X1 U7438 ( .A1(n8531), .A2(n8530), .ZN(n13667) );
  NAND2_X1 U7439 ( .A1(n11048), .A2(n11047), .ZN(n11102) );
  NAND2_X1 U7440 ( .A1(n8514), .A2(n8513), .ZN(n11018) );
  NAND2_X1 U7441 ( .A1(n7771), .A2(n7770), .ZN(n12021) );
  NAND2_X1 U7442 ( .A1(n8486), .A2(n8485), .ZN(n14500) );
  XNOR2_X1 U7443 ( .A(n7785), .B(n7784), .ZN(n9510) );
  XNOR2_X1 U7444 ( .A(n7808), .B(n7807), .ZN(n9514) );
  AOI21_X1 U7445 ( .B1(n7528), .B2(n7820), .A(n7234), .ZN(n7232) );
  NAND2_X1 U7446 ( .A1(n11558), .A2(n11557), .ZN(n12552) );
  NAND2_X1 U7447 ( .A1(n7735), .A2(n7272), .ZN(n7764) );
  NAND2_X1 U7448 ( .A1(n9494), .A2(n9493), .ZN(n9497) );
  AND2_X1 U7449 ( .A1(n7144), .A2(n6669), .ZN(n9598) );
  XNOR2_X1 U7450 ( .A(n7527), .B(n11261), .ZN(n7821) );
  AOI21_X2 U7451 ( .B1(n7733), .B2(n6578), .A(n7270), .ZN(n7527) );
  OR2_X1 U7452 ( .A1(n11552), .A2(P3_REG3_REG_26__SCAN_IN), .ZN(n11563) );
  NAND2_X1 U7453 ( .A1(n7716), .A2(n7715), .ZN(n9097) );
  NAND2_X1 U7454 ( .A1(n7704), .A2(n7703), .ZN(n14788) );
  NOR2_X1 U7455 ( .A1(n8266), .A2(n14283), .ZN(n8268) );
  NAND2_X1 U7456 ( .A1(n7652), .A2(n7651), .ZN(n11973) );
  AND2_X1 U7457 ( .A1(n8398), .A2(n8397), .ZN(n9854) );
  CLKBUF_X1 U7458 ( .A(n12915), .Z(n6541) );
  NAND2_X1 U7459 ( .A1(n7621), .A2(n7620), .ZN(n11946) );
  AND2_X1 U7460 ( .A1(n7023), .A2(n6658), .ZN(n14887) );
  AND3_X1 U7461 ( .A1(n10524), .A2(n10523), .A3(n10522), .ZN(n15004) );
  INV_X1 U7462 ( .A(n15030), .ZN(n12348) );
  INV_X1 U7463 ( .A(n10545), .ZN(n12344) );
  INV_X1 U7464 ( .A(n9866), .ZN(n13769) );
  NAND2_X1 U7465 ( .A1(n9792), .A2(n11672), .ZN(n15046) );
  AND4_X1 U7466 ( .A1(n10389), .A2(n10388), .A3(n10387), .A4(n10386), .ZN(
        n10545) );
  OR3_X2 U7467 ( .A1(n9395), .A2(n9394), .A3(n9393), .ZN(n15039) );
  XNOR2_X1 U7468 ( .A(n13051), .B(n11932), .ZN(n12192) );
  NAND2_X1 U7469 ( .A1(n7237), .A2(n7490), .ZN(n7630) );
  CLKBUF_X2 U7470 ( .A(n11436), .Z(n11570) );
  BUF_X2 U7471 ( .A(n6530), .Z(n6865) );
  NAND4_X1 U7472 ( .A1(n7611), .A2(n7610), .A3(n7609), .A4(n7608), .ZN(n13050)
         );
  NAND2_X2 U7473 ( .A1(n11635), .A2(n8324), .ZN(n8781) );
  NAND2_X1 U7474 ( .A1(n9704), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9706) );
  AND2_X1 U7475 ( .A1(n14830), .A2(P3_REG2_REG_3__SCAN_IN), .ZN(n14831) );
  AOI22_X1 U7476 ( .A1(n8622), .A2(P2_DATAO_REG_2__SCAN_IN), .B1(n8633), .B2(
        n13797), .ZN(n8381) );
  INV_X2 U7477 ( .A(n7596), .ZN(n8157) );
  NAND2_X1 U7478 ( .A1(n9387), .A2(n11339), .ZN(n9740) );
  AOI22_X1 U7479 ( .A1(n7908), .A2(P1_DATAO_REG_2__SCAN_IN), .B1(n7907), .B2(
        n13068), .ZN(n7621) );
  INV_X1 U7480 ( .A(n8325), .ZN(n11635) );
  INV_X2 U7481 ( .A(n8796), .ZN(n8622) );
  XNOR2_X1 U7482 ( .A(n8853), .B(P1_IR_REG_26__SCAN_IN), .ZN(n14265) );
  INV_X1 U7483 ( .A(n11637), .ZN(n8324) );
  CLKBUF_X1 U7484 ( .A(n7612), .Z(n8193) );
  INV_X1 U7485 ( .A(n8785), .ZN(n6533) );
  NAND2_X1 U7486 ( .A1(n11906), .A2(n7467), .ZN(n7607) );
  NAND2_X1 U7487 ( .A1(n7471), .A2(n7467), .ZN(n8041) );
  AND2_X1 U7488 ( .A1(n9632), .A2(n9631), .ZN(n9683) );
  NAND2_X1 U7489 ( .A1(n14257), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8319) );
  XNOR2_X1 U7490 ( .A(n8340), .B(n8339), .ZN(n10459) );
  MUX2_X1 U7491 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8059), .S(
        P2_IR_REG_20__SCAN_IN), .Z(n8062) );
  OR2_X1 U7492 ( .A1(n10580), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n11055) );
  INV_X2 U7493 ( .A(n9273), .ZN(n7907) );
  AND3_X1 U7494 ( .A1(n8356), .A2(n8355), .A3(n8354), .ZN(n8928) );
  NAND2_X1 U7495 ( .A1(n7494), .A2(SI_4_), .ZN(n7496) );
  INV_X1 U7496 ( .A(n8061), .ZN(n8060) );
  INV_X2 U7497 ( .A(n11009), .ZN(n6534) );
  XNOR2_X1 U7498 ( .A(n8346), .B(P1_IR_REG_22__SCAN_IN), .ZN(n14271) );
  NAND2_X1 U7499 ( .A1(n13474), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7463) );
  NAND2_X1 U7500 ( .A1(n6965), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8332) );
  XNOR2_X1 U7501 ( .A(n7574), .B(n7573), .ZN(n13484) );
  AND2_X1 U7502 ( .A1(n7428), .A2(n8321), .ZN(n6790) );
  INV_X2 U7503 ( .A(n11006), .ZN(n6535) );
  AND2_X1 U7504 ( .A1(n7411), .A2(n6864), .ZN(n7410) );
  AND2_X1 U7505 ( .A1(n7061), .A2(n8049), .ZN(n8057) );
  AND2_X1 U7506 ( .A1(n7439), .A2(n6592), .ZN(n6750) );
  AOI22_X1 U7507 ( .A1(n8248), .A2(n6759), .B1(P3_ADDR_REG_1__SCAN_IN), .B2(
        n6758), .ZN(n8246) );
  INV_X1 U7508 ( .A(n9014), .ZN(n6942) );
  AND2_X1 U7509 ( .A1(n6859), .A2(P3_ADDR_REG_0__SCAN_IN), .ZN(n8248) );
  AND4_X1 U7510 ( .A1(n6774), .A2(n8308), .A3(n8429), .A4(n8419), .ZN(n8311)
         );
  AND3_X1 U7511 ( .A1(n7855), .A2(n7854), .A3(n7452), .ZN(n7453) );
  AND3_X1 U7512 ( .A1(n7451), .A2(n7450), .A3(n7856), .ZN(n7454) );
  AND2_X1 U7513 ( .A1(n9374), .A2(n9373), .ZN(n9375) );
  AND3_X1 U7514 ( .A1(n6819), .A2(n6818), .A3(n7456), .ZN(n7458) );
  AND2_X1 U7515 ( .A1(n8860), .A2(n8982), .ZN(n6984) );
  AND2_X1 U7516 ( .A1(n6986), .A2(n6985), .ZN(n8862) );
  AND3_X1 U7517 ( .A1(n8864), .A2(n8863), .A3(n9150), .ZN(n6554) );
  NOR2_X1 U7518 ( .A1(P3_IR_REG_12__SCAN_IN), .A2(P3_IR_REG_10__SCAN_IN), .ZN(
        n8863) );
  INV_X1 U7519 ( .A(P3_IR_REG_6__SCAN_IN), .ZN(n8982) );
  NOR2_X2 U7520 ( .A1(P3_IR_REG_5__SCAN_IN), .A2(P3_IR_REG_7__SCAN_IN), .ZN(
        n8861) );
  INV_X4 U7521 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3088) );
  INV_X1 U7522 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n8309) );
  INV_X1 U7523 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n8337) );
  NOR2_X1 U7524 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_13__SCAN_IN), .ZN(
        n8313) );
  INV_X1 U7525 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n8336) );
  INV_X1 U7526 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n8419) );
  INV_X1 U7527 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n8429) );
  NOR2_X1 U7528 ( .A1(P1_IR_REG_7__SCAN_IN), .A2(P1_IR_REG_3__SCAN_IN), .ZN(
        n6774) );
  INV_X1 U7529 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n8051) );
  INV_X1 U7530 ( .A(P3_IR_REG_3__SCAN_IN), .ZN(n8860) );
  INV_X1 U7531 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n8050) );
  NOR2_X1 U7532 ( .A1(P3_IR_REG_1__SCAN_IN), .A2(P3_IR_REG_0__SCAN_IN), .ZN(
        n9003) );
  INV_X2 U7533 ( .A(P3_STATE_REG_SCAN_IN), .ZN(P3_U3151) );
  NOR2_X1 U7534 ( .A1(P2_IR_REG_13__SCAN_IN), .A2(P2_IR_REG_10__SCAN_IN), .ZN(
        n7856) );
  NOR2_X1 U7535 ( .A1(P2_IR_REG_12__SCAN_IN), .A2(P2_IR_REG_11__SCAN_IN), .ZN(
        n7855) );
  INV_X1 U7536 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n8847) );
  INV_X1 U7537 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n7477) );
  INV_X1 U7538 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n13852) );
  NOR2_X1 U7539 ( .A1(P2_IR_REG_6__SCAN_IN), .A2(P2_IR_REG_4__SCAN_IN), .ZN(
        n6819) );
  NOR2_X1 U7540 ( .A1(P2_IR_REG_5__SCAN_IN), .A2(P2_IR_REG_7__SCAN_IN), .ZN(
        n6818) );
  INV_X4 U7541 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  INV_X1 U7542 ( .A(P3_IR_REG_20__SCAN_IN), .ZN(n9700) );
  INV_X1 U7543 ( .A(P3_IR_REG_13__SCAN_IN), .ZN(n9150) );
  NOR2_X1 U7544 ( .A1(P3_IR_REG_11__SCAN_IN), .A2(P3_IR_REG_4__SCAN_IN), .ZN(
        n8864) );
  OR2_X4 U7545 ( .A1(n9431), .A2(n12230), .ZN(n9445) );
  AOI21_X2 U7546 ( .B1(n11873), .B2(n11872), .A(n12263), .ZN(n12305) );
  NOR2_X2 U7547 ( .A1(n12264), .A2(n12265), .ZN(n12263) );
  NOR2_X2 U7548 ( .A1(n10600), .A2(n14518), .ZN(n14504) );
  NAND2_X1 U7549 ( .A1(n14519), .A2(n14621), .ZN(n14518) );
  OAI21_X2 U7550 ( .B1(n10506), .B2(n7276), .A(n7274), .ZN(n7277) );
  OR2_X1 U7551 ( .A1(n7821), .A2(n7820), .ZN(n7235) );
  XNOR2_X1 U7552 ( .A(n7821), .B(n7820), .ZN(n9593) );
  XNOR2_X2 U7553 ( .A(n7572), .B(n7571), .ZN(n8155) );
  OR2_X1 U7554 ( .A1(n7570), .A2(n13473), .ZN(n7572) );
  OAI21_X1 U7555 ( .B1(n12179), .B2(n6562), .A(n13144), .ZN(n8094) );
  BUF_X8 U7556 ( .A(n13639), .Z(n6536) );
  AND2_X2 U7557 ( .A1(n9246), .A2(n8936), .ZN(n13639) );
  AOI21_X2 U7558 ( .B1(n9863), .B2(n6563), .A(n6627), .ZN(n9864) );
  BUF_X4 U7559 ( .A(n8037), .Z(n6537) );
  NOR2_X2 U7560 ( .A1(n11461), .A2(n11460), .ZN(n11465) );
  XNOR2_X2 U7561 ( .A(n11882), .B(n11884), .ZN(n12254) );
  NOR2_X2 U7562 ( .A1(n13890), .A2(n11391), .ZN(n14112) );
  NAND2_X1 U7563 ( .A1(n8376), .A2(n7499), .ZN(n8785) );
  XNOR2_X2 U7564 ( .A(n8052), .B(P2_IR_REG_22__SCAN_IN), .ZN(n8153) );
  OAI22_X2 U7565 ( .A1(n9661), .A2(n9660), .B1(n14580), .B2(n14556), .ZN(n9758) );
  NOR2_X2 U7566 ( .A1(n10863), .A2(n13667), .ZN(n6972) );
  OAI222_X1 U7567 ( .A1(P1_U3086), .A2(n14264), .B1(n6535), .B2(n14263), .C1(
        n15217), .C2(n14266), .ZN(P1_U3328) );
  CLKBUF_X1 U7568 ( .A(n14565), .Z(n6539) );
  OAI21_X1 U7569 ( .B1(n8951), .B2(n8785), .A(n7278), .ZN(n14565) );
  AOI21_X1 U7570 ( .B1(n6560), .B2(n8617), .A(n6923), .ZN(n6922) );
  INV_X1 U7571 ( .A(n12801), .ZN(n11890) );
  INV_X1 U7572 ( .A(n8979), .ZN(n7350) );
  INV_X1 U7573 ( .A(n8995), .ZN(n8980) );
  AND2_X1 U7574 ( .A1(n13956), .A2(n13885), .ZN(n7295) );
  NAND2_X1 U7575 ( .A1(n7009), .A2(n7008), .ZN(n7007) );
  INV_X1 U7576 ( .A(n12330), .ZN(n7008) );
  AND2_X1 U7577 ( .A1(n11880), .A2(n11879), .ZN(n11881) );
  OR2_X1 U7578 ( .A1(n12847), .A2(n12341), .ZN(n11775) );
  NOR2_X1 U7579 ( .A1(n11924), .A2(n8153), .ZN(n12179) );
  NAND2_X1 U7580 ( .A1(n10178), .A2(n12200), .ZN(n7099) );
  NAND2_X1 U7581 ( .A1(n9273), .A2(n7499), .ZN(n7612) );
  OAI21_X1 U7582 ( .B1(n6844), .B2(n11967), .A(n7303), .ZN(n11984) );
  OR2_X1 U7583 ( .A1(n6845), .A2(n11970), .ZN(n6844) );
  AND2_X1 U7584 ( .A1(n8506), .A2(n7167), .ZN(n7166) );
  INV_X1 U7585 ( .A(n8504), .ZN(n7167) );
  AND2_X1 U7586 ( .A1(n14091), .A2(n8631), .ZN(n8632) );
  OAI21_X1 U7587 ( .B1(n8659), .B2(n8658), .A(n8657), .ZN(n6920) );
  MUX2_X1 U7588 ( .A(n11782), .B(n11781), .S(n11815), .Z(n11786) );
  INV_X1 U7589 ( .A(n7272), .ZN(n7271) );
  INV_X1 U7590 ( .A(n11860), .ZN(n9708) );
  INV_X1 U7591 ( .A(n7266), .ZN(n7265) );
  OAI21_X1 U7592 ( .B1(P1_ADDR_REG_3__SCAN_IN), .B2(n8244), .A(n6586), .ZN(
        n6766) );
  INV_X1 U7593 ( .A(n7043), .ZN(n8212) );
  NAND2_X1 U7594 ( .A1(n7343), .A2(n7342), .ZN(n7341) );
  NAND2_X1 U7595 ( .A1(n11813), .A2(n11814), .ZN(n7342) );
  OR2_X1 U7596 ( .A1(n12532), .A2(n12521), .ZN(n11802) );
  NAND2_X1 U7597 ( .A1(n6888), .A2(n6620), .ZN(n6885) );
  NOR2_X1 U7598 ( .A1(n7441), .A2(n10752), .ZN(n7379) );
  NAND2_X1 U7599 ( .A1(n12532), .A2(n12521), .ZN(n11810) );
  OR2_X1 U7600 ( .A1(n12574), .A2(n6870), .ZN(n6869) );
  XNOR2_X1 U7601 ( .A(n12584), .B(n12592), .ZN(n12574) );
  OR2_X1 U7602 ( .A1(n12825), .A2(n12615), .ZN(n11787) );
  OR2_X1 U7603 ( .A1(n12866), .A2(n12719), .ZN(n11754) );
  INV_X1 U7604 ( .A(n11283), .ZN(n7140) );
  XNOR2_X1 U7605 ( .A(n12174), .B(n13022), .ZN(n12186) );
  INV_X1 U7606 ( .A(n7056), .ZN(n7055) );
  OAI21_X1 U7607 ( .B1(n6549), .B2(n7058), .A(n12188), .ZN(n7056) );
  AND2_X1 U7608 ( .A1(n13334), .A2(n7886), .ZN(n7104) );
  NAND2_X1 U7609 ( .A1(n10763), .A2(n6581), .ZN(n7076) );
  NOR2_X1 U7610 ( .A1(n12206), .A2(n7079), .ZN(n7078) );
  INV_X1 U7611 ( .A(n8120), .ZN(n7079) );
  NOR2_X1 U7612 ( .A1(n10471), .A2(n14795), .ZN(n10470) );
  NAND2_X1 U7613 ( .A1(n13714), .A2(n13569), .ZN(n7227) );
  INV_X1 U7614 ( .A(n13880), .ZN(n7301) );
  NOR2_X1 U7615 ( .A1(n14181), .A2(n14186), .ZN(n6983) );
  OAI21_X1 U7616 ( .B1(n8036), .B2(n8035), .A(n8034), .ZN(n8178) );
  NAND2_X1 U7617 ( .A1(n7976), .A2(n7974), .ZN(n7564) );
  XNOR2_X1 U7618 ( .A(n7533), .B(SI_16_), .ZN(n7851) );
  XNOR2_X1 U7619 ( .A(n6766), .B(P3_ADDR_REG_4__SCAN_IN), .ZN(n8242) );
  XNOR2_X1 U7620 ( .A(n8214), .B(P3_ADDR_REG_5__SCAN_IN), .ZN(n8240) );
  AND2_X1 U7621 ( .A1(n9689), .A2(n9688), .ZN(n9805) );
  NAND2_X1 U7622 ( .A1(n11866), .A2(n12691), .ZN(n6993) );
  NAND2_X1 U7623 ( .A1(n11883), .A2(n11884), .ZN(n7011) );
  OAI22_X1 U7624 ( .A1(n11867), .A2(n6631), .B1(n6989), .B2(n6992), .ZN(n12317) );
  AOI21_X1 U7625 ( .B1(n6542), .B2(n12296), .A(n6647), .ZN(n7009) );
  INV_X1 U7626 ( .A(n12280), .ZN(n7010) );
  INV_X1 U7627 ( .A(n6530), .ZN(n11567) );
  XNOR2_X1 U7629 ( .A(n7030), .B(n14842), .ZN(n14830) );
  OR2_X1 U7630 ( .A1(n14957), .A2(n14956), .ZN(n7022) );
  NAND2_X1 U7631 ( .A1(n6568), .A2(n6707), .ZN(n7016) );
  NAND2_X1 U7632 ( .A1(n7018), .A2(n7019), .ZN(n7017) );
  INV_X1 U7633 ( .A(n12475), .ZN(n7018) );
  AND2_X1 U7634 ( .A1(n12475), .A2(n6727), .ZN(n6568) );
  OR2_X1 U7635 ( .A1(n12455), .A2(n12465), .ZN(n6727) );
  NAND2_X1 U7636 ( .A1(n11615), .A2(n7401), .ZN(n7400) );
  INV_X1 U7637 ( .A(n7399), .ZN(n7398) );
  INV_X1 U7638 ( .A(n7402), .ZN(n7401) );
  NAND2_X1 U7639 ( .A1(n12514), .A2(n11812), .ZN(n7387) );
  NOR2_X1 U7640 ( .A1(n12650), .A2(n7389), .ZN(n7388) );
  INV_X1 U7641 ( .A(n11775), .ZN(n7389) );
  NAND2_X1 U7642 ( .A1(n14303), .A2(n11590), .ZN(n6956) );
  INV_X1 U7643 ( .A(n11662), .ZN(n11493) );
  NAND2_X1 U7644 ( .A1(n11646), .A2(n11645), .ZN(n11655) );
  INV_X1 U7645 ( .A(P3_IR_REG_27__SCAN_IN), .ZN(n7409) );
  NAND2_X1 U7646 ( .A1(n10283), .A2(n10282), .ZN(n10788) );
  NAND2_X1 U7647 ( .A1(n10281), .A2(n10280), .ZN(n10283) );
  XNOR2_X1 U7648 ( .A(n9634), .B(P3_IR_REG_19__SCAN_IN), .ZN(n12489) );
  OR2_X1 U7649 ( .A1(n9073), .A2(n9072), .ZN(n9075) );
  NAND2_X1 U7650 ( .A1(n9020), .A2(n9019), .ZN(n9037) );
  NAND2_X1 U7651 ( .A1(n7347), .A2(n7346), .ZN(n9020) );
  AND2_X1 U7652 ( .A1(n7348), .A2(n6682), .ZN(n7346) );
  NAND2_X1 U7653 ( .A1(n8976), .A2(n8975), .ZN(n8985) );
  NAND2_X1 U7654 ( .A1(n9030), .A2(n8974), .ZN(n8976) );
  NOR2_X1 U7655 ( .A1(n7138), .A2(n14339), .ZN(n7137) );
  INV_X1 U7656 ( .A(n7137), .ZN(n7135) );
  NAND2_X1 U7657 ( .A1(n8060), .A2(n8051), .ZN(n8063) );
  NOR2_X1 U7658 ( .A1(n13159), .A2(n6804), .ZN(n6803) );
  INV_X1 U7659 ( .A(n6805), .ZN(n6804) );
  XNOR2_X1 U7660 ( .A(n13351), .B(n12949), .ZN(n12224) );
  OR2_X1 U7661 ( .A1(n13216), .A2(n13205), .ZN(n13201) );
  OR2_X1 U7662 ( .A1(n13259), .A2(n13385), .ZN(n7436) );
  NAND2_X1 U7663 ( .A1(n11449), .A2(n7104), .ZN(n13322) );
  NAND2_X1 U7664 ( .A1(n7050), .A2(n8125), .ZN(n7049) );
  INV_X1 U7665 ( .A(n14349), .ZN(n7050) );
  NAND2_X1 U7666 ( .A1(n8121), .A2(n7078), .ZN(n7077) );
  NAND2_X1 U7667 ( .A1(n10464), .A2(n12201), .ZN(n7068) );
  OR2_X1 U7668 ( .A1(n9174), .A2(n7592), .ZN(n6714) );
  NOR2_X1 U7669 ( .A1(n12201), .A2(n7098), .ZN(n7097) );
  INV_X1 U7670 ( .A(n7712), .ZN(n7098) );
  NAND2_X1 U7671 ( .A1(n8008), .A2(n8007), .ZN(n13187) );
  INV_X1 U7672 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n7456) );
  INV_X1 U7673 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n7452) );
  AOI21_X1 U7674 ( .B1(n7206), .B2(n7204), .A(n6642), .ZN(n7203) );
  INV_X1 U7675 ( .A(n10607), .ZN(n7204) );
  AND4_X1 U7676 ( .A1(n8571), .A2(n8570), .A3(n8569), .A4(n8568), .ZN(n13517)
         );
  XOR2_X1 U7677 ( .A(n13758), .B(n14136), .Z(n13913) );
  NAND2_X1 U7678 ( .A1(n13962), .A2(n6788), .ZN(n13951) );
  NOR2_X1 U7679 ( .A1(n13948), .A2(n6789), .ZN(n6788) );
  INV_X1 U7680 ( .A(n13909), .ZN(n6789) );
  NAND2_X2 U7681 ( .A1(n8743), .A2(n8742), .ZN(n13956) );
  NAND2_X1 U7682 ( .A1(n13964), .A2(n13963), .ZN(n13962) );
  OR2_X1 U7683 ( .A1(n13754), .A2(n13517), .ZN(n11389) );
  NAND2_X1 U7684 ( .A1(n10317), .A2(n7297), .ZN(n14509) );
  AND2_X1 U7685 ( .A1(n10310), .A2(n10316), .ZN(n7297) );
  NAND2_X1 U7686 ( .A1(n9244), .A2(n9243), .ZN(n14497) );
  AND2_X1 U7687 ( .A1(n8936), .A2(n9187), .ZN(n9056) );
  NAND2_X1 U7688 ( .A1(n7733), .A2(n7732), .ZN(n7735) );
  NAND2_X1 U7689 ( .A1(n6846), .A2(n14420), .ZN(n8278) );
  OAI21_X1 U7690 ( .B1(n14422), .B2(n14421), .A(n7042), .ZN(n6846) );
  INV_X1 U7691 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n7042) );
  INV_X1 U7692 ( .A(n6769), .ZN(n8280) );
  OAI21_X1 U7693 ( .B1(n8233), .B2(n8232), .A(n6770), .ZN(n6769) );
  NAND2_X1 U7694 ( .A1(n14470), .A2(P3_ADDR_REG_12__SCAN_IN), .ZN(n6770) );
  OR2_X1 U7695 ( .A1(n9831), .A2(n9830), .ZN(n7113) );
  XNOR2_X1 U7696 ( .A(n12902), .B(n12901), .ZN(n12924) );
  INV_X1 U7697 ( .A(n12179), .ZN(n8093) );
  NAND2_X1 U7698 ( .A1(n6908), .A2(n6905), .ZN(n6907) );
  NAND2_X1 U7699 ( .A1(n8369), .A2(n8370), .ZN(n6908) );
  AND2_X1 U7700 ( .A1(n11945), .A2(n11944), .ZN(n11957) );
  NAND2_X1 U7701 ( .A1(n6939), .A2(n6938), .ZN(n8456) );
  NAND2_X1 U7702 ( .A1(n8441), .A2(n7163), .ZN(n6938) );
  NAND2_X1 U7703 ( .A1(n11988), .A2(n7316), .ZN(n7315) );
  NAND2_X1 U7704 ( .A1(n7319), .A2(n6613), .ZN(n7318) );
  INV_X1 U7705 ( .A(n11993), .ZN(n6821) );
  INV_X1 U7706 ( .A(n7305), .ZN(n6829) );
  INV_X1 U7707 ( .A(n12025), .ZN(n6828) );
  NAND2_X1 U7708 ( .A1(n6651), .A2(n6826), .ZN(n6825) );
  NAND2_X1 U7709 ( .A1(n6585), .A2(n7306), .ZN(n6826) );
  INV_X1 U7710 ( .A(n6831), .ZN(n6830) );
  NAND2_X1 U7711 ( .A1(n6900), .A2(n6899), .ZN(n8579) );
  NAND2_X1 U7712 ( .A1(n8532), .A2(n8534), .ZN(n6899) );
  INV_X1 U7713 ( .A(n8632), .ZN(n6927) );
  INV_X1 U7714 ( .A(n8617), .ZN(n6926) );
  INV_X1 U7715 ( .A(n12060), .ZN(n6837) );
  NAND2_X1 U7716 ( .A1(n12060), .A2(n6835), .ZN(n6834) );
  INV_X1 U7717 ( .A(n12067), .ZN(n7323) );
  INV_X1 U7718 ( .A(n12066), .ZN(n7322) );
  OAI21_X1 U7719 ( .B1(n11767), .B2(n11766), .A(n11765), .ZN(n11768) );
  INV_X1 U7720 ( .A(n12091), .ZN(n7320) );
  NAND2_X1 U7721 ( .A1(n7314), .A2(n6598), .ZN(n7311) );
  NAND2_X1 U7722 ( .A1(n6919), .A2(n6918), .ZN(n8683) );
  NAND2_X1 U7723 ( .A1(n8670), .A2(n8672), .ZN(n6918) );
  NAND2_X1 U7724 ( .A1(n11793), .A2(n12574), .ZN(n6720) );
  AND2_X1 U7725 ( .A1(n8698), .A2(n7169), .ZN(n7168) );
  INV_X1 U7726 ( .A(n8696), .ZN(n7169) );
  AOI21_X1 U7727 ( .B1(n11805), .B2(n11804), .A(n11803), .ZN(n11806) );
  INV_X1 U7728 ( .A(n12146), .ZN(n7239) );
  INV_X1 U7729 ( .A(n12147), .ZN(n7238) );
  OR2_X1 U7730 ( .A1(n14271), .A2(n8928), .ZN(n8357) );
  INV_X1 U7731 ( .A(n8723), .ZN(n6935) );
  INV_X1 U7732 ( .A(n8744), .ZN(n6917) );
  OR2_X1 U7733 ( .A1(n14405), .A2(n13506), .ZN(n8583) );
  INV_X1 U7734 ( .A(n7268), .ZN(n7267) );
  INV_X1 U7735 ( .A(n7568), .ZN(n7264) );
  AOI21_X1 U7736 ( .B1(n7987), .B2(n7568), .A(n6705), .ZN(n7266) );
  NOR2_X1 U7737 ( .A1(n6694), .A2(n7245), .ZN(n7243) );
  INV_X1 U7738 ( .A(n7949), .ZN(n7245) );
  NOR2_X1 U7739 ( .A1(n7546), .A2(n7545), .ZN(n7547) );
  OR2_X1 U7740 ( .A1(n7431), .A2(n6676), .ZN(n7270) );
  INV_X1 U7741 ( .A(n7750), .ZN(n7513) );
  INV_X1 U7742 ( .A(n7496), .ZN(n7250) );
  INV_X1 U7743 ( .A(n7498), .ZN(n7247) );
  NAND4_X1 U7744 ( .A1(n13852), .A2(n7477), .A3(n7478), .A4(
        P3_ADDR_REG_19__SCAN_IN), .ZN(n7252) );
  INV_X1 U7745 ( .A(P1_RD_REG_SCAN_IN), .ZN(n7478) );
  NAND4_X1 U7746 ( .A1(n8302), .A2(n7479), .A3(P1_ADDR_REG_19__SCAN_IN), .A4(
        P2_ADDR_REG_19__SCAN_IN), .ZN(n7251) );
  INV_X1 U7747 ( .A(P2_RD_REG_SCAN_IN), .ZN(n7479) );
  OAI21_X1 U7748 ( .B1(n8246), .B2(n8245), .A(n7044), .ZN(n7043) );
  NAND2_X1 U7749 ( .A1(n8210), .A2(P3_ADDR_REG_2__SCAN_IN), .ZN(n7044) );
  NAND2_X1 U7750 ( .A1(n14896), .A2(n10905), .ZN(n10906) );
  NAND2_X1 U7751 ( .A1(n14931), .A2(n6891), .ZN(n10908) );
  OR2_X1 U7752 ( .A1(n10947), .A2(n10945), .ZN(n6891) );
  NAND2_X1 U7753 ( .A1(n14970), .A2(n6697), .ZN(n11126) );
  NAND2_X1 U7754 ( .A1(n12364), .A2(n6889), .ZN(n12375) );
  OR2_X1 U7755 ( .A1(n12360), .A2(n11129), .ZN(n6889) );
  INV_X1 U7756 ( .A(n12419), .ZN(n7036) );
  INV_X1 U7757 ( .A(n10094), .ZN(n10095) );
  INV_X1 U7758 ( .A(n6885), .ZN(n6884) );
  AOI21_X1 U7759 ( .B1(n6883), .B2(n6885), .A(n11800), .ZN(n6882) );
  INV_X1 U7760 ( .A(n6886), .ZN(n6883) );
  OR2_X1 U7761 ( .A1(n12819), .A2(n12577), .ZN(n11791) );
  OR2_X1 U7762 ( .A1(n12764), .A2(n12626), .ZN(n11769) );
  OR2_X1 U7763 ( .A1(n11601), .A2(n12703), .ZN(n11760) );
  INV_X1 U7764 ( .A(n11479), .ZN(n7393) );
  AND3_X1 U7765 ( .A1(n8866), .A2(n6567), .A3(n9375), .ZN(n6864) );
  INV_X1 U7766 ( .A(n8869), .ZN(n7411) );
  NAND2_X1 U7767 ( .A1(n9152), .A2(P2_DATAO_REG_13__SCAN_IN), .ZN(n7361) );
  INV_X1 U7768 ( .A(n7363), .ZN(n7362) );
  OAI21_X1 U7769 ( .B1(n6579), .B2(n7364), .A(n9515), .ZN(n7363) );
  INV_X1 U7770 ( .A(n9152), .ZN(n7364) );
  OR2_X1 U7771 ( .A1(n9026), .A2(P3_IR_REG_6__SCAN_IN), .ZN(n8997) );
  NOR2_X1 U7772 ( .A1(n8956), .A2(P3_IR_REG_4__SCAN_IN), .ZN(n9034) );
  NAND2_X1 U7773 ( .A1(n6719), .A2(n10067), .ZN(n7110) );
  NAND2_X1 U7774 ( .A1(n9830), .A2(n9829), .ZN(n6719) );
  AND2_X1 U7775 ( .A1(P2_REG3_REG_24__SCAN_IN), .A2(n7981), .ZN(n7980) );
  INV_X1 U7776 ( .A(n7470), .ZN(n7467) );
  OR2_X1 U7777 ( .A1(n13356), .A2(n8032), .ZN(n8151) );
  INV_X1 U7778 ( .A(n12187), .ZN(n7052) );
  INV_X1 U7779 ( .A(n13402), .ZN(n6798) );
  NOR2_X1 U7780 ( .A1(n13327), .A2(n6523), .ZN(n13308) );
  INV_X1 U7781 ( .A(n8131), .ZN(n7070) );
  OAI21_X1 U7782 ( .B1(n9565), .B2(n7083), .A(n7081), .ZN(n10136) );
  INV_X1 U7783 ( .A(n7678), .ZN(n7083) );
  AOI21_X1 U7784 ( .B1(n7678), .B2(n7082), .A(n6628), .ZN(n7081) );
  NAND2_X1 U7785 ( .A1(n8057), .A2(n8050), .ZN(n8061) );
  INV_X1 U7786 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n7066) );
  INV_X1 U7787 ( .A(n13700), .ZN(n7230) );
  INV_X1 U7788 ( .A(n11022), .ZN(n7202) );
  OR2_X1 U7789 ( .A1(n8746), .A2(n6917), .ZN(n6916) );
  NOR2_X1 U7790 ( .A1(n8762), .A2(n8759), .ZN(n7154) );
  NAND2_X1 U7791 ( .A1(n8759), .A2(n8762), .ZN(n7153) );
  NAND2_X1 U7792 ( .A1(n7413), .A2(n13899), .ZN(n7412) );
  INV_X1 U7793 ( .A(n7414), .ZN(n7413) );
  AND2_X1 U7794 ( .A1(n7415), .A2(n13898), .ZN(n7414) );
  INV_X1 U7795 ( .A(n14049), .ZN(n7415) );
  NOR2_X1 U7796 ( .A1(n14096), .A2(n14109), .ZN(n7423) );
  NOR2_X1 U7797 ( .A1(n7423), .A2(n7420), .ZN(n7419) );
  INV_X1 U7798 ( .A(n7422), .ZN(n7420) );
  AND2_X1 U7799 ( .A1(n8583), .A2(n11295), .ZN(n11212) );
  NAND2_X1 U7800 ( .A1(n9753), .A2(n14545), .ZN(n9762) );
  INV_X1 U7801 ( .A(n13771), .ZN(n9753) );
  AND2_X1 U7802 ( .A1(n10459), .A2(n9242), .ZN(n9246) );
  XNOR2_X1 U7803 ( .A(n14556), .B(n14580), .ZN(n6776) );
  NAND2_X1 U7804 ( .A1(n7262), .A2(n7266), .ZN(n7269) );
  NAND2_X1 U7805 ( .A1(n7988), .A2(n7568), .ZN(n7262) );
  NAND2_X1 U7806 ( .A1(n8003), .A2(n11550), .ZN(n7268) );
  NAND2_X1 U7807 ( .A1(n7554), .A2(n7553), .ZN(n7556) );
  INV_X1 U7808 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n8312) );
  NOR2_X1 U7809 ( .A1(P1_IR_REG_14__SCAN_IN), .A2(P1_IR_REG_12__SCAN_IN), .ZN(
        n8315) );
  NOR2_X1 U7810 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(P1_IR_REG_11__SCAN_IN), .ZN(
        n8314) );
  NAND2_X1 U7811 ( .A1(n8561), .A2(n7173), .ZN(n8605) );
  AND2_X1 U7812 ( .A1(n8336), .A2(n8337), .ZN(n7173) );
  XNOR2_X1 U7813 ( .A(n7529), .B(SI_15_), .ZN(n7837) );
  NAND2_X1 U7814 ( .A1(n7509), .A2(SI_9_), .ZN(n7511) );
  NAND2_X1 U7815 ( .A1(n7506), .A2(SI_8_), .ZN(n7508) );
  INV_X1 U7816 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n8308) );
  NAND2_X1 U7817 ( .A1(n7630), .A2(n7492), .ZN(n7633) );
  INV_X1 U7818 ( .A(n7237), .ZN(n7236) );
  AND2_X2 U7819 ( .A1(n7252), .A2(n7251), .ZN(n7488) );
  INV_X1 U7820 ( .A(n7045), .ZN(n8214) );
  OAI21_X1 U7821 ( .B1(n8242), .B2(P1_ADDR_REG_4__SCAN_IN), .A(n6765), .ZN(
        n7045) );
  INV_X1 U7822 ( .A(n6763), .ZN(n8217) );
  OAI21_X1 U7823 ( .B1(n8262), .B2(n8263), .A(n6688), .ZN(n6763) );
  AND2_X1 U7824 ( .A1(n6768), .A2(n6767), .ZN(n8239) );
  NAND2_X1 U7825 ( .A1(n9131), .A2(P3_ADDR_REG_8__SCAN_IN), .ZN(n6767) );
  OR2_X1 U7826 ( .A1(n8272), .A2(n8271), .ZN(n6768) );
  AOI21_X1 U7827 ( .B1(P3_ADDR_REG_9__SCAN_IN), .B2(n8221), .A(n8220), .ZN(
        n8222) );
  NOR2_X1 U7828 ( .A1(n8239), .A2(n8238), .ZN(n8220) );
  AND2_X1 U7829 ( .A1(n6772), .A2(n6771), .ZN(n8233) );
  NAND2_X1 U7830 ( .A1(n8225), .A2(P3_ADDR_REG_11__SCAN_IN), .ZN(n6771) );
  OR2_X1 U7831 ( .A1(n8235), .A2(n8234), .ZN(n6772) );
  OR2_X1 U7832 ( .A1(n6865), .A2(n11086), .ZN(n11092) );
  INV_X1 U7833 ( .A(n14985), .ZN(n11472) );
  NAND2_X1 U7834 ( .A1(n6723), .A2(n10061), .ZN(n10094) );
  NOR2_X2 U7835 ( .A1(n15386), .A2(n15387), .ZN(n15385) );
  AOI21_X1 U7836 ( .B1(n12288), .B2(n6990), .A(n6614), .ZN(n6989) );
  INV_X1 U7837 ( .A(n6993), .ZN(n6990) );
  AOI21_X1 U7838 ( .B1(n6999), .B2(n11265), .A(n6637), .ZN(n6998) );
  INV_X1 U7839 ( .A(n11169), .ZN(n6999) );
  INV_X1 U7840 ( .A(n11265), .ZN(n7000) );
  NAND2_X1 U7841 ( .A1(n11670), .A2(n11809), .ZN(n7386) );
  NAND2_X1 U7842 ( .A1(n11686), .A2(n9791), .ZN(n11852) );
  NOR2_X1 U7843 ( .A1(n11817), .A2(n11818), .ZN(n7339) );
  OAI211_X1 U7844 ( .C1(n7343), .C2(n11811), .A(n7341), .B(n11809), .ZN(n7340)
         );
  OR2_X1 U7845 ( .A1(n6865), .A2(n11122), .ZN(n11077) );
  NAND2_X1 U7846 ( .A1(n7371), .A2(P3_REG0_REG_0__SCAN_IN), .ZN(n9715) );
  NAND2_X1 U7847 ( .A1(n10889), .A2(n10888), .ZN(n7030) );
  NAND2_X1 U7848 ( .A1(n14898), .A2(n14897), .ZN(n14896) );
  AND2_X1 U7849 ( .A1(n14857), .A2(P3_REG2_REG_4__SCAN_IN), .ZN(n7025) );
  XNOR2_X1 U7850 ( .A(n10906), .B(n10941), .ZN(n14915) );
  OR2_X1 U7851 ( .A1(n14922), .A2(n14921), .ZN(n7028) );
  NAND2_X1 U7852 ( .A1(n14933), .A2(n14932), .ZN(n14931) );
  XNOR2_X1 U7853 ( .A(n10908), .B(n10954), .ZN(n14950) );
  NAND2_X1 U7854 ( .A1(n7028), .A2(n7027), .ZN(n7026) );
  NAND2_X1 U7855 ( .A1(n14928), .A2(P3_REG2_REG_8__SCAN_IN), .ZN(n7027) );
  NAND2_X1 U7856 ( .A1(n14972), .A2(n14971), .ZN(n14970) );
  XNOR2_X1 U7857 ( .A(n11126), .B(n6890), .ZN(n10910) );
  NAND2_X1 U7858 ( .A1(n12366), .A2(n12365), .ZN(n12364) );
  INV_X1 U7859 ( .A(n7020), .ZN(n11119) );
  NAND2_X1 U7860 ( .A1(n6576), .A2(n6724), .ZN(n12362) );
  XNOR2_X1 U7861 ( .A(n12375), .B(n12383), .ZN(n11130) );
  NOR2_X1 U7862 ( .A1(n12432), .A2(n12416), .ZN(n12418) );
  INV_X1 U7863 ( .A(n6741), .ZN(n12416) );
  OR2_X1 U7864 ( .A1(n12397), .A2(n12693), .ZN(n7035) );
  NAND2_X1 U7865 ( .A1(n12423), .A2(n12424), .ZN(n12425) );
  NAND2_X1 U7866 ( .A1(n12425), .A2(n12426), .ZN(n12443) );
  OR2_X1 U7867 ( .A1(n6961), .A2(n12531), .ZN(n6960) );
  NAND2_X1 U7868 ( .A1(n6881), .A2(n6885), .ZN(n6961) );
  NOR2_X1 U7869 ( .A1(n6872), .A2(n6869), .ZN(n6867) );
  NAND2_X1 U7870 ( .A1(n11433), .A2(n15204), .ZN(n11435) );
  AOI21_X1 U7871 ( .B1(n11479), .B2(n14982), .A(n7396), .ZN(n7395) );
  INV_X1 U7872 ( .A(n11737), .ZN(n7396) );
  AND2_X1 U7873 ( .A1(n11076), .A2(n11075), .ZN(n14309) );
  INV_X1 U7874 ( .A(n15388), .ZN(n14320) );
  OR2_X1 U7875 ( .A1(n14980), .A2(n14982), .ZN(n14313) );
  NAND2_X1 U7876 ( .A1(n7374), .A2(n7372), .ZN(n11476) );
  INV_X1 U7877 ( .A(n7373), .ZN(n7372) );
  OAI21_X1 U7878 ( .B1(n7379), .B2(n7376), .A(n11834), .ZN(n7373) );
  NAND2_X1 U7879 ( .A1(n10748), .A2(n10747), .ZN(n7380) );
  AND4_X1 U7880 ( .A1(n10272), .A2(n10271), .A3(n10270), .A4(n10269), .ZN(
        n10708) );
  OR2_X1 U7881 ( .A1(n6530), .A2(n10933), .ZN(n10269) );
  AND4_X1 U7882 ( .A1(n10017), .A2(n10016), .A3(n10015), .A4(n10014), .ZN(
        n10709) );
  AND2_X1 U7883 ( .A1(n11709), .A2(n11708), .ZN(n11826) );
  AND2_X1 U7884 ( .A1(n9788), .A2(n9699), .ZN(n10088) );
  NOR2_X1 U7885 ( .A1(n6988), .A2(n9686), .ZN(n9789) );
  NOR2_X1 U7886 ( .A1(n12529), .A2(n11575), .ZN(n12514) );
  NAND2_X1 U7887 ( .A1(n11680), .A2(n11675), .ZN(n7402) );
  OR2_X1 U7888 ( .A1(n6954), .A2(n6596), .ZN(n6951) );
  NAND2_X1 U7889 ( .A1(n12623), .A2(n6952), .ZN(n6873) );
  NOR2_X1 U7890 ( .A1(n6596), .A2(n6953), .ZN(n6952) );
  INV_X1 U7891 ( .A(n7407), .ZN(n7406) );
  AOI21_X1 U7892 ( .B1(n11509), .B2(n11496), .A(n7408), .ZN(n7407) );
  INV_X1 U7893 ( .A(n11784), .ZN(n7408) );
  XNOR2_X1 U7894 ( .A(n12758), .B(n12627), .ZN(n12614) );
  NAND2_X1 U7895 ( .A1(n12652), .A2(n11769), .ZN(n12634) );
  NAND2_X1 U7896 ( .A1(n11588), .A2(n11587), .ZN(n14303) );
  AND2_X1 U7897 ( .A1(n11811), .A2(n9820), .ZN(n15041) );
  OR2_X1 U7898 ( .A1(n9788), .A2(n9787), .ZN(n10398) );
  AND3_X1 U7899 ( .A1(n11811), .A2(n10396), .A3(n9799), .ZN(n10399) );
  INV_X1 U7900 ( .A(n10089), .ZN(n10396) );
  OR2_X1 U7901 ( .A1(n11815), .A2(n9820), .ZN(n15031) );
  INV_X1 U7902 ( .A(n15046), .ZN(n15027) );
  AND4_X2 U7903 ( .A1(n9744), .A2(n9743), .A3(n9742), .A4(n9741), .ZN(n15028)
         );
  OR2_X1 U7904 ( .A1(n9738), .A2(n9737), .ZN(n9743) );
  AOI21_X1 U7905 ( .B1(P3_IR_REG_31__SCAN_IN), .B2(P3_IR_REG_28__SCAN_IN), .A(
        P3_IR_REG_29__SCAN_IN), .ZN(n6877) );
  NAND2_X1 U7906 ( .A1(n11337), .A2(n11336), .ZN(n11643) );
  NAND2_X1 U7907 ( .A1(n11578), .A2(n11335), .ZN(n11337) );
  NAND2_X1 U7908 ( .A1(n11334), .A2(n11333), .ZN(n11578) );
  NAND2_X1 U7909 ( .A1(n11117), .A2(n11116), .ZN(n11334) );
  NAND2_X1 U7910 ( .A1(n11003), .A2(n11002), .ZN(n11114) );
  NAND2_X1 U7911 ( .A1(n10790), .A2(n10789), .ZN(n10791) );
  OR2_X1 U7912 ( .A1(n10788), .A2(n10787), .ZN(n10790) );
  NAND2_X1 U7913 ( .A1(n7332), .A2(n7330), .ZN(n10281) );
  AOI21_X1 U7914 ( .B1(n7333), .B2(n7335), .A(n7331), .ZN(n7330) );
  INV_X1 U7915 ( .A(n10118), .ZN(n7331) );
  NAND2_X1 U7916 ( .A1(n9680), .A2(n9679), .ZN(n10028) );
  NAND2_X1 U7917 ( .A1(n9629), .A2(n9628), .ZN(n9677) );
  NAND2_X1 U7918 ( .A1(n7326), .A2(n7324), .ZN(n9624) );
  AOI21_X1 U7919 ( .B1(n7327), .B2(n7329), .A(n7325), .ZN(n7324) );
  NAND2_X1 U7920 ( .A1(n9497), .A2(n7327), .ZN(n7326) );
  INV_X1 U7921 ( .A(n9617), .ZN(n7325) );
  NAND2_X1 U7922 ( .A1(n9497), .A2(n9496), .ZN(n9528) );
  AND2_X1 U7923 ( .A1(n8865), .A2(n6946), .ZN(n6945) );
  NOR2_X1 U7924 ( .A1(n6941), .A2(n9014), .ZN(n6947) );
  NAND2_X1 U7925 ( .A1(n9049), .A2(n9048), .ZN(n9073) );
  NAND2_X1 U7926 ( .A1(n7338), .A2(n7336), .ZN(n9049) );
  AOI21_X1 U7927 ( .B1(n8978), .B2(n7349), .A(n6572), .ZN(n7348) );
  NAND2_X1 U7928 ( .A1(n8985), .A2(n7349), .ZN(n7347) );
  XNOR2_X1 U7929 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .ZN(n8995) );
  NAND2_X1 U7930 ( .A1(n9068), .A2(P2_DATAO_REG_6__SCAN_IN), .ZN(n8979) );
  XNOR2_X1 U7931 ( .A(n9066), .B(P1_DATAO_REG_5__SCAN_IN), .ZN(n9029) );
  OAI21_X1 U7932 ( .B1(n9013), .B2(n7355), .A(n7354), .ZN(n9030) );
  NAND2_X1 U7933 ( .A1(n8972), .A2(n7357), .ZN(n7355) );
  AOI21_X1 U7934 ( .B1(n6553), .B2(n8972), .A(n6590), .ZN(n7354) );
  NAND2_X1 U7935 ( .A1(n9016), .A2(n8956), .ZN(n10917) );
  NAND2_X1 U7936 ( .A1(n8954), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n9041) );
  INV_X1 U7937 ( .A(n12965), .ZN(n7146) );
  NAND2_X1 U7938 ( .A1(n12890), .A2(n12891), .ZN(n6746) );
  OAI21_X1 U7939 ( .B1(n7140), .B2(n7135), .A(n7142), .ZN(n7134) );
  INV_X1 U7940 ( .A(n11377), .ZN(n7142) );
  NAND2_X1 U7941 ( .A1(n7127), .A2(n7131), .ZN(n7129) );
  NAND2_X1 U7942 ( .A1(n9458), .A2(n9449), .ZN(n9450) );
  NAND2_X1 U7943 ( .A1(n7980), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n7994) );
  NOR2_X1 U7944 ( .A1(n13013), .A2(n12910), .ZN(n7148) );
  OR3_X1 U7945 ( .A1(n12225), .A2(n12224), .A3(n12223), .ZN(n12229) );
  NAND2_X1 U7946 ( .A1(n11906), .A2(n7470), .ZN(n7625) );
  NAND2_X1 U7947 ( .A1(n13180), .A2(n6736), .ZN(n13169) );
  AND2_X1 U7948 ( .A1(n13170), .A2(n13171), .ZN(n6736) );
  AOI21_X1 U7949 ( .B1(n13224), .B2(n7086), .A(n6630), .ZN(n7085) );
  INV_X1 U7950 ( .A(n7059), .ZN(n7058) );
  AOI21_X1 U7951 ( .B1(n8149), .B2(n6594), .A(n8148), .ZN(n7059) );
  INV_X1 U7952 ( .A(n13223), .ZN(n7088) );
  NAND2_X1 U7953 ( .A1(n13256), .A2(n8143), .ZN(n13240) );
  NAND2_X1 U7954 ( .A1(n13272), .A2(n7080), .ZN(n13256) );
  AND2_X1 U7955 ( .A1(n13250), .A2(n8141), .ZN(n7080) );
  NAND2_X1 U7956 ( .A1(n13272), .A2(n8141), .ZN(n13254) );
  NAND2_X1 U7957 ( .A1(n6738), .A2(n6737), .ZN(n13286) );
  INV_X1 U7958 ( .A(n13289), .ZN(n6737) );
  NAND2_X1 U7959 ( .A1(n8123), .A2(n10984), .ZN(n14349) );
  INV_X1 U7960 ( .A(n7076), .ZN(n7075) );
  NAND2_X1 U7961 ( .A1(n7077), .A2(n6581), .ZN(n10765) );
  AND2_X1 U7962 ( .A1(n12202), .A2(n8116), .ZN(n7067) );
  INV_X1 U7963 ( .A(n12202), .ZN(n10485) );
  NAND2_X1 U7964 ( .A1(n10485), .A2(n10486), .ZN(n10484) );
  INV_X1 U7965 ( .A(n12198), .ZN(n10138) );
  NAND2_X1 U7966 ( .A1(n9569), .A2(n9566), .ZN(n9565) );
  NOR2_X1 U7967 ( .A1(n9532), .A2(n11965), .ZN(n9567) );
  INV_X1 U7968 ( .A(n13335), .ZN(n14351) );
  NAND2_X1 U7969 ( .A1(n8039), .A2(n8038), .ZN(n13351) );
  INV_X1 U7970 ( .A(n14806), .ZN(n14810) );
  AND2_X1 U7971 ( .A1(n7459), .A2(n6665), .ZN(n7108) );
  INV_X1 U7972 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n7571) );
  AND2_X1 U7973 ( .A1(n6599), .A2(n10287), .ZN(n7209) );
  INV_X1 U7974 ( .A(n7183), .ZN(n7182) );
  OAI21_X1 U7975 ( .B1(n11238), .B2(n7184), .A(n13498), .ZN(n7183) );
  INV_X1 U7976 ( .A(n11244), .ZN(n7184) );
  AND2_X1 U7977 ( .A1(n13701), .A2(n13578), .ZN(n13619) );
  INV_X1 U7978 ( .A(n10673), .ZN(n7207) );
  NOR2_X1 U7979 ( .A1(n13537), .A2(n13526), .ZN(n7199) );
  AOI21_X1 U7980 ( .B1(n13709), .B2(n13708), .A(n13553), .ZN(n13651) );
  AOI21_X1 U7981 ( .B1(n13746), .B2(n13745), .A(n7170), .ZN(n13680) );
  NAND2_X1 U7982 ( .A1(n13680), .A2(n13681), .ZN(n13692) );
  NAND2_X1 U7983 ( .A1(n7222), .A2(n7230), .ZN(n7221) );
  INV_X1 U7984 ( .A(n7225), .ZN(n7222) );
  AOI21_X1 U7985 ( .B1(n6546), .B2(n7229), .A(n7226), .ZN(n7225) );
  INV_X1 U7986 ( .A(n13701), .ZN(n7226) );
  AOI21_X1 U7987 ( .B1(n7177), .B2(n8903), .A(n7176), .ZN(n9924) );
  NOR2_X1 U7988 ( .A1(n7178), .A2(n9838), .ZN(n7176) );
  NOR2_X1 U7989 ( .A1(n8934), .A2(n7179), .ZN(n7177) );
  NAND2_X1 U7990 ( .A1(n8902), .A2(n9841), .ZN(n7179) );
  NAND2_X1 U7991 ( .A1(n8636), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n8648) );
  NOR2_X1 U7992 ( .A1(n13724), .A2(n7196), .ZN(n7195) );
  INV_X1 U7993 ( .A(n7198), .ZN(n7196) );
  NOR2_X1 U7994 ( .A1(n9936), .A2(n9937), .ZN(n7212) );
  NAND2_X1 U7995 ( .A1(n6589), .A2(n7178), .ZN(n9925) );
  OAI22_X1 U7996 ( .A1(n8735), .A2(n7156), .B1(n8736), .B2(n7155), .ZN(n8745)
         );
  INV_X1 U7997 ( .A(n8734), .ZN(n7155) );
  NOR2_X1 U7998 ( .A1(n8737), .A2(n8734), .ZN(n7156) );
  INV_X1 U7999 ( .A(n8763), .ZN(n8784) );
  AND2_X1 U8000 ( .A1(n9052), .A2(n8924), .ZN(n8854) );
  AOI21_X1 U8001 ( .B1(n9477), .B2(P1_REG1_REG_10__SCAN_IN), .A(n9476), .ZN(
        n9488) );
  AOI21_X1 U8002 ( .B1(n11194), .B2(P1_REG1_REG_16__SCAN_IN), .A(n11193), .ZN(
        n13824) );
  AND2_X1 U8003 ( .A1(n7290), .A2(n6740), .ZN(n7287) );
  XNOR2_X1 U8004 ( .A(n14168), .B(n13907), .ZN(n13989) );
  NAND2_X1 U8005 ( .A1(n13994), .A2(n13998), .ZN(n7424) );
  NOR2_X1 U8006 ( .A1(n14034), .A2(n7281), .ZN(n7280) );
  NAND2_X1 U8007 ( .A1(n14010), .A2(n14020), .ZN(n14009) );
  NAND2_X1 U8008 ( .A1(n14065), .A2(n7414), .ZN(n14046) );
  NOR2_X1 U8009 ( .A1(n13897), .A2(n13871), .ZN(n6779) );
  NAND2_X1 U8010 ( .A1(n6781), .A2(n14068), .ZN(n6780) );
  INV_X1 U8011 ( .A(n14071), .ZN(n6781) );
  AND2_X1 U8012 ( .A1(n6588), .A2(n13891), .ZN(n7422) );
  NOR2_X1 U8013 ( .A1(n13865), .A2(n7285), .ZN(n7284) );
  INV_X1 U8014 ( .A(n11389), .ZN(n7285) );
  NAND2_X1 U8015 ( .A1(n8603), .A2(n8602), .ZN(n13890) );
  OAI21_X1 U8016 ( .B1(n11147), .B2(n6787), .A(n6641), .ZN(n11397) );
  AND2_X1 U8017 ( .A1(n11387), .A2(n11301), .ZN(n7427) );
  NAND2_X1 U8018 ( .A1(n6786), .A2(n11152), .ZN(n6785) );
  NAND2_X1 U8019 ( .A1(n11211), .A2(n6786), .ZN(n11302) );
  NAND2_X1 U8020 ( .A1(n11147), .A2(n11151), .ZN(n11211) );
  NAND2_X1 U8021 ( .A1(n10813), .A2(n6783), .ZN(n6782) );
  NOR2_X1 U8022 ( .A1(n10869), .A2(n6784), .ZN(n6783) );
  INV_X1 U8023 ( .A(n10812), .ZN(n6784) );
  NAND2_X1 U8024 ( .A1(n9397), .A2(n8417), .ZN(n8514) );
  NAND2_X1 U8025 ( .A1(n10506), .A2(n10504), .ZN(n10807) );
  AND2_X1 U8026 ( .A1(n8931), .A2(n9128), .ZN(n14107) );
  INV_X1 U8027 ( .A(n10504), .ZN(n10810) );
  OR2_X1 U8028 ( .A1(n14572), .A2(n13847), .ZN(n9251) );
  NAND2_X1 U8029 ( .A1(n9864), .A2(n10305), .ZN(n10317) );
  NAND2_X1 U8030 ( .A1(n8695), .A2(n8694), .ZN(n14181) );
  NAND2_X1 U8031 ( .A1(n8608), .A2(n8607), .ZN(n14218) );
  NAND2_X1 U8032 ( .A1(n9664), .A2(n8930), .ZN(n14607) );
  INV_X1 U8033 ( .A(n14497), .ZN(n14560) );
  OR2_X1 U8034 ( .A1(n8184), .A2(n8183), .ZN(n8189) );
  AND2_X1 U8035 ( .A1(n6675), .A2(n8331), .ZN(n7428) );
  OR2_X1 U8036 ( .A1(n8849), .A2(P1_IR_REG_24__SCAN_IN), .ZN(n8852) );
  XNOR2_X1 U8037 ( .A(n8004), .B(n7569), .ZN(n13486) );
  OAI21_X1 U8038 ( .B1(n7988), .B2(n7987), .A(n7568), .ZN(n8004) );
  OR2_X1 U8039 ( .A1(n8605), .A2(P1_IR_REG_17__SCAN_IN), .ZN(n8620) );
  INV_X1 U8040 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n8353) );
  XNOR2_X1 U8041 ( .A(n7923), .B(n7922), .ZN(n10458) );
  NAND2_X1 U8042 ( .A1(n7258), .A2(n7257), .ZN(n7920) );
  NAND2_X1 U8043 ( .A1(n8311), .A2(n8310), .ZN(n8444) );
  NAND2_X1 U8044 ( .A1(n15407), .A2(n8258), .ZN(n8260) );
  XOR2_X1 U8045 ( .A(P3_ADDR_REG_7__SCAN_IN), .B(n8217), .Z(n8267) );
  AND2_X1 U8046 ( .A1(n7039), .A2(n14286), .ZN(n8274) );
  OAI21_X1 U8047 ( .B1(n14288), .B2(n14287), .A(n7040), .ZN(n7039) );
  AOI21_X1 U8048 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(n12408), .A(n8287), .ZN(
        n8291) );
  OAI211_X1 U8049 ( .C1(n7007), .C2(n7011), .A(n7001), .B(n7004), .ZN(n12246)
         );
  AOI21_X1 U8050 ( .B1(n7009), .B2(n7006), .A(n7005), .ZN(n7004) );
  NOR2_X1 U8051 ( .A1(n11891), .A2(n12552), .ZN(n7005) );
  AND3_X1 U8052 ( .A1(n10568), .A2(n10567), .A3(n10566), .ZN(n14988) );
  NAND2_X1 U8053 ( .A1(n11532), .A2(n11531), .ZN(n12745) );
  OR2_X1 U8054 ( .A1(n11662), .A2(n11530), .ZN(n11531) );
  AND3_X1 U8055 ( .A1(n10197), .A2(n10196), .A3(n10195), .ZN(n10633) );
  INV_X1 U8056 ( .A(n11879), .ZN(n11878) );
  INV_X1 U8057 ( .A(n15401), .ZN(n12318) );
  INV_X1 U8058 ( .A(n10709), .ZN(n12347) );
  OAI21_X1 U8059 ( .B1(n12496), .B2(n12495), .A(n6712), .ZN(n6898) );
  NAND2_X1 U8060 ( .A1(n7016), .A2(n6622), .ZN(n7015) );
  NOR2_X1 U8061 ( .A1(n12491), .A2(n12483), .ZN(n7013) );
  NAND2_X1 U8062 ( .A1(n6568), .A2(n6710), .ZN(n7014) );
  NAND2_X1 U8063 ( .A1(n6895), .A2(n6894), .ZN(n6893) );
  INV_X1 U8064 ( .A(n12502), .ZN(n6894) );
  NAND2_X1 U8065 ( .A1(n12503), .A2(n14961), .ZN(n6895) );
  AND2_X1 U8066 ( .A1(n11562), .A2(n11898), .ZN(n12506) );
  NAND2_X1 U8067 ( .A1(n11513), .A2(n11512), .ZN(n12825) );
  OR2_X1 U8068 ( .A1(n11662), .A2(n11511), .ZN(n11512) );
  NAND2_X1 U8069 ( .A1(n11487), .A2(n11486), .ZN(n12847) );
  OR2_X1 U8070 ( .A1(n15086), .A2(n12748), .ZN(n12859) );
  NAND2_X1 U8071 ( .A1(n11263), .A2(n11262), .ZN(n12866) );
  XNOR2_X1 U8072 ( .A(n9703), .B(n9702), .ZN(n11860) );
  OAI21_X1 U8073 ( .B1(n9704), .B2(P3_IR_REG_21__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n9703) );
  OR2_X1 U8074 ( .A1(n9086), .A2(n7592), .ZN(n7704) );
  NAND2_X1 U8075 ( .A1(n7964), .A2(n7963), .ZN(n13385) );
  OR2_X1 U8076 ( .A1(n9097), .A2(n7592), .ZN(n7722) );
  INV_X1 U8077 ( .A(n7117), .ZN(n7116) );
  OAI22_X1 U8078 ( .A1(n7120), .A2(n10620), .B1(n10842), .B2(n10843), .ZN(
        n7117) );
  NAND2_X1 U8079 ( .A1(n12974), .A2(n12907), .ZN(n12966) );
  NAND2_X1 U8080 ( .A1(n12966), .A2(n12965), .ZN(n12964) );
  NAND2_X1 U8081 ( .A1(n9605), .A2(n9604), .ZN(n9831) );
  NAND2_X1 U8082 ( .A1(n8063), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8052) );
  NAND2_X1 U8083 ( .A1(n6800), .A2(n6806), .ZN(n6799) );
  AND2_X1 U8084 ( .A1(n11449), .A2(n7886), .ZN(n13320) );
  NAND2_X1 U8085 ( .A1(n7071), .A2(n8131), .ZN(n13333) );
  NAND2_X1 U8086 ( .A1(n8075), .A2(n14773), .ZN(n13323) );
  INV_X1 U8087 ( .A(n9415), .ZN(n8075) );
  AND3_X1 U8088 ( .A1(n11011), .A2(P2_STATE_REG_SCAN_IN), .A3(n9553), .ZN(
        n14773) );
  NAND2_X1 U8089 ( .A1(n7304), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7574) );
  AND2_X1 U8090 ( .A1(n7454), .A2(n7458), .ZN(n7064) );
  NAND2_X1 U8091 ( .A1(n13610), .A2(n13611), .ZN(n13635) );
  NAND2_X1 U8092 ( .A1(n11638), .A2(n8417), .ZN(n8758) );
  INV_X1 U8093 ( .A(n14061), .ZN(n14197) );
  INV_X1 U8094 ( .A(n13756), .ZN(n14395) );
  NAND2_X1 U8095 ( .A1(n8943), .A2(n14542), .ZN(n14398) );
  NAND2_X1 U8096 ( .A1(n8769), .A2(n8768), .ZN(n14136) );
  NAND2_X1 U8097 ( .A1(n13951), .A2(n13911), .ZN(n13937) );
  NAND2_X1 U8098 ( .A1(n13951), .A2(n7425), .ZN(n13938) );
  NOR2_X1 U8099 ( .A1(n13936), .A2(n7426), .ZN(n7425) );
  INV_X1 U8100 ( .A(n13911), .ZN(n7426) );
  XNOR2_X1 U8101 ( .A(n13928), .B(n6752), .ZN(n6751) );
  INV_X1 U8102 ( .A(n13936), .ZN(n6752) );
  NAND2_X1 U8103 ( .A1(n7291), .A2(n7292), .ZN(n13928) );
  OR2_X1 U8104 ( .A1(n9174), .A2(n8785), .ZN(n8486) );
  NAND2_X1 U8105 ( .A1(n14135), .A2(n14641), .ZN(n6794) );
  INV_X1 U8106 ( .A(n14139), .ZN(n6793) );
  NAND2_X1 U8107 ( .A1(n6863), .A2(n6862), .ZN(n14280) );
  INV_X1 U8108 ( .A(n8254), .ZN(n6862) );
  INV_X1 U8109 ( .A(n8253), .ZN(n6863) );
  NAND2_X1 U8110 ( .A1(n8274), .A2(n8273), .ZN(n14293) );
  NAND2_X1 U8111 ( .A1(n14293), .A2(n14703), .ZN(n14290) );
  NAND2_X1 U8112 ( .A1(n6848), .A2(n6847), .ZN(n14292) );
  INV_X1 U8113 ( .A(n8273), .ZN(n6847) );
  INV_X1 U8114 ( .A(n8274), .ZN(n6848) );
  XNOR2_X1 U8115 ( .A(n8278), .B(n7041), .ZN(n14425) );
  INV_X1 U8116 ( .A(n8277), .ZN(n7041) );
  INV_X1 U8117 ( .A(n14427), .ZN(n6855) );
  NAND2_X1 U8118 ( .A1(n6756), .A2(n6757), .ZN(n6850) );
  INV_X1 U8119 ( .A(n14299), .ZN(n6756) );
  OAI21_X1 U8120 ( .B1(n6850), .B2(n6552), .A(P2_ADDR_REG_18__SCAN_IN), .ZN(
        n6754) );
  XNOR2_X1 U8121 ( .A(n9661), .B(n8788), .ZN(n6904) );
  NAND2_X1 U8122 ( .A1(n13051), .A2(n11977), .ZN(n11931) );
  NAND2_X1 U8123 ( .A1(n8456), .A2(n8457), .ZN(n8455) );
  INV_X1 U8124 ( .A(n8469), .ZN(n7164) );
  OR2_X1 U8125 ( .A1(n11995), .A2(n6821), .ZN(n6820) );
  NOR2_X1 U8126 ( .A1(n11996), .A2(n11993), .ZN(n6822) );
  NAND2_X1 U8127 ( .A1(n6584), .A2(n7307), .ZN(n7305) );
  NOR2_X1 U8128 ( .A1(n6584), .A2(n7307), .ZN(n7306) );
  NAND2_X1 U8129 ( .A1(n6903), .A2(n8515), .ZN(n6902) );
  NAND2_X1 U8130 ( .A1(n8516), .A2(n8517), .ZN(n6903) );
  OR2_X1 U8131 ( .A1(n8516), .A2(n8517), .ZN(n6901) );
  MUX2_X1 U8132 ( .A(n11724), .B(n11723), .S(n11811), .Z(n11729) );
  NAND2_X1 U8133 ( .A1(n7308), .A2(n6626), .ZN(n12037) );
  AOI21_X1 U8134 ( .B1(n6827), .B2(n6830), .A(n6825), .ZN(n6824) );
  INV_X1 U8135 ( .A(n8579), .ZN(n8582) );
  OAI22_X1 U8136 ( .A1(n12047), .A2(n7321), .B1(n12045), .B2(n12046), .ZN(
        n12054) );
  AND2_X1 U8137 ( .A1(n12046), .A2(n12045), .ZN(n7321) );
  OAI21_X1 U8138 ( .B1(n11749), .B2(n11748), .A(n12717), .ZN(n11758) );
  OAI21_X1 U8139 ( .B1(n6927), .B2(n8619), .A(n7434), .ZN(n6923) );
  OR2_X1 U8140 ( .A1(n6925), .A2(n6560), .ZN(n6924) );
  NOR2_X1 U8141 ( .A1(n6927), .A2(n6926), .ZN(n6925) );
  AOI21_X1 U8142 ( .B1(n6561), .B2(n6836), .A(n6649), .ZN(n6832) );
  AND2_X1 U8143 ( .A1(n12062), .A2(n6837), .ZN(n6836) );
  OR2_X1 U8144 ( .A1(n7314), .A2(n6598), .ZN(n7313) );
  AOI21_X1 U8145 ( .B1(n6543), .B2(n6840), .A(n6643), .ZN(n6838) );
  AND2_X1 U8146 ( .A1(n12087), .A2(n6557), .ZN(n6840) );
  NAND2_X1 U8147 ( .A1(n8683), .A2(n8684), .ZN(n8682) );
  INV_X1 U8148 ( .A(n7872), .ZN(n7536) );
  AND2_X1 U8149 ( .A1(n7804), .A2(n7515), .ZN(n7526) );
  NOR2_X1 U8150 ( .A1(n7525), .A2(n7524), .ZN(n7431) );
  INV_X1 U8151 ( .A(P3_IR_REG_25__SCAN_IN), .ZN(n9377) );
  INV_X1 U8152 ( .A(P3_IR_REG_23__SCAN_IN), .ZN(n9374) );
  INV_X1 U8153 ( .A(n7662), .ZN(n7082) );
  INV_X1 U8154 ( .A(n7921), .ZN(n7548) );
  NAND2_X1 U8155 ( .A1(n7257), .A2(n7260), .ZN(n7255) );
  INV_X1 U8156 ( .A(n7257), .ZN(n7256) );
  INV_X1 U8157 ( .A(n7837), .ZN(n7234) );
  NOR2_X1 U8158 ( .A1(n7512), .A2(n7273), .ZN(n7272) );
  INV_X1 U8159 ( .A(n7511), .ZN(n7273) );
  INV_X1 U8160 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n8210) );
  NAND2_X1 U8161 ( .A1(n7345), .A2(n7344), .ZN(n7343) );
  INV_X1 U8162 ( .A(n12516), .ZN(n7344) );
  INV_X1 U8163 ( .A(n12474), .ZN(n7019) );
  OAI21_X1 U8164 ( .B1(n11801), .B2(n11613), .A(n11799), .ZN(n7399) );
  NOR2_X1 U8165 ( .A1(n6962), .A2(n6887), .ZN(n6886) );
  INV_X1 U8166 ( .A(n11614), .ZN(n6887) );
  INV_X1 U8167 ( .A(n11720), .ZN(n7376) );
  NOR2_X1 U8168 ( .A1(n7377), .A2(n7376), .ZN(n7375) );
  INV_X1 U8169 ( .A(n10747), .ZN(n7377) );
  INV_X1 U8170 ( .A(n11608), .ZN(n6953) );
  AND2_X1 U8171 ( .A1(n6955), .A2(n12614), .ZN(n6954) );
  NAND2_X1 U8172 ( .A1(n12633), .A2(n11608), .ZN(n6955) );
  OR2_X1 U8173 ( .A1(n6865), .A2(n10940), .ZN(n10386) );
  INV_X1 U8174 ( .A(n9090), .ZN(n6987) );
  NOR2_X1 U8175 ( .A1(n8869), .A2(P3_IR_REG_16__SCAN_IN), .ZN(n7012) );
  OR2_X1 U8176 ( .A1(n9091), .A2(n9087), .ZN(n9088) );
  INV_X1 U8177 ( .A(n7334), .ZN(n7333) );
  OAI21_X1 U8178 ( .B1(n9679), .B2(n7335), .A(n10116), .ZN(n7334) );
  INV_X1 U8179 ( .A(n10027), .ZN(n7335) );
  INV_X1 U8180 ( .A(n7328), .ZN(n7327) );
  OAI21_X1 U8181 ( .B1(n9496), .B2(n7329), .A(n9615), .ZN(n7328) );
  INV_X1 U8182 ( .A(n9527), .ZN(n7329) );
  AND2_X1 U8183 ( .A1(n7337), .A2(n9045), .ZN(n7336) );
  NAND2_X1 U8184 ( .A1(n6587), .A2(n9038), .ZN(n7337) );
  INV_X1 U8185 ( .A(n8971), .ZN(n7356) );
  INV_X1 U8186 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n8973) );
  INV_X1 U8187 ( .A(P3_IR_REG_2__SCAN_IN), .ZN(n8859) );
  XNOR2_X1 U8188 ( .A(n13406), .B(n6528), .ZN(n12890) );
  OAI21_X1 U8189 ( .B1(n6843), .B2(n12148), .A(n6639), .ZN(n6842) );
  NOR2_X1 U8190 ( .A1(n13351), .A2(n13356), .ZN(n6805) );
  INV_X1 U8191 ( .A(n12216), .ZN(n7106) );
  INV_X1 U8192 ( .A(n7894), .ZN(n7103) );
  NOR2_X1 U8193 ( .A1(n7882), .A2(n15294), .ZN(n7890) );
  NOR2_X1 U8194 ( .A1(n12050), .A2(n14356), .ZN(n6811) );
  INV_X1 U8195 ( .A(n7749), .ZN(n7096) );
  INV_X1 U8196 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n7724) );
  OR2_X1 U8197 ( .A1(n7725), .A2(n7724), .ZN(n7742) );
  INV_X1 U8198 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n7854) );
  INV_X1 U8199 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n8064) );
  INV_X1 U8200 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n7737) );
  INV_X1 U8201 ( .A(n7614), .ZN(n7636) );
  INV_X1 U8202 ( .A(n8715), .ZN(n8716) );
  INV_X1 U8203 ( .A(n8699), .ZN(n8700) );
  NAND2_X1 U8204 ( .A1(P1_REG3_REG_25__SCAN_IN), .A2(n8716), .ZN(n8726) );
  AND2_X1 U8205 ( .A1(n13640), .A2(n14572), .ZN(n13603) );
  NAND2_X1 U8206 ( .A1(n8724), .A2(n6935), .ZN(n6934) );
  NAND2_X1 U8207 ( .A1(n6937), .A2(n8723), .ZN(n6936) );
  NOR2_X1 U8208 ( .A1(n7295), .A2(n7294), .ZN(n7293) );
  INV_X1 U8209 ( .A(n13875), .ZN(n7281) );
  NAND2_X1 U8210 ( .A1(n7435), .A2(n10806), .ZN(n7276) );
  AND2_X1 U8211 ( .A1(n14599), .A2(n14548), .ZN(n9756) );
  NAND2_X1 U8212 ( .A1(n6775), .A2(n6624), .ZN(n9749) );
  NAND2_X1 U8213 ( .A1(n8017), .A2(n8016), .ZN(n8036) );
  OAI21_X1 U8214 ( .B1(n7988), .B2(n7265), .A(n7263), .ZN(n8017) );
  AOI21_X1 U8215 ( .B1(n7266), .B2(n7264), .A(n6703), .ZN(n7263) );
  INV_X1 U8216 ( .A(n7241), .ZN(n7240) );
  AND2_X1 U8217 ( .A1(n7544), .A2(n7901), .ZN(n7919) );
  AND2_X1 U8218 ( .A1(n7261), .A2(n7537), .ZN(n7257) );
  NOR2_X1 U8219 ( .A1(n7540), .A2(n7539), .ZN(n7261) );
  INV_X1 U8220 ( .A(n7902), .ZN(n7540) );
  NOR2_X1 U8221 ( .A1(n7538), .A2(n9619), .ZN(n7539) );
  NAND2_X1 U8222 ( .A1(n7542), .A2(SI_19_), .ZN(n7902) );
  INV_X1 U8223 ( .A(n7160), .ZN(n8598) );
  AND2_X1 U8224 ( .A1(n7781), .A2(n7517), .ZN(n7804) );
  AND2_X1 U8225 ( .A1(n7765), .A2(n7519), .ZN(n7781) );
  NAND2_X1 U8226 ( .A1(n7503), .A2(SI_7_), .ZN(n7505) );
  AOI21_X1 U8227 ( .B1(n7249), .B2(n7250), .A(n7247), .ZN(n7246) );
  INV_X1 U8228 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n6758) );
  NAND2_X1 U8229 ( .A1(n6760), .A2(P1_ADDR_REG_1__SCAN_IN), .ZN(n6759) );
  XNOR2_X1 U8230 ( .A(n8210), .B(P3_ADDR_REG_2__SCAN_IN), .ZN(n8245) );
  XNOR2_X1 U8231 ( .A(n7043), .B(P3_ADDR_REG_3__SCAN_IN), .ZN(n8244) );
  NOR2_X1 U8232 ( .A1(n7007), .A2(n12592), .ZN(n7002) );
  NOR2_X1 U8233 ( .A1(n12330), .A2(n6542), .ZN(n7006) );
  AND2_X1 U8234 ( .A1(n11171), .A2(n11168), .ZN(n11169) );
  NAND2_X1 U8235 ( .A1(n12270), .A2(n11877), .ZN(n11880) );
  AND2_X1 U8236 ( .A1(n11072), .A2(n11071), .ZN(n15398) );
  INV_X1 U8237 ( .A(n12288), .ZN(n6991) );
  INV_X1 U8238 ( .A(n15392), .ZN(n12332) );
  NAND2_X1 U8239 ( .A1(n11819), .A2(n12786), .ZN(n7384) );
  OR2_X1 U8240 ( .A1(n6865), .A2(n10256), .ZN(n6866) );
  OR2_X1 U8241 ( .A1(n6865), .A2(n12631), .ZN(n9384) );
  OR2_X1 U8242 ( .A1(n8874), .A2(n11005), .ZN(n9795) );
  AND2_X1 U8243 ( .A1(n9989), .A2(n10038), .ZN(n10031) );
  NAND2_X1 U8244 ( .A1(n14878), .A2(n10904), .ZN(n14898) );
  OR2_X1 U8245 ( .A1(n14868), .A2(n10928), .ZN(n7023) );
  NAND2_X1 U8246 ( .A1(n6726), .A2(n6725), .ZN(n14884) );
  INV_X1 U8247 ( .A(n14886), .ZN(n6725) );
  INV_X1 U8248 ( .A(n14887), .ZN(n6726) );
  AND2_X1 U8249 ( .A1(n14884), .A2(n10892), .ZN(n10893) );
  NAND2_X1 U8250 ( .A1(n14914), .A2(n10907), .ZN(n14933) );
  NAND2_X1 U8251 ( .A1(n14949), .A2(n10909), .ZN(n14972) );
  NAND2_X1 U8252 ( .A1(n7022), .A2(n7021), .ZN(n7020) );
  NAND2_X1 U8253 ( .A1(n14965), .A2(P3_REG2_REG_10__SCAN_IN), .ZN(n7021) );
  NAND2_X1 U8254 ( .A1(n11127), .A2(n11128), .ZN(n12366) );
  AND2_X1 U8255 ( .A1(n12362), .A2(n11124), .ZN(n12372) );
  NOR2_X1 U8256 ( .A1(n12383), .A2(n12372), .ZN(n12374) );
  NAND2_X1 U8257 ( .A1(n12377), .A2(n12378), .ZN(n12379) );
  NAND2_X1 U8258 ( .A1(n12379), .A2(n12385), .ZN(n12398) );
  NAND2_X1 U8259 ( .A1(n12398), .A2(n12401), .ZN(n12421) );
  NAND2_X1 U8260 ( .A1(n7036), .A2(P3_REG2_REG_15__SCAN_IN), .ZN(n7033) );
  NAND2_X1 U8261 ( .A1(n12418), .A2(n7036), .ZN(n7032) );
  NAND2_X1 U8262 ( .A1(n6568), .A2(P3_REG2_REG_17__SCAN_IN), .ZN(n12476) );
  NAND2_X1 U8263 ( .A1(n12443), .A2(n6708), .ZN(n12460) );
  OR2_X1 U8264 ( .A1(n11518), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n11520) );
  NAND2_X1 U8265 ( .A1(n11504), .A2(n9468), .ZN(n11518) );
  NOR2_X1 U8266 ( .A1(n11270), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n11321) );
  NOR2_X1 U8267 ( .A1(n11055), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n11088) );
  AND4_X1 U8268 ( .A1(n10575), .A2(n10574), .A3(n10573), .A4(n10572), .ZN(
        n15393) );
  INV_X1 U8269 ( .A(n15398), .ZN(n14321) );
  OR2_X1 U8270 ( .A1(n10570), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n10580) );
  INV_X1 U8271 ( .A(P3_REG3_REG_8__SCAN_IN), .ZN(n10798) );
  AND2_X1 U8272 ( .A1(n10532), .A2(n10798), .ZN(n10558) );
  AND2_X1 U8273 ( .A1(n11046), .A2(n11045), .ZN(n11048) );
  NAND2_X1 U8274 ( .A1(n10753), .A2(n10752), .ZN(n11046) );
  NOR2_X1 U8275 ( .A1(n10384), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n10532) );
  OR2_X1 U8276 ( .A1(n10267), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n10384) );
  NOR2_X1 U8277 ( .A1(P3_REG3_REG_3__SCAN_IN), .A2(P3_REG3_REG_4__SCAN_IN), 
        .ZN(n10209) );
  AND2_X1 U8278 ( .A1(n11699), .A2(n11696), .ZN(n11825) );
  OR2_X1 U8279 ( .A1(n6530), .A2(n10915), .ZN(n9972) );
  INV_X1 U8280 ( .A(n11845), .ZN(n11618) );
  NAND2_X1 U8281 ( .A1(n11809), .A2(n11816), .ZN(n11845) );
  NAND2_X1 U8282 ( .A1(n6880), .A2(n6879), .ZN(n12515) );
  AOI21_X1 U8283 ( .B1(n6882), .B2(n6884), .A(n6648), .ZN(n6879) );
  NAND2_X1 U8284 ( .A1(n11814), .A2(n11812), .ZN(n12516) );
  OR2_X1 U8285 ( .A1(n11887), .A2(n12331), .ZN(n11614) );
  INV_X1 U8286 ( .A(n11612), .ZN(n6871) );
  INV_X1 U8287 ( .A(n12574), .ZN(n12572) );
  AND2_X1 U8288 ( .A1(n11791), .A2(n11792), .ZN(n12587) );
  INV_X1 U8289 ( .A(n7405), .ZN(n7404) );
  OAI21_X1 U8290 ( .B1(n7406), .B2(n11509), .A(n11788), .ZN(n7405) );
  NAND2_X1 U8291 ( .A1(n12625), .A2(n11608), .ZN(n12613) );
  NAND2_X1 U8292 ( .A1(n6950), .A2(n6954), .ZN(n12612) );
  NAND2_X1 U8293 ( .A1(n12623), .A2(n11608), .ZN(n6950) );
  AND3_X1 U8294 ( .A1(n11507), .A2(n11506), .A3(n11505), .ZN(n12627) );
  OR2_X1 U8295 ( .A1(n12623), .A2(n12633), .ZN(n12625) );
  AND2_X1 U8296 ( .A1(n11778), .A2(n12610), .ZN(n12633) );
  NAND2_X1 U8297 ( .A1(n12658), .A2(n12662), .ZN(n7390) );
  INV_X1 U8298 ( .A(n12659), .ZN(n12662) );
  AND4_X1 U8299 ( .A1(n11275), .A2(n11274), .A3(n11273), .A4(n11272), .ZN(
        n12678) );
  OR2_X1 U8300 ( .A1(n6865), .A2(n12693), .ZN(n11274) );
  AND2_X1 U8301 ( .A1(n11764), .A2(n11763), .ZN(n12676) );
  NAND2_X1 U8302 ( .A1(n11317), .A2(n11316), .ZN(n11601) );
  AND2_X1 U8303 ( .A1(n11760), .A2(n11759), .ZN(n12689) );
  INV_X1 U8304 ( .A(n7395), .ZN(n7394) );
  AOI21_X1 U8305 ( .B1(n7395), .B2(n7393), .A(n12714), .ZN(n7392) );
  AND4_X1 U8306 ( .A1(n10214), .A2(n10213), .A3(n10212), .A4(n10211), .ZN(
        n10638) );
  OR2_X1 U8307 ( .A1(n6530), .A2(n10928), .ZN(n10211) );
  NAND2_X1 U8308 ( .A1(n9088), .A2(n9089), .ZN(n9090) );
  XNOR2_X1 U8309 ( .A(n9380), .B(P3_IR_REG_29__SCAN_IN), .ZN(n9381) );
  NAND2_X1 U8310 ( .A1(n11114), .A2(n11113), .ZN(n11117) );
  INV_X1 U8311 ( .A(P3_IR_REG_26__SCAN_IN), .ZN(n9373) );
  OR2_X1 U8312 ( .A1(n8876), .A2(P3_IR_REG_24__SCAN_IN), .ZN(n8872) );
  NAND2_X1 U8313 ( .A1(n11000), .A2(n10999), .ZN(n11003) );
  OAI21_X1 U8314 ( .B1(n10791), .B2(n7367), .A(n7366), .ZN(n10884) );
  NAND2_X1 U8315 ( .A1(P1_DATAO_REG_24__SCAN_IN), .A2(n7368), .ZN(n7366) );
  NOR2_X1 U8316 ( .A1(P1_DATAO_REG_24__SCAN_IN), .A2(n7368), .ZN(n7367) );
  NAND2_X1 U8317 ( .A1(n9701), .A2(n9700), .ZN(n9704) );
  NAND2_X1 U8318 ( .A1(n9626), .A2(n9625), .ZN(n9629) );
  NAND2_X1 U8319 ( .A1(n9624), .A2(n9623), .ZN(n9626) );
  NAND2_X1 U8320 ( .A1(n9291), .A2(n9290), .ZN(n9294) );
  NAND2_X1 U8321 ( .A1(n9294), .A2(n9293), .ZN(n9494) );
  NAND2_X1 U8322 ( .A1(n9200), .A2(n9199), .ZN(n9203) );
  OAI21_X1 U8323 ( .B1(n9075), .B2(n7364), .A(n7362), .ZN(n9199) );
  AND2_X1 U8324 ( .A1(n9290), .A2(n9201), .ZN(n9202) );
  NAND2_X1 U8325 ( .A1(n9203), .A2(n9202), .ZN(n9291) );
  AOI21_X1 U8326 ( .B1(n7362), .B2(n7364), .A(n7360), .ZN(n7359) );
  NOR2_X1 U8327 ( .A1(n6579), .A2(n7361), .ZN(n7360) );
  OR2_X1 U8328 ( .A1(n9154), .A2(n15367), .ZN(n9200) );
  NAND2_X1 U8329 ( .A1(n9010), .A2(n9009), .ZN(n14857) );
  AND2_X1 U8330 ( .A1(n8987), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n8970) );
  XNOR2_X1 U8331 ( .A(n8973), .B(P1_DATAO_REG_4__SCAN_IN), .ZN(n9006) );
  NAND2_X1 U8332 ( .A1(n8969), .A2(n8968), .ZN(n9013) );
  AND2_X1 U8333 ( .A1(n11281), .A2(n6745), .ZN(n7138) );
  INV_X1 U8334 ( .A(n11282), .ZN(n6745) );
  NAND2_X1 U8335 ( .A1(n7141), .A2(n7140), .ZN(n7139) );
  INV_X1 U8336 ( .A(n11284), .ZN(n7141) );
  NOR2_X1 U8337 ( .A1(n7742), .A2(n7741), .ZN(n7757) );
  AND2_X1 U8338 ( .A1(n7757), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n7772) );
  NAND2_X1 U8339 ( .A1(n7109), .A2(n7111), .ZN(n10075) );
  NAND2_X1 U8340 ( .A1(n7110), .A2(n6595), .ZN(n7109) );
  AND2_X1 U8341 ( .A1(n9829), .A2(n6595), .ZN(n7112) );
  NAND2_X1 U8342 ( .A1(n10075), .A2(n10074), .ZN(n10242) );
  NOR2_X1 U8343 ( .A1(n10841), .A2(n7121), .ZN(n7120) );
  INV_X1 U8344 ( .A(n10843), .ZN(n7121) );
  INV_X1 U8345 ( .A(n7122), .ZN(n7119) );
  INV_X1 U8346 ( .A(n7120), .ZN(n7118) );
  INV_X1 U8347 ( .A(n7966), .ZN(n7981) );
  XNOR2_X1 U8348 ( .A(n12032), .B(n6528), .ZN(n11281) );
  NOR2_X1 U8349 ( .A1(n7952), .A2(n12998), .ZN(n7967) );
  OR2_X1 U8350 ( .A1(n10621), .A2(n7123), .ZN(n7122) );
  INV_X1 U8351 ( .A(n10328), .ZN(n7123) );
  NOR2_X1 U8352 ( .A1(n7827), .A2(n7826), .ZN(n7843) );
  NAND2_X1 U8353 ( .A1(n11286), .A2(n11285), .ZN(n11373) );
  INV_X1 U8354 ( .A(n8199), .ZN(n8040) );
  OR2_X1 U8355 ( .A1(n14688), .A2(n14687), .ZN(n14690) );
  OR2_X1 U8356 ( .A1(n9318), .A2(n9317), .ZN(n14726) );
  INV_X1 U8357 ( .A(n6803), .ZN(n6800) );
  INV_X1 U8358 ( .A(n7994), .ZN(n7468) );
  NAND2_X1 U8359 ( .A1(n8151), .A2(n8033), .ZN(n13161) );
  INV_X1 U8360 ( .A(n7055), .ZN(n7053) );
  AOI21_X1 U8361 ( .B1(n7055), .B2(n7058), .A(n7052), .ZN(n7051) );
  XNOR2_X1 U8362 ( .A(n13187), .B(n13026), .ZN(n13181) );
  NOR2_X1 U8363 ( .A1(n7436), .A2(n13233), .ZN(n13228) );
  AND2_X1 U8364 ( .A1(n6556), .A2(n13456), .ZN(n6796) );
  NAND2_X1 U8365 ( .A1(n13308), .A2(n6550), .ZN(n13292) );
  AND2_X1 U8366 ( .A1(n7890), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n7910) );
  AND2_X1 U8367 ( .A1(n7910), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n7926) );
  NAND2_X1 U8368 ( .A1(n13308), .A2(n8168), .ZN(n13309) );
  NOR2_X1 U8369 ( .A1(n6583), .A2(n7070), .ZN(n7069) );
  NAND2_X1 U8370 ( .A1(n10990), .A2(n6807), .ZN(n13327) );
  NOR2_X1 U8371 ( .A1(n12065), .A2(n6809), .ZN(n6807) );
  NAND2_X1 U8372 ( .A1(n11342), .A2(n11341), .ZN(n7100) );
  AOI21_X1 U8373 ( .B1(n7048), .B2(n14358), .A(n6633), .ZN(n7047) );
  NAND2_X1 U8374 ( .A1(n10990), .A2(n6811), .ZN(n11406) );
  NAND2_X1 U8375 ( .A1(n10990), .A2(n8167), .ZN(n14360) );
  INV_X1 U8376 ( .A(n7078), .ZN(n7074) );
  NAND2_X1 U8377 ( .A1(n6814), .A2(n6813), .ZN(n10989) );
  AND2_X1 U8378 ( .A1(n6816), .A2(n10782), .ZN(n6813) );
  INV_X1 U8379 ( .A(n14379), .ZN(n6816) );
  INV_X1 U8380 ( .A(n14811), .ZN(n6815) );
  NAND2_X1 U8381 ( .A1(n6814), .A2(n10782), .ZN(n10772) );
  NAND2_X1 U8382 ( .A1(n10470), .A2(n14807), .ZN(n10489) );
  NOR2_X1 U8383 ( .A1(n10172), .A2(n14782), .ZN(n10183) );
  OR2_X1 U8384 ( .A1(n12940), .A2(n13144), .ZN(n9415) );
  NAND2_X1 U8385 ( .A1(n6706), .A2(n6795), .ZN(n10172) );
  NAND2_X1 U8386 ( .A1(n9539), .A2(n9541), .ZN(n9540) );
  AND2_X1 U8387 ( .A1(n13356), .A2(n14810), .ZN(n13357) );
  AND2_X1 U8388 ( .A1(n6538), .A2(n14803), .ZN(n14791) );
  AOI21_X1 U8389 ( .B1(n11257), .B2(n8076), .A(n13488), .ZN(n14765) );
  AND3_X1 U8390 ( .A1(n6555), .A2(n7738), .A3(n7108), .ZN(n7570) );
  AND2_X1 U8391 ( .A1(n7614), .A2(n7063), .ZN(n7062) );
  AND2_X1 U8392 ( .A1(n7066), .A2(n7460), .ZN(n7063) );
  INV_X1 U8393 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n7648) );
  NOR2_X1 U8394 ( .A1(n8934), .A2(n7175), .ZN(n7174) );
  INV_X1 U8395 ( .A(n8902), .ZN(n7175) );
  AOI21_X1 U8396 ( .B1(n13611), .B2(n13608), .A(n13634), .ZN(n7191) );
  INV_X1 U8397 ( .A(n7191), .ZN(n7189) );
  INV_X1 U8398 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n8518) );
  NAND2_X1 U8399 ( .A1(n7214), .A2(n7215), .ZN(n13669) );
  AOI21_X1 U8400 ( .B1(n7217), .B2(n7223), .A(n7216), .ZN(n7215) );
  INV_X1 U8401 ( .A(n13671), .ZN(n7216) );
  NAND2_X1 U8402 ( .A1(n7224), .A2(n6546), .ZN(n13617) );
  NAND2_X1 U8403 ( .A1(n13716), .A2(n7228), .ZN(n7224) );
  NAND2_X1 U8404 ( .A1(n10606), .A2(n10607), .ZN(n10674) );
  OR2_X1 U8405 ( .A1(n8648), .A2(n8647), .ZN(n8661) );
  NAND2_X1 U8406 ( .A1(n11239), .A2(n11238), .ZN(n13661) );
  OR2_X1 U8407 ( .A1(n8661), .A2(n13653), .ZN(n8673) );
  NOR2_X1 U8408 ( .A1(n15322), .A2(n8673), .ZN(n8689) );
  INV_X1 U8409 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n8519) );
  AOI21_X1 U8410 ( .B1(n6629), .B2(n7201), .A(n6732), .ZN(n11024) );
  OAI21_X1 U8411 ( .B1(n7203), .B2(n7202), .A(n6638), .ZN(n6732) );
  NOR2_X1 U8412 ( .A1(n8610), .A2(n8609), .ZN(n8625) );
  AND2_X1 U8413 ( .A1(n8625), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n8636) );
  NAND2_X1 U8414 ( .A1(n13690), .A2(n13536), .ZN(n7198) );
  NAND2_X1 U8415 ( .A1(n13692), .A2(n7199), .ZN(n7197) );
  NAND2_X1 U8416 ( .A1(n13669), .A2(n13599), .ZN(n13732) );
  AND2_X1 U8417 ( .A1(n8555), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n8566) );
  NAND2_X1 U8418 ( .A1(n14394), .A2(n13515), .ZN(n7172) );
  INV_X1 U8419 ( .A(n13603), .ZN(n13548) );
  AND2_X1 U8420 ( .A1(n6916), .A2(n6915), .ZN(n6914) );
  INV_X1 U8421 ( .A(n7154), .ZN(n6915) );
  NAND2_X1 U8422 ( .A1(n6913), .A2(n7153), .ZN(n6912) );
  NAND2_X1 U8423 ( .A1(n6914), .A2(n6558), .ZN(n6913) );
  AOI21_X1 U8424 ( .B1(n7154), .B2(n7153), .A(n7152), .ZN(n7151) );
  NAND2_X1 U8425 ( .A1(n9100), .A2(n13787), .ZN(n13811) );
  CLKBUF_X1 U8426 ( .A(n8378), .Z(n8379) );
  OR2_X1 U8427 ( .A1(n9160), .A2(n9161), .ZN(n9158) );
  NOR2_X1 U8428 ( .A1(n14458), .A2(n14457), .ZN(n14456) );
  OAI22_X1 U8429 ( .A1(n13824), .A2(n13823), .B1(n13822), .B2(n13821), .ZN(
        n13833) );
  AND2_X1 U8430 ( .A1(n7292), .A2(n6655), .ZN(n7290) );
  INV_X1 U8431 ( .A(n7293), .ZN(n7289) );
  NAND2_X1 U8432 ( .A1(n13965), .A2(n7293), .ZN(n7291) );
  OR2_X1 U8433 ( .A1(n13948), .A2(n7295), .ZN(n7292) );
  OR2_X1 U8434 ( .A1(n14143), .A2(n13945), .ZN(n8809) );
  AOI21_X1 U8435 ( .B1(n13965), .B2(n13941), .A(n13884), .ZN(n13944) );
  AND2_X1 U8436 ( .A1(n13989), .A2(n6605), .ZN(n7299) );
  AND2_X1 U8437 ( .A1(n7298), .A2(n6605), .ZN(n13977) );
  AND2_X1 U8438 ( .A1(n13987), .A2(n6569), .ZN(n6981) );
  NAND2_X1 U8439 ( .A1(n6547), .A2(n14070), .ZN(n6778) );
  NAND2_X1 U8440 ( .A1(n14042), .A2(n6983), .ZN(n14013) );
  NAND2_X1 U8441 ( .A1(n14042), .A2(n14033), .ZN(n14028) );
  OR2_X1 U8442 ( .A1(n14113), .A2(n14096), .ZN(n14098) );
  INV_X1 U8443 ( .A(n7418), .ZN(n7417) );
  AOI21_X1 U8444 ( .B1(n13894), .B2(n13893), .A(n7423), .ZN(n7418) );
  NAND2_X1 U8445 ( .A1(n14112), .A2(n14120), .ZN(n14113) );
  NAND2_X1 U8446 ( .A1(n6968), .A2(n6967), .ZN(n11391) );
  INV_X1 U8447 ( .A(n11306), .ZN(n6968) );
  NAND2_X1 U8448 ( .A1(n6970), .A2(n6969), .ZN(n11306) );
  NOR2_X1 U8449 ( .A1(n8536), .A2(n8535), .ZN(n8555) );
  OR3_X1 U8450 ( .A1(n8520), .A2(n8519), .A3(n8518), .ZN(n8536) );
  AND4_X1 U8451 ( .A1(n8560), .A2(n8559), .A3(n8558), .A4(n8557), .ZN(n13506)
         );
  NOR2_X1 U8452 ( .A1(n8474), .A2(n8473), .ZN(n8495) );
  NAND2_X1 U8453 ( .A1(n8495), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n8520) );
  NOR2_X1 U8454 ( .A1(n8411), .A2(n9162), .ZN(n8434) );
  NAND2_X1 U8455 ( .A1(n9756), .A2(n6548), .ZN(n14531) );
  INV_X1 U8456 ( .A(n9860), .ZN(n9852) );
  AND2_X1 U8457 ( .A1(n9756), .A2(n9854), .ZN(n14532) );
  AND2_X1 U8458 ( .A1(n13637), .A2(n9247), .ZN(n9658) );
  NOR2_X1 U8459 ( .A1(n6603), .A2(n6978), .ZN(n6977) );
  NAND2_X1 U8460 ( .A1(n14138), .A2(n14137), .ZN(n6978) );
  AND3_X1 U8461 ( .A1(n8640), .A2(n8639), .A3(n8638), .ZN(n14210) );
  INV_X1 U8462 ( .A(n14607), .ZN(n14638) );
  XNOR2_X1 U8463 ( .A(n8192), .B(n8191), .ZN(n8795) );
  XNOR2_X1 U8464 ( .A(n8178), .B(n8177), .ZN(n11636) );
  INV_X1 U8465 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n8331) );
  XNOR2_X1 U8466 ( .A(n8036), .B(n8035), .ZN(n11638) );
  INV_X1 U8467 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n8333) );
  NOR2_X2 U8468 ( .A1(n8341), .A2(n8307), .ZN(n7439) );
  INV_X1 U8469 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n8306) );
  INV_X1 U8470 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n8317) );
  INV_X1 U8471 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n8316) );
  NAND2_X1 U8472 ( .A1(n7269), .A2(n7268), .ZN(n8014) );
  XNOR2_X1 U8473 ( .A(n7988), .B(n7987), .ZN(n11256) );
  AND2_X1 U8474 ( .A1(n8851), .A2(n8852), .ZN(n8924) );
  OR2_X1 U8475 ( .A1(n7160), .A2(n8341), .ZN(n8345) );
  NAND2_X1 U8476 ( .A1(n7535), .A2(n7534), .ZN(n7874) );
  NAND2_X1 U8477 ( .A1(n7528), .A2(n7235), .ZN(n7838) );
  NAND2_X1 U8478 ( .A1(n7644), .A2(n7496), .ZN(n7664) );
  NAND2_X1 U8479 ( .A1(n7236), .A2(n7490), .ZN(n7619) );
  NAND2_X1 U8480 ( .A1(n7487), .A2(n7490), .ZN(n7617) );
  OAI21_X1 U8481 ( .B1(n7488), .B2(P2_DATAO_REG_0__SCAN_IN), .A(n6748), .ZN(
        n7481) );
  NAND2_X1 U8482 ( .A1(n7488), .A2(n8954), .ZN(n6748) );
  INV_X1 U8483 ( .A(P3_ADDR_REG_0__SCAN_IN), .ZN(n9882) );
  XNOR2_X1 U8484 ( .A(n6860), .B(n8248), .ZN(n8250) );
  NAND2_X1 U8485 ( .A1(n14278), .A2(n14280), .ZN(n8256) );
  XNOR2_X1 U8486 ( .A(n8242), .B(n8241), .ZN(n8243) );
  NAND2_X1 U8487 ( .A1(n15410), .A2(n8261), .ZN(n8265) );
  AND2_X1 U8488 ( .A1(n6764), .A2(n6659), .ZN(n8262) );
  NAND2_X1 U8489 ( .A1(n8240), .A2(n15281), .ZN(n6764) );
  NOR2_X1 U8490 ( .A1(n8218), .A2(n8219), .ZN(n8272) );
  AND2_X1 U8491 ( .A1(n14290), .A2(n14292), .ZN(n8276) );
  NOR2_X1 U8492 ( .A1(n8224), .A2(n8223), .ZN(n8235) );
  NOR2_X1 U8493 ( .A1(n8237), .A2(n8236), .ZN(n8223) );
  OAI22_X1 U8494 ( .A1(P1_ADDR_REG_13__SCAN_IN), .A2(n8228), .B1(n8280), .B2(
        n8227), .ZN(n8282) );
  OR2_X1 U8495 ( .A1(n14427), .A2(n6858), .ZN(n6854) );
  AOI21_X1 U8496 ( .B1(n14427), .B2(n6858), .A(n6762), .ZN(n6761) );
  OAI21_X1 U8497 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(n12429), .A(n8292), .ZN(
        n8295) );
  INV_X1 U8498 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n6852) );
  NAND2_X1 U8499 ( .A1(n11561), .A2(n11560), .ZN(n12532) );
  OR2_X1 U8500 ( .A1(n11559), .A2(n10001), .ZN(n11561) );
  AOI22_X1 U8501 ( .A1(n12246), .A2(n12247), .B1(n12521), .B2(n11895), .ZN(
        n11897) );
  AND4_X1 U8502 ( .A1(n11093), .A2(n11092), .A3(n11091), .A4(n11090), .ZN(
        n11589) );
  INV_X1 U8503 ( .A(n14309), .ZN(n11592) );
  INV_X1 U8504 ( .A(n12552), .ZN(n12283) );
  AND2_X1 U8505 ( .A1(n11428), .A2(n11427), .ZN(n11483) );
  NAND2_X1 U8506 ( .A1(n6996), .A2(n6994), .ZN(n11432) );
  AOI21_X1 U8507 ( .B1(n6559), .B2(n7000), .A(n6995), .ZN(n6994) );
  INV_X1 U8508 ( .A(n11429), .ZN(n6995) );
  AND3_X1 U8509 ( .A1(n10261), .A2(n10260), .A3(n10259), .ZN(n10710) );
  AND4_X1 U8510 ( .A1(n9508), .A2(n9507), .A3(n9506), .A4(n9505), .ZN(n12626)
         );
  OR2_X1 U8511 ( .A1(n6865), .A2(n12472), .ZN(n9507) );
  NAND2_X1 U8512 ( .A1(n12289), .A2(n12288), .ZN(n12287) );
  NAND2_X1 U8513 ( .A1(n11867), .A2(n6993), .ZN(n12289) );
  AND3_X1 U8514 ( .A1(n10556), .A2(n10555), .A3(n10554), .ZN(n11730) );
  OR2_X1 U8515 ( .A1(n10193), .A2(n9728), .ZN(n9732) );
  OR2_X1 U8516 ( .A1(n10395), .A2(n11862), .ZN(n15392) );
  NAND2_X1 U8517 ( .A1(n11170), .A2(n11169), .ZN(n11268) );
  CLKBUF_X1 U8518 ( .A(n10010), .Z(n10006) );
  OAI21_X1 U8519 ( .B1(n11867), .B2(n6991), .A(n6989), .ZN(n12320) );
  NAND2_X1 U8520 ( .A1(n11490), .A2(n11489), .ZN(n12764) );
  NAND2_X1 U8521 ( .A1(n12295), .A2(n6542), .ZN(n7003) );
  NAND2_X1 U8522 ( .A1(n9814), .A2(n10396), .ZN(n15401) );
  AOI21_X1 U8523 ( .B1(n10398), .B2(n15050), .A(n9818), .ZN(n12338) );
  NAND2_X1 U8524 ( .A1(n6997), .A2(n6998), .ZN(n11430) );
  OR2_X1 U8525 ( .A1(n11170), .A2(n7000), .ZN(n6997) );
  AND2_X1 U8526 ( .A1(n10303), .A2(n10225), .ZN(n12520) );
  INV_X1 U8527 ( .A(n12627), .ZN(n12603) );
  INV_X1 U8528 ( .A(n12626), .ZN(n12665) );
  NOR2_X1 U8529 ( .A1(n6865), .A2(n12668), .ZN(n11440) );
  NOR2_X1 U8530 ( .A1(n6865), .A2(n12683), .ZN(n11326) );
  INV_X1 U8531 ( .A(n12678), .ZN(n12703) );
  OR3_X1 U8532 ( .A1(n11178), .A2(n11177), .A3(n11176), .ZN(n12719) );
  NOR2_X1 U8533 ( .A1(n6865), .A2(n12705), .ZN(n11176) );
  INV_X1 U8534 ( .A(n11589), .ZN(n14304) );
  OR3_X1 U8535 ( .A1(n11081), .A2(n11080), .A3(n11079), .ZN(n15388) );
  OR3_X1 U8536 ( .A1(n10588), .A2(n10587), .A3(n10586), .ZN(n14984) );
  NOR2_X1 U8537 ( .A1(n6865), .A2(n10584), .ZN(n10587) );
  INV_X1 U8538 ( .A(n15393), .ZN(n12342) );
  OR3_X1 U8539 ( .A1(n10564), .A2(n10563), .A3(n10562), .ZN(n14985) );
  NOR2_X1 U8540 ( .A1(n6865), .A2(n10953), .ZN(n10563) );
  OR3_X1 U8541 ( .A1(n10538), .A2(n10537), .A3(n10536), .ZN(n12343) );
  NOR2_X1 U8542 ( .A1(n6865), .A2(n10946), .ZN(n10537) );
  INV_X1 U8543 ( .A(n10708), .ZN(n12345) );
  OR2_X1 U8544 ( .A1(n11436), .A2(n9713), .ZN(n9716) );
  NOR2_X1 U8545 ( .A1(n15205), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n9989) );
  INV_X1 U8546 ( .A(n14961), .ZN(n14838) );
  AND2_X1 U8547 ( .A1(n7030), .A2(n10917), .ZN(n7029) );
  INV_X1 U8548 ( .A(n7023), .ZN(n14867) );
  XNOR2_X1 U8549 ( .A(n10893), .B(n10941), .ZN(n14904) );
  NOR2_X1 U8550 ( .A1(n14904), .A2(n10940), .ZN(n14903) );
  INV_X1 U8551 ( .A(n7028), .ZN(n14920) );
  INV_X1 U8552 ( .A(n7026), .ZN(n10895) );
  INV_X1 U8553 ( .A(n7022), .ZN(n14955) );
  XNOR2_X1 U8554 ( .A(n7020), .B(n11132), .ZN(n10897) );
  AND2_X1 U8555 ( .A1(n9083), .A2(n7381), .ZN(n12360) );
  NOR2_X1 U8556 ( .A1(n11125), .A2(n11086), .ZN(n12373) );
  OAI21_X1 U8557 ( .B1(n11125), .B2(n7038), .A(n7037), .ZN(n12396) );
  NAND2_X1 U8558 ( .A1(n12386), .A2(P3_REG2_REG_13__SCAN_IN), .ZN(n7038) );
  NAND2_X1 U8559 ( .A1(n12374), .A2(n12386), .ZN(n7037) );
  XNOR2_X1 U8560 ( .A(n12421), .B(n12432), .ZN(n12399) );
  INV_X1 U8561 ( .A(n7035), .ZN(n12417) );
  INV_X1 U8562 ( .A(n12418), .ZN(n7034) );
  NAND2_X1 U8563 ( .A1(n7032), .A2(n7031), .ZN(n12454) );
  XNOR2_X1 U8564 ( .A(n12460), .B(n6892), .ZN(n12461) );
  AND2_X1 U8565 ( .A1(n12476), .A2(n6744), .ZN(n12478) );
  AND2_X1 U8566 ( .A1(n12475), .A2(n12474), .ZN(n6744) );
  INV_X1 U8567 ( .A(n12497), .ZN(n6897) );
  AOI21_X1 U8568 ( .B1(n12882), .B2(n11664), .A(n11663), .ZN(n12511) );
  OR2_X1 U8569 ( .A1(n12506), .A2(n10355), .ZN(n12525) );
  INV_X1 U8570 ( .A(n6958), .ZN(n6957) );
  NAND2_X1 U8571 ( .A1(n12528), .A2(n6960), .ZN(n6959) );
  AOI22_X1 U8572 ( .A1(n11616), .A2(n15038), .B1(n15041), .B2(n12552), .ZN(
        n6958) );
  NAND2_X1 U8573 ( .A1(n11528), .A2(n11527), .ZN(n12584) );
  NAND2_X1 U8574 ( .A1(n11500), .A2(n11499), .ZN(n12758) );
  OR2_X1 U8575 ( .A1(n11497), .A2(n10001), .ZN(n11500) );
  NAND2_X1 U8576 ( .A1(n14980), .A2(n11479), .ZN(n7391) );
  NAND2_X1 U8577 ( .A1(n14313), .A2(n11479), .ZN(n14315) );
  INV_X1 U8578 ( .A(n7441), .ZN(n7378) );
  NAND2_X1 U8579 ( .A1(n10635), .A2(n10373), .ZN(n10706) );
  OR2_X1 U8580 ( .A1(n15052), .A2(n15010), .ZN(n12725) );
  NAND2_X1 U8581 ( .A1(n11653), .A2(n11652), .ZN(n12730) );
  AND2_X1 U8582 ( .A1(n15096), .A2(n15049), .ZN(n12782) );
  AND2_X2 U8583 ( .A1(n10088), .A2(n9712), .ZN(n15096) );
  INV_X1 U8584 ( .A(n12511), .ZN(n12786) );
  NAND2_X1 U8585 ( .A1(n11584), .A2(n11583), .ZN(n11917) );
  NAND2_X1 U8586 ( .A1(n11580), .A2(n11579), .ZN(n12794) );
  OAI21_X1 U8587 ( .B1(n11549), .B2(n10001), .A(n11551), .ZN(n12801) );
  AND2_X1 U8588 ( .A1(n7397), .A2(n11613), .ZN(n12539) );
  OR2_X1 U8589 ( .A1(n12563), .A2(n7402), .ZN(n7397) );
  NAND2_X1 U8590 ( .A1(n11542), .A2(n11541), .ZN(n12807) );
  OR2_X1 U8591 ( .A1(n11662), .A2(n11540), .ZN(n11541) );
  AND2_X1 U8592 ( .A1(n12554), .A2(n12553), .ZN(n12806) );
  NAND2_X1 U8593 ( .A1(n11517), .A2(n11516), .ZN(n12819) );
  INV_X1 U8594 ( .A(n7403), .ZN(n12599) );
  AOI21_X1 U8595 ( .B1(n12634), .B2(n11509), .A(n7406), .ZN(n7403) );
  AND2_X1 U8596 ( .A1(n11495), .A2(n11494), .ZN(n12835) );
  INV_X1 U8597 ( .A(n11483), .ZN(n12850) );
  INV_X1 U8598 ( .A(n12867), .ZN(n12870) );
  AND2_X1 U8599 ( .A1(n10402), .A2(n10401), .ZN(n15086) );
  OR2_X1 U8600 ( .A1(n15086), .A2(n15018), .ZN(n12867) );
  AOI21_X1 U8601 ( .B1(n6877), .B2(n9718), .A(n9718), .ZN(n6875) );
  XNOR2_X1 U8602 ( .A(n9373), .B(n8873), .ZN(n11005) );
  OAI21_X1 U8603 ( .B1(n8872), .B2(P3_IR_REG_25__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n8873) );
  NAND2_X1 U8604 ( .A1(n7370), .A2(n7369), .ZN(n10881) );
  NAND2_X1 U8605 ( .A1(n10791), .A2(n11228), .ZN(n7369) );
  OR2_X1 U8606 ( .A1(n10791), .A2(n11228), .ZN(n7370) );
  NAND2_X1 U8607 ( .A1(n10028), .A2(n10027), .ZN(n10117) );
  INV_X1 U8608 ( .A(n12489), .ZN(n12501) );
  NAND2_X1 U8609 ( .A1(n9528), .A2(n9527), .ZN(n9616) );
  OR2_X1 U8610 ( .A1(n9198), .A2(n9197), .ZN(n12400) );
  INV_X1 U8611 ( .A(SI_13_), .ZN(n11163) );
  INV_X1 U8612 ( .A(SI_12_), .ZN(n15330) );
  NAND2_X1 U8613 ( .A1(n9075), .A2(n6579), .ZN(n9153) );
  NAND2_X1 U8614 ( .A1(n9075), .A2(n9074), .ZN(n9078) );
  INV_X1 U8615 ( .A(SI_11_), .ZN(n11070) );
  OAI21_X1 U8616 ( .B1(n9037), .B2(n6587), .A(n9038), .ZN(n9046) );
  NAND2_X1 U8617 ( .A1(n8960), .A2(n9022), .ZN(n14928) );
  NAND2_X1 U8618 ( .A1(n7347), .A2(n7348), .ZN(n9018) );
  NAND2_X1 U8619 ( .A1(n7351), .A2(n8979), .ZN(n8996) );
  NAND2_X1 U8620 ( .A1(n7352), .A2(n8984), .ZN(n7351) );
  INV_X1 U8621 ( .A(n8985), .ZN(n7352) );
  INV_X1 U8622 ( .A(n10917), .ZN(n14842) );
  NAND2_X1 U8623 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(P3_IR_REG_0__SCAN_IN), .ZN(
        n8955) );
  INV_X1 U8624 ( .A(SI_0_), .ZN(n9728) );
  INV_X1 U8625 ( .A(P3_IR_REG_0__SCAN_IN), .ZN(n9883) );
  OAI21_X1 U8626 ( .B1(n12966), .B2(n7147), .A(n7145), .ZN(n7149) );
  INV_X1 U8627 ( .A(n7148), .ZN(n7147) );
  AOI21_X1 U8628 ( .B1(n7148), .B2(n7146), .A(n6644), .ZN(n7145) );
  NAND2_X1 U8629 ( .A1(n12919), .A2(n12918), .ZN(n12939) );
  NAND2_X1 U8630 ( .A1(n7139), .A2(n7136), .ZN(n14338) );
  INV_X1 U8631 ( .A(n7138), .ZN(n7136) );
  NAND2_X1 U8632 ( .A1(n10329), .A2(n10328), .ZN(n10622) );
  NAND2_X1 U8633 ( .A1(n7129), .A2(n7130), .ZN(n7128) );
  OAI21_X1 U8634 ( .B1(n12987), .B2(n12983), .A(n12984), .ZN(n12956) );
  AOI21_X1 U8635 ( .B1(n7133), .B2(n7135), .A(n6571), .ZN(n7132) );
  AOI21_X1 U8636 ( .B1(n12924), .B2(n12925), .A(n6749), .ZN(n12976) );
  NAND2_X1 U8637 ( .A1(n12976), .A2(n12975), .ZN(n12974) );
  MUX2_X1 U8638 ( .A(n7603), .B(n13489), .S(n9273), .Z(n11922) );
  NAND2_X1 U8639 ( .A1(n7925), .A2(n7924), .ZN(n13402) );
  NAND2_X1 U8640 ( .A1(n7115), .A2(n10620), .ZN(n10840) );
  OR2_X1 U8641 ( .A1(n7124), .A2(n7122), .ZN(n7115) );
  INV_X1 U8642 ( .A(n10329), .ZN(n7124) );
  AND2_X1 U8643 ( .A1(n9423), .A2(n12235), .ZN(n13016) );
  NAND2_X1 U8644 ( .A1(n12964), .A2(n12911), .ZN(n13012) );
  NAND2_X1 U8645 ( .A1(n7576), .A2(n7575), .ZN(n13205) );
  NAND4_X1 U8646 ( .A1(n7661), .A2(n7660), .A3(n7659), .A4(n7658), .ZN(n13048)
         );
  OR2_X1 U8647 ( .A1(n8157), .A2(n7657), .ZN(n7658) );
  NAND2_X1 U8648 ( .A1(n7605), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n7611) );
  OR2_X1 U8649 ( .A1(n14708), .A2(n14707), .ZN(n14709) );
  AND2_X1 U8650 ( .A1(n9278), .A2(n13484), .ZN(n14759) );
  OR2_X1 U8651 ( .A1(n11907), .A2(n7592), .ZN(n8187) );
  INV_X1 U8652 ( .A(n8164), .ZN(n8165) );
  AOI21_X1 U8653 ( .B1(n13025), .B2(n14334), .A(n7442), .ZN(n8164) );
  CLKBUF_X1 U8654 ( .A(n11921), .Z(n13167) );
  NAND2_X1 U8655 ( .A1(n7084), .A2(n7085), .ZN(n13195) );
  AOI21_X1 U8656 ( .B1(n13225), .B2(n6549), .A(n7058), .ZN(n13197) );
  INV_X1 U8657 ( .A(n13375), .ZN(n13220) );
  NAND2_X1 U8658 ( .A1(n7087), .A2(n7089), .ZN(n13210) );
  NAND2_X1 U8659 ( .A1(n7088), .A2(n7060), .ZN(n7087) );
  NAND2_X1 U8660 ( .A1(n13253), .A2(n7961), .ZN(n13238) );
  AND2_X1 U8661 ( .A1(n13258), .A2(n13257), .ZN(n13389) );
  NAND2_X1 U8662 ( .A1(n13322), .A2(n7894), .ZN(n13301) );
  CLKBUF_X1 U8663 ( .A(n11412), .Z(n13425) );
  NAND2_X1 U8664 ( .A1(n7049), .A2(n7048), .ZN(n11348) );
  AND2_X1 U8665 ( .A1(n7049), .A2(n6606), .ZN(n11349) );
  NAND2_X1 U8666 ( .A1(n7077), .A2(n7075), .ZN(n10768) );
  NAND2_X1 U8667 ( .A1(n8121), .A2(n8120), .ZN(n10644) );
  NAND2_X1 U8668 ( .A1(n10484), .A2(n7749), .ZN(n10414) );
  NAND2_X1 U8669 ( .A1(n7068), .A2(n8116), .ZN(n10480) );
  INV_X1 U8670 ( .A(n14362), .ZN(n13330) );
  NAND2_X1 U8671 ( .A1(n7099), .A2(n7712), .ZN(n10467) );
  NAND2_X1 U8672 ( .A1(n7072), .A2(n8111), .ZN(n10139) );
  NAND2_X1 U8673 ( .A1(n9565), .A2(n7662), .ZN(n10167) );
  NAND2_X1 U8674 ( .A1(n13281), .A2(n9413), .ZN(n13311) );
  AOI22_X1 U8675 ( .A1(n7908), .A2(P1_DATAO_REG_3__SCAN_IN), .B1(n7907), .B2(
        n13081), .ZN(n7638) );
  INV_X1 U8676 ( .A(n14829), .ZN(n14827) );
  NAND2_X1 U8677 ( .A1(n13362), .A2(n13361), .ZN(n13438) );
  NOR2_X1 U8678 ( .A1(n13360), .A2(n13359), .ZN(n13361) );
  OR2_X1 U8679 ( .A1(n13355), .A2(n14791), .ZN(n13362) );
  OR2_X1 U8680 ( .A1(n13358), .A2(n13357), .ZN(n13359) );
  INV_X1 U8681 ( .A(n13187), .ZN(n13442) );
  OR3_X1 U8682 ( .A1(n13417), .A2(n13416), .A3(n13415), .ZN(n13464) );
  NAND2_X1 U8683 ( .A1(n7464), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7465) );
  INV_X1 U8684 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n15170) );
  INV_X1 U8685 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n11013) );
  NOR2_X1 U8686 ( .A1(n8054), .A2(n7438), .ZN(n8055) );
  INV_X1 U8687 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n10497) );
  INV_X1 U8688 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n9961) );
  INV_X1 U8689 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n15181) );
  INV_X1 U8690 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n15325) );
  INV_X1 U8691 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n15367) );
  INV_X1 U8692 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n15272) );
  INV_X1 U8693 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n9173) );
  INV_X1 U8694 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n9096) );
  INV_X1 U8695 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n9068) );
  INV_X1 U8696 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n8987) );
  INV_X1 U8697 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n8967) );
  INV_X1 U8698 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n8963) );
  BUF_X1 U8699 ( .A(P2_IR_REG_0__SCAN_IN), .Z(n15206) );
  NAND2_X1 U8700 ( .A1(n6646), .A2(n10287), .ZN(n7210) );
  AOI21_X1 U8701 ( .B1(n7182), .B2(n7184), .A(n6611), .ZN(n7181) );
  OAI21_X1 U8702 ( .B1(n10606), .B2(n7205), .A(n7203), .ZN(n11023) );
  NAND2_X1 U8703 ( .A1(n8903), .A2(n8902), .ZN(n8935) );
  NAND2_X1 U8704 ( .A1(n7193), .A2(n6565), .ZN(n13629) );
  AND2_X1 U8705 ( .A1(n7200), .A2(n7199), .ZN(n7194) );
  NOR2_X1 U8706 ( .A1(n7279), .A2(n6964), .ZN(n7278) );
  AND2_X1 U8707 ( .A1(n9059), .A2(n6573), .ZN(n6964) );
  NAND2_X1 U8708 ( .A1(n9842), .A2(n9925), .ZN(n9938) );
  AOI21_X1 U8709 ( .B1(n13692), .B2(n13691), .A(n13690), .ZN(n13694) );
  NAND2_X1 U8710 ( .A1(n7218), .A2(n7221), .ZN(n13670) );
  NAND2_X1 U8711 ( .A1(n7220), .A2(n7219), .ZN(n7218) );
  INV_X1 U8712 ( .A(n13716), .ZN(n7220) );
  NAND2_X1 U8713 ( .A1(n10674), .A2(n10673), .ZN(n10828) );
  NAND2_X1 U8714 ( .A1(n13661), .A2(n11244), .ZN(n13499) );
  NAND2_X1 U8715 ( .A1(n7197), .A2(n7198), .ZN(n13725) );
  NAND2_X1 U8716 ( .A1(n7213), .A2(n7211), .ZN(n10286) );
  INV_X1 U8717 ( .A(n7212), .ZN(n7211) );
  NAND2_X1 U8718 ( .A1(n6704), .A2(n9842), .ZN(n7213) );
  NAND2_X1 U8719 ( .A1(n8940), .A2(P1_STATE_REG_SCAN_IN), .ZN(n14401) );
  XNOR2_X1 U8720 ( .A(n7172), .B(n13518), .ZN(n13746) );
  OR2_X1 U8721 ( .A1(n8941), .A2(n8932), .ZN(n13756) );
  NAND2_X1 U8722 ( .A1(n8843), .A2(n7161), .ZN(n6932) );
  OR2_X1 U8723 ( .A1(n8781), .A2(n8385), .ZN(n8387) );
  OR2_X1 U8724 ( .A1(n8781), .A2(n8371), .ZN(n8373) );
  OAI21_X1 U8725 ( .B1(n9217), .B2(n9212), .A(n9109), .ZN(n9215) );
  NOR2_X1 U8726 ( .A1(n9110), .A2(n9111), .ZN(n9143) );
  AND2_X1 U8727 ( .A1(n9488), .A2(n9487), .ZN(n9898) );
  NOR2_X1 U8728 ( .A1(n9901), .A2(n9900), .ZN(n10340) );
  NAND2_X1 U8729 ( .A1(n10691), .A2(n10690), .ZN(n11192) );
  OR2_X1 U8730 ( .A1(n11907), .A2(n8785), .ZN(n8787) );
  AND2_X1 U8731 ( .A1(n6980), .A2(n14546), .ZN(n6979) );
  NAND2_X1 U8732 ( .A1(n13962), .A2(n13909), .ZN(n13949) );
  NAND2_X1 U8733 ( .A1(n7424), .A2(n6623), .ZN(n14167) );
  INV_X1 U8734 ( .A(n13989), .ZN(n13906) );
  NAND2_X1 U8735 ( .A1(n7424), .A2(n13905), .ZN(n13990) );
  AOI211_X1 U8736 ( .C1(n14003), .C2(n14596), .A(n14000), .B(n13999), .ZN(
        n14178) );
  NAND2_X1 U8737 ( .A1(n14009), .A2(n13880), .ZN(n13997) );
  NAND2_X1 U8738 ( .A1(n14046), .A2(n13899), .ZN(n14035) );
  NAND2_X1 U8739 ( .A1(n7282), .A2(n13875), .ZN(n14024) );
  NAND2_X1 U8740 ( .A1(n14065), .A2(n13898), .ZN(n14048) );
  AND2_X1 U8741 ( .A1(n8656), .A2(n8655), .ZN(n14061) );
  AND2_X1 U8742 ( .A1(n6780), .A2(n13896), .ZN(n14064) );
  AOI21_X1 U8743 ( .B1(n13892), .B2(n7422), .A(n7421), .ZN(n14090) );
  NAND2_X1 U8744 ( .A1(n13892), .A2(n13891), .ZN(n14122) );
  AND2_X1 U8745 ( .A1(n7283), .A2(n6597), .ZN(n14105) );
  NAND2_X1 U8746 ( .A1(n11390), .A2(n11389), .ZN(n13866) );
  NAND2_X1 U8747 ( .A1(n11302), .A2(n11301), .ZN(n11304) );
  AND2_X1 U8748 ( .A1(n11211), .A2(n11210), .ZN(n7429) );
  NAND2_X1 U8749 ( .A1(n6782), .A2(n10871), .ZN(n10873) );
  NAND2_X1 U8750 ( .A1(n10807), .A2(n10806), .ZN(n10856) );
  NAND2_X1 U8751 ( .A1(n10813), .A2(n10812), .ZN(n10870) );
  NAND2_X1 U8752 ( .A1(n9222), .A2(n8417), .ZN(n8503) );
  NAND2_X1 U8753 ( .A1(n10317), .A2(n10316), .ZN(n14511) );
  INV_X1 U8754 ( .A(n14566), .ZN(n14119) );
  NAND2_X1 U8755 ( .A1(n8942), .A2(n9056), .ZN(n14542) );
  INV_X1 U8756 ( .A(n13959), .ZN(n14574) );
  NAND2_X1 U8757 ( .A1(n8335), .A2(n9654), .ZN(n9895) );
  OR2_X1 U8758 ( .A1(n8344), .A2(n14553), .ZN(n8335) );
  NAND2_X1 U8759 ( .A1(n8780), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n8363) );
  INV_X1 U8760 ( .A(n14147), .ZN(n14148) );
  AND2_X2 U8761 ( .A1(n9359), .A2(n9657), .ZN(n14645) );
  INV_X1 U8762 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n15297) );
  INV_X1 U8763 ( .A(n8924), .ZN(n11225) );
  NAND2_X1 U8764 ( .A1(n7244), .A2(n7557), .ZN(n7962) );
  NAND2_X1 U8765 ( .A1(n7555), .A2(n7949), .ZN(n7244) );
  OAI21_X1 U8766 ( .B1(n7160), .B2(n7158), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n8346) );
  NAND2_X1 U8767 ( .A1(n8342), .A2(n7159), .ZN(n7158) );
  OAI21_X1 U8768 ( .B1(n8620), .B2(n8338), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n8340) );
  INV_X1 U8769 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n15263) );
  INV_X1 U8770 ( .A(n8928), .ZN(n13847) );
  INV_X1 U8771 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n9915) );
  INV_X1 U8772 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n9785) );
  INV_X1 U8773 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n9398) );
  NAND2_X1 U8774 ( .A1(n6713), .A2(n7510), .ZN(n7734) );
  INV_X1 U8775 ( .A(n7733), .ZN(n6713) );
  INV_X1 U8776 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n9172) );
  INV_X1 U8777 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n9094) );
  INV_X1 U8778 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n9071) );
  INV_X1 U8779 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n9066) );
  INV_X1 U8780 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n8991) );
  INV_X1 U8781 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n8988) );
  XNOR2_X1 U8782 ( .A(n8256), .B(n6861), .ZN(n15419) );
  INV_X1 U8783 ( .A(n8255), .ZN(n6861) );
  XNOR2_X1 U8784 ( .A(n8260), .B(n6728), .ZN(n15412) );
  NAND2_X1 U8785 ( .A1(n15412), .A2(n15411), .ZN(n15410) );
  XNOR2_X1 U8786 ( .A(n8265), .B(n8264), .ZN(n14284) );
  NOR2_X1 U8787 ( .A1(n8270), .A2(n15414), .ZN(n14288) );
  NAND2_X1 U8788 ( .A1(n14288), .A2(n14287), .ZN(n14286) );
  NOR2_X1 U8789 ( .A1(n8276), .A2(n8275), .ZN(n14295) );
  NAND2_X1 U8790 ( .A1(n14296), .A2(n14294), .ZN(n14422) );
  NAND2_X1 U8791 ( .A1(n14422), .A2(n14421), .ZN(n14420) );
  NAND2_X1 U8792 ( .A1(n14430), .A2(n6716), .ZN(n14435) );
  NAND2_X1 U8793 ( .A1(n6718), .A2(n6717), .ZN(n6716) );
  INV_X1 U8794 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n6717) );
  NAND2_X1 U8795 ( .A1(n6857), .A2(n6856), .ZN(n6718) );
  AOI211_X1 U8796 ( .C1(n11858), .C2(n11857), .A(n11856), .B(n11855), .ZN(
        n11865) );
  AOI21_X1 U8797 ( .B1(n6896), .B2(n14973), .A(n6893), .ZN(n12504) );
  OAI211_X1 U8798 ( .C1(n6545), .C2(n12485), .A(n7015), .B(n7014), .ZN(n12505)
         );
  XNOR2_X1 U8799 ( .A(n6898), .B(n6897), .ZN(n6896) );
  NAND2_X1 U8800 ( .A1(n7113), .A2(n9829), .ZN(n10068) );
  NAND2_X1 U8801 ( .A1(n9552), .A2(n9551), .ZN(n9575) );
  AND3_X1 U8802 ( .A1(n12234), .A2(n12233), .A3(n12232), .ZN(n12240) );
  OAI21_X1 U8803 ( .B1(n6806), .B2(n13468), .A(n8205), .ZN(n8206) );
  INV_X1 U8804 ( .A(n6730), .ZN(n6729) );
  OAI21_X1 U8805 ( .B1(n14151), .B2(n13743), .A(n13616), .ZN(n6730) );
  NAND2_X1 U8806 ( .A1(n14237), .A2(n14645), .ZN(n6975) );
  INV_X1 U8807 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n6974) );
  INV_X1 U8808 ( .A(n14280), .ZN(n14279) );
  INV_X1 U8809 ( .A(n14292), .ZN(n14291) );
  NAND2_X1 U8810 ( .A1(n14424), .A2(n8279), .ZN(n14428) );
  AND2_X1 U8811 ( .A1(n14424), .A2(n6690), .ZN(n14426) );
  NOR2_X1 U8812 ( .A1(n14274), .A2(n6849), .ZN(n14275) );
  NOR2_X1 U8813 ( .A1(n6850), .A2(n6552), .ZN(n6849) );
  INV_X1 U8814 ( .A(n6755), .ZN(n14274) );
  XNOR2_X1 U8815 ( .A(n6753), .B(n6601), .ZN(SUB_1596_U4) );
  NAND2_X1 U8816 ( .A1(n6755), .A2(n6754), .ZN(n6753) );
  INV_X1 U8817 ( .A(n12090), .ZN(n12149) );
  AND2_X1 U8818 ( .A1(n6551), .A2(n6582), .ZN(n6542) );
  XNOR2_X1 U8819 ( .A(n13956), .B(n13910), .ZN(n13948) );
  AND2_X1 U8820 ( .A1(n6653), .A2(n6566), .ZN(n6543) );
  AND2_X1 U8821 ( .A1(n14143), .A2(n13886), .ZN(n6544) );
  AND2_X1 U8822 ( .A1(n7017), .A2(n12482), .ZN(n6545) );
  AND2_X1 U8823 ( .A1(n13619), .A2(n7227), .ZN(n6546) );
  AND2_X1 U8824 ( .A1(n6779), .A2(n13899), .ZN(n6547) );
  INV_X1 U8825 ( .A(n9841), .ZN(n7178) );
  AND2_X1 U8826 ( .A1(n14615), .A2(n9854), .ZN(n6548) );
  AND2_X1 U8827 ( .A1(n8149), .A2(n13224), .ZN(n6549) );
  AND2_X1 U8828 ( .A1(n8979), .A2(n8977), .ZN(n8984) );
  AND2_X1 U8829 ( .A1(n8168), .A2(n6798), .ZN(n6550) );
  OR2_X1 U8830 ( .A1(n11886), .A2(n12551), .ZN(n6551) );
  XOR2_X1 U8831 ( .A(n8300), .B(n8299), .Z(n6552) );
  AND2_X1 U8832 ( .A1(n7357), .A2(n7356), .ZN(n6553) );
  OR3_X1 U8833 ( .A1(n11327), .A2(n11326), .A3(n11325), .ZN(n12691) );
  AND3_X1 U8834 ( .A1(n7454), .A2(n7453), .A3(n6602), .ZN(n6555) );
  AND2_X1 U8835 ( .A1(n6550), .A2(n6797), .ZN(n6556) );
  AND2_X1 U8836 ( .A1(n12085), .A2(n12084), .ZN(n6557) );
  AND2_X1 U8837 ( .A1(n8746), .A2(n6917), .ZN(n6558) );
  AND2_X1 U8838 ( .A1(n6998), .A2(n6695), .ZN(n6559) );
  AND2_X1 U8839 ( .A1(n8632), .A2(n8604), .ZN(n6560) );
  AND2_X1 U8840 ( .A1(n6652), .A2(n6834), .ZN(n6561) );
  AND2_X1 U8841 ( .A1(n11924), .A2(n8153), .ZN(n6562) );
  INV_X1 U8842 ( .A(n12065), .ZN(n13469) );
  AND2_X1 U8843 ( .A1(n6640), .A2(n9862), .ZN(n6563) );
  INV_X1 U8844 ( .A(n8773), .ZN(n7152) );
  AND2_X1 U8845 ( .A1(n6747), .A2(n6746), .ZN(n6564) );
  INV_X1 U8846 ( .A(P3_IR_REG_28__SCAN_IN), .ZN(n9719) );
  OR2_X1 U8847 ( .A1(n7195), .A2(n7449), .ZN(n6565) );
  OR2_X1 U8848 ( .A1(n12087), .A2(n6557), .ZN(n6566) );
  AND2_X1 U8849 ( .A1(n9377), .A2(n9376), .ZN(n6567) );
  INV_X1 U8850 ( .A(n13963), .ZN(n6740) );
  AND2_X1 U8851 ( .A1(n6983), .A2(n6982), .ZN(n6569) );
  NAND2_X1 U8852 ( .A1(n6868), .A2(n6948), .ZN(n6570) );
  INV_X1 U8853 ( .A(n6787), .ZN(n6786) );
  NAND2_X1 U8854 ( .A1(n11221), .A2(n11210), .ZN(n6787) );
  OR2_X1 U8855 ( .A1(n11917), .A2(n12520), .ZN(n11809) );
  AND2_X1 U8856 ( .A1(n11375), .A2(n11374), .ZN(n6571) );
  AND2_X1 U8857 ( .A1(P1_DATAO_REG_7__SCAN_IN), .A2(n7353), .ZN(n6572) );
  INV_X1 U8858 ( .A(n8532), .ZN(n7165) );
  INV_X1 U8859 ( .A(n8670), .ZN(n7157) );
  AND2_X1 U8860 ( .A1(n9727), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n6573) );
  NOR2_X1 U8861 ( .A1(n12813), .A2(n12313), .ZN(n6949) );
  AND2_X1 U8862 ( .A1(n8843), .A2(n6660), .ZN(n6574) );
  INV_X1 U8863 ( .A(n8440), .ZN(n7163) );
  INV_X1 U8864 ( .A(n11464), .ZN(n7131) );
  AND2_X1 U8865 ( .A1(n13308), .A2(n6556), .ZN(n6575) );
  OR2_X1 U8866 ( .A1(n11120), .A2(n11121), .ZN(n6576) );
  AND3_X1 U8867 ( .A1(n6687), .A2(n6554), .A3(n6942), .ZN(n9194) );
  NOR2_X1 U8868 ( .A1(n10989), .A2(n12032), .ZN(n10990) );
  INV_X1 U8869 ( .A(n7381), .ZN(n9082) );
  INV_X1 U8870 ( .A(n11132), .ZN(n6890) );
  INV_X1 U8871 ( .A(n6817), .ZN(n6814) );
  NAND2_X1 U8872 ( .A1(n6701), .A2(n7738), .ZN(n6577) );
  NAND2_X1 U8873 ( .A1(n8552), .A2(n8551), .ZN(n14405) );
  INV_X1 U8874 ( .A(n14405), .ZN(n6969) );
  NAND2_X1 U8875 ( .A1(n8561), .A2(n7439), .ZN(n8844) );
  INV_X1 U8876 ( .A(n11980), .ZN(n6795) );
  AND2_X1 U8877 ( .A1(n7738), .A2(n7737), .ZN(n8049) );
  AND2_X1 U8878 ( .A1(n7526), .A2(n7732), .ZN(n6578) );
  INV_X1 U8879 ( .A(n13224), .ZN(n7060) );
  AND2_X1 U8880 ( .A1(n7365), .A2(n9074), .ZN(n6579) );
  NAND4_X1 U8881 ( .A1(n7601), .A2(n7600), .A3(n7599), .A4(n7598), .ZN(n11928)
         );
  NOR2_X1 U8882 ( .A1(n12564), .A2(n12565), .ZN(n12563) );
  NAND2_X1 U8883 ( .A1(n6942), .A2(n8860), .ZN(n8956) );
  NOR2_X1 U8884 ( .A1(n12764), .A2(n12665), .ZN(n6580) );
  NAND2_X1 U8885 ( .A1(n8635), .A2(n8634), .ZN(n14203) );
  OR2_X1 U8886 ( .A1(n10782), .A2(n13040), .ZN(n6581) );
  NAND2_X1 U8887 ( .A1(n11889), .A2(n12331), .ZN(n6582) );
  NOR2_X1 U8888 ( .A1(n6523), .A2(n8132), .ZN(n6583) );
  AND2_X1 U8889 ( .A1(n12016), .A2(n12015), .ZN(n6584) );
  AND2_X1 U8890 ( .A1(n6619), .A2(n7305), .ZN(n6585) );
  INV_X1 U8891 ( .A(P3_ADDR_REG_4__SCAN_IN), .ZN(n15262) );
  OR2_X1 U8892 ( .A1(n8212), .A2(n8211), .ZN(n6586) );
  AND2_X1 U8893 ( .A1(n9173), .A2(P2_DATAO_REG_9__SCAN_IN), .ZN(n6587) );
  OR2_X1 U8894 ( .A1(n14218), .A2(n14088), .ZN(n6588) );
  INV_X1 U8895 ( .A(n10858), .ZN(n10874) );
  AND2_X1 U8896 ( .A1(n9839), .A2(n9838), .ZN(n6589) );
  AND2_X1 U8897 ( .A1(n8973), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n6590) );
  AOI21_X1 U8898 ( .B1(n8795), .B2(n8417), .A(n8797), .ZN(n14128) );
  AND2_X1 U8899 ( .A1(n14042), .A2(n6569), .ZN(n6591) );
  AND4_X1 U8900 ( .A1(n8318), .A2(n8847), .A3(n8317), .A4(n8316), .ZN(n6592)
         );
  AND4_X1 U8901 ( .A1(n8315), .A2(n8314), .A3(n8313), .A4(n8312), .ZN(n6593)
         );
  AND2_X1 U8902 ( .A1(n13233), .A2(n8146), .ZN(n6594) );
  NAND2_X1 U8903 ( .A1(n10066), .A2(n10065), .ZN(n6595) );
  AND2_X1 U8904 ( .A1(n12758), .A2(n12603), .ZN(n6596) );
  NAND2_X1 U8905 ( .A1(n13890), .A2(n13864), .ZN(n6597) );
  AND2_X1 U8906 ( .A1(n12080), .A2(n12079), .ZN(n6598) );
  NAND2_X1 U8907 ( .A1(n9937), .A2(n9936), .ZN(n6599) );
  NAND2_X1 U8908 ( .A1(n12888), .A2(n12889), .ZN(n6600) );
  INV_X1 U8909 ( .A(n11613), .ZN(n11681) );
  NAND2_X1 U8910 ( .A1(n6773), .A2(n13904), .ZN(n13994) );
  XOR2_X1 U8911 ( .A(n8304), .B(n8298), .Z(n6601) );
  INV_X1 U8912 ( .A(n12174), .ZN(n6806) );
  NAND2_X1 U8913 ( .A1(n7231), .A2(n8194), .ZN(n12174) );
  INV_X1 U8914 ( .A(n13941), .ZN(n7294) );
  NAND2_X1 U8915 ( .A1(n12876), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9380) );
  AOI21_X1 U8916 ( .B1(n13716), .B2(n13715), .A(n13714), .ZN(n13618) );
  AND4_X1 U8917 ( .A1(n7455), .A2(n8051), .A3(n8050), .A4(n8064), .ZN(n6602)
         );
  AND2_X1 U8918 ( .A1(n14136), .A2(n14607), .ZN(n6603) );
  AND2_X1 U8919 ( .A1(n14034), .A2(n7412), .ZN(n6604) );
  AND2_X1 U8920 ( .A1(n8644), .A2(n13869), .ZN(n14070) );
  NAND2_X1 U8921 ( .A1(n7458), .A2(n7614), .ZN(n7717) );
  AND3_X1 U8922 ( .A1(n8862), .A2(n8861), .A3(n8982), .ZN(n9033) );
  OR2_X1 U8923 ( .A1(n14176), .A2(n13881), .ZN(n6605) );
  NAND2_X1 U8924 ( .A1(n14356), .A2(n8124), .ZN(n6606) );
  OR2_X1 U8925 ( .A1(n7918), .A2(n7103), .ZN(n6607) );
  AND3_X1 U8926 ( .A1(n11790), .A2(n12587), .A3(n11789), .ZN(n6608) );
  OR2_X1 U8927 ( .A1(n6827), .A2(n6585), .ZN(n6609) );
  OR2_X1 U8928 ( .A1(n12568), .A2(n12578), .ZN(n6610) );
  INV_X1 U8929 ( .A(n13611), .ZN(n7192) );
  AND2_X1 U8930 ( .A1(n13502), .A2(n13501), .ZN(n6611) );
  OR2_X1 U8931 ( .A1(n12054), .A2(n12053), .ZN(n6612) );
  AND2_X1 U8932 ( .A1(n11987), .A2(n11986), .ZN(n6613) );
  AND2_X1 U8933 ( .A1(n11869), .A2(n12341), .ZN(n6614) );
  AND2_X1 U8934 ( .A1(n12089), .A2(n12088), .ZN(n6615) );
  INV_X1 U8935 ( .A(n13893), .ZN(n7421) );
  AND2_X1 U8936 ( .A1(n11972), .A2(n11971), .ZN(n6616) );
  INV_X1 U8937 ( .A(n7206), .ZN(n7205) );
  NOR2_X1 U8938 ( .A1(n10827), .A2(n7207), .ZN(n7206) );
  NAND2_X1 U8939 ( .A1(n8022), .A2(n8021), .ZN(n13356) );
  INV_X1 U8940 ( .A(n12062), .ZN(n6835) );
  NAND2_X1 U8941 ( .A1(n8187), .A2(n8186), .ZN(n13159) );
  AND2_X1 U8942 ( .A1(n14811), .A2(n13041), .ZN(n6617) );
  NAND2_X1 U8943 ( .A1(n11018), .A2(n10857), .ZN(n6618) );
  NOR2_X1 U8944 ( .A1(n8980), .A2(n7350), .ZN(n7349) );
  AND2_X1 U8945 ( .A1(n12020), .A2(n12019), .ZN(n6619) );
  AND2_X1 U8946 ( .A1(n11890), .A2(n12283), .ZN(n6620) );
  AND2_X1 U8947 ( .A1(n12964), .A2(n7148), .ZN(n6621) );
  AND2_X1 U8948 ( .A1(n7017), .A2(n7013), .ZN(n6622) );
  INV_X1 U8949 ( .A(n7223), .ZN(n7219) );
  NAND2_X1 U8950 ( .A1(n6546), .A2(n7230), .ZN(n7223) );
  AND2_X1 U8951 ( .A1(n13906), .A2(n13905), .ZN(n6623) );
  OR2_X1 U8952 ( .A1(n14556), .A2(n6539), .ZN(n6624) );
  INV_X1 U8953 ( .A(n7229), .ZN(n7228) );
  OR2_X1 U8954 ( .A1(n13620), .A2(n13562), .ZN(n7229) );
  AND2_X1 U8955 ( .A1(n7035), .A2(n7034), .ZN(n6625) );
  OR2_X1 U8956 ( .A1(n12028), .A2(n12029), .ZN(n6626) );
  AND2_X1 U8957 ( .A1(n14615), .A2(n13769), .ZN(n6627) );
  AND2_X1 U8958 ( .A1(n12210), .A2(n6606), .ZN(n7048) );
  OR2_X1 U8959 ( .A1(n14190), .A2(n14025), .ZN(n13899) );
  AND2_X1 U8960 ( .A1(n12540), .A2(n12801), .ZN(n6962) );
  OR2_X1 U8961 ( .A1(n12890), .A2(n12891), .ZN(n6747) );
  NOR2_X1 U8962 ( .A1(n11980), .A2(n13047), .ZN(n6628) );
  INV_X1 U8963 ( .A(n12646), .ZN(n12650) );
  AND2_X1 U8964 ( .A1(n11769), .A2(n11777), .ZN(n12646) );
  AND2_X1 U8965 ( .A1(n11022), .A2(n7206), .ZN(n6629) );
  NOR2_X1 U8966 ( .A1(n13375), .A2(n13028), .ZN(n6630) );
  OR2_X1 U8967 ( .A1(n6992), .A2(n6991), .ZN(n6631) );
  OR2_X1 U8968 ( .A1(n11984), .A2(n11983), .ZN(n6632) );
  NOR2_X1 U8969 ( .A1(n12050), .A2(n8126), .ZN(n6633) );
  NOR2_X1 U8970 ( .A1(n14379), .A2(n8122), .ZN(n6634) );
  INV_X1 U8971 ( .A(n7090), .ZN(n7089) );
  NOR2_X1 U8972 ( .A1(n13451), .A2(n8146), .ZN(n7090) );
  INV_X1 U8973 ( .A(n8844), .ZN(n6791) );
  NAND2_X1 U8974 ( .A1(n13446), .A2(n8150), .ZN(n6635) );
  OR2_X1 U8975 ( .A1(n8824), .A2(n6739), .ZN(n6636) );
  AOI21_X1 U8976 ( .B1(n8745), .B2(n6914), .A(n6912), .ZN(n6911) );
  INV_X1 U8977 ( .A(n12714), .ZN(n14308) );
  NOR2_X1 U8978 ( .A1(n11313), .A2(n12719), .ZN(n6637) );
  NAND2_X1 U8979 ( .A1(n11021), .A2(n11020), .ZN(n6638) );
  INV_X1 U8980 ( .A(n7449), .ZN(n7200) );
  INV_X1 U8981 ( .A(n6809), .ZN(n6808) );
  NAND2_X1 U8982 ( .A1(n6811), .A2(n6810), .ZN(n6809) );
  AND2_X1 U8983 ( .A1(n12170), .A2(n12169), .ZN(n6639) );
  OR2_X1 U8984 ( .A1(n14615), .A2(n13769), .ZN(n6640) );
  AND2_X1 U8985 ( .A1(n7427), .A2(n6785), .ZN(n6641) );
  AND2_X1 U8986 ( .A1(n10826), .A2(n10825), .ZN(n6642) );
  AND2_X1 U8987 ( .A1(n7320), .A2(n6615), .ZN(n6643) );
  NOR2_X1 U8988 ( .A1(n12914), .A2(n12913), .ZN(n6644) );
  NAND2_X1 U8989 ( .A1(n12786), .A2(n11667), .ZN(n6645) );
  OR2_X1 U8990 ( .A1(n10285), .A2(n7212), .ZN(n6646) );
  INV_X1 U8991 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n15304) );
  OR2_X1 U8992 ( .A1(n6871), .A2(n6869), .ZN(n6868) );
  OR2_X1 U8993 ( .A1(n9028), .A2(n9027), .ZN(n14875) );
  INV_X1 U8994 ( .A(n14875), .ZN(n7024) );
  AND2_X1 U8995 ( .A1(n7010), .A2(n6582), .ZN(n6647) );
  NAND2_X1 U8996 ( .A1(n12516), .A2(n12517), .ZN(n6648) );
  INV_X1 U8997 ( .A(n12565), .ZN(n6872) );
  NAND2_X1 U8998 ( .A1(n11674), .A2(n11675), .ZN(n12565) );
  AND2_X1 U8999 ( .A1(n7323), .A2(n7322), .ZN(n6649) );
  AND2_X1 U9000 ( .A1(n12565), .A2(n6949), .ZN(n6650) );
  INV_X1 U9001 ( .A(n8984), .ZN(n8978) );
  OR2_X1 U9002 ( .A1(n7310), .A2(n7309), .ZN(n6651) );
  NAND2_X1 U9003 ( .A1(n12067), .A2(n12066), .ZN(n6652) );
  OR2_X1 U9004 ( .A1(n7320), .A2(n6615), .ZN(n6653) );
  INV_X1 U9005 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n9085) );
  INV_X1 U9006 ( .A(n8724), .ZN(n6937) );
  AND3_X1 U9007 ( .A1(n10005), .A2(n10004), .A3(n10003), .ZN(n10369) );
  NOR2_X1 U9008 ( .A1(n12563), .A2(n11678), .ZN(n6654) );
  OR2_X1 U9009 ( .A1(n14143), .A2(n13886), .ZN(n6655) );
  OR2_X1 U9010 ( .A1(n12640), .A2(n6580), .ZN(n6656) );
  OR2_X1 U9011 ( .A1(n6580), .A2(n12642), .ZN(n6657) );
  OR2_X1 U9012 ( .A1(n7024), .A2(n10890), .ZN(n6658) );
  OR2_X1 U9013 ( .A1(n8214), .A2(n8213), .ZN(n6659) );
  OR2_X1 U9014 ( .A1(n8807), .A2(n8830), .ZN(n6660) );
  AND2_X1 U9015 ( .A1(n7085), .A2(n6635), .ZN(n6661) );
  AND2_X1 U9016 ( .A1(n6803), .A2(n12174), .ZN(n6662) );
  AND2_X1 U9017 ( .A1(n14121), .A2(n6597), .ZN(n6663) );
  AND2_X1 U9018 ( .A1(n14807), .A2(n6815), .ZN(n6664) );
  AND2_X1 U9019 ( .A1(n7460), .A2(n7573), .ZN(n6665) );
  AND2_X1 U9020 ( .A1(n12198), .A2(n8111), .ZN(n6666) );
  NOR2_X1 U9021 ( .A1(n13998), .A2(n7301), .ZN(n6667) );
  NAND2_X1 U9022 ( .A1(n7951), .A2(n7950), .ZN(n13263) );
  AND2_X1 U9023 ( .A1(n7012), .A2(n9374), .ZN(n6668) );
  NAND2_X1 U9024 ( .A1(n13941), .A2(n8811), .ZN(n13963) );
  NAND2_X1 U9025 ( .A1(n9578), .A2(n9577), .ZN(n6669) );
  AND2_X1 U9026 ( .A1(n7870), .A2(n7850), .ZN(n6670) );
  AND2_X1 U9027 ( .A1(n13559), .A2(n13558), .ZN(n13562) );
  NOR2_X1 U9028 ( .A1(n8001), .A2(n7090), .ZN(n7086) );
  AND2_X1 U9029 ( .A1(n12073), .A2(n12072), .ZN(n6671) );
  AND2_X1 U9030 ( .A1(n10858), .A2(n10871), .ZN(n6672) );
  NAND2_X1 U9031 ( .A1(n8722), .A2(n8721), .ZN(n14168) );
  AND2_X1 U9032 ( .A1(n10374), .A2(n10373), .ZN(n6673) );
  OR2_X1 U9033 ( .A1(n12794), .A2(n12250), .ZN(n11814) );
  OR2_X1 U9034 ( .A1(n7163), .A2(n8441), .ZN(n6674) );
  AND2_X1 U9035 ( .A1(n7453), .A2(n7454), .ZN(n7061) );
  AND2_X1 U9036 ( .A1(n6592), .A2(n8333), .ZN(n6675) );
  AND2_X1 U9037 ( .A1(n8787), .A2(n8786), .ZN(n14134) );
  AND2_X1 U9038 ( .A1(n7526), .A2(n7271), .ZN(n6676) );
  NAND2_X1 U9039 ( .A1(n8533), .A2(n7165), .ZN(n6677) );
  NAND2_X1 U9040 ( .A1(n8671), .A2(n7157), .ZN(n6678) );
  AND2_X1 U9041 ( .A1(n7239), .A2(n7238), .ZN(n6679) );
  AND2_X1 U9042 ( .A1(n8471), .A2(n7164), .ZN(n6680) );
  AND2_X1 U9043 ( .A1(n7221), .A2(n13588), .ZN(n7217) );
  INV_X1 U9044 ( .A(P3_IR_REG_16__SCAN_IN), .ZN(n8866) );
  INV_X1 U9045 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n7159) );
  OR2_X1 U9046 ( .A1(n7192), .A2(n7190), .ZN(n6681) );
  NAND2_X1 U9047 ( .A1(n9094), .A2(P1_DATAO_REG_8__SCAN_IN), .ZN(n6682) );
  NAND2_X1 U9048 ( .A1(n8565), .A2(n8564), .ZN(n13754) );
  INV_X1 U9049 ( .A(n13754), .ZN(n6967) );
  NAND2_X1 U9050 ( .A1(n8706), .A2(n8705), .ZN(n14176) );
  INV_X1 U9051 ( .A(n14176), .ZN(n6982) );
  NAND2_X1 U9052 ( .A1(n6947), .A2(n6554), .ZN(n9196) );
  NAND2_X1 U9053 ( .A1(n6780), .A2(n6779), .ZN(n14065) );
  AND2_X1 U9054 ( .A1(n7137), .A2(n7139), .ZN(n6683) );
  INV_X1 U9055 ( .A(P3_IR_REG_9__SCAN_IN), .ZN(n6985) );
  NOR2_X1 U9056 ( .A1(n7859), .A2(P2_IR_REG_16__SCAN_IN), .ZN(n7878) );
  NAND2_X1 U9057 ( .A1(n7100), .A2(n7850), .ZN(n11413) );
  NAND2_X1 U9058 ( .A1(n7390), .A2(n11775), .ZN(n12649) );
  NOR2_X1 U9059 ( .A1(n12373), .A2(n12374), .ZN(n6684) );
  AND2_X1 U9060 ( .A1(n11268), .A2(n11265), .ZN(n6685) );
  NAND2_X1 U9061 ( .A1(n10990), .A2(n6808), .ZN(n6812) );
  AND2_X1 U9062 ( .A1(n7197), .A2(n7195), .ZN(n6686) );
  AND3_X1 U9063 ( .A1(n6984), .A2(n8862), .A3(n8861), .ZN(n6687) );
  INV_X1 U9064 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n9515) );
  INV_X1 U9065 ( .A(n7260), .ZN(n7259) );
  NAND2_X1 U9066 ( .A1(n6689), .A2(n7534), .ZN(n7260) );
  OR2_X1 U9067 ( .A1(P1_ADDR_REG_6__SCAN_IN), .A2(n15271), .ZN(n6688) );
  OR2_X1 U9068 ( .A1(n7536), .A2(SI_17_), .ZN(n6689) );
  AND2_X1 U9069 ( .A1(n8279), .A2(n6855), .ZN(n6690) );
  AND2_X1 U9070 ( .A1(n7547), .A2(n7255), .ZN(n6691) );
  OR2_X1 U9071 ( .A1(n12634), .A2(n11496), .ZN(n6692) );
  AND2_X1 U9072 ( .A1(n7128), .A2(n6600), .ZN(n6693) );
  INV_X1 U9073 ( .A(n6949), .ZN(n6948) );
  INV_X1 U9074 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n7368) );
  NAND2_X1 U9075 ( .A1(n7380), .A2(n7379), .ZN(n11043) );
  XOR2_X1 U9076 ( .A(n7558), .B(SI_23_), .Z(n6694) );
  NAND2_X1 U9077 ( .A1(n7862), .A2(n7861), .ZN(n13426) );
  INV_X1 U9078 ( .A(n13426), .ZN(n6810) );
  NAND2_X1 U9079 ( .A1(n7391), .A2(n7395), .ZN(n14307) );
  INV_X1 U9080 ( .A(P3_IR_REG_15__SCAN_IN), .ZN(n6946) );
  NAND2_X1 U9081 ( .A1(n7937), .A2(n7936), .ZN(n13459) );
  INV_X1 U9082 ( .A(n13459), .ZN(n6797) );
  NAND2_X1 U9083 ( .A1(n8546), .A2(n8545), .ZN(n11253) );
  INV_X1 U9084 ( .A(n11253), .ZN(n6971) );
  OR2_X1 U9085 ( .A1(n11318), .A2(n12703), .ZN(n6695) );
  OR2_X1 U9086 ( .A1(n15057), .A2(P3_REG2_REG_29__SCAN_IN), .ZN(n6696) );
  NAND2_X1 U9087 ( .A1(n6972), .A2(n6971), .ZN(n11213) );
  INV_X1 U9088 ( .A(n11213), .ZN(n6970) );
  INV_X1 U9089 ( .A(n6972), .ZN(n11156) );
  OR2_X1 U9090 ( .A1(n10960), .A2(n10958), .ZN(n6697) );
  AND2_X1 U9091 ( .A1(n10255), .A2(n6866), .ZN(n6698) );
  AND2_X1 U9092 ( .A1(n10254), .A2(n6698), .ZN(n6699) );
  NAND2_X1 U9093 ( .A1(n7380), .A2(n7378), .ZN(n6700) );
  AND2_X1 U9094 ( .A1(n7065), .A2(n7061), .ZN(n6701) );
  NAND2_X1 U9095 ( .A1(n9499), .A2(n7012), .ZN(n6702) );
  OR2_X1 U9096 ( .A1(n8013), .A2(n7267), .ZN(n6703) );
  AND2_X1 U9097 ( .A1(n9925), .A2(n6599), .ZN(n6704) );
  NOR2_X1 U9098 ( .A1(n8003), .A2(n11550), .ZN(n6705) );
  INV_X1 U9099 ( .A(n10315), .ZN(n6966) );
  AND2_X1 U9100 ( .A1(n9567), .A2(n10130), .ZN(n6706) );
  AND2_X1 U9101 ( .A1(n7019), .A2(P3_REG2_REG_17__SCAN_IN), .ZN(n6707) );
  OR2_X1 U9102 ( .A1(n12453), .A2(n12770), .ZN(n6708) );
  NAND4_X1 U9103 ( .A1(n9717), .A2(n9716), .A3(n9715), .A4(n9714), .ZN(n15040)
         );
  INV_X1 U9104 ( .A(n15040), .ZN(n6723) );
  OR2_X1 U9105 ( .A1(n12453), .A2(n12683), .ZN(n6709) );
  INV_X1 U9106 ( .A(n12361), .ZN(n6724) );
  AND2_X1 U9107 ( .A1(n6707), .A2(n12491), .ZN(n6710) );
  INV_X1 U9108 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n11228) );
  OR2_X1 U9109 ( .A1(n9698), .A2(n9697), .ZN(n6711) );
  INV_X1 U9110 ( .A(n12465), .ZN(n6892) );
  INV_X1 U9111 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n7040) );
  OR2_X1 U9112 ( .A1(n12494), .A2(n12765), .ZN(n6712) );
  INV_X1 U9113 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n7353) );
  INV_X1 U9114 ( .A(P3_ADDR_REG_1__SCAN_IN), .ZN(n6760) );
  NAND2_X1 U9115 ( .A1(n7485), .A2(n7484), .ZN(n7487) );
  NAND2_X1 U9116 ( .A1(n7682), .A2(n7502), .ZN(n7700) );
  AOI21_X1 U9117 ( .B1(n13027), .B2(n13205), .A(n8002), .ZN(n13179) );
  OAI21_X1 U9118 ( .B1(n10485), .B2(n7096), .A(n7763), .ZN(n7095) );
  NAND2_X2 U9119 ( .A1(n6714), .A2(n7740), .ZN(n12008) );
  NAND2_X1 U9120 ( .A1(n7482), .A2(n7583), .ZN(n7587) );
  NAND2_X1 U9121 ( .A1(n7300), .A2(n7299), .ZN(n13976) );
  NAND2_X1 U9122 ( .A1(n14053), .A2(n13873), .ZN(n14039) );
  NAND2_X1 U9123 ( .A1(n11390), .A2(n7284), .ZN(n7283) );
  OAI21_X2 U9124 ( .B1(n11297), .B2(n11296), .A(n11295), .ZN(n11388) );
  AOI21_X2 U9125 ( .B1(n14087), .B2(n14091), .A(n13868), .ZN(n14069) );
  INV_X1 U9126 ( .A(n7277), .ZN(n10859) );
  INV_X1 U9127 ( .A(n14240), .ZN(n14239) );
  NAND2_X1 U9128 ( .A1(n13878), .A2(n13877), .ZN(n14010) );
  OAI21_X1 U9129 ( .B1(n7276), .B2(n10504), .A(n6618), .ZN(n7275) );
  OR2_X1 U9130 ( .A1(n12098), .A2(n12097), .ZN(n12110) );
  NOR2_X1 U9131 ( .A1(n6735), .A2(n6734), .ZN(n7126) );
  NOR2_X1 U9132 ( .A1(n12995), .A2(n12994), .ZN(n12993) );
  NAND2_X1 U9133 ( .A1(n12931), .A2(n6747), .ZN(n12987) );
  NAND2_X1 U9134 ( .A1(n6839), .A2(n6838), .ZN(n12096) );
  NAND2_X1 U9135 ( .A1(n12055), .A2(n6612), .ZN(n12061) );
  NAND2_X1 U9136 ( .A1(n6842), .A2(n12173), .ZN(n12178) );
  NAND2_X1 U9137 ( .A1(n6833), .A2(n6832), .ZN(n12074) );
  OAI21_X1 U9138 ( .B1(n6671), .B2(n7312), .A(n7311), .ZN(n12086) );
  AOI21_X1 U9139 ( .B1(n12145), .B2(n12144), .A(n6679), .ZN(n6843) );
  AOI21_X1 U9140 ( .B1(n12054), .B2(n12053), .A(n12051), .ZN(n12052) );
  AOI21_X1 U9141 ( .B1(n6831), .B2(n6829), .A(n6828), .ZN(n6827) );
  NAND2_X1 U9142 ( .A1(n10656), .A2(n6537), .ZN(n6715) );
  NAND2_X1 U9143 ( .A1(n7947), .A2(n7946), .ZN(n13251) );
  AOI22_X1 U9144 ( .A1(n13162), .A2(n13161), .B1(n13356), .B2(n13025), .ZN(
        n8048) );
  INV_X2 U9145 ( .A(n7625), .ZN(n7596) );
  OR2_X2 U9146 ( .A1(n13251), .A2(n13250), .ZN(n13253) );
  NAND2_X1 U9147 ( .A1(n14281), .A2(n14282), .ZN(n14278) );
  NAND2_X1 U9148 ( .A1(n6761), .A2(n14424), .ZN(n6853) );
  NOR2_X2 U9149 ( .A1(n12993), .A2(n12900), .ZN(n12902) );
  NAND2_X1 U9150 ( .A1(n6932), .A2(n8846), .ZN(n6931) );
  OR4_X2 U9151 ( .A1(n13998), .A2(n13903), .A3(n14034), .A4(n8823), .ZN(n8824)
         );
  OAI21_X1 U9152 ( .B1(n11284), .B2(n7134), .A(n7132), .ZN(n11378) );
  INV_X1 U9153 ( .A(n7134), .ZN(n7133) );
  OR2_X1 U9154 ( .A1(n9097), .A2(n8785), .ZN(n8468) );
  OR2_X1 U9155 ( .A1(n7714), .A2(n7713), .ZN(n7715) );
  INV_X1 U9156 ( .A(n7275), .ZN(n7274) );
  NAND2_X2 U9157 ( .A1(n7716), .A2(n7508), .ZN(n7733) );
  NAND2_X2 U9158 ( .A1(n7714), .A2(n7713), .ZN(n7716) );
  INV_X1 U9159 ( .A(n7298), .ZN(n13996) );
  NAND2_X1 U9160 ( .A1(n14039), .A2(n14049), .ZN(n7282) );
  OAI21_X1 U9161 ( .B1(n6608), .B2(n6720), .A(n11794), .ZN(n11795) );
  NAND2_X1 U9162 ( .A1(n11796), .A2(n6721), .ZN(n11805) );
  OAI21_X1 U9163 ( .B1(n11822), .B2(n11824), .A(n11847), .ZN(n11823) );
  NOR2_X2 U9164 ( .A1(n8380), .A2(n8310), .ZN(n13797) );
  INV_X1 U9165 ( .A(n11808), .ZN(n7345) );
  NAND3_X1 U9166 ( .A1(n7119), .A2(n7118), .A3(n10329), .ZN(n7114) );
  NAND2_X1 U9167 ( .A1(n15408), .A2(n15409), .ZN(n15407) );
  INV_X1 U9168 ( .A(n8247), .ZN(n6860) );
  OR2_X1 U9169 ( .A1(n8252), .A2(n15420), .ZN(n8253) );
  INV_X1 U9170 ( .A(n6851), .ZN(n6757) );
  INV_X1 U9171 ( .A(n8279), .ZN(n6762) );
  INV_X1 U9172 ( .A(n8259), .ZN(n6728) );
  XNOR2_X1 U9173 ( .A(n8240), .B(P1_ADDR_REG_5__SCAN_IN), .ZN(n8259) );
  NAND2_X1 U9174 ( .A1(n6731), .A2(n6729), .ZN(P1_U3214) );
  NAND2_X1 U9175 ( .A1(n13612), .A2(n14395), .ZN(n6731) );
  NAND2_X1 U9176 ( .A1(n7531), .A2(n7530), .ZN(n7852) );
  AND2_X1 U9177 ( .A1(n7130), .A2(n11464), .ZN(n6734) );
  AND2_X2 U9178 ( .A1(n6733), .A2(n7011), .ZN(n12295) );
  NAND2_X1 U9179 ( .A1(n12254), .A2(n12313), .ZN(n6733) );
  OR2_X1 U9180 ( .A1(n10193), .A2(n15202), .ZN(n9803) );
  NAND2_X1 U9181 ( .A1(n7003), .A2(n7009), .ZN(n12329) );
  INV_X1 U9182 ( .A(n6944), .ZN(n6943) );
  OAI21_X1 U9183 ( .B1(n11066), .B2(n11062), .A(n11063), .ZN(n11068) );
  AND3_X2 U9184 ( .A1(n9499), .A2(n7409), .A3(n7410), .ZN(n9723) );
  NAND2_X1 U9185 ( .A1(n6564), .A2(n6600), .ZN(n6735) );
  NAND2_X1 U9186 ( .A1(n11454), .A2(n12213), .ZN(n7071) );
  NAND2_X1 U9188 ( .A1(n8134), .A2(n8133), .ZN(n13303) );
  INV_X1 U9189 ( .A(n13288), .ZN(n6738) );
  INV_X1 U9190 ( .A(n7057), .ZN(n13212) );
  NAND2_X1 U9191 ( .A1(n8129), .A2(n8128), .ZN(n11454) );
  OAI21_X1 U9192 ( .B1(n8121), .B2(n7076), .A(n7073), .ZN(n10985) );
  NAND4_X1 U9193 ( .A1(n13936), .A2(n6740), .A3(n13989), .A4(n13948), .ZN(
        n6739) );
  OR4_X2 U9194 ( .A1(n8822), .A2(n14068), .A3(n14086), .A4(n14063), .ZN(n8823)
         );
  NOR2_X1 U9195 ( .A1(n6574), .A2(n11007), .ZN(n6930) );
  AOI21_X1 U9196 ( .B1(n14069), .B2(n14070), .A(n13870), .ZN(n14054) );
  NOR2_X1 U9197 ( .A1(n14938), .A2(n10896), .ZN(n14957) );
  NOR2_X1 U9198 ( .A1(n6743), .A2(n12705), .ZN(n6742) );
  INV_X1 U9199 ( .A(n12400), .ZN(n6743) );
  XNOR2_X1 U9200 ( .A(n7026), .B(n14946), .ZN(n14939) );
  NOR2_X1 U9201 ( .A1(n14831), .A2(n7029), .ZN(n14851) );
  NOR2_X1 U9202 ( .A1(n14903), .A2(n10894), .ZN(n14922) );
  NOR2_X1 U9203 ( .A1(n14849), .A2(n7025), .ZN(n10890) );
  XNOR2_X1 U9204 ( .A(n10890), .B(n7024), .ZN(n14868) );
  NAND2_X1 U9205 ( .A1(n7735), .A2(n7511), .ZN(n7752) );
  NAND2_X1 U9206 ( .A1(n6794), .A2(n6792), .ZN(n14237) );
  OAI21_X1 U9207 ( .B1(n14140), .B2(n14560), .A(n6977), .ZN(n6976) );
  NAND2_X1 U9208 ( .A1(n12956), .A2(n12955), .ZN(n12954) );
  OAI21_X1 U9209 ( .B1(n7497), .B2(SI_5_), .A(n7498), .ZN(n7663) );
  NAND2_X1 U9210 ( .A1(n7125), .A2(n7126), .ZN(n12931) );
  NAND2_X2 U9211 ( .A1(n7973), .A2(n12217), .ZN(n13223) );
  NAND2_X2 U9212 ( .A1(n11447), .A2(n11446), .ZN(n11449) );
  INV_X1 U9213 ( .A(n7095), .ZN(n7094) );
  OAI22_X1 U9214 ( .A1(n10988), .A2(n7819), .B1(n14374), .B2(n12034), .ZN(
        n14357) );
  NAND2_X1 U9215 ( .A1(n7093), .A2(n7092), .ZN(n10652) );
  XNOR2_X2 U9216 ( .A(n7898), .B(SI_18_), .ZN(n7895) );
  AND2_X1 U9217 ( .A1(n12902), .A2(n12903), .ZN(n6749) );
  NAND2_X1 U9218 ( .A1(n7248), .A2(n7246), .ZN(n7680) );
  NAND2_X1 U9219 ( .A1(n6750), .A2(n8561), .ZN(n7302) );
  NAND2_X1 U9220 ( .A1(n14509), .A2(n10318), .ZN(n10501) );
  NAND2_X2 U9221 ( .A1(n13976), .A2(n13883), .ZN(n13966) );
  NAND2_X1 U9222 ( .A1(n7282), .A2(n7280), .ZN(n13878) );
  NAND2_X4 U9223 ( .A1(n8376), .A2(n9727), .ZN(n8796) );
  AOI21_X2 U9224 ( .B1(n6751), .B2(n14497), .A(n13929), .ZN(n14149) );
  XNOR2_X2 U9225 ( .A(n14589), .B(n13772), .ZN(n9757) );
  NAND2_X2 U9226 ( .A1(n8381), .A2(n8382), .ZN(n14589) );
  NAND2_X1 U9227 ( .A1(n6766), .A2(P3_ADDR_REG_4__SCAN_IN), .ZN(n6765) );
  NAND2_X1 U9228 ( .A1(n14019), .A2(n13903), .ZN(n6773) );
  NAND4_X4 U9229 ( .A1(n8363), .A2(n8362), .A3(n8361), .A4(n8360), .ZN(n14556)
         );
  INV_X1 U9230 ( .A(n6776), .ZN(n14557) );
  NAND2_X1 U9231 ( .A1(n9748), .A2(n9749), .ZN(n9752) );
  NAND2_X1 U9232 ( .A1(n9654), .A2(n6776), .ZN(n6775) );
  NAND2_X1 U9233 ( .A1(n14071), .A2(n6547), .ZN(n6777) );
  NAND3_X1 U9234 ( .A1(n6777), .A2(n6778), .A3(n6604), .ZN(n13902) );
  NAND2_X1 U9235 ( .A1(n6672), .A2(n6782), .ZN(n11146) );
  NAND2_X1 U9236 ( .A1(n6790), .A2(n6791), .ZN(n14257) );
  NAND2_X1 U9237 ( .A1(n6791), .A2(n7428), .ZN(n8320) );
  NAND2_X1 U9238 ( .A1(n13308), .A2(n6796), .ZN(n13259) );
  AND2_X1 U9239 ( .A1(n13163), .A2(n6805), .ZN(n13155) );
  NAND2_X1 U9240 ( .A1(n13163), .A2(n8169), .ZN(n13164) );
  NAND2_X1 U9241 ( .A1(n13163), .A2(n6803), .ZN(n13154) );
  NAND3_X1 U9242 ( .A1(n6802), .A2(n6801), .A3(n6799), .ZN(n13150) );
  OR2_X1 U9243 ( .A1(n13163), .A2(n12174), .ZN(n6801) );
  NAND2_X1 U9244 ( .A1(n13163), .A2(n6662), .ZN(n6802) );
  INV_X1 U9245 ( .A(n6812), .ZN(n11450) );
  NAND2_X1 U9246 ( .A1(n6664), .A2(n10470), .ZN(n6817) );
  OAI21_X2 U9247 ( .B1(n11994), .B2(n6822), .A(n6820), .ZN(n12001) );
  NOR2_X1 U9248 ( .A1(n12001), .A2(n12000), .ZN(n12002) );
  NAND2_X1 U9249 ( .A1(n6823), .A2(n6824), .ZN(n7308) );
  NAND2_X1 U9250 ( .A1(n12018), .A2(n6609), .ZN(n6823) );
  AOI21_X1 U9251 ( .B1(n7306), .B2(n7305), .A(n6619), .ZN(n6831) );
  NAND2_X1 U9252 ( .A1(n12061), .A2(n6561), .ZN(n6833) );
  NAND2_X1 U9253 ( .A1(n12086), .A2(n6543), .ZN(n6839) );
  NAND2_X1 U9254 ( .A1(n11925), .A2(n11921), .ZN(n6841) );
  NOR2_X4 U9255 ( .A1(n6841), .A2(n11924), .ZN(n11977) );
  NAND2_X1 U9256 ( .A1(n11928), .A2(n11977), .ZN(n11923) );
  NOR2_X1 U9257 ( .A1(n6616), .A2(n11976), .ZN(n6845) );
  AOI21_X1 U9258 ( .B1(n14301), .B2(n14300), .A(n6852), .ZN(n6851) );
  NAND2_X1 U9259 ( .A1(n6853), .A2(n6854), .ZN(n6857) );
  INV_X1 U9260 ( .A(n6857), .ZN(n14431) );
  INV_X1 U9261 ( .A(n14432), .ZN(n6856) );
  INV_X1 U9262 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n6858) );
  INV_X1 U9263 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n6859) );
  NAND2_X1 U9264 ( .A1(n10635), .A2(n6673), .ZN(n10704) );
  NAND2_X2 U9265 ( .A1(n10637), .A2(n10636), .ZN(n10635) );
  AOI21_X2 U9266 ( .B1(n11612), .B2(n6867), .A(n6650), .ZN(n12559) );
  NAND2_X1 U9267 ( .A1(n11612), .A2(n11611), .ZN(n12575) );
  INV_X1 U9268 ( .A(n11611), .ZN(n6870) );
  AND2_X2 U9269 ( .A1(n6874), .A2(n6657), .ZN(n12623) );
  OR2_X2 U9270 ( .A1(n12677), .A2(n6656), .ZN(n6874) );
  NAND2_X1 U9271 ( .A1(n9723), .A2(n6877), .ZN(n6876) );
  NAND2_X1 U9272 ( .A1(n9723), .A2(n9719), .ZN(n12876) );
  NAND2_X1 U9273 ( .A1(n12548), .A2(n6882), .ZN(n6880) );
  NAND2_X1 U9274 ( .A1(n12548), .A2(n6886), .ZN(n6881) );
  NAND2_X1 U9275 ( .A1(n12548), .A2(n11614), .ZN(n12541) );
  OR2_X2 U9276 ( .A1(n12548), .A2(n6884), .ZN(n6878) );
  INV_X1 U9277 ( .A(n6962), .ZN(n6888) );
  NAND3_X1 U9278 ( .A1(n6902), .A2(n6901), .A3(n6677), .ZN(n6900) );
  AOI21_X1 U9279 ( .B1(n9895), .B2(n9246), .A(n6904), .ZN(n6905) );
  NAND2_X1 U9280 ( .A1(n6907), .A2(n6906), .ZN(n6909) );
  NAND2_X1 U9281 ( .A1(n6910), .A2(n6624), .ZN(n6906) );
  NAND2_X1 U9282 ( .A1(n6909), .A2(n9757), .ZN(n8394) );
  INV_X1 U9283 ( .A(n8369), .ZN(n6910) );
  OAI21_X1 U9284 ( .B1(n8745), .B2(n6558), .A(n6916), .ZN(n8760) );
  NAND3_X1 U9285 ( .A1(n8660), .A2(n6920), .A3(n6678), .ZN(n6919) );
  NAND2_X1 U9286 ( .A1(n6921), .A2(n6922), .ZN(n8646) );
  NAND2_X1 U9287 ( .A1(n8618), .A2(n6924), .ZN(n6921) );
  OR2_X1 U9288 ( .A1(n7162), .A2(n6931), .ZN(n6929) );
  NAND3_X1 U9289 ( .A1(n6929), .A2(n6928), .A3(n8857), .ZN(P1_U3242) );
  NAND2_X1 U9290 ( .A1(n7162), .A2(n6930), .ZN(n6928) );
  NAND2_X1 U9291 ( .A1(n6933), .A2(n6936), .ZN(n8735) );
  NAND3_X1 U9292 ( .A1(n8714), .A2(n6934), .A3(n8713), .ZN(n6933) );
  NAND3_X1 U9293 ( .A1(n6940), .A2(n8427), .A3(n6674), .ZN(n6939) );
  OAI21_X1 U9294 ( .B1(n8426), .B2(n8425), .A(n8424), .ZN(n6940) );
  NAND3_X1 U9295 ( .A1(n8348), .A2(n8305), .A3(n8337), .ZN(n8341) );
  NAND4_X1 U9296 ( .A1(n6984), .A2(n8862), .A3(n8861), .A4(n8865), .ZN(n6941)
         );
  AND3_X2 U9297 ( .A1(n6554), .A2(n6943), .A3(n6942), .ZN(n9499) );
  NAND4_X1 U9298 ( .A1(n6984), .A2(n8862), .A3(n8861), .A4(n6945), .ZN(n6944)
         );
  NAND2_X1 U9299 ( .A1(n7410), .A2(n9499), .ZN(n9721) );
  NAND2_X2 U9300 ( .A1(n12550), .A2(n12549), .ZN(n12548) );
  NAND2_X2 U9301 ( .A1(n12559), .A2(n6610), .ZN(n12550) );
  OAI21_X2 U9302 ( .B1(n12690), .B2(n11603), .A(n11602), .ZN(n12677) );
  AND2_X2 U9303 ( .A1(n11102), .A2(n11101), .ZN(n11104) );
  OR2_X2 U9304 ( .A1(n14077), .A2(n14197), .ZN(n14055) );
  OR2_X2 U9305 ( .A1(n14098), .A2(n14203), .ZN(n14077) );
  NAND2_X1 U9306 ( .A1(n14127), .A2(n14546), .ZN(n14131) );
  XNOR2_X1 U9307 ( .A(n6963), .B(n8803), .ZN(n14127) );
  NOR2_X1 U9308 ( .A1(n13916), .A2(n8808), .ZN(n6963) );
  NAND2_X2 U9309 ( .A1(n11640), .A2(n14264), .ZN(n8376) );
  NAND3_X1 U9310 ( .A1(n6675), .A2(n8561), .A3(n7439), .ZN(n6965) );
  AND3_X4 U9311 ( .A1(n6593), .A2(n8311), .A3(n8310), .ZN(n8561) );
  NAND2_X1 U9312 ( .A1(n6975), .A2(n6973), .ZN(P1_U3525) );
  OR2_X1 U9313 ( .A1(n14645), .A2(n6974), .ZN(n6973) );
  NAND2_X1 U9314 ( .A1(n6979), .A2(n13916), .ZN(n14139) );
  OR2_X1 U9315 ( .A1(n13930), .A2(n13917), .ZN(n6980) );
  NAND2_X1 U9316 ( .A1(n14042), .A2(n6981), .ZN(n13984) );
  INV_X1 U9317 ( .A(P3_IR_REG_8__SCAN_IN), .ZN(n6986) );
  NAND3_X1 U9318 ( .A1(n9089), .A2(n9088), .A3(n15180), .ZN(n9689) );
  NAND2_X1 U9319 ( .A1(n6987), .A2(n6711), .ZN(n9790) );
  NOR2_X1 U9320 ( .A1(n9090), .A2(P3_D_REG_1__SCAN_IN), .ZN(n6988) );
  INV_X1 U9321 ( .A(n12321), .ZN(n6992) );
  NAND2_X1 U9322 ( .A1(n11170), .A2(n6559), .ZN(n6996) );
  NAND2_X1 U9323 ( .A1(n12254), .A2(n7002), .ZN(n7001) );
  XNOR2_X1 U9324 ( .A(n10191), .B(n12348), .ZN(n10008) );
  XNOR2_X1 U9325 ( .A(n10525), .B(n10110), .ZN(n10191) );
  AND2_X2 U9326 ( .A1(n9808), .A2(n9807), .ZN(n10525) );
  NAND2_X1 U9327 ( .A1(n9499), .A2(n6668), .ZN(n8876) );
  NAND2_X1 U9328 ( .A1(n9499), .A2(n8866), .ZN(n9524) );
  NAND2_X1 U9329 ( .A1(n7016), .A2(n7017), .ZN(n12484) );
  NAND3_X1 U9330 ( .A1(n7032), .A2(n7031), .A3(n6709), .ZN(n12455) );
  MUX2_X1 U9331 ( .A(n9888), .B(n14966), .S(P3_IR_REG_0__SCAN_IN), .Z(n9889)
         );
  NAND2_X1 U9332 ( .A1(n14349), .A2(n7048), .ZN(n7046) );
  NAND2_X1 U9333 ( .A1(n7046), .A2(n7047), .ZN(n11401) );
  INV_X1 U9334 ( .A(n13225), .ZN(n7054) );
  AOI21_X1 U9335 ( .B1(n13225), .B2(n13224), .A(n6594), .ZN(n7057) );
  OAI21_X2 U9336 ( .B1(n7054), .B2(n7053), .A(n7051), .ZN(n13182) );
  AND2_X1 U9337 ( .A1(n6602), .A2(n7459), .ZN(n7065) );
  NAND4_X1 U9338 ( .A1(n7065), .A2(n7064), .A3(n7453), .A4(n7062), .ZN(n7304)
         );
  AND3_X2 U9339 ( .A1(n7458), .A2(n7614), .A3(n7066), .ZN(n7738) );
  NAND2_X1 U9340 ( .A1(n7068), .A2(n7067), .ZN(n10482) );
  NAND2_X1 U9341 ( .A1(n7071), .A2(n7069), .ZN(n8134) );
  NAND2_X1 U9342 ( .A1(n7072), .A2(n6666), .ZN(n10141) );
  OR2_X1 U9343 ( .A1(n10168), .A2(n8109), .ZN(n7072) );
  AOI21_X1 U9344 ( .B1(n7075), .B2(n7074), .A(n6634), .ZN(n7073) );
  NAND2_X1 U9345 ( .A1(n9544), .A2(n8099), .ZN(n9535) );
  OAI22_X1 U9346 ( .A1(n7592), .A2(n8951), .B1(n9273), .B2(n13058), .ZN(n7593)
         );
  NOR2_X1 U9347 ( .A1(n14440), .A2(n14439), .ZN(n14438) );
  NOR2_X1 U9348 ( .A1(n14436), .A2(n14435), .ZN(n14434) );
  OAI21_X1 U9349 ( .B1(n11066), .B2(n11065), .A(n11064), .ZN(n11067) );
  NAND2_X2 U9350 ( .A1(n9273), .A2(n9727), .ZN(n7592) );
  AOI211_X2 U9351 ( .C1(n13365), .C2(n14378), .A(n13364), .B(n13363), .ZN(
        n13439) );
  INV_X1 U9352 ( .A(n11067), .ZN(n11073) );
  NAND2_X1 U9353 ( .A1(n9812), .A2(n9811), .ZN(n9967) );
  OAI21_X2 U9354 ( .B1(n15385), .B2(n11083), .A(n11082), .ZN(n11170) );
  NAND2_X1 U9355 ( .A1(n9968), .A2(n9969), .ZN(n10010) );
  NOR2_X4 U9356 ( .A1(n14055), .A2(n14190), .ZN(n14042) );
  INV_X2 U9357 ( .A(n8378), .ZN(n8310) );
  NOR2_X1 U9358 ( .A1(n14555), .A2(n14589), .ZN(n14548) );
  XNOR2_X2 U9359 ( .A(n9004), .B(P3_IR_REG_2__SCAN_IN), .ZN(n10046) );
  INV_X1 U9360 ( .A(n7593), .ZN(n7595) );
  OAI22_X2 U9361 ( .A1(n13240), .A2(n8145), .B1(n13247), .B2(n13030), .ZN(
        n13225) );
  NAND2_X1 U9362 ( .A1(n10482), .A2(n8118), .ZN(n10416) );
  OAI22_X1 U9363 ( .A1(n13303), .A2(n8135), .B1(n12189), .B2(n13406), .ZN(
        n13288) );
  NAND2_X2 U9364 ( .A1(n7639), .A2(n7638), .ZN(n11965) );
  NAND2_X1 U9365 ( .A1(n13223), .A2(n7086), .ZN(n7084) );
  AND2_X1 U9366 ( .A1(n7580), .A2(n7579), .ZN(n7091) );
  NAND2_X1 U9367 ( .A1(n13051), .A2(n12090), .ZN(n11934) );
  NAND2_X1 U9368 ( .A1(n10486), .A2(n7094), .ZN(n7093) );
  AOI21_X1 U9369 ( .B1(n7094), .B2(n7096), .A(n6617), .ZN(n7092) );
  NAND2_X1 U9370 ( .A1(n7100), .A2(n6670), .ZN(n11412) );
  OAI21_X1 U9371 ( .B1(n11449), .B2(n6607), .A(n7101), .ZN(n13285) );
  NAND2_X1 U9372 ( .A1(n13253), .A2(n7105), .ZN(n7973) );
  INV_X1 U9373 ( .A(n7961), .ZN(n7107) );
  NAND4_X1 U9374 ( .A1(n6555), .A2(n7108), .A3(n7738), .A4(n7571), .ZN(n7464)
         );
  NAND2_X1 U9375 ( .A1(n9831), .A2(n7112), .ZN(n7111) );
  NAND2_X1 U9376 ( .A1(n7114), .A2(n7116), .ZN(n10976) );
  INV_X1 U9377 ( .A(n11465), .ZN(n7127) );
  NAND2_X1 U9378 ( .A1(n11465), .A2(n7130), .ZN(n7125) );
  INV_X1 U9379 ( .A(n7129), .ZN(n12886) );
  NOR2_X1 U9380 ( .A1(n12886), .A2(n12885), .ZN(n13005) );
  NAND3_X1 U9381 ( .A1(n7143), .A2(n9551), .A3(n9552), .ZN(n7144) );
  NAND2_X1 U9382 ( .A1(n9450), .A2(n9451), .ZN(n9552) );
  INV_X1 U9383 ( .A(n9576), .ZN(n7143) );
  XNOR2_X1 U9384 ( .A(n9578), .B(n9577), .ZN(n9576) );
  XNOR2_X1 U9385 ( .A(n12942), .B(n11965), .ZN(n9578) );
  INV_X1 U9386 ( .A(n7149), .ZN(n12919) );
  NAND2_X1 U9387 ( .A1(n8760), .A2(n7153), .ZN(n7150) );
  NAND2_X1 U9388 ( .A1(n7150), .A2(n7151), .ZN(n8772) );
  NAND4_X1 U9389 ( .A1(n6593), .A2(n8336), .A3(n8310), .A4(n8311), .ZN(n7160)
         );
  OR2_X1 U9390 ( .A1(n8827), .A2(n8829), .ZN(n7161) );
  NAND2_X1 U9391 ( .A1(n8775), .A2(n8774), .ZN(n7162) );
  OAI22_X1 U9392 ( .A1(n8470), .A2(n6680), .B1(n8471), .B2(n7164), .ZN(n8489)
         );
  NAND2_X1 U9393 ( .A1(n8489), .A2(n8490), .ZN(n8488) );
  OAI22_X1 U9394 ( .A1(n8505), .A2(n7166), .B1(n8506), .B2(n7167), .ZN(n8516)
         );
  OAI22_X1 U9395 ( .A1(n8697), .A2(n7168), .B1(n8698), .B2(n7169), .ZN(n8709)
         );
  NAND2_X1 U9396 ( .A1(n8709), .A2(n8710), .ZN(n8708) );
  NOR2_X1 U9397 ( .A1(n7172), .A2(n7171), .ZN(n7170) );
  INV_X1 U9398 ( .A(n13518), .ZN(n7171) );
  NAND2_X1 U9399 ( .A1(n13514), .A2(n13513), .ZN(n14394) );
  NAND2_X1 U9400 ( .A1(n7174), .A2(n8903), .ZN(n9839) );
  NAND2_X1 U9401 ( .A1(n11239), .A2(n7182), .ZN(n7180) );
  NAND2_X1 U9402 ( .A1(n7180), .A2(n7181), .ZN(n14392) );
  NAND2_X1 U9403 ( .A1(n13731), .A2(n13609), .ZN(n13610) );
  OAI211_X1 U9404 ( .C1(n13731), .C2(n6681), .A(n7187), .B(n7185), .ZN(n13649)
         );
  NAND2_X1 U9405 ( .A1(n13731), .A2(n7186), .ZN(n7185) );
  NOR2_X1 U9406 ( .A1(n7189), .A2(n13643), .ZN(n7186) );
  OAI22_X1 U9407 ( .A1(n7189), .A2(n7188), .B1(n13643), .B2(n7191), .ZN(n7187)
         );
  NOR2_X1 U9408 ( .A1(n13643), .A2(n13611), .ZN(n7188) );
  INV_X1 U9409 ( .A(n13643), .ZN(n7190) );
  NAND2_X1 U9410 ( .A1(n13692), .A2(n7194), .ZN(n7193) );
  INV_X1 U9411 ( .A(n10606), .ZN(n7201) );
  NAND2_X1 U9412 ( .A1(n7208), .A2(n7210), .ZN(n10293) );
  NAND3_X1 U9413 ( .A1(n9842), .A2(n7209), .A3(n9925), .ZN(n7208) );
  NAND2_X1 U9414 ( .A1(n13716), .A2(n7217), .ZN(n7214) );
  NAND2_X1 U9415 ( .A1(n8795), .A2(n6537), .ZN(n7231) );
  NAND2_X1 U9416 ( .A1(n7233), .A2(n7232), .ZN(n7531) );
  NAND2_X1 U9417 ( .A1(n7821), .A2(n7528), .ZN(n7233) );
  NAND2_X1 U9418 ( .A1(n7555), .A2(n7243), .ZN(n7242) );
  NAND2_X1 U9419 ( .A1(n7641), .A2(n7249), .ZN(n7248) );
  NAND2_X1 U9420 ( .A1(n7641), .A2(n7495), .ZN(n7644) );
  NAND3_X1 U9421 ( .A1(n7252), .A2(n7251), .A3(P1_DATAO_REG_1__SCAN_IN), .ZN(
        n7253) );
  OAI21_X2 U9422 ( .B1(n7488), .B2(n8950), .A(n7253), .ZN(n7480) );
  NAND2_X1 U9423 ( .A1(n7254), .A2(n6691), .ZN(n7550) );
  NAND2_X2 U9424 ( .A1(n7258), .A2(n7537), .ZN(n7898) );
  INV_X2 U9425 ( .A(n14565), .ZN(n14580) );
  NOR2_X1 U9426 ( .A1(n9059), .A2(n13778), .ZN(n7279) );
  NAND2_X1 U9427 ( .A1(n7283), .A2(n6663), .ZN(n14104) );
  NAND2_X1 U9428 ( .A1(n13966), .A2(n7287), .ZN(n7286) );
  NAND2_X1 U9429 ( .A1(n7286), .A2(n7288), .ZN(n13887) );
  NAND2_X1 U9430 ( .A1(n9863), .A2(n9862), .ZN(n7296) );
  XNOR2_X1 U9431 ( .A(n7296), .B(n14524), .ZN(n14525) );
  NAND2_X1 U9432 ( .A1(n14009), .A2(n6667), .ZN(n7300) );
  CLKBUF_X1 U9433 ( .A(n7300), .Z(n7298) );
  NAND2_X1 U9434 ( .A1(n11976), .A2(n6616), .ZN(n7303) );
  INV_X1 U9435 ( .A(n12017), .ZN(n7307) );
  INV_X1 U9436 ( .A(n12029), .ZN(n7309) );
  INV_X1 U9437 ( .A(n12028), .ZN(n7310) );
  NAND2_X1 U9438 ( .A1(n12078), .A2(n7313), .ZN(n7312) );
  INV_X1 U9439 ( .A(n12081), .ZN(n7314) );
  NAND3_X1 U9440 ( .A1(n11985), .A2(n6632), .A3(n7315), .ZN(n7317) );
  INV_X1 U9441 ( .A(n6613), .ZN(n7316) );
  NAND2_X1 U9442 ( .A1(n7317), .A2(n7318), .ZN(n11994) );
  INV_X1 U9443 ( .A(n11988), .ZN(n7319) );
  NAND2_X1 U9444 ( .A1(n9680), .A2(n7333), .ZN(n7332) );
  NAND2_X1 U9445 ( .A1(n9037), .A2(n9038), .ZN(n7338) );
  NAND2_X1 U9446 ( .A1(n11004), .A2(n11114), .ZN(n11549) );
  OAI21_X1 U9447 ( .B1(n9013), .B2(n8970), .A(n8971), .ZN(n9007) );
  NAND2_X1 U9448 ( .A1(n8970), .A2(n8971), .ZN(n7357) );
  NAND2_X1 U9449 ( .A1(n9075), .A2(n7362), .ZN(n7358) );
  OAI211_X1 U9450 ( .C1(n9075), .C2(n7361), .A(n7358), .B(n7359), .ZN(n9154)
         );
  INV_X1 U9451 ( .A(n9077), .ZN(n7365) );
  NAND2_X1 U9452 ( .A1(n7371), .A2(P3_REG0_REG_3__SCAN_IN), .ZN(n9974) );
  NAND2_X1 U9453 ( .A1(n7371), .A2(P3_REG0_REG_7__SCAN_IN), .ZN(n10389) );
  NAND2_X1 U9454 ( .A1(n7371), .A2(P3_REG0_REG_6__SCAN_IN), .ZN(n10272) );
  NAND2_X1 U9455 ( .A1(n7371), .A2(P3_REG0_REG_5__SCAN_IN), .ZN(n10214) );
  NAND2_X1 U9456 ( .A1(n7371), .A2(P3_REG0_REG_13__SCAN_IN), .ZN(n11093) );
  NAND2_X1 U9457 ( .A1(n7371), .A2(P3_REG0_REG_15__SCAN_IN), .ZN(n11275) );
  NAND2_X1 U9458 ( .A1(n7371), .A2(P3_REG0_REG_23__SCAN_IN), .ZN(n9636) );
  NAND2_X1 U9459 ( .A1(n7371), .A2(P3_REG0_REG_24__SCAN_IN), .ZN(n11535) );
  NAND2_X1 U9460 ( .A1(n7371), .A2(P3_REG0_REG_25__SCAN_IN), .ZN(n11547) );
  NAND2_X1 U9461 ( .A1(n7371), .A2(P3_REG0_REG_27__SCAN_IN), .ZN(n11568) );
  NAND2_X1 U9462 ( .A1(n7371), .A2(P3_REG0_REG_26__SCAN_IN), .ZN(n11554) );
  NAND2_X1 U9463 ( .A1(n7371), .A2(P3_REG0_REG_28__SCAN_IN), .ZN(n10356) );
  NAND2_X1 U9464 ( .A1(n7371), .A2(P3_REG0_REG_29__SCAN_IN), .ZN(n10222) );
  NAND2_X1 U9465 ( .A1(n7371), .A2(P3_REG0_REG_30__SCAN_IN), .ZN(n10298) );
  AOI22_X1 U9466 ( .A1(n11567), .A2(P3_REG2_REG_21__SCAN_IN), .B1(
        P3_REG0_REG_21__SCAN_IN), .B2(n7371), .ZN(n9471) );
  AOI22_X1 U9467 ( .A1(n11567), .A2(P3_REG2_REG_22__SCAN_IN), .B1(
        P3_REG0_REG_22__SCAN_IN), .B2(n7371), .ZN(n11523) );
  AOI22_X1 U9468 ( .A1(n11567), .A2(P3_REG2_REG_20__SCAN_IN), .B1(
        P3_REG0_REG_20__SCAN_IN), .B2(n7371), .ZN(n11506) );
  INV_X2 U9469 ( .A(n9738), .ZN(n7371) );
  NAND2_X1 U9470 ( .A1(n10748), .A2(n7375), .ZN(n7374) );
  AND2_X1 U9471 ( .A1(n8864), .A2(n8863), .ZN(n7382) );
  NAND3_X1 U9472 ( .A1(n6687), .A2(n7382), .A3(n6942), .ZN(n7381) );
  NOR2_X1 U9473 ( .A1(n11821), .A2(n11669), .ZN(n7385) );
  NAND2_X1 U9474 ( .A1(n7390), .A2(n7388), .ZN(n12652) );
  OAI21_X1 U9475 ( .B1(n14980), .B2(n7394), .A(n7392), .ZN(n11480) );
  OAI21_X1 U9476 ( .B1(n7400), .B2(n12563), .A(n7398), .ZN(n12530) );
  OAI21_X1 U9477 ( .B1(n12634), .B2(n7406), .A(n7404), .ZN(n11514) );
  NAND2_X1 U9478 ( .A1(n7417), .A2(n7416), .ZN(n14071) );
  NAND2_X1 U9479 ( .A1(n7419), .A2(n13892), .ZN(n7416) );
  INV_X1 U9480 ( .A(n13938), .ZN(n14146) );
  BUF_X8 U9481 ( .A(n10531), .Z(n11892) );
  INV_X2 U9482 ( .A(n11521), .ZN(n11436) );
  NAND2_X1 U9483 ( .A1(n11915), .A2(n15057), .ZN(n11912) );
  INV_X1 U9484 ( .A(n12192), .ZN(n9539) );
  AOI21_X2 U9485 ( .B1(n11871), .B2(n12665), .A(n12317), .ZN(n12264) );
  NAND2_X1 U9486 ( .A1(n7550), .A2(n7549), .ZN(n7935) );
  NAND2_X1 U9487 ( .A1(n8189), .A2(n8188), .ZN(n8192) );
  AOI21_X2 U9488 ( .B1(n10501), .B2(n10500), .A(n10499), .ZN(n14490) );
  MUX2_X1 U9489 ( .A(n8384), .B(n8383), .S(n14589), .Z(n8393) );
  NAND2_X1 U9490 ( .A1(n8181), .A2(n8180), .ZN(n8184) );
  AOI21_X2 U9491 ( .B1(n10976), .B2(n10975), .A(n10974), .ZN(n11284) );
  NAND2_X2 U9492 ( .A1(n11432), .A2(n11431), .ZN(n11867) );
  OR2_X1 U9493 ( .A1(n7612), .A2(n8963), .ZN(n7594) );
  OAI21_X2 U9494 ( .B1(n10764), .B2(n7803), .A(n7802), .ZN(n10988) );
  NAND2_X1 U9495 ( .A1(n12178), .A2(n12177), .ZN(n12231) );
  INV_X1 U9496 ( .A(n12037), .ZN(n12040) );
  XNOR2_X2 U9497 ( .A(n10038), .B(n8955), .ZN(n9999) );
  OR2_X1 U9498 ( .A1(n12003), .A2(n12002), .ZN(n12007) );
  INV_X1 U9499 ( .A(n8842), .ZN(n8843) );
  NAND2_X1 U9500 ( .A1(n10632), .A2(n11830), .ZN(n10631) );
  NOR2_X2 U9501 ( .A1(n14635), .A2(n14503), .ZN(n10816) );
  NAND2_X1 U9502 ( .A1(n15017), .A2(n15025), .ZN(n11683) );
  INV_X1 U9503 ( .A(n9381), .ZN(n11339) );
  MUX2_X1 U9504 ( .A(n11688), .B(n10097), .S(n10525), .Z(n9812) );
  NAND2_X2 U9505 ( .A1(n7471), .A2(n7470), .ZN(n8199) );
  INV_X1 U9506 ( .A(n7471), .ZN(n11906) );
  NOR2_X2 U9507 ( .A1(n12530), .A2(n12531), .ZN(n12529) );
  AND2_X1 U9508 ( .A1(n11212), .A2(n11253), .ZN(n7430) );
  OR2_X1 U9509 ( .A1(n12838), .A2(n12837), .ZN(P3_U3446) );
  OR2_X1 U9510 ( .A1(n12762), .A2(n12761), .ZN(P3_U3478) );
  AND2_X1 U9511 ( .A1(n14070), .A2(n8643), .ZN(n7434) );
  INV_X1 U9512 ( .A(n13406), .ZN(n8168) );
  OR2_X1 U9513 ( .A1(n11018), .A2(n10857), .ZN(n7435) );
  AND3_X1 U9514 ( .A1(n12229), .A2(n13167), .A3(n8092), .ZN(n7437) );
  AND2_X1 U9515 ( .A1(n13473), .A2(n8051), .ZN(n7438) );
  AND2_X1 U9516 ( .A1(n14985), .A2(n11474), .ZN(n7440) );
  NOR2_X1 U9517 ( .A1(n11718), .A2(n11831), .ZN(n7441) );
  INV_X1 U9518 ( .A(n14063), .ZN(n13871) );
  INV_X1 U9519 ( .A(n15041), .ZN(n15029) );
  AND2_X1 U9520 ( .A1(n13023), .A2(n8200), .ZN(n7442) );
  INV_X1 U9521 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n7460) );
  NOR3_X1 U9522 ( .A1(n12229), .A2(n12226), .A3(n13167), .ZN(n12227) );
  INV_X1 U9523 ( .A(n11007), .ZN(n8846) );
  INV_X1 U9524 ( .A(n13250), .ZN(n7960) );
  OR2_X1 U9525 ( .A1(n13353), .A2(n14367), .ZN(n7443) );
  AND3_X1 U9526 ( .A1(n8587), .A2(n8586), .A3(n8585), .ZN(n7444) );
  AND2_X1 U9527 ( .A1(n10104), .A2(n10103), .ZN(n7445) );
  AND2_X1 U9528 ( .A1(n12090), .A2(n11928), .ZN(n7446) );
  INV_X1 U9529 ( .A(n13163), .ZN(n13186) );
  INV_X1 U9530 ( .A(n10310), .ZN(n14512) );
  INV_X1 U9531 ( .A(n12341), .ZN(n12679) );
  AOI21_X1 U9532 ( .B1(n12525), .B2(n11566), .A(n10358), .ZN(n12250) );
  INV_X1 U9533 ( .A(n12615), .ZN(n12591) );
  AND2_X1 U9534 ( .A1(n12125), .A2(n12124), .ZN(n7447) );
  AND2_X1 U9535 ( .A1(n9862), .A2(n8404), .ZN(n7448) );
  AND2_X1 U9536 ( .A1(n13543), .A2(n13542), .ZN(n7449) );
  INV_X1 U9537 ( .A(n11995), .ZN(n11996) );
  INV_X1 U9538 ( .A(n11295), .ZN(n8572) );
  NOR2_X1 U9539 ( .A1(n8573), .A2(n8572), .ZN(n8574) );
  INV_X1 U9540 ( .A(n12038), .ZN(n12039) );
  NAND2_X1 U9541 ( .A1(n8630), .A2(n6588), .ZN(n8631) );
  NAND2_X1 U9542 ( .A1(n12186), .A2(n12135), .ZN(n12148) );
  INV_X1 U9543 ( .A(P3_IR_REG_24__SCAN_IN), .ZN(n9376) );
  AND2_X1 U9544 ( .A1(n14556), .A2(n14580), .ZN(n9660) );
  INV_X1 U9545 ( .A(n12250), .ZN(n11616) );
  INV_X1 U9546 ( .A(n11834), .ZN(n11047) );
  INV_X1 U9547 ( .A(P3_IR_REG_14__SCAN_IN), .ZN(n8865) );
  INV_X1 U9548 ( .A(n14358), .ZN(n8125) );
  INV_X1 U9549 ( .A(n7919), .ZN(n7546) );
  NOR2_X1 U9550 ( .A1(n7513), .A2(n9039), .ZN(n7512) );
  INV_X1 U9551 ( .A(P3_REG3_REG_9__SCAN_IN), .ZN(n10557) );
  OR2_X1 U9552 ( .A1(n11596), .A2(n11595), .ZN(n12699) );
  INV_X1 U9553 ( .A(n11835), .ZN(n11103) );
  INV_X1 U9554 ( .A(P3_IR_REG_19__SCAN_IN), .ZN(n9682) );
  NAND2_X1 U9555 ( .A1(n12894), .A2(n12896), .ZN(n12897) );
  INV_X1 U9556 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n7741) );
  INV_X1 U9557 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n7686) );
  INV_X1 U9558 ( .A(n14356), .ZN(n8167) );
  INV_X1 U9559 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n7457) );
  INV_X1 U9560 ( .A(n8726), .ZN(n8725) );
  INV_X1 U9561 ( .A(n7948), .ZN(n7555) );
  INV_X1 U9562 ( .A(n12807), .ZN(n11887) );
  NAND2_X1 U9563 ( .A1(n11876), .A2(n12615), .ZN(n11877) );
  AND2_X1 U9564 ( .A1(n11266), .A2(n11267), .ZN(n11265) );
  NOR2_X1 U9565 ( .A1(n9504), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n11502) );
  INV_X1 U9566 ( .A(n6527), .ZN(n9736) );
  NAND2_X1 U9567 ( .A1(n10558), .A2(n10557), .ZN(n10570) );
  NAND2_X1 U9568 ( .A1(n10703), .A2(n11826), .ZN(n10748) );
  AND2_X1 U9569 ( .A1(n9817), .A2(n12501), .ZN(n9799) );
  XNOR2_X1 U9570 ( .A(n9444), .B(n11932), .ZN(n9446) );
  NAND2_X1 U9571 ( .A1(n7468), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n8024) );
  NAND2_X1 U9572 ( .A1(n7938), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n7952) );
  OR2_X1 U9573 ( .A1(n7795), .A2(n7794), .ZN(n7813) );
  OR2_X1 U9574 ( .A1(n8041), .A2(n7597), .ZN(n7599) );
  OR2_X1 U9575 ( .A1(n14693), .A2(n14692), .ZN(n14695) );
  INV_X1 U9576 ( .A(n13356), .ZN(n8169) );
  INV_X1 U9577 ( .A(n12211), .ZN(n7870) );
  NAND2_X1 U9578 ( .A1(n7772), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n7795) );
  NOR2_X1 U9579 ( .A1(n7687), .A2(n7686), .ZN(n7705) );
  AND2_X1 U9580 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n7672) );
  INV_X2 U9581 ( .A(n7612), .ZN(n7908) );
  INV_X1 U9582 ( .A(n10470), .ZN(n10487) );
  INV_X1 U9583 ( .A(n14391), .ZN(n13513) );
  AND2_X1 U9584 ( .A1(n13552), .A2(n13551), .ZN(n13553) );
  INV_X1 U9585 ( .A(n13664), .ZN(n11238) );
  INV_X1 U9586 ( .A(n13548), .ZN(n13636) );
  NAND2_X1 U9587 ( .A1(n8566), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n8592) );
  NAND2_X1 U9588 ( .A1(n8725), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n8748) );
  NAND2_X1 U9589 ( .A1(n8700), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n8715) );
  OR2_X1 U9590 ( .A1(n8592), .A2(n8591), .ZN(n8610) );
  OR2_X1 U9591 ( .A1(n8448), .A2(n9208), .ZN(n8474) );
  INV_X1 U9592 ( .A(n14271), .ZN(n8929) );
  NAND2_X1 U9593 ( .A1(n7527), .A2(n11261), .ZN(n7528) );
  INV_X1 U9594 ( .A(n7616), .ZN(n7489) );
  NOR2_X1 U9595 ( .A1(P1_ADDR_REG_7__SCAN_IN), .A2(n8267), .ZN(n8218) );
  NOR2_X1 U9596 ( .A1(n8283), .A2(n8282), .ZN(n8229) );
  OR2_X1 U9597 ( .A1(n11662), .A2(n15188), .ZN(n11560) );
  INV_X1 U9598 ( .A(n12691), .ZN(n11868) );
  INV_X1 U9599 ( .A(n12592), .ZN(n12313) );
  OR2_X1 U9600 ( .A1(n11435), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n9504) );
  OR2_X1 U9601 ( .A1(n10395), .A2(n9819), .ZN(n12336) );
  INV_X1 U9602 ( .A(n9799), .ZN(n11853) );
  AND3_X1 U9603 ( .A1(n9472), .A2(n9471), .A3(n9470), .ZN(n12615) );
  OAI21_X1 U9604 ( .B1(n11436), .B2(n10044), .A(n9391), .ZN(n9395) );
  OR2_X1 U9605 ( .A1(n11520), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n11533) );
  AND2_X1 U9606 ( .A1(n11502), .A2(n11501), .ZN(n11504) );
  AND2_X1 U9607 ( .A1(n11321), .A2(n11320), .ZN(n11433) );
  OR2_X1 U9608 ( .A1(n10109), .A2(n15022), .ZN(n12535) );
  INV_X1 U9609 ( .A(n9805), .ZN(n10085) );
  OAI21_X1 U9610 ( .B1(n12250), .B2(n15029), .A(n11622), .ZN(n11623) );
  OR2_X1 U9611 ( .A1(n12677), .A2(n12676), .ZN(n12681) );
  NAND2_X1 U9612 ( .A1(n11738), .A2(n11733), .ZN(n14982) );
  INV_X1 U9613 ( .A(n15018), .ZN(n15049) );
  NAND2_X1 U9614 ( .A1(n10884), .A2(n10883), .ZN(n11000) );
  NAND2_X1 U9615 ( .A1(n9677), .A2(n9676), .ZN(n9680) );
  OR2_X1 U9616 ( .A1(n7813), .A2(n7812), .ZN(n7827) );
  OR2_X1 U9617 ( .A1(n8092), .A2(n11925), .ZN(n9421) );
  AND2_X1 U9618 ( .A1(n7926), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n7938) );
  OR2_X1 U9619 ( .A1(n7864), .A2(n7863), .ZN(n7882) );
  AND2_X1 U9620 ( .A1(n14720), .A2(n14719), .ZN(n14722) );
  OR2_X1 U9621 ( .A1(n14821), .A2(n8204), .ZN(n8205) );
  NAND2_X1 U9622 ( .A1(n9540), .A2(n7604), .ZN(n9531) );
  AND2_X1 U9623 ( .A1(n9415), .A2(n14772), .ZN(n8201) );
  AND2_X1 U9624 ( .A1(n13599), .A2(n13598), .ZN(n13671) );
  NAND2_X1 U9625 ( .A1(n13545), .A2(n13546), .ZN(n13547) );
  INV_X1 U9626 ( .A(n8399), .ZN(n8674) );
  INV_X1 U9627 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n9162) );
  INV_X1 U9628 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n9208) );
  INV_X1 U9629 ( .A(n13913), .ZN(n13914) );
  INV_X1 U9630 ( .A(n13869), .ZN(n13870) );
  INV_X1 U9631 ( .A(n14107), .ZN(n14561) );
  OR2_X1 U9632 ( .A1(n9058), .A2(n9128), .ZN(n14581) );
  AND2_X1 U9633 ( .A1(n8912), .A2(n8911), .ZN(n9655) );
  OR2_X1 U9634 ( .A1(n8542), .A2(P1_IR_REG_12__SCAN_IN), .ZN(n8543) );
  OR2_X1 U9635 ( .A1(n8511), .A2(P1_IR_REG_10__SCAN_IN), .ZN(n8526) );
  AOI21_X1 U9636 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(n8230), .A(n8229), .ZN(
        n8286) );
  OR2_X1 U9637 ( .A1(n9881), .A2(n9880), .ZN(n14834) );
  INV_X1 U9638 ( .A(n12336), .ZN(n15389) );
  INV_X1 U9639 ( .A(n15395), .ZN(n12333) );
  AND2_X1 U9640 ( .A1(n11574), .A2(n11573), .ZN(n12521) );
  AND3_X1 U9641 ( .A1(n11524), .A2(n11523), .A3(n11522), .ZN(n12577) );
  INV_X1 U9642 ( .A(n12498), .ZN(n14973) );
  INV_X1 U9643 ( .A(n15031), .ZN(n15038) );
  NAND2_X1 U9644 ( .A1(n9795), .A2(n9800), .ZN(n10089) );
  INV_X1 U9645 ( .A(n15020), .ZN(n15055) );
  AND2_X1 U9646 ( .A1(n12667), .A2(n12666), .ZN(n12843) );
  INV_X1 U9647 ( .A(n15083), .ZN(n12748) );
  NAND2_X1 U9648 ( .A1(n15043), .A2(n15058), .ZN(n15083) );
  NAND2_X1 U9649 ( .A1(n11860), .A2(n6527), .ZN(n15018) );
  INV_X1 U9650 ( .A(n14342), .ZN(n12973) );
  NAND2_X1 U9651 ( .A1(n9414), .A2(n13323), .ZN(n13019) );
  OR2_X1 U9652 ( .A1(n7995), .A2(n13166), .ZN(n8029) );
  OR2_X1 U9653 ( .A1(n14712), .A2(n14713), .ZN(n14714) );
  INV_X1 U9654 ( .A(n14739), .ZN(n14754) );
  INV_X1 U9655 ( .A(n14745), .ZN(n14756) );
  INV_X1 U9656 ( .A(n13311), .ZN(n14355) );
  OR2_X1 U9657 ( .A1(n9433), .A2(n8091), .ZN(n8170) );
  INV_X1 U9658 ( .A(n14791), .ZN(n14378) );
  AND2_X1 U9659 ( .A1(n8080), .A2(n8079), .ZN(n9409) );
  OR2_X1 U9660 ( .A1(n8068), .A2(P2_IR_REG_24__SCAN_IN), .ZN(n8070) );
  AND2_X1 U9661 ( .A1(n7669), .A2(n7701), .ZN(n14681) );
  NAND2_X1 U9662 ( .A1(n10293), .A2(n10292), .ZN(n10605) );
  INV_X1 U9663 ( .A(n14401), .ZN(n13740) );
  OR2_X1 U9664 ( .A1(n8752), .A2(n13954), .ZN(n8738) );
  AND2_X1 U9665 ( .A1(n8654), .A2(n8653), .ZN(n14074) );
  OR2_X1 U9666 ( .A1(n9056), .A2(n8846), .ZN(n9113) );
  INV_X1 U9667 ( .A(n14464), .ZN(n14478) );
  INV_X1 U9668 ( .A(n11212), .ZN(n11221) );
  INV_X1 U9669 ( .A(n14542), .ZN(n14567) );
  NAND2_X1 U9670 ( .A1(n13921), .A2(n14542), .ZN(n14543) );
  AND2_X1 U9671 ( .A1(n8925), .A2(n9353), .ZN(n9253) );
  INV_X1 U9672 ( .A(n14581), .ZN(n14108) );
  INV_X1 U9673 ( .A(n14641), .ZN(n14611) );
  AND2_X1 U9674 ( .A1(n9358), .A2(n9357), .ZN(n9657) );
  OAI211_X1 U9675 ( .C1(P1_B_REG_SCAN_IN), .C2(n11225), .A(n8910), .B(n14265), 
        .ZN(n9356) );
  XNOR2_X1 U9676 ( .A(n8343), .B(P1_IR_REG_21__SCAN_IN), .ZN(n9242) );
  INV_X1 U9677 ( .A(n14834), .ZN(n14969) );
  AND2_X1 U9678 ( .A1(n10021), .A2(n10020), .ZN(n15395) );
  INV_X1 U9679 ( .A(n12338), .ZN(n12327) );
  INV_X1 U9680 ( .A(n12577), .ZN(n12604) );
  OR3_X1 U9681 ( .A1(n11441), .A2(n11440), .A3(n11439), .ZN(n12341) );
  OR2_X1 U9682 ( .A1(n9795), .A2(n8878), .ZN(n12350) );
  OR2_X1 U9683 ( .A1(n9887), .A2(n12490), .ZN(n12498) );
  OR2_X1 U9684 ( .A1(n9887), .A2(n9878), .ZN(n14977) );
  AND2_X1 U9685 ( .A1(n10109), .A2(n15020), .ZN(n15052) );
  OR2_X1 U9686 ( .A1(n10090), .A2(n10089), .ZN(n15020) );
  INV_X1 U9687 ( .A(n12782), .ZN(n12780) );
  INV_X1 U9688 ( .A(n15096), .ZN(n15094) );
  INV_X1 U9689 ( .A(n12730), .ZN(n12791) );
  INV_X2 U9690 ( .A(n15086), .ZN(n15085) );
  AND2_X1 U9691 ( .A1(n9877), .A2(P3_STATE_REG_SCAN_IN), .ZN(n9800) );
  NAND2_X1 U9692 ( .A1(n9090), .A2(n9800), .ZN(n9156) );
  INV_X1 U9693 ( .A(SI_14_), .ZN(n11261) );
  INV_X1 U9694 ( .A(SI_10_), .ZN(n9039) );
  NAND2_X1 U9695 ( .A1(n9557), .A2(P2_STATE_REG_SCAN_IN), .ZN(n14348) );
  NAND2_X1 U9696 ( .A1(n9423), .A2(n9422), .ZN(n14342) );
  OR2_X1 U9697 ( .A1(n7849), .A2(n7848), .ZN(n14337) );
  INV_X1 U9698 ( .A(n14752), .ZN(n14736) );
  AND2_X1 U9699 ( .A1(n10771), .A2(n10770), .ZN(n14385) );
  NAND2_X1 U9700 ( .A1(n13281), .A2(n8096), .ZN(n13342) );
  AND2_X2 U9701 ( .A1(n13323), .A2(n8170), .ZN(n14367) );
  AND2_X2 U9702 ( .A1(n9435), .A2(n9434), .ZN(n14829) );
  INV_X1 U9703 ( .A(n13159), .ZN(n13436) );
  INV_X1 U9704 ( .A(n13263), .ZN(n13456) );
  AND2_X1 U9705 ( .A1(n14385), .A2(n14384), .ZN(n14390) );
  INV_X1 U9706 ( .A(n14821), .ZN(n14819) );
  AND2_X2 U9707 ( .A1(n9435), .A2(n8202), .ZN(n14821) );
  INV_X1 U9708 ( .A(n14766), .ZN(n14767) );
  INV_X1 U9709 ( .A(n14203), .ZN(n14079) );
  INV_X1 U9710 ( .A(n14186), .ZN(n14033) );
  INV_X1 U9711 ( .A(n14398), .ZN(n13743) );
  NAND4_X1 U9712 ( .A1(n8741), .A2(n8740), .A3(n8739), .A4(n8738), .ZN(n13910)
         );
  INV_X1 U9713 ( .A(n14083), .ZN(n14123) );
  AND2_X2 U9714 ( .A1(n9359), .A2(n9253), .ZN(n14658) );
  INV_X1 U9715 ( .A(n14645), .ZN(n14643) );
  AND2_X1 U9716 ( .A1(n8939), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9187) );
  INV_X1 U9717 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n15293) );
  INV_X1 U9718 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n9959) );
  INV_X1 U9719 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n9512) );
  XNOR2_X1 U9720 ( .A(n8303), .B(n8302), .ZN(n8304) );
  INV_X2 U9721 ( .A(n12350), .ZN(P3_U3897) );
  AND2_X1 U9722 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9272), .ZN(P2_U3947) );
  NOR2_X1 U9723 ( .A1(P2_IR_REG_16__SCAN_IN), .A2(P2_IR_REG_15__SCAN_IN), .ZN(
        n7451) );
  NOR2_X1 U9724 ( .A1(P2_IR_REG_17__SCAN_IN), .A2(P2_IR_REG_19__SCAN_IN), .ZN(
        n7450) );
  INV_X1 U9725 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n7455) );
  NOR2_X2 U9726 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n7589) );
  AND2_X2 U9727 ( .A1(n7589), .A2(n7457), .ZN(n7614) );
  NOR3_X1 U9728 ( .A1(P2_IR_REG_24__SCAN_IN), .A2(P2_IR_REG_9__SCAN_IN), .A3(
        P2_IR_REG_25__SCAN_IN), .ZN(n7459) );
  INV_X1 U9729 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n7461) );
  AND2_X1 U9730 ( .A1(n7461), .A2(n7571), .ZN(n7462) );
  NAND2_X1 U9731 ( .A1(n7570), .A2(n7462), .ZN(n13474) );
  XNOR2_X2 U9732 ( .A(n7463), .B(P2_IR_REG_30__SCAN_IN), .ZN(n7471) );
  NAND2_X1 U9733 ( .A1(n8195), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n7476) );
  INV_X1 U9734 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n7466) );
  OR2_X1 U9735 ( .A1(n8157), .A2(n7466), .ZN(n7475) );
  NAND2_X1 U9736 ( .A1(n7672), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n7687) );
  NAND2_X1 U9737 ( .A1(n7705), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n7725) );
  INV_X1 U9738 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n7794) );
  INV_X1 U9739 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n7812) );
  INV_X1 U9740 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n7826) );
  NAND2_X1 U9741 ( .A1(n7843), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n7864) );
  INV_X1 U9742 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n7863) );
  INV_X1 U9743 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n15294) );
  INV_X1 U9744 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n12998) );
  NAND2_X1 U9745 ( .A1(n7967), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n7966) );
  INV_X1 U9746 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n15355) );
  NAND2_X1 U9747 ( .A1(n7994), .A2(n15355), .ZN(n7469) );
  NAND2_X1 U9748 ( .A1(n8024), .A2(n7469), .ZN(n13203) );
  OR2_X1 U9749 ( .A1(n8041), .A2(n13203), .ZN(n7474) );
  INV_X1 U9750 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n7472) );
  OR2_X1 U9751 ( .A1(n8199), .A2(n7472), .ZN(n7473) );
  NAND4_X1 U9752 ( .A1(n7476), .A2(n7475), .A3(n7474), .A4(n7473), .ZN(n13027)
         );
  NAND2_X1 U9753 ( .A1(n7480), .A2(SI_1_), .ZN(n7483) );
  OAI21_X1 U9754 ( .B1(SI_1_), .B2(n7480), .A(n7483), .ZN(n7585) );
  INV_X1 U9755 ( .A(n7585), .ZN(n7482) );
  INV_X1 U9756 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n8954) );
  NOR2_X1 U9757 ( .A1(n7481), .A2(n9728), .ZN(n7583) );
  NAND2_X1 U9758 ( .A1(n7587), .A2(n7483), .ZN(n7486) );
  INV_X1 U9759 ( .A(n7486), .ZN(n7485) );
  INV_X1 U9760 ( .A(SI_2_), .ZN(n7484) );
  NAND2_X1 U9761 ( .A1(n7486), .A2(SI_2_), .ZN(n7490) );
  MUX2_X1 U9762 ( .A(n8988), .B(n8967), .S(n9729), .Z(n7616) );
  MUX2_X1 U9763 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(P1_DATAO_REG_3__SCAN_IN), 
        .S(n9729), .Z(n7491) );
  NAND2_X1 U9764 ( .A1(n7491), .A2(SI_3_), .ZN(n7493) );
  OAI21_X1 U9765 ( .B1(n7491), .B2(SI_3_), .A(n7493), .ZN(n7631) );
  INV_X1 U9766 ( .A(n7631), .ZN(n7492) );
  NAND2_X1 U9767 ( .A1(n7633), .A2(n7493), .ZN(n7641) );
  MUX2_X1 U9768 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(P1_DATAO_REG_4__SCAN_IN), 
        .S(n9729), .Z(n7494) );
  INV_X1 U9769 ( .A(n7642), .ZN(n7495) );
  MUX2_X1 U9770 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(P1_DATAO_REG_5__SCAN_IN), 
        .S(n9729), .Z(n7497) );
  NAND2_X1 U9771 ( .A1(n7497), .A2(SI_5_), .ZN(n7498) );
  INV_X8 U9772 ( .A(n7499), .ZN(n9727) );
  MUX2_X1 U9773 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(P1_DATAO_REG_6__SCAN_IN), 
        .S(n9727), .Z(n7500) );
  NAND2_X1 U9774 ( .A1(n7500), .A2(SI_6_), .ZN(n7502) );
  OAI21_X1 U9775 ( .B1(n7500), .B2(SI_6_), .A(n7502), .ZN(n7501) );
  INV_X1 U9776 ( .A(n7501), .ZN(n7679) );
  NAND2_X1 U9777 ( .A1(n7680), .A2(n7679), .ZN(n7682) );
  MUX2_X1 U9778 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(P1_DATAO_REG_7__SCAN_IN), 
        .S(n9727), .Z(n7503) );
  OAI21_X1 U9779 ( .B1(n7503), .B2(SI_7_), .A(n7505), .ZN(n7504) );
  INV_X1 U9780 ( .A(n7504), .ZN(n7699) );
  NAND2_X1 U9781 ( .A1(n7698), .A2(n7505), .ZN(n7714) );
  MUX2_X1 U9782 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(P1_DATAO_REG_8__SCAN_IN), 
        .S(n9727), .Z(n7506) );
  OAI21_X1 U9783 ( .B1(n7506), .B2(SI_8_), .A(n7508), .ZN(n7507) );
  INV_X1 U9784 ( .A(n7507), .ZN(n7713) );
  MUX2_X1 U9785 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(P1_DATAO_REG_9__SCAN_IN), 
        .S(n9727), .Z(n7509) );
  OAI21_X1 U9786 ( .B1(n7509), .B2(SI_9_), .A(n7511), .ZN(n7510) );
  INV_X1 U9787 ( .A(n7510), .ZN(n7732) );
  MUX2_X1 U9788 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(P1_DATAO_REG_10__SCAN_IN), 
        .S(n9727), .Z(n7750) );
  NAND2_X1 U9789 ( .A1(n7513), .A2(n9039), .ZN(n7765) );
  MUX2_X1 U9790 ( .A(n9398), .B(n15272), .S(n9727), .Z(n7520) );
  NAND2_X1 U9791 ( .A1(n7520), .A2(n11070), .ZN(n7519) );
  MUX2_X1 U9792 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(P1_DATAO_REG_12__SCAN_IN), 
        .S(n9727), .Z(n7518) );
  INV_X1 U9793 ( .A(n7518), .ZN(n7514) );
  NAND2_X1 U9794 ( .A1(n7514), .A2(n15330), .ZN(n7517) );
  MUX2_X1 U9795 ( .A(n9515), .B(n15367), .S(n9727), .Z(n7516) );
  NAND2_X1 U9796 ( .A1(n7516), .A2(n11163), .ZN(n7515) );
  INV_X1 U9797 ( .A(n7515), .ZN(n7525) );
  XNOR2_X1 U9798 ( .A(n7516), .B(SI_13_), .ZN(n7807) );
  INV_X1 U9799 ( .A(n7517), .ZN(n7523) );
  XNOR2_X1 U9800 ( .A(n7518), .B(n15330), .ZN(n7784) );
  INV_X1 U9801 ( .A(n7519), .ZN(n7521) );
  XNOR2_X1 U9802 ( .A(n7520), .B(SI_11_), .ZN(n7766) );
  OR2_X2 U9803 ( .A1(n7521), .A2(n7766), .ZN(n7782) );
  OR2_X2 U9804 ( .A1(n7523), .A2(n7522), .ZN(n7805) );
  AND2_X2 U9805 ( .A1(n7807), .A2(n7805), .ZN(n7524) );
  MUX2_X1 U9806 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(P1_DATAO_REG_14__SCAN_IN), 
        .S(n9727), .Z(n7820) );
  MUX2_X1 U9807 ( .A(n9785), .B(n15325), .S(n9727), .Z(n7529) );
  INV_X1 U9808 ( .A(SI_15_), .ZN(n11315) );
  NAND2_X1 U9809 ( .A1(n7529), .A2(n11315), .ZN(n7530) );
  MUX2_X1 U9810 ( .A(n9915), .B(n15181), .S(n9727), .Z(n7533) );
  NAND2_X2 U9811 ( .A1(n7852), .A2(n7851), .ZN(n7535) );
  INV_X1 U9812 ( .A(SI_16_), .ZN(n7532) );
  NAND2_X1 U9813 ( .A1(n7533), .A2(n7532), .ZN(n7534) );
  MUX2_X1 U9814 ( .A(n9959), .B(n9961), .S(n9729), .Z(n7872) );
  NAND2_X1 U9815 ( .A1(n7536), .A2(SI_17_), .ZN(n7537) );
  MUX2_X1 U9816 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(P1_DATAO_REG_19__SCAN_IN), 
        .S(n9727), .Z(n7542) );
  MUX2_X1 U9817 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(P1_DATAO_REG_18__SCAN_IN), 
        .S(n9727), .Z(n7896) );
  INV_X1 U9818 ( .A(n7896), .ZN(n7538) );
  INV_X1 U9819 ( .A(SI_18_), .ZN(n9619) );
  NOR2_X1 U9820 ( .A1(n7896), .A2(SI_18_), .ZN(n7541) );
  NAND2_X1 U9821 ( .A1(n7902), .A2(n7541), .ZN(n7544) );
  INV_X1 U9822 ( .A(n7542), .ZN(n7543) );
  INV_X1 U9823 ( .A(SI_19_), .ZN(n15312) );
  NAND2_X1 U9824 ( .A1(n7543), .A2(n15312), .ZN(n7901) );
  MUX2_X1 U9825 ( .A(n15263), .B(n10497), .S(n9727), .Z(n7921) );
  NOR2_X1 U9826 ( .A1(n7548), .A2(SI_20_), .ZN(n7545) );
  NAND2_X1 U9827 ( .A1(n7548), .A2(SI_20_), .ZN(n7549) );
  MUX2_X1 U9828 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(P1_DATAO_REG_21__SCAN_IN), 
        .S(n9727), .Z(n7552) );
  XNOR2_X1 U9829 ( .A(n7552), .B(SI_21_), .ZN(n7934) );
  INV_X1 U9830 ( .A(n7934), .ZN(n7551) );
  NAND2_X1 U9831 ( .A1(n7935), .A2(n7551), .ZN(n7554) );
  NAND2_X1 U9832 ( .A1(n7552), .A2(SI_21_), .ZN(n7553) );
  MUX2_X1 U9833 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(P1_DATAO_REG_22__SCAN_IN), 
        .S(n9729), .Z(n7949) );
  NAND2_X1 U9834 ( .A1(n7556), .A2(SI_22_), .ZN(n7557) );
  MUX2_X1 U9835 ( .A(n15293), .B(n11013), .S(n9727), .Z(n7558) );
  INV_X1 U9836 ( .A(n7558), .ZN(n7559) );
  NAND2_X1 U9837 ( .A1(n7559), .A2(SI_23_), .ZN(n7560) );
  MUX2_X1 U9838 ( .A(n7368), .B(n11228), .S(n9727), .Z(n7561) );
  XNOR2_X1 U9839 ( .A(n7561), .B(SI_24_), .ZN(n7974) );
  INV_X1 U9840 ( .A(n7561), .ZN(n7562) );
  NAND2_X1 U9841 ( .A1(n7562), .A2(SI_24_), .ZN(n7563) );
  MUX2_X1 U9842 ( .A(n15297), .B(n15170), .S(n9727), .Z(n7565) );
  INV_X1 U9843 ( .A(SI_25_), .ZN(n11540) );
  NAND2_X1 U9844 ( .A1(n7565), .A2(n11540), .ZN(n7568) );
  INV_X1 U9845 ( .A(n7565), .ZN(n7566) );
  NAND2_X1 U9846 ( .A1(n7566), .A2(SI_25_), .ZN(n7567) );
  NAND2_X1 U9847 ( .A1(n7568), .A2(n7567), .ZN(n7987) );
  INV_X1 U9848 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n14267) );
  INV_X1 U9849 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n13487) );
  MUX2_X1 U9850 ( .A(n14267), .B(n13487), .S(n9727), .Z(n8003) );
  XNOR2_X1 U9851 ( .A(n8003), .B(SI_26_), .ZN(n7569) );
  INV_X1 U9852 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n7573) );
  NAND2_X2 U9853 ( .A1(n8155), .A2(n13484), .ZN(n9273) );
  NAND2_X1 U9854 ( .A1(n13486), .A2(n6537), .ZN(n7576) );
  OR2_X1 U9855 ( .A1(n8193), .A2(n13487), .ZN(n7575) );
  INV_X1 U9856 ( .A(n13027), .ZN(n8150) );
  INV_X1 U9857 ( .A(n13205), .ZN(n13446) );
  NAND2_X1 U9858 ( .A1(n7605), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n7582) );
  INV_X1 U9859 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n7577) );
  OR2_X1 U9860 ( .A1(n7625), .A2(n7577), .ZN(n7581) );
  INV_X1 U9861 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n9322) );
  OR2_X1 U9862 ( .A1(n7607), .A2(n9322), .ZN(n7580) );
  INV_X1 U9863 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n7578) );
  OR2_X1 U9864 ( .A1(n8041), .A2(n7578), .ZN(n7579) );
  INV_X1 U9865 ( .A(n7583), .ZN(n7584) );
  NAND2_X1 U9866 ( .A1(n7585), .A2(n7584), .ZN(n7586) );
  NAND2_X1 U9867 ( .A1(n7587), .A2(n7586), .ZN(n8951) );
  NAND2_X1 U9868 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(n15206), .ZN(n7588) );
  MUX2_X1 U9869 ( .A(P2_IR_REG_31__SCAN_IN), .B(n7588), .S(
        P2_IR_REG_1__SCAN_IN), .Z(n7591) );
  INV_X1 U9870 ( .A(n7589), .ZN(n7590) );
  NAND2_X1 U9871 ( .A1(n7591), .A2(n7590), .ZN(n13058) );
  NAND2_X1 U9872 ( .A1(n7596), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n7601) );
  NAND2_X1 U9873 ( .A1(n7605), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n7600) );
  INV_X1 U9874 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n7597) );
  INV_X1 U9875 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n9279) );
  OR2_X1 U9876 ( .A1(n7607), .A2(n9279), .ZN(n7598) );
  INV_X1 U9877 ( .A(n15206), .ZN(n7603) );
  NAND2_X1 U9878 ( .A1(n9729), .A2(SI_0_), .ZN(n7602) );
  XNOR2_X1 U9879 ( .A(n7602), .B(n8954), .ZN(n13489) );
  INV_X1 U9880 ( .A(n11922), .ZN(n11935) );
  NAND2_X1 U9881 ( .A1(n11928), .A2(n11935), .ZN(n9541) );
  INV_X1 U9882 ( .A(n13051), .ZN(n8098) );
  INV_X1 U9883 ( .A(n11932), .ZN(n10444) );
  NAND2_X1 U9884 ( .A1(n8098), .A2(n10444), .ZN(n7604) );
  INV_X1 U9885 ( .A(n8041), .ZN(n7940) );
  NAND2_X1 U9886 ( .A1(n7940), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n7610) );
  INV_X1 U9887 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n7606) );
  OR2_X1 U9888 ( .A1(n7625), .A2(n7606), .ZN(n7609) );
  INV_X1 U9889 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n9321) );
  OR2_X1 U9890 ( .A1(n7607), .A2(n9321), .ZN(n7608) );
  NOR2_X1 U9891 ( .A1(n7589), .A2(n6522), .ZN(n7613) );
  MUX2_X1 U9892 ( .A(n13473), .B(n7613), .S(P2_IR_REG_2__SCAN_IN), .Z(n7615)
         );
  NOR2_X1 U9893 ( .A1(n7615), .A2(n7614), .ZN(n13068) );
  NAND2_X1 U9894 ( .A1(n7617), .A2(n7616), .ZN(n7618) );
  AND2_X1 U9895 ( .A1(n7619), .A2(n7618), .ZN(n8952) );
  NAND2_X1 U9896 ( .A1(n8952), .A2(n8037), .ZN(n7620) );
  NAND2_X1 U9897 ( .A1(n9531), .A2(n9534), .ZN(n9530) );
  INV_X1 U9898 ( .A(n13050), .ZN(n8100) );
  INV_X1 U9899 ( .A(n6524), .ZN(n10453) );
  NAND2_X1 U9900 ( .A1(n8100), .A2(n10453), .ZN(n7622) );
  NAND2_X1 U9901 ( .A1(n9530), .A2(n7622), .ZN(n9518) );
  INV_X1 U9902 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n7623) );
  OR2_X1 U9903 ( .A1(n8156), .A2(n7623), .ZN(n7629) );
  OR2_X1 U9904 ( .A1(n8041), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n7628) );
  INV_X1 U9905 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n7624) );
  OR2_X1 U9906 ( .A1(n7625), .A2(n7624), .ZN(n7627) );
  INV_X1 U9907 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n9301) );
  OR2_X1 U9908 ( .A1(n8199), .A2(n9301), .ZN(n7626) );
  INV_X1 U9909 ( .A(n7630), .ZN(n7632) );
  NAND2_X1 U9910 ( .A1(n7632), .A2(n7631), .ZN(n7634) );
  AND2_X1 U9911 ( .A1(n7633), .A2(n7634), .ZN(n8986) );
  NAND2_X1 U9912 ( .A1(n8986), .A2(n6537), .ZN(n7639) );
  NAND2_X1 U9913 ( .A1(n7636), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7635) );
  MUX2_X1 U9914 ( .A(P2_IR_REG_31__SCAN_IN), .B(n7635), .S(
        P2_IR_REG_3__SCAN_IN), .Z(n7637) );
  OR2_X1 U9915 ( .A1(n7636), .A2(P2_IR_REG_3__SCAN_IN), .ZN(n7647) );
  AND2_X1 U9916 ( .A1(n7637), .A2(n7647), .ZN(n13081) );
  NAND2_X1 U9917 ( .A1(n9518), .A2(n12194), .ZN(n9517) );
  INV_X1 U9918 ( .A(n11965), .ZN(n10228) );
  NAND2_X1 U9919 ( .A1(n10228), .A2(n8104), .ZN(n7640) );
  NAND2_X1 U9920 ( .A1(n9517), .A2(n7640), .ZN(n9566) );
  INV_X1 U9921 ( .A(n7641), .ZN(n7643) );
  NAND2_X1 U9922 ( .A1(n7643), .A2(n7642), .ZN(n7645) );
  NAND2_X1 U9923 ( .A1(n7645), .A2(n7644), .ZN(n8993) );
  OR2_X1 U9924 ( .A1(n8993), .A2(n7592), .ZN(n7652) );
  NAND2_X1 U9925 ( .A1(n7647), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7646) );
  MUX2_X1 U9926 ( .A(n7646), .B(P2_IR_REG_31__SCAN_IN), .S(n7648), .Z(n7650)
         );
  INV_X1 U9927 ( .A(n7647), .ZN(n7649) );
  NAND2_X1 U9928 ( .A1(n7649), .A2(n7648), .ZN(n7666) );
  NAND2_X1 U9929 ( .A1(n7650), .A2(n7666), .ZN(n14660) );
  INV_X1 U9930 ( .A(n14660), .ZN(n14668) );
  AOI22_X1 U9931 ( .A1(n7908), .A2(P1_DATAO_REG_4__SCAN_IN), .B1(n7907), .B2(
        n14668), .ZN(n7651) );
  NAND2_X1 U9932 ( .A1(n8195), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n7661) );
  INV_X1 U9933 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n10128) );
  OR2_X1 U9934 ( .A1(n8199), .A2(n10128), .ZN(n7660) );
  INV_X1 U9935 ( .A(n7672), .ZN(n7656) );
  INV_X1 U9936 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n7654) );
  INV_X1 U9937 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n7653) );
  NAND2_X1 U9938 ( .A1(n7654), .A2(n7653), .ZN(n7655) );
  NAND2_X1 U9939 ( .A1(n7656), .A2(n7655), .ZN(n10129) );
  OR2_X1 U9940 ( .A1(n7995), .A2(n10129), .ZN(n7659) );
  INV_X1 U9941 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n7657) );
  XNOR2_X1 U9942 ( .A(n11973), .B(n13048), .ZN(n12195) );
  INV_X1 U9943 ( .A(n12195), .ZN(n9569) );
  INV_X1 U9944 ( .A(n11973), .ZN(n10130) );
  INV_X1 U9945 ( .A(n13048), .ZN(n11975) );
  NAND2_X1 U9946 ( .A1(n10130), .A2(n11975), .ZN(n7662) );
  XNOR2_X1 U9947 ( .A(n7664), .B(n7663), .ZN(n9062) );
  NAND2_X1 U9948 ( .A1(n9062), .A2(n6537), .ZN(n7671) );
  NAND2_X1 U9949 ( .A1(n7666), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7665) );
  MUX2_X1 U9950 ( .A(P2_IR_REG_31__SCAN_IN), .B(n7665), .S(
        P2_IR_REG_5__SCAN_IN), .Z(n7669) );
  INV_X1 U9951 ( .A(n7666), .ZN(n7668) );
  INV_X1 U9952 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n7667) );
  NAND2_X1 U9953 ( .A1(n7668), .A2(n7667), .ZN(n7701) );
  AOI22_X1 U9954 ( .A1(n7908), .A2(P1_DATAO_REG_5__SCAN_IN), .B1(n7907), .B2(
        n14681), .ZN(n7670) );
  NAND2_X1 U9955 ( .A1(n7671), .A2(n7670), .ZN(n11980) );
  NAND2_X1 U9956 ( .A1(n8040), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n7677) );
  INV_X1 U9957 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n9329) );
  OR2_X1 U9958 ( .A1(n8156), .A2(n9329), .ZN(n7676) );
  OAI21_X1 U9959 ( .B1(n7672), .B2(P2_REG3_REG_5__SCAN_IN), .A(n7687), .ZN(
        n10173) );
  OR2_X1 U9960 ( .A1(n7995), .A2(n10173), .ZN(n7675) );
  INV_X1 U9961 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n7673) );
  OR2_X1 U9962 ( .A1(n8157), .A2(n7673), .ZN(n7674) );
  NAND4_X1 U9963 ( .A1(n7677), .A2(n7676), .A3(n7675), .A4(n7674), .ZN(n13047)
         );
  NAND2_X1 U9964 ( .A1(n11980), .A2(n13047), .ZN(n7678) );
  OR2_X1 U9965 ( .A1(n7680), .A2(n7679), .ZN(n7681) );
  AND2_X1 U9966 ( .A1(n7682), .A2(n7681), .ZN(n9067) );
  NAND2_X1 U9967 ( .A1(n9067), .A2(n6537), .ZN(n7685) );
  NAND2_X1 U9968 ( .A1(n7701), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7683) );
  XNOR2_X1 U9969 ( .A(n7683), .B(P2_IR_REG_6__SCAN_IN), .ZN(n9370) );
  AOI22_X1 U9970 ( .A1(n7908), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n7907), .B2(
        n9370), .ZN(n7684) );
  NAND2_X1 U9971 ( .A1(n7685), .A2(n7684), .ZN(n14782) );
  NAND2_X1 U9972 ( .A1(n8040), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n7693) );
  NAND2_X1 U9973 ( .A1(n8195), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n7692) );
  AND2_X1 U9974 ( .A1(n7687), .A2(n7686), .ZN(n7688) );
  OR2_X1 U9975 ( .A1(n7688), .A2(n7705), .ZN(n10146) );
  OR2_X1 U9976 ( .A1(n7995), .A2(n10146), .ZN(n7691) );
  INV_X1 U9977 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n7689) );
  OR2_X1 U9978 ( .A1(n8157), .A2(n7689), .ZN(n7690) );
  NAND4_X1 U9979 ( .A1(n7693), .A2(n7692), .A3(n7691), .A4(n7690), .ZN(n13046)
         );
  INV_X1 U9980 ( .A(n13046), .ZN(n7694) );
  OR2_X1 U9981 ( .A1(n14782), .A2(n7694), .ZN(n7695) );
  NAND2_X1 U9982 ( .A1(n14782), .A2(n7694), .ZN(n8112) );
  AND2_X1 U9983 ( .A1(n7695), .A2(n8112), .ZN(n12198) );
  NAND2_X1 U9984 ( .A1(n10136), .A2(n10138), .ZN(n7697) );
  OR2_X1 U9985 ( .A1(n14782), .A2(n13046), .ZN(n7696) );
  NAND2_X1 U9986 ( .A1(n7697), .A2(n7696), .ZN(n10178) );
  OAI21_X1 U9987 ( .B1(n7700), .B2(n7699), .A(n7698), .ZN(n9086) );
  OAI21_X1 U9988 ( .B1(n7701), .B2(P2_IR_REG_6__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n7702) );
  XNOR2_X1 U9989 ( .A(n7702), .B(P2_IR_REG_7__SCAN_IN), .ZN(n13096) );
  AOI22_X1 U9990 ( .A1(n7908), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n7907), .B2(
        n13096), .ZN(n7703) );
  NAND2_X1 U9991 ( .A1(n8195), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n7711) );
  INV_X1 U9992 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n10182) );
  OR2_X1 U9993 ( .A1(n8199), .A2(n10182), .ZN(n7710) );
  OR2_X1 U9994 ( .A1(n7705), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n7706) );
  NAND2_X1 U9995 ( .A1(n7725), .A2(n7706), .ZN(n10186) );
  OR2_X1 U9996 ( .A1(n7995), .A2(n10186), .ZN(n7709) );
  INV_X1 U9997 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n7707) );
  OR2_X1 U9998 ( .A1(n8157), .A2(n7707), .ZN(n7708) );
  NAND4_X1 U9999 ( .A1(n7711), .A2(n7710), .A3(n7709), .A4(n7708), .ZN(n13045)
         );
  INV_X1 U10000 ( .A(n13045), .ZN(n11992) );
  XNOR2_X1 U10001 ( .A(n14788), .B(n11992), .ZN(n12200) );
  INV_X1 U10002 ( .A(n14788), .ZN(n10187) );
  NAND2_X1 U10003 ( .A1(n10187), .A2(n11992), .ZN(n7712) );
  NAND2_X1 U10004 ( .A1(n7717), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7718) );
  MUX2_X1 U10005 ( .A(P2_IR_REG_31__SCAN_IN), .B(n7718), .S(
        P2_IR_REG_8__SCAN_IN), .Z(n7719) );
  INV_X1 U10006 ( .A(n7719), .ZN(n7720) );
  NOR2_X1 U10007 ( .A1(n7720), .A2(n7738), .ZN(n13111) );
  AOI22_X1 U10008 ( .A1(n7908), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n7907), .B2(
        n13111), .ZN(n7721) );
  NAND2_X1 U10009 ( .A1(n8195), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n7730) );
  INV_X1 U10010 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n7723) );
  OR2_X1 U10011 ( .A1(n8157), .A2(n7723), .ZN(n7729) );
  NAND2_X1 U10012 ( .A1(n7725), .A2(n7724), .ZN(n7726) );
  NAND2_X1 U10013 ( .A1(n7742), .A2(n7726), .ZN(n10473) );
  OR2_X1 U10014 ( .A1(n7995), .A2(n10473), .ZN(n7728) );
  INV_X1 U10015 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n10474) );
  OR2_X1 U10016 ( .A1(n8199), .A2(n10474), .ZN(n7727) );
  NAND4_X1 U10017 ( .A1(n7730), .A2(n7729), .A3(n7728), .A4(n7727), .ZN(n13044) );
  XNOR2_X1 U10018 ( .A(n14795), .B(n13044), .ZN(n12201) );
  NAND2_X1 U10019 ( .A1(n14795), .A2(n13044), .ZN(n7731) );
  NAND2_X1 U10020 ( .A1(n7735), .A2(n7734), .ZN(n9174) );
  NOR2_X1 U10021 ( .A1(n7738), .A2(n13473), .ZN(n7736) );
  MUX2_X1 U10022 ( .A(n13473), .B(n7736), .S(P2_IR_REG_9__SCAN_IN), .Z(n7739)
         );
  NOR2_X1 U10023 ( .A1(n7739), .A2(n8049), .ZN(n9341) );
  AOI22_X1 U10024 ( .A1(n7908), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n7907), .B2(
        n9341), .ZN(n7740) );
  NAND2_X1 U10025 ( .A1(n8040), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n7748) );
  NAND2_X1 U10026 ( .A1(n8195), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n7747) );
  AND2_X1 U10027 ( .A1(n7742), .A2(n7741), .ZN(n7743) );
  OR2_X1 U10028 ( .A1(n7743), .A2(n7757), .ZN(n10246) );
  OR2_X1 U10029 ( .A1(n7995), .A2(n10246), .ZN(n7746) );
  INV_X1 U10030 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n7744) );
  OR2_X1 U10031 ( .A1(n8157), .A2(n7744), .ZN(n7745) );
  NAND4_X1 U10032 ( .A1(n7748), .A2(n7747), .A3(n7746), .A4(n7745), .ZN(n13042) );
  XNOR2_X1 U10033 ( .A(n12008), .B(n13042), .ZN(n12202) );
  NAND2_X1 U10034 ( .A1(n12008), .A2(n13042), .ZN(n7749) );
  XNOR2_X1 U10035 ( .A(n7750), .B(SI_10_), .ZN(n7751) );
  XNOR2_X1 U10036 ( .A(n7752), .B(n7751), .ZN(n9222) );
  NAND2_X1 U10037 ( .A1(n9222), .A2(n6537), .ZN(n7755) );
  OR2_X1 U10038 ( .A1(n8049), .A2(n13473), .ZN(n7753) );
  XNOR2_X1 U10039 ( .A(n7753), .B(P2_IR_REG_10__SCAN_IN), .ZN(n9343) );
  AOI22_X1 U10040 ( .A1(n7908), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n7907), 
        .B2(n9343), .ZN(n7754) );
  NAND2_X1 U10041 ( .A1(n7596), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n7762) );
  INV_X1 U10042 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n7756) );
  OR2_X1 U10043 ( .A1(n8156), .A2(n7756), .ZN(n7761) );
  NOR2_X1 U10044 ( .A1(n7757), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n7758) );
  OR2_X1 U10045 ( .A1(n7772), .A2(n7758), .ZN(n10424) );
  OR2_X1 U10046 ( .A1(n7995), .A2(n10424), .ZN(n7760) );
  INV_X1 U10047 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n10425) );
  OR2_X1 U10048 ( .A1(n8199), .A2(n10425), .ZN(n7759) );
  NAND4_X1 U10049 ( .A1(n7762), .A2(n7761), .A3(n7760), .A4(n7759), .ZN(n13041) );
  OR2_X1 U10050 ( .A1(n14811), .A2(n13041), .ZN(n7763) );
  NAND2_X1 U10051 ( .A1(n7764), .A2(n7765), .ZN(n7767) );
  XNOR2_X1 U10052 ( .A(n7767), .B(n7766), .ZN(n9397) );
  NAND2_X1 U10053 ( .A1(n9397), .A2(n6537), .ZN(n7771) );
  INV_X1 U10054 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n7768) );
  NAND2_X1 U10055 ( .A1(n8049), .A2(n7768), .ZN(n7786) );
  NAND2_X1 U10056 ( .A1(n7786), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7769) );
  XNOR2_X1 U10057 ( .A(n7769), .B(P2_IR_REG_11__SCAN_IN), .ZN(n10157) );
  AOI22_X1 U10058 ( .A1(n7908), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n7907), 
        .B2(n10157), .ZN(n7770) );
  NAND2_X1 U10059 ( .A1(n8040), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n7778) );
  INV_X1 U10060 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n9344) );
  OR2_X1 U10061 ( .A1(n8156), .A2(n9344), .ZN(n7777) );
  OR2_X1 U10062 ( .A1(n7772), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n7773) );
  NAND2_X1 U10063 ( .A1(n7795), .A2(n7773), .ZN(n10648) );
  OR2_X1 U10064 ( .A1(n8041), .A2(n10648), .ZN(n7776) );
  INV_X1 U10065 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n7774) );
  OR2_X1 U10066 ( .A1(n8157), .A2(n7774), .ZN(n7775) );
  NAND4_X1 U10067 ( .A1(n7778), .A2(n7777), .A3(n7776), .A4(n7775), .ZN(n13040) );
  INV_X1 U10068 ( .A(n13040), .ZN(n12024) );
  XNOR2_X1 U10069 ( .A(n12021), .B(n12024), .ZN(n12206) );
  NAND2_X1 U10070 ( .A1(n10652), .A2(n12206), .ZN(n7780) );
  NAND2_X1 U10071 ( .A1(n12021), .A2(n13040), .ZN(n7779) );
  NAND2_X1 U10072 ( .A1(n7780), .A2(n7779), .ZN(n10764) );
  NAND2_X1 U10073 ( .A1(n7764), .A2(n7781), .ZN(n7783) );
  AND2_X1 U10074 ( .A1(n7783), .A2(n7782), .ZN(n7785) );
  NAND2_X1 U10075 ( .A1(n9510), .A2(n6537), .ZN(n7793) );
  NOR2_X1 U10076 ( .A1(n7786), .A2(P2_IR_REG_11__SCAN_IN), .ZN(n7790) );
  INV_X1 U10077 ( .A(n7790), .ZN(n7787) );
  NAND2_X1 U10078 ( .A1(n7787), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7788) );
  MUX2_X1 U10079 ( .A(P2_IR_REG_31__SCAN_IN), .B(n7788), .S(
        P2_IR_REG_12__SCAN_IN), .Z(n7791) );
  INV_X1 U10080 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n7789) );
  NAND2_X1 U10081 ( .A1(n7790), .A2(n7789), .ZN(n7822) );
  NAND2_X1 U10082 ( .A1(n7791), .A2(n7822), .ZN(n14732) );
  INV_X1 U10083 ( .A(n14732), .ZN(n10159) );
  AOI22_X1 U10084 ( .A1(n7908), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n7907), 
        .B2(n10159), .ZN(n7792) );
  NAND2_X1 U10085 ( .A1(n8195), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n7801) );
  INV_X1 U10086 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n10774) );
  OR2_X1 U10087 ( .A1(n8199), .A2(n10774), .ZN(n7800) );
  NAND2_X1 U10088 ( .A1(n7795), .A2(n7794), .ZN(n7796) );
  NAND2_X1 U10089 ( .A1(n7813), .A2(n7796), .ZN(n10852) );
  OR2_X1 U10090 ( .A1(n7995), .A2(n10852), .ZN(n7799) );
  INV_X1 U10091 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n7797) );
  OR2_X1 U10092 ( .A1(n8157), .A2(n7797), .ZN(n7798) );
  NAND4_X1 U10093 ( .A1(n7801), .A2(n7800), .A3(n7799), .A4(n7798), .ZN(n13039) );
  AND2_X1 U10094 ( .A1(n14379), .A2(n13039), .ZN(n7803) );
  OR2_X1 U10095 ( .A1(n14379), .A2(n13039), .ZN(n7802) );
  NAND2_X1 U10096 ( .A1(n7764), .A2(n7804), .ZN(n7806) );
  AND2_X1 U10097 ( .A1(n7806), .A2(n7805), .ZN(n7808) );
  NAND2_X1 U10098 ( .A1(n9514), .A2(n6537), .ZN(n7811) );
  NAND2_X1 U10099 ( .A1(n7822), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7809) );
  XNOR2_X1 U10100 ( .A(n7809), .B(P2_IR_REG_13__SCAN_IN), .ZN(n10160) );
  AOI22_X1 U10101 ( .A1(n7908), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n7907), 
        .B2(n10160), .ZN(n7810) );
  NAND2_X2 U10102 ( .A1(n7811), .A2(n7810), .ZN(n12032) );
  NAND2_X1 U10103 ( .A1(n7596), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n7818) );
  NAND2_X1 U10104 ( .A1(n7813), .A2(n7812), .ZN(n7814) );
  NAND2_X1 U10105 ( .A1(n7827), .A2(n7814), .ZN(n10992) );
  OR2_X1 U10106 ( .A1(n7995), .A2(n10992), .ZN(n7817) );
  INV_X1 U10107 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n10153) );
  OR2_X1 U10108 ( .A1(n8156), .A2(n10153), .ZN(n7816) );
  INV_X1 U10109 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n10993) );
  OR2_X1 U10110 ( .A1(n8199), .A2(n10993), .ZN(n7815) );
  NAND4_X1 U10111 ( .A1(n7818), .A2(n7817), .A3(n7816), .A4(n7815), .ZN(n14335) );
  NOR2_X1 U10112 ( .A1(n12032), .A2(n14335), .ZN(n7819) );
  INV_X1 U10113 ( .A(n12032), .ZN(n14374) );
  INV_X1 U10114 ( .A(n14335), .ZN(n12034) );
  NAND2_X1 U10115 ( .A1(n9593), .A2(n6537), .ZN(n7825) );
  OR2_X1 U10116 ( .A1(n7822), .A2(P2_IR_REG_13__SCAN_IN), .ZN(n7839) );
  NAND2_X1 U10117 ( .A1(n7839), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7823) );
  XNOR2_X1 U10118 ( .A(n7823), .B(P2_IR_REG_14__SCAN_IN), .ZN(n10163) );
  AOI22_X1 U10119 ( .A1(n7908), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n10163), 
        .B2(n7907), .ZN(n7824) );
  AND2_X1 U10120 ( .A1(n7827), .A2(n7826), .ZN(n7828) );
  OR2_X1 U10121 ( .A1(n7828), .A2(n7843), .ZN(n14347) );
  INV_X1 U10122 ( .A(n14347), .ZN(n14353) );
  NAND2_X1 U10123 ( .A1(n14353), .A2(n7940), .ZN(n7834) );
  NAND2_X1 U10124 ( .A1(n8195), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n7833) );
  INV_X1 U10125 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n7829) );
  OR2_X1 U10126 ( .A1(n8157), .A2(n7829), .ZN(n7832) );
  INV_X1 U10127 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n7830) );
  OR2_X1 U10128 ( .A1(n8199), .A2(n7830), .ZN(n7831) );
  NAND4_X1 U10129 ( .A1(n7834), .A2(n7833), .A3(n7832), .A4(n7831), .ZN(n13038) );
  AND2_X1 U10130 ( .A1(n14356), .A2(n13038), .ZN(n7836) );
  OR2_X1 U10131 ( .A1(n14356), .A2(n13038), .ZN(n7835) );
  OAI21_X2 U10132 ( .B1(n14357), .B2(n7836), .A(n7835), .ZN(n11342) );
  XNOR2_X1 U10133 ( .A(n7838), .B(n7837), .ZN(n9784) );
  NAND2_X1 U10134 ( .A1(n9784), .A2(n6537), .ZN(n7842) );
  OAI21_X1 U10135 ( .B1(n7839), .B2(P2_IR_REG_14__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n7840) );
  XNOR2_X1 U10136 ( .A(n7840), .B(P2_IR_REG_15__SCAN_IN), .ZN(n14753) );
  AOI22_X1 U10137 ( .A1(n14753), .A2(n7907), .B1(n7908), .B2(
        P1_DATAO_REG_15__SCAN_IN), .ZN(n7841) );
  OR2_X1 U10138 ( .A1(n7843), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n7844) );
  NAND2_X1 U10139 ( .A1(n7864), .A2(n7844), .ZN(n11345) );
  NAND2_X1 U10140 ( .A1(n7596), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n7845) );
  OAI21_X1 U10141 ( .B1(n11345), .B2(n7995), .A(n7845), .ZN(n7849) );
  INV_X1 U10142 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n7847) );
  INV_X1 U10143 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n7846) );
  OAI22_X1 U10144 ( .A1(n8199), .A2(n7847), .B1(n8156), .B2(n7846), .ZN(n7848)
         );
  XNOR2_X1 U10145 ( .A(n12050), .B(n14337), .ZN(n12210) );
  INV_X1 U10146 ( .A(n12210), .ZN(n11341) );
  OR2_X1 U10147 ( .A1(n12050), .A2(n14337), .ZN(n7850) );
  XNOR2_X1 U10148 ( .A(n7852), .B(n7851), .ZN(n9914) );
  NAND2_X1 U10149 ( .A1(n9914), .A2(n6537), .ZN(n7862) );
  INV_X1 U10150 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n7853) );
  AND4_X1 U10151 ( .A1(n7856), .A2(n7855), .A3(n7854), .A4(n7853), .ZN(n7857)
         );
  NAND2_X1 U10152 ( .A1(n8049), .A2(n7857), .ZN(n7859) );
  NAND2_X1 U10153 ( .A1(n7859), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7858) );
  MUX2_X1 U10154 ( .A(P2_IR_REG_31__SCAN_IN), .B(n7858), .S(
        P2_IR_REG_16__SCAN_IN), .Z(n7860) );
  INV_X1 U10155 ( .A(n7878), .ZN(n7875) );
  AND2_X1 U10156 ( .A1(n7860), .A2(n7875), .ZN(n10743) );
  AOI22_X1 U10157 ( .A1(n7908), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n7907), 
        .B2(n10743), .ZN(n7861) );
  NAND2_X1 U10158 ( .A1(n7864), .A2(n7863), .ZN(n7865) );
  NAND2_X1 U10159 ( .A1(n7882), .A2(n7865), .ZN(n11381) );
  INV_X1 U10160 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n11409) );
  OR2_X1 U10161 ( .A1(n8199), .A2(n11409), .ZN(n7867) );
  INV_X1 U10162 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n15259) );
  OR2_X1 U10163 ( .A1(n8156), .A2(n15259), .ZN(n7866) );
  AND2_X1 U10164 ( .A1(n7867), .A2(n7866), .ZN(n7869) );
  NAND2_X1 U10165 ( .A1(n7596), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n7868) );
  OAI211_X1 U10166 ( .C1(n11381), .C2(n7995), .A(n7869), .B(n7868), .ZN(n13037) );
  XNOR2_X1 U10167 ( .A(n13426), .B(n13037), .ZN(n12211) );
  NAND2_X1 U10168 ( .A1(n13426), .A2(n13037), .ZN(n7871) );
  NAND2_X1 U10169 ( .A1(n11412), .A2(n7871), .ZN(n11447) );
  XNOR2_X1 U10170 ( .A(n7872), .B(SI_17_), .ZN(n7873) );
  XNOR2_X1 U10171 ( .A(n7874), .B(n7873), .ZN(n9958) );
  NAND2_X1 U10172 ( .A1(n9958), .A2(n6537), .ZN(n7881) );
  NAND2_X1 U10173 ( .A1(n7875), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7876) );
  MUX2_X1 U10174 ( .A(P2_IR_REG_31__SCAN_IN), .B(n7876), .S(
        P2_IR_REG_17__SCAN_IN), .Z(n7879) );
  INV_X1 U10175 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n7877) );
  NAND2_X1 U10176 ( .A1(n7878), .A2(n7877), .ZN(n7905) );
  NAND2_X1 U10177 ( .A1(n7879), .A2(n7905), .ZN(n13124) );
  INV_X1 U10178 ( .A(n13124), .ZN(n11361) );
  AOI22_X1 U10179 ( .A1(n7908), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n7907), 
        .B2(n11361), .ZN(n7880) );
  AND2_X1 U10180 ( .A1(n7882), .A2(n15294), .ZN(n7883) );
  OR2_X1 U10181 ( .A1(n7883), .A2(n7890), .ZN(n11466) );
  AOI22_X1 U10182 ( .A1(n8040), .A2(P2_REG2_REG_17__SCAN_IN), .B1(n8195), .B2(
        P2_REG1_REG_17__SCAN_IN), .ZN(n7885) );
  NAND2_X1 U10183 ( .A1(n7596), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n7884) );
  OAI211_X1 U10184 ( .C1(n11466), .C2(n7995), .A(n7885), .B(n7884), .ZN(n13036) );
  XNOR2_X1 U10185 ( .A(n12065), .B(n13036), .ZN(n12213) );
  INV_X1 U10186 ( .A(n12213), .ZN(n11446) );
  NAND2_X1 U10187 ( .A1(n12065), .A2(n13036), .ZN(n7886) );
  XNOR2_X1 U10188 ( .A(n7895), .B(n7896), .ZN(n10460) );
  NAND2_X1 U10189 ( .A1(n10460), .A2(n6537), .ZN(n7889) );
  NAND2_X1 U10190 ( .A1(n7905), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7887) );
  XNOR2_X1 U10191 ( .A(n7887), .B(P2_IR_REG_18__SCAN_IN), .ZN(n13135) );
  AOI22_X1 U10192 ( .A1(n7908), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n7907), 
        .B2(n13135), .ZN(n7888) );
  NOR2_X1 U10193 ( .A1(n7890), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n7891) );
  OR2_X1 U10194 ( .A1(n7910), .A2(n7891), .ZN(n13324) );
  AOI22_X1 U10195 ( .A1(n8195), .A2(P2_REG1_REG_18__SCAN_IN), .B1(n7596), .B2(
        P2_REG0_REG_18__SCAN_IN), .ZN(n7893) );
  NAND2_X1 U10196 ( .A1(n8040), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n7892) );
  OAI211_X1 U10197 ( .C1(n13324), .C2(n7995), .A(n7893), .B(n7892), .ZN(n13035) );
  INV_X1 U10198 ( .A(n13035), .ZN(n8132) );
  XNOR2_X1 U10199 ( .A(n6523), .B(n8132), .ZN(n13334) );
  OR2_X1 U10200 ( .A1(n6523), .A2(n13035), .ZN(n7894) );
  INV_X1 U10201 ( .A(n7895), .ZN(n7897) );
  NAND2_X1 U10202 ( .A1(n7897), .A2(n7896), .ZN(n7900) );
  NAND2_X1 U10203 ( .A1(n7898), .A2(SI_18_), .ZN(n7899) );
  NAND2_X1 U10204 ( .A1(n7900), .A2(n7899), .ZN(n7904) );
  NAND2_X1 U10205 ( .A1(n7902), .A2(n7901), .ZN(n7903) );
  XNOR2_X2 U10206 ( .A(n7904), .B(n7903), .ZN(n10656) );
  AOI22_X1 U10207 ( .A1(n7908), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n13167), 
        .B2(n7907), .ZN(n7909) );
  NOR2_X1 U10208 ( .A1(n7910), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n7911) );
  OR2_X1 U10209 ( .A1(n7926), .A2(n7911), .ZN(n13313) );
  INV_X1 U10210 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n13312) );
  NAND2_X1 U10211 ( .A1(n8195), .A2(P2_REG1_REG_19__SCAN_IN), .ZN(n7914) );
  INV_X1 U10212 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n7912) );
  OR2_X1 U10213 ( .A1(n8157), .A2(n7912), .ZN(n7913) );
  OAI211_X1 U10214 ( .C1(n8199), .C2(n13312), .A(n7914), .B(n7913), .ZN(n7915)
         );
  INV_X1 U10215 ( .A(n7915), .ZN(n7916) );
  OAI21_X1 U10216 ( .B1(n13313), .B2(n7995), .A(n7916), .ZN(n13034) );
  NOR2_X1 U10217 ( .A1(n13406), .A2(n13034), .ZN(n7918) );
  NAND2_X1 U10218 ( .A1(n13406), .A2(n13034), .ZN(n7917) );
  NAND2_X1 U10219 ( .A1(n7920), .A2(n7919), .ZN(n7923) );
  XNOR2_X1 U10220 ( .A(n7921), .B(SI_20_), .ZN(n7922) );
  NAND2_X1 U10221 ( .A1(n10458), .A2(n6537), .ZN(n7925) );
  OR2_X1 U10222 ( .A1(n8193), .A2(n10497), .ZN(n7924) );
  NOR2_X1 U10223 ( .A1(n7926), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n7927) );
  OR2_X1 U10224 ( .A1(n7938), .A2(n7927), .ZN(n13295) );
  INV_X1 U10225 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n13294) );
  NAND2_X1 U10226 ( .A1(n7596), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n7929) );
  NAND2_X1 U10227 ( .A1(n8195), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n7928) );
  OAI211_X1 U10228 ( .C1(n8199), .C2(n13294), .A(n7929), .B(n7928), .ZN(n7930)
         );
  INV_X1 U10229 ( .A(n7930), .ZN(n7931) );
  OAI21_X1 U10230 ( .B1(n13295), .B2(n7995), .A(n7931), .ZN(n13033) );
  AND2_X1 U10231 ( .A1(n13402), .A2(n13033), .ZN(n7933) );
  OR2_X1 U10232 ( .A1(n13402), .A2(n13033), .ZN(n7932) );
  OAI21_X2 U10233 ( .B1(n13285), .B2(n7933), .A(n7932), .ZN(n13268) );
  XNOR2_X1 U10234 ( .A(n7935), .B(n7934), .ZN(n10667) );
  NAND2_X1 U10235 ( .A1(n10667), .A2(n6537), .ZN(n7937) );
  INV_X1 U10236 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n11911) );
  OR2_X1 U10237 ( .A1(n8193), .A2(n11911), .ZN(n7936) );
  OR2_X1 U10238 ( .A1(n7938), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n7939) );
  AND2_X1 U10239 ( .A1(n7952), .A2(n7939), .ZN(n13277) );
  NAND2_X1 U10240 ( .A1(n13277), .A2(n7940), .ZN(n7945) );
  INV_X1 U10241 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n15233) );
  NAND2_X1 U10242 ( .A1(n8040), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n7942) );
  NAND2_X1 U10243 ( .A1(n8195), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n7941) );
  OAI211_X1 U10244 ( .C1(n15233), .C2(n8157), .A(n7942), .B(n7941), .ZN(n7943)
         );
  INV_X1 U10245 ( .A(n7943), .ZN(n7944) );
  NAND2_X1 U10246 ( .A1(n7945), .A2(n7944), .ZN(n13032) );
  INV_X1 U10247 ( .A(n13032), .ZN(n8140) );
  XNOR2_X1 U10248 ( .A(n13459), .B(n8140), .ZN(n13270) );
  NAND2_X1 U10249 ( .A1(n13268), .A2(n13270), .ZN(n7947) );
  OR2_X1 U10250 ( .A1(n13459), .A2(n13032), .ZN(n7946) );
  XNOR2_X1 U10251 ( .A(n7948), .B(n7949), .ZN(n10878) );
  NAND2_X1 U10252 ( .A1(n10878), .A2(n6537), .ZN(n7951) );
  INV_X1 U10253 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n10880) );
  OR2_X1 U10254 ( .A1(n8193), .A2(n10880), .ZN(n7950) );
  NAND2_X1 U10255 ( .A1(n7952), .A2(n12998), .ZN(n7954) );
  INV_X1 U10256 ( .A(n7967), .ZN(n7953) );
  NAND2_X1 U10257 ( .A1(n7954), .A2(n7953), .ZN(n13261) );
  OR2_X1 U10258 ( .A1(n13261), .A2(n7995), .ZN(n7959) );
  INV_X1 U10259 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n13260) );
  NAND2_X1 U10260 ( .A1(n7596), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n7956) );
  INV_X1 U10261 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n15345) );
  OR2_X1 U10262 ( .A1(n8156), .A2(n15345), .ZN(n7955) );
  OAI211_X1 U10263 ( .C1(n8199), .C2(n13260), .A(n7956), .B(n7955), .ZN(n7957)
         );
  INV_X1 U10264 ( .A(n7957), .ZN(n7958) );
  NAND2_X1 U10265 ( .A1(n7959), .A2(n7958), .ZN(n13031) );
  XNOR2_X1 U10266 ( .A(n13263), .B(n13031), .ZN(n13250) );
  NAND2_X1 U10267 ( .A1(n13263), .A2(n13031), .ZN(n7961) );
  XNOR2_X1 U10268 ( .A(n7962), .B(n6694), .ZN(n11010) );
  NAND2_X1 U10269 ( .A1(n11010), .A2(n6537), .ZN(n7964) );
  OR2_X1 U10270 ( .A1(n8193), .A2(n11013), .ZN(n7963) );
  NAND2_X1 U10271 ( .A1(n8040), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n7972) );
  INV_X1 U10272 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n7965) );
  OR2_X1 U10273 ( .A1(n8156), .A2(n7965), .ZN(n7971) );
  OAI21_X1 U10274 ( .B1(P2_REG3_REG_23__SCAN_IN), .B2(n7967), .A(n7966), .ZN(
        n12926) );
  OR2_X1 U10275 ( .A1(n8041), .A2(n12926), .ZN(n7970) );
  INV_X1 U10276 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n7968) );
  OR2_X1 U10277 ( .A1(n8157), .A2(n7968), .ZN(n7969) );
  NAND4_X1 U10278 ( .A1(n7972), .A2(n7971), .A3(n7970), .A4(n7969), .ZN(n13030) );
  NAND2_X1 U10279 ( .A1(n13385), .A2(n13030), .ZN(n12216) );
  OR2_X1 U10280 ( .A1(n13385), .A2(n13030), .ZN(n12217) );
  INV_X1 U10281 ( .A(n7974), .ZN(n7975) );
  XNOR2_X1 U10282 ( .A(n7976), .B(n7975), .ZN(n11224) );
  NAND2_X1 U10283 ( .A1(n11224), .A2(n6537), .ZN(n7978) );
  OR2_X1 U10284 ( .A1(n8193), .A2(n11228), .ZN(n7977) );
  NAND2_X1 U10285 ( .A1(n8195), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n7986) );
  INV_X1 U10286 ( .A(P2_REG2_REG_24__SCAN_IN), .ZN(n7979) );
  OR2_X1 U10287 ( .A1(n8199), .A2(n7979), .ZN(n7985) );
  INV_X1 U10288 ( .A(n7980), .ZN(n7992) );
  OAI21_X1 U10289 ( .B1(P2_REG3_REG_24__SCAN_IN), .B2(n7981), .A(n7992), .ZN(
        n13231) );
  OR2_X1 U10290 ( .A1(n7995), .A2(n13231), .ZN(n7984) );
  INV_X1 U10291 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n7982) );
  OR2_X1 U10292 ( .A1(n8157), .A2(n7982), .ZN(n7983) );
  NAND4_X1 U10293 ( .A1(n7986), .A2(n7985), .A3(n7984), .A4(n7983), .ZN(n13029) );
  XNOR2_X1 U10294 ( .A(n13233), .B(n13029), .ZN(n13224) );
  INV_X1 U10295 ( .A(n13233), .ZN(n13451) );
  INV_X1 U10296 ( .A(n13029), .ZN(n8146) );
  NAND2_X1 U10297 ( .A1(n11256), .A2(n6537), .ZN(n7990) );
  OR2_X1 U10298 ( .A1(n8193), .A2(n15170), .ZN(n7989) );
  NAND2_X1 U10299 ( .A1(n8195), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n8000) );
  INV_X1 U10300 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n7991) );
  OR2_X1 U10301 ( .A1(n8157), .A2(n7991), .ZN(n7999) );
  INV_X1 U10302 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n15148) );
  NAND2_X1 U10303 ( .A1(n15148), .A2(n7992), .ZN(n7993) );
  NAND2_X1 U10304 ( .A1(n7994), .A2(n7993), .ZN(n12967) );
  OR2_X1 U10305 ( .A1(n7995), .A2(n12967), .ZN(n7998) );
  INV_X1 U10306 ( .A(P2_REG2_REG_25__SCAN_IN), .ZN(n7996) );
  OR2_X1 U10307 ( .A1(n8199), .A2(n7996), .ZN(n7997) );
  NAND4_X1 U10308 ( .A1(n8000), .A2(n7999), .A3(n7998), .A4(n7997), .ZN(n13028) );
  AND2_X1 U10309 ( .A1(n13375), .A2(n13028), .ZN(n8001) );
  INV_X1 U10310 ( .A(SI_26_), .ZN(n11550) );
  MUX2_X1 U10311 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(P1_DATAO_REG_27__SCAN_IN), 
        .S(n9727), .Z(n8015) );
  INV_X1 U10312 ( .A(n8015), .ZN(n8005) );
  XNOR2_X1 U10313 ( .A(n8005), .B(SI_27_), .ZN(n8006) );
  NAND2_X1 U10314 ( .A1(n13483), .A2(n6537), .ZN(n8008) );
  INV_X1 U10315 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n13485) );
  OR2_X1 U10316 ( .A1(n8193), .A2(n13485), .ZN(n8007) );
  NAND2_X1 U10317 ( .A1(n8040), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n8012) );
  INV_X1 U10318 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n13366) );
  OR2_X1 U10319 ( .A1(n8156), .A2(n13366), .ZN(n8011) );
  INV_X1 U10320 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n15265) );
  XNOR2_X1 U10321 ( .A(n8024), .B(n15265), .ZN(n12920) );
  OR2_X1 U10322 ( .A1(n7995), .A2(n12920), .ZN(n8010) );
  INV_X1 U10323 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n13440) );
  OR2_X1 U10324 ( .A1(n8157), .A2(n13440), .ZN(n8009) );
  NAND4_X1 U10325 ( .A1(n8012), .A2(n8011), .A3(n8010), .A4(n8009), .ZN(n13026) );
  INV_X1 U10326 ( .A(n13026), .ZN(n12947) );
  OAI22_X1 U10327 ( .A1(n13179), .A2(n13181), .B1(n13442), .B2(n12947), .ZN(
        n13162) );
  NOR2_X1 U10328 ( .A1(n8015), .A2(SI_27_), .ZN(n8013) );
  NAND2_X1 U10329 ( .A1(n8015), .A2(SI_27_), .ZN(n8016) );
  INV_X1 U10330 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n11639) );
  INV_X1 U10331 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n11576) );
  MUX2_X1 U10332 ( .A(n11639), .B(n11576), .S(n9727), .Z(n8018) );
  INV_X1 U10333 ( .A(SI_28_), .ZN(n12243) );
  NAND2_X1 U10334 ( .A1(n8018), .A2(n12243), .ZN(n8034) );
  INV_X1 U10335 ( .A(n8018), .ZN(n8019) );
  NAND2_X1 U10336 ( .A1(n8019), .A2(SI_28_), .ZN(n8020) );
  NAND2_X1 U10337 ( .A1(n8034), .A2(n8020), .ZN(n8035) );
  NAND2_X1 U10338 ( .A1(n11638), .A2(n6537), .ZN(n8022) );
  OR2_X1 U10339 ( .A1(n8193), .A2(n11576), .ZN(n8021) );
  NAND2_X1 U10340 ( .A1(n8040), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n8031) );
  INV_X1 U10341 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n15288) );
  OR2_X1 U10342 ( .A1(n8156), .A2(n15288), .ZN(n8030) );
  INV_X1 U10343 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n8023) );
  OAI21_X1 U10344 ( .B1(n8024), .B2(n15265), .A(n8023), .ZN(n8027) );
  INV_X1 U10345 ( .A(n8024), .ZN(n8026) );
  AND2_X1 U10346 ( .A1(P2_REG3_REG_27__SCAN_IN), .A2(P2_REG3_REG_28__SCAN_IN), 
        .ZN(n8025) );
  NAND2_X1 U10347 ( .A1(n8026), .A2(n8025), .ZN(n8171) );
  NAND2_X1 U10348 ( .A1(n8027), .A2(n8171), .ZN(n13166) );
  INV_X1 U10349 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n15280) );
  OR2_X1 U10350 ( .A1(n8157), .A2(n15280), .ZN(n8028) );
  NAND4_X1 U10351 ( .A1(n8031), .A2(n8030), .A3(n8029), .A4(n8028), .ZN(n13025) );
  INV_X1 U10352 ( .A(n13025), .ZN(n8032) );
  NAND2_X1 U10353 ( .A1(n13356), .A2(n8032), .ZN(n8033) );
  INV_X1 U10354 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n11644) );
  INV_X1 U10355 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n13477) );
  MUX2_X1 U10356 ( .A(n11644), .B(n13477), .S(n9727), .Z(n8179) );
  XNOR2_X1 U10357 ( .A(n8179), .B(SI_29_), .ZN(n8177) );
  NAND2_X1 U10358 ( .A1(n11636), .A2(n6537), .ZN(n8039) );
  OR2_X1 U10359 ( .A1(n8193), .A2(n13477), .ZN(n8038) );
  NAND2_X1 U10360 ( .A1(n8195), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n8046) );
  NAND2_X1 U10361 ( .A1(n8040), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n8045) );
  OR2_X1 U10362 ( .A1(n8041), .A2(n8171), .ZN(n8044) );
  INV_X1 U10363 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n8042) );
  OR2_X1 U10364 ( .A1(n8157), .A2(n8042), .ZN(n8043) );
  NAND4_X1 U10365 ( .A1(n8046), .A2(n8045), .A3(n8044), .A4(n8043), .ZN(n13024) );
  INV_X1 U10366 ( .A(n13024), .ZN(n12949) );
  INV_X1 U10367 ( .A(n12224), .ZN(n8047) );
  XNOR2_X1 U10368 ( .A(n8048), .B(n8047), .ZN(n13354) );
  NOR2_X1 U10369 ( .A1(n8060), .A2(n13473), .ZN(n8053) );
  INV_X1 U10370 ( .A(n8063), .ZN(n8054) );
  NAND2_X2 U10371 ( .A1(n8056), .A2(n8055), .ZN(n8092) );
  NAND2_X1 U10372 ( .A1(n11925), .A2(n8092), .ZN(n9431) );
  INV_X1 U10373 ( .A(n8057), .ZN(n8058) );
  NAND2_X1 U10374 ( .A1(n8058), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8059) );
  AND2_X2 U10375 ( .A1(n8062), .A2(n8061), .ZN(n12230) );
  INV_X4 U10376 ( .A(n9550), .ZN(n13326) );
  INV_X1 U10377 ( .A(n11921), .ZN(n13144) );
  OAI21_X1 U10378 ( .B1(n8063), .B2(P2_IR_REG_22__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n8065) );
  XNOR2_X1 U10379 ( .A(n8065), .B(n8064), .ZN(n11011) );
  NAND2_X1 U10380 ( .A1(n8049), .A2(n6555), .ZN(n8068) );
  NAND2_X1 U10381 ( .A1(n8070), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8066) );
  MUX2_X1 U10382 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8066), .S(
        P2_IR_REG_25__SCAN_IN), .Z(n8067) );
  NAND2_X1 U10383 ( .A1(n8067), .A2(n6577), .ZN(n11257) );
  INV_X1 U10384 ( .A(n11257), .ZN(n8074) );
  NAND2_X1 U10385 ( .A1(n8068), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8069) );
  MUX2_X1 U10386 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8069), .S(
        P2_IR_REG_24__SCAN_IN), .Z(n8071) );
  NAND2_X1 U10387 ( .A1(n8071), .A2(n8070), .ZN(n11226) );
  NAND2_X1 U10388 ( .A1(n6577), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8072) );
  XNOR2_X1 U10389 ( .A(n8072), .B(n7460), .ZN(n13488) );
  NOR2_X1 U10390 ( .A1(n11226), .A2(n13488), .ZN(n8073) );
  NAND2_X1 U10391 ( .A1(n8074), .A2(n8073), .ZN(n9553) );
  INV_X1 U10392 ( .A(n9421), .ZN(n8161) );
  NAND2_X1 U10393 ( .A1(n8161), .A2(n12180), .ZN(n9554) );
  NAND2_X1 U10394 ( .A1(n9554), .A2(n14773), .ZN(n9433) );
  INV_X1 U10395 ( .A(P2_B_REG_SCAN_IN), .ZN(n8162) );
  XOR2_X1 U10396 ( .A(n11226), .B(n8162), .Z(n8076) );
  INV_X1 U10397 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n14768) );
  NAND2_X1 U10398 ( .A1(n14765), .A2(n14768), .ZN(n8078) );
  NAND2_X1 U10399 ( .A1(n11226), .A2(n13488), .ZN(n8077) );
  NAND2_X1 U10400 ( .A1(n8078), .A2(n8077), .ZN(n14769) );
  INV_X1 U10401 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n14771) );
  NAND2_X1 U10402 ( .A1(n14765), .A2(n14771), .ZN(n8080) );
  NAND2_X1 U10403 ( .A1(n11257), .A2(n13488), .ZN(n8079) );
  NOR4_X1 U10404 ( .A1(P2_D_REG_14__SCAN_IN), .A2(P2_D_REG_16__SCAN_IN), .A3(
        P2_D_REG_17__SCAN_IN), .A4(P2_D_REG_19__SCAN_IN), .ZN(n8084) );
  NOR4_X1 U10405 ( .A1(P2_D_REG_11__SCAN_IN), .A2(P2_D_REG_12__SCAN_IN), .A3(
        P2_D_REG_15__SCAN_IN), .A4(P2_D_REG_13__SCAN_IN), .ZN(n8083) );
  NOR4_X1 U10406 ( .A1(P2_D_REG_24__SCAN_IN), .A2(P2_D_REG_26__SCAN_IN), .A3(
        P2_D_REG_27__SCAN_IN), .A4(P2_D_REG_29__SCAN_IN), .ZN(n8082) );
  NOR4_X1 U10407 ( .A1(P2_D_REG_20__SCAN_IN), .A2(P2_D_REG_23__SCAN_IN), .A3(
        P2_D_REG_21__SCAN_IN), .A4(P2_D_REG_22__SCAN_IN), .ZN(n8081) );
  NAND4_X1 U10408 ( .A1(n8084), .A2(n8083), .A3(n8082), .A4(n8081), .ZN(n8089)
         );
  NOR2_X1 U10409 ( .A1(P2_D_REG_25__SCAN_IN), .A2(P2_D_REG_28__SCAN_IN), .ZN(
        n15104) );
  NOR4_X1 U10410 ( .A1(P2_D_REG_30__SCAN_IN), .A2(P2_D_REG_31__SCAN_IN), .A3(
        P2_D_REG_10__SCAN_IN), .A4(P2_D_REG_18__SCAN_IN), .ZN(n8087) );
  NOR4_X1 U10411 ( .A1(P2_D_REG_5__SCAN_IN), .A2(P2_D_REG_6__SCAN_IN), .A3(
        P2_D_REG_8__SCAN_IN), .A4(P2_D_REG_9__SCAN_IN), .ZN(n8086) );
  NOR4_X1 U10412 ( .A1(P2_D_REG_7__SCAN_IN), .A2(P2_D_REG_2__SCAN_IN), .A3(
        P2_D_REG_3__SCAN_IN), .A4(P2_D_REG_4__SCAN_IN), .ZN(n8085) );
  NAND4_X1 U10413 ( .A1(n15104), .A2(n8087), .A3(n8086), .A4(n8085), .ZN(n8088) );
  OAI21_X1 U10414 ( .B1(n8089), .B2(n8088), .A(n14765), .ZN(n9412) );
  AND2_X1 U10415 ( .A1(n9409), .A2(n9412), .ZN(n8090) );
  NAND2_X1 U10416 ( .A1(n14769), .A2(n8090), .ZN(n8091) );
  INV_X2 U10417 ( .A(n14367), .ZN(n13281) );
  NAND2_X1 U10418 ( .A1(n6538), .A2(n13144), .ZN(n8095) );
  AND2_X1 U10419 ( .A1(n6528), .A2(n8095), .ZN(n8096) );
  INV_X1 U10420 ( .A(n11928), .ZN(n9419) );
  NAND2_X1 U10421 ( .A1(n9419), .A2(n11935), .ZN(n9546) );
  INV_X1 U10422 ( .A(n9546), .ZN(n8097) );
  NAND2_X1 U10423 ( .A1(n8097), .A2(n12192), .ZN(n9544) );
  NAND2_X1 U10424 ( .A1(n8098), .A2(n11932), .ZN(n8099) );
  NAND2_X1 U10425 ( .A1(n9535), .A2(n12191), .ZN(n8102) );
  NAND2_X1 U10426 ( .A1(n8100), .A2(n6524), .ZN(n8101) );
  NAND2_X1 U10427 ( .A1(n8102), .A2(n8101), .ZN(n9519) );
  INV_X1 U10428 ( .A(n12194), .ZN(n8103) );
  NAND2_X1 U10429 ( .A1(n9519), .A2(n8103), .ZN(n8106) );
  NAND2_X1 U10430 ( .A1(n11965), .A2(n8104), .ZN(n8105) );
  NAND2_X1 U10431 ( .A1(n8106), .A2(n8105), .ZN(n9570) );
  NAND2_X1 U10432 ( .A1(n9570), .A2(n12195), .ZN(n8108) );
  NAND2_X1 U10433 ( .A1(n11973), .A2(n11975), .ZN(n8107) );
  NAND2_X1 U10434 ( .A1(n8108), .A2(n8107), .ZN(n10168) );
  INV_X1 U10435 ( .A(n13047), .ZN(n8110) );
  AND2_X1 U10436 ( .A1(n11980), .A2(n8110), .ZN(n8109) );
  OR2_X1 U10437 ( .A1(n11980), .A2(n8110), .ZN(n8111) );
  NAND2_X1 U10438 ( .A1(n10141), .A2(n8112), .ZN(n10179) );
  NAND2_X1 U10439 ( .A1(n10187), .A2(n13045), .ZN(n8113) );
  NAND2_X1 U10440 ( .A1(n10179), .A2(n8113), .ZN(n8115) );
  NAND2_X1 U10441 ( .A1(n14788), .A2(n11992), .ZN(n8114) );
  NAND2_X1 U10442 ( .A1(n8115), .A2(n8114), .ZN(n10464) );
  INV_X1 U10443 ( .A(n13044), .ZN(n10248) );
  NAND2_X1 U10444 ( .A1(n14795), .A2(n10248), .ZN(n8116) );
  INV_X1 U10445 ( .A(n13042), .ZN(n8117) );
  OR2_X1 U10446 ( .A1(n12008), .A2(n8117), .ZN(n8118) );
  INV_X1 U10447 ( .A(n13041), .ZN(n10247) );
  NAND2_X1 U10448 ( .A1(n14811), .A2(n10247), .ZN(n8119) );
  NAND2_X1 U10449 ( .A1(n10416), .A2(n8119), .ZN(n8121) );
  OR2_X1 U10450 ( .A1(n14811), .A2(n10247), .ZN(n8120) );
  INV_X1 U10451 ( .A(n13039), .ZN(n8122) );
  XNOR2_X1 U10452 ( .A(n14379), .B(n8122), .ZN(n12207) );
  NAND2_X1 U10453 ( .A1(n12032), .A2(n12034), .ZN(n10983) );
  NAND2_X1 U10454 ( .A1(n10985), .A2(n10983), .ZN(n8123) );
  OR2_X1 U10455 ( .A1(n12032), .A2(n12034), .ZN(n10984) );
  INV_X1 U10456 ( .A(n13038), .ZN(n8124) );
  XNOR2_X1 U10457 ( .A(n14356), .B(n8124), .ZN(n14358) );
  INV_X1 U10458 ( .A(n14337), .ZN(n8126) );
  INV_X1 U10459 ( .A(n13037), .ZN(n12059) );
  NAND2_X1 U10460 ( .A1(n13426), .A2(n12059), .ZN(n8127) );
  NAND2_X1 U10461 ( .A1(n11401), .A2(n8127), .ZN(n8129) );
  OR2_X1 U10462 ( .A1(n13426), .A2(n12059), .ZN(n8128) );
  INV_X1 U10463 ( .A(n13036), .ZN(n8130) );
  OR2_X1 U10464 ( .A1(n12065), .A2(n8130), .ZN(n8131) );
  NAND2_X1 U10465 ( .A1(n6523), .A2(n8132), .ZN(n8133) );
  INV_X1 U10466 ( .A(n13034), .ZN(n12189) );
  AND2_X1 U10467 ( .A1(n12189), .A2(n13406), .ZN(n8135) );
  INV_X1 U10468 ( .A(n13033), .ZN(n8136) );
  NAND2_X1 U10469 ( .A1(n13402), .A2(n8136), .ZN(n13269) );
  OR2_X1 U10470 ( .A1(n13402), .A2(n8136), .ZN(n8137) );
  NAND2_X1 U10471 ( .A1(n13269), .A2(n8137), .ZN(n13289) );
  NAND2_X1 U10472 ( .A1(n13286), .A2(n13269), .ZN(n8139) );
  INV_X1 U10473 ( .A(n13270), .ZN(n8138) );
  NAND2_X1 U10474 ( .A1(n13459), .A2(n8140), .ZN(n8141) );
  INV_X1 U10475 ( .A(n13031), .ZN(n8142) );
  OR2_X1 U10476 ( .A1(n13263), .A2(n8142), .ZN(n8143) );
  INV_X1 U10477 ( .A(n13030), .ZN(n8144) );
  NOR2_X1 U10478 ( .A1(n13385), .A2(n8144), .ZN(n8145) );
  INV_X1 U10479 ( .A(n13385), .ZN(n13247) );
  INV_X1 U10480 ( .A(n13028), .ZN(n8147) );
  XNOR2_X1 U10481 ( .A(n13375), .B(n8147), .ZN(n13211) );
  INV_X1 U10482 ( .A(n13211), .ZN(n8149) );
  AND2_X1 U10483 ( .A1(n13375), .A2(n8147), .ZN(n8148) );
  OR2_X1 U10484 ( .A1(n13205), .A2(n8150), .ZN(n12188) );
  NAND2_X1 U10485 ( .A1(n13205), .A2(n8150), .ZN(n12187) );
  INV_X1 U10486 ( .A(n13161), .ZN(n13170) );
  NAND2_X1 U10487 ( .A1(n13187), .A2(n12947), .ZN(n13171) );
  NAND2_X1 U10488 ( .A1(n13169), .A2(n8151), .ZN(n8152) );
  XNOR2_X1 U10489 ( .A(n8152), .B(n12224), .ZN(n8166) );
  NAND2_X1 U10490 ( .A1(n11921), .A2(n8153), .ZN(n12152) );
  INV_X1 U10491 ( .A(n12230), .ZN(n12183) );
  OR2_X1 U10492 ( .A1(n8092), .A2(n12183), .ZN(n8154) );
  NAND2_X1 U10493 ( .A1(n12152), .A2(n8154), .ZN(n13335) );
  OR2_X1 U10494 ( .A1(n9421), .A2(n8155), .ZN(n12946) );
  INV_X1 U10495 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n13348) );
  OR2_X1 U10496 ( .A1(n8156), .A2(n13348), .ZN(n8160) );
  INV_X1 U10497 ( .A(P2_REG2_REG_30__SCAN_IN), .ZN(n13156) );
  OR2_X1 U10498 ( .A1(n8199), .A2(n13156), .ZN(n8159) );
  INV_X1 U10499 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n13434) );
  OR2_X1 U10500 ( .A1(n8157), .A2(n13434), .ZN(n8158) );
  AND3_X1 U10501 ( .A1(n8160), .A2(n8159), .A3(n8158), .ZN(n12154) );
  INV_X1 U10502 ( .A(n12154), .ZN(n13023) );
  NAND2_X1 U10503 ( .A1(n8161), .A2(n8155), .ZN(n12948) );
  NOR2_X1 U10504 ( .A1(n13484), .A2(n8162), .ZN(n8163) );
  NOR2_X1 U10505 ( .A1(n12948), .A2(n8163), .ZN(n8200) );
  INV_X1 U10506 ( .A(n12008), .ZN(n14807) );
  NAND2_X1 U10507 ( .A1(n10444), .A2(n11922), .ZN(n9542) );
  OR2_X1 U10508 ( .A1(n6524), .A2(n9542), .ZN(n9532) );
  NAND2_X1 U10509 ( .A1(n10187), .A2(n10183), .ZN(n10471) );
  NAND2_X1 U10510 ( .A1(n13220), .A2(n13228), .ZN(n13216) );
  NOR2_X2 U10511 ( .A1(n13201), .A2(n13187), .ZN(n13163) );
  AOI211_X1 U10512 ( .C1(n13351), .C2(n13164), .A(n9445), .B(n13155), .ZN(
        n13350) );
  NOR2_X2 U10513 ( .A1(n8170), .A2(n13167), .ZN(n14362) );
  INV_X1 U10514 ( .A(n13351), .ZN(n8174) );
  NOR2_X1 U10515 ( .A1(n9431), .A2(n12183), .ZN(n9413) );
  INV_X1 U10516 ( .A(n13323), .ZN(n14354) );
  INV_X1 U10517 ( .A(n8171), .ZN(n8172) );
  AOI22_X1 U10518 ( .A1(n14367), .A2(P2_REG2_REG_29__SCAN_IN), .B1(n14354), 
        .B2(n8172), .ZN(n8173) );
  OAI21_X1 U10519 ( .B1(n8174), .B2(n13311), .A(n8173), .ZN(n8175) );
  AOI21_X1 U10520 ( .B1(n13350), .B2(n14362), .A(n8175), .ZN(n8176) );
  OAI211_X1 U10521 ( .C1(n13354), .C2(n13342), .A(n7443), .B(n8176), .ZN(
        P2_U3236) );
  NAND2_X1 U10522 ( .A1(n8178), .A2(n8177), .ZN(n8181) );
  INV_X1 U10523 ( .A(SI_29_), .ZN(n11582) );
  NAND2_X1 U10524 ( .A1(n8179), .A2(n11582), .ZN(n8180) );
  MUX2_X1 U10525 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(P1_DATAO_REG_30__SCAN_IN), 
        .S(n9727), .Z(n8182) );
  NAND2_X1 U10526 ( .A1(n8182), .A2(SI_30_), .ZN(n8188) );
  OAI21_X1 U10527 ( .B1(n8182), .B2(SI_30_), .A(n8188), .ZN(n8183) );
  NAND2_X1 U10528 ( .A1(n8184), .A2(n8183), .ZN(n8185) );
  INV_X1 U10529 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n11905) );
  OR2_X1 U10530 ( .A1(n8193), .A2(n11905), .ZN(n8186) );
  MUX2_X1 U10531 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n9727), .Z(n8190) );
  XNOR2_X1 U10532 ( .A(n8190), .B(SI_31_), .ZN(n8191) );
  INV_X1 U10533 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n11659) );
  OR2_X1 U10534 ( .A1(n8193), .A2(n11659), .ZN(n8194) );
  INV_X1 U10535 ( .A(P2_REG2_REG_31__SCAN_IN), .ZN(n8198) );
  NAND2_X1 U10536 ( .A1(n8195), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n8197) );
  NAND2_X1 U10537 ( .A1(n7596), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n8196) );
  OAI211_X1 U10538 ( .C1(n8199), .C2(n8198), .A(n8197), .B(n8196), .ZN(n13022)
         );
  AND2_X1 U10539 ( .A1(n8200), .A2(n13022), .ZN(n13151) );
  AOI21_X1 U10540 ( .B1(n13150), .B2(n9550), .A(n13151), .ZN(n13343) );
  INV_X1 U10541 ( .A(n9409), .ZN(n14772) );
  AND2_X1 U10542 ( .A1(n9412), .A2(n8201), .ZN(n9435) );
  INV_X1 U10543 ( .A(n14769), .ZN(n9410) );
  NOR2_X1 U10544 ( .A1(n9433), .A2(n9410), .ZN(n8202) );
  OR2_X1 U10545 ( .A1(n13343), .A2(n14819), .ZN(n8208) );
  INV_X1 U10546 ( .A(n9431), .ZN(n8203) );
  NAND2_X1 U10547 ( .A1(n8203), .A2(n12180), .ZN(n14806) );
  NAND2_X1 U10548 ( .A1(n14821), .A2(n14810), .ZN(n13468) );
  INV_X1 U10549 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n8204) );
  INV_X1 U10550 ( .A(n8206), .ZN(n8207) );
  NAND2_X1 U10551 ( .A1(n8208), .A2(n8207), .ZN(P2_U3498) );
  INV_X1 U10552 ( .A(P3_ADDR_REG_14__SCAN_IN), .ZN(n8230) );
  INV_X1 U10553 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n8209) );
  XOR2_X1 U10554 ( .A(n8230), .B(n8209), .Z(n8283) );
  INV_X1 U10555 ( .A(P3_ADDR_REG_13__SCAN_IN), .ZN(n8228) );
  INV_X1 U10556 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n14470) );
  INV_X1 U10557 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n8225) );
  INV_X1 U10558 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n8221) );
  INV_X1 U10559 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n9131) );
  INV_X1 U10560 ( .A(P3_ADDR_REG_6__SCAN_IN), .ZN(n15271) );
  INV_X1 U10561 ( .A(P3_ADDR_REG_3__SCAN_IN), .ZN(n8211) );
  INV_X1 U10562 ( .A(P3_ADDR_REG_5__SCAN_IN), .ZN(n8213) );
  INV_X1 U10563 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n15281) );
  INV_X1 U10564 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n8215) );
  AOI22_X1 U10565 ( .A1(P3_ADDR_REG_6__SCAN_IN), .A2(P1_ADDR_REG_6__SCAN_IN), 
        .B1(n8215), .B2(n15271), .ZN(n8263) );
  INV_X1 U10566 ( .A(P3_ADDR_REG_7__SCAN_IN), .ZN(n8216) );
  NOR2_X1 U10567 ( .A1(n8217), .A2(n8216), .ZN(n8219) );
  XOR2_X1 U10568 ( .A(P3_ADDR_REG_8__SCAN_IN), .B(P1_ADDR_REG_8__SCAN_IN), .Z(
        n8271) );
  XOR2_X1 U10569 ( .A(P3_ADDR_REG_9__SCAN_IN), .B(P1_ADDR_REG_9__SCAN_IN), .Z(
        n8238) );
  NOR2_X1 U10570 ( .A1(P1_ADDR_REG_10__SCAN_IN), .A2(n8222), .ZN(n8224) );
  INV_X1 U10571 ( .A(P3_ADDR_REG_10__SCAN_IN), .ZN(n8237) );
  XNOR2_X1 U10572 ( .A(P1_ADDR_REG_10__SCAN_IN), .B(n8222), .ZN(n8236) );
  INV_X1 U10573 ( .A(P3_ADDR_REG_11__SCAN_IN), .ZN(n10912) );
  XOR2_X1 U10574 ( .A(n10912), .B(n8225), .Z(n8234) );
  XNOR2_X1 U10575 ( .A(P3_ADDR_REG_12__SCAN_IN), .B(n14470), .ZN(n8232) );
  INV_X1 U10576 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n8226) );
  NOR2_X1 U10577 ( .A1(P3_ADDR_REG_13__SCAN_IN), .A2(n8226), .ZN(n8227) );
  INV_X1 U10578 ( .A(P3_ADDR_REG_15__SCAN_IN), .ZN(n12408) );
  NAND2_X1 U10579 ( .A1(P1_ADDR_REG_15__SCAN_IN), .A2(n12408), .ZN(n8231) );
  OAI21_X1 U10580 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(n12408), .A(n8231), .ZN(
        n8285) );
  XNOR2_X1 U10581 ( .A(n8286), .B(n8285), .ZN(n14436) );
  XOR2_X1 U10582 ( .A(n8233), .B(n8232), .Z(n8277) );
  XOR2_X1 U10583 ( .A(n8235), .B(n8234), .Z(n14421) );
  XNOR2_X1 U10584 ( .A(n8237), .B(n8236), .ZN(n8275) );
  XNOR2_X1 U10585 ( .A(n8239), .B(n8238), .ZN(n8273) );
  INV_X1 U10586 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n8241) );
  INV_X1 U10587 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n15156) );
  NAND2_X1 U10588 ( .A1(n8243), .A2(n15156), .ZN(n8258) );
  XNOR2_X1 U10589 ( .A(P2_ADDR_REG_4__SCAN_IN), .B(n8243), .ZN(n15409) );
  XOR2_X1 U10590 ( .A(n8244), .B(P1_ADDR_REG_3__SCAN_IN), .Z(n8255) );
  XNOR2_X1 U10591 ( .A(n8246), .B(n8245), .ZN(n8254) );
  XNOR2_X1 U10592 ( .A(P1_ADDR_REG_1__SCAN_IN), .B(P3_ADDR_REG_1__SCAN_IN), 
        .ZN(n8247) );
  INV_X1 U10593 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n8251) );
  NOR2_X1 U10594 ( .A1(n8250), .A2(n8251), .ZN(n8252) );
  AOI21_X1 U10595 ( .B1(n9882), .B2(P1_ADDR_REG_0__SCAN_IN), .A(n8248), .ZN(
        n8249) );
  INV_X1 U10596 ( .A(n8249), .ZN(n15413) );
  NAND2_X1 U10597 ( .A1(P2_ADDR_REG_0__SCAN_IN), .A2(n15413), .ZN(n15422) );
  XNOR2_X1 U10598 ( .A(n8251), .B(n8250), .ZN(n15421) );
  NOR2_X1 U10599 ( .A1(n15422), .A2(n15421), .ZN(n15420) );
  INV_X1 U10600 ( .A(P2_ADDR_REG_2__SCAN_IN), .ZN(n14282) );
  NAND2_X1 U10601 ( .A1(n8254), .A2(n8253), .ZN(n14281) );
  NAND2_X1 U10602 ( .A1(n8255), .A2(n8256), .ZN(n8257) );
  INV_X1 U10603 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n15418) );
  NAND2_X1 U10604 ( .A1(n15419), .A2(n15418), .ZN(n15417) );
  NAND2_X1 U10605 ( .A1(n8257), .A2(n15417), .ZN(n15408) );
  NAND2_X1 U10606 ( .A1(n8259), .A2(n8260), .ZN(n8261) );
  INV_X1 U10607 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n15411) );
  INV_X1 U10608 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n8264) );
  NOR2_X1 U10609 ( .A1(n8265), .A2(n8264), .ZN(n8266) );
  XOR2_X1 U10610 ( .A(n8263), .B(n8262), .Z(n14285) );
  NOR2_X1 U10611 ( .A1(n14285), .A2(n14284), .ZN(n14283) );
  INV_X1 U10612 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n8269) );
  NOR2_X1 U10613 ( .A1(n8268), .A2(n8269), .ZN(n8270) );
  XOR2_X1 U10614 ( .A(n8267), .B(P1_ADDR_REG_7__SCAN_IN), .Z(n15416) );
  XNOR2_X1 U10615 ( .A(n8269), .B(n8268), .ZN(n15415) );
  NOR2_X1 U10616 ( .A1(n15416), .A2(n15415), .ZN(n15414) );
  XOR2_X1 U10617 ( .A(n8272), .B(n8271), .Z(n14287) );
  INV_X1 U10618 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n14703) );
  INV_X1 U10619 ( .A(n14295), .ZN(n14296) );
  INV_X1 U10620 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n14298) );
  NAND2_X1 U10621 ( .A1(n8276), .A2(n8275), .ZN(n14297) );
  NAND2_X1 U10622 ( .A1(n14298), .A2(n14297), .ZN(n14294) );
  NAND2_X1 U10623 ( .A1(n8277), .A2(n8278), .ZN(n8279) );
  INV_X1 U10624 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n15365) );
  NAND2_X1 U10625 ( .A1(n14425), .A2(n15365), .ZN(n14424) );
  XNOR2_X1 U10626 ( .A(P3_ADDR_REG_13__SCAN_IN), .B(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n8281) );
  XNOR2_X1 U10627 ( .A(n8281), .B(n8280), .ZN(n14427) );
  XNOR2_X1 U10628 ( .A(n8283), .B(n8282), .ZN(n14432) );
  NAND2_X1 U10629 ( .A1(n14431), .A2(n14432), .ZN(n14430) );
  NAND2_X1 U10630 ( .A1(n14436), .A2(n14435), .ZN(n8284) );
  NOR2_X1 U10631 ( .A1(n8286), .A2(n8285), .ZN(n8287) );
  INV_X1 U10632 ( .A(P3_ADDR_REG_16__SCAN_IN), .ZN(n12429) );
  NOR2_X1 U10633 ( .A1(P1_ADDR_REG_16__SCAN_IN), .A2(n12429), .ZN(n8288) );
  AOI21_X1 U10634 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(n12429), .A(n8288), .ZN(
        n8290) );
  XOR2_X1 U10635 ( .A(n8291), .B(n8290), .Z(n14439) );
  NAND2_X1 U10636 ( .A1(n14440), .A2(n14439), .ZN(n8289) );
  NAND2_X1 U10637 ( .A1(n8291), .A2(n8290), .ZN(n8292) );
  INV_X1 U10638 ( .A(P3_ADDR_REG_17__SCAN_IN), .ZN(n12445) );
  NAND2_X1 U10639 ( .A1(P1_ADDR_REG_17__SCAN_IN), .A2(n12445), .ZN(n8293) );
  OAI21_X1 U10640 ( .B1(P1_ADDR_REG_17__SCAN_IN), .B2(n12445), .A(n8293), .ZN(
        n8294) );
  XNOR2_X1 U10641 ( .A(n8295), .B(n8294), .ZN(n14300) );
  NOR2_X1 U10642 ( .A1(n8295), .A2(n8294), .ZN(n8296) );
  AOI21_X1 U10643 ( .B1(P1_ADDR_REG_17__SCAN_IN), .B2(n12445), .A(n8296), .ZN(
        n8300) );
  INV_X1 U10644 ( .A(P3_ADDR_REG_18__SCAN_IN), .ZN(n15142) );
  NAND2_X1 U10645 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(n15142), .ZN(n8297) );
  OAI21_X1 U10646 ( .B1(P1_ADDR_REG_18__SCAN_IN), .B2(n15142), .A(n8297), .ZN(
        n8299) );
  XNOR2_X1 U10647 ( .A(P2_ADDR_REG_19__SCAN_IN), .B(P1_ADDR_REG_19__SCAN_IN), 
        .ZN(n8298) );
  NOR2_X1 U10648 ( .A1(n8300), .A2(n8299), .ZN(n8301) );
  AOI21_X1 U10649 ( .B1(P1_ADDR_REG_18__SCAN_IN), .B2(n15142), .A(n8301), .ZN(
        n8303) );
  NOR2_X2 U10650 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P1_IR_REG_17__SCAN_IN), 
        .ZN(n8348) );
  NOR2_X1 U10651 ( .A1(P1_IR_REG_18__SCAN_IN), .A2(P1_IR_REG_20__SCAN_IN), 
        .ZN(n8305) );
  NAND3_X1 U10652 ( .A1(n8336), .A2(n7159), .A3(n8306), .ZN(n8307) );
  NAND2_X1 U10653 ( .A1(n8365), .A2(n8309), .ZN(n8378) );
  INV_X1 U10654 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n8318) );
  XNOR2_X2 U10655 ( .A(n8319), .B(P1_IR_REG_30__SCAN_IN), .ZN(n8325) );
  INV_X1 U10656 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n8321) );
  XNOR2_X2 U10657 ( .A(n8322), .B(n8321), .ZN(n11637) );
  AND2_X4 U10658 ( .A1(n8325), .A2(n11637), .ZN(n8780) );
  NAND2_X1 U10659 ( .A1(n8780), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n8329) );
  AND2_X4 U10660 ( .A1(n11635), .A2(n11637), .ZN(n8763) );
  NAND2_X1 U10661 ( .A1(n8763), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n8328) );
  INV_X1 U10662 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n8323) );
  OR2_X1 U10663 ( .A1(n8781), .A2(n8323), .ZN(n8327) );
  NAND2_X1 U10664 ( .A1(n8674), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n8326) );
  NAND4_X4 U10665 ( .A1(n8329), .A2(n8328), .A3(n8327), .A4(n8326), .ZN(n8344)
         );
  INV_X1 U10666 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n14445) );
  NOR2_X1 U10667 ( .A1(n9727), .A2(n9728), .ZN(n8330) );
  XNOR2_X1 U10668 ( .A(n8330), .B(P2_DATAO_REG_0__SCAN_IN), .ZN(n14272) );
  XNOR2_X2 U10669 ( .A(n8332), .B(n8331), .ZN(n11640) );
  XNOR2_X2 U10670 ( .A(n8334), .B(n8333), .ZN(n14264) );
  MUX2_X1 U10671 ( .A(n14445), .B(n14272), .S(n9059), .Z(n9669) );
  INV_X1 U10672 ( .A(n9669), .ZN(n14553) );
  NAND2_X1 U10673 ( .A1(n8344), .A2(n14553), .ZN(n9654) );
  INV_X1 U10674 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n8347) );
  NAND2_X1 U10675 ( .A1(n8347), .A2(n8353), .ZN(n8338) );
  INV_X1 U10676 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n8339) );
  INV_X1 U10677 ( .A(n8341), .ZN(n8342) );
  NAND2_X1 U10678 ( .A1(n8345), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8343) );
  OR2_X2 U10679 ( .A1(n8344), .A2(n9669), .ZN(n9661) );
  NAND2_X1 U10680 ( .A1(n8348), .A2(n8347), .ZN(n8349) );
  OR2_X1 U10681 ( .A1(n8605), .A2(n8349), .ZN(n8356) );
  AND2_X1 U10682 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_19__SCAN_IN), 
        .ZN(n8350) );
  NAND2_X1 U10683 ( .A1(n8605), .A2(n8350), .ZN(n8355) );
  OAI21_X1 U10684 ( .B1(P1_IR_REG_18__SCAN_IN), .B2(P1_IR_REG_17__SCAN_IN), 
        .A(P1_IR_REG_19__SCAN_IN), .ZN(n8351) );
  NAND2_X1 U10685 ( .A1(n8351), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8352) );
  OAI21_X1 U10686 ( .B1(P1_IR_REG_31__SCAN_IN), .B2(n8353), .A(n8352), .ZN(
        n8354) );
  NAND2_X1 U10687 ( .A1(n14271), .A2(n8928), .ZN(n9243) );
  NAND2_X1 U10688 ( .A1(n9243), .A2(n8357), .ZN(n8791) );
  MUX2_X1 U10689 ( .A(n9242), .B(n10459), .S(n8791), .Z(n8368) );
  NAND2_X1 U10690 ( .A1(n8763), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n8362) );
  INV_X1 U10691 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n8358) );
  OR2_X1 U10692 ( .A1(n8781), .A2(n8358), .ZN(n8361) );
  INV_X1 U10693 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n8359) );
  OR2_X1 U10694 ( .A1(n8399), .A2(n8359), .ZN(n8360) );
  NAND2_X1 U10695 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), 
        .ZN(n8364) );
  MUX2_X1 U10696 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8364), .S(
        P1_IR_REG_1__SCAN_IN), .Z(n8367) );
  INV_X1 U10697 ( .A(n8365), .ZN(n8366) );
  NAND2_X1 U10698 ( .A1(n8367), .A2(n8366), .ZN(n13778) );
  INV_X1 U10699 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n8950) );
  INV_X4 U10700 ( .A(n8368), .ZN(n8788) );
  MUX2_X1 U10701 ( .A(n6539), .B(n14556), .S(n8788), .Z(n8369) );
  NAND2_X1 U10702 ( .A1(n14556), .A2(n6539), .ZN(n8370) );
  NAND2_X1 U10703 ( .A1(n8780), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n8375) );
  NAND2_X1 U10704 ( .A1(n8763), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n8374) );
  INV_X1 U10705 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n8371) );
  INV_X1 U10706 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n9666) );
  OR2_X1 U10707 ( .A1(n8399), .A2(n9666), .ZN(n8372) );
  INV_X2 U10708 ( .A(n8785), .ZN(n8417) );
  NAND2_X1 U10709 ( .A1(n8952), .A2(n6533), .ZN(n8382) );
  INV_X2 U10710 ( .A(n8376), .ZN(n8633) );
  INV_X1 U10711 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n14258) );
  NOR2_X1 U10712 ( .A1(n8365), .A2(n14258), .ZN(n8377) );
  MUX2_X1 U10713 ( .A(n14258), .B(n8377), .S(P1_IR_REG_2__SCAN_IN), .Z(n8380)
         );
  NAND2_X1 U10714 ( .A1(n13772), .A2(n8770), .ZN(n8384) );
  INV_X1 U10715 ( .A(n13772), .ZN(n14582) );
  NAND2_X1 U10716 ( .A1(n14582), .A2(n8788), .ZN(n8383) );
  NAND2_X1 U10717 ( .A1(n8780), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n8389) );
  NAND2_X1 U10718 ( .A1(n8763), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n8388) );
  INV_X1 U10719 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n8385) );
  OR2_X1 U10720 ( .A1(n8399), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n8386) );
  NAND4_X1 U10721 ( .A1(n8389), .A2(n8388), .A3(n8387), .A4(n8386), .ZN(n13771) );
  NAND2_X1 U10722 ( .A1(n8986), .A2(n6533), .ZN(n8392) );
  NAND2_X1 U10723 ( .A1(n8379), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8390) );
  XNOR2_X1 U10724 ( .A(n8390), .B(P1_IR_REG_3__SCAN_IN), .ZN(n13808) );
  AOI22_X1 U10725 ( .A1(n8622), .A2(P2_DATAO_REG_3__SCAN_IN), .B1(n8633), .B2(
        n13808), .ZN(n8391) );
  INV_X1 U10726 ( .A(n14599), .ZN(n14545) );
  NAND2_X1 U10727 ( .A1(n14599), .A2(n13771), .ZN(n8395) );
  AND2_X1 U10728 ( .A1(n9762), .A2(n8395), .ZN(n9761) );
  NAND3_X1 U10729 ( .A1(n8394), .A2(n8393), .A3(n9761), .ZN(n8406) );
  MUX2_X1 U10730 ( .A(n8395), .B(n9762), .S(n8770), .Z(n8405) );
  OR2_X1 U10731 ( .A1(n8993), .A2(n8785), .ZN(n8398) );
  OR2_X1 U10732 ( .A1(n8379), .A2(P1_IR_REG_3__SCAN_IN), .ZN(n8418) );
  NAND2_X1 U10733 ( .A1(n8418), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8396) );
  XNOR2_X1 U10734 ( .A(n8396), .B(P1_IR_REG_4__SCAN_IN), .ZN(n9232) );
  AOI22_X1 U10735 ( .A1(n8622), .A2(P2_DATAO_REG_4__SCAN_IN), .B1(n8633), .B2(
        n9232), .ZN(n8397) );
  NAND2_X1 U10736 ( .A1(n8776), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n8403) );
  NAND2_X1 U10737 ( .A1(n8780), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n8402) );
  NAND2_X1 U10738 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n8411) );
  OAI21_X1 U10739 ( .B1(P1_REG3_REG_4__SCAN_IN), .B2(P1_REG3_REG_3__SCAN_IN), 
        .A(n8411), .ZN(n9932) );
  OR2_X1 U10740 ( .A1(n8752), .A2(n9932), .ZN(n8401) );
  NAND2_X1 U10741 ( .A1(n8763), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n8400) );
  NAND4_X1 U10742 ( .A1(n8403), .A2(n8402), .A3(n8401), .A4(n8400), .ZN(n8944)
         );
  NAND2_X1 U10743 ( .A1(n14608), .A2(n13770), .ZN(n9862) );
  NAND2_X1 U10744 ( .A1(n9854), .A2(n8944), .ZN(n8404) );
  NAND3_X1 U10745 ( .A1(n8406), .A2(n8405), .A3(n7448), .ZN(n8410) );
  AND2_X1 U10746 ( .A1(n8944), .A2(n8770), .ZN(n8408) );
  OAI21_X1 U10747 ( .B1(n8770), .B2(n8944), .A(n14608), .ZN(n8407) );
  OAI21_X1 U10748 ( .B1(n8408), .B2(n14608), .A(n8407), .ZN(n8409) );
  NAND2_X1 U10749 ( .A1(n8410), .A2(n8409), .ZN(n8426) );
  NAND2_X1 U10750 ( .A1(n8763), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n8416) );
  INV_X1 U10751 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n9107) );
  OR2_X1 U10752 ( .A1(n8781), .A2(n9107), .ZN(n8415) );
  INV_X1 U10753 ( .A(n8780), .ZN(n8553) );
  INV_X1 U10754 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n9119) );
  OR2_X1 U10755 ( .A1(n8553), .A2(n9119), .ZN(n8414) );
  AND2_X1 U10756 ( .A1(n8411), .A2(n9162), .ZN(n8412) );
  OR2_X1 U10757 ( .A1(n8412), .A2(n8434), .ZN(n14528) );
  OR2_X1 U10758 ( .A1(n8752), .A2(n14528), .ZN(n8413) );
  NAND2_X1 U10759 ( .A1(n9062), .A2(n8417), .ZN(n8423) );
  INV_X1 U10760 ( .A(n8418), .ZN(n8420) );
  NAND2_X1 U10761 ( .A1(n8420), .A2(n8419), .ZN(n8428) );
  NAND2_X1 U10762 ( .A1(n8428), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8421) );
  XNOR2_X1 U10763 ( .A(n8421), .B(P1_IR_REG_5__SCAN_IN), .ZN(n9164) );
  AOI22_X1 U10764 ( .A1(n8622), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n8633), .B2(
        n9164), .ZN(n8422) );
  MUX2_X1 U10765 ( .A(n9866), .B(n14615), .S(n8770), .Z(n8425) );
  INV_X1 U10766 ( .A(n14615), .ZN(n14530) );
  MUX2_X1 U10767 ( .A(n13769), .B(n14530), .S(n8788), .Z(n8424) );
  NAND2_X1 U10768 ( .A1(n8426), .A2(n8425), .ZN(n8427) );
  NAND2_X1 U10769 ( .A1(n9067), .A2(n8417), .ZN(n8433) );
  INV_X1 U10770 ( .A(n8428), .ZN(n8430) );
  NAND2_X1 U10771 ( .A1(n8430), .A2(n8429), .ZN(n8442) );
  NAND2_X1 U10772 ( .A1(n8442), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8431) );
  XNOR2_X1 U10773 ( .A(n8431), .B(P1_IR_REG_6__SCAN_IN), .ZN(n9121) );
  AOI22_X1 U10774 ( .A1(n8622), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n8633), .B2(
        n9121), .ZN(n8432) );
  NAND2_X1 U10775 ( .A1(n8433), .A2(n8432), .ZN(n10315) );
  NAND2_X1 U10776 ( .A1(n8776), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n8439) );
  NAND2_X1 U10777 ( .A1(n8780), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n8438) );
  NAND2_X1 U10778 ( .A1(n8763), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n8437) );
  NAND2_X1 U10779 ( .A1(n8434), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n8448) );
  OR2_X1 U10780 ( .A1(n8434), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n8435) );
  NAND2_X1 U10781 ( .A1(n8448), .A2(n8435), .ZN(n9954) );
  OR2_X1 U10782 ( .A1(n8752), .A2(n9954), .ZN(n8436) );
  NAND4_X1 U10783 ( .A1(n8439), .A2(n8438), .A3(n8437), .A4(n8436), .ZN(n13768) );
  MUX2_X1 U10784 ( .A(n10315), .B(n13768), .S(n8770), .Z(n8440) );
  MUX2_X1 U10785 ( .A(n10315), .B(n13768), .S(n8788), .Z(n8441) );
  OR2_X1 U10786 ( .A1(n9086), .A2(n8785), .ZN(n8447) );
  OAI21_X1 U10787 ( .B1(n8442), .B2(P1_IR_REG_6__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n8443) );
  MUX2_X1 U10788 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8443), .S(
        P1_IR_REG_7__SCAN_IN), .Z(n8445) );
  AND2_X1 U10789 ( .A1(n8445), .A2(n8444), .ZN(n9211) );
  AOI22_X1 U10790 ( .A1(n8622), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n8633), .B2(
        n9211), .ZN(n8446) );
  NAND2_X1 U10791 ( .A1(n8447), .A2(n8446), .ZN(n14517) );
  NAND2_X1 U10792 ( .A1(n8776), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n8453) );
  NAND2_X1 U10793 ( .A1(n8780), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n8452) );
  NAND2_X1 U10794 ( .A1(n8763), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n8451) );
  NAND2_X1 U10795 ( .A1(n8448), .A2(n9208), .ZN(n8449) );
  NAND2_X1 U10796 ( .A1(n8474), .A2(n8449), .ZN(n14515) );
  OR2_X1 U10797 ( .A1(n8752), .A2(n14515), .ZN(n8450) );
  NAND4_X1 U10798 ( .A1(n8453), .A2(n8452), .A3(n8451), .A4(n8450), .ZN(n13767) );
  MUX2_X1 U10799 ( .A(n14517), .B(n13767), .S(n8788), .Z(n8457) );
  MUX2_X1 U10800 ( .A(n14517), .B(n13767), .S(n8770), .Z(n8454) );
  NAND2_X1 U10801 ( .A1(n8455), .A2(n8454), .ZN(n8461) );
  INV_X1 U10802 ( .A(n8456), .ZN(n8459) );
  INV_X1 U10803 ( .A(n8457), .ZN(n8458) );
  NAND2_X1 U10804 ( .A1(n8459), .A2(n8458), .ZN(n8460) );
  NAND2_X1 U10805 ( .A1(n8461), .A2(n8460), .ZN(n8470) );
  NAND2_X1 U10806 ( .A1(n8776), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n8465) );
  NAND2_X1 U10807 ( .A1(n8780), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n8464) );
  NAND2_X1 U10808 ( .A1(n8763), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n8463) );
  INV_X1 U10809 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n10609) );
  XNOR2_X1 U10810 ( .A(n8474), .B(n10609), .ZN(n10360) );
  OR2_X1 U10811 ( .A1(n8752), .A2(n10360), .ZN(n8462) );
  NAND4_X1 U10812 ( .A1(n8465), .A2(n8464), .A3(n8463), .A4(n8462), .ZN(n13766) );
  NAND2_X1 U10813 ( .A1(n8444), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8466) );
  XNOR2_X1 U10814 ( .A(n8466), .B(P1_IR_REG_8__SCAN_IN), .ZN(n9140) );
  AOI22_X1 U10815 ( .A1(n8622), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n8633), .B2(
        n9140), .ZN(n8467) );
  MUX2_X1 U10816 ( .A(n13766), .B(n10600), .S(n8788), .Z(n8471) );
  MUX2_X1 U10817 ( .A(n10600), .B(n13766), .S(n8788), .Z(n8469) );
  NAND2_X1 U10818 ( .A1(n8776), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n8479) );
  NAND2_X1 U10819 ( .A1(n8780), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n8478) );
  NAND2_X1 U10820 ( .A1(n8763), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n8477) );
  INV_X1 U10821 ( .A(n8474), .ZN(n8472) );
  AOI21_X1 U10822 ( .B1(n8472), .B2(P1_REG3_REG_8__SCAN_IN), .A(
        P1_REG3_REG_9__SCAN_IN), .ZN(n8475) );
  NAND2_X1 U10823 ( .A1(P1_REG3_REG_9__SCAN_IN), .A2(P1_REG3_REG_8__SCAN_IN), 
        .ZN(n8473) );
  OR2_X1 U10824 ( .A1(n8475), .A2(n8495), .ZN(n14498) );
  OR2_X1 U10825 ( .A1(n8752), .A2(n14498), .ZN(n8476) );
  NAND4_X1 U10826 ( .A1(n8479), .A2(n8478), .A3(n8477), .A4(n8476), .ZN(n13765) );
  NOR2_X1 U10827 ( .A1(n8444), .A2(P1_IR_REG_8__SCAN_IN), .ZN(n8483) );
  INV_X1 U10828 ( .A(n8483), .ZN(n8480) );
  NAND2_X1 U10829 ( .A1(n8480), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8481) );
  MUX2_X1 U10830 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8481), .S(
        P1_IR_REG_9__SCAN_IN), .Z(n8484) );
  INV_X1 U10831 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n8482) );
  NAND2_X1 U10832 ( .A1(n8483), .A2(n8482), .ZN(n8511) );
  NAND2_X1 U10833 ( .A1(n8484), .A2(n8511), .ZN(n9260) );
  INV_X1 U10834 ( .A(n9260), .ZN(n9256) );
  AOI22_X1 U10835 ( .A1(n8622), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n8633), .B2(
        n9256), .ZN(n8485) );
  MUX2_X1 U10836 ( .A(n13765), .B(n14500), .S(n8770), .Z(n8490) );
  MUX2_X1 U10837 ( .A(n13765), .B(n14500), .S(n8788), .Z(n8487) );
  NAND2_X1 U10838 ( .A1(n8488), .A2(n8487), .ZN(n8494) );
  INV_X1 U10839 ( .A(n8489), .ZN(n8492) );
  INV_X1 U10840 ( .A(n8490), .ZN(n8491) );
  NAND2_X1 U10841 ( .A1(n8492), .A2(n8491), .ZN(n8493) );
  NAND2_X1 U10842 ( .A1(n8494), .A2(n8493), .ZN(n8505) );
  NAND2_X1 U10843 ( .A1(n8780), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n8500) );
  NAND2_X1 U10844 ( .A1(n8763), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n8499) );
  NAND2_X1 U10845 ( .A1(n8776), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n8498) );
  OR2_X1 U10846 ( .A1(n8495), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n8496) );
  NAND2_X1 U10847 ( .A1(n8520), .A2(n8496), .ZN(n10836) );
  OR2_X1 U10848 ( .A1(n8752), .A2(n10836), .ZN(n8497) );
  NAND4_X1 U10849 ( .A1(n8500), .A2(n8499), .A3(n8498), .A4(n8497), .ZN(n13764) );
  NAND2_X1 U10850 ( .A1(n8511), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8501) );
  XNOR2_X1 U10851 ( .A(n8501), .B(P1_IR_REG_10__SCAN_IN), .ZN(n9477) );
  AOI22_X1 U10852 ( .A1(n8622), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n8633), 
        .B2(n9477), .ZN(n8502) );
  MUX2_X1 U10853 ( .A(n13764), .B(n14635), .S(n8788), .Z(n8506) );
  MUX2_X1 U10854 ( .A(n13764), .B(n14635), .S(n8770), .Z(n8504) );
  NAND2_X1 U10855 ( .A1(n8776), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n8510) );
  INV_X1 U10856 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n10817) );
  OR2_X1 U10857 ( .A1(n8553), .A2(n10817), .ZN(n8509) );
  XNOR2_X1 U10858 ( .A(n8520), .B(n8519), .ZN(n11027) );
  OR2_X1 U10859 ( .A1(n8752), .A2(n11027), .ZN(n8508) );
  NAND2_X1 U10860 ( .A1(n8763), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n8507) );
  NAND4_X1 U10861 ( .A1(n8510), .A2(n8509), .A3(n8508), .A4(n8507), .ZN(n13763) );
  NAND2_X1 U10862 ( .A1(n8526), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8512) );
  INV_X1 U10863 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n8527) );
  XNOR2_X1 U10864 ( .A(n8512), .B(n8527), .ZN(n9907) );
  INV_X1 U10865 ( .A(n9907), .ZN(n9486) );
  AOI22_X1 U10866 ( .A1(n8622), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n8633), 
        .B2(n9486), .ZN(n8513) );
  MUX2_X1 U10867 ( .A(n13763), .B(n11018), .S(n8770), .Z(n8517) );
  MUX2_X1 U10868 ( .A(n13763), .B(n11018), .S(n8788), .Z(n8515) );
  INV_X1 U10869 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n10865) );
  OR2_X1 U10870 ( .A1(n8553), .A2(n10865), .ZN(n8525) );
  NAND2_X1 U10871 ( .A1(n8763), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n8524) );
  OAI21_X1 U10872 ( .B1(n8520), .B2(n8519), .A(n8518), .ZN(n8521) );
  NAND2_X1 U10873 ( .A1(n8521), .A2(n8536), .ZN(n13660) );
  OR2_X1 U10874 ( .A1(n8752), .A2(n13660), .ZN(n8523) );
  NAND2_X1 U10875 ( .A1(n8776), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n8522) );
  NAND4_X1 U10876 ( .A1(n8525), .A2(n8524), .A3(n8523), .A4(n8522), .ZN(n13762) );
  NAND2_X1 U10877 ( .A1(n9510), .A2(n8417), .ZN(n8531) );
  INV_X1 U10878 ( .A(n8526), .ZN(n8528) );
  NAND2_X1 U10879 ( .A1(n8528), .A2(n8527), .ZN(n8542) );
  NAND2_X1 U10880 ( .A1(n8542), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8529) );
  XNOR2_X1 U10881 ( .A(n8529), .B(P1_IR_REG_12__SCAN_IN), .ZN(n14461) );
  AOI22_X1 U10882 ( .A1(n8622), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n8633), 
        .B2(n14461), .ZN(n8530) );
  MUX2_X1 U10883 ( .A(n13762), .B(n13667), .S(n8788), .Z(n8533) );
  MUX2_X1 U10884 ( .A(n13762), .B(n13667), .S(n8770), .Z(n8532) );
  INV_X1 U10885 ( .A(n8533), .ZN(n8534) );
  NAND2_X1 U10886 ( .A1(n8780), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n8541) );
  NAND2_X1 U10887 ( .A1(n8763), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n8540) );
  NAND2_X1 U10888 ( .A1(n8776), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n8539) );
  INV_X1 U10889 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n8535) );
  AND2_X1 U10890 ( .A1(n8536), .A2(n8535), .ZN(n8537) );
  OR2_X1 U10891 ( .A1(n8537), .A2(n8555), .ZN(n11251) );
  OR2_X1 U10892 ( .A1(n8752), .A2(n11251), .ZN(n8538) );
  NAND4_X1 U10893 ( .A1(n8541), .A2(n8540), .A3(n8539), .A4(n8538), .ZN(n13761) );
  NAND2_X1 U10894 ( .A1(n9514), .A2(n8417), .ZN(n8546) );
  NAND2_X1 U10895 ( .A1(n8543), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8548) );
  INV_X1 U10896 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n8547) );
  XNOR2_X1 U10897 ( .A(n8548), .B(n8547), .ZN(n14471) );
  OAI22_X1 U10898 ( .A1(n8796), .A2(n9515), .B1(n14471), .B2(n9059), .ZN(n8544) );
  INV_X1 U10899 ( .A(n8544), .ZN(n8545) );
  MUX2_X1 U10900 ( .A(n13761), .B(n11253), .S(n8770), .Z(n8580) );
  NAND2_X1 U10901 ( .A1(n8579), .A2(n8580), .ZN(n8578) );
  NAND2_X1 U10902 ( .A1(n9593), .A2(n8417), .ZN(n8552) );
  NAND2_X1 U10903 ( .A1(n8548), .A2(n8547), .ZN(n8549) );
  NAND2_X1 U10904 ( .A1(n8549), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8550) );
  XNOR2_X1 U10905 ( .A(n8550), .B(P1_IR_REG_14__SCAN_IN), .ZN(n10336) );
  AOI22_X1 U10906 ( .A1(n10336), .A2(n8633), .B1(n8622), .B2(
        P2_DATAO_REG_14__SCAN_IN), .ZN(n8551) );
  NAND2_X1 U10907 ( .A1(n8763), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n8560) );
  INV_X1 U10908 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n11214) );
  OR2_X1 U10909 ( .A1(n8553), .A2(n11214), .ZN(n8559) );
  INV_X1 U10910 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n8554) );
  OR2_X1 U10911 ( .A1(n8781), .A2(n8554), .ZN(n8558) );
  NOR2_X1 U10912 ( .A1(n8555), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n8556) );
  OR2_X1 U10913 ( .A1(n8566), .A2(n8556), .ZN(n14402) );
  OR2_X1 U10914 ( .A1(n8752), .A2(n14402), .ZN(n8557) );
  NAND2_X1 U10915 ( .A1(n14405), .A2(n13506), .ZN(n11295) );
  NAND2_X1 U10916 ( .A1(n8578), .A2(n7430), .ZN(n8575) );
  NAND2_X1 U10917 ( .A1(n9784), .A2(n8417), .ZN(n8565) );
  NOR2_X1 U10918 ( .A1(n8561), .A2(n14258), .ZN(n8562) );
  MUX2_X1 U10919 ( .A(n14258), .B(n8562), .S(P1_IR_REG_15__SCAN_IN), .Z(n8563)
         );
  NOR2_X1 U10920 ( .A1(n8563), .A2(n8598), .ZN(n10342) );
  AOI22_X1 U10921 ( .A1(n8622), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n8633), 
        .B2(n10342), .ZN(n8564) );
  NAND2_X1 U10922 ( .A1(n8780), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n8571) );
  INV_X1 U10923 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n15145) );
  OR2_X1 U10924 ( .A1(n8781), .A2(n15145), .ZN(n8570) );
  OR2_X1 U10925 ( .A1(n8566), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n8567) );
  NAND2_X1 U10926 ( .A1(n8592), .A2(n8567), .ZN(n13752) );
  OR2_X1 U10927 ( .A1(n8752), .A2(n13752), .ZN(n8569) );
  INV_X1 U10928 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n14255) );
  OR2_X1 U10929 ( .A1(n8784), .A2(n14255), .ZN(n8568) );
  NAND2_X1 U10930 ( .A1(n13754), .A2(n13517), .ZN(n8813) );
  INV_X1 U10931 ( .A(n8813), .ZN(n8573) );
  NAND2_X1 U10932 ( .A1(n8575), .A2(n8574), .ZN(n8576) );
  NAND2_X1 U10933 ( .A1(n8576), .A2(n8788), .ZN(n8588) );
  AND4_X1 U10934 ( .A1(n11212), .A2(n8813), .A3(n8770), .A4(n13761), .ZN(n8577) );
  NAND2_X1 U10935 ( .A1(n8578), .A2(n8577), .ZN(n8587) );
  INV_X1 U10936 ( .A(n8580), .ZN(n8581) );
  NAND4_X1 U10937 ( .A1(n8582), .A2(n8581), .A3(n11212), .A4(n8813), .ZN(n8586) );
  INV_X1 U10938 ( .A(n8583), .ZN(n11296) );
  INV_X1 U10939 ( .A(n13517), .ZN(n13759) );
  OAI21_X1 U10940 ( .B1(n8583), .B2(n13517), .A(n13754), .ZN(n8584) );
  OAI211_X1 U10941 ( .C1(n11296), .C2(n13759), .A(n8584), .B(n8770), .ZN(n8585) );
  NAND2_X1 U10942 ( .A1(n8588), .A2(n7444), .ZN(n8590) );
  OR2_X1 U10943 ( .A1(n11389), .A2(n8770), .ZN(n8589) );
  NAND2_X1 U10944 ( .A1(n8590), .A2(n8589), .ZN(n8618) );
  NAND2_X1 U10945 ( .A1(n8776), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n8597) );
  NAND2_X1 U10946 ( .A1(n8780), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n8596) );
  NAND2_X1 U10947 ( .A1(n8763), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n8595) );
  INV_X1 U10948 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n8591) );
  NAND2_X1 U10949 ( .A1(n8592), .A2(n8591), .ZN(n8593) );
  NAND2_X1 U10950 ( .A1(n8610), .A2(n8593), .ZN(n13685) );
  OR2_X1 U10951 ( .A1(n8752), .A2(n13685), .ZN(n8594) );
  NAND4_X1 U10952 ( .A1(n8597), .A2(n8596), .A3(n8595), .A4(n8594), .ZN(n14106) );
  NAND2_X1 U10953 ( .A1(n9914), .A2(n8417), .ZN(n8603) );
  NOR2_X1 U10954 ( .A1(n8598), .A2(n14258), .ZN(n8599) );
  MUX2_X1 U10955 ( .A(n14258), .B(n8599), .S(P1_IR_REG_16__SCAN_IN), .Z(n8601)
         );
  INV_X1 U10956 ( .A(n8605), .ZN(n8600) );
  NOR2_X1 U10957 ( .A1(n8601), .A2(n8600), .ZN(n11194) );
  AOI22_X1 U10958 ( .A1(n8622), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n8633), 
        .B2(n11194), .ZN(n8602) );
  MUX2_X1 U10959 ( .A(n14106), .B(n13890), .S(n8770), .Z(n8617) );
  INV_X1 U10960 ( .A(n14106), .ZN(n13864) );
  INV_X1 U10961 ( .A(n13890), .ZN(n14223) );
  MUX2_X1 U10962 ( .A(n13864), .B(n14223), .S(n8788), .Z(n8604) );
  NAND2_X1 U10963 ( .A1(n9958), .A2(n8417), .ZN(n8608) );
  NAND2_X1 U10964 ( .A1(n8605), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8606) );
  XNOR2_X1 U10965 ( .A(n8606), .B(P1_IR_REG_17__SCAN_IN), .ZN(n11195) );
  AOI22_X1 U10966 ( .A1(n8622), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n8633), 
        .B2(n11195), .ZN(n8607) );
  INV_X1 U10967 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n8609) );
  AND2_X1 U10968 ( .A1(n8610), .A2(n8609), .ZN(n8611) );
  OR2_X1 U10969 ( .A1(n8611), .A2(n8625), .ZN(n14116) );
  NAND2_X1 U10970 ( .A1(n8776), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n8613) );
  NAND2_X1 U10971 ( .A1(n8780), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n8612) );
  AND2_X1 U10972 ( .A1(n8613), .A2(n8612), .ZN(n8615) );
  NAND2_X1 U10973 ( .A1(n8763), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n8614) );
  OAI211_X1 U10974 ( .C1(n14116), .C2(n8752), .A(n8615), .B(n8614), .ZN(n14088) );
  INV_X1 U10975 ( .A(n14088), .ZN(n13684) );
  NAND2_X1 U10976 ( .A1(n14218), .A2(n13684), .ZN(n8616) );
  OR2_X1 U10977 ( .A1(n14218), .A2(n13684), .ZN(n13867) );
  MUX2_X1 U10978 ( .A(n8616), .B(n13867), .S(n8788), .Z(n8619) );
  NAND2_X1 U10979 ( .A1(n10460), .A2(n8417), .ZN(n8624) );
  NAND2_X1 U10980 ( .A1(n8620), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8621) );
  XNOR2_X1 U10981 ( .A(n8621), .B(P1_IR_REG_18__SCAN_IN), .ZN(n13839) );
  AOI22_X1 U10982 ( .A1(n8622), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n8633), 
        .B2(n13839), .ZN(n8623) );
  NAND2_X2 U10983 ( .A1(n8624), .A2(n8623), .ZN(n14096) );
  NOR2_X1 U10984 ( .A1(n8625), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n8626) );
  OR2_X1 U10985 ( .A1(n8636), .A2(n8626), .ZN(n14092) );
  AOI22_X1 U10986 ( .A1(n8776), .A2(P1_REG1_REG_18__SCAN_IN), .B1(n8780), .B2(
        P1_REG2_REG_18__SCAN_IN), .ZN(n8628) );
  NAND2_X1 U10987 ( .A1(n8763), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n8627) );
  OAI211_X1 U10988 ( .C1(n14092), .C2(n8752), .A(n8628), .B(n8627), .ZN(n14109) );
  XNOR2_X1 U10989 ( .A(n14096), .B(n14109), .ZN(n14091) );
  MUX2_X1 U10990 ( .A(n14088), .B(n14218), .S(n8770), .Z(n8629) );
  INV_X1 U10991 ( .A(n8629), .ZN(n8630) );
  NAND2_X1 U10992 ( .A1(n10656), .A2(n8417), .ZN(n8635) );
  AOI22_X1 U10993 ( .A1(n8622), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n8928), 
        .B2(n8633), .ZN(n8634) );
  OR2_X1 U10994 ( .A1(n8636), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n8637) );
  AND2_X1 U10995 ( .A1(n8648), .A2(n8637), .ZN(n14072) );
  NAND2_X1 U10996 ( .A1(n14072), .A2(n8674), .ZN(n8640) );
  AOI22_X1 U10997 ( .A1(n8776), .A2(P1_REG1_REG_19__SCAN_IN), .B1(n8780), .B2(
        P1_REG2_REG_19__SCAN_IN), .ZN(n8639) );
  INV_X1 U10998 ( .A(P1_REG0_REG_19__SCAN_IN), .ZN(n15370) );
  OR2_X1 U10999 ( .A1(n8784), .A2(n15370), .ZN(n8638) );
  OR2_X1 U11000 ( .A1(n14203), .A2(n14210), .ZN(n8644) );
  NAND2_X1 U11001 ( .A1(n14203), .A2(n14210), .ZN(n13869) );
  AND2_X1 U11002 ( .A1(n14109), .A2(n8788), .ZN(n8642) );
  OAI21_X1 U11003 ( .B1(n8788), .B2(n14109), .A(n14096), .ZN(n8641) );
  OAI21_X1 U11004 ( .B1(n8642), .B2(n14096), .A(n8641), .ZN(n8643) );
  MUX2_X1 U11005 ( .A(n13869), .B(n8644), .S(n8770), .Z(n8645) );
  NAND2_X1 U11006 ( .A1(n8646), .A2(n8645), .ZN(n8659) );
  INV_X1 U11007 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n8647) );
  NAND2_X1 U11008 ( .A1(n8648), .A2(n8647), .ZN(n8649) );
  NAND2_X1 U11009 ( .A1(n8661), .A2(n8649), .ZN(n14057) );
  OR2_X1 U11010 ( .A1(n14057), .A2(n8752), .ZN(n8654) );
  INV_X1 U11011 ( .A(P1_REG0_REG_20__SCAN_IN), .ZN(n15372) );
  NAND2_X1 U11012 ( .A1(n8776), .A2(P1_REG1_REG_20__SCAN_IN), .ZN(n8651) );
  NAND2_X1 U11013 ( .A1(n8780), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n8650) );
  OAI211_X1 U11014 ( .C1(n15372), .C2(n8784), .A(n8651), .B(n8650), .ZN(n8652)
         );
  INV_X1 U11015 ( .A(n8652), .ZN(n8653) );
  NAND2_X1 U11016 ( .A1(n10458), .A2(n8417), .ZN(n8656) );
  OR2_X1 U11017 ( .A1(n8796), .A2(n15263), .ZN(n8655) );
  MUX2_X1 U11018 ( .A(n14074), .B(n14061), .S(n8770), .Z(n8658) );
  INV_X1 U11019 ( .A(n14074), .ZN(n13872) );
  MUX2_X1 U11020 ( .A(n13872), .B(n14197), .S(n8788), .Z(n8657) );
  NAND2_X1 U11021 ( .A1(n8659), .A2(n8658), .ZN(n8660) );
  INV_X1 U11022 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n13653) );
  NAND2_X1 U11023 ( .A1(n8661), .A2(n13653), .ZN(n8662) );
  AND2_X1 U11024 ( .A1(n8673), .A2(n8662), .ZN(n14043) );
  NAND2_X1 U11025 ( .A1(n14043), .A2(n8674), .ZN(n8667) );
  INV_X1 U11026 ( .A(P1_REG0_REG_21__SCAN_IN), .ZN(n15171) );
  NAND2_X1 U11027 ( .A1(n8776), .A2(P1_REG1_REG_21__SCAN_IN), .ZN(n8664) );
  NAND2_X1 U11028 ( .A1(n8780), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n8663) );
  OAI211_X1 U11029 ( .C1(n15171), .C2(n8784), .A(n8664), .B(n8663), .ZN(n8665)
         );
  INV_X1 U11030 ( .A(n8665), .ZN(n8666) );
  NAND2_X1 U11031 ( .A1(n8667), .A2(n8666), .ZN(n14025) );
  NAND2_X1 U11032 ( .A1(n10667), .A2(n8417), .ZN(n8669) );
  INV_X1 U11033 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n10668) );
  OR2_X1 U11034 ( .A1(n8796), .A2(n10668), .ZN(n8668) );
  MUX2_X1 U11035 ( .A(n14025), .B(n14190), .S(n8788), .Z(n8671) );
  MUX2_X1 U11036 ( .A(n14025), .B(n14190), .S(n8770), .Z(n8670) );
  INV_X1 U11037 ( .A(n8671), .ZN(n8672) );
  INV_X1 U11038 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n15322) );
  AOI21_X1 U11039 ( .B1(n8673), .B2(n15322), .A(n8689), .ZN(n14031) );
  NAND2_X1 U11040 ( .A1(n14031), .A2(n8674), .ZN(n8679) );
  INV_X1 U11041 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n15221) );
  NAND2_X1 U11042 ( .A1(n8763), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n8676) );
  NAND2_X1 U11043 ( .A1(n8780), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n8675) );
  OAI211_X1 U11044 ( .C1(n8781), .C2(n15221), .A(n8676), .B(n8675), .ZN(n8677)
         );
  INV_X1 U11045 ( .A(n8677), .ZN(n8678) );
  NAND2_X1 U11046 ( .A1(n8679), .A2(n8678), .ZN(n13900) );
  OR2_X1 U11047 ( .A1(n7948), .A2(n9727), .ZN(n8680) );
  XNOR2_X1 U11048 ( .A(n8680), .B(P2_DATAO_REG_22__SCAN_IN), .ZN(n14270) );
  MUX2_X1 U11049 ( .A(n13900), .B(n14186), .S(n8770), .Z(n8684) );
  MUX2_X1 U11050 ( .A(n13900), .B(n14186), .S(n8788), .Z(n8681) );
  NAND2_X1 U11051 ( .A1(n8682), .A2(n8681), .ZN(n8688) );
  INV_X1 U11052 ( .A(n8683), .ZN(n8686) );
  INV_X1 U11053 ( .A(n8684), .ZN(n8685) );
  NAND2_X1 U11054 ( .A1(n8686), .A2(n8685), .ZN(n8687) );
  NAND2_X1 U11055 ( .A1(n8688), .A2(n8687), .ZN(n8697) );
  NAND2_X1 U11056 ( .A1(n8776), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n8693) );
  NAND2_X1 U11057 ( .A1(n8780), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n8692) );
  NAND2_X1 U11058 ( .A1(n8689), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n8699) );
  OAI21_X1 U11059 ( .B1(P1_REG3_REG_23__SCAN_IN), .B2(n8689), .A(n8699), .ZN(
        n14015) );
  OR2_X1 U11060 ( .A1(n8752), .A2(n14015), .ZN(n8691) );
  NAND2_X1 U11061 ( .A1(n8763), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n8690) );
  NAND4_X1 U11062 ( .A1(n8693), .A2(n8692), .A3(n8691), .A4(n8690), .ZN(n14026) );
  NAND2_X1 U11063 ( .A1(n11010), .A2(n8417), .ZN(n8695) );
  OR2_X1 U11064 ( .A1(n8796), .A2(n15293), .ZN(n8694) );
  MUX2_X1 U11065 ( .A(n14026), .B(n14181), .S(n8788), .Z(n8698) );
  MUX2_X1 U11066 ( .A(n14026), .B(n14181), .S(n8770), .Z(n8696) );
  NAND2_X1 U11067 ( .A1(n8776), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n8704) );
  NAND2_X1 U11068 ( .A1(n8780), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n8703) );
  OAI21_X1 U11069 ( .B1(P1_REG3_REG_24__SCAN_IN), .B2(n8700), .A(n8715), .ZN(
        n13703) );
  OR2_X1 U11070 ( .A1(n8752), .A2(n13703), .ZN(n8702) );
  NAND2_X1 U11071 ( .A1(n8763), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n8701) );
  NAND4_X1 U11072 ( .A1(n8704), .A2(n8703), .A3(n8702), .A4(n8701), .ZN(n13980) );
  NAND2_X1 U11073 ( .A1(n11224), .A2(n8417), .ZN(n8706) );
  OR2_X1 U11074 ( .A1(n8796), .A2(n7368), .ZN(n8705) );
  MUX2_X1 U11075 ( .A(n13980), .B(n14176), .S(n8770), .Z(n8710) );
  MUX2_X1 U11076 ( .A(n13980), .B(n14176), .S(n8788), .Z(n8707) );
  NAND2_X1 U11077 ( .A1(n8708), .A2(n8707), .ZN(n8714) );
  INV_X1 U11078 ( .A(n8709), .ZN(n8712) );
  INV_X1 U11079 ( .A(n8710), .ZN(n8711) );
  NAND2_X1 U11080 ( .A1(n8712), .A2(n8711), .ZN(n8713) );
  NAND2_X1 U11081 ( .A1(n8780), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n8720) );
  INV_X1 U11082 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n15337) );
  OR2_X1 U11083 ( .A1(n8781), .A2(n15337), .ZN(n8719) );
  OAI21_X1 U11084 ( .B1(P1_REG3_REG_25__SCAN_IN), .B2(n8716), .A(n8726), .ZN(
        n13675) );
  OR2_X1 U11085 ( .A1(n8752), .A2(n13675), .ZN(n8718) );
  NAND2_X1 U11086 ( .A1(n8763), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n8717) );
  NAND4_X1 U11087 ( .A1(n8720), .A2(n8719), .A3(n8718), .A4(n8717), .ZN(n13907) );
  NAND2_X1 U11088 ( .A1(n11256), .A2(n8417), .ZN(n8722) );
  OR2_X1 U11089 ( .A1(n8796), .A2(n15297), .ZN(n8721) );
  MUX2_X1 U11090 ( .A(n13907), .B(n14168), .S(n8788), .Z(n8724) );
  MUX2_X1 U11091 ( .A(n13907), .B(n14168), .S(n8770), .Z(n8723) );
  NAND2_X1 U11092 ( .A1(n8780), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n8731) );
  NAND2_X1 U11093 ( .A1(n8763), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n8730) );
  INV_X1 U11094 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n15274) );
  NAND2_X1 U11095 ( .A1(n15274), .A2(n8726), .ZN(n8727) );
  NAND2_X1 U11096 ( .A1(n8748), .A2(n8727), .ZN(n13735) );
  OR2_X1 U11097 ( .A1(n8752), .A2(n13735), .ZN(n8729) );
  NAND2_X1 U11098 ( .A1(n8776), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n8728) );
  NAND4_X1 U11099 ( .A1(n8731), .A2(n8730), .A3(n8729), .A4(n8728), .ZN(n13979) );
  NAND2_X1 U11100 ( .A1(n13486), .A2(n8417), .ZN(n8733) );
  OR2_X1 U11101 ( .A1(n8796), .A2(n14267), .ZN(n8732) );
  MUX2_X1 U11102 ( .A(n13979), .B(n14162), .S(n8770), .Z(n8736) );
  MUX2_X1 U11103 ( .A(n13979), .B(n14162), .S(n8788), .Z(n8734) );
  INV_X1 U11104 ( .A(n8736), .ZN(n8737) );
  NAND2_X1 U11105 ( .A1(n8780), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n8741) );
  NAND2_X1 U11106 ( .A1(n8763), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n8740) );
  NAND2_X1 U11107 ( .A1(n8776), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n8739) );
  INV_X1 U11108 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n13613) );
  XNOR2_X1 U11109 ( .A(n8748), .B(n13613), .ZN(n13954) );
  NAND2_X1 U11110 ( .A1(n13483), .A2(n8417), .ZN(n8743) );
  INV_X1 U11111 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n15217) );
  OR2_X1 U11112 ( .A1(n8796), .A2(n15217), .ZN(n8742) );
  MUX2_X1 U11113 ( .A(n13910), .B(n13956), .S(n8788), .Z(n8746) );
  MUX2_X1 U11114 ( .A(n13910), .B(n13956), .S(n8770), .Z(n8744) );
  NAND2_X1 U11115 ( .A1(n8776), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n8756) );
  NAND2_X1 U11116 ( .A1(n8780), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n8755) );
  NAND2_X1 U11117 ( .A1(n8763), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n8754) );
  INV_X1 U11118 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n8747) );
  OAI21_X1 U11119 ( .B1(n8748), .B2(n13613), .A(n8747), .ZN(n8751) );
  INV_X1 U11120 ( .A(n8748), .ZN(n8750) );
  AND2_X1 U11121 ( .A1(P1_REG3_REG_27__SCAN_IN), .A2(P1_REG3_REG_28__SCAN_IN), 
        .ZN(n8749) );
  NAND2_X1 U11122 ( .A1(n8750), .A2(n8749), .ZN(n13920) );
  NAND2_X1 U11123 ( .A1(n8751), .A2(n13920), .ZN(n13931) );
  OR2_X1 U11124 ( .A1(n8752), .A2(n13931), .ZN(n8753) );
  NAND4_X1 U11125 ( .A1(n8756), .A2(n8755), .A3(n8754), .A4(n8753), .ZN(n13945) );
  OR2_X1 U11126 ( .A1(n8796), .A2(n11639), .ZN(n8757) );
  MUX2_X1 U11127 ( .A(n13945), .B(n14143), .S(n8770), .Z(n8761) );
  MUX2_X1 U11128 ( .A(n13945), .B(n14143), .S(n8788), .Z(n8759) );
  INV_X1 U11129 ( .A(n8761), .ZN(n8762) );
  NAND2_X1 U11130 ( .A1(n8780), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n8767) );
  NAND2_X1 U11131 ( .A1(n8763), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n8766) );
  OR2_X1 U11132 ( .A1(n8752), .A2(n13920), .ZN(n8765) );
  INV_X1 U11133 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n15146) );
  OR2_X1 U11134 ( .A1(n8781), .A2(n15146), .ZN(n8764) );
  NAND4_X1 U11135 ( .A1(n8767), .A2(n8766), .A3(n8765), .A4(n8764), .ZN(n13758) );
  NAND2_X1 U11136 ( .A1(n11636), .A2(n8417), .ZN(n8769) );
  OR2_X1 U11137 ( .A1(n8796), .A2(n11644), .ZN(n8768) );
  MUX2_X1 U11138 ( .A(n13758), .B(n14136), .S(n8788), .Z(n8773) );
  MUX2_X1 U11139 ( .A(n13758), .B(n14136), .S(n8770), .Z(n8771) );
  NAND2_X1 U11140 ( .A1(n8772), .A2(n8771), .ZN(n8775) );
  NAND2_X1 U11141 ( .A1(n6911), .A2(n7152), .ZN(n8774) );
  INV_X1 U11142 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n8779) );
  NAND2_X1 U11143 ( .A1(n8780), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n8778) );
  NAND2_X1 U11144 ( .A1(n8776), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n8777) );
  OAI211_X1 U11145 ( .C1(n8784), .C2(n8779), .A(n8778), .B(n8777), .ZN(n13855)
         );
  INV_X1 U11146 ( .A(n10459), .ZN(n8801) );
  NAND2_X1 U11147 ( .A1(n8801), .A2(n9242), .ZN(n9244) );
  INV_X1 U11148 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n15346) );
  NAND2_X1 U11149 ( .A1(n8780), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n8783) );
  INV_X1 U11150 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n15159) );
  OR2_X1 U11151 ( .A1(n8781), .A2(n15159), .ZN(n8782) );
  OAI211_X1 U11152 ( .C1(n8784), .C2(n15346), .A(n8783), .B(n8782), .ZN(n13919) );
  OAI21_X1 U11153 ( .B1(n13855), .B2(n9244), .A(n13919), .ZN(n8789) );
  INV_X1 U11154 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n11656) );
  OR2_X1 U11155 ( .A1(n8796), .A2(n11656), .ZN(n8786) );
  MUX2_X1 U11156 ( .A(n8789), .B(n14134), .S(n8788), .Z(n8806) );
  INV_X1 U11157 ( .A(n14134), .ZN(n8808) );
  NAND2_X1 U11158 ( .A1(n8808), .A2(n8770), .ZN(n8794) );
  NAND2_X1 U11159 ( .A1(n13855), .A2(n8788), .ZN(n8790) );
  OAI21_X1 U11160 ( .B1(n9242), .B2(n8791), .A(n8790), .ZN(n8792) );
  NAND2_X1 U11161 ( .A1(n8792), .A2(n13919), .ZN(n8793) );
  NAND2_X1 U11162 ( .A1(n8794), .A2(n8793), .ZN(n8805) );
  AND2_X1 U11163 ( .A1(n8806), .A2(n8805), .ZN(n8829) );
  INV_X1 U11164 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n15260) );
  NOR2_X1 U11165 ( .A1(n8796), .A2(n15260), .ZN(n8797) );
  NAND2_X1 U11166 ( .A1(n14128), .A2(n13855), .ZN(n8799) );
  OR2_X1 U11167 ( .A1(n14128), .A2(n13855), .ZN(n8798) );
  MUX2_X1 U11168 ( .A(n8799), .B(n8798), .S(n8788), .Z(n8835) );
  INV_X1 U11169 ( .A(n9246), .ZN(n8879) );
  OR2_X1 U11170 ( .A1(n8879), .A2(n13847), .ZN(n14004) );
  NAND2_X1 U11171 ( .A1(n10459), .A2(n8929), .ZN(n9248) );
  NAND2_X1 U11172 ( .A1(n14271), .A2(n9242), .ZN(n9058) );
  NAND2_X1 U11173 ( .A1(n9248), .A2(n9058), .ZN(n8800) );
  AND2_X1 U11174 ( .A1(n14004), .A2(n8800), .ZN(n8832) );
  INV_X1 U11175 ( .A(n9242), .ZN(n10669) );
  AND2_X1 U11176 ( .A1(n8801), .A2(n10669), .ZN(n8927) );
  NOR2_X1 U11177 ( .A1(n8832), .A2(n8927), .ZN(n8833) );
  NAND2_X1 U11178 ( .A1(n8835), .A2(n8833), .ZN(n8827) );
  INV_X1 U11179 ( .A(n14128), .ZN(n8803) );
  INV_X1 U11180 ( .A(n13855), .ZN(n8802) );
  XNOR2_X1 U11181 ( .A(n8803), .B(n8802), .ZN(n8834) );
  INV_X1 U11182 ( .A(n8834), .ZN(n8804) );
  INV_X1 U11183 ( .A(n8828), .ZN(n8807) );
  NOR2_X1 U11184 ( .A1(n8806), .A2(n8805), .ZN(n8830) );
  XOR2_X1 U11185 ( .A(n13919), .B(n8808), .Z(n8825) );
  NAND2_X1 U11186 ( .A1(n14143), .A2(n13945), .ZN(n13912) );
  INV_X1 U11187 ( .A(n13979), .ZN(n8810) );
  NAND2_X1 U11188 ( .A1(n14162), .A2(n8810), .ZN(n13941) );
  OR2_X1 U11189 ( .A1(n14162), .A2(n8810), .ZN(n8811) );
  INV_X1 U11190 ( .A(n13980), .ZN(n13881) );
  XNOR2_X1 U11191 ( .A(n14176), .B(n13881), .ZN(n13998) );
  INV_X1 U11192 ( .A(n14026), .ZN(n13879) );
  XNOR2_X1 U11193 ( .A(n14181), .B(n13879), .ZN(n13903) );
  XNOR2_X1 U11194 ( .A(n14033), .B(n13900), .ZN(n14034) );
  NAND2_X1 U11195 ( .A1(n14190), .A2(n14025), .ZN(n8812) );
  NAND2_X1 U11196 ( .A1(n13899), .A2(n8812), .ZN(n14049) );
  NAND2_X1 U11197 ( .A1(n11389), .A2(n8813), .ZN(n11387) );
  INV_X1 U11198 ( .A(n13761), .ZN(n11218) );
  XNOR2_X1 U11199 ( .A(n11253), .B(n11218), .ZN(n11151) );
  INV_X1 U11200 ( .A(n13762), .ZN(n10809) );
  OR2_X1 U11201 ( .A1(n13667), .A2(n10809), .ZN(n11149) );
  NAND2_X1 U11202 ( .A1(n13667), .A2(n10809), .ZN(n8814) );
  NAND2_X1 U11203 ( .A1(n11149), .A2(n8814), .ZN(n10858) );
  OR2_X1 U11204 ( .A1(n11018), .A2(n13763), .ZN(n10868) );
  NAND2_X1 U11205 ( .A1(n11018), .A2(n13763), .ZN(n10871) );
  NAND2_X1 U11206 ( .A1(n10868), .A2(n10871), .ZN(n10814) );
  INV_X1 U11207 ( .A(n13766), .ZN(n10498) );
  XNOR2_X1 U11208 ( .A(n10600), .B(n10498), .ZN(n10512) );
  XNOR2_X1 U11209 ( .A(n14517), .B(n13767), .ZN(n10310) );
  NAND4_X1 U11210 ( .A1(n9761), .A2(n9757), .A3(n9895), .A4(n14557), .ZN(n8815) );
  XNOR2_X1 U11211 ( .A(n14608), .B(n8944), .ZN(n9860) );
  NOR2_X1 U11212 ( .A1(n8815), .A2(n9852), .ZN(n8816) );
  XNOR2_X1 U11213 ( .A(n14530), .B(n13769), .ZN(n9857) );
  XNOR2_X1 U11214 ( .A(n10315), .B(n13768), .ZN(n10305) );
  NAND4_X1 U11215 ( .A1(n10310), .A2(n8816), .A3(n9857), .A4(n10305), .ZN(
        n8817) );
  NOR2_X1 U11216 ( .A1(n10512), .A2(n8817), .ZN(n8818) );
  XNOR2_X1 U11217 ( .A(n14635), .B(n13764), .ZN(n10504) );
  XNOR2_X1 U11218 ( .A(n14500), .B(n13765), .ZN(n14491) );
  NAND4_X1 U11219 ( .A1(n10814), .A2(n8818), .A3(n10504), .A4(n14491), .ZN(
        n8819) );
  OR4_X1 U11220 ( .A1(n11221), .A2(n11151), .A3(n10858), .A4(n8819), .ZN(n8820) );
  NOR2_X1 U11221 ( .A1(n11387), .A2(n8820), .ZN(n8821) );
  XNOR2_X1 U11222 ( .A(n13890), .B(n14106), .ZN(n11398) );
  NAND2_X1 U11223 ( .A1(n14218), .A2(n14088), .ZN(n13893) );
  NAND2_X1 U11224 ( .A1(n6588), .A2(n13893), .ZN(n14121) );
  NAND4_X1 U11225 ( .A1(n14049), .A2(n8821), .A3(n11398), .A4(n14121), .ZN(
        n8822) );
  INV_X1 U11226 ( .A(n14070), .ZN(n14068) );
  INV_X1 U11227 ( .A(n14091), .ZN(n14086) );
  XNOR2_X1 U11228 ( .A(n14197), .B(n14074), .ZN(n14063) );
  NOR4_X1 U11229 ( .A1(n8834), .A2(n8825), .A3(n13913), .A4(n6636), .ZN(n8826)
         );
  XNOR2_X1 U11230 ( .A(n8826), .B(n8928), .ZN(n8841) );
  INV_X1 U11231 ( .A(n8927), .ZN(n8840) );
  INV_X1 U11232 ( .A(n8827), .ZN(n8831) );
  AOI22_X1 U11233 ( .A1(n8831), .A2(n8830), .B1(n8829), .B2(n8828), .ZN(n8839)
         );
  INV_X1 U11234 ( .A(n8832), .ZN(n8837) );
  NAND2_X1 U11235 ( .A1(n8834), .A2(n8833), .ZN(n8836) );
  MUX2_X1 U11236 ( .A(n8837), .B(n8836), .S(n8835), .Z(n8838) );
  OAI211_X1 U11237 ( .C1(n8841), .C2(n8840), .A(n8839), .B(n8838), .ZN(n8842)
         );
  NAND2_X1 U11238 ( .A1(n8844), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8845) );
  XNOR2_X1 U11239 ( .A(n8845), .B(n8847), .ZN(n8939) );
  INV_X1 U11240 ( .A(n8939), .ZN(n9057) );
  NAND2_X1 U11241 ( .A1(n9057), .A2(P1_STATE_REG_SCAN_IN), .ZN(n11007) );
  NAND2_X1 U11242 ( .A1(n6791), .A2(n8847), .ZN(n8849) );
  NAND2_X1 U11243 ( .A1(n8852), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8848) );
  XNOR2_X1 U11244 ( .A(n8848), .B(P1_IR_REG_25__SCAN_IN), .ZN(n9052) );
  NAND2_X1 U11245 ( .A1(n8849), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8850) );
  MUX2_X1 U11246 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8850), .S(
        P1_IR_REG_24__SCAN_IN), .Z(n8851) );
  NAND2_X2 U11247 ( .A1(n8854), .A2(n14265), .ZN(n8936) );
  NAND2_X1 U11248 ( .A1(n10459), .A2(n13847), .ZN(n8855) );
  INV_X1 U11249 ( .A(n9058), .ZN(n8931) );
  NAND2_X1 U11250 ( .A1(n8855), .A2(n8931), .ZN(n8937) );
  AND2_X1 U11251 ( .A1(n9056), .A2(n8937), .ZN(n9656) );
  INV_X1 U11252 ( .A(n14264), .ZN(n14442) );
  INV_X1 U11253 ( .A(n11640), .ZN(n9128) );
  NAND3_X1 U11254 ( .A1(n9656), .A2(n14442), .A3(n14107), .ZN(n8856) );
  OAI211_X1 U11255 ( .C1(n14271), .C2(n11007), .A(n8856), .B(P1_B_REG_SCAN_IN), 
        .ZN(n8857) );
  INV_X1 U11256 ( .A(n9553), .ZN(n8858) );
  AND2_X1 U11257 ( .A1(n8858), .A2(n11011), .ZN(n9272) );
  NAND2_X1 U11258 ( .A1(n9003), .A2(n8859), .ZN(n9014) );
  NOR2_X1 U11259 ( .A1(P3_IR_REG_22__SCAN_IN), .A2(P3_IR_REG_21__SCAN_IN), 
        .ZN(n8868) );
  NOR2_X1 U11260 ( .A1(P3_IR_REG_18__SCAN_IN), .A2(P3_IR_REG_17__SCAN_IN), 
        .ZN(n8867) );
  NAND4_X1 U11261 ( .A1(n8868), .A2(n8867), .A3(n9700), .A4(n9682), .ZN(n8869)
         );
  NAND2_X1 U11262 ( .A1(n8872), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8870) );
  XNOR2_X1 U11263 ( .A(n8870), .B(P3_IR_REG_25__SCAN_IN), .ZN(n9091) );
  NAND2_X1 U11264 ( .A1(n8876), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8871) );
  XNOR2_X1 U11265 ( .A(n8871), .B(P3_IR_REG_24__SCAN_IN), .ZN(n9092) );
  NAND2_X1 U11266 ( .A1(n9091), .A2(n9092), .ZN(n8874) );
  NAND2_X1 U11267 ( .A1(n6702), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8875) );
  MUX2_X1 U11268 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8875), .S(
        P3_IR_REG_23__SCAN_IN), .Z(n8877) );
  NAND2_X1 U11269 ( .A1(n8877), .A2(n8876), .ZN(n9877) );
  INV_X1 U11270 ( .A(n9800), .ZN(n8878) );
  INV_X1 U11271 ( .A(n9187), .ZN(n9051) );
  OR2_X2 U11272 ( .A1(n8936), .A2(n9051), .ZN(n13773) );
  INV_X1 U11273 ( .A(n13773), .ZN(P1_U4016) );
  NAND2_X1 U11274 ( .A1(n14556), .A2(n6536), .ZN(n8881) );
  AND2_X2 U11275 ( .A1(n8879), .A2(n8936), .ZN(n13640) );
  NAND2_X1 U11276 ( .A1(n13640), .A2(n6539), .ZN(n8880) );
  NAND2_X1 U11277 ( .A1(n8881), .A2(n8880), .ZN(n8882) );
  AND2_X1 U11278 ( .A1(n14271), .A2(n13847), .ZN(n9245) );
  OR2_X2 U11279 ( .A1(n9246), .A2(n9245), .ZN(n13637) );
  XNOR2_X1 U11280 ( .A(n8882), .B(n13637), .ZN(n8889) );
  AND2_X1 U11281 ( .A1(n6539), .A2(n6536), .ZN(n8883) );
  AOI21_X1 U11282 ( .B1(n14556), .B2(n13603), .A(n8883), .ZN(n8890) );
  XNOR2_X1 U11283 ( .A(n8889), .B(n8890), .ZN(n9296) );
  OAI22_X1 U11284 ( .A1(n9669), .A2(n13549), .B1(n8936), .B2(n14445), .ZN(
        n8884) );
  AOI21_X1 U11285 ( .B1(n8344), .B2(n13603), .A(n8884), .ZN(n9191) );
  NAND2_X1 U11286 ( .A1(n8344), .A2(n6536), .ZN(n8887) );
  INV_X1 U11287 ( .A(n8936), .ZN(n8885) );
  AOI22_X1 U11288 ( .A1(n14553), .A2(n13640), .B1(n8885), .B2(
        P1_REG1_REG_0__SCAN_IN), .ZN(n8886) );
  NAND2_X1 U11289 ( .A1(n8887), .A2(n8886), .ZN(n9190) );
  NAND2_X1 U11290 ( .A1(n9191), .A2(n9190), .ZN(n9189) );
  OR2_X1 U11291 ( .A1(n9190), .A2(n13591), .ZN(n8888) );
  NAND2_X1 U11292 ( .A1(n9189), .A2(n8888), .ZN(n9295) );
  NAND2_X1 U11293 ( .A1(n9296), .A2(n9295), .ZN(n8893) );
  INV_X1 U11294 ( .A(n8889), .ZN(n8891) );
  NAND2_X1 U11295 ( .A1(n8891), .A2(n8890), .ZN(n8892) );
  NAND2_X1 U11296 ( .A1(n8893), .A2(n8892), .ZN(n9402) );
  NAND2_X1 U11297 ( .A1(n13772), .A2(n6536), .ZN(n8895) );
  NAND2_X1 U11298 ( .A1(n14589), .A2(n13640), .ZN(n8894) );
  NAND2_X1 U11299 ( .A1(n8895), .A2(n8894), .ZN(n8896) );
  XNOR2_X1 U11300 ( .A(n8896), .B(n13591), .ZN(n8901) );
  NAND2_X1 U11301 ( .A1(n13772), .A2(n13603), .ZN(n8898) );
  NAND2_X1 U11302 ( .A1(n14589), .A2(n6536), .ZN(n8897) );
  NAND2_X1 U11303 ( .A1(n8898), .A2(n8897), .ZN(n8899) );
  XNOR2_X1 U11304 ( .A(n8901), .B(n8899), .ZN(n9401) );
  NAND2_X1 U11305 ( .A1(n9402), .A2(n9401), .ZN(n8903) );
  INV_X1 U11306 ( .A(n8899), .ZN(n8900) );
  NAND2_X1 U11307 ( .A1(n8901), .A2(n8900), .ZN(n8902) );
  INV_X1 U11308 ( .A(n13640), .ZN(n9939) );
  INV_X2 U11309 ( .A(n13639), .ZN(n13549) );
  OAI22_X1 U11310 ( .A1(n14599), .A2(n9939), .B1(n9753), .B2(n13549), .ZN(
        n8904) );
  XNOR2_X1 U11311 ( .A(n8904), .B(n13637), .ZN(n8905) );
  OAI22_X1 U11312 ( .A1(n14599), .A2(n13549), .B1(n9753), .B2(n13548), .ZN(
        n8906) );
  NAND2_X1 U11313 ( .A1(n8905), .A2(n8906), .ZN(n9838) );
  INV_X1 U11314 ( .A(n8905), .ZN(n8908) );
  INV_X1 U11315 ( .A(n8906), .ZN(n8907) );
  NAND2_X1 U11316 ( .A1(n8908), .A2(n8907), .ZN(n8909) );
  NAND2_X1 U11317 ( .A1(n9838), .A2(n8909), .ZN(n8934) );
  INV_X1 U11318 ( .A(n9052), .ZN(n11259) );
  NAND3_X1 U11319 ( .A1(n11259), .A2(P1_B_REG_SCAN_IN), .A3(n11225), .ZN(n8910) );
  OR2_X1 U11320 ( .A1(n9356), .A2(P1_D_REG_1__SCAN_IN), .ZN(n8912) );
  OR2_X1 U11321 ( .A1(n14265), .A2(n9052), .ZN(n8911) );
  NOR4_X1 U11322 ( .A1(P1_D_REG_16__SCAN_IN), .A2(P1_D_REG_17__SCAN_IN), .A3(
        P1_D_REG_19__SCAN_IN), .A4(P1_D_REG_20__SCAN_IN), .ZN(n8916) );
  NOR4_X1 U11323 ( .A1(P1_D_REG_14__SCAN_IN), .A2(P1_D_REG_12__SCAN_IN), .A3(
        P1_D_REG_13__SCAN_IN), .A4(P1_D_REG_15__SCAN_IN), .ZN(n8915) );
  NOR4_X1 U11324 ( .A1(P1_D_REG_25__SCAN_IN), .A2(P1_D_REG_26__SCAN_IN), .A3(
        P1_D_REG_27__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n8914) );
  NOR4_X1 U11325 ( .A1(P1_D_REG_21__SCAN_IN), .A2(P1_D_REG_22__SCAN_IN), .A3(
        P1_D_REG_23__SCAN_IN), .A4(P1_D_REG_24__SCAN_IN), .ZN(n8913) );
  AND4_X1 U11326 ( .A1(n8916), .A2(n8915), .A3(n8914), .A4(n8913), .ZN(n8922)
         );
  NOR2_X1 U11327 ( .A1(P1_D_REG_18__SCAN_IN), .A2(P1_D_REG_28__SCAN_IN), .ZN(
        n8920) );
  NOR4_X1 U11328 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        P1_D_REG_11__SCAN_IN), .A4(P1_D_REG_2__SCAN_IN), .ZN(n8919) );
  NOR4_X1 U11329 ( .A1(P1_D_REG_7__SCAN_IN), .A2(P1_D_REG_8__SCAN_IN), .A3(
        P1_D_REG_9__SCAN_IN), .A4(P1_D_REG_10__SCAN_IN), .ZN(n8918) );
  NOR4_X1 U11330 ( .A1(P1_D_REG_3__SCAN_IN), .A2(P1_D_REG_4__SCAN_IN), .A3(
        P1_D_REG_5__SCAN_IN), .A4(P1_D_REG_6__SCAN_IN), .ZN(n8917) );
  AND4_X1 U11331 ( .A1(n8920), .A2(n8919), .A3(n8918), .A4(n8917), .ZN(n8921)
         );
  NAND2_X1 U11332 ( .A1(n8922), .A2(n8921), .ZN(n9354) );
  INV_X1 U11333 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n15290) );
  NOR2_X1 U11334 ( .A1(n9354), .A2(n15290), .ZN(n8923) );
  OR2_X1 U11335 ( .A1(n9356), .A2(n8923), .ZN(n8925) );
  OR2_X1 U11336 ( .A1(n8924), .A2(n14265), .ZN(n9353) );
  NAND2_X1 U11337 ( .A1(n9655), .A2(n9253), .ZN(n8946) );
  INV_X1 U11338 ( .A(n8946), .ZN(n8926) );
  NAND2_X1 U11339 ( .A1(n8926), .A2(n9056), .ZN(n8941) );
  NAND2_X1 U11340 ( .A1(n8927), .A2(n8929), .ZN(n9664) );
  NAND3_X1 U11341 ( .A1(n8929), .A2(n8928), .A3(n10669), .ZN(n8930) );
  OR2_X1 U11342 ( .A1(n14607), .A2(n8931), .ZN(n8932) );
  INV_X1 U11343 ( .A(n9839), .ZN(n8933) );
  AOI211_X1 U11344 ( .C1(n8935), .C2(n8934), .A(n13756), .B(n8933), .ZN(n8949)
         );
  NAND2_X1 U11345 ( .A1(n8937), .A2(n8936), .ZN(n8938) );
  AOI21_X1 U11346 ( .B1(n8946), .B2(n9251), .A(n8938), .ZN(n9188) );
  NAND2_X1 U11347 ( .A1(n9188), .A2(n8939), .ZN(n8940) );
  MUX2_X1 U11348 ( .A(n13740), .B(P1_U3086), .S(P1_REG3_REG_3__SCAN_IN), .Z(
        n8948) );
  OR2_X1 U11349 ( .A1(n8941), .A2(n9664), .ZN(n8943) );
  INV_X1 U11350 ( .A(n9251), .ZN(n8942) );
  AOI22_X1 U11351 ( .A1(n14108), .A2(n8944), .B1(n13772), .B2(n14107), .ZN(
        n14539) );
  INV_X1 U11352 ( .A(n9656), .ZN(n8945) );
  NOR2_X2 U11353 ( .A1(n8946), .A2(n8945), .ZN(n14397) );
  INV_X1 U11354 ( .A(n14397), .ZN(n13738) );
  OAI22_X1 U11355 ( .A1(n13743), .A2(n14599), .B1(n14539), .B2(n13738), .ZN(
        n8947) );
  OR3_X1 U11356 ( .A1(n8949), .A2(n8948), .A3(n8947), .ZN(P1_U3218) );
  AND2_X1 U11357 ( .A1(n7499), .A2(P1_U3086), .ZN(n11006) );
  OAI222_X1 U11358 ( .A1(P1_U3086), .A2(n13778), .B1(n6535), .B2(n8951), .C1(
        n8950), .C2(n14266), .ZN(P1_U3354) );
  AND2_X1 U11359 ( .A1(n9727), .A2(P2_U3088), .ZN(n11009) );
  NOR2_X1 U11360 ( .A1(n9727), .A2(P2_STATE_REG_SCAN_IN), .ZN(n13480) );
  INV_X2 U11361 ( .A(n13480), .ZN(n11904) );
  OAI222_X1 U11362 ( .A1(P2_U3088), .A2(n13058), .B1(n6534), .B2(n8951), .C1(
        n8963), .C2(n11904), .ZN(P2_U3326) );
  INV_X1 U11363 ( .A(n13068), .ZN(n8953) );
  INV_X1 U11364 ( .A(n8952), .ZN(n8989) );
  OAI222_X1 U11365 ( .A1(P2_U3088), .A2(n8953), .B1(n6534), .B2(n8989), .C1(
        n8967), .C2(n11904), .ZN(P2_U3325) );
  NOR2_X1 U11366 ( .A1(n9727), .A2(P3_STATE_REG_SCAN_IN), .ZN(n12881) );
  INV_X1 U11367 ( .A(n12881), .ZN(n12245) );
  XNOR2_X1 U11368 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .ZN(n8962) );
  XNOR2_X1 U11369 ( .A(n8962), .B(n9041), .ZN(n9801) );
  INV_X1 U11370 ( .A(SI_1_), .ZN(n15202) );
  INV_X1 U11371 ( .A(P3_IR_REG_1__SCAN_IN), .ZN(n10038) );
  OAI222_X1 U11372 ( .A1(n12245), .A2(n9801), .B1(n11338), .B2(n15202), .C1(
        P3_U3151), .C2(n9999), .ZN(P3_U3294) );
  INV_X1 U11373 ( .A(P3_IR_REG_5__SCAN_IN), .ZN(n8957) );
  NAND2_X1 U11374 ( .A1(n9034), .A2(n8957), .ZN(n9026) );
  NOR2_X1 U11375 ( .A1(n8997), .A2(P3_IR_REG_7__SCAN_IN), .ZN(n8959) );
  OR2_X1 U11376 ( .A1(n8959), .A2(n9718), .ZN(n8958) );
  MUX2_X1 U11377 ( .A(n8958), .B(P3_IR_REG_31__SCAN_IN), .S(n6986), .Z(n8960)
         );
  NAND2_X1 U11378 ( .A1(n8959), .A2(n6986), .ZN(n9022) );
  INV_X1 U11379 ( .A(SI_8_), .ZN(n10527) );
  INV_X1 U11380 ( .A(n9041), .ZN(n8961) );
  NAND2_X1 U11381 ( .A1(n8962), .A2(n8961), .ZN(n8965) );
  NAND2_X1 U11382 ( .A1(n8963), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n8964) );
  NAND2_X1 U11383 ( .A1(n8965), .A2(n8964), .ZN(n9002) );
  NAND2_X1 U11384 ( .A1(n8988), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n8966) );
  NAND2_X1 U11385 ( .A1(n9002), .A2(n8966), .ZN(n8969) );
  NAND2_X1 U11386 ( .A1(n8967), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n8968) );
  NAND2_X1 U11387 ( .A1(n8991), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n8971) );
  INV_X1 U11388 ( .A(n9006), .ZN(n8972) );
  INV_X1 U11389 ( .A(n9029), .ZN(n8974) );
  NAND2_X1 U11390 ( .A1(n9066), .A2(P1_DATAO_REG_5__SCAN_IN), .ZN(n8975) );
  NAND2_X1 U11391 ( .A1(n9071), .A2(P1_DATAO_REG_6__SCAN_IN), .ZN(n8977) );
  XNOR2_X1 U11392 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(P2_DATAO_REG_8__SCAN_IN), 
        .ZN(n8981) );
  XNOR2_X1 U11393 ( .A(n9018), .B(n8981), .ZN(n10526) );
  OAI222_X1 U11394 ( .A1(P3_U3151), .A2(n14928), .B1(n11338), .B2(n10527), 
        .C1(n12245), .C2(n10526), .ZN(P3_U3287) );
  NAND2_X1 U11395 ( .A1(n9026), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8983) );
  XNOR2_X1 U11396 ( .A(n8983), .B(n8982), .ZN(n14893) );
  XNOR2_X1 U11397 ( .A(n8985), .B(n8984), .ZN(n10376) );
  INV_X1 U11398 ( .A(SI_6_), .ZN(n10375) );
  OAI222_X1 U11399 ( .A1(P3_U3151), .A2(n14893), .B1(n12245), .B2(n10376), 
        .C1(n10375), .C2(n11338), .ZN(P3_U3289) );
  INV_X1 U11400 ( .A(n13081), .ZN(n13074) );
  INV_X1 U11401 ( .A(n8986), .ZN(n8992) );
  OAI222_X1 U11402 ( .A1(P2_U3088), .A2(n13074), .B1(n6534), .B2(n8992), .C1(
        n8987), .C2(n11904), .ZN(P2_U3324) );
  INV_X1 U11403 ( .A(n13797), .ZN(n8990) );
  OAI222_X1 U11404 ( .A1(P1_U3086), .A2(n8990), .B1(n6535), .B2(n8989), .C1(
        n8988), .C2(n14266), .ZN(P1_U3353) );
  INV_X1 U11405 ( .A(n13808), .ZN(n9117) );
  OAI222_X1 U11406 ( .A1(P1_U3086), .A2(n9117), .B1(n6535), .B2(n8992), .C1(
        n8991), .C2(n14266), .ZN(P1_U3352) );
  INV_X1 U11407 ( .A(n14266), .ZN(n14260) );
  AOI22_X1 U11408 ( .A1(n9232), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_4__SCAN_IN), .B2(n14260), .ZN(n8994) );
  OAI21_X1 U11409 ( .B1(n8993), .B2(n6535), .A(n8994), .ZN(P1_U3351) );
  XNOR2_X1 U11410 ( .A(n8996), .B(n8995), .ZN(n10521) );
  NAND2_X1 U11411 ( .A1(n8997), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8999) );
  INV_X1 U11412 ( .A(P3_IR_REG_7__SCAN_IN), .ZN(n8998) );
  XNOR2_X1 U11413 ( .A(n8999), .B(n8998), .ZN(n14911) );
  INV_X1 U11414 ( .A(n14911), .ZN(n10941) );
  INV_X1 U11415 ( .A(n11338), .ZN(n10122) );
  AOI222_X1 U11416 ( .A1(n10521), .A2(n12881), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n10941), .C1(SI_7_), .C2(n10122), .ZN(n9000) );
  INV_X1 U11417 ( .A(n9000), .ZN(P3_U3288) );
  XNOR2_X1 U11418 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(P2_DATAO_REG_2__SCAN_IN), 
        .ZN(n9001) );
  XNOR2_X1 U11419 ( .A(n9002), .B(n9001), .ZN(n9962) );
  AOI222_X1 U11420 ( .A1(n9962), .A2(n12881), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n10046), .C1(SI_2_), .C2(n10122), .ZN(n9005) );
  INV_X1 U11421 ( .A(n9005), .ZN(P3_U3293) );
  XNOR2_X1 U11422 ( .A(n9007), .B(n9006), .ZN(n10194) );
  INV_X1 U11423 ( .A(n9034), .ZN(n9010) );
  NAND2_X1 U11424 ( .A1(n8956), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9008) );
  MUX2_X1 U11425 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9008), .S(
        P3_IR_REG_4__SCAN_IN), .Z(n9009) );
  INV_X1 U11426 ( .A(n14857), .ZN(n10922) );
  AOI222_X1 U11427 ( .A1(n10194), .A2(n12881), .B1(n10922), .B2(
        P3_STATE_REG_SCAN_IN), .C1(SI_4_), .C2(n10122), .ZN(n9011) );
  INV_X1 U11428 ( .A(n9011), .ZN(P3_U3291) );
  XNOR2_X1 U11429 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(P2_DATAO_REG_3__SCAN_IN), 
        .ZN(n9012) );
  XNOR2_X1 U11430 ( .A(n9013), .B(n9012), .ZN(n10002) );
  NAND2_X1 U11431 ( .A1(n9014), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9015) );
  MUX2_X1 U11432 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9015), .S(
        P3_IR_REG_3__SCAN_IN), .Z(n9016) );
  AOI222_X1 U11433 ( .A1(n10002), .A2(n12881), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n14842), .C1(SI_3_), .C2(n10122), .ZN(n9017) );
  INV_X1 U11434 ( .A(n9017), .ZN(P3_U3292) );
  NAND2_X1 U11435 ( .A1(n9096), .A2(P2_DATAO_REG_8__SCAN_IN), .ZN(n9019) );
  XNOR2_X1 U11436 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(P2_DATAO_REG_9__SCAN_IN), 
        .ZN(n9021) );
  XNOR2_X1 U11437 ( .A(n9037), .B(n9021), .ZN(n10553) );
  NAND2_X1 U11438 ( .A1(n9022), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9023) );
  XNOR2_X1 U11439 ( .A(n9023), .B(n6985), .ZN(n14946) );
  INV_X1 U11440 ( .A(n14946), .ZN(n10954) );
  AOI222_X1 U11441 ( .A1(n10553), .A2(n12881), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n10954), .C1(SI_9_), .C2(n10122), .ZN(n9024) );
  INV_X1 U11442 ( .A(n9024), .ZN(P3_U3286) );
  NOR2_X1 U11443 ( .A1(n9034), .A2(n9718), .ZN(n9025) );
  MUX2_X1 U11444 ( .A(n9718), .B(n9025), .S(P3_IR_REG_5__SCAN_IN), .Z(n9028)
         );
  INV_X1 U11445 ( .A(n9026), .ZN(n9027) );
  XNOR2_X1 U11446 ( .A(n9030), .B(n9029), .ZN(n10258) );
  AOI222_X1 U11447 ( .A1(n7024), .A2(P3_STATE_REG_SCAN_IN), .B1(n10258), .B2(
        n12881), .C1(SI_5_), .C2(n10122), .ZN(n9031) );
  INV_X1 U11448 ( .A(n9031), .ZN(P3_U3290) );
  INV_X1 U11449 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n9032) );
  OAI222_X1 U11450 ( .A1(P2_U3088), .A2(n14660), .B1(n6534), .B2(n8993), .C1(
        n9032), .C2(n11904), .ZN(P2_U3323) );
  NAND2_X1 U11451 ( .A1(n9034), .A2(n9033), .ZN(n9042) );
  NAND2_X1 U11452 ( .A1(n9042), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9036) );
  INV_X1 U11453 ( .A(P3_IR_REG_10__SCAN_IN), .ZN(n9035) );
  XNOR2_X1 U11454 ( .A(n9036), .B(n9035), .ZN(n14965) );
  NAND2_X1 U11455 ( .A1(n9172), .A2(P1_DATAO_REG_9__SCAN_IN), .ZN(n9038) );
  XNOR2_X1 U11456 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(P2_DATAO_REG_10__SCAN_IN), 
        .ZN(n9045) );
  XNOR2_X1 U11457 ( .A(n9046), .B(n9045), .ZN(n10565) );
  OAI222_X1 U11458 ( .A1(P3_U3151), .A2(n14965), .B1(n11338), .B2(n9039), .C1(
        n12245), .C2(n10565), .ZN(P3_U3285) );
  NAND2_X1 U11459 ( .A1(n15304), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n9040) );
  AND2_X1 U11460 ( .A1(n9041), .A2(n9040), .ZN(n9730) );
  OAI222_X1 U11461 ( .A1(P3_U3151), .A2(n9883), .B1(n12245), .B2(n9730), .C1(
        n9728), .C2(n11338), .ZN(P3_U3295) );
  OR2_X1 U11462 ( .A1(n9042), .A2(P3_IR_REG_10__SCAN_IN), .ZN(n9080) );
  NAND2_X1 U11463 ( .A1(n9080), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9044) );
  INV_X1 U11464 ( .A(P3_IR_REG_11__SCAN_IN), .ZN(n9043) );
  XNOR2_X1 U11465 ( .A(n9044), .B(n9043), .ZN(n11132) );
  INV_X1 U11466 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n9047) );
  NAND2_X1 U11467 ( .A1(n9047), .A2(P1_DATAO_REG_10__SCAN_IN), .ZN(n9048) );
  XNOR2_X1 U11468 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(P2_DATAO_REG_11__SCAN_IN), 
        .ZN(n9050) );
  XNOR2_X1 U11469 ( .A(n9073), .B(n9050), .ZN(n11069) );
  OAI222_X1 U11470 ( .A1(P3_U3151), .A2(n11132), .B1(n11338), .B2(n11070), 
        .C1(n12245), .C2(n11069), .ZN(P3_U3284) );
  NAND2_X1 U11471 ( .A1(n9056), .A2(n9356), .ZN(n14579) );
  INV_X1 U11472 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n9054) );
  NOR3_X1 U11473 ( .A1(n14265), .A2(n9052), .A3(n9051), .ZN(n9053) );
  AOI21_X1 U11474 ( .B1(n14579), .B2(n9054), .A(n9053), .ZN(P1_U3446) );
  INV_X1 U11475 ( .A(n9353), .ZN(n9055) );
  AOI22_X1 U11476 ( .A1(n14579), .A2(n15290), .B1(n9187), .B2(n9055), .ZN(
        P1_U3445) );
  OR2_X1 U11477 ( .A1(n9058), .A2(n9057), .ZN(n9060) );
  AND2_X1 U11478 ( .A1(n9060), .A2(n9059), .ZN(n9112) );
  INV_X1 U11479 ( .A(n9112), .ZN(n9061) );
  AND2_X1 U11480 ( .A1(n9113), .A2(n9061), .ZN(n14472) );
  NOR2_X1 U11481 ( .A1(n14472), .A2(P1_U4016), .ZN(P1_U3085) );
  INV_X1 U11482 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n9064) );
  INV_X1 U11483 ( .A(n9062), .ZN(n9065) );
  INV_X1 U11484 ( .A(n14681), .ZN(n9063) );
  OAI222_X1 U11485 ( .A1(n11904), .A2(n9064), .B1(n6534), .B2(n9065), .C1(
        P2_U3088), .C2(n9063), .ZN(P2_U3322) );
  INV_X1 U11486 ( .A(n9164), .ZN(n9120) );
  OAI222_X1 U11487 ( .A1(n14266), .A2(n9066), .B1(n6535), .B2(n9065), .C1(
        n9120), .C2(P1_U3086), .ZN(P1_U3350) );
  INV_X1 U11488 ( .A(n9370), .ZN(n9069) );
  INV_X1 U11489 ( .A(n9067), .ZN(n9070) );
  OAI222_X1 U11490 ( .A1(P2_U3088), .A2(n9069), .B1(n6534), .B2(n9070), .C1(
        n9068), .C2(n11904), .ZN(P2_U3321) );
  INV_X1 U11491 ( .A(n9121), .ZN(n9183) );
  OAI222_X1 U11492 ( .A1(n14266), .A2(n9071), .B1(n6535), .B2(n9070), .C1(
        P1_U3086), .C2(n9183), .ZN(P1_U3349) );
  AND2_X1 U11493 ( .A1(n9398), .A2(P1_DATAO_REG_11__SCAN_IN), .ZN(n9072) );
  NAND2_X1 U11494 ( .A1(n15272), .A2(P2_DATAO_REG_11__SCAN_IN), .ZN(n9074) );
  NAND2_X1 U11495 ( .A1(n9512), .A2(P1_DATAO_REG_12__SCAN_IN), .ZN(n9152) );
  INV_X1 U11496 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n9511) );
  NAND2_X1 U11497 ( .A1(n9511), .A2(P2_DATAO_REG_12__SCAN_IN), .ZN(n9076) );
  NAND2_X1 U11498 ( .A1(n9152), .A2(n9076), .ZN(n9077) );
  NAND2_X1 U11499 ( .A1(n9078), .A2(n9077), .ZN(n9079) );
  AND2_X1 U11500 ( .A1(n9153), .A2(n9079), .ZN(n11074) );
  INV_X1 U11501 ( .A(n11074), .ZN(n9084) );
  OAI21_X1 U11502 ( .B1(n9080), .B2(P3_IR_REG_11__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n9081) );
  MUX2_X1 U11503 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9081), .S(
        P3_IR_REG_12__SCAN_IN), .Z(n9083) );
  INV_X1 U11504 ( .A(n12360), .ZN(n11123) );
  OAI222_X1 U11505 ( .A1(n11338), .A2(n15330), .B1(n12245), .B2(n9084), .C1(
        n11123), .C2(P3_U3151), .ZN(P3_U3283) );
  INV_X1 U11506 ( .A(n13096), .ZN(n13090) );
  OAI222_X1 U11507 ( .A1(P2_U3088), .A2(n13090), .B1(n6534), .B2(n9086), .C1(
        n9085), .C2(n11904), .ZN(P2_U3320) );
  INV_X1 U11508 ( .A(n9211), .ZN(n9209) );
  OAI222_X1 U11509 ( .A1(P1_U3086), .A2(n9209), .B1(n6535), .B2(n9086), .C1(
        n7353), .C2(n14266), .ZN(P1_U3348) );
  INV_X1 U11510 ( .A(n11005), .ZN(n9089) );
  XNOR2_X1 U11511 ( .A(n9092), .B(P3_B_REG_SCAN_IN), .ZN(n9087) );
  INV_X1 U11512 ( .A(P3_D_REG_1__SCAN_IN), .ZN(n9687) );
  INV_X1 U11513 ( .A(n9091), .ZN(n10886) );
  AND2_X1 U11514 ( .A1(n10886), .A2(n11005), .ZN(n9686) );
  AOI22_X1 U11515 ( .A1(n9156), .A2(n9687), .B1(n9800), .B2(n9686), .ZN(
        P3_U3377) );
  INV_X1 U11516 ( .A(P3_D_REG_0__SCAN_IN), .ZN(n15180) );
  INV_X1 U11517 ( .A(n9092), .ZN(n10793) );
  NAND2_X1 U11518 ( .A1(n11005), .A2(n10793), .ZN(n9688) );
  INV_X1 U11519 ( .A(n9688), .ZN(n9093) );
  AOI22_X1 U11520 ( .A1(n9156), .A2(n15180), .B1(n9093), .B2(n9800), .ZN(
        P3_U3376) );
  INV_X1 U11521 ( .A(n9140), .ZN(n9095) );
  OAI222_X1 U11522 ( .A1(P1_U3086), .A2(n9095), .B1(n6535), .B2(n9097), .C1(
        n9094), .C2(n14266), .ZN(P1_U3347) );
  INV_X1 U11523 ( .A(n13111), .ZN(n9098) );
  OAI222_X1 U11524 ( .A1(P2_U3088), .A2(n9098), .B1(n6534), .B2(n9097), .C1(
        n9096), .C2(n11904), .ZN(P2_U3319) );
  AND2_X1 U11525 ( .A1(n9156), .A2(P3_D_REG_18__SCAN_IN), .ZN(P3_U3247) );
  AND2_X1 U11526 ( .A1(n9156), .A2(P3_D_REG_27__SCAN_IN), .ZN(P3_U3238) );
  AND2_X1 U11527 ( .A1(n9156), .A2(P3_D_REG_23__SCAN_IN), .ZN(P3_U3242) );
  AND2_X1 U11528 ( .A1(n9156), .A2(P3_D_REG_28__SCAN_IN), .ZN(P3_U3237) );
  AND2_X1 U11529 ( .A1(n9156), .A2(P3_D_REG_26__SCAN_IN), .ZN(P3_U3239) );
  AND2_X1 U11530 ( .A1(n9156), .A2(P3_D_REG_21__SCAN_IN), .ZN(P3_U3244) );
  AND2_X1 U11531 ( .A1(n9156), .A2(P3_D_REG_31__SCAN_IN), .ZN(P3_U3234) );
  AND2_X1 U11532 ( .A1(n9156), .A2(P3_D_REG_19__SCAN_IN), .ZN(P3_U3246) );
  AND2_X1 U11533 ( .A1(n9156), .A2(P3_D_REG_20__SCAN_IN), .ZN(P3_U3245) );
  AND2_X1 U11534 ( .A1(n9156), .A2(P3_D_REG_24__SCAN_IN), .ZN(P3_U3241) );
  AND2_X1 U11535 ( .A1(n9156), .A2(P3_D_REG_17__SCAN_IN), .ZN(P3_U3248) );
  AND2_X1 U11536 ( .A1(n9156), .A2(P3_D_REG_16__SCAN_IN), .ZN(P3_U3249) );
  AND2_X1 U11537 ( .A1(n9156), .A2(P3_D_REG_22__SCAN_IN), .ZN(P3_U3243) );
  AND2_X1 U11538 ( .A1(n9156), .A2(P3_D_REG_10__SCAN_IN), .ZN(P3_U3255) );
  AND2_X1 U11539 ( .A1(n9156), .A2(P3_D_REG_25__SCAN_IN), .ZN(P3_U3240) );
  AND2_X1 U11540 ( .A1(n9156), .A2(P3_D_REG_14__SCAN_IN), .ZN(P3_U3251) );
  AND2_X1 U11541 ( .A1(n9156), .A2(P3_D_REG_13__SCAN_IN), .ZN(P3_U3252) );
  AND2_X1 U11542 ( .A1(n9156), .A2(P3_D_REG_11__SCAN_IN), .ZN(P3_U3254) );
  AND2_X1 U11543 ( .A1(n9156), .A2(P3_D_REG_30__SCAN_IN), .ZN(P3_U3235) );
  AND2_X1 U11544 ( .A1(n9156), .A2(P3_D_REG_29__SCAN_IN), .ZN(P3_U3236) );
  AND2_X1 U11545 ( .A1(n9156), .A2(P3_D_REG_9__SCAN_IN), .ZN(P3_U3256) );
  AND2_X1 U11546 ( .A1(n9156), .A2(P3_D_REG_7__SCAN_IN), .ZN(P3_U3258) );
  AND2_X1 U11547 ( .A1(n9156), .A2(P3_D_REG_4__SCAN_IN), .ZN(P3_U3261) );
  AND2_X1 U11548 ( .A1(n9156), .A2(P3_D_REG_3__SCAN_IN), .ZN(P3_U3262) );
  AND2_X1 U11549 ( .A1(n9156), .A2(P3_D_REG_2__SCAN_IN), .ZN(P3_U3263) );
  INV_X1 U11550 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n9099) );
  MUX2_X1 U11551 ( .A(n9099), .B(P1_REG1_REG_8__SCAN_IN), .S(n9140), .Z(n9111)
         );
  INV_X1 U11552 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n14651) );
  MUX2_X1 U11553 ( .A(P1_REG1_REG_2__SCAN_IN), .B(n8371), .S(n13797), .Z(n9100) );
  MUX2_X1 U11554 ( .A(n8358), .B(P1_REG1_REG_1__SCAN_IN), .S(n13778), .Z(
        n13781) );
  AND2_X1 U11555 ( .A1(P1_REG1_REG_0__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), 
        .ZN(n13782) );
  NAND2_X1 U11556 ( .A1(n13781), .A2(n13782), .ZN(n13780) );
  OAI21_X1 U11557 ( .B1(n8358), .B2(n13778), .A(n13780), .ZN(n13787) );
  NAND2_X1 U11558 ( .A1(n13797), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n13810) );
  NAND2_X1 U11559 ( .A1(n13811), .A2(n13810), .ZN(n9102) );
  MUX2_X1 U11560 ( .A(P1_REG1_REG_3__SCAN_IN), .B(n8385), .S(n13808), .Z(n9101) );
  NAND2_X1 U11561 ( .A1(n9102), .A2(n9101), .ZN(n13813) );
  NAND2_X1 U11562 ( .A1(n13808), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n9234) );
  NAND2_X1 U11563 ( .A1(n13813), .A2(n9234), .ZN(n9105) );
  INV_X1 U11564 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n9103) );
  MUX2_X1 U11565 ( .A(P1_REG1_REG_4__SCAN_IN), .B(n9103), .S(n9232), .Z(n9104)
         );
  NAND2_X1 U11566 ( .A1(n9105), .A2(n9104), .ZN(n9236) );
  NAND2_X1 U11567 ( .A1(n9232), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n9106) );
  NAND2_X1 U11568 ( .A1(n9236), .A2(n9106), .ZN(n9160) );
  MUX2_X1 U11569 ( .A(n9107), .B(P1_REG1_REG_5__SCAN_IN), .S(n9164), .Z(n9161)
         );
  OR2_X1 U11570 ( .A1(n9164), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n9108) );
  NAND2_X1 U11571 ( .A1(n9158), .A2(n9108), .ZN(n9176) );
  INV_X1 U11572 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n9871) );
  MUX2_X1 U11573 ( .A(n9871), .B(P1_REG1_REG_6__SCAN_IN), .S(n9121), .Z(n9175)
         );
  NOR2_X1 U11574 ( .A1(n9176), .A2(n9175), .ZN(n9217) );
  NOR2_X1 U11575 ( .A1(n9183), .A2(n9871), .ZN(n9212) );
  MUX2_X1 U11576 ( .A(P1_REG1_REG_7__SCAN_IN), .B(n14651), .S(n9211), .Z(n9109) );
  OAI21_X1 U11577 ( .B1(n14651), .B2(n9209), .A(n9215), .ZN(n9110) );
  AOI21_X1 U11578 ( .B1(n9111), .B2(n9110), .A(n9143), .ZN(n9135) );
  NAND2_X1 U11579 ( .A1(n9113), .A2(n9112), .ZN(n14452) );
  NOR2_X2 U11580 ( .A1(n14452), .A2(n14442), .ZN(n14483) );
  INV_X1 U11581 ( .A(n14483), .ZN(n14459) );
  INV_X1 U11582 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n15232) );
  MUX2_X1 U11583 ( .A(P1_REG2_REG_2__SCAN_IN), .B(n15232), .S(n13797), .Z(
        n9115) );
  INV_X1 U11584 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n9114) );
  MUX2_X1 U11585 ( .A(n9114), .B(P1_REG2_REG_1__SCAN_IN), .S(n13778), .Z(
        n13776) );
  NAND3_X1 U11586 ( .A1(n13776), .A2(P1_IR_REG_0__SCAN_IN), .A3(
        P1_REG2_REG_0__SCAN_IN), .ZN(n13775) );
  OAI21_X1 U11587 ( .B1(n9114), .B2(n13778), .A(n13775), .ZN(n13791) );
  NAND2_X1 U11588 ( .A1(n9115), .A2(n13791), .ZN(n13805) );
  NAND2_X1 U11589 ( .A1(n13797), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n13804) );
  INV_X1 U11590 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n9116) );
  MUX2_X1 U11591 ( .A(n9116), .B(P1_REG2_REG_3__SCAN_IN), .S(n13808), .Z(
        n13803) );
  AOI21_X1 U11592 ( .B1(n13805), .B2(n13804), .A(n13803), .ZN(n13802) );
  NOR2_X1 U11593 ( .A1(n9117), .A2(n9116), .ZN(n9227) );
  INV_X1 U11594 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n9768) );
  MUX2_X1 U11595 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n9768), .S(n9232), .Z(n9118)
         );
  OAI21_X1 U11596 ( .B1(n13802), .B2(n9227), .A(n9118), .ZN(n9230) );
  NAND2_X1 U11597 ( .A1(n9232), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n9166) );
  MUX2_X1 U11598 ( .A(n9119), .B(P1_REG2_REG_5__SCAN_IN), .S(n9164), .Z(n9165)
         );
  AOI21_X1 U11599 ( .B1(n9230), .B2(n9166), .A(n9165), .ZN(n9179) );
  NOR2_X1 U11600 ( .A1(n9120), .A2(n9119), .ZN(n9178) );
  INV_X1 U11601 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n9918) );
  MUX2_X1 U11602 ( .A(P1_REG2_REG_6__SCAN_IN), .B(n9918), .S(n9121), .Z(n9177)
         );
  OAI21_X1 U11603 ( .B1(n9179), .B2(n9178), .A(n9177), .ZN(n9206) );
  NAND2_X1 U11604 ( .A1(n9121), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n9205) );
  INV_X1 U11605 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n9122) );
  MUX2_X1 U11606 ( .A(n9122), .B(P1_REG2_REG_7__SCAN_IN), .S(n9211), .Z(n9204)
         );
  AOI21_X1 U11607 ( .B1(n9206), .B2(n9205), .A(n9204), .ZN(n9221) );
  NOR2_X1 U11608 ( .A1(n9209), .A2(n9122), .ZN(n9127) );
  INV_X1 U11609 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n10364) );
  MUX2_X1 U11610 ( .A(P1_REG2_REG_8__SCAN_IN), .B(n10364), .S(n9140), .Z(n9126) );
  NOR3_X1 U11611 ( .A1(n9221), .A2(n9127), .A3(n9126), .ZN(n9125) );
  INV_X1 U11612 ( .A(n14452), .ZN(n9124) );
  NOR2_X1 U11613 ( .A1(n11640), .A2(n14264), .ZN(n9123) );
  NAND2_X1 U11614 ( .A1(n9124), .A2(n9123), .ZN(n14464) );
  NOR2_X1 U11615 ( .A1(n9125), .A2(n14464), .ZN(n9133) );
  OAI21_X1 U11616 ( .B1(n9221), .B2(n9127), .A(n9126), .ZN(n9138) );
  INV_X1 U11617 ( .A(n14472), .ZN(n14469) );
  NOR2_X2 U11618 ( .A1(n14452), .A2(n9128), .ZN(n14476) );
  NAND2_X1 U11619 ( .A1(n14476), .A2(n9140), .ZN(n9130) );
  NAND2_X1 U11620 ( .A1(P1_REG3_REG_8__SCAN_IN), .A2(P1_U3086), .ZN(n9129) );
  OAI211_X1 U11621 ( .C1(n9131), .C2(n14469), .A(n9130), .B(n9129), .ZN(n9132)
         );
  AOI21_X1 U11622 ( .B1(n9133), .B2(n9138), .A(n9132), .ZN(n9134) );
  OAI21_X1 U11623 ( .B1(n9135), .B2(n14459), .A(n9134), .ZN(P1_U3251) );
  NAND2_X1 U11624 ( .A1(n9140), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n9137) );
  INV_X1 U11625 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n9259) );
  MUX2_X1 U11626 ( .A(P1_REG2_REG_9__SCAN_IN), .B(n9259), .S(n9260), .Z(n9136)
         );
  AOI21_X1 U11627 ( .B1(n9138), .B2(n9137), .A(n9136), .ZN(n9263) );
  NAND3_X1 U11628 ( .A1(n9138), .A2(n9137), .A3(n9136), .ZN(n9139) );
  NAND2_X1 U11629 ( .A1(n9139), .A2(n14478), .ZN(n9149) );
  NOR2_X1 U11630 ( .A1(n9140), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n9141) );
  INV_X1 U11631 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n14653) );
  MUX2_X1 U11632 ( .A(n14653), .B(P1_REG1_REG_9__SCAN_IN), .S(n9260), .Z(n9142) );
  OAI21_X1 U11633 ( .B1(n9143), .B2(n9141), .A(n9142), .ZN(n9255) );
  INV_X1 U11634 ( .A(n9255), .ZN(n9145) );
  NOR3_X1 U11635 ( .A1(n9143), .A2(n9142), .A3(n9141), .ZN(n9144) );
  OAI21_X1 U11636 ( .B1(n9145), .B2(n9144), .A(n14483), .ZN(n9148) );
  NAND2_X1 U11637 ( .A1(P1_U3086), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n10683) );
  OAI21_X1 U11638 ( .B1(n14469), .B2(n8221), .A(n10683), .ZN(n9146) );
  AOI21_X1 U11639 ( .B1(n9256), .B2(n14476), .A(n9146), .ZN(n9147) );
  OAI211_X1 U11640 ( .C1(n9263), .C2(n9149), .A(n9148), .B(n9147), .ZN(
        P1_U3252) );
  OR2_X1 U11641 ( .A1(n9082), .A2(n9718), .ZN(n9151) );
  XNOR2_X1 U11642 ( .A(n9151), .B(n9150), .ZN(n12376) );
  NAND2_X1 U11643 ( .A1(n9154), .A2(n15367), .ZN(n9155) );
  NAND2_X1 U11644 ( .A1(n9200), .A2(n9155), .ZN(n11162) );
  OAI222_X1 U11645 ( .A1(P3_U3151), .A2(n12376), .B1(n11338), .B2(n11163), 
        .C1(n12245), .C2(n11162), .ZN(P3_U3282) );
  INV_X1 U11646 ( .A(n9156), .ZN(n9157) );
  INV_X1 U11647 ( .A(P3_D_REG_15__SCAN_IN), .ZN(n15329) );
  NOR2_X1 U11648 ( .A1(n9157), .A2(n15329), .ZN(P3_U3250) );
  INV_X1 U11649 ( .A(P3_D_REG_8__SCAN_IN), .ZN(n15216) );
  NOR2_X1 U11650 ( .A1(n9157), .A2(n15216), .ZN(P3_U3257) );
  INV_X1 U11651 ( .A(P3_D_REG_6__SCAN_IN), .ZN(n15229) );
  NOR2_X1 U11652 ( .A1(n9157), .A2(n15229), .ZN(P3_U3259) );
  INV_X1 U11653 ( .A(P3_D_REG_5__SCAN_IN), .ZN(n15187) );
  NOR2_X1 U11654 ( .A1(n9157), .A2(n15187), .ZN(P3_U3260) );
  INV_X1 U11655 ( .A(P3_D_REG_12__SCAN_IN), .ZN(n15338) );
  NOR2_X1 U11656 ( .A1(n9157), .A2(n15338), .ZN(P3_U3253) );
  INV_X1 U11657 ( .A(n9158), .ZN(n9159) );
  AOI21_X1 U11658 ( .B1(n9161), .B2(n9160), .A(n9159), .ZN(n9171) );
  NOR2_X1 U11659 ( .A1(n9162), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9847) );
  NOR2_X1 U11660 ( .A1(n14469), .A2(n15281), .ZN(n9163) );
  AOI211_X1 U11661 ( .C1(n14476), .C2(n9164), .A(n9847), .B(n9163), .ZN(n9170)
         );
  INV_X1 U11662 ( .A(n9179), .ZN(n9168) );
  NAND3_X1 U11663 ( .A1(n9230), .A2(n9166), .A3(n9165), .ZN(n9167) );
  NAND3_X1 U11664 ( .A1(n14478), .A2(n9168), .A3(n9167), .ZN(n9169) );
  OAI211_X1 U11665 ( .C1(n9171), .C2(n14459), .A(n9170), .B(n9169), .ZN(
        P1_U3248) );
  OAI222_X1 U11666 ( .A1(P1_U3086), .A2(n9260), .B1(n6535), .B2(n9174), .C1(
        n9172), .C2(n14266), .ZN(P1_U3346) );
  INV_X1 U11667 ( .A(n9341), .ZN(n14699) );
  OAI222_X1 U11668 ( .A1(P2_U3088), .A2(n14699), .B1(n6534), .B2(n9174), .C1(
        n9173), .C2(n11904), .ZN(P2_U3318) );
  AOI211_X1 U11669 ( .C1(n9176), .C2(n9175), .A(n9217), .B(n14459), .ZN(n9186)
         );
  INV_X1 U11670 ( .A(n9206), .ZN(n9181) );
  NOR3_X1 U11671 ( .A1(n9179), .A2(n9178), .A3(n9177), .ZN(n9180) );
  NOR3_X1 U11672 ( .A1(n14464), .A2(n9181), .A3(n9180), .ZN(n9185) );
  INV_X1 U11673 ( .A(n14476), .ZN(n13832) );
  NAND2_X1 U11674 ( .A1(P1_U3086), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n9951) );
  NAND2_X1 U11675 ( .A1(n14472), .A2(P1_ADDR_REG_6__SCAN_IN), .ZN(n9182) );
  OAI211_X1 U11676 ( .C1(n13832), .C2(n9183), .A(n9951), .B(n9182), .ZN(n9184)
         );
  OR3_X1 U11677 ( .A1(n9186), .A2(n9185), .A3(n9184), .ZN(P1_U3249) );
  NAND2_X1 U11678 ( .A1(n14397), .A2(n14108), .ZN(n13748) );
  INV_X1 U11679 ( .A(n13748), .ZN(n13718) );
  NAND2_X1 U11680 ( .A1(n9188), .A2(n9187), .ZN(n9406) );
  AOI22_X1 U11681 ( .A1(n13718), .A2(n14556), .B1(P1_REG3_REG_0__SCAN_IN), 
        .B2(n9406), .ZN(n9193) );
  OAI21_X1 U11682 ( .B1(n9191), .B2(n9190), .A(n9189), .ZN(n9224) );
  NAND2_X1 U11683 ( .A1(n9224), .A2(n14395), .ZN(n9192) );
  OAI211_X1 U11684 ( .C1(n13743), .C2(n9669), .A(n9193), .B(n9192), .ZN(
        P1_U3232) );
  NOR2_X1 U11685 ( .A1(n9194), .A2(n9718), .ZN(n9195) );
  MUX2_X1 U11686 ( .A(n9718), .B(n9195), .S(P3_IR_REG_14__SCAN_IN), .Z(n9198)
         );
  INV_X1 U11687 ( .A(n9196), .ZN(n9197) );
  INV_X1 U11688 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n9595) );
  NAND2_X1 U11689 ( .A1(n9595), .A2(P1_DATAO_REG_14__SCAN_IN), .ZN(n9290) );
  INV_X1 U11690 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n9594) );
  NAND2_X1 U11691 ( .A1(n9594), .A2(P2_DATAO_REG_14__SCAN_IN), .ZN(n9201) );
  OAI21_X1 U11692 ( .B1(n9203), .B2(n9202), .A(n9291), .ZN(n11260) );
  OAI222_X1 U11693 ( .A1(P3_U3151), .A2(n12400), .B1(n11338), .B2(n11261), 
        .C1(n12245), .C2(n11260), .ZN(P3_U3281) );
  NAND3_X1 U11694 ( .A1(n9206), .A2(n9205), .A3(n9204), .ZN(n9207) );
  NAND2_X1 U11695 ( .A1(n14478), .A2(n9207), .ZN(n9220) );
  NOR2_X1 U11696 ( .A1(n9208), .A2(P1_STATE_REG_SCAN_IN), .ZN(n10295) );
  NOR2_X1 U11697 ( .A1(n13832), .A2(n9209), .ZN(n9210) );
  AOI211_X1 U11698 ( .C1(n14472), .C2(P1_ADDR_REG_7__SCAN_IN), .A(n10295), .B(
        n9210), .ZN(n9219) );
  MUX2_X1 U11699 ( .A(n14651), .B(P1_REG1_REG_7__SCAN_IN), .S(n9211), .Z(n9214) );
  INV_X1 U11700 ( .A(n9212), .ZN(n9213) );
  NAND2_X1 U11701 ( .A1(n9214), .A2(n9213), .ZN(n9216) );
  OAI211_X1 U11702 ( .C1(n9217), .C2(n9216), .A(n9215), .B(n14483), .ZN(n9218)
         );
  OAI211_X1 U11703 ( .C1(n9221), .C2(n9220), .A(n9219), .B(n9218), .ZN(
        P1_U3250) );
  INV_X1 U11704 ( .A(n9222), .ZN(n9270) );
  AOI22_X1 U11705 ( .A1(n9477), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n14260), .ZN(n9223) );
  OAI21_X1 U11706 ( .B1(n9270), .B2(n6535), .A(n9223), .ZN(P1_U3345) );
  NAND2_X1 U11707 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n13774) );
  MUX2_X1 U11708 ( .A(n13774), .B(n9224), .S(n14264), .Z(n9226) );
  NOR2_X1 U11709 ( .A1(n14264), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n9225) );
  OR2_X1 U11710 ( .A1(n11640), .A2(n9225), .ZN(n14443) );
  NAND2_X1 U11711 ( .A1(n14443), .A2(n14445), .ZN(n14448) );
  OAI211_X1 U11712 ( .C1(n9226), .C2(n11640), .A(P1_U4016), .B(n14448), .ZN(
        n13801) );
  INV_X1 U11713 ( .A(n9227), .ZN(n9229) );
  MUX2_X1 U11714 ( .A(n9768), .B(P1_REG2_REG_4__SCAN_IN), .S(n9232), .Z(n9228)
         );
  NAND2_X1 U11715 ( .A1(n9229), .A2(n9228), .ZN(n9231) );
  OAI211_X1 U11716 ( .C1(n13802), .C2(n9231), .A(n14478), .B(n9230), .ZN(n9240) );
  AND2_X1 U11717 ( .A1(P1_U3086), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n9928) );
  AOI21_X1 U11718 ( .B1(n14472), .B2(P1_ADDR_REG_4__SCAN_IN), .A(n9928), .ZN(
        n9239) );
  NAND2_X1 U11719 ( .A1(n14476), .A2(n9232), .ZN(n9238) );
  MUX2_X1 U11720 ( .A(n9103), .B(P1_REG1_REG_4__SCAN_IN), .S(n9232), .Z(n9233)
         );
  NAND3_X1 U11721 ( .A1(n13813), .A2(n9234), .A3(n9233), .ZN(n9235) );
  NAND3_X1 U11722 ( .A1(n14483), .A2(n9236), .A3(n9235), .ZN(n9237) );
  AND4_X1 U11723 ( .A1(n9240), .A2(n9239), .A3(n9238), .A4(n9237), .ZN(n9241)
         );
  NAND2_X1 U11724 ( .A1(n13801), .A2(n9241), .ZN(P1_U3247) );
  NOR3_X1 U11725 ( .A1(n9669), .A2(n14271), .A3(n9242), .ZN(n9250) );
  NAND2_X1 U11726 ( .A1(n9246), .A2(n9245), .ZN(n9247) );
  NAND2_X1 U11727 ( .A1(n9658), .A2(n13847), .ZN(n14493) );
  OR2_X1 U11728 ( .A1(n9248), .A2(n13847), .ZN(n14592) );
  NAND2_X1 U11729 ( .A1(n14493), .A2(n14592), .ZN(n14641) );
  AOI21_X1 U11730 ( .B1(n14560), .B2(n14611), .A(n9895), .ZN(n9249) );
  AOI211_X1 U11731 ( .C1(n14108), .C2(n14556), .A(n9250), .B(n9249), .ZN(n9360) );
  NAND2_X1 U11732 ( .A1(n9656), .A2(n9251), .ZN(n9252) );
  NOR2_X1 U11733 ( .A1(n9252), .A2(n9655), .ZN(n9359) );
  INV_X1 U11734 ( .A(n14658), .ZN(n14655) );
  NAND2_X1 U11735 ( .A1(n14655), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n9254) );
  OAI21_X1 U11736 ( .B1(n9360), .B2(n14655), .A(n9254), .ZN(P1_U3528) );
  OAI21_X1 U11737 ( .B1(n9256), .B2(P1_REG1_REG_9__SCAN_IN), .A(n9255), .ZN(
        n9258) );
  INV_X1 U11738 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n14656) );
  MUX2_X1 U11739 ( .A(n14656), .B(P1_REG1_REG_10__SCAN_IN), .S(n9477), .Z(
        n9257) );
  NOR2_X1 U11740 ( .A1(n9258), .A2(n9257), .ZN(n9476) );
  AOI211_X1 U11741 ( .C1(n9258), .C2(n9257), .A(n14459), .B(n9476), .ZN(n9269)
         );
  INV_X1 U11742 ( .A(n9477), .ZN(n9475) );
  NOR2_X1 U11743 ( .A1(n9260), .A2(n9259), .ZN(n9262) );
  INV_X1 U11744 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n10508) );
  MUX2_X1 U11745 ( .A(P1_REG2_REG_10__SCAN_IN), .B(n10508), .S(n9477), .Z(
        n9261) );
  OAI21_X1 U11746 ( .B1(n9263), .B2(n9262), .A(n9261), .ZN(n9474) );
  OR3_X1 U11747 ( .A1(n9263), .A2(n9262), .A3(n9261), .ZN(n9264) );
  NAND3_X1 U11748 ( .A1(n9474), .A2(n14478), .A3(n9264), .ZN(n9267) );
  INV_X1 U11749 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n9265) );
  NOR2_X1 U11750 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n9265), .ZN(n10834) );
  AOI21_X1 U11751 ( .B1(n14472), .B2(P1_ADDR_REG_10__SCAN_IN), .A(n10834), 
        .ZN(n9266) );
  OAI211_X1 U11752 ( .C1(n13832), .C2(n9475), .A(n9267), .B(n9266), .ZN(n9268)
         );
  OR2_X1 U11753 ( .A1(n9269), .A2(n9268), .ZN(P1_U3253) );
  INV_X1 U11754 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n9271) );
  INV_X1 U11755 ( .A(n9343), .ZN(n14704) );
  OAI222_X1 U11756 ( .A1(n11904), .A2(n9271), .B1(n6534), .B2(n9270), .C1(
        P2_U3088), .C2(n14704), .ZN(P2_U3317) );
  INV_X1 U11757 ( .A(n9272), .ZN(n9276) );
  INV_X1 U11758 ( .A(n11011), .ZN(n9274) );
  OAI21_X1 U11759 ( .B1(n9274), .B2(n9421), .A(n9273), .ZN(n9275) );
  AND2_X1 U11760 ( .A1(n9276), .A2(n9275), .ZN(n9286) );
  INV_X1 U11761 ( .A(n9286), .ZN(n9281) );
  NOR2_X1 U11762 ( .A1(n8155), .A2(P2_U3088), .ZN(n13479) );
  AND2_X1 U11763 ( .A1(n9281), .A2(n13479), .ZN(n9278) );
  INV_X1 U11764 ( .A(n9278), .ZN(n9277) );
  OR2_X1 U11765 ( .A1(n9277), .A2(n13484), .ZN(n14745) );
  AOI22_X1 U11766 ( .A1(P2_REG2_REG_0__SCAN_IN), .A2(n14756), .B1(n14759), 
        .B2(P2_REG1_REG_0__SCAN_IN), .ZN(n9285) );
  NAND2_X1 U11767 ( .A1(n14759), .A2(n9279), .ZN(n9282) );
  AND2_X1 U11768 ( .A1(n8155), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9280) );
  NAND2_X1 U11769 ( .A1(n9281), .A2(n9280), .ZN(n14739) );
  OAI211_X1 U11770 ( .C1(P2_REG2_REG_0__SCAN_IN), .C2(n14745), .A(n9282), .B(
        n14739), .ZN(n9283) );
  INV_X1 U11771 ( .A(n9283), .ZN(n9284) );
  MUX2_X1 U11772 ( .A(n9285), .B(n9284), .S(n15206), .Z(n9288) );
  AND2_X1 U11773 ( .A1(n9286), .A2(P2_STATE_REG_SCAN_IN), .ZN(n14752) );
  AOI22_X1 U11774 ( .A1(n14752), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3088), .ZN(n9287) );
  NAND2_X1 U11775 ( .A1(n9288), .A2(n9287), .ZN(P2_U3214) );
  NAND2_X1 U11776 ( .A1(n9196), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9289) );
  XNOR2_X1 U11777 ( .A(n9289), .B(n6946), .ZN(n12422) );
  NAND2_X1 U11778 ( .A1(n9785), .A2(P1_DATAO_REG_15__SCAN_IN), .ZN(n9493) );
  NAND2_X1 U11779 ( .A1(n15325), .A2(P2_DATAO_REG_15__SCAN_IN), .ZN(n9292) );
  AND2_X1 U11780 ( .A1(n9493), .A2(n9292), .ZN(n9293) );
  OAI21_X1 U11781 ( .B1(n9294), .B2(n9293), .A(n9494), .ZN(n11314) );
  OAI222_X1 U11782 ( .A1(P3_U3151), .A2(n12422), .B1(n11338), .B2(n11315), 
        .C1(n12245), .C2(n11314), .ZN(P3_U3280) );
  XOR2_X1 U11783 ( .A(n9296), .B(n9295), .Z(n9299) );
  NOR2_X1 U11784 ( .A1(n13738), .A2(n14561), .ZN(n13750) );
  AOI22_X1 U11785 ( .A1(n13750), .A2(n8344), .B1(n13718), .B2(n13772), .ZN(
        n9298) );
  AOI22_X1 U11786 ( .A1(n14398), .A2(n6539), .B1(n9406), .B2(
        P1_REG3_REG_1__SCAN_IN), .ZN(n9297) );
  OAI211_X1 U11787 ( .C1(n9299), .C2(n13756), .A(n9298), .B(n9297), .ZN(
        P1_U3222) );
  INV_X1 U11788 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n9300) );
  MUX2_X1 U11789 ( .A(P2_REG2_REG_2__SCAN_IN), .B(n9300), .S(n13068), .Z(
        n13065) );
  INV_X1 U11790 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n15230) );
  MUX2_X1 U11791 ( .A(n15230), .B(P2_REG2_REG_1__SCAN_IN), .S(n13058), .Z(
        n13053) );
  AND2_X1 U11792 ( .A1(P2_REG2_REG_0__SCAN_IN), .A2(n15206), .ZN(n13054) );
  NAND2_X1 U11793 ( .A1(n13053), .A2(n13054), .ZN(n13052) );
  OAI21_X1 U11794 ( .B1(n15230), .B2(n13058), .A(n13052), .ZN(n13064) );
  NAND2_X1 U11795 ( .A1(n13065), .A2(n13064), .ZN(n13078) );
  NAND2_X1 U11796 ( .A1(n13068), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n13077) );
  NAND2_X1 U11797 ( .A1(n13078), .A2(n13077), .ZN(n9303) );
  MUX2_X1 U11798 ( .A(P2_REG2_REG_3__SCAN_IN), .B(n9301), .S(n13081), .Z(n9302) );
  NAND2_X1 U11799 ( .A1(n9303), .A2(n9302), .ZN(n13080) );
  NAND2_X1 U11800 ( .A1(n13081), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n9304) );
  NAND2_X1 U11801 ( .A1(n13080), .A2(n9304), .ZN(n14670) );
  MUX2_X1 U11802 ( .A(n10128), .B(P2_REG2_REG_4__SCAN_IN), .S(n14660), .Z(
        n14669) );
  NAND2_X1 U11803 ( .A1(n14670), .A2(n14669), .ZN(n14676) );
  NAND2_X1 U11804 ( .A1(n14668), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n14675) );
  NAND2_X1 U11805 ( .A1(n14676), .A2(n14675), .ZN(n9306) );
  INV_X1 U11806 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n10171) );
  MUX2_X1 U11807 ( .A(P2_REG2_REG_5__SCAN_IN), .B(n10171), .S(n14681), .Z(
        n9305) );
  NAND2_X1 U11808 ( .A1(n9306), .A2(n9305), .ZN(n14678) );
  NAND2_X1 U11809 ( .A1(n14681), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n9307) );
  NAND2_X1 U11810 ( .A1(n14678), .A2(n9307), .ZN(n9367) );
  INV_X1 U11811 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n10145) );
  MUX2_X1 U11812 ( .A(P2_REG2_REG_6__SCAN_IN), .B(n10145), .S(n9370), .Z(n9366) );
  NAND2_X1 U11813 ( .A1(n9367), .A2(n9366), .ZN(n13094) );
  NAND2_X1 U11814 ( .A1(n9370), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n13093) );
  NAND2_X1 U11815 ( .A1(n13094), .A2(n13093), .ZN(n9309) );
  MUX2_X1 U11816 ( .A(P2_REG2_REG_7__SCAN_IN), .B(n10182), .S(n13096), .Z(
        n9308) );
  NAND2_X1 U11817 ( .A1(n9309), .A2(n9308), .ZN(n13108) );
  NAND2_X1 U11818 ( .A1(n13096), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n13107) );
  NAND2_X1 U11819 ( .A1(n13108), .A2(n13107), .ZN(n9311) );
  MUX2_X1 U11820 ( .A(P2_REG2_REG_8__SCAN_IN), .B(n10474), .S(n13111), .Z(
        n9310) );
  NAND2_X1 U11821 ( .A1(n9311), .A2(n9310), .ZN(n13110) );
  NAND2_X1 U11822 ( .A1(n13111), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n9312) );
  NAND2_X1 U11823 ( .A1(n13110), .A2(n9312), .ZN(n14688) );
  INV_X1 U11824 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n9313) );
  MUX2_X1 U11825 ( .A(n9313), .B(P2_REG2_REG_9__SCAN_IN), .S(n9341), .Z(n14687) );
  OR2_X1 U11826 ( .A1(n9341), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n9314) );
  NAND2_X1 U11827 ( .A1(n14690), .A2(n9314), .ZN(n14708) );
  MUX2_X1 U11828 ( .A(n10425), .B(P2_REG2_REG_10__SCAN_IN), .S(n9343), .Z(
        n14707) );
  NAND2_X1 U11829 ( .A1(n9343), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n9315) );
  NAND2_X1 U11830 ( .A1(n14709), .A2(n9315), .ZN(n9318) );
  INV_X1 U11831 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n10649) );
  MUX2_X1 U11832 ( .A(n10649), .B(P2_REG2_REG_11__SCAN_IN), .S(n10157), .Z(
        n9317) );
  INV_X1 U11833 ( .A(n14726), .ZN(n9316) );
  AOI21_X1 U11834 ( .B1(n9318), .B2(n9317), .A(n9316), .ZN(n9352) );
  INV_X1 U11835 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n10626) );
  NOR2_X1 U11836 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10626), .ZN(n9320) );
  INV_X1 U11837 ( .A(n10157), .ZN(n9400) );
  NOR2_X1 U11838 ( .A1(n14739), .A2(n9400), .ZN(n9319) );
  AOI211_X1 U11839 ( .C1(P2_ADDR_REG_11__SCAN_IN), .C2(n14752), .A(n9320), .B(
        n9319), .ZN(n9351) );
  MUX2_X1 U11840 ( .A(P2_REG1_REG_2__SCAN_IN), .B(n9321), .S(n13068), .Z(
        n13067) );
  MUX2_X1 U11841 ( .A(n9322), .B(P2_REG1_REG_1__SCAN_IN), .S(n13058), .Z(
        n13056) );
  AND2_X1 U11842 ( .A1(P2_REG1_REG_0__SCAN_IN), .A2(n15206), .ZN(n13057) );
  NAND2_X1 U11843 ( .A1(n13056), .A2(n13057), .ZN(n13055) );
  OAI21_X1 U11844 ( .B1(n9322), .B2(n13058), .A(n13055), .ZN(n13066) );
  NAND2_X1 U11845 ( .A1(n13067), .A2(n13066), .ZN(n13084) );
  NAND2_X1 U11846 ( .A1(n13068), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n13083) );
  NAND2_X1 U11847 ( .A1(n13084), .A2(n13083), .ZN(n9324) );
  MUX2_X1 U11848 ( .A(P2_REG1_REG_3__SCAN_IN), .B(n7623), .S(n13081), .Z(n9323) );
  NAND2_X1 U11849 ( .A1(n9324), .A2(n9323), .ZN(n14663) );
  NAND2_X1 U11850 ( .A1(n13081), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n14662) );
  NAND2_X1 U11851 ( .A1(n14663), .A2(n14662), .ZN(n9327) );
  INV_X1 U11852 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n9325) );
  MUX2_X1 U11853 ( .A(n9325), .B(P2_REG1_REG_4__SCAN_IN), .S(n14660), .Z(n9326) );
  NAND2_X1 U11854 ( .A1(n9327), .A2(n9326), .ZN(n14665) );
  NAND2_X1 U11855 ( .A1(n14668), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n9328) );
  NAND2_X1 U11856 ( .A1(n14665), .A2(n9328), .ZN(n14684) );
  MUX2_X1 U11857 ( .A(P2_REG1_REG_5__SCAN_IN), .B(n9329), .S(n14681), .Z(
        n14683) );
  NAND2_X1 U11858 ( .A1(n14684), .A2(n14683), .ZN(n14682) );
  NAND2_X1 U11859 ( .A1(n14681), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n9364) );
  NAND2_X1 U11860 ( .A1(n14682), .A2(n9364), .ZN(n9332) );
  INV_X1 U11861 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n9330) );
  MUX2_X1 U11862 ( .A(P2_REG1_REG_6__SCAN_IN), .B(n9330), .S(n9370), .Z(n9331)
         );
  NAND2_X1 U11863 ( .A1(n9332), .A2(n9331), .ZN(n13099) );
  NAND2_X1 U11864 ( .A1(n9370), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n13098) );
  NAND2_X1 U11865 ( .A1(n13099), .A2(n13098), .ZN(n9335) );
  INV_X1 U11866 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n9333) );
  MUX2_X1 U11867 ( .A(P2_REG1_REG_7__SCAN_IN), .B(n9333), .S(n13096), .Z(n9334) );
  NAND2_X1 U11868 ( .A1(n9335), .A2(n9334), .ZN(n13114) );
  NAND2_X1 U11869 ( .A1(n13096), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n13113) );
  NAND2_X1 U11870 ( .A1(n13114), .A2(n13113), .ZN(n9338) );
  INV_X1 U11871 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n9336) );
  MUX2_X1 U11872 ( .A(P2_REG1_REG_8__SCAN_IN), .B(n9336), .S(n13111), .Z(n9337) );
  NAND2_X1 U11873 ( .A1(n9338), .A2(n9337), .ZN(n13116) );
  NAND2_X1 U11874 ( .A1(n13111), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n9339) );
  NAND2_X1 U11875 ( .A1(n13116), .A2(n9339), .ZN(n14693) );
  INV_X1 U11876 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n9340) );
  MUX2_X1 U11877 ( .A(n9340), .B(P2_REG1_REG_9__SCAN_IN), .S(n9341), .Z(n14692) );
  OR2_X1 U11878 ( .A1(n9341), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n9342) );
  NAND2_X1 U11879 ( .A1(n14695), .A2(n9342), .ZN(n14712) );
  MUX2_X1 U11880 ( .A(n7756), .B(P2_REG1_REG_10__SCAN_IN), .S(n9343), .Z(
        n14713) );
  NAND2_X1 U11881 ( .A1(n9343), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n9348) );
  NAND2_X1 U11882 ( .A1(n14714), .A2(n9348), .ZN(n9346) );
  MUX2_X1 U11883 ( .A(P2_REG1_REG_11__SCAN_IN), .B(n9344), .S(n10157), .Z(
        n9345) );
  NAND2_X1 U11884 ( .A1(n9346), .A2(n9345), .ZN(n10152) );
  MUX2_X1 U11885 ( .A(n9344), .B(P2_REG1_REG_11__SCAN_IN), .S(n10157), .Z(
        n9347) );
  NAND3_X1 U11886 ( .A1(n14714), .A2(n9348), .A3(n9347), .ZN(n9349) );
  NAND3_X1 U11887 ( .A1(n10152), .A2(n14759), .A3(n9349), .ZN(n9350) );
  OAI211_X1 U11888 ( .C1(n9352), .C2(n14745), .A(n9351), .B(n9350), .ZN(
        P2_U3225) );
  OAI21_X1 U11889 ( .B1(n9356), .B2(P1_D_REG_0__SCAN_IN), .A(n9353), .ZN(n9358) );
  INV_X1 U11890 ( .A(n9354), .ZN(n9355) );
  OR2_X1 U11891 ( .A1(n9356), .A2(n9355), .ZN(n9357) );
  INV_X1 U11892 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n9362) );
  OR2_X1 U11893 ( .A1(n9360), .A2(n14643), .ZN(n9361) );
  OAI21_X1 U11894 ( .B1(n14645), .B2(n9362), .A(n9361), .ZN(P1_U3459) );
  MUX2_X1 U11895 ( .A(n9330), .B(P2_REG1_REG_6__SCAN_IN), .S(n9370), .Z(n9363)
         );
  NAND3_X1 U11896 ( .A1(n14682), .A2(n9364), .A3(n9363), .ZN(n9365) );
  NAND3_X1 U11897 ( .A1(n14759), .A2(n13099), .A3(n9365), .ZN(n9372) );
  NAND2_X1 U11898 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_U3088), .ZN(n9608) );
  OAI211_X1 U11899 ( .C1(n9367), .C2(n9366), .A(n14756), .B(n13094), .ZN(n9368) );
  NAND2_X1 U11900 ( .A1(n9608), .A2(n9368), .ZN(n9369) );
  AOI21_X1 U11901 ( .B1(n14754), .B2(n9370), .A(n9369), .ZN(n9371) );
  OAI211_X1 U11902 ( .C1(n14736), .C2(n8264), .A(n9372), .B(n9371), .ZN(
        P2_U3220) );
  INV_X1 U11903 ( .A(P3_DATAO_REG_19__SCAN_IN), .ZN(n15277) );
  INV_X1 U11904 ( .A(P3_IR_REG_29__SCAN_IN), .ZN(n9378) );
  INV_X1 U11905 ( .A(P3_IR_REG_30__SCAN_IN), .ZN(n12877) );
  XNOR2_X2 U11906 ( .A(n9379), .B(n12877), .ZN(n11649) );
  AND2_X2 U11907 ( .A1(n11649), .A2(n9386), .ZN(n11521) );
  INV_X1 U11908 ( .A(P3_REG1_REG_19__SCAN_IN), .ZN(n12488) );
  INV_X1 U11909 ( .A(P3_REG2_REG_19__SCAN_IN), .ZN(n12631) );
  NAND2_X1 U11910 ( .A1(n11649), .A2(n11339), .ZN(n9738) );
  INV_X1 U11911 ( .A(P3_REG0_REG_19__SCAN_IN), .ZN(n9382) );
  OR2_X1 U11912 ( .A1(n11438), .A2(n9382), .ZN(n9383) );
  AND2_X1 U11913 ( .A1(n9384), .A2(n9383), .ZN(n9389) );
  INV_X1 U11914 ( .A(P3_REG3_REG_5__SCAN_IN), .ZN(n10208) );
  NAND2_X1 U11915 ( .A1(n10209), .A2(n10208), .ZN(n10267) );
  INV_X1 U11916 ( .A(P3_REG3_REG_13__SCAN_IN), .ZN(n11087) );
  NAND2_X1 U11917 ( .A1(n11088), .A2(n11087), .ZN(n11173) );
  OR2_X2 U11918 ( .A1(n11173), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n11270) );
  INV_X1 U11919 ( .A(P3_REG3_REG_16__SCAN_IN), .ZN(n11320) );
  INV_X1 U11920 ( .A(P3_REG3_REG_17__SCAN_IN), .ZN(n15204) );
  AND2_X1 U11921 ( .A1(n9504), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n9385) );
  OR2_X1 U11922 ( .A1(n9385), .A2(n11502), .ZN(n12260) );
  NAND2_X4 U11923 ( .A1(n9387), .A2(n9386), .ZN(n10012) );
  INV_X2 U11924 ( .A(n10012), .ZN(n11566) );
  NAND2_X1 U11925 ( .A1(n12260), .A2(n11566), .ZN(n9388) );
  OAI211_X1 U11926 ( .C1(n11570), .C2(n12488), .A(n9389), .B(n9388), .ZN(
        n11872) );
  NAND2_X1 U11927 ( .A1(n11872), .A2(P3_U3897), .ZN(n9390) );
  OAI21_X1 U11928 ( .B1(P3_U3897), .B2(n15277), .A(n9390), .ZN(P3_U3510) );
  INV_X1 U11929 ( .A(P3_DATAO_REG_2__SCAN_IN), .ZN(n15173) );
  INV_X1 U11930 ( .A(P3_REG1_REG_2__SCAN_IN), .ZN(n10044) );
  INV_X1 U11931 ( .A(P3_REG2_REG_2__SCAN_IN), .ZN(n10045) );
  OR2_X1 U11932 ( .A1(n6529), .A2(n10045), .ZN(n9391) );
  INV_X1 U11933 ( .A(P3_REG3_REG_2__SCAN_IN), .ZN(n15021) );
  NOR2_X1 U11934 ( .A1(n10012), .A2(n15021), .ZN(n9394) );
  INV_X1 U11935 ( .A(P3_REG0_REG_2__SCAN_IN), .ZN(n9392) );
  NOR2_X1 U11936 ( .A1(n9738), .A2(n9392), .ZN(n9393) );
  NAND2_X1 U11937 ( .A1(n15039), .A2(P3_U3897), .ZN(n9396) );
  OAI21_X1 U11938 ( .B1(P3_U3897), .B2(n15173), .A(n9396), .ZN(P3_U3493) );
  INV_X1 U11939 ( .A(n9397), .ZN(n9399) );
  OAI222_X1 U11940 ( .A1(P1_U3086), .A2(n9907), .B1(n6535), .B2(n9399), .C1(
        n9398), .C2(n14266), .ZN(P1_U3344) );
  OAI222_X1 U11941 ( .A1(P2_U3088), .A2(n9400), .B1(n6534), .B2(n9399), .C1(
        n15272), .C2(n11904), .ZN(P2_U3316) );
  INV_X1 U11942 ( .A(n14589), .ZN(n9750) );
  XNOR2_X1 U11943 ( .A(n9402), .B(n9401), .ZN(n9403) );
  NAND2_X1 U11944 ( .A1(n9403), .A2(n14395), .ZN(n9408) );
  NAND2_X1 U11945 ( .A1(n14556), .A2(n14107), .ZN(n9405) );
  NAND2_X1 U11946 ( .A1(n13771), .A2(n14108), .ZN(n9404) );
  NAND2_X1 U11947 ( .A1(n9405), .A2(n9404), .ZN(n9662) );
  AOI22_X1 U11948 ( .A1(n9406), .A2(P1_REG3_REG_2__SCAN_IN), .B1(n14397), .B2(
        n9662), .ZN(n9407) );
  OAI211_X1 U11949 ( .C1(n9750), .C2(n13743), .A(n9408), .B(n9407), .ZN(
        P1_U3237) );
  AND2_X1 U11950 ( .A1(n9410), .A2(n9409), .ZN(n9411) );
  NAND2_X1 U11951 ( .A1(n9412), .A2(n9411), .ZN(n9416) );
  INV_X1 U11952 ( .A(n14773), .ZN(n14770) );
  NOR2_X1 U11953 ( .A1(n9416), .A2(n14770), .ZN(n9423) );
  NAND2_X1 U11954 ( .A1(n9423), .A2(n9413), .ZN(n9414) );
  INV_X1 U11955 ( .A(n13019), .ZN(n14340) );
  INV_X1 U11956 ( .A(n12180), .ZN(n12235) );
  INV_X2 U11957 ( .A(n12948), .ZN(n14336) );
  NAND2_X1 U11958 ( .A1(n13051), .A2(n14336), .ZN(n9428) );
  INV_X1 U11959 ( .A(n9428), .ZN(n9418) );
  NAND2_X1 U11960 ( .A1(n9416), .A2(n9415), .ZN(n9556) );
  INV_X1 U11961 ( .A(n9433), .ZN(n9417) );
  NAND2_X1 U11962 ( .A1(n9556), .A2(n9417), .ZN(n9464) );
  AOI22_X1 U11963 ( .A1(n13016), .A2(n9418), .B1(P2_REG3_REG_0__SCAN_IN), .B2(
        n9464), .ZN(n9427) );
  NOR3_X1 U11964 ( .A1(n9419), .A2(n9550), .A3(n11935), .ZN(n9425) );
  OR2_X1 U11965 ( .A1(n9445), .A2(n11922), .ZN(n9420) );
  AND2_X1 U11966 ( .A1(n9546), .A2(n9420), .ZN(n9443) );
  INV_X1 U11967 ( .A(n9443), .ZN(n9424) );
  AND2_X1 U11968 ( .A1(n14806), .A2(n9421), .ZN(n9422) );
  OAI21_X1 U11969 ( .B1(n9425), .B2(n9424), .A(n12973), .ZN(n9426) );
  OAI211_X1 U11970 ( .C1(n14340), .C2(n11922), .A(n9427), .B(n9426), .ZN(
        P2_U3204) );
  INV_X1 U11971 ( .A(n6538), .ZN(n13307) );
  NOR2_X1 U11972 ( .A1(n13307), .A2(n13335), .ZN(n9429) );
  OAI21_X1 U11973 ( .B1(n11928), .B2(n11935), .A(n9541), .ZN(n12190) );
  OAI21_X1 U11974 ( .B1(n9429), .B2(n12190), .A(n9428), .ZN(n10353) );
  NOR2_X1 U11975 ( .A1(n8153), .A2(n12230), .ZN(n9430) );
  NAND2_X1 U11976 ( .A1(n9430), .A2(n13167), .ZN(n14803) );
  OAI22_X1 U11977 ( .A1(n12190), .A2(n14803), .B1(n9431), .B2(n11922), .ZN(
        n9432) );
  NOR2_X1 U11978 ( .A1(n10353), .A2(n9432), .ZN(n14775) );
  NOR2_X1 U11979 ( .A1(n9433), .A2(n14769), .ZN(n9434) );
  NAND2_X1 U11980 ( .A1(n14827), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n9436) );
  OAI21_X1 U11981 ( .B1(n14775), .B2(n14827), .A(n9436), .ZN(P2_U3499) );
  XNOR2_X1 U11982 ( .A(n9444), .B(n10453), .ZN(n9437) );
  NAND2_X1 U11983 ( .A1(n13050), .A2(n9445), .ZN(n9438) );
  NAND2_X1 U11984 ( .A1(n9437), .A2(n9438), .ZN(n9551) );
  INV_X1 U11985 ( .A(n9437), .ZN(n9440) );
  INV_X1 U11986 ( .A(n9438), .ZN(n9439) );
  NAND2_X1 U11987 ( .A1(n9440), .A2(n9439), .ZN(n9441) );
  AND2_X1 U11988 ( .A1(n9551), .A2(n9441), .ZN(n9451) );
  NAND2_X1 U11989 ( .A1(n12942), .A2(n11922), .ZN(n9442) );
  NAND2_X1 U11990 ( .A1(n9443), .A2(n9442), .ZN(n9459) );
  NAND2_X1 U11991 ( .A1(n13051), .A2(n9445), .ZN(n9447) );
  XNOR2_X1 U11992 ( .A(n9446), .B(n9447), .ZN(n9460) );
  NAND2_X1 U11993 ( .A1(n9459), .A2(n9460), .ZN(n9458) );
  INV_X1 U11994 ( .A(n9446), .ZN(n9448) );
  NAND2_X1 U11995 ( .A1(n9448), .A2(n9447), .ZN(n9449) );
  OAI21_X1 U11996 ( .B1(n9451), .B2(n9450), .A(n9552), .ZN(n9452) );
  NAND2_X1 U11997 ( .A1(n9452), .A2(n12973), .ZN(n9457) );
  INV_X2 U11998 ( .A(n12946), .ZN(n14334) );
  NAND2_X1 U11999 ( .A1(n13051), .A2(n14334), .ZN(n9454) );
  NAND2_X1 U12000 ( .A1(n13049), .A2(n14336), .ZN(n9453) );
  AND2_X1 U12001 ( .A1(n9454), .A2(n9453), .ZN(n9536) );
  INV_X1 U12002 ( .A(n9536), .ZN(n9455) );
  INV_X1 U12003 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n15227) );
  AOI22_X1 U12004 ( .A1(n13016), .A2(n9455), .B1(P2_REG3_REG_2__SCAN_IN), .B2(
        n9464), .ZN(n9456) );
  OAI211_X1 U12005 ( .C1(n10453), .C2(n14340), .A(n9457), .B(n9456), .ZN(
        P2_U3209) );
  OAI21_X1 U12006 ( .B1(n9460), .B2(n9459), .A(n9458), .ZN(n9461) );
  NAND2_X1 U12007 ( .A1(n9461), .A2(n12973), .ZN(n9467) );
  NAND2_X1 U12008 ( .A1(n11928), .A2(n14334), .ZN(n9463) );
  NAND2_X1 U12009 ( .A1(n13050), .A2(n14336), .ZN(n9462) );
  AND2_X1 U12010 ( .A1(n9463), .A2(n9462), .ZN(n9547) );
  INV_X1 U12011 ( .A(n9547), .ZN(n9465) );
  AOI22_X1 U12012 ( .A1(n13016), .A2(n9465), .B1(n9464), .B2(
        P2_REG3_REG_1__SCAN_IN), .ZN(n9466) );
  OAI211_X1 U12013 ( .C1(n10444), .C2(n14340), .A(n9467), .B(n9466), .ZN(
        P2_U3194) );
  INV_X1 U12014 ( .A(P3_DATAO_REG_21__SCAN_IN), .ZN(n15303) );
  INV_X1 U12015 ( .A(P3_REG3_REG_20__SCAN_IN), .ZN(n11501) );
  INV_X1 U12016 ( .A(P3_REG3_REG_21__SCAN_IN), .ZN(n9468) );
  OR2_X1 U12017 ( .A1(n11504), .A2(n9468), .ZN(n9469) );
  NAND2_X1 U12018 ( .A1(n11518), .A2(n9469), .ZN(n12607) );
  NAND2_X1 U12019 ( .A1(n12607), .A2(n11566), .ZN(n9472) );
  NAND2_X1 U12020 ( .A1(n11521), .A2(P3_REG1_REG_21__SCAN_IN), .ZN(n9470) );
  NAND2_X1 U12021 ( .A1(n12591), .A2(P3_U3897), .ZN(n9473) );
  OAI21_X1 U12022 ( .B1(P3_U3897), .B2(n15303), .A(n9473), .ZN(P3_U3512) );
  OAI21_X1 U12023 ( .B1(n9475), .B2(n10508), .A(n9474), .ZN(n9482) );
  INV_X1 U12024 ( .A(n9482), .ZN(n9480) );
  NOR2_X1 U12025 ( .A1(n14464), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n9479) );
  INV_X1 U12026 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n14415) );
  NOR3_X1 U12027 ( .A1(n9488), .A2(n14415), .A3(n14459), .ZN(n9478) );
  AOI211_X1 U12028 ( .C1(n9480), .C2(n9479), .A(n14476), .B(n9478), .ZN(n9492)
         );
  AND2_X1 U12029 ( .A1(P1_U3086), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n11028) );
  AOI21_X1 U12030 ( .B1(n9907), .B2(P1_REG2_REG_11__SCAN_IN), .A(n9482), .ZN(
        n9484) );
  MUX2_X1 U12031 ( .A(n10817), .B(P1_REG2_REG_11__SCAN_IN), .S(n9907), .Z(
        n9481) );
  NAND2_X1 U12032 ( .A1(n9482), .A2(n9481), .ZN(n9906) );
  INV_X1 U12033 ( .A(n9906), .ZN(n9483) );
  NOR3_X1 U12034 ( .A1(n9484), .A2(n9483), .A3(n14464), .ZN(n9485) );
  AOI211_X1 U12035 ( .C1(n14472), .C2(P1_ADDR_REG_11__SCAN_IN), .A(n11028), 
        .B(n9485), .ZN(n9491) );
  NOR3_X1 U12036 ( .A1(n9488), .A2(n9486), .A3(P1_REG1_REG_11__SCAN_IN), .ZN(
        n9489) );
  MUX2_X1 U12037 ( .A(n14415), .B(P1_REG1_REG_11__SCAN_IN), .S(n9907), .Z(
        n9487) );
  OAI21_X1 U12038 ( .B1(n9489), .B2(n9898), .A(n14483), .ZN(n9490) );
  OAI211_X1 U12039 ( .C1(n9492), .C2(n9907), .A(n9491), .B(n9490), .ZN(
        P1_U3254) );
  NAND2_X1 U12040 ( .A1(n9915), .A2(P1_DATAO_REG_16__SCAN_IN), .ZN(n9527) );
  NAND2_X1 U12041 ( .A1(n15181), .A2(P2_DATAO_REG_16__SCAN_IN), .ZN(n9495) );
  AND2_X1 U12042 ( .A1(n9527), .A2(n9495), .ZN(n9496) );
  OR2_X1 U12043 ( .A1(n9497), .A2(n9496), .ZN(n9498) );
  AND2_X1 U12044 ( .A1(n9498), .A2(n9528), .ZN(n11426) );
  INV_X1 U12045 ( .A(n9499), .ZN(n9500) );
  NAND2_X1 U12046 ( .A1(n9500), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9501) );
  XNOR2_X1 U12047 ( .A(n9501), .B(P3_IR_REG_16__SCAN_IN), .ZN(n12453) );
  AOI222_X1 U12048 ( .A1(n11426), .A2(n12881), .B1(n12453), .B2(
        P3_STATE_REG_SCAN_IN), .C1(SI_16_), .C2(n10122), .ZN(n9502) );
  INV_X1 U12049 ( .A(n9502), .ZN(P3_U3279) );
  INV_X1 U12050 ( .A(P3_DATAO_REG_18__SCAN_IN), .ZN(n15310) );
  NAND2_X1 U12051 ( .A1(n11435), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n9503) );
  NAND2_X1 U12052 ( .A1(n9504), .A2(n9503), .ZN(n12653) );
  NAND2_X1 U12053 ( .A1(n11566), .A2(n12653), .ZN(n9508) );
  INV_X1 U12054 ( .A(P3_REG2_REG_18__SCAN_IN), .ZN(n12472) );
  INV_X1 U12055 ( .A(P3_REG0_REG_18__SCAN_IN), .ZN(n15154) );
  OR2_X1 U12056 ( .A1(n11438), .A2(n15154), .ZN(n9506) );
  INV_X1 U12057 ( .A(P3_REG1_REG_18__SCAN_IN), .ZN(n12765) );
  OR2_X1 U12058 ( .A1(n11570), .A2(n12765), .ZN(n9505) );
  NAND2_X1 U12059 ( .A1(n12665), .A2(P3_U3897), .ZN(n9509) );
  OAI21_X1 U12060 ( .B1(P3_U3897), .B2(n15310), .A(n9509), .ZN(P3_U3509) );
  INV_X1 U12061 ( .A(n9510), .ZN(n9513) );
  OAI222_X1 U12062 ( .A1(P2_U3088), .A2(n14732), .B1(n6534), .B2(n9513), .C1(
        n9511), .C2(n11904), .ZN(P2_U3315) );
  INV_X1 U12063 ( .A(n14461), .ZN(n9905) );
  OAI222_X1 U12064 ( .A1(P1_U3086), .A2(n9905), .B1(n6535), .B2(n9513), .C1(
        n9512), .C2(n14266), .ZN(P1_U3343) );
  INV_X1 U12065 ( .A(n9514), .ZN(n9516) );
  OAI222_X1 U12066 ( .A1(P1_U3086), .A2(n14471), .B1(n6535), .B2(n9516), .C1(
        n9515), .C2(n14266), .ZN(P1_U3342) );
  INV_X1 U12067 ( .A(n10160), .ZN(n14738) );
  OAI222_X1 U12068 ( .A1(P2_U3088), .A2(n14738), .B1(n6534), .B2(n9516), .C1(
        n15367), .C2(n11904), .ZN(P2_U3314) );
  OAI21_X1 U12069 ( .B1(n9518), .B2(n12194), .A(n9517), .ZN(n10227) );
  AOI211_X1 U12070 ( .C1(n11965), .C2(n9532), .A(n9445), .B(n9567), .ZN(n10231) );
  XNOR2_X1 U12071 ( .A(n9519), .B(n12194), .ZN(n9522) );
  NAND2_X1 U12072 ( .A1(n13050), .A2(n14334), .ZN(n9521) );
  NAND2_X1 U12073 ( .A1(n13048), .A2(n14336), .ZN(n9520) );
  AND2_X1 U12074 ( .A1(n9521), .A2(n9520), .ZN(n9558) );
  OAI21_X1 U12075 ( .B1(n9522), .B2(n14351), .A(n9558), .ZN(n10232) );
  AOI211_X1 U12076 ( .C1(n14378), .C2(n10227), .A(n10231), .B(n10232), .ZN(
        n9650) );
  NAND2_X1 U12077 ( .A1(n14829), .A2(n14810), .ZN(n13423) );
  INV_X1 U12078 ( .A(n13423), .ZN(n13398) );
  AOI22_X1 U12079 ( .A1(n13398), .A2(n11965), .B1(n14827), .B2(
        P2_REG1_REG_3__SCAN_IN), .ZN(n9523) );
  OAI21_X1 U12080 ( .B1(n9650), .B2(n14827), .A(n9523), .ZN(P2_U3502) );
  NAND2_X1 U12081 ( .A1(n9524), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9526) );
  INV_X1 U12082 ( .A(P3_IR_REG_17__SCAN_IN), .ZN(n9525) );
  XNOR2_X1 U12083 ( .A(n9526), .B(n9525), .ZN(n12465) );
  NAND2_X1 U12084 ( .A1(n9959), .A2(P1_DATAO_REG_17__SCAN_IN), .ZN(n9617) );
  NAND2_X1 U12085 ( .A1(n9961), .A2(P2_DATAO_REG_17__SCAN_IN), .ZN(n9529) );
  AND2_X1 U12086 ( .A1(n9617), .A2(n9529), .ZN(n9615) );
  XNOR2_X1 U12087 ( .A(n9616), .B(n9615), .ZN(n11484) );
  INV_X1 U12088 ( .A(SI_17_), .ZN(n11485) );
  OAI222_X1 U12089 ( .A1(n12465), .A2(P3_U3151), .B1(n12245), .B2(n11484), 
        .C1(n11485), .C2(n11338), .ZN(P3_U3278) );
  OAI21_X1 U12090 ( .B1(n9531), .B2(n9534), .A(n9530), .ZN(n10455) );
  INV_X1 U12091 ( .A(n9532), .ZN(n9533) );
  AOI211_X1 U12092 ( .C1(n6524), .C2(n9542), .A(n9445), .B(n9533), .ZN(n10450)
         );
  XNOR2_X1 U12093 ( .A(n9535), .B(n9534), .ZN(n9537) );
  OAI21_X1 U12094 ( .B1(n9537), .B2(n14351), .A(n9536), .ZN(n10449) );
  AOI211_X1 U12095 ( .C1(n14378), .C2(n10455), .A(n10450), .B(n10449), .ZN(
        n9647) );
  AOI22_X1 U12096 ( .A1(n13398), .A2(n6524), .B1(n14827), .B2(
        P2_REG1_REG_2__SCAN_IN), .ZN(n9538) );
  OAI21_X1 U12097 ( .B1(n9647), .B2(n14827), .A(n9538), .ZN(P2_U3501) );
  OAI21_X1 U12098 ( .B1(n9539), .B2(n9541), .A(n9540), .ZN(n10446) );
  AOI21_X1 U12099 ( .B1(n11935), .B2(n11932), .A(n9445), .ZN(n9543) );
  AND2_X1 U12100 ( .A1(n9543), .A2(n9542), .ZN(n10442) );
  INV_X1 U12101 ( .A(n9544), .ZN(n9545) );
  AOI21_X1 U12102 ( .B1(n9539), .B2(n9546), .A(n9545), .ZN(n9548) );
  OAI21_X1 U12103 ( .B1(n9548), .B2(n14351), .A(n9547), .ZN(n10440) );
  AOI211_X1 U12104 ( .C1(n14378), .C2(n10446), .A(n10442), .B(n10440), .ZN(
        n9653) );
  AOI22_X1 U12105 ( .A1(n13398), .A2(n11932), .B1(n14827), .B2(
        P2_REG1_REG_1__SCAN_IN), .ZN(n9549) );
  OAI21_X1 U12106 ( .B1(n9653), .B2(n14827), .A(n9549), .ZN(P2_U3500) );
  AND2_X1 U12107 ( .A1(n13049), .A2(n9445), .ZN(n9577) );
  XNOR2_X1 U12108 ( .A(n9576), .B(n9575), .ZN(n9564) );
  AND3_X1 U12109 ( .A1(n9554), .A2(n11011), .A3(n9553), .ZN(n9555) );
  NAND2_X1 U12110 ( .A1(n9556), .A2(n9555), .ZN(n9557) );
  INV_X1 U12111 ( .A(n14348), .ZN(n13000) );
  NAND2_X1 U12112 ( .A1(n13019), .A2(n11965), .ZN(n9561) );
  NAND2_X1 U12113 ( .A1(P2_U3088), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n13073) );
  INV_X1 U12114 ( .A(n9558), .ZN(n9559) );
  NAND2_X1 U12115 ( .A1(n13016), .A2(n9559), .ZN(n9560) );
  NAND3_X1 U12116 ( .A1(n9561), .A2(n13073), .A3(n9560), .ZN(n9562) );
  AOI21_X1 U12117 ( .B1(n13000), .B2(n7654), .A(n9562), .ZN(n9563) );
  OAI21_X1 U12118 ( .B1(n9564), .B2(n14342), .A(n9563), .ZN(P2_U3190) );
  OAI21_X1 U12119 ( .B1(n9566), .B2(n9569), .A(n9565), .ZN(n10125) );
  INV_X1 U12120 ( .A(n9567), .ZN(n9568) );
  AOI211_X1 U12121 ( .C1(n11973), .C2(n9568), .A(n9445), .B(n6706), .ZN(n10132) );
  XNOR2_X1 U12122 ( .A(n9570), .B(n9569), .ZN(n9573) );
  NAND2_X1 U12123 ( .A1(n13049), .A2(n14334), .ZN(n9572) );
  NAND2_X1 U12124 ( .A1(n13047), .A2(n14336), .ZN(n9571) );
  AND2_X1 U12125 ( .A1(n9572), .A2(n9571), .ZN(n9586) );
  OAI21_X1 U12126 ( .B1(n9573), .B2(n14351), .A(n9586), .ZN(n10126) );
  AOI211_X1 U12127 ( .C1(n14378), .C2(n10125), .A(n10132), .B(n10126), .ZN(
        n9644) );
  AOI22_X1 U12128 ( .A1(n13398), .A2(n11973), .B1(n14827), .B2(
        P2_REG1_REG_4__SCAN_IN), .ZN(n9574) );
  OAI21_X1 U12129 ( .B1(n9644), .B2(n14827), .A(n9574), .ZN(P2_U3503) );
  INV_X1 U12130 ( .A(n9598), .ZN(n9585) );
  XNOR2_X1 U12131 ( .A(n11973), .B(n6528), .ZN(n9582) );
  INV_X1 U12132 ( .A(n9582), .ZN(n9580) );
  AND2_X1 U12133 ( .A1(n13048), .A2(n12940), .ZN(n9581) );
  INV_X1 U12134 ( .A(n9581), .ZN(n9579) );
  AND2_X1 U12135 ( .A1(n9580), .A2(n9579), .ZN(n9774) );
  INV_X1 U12136 ( .A(n9774), .ZN(n9583) );
  NAND2_X1 U12137 ( .A1(n9582), .A2(n9581), .ZN(n9597) );
  NAND2_X1 U12138 ( .A1(n9583), .A2(n9597), .ZN(n9584) );
  NOR2_X1 U12139 ( .A1(n9585), .A2(n9584), .ZN(n9775) );
  AOI21_X1 U12140 ( .B1(n9585), .B2(n9584), .A(n9775), .ZN(n9592) );
  NOR2_X1 U12141 ( .A1(n14348), .A2(n10129), .ZN(n9590) );
  INV_X1 U12142 ( .A(n9586), .ZN(n9587) );
  NAND2_X1 U12143 ( .A1(n13016), .A2(n9587), .ZN(n9588) );
  NAND2_X1 U12144 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_U3088), .ZN(n14659) );
  NAND2_X1 U12145 ( .A1(n9588), .A2(n14659), .ZN(n9589) );
  AOI211_X1 U12146 ( .C1(n11973), .C2(n13019), .A(n9590), .B(n9589), .ZN(n9591) );
  OAI21_X1 U12147 ( .B1(n9592), .B2(n14342), .A(n9591), .ZN(P2_U3202) );
  INV_X1 U12148 ( .A(n10163), .ZN(n10736) );
  INV_X1 U12149 ( .A(n9593), .ZN(n9596) );
  OAI222_X1 U12150 ( .A1(P2_U3088), .A2(n10736), .B1(n6534), .B2(n9596), .C1(
        n9594), .C2(n11904), .ZN(P2_U3313) );
  INV_X1 U12151 ( .A(n10336), .ZN(n10341) );
  OAI222_X1 U12152 ( .A1(P1_U3086), .A2(n10341), .B1(n6535), .B2(n9596), .C1(
        n9595), .C2(n14266), .ZN(P1_U3341) );
  XNOR2_X1 U12153 ( .A(n11980), .B(n6528), .ZN(n9599) );
  AND2_X1 U12154 ( .A1(n13047), .A2(n13326), .ZN(n9600) );
  NAND2_X1 U12155 ( .A1(n9599), .A2(n9600), .ZN(n9773) );
  NAND3_X1 U12156 ( .A1(n9598), .A2(n9773), .A3(n9597), .ZN(n9605) );
  NAND2_X1 U12157 ( .A1(n9773), .A2(n9774), .ZN(n9603) );
  INV_X1 U12158 ( .A(n9599), .ZN(n9602) );
  INV_X1 U12159 ( .A(n9600), .ZN(n9601) );
  NAND2_X1 U12160 ( .A1(n9602), .A2(n9601), .ZN(n9772) );
  AND2_X1 U12161 ( .A1(n9603), .A2(n9772), .ZN(n9604) );
  XNOR2_X1 U12162 ( .A(n14782), .B(n12915), .ZN(n9825) );
  NAND2_X1 U12163 ( .A1(n13046), .A2(n13326), .ZN(n9826) );
  XNOR2_X1 U12164 ( .A(n9825), .B(n9826), .ZN(n9830) );
  XNOR2_X1 U12165 ( .A(n9831), .B(n9830), .ZN(n9612) );
  NAND2_X1 U12166 ( .A1(n13047), .A2(n14334), .ZN(n9607) );
  NAND2_X1 U12167 ( .A1(n13045), .A2(n14336), .ZN(n9606) );
  NAND2_X1 U12168 ( .A1(n9607), .A2(n9606), .ZN(n10143) );
  NAND2_X1 U12169 ( .A1(n13016), .A2(n10143), .ZN(n9609) );
  OAI211_X1 U12170 ( .C1(n14348), .C2(n10146), .A(n9609), .B(n9608), .ZN(n9610) );
  AOI21_X1 U12171 ( .B1(n14782), .B2(n13019), .A(n9610), .ZN(n9611) );
  OAI21_X1 U12172 ( .B1(n9612), .B2(n14342), .A(n9611), .ZN(P2_U3211) );
  NOR2_X2 U12173 ( .A1(n9524), .A2(P3_IR_REG_17__SCAN_IN), .ZN(n9632) );
  INV_X1 U12174 ( .A(n9632), .ZN(n9613) );
  NAND2_X1 U12175 ( .A1(n9613), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9614) );
  XNOR2_X1 U12176 ( .A(n9614), .B(P3_IR_REG_18__SCAN_IN), .ZN(n12494) );
  INV_X1 U12177 ( .A(n12494), .ZN(n9621) );
  INV_X1 U12178 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n10461) );
  NAND2_X1 U12179 ( .A1(n10461), .A2(P1_DATAO_REG_18__SCAN_IN), .ZN(n9625) );
  INV_X1 U12180 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n10463) );
  NAND2_X1 U12181 ( .A1(n10463), .A2(P2_DATAO_REG_18__SCAN_IN), .ZN(n9618) );
  NAND2_X1 U12182 ( .A1(n9625), .A2(n9618), .ZN(n9622) );
  XNOR2_X1 U12183 ( .A(n9624), .B(n9622), .ZN(n11488) );
  INV_X1 U12184 ( .A(n11488), .ZN(n9620) );
  OAI222_X1 U12185 ( .A1(n9621), .A2(P3_U3151), .B1(n12245), .B2(n9620), .C1(
        n9619), .C2(n11338), .ZN(P3_U3277) );
  INV_X1 U12186 ( .A(n9622), .ZN(n9623) );
  INV_X1 U12187 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n10657) );
  NAND2_X1 U12188 ( .A1(n10657), .A2(P1_DATAO_REG_19__SCAN_IN), .ZN(n9676) );
  INV_X1 U12189 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n11909) );
  NAND2_X1 U12190 ( .A1(n11909), .A2(P2_DATAO_REG_19__SCAN_IN), .ZN(n9627) );
  AND2_X1 U12191 ( .A1(n9676), .A2(n9627), .ZN(n9628) );
  OR2_X1 U12192 ( .A1(n9629), .A2(n9628), .ZN(n9630) );
  NAND2_X1 U12193 ( .A1(n9677), .A2(n9630), .ZN(n11491) );
  INV_X1 U12194 ( .A(P3_IR_REG_18__SCAN_IN), .ZN(n9631) );
  INV_X1 U12195 ( .A(n9683), .ZN(n9633) );
  NAND2_X1 U12196 ( .A1(n9633), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9634) );
  OAI222_X1 U12197 ( .A1(n12245), .A2(n11491), .B1(n11338), .B2(n15312), .C1(
        P3_U3151), .C2(n12501), .ZN(P3_U3276) );
  INV_X1 U12198 ( .A(P3_DATAO_REG_23__SCAN_IN), .ZN(n15235) );
  NAND2_X1 U12199 ( .A1(n11520), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n9635) );
  NAND2_X1 U12200 ( .A1(n11533), .A2(n9635), .ZN(n12583) );
  NAND2_X1 U12201 ( .A1(n12583), .A2(n11566), .ZN(n9640) );
  INV_X1 U12202 ( .A(P3_REG1_REG_23__SCAN_IN), .ZN(n15174) );
  NAND2_X1 U12203 ( .A1(n11567), .A2(P3_REG2_REG_23__SCAN_IN), .ZN(n9637) );
  OAI211_X1 U12204 ( .C1(n15174), .C2(n11570), .A(n9637), .B(n9636), .ZN(n9638) );
  INV_X1 U12205 ( .A(n9638), .ZN(n9639) );
  NAND2_X1 U12206 ( .A1(n12592), .A2(P3_U3897), .ZN(n9641) );
  OAI21_X1 U12207 ( .B1(P3_U3897), .B2(n15235), .A(n9641), .ZN(P3_U3514) );
  OAI22_X1 U12208 ( .A1(n13468), .A2(n10130), .B1(n14821), .B2(n7657), .ZN(
        n9642) );
  INV_X1 U12209 ( .A(n9642), .ZN(n9643) );
  OAI21_X1 U12210 ( .B1(n9644), .B2(n14819), .A(n9643), .ZN(P2_U3442) );
  OAI22_X1 U12211 ( .A1(n13468), .A2(n10453), .B1(n14821), .B2(n7606), .ZN(
        n9645) );
  INV_X1 U12212 ( .A(n9645), .ZN(n9646) );
  OAI21_X1 U12213 ( .B1(n9647), .B2(n14819), .A(n9646), .ZN(P2_U3436) );
  OAI22_X1 U12214 ( .A1(n13468), .A2(n10228), .B1(n14821), .B2(n7624), .ZN(
        n9648) );
  INV_X1 U12215 ( .A(n9648), .ZN(n9649) );
  OAI21_X1 U12216 ( .B1(n9650), .B2(n14819), .A(n9649), .ZN(P2_U3439) );
  OAI22_X1 U12217 ( .A1(n13468), .A2(n10444), .B1(n14821), .B2(n7577), .ZN(
        n9651) );
  INV_X1 U12218 ( .A(n9651), .ZN(n9652) );
  OAI21_X1 U12219 ( .B1(n9653), .B2(n14819), .A(n9652), .ZN(P2_U3433) );
  INV_X1 U12220 ( .A(n9654), .ZN(n14552) );
  XNOR2_X1 U12221 ( .A(n9749), .B(n9757), .ZN(n14593) );
  INV_X1 U12222 ( .A(n14593), .ZN(n14595) );
  NAND3_X1 U12223 ( .A1(n9657), .A2(n9656), .A3(n9655), .ZN(n13921) );
  INV_X1 U12224 ( .A(n9658), .ZN(n9659) );
  NOR2_X2 U12225 ( .A1(n6531), .A2(n9659), .ZN(n14083) );
  XNOR2_X1 U12226 ( .A(n9758), .B(n9757), .ZN(n9663) );
  AOI21_X1 U12227 ( .B1(n9663), .B2(n14497), .A(n9662), .ZN(n14591) );
  NOR2_X2 U12228 ( .A1(n6531), .A2(n9664), .ZN(n14566) );
  NAND2_X1 U12229 ( .A1(n6531), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n9665) );
  OAI21_X1 U12230 ( .B1(n14542), .B2(n9666), .A(n9665), .ZN(n9667) );
  AOI21_X1 U12231 ( .B1(n14566), .B2(n14589), .A(n9667), .ZN(n9673) );
  INV_X1 U12232 ( .A(n13921), .ZN(n9668) );
  NAND2_X1 U12233 ( .A1(n9668), .A2(n13847), .ZN(n13959) );
  NAND2_X1 U12234 ( .A1(n14580), .A2(n9669), .ZN(n14555) );
  NAND2_X1 U12235 ( .A1(n14555), .A2(n14589), .ZN(n9670) );
  INV_X1 U12236 ( .A(n14572), .ZN(n14546) );
  NAND2_X1 U12237 ( .A1(n9670), .A2(n14546), .ZN(n9671) );
  NOR2_X1 U12238 ( .A1(n14548), .A2(n9671), .ZN(n14588) );
  NAND2_X1 U12239 ( .A1(n14574), .A2(n14588), .ZN(n9672) );
  OAI211_X1 U12240 ( .C1(n14591), .C2(n6531), .A(n9673), .B(n9672), .ZN(n9674)
         );
  AOI21_X1 U12241 ( .B1(n14595), .B2(n14083), .A(n9674), .ZN(n9675) );
  INV_X1 U12242 ( .A(n9675), .ZN(P1_U3291) );
  NAND2_X1 U12243 ( .A1(n15263), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n10027) );
  NAND2_X1 U12244 ( .A1(n10497), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n9678) );
  AND2_X1 U12245 ( .A1(n10027), .A2(n9678), .ZN(n9679) );
  OR2_X1 U12246 ( .A1(n9680), .A2(n9679), .ZN(n9681) );
  NAND2_X1 U12247 ( .A1(n10028), .A2(n9681), .ZN(n11497) );
  INV_X1 U12248 ( .A(SI_20_), .ZN(n11498) );
  INV_X1 U12249 ( .A(n9701), .ZN(n9684) );
  NAND2_X1 U12250 ( .A1(n9684), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9685) );
  XNOR2_X2 U12251 ( .A(n9685), .B(n9700), .ZN(n9817) );
  OAI222_X1 U12252 ( .A1(n12245), .A2(n11497), .B1(n11338), .B2(n11498), .C1(
        P3_U3151), .C2(n9817), .ZN(P3_U3275) );
  NAND2_X1 U12253 ( .A1(n9789), .A2(n9805), .ZN(n9788) );
  NOR2_X1 U12254 ( .A1(P3_D_REG_5__SCAN_IN), .A2(P3_D_REG_12__SCAN_IN), .ZN(
        n15105) );
  NOR4_X1 U12255 ( .A1(P3_D_REG_2__SCAN_IN), .A2(P3_D_REG_7__SCAN_IN), .A3(
        P3_D_REG_8__SCAN_IN), .A4(P3_D_REG_15__SCAN_IN), .ZN(n9692) );
  NOR4_X1 U12256 ( .A1(P3_D_REG_20__SCAN_IN), .A2(P3_D_REG_19__SCAN_IN), .A3(
        P3_D_REG_18__SCAN_IN), .A4(P3_D_REG_27__SCAN_IN), .ZN(n9691) );
  NOR4_X1 U12257 ( .A1(P3_D_REG_6__SCAN_IN), .A2(P3_D_REG_17__SCAN_IN), .A3(
        P3_D_REG_22__SCAN_IN), .A4(P3_D_REG_25__SCAN_IN), .ZN(n9690) );
  NAND4_X1 U12258 ( .A1(n15105), .A2(n9692), .A3(n9691), .A4(n9690), .ZN(n9698) );
  NOR4_X1 U12259 ( .A1(P3_D_REG_31__SCAN_IN), .A2(P3_D_REG_21__SCAN_IN), .A3(
        P3_D_REG_11__SCAN_IN), .A4(P3_D_REG_26__SCAN_IN), .ZN(n9696) );
  NOR4_X1 U12260 ( .A1(P3_D_REG_24__SCAN_IN), .A2(P3_D_REG_29__SCAN_IN), .A3(
        P3_D_REG_14__SCAN_IN), .A4(P3_D_REG_10__SCAN_IN), .ZN(n9695) );
  NOR4_X1 U12261 ( .A1(P3_D_REG_28__SCAN_IN), .A2(P3_D_REG_23__SCAN_IN), .A3(
        P3_D_REG_3__SCAN_IN), .A4(P3_D_REG_4__SCAN_IN), .ZN(n9694) );
  NOR4_X1 U12262 ( .A1(P3_D_REG_9__SCAN_IN), .A2(P3_D_REG_13__SCAN_IN), .A3(
        P3_D_REG_16__SCAN_IN), .A4(P3_D_REG_30__SCAN_IN), .ZN(n9693) );
  NAND4_X1 U12263 ( .A1(n9696), .A2(n9695), .A3(n9694), .A4(n9693), .ZN(n9697)
         );
  AND2_X1 U12264 ( .A1(n9790), .A2(n10396), .ZN(n9699) );
  INV_X1 U12265 ( .A(P3_IR_REG_22__SCAN_IN), .ZN(n9702) );
  NAND2_X1 U12266 ( .A1(n9708), .A2(n12489), .ZN(n9792) );
  NAND2_X1 U12267 ( .A1(n9792), .A2(n11853), .ZN(n9707) );
  INV_X1 U12268 ( .A(P3_IR_REG_21__SCAN_IN), .ZN(n9705) );
  NAND2_X1 U12269 ( .A1(n6527), .A2(n9817), .ZN(n9733) );
  AOI22_X1 U12270 ( .A1(n9707), .A2(n6527), .B1(n11860), .B2(n9733), .ZN(n9711) );
  NAND2_X2 U12271 ( .A1(n9708), .A2(n9736), .ZN(n11815) );
  OR2_X1 U12272 ( .A1(n11815), .A2(n9799), .ZN(n9794) );
  OR3_X1 U12273 ( .A1(n11860), .A2(n9817), .A3(n12489), .ZN(n10092) );
  NAND2_X1 U12274 ( .A1(n11815), .A2(n10092), .ZN(n10083) );
  NAND2_X1 U12275 ( .A1(n9794), .A2(n10083), .ZN(n10086) );
  INV_X1 U12276 ( .A(n10086), .ZN(n9709) );
  NAND2_X1 U12277 ( .A1(n9709), .A2(n9789), .ZN(n9710) );
  OAI21_X1 U12278 ( .B1(n10085), .B2(n9711), .A(n9710), .ZN(n9712) );
  NAND2_X1 U12279 ( .A1(n11566), .A2(P3_REG3_REG_0__SCAN_IN), .ZN(n9717) );
  INV_X1 U12280 ( .A(P3_REG1_REG_0__SCAN_IN), .ZN(n9713) );
  INV_X1 U12281 ( .A(P3_REG2_REG_0__SCAN_IN), .ZN(n15205) );
  OR2_X1 U12282 ( .A1(n6530), .A2(n15205), .ZN(n9714) );
  OR2_X1 U12283 ( .A1(n9723), .A2(n9718), .ZN(n9720) );
  NAND2_X1 U12284 ( .A1(n9721), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9722) );
  MUX2_X2 U12285 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9722), .S(
        P3_IR_REG_27__SCAN_IN), .Z(n9725) );
  INV_X1 U12286 ( .A(n9723), .ZN(n9724) );
  NAND2_X4 U12287 ( .A1(n9725), .A2(n9724), .ZN(n12463) );
  OR2_X1 U12288 ( .A1(n10001), .A2(n9730), .ZN(n9731) );
  OAI211_X1 U12289 ( .C1(n9883), .C2(n10530), .A(n9732), .B(n9731), .ZN(n10061) );
  INV_X1 U12290 ( .A(n10061), .ZN(n11634) );
  NAND2_X1 U12291 ( .A1(n15040), .A2(n11634), .ZN(n11684) );
  AND2_X1 U12292 ( .A1(n10094), .A2(n11684), .ZN(n11829) );
  XNOR2_X1 U12293 ( .A(n11860), .B(n9733), .ZN(n9735) );
  AND2_X1 U12294 ( .A1(n6527), .A2(n12501), .ZN(n9734) );
  OR2_X1 U12295 ( .A1(n9735), .A2(n9734), .ZN(n10392) );
  NAND2_X1 U12296 ( .A1(n10392), .A2(n15018), .ZN(n10091) );
  INV_X1 U12297 ( .A(n9817), .ZN(n9791) );
  NAND2_X1 U12298 ( .A1(n9736), .A2(n9791), .ZN(n11672) );
  AND2_X1 U12299 ( .A1(n10091), .A2(n15027), .ZN(n9745) );
  NAND2_X1 U12300 ( .A1(n11521), .A2(P3_REG1_REG_1__SCAN_IN), .ZN(n9744) );
  INV_X1 U12301 ( .A(P3_REG0_REG_1__SCAN_IN), .ZN(n9737) );
  INV_X1 U12302 ( .A(P3_REG2_REG_1__SCAN_IN), .ZN(n9739) );
  OR2_X1 U12303 ( .A1(n6529), .A2(n9739), .ZN(n9742) );
  INV_X1 U12304 ( .A(P3_REG3_REG_1__SCAN_IN), .ZN(n9982) );
  OR2_X1 U12305 ( .A1(n10012), .A2(n9982), .ZN(n9741) );
  INV_X1 U12306 ( .A(n12242), .ZN(n11620) );
  INV_X1 U12307 ( .A(n12463), .ZN(n12490) );
  NAND2_X1 U12308 ( .A1(n11620), .A2(n12490), .ZN(n9878) );
  AND2_X1 U12309 ( .A1(n10530), .A2(n9878), .ZN(n9820) );
  OAI22_X1 U12310 ( .A1(n11829), .A2(n9745), .B1(n15028), .B2(n15031), .ZN(
        n11631) );
  OAI22_X1 U12311 ( .A1(n12780), .A2(n11634), .B1(n15096), .B2(n9713), .ZN(
        n9746) );
  AOI21_X1 U12312 ( .B1(n15096), .B2(n11631), .A(n9746), .ZN(n9747) );
  INV_X1 U12313 ( .A(n9747), .ZN(P3_U3459) );
  INV_X1 U12314 ( .A(n9757), .ZN(n9748) );
  NAND2_X1 U12315 ( .A1(n14582), .A2(n9750), .ZN(n9751) );
  NAND2_X1 U12316 ( .A1(n9752), .A2(n9751), .ZN(n14536) );
  INV_X1 U12317 ( .A(n9761), .ZN(n14538) );
  NAND2_X1 U12318 ( .A1(n14536), .A2(n14538), .ZN(n9755) );
  NAND2_X1 U12319 ( .A1(n14599), .A2(n9753), .ZN(n9754) );
  NAND2_X1 U12320 ( .A1(n9755), .A2(n9754), .ZN(n9853) );
  XNOR2_X1 U12321 ( .A(n9853), .B(n9860), .ZN(n14610) );
  INV_X1 U12322 ( .A(n9756), .ZN(n14547) );
  AOI211_X1 U12323 ( .C1(n14608), .C2(n14547), .A(n14572), .B(n14532), .ZN(
        n14606) );
  NAND2_X1 U12324 ( .A1(n9758), .A2(n9757), .ZN(n9760) );
  NAND2_X1 U12325 ( .A1(n14582), .A2(n14589), .ZN(n9759) );
  NAND2_X1 U12326 ( .A1(n9760), .A2(n9759), .ZN(n14537) );
  NAND2_X1 U12327 ( .A1(n14537), .A2(n9761), .ZN(n9763) );
  NAND2_X1 U12328 ( .A1(n9763), .A2(n9762), .ZN(n9861) );
  XNOR2_X1 U12329 ( .A(n9861), .B(n9852), .ZN(n9766) );
  NAND2_X1 U12330 ( .A1(n13771), .A2(n14107), .ZN(n9764) );
  OAI21_X1 U12331 ( .B1(n9866), .B2(n14581), .A(n9764), .ZN(n9929) );
  INV_X1 U12332 ( .A(n9929), .ZN(n9765) );
  OAI21_X1 U12333 ( .B1(n9766), .B2(n14560), .A(n9765), .ZN(n14605) );
  AOI21_X1 U12334 ( .B1(n14606), .B2(n13847), .A(n14605), .ZN(n9767) );
  MUX2_X1 U12335 ( .A(n9768), .B(n9767), .S(n14543), .Z(n9771) );
  INV_X1 U12336 ( .A(n9932), .ZN(n9769) );
  AOI22_X1 U12337 ( .A1(n14566), .A2(n14608), .B1(n14567), .B2(n9769), .ZN(
        n9770) );
  OAI211_X1 U12338 ( .C1(n14123), .C2(n14610), .A(n9771), .B(n9770), .ZN(
        P1_U3289) );
  NAND2_X1 U12339 ( .A1(n9773), .A2(n9772), .ZN(n9777) );
  NOR2_X1 U12340 ( .A1(n9775), .A2(n9774), .ZN(n9776) );
  XOR2_X1 U12341 ( .A(n9777), .B(n9776), .Z(n9783) );
  NAND2_X1 U12342 ( .A1(n13046), .A2(n14336), .ZN(n9779) );
  NAND2_X1 U12343 ( .A1(n13048), .A2(n14334), .ZN(n9778) );
  NAND2_X1 U12344 ( .A1(n9779), .A2(n9778), .ZN(n10169) );
  NAND2_X1 U12345 ( .A1(n13016), .A2(n10169), .ZN(n9780) );
  NAND2_X1 U12346 ( .A1(P2_REG3_REG_5__SCAN_IN), .A2(P2_U3088), .ZN(n14673) );
  OAI211_X1 U12347 ( .C1(n14348), .C2(n10173), .A(n9780), .B(n14673), .ZN(
        n9781) );
  AOI21_X1 U12348 ( .B1(n11980), .B2(n13019), .A(n9781), .ZN(n9782) );
  OAI21_X1 U12349 ( .B1(n9783), .B2(n14342), .A(n9782), .ZN(P2_U3199) );
  INV_X1 U12350 ( .A(n10342), .ZN(n10695) );
  INV_X1 U12351 ( .A(n9784), .ZN(n9786) );
  OAI222_X1 U12352 ( .A1(P1_U3086), .A2(n10695), .B1(n6535), .B2(n9786), .C1(
        n9785), .C2(n14266), .ZN(P1_U3340) );
  INV_X1 U12353 ( .A(n14753), .ZN(n10737) );
  OAI222_X1 U12354 ( .A1(P2_U3088), .A2(n10737), .B1(n6534), .B2(n9786), .C1(
        n15325), .C2(n11904), .ZN(P2_U3312) );
  INV_X1 U12355 ( .A(n9790), .ZN(n9787) );
  NAND2_X1 U12356 ( .A1(n10398), .A2(n10392), .ZN(n9797) );
  INV_X1 U12357 ( .A(n9789), .ZN(n10084) );
  NAND3_X1 U12358 ( .A1(n10084), .A2(n10085), .A3(n9790), .ZN(n10395) );
  OR2_X1 U12359 ( .A1(n9792), .A2(n11852), .ZN(n10393) );
  INV_X1 U12360 ( .A(n10393), .ZN(n9793) );
  NAND2_X1 U12361 ( .A1(n10395), .A2(n9793), .ZN(n9796) );
  NAND4_X1 U12362 ( .A1(n9797), .A2(n9796), .A3(n9795), .A4(n9794), .ZN(n9798)
         );
  NAND2_X1 U12363 ( .A1(n9798), .A2(P3_STATE_REG_SCAN_IN), .ZN(n10021) );
  NAND2_X1 U12364 ( .A1(n10395), .A2(n10399), .ZN(n10019) );
  AND3_X1 U12365 ( .A1(n10021), .A2(n9800), .A3(n10019), .ZN(n10059) );
  OR2_X1 U12366 ( .A1(n10001), .A2(n9801), .ZN(n9802) );
  NAND2_X1 U12367 ( .A1(n15028), .A2(n15048), .ZN(n11688) );
  INV_X1 U12368 ( .A(n15028), .ZN(n12349) );
  INV_X1 U12369 ( .A(n15048), .ZN(n10098) );
  NAND2_X2 U12370 ( .A1(n11685), .A2(n11688), .ZN(n10097) );
  INV_X1 U12371 ( .A(n11852), .ZN(n9804) );
  NAND2_X1 U12372 ( .A1(n9805), .A2(n9804), .ZN(n9808) );
  NAND2_X1 U12373 ( .A1(n6527), .A2(n12489), .ZN(n9806) );
  NAND2_X1 U12374 ( .A1(n9806), .A2(n9817), .ZN(n9807) );
  NAND2_X1 U12375 ( .A1(n11685), .A2(n10061), .ZN(n9809) );
  NAND2_X1 U12376 ( .A1(n9809), .A2(n10531), .ZN(n9810) );
  NAND2_X1 U12377 ( .A1(n15040), .A2(n10061), .ZN(n15035) );
  AND2_X1 U12378 ( .A1(n9810), .A2(n15035), .ZN(n9811) );
  INV_X1 U12379 ( .A(n9967), .ZN(n9816) );
  NAND2_X1 U12380 ( .A1(n10097), .A2(n10094), .ZN(n15036) );
  OAI22_X1 U12381 ( .A1(n9812), .A2(n15035), .B1(n10525), .B2(n15036), .ZN(
        n9815) );
  OR2_X1 U12382 ( .A1(n10395), .A2(n10393), .ZN(n9813) );
  OAI21_X1 U12383 ( .B1(n10091), .B2(n10398), .A(n9813), .ZN(n9814) );
  OAI21_X1 U12384 ( .B1(n9816), .B2(n9815), .A(n12318), .ZN(n9824) );
  NAND2_X1 U12385 ( .A1(n9817), .A2(n12489), .ZN(n15050) );
  NAND2_X1 U12386 ( .A1(n15049), .A2(n10396), .ZN(n9818) );
  INV_X1 U12387 ( .A(n15039), .ZN(n10102) );
  NOR2_X1 U12388 ( .A1(n10089), .A2(n11853), .ZN(n9821) );
  NAND2_X1 U12389 ( .A1(n15038), .A2(n9821), .ZN(n9819) );
  NAND2_X1 U12390 ( .A1(n15041), .A2(n9821), .ZN(n11862) );
  OAI22_X1 U12391 ( .A1(n10102), .A2(n12336), .B1(n15392), .B2(n6723), .ZN(
        n9822) );
  AOI21_X1 U12392 ( .B1(n12338), .B2(n15048), .A(n9822), .ZN(n9823) );
  OAI211_X1 U12393 ( .C1(n10059), .C2(n9982), .A(n9824), .B(n9823), .ZN(
        P3_U3162) );
  INV_X1 U12394 ( .A(n9825), .ZN(n9828) );
  INV_X1 U12395 ( .A(n9826), .ZN(n9827) );
  NAND2_X1 U12396 ( .A1(n9828), .A2(n9827), .ZN(n9829) );
  XNOR2_X1 U12397 ( .A(n14788), .B(n6528), .ZN(n10066) );
  NAND2_X1 U12398 ( .A1(n13045), .A2(n13326), .ZN(n10064) );
  XNOR2_X1 U12399 ( .A(n10066), .B(n10064), .ZN(n10067) );
  XNOR2_X1 U12400 ( .A(n10067), .B(n10068), .ZN(n9837) );
  NAND2_X1 U12401 ( .A1(n13046), .A2(n14334), .ZN(n9833) );
  NAND2_X1 U12402 ( .A1(n13044), .A2(n14336), .ZN(n9832) );
  NAND2_X1 U12403 ( .A1(n9833), .A2(n9832), .ZN(n10180) );
  NAND2_X1 U12404 ( .A1(n13016), .A2(n10180), .ZN(n9834) );
  NAND2_X1 U12405 ( .A1(P2_U3088), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n13089) );
  OAI211_X1 U12406 ( .C1(n14348), .C2(n10186), .A(n9834), .B(n13089), .ZN(
        n9835) );
  AOI21_X1 U12407 ( .B1(n14788), .B2(n13019), .A(n9835), .ZN(n9836) );
  OAI21_X1 U12408 ( .B1(n9837), .B2(n14342), .A(n9836), .ZN(P2_U3185) );
  OAI22_X1 U12409 ( .A1(n9854), .A2(n13549), .B1(n13770), .B2(n13548), .ZN(
        n9841) );
  OAI22_X1 U12410 ( .A1(n9854), .A2(n9939), .B1(n13770), .B2(n13549), .ZN(
        n9840) );
  XNOR2_X1 U12411 ( .A(n9840), .B(n13591), .ZN(n9927) );
  NAND2_X1 U12412 ( .A1(n9924), .A2(n9927), .ZN(n9842) );
  OAI22_X1 U12413 ( .A1(n14615), .A2(n9939), .B1(n9866), .B2(n13549), .ZN(
        n9843) );
  XNOR2_X1 U12414 ( .A(n9843), .B(n13591), .ZN(n9937) );
  OR2_X1 U12415 ( .A1(n14615), .A2(n13549), .ZN(n9845) );
  NAND2_X1 U12416 ( .A1(n13769), .A2(n13636), .ZN(n9844) );
  AND2_X1 U12417 ( .A1(n9845), .A2(n9844), .ZN(n9936) );
  XNOR2_X1 U12418 ( .A(n9937), .B(n9936), .ZN(n9846) );
  XNOR2_X1 U12419 ( .A(n9938), .B(n9846), .ZN(n9851) );
  INV_X1 U12420 ( .A(n13768), .ZN(n10314) );
  OAI22_X1 U12421 ( .A1(n13770), .A2(n14561), .B1(n10314), .B2(n14581), .ZN(
        n14527) );
  AOI21_X1 U12422 ( .B1(n14527), .B2(n14397), .A(n9847), .ZN(n9848) );
  OAI21_X1 U12423 ( .B1(n14528), .B2(n14401), .A(n9848), .ZN(n9849) );
  AOI21_X1 U12424 ( .B1(n14530), .B2(n14398), .A(n9849), .ZN(n9850) );
  OAI21_X1 U12425 ( .B1(n9851), .B2(n13756), .A(n9850), .ZN(P1_U3227) );
  NAND2_X1 U12426 ( .A1(n9853), .A2(n9852), .ZN(n9856) );
  NAND2_X1 U12427 ( .A1(n9854), .A2(n13770), .ZN(n9855) );
  NAND2_X1 U12428 ( .A1(n9856), .A2(n9855), .ZN(n14523) );
  INV_X1 U12429 ( .A(n9857), .ZN(n14524) );
  NAND2_X1 U12430 ( .A1(n14523), .A2(n14524), .ZN(n9859) );
  NAND2_X1 U12431 ( .A1(n14615), .A2(n9866), .ZN(n9858) );
  NAND2_X1 U12432 ( .A1(n9859), .A2(n9858), .ZN(n10307) );
  XNOR2_X1 U12433 ( .A(n10307), .B(n10305), .ZN(n9923) );
  NAND2_X1 U12434 ( .A1(n9861), .A2(n9860), .ZN(n9863) );
  OAI21_X1 U12435 ( .B1(n9864), .B2(n10305), .A(n10317), .ZN(n9868) );
  NAND2_X1 U12436 ( .A1(n13767), .A2(n14108), .ZN(n9865) );
  OAI21_X1 U12437 ( .B1(n9866), .B2(n14561), .A(n9865), .ZN(n9867) );
  AOI21_X1 U12438 ( .B1(n9868), .B2(n14497), .A(n9867), .ZN(n9917) );
  AOI21_X1 U12439 ( .B1(n10315), .B2(n14531), .A(n14519), .ZN(n9920) );
  AOI22_X1 U12440 ( .A1(n9920), .A2(n14546), .B1(n10315), .B2(n14607), .ZN(
        n9869) );
  OAI211_X1 U12441 ( .C1(n14611), .C2(n9923), .A(n9917), .B(n9869), .ZN(n9872)
         );
  NAND2_X1 U12442 ( .A1(n9872), .A2(n14658), .ZN(n9870) );
  OAI21_X1 U12443 ( .B1(n14658), .B2(n9871), .A(n9870), .ZN(P1_U3534) );
  INV_X1 U12444 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n9874) );
  NAND2_X1 U12445 ( .A1(n9872), .A2(n14645), .ZN(n9873) );
  OAI21_X1 U12446 ( .B1(n14645), .B2(n9874), .A(n9873), .ZN(P1_U3477) );
  INV_X1 U12447 ( .A(n9877), .ZN(n9875) );
  OR2_X1 U12448 ( .A1(n11815), .A2(n9875), .ZN(n9876) );
  AND2_X1 U12449 ( .A1(n9876), .A2(n9726), .ZN(n9881) );
  NOR2_X1 U12450 ( .A1(n9877), .A2(P3_U3151), .ZN(n11859) );
  INV_X1 U12451 ( .A(n11859), .ZN(n11864) );
  NAND2_X1 U12452 ( .A1(n10089), .A2(n11864), .ZN(n9879) );
  NAND2_X1 U12453 ( .A1(n9881), .A2(n9879), .ZN(n9887) );
  INV_X1 U12454 ( .A(n14977), .ZN(n12477) );
  AND2_X1 U12455 ( .A1(n12242), .A2(P3_U3897), .ZN(n14961) );
  NOR3_X1 U12456 ( .A1(n12477), .A2(n14973), .A3(n14961), .ZN(n9891) );
  MUX2_X1 U12457 ( .A(P3_REG2_REG_0__SCAN_IN), .B(P3_REG1_REG_0__SCAN_IN), .S(
        n12463), .Z(n9886) );
  NOR2_X1 U12458 ( .A1(n9886), .A2(n9883), .ZN(n9984) );
  INV_X1 U12459 ( .A(n9984), .ZN(n9988) );
  INV_X1 U12460 ( .A(n9879), .ZN(n9880) );
  INV_X1 U12461 ( .A(P3_REG3_REG_0__SCAN_IN), .ZN(n15296) );
  OAI22_X1 U12462 ( .A1(n14834), .A2(n9882), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n15296), .ZN(n9885) );
  NAND2_X1 U12463 ( .A1(P3_REG1_REG_0__SCAN_IN), .A2(n9883), .ZN(n9979) );
  INV_X1 U12464 ( .A(n9979), .ZN(n10037) );
  AND2_X1 U12465 ( .A1(n14973), .A2(n10037), .ZN(n9884) );
  AOI211_X1 U12466 ( .C1(n9989), .C2(n12477), .A(n9885), .B(n9884), .ZN(n9890)
         );
  NAND2_X1 U12467 ( .A1(n14961), .A2(n9886), .ZN(n9888) );
  MUX2_X1 U12468 ( .A(n12350), .B(n9887), .S(n12242), .Z(n14966) );
  OAI211_X1 U12469 ( .C1(n9891), .C2(n9988), .A(n9890), .B(n9889), .ZN(
        P3_U3182) );
  INV_X1 U12470 ( .A(n14556), .ZN(n9894) );
  NAND2_X1 U12471 ( .A1(n14543), .A2(n14108), .ZN(n14570) );
  OR2_X1 U12472 ( .A1(n13959), .A2(n14572), .ZN(n14080) );
  INV_X1 U12473 ( .A(n14080), .ZN(n14099) );
  OAI21_X1 U12474 ( .B1(n14099), .B2(n14566), .A(n14553), .ZN(n9893) );
  AOI22_X1 U12475 ( .A1(n6531), .A2(P1_REG2_REG_0__SCAN_IN), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(n14567), .ZN(n9892) );
  OAI211_X1 U12476 ( .C1(n9894), .C2(n14570), .A(n9893), .B(n9892), .ZN(n9897)
         );
  NAND2_X1 U12477 ( .A1(n14543), .A2(n14497), .ZN(n14085) );
  AOI21_X1 U12478 ( .B1(n14123), .B2(n14085), .A(n9895), .ZN(n9896) );
  OR2_X1 U12479 ( .A1(n9897), .A2(n9896), .ZN(P1_U3293) );
  AOI22_X1 U12480 ( .A1(n10336), .A2(n8554), .B1(P1_REG1_REG_14__SCAN_IN), 
        .B2(n10341), .ZN(n9901) );
  INV_X1 U12481 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n11206) );
  AOI21_X1 U12482 ( .B1(n14415), .B2(n9907), .A(n9898), .ZN(n14458) );
  INV_X1 U12483 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n11040) );
  AOI22_X1 U12484 ( .A1(n14461), .A2(n11040), .B1(P1_REG1_REG_12__SCAN_IN), 
        .B2(n9905), .ZN(n14457) );
  NOR2_X1 U12485 ( .A1(n14461), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n9899) );
  NOR2_X1 U12486 ( .A1(n14456), .A2(n9899), .ZN(n14485) );
  MUX2_X1 U12487 ( .A(n11206), .B(P1_REG1_REG_13__SCAN_IN), .S(n14471), .Z(
        n14484) );
  NAND2_X1 U12488 ( .A1(n14485), .A2(n14484), .ZN(n14482) );
  OAI21_X1 U12489 ( .B1(n11206), .B2(n14471), .A(n14482), .ZN(n9900) );
  AOI21_X1 U12490 ( .B1(n9901), .B2(n9900), .A(n10340), .ZN(n9913) );
  NAND2_X1 U12491 ( .A1(n14472), .A2(P1_ADDR_REG_14__SCAN_IN), .ZN(n9902) );
  NAND2_X1 U12492 ( .A1(P1_REG3_REG_14__SCAN_IN), .A2(P1_U3086), .ZN(n14399)
         );
  NAND2_X1 U12493 ( .A1(n9902), .A2(n14399), .ZN(n9903) );
  AOI21_X1 U12494 ( .B1(n10336), .B2(n14476), .A(n9903), .ZN(n9912) );
  MUX2_X1 U12495 ( .A(n11214), .B(P1_REG2_REG_14__SCAN_IN), .S(n10336), .Z(
        n9904) );
  INV_X1 U12496 ( .A(n9904), .ZN(n9910) );
  INV_X1 U12497 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n11157) );
  MUX2_X1 U12498 ( .A(n11157), .B(P1_REG2_REG_13__SCAN_IN), .S(n14471), .Z(
        n14480) );
  AOI22_X1 U12499 ( .A1(n14461), .A2(n10865), .B1(P1_REG2_REG_12__SCAN_IN), 
        .B2(n9905), .ZN(n14455) );
  OAI21_X1 U12500 ( .B1(n9907), .B2(n10817), .A(n9906), .ZN(n14454) );
  NOR2_X1 U12501 ( .A1(n14455), .A2(n14454), .ZN(n14453) );
  NOR2_X1 U12502 ( .A1(n14461), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n9908) );
  NOR2_X1 U12503 ( .A1(n14453), .A2(n9908), .ZN(n14481) );
  NAND2_X1 U12504 ( .A1(n14480), .A2(n14481), .ZN(n14479) );
  OAI21_X1 U12505 ( .B1(n14471), .B2(n11157), .A(n14479), .ZN(n9909) );
  NAND2_X1 U12506 ( .A1(n9910), .A2(n9909), .ZN(n10337) );
  OAI211_X1 U12507 ( .C1(n9910), .C2(n9909), .A(n14478), .B(n10337), .ZN(n9911) );
  OAI211_X1 U12508 ( .C1(n9913), .C2(n14459), .A(n9912), .B(n9911), .ZN(
        P1_U3257) );
  INV_X1 U12509 ( .A(n10743), .ZN(n11363) );
  INV_X1 U12510 ( .A(n9914), .ZN(n9916) );
  OAI222_X1 U12511 ( .A1(P2_U3088), .A2(n11363), .B1(n6534), .B2(n9916), .C1(
        n15181), .C2(n11904), .ZN(P2_U3311) );
  INV_X1 U12512 ( .A(n11194), .ZN(n11187) );
  OAI222_X1 U12513 ( .A1(P1_U3086), .A2(n11187), .B1(n6535), .B2(n9916), .C1(
        n9915), .C2(n14266), .ZN(P1_U3339) );
  MUX2_X1 U12514 ( .A(n9918), .B(n9917), .S(n14543), .Z(n9922) );
  OAI22_X1 U12515 ( .A1(n6966), .A2(n14119), .B1(n9954), .B2(n14542), .ZN(
        n9919) );
  AOI21_X1 U12516 ( .B1(n9920), .B2(n14099), .A(n9919), .ZN(n9921) );
  OAI211_X1 U12517 ( .C1(n9923), .C2(n14123), .A(n9922), .B(n9921), .ZN(
        P1_U3287) );
  NAND2_X1 U12518 ( .A1(n9925), .A2(n9924), .ZN(n9926) );
  XOR2_X1 U12519 ( .A(n9927), .B(n9926), .Z(n9934) );
  NAND2_X1 U12520 ( .A1(n14608), .A2(n14398), .ZN(n9931) );
  AOI21_X1 U12521 ( .B1(n9929), .B2(n14397), .A(n9928), .ZN(n9930) );
  OAI211_X1 U12522 ( .C1(n14401), .C2(n9932), .A(n9931), .B(n9930), .ZN(n9933)
         );
  AOI21_X1 U12523 ( .B1(n9934), .B2(n14395), .A(n9933), .ZN(n9935) );
  INV_X1 U12524 ( .A(n9935), .ZN(P1_U3230) );
  NAND2_X1 U12525 ( .A1(n10315), .A2(n13640), .ZN(n9941) );
  NAND2_X1 U12526 ( .A1(n13768), .A2(n6536), .ZN(n9940) );
  NAND2_X1 U12527 ( .A1(n9941), .A2(n9940), .ZN(n9942) );
  XNOR2_X1 U12528 ( .A(n9942), .B(n13637), .ZN(n9948) );
  INV_X1 U12529 ( .A(n9948), .ZN(n9946) );
  NAND2_X1 U12530 ( .A1(n10315), .A2(n6536), .ZN(n9944) );
  NAND2_X1 U12531 ( .A1(n13768), .A2(n13636), .ZN(n9943) );
  NAND2_X1 U12532 ( .A1(n9944), .A2(n9943), .ZN(n9947) );
  INV_X1 U12533 ( .A(n9947), .ZN(n9945) );
  NAND2_X1 U12534 ( .A1(n9946), .A2(n9945), .ZN(n10287) );
  INV_X1 U12535 ( .A(n10287), .ZN(n9949) );
  AND2_X1 U12536 ( .A1(n9948), .A2(n9947), .ZN(n10285) );
  NOR2_X1 U12537 ( .A1(n9949), .A2(n10285), .ZN(n9950) );
  XNOR2_X1 U12538 ( .A(n10286), .B(n9950), .ZN(n9957) );
  INV_X1 U12539 ( .A(n13767), .ZN(n10311) );
  OAI21_X1 U12540 ( .B1(n13748), .B2(n10311), .A(n9951), .ZN(n9952) );
  AOI21_X1 U12541 ( .B1(n13750), .B2(n13769), .A(n9952), .ZN(n9953) );
  OAI21_X1 U12542 ( .B1(n9954), .B2(n14401), .A(n9953), .ZN(n9955) );
  AOI21_X1 U12543 ( .B1(n10315), .B2(n14398), .A(n9955), .ZN(n9956) );
  OAI21_X1 U12544 ( .B1(n9957), .B2(n13756), .A(n9956), .ZN(P1_U3239) );
  INV_X1 U12545 ( .A(n11195), .ZN(n13821) );
  INV_X1 U12546 ( .A(n9958), .ZN(n9960) );
  OAI222_X1 U12547 ( .A1(P1_U3086), .A2(n13821), .B1(n6535), .B2(n9960), .C1(
        n9959), .C2(n14266), .ZN(P1_U3338) );
  OAI222_X1 U12548 ( .A1(n11904), .A2(n9961), .B1(n6534), .B2(n9960), .C1(
        n13124), .C2(P2_U3088), .ZN(P2_U3310) );
  OR2_X1 U12549 ( .A1(n10001), .A2(n9962), .ZN(n9964) );
  OR2_X1 U12550 ( .A1(n10193), .A2(SI_2_), .ZN(n9963) );
  OAI211_X1 U12551 ( .C1(n10046), .C2(n9726), .A(n9964), .B(n9963), .ZN(n15019) );
  INV_X1 U12552 ( .A(n15019), .ZN(n10096) );
  XNOR2_X1 U12553 ( .A(n10531), .B(n10096), .ZN(n10000) );
  XNOR2_X1 U12554 ( .A(n10000), .B(n15039), .ZN(n9969) );
  XNOR2_X1 U12555 ( .A(n15048), .B(n10531), .ZN(n9965) );
  NAND2_X1 U12556 ( .A1(n9965), .A2(n15028), .ZN(n9966) );
  NAND2_X1 U12557 ( .A1(n9967), .A2(n9966), .ZN(n9968) );
  OAI21_X1 U12558 ( .B1(n9969), .B2(n9968), .A(n10006), .ZN(n9970) );
  NAND2_X1 U12559 ( .A1(n9970), .A2(n12318), .ZN(n9977) );
  INV_X1 U12560 ( .A(P3_REG1_REG_3__SCAN_IN), .ZN(n10914) );
  OR2_X1 U12561 ( .A1(n11436), .A2(n10914), .ZN(n9973) );
  INV_X1 U12562 ( .A(P3_REG2_REG_3__SCAN_IN), .ZN(n10915) );
  OR2_X1 U12563 ( .A1(n10012), .A2(P3_REG3_REG_3__SCAN_IN), .ZN(n9971) );
  OAI22_X1 U12564 ( .A1(n15028), .A2(n15392), .B1(n12336), .B2(n15030), .ZN(
        n9975) );
  AOI21_X1 U12565 ( .B1(n10096), .B2(n12338), .A(n9975), .ZN(n9976) );
  OAI211_X1 U12566 ( .C1(n10059), .C2(n15021), .A(n9977), .B(n9976), .ZN(
        P3_U3177) );
  INV_X1 U12567 ( .A(n9999), .ZN(n9980) );
  NOR2_X1 U12568 ( .A1(P3_IR_REG_1__SCAN_IN), .A2(n9979), .ZN(n9978) );
  AOI21_X1 U12569 ( .B1(n9980), .B2(n9979), .A(n9978), .ZN(n9981) );
  NAND2_X1 U12570 ( .A1(n9981), .A2(P3_REG1_REG_1__SCAN_IN), .ZN(n10035) );
  OAI21_X1 U12571 ( .B1(P3_REG1_REG_1__SCAN_IN), .B2(n9981), .A(n10035), .ZN(
        n9997) );
  OAI22_X1 U12572 ( .A1(n14834), .A2(n6760), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n9982), .ZN(n9996) );
  MUX2_X1 U12573 ( .A(P3_REG2_REG_1__SCAN_IN), .B(P3_REG1_REG_1__SCAN_IN), .S(
        n12463), .Z(n9983) );
  NOR2_X1 U12574 ( .A1(n9983), .A2(n9999), .ZN(n10043) );
  AOI21_X1 U12575 ( .B1(n9983), .B2(n9999), .A(n10043), .ZN(n9985) );
  INV_X1 U12576 ( .A(n9985), .ZN(n9987) );
  NAND2_X1 U12577 ( .A1(n9985), .A2(n9984), .ZN(n10052) );
  INV_X1 U12578 ( .A(n10052), .ZN(n9986) );
  AOI21_X1 U12579 ( .B1(n9988), .B2(n9987), .A(n9986), .ZN(n9994) );
  OR2_X1 U12580 ( .A1(n9999), .A2(n9989), .ZN(n9991) );
  INV_X1 U12581 ( .A(n10031), .ZN(n9990) );
  NAND2_X1 U12582 ( .A1(n9991), .A2(n9990), .ZN(n9992) );
  NOR2_X1 U12583 ( .A1(n9992), .A2(n9739), .ZN(n10032) );
  AOI21_X1 U12584 ( .B1(n9739), .B2(n9992), .A(n10032), .ZN(n9993) );
  OAI22_X1 U12585 ( .A1(n9994), .A2(n14838), .B1(n9993), .B2(n14977), .ZN(
        n9995) );
  AOI211_X1 U12586 ( .C1(n14973), .C2(n9997), .A(n9996), .B(n9995), .ZN(n9998)
         );
  OAI21_X1 U12587 ( .B1(n9999), .B2(n14966), .A(n9998), .ZN(P3_U3183) );
  NAND2_X1 U12588 ( .A1(n10000), .A2(n10102), .ZN(n10007) );
  OR2_X1 U12589 ( .A1(n10193), .A2(SI_3_), .ZN(n10005) );
  OR2_X1 U12590 ( .A1(n10001), .A2(n10002), .ZN(n10004) );
  NAND2_X1 U12591 ( .A1(n11492), .A2(n10917), .ZN(n10003) );
  AOI21_X1 U12592 ( .B1(n10006), .B2(n10007), .A(n10008), .ZN(n10026) );
  AND2_X1 U12593 ( .A1(n10008), .A2(n10007), .ZN(n10009) );
  NAND2_X1 U12594 ( .A1(n10010), .A2(n10009), .ZN(n10204) );
  NAND2_X1 U12595 ( .A1(n10204), .A2(n12318), .ZN(n10025) );
  INV_X1 U12596 ( .A(n12327), .ZN(n15399) );
  NAND2_X1 U12597 ( .A1(n11567), .A2(P3_REG2_REG_4__SCAN_IN), .ZN(n10017) );
  INV_X1 U12598 ( .A(P3_REG0_REG_4__SCAN_IN), .ZN(n10011) );
  OR2_X1 U12599 ( .A1(n11438), .A2(n10011), .ZN(n10016) );
  AND2_X1 U12600 ( .A1(P3_REG3_REG_3__SCAN_IN), .A2(P3_REG3_REG_4__SCAN_IN), 
        .ZN(n10013) );
  NOR2_X1 U12601 ( .A1(n10209), .A2(n10013), .ZN(n10634) );
  OR2_X1 U12602 ( .A1(n10012), .A2(n10634), .ZN(n10015) );
  INV_X1 U12603 ( .A(P3_REG1_REG_4__SCAN_IN), .ZN(n10920) );
  OR2_X1 U12604 ( .A1(n11570), .A2(n10920), .ZN(n10014) );
  NAND2_X1 U12605 ( .A1(n12332), .A2(n15039), .ZN(n10018) );
  INV_X1 U12606 ( .A(P3_REG3_REG_3__SCAN_IN), .ZN(n10111) );
  OR2_X1 U12607 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n10111), .ZN(n14833) );
  OAI211_X1 U12608 ( .C1(n10709), .C2(n12336), .A(n10018), .B(n14833), .ZN(
        n10023) );
  AND2_X1 U12609 ( .A1(n10019), .A2(n11864), .ZN(n10020) );
  NOR2_X1 U12610 ( .A1(n15395), .A2(P3_REG3_REG_3__SCAN_IN), .ZN(n10022) );
  AOI211_X1 U12611 ( .C1(n15399), .C2(n10369), .A(n10023), .B(n10022), .ZN(
        n10024) );
  OAI21_X1 U12612 ( .B1(n10026), .B2(n10025), .A(n10024), .ZN(P3_U3158) );
  NAND2_X1 U12613 ( .A1(n10668), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n10118) );
  NAND2_X1 U12614 ( .A1(n11911), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n10029) );
  NAND2_X1 U12615 ( .A1(n10118), .A2(n10029), .ZN(n10115) );
  XNOR2_X1 U12616 ( .A(n10117), .B(n10115), .ZN(n11510) );
  INV_X1 U12617 ( .A(n11510), .ZN(n10030) );
  INV_X1 U12618 ( .A(SI_21_), .ZN(n11511) );
  OAI222_X1 U12619 ( .A1(n6527), .A2(P3_U3151), .B1(n12245), .B2(n10030), .C1(
        n11511), .C2(n11338), .ZN(P3_U3274) );
  INV_X1 U12620 ( .A(n10046), .ZN(n10899) );
  MUX2_X1 U12621 ( .A(n10045), .B(P3_REG2_REG_2__SCAN_IN), .S(n10046), .Z(
        n10034) );
  OR2_X1 U12622 ( .A1(n10032), .A2(n10031), .ZN(n10033) );
  NAND2_X1 U12623 ( .A1(n10034), .A2(n10033), .ZN(n10889) );
  OAI21_X1 U12624 ( .B1(n10034), .B2(n10033), .A(n10889), .ZN(n10057) );
  MUX2_X1 U12625 ( .A(P3_REG1_REG_2__SCAN_IN), .B(n10044), .S(n10046), .Z(
        n10040) );
  INV_X1 U12626 ( .A(n10035), .ZN(n10036) );
  AOI21_X1 U12627 ( .B1(n10038), .B2(n10037), .A(n10036), .ZN(n10039) );
  NOR2_X1 U12628 ( .A1(n10039), .A2(n10040), .ZN(n10898) );
  AOI21_X1 U12629 ( .B1(n10040), .B2(n10039), .A(n10898), .ZN(n10042) );
  AOI22_X1 U12630 ( .A1(n14969), .A2(P3_ADDR_REG_2__SCAN_IN), .B1(
        P3_REG3_REG_2__SCAN_IN), .B2(P3_U3151), .ZN(n10041) );
  OAI21_X1 U12631 ( .B1(n10042), .B2(n12498), .A(n10041), .ZN(n10056) );
  INV_X1 U12632 ( .A(n10043), .ZN(n10051) );
  MUX2_X1 U12633 ( .A(n10045), .B(n10044), .S(n12463), .Z(n10047) );
  NAND2_X1 U12634 ( .A1(n10047), .A2(n10046), .ZN(n10913) );
  INV_X1 U12635 ( .A(n10047), .ZN(n10048) );
  NAND2_X1 U12636 ( .A1(n10048), .A2(n10899), .ZN(n10049) );
  NAND2_X1 U12637 ( .A1(n10913), .A2(n10049), .ZN(n10050) );
  AOI21_X1 U12638 ( .B1(n10052), .B2(n10051), .A(n10050), .ZN(n14837) );
  INV_X1 U12639 ( .A(n14837), .ZN(n10054) );
  NAND3_X1 U12640 ( .A1(n10052), .A2(n10051), .A3(n10050), .ZN(n10053) );
  AOI21_X1 U12641 ( .B1(n10054), .B2(n10053), .A(n14838), .ZN(n10055) );
  AOI211_X1 U12642 ( .C1(n12477), .C2(n10057), .A(n10056), .B(n10055), .ZN(
        n10058) );
  OAI21_X1 U12643 ( .B1(n10899), .B2(n14966), .A(n10058), .ZN(P3_U3184) );
  INV_X1 U12644 ( .A(n10059), .ZN(n10060) );
  NAND2_X1 U12645 ( .A1(n10060), .A2(P3_REG3_REG_0__SCAN_IN), .ZN(n10063) );
  AOI22_X1 U12646 ( .A1(n15389), .A2(n12349), .B1(n15399), .B2(n10061), .ZN(
        n10062) );
  OAI211_X1 U12647 ( .C1(n11829), .C2(n15401), .A(n10063), .B(n10062), .ZN(
        P3_U3172) );
  INV_X1 U12648 ( .A(n14795), .ZN(n10082) );
  INV_X1 U12649 ( .A(n10064), .ZN(n10065) );
  XNOR2_X1 U12650 ( .A(n14795), .B(n6540), .ZN(n10069) );
  NAND2_X1 U12651 ( .A1(n13044), .A2(n13326), .ZN(n10070) );
  NAND2_X1 U12652 ( .A1(n10069), .A2(n10070), .ZN(n10241) );
  INV_X1 U12653 ( .A(n10069), .ZN(n10072) );
  INV_X1 U12654 ( .A(n10070), .ZN(n10071) );
  NAND2_X1 U12655 ( .A1(n10072), .A2(n10071), .ZN(n10073) );
  AND2_X1 U12656 ( .A1(n10241), .A2(n10073), .ZN(n10074) );
  OAI21_X1 U12657 ( .B1(n10075), .B2(n10074), .A(n10242), .ZN(n10076) );
  NAND2_X1 U12658 ( .A1(n10076), .A2(n12973), .ZN(n10081) );
  NAND2_X1 U12659 ( .A1(n13042), .A2(n14336), .ZN(n10078) );
  NAND2_X1 U12660 ( .A1(n13045), .A2(n14334), .ZN(n10077) );
  NAND2_X1 U12661 ( .A1(n10078), .A2(n10077), .ZN(n10465) );
  AND2_X1 U12662 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(P2_U3088), .ZN(n13105) );
  NOR2_X1 U12663 ( .A1(n14348), .A2(n10473), .ZN(n10079) );
  AOI211_X1 U12664 ( .C1(n13016), .C2(n10465), .A(n13105), .B(n10079), .ZN(
        n10080) );
  OAI211_X1 U12665 ( .C1(n10082), .C2(n14340), .A(n10081), .B(n10080), .ZN(
        P2_U3193) );
  OAI22_X1 U12666 ( .A1(n10086), .A2(n10085), .B1(n10084), .B2(n10083), .ZN(
        n10087) );
  NAND2_X1 U12667 ( .A1(n10088), .A2(n10087), .ZN(n10109) );
  OR2_X1 U12668 ( .A1(n15018), .A2(n15050), .ZN(n10090) );
  OR2_X1 U12669 ( .A1(n10091), .A2(n11853), .ZN(n10093) );
  NAND2_X1 U12670 ( .A1(n10093), .A2(n10092), .ZN(n10408) );
  NOR2_X1 U12671 ( .A1(n6527), .A2(n15050), .ZN(n15051) );
  NOR2_X1 U12672 ( .A1(n10408), .A2(n15051), .ZN(n15010) );
  INV_X1 U12673 ( .A(n10097), .ZN(n11828) );
  NAND2_X1 U12674 ( .A1(n11828), .A2(n10095), .ZN(n15037) );
  NAND2_X1 U12675 ( .A1(n15037), .A2(n11688), .ZN(n15017) );
  XNOR2_X1 U12676 ( .A(n15039), .B(n15019), .ZN(n10101) );
  INV_X1 U12677 ( .A(n10101), .ZN(n15025) );
  NAND2_X1 U12678 ( .A1(n10102), .A2(n10096), .ZN(n11698) );
  NAND2_X1 U12679 ( .A1(n11683), .A2(n11698), .ZN(n10403) );
  NAND2_X1 U12680 ( .A1(n15030), .A2(n10369), .ZN(n11699) );
  INV_X1 U12681 ( .A(n10369), .ZN(n10110) );
  NAND2_X1 U12682 ( .A1(n12348), .A2(n10110), .ZN(n11696) );
  XNOR2_X1 U12683 ( .A(n10403), .B(n11825), .ZN(n15069) );
  INV_X1 U12684 ( .A(n15069), .ZN(n10114) );
  NAND2_X1 U12685 ( .A1(n15035), .A2(n10097), .ZN(n10100) );
  NAND2_X1 U12686 ( .A1(n15028), .A2(n10098), .ZN(n10099) );
  NAND2_X1 U12687 ( .A1(n10100), .A2(n10099), .ZN(n15024) );
  NAND2_X1 U12688 ( .A1(n15024), .A2(n10101), .ZN(n10104) );
  NAND2_X1 U12689 ( .A1(n10102), .A2(n15019), .ZN(n10103) );
  INV_X1 U12690 ( .A(n11825), .ZN(n10105) );
  NAND2_X1 U12691 ( .A1(n7445), .A2(n10105), .ZN(n10371) );
  OAI211_X1 U12692 ( .C1(n7445), .C2(n10105), .A(n15046), .B(n10371), .ZN(
        n10107) );
  AOI22_X1 U12693 ( .A1(n12347), .A2(n15038), .B1(n15041), .B2(n15039), .ZN(
        n10106) );
  NAND2_X1 U12694 ( .A1(n10107), .A2(n10106), .ZN(n15067) );
  INV_X1 U12695 ( .A(n15067), .ZN(n10108) );
  INV_X2 U12696 ( .A(n15052), .ZN(n15057) );
  MUX2_X1 U12697 ( .A(n10915), .B(n10108), .S(n15057), .Z(n10113) );
  INV_X1 U12698 ( .A(n15050), .ZN(n15022) );
  INV_X1 U12699 ( .A(n12535), .ZN(n14991) );
  NOR2_X1 U12700 ( .A1(n10110), .A2(n15018), .ZN(n15068) );
  AOI22_X1 U12701 ( .A1(n14991), .A2(n15068), .B1(n15055), .B2(n10111), .ZN(
        n10112) );
  OAI211_X1 U12702 ( .C1(n12725), .C2(n10114), .A(n10113), .B(n10112), .ZN(
        P3_U3230) );
  INV_X1 U12703 ( .A(n10115), .ZN(n10116) );
  INV_X1 U12704 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n10119) );
  NAND2_X1 U12705 ( .A1(n10119), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n10282) );
  NAND2_X1 U12706 ( .A1(n10880), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n10120) );
  NAND2_X1 U12707 ( .A1(n10282), .A2(n10120), .ZN(n10279) );
  XNOR2_X1 U12708 ( .A(n10281), .B(n10279), .ZN(n11515) );
  INV_X1 U12709 ( .A(SI_22_), .ZN(n10121) );
  AOI22_X1 U12710 ( .A1(n11860), .A2(P3_STATE_REG_SCAN_IN), .B1(n10122), .B2(
        n10121), .ZN(n10123) );
  OAI21_X1 U12711 ( .B1(n11515), .B2(n12245), .A(n10123), .ZN(n10124) );
  INV_X1 U12712 ( .A(n10124), .ZN(P3_U3273) );
  INV_X1 U12713 ( .A(n10125), .ZN(n10135) );
  INV_X1 U12714 ( .A(n10126), .ZN(n10127) );
  MUX2_X1 U12715 ( .A(n10128), .B(n10127), .S(n13281), .Z(n10134) );
  OAI22_X1 U12716 ( .A1(n13311), .A2(n10130), .B1(n10129), .B2(n13323), .ZN(
        n10131) );
  AOI21_X1 U12717 ( .B1(n10132), .B2(n14362), .A(n10131), .ZN(n10133) );
  OAI211_X1 U12718 ( .C1(n13342), .C2(n10135), .A(n10134), .B(n10133), .ZN(
        P2_U3261) );
  XNOR2_X1 U12719 ( .A(n10136), .B(n10138), .ZN(n10144) );
  INV_X1 U12720 ( .A(n10144), .ZN(n14785) );
  NOR2_X1 U12721 ( .A1(n13144), .A2(n11924), .ZN(n10137) );
  NAND2_X1 U12722 ( .A1(n13281), .A2(n10137), .ZN(n10421) );
  NAND2_X1 U12723 ( .A1(n10139), .A2(n10138), .ZN(n10140) );
  AOI21_X1 U12724 ( .B1(n10141), .B2(n10140), .A(n14351), .ZN(n10142) );
  AOI211_X1 U12725 ( .C1(n13307), .C2(n10144), .A(n10143), .B(n10142), .ZN(
        n14784) );
  MUX2_X1 U12726 ( .A(n10145), .B(n14784), .S(n13281), .Z(n10150) );
  AOI211_X1 U12727 ( .C1(n14782), .C2(n10172), .A(n9445), .B(n10183), .ZN(
        n14781) );
  INV_X1 U12728 ( .A(n14782), .ZN(n10147) );
  OAI22_X1 U12729 ( .A1(n10147), .A2(n13311), .B1(n13323), .B2(n10146), .ZN(
        n10148) );
  AOI21_X1 U12730 ( .B1(n14781), .B2(n14362), .A(n10148), .ZN(n10149) );
  OAI211_X1 U12731 ( .C1(n14785), .C2(n10421), .A(n10150), .B(n10149), .ZN(
        P2_U3259) );
  INV_X1 U12732 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n14386) );
  NAND2_X1 U12733 ( .A1(n10157), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n10151) );
  AND2_X1 U12734 ( .A1(n10152), .A2(n10151), .ZN(n14720) );
  MUX2_X1 U12735 ( .A(n14386), .B(P2_REG1_REG_12__SCAN_IN), .S(n14732), .Z(
        n14719) );
  AOI21_X1 U12736 ( .B1(n14386), .B2(n14732), .A(n14722), .ZN(n14743) );
  MUX2_X1 U12737 ( .A(P2_REG1_REG_13__SCAN_IN), .B(n10153), .S(n10160), .Z(
        n14742) );
  NAND2_X1 U12738 ( .A1(n14743), .A2(n14742), .ZN(n14741) );
  NAND2_X1 U12739 ( .A1(n10160), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n10155) );
  INV_X1 U12740 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n14372) );
  MUX2_X1 U12741 ( .A(n14372), .B(P2_REG1_REG_14__SCAN_IN), .S(n10163), .Z(
        n10154) );
  AOI21_X1 U12742 ( .B1(n14741), .B2(n10155), .A(n10154), .ZN(n10734) );
  NAND3_X1 U12743 ( .A1(n14741), .A2(n10155), .A3(n10154), .ZN(n10156) );
  NAND2_X1 U12744 ( .A1(n10156), .A2(n14759), .ZN(n10166) );
  NAND2_X1 U12745 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(P2_U3088), .ZN(n14345)
         );
  OR2_X1 U12746 ( .A1(n10157), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n14724) );
  NAND2_X1 U12747 ( .A1(n14726), .A2(n14724), .ZN(n10158) );
  MUX2_X1 U12748 ( .A(n10774), .B(P2_REG2_REG_12__SCAN_IN), .S(n14732), .Z(
        n14723) );
  NAND2_X1 U12749 ( .A1(n10158), .A2(n14723), .ZN(n14728) );
  OAI21_X1 U12750 ( .B1(n10159), .B2(P2_REG2_REG_12__SCAN_IN), .A(n14728), 
        .ZN(n14746) );
  MUX2_X1 U12751 ( .A(n10993), .B(P2_REG2_REG_13__SCAN_IN), .S(n10160), .Z(
        n14747) );
  NOR2_X1 U12752 ( .A1(n14746), .A2(n14747), .ZN(n14744) );
  AOI21_X1 U12753 ( .B1(P2_REG2_REG_13__SCAN_IN), .B2(n10160), .A(n14744), 
        .ZN(n10725) );
  XNOR2_X1 U12754 ( .A(n10725), .B(n10163), .ZN(n10161) );
  NAND2_X1 U12755 ( .A1(n10161), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n10726) );
  OAI211_X1 U12756 ( .C1(n10161), .C2(P2_REG2_REG_14__SCAN_IN), .A(n10726), 
        .B(n14756), .ZN(n10162) );
  AND2_X1 U12757 ( .A1(n14345), .A2(n10162), .ZN(n10165) );
  AOI22_X1 U12758 ( .A1(n14752), .A2(P2_ADDR_REG_14__SCAN_IN), .B1(n14754), 
        .B2(n10163), .ZN(n10164) );
  OAI211_X1 U12759 ( .C1(n10734), .C2(n10166), .A(n10165), .B(n10164), .ZN(
        P2_U3228) );
  XNOR2_X1 U12760 ( .A(n11980), .B(n13047), .ZN(n12196) );
  XNOR2_X1 U12761 ( .A(n10167), .B(n12196), .ZN(n14776) );
  XNOR2_X1 U12762 ( .A(n10168), .B(n12196), .ZN(n10170) );
  AOI21_X1 U12763 ( .B1(n10170), .B2(n13335), .A(n10169), .ZN(n14778) );
  MUX2_X1 U12764 ( .A(n10171), .B(n14778), .S(n13281), .Z(n10177) );
  OAI211_X1 U12765 ( .C1(n6795), .C2(n6706), .A(n9550), .B(n10172), .ZN(n14777) );
  INV_X1 U12766 ( .A(n14777), .ZN(n10175) );
  OAI22_X1 U12767 ( .A1(n6795), .A2(n13311), .B1(n13323), .B2(n10173), .ZN(
        n10174) );
  AOI21_X1 U12768 ( .B1(n10175), .B2(n14362), .A(n10174), .ZN(n10176) );
  OAI211_X1 U12769 ( .C1(n13342), .C2(n14776), .A(n10177), .B(n10176), .ZN(
        P2_U3260) );
  XOR2_X1 U12770 ( .A(n10178), .B(n12200), .Z(n14792) );
  XOR2_X1 U12771 ( .A(n10179), .B(n12200), .Z(n10181) );
  AOI21_X1 U12772 ( .B1(n10181), .B2(n13335), .A(n10180), .ZN(n14790) );
  MUX2_X1 U12773 ( .A(n14790), .B(n10182), .S(n14367), .Z(n10190) );
  INV_X1 U12774 ( .A(n10183), .ZN(n10185) );
  INV_X1 U12775 ( .A(n10471), .ZN(n10184) );
  AOI211_X1 U12776 ( .C1(n14788), .C2(n10185), .A(n9445), .B(n10184), .ZN(
        n14787) );
  OAI22_X1 U12777 ( .A1(n10187), .A2(n13311), .B1(n13323), .B2(n10186), .ZN(
        n10188) );
  AOI21_X1 U12778 ( .B1(n14787), .B2(n14362), .A(n10188), .ZN(n10189) );
  OAI211_X1 U12779 ( .C1(n13342), .C2(n14792), .A(n10190), .B(n10189), .ZN(
        P2_U3258) );
  INV_X1 U12780 ( .A(n10191), .ZN(n10192) );
  NAND2_X1 U12781 ( .A1(n10192), .A2(n12348), .ZN(n10201) );
  NAND2_X1 U12782 ( .A1(n10204), .A2(n10201), .ZN(n10207) );
  OR2_X1 U12783 ( .A1(n11662), .A2(SI_4_), .ZN(n10197) );
  OR2_X1 U12784 ( .A1(n10001), .A2(n10194), .ZN(n10196) );
  NAND2_X1 U12785 ( .A1(n11492), .A2(n14857), .ZN(n10195) );
  XNOR2_X1 U12786 ( .A(n10531), .B(n10633), .ZN(n10198) );
  NAND2_X1 U12787 ( .A1(n10198), .A2(n10709), .ZN(n10262) );
  INV_X1 U12788 ( .A(n10198), .ZN(n10199) );
  NAND2_X1 U12789 ( .A1(n10199), .A2(n12347), .ZN(n10200) );
  NAND2_X1 U12790 ( .A1(n10262), .A2(n10200), .ZN(n10206) );
  INV_X1 U12791 ( .A(n10206), .ZN(n10202) );
  AND2_X1 U12792 ( .A1(n10202), .A2(n10201), .ZN(n10203) );
  NAND2_X1 U12793 ( .A1(n10204), .A2(n10203), .ZN(n10263) );
  INV_X1 U12794 ( .A(n10263), .ZN(n10205) );
  AOI21_X1 U12795 ( .B1(n10207), .B2(n10206), .A(n10205), .ZN(n10221) );
  INV_X1 U12796 ( .A(P3_REG1_REG_5__SCAN_IN), .ZN(n10927) );
  OR2_X1 U12797 ( .A1(n11436), .A2(n10927), .ZN(n10213) );
  OR2_X1 U12798 ( .A1(n10209), .A2(n10208), .ZN(n10210) );
  AND2_X1 U12799 ( .A1(n10267), .A2(n10210), .ZN(n10711) );
  OR2_X1 U12800 ( .A1(n10012), .A2(n10711), .ZN(n10212) );
  INV_X1 U12801 ( .A(P3_REG2_REG_5__SCAN_IN), .ZN(n10928) );
  INV_X1 U12802 ( .A(n10638), .ZN(n12346) );
  NAND2_X1 U12803 ( .A1(n15389), .A2(n12346), .ZN(n10217) );
  INV_X1 U12804 ( .A(P3_REG3_REG_4__SCAN_IN), .ZN(n10215) );
  NOR2_X1 U12805 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n10215), .ZN(n14859) );
  INV_X1 U12806 ( .A(n14859), .ZN(n10216) );
  OAI211_X1 U12807 ( .C1(n15030), .C2(n15392), .A(n10217), .B(n10216), .ZN(
        n10219) );
  NOR2_X1 U12808 ( .A1(n15395), .A2(n10634), .ZN(n10218) );
  AOI211_X1 U12809 ( .C1(n15399), .C2(n10633), .A(n10219), .B(n10218), .ZN(
        n10220) );
  OAI21_X1 U12810 ( .B1(n10221), .B2(n15401), .A(n10220), .ZN(P3_U3170) );
  INV_X1 U12811 ( .A(P3_REG3_REG_25__SCAN_IN), .ZN(n11543) );
  NAND2_X1 U12812 ( .A1(n11544), .A2(n11543), .ZN(n11552) );
  INV_X1 U12813 ( .A(P3_REG3_REG_28__SCAN_IN), .ZN(n11898) );
  NAND2_X1 U12814 ( .A1(n12506), .A2(n11566), .ZN(n10303) );
  INV_X1 U12815 ( .A(P3_REG1_REG_29__SCAN_IN), .ZN(n11625) );
  NAND2_X1 U12816 ( .A1(n11567), .A2(P3_REG2_REG_29__SCAN_IN), .ZN(n10223) );
  OAI211_X1 U12817 ( .C1(n11625), .C2(n11570), .A(n10223), .B(n10222), .ZN(
        n10224) );
  INV_X1 U12818 ( .A(n10224), .ZN(n10225) );
  NAND2_X1 U12819 ( .A1(n12350), .A2(P3_DATAO_REG_29__SCAN_IN), .ZN(n10226) );
  OAI21_X1 U12820 ( .B1(n12520), .B2(n12350), .A(n10226), .ZN(P3_U3520) );
  INV_X1 U12821 ( .A(n10227), .ZN(n10235) );
  NOR2_X1 U12822 ( .A1(n13311), .A2(n10228), .ZN(n10230) );
  OAI22_X1 U12823 ( .A1(n13281), .A2(n9301), .B1(P2_REG3_REG_3__SCAN_IN), .B2(
        n13323), .ZN(n10229) );
  AOI211_X1 U12824 ( .C1(n10231), .C2(n14362), .A(n10230), .B(n10229), .ZN(
        n10234) );
  NAND2_X1 U12825 ( .A1(n10232), .A2(n13281), .ZN(n10233) );
  OAI211_X1 U12826 ( .C1(n10235), .C2(n13342), .A(n10234), .B(n10233), .ZN(
        P2_U3262) );
  XNOR2_X1 U12827 ( .A(n12008), .B(n6540), .ZN(n10236) );
  NAND2_X1 U12828 ( .A1(n13042), .A2(n13326), .ZN(n10237) );
  NAND2_X1 U12829 ( .A1(n10236), .A2(n10237), .ZN(n10328) );
  INV_X1 U12830 ( .A(n10236), .ZN(n10239) );
  INV_X1 U12831 ( .A(n10237), .ZN(n10238) );
  NAND2_X1 U12832 ( .A1(n10239), .A2(n10238), .ZN(n10240) );
  AND2_X1 U12833 ( .A1(n10328), .A2(n10240), .ZN(n10244) );
  OAI21_X1 U12834 ( .B1(n10244), .B2(n10243), .A(n10329), .ZN(n10245) );
  NAND2_X1 U12835 ( .A1(n10245), .A2(n12973), .ZN(n10252) );
  INV_X1 U12836 ( .A(n10246), .ZN(n10490) );
  INV_X1 U12837 ( .A(n13016), .ZN(n14343) );
  OAI22_X1 U12838 ( .A1(n10248), .A2(n12946), .B1(n10247), .B2(n12948), .ZN(
        n10481) );
  INV_X1 U12839 ( .A(n10481), .ZN(n10249) );
  NAND2_X1 U12840 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(P2_U3088), .ZN(n14701) );
  OAI21_X1 U12841 ( .B1(n14343), .B2(n10249), .A(n14701), .ZN(n10250) );
  AOI21_X1 U12842 ( .B1(n10490), .B2(n13000), .A(n10250), .ZN(n10251) );
  OAI211_X1 U12843 ( .C1(n14807), .C2(n14340), .A(n10252), .B(n10251), .ZN(
        P2_U3203) );
  INV_X1 U12844 ( .A(P3_DATAO_REG_31__SCAN_IN), .ZN(n15336) );
  INV_X1 U12845 ( .A(P3_REG2_REG_31__SCAN_IN), .ZN(n10256) );
  NAND2_X1 U12846 ( .A1(n11521), .A2(P3_REG1_REG_31__SCAN_IN), .ZN(n10255) );
  INV_X1 U12847 ( .A(P3_REG0_REG_31__SCAN_IN), .ZN(n10253) );
  OR2_X1 U12848 ( .A1(n11438), .A2(n10253), .ZN(n10254) );
  NAND2_X1 U12849 ( .A1(n10303), .A2(n6699), .ZN(n12508) );
  NAND2_X1 U12850 ( .A1(n12508), .A2(P3_U3897), .ZN(n10257) );
  OAI21_X1 U12851 ( .B1(P3_U3897), .B2(n15336), .A(n10257), .ZN(P3_U3522) );
  OR2_X1 U12852 ( .A1(n11662), .A2(SI_5_), .ZN(n10261) );
  OR2_X1 U12853 ( .A1(n10001), .A2(n10258), .ZN(n10260) );
  NAND2_X1 U12854 ( .A1(n11492), .A2(n14875), .ZN(n10259) );
  XNOR2_X1 U12855 ( .A(n11892), .B(n10710), .ZN(n10430) );
  XNOR2_X1 U12856 ( .A(n10430), .B(n12346), .ZN(n10265) );
  NAND2_X1 U12857 ( .A1(n10263), .A2(n10262), .ZN(n10264) );
  NAND2_X1 U12858 ( .A1(n10264), .A2(n10265), .ZN(n10542) );
  OAI21_X1 U12859 ( .B1(n10265), .B2(n10264), .A(n10542), .ZN(n10266) );
  NAND2_X1 U12860 ( .A1(n10266), .A2(n12318), .ZN(n10278) );
  INV_X1 U12861 ( .A(P3_REG1_REG_6__SCAN_IN), .ZN(n10932) );
  OR2_X1 U12862 ( .A1(n11436), .A2(n10932), .ZN(n10271) );
  NAND2_X1 U12863 ( .A1(n10267), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n10268) );
  AND2_X1 U12864 ( .A1(n10384), .A2(n10268), .ZN(n15016) );
  OR2_X1 U12865 ( .A1(n10012), .A2(n15016), .ZN(n10270) );
  INV_X1 U12866 ( .A(P3_REG2_REG_6__SCAN_IN), .ZN(n10933) );
  NAND2_X1 U12867 ( .A1(n15389), .A2(n12345), .ZN(n10274) );
  AND2_X1 U12868 ( .A1(P3_U3151), .A2(P3_REG3_REG_5__SCAN_IN), .ZN(n14877) );
  INV_X1 U12869 ( .A(n14877), .ZN(n10273) );
  OAI211_X1 U12870 ( .C1(n10709), .C2(n15392), .A(n10274), .B(n10273), .ZN(
        n10276) );
  NOR2_X1 U12871 ( .A1(n15395), .A2(n10711), .ZN(n10275) );
  AOI211_X1 U12872 ( .C1(n15399), .C2(n10710), .A(n10276), .B(n10275), .ZN(
        n10277) );
  NAND2_X1 U12873 ( .A1(n10278), .A2(n10277), .ZN(P3_U3167) );
  INV_X1 U12874 ( .A(SI_23_), .ZN(n15291) );
  INV_X1 U12875 ( .A(n10279), .ZN(n10280) );
  XNOR2_X1 U12876 ( .A(n11013), .B(P2_DATAO_REG_23__SCAN_IN), .ZN(n10787) );
  XNOR2_X1 U12877 ( .A(n10788), .B(n10787), .ZN(n11526) );
  NAND2_X1 U12878 ( .A1(n11526), .A2(n12881), .ZN(n10284) );
  OAI211_X1 U12879 ( .C1(n15291), .C2(n11338), .A(n10284), .B(n11864), .ZN(
        P3_U3272) );
  INV_X1 U12880 ( .A(n14517), .ZN(n14621) );
  NAND2_X1 U12881 ( .A1(n14517), .A2(n13640), .ZN(n10289) );
  NAND2_X1 U12882 ( .A1(n13767), .A2(n6536), .ZN(n10288) );
  NAND2_X1 U12883 ( .A1(n10289), .A2(n10288), .ZN(n10290) );
  XNOR2_X1 U12884 ( .A(n10290), .B(n13637), .ZN(n10603) );
  AND2_X1 U12885 ( .A1(n13767), .A2(n13636), .ZN(n10291) );
  AOI21_X1 U12886 ( .B1(n14517), .B2(n6536), .A(n10291), .ZN(n10601) );
  XNOR2_X1 U12887 ( .A(n10603), .B(n10601), .ZN(n10292) );
  OAI211_X1 U12888 ( .C1(n10293), .C2(n10292), .A(n10605), .B(n14395), .ZN(
        n10297) );
  OAI22_X1 U12889 ( .A1(n10314), .A2(n14561), .B1(n10498), .B2(n14581), .ZN(
        n14514) );
  NOR2_X1 U12890 ( .A1(n14401), .A2(n14515), .ZN(n10294) );
  AOI211_X1 U12891 ( .C1(n14397), .C2(n14514), .A(n10295), .B(n10294), .ZN(
        n10296) );
  OAI211_X1 U12892 ( .C1(n14621), .C2(n13743), .A(n10297), .B(n10296), .ZN(
        P1_U3213) );
  INV_X1 U12893 ( .A(P3_DATAO_REG_30__SCAN_IN), .ZN(n15198) );
  INV_X1 U12894 ( .A(P3_REG1_REG_30__SCAN_IN), .ZN(n10300) );
  NAND2_X1 U12895 ( .A1(n11567), .A2(P3_REG2_REG_30__SCAN_IN), .ZN(n10299) );
  OAI211_X1 U12896 ( .C1(n10300), .C2(n11570), .A(n10299), .B(n10298), .ZN(
        n10301) );
  INV_X1 U12897 ( .A(n10301), .ZN(n10302) );
  NAND2_X1 U12898 ( .A1(n10303), .A2(n10302), .ZN(n11665) );
  NAND2_X1 U12899 ( .A1(n11665), .A2(P3_U3897), .ZN(n10304) );
  OAI21_X1 U12900 ( .B1(P3_U3897), .B2(n15198), .A(n10304), .ZN(P3_U3521) );
  INV_X1 U12901 ( .A(n10305), .ZN(n10306) );
  NAND2_X1 U12902 ( .A1(n10307), .A2(n10306), .ZN(n10309) );
  OR2_X1 U12903 ( .A1(n10315), .A2(n13768), .ZN(n10308) );
  NAND2_X1 U12904 ( .A1(n10309), .A2(n10308), .ZN(n14508) );
  NAND2_X1 U12905 ( .A1(n14508), .A2(n14512), .ZN(n10313) );
  NAND2_X1 U12906 ( .A1(n14621), .A2(n10311), .ZN(n10312) );
  NAND2_X1 U12907 ( .A1(n10313), .A2(n10312), .ZN(n10513) );
  INV_X1 U12908 ( .A(n10512), .ZN(n10500) );
  XNOR2_X1 U12909 ( .A(n10500), .B(n10513), .ZN(n10368) );
  AOI211_X1 U12910 ( .C1(n10600), .C2(n14518), .A(n14572), .B(n14504), .ZN(
        n10365) );
  AOI21_X1 U12911 ( .B1(n10600), .B2(n14607), .A(n10365), .ZN(n10323) );
  NAND2_X1 U12912 ( .A1(n10315), .A2(n10314), .ZN(n10316) );
  NAND2_X1 U12913 ( .A1(n14621), .A2(n13767), .ZN(n10318) );
  XNOR2_X1 U12914 ( .A(n10501), .B(n10512), .ZN(n10322) );
  NAND2_X1 U12915 ( .A1(n13767), .A2(n14107), .ZN(n10320) );
  NAND2_X1 U12916 ( .A1(n13765), .A2(n14108), .ZN(n10319) );
  AND2_X1 U12917 ( .A1(n10320), .A2(n10319), .ZN(n10610) );
  INV_X1 U12918 ( .A(n10610), .ZN(n10321) );
  AOI21_X1 U12919 ( .B1(n10322), .B2(n14497), .A(n10321), .ZN(n10361) );
  OAI211_X1 U12920 ( .C1(n14611), .C2(n10368), .A(n10323), .B(n10361), .ZN(
        n10325) );
  NAND2_X1 U12921 ( .A1(n10325), .A2(n14658), .ZN(n10324) );
  OAI21_X1 U12922 ( .B1(n14658), .B2(n9099), .A(n10324), .ZN(P1_U3536) );
  INV_X1 U12923 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n10327) );
  NAND2_X1 U12924 ( .A1(n10325), .A2(n14645), .ZN(n10326) );
  OAI21_X1 U12925 ( .B1(n14645), .B2(n10327), .A(n10326), .ZN(P1_U3483) );
  XNOR2_X1 U12926 ( .A(n14811), .B(n6541), .ZN(n10616) );
  NAND2_X1 U12927 ( .A1(n13041), .A2(n13326), .ZN(n10617) );
  XNOR2_X1 U12928 ( .A(n10616), .B(n10617), .ZN(n10621) );
  XNOR2_X1 U12929 ( .A(n10621), .B(n10622), .ZN(n10335) );
  NAND2_X1 U12930 ( .A1(n13042), .A2(n14334), .ZN(n10331) );
  NAND2_X1 U12931 ( .A1(n13040), .A2(n14336), .ZN(n10330) );
  NAND2_X1 U12932 ( .A1(n10331), .A2(n10330), .ZN(n10417) );
  AND2_X1 U12933 ( .A1(P2_U3088), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n14706) );
  AOI21_X1 U12934 ( .B1(n13016), .B2(n10417), .A(n14706), .ZN(n10332) );
  OAI21_X1 U12935 ( .B1(n10424), .B2(n14348), .A(n10332), .ZN(n10333) );
  AOI21_X1 U12936 ( .B1(n14811), .B2(n13019), .A(n10333), .ZN(n10334) );
  OAI21_X1 U12937 ( .B1(n10335), .B2(n14342), .A(n10334), .ZN(P2_U3189) );
  NAND2_X1 U12938 ( .A1(n10336), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n10338) );
  NAND2_X1 U12939 ( .A1(n10338), .A2(n10337), .ZN(n10692) );
  XNOR2_X1 U12940 ( .A(n10692), .B(n10342), .ZN(n10339) );
  NOR2_X1 U12941 ( .A1(P1_REG2_REG_15__SCAN_IN), .A2(n10339), .ZN(n10693) );
  AOI21_X1 U12942 ( .B1(n10339), .B2(P1_REG2_REG_15__SCAN_IN), .A(n10693), 
        .ZN(n10349) );
  AOI21_X1 U12943 ( .B1(n8554), .B2(n10341), .A(n10340), .ZN(n10687) );
  XNOR2_X1 U12944 ( .A(n10687), .B(n10342), .ZN(n10343) );
  AND2_X1 U12945 ( .A1(n10343), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n10344) );
  NOR2_X1 U12946 ( .A1(P1_REG1_REG_15__SCAN_IN), .A2(n10343), .ZN(n10688) );
  OAI21_X1 U12947 ( .B1(n10344), .B2(n10688), .A(n14483), .ZN(n10348) );
  INV_X1 U12948 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n13747) );
  NOR2_X1 U12949 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n13747), .ZN(n10346) );
  NOR2_X1 U12950 ( .A1(n13832), .A2(n10695), .ZN(n10345) );
  AOI211_X1 U12951 ( .C1(n14472), .C2(P1_ADDR_REG_15__SCAN_IN), .A(n10346), 
        .B(n10345), .ZN(n10347) );
  OAI211_X1 U12952 ( .C1(n10349), .C2(n14464), .A(n10348), .B(n10347), .ZN(
        P1_U3258) );
  AND2_X1 U12953 ( .A1(n14362), .A2(n9550), .ZN(n13316) );
  OAI21_X1 U12954 ( .B1(n14355), .B2(n13316), .A(n11935), .ZN(n10351) );
  AOI22_X1 U12955 ( .A1(n14367), .A2(P2_REG2_REG_0__SCAN_IN), .B1(n14354), 
        .B2(P2_REG3_REG_0__SCAN_IN), .ZN(n10350) );
  OAI211_X1 U12956 ( .C1(n10421), .C2(n12190), .A(n10351), .B(n10350), .ZN(
        n10352) );
  AOI21_X1 U12957 ( .B1(n13281), .B2(n10353), .A(n10352), .ZN(n10354) );
  INV_X1 U12958 ( .A(n10354), .ZN(P2_U3265) );
  INV_X1 U12959 ( .A(P3_DATAO_REG_28__SCAN_IN), .ZN(n15257) );
  NOR2_X1 U12960 ( .A1(n11562), .A2(n11898), .ZN(n10355) );
  INV_X1 U12961 ( .A(P3_REG1_REG_28__SCAN_IN), .ZN(n12733) );
  NAND2_X1 U12962 ( .A1(n11567), .A2(P3_REG2_REG_28__SCAN_IN), .ZN(n10357) );
  OAI211_X1 U12963 ( .C1(n12733), .C2(n11570), .A(n10357), .B(n10356), .ZN(
        n10358) );
  NAND2_X1 U12964 ( .A1(n11616), .A2(P3_U3897), .ZN(n10359) );
  OAI21_X1 U12965 ( .B1(P3_U3897), .B2(n15257), .A(n10359), .ZN(P3_U3519) );
  INV_X1 U12966 ( .A(n10360), .ZN(n10612) );
  INV_X1 U12967 ( .A(n10361), .ZN(n10362) );
  AOI21_X1 U12968 ( .B1(n10612), .B2(n14567), .A(n10362), .ZN(n10363) );
  MUX2_X1 U12969 ( .A(n10364), .B(n10363), .S(n14543), .Z(n10367) );
  AOI22_X1 U12970 ( .A1(n10365), .A2(n14574), .B1(n14566), .B2(n10600), .ZN(
        n10366) );
  OAI211_X1 U12971 ( .C1(n14123), .C2(n10368), .A(n10367), .B(n10366), .ZN(
        P1_U3285) );
  NAND2_X1 U12972 ( .A1(n12348), .A2(n10369), .ZN(n10370) );
  NAND2_X1 U12973 ( .A1(n10371), .A2(n10370), .ZN(n10637) );
  NAND2_X1 U12974 ( .A1(n10709), .A2(n10633), .ZN(n11704) );
  INV_X1 U12975 ( .A(n10633), .ZN(n10372) );
  NAND2_X1 U12976 ( .A1(n12347), .A2(n10372), .ZN(n11705) );
  NAND2_X1 U12977 ( .A1(n11704), .A2(n11705), .ZN(n10636) );
  NAND2_X1 U12978 ( .A1(n12347), .A2(n10633), .ZN(n10373) );
  NAND2_X1 U12979 ( .A1(n10638), .A2(n10710), .ZN(n11709) );
  INV_X1 U12980 ( .A(n10710), .ZN(n10379) );
  NAND2_X1 U12981 ( .A1(n12346), .A2(n10379), .ZN(n11708) );
  INV_X1 U12982 ( .A(n11826), .ZN(n10374) );
  OR2_X1 U12983 ( .A1(n11662), .A2(n10375), .ZN(n10378) );
  OR2_X1 U12984 ( .A1(n10001), .A2(n10376), .ZN(n10377) );
  OAI211_X1 U12985 ( .C1(n9726), .C2(n14893), .A(n10378), .B(n10377), .ZN(
        n15013) );
  NAND2_X1 U12986 ( .A1(n10708), .A2(n15013), .ZN(n11710) );
  INV_X1 U12987 ( .A(n15013), .ZN(n10411) );
  NAND2_X1 U12988 ( .A1(n12345), .A2(n10411), .ZN(n11719) );
  NAND2_X1 U12989 ( .A1(n11710), .A2(n11719), .ZN(n10405) );
  NAND2_X1 U12990 ( .A1(n10638), .A2(n10379), .ZN(n10381) );
  AND2_X1 U12991 ( .A1(n10405), .A2(n10381), .ZN(n10380) );
  NAND2_X1 U12992 ( .A1(n10704), .A2(n10380), .ZN(n10751) );
  INV_X1 U12993 ( .A(n10751), .ZN(n10383) );
  AOI21_X1 U12994 ( .B1(n10704), .B2(n10381), .A(n10405), .ZN(n10382) );
  NOR3_X1 U12995 ( .A1(n10383), .A2(n10382), .A3(n15027), .ZN(n10391) );
  AND2_X1 U12996 ( .A1(n10384), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n10385) );
  NOR2_X1 U12997 ( .A1(n10532), .A2(n10385), .ZN(n15006) );
  OR2_X1 U12998 ( .A1(n10012), .A2(n15006), .ZN(n10388) );
  INV_X1 U12999 ( .A(P3_REG1_REG_7__SCAN_IN), .ZN(n10939) );
  OR2_X1 U13000 ( .A1(n11436), .A2(n10939), .ZN(n10387) );
  INV_X1 U13001 ( .A(P3_REG2_REG_7__SCAN_IN), .ZN(n10940) );
  OAI22_X1 U13002 ( .A1(n10545), .A2(n15031), .B1(n10638), .B2(n15029), .ZN(
        n10390) );
  NOR2_X1 U13003 ( .A1(n10391), .A2(n10390), .ZN(n15008) );
  INV_X1 U13004 ( .A(n10392), .ZN(n10394) );
  OAI22_X1 U13005 ( .A1(n10395), .A2(n10394), .B1(n10398), .B2(n10393), .ZN(
        n10397) );
  NAND2_X1 U13006 ( .A1(n10397), .A2(n10396), .ZN(n10402) );
  INV_X1 U13007 ( .A(n10398), .ZN(n10400) );
  NAND2_X1 U13008 ( .A1(n10400), .A2(n10399), .ZN(n10401) );
  NAND2_X1 U13009 ( .A1(n10403), .A2(n11825), .ZN(n10404) );
  NAND2_X1 U13010 ( .A1(n10404), .A2(n11699), .ZN(n10632) );
  INV_X1 U13011 ( .A(n10636), .ZN(n11830) );
  NAND2_X1 U13012 ( .A1(n10631), .A2(n11704), .ZN(n10703) );
  NAND2_X1 U13013 ( .A1(n10748), .A2(n11709), .ZN(n10407) );
  INV_X1 U13014 ( .A(n10405), .ZN(n11831) );
  NAND2_X1 U13015 ( .A1(n10407), .A2(n11831), .ZN(n10406) );
  OAI21_X1 U13016 ( .B1(n10407), .B2(n11831), .A(n10406), .ZN(n15007) );
  INV_X1 U13017 ( .A(n10408), .ZN(n15043) );
  NAND2_X1 U13018 ( .A1(n11860), .A2(n15022), .ZN(n15058) );
  INV_X1 U13019 ( .A(n12859), .ZN(n12872) );
  INV_X1 U13020 ( .A(P3_REG0_REG_6__SCAN_IN), .ZN(n15278) );
  OAI22_X1 U13021 ( .A1(n10411), .A2(n12867), .B1(n15085), .B2(n15278), .ZN(
        n10409) );
  AOI21_X1 U13022 ( .B1(n15007), .B2(n12872), .A(n10409), .ZN(n10410) );
  OAI21_X1 U13023 ( .B1(n15008), .B2(n15086), .A(n10410), .ZN(P3_U3408) );
  NAND2_X1 U13024 ( .A1(n15083), .A2(n15096), .ZN(n12776) );
  INV_X1 U13025 ( .A(n12776), .ZN(n12783) );
  OAI22_X1 U13026 ( .A1(n12780), .A2(n10411), .B1(n15096), .B2(n10932), .ZN(
        n10412) );
  AOI21_X1 U13027 ( .B1(n15007), .B2(n12783), .A(n10412), .ZN(n10413) );
  OAI21_X1 U13028 ( .B1(n15008), .B2(n15094), .A(n10413), .ZN(P3_U3465) );
  XNOR2_X1 U13029 ( .A(n14811), .B(n13041), .ZN(n12204) );
  XNOR2_X1 U13030 ( .A(n10414), .B(n12204), .ZN(n14816) );
  NAND2_X1 U13031 ( .A1(n14816), .A2(n13307), .ZN(n10420) );
  INV_X1 U13032 ( .A(n12204), .ZN(n10415) );
  XNOR2_X1 U13033 ( .A(n10416), .B(n10415), .ZN(n10418) );
  AOI21_X1 U13034 ( .B1(n10418), .B2(n13335), .A(n10417), .ZN(n10419) );
  AND2_X1 U13035 ( .A1(n10420), .A2(n10419), .ZN(n14818) );
  INV_X1 U13036 ( .A(n10421), .ZN(n13317) );
  NAND2_X1 U13037 ( .A1(n14811), .A2(n10489), .ZN(n10422) );
  NAND2_X1 U13038 ( .A1(n10422), .A2(n9550), .ZN(n10423) );
  OR2_X1 U13039 ( .A1(n6814), .A2(n10423), .ZN(n14813) );
  OAI22_X1 U13040 ( .A1(n13281), .A2(n10425), .B1(n10424), .B2(n13323), .ZN(
        n10426) );
  AOI21_X1 U13041 ( .B1(n14811), .B2(n14355), .A(n10426), .ZN(n10427) );
  OAI21_X1 U13042 ( .B1(n14813), .B2(n13330), .A(n10427), .ZN(n10428) );
  AOI21_X1 U13043 ( .B1(n14816), .B2(n13317), .A(n10428), .ZN(n10429) );
  OAI21_X1 U13044 ( .B1(n14818), .B2(n14367), .A(n10429), .ZN(P2_U3255) );
  NAND2_X1 U13045 ( .A1(n10430), .A2(n10638), .ZN(n10540) );
  AND2_X1 U13046 ( .A1(n10542), .A2(n10540), .ZN(n10432) );
  XNOR2_X1 U13047 ( .A(n11892), .B(n15013), .ZN(n10543) );
  XNOR2_X1 U13048 ( .A(n10543), .B(n12345), .ZN(n10431) );
  NAND2_X1 U13049 ( .A1(n10432), .A2(n10431), .ZN(n10659) );
  OAI211_X1 U13050 ( .C1(n10432), .C2(n10431), .A(n10659), .B(n12318), .ZN(
        n10439) );
  NAND2_X1 U13051 ( .A1(n15389), .A2(n12344), .ZN(n10435) );
  INV_X1 U13052 ( .A(P3_REG3_REG_6__SCAN_IN), .ZN(n10433) );
  NOR2_X1 U13053 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n10433), .ZN(n14895) );
  INV_X1 U13054 ( .A(n14895), .ZN(n10434) );
  OAI211_X1 U13055 ( .C1(n10638), .C2(n15392), .A(n10435), .B(n10434), .ZN(
        n10437) );
  NOR2_X1 U13056 ( .A1(n15395), .A2(n15016), .ZN(n10436) );
  AOI211_X1 U13057 ( .C1(n15399), .C2(n15013), .A(n10437), .B(n10436), .ZN(
        n10438) );
  NAND2_X1 U13058 ( .A1(n10439), .A2(n10438), .ZN(P3_U3179) );
  INV_X1 U13059 ( .A(n10440), .ZN(n10448) );
  INV_X1 U13060 ( .A(n13342), .ZN(n14363) );
  OAI22_X1 U13061 ( .A1(n13281), .A2(n15230), .B1(n7578), .B2(n13323), .ZN(
        n10441) );
  AOI21_X1 U13062 ( .B1(n14362), .B2(n10442), .A(n10441), .ZN(n10443) );
  OAI21_X1 U13063 ( .B1(n10444), .B2(n13311), .A(n10443), .ZN(n10445) );
  AOI21_X1 U13064 ( .B1(n14363), .B2(n10446), .A(n10445), .ZN(n10447) );
  OAI21_X1 U13065 ( .B1(n14367), .B2(n10448), .A(n10447), .ZN(P2_U3264) );
  INV_X1 U13066 ( .A(n10449), .ZN(n10457) );
  NAND2_X1 U13067 ( .A1(n10450), .A2(n14362), .ZN(n10452) );
  AOI22_X1 U13068 ( .A1(n14367), .A2(P2_REG2_REG_2__SCAN_IN), .B1(n14354), 
        .B2(P2_REG3_REG_2__SCAN_IN), .ZN(n10451) );
  OAI211_X1 U13069 ( .C1(n10453), .C2(n13311), .A(n10452), .B(n10451), .ZN(
        n10454) );
  AOI21_X1 U13070 ( .B1(n14363), .B2(n10455), .A(n10454), .ZN(n10456) );
  OAI21_X1 U13071 ( .B1(n14367), .B2(n10457), .A(n10456), .ZN(P2_U3263) );
  INV_X1 U13072 ( .A(n10458), .ZN(n10496) );
  OAI222_X1 U13073 ( .A1(n10459), .A2(P1_U3086), .B1(n6535), .B2(n10496), .C1(
        n15263), .C2(n14266), .ZN(P1_U3335) );
  INV_X1 U13074 ( .A(n10460), .ZN(n10462) );
  INV_X1 U13075 ( .A(n13839), .ZN(n13831) );
  OAI222_X1 U13076 ( .A1(n14266), .A2(n10461), .B1(n6535), .B2(n10462), .C1(
        n13831), .C2(P1_U3086), .ZN(P1_U3337) );
  INV_X1 U13077 ( .A(n13135), .ZN(n11366) );
  OAI222_X1 U13078 ( .A1(n11904), .A2(n10463), .B1(n6534), .B2(n10462), .C1(
        P2_U3088), .C2(n11366), .ZN(P2_U3309) );
  XNOR2_X1 U13079 ( .A(n10464), .B(n12201), .ZN(n10466) );
  AOI21_X1 U13080 ( .B1(n10466), .B2(n13335), .A(n10465), .ZN(n14799) );
  NAND2_X1 U13081 ( .A1(n10467), .A2(n12201), .ZN(n10468) );
  NAND2_X1 U13082 ( .A1(n10469), .A2(n10468), .ZN(n14794) );
  INV_X1 U13083 ( .A(n14794), .ZN(n10478) );
  NAND2_X1 U13084 ( .A1(n14795), .A2(n10471), .ZN(n10472) );
  NAND3_X1 U13085 ( .A1(n10487), .A2(n9550), .A3(n10472), .ZN(n14797) );
  OAI22_X1 U13086 ( .A1(n13281), .A2(n10474), .B1(n10473), .B2(n13323), .ZN(
        n10475) );
  AOI21_X1 U13087 ( .B1(n14795), .B2(n14355), .A(n10475), .ZN(n10476) );
  OAI21_X1 U13088 ( .B1(n14797), .B2(n13330), .A(n10476), .ZN(n10477) );
  AOI21_X1 U13089 ( .B1(n10478), .B2(n14363), .A(n10477), .ZN(n10479) );
  OAI21_X1 U13090 ( .B1(n14367), .B2(n14799), .A(n10479), .ZN(P2_U3257) );
  AOI21_X1 U13091 ( .B1(n10480), .B2(n10485), .A(n14351), .ZN(n10483) );
  AOI21_X1 U13092 ( .B1(n10483), .B2(n10482), .A(n10481), .ZN(n14805) );
  OAI21_X1 U13093 ( .B1(n10486), .B2(n10485), .A(n10484), .ZN(n14802) );
  INV_X1 U13094 ( .A(n14802), .ZN(n10494) );
  AOI21_X1 U13095 ( .B1(n12008), .B2(n10487), .A(n9445), .ZN(n10488) );
  NAND2_X1 U13096 ( .A1(n10489), .A2(n10488), .ZN(n14804) );
  AOI22_X1 U13097 ( .A1(n14367), .A2(P2_REG2_REG_9__SCAN_IN), .B1(n14354), 
        .B2(n10490), .ZN(n10492) );
  NAND2_X1 U13098 ( .A1(n12008), .A2(n14355), .ZN(n10491) );
  OAI211_X1 U13099 ( .C1(n14804), .C2(n13330), .A(n10492), .B(n10491), .ZN(
        n10493) );
  AOI21_X1 U13100 ( .B1(n10494), .B2(n14363), .A(n10493), .ZN(n10495) );
  OAI21_X1 U13101 ( .B1(n14367), .B2(n14805), .A(n10495), .ZN(P2_U3256) );
  OAI222_X1 U13102 ( .A1(n11904), .A2(n10497), .B1(P2_U3088), .B2(n12183), 
        .C1(n6534), .C2(n10496), .ZN(P2_U3307) );
  NOR2_X1 U13103 ( .A1(n10600), .A2(n10498), .ZN(n10499) );
  NAND2_X1 U13104 ( .A1(n14490), .A2(n14491), .ZN(n14489) );
  INV_X1 U13105 ( .A(n13765), .ZN(n10502) );
  NAND2_X1 U13106 ( .A1(n14500), .A2(n10502), .ZN(n10503) );
  NAND2_X1 U13107 ( .A1(n14489), .A2(n10503), .ZN(n10505) );
  AOI21_X1 U13108 ( .B1(n10505), .B2(n10810), .A(n14560), .ZN(n10507) );
  INV_X1 U13109 ( .A(n10505), .ZN(n10506) );
  AOI22_X1 U13110 ( .A1(n10507), .A2(n10807), .B1(n14107), .B2(n13765), .ZN(
        n14636) );
  OAI22_X1 U13111 ( .A1(n14543), .A2(n10508), .B1(n10836), .B2(n14542), .ZN(
        n10511) );
  INV_X1 U13112 ( .A(n14500), .ZN(n14628) );
  NAND2_X1 U13113 ( .A1(n14628), .A2(n14504), .ZN(n14503) );
  AOI211_X1 U13114 ( .C1(n14635), .C2(n14503), .A(n14572), .B(n10816), .ZN(
        n10509) );
  AOI21_X1 U13115 ( .B1(n14108), .B2(n13763), .A(n10509), .ZN(n14637) );
  NOR2_X1 U13116 ( .A1(n14637), .A2(n13959), .ZN(n10510) );
  AOI211_X1 U13117 ( .C1(n14566), .C2(n14635), .A(n10511), .B(n10510), .ZN(
        n10520) );
  NAND2_X1 U13118 ( .A1(n10513), .A2(n10512), .ZN(n10515) );
  OR2_X1 U13119 ( .A1(n10600), .A2(n13766), .ZN(n10514) );
  NAND2_X1 U13120 ( .A1(n10515), .A2(n10514), .ZN(n14492) );
  INV_X1 U13121 ( .A(n14491), .ZN(n10516) );
  NAND2_X1 U13122 ( .A1(n14492), .A2(n10516), .ZN(n10518) );
  OR2_X1 U13123 ( .A1(n14500), .A2(n13765), .ZN(n10517) );
  NAND2_X1 U13124 ( .A1(n10518), .A2(n10517), .ZN(n10811) );
  XNOR2_X1 U13125 ( .A(n10811), .B(n10810), .ZN(n14642) );
  NAND2_X1 U13126 ( .A1(n14642), .A2(n14083), .ZN(n10519) );
  OAI211_X1 U13127 ( .C1(n6531), .C2(n14636), .A(n10520), .B(n10519), .ZN(
        P1_U3283) );
  OR2_X1 U13128 ( .A1(n11662), .A2(SI_7_), .ZN(n10524) );
  OR2_X1 U13129 ( .A1(n10001), .A2(n10521), .ZN(n10523) );
  NAND2_X1 U13130 ( .A1(n11492), .A2(n14911), .ZN(n10522) );
  NAND2_X1 U13131 ( .A1(n10545), .A2(n15004), .ZN(n11720) );
  INV_X1 U13132 ( .A(n15004), .ZN(n10759) );
  NAND2_X1 U13133 ( .A1(n12344), .A2(n10759), .ZN(n11717) );
  XNOR2_X1 U13134 ( .A(n10752), .B(n10525), .ZN(n10660) );
  OR2_X1 U13135 ( .A1(n10001), .A2(n10526), .ZN(n10529) );
  OR2_X1 U13136 ( .A1(n11662), .A2(n10527), .ZN(n10528) );
  OAI211_X1 U13137 ( .C1(n10530), .C2(n14928), .A(n10529), .B(n10528), .ZN(
        n14996) );
  XNOR2_X1 U13138 ( .A(n10531), .B(n14996), .ZN(n10547) );
  NOR2_X1 U13139 ( .A1(n10532), .A2(n10798), .ZN(n10533) );
  OR2_X1 U13140 ( .A1(n10558), .A2(n10533), .ZN(n14997) );
  INV_X1 U13141 ( .A(n14997), .ZN(n10801) );
  INV_X1 U13142 ( .A(P3_REG1_REG_8__SCAN_IN), .ZN(n10945) );
  OR2_X1 U13143 ( .A1(n11436), .A2(n10945), .ZN(n10534) );
  OAI21_X1 U13144 ( .B1(n10012), .B2(n10801), .A(n10534), .ZN(n10538) );
  INV_X1 U13145 ( .A(P3_REG2_REG_8__SCAN_IN), .ZN(n10946) );
  INV_X1 U13146 ( .A(P3_REG0_REG_8__SCAN_IN), .ZN(n10535) );
  NOR2_X1 U13147 ( .A1(n11438), .A2(n10535), .ZN(n10536) );
  XNOR2_X1 U13148 ( .A(n10547), .B(n12343), .ZN(n10796) );
  NAND2_X1 U13149 ( .A1(n10543), .A2(n10708), .ZN(n10539) );
  AND4_X1 U13150 ( .A1(n10660), .A2(n10796), .A3(n10540), .A4(n10539), .ZN(
        n10541) );
  NAND2_X1 U13151 ( .A1(n10542), .A2(n10541), .ZN(n10552) );
  INV_X1 U13152 ( .A(n10796), .ZN(n10546) );
  INV_X1 U13153 ( .A(n10543), .ZN(n10544) );
  NAND2_X1 U13154 ( .A1(n10544), .A2(n12345), .ZN(n10658) );
  OAI21_X1 U13155 ( .B1(n10546), .B2(n10658), .A(n10660), .ZN(n10550) );
  INV_X1 U13156 ( .A(n10660), .ZN(n10794) );
  OAI21_X1 U13157 ( .B1(n10546), .B2(n10545), .A(n10794), .ZN(n10549) );
  INV_X1 U13158 ( .A(n10547), .ZN(n10548) );
  AOI22_X1 U13159 ( .A1(n10550), .A2(n10549), .B1(n10548), .B2(n12343), .ZN(
        n10551) );
  OR2_X1 U13160 ( .A1(n10001), .A2(n10553), .ZN(n10556) );
  OR2_X1 U13161 ( .A1(n11662), .A2(SI_9_), .ZN(n10555) );
  NAND2_X1 U13162 ( .A1(n11492), .A2(n14946), .ZN(n10554) );
  XNOR2_X1 U13163 ( .A(n11892), .B(n11730), .ZN(n10576) );
  OR2_X1 U13164 ( .A1(n10558), .A2(n10557), .ZN(n10559) );
  AND2_X1 U13165 ( .A1(n10570), .A2(n10559), .ZN(n11107) );
  INV_X1 U13166 ( .A(P3_REG1_REG_9__SCAN_IN), .ZN(n10952) );
  OR2_X1 U13167 ( .A1(n11436), .A2(n10952), .ZN(n10560) );
  OAI21_X1 U13168 ( .B1(n10012), .B2(n11107), .A(n10560), .ZN(n10564) );
  INV_X1 U13169 ( .A(P3_REG2_REG_9__SCAN_IN), .ZN(n10953) );
  INV_X1 U13170 ( .A(P3_REG0_REG_9__SCAN_IN), .ZN(n10561) );
  NOR2_X1 U13171 ( .A1(n11438), .A2(n10561), .ZN(n10562) );
  XNOR2_X1 U13172 ( .A(n10576), .B(n11472), .ZN(n11059) );
  OR2_X1 U13173 ( .A1(n11066), .A2(n11059), .ZN(n10717) );
  NAND2_X1 U13174 ( .A1(n10565), .A2(n11664), .ZN(n10568) );
  NAND2_X1 U13175 ( .A1(n11492), .A2(n14965), .ZN(n10567) );
  OR2_X1 U13176 ( .A1(n11662), .A2(SI_10_), .ZN(n10566) );
  XNOR2_X1 U13177 ( .A(n11892), .B(n14988), .ZN(n11057) );
  NAND2_X1 U13178 ( .A1(n11567), .A2(P3_REG2_REG_10__SCAN_IN), .ZN(n10575) );
  INV_X1 U13179 ( .A(P3_REG0_REG_10__SCAN_IN), .ZN(n10569) );
  OR2_X1 U13180 ( .A1(n11438), .A2(n10569), .ZN(n10574) );
  NAND2_X1 U13181 ( .A1(n10570), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n10571) );
  AND2_X1 U13182 ( .A1(n10580), .A2(n10571), .ZN(n14989) );
  OR2_X1 U13183 ( .A1(n10012), .A2(n14989), .ZN(n10573) );
  INV_X1 U13184 ( .A(P3_REG1_REG_10__SCAN_IN), .ZN(n10958) );
  OR2_X1 U13185 ( .A1(n11436), .A2(n10958), .ZN(n10572) );
  XNOR2_X1 U13186 ( .A(n11057), .B(n12342), .ZN(n10578) );
  NAND2_X1 U13187 ( .A1(n10576), .A2(n11472), .ZN(n10579) );
  NAND2_X1 U13188 ( .A1(n10717), .A2(n11060), .ZN(n10577) );
  NAND2_X1 U13189 ( .A1(n10577), .A2(n12318), .ZN(n10595) );
  AOI21_X1 U13190 ( .B1(n10717), .B2(n10579), .A(n10578), .ZN(n10594) );
  NAND2_X1 U13191 ( .A1(n10580), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n10581) );
  AND2_X1 U13192 ( .A1(n11055), .A2(n10581), .ZN(n15394) );
  INV_X1 U13193 ( .A(P3_REG1_REG_11__SCAN_IN), .ZN(n10582) );
  OR2_X1 U13194 ( .A1(n11436), .A2(n10582), .ZN(n10583) );
  OAI21_X1 U13195 ( .B1(n10012), .B2(n15394), .A(n10583), .ZN(n10588) );
  INV_X1 U13196 ( .A(P3_REG2_REG_11__SCAN_IN), .ZN(n10584) );
  INV_X1 U13197 ( .A(P3_REG0_REG_11__SCAN_IN), .ZN(n10585) );
  NOR2_X1 U13198 ( .A1(n11438), .A2(n10585), .ZN(n10586) );
  INV_X1 U13199 ( .A(n14984), .ZN(n11478) );
  NAND2_X1 U13200 ( .A1(n12332), .A2(n14985), .ZN(n10590) );
  INV_X1 U13201 ( .A(P3_REG3_REG_10__SCAN_IN), .ZN(n15199) );
  NOR2_X1 U13202 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n15199), .ZN(n14968) );
  INV_X1 U13203 ( .A(n14968), .ZN(n10589) );
  OAI211_X1 U13204 ( .C1(n11478), .C2(n12336), .A(n10590), .B(n10589), .ZN(
        n10592) );
  NOR2_X1 U13205 ( .A1(n15395), .A2(n14989), .ZN(n10591) );
  AOI211_X1 U13206 ( .C1(n15399), .C2(n14988), .A(n10592), .B(n10591), .ZN(
        n10593) );
  OAI21_X1 U13207 ( .B1(n10595), .B2(n10594), .A(n10593), .ZN(P3_U3157) );
  INV_X1 U13208 ( .A(n10600), .ZN(n10615) );
  NAND2_X1 U13209 ( .A1(n10600), .A2(n13640), .ZN(n10597) );
  NAND2_X1 U13210 ( .A1(n13766), .A2(n6536), .ZN(n10596) );
  NAND2_X1 U13211 ( .A1(n10597), .A2(n10596), .ZN(n10598) );
  XNOR2_X1 U13212 ( .A(n10598), .B(n13637), .ZN(n10670) );
  AND2_X1 U13213 ( .A1(n13766), .A2(n13603), .ZN(n10599) );
  AOI21_X1 U13214 ( .B1(n10600), .B2(n6536), .A(n10599), .ZN(n10671) );
  XNOR2_X1 U13215 ( .A(n10670), .B(n10671), .ZN(n10607) );
  INV_X1 U13216 ( .A(n10601), .ZN(n10602) );
  NAND2_X1 U13217 ( .A1(n10603), .A2(n10602), .ZN(n10604) );
  AND2_X2 U13218 ( .A1(n10605), .A2(n10604), .ZN(n10606) );
  OAI21_X1 U13219 ( .B1(n10607), .B2(n10606), .A(n10674), .ZN(n10608) );
  NAND2_X1 U13220 ( .A1(n10608), .A2(n14395), .ZN(n10614) );
  OAI22_X1 U13221 ( .A1(n13738), .A2(n10610), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n10609), .ZN(n10611) );
  AOI21_X1 U13222 ( .B1(n10612), .B2(n13740), .A(n10611), .ZN(n10613) );
  OAI211_X1 U13223 ( .C1(n10615), .C2(n13743), .A(n10614), .B(n10613), .ZN(
        P1_U3221) );
  INV_X1 U13224 ( .A(n10616), .ZN(n10619) );
  INV_X1 U13225 ( .A(n10617), .ZN(n10618) );
  NAND2_X1 U13226 ( .A1(n10619), .A2(n10618), .ZN(n10620) );
  XNOR2_X1 U13227 ( .A(n12021), .B(n6528), .ZN(n10841) );
  NAND2_X1 U13228 ( .A1(n13040), .A2(n13326), .ZN(n10843) );
  XNOR2_X1 U13229 ( .A(n10841), .B(n10843), .ZN(n10623) );
  XNOR2_X1 U13230 ( .A(n10840), .B(n10623), .ZN(n10630) );
  NOR2_X1 U13231 ( .A1(n14348), .A2(n10648), .ZN(n10628) );
  NAND2_X1 U13232 ( .A1(n13041), .A2(n14334), .ZN(n10625) );
  NAND2_X1 U13233 ( .A1(n13039), .A2(n14336), .ZN(n10624) );
  AND2_X1 U13234 ( .A1(n10625), .A2(n10624), .ZN(n10645) );
  OAI22_X1 U13235 ( .A1(n14343), .A2(n10645), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10626), .ZN(n10627) );
  AOI211_X1 U13236 ( .C1(n12021), .C2(n13019), .A(n10628), .B(n10627), .ZN(
        n10629) );
  OAI21_X1 U13237 ( .B1(n10630), .B2(n14342), .A(n10629), .ZN(P2_U3208) );
  INV_X1 U13238 ( .A(n12725), .ZN(n14310) );
  OAI21_X1 U13239 ( .B1(n10632), .B2(n11830), .A(n10631), .ZN(n15074) );
  NAND2_X1 U13240 ( .A1(n10633), .A2(n15049), .ZN(n15071) );
  OAI22_X1 U13241 ( .A1(n12535), .A2(n15071), .B1(n10634), .B2(n15020), .ZN(
        n10642) );
  OAI211_X1 U13242 ( .C1(n10637), .C2(n10636), .A(n10635), .B(n15046), .ZN(
        n10640) );
  OR2_X1 U13243 ( .A1(n10638), .A2(n15031), .ZN(n10639) );
  OAI211_X1 U13244 ( .C1(n15030), .C2(n15029), .A(n10640), .B(n10639), .ZN(
        n15072) );
  MUX2_X1 U13245 ( .A(n15072), .B(P3_REG2_REG_4__SCAN_IN), .S(n15052), .Z(
        n10641) );
  AOI211_X1 U13246 ( .C1(n14310), .C2(n15074), .A(n10642), .B(n10641), .ZN(
        n10643) );
  INV_X1 U13247 ( .A(n10643), .ZN(P3_U3229) );
  XOR2_X1 U13248 ( .A(n12206), .B(n10644), .Z(n10646) );
  OAI21_X1 U13249 ( .B1(n10646), .B2(n14351), .A(n10645), .ZN(n10779) );
  INV_X1 U13250 ( .A(n10779), .ZN(n10655) );
  INV_X1 U13251 ( .A(n10772), .ZN(n10647) );
  AOI211_X1 U13252 ( .C1(n12021), .C2(n6817), .A(n9445), .B(n10647), .ZN(
        n10780) );
  NOR2_X1 U13253 ( .A1(n10782), .A2(n13311), .ZN(n10651) );
  OAI22_X1 U13254 ( .A1(n13281), .A2(n10649), .B1(n10648), .B2(n13323), .ZN(
        n10650) );
  AOI211_X1 U13255 ( .C1(n10780), .C2(n14362), .A(n10651), .B(n10650), .ZN(
        n10654) );
  XOR2_X1 U13256 ( .A(n10652), .B(n12206), .Z(n10781) );
  NAND2_X1 U13257 ( .A1(n10781), .A2(n14363), .ZN(n10653) );
  OAI211_X1 U13258 ( .C1(n10655), .C2(n14367), .A(n10654), .B(n10653), .ZN(
        P2_U3254) );
  INV_X1 U13259 ( .A(n10656), .ZN(n11908) );
  OAI222_X1 U13260 ( .A1(P1_U3086), .A2(n13847), .B1(n6535), .B2(n11908), .C1(
        n10657), .C2(n14266), .ZN(P1_U3336) );
  NAND2_X1 U13261 ( .A1(n10659), .A2(n10658), .ZN(n10795) );
  XNOR2_X1 U13262 ( .A(n10795), .B(n10660), .ZN(n10666) );
  NAND2_X1 U13263 ( .A1(n15389), .A2(n12343), .ZN(n10662) );
  INV_X1 U13264 ( .A(P3_REG3_REG_7__SCAN_IN), .ZN(n15275) );
  NOR2_X1 U13265 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n15275), .ZN(n14913) );
  INV_X1 U13266 ( .A(n14913), .ZN(n10661) );
  OAI211_X1 U13267 ( .C1(n10708), .C2(n15392), .A(n10662), .B(n10661), .ZN(
        n10664) );
  NOR2_X1 U13268 ( .A1(n15395), .A2(n15006), .ZN(n10663) );
  AOI211_X1 U13269 ( .C1(n15399), .C2(n15004), .A(n10664), .B(n10663), .ZN(
        n10665) );
  OAI21_X1 U13270 ( .B1(n10666), .B2(n15401), .A(n10665), .ZN(P3_U3153) );
  INV_X1 U13271 ( .A(n10667), .ZN(n11910) );
  OAI222_X1 U13272 ( .A1(P1_U3086), .A2(n10669), .B1(n6535), .B2(n11910), .C1(
        n10668), .C2(n14266), .ZN(P1_U3334) );
  INV_X1 U13273 ( .A(n10670), .ZN(n10672) );
  NAND2_X1 U13274 ( .A1(n10672), .A2(n10671), .ZN(n10673) );
  NAND2_X1 U13275 ( .A1(n14500), .A2(n13640), .ZN(n10676) );
  NAND2_X1 U13276 ( .A1(n13765), .A2(n6536), .ZN(n10675) );
  NAND2_X1 U13277 ( .A1(n10676), .A2(n10675), .ZN(n10677) );
  XNOR2_X1 U13278 ( .A(n10677), .B(n13591), .ZN(n10823) );
  AND2_X1 U13279 ( .A1(n13765), .A2(n13636), .ZN(n10678) );
  AOI21_X1 U13280 ( .B1(n14500), .B2(n6536), .A(n10678), .ZN(n10824) );
  XNOR2_X1 U13281 ( .A(n10823), .B(n10824), .ZN(n10679) );
  XNOR2_X1 U13282 ( .A(n10828), .B(n10679), .ZN(n10686) );
  NAND2_X1 U13283 ( .A1(n13766), .A2(n14107), .ZN(n10681) );
  NAND2_X1 U13284 ( .A1(n13764), .A2(n14108), .ZN(n10680) );
  NAND2_X1 U13285 ( .A1(n10681), .A2(n10680), .ZN(n14495) );
  NAND2_X1 U13286 ( .A1(n14397), .A2(n14495), .ZN(n10682) );
  OAI211_X1 U13287 ( .C1(n14401), .C2(n14498), .A(n10683), .B(n10682), .ZN(
        n10684) );
  AOI21_X1 U13288 ( .B1(n14500), .B2(n14398), .A(n10684), .ZN(n10685) );
  OAI21_X1 U13289 ( .B1(n10686), .B2(n13756), .A(n10685), .ZN(P1_U3231) );
  INV_X1 U13290 ( .A(n10687), .ZN(n10689) );
  AOI21_X1 U13291 ( .B1(n10689), .B2(n10695), .A(n10688), .ZN(n10691) );
  XOR2_X1 U13292 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n11194), .Z(n10690) );
  OAI211_X1 U13293 ( .C1(n10691), .C2(n10690), .A(n14483), .B(n11192), .ZN(
        n10702) );
  NAND2_X1 U13294 ( .A1(P1_U3086), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n13683)
         );
  INV_X1 U13295 ( .A(n10692), .ZN(n10694) );
  AOI21_X1 U13296 ( .B1(n10695), .B2(n10694), .A(n10693), .ZN(n10698) );
  INV_X1 U13297 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n11186) );
  NOR2_X1 U13298 ( .A1(n11186), .A2(n11187), .ZN(n10696) );
  AOI21_X1 U13299 ( .B1(n11186), .B2(n11187), .A(n10696), .ZN(n10697) );
  NAND2_X1 U13300 ( .A1(n10697), .A2(n10698), .ZN(n11185) );
  OAI211_X1 U13301 ( .C1(n10698), .C2(n10697), .A(n14478), .B(n11185), .ZN(
        n10699) );
  NAND2_X1 U13302 ( .A1(n13683), .A2(n10699), .ZN(n10700) );
  AOI21_X1 U13303 ( .B1(n14472), .B2(P1_ADDR_REG_16__SCAN_IN), .A(n10700), 
        .ZN(n10701) );
  OAI211_X1 U13304 ( .C1(n13832), .C2(n11187), .A(n10702), .B(n10701), .ZN(
        P1_U3259) );
  XNOR2_X1 U13305 ( .A(n10703), .B(n11826), .ZN(n15077) );
  INV_X1 U13306 ( .A(n15077), .ZN(n10716) );
  INV_X1 U13307 ( .A(n10704), .ZN(n10705) );
  AOI21_X1 U13308 ( .B1(n11826), .B2(n10706), .A(n10705), .ZN(n10707) );
  OAI222_X1 U13309 ( .A1(n15029), .A2(n10709), .B1(n15031), .B2(n10708), .C1(
        n15027), .C2(n10707), .ZN(n15075) );
  NOR2_X1 U13310 ( .A1(n15057), .A2(n10928), .ZN(n10714) );
  AND2_X1 U13311 ( .A1(n10710), .A2(n15049), .ZN(n15076) );
  INV_X1 U13312 ( .A(n15076), .ZN(n10712) );
  OAI22_X1 U13313 ( .A1(n12535), .A2(n10712), .B1(n10711), .B2(n15020), .ZN(
        n10713) );
  AOI211_X1 U13314 ( .C1(n15075), .C2(n15057), .A(n10714), .B(n10713), .ZN(
        n10715) );
  OAI21_X1 U13315 ( .B1(n12725), .B2(n10716), .A(n10715), .ZN(P3_U3228) );
  INV_X1 U13316 ( .A(n10717), .ZN(n10718) );
  AOI21_X1 U13317 ( .B1(n11059), .B2(n11066), .A(n10718), .ZN(n10724) );
  NAND2_X1 U13318 ( .A1(n12332), .A2(n12343), .ZN(n10720) );
  NOR2_X1 U13319 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n10557), .ZN(n14948) );
  INV_X1 U13320 ( .A(n14948), .ZN(n10719) );
  OAI211_X1 U13321 ( .C1(n15393), .C2(n12336), .A(n10720), .B(n10719), .ZN(
        n10722) );
  NOR2_X1 U13322 ( .A1(n15395), .A2(n11107), .ZN(n10721) );
  AOI211_X1 U13323 ( .C1(n15399), .C2(n11730), .A(n10722), .B(n10721), .ZN(
        n10723) );
  OAI21_X1 U13324 ( .B1(n10724), .B2(n15401), .A(n10723), .ZN(P3_U3171) );
  INV_X1 U13325 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n10746) );
  OR2_X1 U13326 ( .A1(n10725), .A2(n10736), .ZN(n10727) );
  NAND2_X1 U13327 ( .A1(n10727), .A2(n10726), .ZN(n10728) );
  NAND2_X1 U13328 ( .A1(n14753), .A2(n10728), .ZN(n10729) );
  XNOR2_X1 U13329 ( .A(n10737), .B(n10728), .ZN(n14757) );
  NAND2_X1 U13330 ( .A1(P2_REG2_REG_15__SCAN_IN), .A2(n14757), .ZN(n14755) );
  NAND2_X1 U13331 ( .A1(n10729), .A2(n14755), .ZN(n10733) );
  NAND2_X1 U13332 ( .A1(n10743), .A2(n11409), .ZN(n10730) );
  OAI21_X1 U13333 ( .B1(n10743), .B2(n11409), .A(n10730), .ZN(n10732) );
  NAND2_X1 U13334 ( .A1(n11363), .A2(n11409), .ZN(n10731) );
  OAI211_X1 U13335 ( .C1(n11409), .C2(n11363), .A(n10733), .B(n10731), .ZN(
        n11355) );
  OAI211_X1 U13336 ( .C1(n10733), .C2(n10732), .A(n11355), .B(n14756), .ZN(
        n10745) );
  NAND2_X1 U13337 ( .A1(P2_U3088), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n11382)
         );
  INV_X1 U13338 ( .A(n10734), .ZN(n10735) );
  OAI21_X1 U13339 ( .B1(n14372), .B2(n10736), .A(n10735), .ZN(n10738) );
  NAND2_X1 U13340 ( .A1(n14753), .A2(n10738), .ZN(n10739) );
  XNOR2_X1 U13341 ( .A(n10738), .B(n10737), .ZN(n14760) );
  NAND2_X1 U13342 ( .A1(P2_REG1_REG_15__SCAN_IN), .A2(n14760), .ZN(n14758) );
  NAND2_X1 U13343 ( .A1(n10739), .A2(n14758), .ZN(n11362) );
  XNOR2_X1 U13344 ( .A(n10743), .B(P2_REG1_REG_16__SCAN_IN), .ZN(n11364) );
  XNOR2_X1 U13345 ( .A(n11362), .B(n11364), .ZN(n10740) );
  NAND2_X1 U13346 ( .A1(n14759), .A2(n10740), .ZN(n10741) );
  NAND2_X1 U13347 ( .A1(n11382), .A2(n10741), .ZN(n10742) );
  AOI21_X1 U13348 ( .B1(n14754), .B2(n10743), .A(n10742), .ZN(n10744) );
  OAI211_X1 U13349 ( .C1(n14736), .C2(n10746), .A(n10745), .B(n10744), .ZN(
        P2_U3230) );
  AND2_X1 U13350 ( .A1(n11709), .A2(n11710), .ZN(n10747) );
  INV_X1 U13351 ( .A(n11710), .ZN(n11718) );
  INV_X1 U13352 ( .A(n10752), .ZN(n11827) );
  INV_X1 U13353 ( .A(n11043), .ZN(n10749) );
  AOI21_X1 U13354 ( .B1(n6700), .B2(n10752), .A(n10749), .ZN(n15001) );
  NAND2_X1 U13355 ( .A1(n12345), .A2(n15013), .ZN(n10750) );
  NAND2_X1 U13356 ( .A1(n10751), .A2(n10750), .ZN(n10753) );
  OAI211_X1 U13357 ( .C1(n10753), .C2(n10752), .A(n11046), .B(n15046), .ZN(
        n10755) );
  AOI22_X1 U13358 ( .A1(n12345), .A2(n15041), .B1(n15038), .B2(n12343), .ZN(
        n10754) );
  AND2_X1 U13359 ( .A1(n10755), .A2(n10754), .ZN(n15000) );
  OAI21_X1 U13360 ( .B1(n15001), .B2(n12748), .A(n15000), .ZN(n10761) );
  INV_X1 U13361 ( .A(n10761), .ZN(n10757) );
  AOI22_X1 U13362 ( .A1(n12782), .A2(n15004), .B1(n15094), .B2(
        P3_REG1_REG_7__SCAN_IN), .ZN(n10756) );
  OAI21_X1 U13363 ( .B1(n10757), .B2(n15094), .A(n10756), .ZN(P3_U3466) );
  INV_X1 U13364 ( .A(P3_REG0_REG_7__SCAN_IN), .ZN(n10758) );
  OAI22_X1 U13365 ( .A1(n10759), .A2(n12867), .B1(n15085), .B2(n10758), .ZN(
        n10760) );
  AOI21_X1 U13366 ( .B1(n10761), .B2(n15085), .A(n10760), .ZN(n10762) );
  INV_X1 U13367 ( .A(n10762), .ZN(P3_U3411) );
  INV_X1 U13368 ( .A(n12207), .ZN(n10763) );
  XNOR2_X1 U13369 ( .A(n10764), .B(n10763), .ZN(n14383) );
  NAND2_X1 U13370 ( .A1(n14383), .A2(n13307), .ZN(n10771) );
  AOI21_X1 U13371 ( .B1(n10765), .B2(n12207), .A(n14351), .ZN(n10769) );
  NAND2_X1 U13372 ( .A1(n13040), .A2(n14334), .ZN(n10767) );
  NAND2_X1 U13373 ( .A1(n14335), .A2(n14336), .ZN(n10766) );
  NAND2_X1 U13374 ( .A1(n10767), .A2(n10766), .ZN(n10850) );
  AOI21_X1 U13375 ( .B1(n10769), .B2(n10768), .A(n10850), .ZN(n10770) );
  AOI21_X1 U13376 ( .B1(n10772), .B2(n14379), .A(n9445), .ZN(n10773) );
  NAND2_X1 U13377 ( .A1(n10773), .A2(n10989), .ZN(n14381) );
  OAI22_X1 U13378 ( .A1(n13281), .A2(n10774), .B1(n10852), .B2(n13323), .ZN(
        n10775) );
  AOI21_X1 U13379 ( .B1(n14379), .B2(n14355), .A(n10775), .ZN(n10776) );
  OAI21_X1 U13380 ( .B1(n14381), .B2(n13330), .A(n10776), .ZN(n10777) );
  AOI21_X1 U13381 ( .B1(n14383), .B2(n13317), .A(n10777), .ZN(n10778) );
  OAI21_X1 U13382 ( .B1(n14385), .B2(n14367), .A(n10778), .ZN(P2_U3253) );
  AOI211_X1 U13383 ( .C1(n14378), .C2(n10781), .A(n10780), .B(n10779), .ZN(
        n10786) );
  OAI22_X1 U13384 ( .A1(n10782), .A2(n13468), .B1(n14821), .B2(n7774), .ZN(
        n10783) );
  INV_X1 U13385 ( .A(n10783), .ZN(n10784) );
  OAI21_X1 U13386 ( .B1(n10786), .B2(n14819), .A(n10784), .ZN(P2_U3463) );
  AOI22_X1 U13387 ( .A1(n12021), .A2(n13398), .B1(n14827), .B2(
        P2_REG1_REG_11__SCAN_IN), .ZN(n10785) );
  OAI21_X1 U13388 ( .B1(n10786), .B2(n14827), .A(n10785), .ZN(P2_U3510) );
  NAND2_X1 U13389 ( .A1(n11013), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n10789) );
  XNOR2_X1 U13390 ( .A(n10881), .B(n7368), .ZN(n11529) );
  INV_X1 U13391 ( .A(n11529), .ZN(n10792) );
  INV_X1 U13392 ( .A(SI_24_), .ZN(n11530) );
  OAI222_X1 U13393 ( .A1(P3_U3151), .A2(n10793), .B1(n12245), .B2(n10792), 
        .C1(n11530), .C2(n11338), .ZN(P3_U3271) );
  MUX2_X1 U13394 ( .A(n10795), .B(n12344), .S(n10794), .Z(n10797) );
  XNOR2_X1 U13395 ( .A(n10797), .B(n10796), .ZN(n10805) );
  NAND2_X1 U13396 ( .A1(n12332), .A2(n12344), .ZN(n10800) );
  NOR2_X1 U13397 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n10798), .ZN(n14930) );
  INV_X1 U13398 ( .A(n14930), .ZN(n10799) );
  OAI211_X1 U13399 ( .C1(n11472), .C2(n12336), .A(n10800), .B(n10799), .ZN(
        n10803) );
  NOR2_X1 U13400 ( .A1(n15395), .A2(n10801), .ZN(n10802) );
  AOI211_X1 U13401 ( .C1(n15399), .C2(n14996), .A(n10803), .B(n10802), .ZN(
        n10804) );
  OAI21_X1 U13402 ( .B1(n10805), .B2(n15401), .A(n10804), .ZN(P3_U3161) );
  INV_X1 U13403 ( .A(n13764), .ZN(n11030) );
  OR2_X1 U13404 ( .A1(n14635), .A2(n11030), .ZN(n10806) );
  XNOR2_X1 U13405 ( .A(n10856), .B(n10814), .ZN(n10808) );
  OAI222_X1 U13406 ( .A1(n14581), .A2(n10809), .B1(n10808), .B2(n14560), .C1(
        n14561), .C2(n11030), .ZN(n14412) );
  INV_X1 U13407 ( .A(n14412), .ZN(n10822) );
  NAND2_X1 U13408 ( .A1(n10811), .A2(n10810), .ZN(n10813) );
  OR2_X1 U13409 ( .A1(n14635), .A2(n13764), .ZN(n10812) );
  INV_X1 U13410 ( .A(n10814), .ZN(n10815) );
  XNOR2_X1 U13411 ( .A(n10870), .B(n10815), .ZN(n14414) );
  INV_X1 U13412 ( .A(n11018), .ZN(n14411) );
  NAND2_X1 U13413 ( .A1(n14411), .A2(n10816), .ZN(n10863) );
  OAI211_X1 U13414 ( .C1(n14411), .C2(n10816), .A(n14546), .B(n10863), .ZN(
        n14410) );
  OAI22_X1 U13415 ( .A1(n14543), .A2(n10817), .B1(n11027), .B2(n14542), .ZN(
        n10818) );
  AOI21_X1 U13416 ( .B1(n11018), .B2(n14566), .A(n10818), .ZN(n10819) );
  OAI21_X1 U13417 ( .B1(n14410), .B2(n13959), .A(n10819), .ZN(n10820) );
  AOI21_X1 U13418 ( .B1(n14414), .B2(n14083), .A(n10820), .ZN(n10821) );
  OAI21_X1 U13419 ( .B1(n10822), .B2(n6531), .A(n10821), .ZN(P1_U3282) );
  AND2_X1 U13420 ( .A1(n10823), .A2(n10824), .ZN(n10827) );
  INV_X1 U13421 ( .A(n10823), .ZN(n10826) );
  INV_X1 U13422 ( .A(n10824), .ZN(n10825) );
  NAND2_X1 U13423 ( .A1(n14635), .A2(n13640), .ZN(n10830) );
  NAND2_X1 U13424 ( .A1(n13764), .A2(n6536), .ZN(n10829) );
  NAND2_X1 U13425 ( .A1(n10830), .A2(n10829), .ZN(n10831) );
  XNOR2_X1 U13426 ( .A(n10831), .B(n13637), .ZN(n11021) );
  AND2_X1 U13427 ( .A1(n13764), .A2(n13636), .ZN(n10832) );
  AOI21_X1 U13428 ( .B1(n14635), .B2(n6536), .A(n10832), .ZN(n11019) );
  XNOR2_X1 U13429 ( .A(n11021), .B(n11019), .ZN(n11022) );
  XNOR2_X1 U13430 ( .A(n11023), .B(n11022), .ZN(n10839) );
  INV_X1 U13431 ( .A(n13763), .ZN(n10857) );
  NOR2_X1 U13432 ( .A1(n13748), .A2(n10857), .ZN(n10833) );
  AOI211_X1 U13433 ( .C1(n13750), .C2(n13765), .A(n10834), .B(n10833), .ZN(
        n10835) );
  OAI21_X1 U13434 ( .B1(n10836), .B2(n14401), .A(n10835), .ZN(n10837) );
  AOI21_X1 U13435 ( .B1(n14635), .B2(n14398), .A(n10837), .ZN(n10838) );
  OAI21_X1 U13436 ( .B1(n10839), .B2(n13756), .A(n10838), .ZN(P1_U3217) );
  INV_X1 U13437 ( .A(n10841), .ZN(n10842) );
  XNOR2_X1 U13438 ( .A(n14379), .B(n6528), .ZN(n10847) );
  INV_X1 U13439 ( .A(n10847), .ZN(n10845) );
  AND2_X1 U13440 ( .A1(n13039), .A2(n13326), .ZN(n10846) );
  INV_X1 U13441 ( .A(n10846), .ZN(n10844) );
  NAND2_X1 U13442 ( .A1(n10845), .A2(n10844), .ZN(n10975) );
  INV_X1 U13443 ( .A(n10975), .ZN(n10848) );
  AND2_X1 U13444 ( .A1(n10847), .A2(n10846), .ZN(n10974) );
  NOR2_X1 U13445 ( .A1(n10848), .A2(n10974), .ZN(n10849) );
  XNOR2_X1 U13446 ( .A(n10976), .B(n10849), .ZN(n10855) );
  NAND2_X1 U13447 ( .A1(n13016), .A2(n10850), .ZN(n10851) );
  NAND2_X1 U13448 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(P2_U3088), .ZN(n14734)
         );
  OAI211_X1 U13449 ( .C1(n14348), .C2(n10852), .A(n10851), .B(n14734), .ZN(
        n10853) );
  AOI21_X1 U13450 ( .B1(n14379), .B2(n13019), .A(n10853), .ZN(n10854) );
  OAI21_X1 U13451 ( .B1(n10855), .B2(n14342), .A(n10854), .ZN(P2_U3196) );
  AOI21_X1 U13452 ( .B1(n7277), .B2(n10858), .A(n14560), .ZN(n10862) );
  NAND2_X1 U13453 ( .A1(n10859), .A2(n10874), .ZN(n11150) );
  NAND2_X1 U13454 ( .A1(n13763), .A2(n14107), .ZN(n10861) );
  NAND2_X1 U13455 ( .A1(n13761), .A2(n14108), .ZN(n10860) );
  NAND2_X1 U13456 ( .A1(n10861), .A2(n10860), .ZN(n13658) );
  AOI21_X1 U13457 ( .B1(n10862), .B2(n11150), .A(n13658), .ZN(n11037) );
  AOI211_X1 U13458 ( .C1(n13667), .C2(n10863), .A(n14572), .B(n6972), .ZN(
        n11035) );
  INV_X1 U13459 ( .A(n13667), .ZN(n10864) );
  NOR2_X1 U13460 ( .A1(n10864), .A2(n14119), .ZN(n10867) );
  OAI22_X1 U13461 ( .A1(n14543), .A2(n10865), .B1(n13660), .B2(n14542), .ZN(
        n10866) );
  AOI211_X1 U13462 ( .C1(n11035), .C2(n14574), .A(n10867), .B(n10866), .ZN(
        n10877) );
  INV_X1 U13463 ( .A(n10868), .ZN(n10869) );
  INV_X1 U13464 ( .A(n11146), .ZN(n10872) );
  AOI21_X1 U13465 ( .B1(n10874), .B2(n10873), .A(n10872), .ZN(n11038) );
  INV_X1 U13466 ( .A(n11038), .ZN(n10875) );
  NAND2_X1 U13467 ( .A1(n10875), .A2(n14083), .ZN(n10876) );
  OAI211_X1 U13468 ( .C1(n11037), .C2(n6531), .A(n10877), .B(n10876), .ZN(
        P1_U3281) );
  INV_X1 U13469 ( .A(n10878), .ZN(n10879) );
  OAI222_X1 U13470 ( .A1(n11904), .A2(n10880), .B1(n6534), .B2(n10879), .C1(
        n11925), .C2(P2_U3088), .ZN(P2_U3305) );
  NAND2_X1 U13471 ( .A1(n15297), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n10999) );
  NAND2_X1 U13472 ( .A1(n15170), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n10882) );
  AND2_X1 U13473 ( .A1(n10999), .A2(n10882), .ZN(n10883) );
  OR2_X1 U13474 ( .A1(n10884), .A2(n10883), .ZN(n10885) );
  AND2_X1 U13475 ( .A1(n11000), .A2(n10885), .ZN(n11539) );
  INV_X1 U13476 ( .A(n11539), .ZN(n10887) );
  OAI222_X1 U13477 ( .A1(n12245), .A2(n10887), .B1(n11338), .B2(n11540), .C1(
        P3_U3151), .C2(n10886), .ZN(P3_U3270) );
  NAND2_X1 U13478 ( .A1(n10899), .A2(P3_REG2_REG_2__SCAN_IN), .ZN(n10888) );
  XNOR2_X1 U13479 ( .A(n14857), .B(P3_REG2_REG_4__SCAN_IN), .ZN(n14850) );
  NOR2_X1 U13480 ( .A1(n14851), .A2(n14850), .ZN(n14849) );
  NAND2_X1 U13481 ( .A1(n14893), .A2(P3_REG2_REG_6__SCAN_IN), .ZN(n10892) );
  OR2_X1 U13482 ( .A1(n14893), .A2(P3_REG2_REG_6__SCAN_IN), .ZN(n10891) );
  NAND2_X1 U13483 ( .A1(n10892), .A2(n10891), .ZN(n14886) );
  NOR2_X1 U13484 ( .A1(n10941), .A2(n10893), .ZN(n10894) );
  MUX2_X1 U13485 ( .A(n10946), .B(P3_REG2_REG_8__SCAN_IN), .S(n14928), .Z(
        n14921) );
  NOR2_X1 U13486 ( .A1(n10954), .A2(n10895), .ZN(n10896) );
  NOR2_X1 U13487 ( .A1(n10953), .A2(n14939), .ZN(n14938) );
  INV_X1 U13488 ( .A(P3_REG2_REG_10__SCAN_IN), .ZN(n10959) );
  MUX2_X1 U13489 ( .A(n10959), .B(P3_REG2_REG_10__SCAN_IN), .S(n14965), .Z(
        n14956) );
  NOR2_X1 U13490 ( .A1(n10584), .A2(n10897), .ZN(n11120) );
  AOI21_X1 U13491 ( .B1(n10584), .B2(n10897), .A(n11120), .ZN(n10973) );
  INV_X1 U13492 ( .A(n14965), .ZN(n10960) );
  INV_X1 U13493 ( .A(n14928), .ZN(n10947) );
  NAND2_X1 U13494 ( .A1(n14893), .A2(P3_REG1_REG_6__SCAN_IN), .ZN(n10905) );
  MUX2_X1 U13495 ( .A(P3_REG1_REG_6__SCAN_IN), .B(n10932), .S(n14893), .Z(
        n14897) );
  NAND2_X1 U13496 ( .A1(n14857), .A2(P3_REG1_REG_4__SCAN_IN), .ZN(n10902) );
  MUX2_X1 U13497 ( .A(P3_REG1_REG_4__SCAN_IN), .B(n10920), .S(n14857), .Z(
        n14861) );
  AOI21_X1 U13498 ( .B1(n10899), .B2(P3_REG1_REG_2__SCAN_IN), .A(n10898), .ZN(
        n10900) );
  XNOR2_X1 U13499 ( .A(n10900), .B(n10917), .ZN(n14844) );
  INV_X1 U13500 ( .A(n14844), .ZN(n10901) );
  OAI22_X1 U13501 ( .A1(n10901), .A2(n10914), .B1(n14842), .B2(n10900), .ZN(
        n14862) );
  NAND2_X1 U13502 ( .A1(n14861), .A2(n14862), .ZN(n14860) );
  NAND2_X1 U13503 ( .A1(n10902), .A2(n14860), .ZN(n10903) );
  NAND2_X1 U13504 ( .A1(n14875), .A2(n10903), .ZN(n10904) );
  XNOR2_X1 U13505 ( .A(n10903), .B(n7024), .ZN(n14879) );
  NAND2_X1 U13506 ( .A1(P3_REG1_REG_5__SCAN_IN), .A2(n14879), .ZN(n14878) );
  NAND2_X1 U13507 ( .A1(n14911), .A2(n10906), .ZN(n10907) );
  NAND2_X1 U13508 ( .A1(P3_REG1_REG_7__SCAN_IN), .A2(n14915), .ZN(n14914) );
  MUX2_X1 U13509 ( .A(P3_REG1_REG_8__SCAN_IN), .B(n10945), .S(n14928), .Z(
        n14932) );
  NAND2_X1 U13510 ( .A1(n14946), .A2(n10908), .ZN(n10909) );
  NAND2_X1 U13511 ( .A1(P3_REG1_REG_9__SCAN_IN), .A2(n14950), .ZN(n14949) );
  MUX2_X1 U13512 ( .A(P3_REG1_REG_10__SCAN_IN), .B(n10958), .S(n14965), .Z(
        n14971) );
  NAND2_X1 U13513 ( .A1(P3_REG1_REG_11__SCAN_IN), .A2(n10910), .ZN(n11127) );
  OAI21_X1 U13514 ( .B1(P3_REG1_REG_11__SCAN_IN), .B2(n10910), .A(n11127), 
        .ZN(n10971) );
  INV_X1 U13515 ( .A(n14966), .ZN(n14843) );
  NAND2_X1 U13516 ( .A1(n14843), .A2(n6890), .ZN(n10911) );
  NAND2_X1 U13517 ( .A1(P3_U3151), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n15390)
         );
  OAI211_X1 U13518 ( .C1(n10912), .C2(n14834), .A(n10911), .B(n15390), .ZN(
        n10970) );
  INV_X1 U13519 ( .A(n10913), .ZN(n14836) );
  MUX2_X1 U13520 ( .A(n10915), .B(n10914), .S(n12463), .Z(n10916) );
  NAND2_X1 U13521 ( .A1(n10916), .A2(n14842), .ZN(n14853) );
  INV_X1 U13522 ( .A(n10916), .ZN(n10918) );
  NAND2_X1 U13523 ( .A1(n10918), .A2(n10917), .ZN(n10919) );
  AND2_X1 U13524 ( .A1(n14853), .A2(n10919), .ZN(n14835) );
  OAI21_X1 U13525 ( .B1(n14837), .B2(n14836), .A(n14835), .ZN(n14854) );
  INV_X1 U13526 ( .A(P3_REG2_REG_4__SCAN_IN), .ZN(n10921) );
  MUX2_X1 U13527 ( .A(n10921), .B(n10920), .S(n12463), .Z(n10923) );
  NAND2_X1 U13528 ( .A1(n10923), .A2(n10922), .ZN(n10926) );
  INV_X1 U13529 ( .A(n10923), .ZN(n10924) );
  NAND2_X1 U13530 ( .A1(n10924), .A2(n14857), .ZN(n10925) );
  NAND2_X1 U13531 ( .A1(n10926), .A2(n10925), .ZN(n14852) );
  AOI21_X1 U13532 ( .B1(n14854), .B2(n14853), .A(n14852), .ZN(n14871) );
  INV_X1 U13533 ( .A(n10926), .ZN(n14870) );
  MUX2_X1 U13534 ( .A(n10928), .B(n10927), .S(n12463), .Z(n10929) );
  NAND2_X1 U13535 ( .A1(n10929), .A2(n7024), .ZN(n14889) );
  INV_X1 U13536 ( .A(n10929), .ZN(n10930) );
  NAND2_X1 U13537 ( .A1(n10930), .A2(n14875), .ZN(n10931) );
  AND2_X1 U13538 ( .A1(n14889), .A2(n10931), .ZN(n14869) );
  OAI21_X1 U13539 ( .B1(n14871), .B2(n14870), .A(n14869), .ZN(n14890) );
  MUX2_X1 U13540 ( .A(n10933), .B(n10932), .S(n12463), .Z(n10935) );
  INV_X1 U13541 ( .A(n14893), .ZN(n10934) );
  NAND2_X1 U13542 ( .A1(n10935), .A2(n10934), .ZN(n10938) );
  INV_X1 U13543 ( .A(n10935), .ZN(n10936) );
  NAND2_X1 U13544 ( .A1(n10936), .A2(n14893), .ZN(n10937) );
  NAND2_X1 U13545 ( .A1(n10938), .A2(n10937), .ZN(n14888) );
  AOI21_X1 U13546 ( .B1(n14890), .B2(n14889), .A(n14888), .ZN(n14907) );
  INV_X1 U13547 ( .A(n10938), .ZN(n14906) );
  MUX2_X1 U13548 ( .A(n10940), .B(n10939), .S(n12463), .Z(n10942) );
  NAND2_X1 U13549 ( .A1(n10942), .A2(n10941), .ZN(n14924) );
  INV_X1 U13550 ( .A(n10942), .ZN(n10943) );
  NAND2_X1 U13551 ( .A1(n10943), .A2(n14911), .ZN(n10944) );
  AND2_X1 U13552 ( .A1(n14924), .A2(n10944), .ZN(n14905) );
  OAI21_X1 U13553 ( .B1(n14907), .B2(n14906), .A(n14905), .ZN(n14925) );
  MUX2_X1 U13554 ( .A(n10946), .B(n10945), .S(n12463), .Z(n10948) );
  NAND2_X1 U13555 ( .A1(n10948), .A2(n10947), .ZN(n10951) );
  INV_X1 U13556 ( .A(n10948), .ZN(n10949) );
  NAND2_X1 U13557 ( .A1(n10949), .A2(n14928), .ZN(n10950) );
  NAND2_X1 U13558 ( .A1(n10951), .A2(n10950), .ZN(n14923) );
  AOI21_X1 U13559 ( .B1(n14925), .B2(n14924), .A(n14923), .ZN(n14942) );
  INV_X1 U13560 ( .A(n10951), .ZN(n14941) );
  MUX2_X1 U13561 ( .A(n10953), .B(n10952), .S(n12463), .Z(n10955) );
  NAND2_X1 U13562 ( .A1(n10955), .A2(n10954), .ZN(n14959) );
  INV_X1 U13563 ( .A(n10955), .ZN(n10956) );
  NAND2_X1 U13564 ( .A1(n10956), .A2(n14946), .ZN(n10957) );
  AND2_X1 U13565 ( .A1(n14959), .A2(n10957), .ZN(n14940) );
  OAI21_X1 U13566 ( .B1(n14942), .B2(n14941), .A(n14940), .ZN(n14960) );
  MUX2_X1 U13567 ( .A(n10959), .B(n10958), .S(n12463), .Z(n10961) );
  NAND2_X1 U13568 ( .A1(n10961), .A2(n10960), .ZN(n10964) );
  INV_X1 U13569 ( .A(n10961), .ZN(n10962) );
  NAND2_X1 U13570 ( .A1(n10962), .A2(n14965), .ZN(n10963) );
  NAND2_X1 U13571 ( .A1(n10964), .A2(n10963), .ZN(n14958) );
  AOI21_X1 U13572 ( .B1(n14960), .B2(n14959), .A(n14958), .ZN(n14963) );
  INV_X1 U13573 ( .A(n10964), .ZN(n10965) );
  NOR2_X1 U13574 ( .A1(n14963), .A2(n10965), .ZN(n10967) );
  MUX2_X1 U13575 ( .A(P3_REG2_REG_11__SCAN_IN), .B(P3_REG1_REG_11__SCAN_IN), 
        .S(n12463), .Z(n11133) );
  XNOR2_X1 U13576 ( .A(n11133), .B(n11132), .ZN(n10966) );
  NOR2_X1 U13577 ( .A1(n10967), .A2(n10966), .ZN(n12354) );
  AOI21_X1 U13578 ( .B1(n10967), .B2(n10966), .A(n12354), .ZN(n10968) );
  NOR2_X1 U13579 ( .A1(n10968), .A2(n14838), .ZN(n10969) );
  AOI211_X1 U13580 ( .C1(n14973), .C2(n10971), .A(n10970), .B(n10969), .ZN(
        n10972) );
  OAI21_X1 U13581 ( .B1(n10973), .B2(n14977), .A(n10972), .ZN(P3_U3193) );
  NAND2_X1 U13582 ( .A1(n14335), .A2(n13326), .ZN(n11282) );
  XOR2_X1 U13583 ( .A(n11282), .B(n11281), .Z(n11283) );
  XNOR2_X1 U13584 ( .A(n11284), .B(n11283), .ZN(n10982) );
  NOR2_X1 U13585 ( .A1(n14348), .A2(n10992), .ZN(n10980) );
  NAND2_X1 U13586 ( .A1(n13038), .A2(n14336), .ZN(n10978) );
  NAND2_X1 U13587 ( .A1(n13039), .A2(n14334), .ZN(n10977) );
  AND2_X1 U13588 ( .A1(n10978), .A2(n10977), .ZN(n10986) );
  NAND2_X1 U13589 ( .A1(P2_U3088), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n14737)
         );
  OAI21_X1 U13590 ( .B1(n14343), .B2(n10986), .A(n14737), .ZN(n10979) );
  AOI211_X1 U13591 ( .C1(n12032), .C2(n13019), .A(n10980), .B(n10979), .ZN(
        n10981) );
  OAI21_X1 U13592 ( .B1(n10982), .B2(n14342), .A(n10981), .ZN(P2_U3206) );
  NAND2_X1 U13593 ( .A1(n10984), .A2(n10983), .ZN(n12208) );
  XOR2_X1 U13594 ( .A(n10985), .B(n12208), .Z(n10987) );
  OAI21_X1 U13595 ( .B1(n10987), .B2(n14351), .A(n10986), .ZN(n14375) );
  INV_X1 U13596 ( .A(n14375), .ZN(n10998) );
  XNOR2_X1 U13597 ( .A(n10988), .B(n12208), .ZN(n14377) );
  INV_X1 U13598 ( .A(n10989), .ZN(n10991) );
  INV_X1 U13599 ( .A(n10990), .ZN(n14359) );
  OAI211_X1 U13600 ( .C1(n14374), .C2(n10991), .A(n9550), .B(n14359), .ZN(
        n14373) );
  OAI22_X1 U13601 ( .A1(n13281), .A2(n10993), .B1(n10992), .B2(n13323), .ZN(
        n10994) );
  AOI21_X1 U13602 ( .B1(n12032), .B2(n14355), .A(n10994), .ZN(n10995) );
  OAI21_X1 U13603 ( .B1(n14373), .B2(n13330), .A(n10995), .ZN(n10996) );
  AOI21_X1 U13604 ( .B1(n14377), .B2(n14363), .A(n10996), .ZN(n10997) );
  OAI21_X1 U13605 ( .B1(n10998), .B2(n14367), .A(n10997), .ZN(P2_U3252) );
  NAND2_X1 U13606 ( .A1(n14267), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n11113) );
  NAND2_X1 U13607 ( .A1(n13487), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n11001) );
  AND2_X1 U13608 ( .A1(n11113), .A2(n11001), .ZN(n11002) );
  OR2_X1 U13609 ( .A1(n11003), .A2(n11002), .ZN(n11004) );
  OAI222_X1 U13610 ( .A1(n12245), .A2(n11549), .B1(n11338), .B2(n11550), .C1(
        P3_U3151), .C2(n11005), .ZN(P3_U3269) );
  NAND2_X1 U13611 ( .A1(n11010), .A2(n11006), .ZN(n11008) );
  OAI211_X1 U13612 ( .C1(n15293), .C2(n14266), .A(n11008), .B(n11007), .ZN(
        P1_U3332) );
  NAND2_X1 U13613 ( .A1(n11010), .A2(n11009), .ZN(n11012) );
  OR2_X1 U13614 ( .A1(n11011), .A2(P2_U3088), .ZN(n12239) );
  OAI211_X1 U13615 ( .C1(n11013), .C2(n11904), .A(n11012), .B(n12239), .ZN(
        P2_U3304) );
  NAND2_X1 U13616 ( .A1(n11018), .A2(n13640), .ZN(n11015) );
  NAND2_X1 U13617 ( .A1(n13763), .A2(n6536), .ZN(n11014) );
  NAND2_X1 U13618 ( .A1(n11015), .A2(n11014), .ZN(n11016) );
  XNOR2_X1 U13619 ( .A(n11016), .B(n13637), .ZN(n11229) );
  AND2_X1 U13620 ( .A1(n13763), .A2(n13636), .ZN(n11017) );
  AOI21_X1 U13621 ( .B1(n11018), .B2(n6536), .A(n11017), .ZN(n11230) );
  XNOR2_X1 U13622 ( .A(n11229), .B(n11230), .ZN(n11025) );
  INV_X1 U13623 ( .A(n11019), .ZN(n11020) );
  NAND2_X1 U13624 ( .A1(n11024), .A2(n11025), .ZN(n11233) );
  OAI21_X1 U13625 ( .B1(n11025), .B2(n11024), .A(n11233), .ZN(n11026) );
  NAND2_X1 U13626 ( .A1(n11026), .A2(n14395), .ZN(n11034) );
  INV_X1 U13627 ( .A(n11027), .ZN(n11032) );
  INV_X1 U13628 ( .A(n13750), .ZN(n13720) );
  AOI21_X1 U13629 ( .B1(n13718), .B2(n13762), .A(n11028), .ZN(n11029) );
  OAI21_X1 U13630 ( .B1(n13720), .B2(n11030), .A(n11029), .ZN(n11031) );
  AOI21_X1 U13631 ( .B1(n11032), .B2(n13740), .A(n11031), .ZN(n11033) );
  OAI211_X1 U13632 ( .C1(n14411), .C2(n13743), .A(n11034), .B(n11033), .ZN(
        P1_U3236) );
  AOI21_X1 U13633 ( .B1(n13667), .B2(n14607), .A(n11035), .ZN(n11036) );
  OAI211_X1 U13634 ( .C1(n14611), .C2(n11038), .A(n11037), .B(n11036), .ZN(
        n11041) );
  NAND2_X1 U13635 ( .A1(n11041), .A2(n14658), .ZN(n11039) );
  OAI21_X1 U13636 ( .B1(n14658), .B2(n11040), .A(n11039), .ZN(P1_U3540) );
  INV_X1 U13637 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n15327) );
  NAND2_X1 U13638 ( .A1(n11041), .A2(n14645), .ZN(n11042) );
  OAI21_X1 U13639 ( .B1(n14645), .B2(n15327), .A(n11042), .ZN(P1_U3495) );
  XNOR2_X1 U13640 ( .A(n12343), .B(n14996), .ZN(n11834) );
  NAND3_X1 U13641 ( .A1(n11043), .A2(n11047), .A3(n11720), .ZN(n11044) );
  AND2_X1 U13642 ( .A1(n11476), .A2(n11044), .ZN(n14995) );
  NAND2_X1 U13643 ( .A1(n12344), .A2(n15004), .ZN(n11045) );
  OAI21_X1 U13644 ( .B1(n11048), .B2(n11047), .A(n11102), .ZN(n11049) );
  AOI222_X1 U13645 ( .A1(n15046), .A2(n11049), .B1(n14985), .B2(n15038), .C1(
        n12344), .C2(n15041), .ZN(n14994) );
  OAI21_X1 U13646 ( .B1(n12748), .B2(n14995), .A(n14994), .ZN(n11053) );
  INV_X1 U13647 ( .A(n14996), .ZN(n11725) );
  OAI22_X1 U13648 ( .A1(n12780), .A2(n11725), .B1(n15096), .B2(n10945), .ZN(
        n11050) );
  AOI21_X1 U13649 ( .B1(n11053), .B2(n15096), .A(n11050), .ZN(n11051) );
  INV_X1 U13650 ( .A(n11051), .ZN(P3_U3467) );
  OAI22_X1 U13651 ( .A1(n11725), .A2(n12867), .B1(n15085), .B2(n10535), .ZN(
        n11052) );
  AOI21_X1 U13652 ( .B1(n11053), .B2(n15085), .A(n11052), .ZN(n11054) );
  INV_X1 U13653 ( .A(n11054), .ZN(P3_U3414) );
  AND2_X1 U13654 ( .A1(n11055), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n11056) );
  OR2_X1 U13655 ( .A1(n11056), .A2(n11088), .ZN(n14306) );
  INV_X1 U13656 ( .A(n14306), .ZN(n11099) );
  INV_X1 U13657 ( .A(n11057), .ZN(n11058) );
  AND2_X1 U13658 ( .A1(n11058), .A2(n12342), .ZN(n11061) );
  OR2_X1 U13659 ( .A1(n11059), .A2(n11061), .ZN(n11062) );
  OR2_X1 U13660 ( .A1(n11061), .A2(n11060), .ZN(n11063) );
  OR2_X1 U13661 ( .A1(n11062), .A2(n14984), .ZN(n11065) );
  OR2_X1 U13662 ( .A1(n14984), .A2(n11063), .ZN(n11064) );
  OAI21_X1 U13663 ( .B1(n11068), .B2(n11478), .A(n11073), .ZN(n15386) );
  NAND2_X1 U13664 ( .A1(n11069), .A2(n11664), .ZN(n11072) );
  AOI22_X1 U13665 ( .A1(n11493), .A2(n11070), .B1(n11492), .B2(n11132), .ZN(
        n11071) );
  XNOR2_X1 U13666 ( .A(n14321), .B(n11892), .ZN(n15387) );
  INV_X1 U13667 ( .A(n11073), .ZN(n11083) );
  NAND2_X1 U13668 ( .A1(n11074), .A2(n11664), .ZN(n11076) );
  AOI22_X1 U13669 ( .A1(n11493), .A2(SI_12_), .B1(n11492), .B2(n12360), .ZN(
        n11075) );
  XNOR2_X1 U13670 ( .A(n14309), .B(n11892), .ZN(n11166) );
  INV_X1 U13671 ( .A(P3_REG1_REG_12__SCAN_IN), .ZN(n11129) );
  INV_X1 U13672 ( .A(P3_REG2_REG_12__SCAN_IN), .ZN(n11122) );
  OAI21_X1 U13673 ( .B1(n11570), .B2(n11129), .A(n11077), .ZN(n11081) );
  NOR2_X1 U13674 ( .A1(n10012), .A2(n11099), .ZN(n11080) );
  INV_X1 U13675 ( .A(P3_REG0_REG_12__SCAN_IN), .ZN(n11078) );
  NOR2_X1 U13676 ( .A1(n11438), .A2(n11078), .ZN(n11079) );
  XNOR2_X1 U13677 ( .A(n11166), .B(n14320), .ZN(n11082) );
  INV_X1 U13678 ( .A(n11170), .ZN(n11085) );
  NOR3_X1 U13679 ( .A1(n15385), .A2(n11083), .A3(n11082), .ZN(n11084) );
  OAI21_X1 U13680 ( .B1(n11085), .B2(n11084), .A(n12318), .ZN(n11098) );
  INV_X1 U13681 ( .A(P3_REG2_REG_13__SCAN_IN), .ZN(n11086) );
  OR2_X1 U13682 ( .A1(n11088), .A2(n11087), .ZN(n11089) );
  AND2_X1 U13683 ( .A1(n11089), .A2(n11173), .ZN(n12721) );
  OR2_X1 U13684 ( .A1(n10012), .A2(n12721), .ZN(n11091) );
  INV_X1 U13685 ( .A(P3_REG1_REG_13__SCAN_IN), .ZN(n12781) );
  OR2_X1 U13686 ( .A1(n11436), .A2(n12781), .ZN(n11090) );
  INV_X1 U13687 ( .A(P3_REG3_REG_12__SCAN_IN), .ZN(n11094) );
  NOR2_X1 U13688 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11094), .ZN(n12359) );
  AOI21_X1 U13689 ( .B1(n12332), .B2(n14984), .A(n12359), .ZN(n11095) );
  OAI21_X1 U13690 ( .B1(n11589), .B2(n12336), .A(n11095), .ZN(n11096) );
  AOI21_X1 U13691 ( .B1(n12338), .B2(n11592), .A(n11096), .ZN(n11097) );
  OAI211_X1 U13692 ( .C1(n11099), .C2(n15395), .A(n11098), .B(n11097), .ZN(
        P3_U3164) );
  OR2_X1 U13693 ( .A1(n12343), .A2(n11725), .ZN(n11727) );
  NAND2_X1 U13694 ( .A1(n11476), .A2(n11727), .ZN(n11100) );
  XNOR2_X1 U13695 ( .A(n14985), .B(n11730), .ZN(n11835) );
  XNOR2_X1 U13696 ( .A(n11100), .B(n11835), .ZN(n15080) );
  INV_X1 U13697 ( .A(n15080), .ZN(n11112) );
  OR2_X1 U13698 ( .A1(n12343), .A2(n14996), .ZN(n11101) );
  NAND2_X1 U13699 ( .A1(n11104), .A2(n11103), .ZN(n11585) );
  OAI211_X1 U13700 ( .C1(n11104), .C2(n11103), .A(n15046), .B(n11585), .ZN(
        n11106) );
  AOI22_X1 U13701 ( .A1(n12342), .A2(n15038), .B1(n15041), .B2(n12343), .ZN(
        n11105) );
  NAND2_X1 U13702 ( .A1(n11106), .A2(n11105), .ZN(n15078) );
  AND2_X1 U13703 ( .A1(n15052), .A2(P3_REG2_REG_9__SCAN_IN), .ZN(n11110) );
  AND2_X1 U13704 ( .A1(n11730), .A2(n15049), .ZN(n15079) );
  INV_X1 U13705 ( .A(n15079), .ZN(n11108) );
  OAI22_X1 U13706 ( .A1(n12535), .A2(n11108), .B1(n11107), .B2(n15020), .ZN(
        n11109) );
  AOI211_X1 U13707 ( .C1(n15078), .C2(n15057), .A(n11110), .B(n11109), .ZN(
        n11111) );
  OAI21_X1 U13708 ( .B1(n12725), .B2(n11112), .A(n11111), .ZN(P3_U3224) );
  NAND2_X1 U13709 ( .A1(n15217), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n11333) );
  NAND2_X1 U13710 ( .A1(n13485), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n11115) );
  AND2_X1 U13711 ( .A1(n11333), .A2(n11115), .ZN(n11116) );
  OR2_X1 U13712 ( .A1(n11117), .A2(n11116), .ZN(n11118) );
  NAND2_X1 U13713 ( .A1(n11334), .A2(n11118), .ZN(n11559) );
  INV_X1 U13714 ( .A(SI_27_), .ZN(n15188) );
  OAI222_X1 U13715 ( .A1(n12245), .A2(n11559), .B1(n11338), .B2(n15188), .C1(
        P3_U3151), .C2(n12463), .ZN(P3_U3268) );
  INV_X1 U13716 ( .A(n12376), .ZN(n12383) );
  NOR2_X1 U13717 ( .A1(n6890), .A2(n11119), .ZN(n11121) );
  MUX2_X1 U13718 ( .A(P3_REG2_REG_12__SCAN_IN), .B(n11122), .S(n12360), .Z(
        n12361) );
  NAND2_X1 U13719 ( .A1(n11123), .A2(P3_REG2_REG_12__SCAN_IN), .ZN(n11124) );
  AOI21_X1 U13720 ( .B1(n11086), .B2(n11125), .A(n12373), .ZN(n11144) );
  NAND2_X1 U13721 ( .A1(n11132), .A2(n11126), .ZN(n11128) );
  MUX2_X1 U13722 ( .A(n11129), .B(P3_REG1_REG_12__SCAN_IN), .S(n12360), .Z(
        n12365) );
  NAND2_X1 U13723 ( .A1(P3_REG1_REG_13__SCAN_IN), .A2(n11130), .ZN(n12377) );
  OAI21_X1 U13724 ( .B1(P3_REG1_REG_13__SCAN_IN), .B2(n11130), .A(n12377), 
        .ZN(n11142) );
  AND2_X1 U13725 ( .A1(P3_U3151), .A2(P3_REG3_REG_13__SCAN_IN), .ZN(n11179) );
  AOI21_X1 U13726 ( .B1(n14969), .B2(P3_ADDR_REG_13__SCAN_IN), .A(n11179), 
        .ZN(n11131) );
  OAI21_X1 U13727 ( .B1(n14966), .B2(n12376), .A(n11131), .ZN(n11141) );
  NOR2_X1 U13728 ( .A1(n11133), .A2(n11132), .ZN(n12353) );
  MUX2_X1 U13729 ( .A(P3_REG2_REG_12__SCAN_IN), .B(P3_REG1_REG_12__SCAN_IN), 
        .S(n12463), .Z(n11134) );
  XOR2_X1 U13730 ( .A(n12360), .B(n11134), .Z(n12352) );
  NOR3_X1 U13731 ( .A1(n12354), .A2(n12353), .A3(n12352), .ZN(n12351) );
  INV_X1 U13732 ( .A(n11134), .ZN(n11135) );
  NOR2_X1 U13733 ( .A1(n11135), .A2(n12360), .ZN(n11137) );
  MUX2_X1 U13734 ( .A(P3_REG2_REG_13__SCAN_IN), .B(P3_REG1_REG_13__SCAN_IN), 
        .S(n12463), .Z(n12380) );
  XNOR2_X1 U13735 ( .A(n12380), .B(n12376), .ZN(n11136) );
  NOR3_X1 U13736 ( .A1(n12351), .A2(n11137), .A3(n11136), .ZN(n12381) );
  INV_X1 U13737 ( .A(n12381), .ZN(n11139) );
  OAI21_X1 U13738 ( .B1(n12351), .B2(n11137), .A(n11136), .ZN(n11138) );
  AOI21_X1 U13739 ( .B1(n11139), .B2(n11138), .A(n14838), .ZN(n11140) );
  AOI211_X1 U13740 ( .C1(n11142), .C2(n14973), .A(n11141), .B(n11140), .ZN(
        n11143) );
  OAI21_X1 U13741 ( .B1(n11144), .B2(n14977), .A(n11143), .ZN(P3_U3195) );
  OR2_X1 U13742 ( .A1(n13667), .A2(n13762), .ZN(n11145) );
  NAND2_X1 U13743 ( .A1(n11146), .A2(n11145), .ZN(n11147) );
  OAI21_X1 U13744 ( .B1(n11147), .B2(n11151), .A(n11211), .ZN(n11148) );
  INV_X1 U13745 ( .A(n11148), .ZN(n11204) );
  NAND2_X1 U13746 ( .A1(n11150), .A2(n11149), .ZN(n11153) );
  INV_X1 U13747 ( .A(n11151), .ZN(n11152) );
  NAND2_X1 U13748 ( .A1(n11153), .A2(n11152), .ZN(n11220) );
  OAI211_X1 U13749 ( .C1(n11153), .C2(n11152), .A(n11220), .B(n14497), .ZN(
        n11202) );
  INV_X1 U13750 ( .A(n11202), .ZN(n11155) );
  NAND2_X1 U13751 ( .A1(n13762), .A2(n14107), .ZN(n11154) );
  OAI21_X1 U13752 ( .B1(n13506), .B2(n14581), .A(n11154), .ZN(n11249) );
  OAI21_X1 U13753 ( .B1(n11155), .B2(n11249), .A(n14543), .ZN(n11161) );
  AOI211_X1 U13754 ( .C1(n11253), .C2(n11156), .A(n14572), .B(n6970), .ZN(
        n11201) );
  NOR2_X1 U13755 ( .A1(n6971), .A2(n14119), .ZN(n11159) );
  OAI22_X1 U13756 ( .A1(n14543), .A2(n11157), .B1(n11251), .B2(n14542), .ZN(
        n11158) );
  AOI211_X1 U13757 ( .C1(n11201), .C2(n14574), .A(n11159), .B(n11158), .ZN(
        n11160) );
  OAI211_X1 U13758 ( .C1(n11204), .C2(n14123), .A(n11161), .B(n11160), .ZN(
        P1_U3280) );
  NAND2_X1 U13759 ( .A1(n11162), .A2(n11664), .ZN(n11165) );
  AOI22_X1 U13760 ( .A1(n11493), .A2(n11163), .B1(n11492), .B2(n12376), .ZN(
        n11164) );
  NAND2_X1 U13761 ( .A1(n11165), .A2(n11164), .ZN(n11593) );
  INV_X1 U13762 ( .A(n11166), .ZN(n11167) );
  NAND2_X1 U13763 ( .A1(n11167), .A2(n14320), .ZN(n11168) );
  AND2_X1 U13764 ( .A1(n11170), .A2(n11168), .ZN(n11172) );
  XNOR2_X1 U13765 ( .A(n11593), .B(n11892), .ZN(n11264) );
  XNOR2_X1 U13766 ( .A(n11264), .B(n11589), .ZN(n11171) );
  OAI211_X1 U13767 ( .C1(n11172), .C2(n11171), .A(n12318), .B(n11268), .ZN(
        n11184) );
  INV_X1 U13768 ( .A(n12721), .ZN(n11182) );
  NAND2_X1 U13769 ( .A1(n11173), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n11174) );
  AND2_X1 U13770 ( .A1(n11270), .A2(n11174), .ZN(n12708) );
  INV_X1 U13771 ( .A(P3_REG1_REG_14__SCAN_IN), .ZN(n12777) );
  OR2_X1 U13772 ( .A1(n11436), .A2(n12777), .ZN(n11175) );
  OAI21_X1 U13773 ( .B1(n10012), .B2(n12708), .A(n11175), .ZN(n11178) );
  INV_X1 U13774 ( .A(P3_REG0_REG_14__SCAN_IN), .ZN(n12862) );
  NOR2_X1 U13775 ( .A1(n11438), .A2(n12862), .ZN(n11177) );
  INV_X1 U13776 ( .A(P3_REG2_REG_14__SCAN_IN), .ZN(n12705) );
  AOI21_X1 U13777 ( .B1(n15389), .B2(n12719), .A(n11179), .ZN(n11180) );
  OAI21_X1 U13778 ( .B1(n14320), .B2(n15392), .A(n11180), .ZN(n11181) );
  AOI21_X1 U13779 ( .B1(n12333), .B2(n11182), .A(n11181), .ZN(n11183) );
  OAI211_X1 U13780 ( .C1(n12327), .C2(n11593), .A(n11184), .B(n11183), .ZN(
        P3_U3174) );
  OAI21_X1 U13781 ( .B1(n11187), .B2(n11186), .A(n11185), .ZN(n11191) );
  NAND2_X1 U13782 ( .A1(n13821), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n11188) );
  OAI21_X1 U13783 ( .B1(n13821), .B2(P1_REG2_REG_17__SCAN_IN), .A(n11188), 
        .ZN(n11190) );
  NAND2_X1 U13784 ( .A1(n11195), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n11189) );
  OAI211_X1 U13785 ( .C1(n11195), .C2(P1_REG2_REG_17__SCAN_IN), .A(n11191), 
        .B(n11189), .ZN(n13818) );
  OAI211_X1 U13786 ( .C1(n11191), .C2(n11190), .A(n14478), .B(n13818), .ZN(
        n11200) );
  NAND2_X1 U13787 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n13695)
         );
  INV_X1 U13788 ( .A(n11192), .ZN(n11193) );
  XNOR2_X1 U13789 ( .A(n11195), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n13823) );
  XOR2_X1 U13790 ( .A(n13824), .B(n13823), .Z(n11196) );
  NAND2_X1 U13791 ( .A1(n14483), .A2(n11196), .ZN(n11197) );
  NAND2_X1 U13792 ( .A1(n13695), .A2(n11197), .ZN(n11198) );
  AOI21_X1 U13793 ( .B1(n14472), .B2(P1_ADDR_REG_17__SCAN_IN), .A(n11198), 
        .ZN(n11199) );
  OAI211_X1 U13794 ( .C1(n13832), .C2(n13821), .A(n11200), .B(n11199), .ZN(
        P1_U3260) );
  AOI211_X1 U13795 ( .C1(n11253), .C2(n14607), .A(n11249), .B(n11201), .ZN(
        n11203) );
  OAI211_X1 U13796 ( .C1(n14611), .C2(n11204), .A(n11203), .B(n11202), .ZN(
        n11207) );
  NAND2_X1 U13797 ( .A1(n11207), .A2(n14658), .ZN(n11205) );
  OAI21_X1 U13798 ( .B1(n14658), .B2(n11206), .A(n11205), .ZN(P1_U3541) );
  INV_X1 U13799 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n11209) );
  NAND2_X1 U13800 ( .A1(n11207), .A2(n14645), .ZN(n11208) );
  OAI21_X1 U13801 ( .B1(n14645), .B2(n11209), .A(n11208), .ZN(P1_U3498) );
  OR2_X1 U13802 ( .A1(n11253), .A2(n13761), .ZN(n11210) );
  OAI21_X1 U13803 ( .B1(n11221), .B2(n7429), .A(n11302), .ZN(n14407) );
  AOI211_X1 U13804 ( .C1(n14405), .C2(n11213), .A(n14572), .B(n6968), .ZN(
        n14403) );
  OAI22_X1 U13805 ( .A1(n11218), .A2(n14561), .B1(n13517), .B2(n14581), .ZN(
        n14404) );
  OAI22_X1 U13806 ( .A1(n14543), .A2(n11214), .B1(n14402), .B2(n14542), .ZN(
        n11215) );
  AOI21_X1 U13807 ( .B1(n14543), .B2(n14404), .A(n11215), .ZN(n11216) );
  OAI21_X1 U13808 ( .B1(n6969), .B2(n14119), .A(n11216), .ZN(n11217) );
  AOI21_X1 U13809 ( .B1(n14403), .B2(n14574), .A(n11217), .ZN(n11223) );
  OR2_X1 U13810 ( .A1(n11253), .A2(n11218), .ZN(n11219) );
  NAND2_X1 U13811 ( .A1(n11220), .A2(n11219), .ZN(n11297) );
  XNOR2_X1 U13812 ( .A(n11297), .B(n11221), .ZN(n14409) );
  INV_X1 U13813 ( .A(n14085), .ZN(n13967) );
  NAND2_X1 U13814 ( .A1(n14409), .A2(n13967), .ZN(n11222) );
  OAI211_X1 U13815 ( .C1(n14407), .C2(n14123), .A(n11223), .B(n11222), .ZN(
        P1_U3279) );
  INV_X1 U13816 ( .A(n11224), .ZN(n11227) );
  OAI222_X1 U13817 ( .A1(P1_U3086), .A2(n11225), .B1(n6535), .B2(n11227), .C1(
        n7368), .C2(n14266), .ZN(P1_U3331) );
  OAI222_X1 U13818 ( .A1(n11904), .A2(n11228), .B1(n6534), .B2(n11227), .C1(
        n11226), .C2(P2_U3088), .ZN(P2_U3303) );
  INV_X1 U13819 ( .A(n11229), .ZN(n11231) );
  NAND2_X1 U13820 ( .A1(n11231), .A2(n11230), .ZN(n11232) );
  NAND2_X1 U13821 ( .A1(n11233), .A2(n11232), .ZN(n13663) );
  INV_X1 U13822 ( .A(n13663), .ZN(n11239) );
  NAND2_X1 U13823 ( .A1(n13667), .A2(n13640), .ZN(n11235) );
  NAND2_X1 U13824 ( .A1(n13762), .A2(n6536), .ZN(n11234) );
  NAND2_X1 U13825 ( .A1(n11235), .A2(n11234), .ZN(n11236) );
  XNOR2_X1 U13826 ( .A(n11236), .B(n13591), .ZN(n11240) );
  AND2_X1 U13827 ( .A1(n13762), .A2(n13636), .ZN(n11237) );
  AOI21_X1 U13828 ( .B1(n13667), .B2(n6536), .A(n11237), .ZN(n11241) );
  XNOR2_X1 U13829 ( .A(n11240), .B(n11241), .ZN(n13664) );
  INV_X1 U13830 ( .A(n11240), .ZN(n11243) );
  INV_X1 U13831 ( .A(n11241), .ZN(n11242) );
  NAND2_X1 U13832 ( .A1(n11243), .A2(n11242), .ZN(n11244) );
  NAND2_X1 U13833 ( .A1(n11253), .A2(n13640), .ZN(n11246) );
  NAND2_X1 U13834 ( .A1(n13761), .A2(n6536), .ZN(n11245) );
  NAND2_X1 U13835 ( .A1(n11246), .A2(n11245), .ZN(n11247) );
  XNOR2_X1 U13836 ( .A(n11247), .B(n13637), .ZN(n13502) );
  AND2_X1 U13837 ( .A1(n13761), .A2(n13636), .ZN(n11248) );
  AOI21_X1 U13838 ( .B1(n11253), .B2(n6536), .A(n11248), .ZN(n13500) );
  XNOR2_X1 U13839 ( .A(n13502), .B(n13500), .ZN(n13498) );
  XNOR2_X1 U13840 ( .A(n13499), .B(n13498), .ZN(n11255) );
  NAND2_X1 U13841 ( .A1(P1_U3086), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n14473)
         );
  NAND2_X1 U13842 ( .A1(n11249), .A2(n14397), .ZN(n11250) );
  OAI211_X1 U13843 ( .C1(n14401), .C2(n11251), .A(n14473), .B(n11250), .ZN(
        n11252) );
  AOI21_X1 U13844 ( .B1(n11253), .B2(n14398), .A(n11252), .ZN(n11254) );
  OAI21_X1 U13845 ( .B1(n11255), .B2(n13756), .A(n11254), .ZN(P1_U3234) );
  INV_X1 U13846 ( .A(n11256), .ZN(n11258) );
  OAI222_X1 U13847 ( .A1(n11904), .A2(n15170), .B1(n6534), .B2(n11258), .C1(
        n11257), .C2(P2_U3088), .ZN(P2_U3302) );
  OAI222_X1 U13848 ( .A1(P1_U3086), .A2(n11259), .B1(n6535), .B2(n11258), .C1(
        n15297), .C2(n14266), .ZN(P1_U3330) );
  NAND2_X1 U13849 ( .A1(n11260), .A2(n11664), .ZN(n11263) );
  AOI22_X1 U13850 ( .A1(n11493), .A2(n11261), .B1(n11492), .B2(n12400), .ZN(
        n11262) );
  XNOR2_X1 U13851 ( .A(n12866), .B(n11892), .ZN(n11313) );
  INV_X1 U13852 ( .A(n12719), .ZN(n11597) );
  XNOR2_X1 U13853 ( .A(n11313), .B(n11597), .ZN(n11266) );
  NAND2_X1 U13854 ( .A1(n11264), .A2(n14304), .ZN(n11267) );
  AOI21_X1 U13855 ( .B1(n11268), .B2(n11267), .A(n11266), .ZN(n11269) );
  OAI21_X1 U13856 ( .B1(n6685), .B2(n11269), .A(n12318), .ZN(n11280) );
  INV_X1 U13857 ( .A(n12708), .ZN(n11278) );
  INV_X1 U13858 ( .A(P3_REG2_REG_15__SCAN_IN), .ZN(n12693) );
  AND2_X1 U13859 ( .A1(n11270), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n11271) );
  NOR2_X1 U13860 ( .A1(n11321), .A2(n11271), .ZN(n12694) );
  OR2_X1 U13861 ( .A1(n10012), .A2(n12694), .ZN(n11273) );
  INV_X1 U13862 ( .A(P3_REG1_REG_15__SCAN_IN), .ZN(n12773) );
  OR2_X1 U13863 ( .A1(n11570), .A2(n12773), .ZN(n11272) );
  AND2_X1 U13864 ( .A1(P3_U3151), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n12389) );
  AOI21_X1 U13865 ( .B1(n12332), .B2(n14304), .A(n12389), .ZN(n11276) );
  OAI21_X1 U13866 ( .B1(n12678), .B2(n12336), .A(n11276), .ZN(n11277) );
  AOI21_X1 U13867 ( .B1(n12333), .B2(n11278), .A(n11277), .ZN(n11279) );
  OAI211_X1 U13868 ( .C1(n12327), .C2(n12866), .A(n11280), .B(n11279), .ZN(
        P3_U3155) );
  XNOR2_X1 U13869 ( .A(n14356), .B(n6541), .ZN(n11286) );
  NAND2_X1 U13870 ( .A1(n13038), .A2(n13326), .ZN(n11285) );
  OAI21_X1 U13871 ( .B1(n11286), .B2(n11285), .A(n11373), .ZN(n14339) );
  INV_X1 U13872 ( .A(n11373), .ZN(n11287) );
  NOR2_X1 U13873 ( .A1(n6683), .A2(n11287), .ZN(n11289) );
  XNOR2_X1 U13874 ( .A(n12050), .B(n6528), .ZN(n11375) );
  AND2_X1 U13875 ( .A1(n14337), .A2(n13326), .ZN(n11374) );
  INV_X1 U13876 ( .A(n11374), .ZN(n11376) );
  XNOR2_X1 U13877 ( .A(n11375), .B(n11376), .ZN(n11288) );
  XNOR2_X1 U13878 ( .A(n11289), .B(n11288), .ZN(n11294) );
  AOI22_X1 U13879 ( .A1(n13037), .A2(n14336), .B1(n14334), .B2(n13038), .ZN(
        n11350) );
  INV_X1 U13880 ( .A(n11350), .ZN(n11290) );
  AOI22_X1 U13881 ( .A1(n13016), .A2(n11290), .B1(P2_REG3_REG_15__SCAN_IN), 
        .B2(P2_U3088), .ZN(n11291) );
  OAI21_X1 U13882 ( .B1(n11345), .B2(n14348), .A(n11291), .ZN(n11292) );
  AOI21_X1 U13883 ( .B1(n12050), .B2(n13019), .A(n11292), .ZN(n11293) );
  OAI21_X1 U13884 ( .B1(n11294), .B2(n14342), .A(n11293), .ZN(P2_U3213) );
  INV_X1 U13885 ( .A(n11387), .ZN(n11303) );
  XNOR2_X1 U13886 ( .A(n11388), .B(n11303), .ZN(n11300) );
  NAND2_X1 U13887 ( .A1(n14106), .A2(n14108), .ZN(n11298) );
  OAI21_X1 U13888 ( .B1(n13506), .B2(n14561), .A(n11298), .ZN(n11299) );
  AOI21_X1 U13889 ( .B1(n11300), .B2(n14497), .A(n11299), .ZN(n14233) );
  INV_X1 U13890 ( .A(n13506), .ZN(n13760) );
  NAND2_X1 U13891 ( .A1(n14405), .A2(n13760), .ZN(n11301) );
  NAND2_X1 U13892 ( .A1(n11304), .A2(n11303), .ZN(n11305) );
  NAND2_X1 U13893 ( .A1(n11397), .A2(n11305), .ZN(n14231) );
  AOI21_X1 U13894 ( .B1(n13754), .B2(n11306), .A(n14572), .ZN(n11307) );
  NAND2_X1 U13895 ( .A1(n11307), .A2(n11391), .ZN(n14229) );
  INV_X1 U13896 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n11308) );
  OAI22_X1 U13897 ( .A1(n14543), .A2(n11308), .B1(n13752), .B2(n14542), .ZN(
        n11309) );
  AOI21_X1 U13898 ( .B1(n13754), .B2(n14566), .A(n11309), .ZN(n11310) );
  OAI21_X1 U13899 ( .B1(n14229), .B2(n13959), .A(n11310), .ZN(n11311) );
  AOI21_X1 U13900 ( .B1(n14231), .B2(n14083), .A(n11311), .ZN(n11312) );
  OAI21_X1 U13901 ( .B1(n14233), .B2(n6531), .A(n11312), .ZN(P1_U3278) );
  NAND2_X1 U13902 ( .A1(n11314), .A2(n11664), .ZN(n11317) );
  AOI22_X1 U13903 ( .A1(n11493), .A2(n11315), .B1(n11492), .B2(n12422), .ZN(
        n11316) );
  XNOR2_X1 U13904 ( .A(n11601), .B(n11892), .ZN(n11318) );
  NAND2_X1 U13905 ( .A1(n11318), .A2(n12703), .ZN(n11429) );
  NAND2_X1 U13906 ( .A1(n6695), .A2(n11429), .ZN(n11319) );
  XNOR2_X1 U13907 ( .A(n11430), .B(n11319), .ZN(n11332) );
  INV_X1 U13908 ( .A(n11601), .ZN(n12856) );
  NOR2_X1 U13909 ( .A1(n11321), .A2(n11320), .ZN(n11322) );
  OR2_X1 U13910 ( .A1(n11433), .A2(n11322), .ZN(n12684) );
  INV_X1 U13911 ( .A(n12684), .ZN(n11324) );
  INV_X1 U13912 ( .A(P3_REG1_REG_16__SCAN_IN), .ZN(n12770) );
  OR2_X1 U13913 ( .A1(n11570), .A2(n12770), .ZN(n11323) );
  OAI21_X1 U13914 ( .B1(n10012), .B2(n11324), .A(n11323), .ZN(n11327) );
  INV_X1 U13915 ( .A(P3_REG2_REG_16__SCAN_IN), .ZN(n12683) );
  INV_X1 U13916 ( .A(P3_REG0_REG_16__SCAN_IN), .ZN(n12849) );
  NOR2_X1 U13917 ( .A1(n11438), .A2(n12849), .ZN(n11325) );
  NAND2_X1 U13918 ( .A1(P3_U3151), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n12407)
         );
  OAI21_X1 U13919 ( .B1(n15392), .B2(n11597), .A(n12407), .ZN(n11328) );
  AOI21_X1 U13920 ( .B1(n15389), .B2(n12691), .A(n11328), .ZN(n11329) );
  OAI21_X1 U13921 ( .B1(n15395), .B2(n12694), .A(n11329), .ZN(n11330) );
  AOI21_X1 U13922 ( .B1(n12856), .B2(n12338), .A(n11330), .ZN(n11331) );
  OAI21_X1 U13923 ( .B1(n11332), .B2(n15401), .A(n11331), .ZN(P3_U3181) );
  NAND2_X1 U13924 ( .A1(n11576), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n11335) );
  NAND2_X1 U13925 ( .A1(n11639), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n11336) );
  XNOR2_X1 U13926 ( .A(n13477), .B(P2_DATAO_REG_29__SCAN_IN), .ZN(n11641) );
  XNOR2_X1 U13927 ( .A(n11643), .B(n11641), .ZN(n11581) );
  INV_X1 U13928 ( .A(n11581), .ZN(n11340) );
  OAI222_X1 U13929 ( .A1(n12245), .A2(n11340), .B1(P3_U3151), .B2(n11339), 
        .C1(n11582), .C2(n11338), .ZN(P3_U3266) );
  XNOR2_X1 U13930 ( .A(n11342), .B(n11341), .ZN(n11417) );
  AOI21_X1 U13931 ( .B1(n12050), .B2(n14360), .A(n9445), .ZN(n11343) );
  NAND2_X1 U13932 ( .A1(n11343), .A2(n11406), .ZN(n11418) );
  NAND2_X1 U13933 ( .A1(n14367), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n11344) );
  OAI21_X1 U13934 ( .B1(n13323), .B2(n11345), .A(n11344), .ZN(n11346) );
  AOI21_X1 U13935 ( .B1(n12050), .B2(n14355), .A(n11346), .ZN(n11347) );
  OAI21_X1 U13936 ( .B1(n11418), .B2(n13330), .A(n11347), .ZN(n11353) );
  OAI211_X1 U13937 ( .C1(n11349), .C2(n12210), .A(n11348), .B(n13335), .ZN(
        n11351) );
  AND2_X1 U13938 ( .A1(n11351), .A2(n11350), .ZN(n11420) );
  NOR2_X1 U13939 ( .A1(n11420), .A2(n14367), .ZN(n11352) );
  AOI211_X1 U13940 ( .C1(n11417), .C2(n14363), .A(n11353), .B(n11352), .ZN(
        n11354) );
  INV_X1 U13941 ( .A(n11354), .ZN(P2_U3250) );
  INV_X1 U13942 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n11356) );
  AOI22_X1 U13943 ( .A1(P2_REG2_REG_17__SCAN_IN), .A2(n11361), .B1(n13124), 
        .B2(n11356), .ZN(n13121) );
  OAI21_X1 U13944 ( .B1(n11409), .B2(n11363), .A(n11355), .ZN(n13122) );
  NAND2_X1 U13945 ( .A1(n13121), .A2(n13122), .ZN(n13120) );
  OAI21_X1 U13946 ( .B1(n13124), .B2(n11356), .A(n13120), .ZN(n11357) );
  NOR2_X1 U13947 ( .A1(n11357), .A2(n13135), .ZN(n13132) );
  AOI21_X1 U13948 ( .B1(n13135), .B2(n11357), .A(n13132), .ZN(n11358) );
  INV_X1 U13949 ( .A(n11358), .ZN(n11359) );
  NOR2_X1 U13950 ( .A1(P2_REG2_REG_18__SCAN_IN), .A2(n11359), .ZN(n13133) );
  AOI21_X1 U13951 ( .B1(n11359), .B2(P2_REG2_REG_18__SCAN_IN), .A(n13133), 
        .ZN(n11370) );
  NAND2_X1 U13952 ( .A1(P2_U3088), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n13007)
         );
  OAI21_X1 U13953 ( .B1(n14739), .B2(n11366), .A(n13007), .ZN(n11360) );
  AOI21_X1 U13954 ( .B1(n14752), .B2(P2_ADDR_REG_18__SCAN_IN), .A(n11360), 
        .ZN(n11369) );
  INV_X1 U13955 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n13421) );
  AOI22_X1 U13956 ( .A1(P2_REG1_REG_17__SCAN_IN), .A2(n11361), .B1(n13124), 
        .B2(n13421), .ZN(n13127) );
  INV_X1 U13957 ( .A(n11362), .ZN(n11365) );
  OAI22_X1 U13958 ( .A1(n11365), .A2(n11364), .B1(n11363), .B2(n15259), .ZN(
        n13128) );
  NAND2_X1 U13959 ( .A1(n13127), .A2(n13128), .ZN(n13126) );
  OAI21_X1 U13960 ( .B1(n13124), .B2(n13421), .A(n13126), .ZN(n13136) );
  XNOR2_X1 U13961 ( .A(n13136), .B(n11366), .ZN(n11367) );
  NAND2_X1 U13962 ( .A1(P2_REG1_REG_18__SCAN_IN), .A2(n11367), .ZN(n13138) );
  OAI211_X1 U13963 ( .C1(P2_REG1_REG_18__SCAN_IN), .C2(n11367), .A(n14759), 
        .B(n13138), .ZN(n11368) );
  OAI211_X1 U13964 ( .C1(n11370), .C2(n14745), .A(n11369), .B(n11368), .ZN(
        P2_U3232) );
  XNOR2_X1 U13965 ( .A(n13426), .B(n6540), .ZN(n11372) );
  NAND2_X1 U13966 ( .A1(n13037), .A2(n13326), .ZN(n11371) );
  NAND2_X1 U13967 ( .A1(n11372), .A2(n11371), .ZN(n11459) );
  OAI21_X1 U13968 ( .B1(n11372), .B2(n11371), .A(n11459), .ZN(n11379) );
  OAI21_X1 U13969 ( .B1(n11375), .B2(n11374), .A(n11373), .ZN(n11377) );
  AOI21_X1 U13970 ( .B1(n11379), .B2(n11378), .A(n11461), .ZN(n11386) );
  AND2_X1 U13971 ( .A1(n14337), .A2(n14334), .ZN(n11380) );
  AOI21_X1 U13972 ( .B1(n13036), .B2(n14336), .A(n11380), .ZN(n11403) );
  INV_X1 U13973 ( .A(n11381), .ZN(n11405) );
  NAND2_X1 U13974 ( .A1(n13000), .A2(n11405), .ZN(n11383) );
  OAI211_X1 U13975 ( .C1(n14343), .C2(n11403), .A(n11383), .B(n11382), .ZN(
        n11384) );
  AOI21_X1 U13976 ( .B1(n13426), .B2(n13019), .A(n11384), .ZN(n11385) );
  OAI21_X1 U13977 ( .B1(n11386), .B2(n14342), .A(n11385), .ZN(P2_U3198) );
  OR2_X1 U13978 ( .A1(n11388), .A2(n11387), .ZN(n11390) );
  XNOR2_X1 U13979 ( .A(n13866), .B(n11398), .ZN(n14228) );
  AOI211_X1 U13980 ( .C1(n13890), .C2(n11391), .A(n14572), .B(n14112), .ZN(
        n14224) );
  AOI22_X1 U13981 ( .A1(n13759), .A2(n14107), .B1(n14088), .B2(n14108), .ZN(
        n14222) );
  NAND2_X1 U13982 ( .A1(n13890), .A2(n14566), .ZN(n11394) );
  INV_X1 U13983 ( .A(n13685), .ZN(n11392) );
  AOI22_X1 U13984 ( .A1(n6531), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n11392), 
        .B2(n14567), .ZN(n11393) );
  OAI211_X1 U13985 ( .C1(n6531), .C2(n14222), .A(n11394), .B(n11393), .ZN(
        n11395) );
  AOI21_X1 U13986 ( .B1(n14224), .B2(n14574), .A(n11395), .ZN(n11400) );
  OR2_X1 U13987 ( .A1(n13754), .A2(n13759), .ZN(n11396) );
  NAND2_X1 U13988 ( .A1(n11397), .A2(n11396), .ZN(n13889) );
  INV_X1 U13989 ( .A(n11398), .ZN(n13865) );
  XNOR2_X1 U13990 ( .A(n13889), .B(n13865), .ZN(n14226) );
  NAND2_X1 U13991 ( .A1(n14226), .A2(n14083), .ZN(n11399) );
  OAI211_X1 U13992 ( .C1(n14228), .C2(n14085), .A(n11400), .B(n11399), .ZN(
        P1_U3277) );
  XNOR2_X1 U13993 ( .A(n11401), .B(n7870), .ZN(n11402) );
  NAND2_X1 U13994 ( .A1(n11402), .A2(n13335), .ZN(n11404) );
  NAND2_X1 U13995 ( .A1(n11404), .A2(n11403), .ZN(n13431) );
  AOI21_X1 U13996 ( .B1(n11405), .B2(n14354), .A(n13431), .ZN(n11416) );
  NAND2_X1 U13997 ( .A1(n13426), .A2(n11406), .ZN(n11407) );
  NAND2_X1 U13998 ( .A1(n11407), .A2(n9550), .ZN(n11408) );
  OR2_X1 U13999 ( .A1(n11450), .A2(n11408), .ZN(n13428) );
  INV_X1 U14000 ( .A(n13428), .ZN(n11411) );
  OAI22_X1 U14001 ( .A1(n6810), .A2(n13311), .B1(n13281), .B2(n11409), .ZN(
        n11410) );
  AOI21_X1 U14002 ( .B1(n11411), .B2(n14362), .A(n11410), .ZN(n11415) );
  NAND2_X1 U14003 ( .A1(n11413), .A2(n12211), .ZN(n13424) );
  NAND3_X1 U14004 ( .A1(n13425), .A2(n13424), .A3(n14363), .ZN(n11414) );
  OAI211_X1 U14005 ( .C1(n11416), .C2(n14367), .A(n11415), .B(n11414), .ZN(
        P2_U3249) );
  INV_X1 U14006 ( .A(n13468), .ZN(n13460) );
  NAND2_X1 U14007 ( .A1(n11417), .A2(n14378), .ZN(n11419) );
  NAND3_X1 U14008 ( .A1(n11420), .A2(n11419), .A3(n11418), .ZN(n11423) );
  MUX2_X1 U14009 ( .A(P2_REG0_REG_15__SCAN_IN), .B(n11423), .S(n14821), .Z(
        n11421) );
  AOI21_X1 U14010 ( .B1(n13460), .B2(n12050), .A(n11421), .ZN(n11422) );
  INV_X1 U14011 ( .A(n11422), .ZN(P2_U3475) );
  MUX2_X1 U14012 ( .A(P2_REG1_REG_15__SCAN_IN), .B(n11423), .S(n14829), .Z(
        n11424) );
  AOI21_X1 U14013 ( .B1(n13398), .B2(n12050), .A(n11424), .ZN(n11425) );
  INV_X1 U14014 ( .A(n11425), .ZN(P2_U3514) );
  NAND2_X1 U14015 ( .A1(n11426), .A2(n11664), .ZN(n11428) );
  AOI22_X1 U14016 ( .A1(n11493), .A2(SI_16_), .B1(n11492), .B2(n12453), .ZN(
        n11427) );
  XNOR2_X1 U14017 ( .A(n11483), .B(n11892), .ZN(n11866) );
  XNOR2_X1 U14018 ( .A(n11866), .B(n11868), .ZN(n11431) );
  OAI211_X1 U14019 ( .C1(n11432), .C2(n11431), .A(n11867), .B(n12318), .ZN(
        n11445) );
  OR2_X1 U14020 ( .A1(n11433), .A2(n15204), .ZN(n11434) );
  AND2_X1 U14021 ( .A1(n11435), .A2(n11434), .ZN(n12290) );
  INV_X1 U14022 ( .A(P3_REG1_REG_17__SCAN_IN), .ZN(n12767) );
  OR2_X1 U14023 ( .A1(n11436), .A2(n12767), .ZN(n11437) );
  OAI21_X1 U14024 ( .B1(n10012), .B2(n12290), .A(n11437), .ZN(n11441) );
  INV_X1 U14025 ( .A(P3_REG2_REG_17__SCAN_IN), .ZN(n12668) );
  INV_X1 U14026 ( .A(P3_REG0_REG_17__SCAN_IN), .ZN(n12842) );
  NOR2_X1 U14027 ( .A1(n11438), .A2(n12842), .ZN(n11439) );
  NAND2_X1 U14028 ( .A1(n12332), .A2(n12703), .ZN(n11442) );
  NAND2_X1 U14029 ( .A1(P3_U3151), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n12427)
         );
  OAI211_X1 U14030 ( .C1(n12679), .C2(n12336), .A(n11442), .B(n12427), .ZN(
        n11443) );
  AOI21_X1 U14031 ( .B1(n12333), .B2(n12684), .A(n11443), .ZN(n11444) );
  OAI211_X1 U14032 ( .C1(n11483), .C2(n12327), .A(n11445), .B(n11444), .ZN(
        P3_U3166) );
  OR2_X1 U14033 ( .A1(n11447), .A2(n11446), .ZN(n11448) );
  AND2_X1 U14034 ( .A1(n11449), .A2(n11448), .ZN(n13420) );
  INV_X1 U14035 ( .A(n13420), .ZN(n11458) );
  INV_X1 U14036 ( .A(n13327), .ZN(n11451) );
  AOI211_X1 U14037 ( .C1(n12065), .C2(n6812), .A(n12940), .B(n11451), .ZN(
        n13418) );
  NOR2_X1 U14038 ( .A1(n13469), .A2(n13311), .ZN(n11453) );
  OAI22_X1 U14039 ( .A1(n13281), .A2(n11356), .B1(n11466), .B2(n13323), .ZN(
        n11452) );
  AOI211_X1 U14040 ( .C1(n13418), .C2(n14362), .A(n11453), .B(n11452), .ZN(
        n11457) );
  XNOR2_X1 U14041 ( .A(n11454), .B(n12213), .ZN(n11455) );
  AOI22_X1 U14042 ( .A1(n13035), .A2(n14336), .B1(n14334), .B2(n13037), .ZN(
        n11467) );
  OAI21_X1 U14043 ( .B1(n11455), .B2(n14351), .A(n11467), .ZN(n13419) );
  NAND2_X1 U14044 ( .A1(n13419), .A2(n13281), .ZN(n11456) );
  OAI211_X1 U14045 ( .C1(n11458), .C2(n13342), .A(n11457), .B(n11456), .ZN(
        P2_U3248) );
  INV_X1 U14046 ( .A(n11459), .ZN(n11460) );
  XNOR2_X1 U14047 ( .A(n12065), .B(n6541), .ZN(n11463) );
  NAND2_X1 U14048 ( .A1(n13036), .A2(n13326), .ZN(n11462) );
  NAND2_X1 U14049 ( .A1(n11463), .A2(n11462), .ZN(n12884) );
  OAI21_X1 U14050 ( .B1(n11463), .B2(n11462), .A(n12884), .ZN(n11464) );
  AOI21_X1 U14051 ( .B1(n11465), .B2(n11464), .A(n12886), .ZN(n11471) );
  NOR2_X1 U14052 ( .A1(n14348), .A2(n11466), .ZN(n11469) );
  NAND2_X1 U14053 ( .A1(P2_U3088), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n13123)
         );
  OAI21_X1 U14054 ( .B1(n11467), .B2(n14343), .A(n13123), .ZN(n11468) );
  AOI211_X1 U14055 ( .C1(n12065), .C2(n13019), .A(n11469), .B(n11468), .ZN(
        n11470) );
  OAI21_X1 U14056 ( .B1(n11471), .B2(n14342), .A(n11470), .ZN(P2_U3200) );
  NAND2_X1 U14057 ( .A1(n11472), .A2(n11730), .ZN(n11473) );
  AND2_X1 U14058 ( .A1(n11727), .A2(n11473), .ZN(n11475) );
  INV_X1 U14059 ( .A(n11730), .ZN(n11474) );
  NAND2_X1 U14060 ( .A1(n15393), .A2(n14988), .ZN(n11738) );
  INV_X1 U14061 ( .A(n14988), .ZN(n11477) );
  NAND2_X1 U14062 ( .A1(n12342), .A2(n11477), .ZN(n11733) );
  NAND2_X1 U14063 ( .A1(n11478), .A2(n15398), .ZN(n11737) );
  NAND2_X1 U14064 ( .A1(n14984), .A2(n14321), .ZN(n11742) );
  NAND2_X1 U14065 ( .A1(n11737), .A2(n11742), .ZN(n14317) );
  INV_X1 U14066 ( .A(n11733), .ZN(n14314) );
  NOR2_X1 U14067 ( .A1(n14317), .A2(n14314), .ZN(n11479) );
  NAND2_X1 U14068 ( .A1(n14309), .A2(n15388), .ZN(n11744) );
  NAND2_X1 U14069 ( .A1(n11592), .A2(n14320), .ZN(n11746) );
  NAND2_X1 U14070 ( .A1(n11744), .A2(n11746), .ZN(n12714) );
  NAND2_X1 U14071 ( .A1(n11480), .A2(n11746), .ZN(n12713) );
  NOR2_X1 U14072 ( .A1(n11593), .A2(n14304), .ZN(n11750) );
  NAND2_X1 U14073 ( .A1(n11593), .A2(n14304), .ZN(n11747) );
  OAI21_X1 U14074 ( .B1(n12713), .B2(n11750), .A(n11747), .ZN(n12706) );
  NAND2_X1 U14075 ( .A1(n12866), .A2(n12719), .ZN(n11753) );
  INV_X1 U14076 ( .A(n11753), .ZN(n11481) );
  OAI21_X1 U14077 ( .B1(n12706), .B2(n11481), .A(n11754), .ZN(n12688) );
  NAND2_X1 U14078 ( .A1(n11601), .A2(n12703), .ZN(n11759) );
  NAND2_X1 U14079 ( .A1(n12688), .A2(n12689), .ZN(n11482) );
  NAND2_X1 U14080 ( .A1(n11482), .A2(n11760), .ZN(n12675) );
  NAND2_X1 U14081 ( .A1(n11483), .A2(n12691), .ZN(n11764) );
  NAND2_X1 U14082 ( .A1(n12850), .A2(n11868), .ZN(n11763) );
  NAND2_X1 U14083 ( .A1(n12675), .A2(n12676), .ZN(n12674) );
  NAND2_X1 U14084 ( .A1(n12674), .A2(n11763), .ZN(n12658) );
  NAND2_X1 U14085 ( .A1(n11484), .A2(n11664), .ZN(n11487) );
  AOI22_X1 U14086 ( .A1(n11493), .A2(n11485), .B1(n11492), .B2(n12465), .ZN(
        n11486) );
  NAND2_X1 U14087 ( .A1(n12847), .A2(n12341), .ZN(n11770) );
  NAND2_X1 U14088 ( .A1(n11775), .A2(n11770), .ZN(n12659) );
  NAND2_X1 U14089 ( .A1(n11488), .A2(n11664), .ZN(n11490) );
  AOI22_X1 U14090 ( .A1(n11493), .A2(SI_18_), .B1(n11492), .B2(n12494), .ZN(
        n11489) );
  NAND2_X1 U14091 ( .A1(n12764), .A2(n12626), .ZN(n11777) );
  OR2_X1 U14092 ( .A1(n11491), .A2(n10001), .ZN(n11495) );
  AOI22_X1 U14093 ( .A1(n11493), .A2(SI_19_), .B1(n11492), .B2(n12489), .ZN(
        n11494) );
  NAND2_X1 U14094 ( .A1(n12835), .A2(n11872), .ZN(n11778) );
  INV_X1 U14095 ( .A(n11778), .ZN(n11496) );
  OR2_X1 U14096 ( .A1(n11662), .A2(n11498), .ZN(n11499) );
  NOR2_X1 U14097 ( .A1(n11502), .A2(n11501), .ZN(n11503) );
  OR2_X1 U14098 ( .A1(n11504), .A2(n11503), .ZN(n12620) );
  NAND2_X1 U14099 ( .A1(n12620), .A2(n11566), .ZN(n11507) );
  NAND2_X1 U14100 ( .A1(n11521), .A2(P3_REG1_REG_20__SCAN_IN), .ZN(n11505) );
  INV_X1 U14101 ( .A(n12614), .ZN(n11508) );
  INV_X1 U14102 ( .A(n12835), .ZN(n12268) );
  INV_X1 U14103 ( .A(n11872), .ZN(n12648) );
  NAND2_X1 U14104 ( .A1(n12268), .A2(n12648), .ZN(n12610) );
  AND2_X1 U14105 ( .A1(n11508), .A2(n12610), .ZN(n11509) );
  OR2_X1 U14106 ( .A1(n12758), .A2(n12627), .ZN(n11784) );
  NAND2_X1 U14107 ( .A1(n11510), .A2(n11664), .ZN(n11513) );
  NAND2_X1 U14108 ( .A1(n12825), .A2(n12615), .ZN(n11788) );
  NAND2_X1 U14109 ( .A1(n11514), .A2(n11787), .ZN(n12588) );
  NAND2_X1 U14110 ( .A1(n11515), .A2(n11664), .ZN(n11517) );
  OR2_X1 U14111 ( .A1(n11662), .A2(n10121), .ZN(n11516) );
  NAND2_X1 U14112 ( .A1(n11518), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n11519) );
  NAND2_X1 U14113 ( .A1(n11520), .A2(n11519), .ZN(n12595) );
  NAND2_X1 U14114 ( .A1(n12595), .A2(n11566), .ZN(n11524) );
  NAND2_X1 U14115 ( .A1(n11521), .A2(P3_REG1_REG_22__SCAN_IN), .ZN(n11522) );
  NAND2_X1 U14116 ( .A1(n12819), .A2(n12577), .ZN(n11792) );
  INV_X1 U14117 ( .A(n11791), .ZN(n11525) );
  NAND2_X1 U14118 ( .A1(n11526), .A2(n11664), .ZN(n11528) );
  OR2_X1 U14119 ( .A1(n11662), .A2(n15291), .ZN(n11527) );
  OR2_X1 U14120 ( .A1(n12584), .A2(n12313), .ZN(n11673) );
  OAI21_X1 U14121 ( .B1(n12573), .B2(n12572), .A(n11673), .ZN(n12564) );
  NAND2_X1 U14122 ( .A1(n11529), .A2(n11664), .ZN(n11532) );
  AND2_X1 U14123 ( .A1(n11533), .A2(P3_REG3_REG_24__SCAN_IN), .ZN(n11534) );
  OR2_X1 U14124 ( .A1(n11534), .A2(n11544), .ZN(n12566) );
  INV_X1 U14125 ( .A(P3_REG1_REG_24__SCAN_IN), .ZN(n11537) );
  NAND2_X1 U14126 ( .A1(n11567), .A2(P3_REG2_REG_24__SCAN_IN), .ZN(n11536) );
  OAI211_X1 U14127 ( .C1(n11537), .C2(n11570), .A(n11536), .B(n11535), .ZN(
        n11538) );
  AOI21_X2 U14128 ( .B1(n12566), .B2(n11566), .A(n11538), .ZN(n12578) );
  OR2_X1 U14129 ( .A1(n12745), .A2(n12578), .ZN(n11674) );
  NAND2_X1 U14130 ( .A1(n12745), .A2(n12578), .ZN(n11675) );
  INV_X1 U14131 ( .A(n11675), .ZN(n11678) );
  NAND2_X1 U14132 ( .A1(n11539), .A2(n11664), .ZN(n11542) );
  OR2_X1 U14133 ( .A1(n11544), .A2(n11543), .ZN(n11545) );
  NAND2_X1 U14134 ( .A1(n11552), .A2(n11545), .ZN(n12556) );
  INV_X1 U14135 ( .A(P3_REG1_REG_25__SCAN_IN), .ZN(n12742) );
  NAND2_X1 U14136 ( .A1(n11567), .A2(P3_REG2_REG_25__SCAN_IN), .ZN(n11546) );
  OAI211_X1 U14137 ( .C1(n12742), .C2(n11570), .A(n11547), .B(n11546), .ZN(
        n11548) );
  AOI21_X2 U14138 ( .B1(n12556), .B2(n11566), .A(n11548), .ZN(n12331) );
  NAND2_X1 U14139 ( .A1(n12807), .A2(n12331), .ZN(n11680) );
  OR2_X1 U14140 ( .A1(n11662), .A2(n11550), .ZN(n11551) );
  NAND2_X1 U14141 ( .A1(n11552), .A2(P3_REG3_REG_26__SCAN_IN), .ZN(n11553) );
  NAND2_X1 U14142 ( .A1(n11563), .A2(n11553), .ZN(n12545) );
  NAND2_X1 U14143 ( .A1(n12545), .A2(n11566), .ZN(n11558) );
  INV_X1 U14144 ( .A(P3_REG1_REG_26__SCAN_IN), .ZN(n12739) );
  NAND2_X1 U14145 ( .A1(n11567), .A2(P3_REG2_REG_26__SCAN_IN), .ZN(n11555) );
  OAI211_X1 U14146 ( .C1(n12739), .C2(n11570), .A(n11555), .B(n11554), .ZN(
        n11556) );
  INV_X1 U14147 ( .A(n11556), .ZN(n11557) );
  NAND2_X1 U14148 ( .A1(n12801), .A2(n12283), .ZN(n11615) );
  INV_X1 U14149 ( .A(n11615), .ZN(n11801) );
  NAND2_X1 U14150 ( .A1(n11890), .A2(n12552), .ZN(n11799) );
  INV_X1 U14151 ( .A(n11562), .ZN(n11565) );
  NAND2_X1 U14152 ( .A1(n11563), .A2(P3_REG3_REG_27__SCAN_IN), .ZN(n11564) );
  NAND2_X1 U14153 ( .A1(n11565), .A2(n11564), .ZN(n12533) );
  NAND2_X1 U14154 ( .A1(n12533), .A2(n11566), .ZN(n11574) );
  INV_X1 U14155 ( .A(P3_REG1_REG_27__SCAN_IN), .ZN(n11571) );
  NAND2_X1 U14156 ( .A1(n11567), .A2(P3_REG2_REG_27__SCAN_IN), .ZN(n11569) );
  OAI211_X1 U14157 ( .C1(n11571), .C2(n11570), .A(n11569), .B(n11568), .ZN(
        n11572) );
  INV_X1 U14158 ( .A(n11572), .ZN(n11573) );
  INV_X1 U14159 ( .A(n11810), .ZN(n11575) );
  XNOR2_X1 U14160 ( .A(n11576), .B(P2_DATAO_REG_28__SCAN_IN), .ZN(n11577) );
  XNOR2_X1 U14161 ( .A(n11578), .B(n11577), .ZN(n12241) );
  NAND2_X1 U14162 ( .A1(n12241), .A2(n11664), .ZN(n11580) );
  OR2_X1 U14163 ( .A1(n11662), .A2(n12243), .ZN(n11579) );
  NAND2_X1 U14164 ( .A1(n12794), .A2(n12250), .ZN(n11812) );
  NAND2_X1 U14165 ( .A1(n11581), .A2(n11664), .ZN(n11584) );
  OR2_X1 U14166 ( .A1(n11662), .A2(n11582), .ZN(n11583) );
  NAND2_X1 U14167 ( .A1(n11917), .A2(n12520), .ZN(n11816) );
  XNOR2_X1 U14168 ( .A(n11670), .B(n11845), .ZN(n11920) );
  INV_X1 U14169 ( .A(n12745), .ZN(n12568) );
  INV_X1 U14170 ( .A(n12584), .ZN(n12813) );
  NAND2_X1 U14171 ( .A1(n14985), .A2(n11730), .ZN(n11732) );
  NAND2_X1 U14172 ( .A1(n11585), .A2(n11732), .ZN(n14983) );
  NAND2_X1 U14173 ( .A1(n14983), .A2(n14982), .ZN(n14981) );
  NAND2_X1 U14174 ( .A1(n12342), .A2(n14988), .ZN(n11586) );
  NAND2_X1 U14175 ( .A1(n14981), .A2(n11586), .ZN(n14318) );
  OAI21_X1 U14176 ( .B1(n14318), .B2(n14984), .A(n15398), .ZN(n11588) );
  NAND2_X1 U14177 ( .A1(n14318), .A2(n14984), .ZN(n11587) );
  NAND2_X1 U14178 ( .A1(n11593), .A2(n11589), .ZN(n11591) );
  AND2_X1 U14179 ( .A1(n12714), .A2(n11591), .ZN(n12698) );
  NAND2_X1 U14180 ( .A1(n11754), .A2(n11753), .ZN(n12707) );
  AND2_X1 U14181 ( .A1(n12698), .A2(n12707), .ZN(n11590) );
  INV_X1 U14182 ( .A(n12707), .ZN(n12701) );
  INV_X1 U14183 ( .A(n11591), .ZN(n11596) );
  NAND2_X1 U14184 ( .A1(n11592), .A2(n15388), .ZN(n12715) );
  INV_X1 U14185 ( .A(n11593), .ZN(n12871) );
  NAND2_X1 U14186 ( .A1(n12871), .A2(n14304), .ZN(n11594) );
  AND2_X1 U14187 ( .A1(n12715), .A2(n11594), .ZN(n11595) );
  OR2_X1 U14188 ( .A1(n12701), .A2(n12699), .ZN(n11599) );
  OR2_X1 U14189 ( .A1(n12866), .A2(n11597), .ZN(n11598) );
  AND2_X1 U14190 ( .A1(n11599), .A2(n11598), .ZN(n11600) );
  NOR2_X1 U14191 ( .A1(n11601), .A2(n12678), .ZN(n11603) );
  NAND2_X1 U14192 ( .A1(n11601), .A2(n12678), .ZN(n11602) );
  OR2_X1 U14193 ( .A1(n12847), .A2(n12679), .ZN(n11605) );
  INV_X1 U14194 ( .A(n11605), .ZN(n11604) );
  NOR2_X1 U14195 ( .A1(n11604), .A2(n12659), .ZN(n11607) );
  OR2_X1 U14196 ( .A1(n12676), .A2(n11607), .ZN(n12640) );
  NAND2_X1 U14197 ( .A1(n12850), .A2(n12691), .ZN(n12661) );
  AND2_X1 U14198 ( .A1(n12661), .A2(n11605), .ZN(n11606) );
  OR2_X1 U14199 ( .A1(n11607), .A2(n11606), .ZN(n12641) );
  AND2_X1 U14200 ( .A1(n12650), .A2(n12641), .ZN(n12642) );
  NAND2_X1 U14201 ( .A1(n12268), .A2(n11872), .ZN(n11608) );
  NAND2_X1 U14202 ( .A1(n11787), .A2(n11788), .ZN(n12601) );
  NAND2_X1 U14203 ( .A1(n12602), .A2(n12601), .ZN(n12600) );
  OR2_X1 U14204 ( .A1(n12825), .A2(n12591), .ZN(n11609) );
  NAND2_X1 U14205 ( .A1(n12600), .A2(n11609), .ZN(n12590) );
  NAND2_X1 U14206 ( .A1(n11791), .A2(n12604), .ZN(n11610) );
  NAND2_X1 U14207 ( .A1(n12590), .A2(n11610), .ZN(n11612) );
  OR2_X1 U14208 ( .A1(n12819), .A2(n12604), .ZN(n11611) );
  NAND2_X1 U14209 ( .A1(n11613), .A2(n11680), .ZN(n12549) );
  INV_X1 U14210 ( .A(n12532), .ZN(n11893) );
  NAND2_X1 U14211 ( .A1(n11893), .A2(n12521), .ZN(n12517) );
  NAND2_X1 U14212 ( .A1(n12794), .A2(n11616), .ZN(n11617) );
  NAND2_X1 U14213 ( .A1(n12515), .A2(n11617), .ZN(n11619) );
  AND2_X1 U14214 ( .A1(n11620), .A2(P3_B_REG_SCAN_IN), .ZN(n11621) );
  NOR2_X1 U14215 ( .A1(n15031), .A2(n11621), .ZN(n12507) );
  NAND2_X1 U14216 ( .A1(n11665), .A2(n12507), .ZN(n11622) );
  MUX2_X1 U14217 ( .A(n11625), .B(n11915), .S(n15096), .Z(n11627) );
  NAND2_X1 U14218 ( .A1(n11917), .A2(n12782), .ZN(n11626) );
  OAI211_X1 U14219 ( .C1(n11920), .C2(n12776), .A(n11627), .B(n11626), .ZN(
        P3_U3488) );
  INV_X1 U14220 ( .A(P3_REG0_REG_0__SCAN_IN), .ZN(n11628) );
  NOR2_X1 U14221 ( .A1(n15085), .A2(n11628), .ZN(n11629) );
  AOI21_X1 U14222 ( .B1(n15085), .B2(n11631), .A(n11629), .ZN(n11630) );
  OAI21_X1 U14223 ( .B1(n11634), .B2(n12867), .A(n11630), .ZN(P3_U3390) );
  NOR2_X2 U14224 ( .A1(n12535), .A2(n15018), .ZN(n15014) );
  INV_X1 U14225 ( .A(n15014), .ZN(n12709) );
  AOI21_X1 U14226 ( .B1(P3_REG3_REG_0__SCAN_IN), .B2(n15055), .A(n11631), .ZN(
        n11632) );
  MUX2_X1 U14227 ( .A(n15205), .B(n11632), .S(n15057), .Z(n11633) );
  OAI21_X1 U14228 ( .B1(n11634), .B2(n12709), .A(n11633), .ZN(P3_U3233) );
  OAI222_X1 U14229 ( .A1(n6535), .A2(n11907), .B1(n11635), .B2(P1_U3086), .C1(
        n11656), .C2(n14266), .ZN(P1_U3325) );
  INV_X1 U14230 ( .A(n11636), .ZN(n13478) );
  OAI222_X1 U14231 ( .A1(n6535), .A2(n13478), .B1(n11637), .B2(P1_U3086), .C1(
        n11644), .C2(n14266), .ZN(P1_U3326) );
  INV_X1 U14232 ( .A(n11638), .ZN(n13482) );
  OAI222_X1 U14233 ( .A1(n11640), .A2(P1_U3086), .B1(n6535), .B2(n13482), .C1(
        n11639), .C2(n14266), .ZN(P1_U3327) );
  INV_X1 U14234 ( .A(SI_30_), .ZN(n11651) );
  INV_X1 U14235 ( .A(n11641), .ZN(n11642) );
  NAND2_X1 U14236 ( .A1(n11643), .A2(n11642), .ZN(n11646) );
  NAND2_X1 U14237 ( .A1(n11644), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n11645) );
  XNOR2_X1 U14238 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(P2_DATAO_REG_30__SCAN_IN), 
        .ZN(n11654) );
  INV_X1 U14239 ( .A(n11654), .ZN(n11647) );
  XNOR2_X1 U14240 ( .A(n11655), .B(n11647), .ZN(n11650) );
  INV_X1 U14241 ( .A(n11650), .ZN(n11648) );
  OAI222_X1 U14242 ( .A1(n11649), .A2(P3_U3151), .B1(n11338), .B2(n11651), 
        .C1(n12245), .C2(n11648), .ZN(P3_U3265) );
  NAND2_X1 U14243 ( .A1(n11650), .A2(n11664), .ZN(n11653) );
  OR2_X1 U14244 ( .A1(n11662), .A2(n11651), .ZN(n11652) );
  AND2_X1 U14245 ( .A1(n12791), .A2(n11665), .ZN(n11819) );
  NAND2_X1 U14246 ( .A1(n11655), .A2(n11654), .ZN(n11658) );
  NAND2_X1 U14247 ( .A1(n11656), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n11657) );
  NAND2_X1 U14248 ( .A1(n11658), .A2(n11657), .ZN(n11661) );
  XNOR2_X1 U14249 ( .A(n11659), .B(P2_DATAO_REG_31__SCAN_IN), .ZN(n11660) );
  XNOR2_X1 U14250 ( .A(n11661), .B(n11660), .ZN(n12882) );
  INV_X1 U14251 ( .A(SI_31_), .ZN(n12878) );
  NOR2_X1 U14252 ( .A1(n11662), .A2(n12878), .ZN(n11663) );
  INV_X1 U14253 ( .A(n12508), .ZN(n11667) );
  AND2_X1 U14254 ( .A1(n12511), .A2(n12508), .ZN(n11821) );
  INV_X1 U14255 ( .A(n11665), .ZN(n11666) );
  NAND2_X1 U14256 ( .A1(n12730), .A2(n11666), .ZN(n11846) );
  NAND2_X1 U14257 ( .A1(n12730), .A2(n11667), .ZN(n11668) );
  NAND3_X1 U14258 ( .A1(n11846), .A2(n11816), .A3(n11668), .ZN(n11669) );
  XNOR2_X1 U14259 ( .A(n11671), .B(n12501), .ZN(n11858) );
  INV_X1 U14260 ( .A(n11672), .ZN(n11857) );
  NAND2_X1 U14261 ( .A1(n11674), .A2(n11673), .ZN(n11676) );
  AND2_X1 U14262 ( .A1(n11676), .A2(n11675), .ZN(n11677) );
  MUX2_X1 U14263 ( .A(n11678), .B(n11677), .S(n11815), .Z(n11679) );
  NOR2_X1 U14264 ( .A1(n11679), .A2(n12549), .ZN(n11798) );
  INV_X1 U14265 ( .A(n11680), .ZN(n11682) );
  MUX2_X1 U14266 ( .A(n11682), .B(n11681), .S(n11811), .Z(n11797) );
  NAND2_X1 U14267 ( .A1(n11685), .A2(n11684), .ZN(n11689) );
  OAI21_X1 U14268 ( .B1(n11689), .B2(n6527), .A(n11815), .ZN(n11687) );
  NAND2_X1 U14269 ( .A1(n11687), .A2(n15025), .ZN(n11693) );
  NAND2_X1 U14270 ( .A1(n11689), .A2(n11688), .ZN(n11690) );
  NAND2_X1 U14271 ( .A1(n11690), .A2(n11811), .ZN(n11691) );
  NAND2_X1 U14272 ( .A1(n11825), .A2(n11691), .ZN(n11692) );
  AOI21_X1 U14273 ( .B1(n11683), .B2(n11693), .A(n11692), .ZN(n11703) );
  NAND2_X1 U14274 ( .A1(n15039), .A2(n15019), .ZN(n11694) );
  NAND2_X1 U14275 ( .A1(n11696), .A2(n11694), .ZN(n11695) );
  AND2_X1 U14276 ( .A1(n11699), .A2(n11695), .ZN(n11701) );
  INV_X1 U14277 ( .A(n11696), .ZN(n11697) );
  AOI21_X1 U14278 ( .B1(n11699), .B2(n11698), .A(n11697), .ZN(n11700) );
  MUX2_X1 U14279 ( .A(n11701), .B(n11700), .S(n11815), .Z(n11702) );
  OAI21_X1 U14280 ( .B1(n11703), .B2(n11702), .A(n11830), .ZN(n11707) );
  MUX2_X1 U14281 ( .A(n11705), .B(n11704), .S(n11815), .Z(n11706) );
  NAND3_X1 U14282 ( .A1(n11707), .A2(n11826), .A3(n11706), .ZN(n11715) );
  NAND2_X1 U14283 ( .A1(n11719), .A2(n11708), .ZN(n11712) );
  NAND2_X1 U14284 ( .A1(n11710), .A2(n11709), .ZN(n11711) );
  MUX2_X1 U14285 ( .A(n11712), .B(n11711), .S(n11811), .Z(n11713) );
  INV_X1 U14286 ( .A(n11713), .ZN(n11714) );
  NAND2_X1 U14287 ( .A1(n11715), .A2(n11714), .ZN(n11716) );
  NAND2_X1 U14288 ( .A1(n11716), .A2(n11827), .ZN(n11722) );
  OAI21_X1 U14289 ( .B1(n11722), .B2(n11718), .A(n11717), .ZN(n11724) );
  INV_X1 U14290 ( .A(n11719), .ZN(n11721) );
  OAI21_X1 U14291 ( .B1(n11722), .B2(n11721), .A(n11720), .ZN(n11723) );
  NAND2_X1 U14292 ( .A1(n12343), .A2(n11725), .ZN(n11726) );
  MUX2_X1 U14293 ( .A(n11727), .B(n11726), .S(n11811), .Z(n11728) );
  OAI211_X1 U14294 ( .C1(n11729), .C2(n11047), .A(n11835), .B(n11728), .ZN(
        n11736) );
  MUX2_X1 U14295 ( .A(n14985), .B(n11730), .S(n11811), .Z(n11731) );
  AOI21_X1 U14296 ( .B1(n11732), .B2(n11731), .A(n14982), .ZN(n11735) );
  NOR2_X1 U14297 ( .A1(n11733), .A2(n11815), .ZN(n11734) );
  AOI21_X1 U14298 ( .B1(n11736), .B2(n11735), .A(n11734), .ZN(n11741) );
  OAI211_X1 U14299 ( .C1(n14317), .C2(n11738), .A(n11746), .B(n11737), .ZN(
        n11739) );
  NAND2_X1 U14300 ( .A1(n11739), .A2(n11815), .ZN(n11740) );
  OAI21_X1 U14301 ( .B1(n11741), .B2(n14317), .A(n11740), .ZN(n11745) );
  AOI21_X1 U14302 ( .B1(n11744), .B2(n11742), .A(n11815), .ZN(n11743) );
  AOI21_X1 U14303 ( .B1(n11745), .B2(n11744), .A(n11743), .ZN(n11749) );
  NOR2_X1 U14304 ( .A1(n11746), .A2(n11815), .ZN(n11748) );
  INV_X1 U14305 ( .A(n11747), .ZN(n11751) );
  OR2_X1 U14306 ( .A1(n11751), .A2(n11750), .ZN(n11837) );
  INV_X1 U14307 ( .A(n11837), .ZN(n12717) );
  MUX2_X1 U14308 ( .A(n11751), .B(n11750), .S(n11811), .Z(n11752) );
  NOR2_X1 U14309 ( .A1(n12707), .A2(n11752), .ZN(n11757) );
  MUX2_X1 U14310 ( .A(n11754), .B(n11753), .S(n11811), .Z(n11755) );
  NAND2_X1 U14311 ( .A1(n12689), .A2(n11755), .ZN(n11756) );
  AOI21_X1 U14312 ( .B1(n11758), .B2(n11757), .A(n11756), .ZN(n11767) );
  NAND2_X1 U14313 ( .A1(n11764), .A2(n11759), .ZN(n11762) );
  NAND2_X1 U14314 ( .A1(n11763), .A2(n11760), .ZN(n11761) );
  MUX2_X1 U14315 ( .A(n11762), .B(n11761), .S(n11811), .Z(n11766) );
  MUX2_X1 U14316 ( .A(n11764), .B(n11763), .S(n11815), .Z(n11765) );
  NAND2_X1 U14317 ( .A1(n11768), .A2(n12662), .ZN(n11776) );
  INV_X1 U14318 ( .A(n11777), .ZN(n11771) );
  OAI211_X1 U14319 ( .C1(n11771), .C2(n11770), .A(n11778), .B(n11769), .ZN(
        n11772) );
  INV_X1 U14320 ( .A(n11772), .ZN(n11773) );
  OAI21_X1 U14321 ( .B1(n11776), .B2(n12650), .A(n11773), .ZN(n11774) );
  NAND2_X1 U14322 ( .A1(n11774), .A2(n12610), .ZN(n11782) );
  AOI21_X1 U14323 ( .B1(n11776), .B2(n11775), .A(n12650), .ZN(n11780) );
  NAND2_X1 U14324 ( .A1(n12610), .A2(n11777), .ZN(n11779) );
  OAI21_X1 U14325 ( .B1(n11780), .B2(n11779), .A(n11778), .ZN(n11781) );
  INV_X1 U14326 ( .A(n12601), .ZN(n12598) );
  NAND2_X1 U14327 ( .A1(n12758), .A2(n12627), .ZN(n11783) );
  MUX2_X1 U14328 ( .A(n11784), .B(n11783), .S(n11815), .Z(n11785) );
  OAI211_X1 U14329 ( .C1(n11786), .C2(n12614), .A(n12598), .B(n11785), .ZN(
        n11790) );
  MUX2_X1 U14330 ( .A(n11788), .B(n11787), .S(n11815), .Z(n11789) );
  MUX2_X1 U14331 ( .A(n11792), .B(n11791), .S(n11811), .Z(n11793) );
  NAND3_X1 U14332 ( .A1(n12584), .A2(n12313), .A3(n11811), .ZN(n11794) );
  NOR2_X1 U14333 ( .A1(n12549), .A2(n12565), .ZN(n11843) );
  NAND2_X1 U14334 ( .A1(n11795), .A2(n11843), .ZN(n11796) );
  INV_X1 U14335 ( .A(n12531), .ZN(n11800) );
  NAND3_X1 U14336 ( .A1(n11805), .A2(n11800), .A3(n11799), .ZN(n11807) );
  NOR2_X1 U14337 ( .A1(n12531), .A2(n11801), .ZN(n11804) );
  INV_X1 U14338 ( .A(n11802), .ZN(n11803) );
  MUX2_X1 U14339 ( .A(n11807), .B(n11806), .S(n11815), .Z(n11808) );
  NAND3_X1 U14340 ( .A1(n11812), .A2(n11811), .A3(n11810), .ZN(n11813) );
  INV_X1 U14341 ( .A(n11816), .ZN(n11818) );
  INV_X1 U14342 ( .A(n11846), .ZN(n11817) );
  INV_X1 U14343 ( .A(n11819), .ZN(n11820) );
  NAND2_X1 U14344 ( .A1(n6645), .A2(n11820), .ZN(n11824) );
  INV_X1 U14345 ( .A(n11821), .ZN(n11847) );
  NOR2_X1 U14346 ( .A1(n11823), .A2(n15050), .ZN(n11856) );
  INV_X1 U14347 ( .A(n11823), .ZN(n11854) );
  INV_X1 U14348 ( .A(n11824), .ZN(n11849) );
  INV_X1 U14349 ( .A(n12587), .ZN(n12589) );
  NAND4_X1 U14350 ( .A1(n11828), .A2(n11827), .A3(n11826), .A4(n11825), .ZN(
        n11833) );
  NAND3_X1 U14351 ( .A1(n11831), .A2(n11830), .A3(n11829), .ZN(n11832) );
  NOR3_X1 U14352 ( .A1(n11833), .A2(n11832), .A3(n14982), .ZN(n11836) );
  NAND4_X1 U14353 ( .A1(n11836), .A2(n11835), .A3(n15025), .A4(n11834), .ZN(
        n11838) );
  NOR4_X1 U14354 ( .A1(n11838), .A2(n11837), .A3(n12714), .A4(n14317), .ZN(
        n11839) );
  AND4_X1 U14355 ( .A1(n12676), .A2(n12701), .A3(n12689), .A4(n11839), .ZN(
        n11840) );
  NAND4_X1 U14356 ( .A1(n12633), .A2(n12646), .A3(n12662), .A4(n11840), .ZN(
        n11841) );
  NOR4_X1 U14357 ( .A1(n12589), .A2(n12601), .A3(n12614), .A4(n11841), .ZN(
        n11842) );
  NAND4_X1 U14358 ( .A1(n12540), .A2(n11843), .A3(n11842), .A4(n12574), .ZN(
        n11844) );
  NOR4_X1 U14359 ( .A1(n11845), .A2(n12516), .A3(n12531), .A4(n11844), .ZN(
        n11848) );
  NAND4_X1 U14360 ( .A1(n11849), .A2(n11848), .A3(n11847), .A4(n11846), .ZN(
        n11850) );
  XNOR2_X1 U14361 ( .A(n11850), .B(n12501), .ZN(n11851) );
  OAI22_X1 U14362 ( .A1(n11854), .A2(n11853), .B1(n11852), .B2(n11851), .ZN(
        n11855) );
  NAND2_X1 U14363 ( .A1(n11860), .A2(n11859), .ZN(n11861) );
  OAI211_X1 U14364 ( .C1(n11862), .C2(n12242), .A(P3_B_REG_SCAN_IN), .B(n11861), .ZN(n11863) );
  OAI21_X1 U14365 ( .B1(n11865), .B2(n11864), .A(n11863), .ZN(P3_U3296) );
  XNOR2_X1 U14366 ( .A(n12758), .B(n11892), .ZN(n11874) );
  INV_X1 U14367 ( .A(n11874), .ZN(n11875) );
  XNOR2_X1 U14368 ( .A(n12835), .B(n11892), .ZN(n11873) );
  XNOR2_X1 U14369 ( .A(n12764), .B(n11892), .ZN(n11870) );
  INV_X1 U14370 ( .A(n11870), .ZN(n11871) );
  XNOR2_X1 U14371 ( .A(n12847), .B(n11892), .ZN(n11869) );
  XNOR2_X1 U14372 ( .A(n11869), .B(n12679), .ZN(n12288) );
  XNOR2_X1 U14373 ( .A(n11870), .B(n12665), .ZN(n12321) );
  XNOR2_X1 U14374 ( .A(n11873), .B(n11872), .ZN(n12265) );
  XNOR2_X1 U14375 ( .A(n11874), .B(n12627), .ZN(n12306) );
  NOR2_X1 U14376 ( .A1(n12305), .A2(n12306), .ZN(n12304) );
  AOI21_X1 U14377 ( .B1(n11875), .B2(n12603), .A(n12304), .ZN(n12272) );
  XNOR2_X1 U14378 ( .A(n12825), .B(n11892), .ZN(n11876) );
  XNOR2_X1 U14379 ( .A(n11876), .B(n12591), .ZN(n12271) );
  NAND2_X1 U14380 ( .A1(n12272), .A2(n12271), .ZN(n12270) );
  XNOR2_X1 U14381 ( .A(n12819), .B(n11892), .ZN(n11879) );
  AOI21_X2 U14382 ( .B1(n12310), .B2(n12577), .A(n11881), .ZN(n11882) );
  XNOR2_X1 U14383 ( .A(n12584), .B(n11892), .ZN(n11884) );
  INV_X1 U14384 ( .A(n11882), .ZN(n11883) );
  XNOR2_X1 U14385 ( .A(n12745), .B(n11892), .ZN(n11885) );
  XNOR2_X1 U14386 ( .A(n11885), .B(n12578), .ZN(n12296) );
  INV_X1 U14387 ( .A(n11885), .ZN(n11886) );
  INV_X1 U14388 ( .A(n12578), .ZN(n12551) );
  XNOR2_X1 U14389 ( .A(n11887), .B(n11892), .ZN(n11888) );
  XNOR2_X1 U14390 ( .A(n11888), .B(n12331), .ZN(n12280) );
  INV_X1 U14391 ( .A(n11888), .ZN(n11889) );
  XNOR2_X1 U14392 ( .A(n11890), .B(n11892), .ZN(n11891) );
  XNOR2_X1 U14393 ( .A(n11891), .B(n12552), .ZN(n12330) );
  XNOR2_X1 U14394 ( .A(n11893), .B(n11892), .ZN(n11894) );
  XNOR2_X1 U14395 ( .A(n11894), .B(n12521), .ZN(n12247) );
  INV_X1 U14396 ( .A(n11894), .ZN(n11895) );
  XOR2_X1 U14397 ( .A(n11892), .B(n12516), .Z(n11896) );
  XNOR2_X1 U14398 ( .A(n11897), .B(n11896), .ZN(n11903) );
  OAI22_X1 U14399 ( .A1(n12521), .A2(n15392), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n11898), .ZN(n11901) );
  INV_X1 U14400 ( .A(n12525), .ZN(n11899) );
  OAI22_X1 U14401 ( .A1(n12520), .A2(n12336), .B1(n11899), .B2(n15395), .ZN(
        n11900) );
  AOI211_X1 U14402 ( .C1(n12794), .C2(n15399), .A(n11901), .B(n11900), .ZN(
        n11902) );
  OAI21_X1 U14403 ( .B1(n11903), .B2(n15401), .A(n11902), .ZN(P3_U3160) );
  OAI222_X1 U14404 ( .A1(n6534), .A2(n11907), .B1(P2_U3088), .B2(n11906), .C1(
        n11905), .C2(n11904), .ZN(P2_U3297) );
  OAI222_X1 U14405 ( .A1(n11904), .A2(n11909), .B1(n6534), .B2(n11908), .C1(
        n13144), .C2(P2_U3088), .ZN(P2_U3308) );
  OAI222_X1 U14406 ( .A1(n11904), .A2(n11911), .B1(n6534), .B2(n11910), .C1(
        n8092), .C2(P2_U3088), .ZN(P2_U3306) );
  NAND2_X1 U14407 ( .A1(n11912), .A2(n6696), .ZN(n11914) );
  AOI22_X1 U14408 ( .A1(n11917), .A2(n15014), .B1(n12506), .B2(n15055), .ZN(
        n11913) );
  OAI211_X1 U14409 ( .C1(n11920), .C2(n12725), .A(n11914), .B(n11913), .ZN(
        P3_U3204) );
  INV_X1 U14410 ( .A(P3_REG0_REG_29__SCAN_IN), .ZN(n11916) );
  MUX2_X1 U14411 ( .A(n11916), .B(n11915), .S(n15085), .Z(n11919) );
  NAND2_X1 U14412 ( .A1(n11917), .A2(n12870), .ZN(n11918) );
  OAI211_X1 U14413 ( .C1(n11920), .C2(n12859), .A(n11919), .B(n11918), .ZN(
        P3_U3456) );
  NAND2_X1 U14414 ( .A1(n11923), .A2(n11922), .ZN(n11937) );
  INV_X1 U14415 ( .A(n11924), .ZN(n11927) );
  NAND2_X1 U14416 ( .A1(n13167), .A2(n11925), .ZN(n11926) );
  AND2_X1 U14417 ( .A1(n11927), .A2(n11926), .ZN(n11938) );
  NAND2_X1 U14418 ( .A1(n11937), .A2(n11938), .ZN(n11929) );
  NAND3_X4 U14419 ( .A1(n12152), .A2(n11927), .A3(n12180), .ZN(n12090) );
  NAND2_X1 U14420 ( .A1(n11929), .A2(n7446), .ZN(n11943) );
  NAND2_X1 U14421 ( .A1(n12090), .A2(n11932), .ZN(n11930) );
  AND2_X1 U14422 ( .A1(n11931), .A2(n11930), .ZN(n11950) );
  NAND2_X1 U14423 ( .A1(n11977), .A2(n11932), .ZN(n11933) );
  NAND2_X1 U14424 ( .A1(n11934), .A2(n11933), .ZN(n11949) );
  NAND2_X1 U14425 ( .A1(n11950), .A2(n11949), .ZN(n11942) );
  NAND2_X1 U14426 ( .A1(n6532), .A2(n11935), .ZN(n11936) );
  INV_X1 U14427 ( .A(n11937), .ZN(n11940) );
  INV_X1 U14428 ( .A(n11938), .ZN(n11939) );
  NAND2_X1 U14429 ( .A1(n11940), .A2(n11939), .ZN(n11941) );
  NAND4_X1 U14430 ( .A1(n11943), .A2(n11942), .A3(n11936), .A4(n11941), .ZN(
        n11955) );
  NAND2_X1 U14431 ( .A1(n13050), .A2(n12090), .ZN(n11945) );
  NAND2_X1 U14432 ( .A1(n6532), .A2(n6524), .ZN(n11944) );
  NAND2_X1 U14433 ( .A1(n13050), .A2(n6532), .ZN(n11948) );
  NAND2_X1 U14434 ( .A1(n6524), .A2(n12090), .ZN(n11947) );
  NAND2_X1 U14435 ( .A1(n11948), .A2(n11947), .ZN(n11956) );
  NAND2_X1 U14436 ( .A1(n11957), .A2(n11956), .ZN(n11954) );
  INV_X1 U14437 ( .A(n11949), .ZN(n11952) );
  INV_X1 U14438 ( .A(n11950), .ZN(n11951) );
  NAND2_X1 U14439 ( .A1(n11952), .A2(n11951), .ZN(n11953) );
  NAND3_X1 U14440 ( .A1(n11955), .A2(n11954), .A3(n11953), .ZN(n11961) );
  INV_X1 U14441 ( .A(n11956), .ZN(n11959) );
  INV_X1 U14442 ( .A(n11957), .ZN(n11958) );
  NAND2_X1 U14443 ( .A1(n11959), .A2(n11958), .ZN(n11960) );
  NAND2_X1 U14444 ( .A1(n11961), .A2(n11960), .ZN(n11969) );
  INV_X1 U14445 ( .A(n11977), .ZN(n12023) );
  INV_X1 U14446 ( .A(n12023), .ZN(n11964) );
  NAND2_X1 U14447 ( .A1(n11965), .A2(n12137), .ZN(n11963) );
  NAND2_X1 U14448 ( .A1(n13049), .A2(n12090), .ZN(n11962) );
  NAND2_X1 U14449 ( .A1(n11963), .A2(n11962), .ZN(n11968) );
  AOI22_X1 U14450 ( .A1(n11965), .A2(n12090), .B1(n11964), .B2(n13049), .ZN(
        n11966) );
  AOI21_X1 U14451 ( .B1(n11969), .B2(n11968), .A(n11966), .ZN(n11967) );
  NOR2_X1 U14452 ( .A1(n11969), .A2(n11968), .ZN(n11970) );
  NAND2_X1 U14453 ( .A1(n11973), .A2(n12090), .ZN(n11972) );
  NAND2_X1 U14454 ( .A1(n13048), .A2(n6525), .ZN(n11971) );
  NAND2_X1 U14455 ( .A1(n11973), .A2(n6526), .ZN(n11974) );
  OAI21_X1 U14456 ( .B1(n11975), .B2(n12149), .A(n11974), .ZN(n11976) );
  NAND2_X1 U14457 ( .A1(n11980), .A2(n11964), .ZN(n11979) );
  NAND2_X1 U14458 ( .A1(n13047), .A2(n12157), .ZN(n11978) );
  NAND2_X1 U14459 ( .A1(n11979), .A2(n11978), .ZN(n11983) );
  AOI22_X1 U14460 ( .A1(n11980), .A2(n12157), .B1(n11964), .B2(n13047), .ZN(
        n11981) );
  AOI21_X1 U14461 ( .B1(n11984), .B2(n11983), .A(n11981), .ZN(n11982) );
  INV_X1 U14462 ( .A(n11982), .ZN(n11985) );
  NAND2_X1 U14463 ( .A1(n14782), .A2(n12157), .ZN(n11987) );
  NAND2_X1 U14464 ( .A1(n13046), .A2(n11964), .ZN(n11986) );
  AOI22_X1 U14465 ( .A1(n14782), .A2(n6525), .B1(n13046), .B2(n12157), .ZN(
        n11988) );
  NAND2_X1 U14466 ( .A1(n14788), .A2(n11964), .ZN(n11990) );
  NAND2_X1 U14467 ( .A1(n13045), .A2(n12157), .ZN(n11989) );
  NAND2_X1 U14468 ( .A1(n11990), .A2(n11989), .ZN(n11995) );
  NAND2_X1 U14469 ( .A1(n14788), .A2(n12090), .ZN(n11991) );
  OAI21_X1 U14470 ( .B1(n11992), .B2(n12023), .A(n11991), .ZN(n11993) );
  NAND2_X1 U14471 ( .A1(n14795), .A2(n12090), .ZN(n11998) );
  NAND2_X1 U14472 ( .A1(n13044), .A2(n12137), .ZN(n11997) );
  NAND2_X1 U14473 ( .A1(n11998), .A2(n11997), .ZN(n12000) );
  AOI22_X1 U14474 ( .A1(n14795), .A2(n6525), .B1(n13044), .B2(n12157), .ZN(
        n11999) );
  AOI21_X1 U14475 ( .B1(n12001), .B2(n12000), .A(n11999), .ZN(n12003) );
  NAND2_X1 U14476 ( .A1(n12008), .A2(n6525), .ZN(n12005) );
  NAND2_X1 U14477 ( .A1(n13042), .A2(n12157), .ZN(n12004) );
  NAND2_X1 U14478 ( .A1(n12005), .A2(n12004), .ZN(n12006) );
  OR2_X1 U14479 ( .A1(n12007), .A2(n12006), .ZN(n12014) );
  NAND2_X1 U14480 ( .A1(n12007), .A2(n12006), .ZN(n12012) );
  NAND2_X1 U14481 ( .A1(n12008), .A2(n12157), .ZN(n12010) );
  NAND2_X1 U14482 ( .A1(n13042), .A2(n12137), .ZN(n12009) );
  NAND2_X1 U14483 ( .A1(n12010), .A2(n12009), .ZN(n12011) );
  NAND2_X1 U14484 ( .A1(n12012), .A2(n12011), .ZN(n12013) );
  NAND2_X1 U14485 ( .A1(n12014), .A2(n12013), .ZN(n12018) );
  NAND2_X1 U14486 ( .A1(n14811), .A2(n12090), .ZN(n12016) );
  NAND2_X1 U14487 ( .A1(n13041), .A2(n11964), .ZN(n12015) );
  AOI22_X1 U14488 ( .A1(n14811), .A2(n6525), .B1(n13041), .B2(n12157), .ZN(
        n12017) );
  NAND2_X1 U14489 ( .A1(n12021), .A2(n11964), .ZN(n12020) );
  NAND2_X1 U14490 ( .A1(n13040), .A2(n12090), .ZN(n12019) );
  NAND2_X1 U14491 ( .A1(n12021), .A2(n12157), .ZN(n12022) );
  OAI21_X1 U14492 ( .B1(n12024), .B2(n12023), .A(n12022), .ZN(n12025) );
  NAND2_X1 U14493 ( .A1(n14379), .A2(n12157), .ZN(n12027) );
  NAND2_X1 U14494 ( .A1(n13039), .A2(n12137), .ZN(n12026) );
  NAND2_X1 U14495 ( .A1(n12027), .A2(n12026), .ZN(n12029) );
  AOI22_X1 U14496 ( .A1(n14379), .A2(n6526), .B1(n13039), .B2(n12157), .ZN(
        n12028) );
  NAND2_X1 U14497 ( .A1(n12032), .A2(n6526), .ZN(n12031) );
  NAND2_X1 U14498 ( .A1(n14335), .A2(n12090), .ZN(n12030) );
  NAND2_X1 U14499 ( .A1(n12031), .A2(n12030), .ZN(n12038) );
  NAND2_X1 U14500 ( .A1(n12037), .A2(n12038), .ZN(n12036) );
  NAND2_X1 U14501 ( .A1(n12032), .A2(n12090), .ZN(n12033) );
  OAI21_X1 U14502 ( .B1(n12034), .B2(n12023), .A(n12033), .ZN(n12035) );
  NAND2_X1 U14503 ( .A1(n12036), .A2(n12035), .ZN(n12042) );
  NAND2_X1 U14504 ( .A1(n12040), .A2(n12039), .ZN(n12041) );
  NAND2_X1 U14505 ( .A1(n12042), .A2(n12041), .ZN(n12047) );
  NAND2_X1 U14506 ( .A1(n14356), .A2(n12157), .ZN(n12044) );
  NAND2_X1 U14507 ( .A1(n13038), .A2(n12137), .ZN(n12043) );
  NAND2_X1 U14508 ( .A1(n12044), .A2(n12043), .ZN(n12046) );
  AOI22_X1 U14509 ( .A1(n14356), .A2(n11964), .B1(n13038), .B2(n12157), .ZN(
        n12045) );
  NAND2_X1 U14510 ( .A1(n12050), .A2(n6526), .ZN(n12049) );
  NAND2_X1 U14511 ( .A1(n14337), .A2(n12090), .ZN(n12048) );
  NAND2_X1 U14512 ( .A1(n12049), .A2(n12048), .ZN(n12053) );
  AOI22_X1 U14513 ( .A1(n12050), .A2(n12157), .B1(n12137), .B2(n14337), .ZN(
        n12051) );
  INV_X1 U14514 ( .A(n12052), .ZN(n12055) );
  NAND2_X1 U14515 ( .A1(n13426), .A2(n12090), .ZN(n12057) );
  NAND2_X1 U14516 ( .A1(n13037), .A2(n6525), .ZN(n12056) );
  NAND2_X1 U14517 ( .A1(n12057), .A2(n12056), .ZN(n12062) );
  NAND2_X1 U14518 ( .A1(n13426), .A2(n11964), .ZN(n12058) );
  OAI21_X1 U14519 ( .B1(n12059), .B2(n12149), .A(n12058), .ZN(n12060) );
  NAND2_X1 U14520 ( .A1(n12065), .A2(n12137), .ZN(n12064) );
  NAND2_X1 U14521 ( .A1(n13036), .A2(n12157), .ZN(n12063) );
  NAND2_X1 U14522 ( .A1(n12064), .A2(n12063), .ZN(n12067) );
  AOI22_X1 U14523 ( .A1(n12065), .A2(n12157), .B1(n6526), .B2(n13036), .ZN(
        n12066) );
  NAND2_X1 U14524 ( .A1(n6523), .A2(n12090), .ZN(n12069) );
  NAND2_X1 U14525 ( .A1(n13035), .A2(n12137), .ZN(n12068) );
  NAND2_X1 U14526 ( .A1(n12069), .A2(n12068), .ZN(n12075) );
  NAND2_X1 U14527 ( .A1(n12074), .A2(n12075), .ZN(n12073) );
  NAND2_X1 U14528 ( .A1(n6523), .A2(n12137), .ZN(n12071) );
  NAND2_X1 U14529 ( .A1(n13035), .A2(n12090), .ZN(n12070) );
  NAND2_X1 U14530 ( .A1(n12071), .A2(n12070), .ZN(n12072) );
  INV_X1 U14531 ( .A(n12074), .ZN(n12077) );
  INV_X1 U14532 ( .A(n12075), .ZN(n12076) );
  NAND2_X1 U14533 ( .A1(n12077), .A2(n12076), .ZN(n12078) );
  NAND2_X1 U14534 ( .A1(n13406), .A2(n6526), .ZN(n12080) );
  NAND2_X1 U14535 ( .A1(n13034), .A2(n12157), .ZN(n12079) );
  AOI22_X1 U14536 ( .A1(n13406), .A2(n12090), .B1(n6532), .B2(n13034), .ZN(
        n12081) );
  NAND2_X1 U14537 ( .A1(n13402), .A2(n12157), .ZN(n12083) );
  NAND2_X1 U14538 ( .A1(n13033), .A2(n6532), .ZN(n12082) );
  NAND2_X1 U14539 ( .A1(n12083), .A2(n12082), .ZN(n12087) );
  NAND2_X1 U14540 ( .A1(n13402), .A2(n6526), .ZN(n12085) );
  NAND2_X1 U14541 ( .A1(n13033), .A2(n12157), .ZN(n12084) );
  NAND2_X1 U14542 ( .A1(n13459), .A2(n11964), .ZN(n12089) );
  NAND2_X1 U14543 ( .A1(n13032), .A2(n12157), .ZN(n12088) );
  AOI22_X1 U14544 ( .A1(n13459), .A2(n12090), .B1(n6525), .B2(n13032), .ZN(
        n12091) );
  NAND2_X1 U14545 ( .A1(n13263), .A2(n12090), .ZN(n12093) );
  NAND2_X1 U14546 ( .A1(n13031), .A2(n6532), .ZN(n12092) );
  NAND2_X1 U14547 ( .A1(n12093), .A2(n12092), .ZN(n12095) );
  AOI22_X1 U14548 ( .A1(n13263), .A2(n12137), .B1(n13031), .B2(n12090), .ZN(
        n12094) );
  AOI21_X1 U14549 ( .B1(n12096), .B2(n12095), .A(n12094), .ZN(n12098) );
  NOR2_X1 U14550 ( .A1(n12096), .A2(n12095), .ZN(n12097) );
  NAND2_X1 U14551 ( .A1(n13385), .A2(n11977), .ZN(n12100) );
  NAND2_X1 U14552 ( .A1(n13030), .A2(n12157), .ZN(n12099) );
  NAND2_X1 U14553 ( .A1(n12100), .A2(n12099), .ZN(n12109) );
  AND2_X1 U14554 ( .A1(n13028), .A2(n12157), .ZN(n12101) );
  AOI21_X1 U14555 ( .B1(n13375), .B2(n6526), .A(n12101), .ZN(n12119) );
  NAND2_X1 U14556 ( .A1(n13375), .A2(n12157), .ZN(n12103) );
  NAND2_X1 U14557 ( .A1(n13028), .A2(n11977), .ZN(n12102) );
  NAND2_X1 U14558 ( .A1(n12103), .A2(n12102), .ZN(n12118) );
  NAND2_X1 U14559 ( .A1(n12119), .A2(n12118), .ZN(n12123) );
  AND2_X1 U14560 ( .A1(n13029), .A2(n12157), .ZN(n12104) );
  AOI21_X1 U14561 ( .B1(n13233), .B2(n11964), .A(n12104), .ZN(n12115) );
  NAND2_X1 U14562 ( .A1(n13233), .A2(n12157), .ZN(n12106) );
  NAND2_X1 U14563 ( .A1(n13029), .A2(n12137), .ZN(n12105) );
  NAND2_X1 U14564 ( .A1(n12106), .A2(n12105), .ZN(n12114) );
  NAND2_X1 U14565 ( .A1(n12115), .A2(n12114), .ZN(n12107) );
  OAI211_X1 U14566 ( .C1(n12110), .C2(n12109), .A(n12123), .B(n12107), .ZN(
        n12127) );
  AOI22_X1 U14567 ( .A1(n13385), .A2(n12157), .B1(n12137), .B2(n13030), .ZN(
        n12108) );
  AOI21_X1 U14568 ( .B1(n12110), .B2(n12109), .A(n12108), .ZN(n12126) );
  AND2_X1 U14569 ( .A1(n13027), .A2(n6525), .ZN(n12111) );
  AOI21_X1 U14570 ( .B1(n13205), .B2(n12090), .A(n12111), .ZN(n12141) );
  NAND2_X1 U14571 ( .A1(n13205), .A2(n6526), .ZN(n12113) );
  NAND2_X1 U14572 ( .A1(n13027), .A2(n12157), .ZN(n12112) );
  NAND2_X1 U14573 ( .A1(n12113), .A2(n12112), .ZN(n12140) );
  NAND2_X1 U14574 ( .A1(n12141), .A2(n12140), .ZN(n12125) );
  INV_X1 U14575 ( .A(n12114), .ZN(n12117) );
  INV_X1 U14576 ( .A(n12115), .ZN(n12116) );
  AND2_X1 U14577 ( .A1(n12117), .A2(n12116), .ZN(n12122) );
  INV_X1 U14578 ( .A(n12118), .ZN(n12121) );
  INV_X1 U14579 ( .A(n12119), .ZN(n12120) );
  AOI22_X1 U14580 ( .A1(n12123), .A2(n12122), .B1(n12121), .B2(n12120), .ZN(
        n12124) );
  OAI21_X1 U14581 ( .B1(n12127), .B2(n12126), .A(n7447), .ZN(n12145) );
  AND2_X1 U14582 ( .A1(n13024), .A2(n12157), .ZN(n12128) );
  AOI21_X1 U14583 ( .B1(n13351), .B2(n11977), .A(n12128), .ZN(n12161) );
  NAND2_X1 U14584 ( .A1(n13351), .A2(n12157), .ZN(n12130) );
  NAND2_X1 U14585 ( .A1(n13024), .A2(n6526), .ZN(n12129) );
  NAND2_X1 U14586 ( .A1(n12130), .A2(n12129), .ZN(n12160) );
  NAND2_X1 U14587 ( .A1(n12161), .A2(n12160), .ZN(n12167) );
  AND2_X1 U14588 ( .A1(n13025), .A2(n12090), .ZN(n12131) );
  AOI21_X1 U14589 ( .B1(n13356), .B2(n11977), .A(n12131), .ZN(n12165) );
  NAND2_X1 U14590 ( .A1(n13356), .A2(n12157), .ZN(n12133) );
  NAND2_X1 U14591 ( .A1(n13025), .A2(n12137), .ZN(n12132) );
  NAND2_X1 U14592 ( .A1(n12133), .A2(n12132), .ZN(n12164) );
  NAND2_X1 U14593 ( .A1(n12165), .A2(n12164), .ZN(n12134) );
  AND2_X1 U14594 ( .A1(n12167), .A2(n12134), .ZN(n12135) );
  AND2_X1 U14595 ( .A1(n13026), .A2(n12157), .ZN(n12136) );
  AOI21_X1 U14596 ( .B1(n13187), .B2(n6526), .A(n12136), .ZN(n12147) );
  NAND2_X1 U14597 ( .A1(n13187), .A2(n12090), .ZN(n12139) );
  NAND2_X1 U14598 ( .A1(n13026), .A2(n6526), .ZN(n12138) );
  NAND2_X1 U14599 ( .A1(n12139), .A2(n12138), .ZN(n12146) );
  INV_X1 U14600 ( .A(n12140), .ZN(n12143) );
  INV_X1 U14601 ( .A(n12141), .ZN(n12142) );
  AOI22_X1 U14602 ( .A1(n12147), .A2(n12146), .B1(n12143), .B2(n12142), .ZN(
        n12144) );
  MUX2_X1 U14603 ( .A(n13022), .B(n12149), .S(n12174), .Z(n12151) );
  NAND2_X1 U14604 ( .A1(n6526), .A2(n13022), .ZN(n12150) );
  NAND2_X1 U14605 ( .A1(n12151), .A2(n12150), .ZN(n12163) );
  NAND2_X1 U14606 ( .A1(n13022), .A2(n12157), .ZN(n12175) );
  INV_X1 U14607 ( .A(n8092), .ZN(n12226) );
  OAI211_X1 U14608 ( .C1(n12152), .C2(n12230), .A(n12226), .B(n12180), .ZN(
        n12153) );
  INV_X1 U14609 ( .A(n12153), .ZN(n12155) );
  AOI21_X1 U14610 ( .B1(n12175), .B2(n12155), .A(n12154), .ZN(n12156) );
  AOI21_X1 U14611 ( .B1(n13159), .B2(n11977), .A(n12156), .ZN(n12172) );
  NAND2_X1 U14612 ( .A1(n13159), .A2(n12157), .ZN(n12159) );
  NAND2_X1 U14613 ( .A1(n12137), .A2(n13023), .ZN(n12158) );
  NAND2_X1 U14614 ( .A1(n12159), .A2(n12158), .ZN(n12171) );
  OAI22_X1 U14615 ( .A1(n12172), .A2(n12171), .B1(n12161), .B2(n12160), .ZN(
        n12162) );
  NAND2_X1 U14616 ( .A1(n12163), .A2(n12162), .ZN(n12170) );
  INV_X1 U14617 ( .A(n12164), .ZN(n12168) );
  INV_X1 U14618 ( .A(n12165), .ZN(n12166) );
  NAND4_X1 U14619 ( .A1(n12186), .A2(n12168), .A3(n12167), .A4(n12166), .ZN(
        n12169) );
  NAND2_X1 U14620 ( .A1(n12172), .A2(n12171), .ZN(n12173) );
  MUX2_X1 U14621 ( .A(n13022), .B(n12023), .S(n12174), .Z(n12176) );
  NAND2_X1 U14622 ( .A1(n12176), .A2(n12175), .ZN(n12177) );
  INV_X1 U14623 ( .A(n12231), .ZN(n12182) );
  OAI211_X1 U14624 ( .C1(n13167), .C2(n8092), .A(n8093), .B(n12180), .ZN(
        n12181) );
  NAND2_X1 U14625 ( .A1(n12182), .A2(n12181), .ZN(n12234) );
  MUX2_X1 U14626 ( .A(n12226), .B(n8153), .S(n12183), .Z(n12184) );
  INV_X1 U14627 ( .A(n12184), .ZN(n12185) );
  NOR2_X1 U14628 ( .A1(n12185), .A2(n13144), .ZN(n12228) );
  INV_X1 U14629 ( .A(n12186), .ZN(n12225) );
  XNOR2_X1 U14630 ( .A(n13159), .B(n13023), .ZN(n12222) );
  NAND2_X1 U14631 ( .A1(n12188), .A2(n12187), .ZN(n13196) );
  XNOR2_X1 U14632 ( .A(n13406), .B(n12189), .ZN(n13302) );
  NAND4_X1 U14633 ( .A1(n12192), .A2(n12191), .A3(n12190), .A4(n12230), .ZN(
        n12193) );
  NOR2_X1 U14634 ( .A1(n12194), .A2(n12193), .ZN(n12197) );
  NAND4_X1 U14635 ( .A1(n12198), .A2(n12197), .A3(n12196), .A4(n12195), .ZN(
        n12199) );
  NOR2_X1 U14636 ( .A1(n12200), .A2(n12199), .ZN(n12203) );
  NAND4_X1 U14637 ( .A1(n12204), .A2(n12203), .A3(n12202), .A4(n12201), .ZN(
        n12205) );
  OR4_X1 U14638 ( .A1(n12208), .A2(n12207), .A3(n12206), .A4(n12205), .ZN(
        n12209) );
  NOR2_X1 U14639 ( .A1(n14358), .A2(n12209), .ZN(n12212) );
  NAND4_X1 U14640 ( .A1(n12213), .A2(n12212), .A3(n12211), .A4(n12210), .ZN(
        n12214) );
  OR4_X1 U14641 ( .A1(n13270), .A2(n13334), .A3(n13289), .A4(n12214), .ZN(
        n12215) );
  NOR2_X1 U14642 ( .A1(n13302), .A2(n12215), .ZN(n12218) );
  NAND2_X1 U14643 ( .A1(n12217), .A2(n12216), .ZN(n13239) );
  NAND4_X1 U14644 ( .A1(n13224), .A2(n12218), .A3(n13250), .A4(n13239), .ZN(
        n12219) );
  OR3_X1 U14645 ( .A1(n13196), .A2(n13211), .A3(n12219), .ZN(n12220) );
  NOR2_X1 U14646 ( .A1(n13161), .A2(n12220), .ZN(n12221) );
  NAND3_X1 U14647 ( .A1(n12222), .A2(n12221), .A3(n13181), .ZN(n12223) );
  AOI21_X1 U14648 ( .B1(n12231), .B2(n12228), .A(n12227), .ZN(n12233) );
  OAI21_X1 U14649 ( .B1(n12231), .B2(n12230), .A(n7437), .ZN(n12232) );
  INV_X1 U14650 ( .A(n13484), .ZN(n12236) );
  NAND4_X1 U14651 ( .A1(n14334), .A2(n12236), .A3(n14773), .A4(n12235), .ZN(
        n12237) );
  OAI211_X1 U14652 ( .C1(n8153), .C2(n12239), .A(n12237), .B(P2_B_REG_SCAN_IN), 
        .ZN(n12238) );
  OAI21_X1 U14653 ( .B1(n12240), .B2(n12239), .A(n12238), .ZN(P2_U3328) );
  INV_X1 U14654 ( .A(n12241), .ZN(n12244) );
  OAI222_X1 U14655 ( .A1(n12245), .A2(n12244), .B1(n11338), .B2(n12243), .C1(
        P3_U3151), .C2(n12242), .ZN(P3_U3267) );
  XOR2_X1 U14656 ( .A(n12247), .B(n12246), .Z(n12253) );
  AOI22_X1 U14657 ( .A1(n12552), .A2(n12332), .B1(P3_REG3_REG_27__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12249) );
  NAND2_X1 U14658 ( .A1(n12533), .A2(n12333), .ZN(n12248) );
  OAI211_X1 U14659 ( .C1(n12250), .C2(n12336), .A(n12249), .B(n12248), .ZN(
        n12251) );
  AOI21_X1 U14660 ( .B1(n12532), .B2(n12338), .A(n12251), .ZN(n12252) );
  OAI21_X1 U14661 ( .B1(n12253), .B2(n15401), .A(n12252), .ZN(P3_U3154) );
  XNOR2_X1 U14662 ( .A(n12254), .B(n12592), .ZN(n12259) );
  AOI22_X1 U14663 ( .A1(n12551), .A2(n15389), .B1(P3_REG3_REG_23__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12256) );
  NAND2_X1 U14664 ( .A1(n12333), .A2(n12583), .ZN(n12255) );
  OAI211_X1 U14665 ( .C1(n12577), .C2(n15392), .A(n12256), .B(n12255), .ZN(
        n12257) );
  AOI21_X1 U14666 ( .B1(n12584), .B2(n12338), .A(n12257), .ZN(n12258) );
  OAI21_X1 U14667 ( .B1(n12259), .B2(n15401), .A(n12258), .ZN(P3_U3156) );
  INV_X1 U14668 ( .A(n12260), .ZN(n12635) );
  INV_X1 U14669 ( .A(P3_REG3_REG_19__SCAN_IN), .ZN(n15353) );
  NOR2_X1 U14670 ( .A1(n15353), .A2(P3_STATE_REG_SCAN_IN), .ZN(n12499) );
  NOR2_X1 U14671 ( .A1(n15392), .A2(n12626), .ZN(n12261) );
  AOI211_X1 U14672 ( .C1(n15389), .C2(n12603), .A(n12499), .B(n12261), .ZN(
        n12262) );
  OAI21_X1 U14673 ( .B1(n12635), .B2(n15395), .A(n12262), .ZN(n12267) );
  AOI211_X1 U14674 ( .C1(n12265), .C2(n12264), .A(n15401), .B(n12263), .ZN(
        n12266) );
  AOI211_X1 U14675 ( .C1(n15399), .C2(n12268), .A(n12267), .B(n12266), .ZN(
        n12269) );
  INV_X1 U14676 ( .A(n12269), .ZN(P3_U3159) );
  INV_X1 U14677 ( .A(n12825), .ZN(n12278) );
  OAI21_X1 U14678 ( .B1(n12272), .B2(n12271), .A(n12270), .ZN(n12273) );
  NAND2_X1 U14679 ( .A1(n12273), .A2(n12318), .ZN(n12277) );
  AOI22_X1 U14680 ( .A1(n12603), .A2(n12332), .B1(P3_REG3_REG_21__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12274) );
  OAI21_X1 U14681 ( .B1(n12577), .B2(n12336), .A(n12274), .ZN(n12275) );
  AOI21_X1 U14682 ( .B1(n12607), .B2(n12333), .A(n12275), .ZN(n12276) );
  OAI211_X1 U14683 ( .C1(n12278), .C2(n12327), .A(n12277), .B(n12276), .ZN(
        P3_U3163) );
  XOR2_X1 U14684 ( .A(n12280), .B(n12279), .Z(n12286) );
  AOI22_X1 U14685 ( .A1(n12551), .A2(n12332), .B1(P3_REG3_REG_25__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12282) );
  NAND2_X1 U14686 ( .A1(n12333), .A2(n12556), .ZN(n12281) );
  OAI211_X1 U14687 ( .C1(n12283), .C2(n12336), .A(n12282), .B(n12281), .ZN(
        n12284) );
  AOI21_X1 U14688 ( .B1(n12807), .B2(n12338), .A(n12284), .ZN(n12285) );
  OAI21_X1 U14689 ( .B1(n12286), .B2(n15401), .A(n12285), .ZN(P3_U3165) );
  OAI211_X1 U14690 ( .C1(n12289), .C2(n12288), .A(n12287), .B(n12318), .ZN(
        n12294) );
  INV_X1 U14691 ( .A(n12290), .ZN(n12669) );
  NAND2_X1 U14692 ( .A1(n12332), .A2(n12691), .ZN(n12291) );
  NAND2_X1 U14693 ( .A1(P3_U3151), .A2(P3_REG3_REG_17__SCAN_IN), .ZN(n12444)
         );
  OAI211_X1 U14694 ( .C1(n12626), .C2(n12336), .A(n12291), .B(n12444), .ZN(
        n12292) );
  AOI21_X1 U14695 ( .B1(n12333), .B2(n12669), .A(n12292), .ZN(n12293) );
  OAI211_X1 U14696 ( .C1(n12327), .C2(n12847), .A(n12294), .B(n12293), .ZN(
        P3_U3168) );
  XOR2_X1 U14697 ( .A(n12296), .B(n12295), .Z(n12301) );
  AOI22_X1 U14698 ( .A1(n12592), .A2(n12332), .B1(P3_REG3_REG_24__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12298) );
  NAND2_X1 U14699 ( .A1(n12333), .A2(n12566), .ZN(n12297) );
  OAI211_X1 U14700 ( .C1(n12331), .C2(n12336), .A(n12298), .B(n12297), .ZN(
        n12299) );
  AOI21_X1 U14701 ( .B1(n12745), .B2(n12338), .A(n12299), .ZN(n12300) );
  OAI21_X1 U14702 ( .B1(n12301), .B2(n15401), .A(n12300), .ZN(P3_U3169) );
  NAND2_X1 U14703 ( .A1(n12333), .A2(n12620), .ZN(n12303) );
  AOI22_X1 U14704 ( .A1(n12591), .A2(n15389), .B1(P3_REG3_REG_20__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12302) );
  OAI211_X1 U14705 ( .C1(n12648), .C2(n15392), .A(n12303), .B(n12302), .ZN(
        n12308) );
  AOI211_X1 U14706 ( .C1(n12306), .C2(n12305), .A(n15401), .B(n12304), .ZN(
        n12307) );
  AOI211_X1 U14707 ( .C1(n15399), .C2(n12758), .A(n12308), .B(n12307), .ZN(
        n12309) );
  INV_X1 U14708 ( .A(n12309), .ZN(P3_U3173) );
  XNOR2_X1 U14709 ( .A(n12310), .B(n12604), .ZN(n12316) );
  NAND2_X1 U14710 ( .A1(n12333), .A2(n12595), .ZN(n12312) );
  AOI22_X1 U14711 ( .A1(n12591), .A2(n12332), .B1(P3_REG3_REG_22__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12311) );
  OAI211_X1 U14712 ( .C1(n12313), .C2(n12336), .A(n12312), .B(n12311), .ZN(
        n12314) );
  AOI21_X1 U14713 ( .B1(n12819), .B2(n12338), .A(n12314), .ZN(n12315) );
  OAI21_X1 U14714 ( .B1(n12316), .B2(n15401), .A(n12315), .ZN(P3_U3175) );
  INV_X1 U14715 ( .A(n12764), .ZN(n12328) );
  INV_X1 U14716 ( .A(n12317), .ZN(n12319) );
  OAI211_X1 U14717 ( .C1(n12321), .C2(n12320), .A(n12319), .B(n12318), .ZN(
        n12326) );
  NAND2_X1 U14718 ( .A1(n12332), .A2(n12341), .ZN(n12323) );
  NAND2_X1 U14719 ( .A1(P3_U3151), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n12462)
         );
  OAI211_X1 U14720 ( .C1(n12648), .C2(n12336), .A(n12323), .B(n12462), .ZN(
        n12324) );
  AOI21_X1 U14721 ( .B1(n12333), .B2(n12653), .A(n12324), .ZN(n12325) );
  OAI211_X1 U14722 ( .C1(n12328), .C2(n12327), .A(n12326), .B(n12325), .ZN(
        P3_U3178) );
  XOR2_X1 U14723 ( .A(n12330), .B(n12329), .Z(n12340) );
  INV_X1 U14724 ( .A(n12331), .ZN(n12560) );
  AOI22_X1 U14725 ( .A1(n12560), .A2(n12332), .B1(P3_REG3_REG_26__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12335) );
  NAND2_X1 U14726 ( .A1(n12545), .A2(n12333), .ZN(n12334) );
  OAI211_X1 U14727 ( .C1(n12521), .C2(n12336), .A(n12335), .B(n12334), .ZN(
        n12337) );
  AOI21_X1 U14728 ( .B1(n12801), .B2(n12338), .A(n12337), .ZN(n12339) );
  OAI21_X1 U14729 ( .B1(n12340), .B2(n15401), .A(n12339), .ZN(P3_U3180) );
  INV_X1 U14730 ( .A(n12521), .ZN(n12542) );
  MUX2_X1 U14731 ( .A(P3_DATAO_REG_27__SCAN_IN), .B(n12542), .S(P3_U3897), .Z(
        P3_U3518) );
  MUX2_X1 U14732 ( .A(n12552), .B(P3_DATAO_REG_26__SCAN_IN), .S(n12350), .Z(
        P3_U3517) );
  MUX2_X1 U14733 ( .A(n12560), .B(P3_DATAO_REG_25__SCAN_IN), .S(n12350), .Z(
        P3_U3516) );
  MUX2_X1 U14734 ( .A(P3_DATAO_REG_24__SCAN_IN), .B(n12551), .S(P3_U3897), .Z(
        P3_U3515) );
  MUX2_X1 U14735 ( .A(P3_DATAO_REG_22__SCAN_IN), .B(n12604), .S(P3_U3897), .Z(
        P3_U3513) );
  MUX2_X1 U14736 ( .A(P3_DATAO_REG_20__SCAN_IN), .B(n12603), .S(P3_U3897), .Z(
        P3_U3511) );
  MUX2_X1 U14737 ( .A(n12341), .B(P3_DATAO_REG_17__SCAN_IN), .S(n12350), .Z(
        P3_U3508) );
  MUX2_X1 U14738 ( .A(n12691), .B(P3_DATAO_REG_16__SCAN_IN), .S(n12350), .Z(
        P3_U3507) );
  MUX2_X1 U14739 ( .A(P3_DATAO_REG_15__SCAN_IN), .B(n12703), .S(P3_U3897), .Z(
        P3_U3506) );
  MUX2_X1 U14740 ( .A(n12719), .B(P3_DATAO_REG_14__SCAN_IN), .S(n12350), .Z(
        P3_U3505) );
  MUX2_X1 U14741 ( .A(P3_DATAO_REG_13__SCAN_IN), .B(n14304), .S(P3_U3897), .Z(
        P3_U3504) );
  MUX2_X1 U14742 ( .A(n15388), .B(P3_DATAO_REG_12__SCAN_IN), .S(n12350), .Z(
        P3_U3503) );
  MUX2_X1 U14743 ( .A(n14984), .B(P3_DATAO_REG_11__SCAN_IN), .S(n12350), .Z(
        P3_U3502) );
  MUX2_X1 U14744 ( .A(P3_DATAO_REG_10__SCAN_IN), .B(n12342), .S(P3_U3897), .Z(
        P3_U3501) );
  MUX2_X1 U14745 ( .A(n14985), .B(P3_DATAO_REG_9__SCAN_IN), .S(n12350), .Z(
        P3_U3500) );
  MUX2_X1 U14746 ( .A(n12343), .B(P3_DATAO_REG_8__SCAN_IN), .S(n12350), .Z(
        P3_U3499) );
  MUX2_X1 U14747 ( .A(P3_DATAO_REG_7__SCAN_IN), .B(n12344), .S(P3_U3897), .Z(
        P3_U3498) );
  MUX2_X1 U14748 ( .A(P3_DATAO_REG_6__SCAN_IN), .B(n12345), .S(P3_U3897), .Z(
        P3_U3497) );
  MUX2_X1 U14749 ( .A(P3_DATAO_REG_5__SCAN_IN), .B(n12346), .S(P3_U3897), .Z(
        P3_U3496) );
  MUX2_X1 U14750 ( .A(P3_DATAO_REG_4__SCAN_IN), .B(n12347), .S(P3_U3897), .Z(
        P3_U3495) );
  MUX2_X1 U14751 ( .A(P3_DATAO_REG_3__SCAN_IN), .B(n12348), .S(P3_U3897), .Z(
        P3_U3494) );
  MUX2_X1 U14752 ( .A(P3_DATAO_REG_1__SCAN_IN), .B(n12349), .S(P3_U3897), .Z(
        P3_U3492) );
  MUX2_X1 U14753 ( .A(n15040), .B(P3_DATAO_REG_0__SCAN_IN), .S(n12350), .Z(
        P3_U3491) );
  INV_X1 U14754 ( .A(n12351), .ZN(n12356) );
  OAI21_X1 U14755 ( .B1(n12354), .B2(n12353), .A(n12352), .ZN(n12355) );
  NAND3_X1 U14756 ( .A1(n12356), .A2(n14961), .A3(n12355), .ZN(n12371) );
  INV_X1 U14757 ( .A(P3_ADDR_REG_12__SCAN_IN), .ZN(n12357) );
  NOR2_X1 U14758 ( .A1(n14834), .A2(n12357), .ZN(n12358) );
  AOI211_X1 U14759 ( .C1(n14843), .C2(n12360), .A(n12359), .B(n12358), .ZN(
        n12370) );
  OAI21_X1 U14760 ( .B1(n6576), .B2(n6724), .A(n12362), .ZN(n12363) );
  NAND2_X1 U14761 ( .A1(n12363), .A2(n12477), .ZN(n12369) );
  OAI21_X1 U14762 ( .B1(n12366), .B2(n12365), .A(n12364), .ZN(n12367) );
  NAND2_X1 U14763 ( .A1(n12367), .A2(n14973), .ZN(n12368) );
  NAND4_X1 U14764 ( .A1(n12371), .A2(n12370), .A3(n12369), .A4(n12368), .ZN(
        P3_U3194) );
  XNOR2_X1 U14765 ( .A(n12400), .B(P3_REG2_REG_14__SCAN_IN), .ZN(n12384) );
  AOI21_X1 U14766 ( .B1(n6684), .B2(n12384), .A(n12396), .ZN(n12395) );
  NAND2_X1 U14767 ( .A1(n12376), .A2(n12375), .ZN(n12378) );
  XNOR2_X1 U14768 ( .A(n12400), .B(n12777), .ZN(n12385) );
  OAI21_X1 U14769 ( .B1(n12379), .B2(n12385), .A(n12398), .ZN(n12393) );
  INV_X1 U14770 ( .A(n12380), .ZN(n12382) );
  AOI21_X1 U14771 ( .B1(n12383), .B2(n12382), .A(n12381), .ZN(n12388) );
  INV_X1 U14772 ( .A(n12384), .ZN(n12386) );
  MUX2_X1 U14773 ( .A(n12386), .B(n12385), .S(n12463), .Z(n12387) );
  NAND2_X1 U14774 ( .A1(n12388), .A2(n12387), .ZN(n12404) );
  OAI211_X1 U14775 ( .C1(n12388), .C2(n12387), .A(n12404), .B(n14961), .ZN(
        n12391) );
  AOI21_X1 U14776 ( .B1(n14969), .B2(P3_ADDR_REG_14__SCAN_IN), .A(n12389), 
        .ZN(n12390) );
  OAI211_X1 U14777 ( .C1(n14966), .C2(n12400), .A(n12391), .B(n12390), .ZN(
        n12392) );
  AOI21_X1 U14778 ( .B1(n14973), .B2(n12393), .A(n12392), .ZN(n12394) );
  OAI21_X1 U14779 ( .B1(n12395), .B2(n14977), .A(n12394), .ZN(P3_U3196) );
  INV_X1 U14780 ( .A(n12422), .ZN(n12432) );
  AOI21_X1 U14781 ( .B1(n12693), .B2(n12397), .A(n12417), .ZN(n12415) );
  NAND2_X1 U14782 ( .A1(n12400), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n12401) );
  NAND2_X1 U14783 ( .A1(P3_REG1_REG_15__SCAN_IN), .A2(n12399), .ZN(n12423) );
  OAI21_X1 U14784 ( .B1(P3_REG1_REG_15__SCAN_IN), .B2(n12399), .A(n12423), 
        .ZN(n12413) );
  NAND2_X1 U14785 ( .A1(n12400), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n12402) );
  MUX2_X1 U14786 ( .A(n12402), .B(n12401), .S(n12463), .Z(n12403) );
  NAND2_X1 U14787 ( .A1(n12404), .A2(n12403), .ZN(n12430) );
  XNOR2_X1 U14788 ( .A(n12430), .B(n12422), .ZN(n12406) );
  MUX2_X1 U14789 ( .A(P3_REG2_REG_15__SCAN_IN), .B(P3_REG1_REG_15__SCAN_IN), 
        .S(n12463), .Z(n12405) );
  NOR2_X1 U14790 ( .A1(n12406), .A2(n12405), .ZN(n12431) );
  AOI21_X1 U14791 ( .B1(n12406), .B2(n12405), .A(n12431), .ZN(n12411) );
  OAI21_X1 U14792 ( .B1(n14834), .B2(n12408), .A(n12407), .ZN(n12409) );
  AOI21_X1 U14793 ( .B1(n14843), .B2(n12432), .A(n12409), .ZN(n12410) );
  OAI21_X1 U14794 ( .B1(n12411), .B2(n14838), .A(n12410), .ZN(n12412) );
  AOI21_X1 U14795 ( .B1(n14973), .B2(n12413), .A(n12412), .ZN(n12414) );
  OAI21_X1 U14796 ( .B1(n12415), .B2(n14977), .A(n12414), .ZN(P3_U3197) );
  INV_X1 U14797 ( .A(n12453), .ZN(n12420) );
  AOI22_X1 U14798 ( .A1(P3_REG2_REG_16__SCAN_IN), .A2(n12453), .B1(n12420), 
        .B2(n12683), .ZN(n12419) );
  AOI21_X1 U14799 ( .B1(n6625), .B2(n12419), .A(n12454), .ZN(n12442) );
  AOI22_X1 U14800 ( .A1(P3_REG1_REG_16__SCAN_IN), .A2(n12420), .B1(n12453), 
        .B2(n12770), .ZN(n12426) );
  NAND2_X1 U14801 ( .A1(n12422), .A2(n12421), .ZN(n12424) );
  OAI21_X1 U14802 ( .B1(n12426), .B2(n12425), .A(n12443), .ZN(n12440) );
  NAND2_X1 U14803 ( .A1(n14843), .A2(n12453), .ZN(n12428) );
  OAI211_X1 U14804 ( .C1(n12429), .C2(n14834), .A(n12428), .B(n12427), .ZN(
        n12439) );
  INV_X1 U14805 ( .A(n12430), .ZN(n12433) );
  AOI21_X1 U14806 ( .B1(n12433), .B2(n12432), .A(n12431), .ZN(n12448) );
  MUX2_X1 U14807 ( .A(n12683), .B(n12770), .S(n12463), .Z(n12434) );
  NOR2_X1 U14808 ( .A1(n12434), .A2(n12453), .ZN(n12447) );
  NAND2_X1 U14809 ( .A1(n12434), .A2(n12453), .ZN(n12446) );
  INV_X1 U14810 ( .A(n12446), .ZN(n12435) );
  NOR2_X1 U14811 ( .A1(n12447), .A2(n12435), .ZN(n12436) );
  XNOR2_X1 U14812 ( .A(n12448), .B(n12436), .ZN(n12437) );
  NOR2_X1 U14813 ( .A1(n12437), .A2(n14838), .ZN(n12438) );
  AOI211_X1 U14814 ( .C1(n14973), .C2(n12440), .A(n12439), .B(n12438), .ZN(
        n12441) );
  OAI21_X1 U14815 ( .B1(n12442), .B2(n14977), .A(n12441), .ZN(P3_U3198) );
  XOR2_X1 U14816 ( .A(P3_REG1_REG_17__SCAN_IN), .B(n12461), .Z(n12459) );
  OAI21_X1 U14817 ( .B1(n14834), .B2(n12445), .A(n12444), .ZN(n12452) );
  MUX2_X1 U14818 ( .A(P3_REG2_REG_17__SCAN_IN), .B(P3_REG1_REG_17__SCAN_IN), 
        .S(n12463), .Z(n12466) );
  XNOR2_X1 U14819 ( .A(n12466), .B(n12465), .ZN(n12450) );
  OAI21_X1 U14820 ( .B1(n12448), .B2(n12447), .A(n12446), .ZN(n12449) );
  NOR2_X1 U14821 ( .A1(n12449), .A2(n12450), .ZN(n12464) );
  AOI211_X1 U14822 ( .C1(n12450), .C2(n12449), .A(n14838), .B(n12464), .ZN(
        n12451) );
  AOI211_X1 U14823 ( .C1(n14843), .C2(n6892), .A(n12452), .B(n12451), .ZN(
        n12458) );
  NAND2_X1 U14824 ( .A1(n12455), .A2(n12465), .ZN(n12475) );
  OAI21_X1 U14825 ( .B1(n6568), .B2(P3_REG2_REG_17__SCAN_IN), .A(n12476), .ZN(
        n12456) );
  NAND2_X1 U14826 ( .A1(n12456), .A2(n12477), .ZN(n12457) );
  OAI211_X1 U14827 ( .C1(n12459), .C2(n12498), .A(n12458), .B(n12457), .ZN(
        P3_U3199) );
  XOR2_X1 U14828 ( .A(P3_REG1_REG_18__SCAN_IN), .B(n12494), .Z(n12495) );
  AOI22_X1 U14829 ( .A1(n12461), .A2(P3_REG1_REG_17__SCAN_IN), .B1(n12465), 
        .B2(n12460), .ZN(n12496) );
  XOR2_X1 U14830 ( .A(n12495), .B(n12496), .Z(n12481) );
  OAI21_X1 U14831 ( .B1(n14834), .B2(n15142), .A(n12462), .ZN(n12471) );
  MUX2_X1 U14832 ( .A(P3_REG2_REG_18__SCAN_IN), .B(P3_REG1_REG_18__SCAN_IN), 
        .S(n12463), .Z(n12468) );
  AOI21_X1 U14833 ( .B1(n12466), .B2(n12465), .A(n12464), .ZN(n12487) );
  XNOR2_X1 U14834 ( .A(n12487), .B(n12494), .ZN(n12467) );
  NOR2_X1 U14835 ( .A1(n12467), .A2(n12468), .ZN(n12486) );
  AOI21_X1 U14836 ( .B1(n12468), .B2(n12467), .A(n12486), .ZN(n12469) );
  NOR2_X1 U14837 ( .A1(n12469), .A2(n14838), .ZN(n12470) );
  AOI211_X1 U14838 ( .C1(n14843), .C2(n12494), .A(n12471), .B(n12470), .ZN(
        n12480) );
  OR2_X1 U14839 ( .A1(n12494), .A2(n12472), .ZN(n12482) );
  NAND2_X1 U14840 ( .A1(n12494), .A2(n12472), .ZN(n12473) );
  NAND2_X1 U14841 ( .A1(n12482), .A2(n12473), .ZN(n12474) );
  OAI21_X1 U14842 ( .B1(n12484), .B2(n12478), .A(n12477), .ZN(n12479) );
  OAI211_X1 U14843 ( .C1(n12481), .C2(n12498), .A(n12480), .B(n12479), .ZN(
        P3_U3200) );
  INV_X1 U14844 ( .A(n12482), .ZN(n12483) );
  XNOR2_X1 U14845 ( .A(n12489), .B(n12631), .ZN(n12491) );
  INV_X1 U14846 ( .A(n12491), .ZN(n12485) );
  AOI21_X1 U14847 ( .B1(n12487), .B2(n12494), .A(n12486), .ZN(n12493) );
  XNOR2_X1 U14848 ( .A(n12489), .B(n12488), .ZN(n12497) );
  MUX2_X1 U14849 ( .A(n12497), .B(n12491), .S(n12490), .Z(n12492) );
  XNOR2_X1 U14850 ( .A(n12493), .B(n12492), .ZN(n12503) );
  AOI21_X1 U14851 ( .B1(n14969), .B2(P3_ADDR_REG_19__SCAN_IN), .A(n12499), 
        .ZN(n12500) );
  OAI21_X1 U14852 ( .B1(n14966), .B2(n12501), .A(n12500), .ZN(n12502) );
  OAI21_X1 U14853 ( .B1(n12505), .B2(n14977), .A(n12504), .ZN(P3_U3201) );
  NAND2_X1 U14854 ( .A1(n12506), .A2(n15055), .ZN(n12509) );
  NAND2_X1 U14855 ( .A1(n12508), .A2(n12507), .ZN(n12727) );
  AOI21_X1 U14856 ( .B1(n12509), .B2(n12727), .A(n15052), .ZN(n12512) );
  AOI21_X1 U14857 ( .B1(P3_REG2_REG_31__SCAN_IN), .B2(n15052), .A(n12512), 
        .ZN(n12510) );
  OAI21_X1 U14858 ( .B1(n12511), .B2(n12709), .A(n12510), .ZN(P3_U3202) );
  AOI21_X1 U14859 ( .B1(n15052), .B2(P3_REG2_REG_30__SCAN_IN), .A(n12512), 
        .ZN(n12513) );
  OAI21_X1 U14860 ( .B1(n12791), .B2(n12709), .A(n12513), .ZN(P3_U3203) );
  XOR2_X1 U14861 ( .A(n12516), .B(n12514), .Z(n12797) );
  INV_X1 U14862 ( .A(P3_REG2_REG_28__SCAN_IN), .ZN(n12524) );
  INV_X1 U14863 ( .A(n12515), .ZN(n12519) );
  AOI21_X1 U14864 ( .B1(n12528), .B2(n12517), .A(n12516), .ZN(n12518) );
  OAI22_X1 U14865 ( .A1(n12521), .A2(n15029), .B1(n12520), .B2(n15031), .ZN(
        n12522) );
  NOR2_X1 U14866 ( .A1(n12523), .A2(n12522), .ZN(n12792) );
  MUX2_X1 U14867 ( .A(n12524), .B(n12792), .S(n15057), .Z(n12527) );
  AOI22_X1 U14868 ( .A1(n12794), .A2(n15014), .B1(n15055), .B2(n12525), .ZN(
        n12526) );
  OAI211_X1 U14869 ( .C1(n12797), .C2(n12725), .A(n12527), .B(n12526), .ZN(
        P3_U3205) );
  AOI21_X1 U14870 ( .B1(n12531), .B2(n12530), .A(n12529), .ZN(n12738) );
  INV_X1 U14871 ( .A(n12738), .ZN(n12537) );
  NAND2_X1 U14872 ( .A1(n12532), .A2(n15049), .ZN(n12736) );
  AOI22_X1 U14873 ( .A1(n12533), .A2(n15055), .B1(n15052), .B2(
        P3_REG2_REG_27__SCAN_IN), .ZN(n12534) );
  OAI21_X1 U14874 ( .B1(n12736), .B2(n12535), .A(n12534), .ZN(n12536) );
  AOI21_X1 U14875 ( .B1(n12537), .B2(n14310), .A(n12536), .ZN(n12538) );
  OAI21_X1 U14876 ( .B1(n12737), .B2(n15052), .A(n12538), .ZN(P3_U3206) );
  XOR2_X1 U14877 ( .A(n12540), .B(n12539), .Z(n12804) );
  INV_X1 U14878 ( .A(P3_REG2_REG_26__SCAN_IN), .ZN(n12544) );
  XNOR2_X1 U14879 ( .A(n12541), .B(n12540), .ZN(n12543) );
  AOI222_X1 U14880 ( .A1(n15046), .A2(n12543), .B1(n12560), .B2(n15041), .C1(
        n12542), .C2(n15038), .ZN(n12799) );
  MUX2_X1 U14881 ( .A(n12544), .B(n12799), .S(n15057), .Z(n12547) );
  AOI22_X1 U14882 ( .A1(n12801), .A2(n15014), .B1(n15055), .B2(n12545), .ZN(
        n12546) );
  OAI211_X1 U14883 ( .C1(n12804), .C2(n12725), .A(n12547), .B(n12546), .ZN(
        P3_U3207) );
  XOR2_X1 U14884 ( .A(n6654), .B(n12549), .Z(n12810) );
  OAI211_X1 U14885 ( .C1(n12550), .C2(n12549), .A(n12548), .B(n15046), .ZN(
        n12554) );
  AOI22_X1 U14886 ( .A1(n12552), .A2(n15038), .B1(n12551), .B2(n15041), .ZN(
        n12553) );
  INV_X1 U14887 ( .A(P3_REG2_REG_25__SCAN_IN), .ZN(n12555) );
  MUX2_X1 U14888 ( .A(n12806), .B(n12555), .S(n15052), .Z(n12558) );
  AOI22_X1 U14889 ( .A1(n12807), .A2(n15014), .B1(n15055), .B2(n12556), .ZN(
        n12557) );
  OAI211_X1 U14890 ( .C1(n12810), .C2(n12725), .A(n12558), .B(n12557), .ZN(
        P3_U3208) );
  OAI211_X1 U14891 ( .C1(n6570), .C2(n12565), .A(n12559), .B(n15046), .ZN(
        n12562) );
  AOI22_X1 U14892 ( .A1(n12560), .A2(n15038), .B1(n15041), .B2(n12592), .ZN(
        n12561) );
  AND2_X1 U14893 ( .A1(n12562), .A2(n12561), .ZN(n12747) );
  AOI21_X1 U14894 ( .B1(n12565), .B2(n12564), .A(n12563), .ZN(n12749) );
  INV_X1 U14895 ( .A(n12749), .ZN(n12570) );
  AOI22_X1 U14896 ( .A1(n12566), .A2(n15055), .B1(n15052), .B2(
        P3_REG2_REG_24__SCAN_IN), .ZN(n12567) );
  OAI21_X1 U14897 ( .B1(n12568), .B2(n12709), .A(n12567), .ZN(n12569) );
  AOI21_X1 U14898 ( .B1(n12570), .B2(n14310), .A(n12569), .ZN(n12571) );
  OAI21_X1 U14899 ( .B1(n15052), .B2(n12747), .A(n12571), .ZN(P3_U3209) );
  XNOR2_X1 U14900 ( .A(n12573), .B(n12572), .ZN(n12814) );
  NAND2_X1 U14901 ( .A1(n12575), .A2(n12574), .ZN(n12576) );
  NAND3_X1 U14902 ( .A1(n6868), .A2(n15046), .A3(n12576), .ZN(n12581) );
  OAI22_X1 U14903 ( .A1(n12578), .A2(n15031), .B1(n12577), .B2(n15029), .ZN(
        n12579) );
  INV_X1 U14904 ( .A(n12579), .ZN(n12580) );
  NAND2_X1 U14905 ( .A1(n12581), .A2(n12580), .ZN(n12812) );
  MUX2_X1 U14906 ( .A(n12812), .B(P3_REG2_REG_23__SCAN_IN), .S(n15052), .Z(
        n12582) );
  INV_X1 U14907 ( .A(n12582), .ZN(n12586) );
  AOI22_X1 U14908 ( .A1(n12584), .A2(n15014), .B1(n15055), .B2(n12583), .ZN(
        n12585) );
  OAI211_X1 U14909 ( .C1(n12814), .C2(n12725), .A(n12586), .B(n12585), .ZN(
        P3_U3210) );
  XNOR2_X1 U14910 ( .A(n12588), .B(n12587), .ZN(n12822) );
  INV_X1 U14911 ( .A(P3_REG2_REG_22__SCAN_IN), .ZN(n12594) );
  XNOR2_X1 U14912 ( .A(n12590), .B(n12589), .ZN(n12593) );
  AOI222_X1 U14913 ( .A1(n15046), .A2(n12593), .B1(n12592), .B2(n15038), .C1(
        n12591), .C2(n15041), .ZN(n12817) );
  MUX2_X1 U14914 ( .A(n12594), .B(n12817), .S(n15057), .Z(n12597) );
  AOI22_X1 U14915 ( .A1(n12819), .A2(n15014), .B1(n15055), .B2(n12595), .ZN(
        n12596) );
  OAI211_X1 U14916 ( .C1(n12822), .C2(n12725), .A(n12597), .B(n12596), .ZN(
        P3_U3211) );
  XNOR2_X1 U14917 ( .A(n12599), .B(n12598), .ZN(n12828) );
  INV_X1 U14918 ( .A(P3_REG2_REG_21__SCAN_IN), .ZN(n12606) );
  OAI21_X1 U14919 ( .B1(n12602), .B2(n12601), .A(n12600), .ZN(n12605) );
  AOI222_X1 U14920 ( .A1(n15046), .A2(n12605), .B1(n12604), .B2(n15038), .C1(
        n12603), .C2(n15041), .ZN(n12823) );
  MUX2_X1 U14921 ( .A(n12606), .B(n12823), .S(n15057), .Z(n12609) );
  AOI22_X1 U14922 ( .A1(n12825), .A2(n15014), .B1(n15055), .B2(n12607), .ZN(
        n12608) );
  OAI211_X1 U14923 ( .C1(n12828), .C2(n12725), .A(n12609), .B(n12608), .ZN(
        P3_U3212) );
  NAND2_X1 U14924 ( .A1(n6692), .A2(n12610), .ZN(n12611) );
  XNOR2_X1 U14925 ( .A(n12611), .B(n12614), .ZN(n12831) );
  OAI211_X1 U14926 ( .C1(n12614), .C2(n12613), .A(n12612), .B(n15046), .ZN(
        n12618) );
  OAI22_X1 U14927 ( .A1(n12615), .A2(n15031), .B1(n12648), .B2(n15029), .ZN(
        n12616) );
  INV_X1 U14928 ( .A(n12616), .ZN(n12617) );
  NAND2_X1 U14929 ( .A1(n12618), .A2(n12617), .ZN(n12829) );
  MUX2_X1 U14930 ( .A(n12829), .B(P3_REG2_REG_20__SCAN_IN), .S(n15052), .Z(
        n12619) );
  INV_X1 U14931 ( .A(n12619), .ZN(n12622) );
  AOI22_X1 U14932 ( .A1(n12758), .A2(n15014), .B1(n15055), .B2(n12620), .ZN(
        n12621) );
  OAI211_X1 U14933 ( .C1(n12831), .C2(n12725), .A(n12622), .B(n12621), .ZN(
        P3_U3213) );
  NAND2_X1 U14934 ( .A1(n12623), .A2(n12633), .ZN(n12624) );
  NAND3_X1 U14935 ( .A1(n12625), .A2(n15046), .A3(n12624), .ZN(n12630) );
  OAI22_X1 U14936 ( .A1(n12627), .A2(n15031), .B1(n12626), .B2(n15029), .ZN(
        n12628) );
  INV_X1 U14937 ( .A(n12628), .ZN(n12629) );
  NAND2_X1 U14938 ( .A1(n12630), .A2(n12629), .ZN(n12834) );
  INV_X1 U14939 ( .A(n12834), .ZN(n12632) );
  MUX2_X1 U14940 ( .A(n12632), .B(n12631), .S(n15052), .Z(n12639) );
  XNOR2_X1 U14941 ( .A(n12634), .B(n12633), .ZN(n12836) );
  INV_X1 U14942 ( .A(n12836), .ZN(n12637) );
  OAI22_X1 U14943 ( .A1(n12835), .A2(n12709), .B1(n12635), .B2(n15020), .ZN(
        n12636) );
  AOI21_X1 U14944 ( .B1(n12637), .B2(n14310), .A(n12636), .ZN(n12638) );
  NAND2_X1 U14945 ( .A1(n12639), .A2(n12638), .ZN(P3_U3214) );
  OR2_X1 U14946 ( .A1(n12677), .A2(n12640), .ZN(n12643) );
  NAND2_X1 U14947 ( .A1(n12643), .A2(n12641), .ZN(n12645) );
  AND2_X1 U14948 ( .A1(n12643), .A2(n12642), .ZN(n12644) );
  AOI21_X1 U14949 ( .B1(n12646), .B2(n12645), .A(n12644), .ZN(n12647) );
  OAI222_X1 U14950 ( .A1(n15031), .A2(n12648), .B1(n15029), .B2(n12679), .C1(
        n15027), .C2(n12647), .ZN(n12763) );
  NAND2_X1 U14951 ( .A1(n12649), .A2(n12650), .ZN(n12651) );
  NAND2_X1 U14952 ( .A1(n12652), .A2(n12651), .ZN(n12841) );
  AOI22_X1 U14953 ( .A1(n15052), .A2(P3_REG2_REG_18__SCAN_IN), .B1(n15055), 
        .B2(n12653), .ZN(n12655) );
  NAND2_X1 U14954 ( .A1(n12764), .A2(n15014), .ZN(n12654) );
  OAI211_X1 U14955 ( .C1(n12841), .C2(n12725), .A(n12655), .B(n12654), .ZN(
        n12656) );
  AOI21_X1 U14956 ( .B1(n12763), .B2(n15057), .A(n12656), .ZN(n12657) );
  INV_X1 U14957 ( .A(n12657), .ZN(P3_U3215) );
  XNOR2_X1 U14958 ( .A(n12658), .B(n12662), .ZN(n12844) );
  INV_X1 U14959 ( .A(n12844), .ZN(n12673) );
  NAND2_X1 U14960 ( .A1(n12681), .A2(n12661), .ZN(n12660) );
  NAND2_X1 U14961 ( .A1(n12660), .A2(n12659), .ZN(n12664) );
  NAND3_X1 U14962 ( .A1(n12681), .A2(n12662), .A3(n12661), .ZN(n12663) );
  NAND3_X1 U14963 ( .A1(n12664), .A2(n15046), .A3(n12663), .ZN(n12667) );
  AOI22_X1 U14964 ( .A1(n12665), .A2(n15038), .B1(n15041), .B2(n12691), .ZN(
        n12666) );
  MUX2_X1 U14965 ( .A(n12843), .B(n12668), .S(n15052), .Z(n12672) );
  INV_X1 U14966 ( .A(n12847), .ZN(n12670) );
  AOI22_X1 U14967 ( .A1(n12670), .A2(n15014), .B1(n15055), .B2(n12669), .ZN(
        n12671) );
  OAI211_X1 U14968 ( .C1(n12673), .C2(n12725), .A(n12672), .B(n12671), .ZN(
        P3_U3216) );
  OAI21_X1 U14969 ( .B1(n12675), .B2(n12676), .A(n12674), .ZN(n12851) );
  INV_X1 U14970 ( .A(n12851), .ZN(n12687) );
  AOI21_X1 U14971 ( .B1(n12677), .B2(n12676), .A(n15027), .ZN(n12682) );
  OAI22_X1 U14972 ( .A1(n12679), .A2(n15031), .B1(n12678), .B2(n15029), .ZN(
        n12680) );
  AOI21_X1 U14973 ( .B1(n12682), .B2(n12681), .A(n12680), .ZN(n12848) );
  MUX2_X1 U14974 ( .A(n12683), .B(n12848), .S(n15057), .Z(n12686) );
  AOI22_X1 U14975 ( .A1(n12850), .A2(n15014), .B1(n15055), .B2(n12684), .ZN(
        n12685) );
  OAI211_X1 U14976 ( .C1(n12687), .C2(n12725), .A(n12686), .B(n12685), .ZN(
        P3_U3217) );
  XOR2_X1 U14977 ( .A(n12688), .B(n12689), .Z(n12860) );
  XNOR2_X1 U14978 ( .A(n12690), .B(n12689), .ZN(n12692) );
  AOI222_X1 U14979 ( .A1(n15046), .A2(n12692), .B1(n12691), .B2(n15038), .C1(
        n12719), .C2(n15041), .ZN(n12854) );
  MUX2_X1 U14980 ( .A(n12693), .B(n12854), .S(n15057), .Z(n12697) );
  INV_X1 U14981 ( .A(n12694), .ZN(n12695) );
  AOI22_X1 U14982 ( .A1(n12856), .A2(n15014), .B1(n15055), .B2(n12695), .ZN(
        n12696) );
  OAI211_X1 U14983 ( .C1(n12860), .C2(n12725), .A(n12697), .B(n12696), .ZN(
        P3_U3218) );
  NAND2_X1 U14984 ( .A1(n14303), .A2(n12698), .ZN(n12700) );
  NAND2_X1 U14985 ( .A1(n12700), .A2(n12699), .ZN(n12702) );
  XNOR2_X1 U14986 ( .A(n12702), .B(n12701), .ZN(n12704) );
  AOI222_X1 U14987 ( .A1(n15046), .A2(n12704), .B1(n12703), .B2(n15038), .C1(
        n14304), .C2(n15041), .ZN(n12861) );
  MUX2_X1 U14988 ( .A(n12705), .B(n12861), .S(n15057), .Z(n12712) );
  XNOR2_X1 U14989 ( .A(n12706), .B(n12707), .ZN(n12863) );
  OAI22_X1 U14990 ( .A1(n12866), .A2(n12709), .B1(n12708), .B2(n15020), .ZN(
        n12710) );
  AOI21_X1 U14991 ( .B1(n12863), .B2(n14310), .A(n12710), .ZN(n12711) );
  NAND2_X1 U14992 ( .A1(n12712), .A2(n12711), .ZN(P3_U3219) );
  XNOR2_X1 U14993 ( .A(n12713), .B(n12717), .ZN(n12873) );
  INV_X1 U14994 ( .A(n12873), .ZN(n12726) );
  NAND2_X1 U14995 ( .A1(n14303), .A2(n12714), .ZN(n12716) );
  NAND2_X1 U14996 ( .A1(n12716), .A2(n12715), .ZN(n12718) );
  XNOR2_X1 U14997 ( .A(n12718), .B(n12717), .ZN(n12720) );
  AOI222_X1 U14998 ( .A1(n15046), .A2(n12720), .B1(n15388), .B2(n15041), .C1(
        n12719), .C2(n15038), .ZN(n12868) );
  MUX2_X1 U14999 ( .A(n11086), .B(n12868), .S(n15057), .Z(n12724) );
  NOR2_X1 U15000 ( .A1(n15020), .A2(n12721), .ZN(n12722) );
  AOI21_X1 U15001 ( .B1(n12871), .B2(n15014), .A(n12722), .ZN(n12723) );
  OAI211_X1 U15002 ( .C1(n12726), .C2(n12725), .A(n12724), .B(n12723), .ZN(
        P3_U3220) );
  INV_X1 U15003 ( .A(P3_REG1_REG_31__SCAN_IN), .ZN(n12729) );
  NAND2_X1 U15004 ( .A1(n12786), .A2(n12782), .ZN(n12728) );
  INV_X1 U15005 ( .A(n12727), .ZN(n12787) );
  NAND2_X1 U15006 ( .A1(n12787), .A2(n15096), .ZN(n12731) );
  OAI211_X1 U15007 ( .C1(n15096), .C2(n12729), .A(n12728), .B(n12731), .ZN(
        P3_U3490) );
  NAND2_X1 U15008 ( .A1(n12730), .A2(n12782), .ZN(n12732) );
  OAI211_X1 U15009 ( .C1(n15096), .C2(n10300), .A(n12732), .B(n12731), .ZN(
        P3_U3489) );
  MUX2_X1 U15010 ( .A(n12733), .B(n12792), .S(n15096), .Z(n12735) );
  NAND2_X1 U15011 ( .A1(n12794), .A2(n12782), .ZN(n12734) );
  OAI211_X1 U15012 ( .C1(n12776), .C2(n12797), .A(n12735), .B(n12734), .ZN(
        P3_U3487) );
  OAI211_X1 U15013 ( .C1(n12748), .C2(n12738), .A(n12737), .B(n12736), .ZN(
        n12798) );
  MUX2_X1 U15014 ( .A(P3_REG1_REG_27__SCAN_IN), .B(n12798), .S(n15096), .Z(
        P3_U3486) );
  MUX2_X1 U15015 ( .A(n12739), .B(n12799), .S(n15096), .Z(n12741) );
  NAND2_X1 U15016 ( .A1(n12801), .A2(n12782), .ZN(n12740) );
  OAI211_X1 U15017 ( .C1(n12804), .C2(n12776), .A(n12741), .B(n12740), .ZN(
        P3_U3485) );
  MUX2_X1 U15018 ( .A(n12806), .B(n12742), .S(n15094), .Z(n12744) );
  NAND2_X1 U15019 ( .A1(n12807), .A2(n12782), .ZN(n12743) );
  OAI211_X1 U15020 ( .C1(n12776), .C2(n12810), .A(n12744), .B(n12743), .ZN(
        P3_U3484) );
  NAND2_X1 U15021 ( .A1(n12745), .A2(n15049), .ZN(n12746) );
  OAI211_X1 U15022 ( .C1(n12749), .C2(n12748), .A(n12747), .B(n12746), .ZN(
        n12811) );
  MUX2_X1 U15023 ( .A(n12811), .B(P3_REG1_REG_24__SCAN_IN), .S(n15094), .Z(
        P3_U3483) );
  MUX2_X1 U15024 ( .A(P3_REG1_REG_23__SCAN_IN), .B(n12812), .S(n15096), .Z(
        n12751) );
  OAI22_X1 U15025 ( .A1(n12814), .A2(n12776), .B1(n12813), .B2(n12780), .ZN(
        n12750) );
  OR2_X1 U15026 ( .A1(n12751), .A2(n12750), .ZN(P3_U3482) );
  INV_X1 U15027 ( .A(P3_REG1_REG_22__SCAN_IN), .ZN(n12752) );
  MUX2_X1 U15028 ( .A(n12752), .B(n12817), .S(n15096), .Z(n12754) );
  NAND2_X1 U15029 ( .A1(n12819), .A2(n12782), .ZN(n12753) );
  OAI211_X1 U15030 ( .C1(n12822), .C2(n12776), .A(n12754), .B(n12753), .ZN(
        P3_U3481) );
  INV_X1 U15031 ( .A(P3_REG1_REG_21__SCAN_IN), .ZN(n12755) );
  MUX2_X1 U15032 ( .A(n12755), .B(n12823), .S(n15096), .Z(n12757) );
  NAND2_X1 U15033 ( .A1(n12825), .A2(n12782), .ZN(n12756) );
  OAI211_X1 U15034 ( .C1(n12828), .C2(n12776), .A(n12757), .B(n12756), .ZN(
        P3_U3480) );
  MUX2_X1 U15035 ( .A(n12829), .B(P3_REG1_REG_20__SCAN_IN), .S(n15094), .Z(
        n12760) );
  INV_X1 U15036 ( .A(n12758), .ZN(n12830) );
  OAI22_X1 U15037 ( .A1(n12831), .A2(n12776), .B1(n12830), .B2(n12780), .ZN(
        n12759) );
  OR2_X1 U15038 ( .A1(n12760), .A2(n12759), .ZN(P3_U3479) );
  MUX2_X1 U15039 ( .A(P3_REG1_REG_19__SCAN_IN), .B(n12834), .S(n15096), .Z(
        n12762) );
  OAI22_X1 U15040 ( .A1(n12836), .A2(n12776), .B1(n12835), .B2(n12780), .ZN(
        n12761) );
  AOI21_X1 U15041 ( .B1(n15049), .B2(n12764), .A(n12763), .ZN(n12839) );
  MUX2_X1 U15042 ( .A(n12765), .B(n12839), .S(n15096), .Z(n12766) );
  OAI21_X1 U15043 ( .B1(n12776), .B2(n12841), .A(n12766), .ZN(P3_U3477) );
  MUX2_X1 U15044 ( .A(n12843), .B(n12767), .S(n15094), .Z(n12769) );
  NAND2_X1 U15045 ( .A1(n12844), .A2(n12783), .ZN(n12768) );
  OAI211_X1 U15046 ( .C1(n12780), .C2(n12847), .A(n12769), .B(n12768), .ZN(
        P3_U3476) );
  MUX2_X1 U15047 ( .A(n12770), .B(n12848), .S(n15096), .Z(n12772) );
  AOI22_X1 U15048 ( .A1(n12851), .A2(n12783), .B1(n12782), .B2(n12850), .ZN(
        n12771) );
  NAND2_X1 U15049 ( .A1(n12772), .A2(n12771), .ZN(P3_U3475) );
  MUX2_X1 U15050 ( .A(n12773), .B(n12854), .S(n15096), .Z(n12775) );
  NAND2_X1 U15051 ( .A1(n12856), .A2(n12782), .ZN(n12774) );
  OAI211_X1 U15052 ( .C1(n12776), .C2(n12860), .A(n12775), .B(n12774), .ZN(
        P3_U3474) );
  MUX2_X1 U15053 ( .A(n12777), .B(n12861), .S(n15096), .Z(n12779) );
  NAND2_X1 U15054 ( .A1(n12863), .A2(n12783), .ZN(n12778) );
  OAI211_X1 U15055 ( .C1(n12780), .C2(n12866), .A(n12779), .B(n12778), .ZN(
        P3_U3473) );
  MUX2_X1 U15056 ( .A(n12781), .B(n12868), .S(n15096), .Z(n12785) );
  AOI22_X1 U15057 ( .A1(n12873), .A2(n12783), .B1(n12871), .B2(n12782), .ZN(
        n12784) );
  NAND2_X1 U15058 ( .A1(n12785), .A2(n12784), .ZN(P3_U3472) );
  NAND2_X1 U15059 ( .A1(n12786), .A2(n12870), .ZN(n12788) );
  NAND2_X1 U15060 ( .A1(n12787), .A2(n15085), .ZN(n12790) );
  OAI211_X1 U15061 ( .C1(n10253), .C2(n15085), .A(n12788), .B(n12790), .ZN(
        P3_U3458) );
  NAND2_X1 U15062 ( .A1(n15086), .A2(P3_REG0_REG_30__SCAN_IN), .ZN(n12789) );
  OAI211_X1 U15063 ( .C1(n12791), .C2(n12867), .A(n12790), .B(n12789), .ZN(
        P3_U3457) );
  INV_X1 U15064 ( .A(P3_REG0_REG_28__SCAN_IN), .ZN(n12793) );
  MUX2_X1 U15065 ( .A(n12793), .B(n12792), .S(n15085), .Z(n12796) );
  NAND2_X1 U15066 ( .A1(n12794), .A2(n12870), .ZN(n12795) );
  OAI211_X1 U15067 ( .C1(n12797), .C2(n12859), .A(n12796), .B(n12795), .ZN(
        P3_U3455) );
  MUX2_X1 U15068 ( .A(P3_REG0_REG_27__SCAN_IN), .B(n12798), .S(n15085), .Z(
        P3_U3454) );
  INV_X1 U15069 ( .A(P3_REG0_REG_26__SCAN_IN), .ZN(n12800) );
  MUX2_X1 U15070 ( .A(n12800), .B(n12799), .S(n15085), .Z(n12803) );
  NAND2_X1 U15071 ( .A1(n12801), .A2(n12870), .ZN(n12802) );
  OAI211_X1 U15072 ( .C1(n12804), .C2(n12859), .A(n12803), .B(n12802), .ZN(
        P3_U3453) );
  INV_X1 U15073 ( .A(P3_REG0_REG_25__SCAN_IN), .ZN(n12805) );
  MUX2_X1 U15074 ( .A(n12806), .B(n12805), .S(n15086), .Z(n12809) );
  NAND2_X1 U15075 ( .A1(n12807), .A2(n12870), .ZN(n12808) );
  OAI211_X1 U15076 ( .C1(n12810), .C2(n12859), .A(n12809), .B(n12808), .ZN(
        P3_U3452) );
  MUX2_X1 U15077 ( .A(n12811), .B(P3_REG0_REG_24__SCAN_IN), .S(n15086), .Z(
        P3_U3451) );
  MUX2_X1 U15078 ( .A(n12812), .B(P3_REG0_REG_23__SCAN_IN), .S(n15086), .Z(
        n12816) );
  OAI22_X1 U15079 ( .A1(n12814), .A2(n12859), .B1(n12813), .B2(n12867), .ZN(
        n12815) );
  OR2_X1 U15080 ( .A1(n12816), .A2(n12815), .ZN(P3_U3450) );
  INV_X1 U15081 ( .A(P3_REG0_REG_22__SCAN_IN), .ZN(n12818) );
  MUX2_X1 U15082 ( .A(n12818), .B(n12817), .S(n15085), .Z(n12821) );
  NAND2_X1 U15083 ( .A1(n12819), .A2(n12870), .ZN(n12820) );
  OAI211_X1 U15084 ( .C1(n12822), .C2(n12859), .A(n12821), .B(n12820), .ZN(
        P3_U3449) );
  INV_X1 U15085 ( .A(P3_REG0_REG_21__SCAN_IN), .ZN(n12824) );
  MUX2_X1 U15086 ( .A(n12824), .B(n12823), .S(n15085), .Z(n12827) );
  NAND2_X1 U15087 ( .A1(n12825), .A2(n12870), .ZN(n12826) );
  OAI211_X1 U15088 ( .C1(n12828), .C2(n12859), .A(n12827), .B(n12826), .ZN(
        P3_U3448) );
  MUX2_X1 U15089 ( .A(n12829), .B(P3_REG0_REG_20__SCAN_IN), .S(n15086), .Z(
        n12833) );
  OAI22_X1 U15090 ( .A1(n12831), .A2(n12859), .B1(n12830), .B2(n12867), .ZN(
        n12832) );
  OR2_X1 U15091 ( .A1(n12833), .A2(n12832), .ZN(P3_U3447) );
  MUX2_X1 U15092 ( .A(n12834), .B(P3_REG0_REG_19__SCAN_IN), .S(n15086), .Z(
        n12838) );
  OAI22_X1 U15093 ( .A1(n12836), .A2(n12859), .B1(n12835), .B2(n12867), .ZN(
        n12837) );
  MUX2_X1 U15094 ( .A(n15154), .B(n12839), .S(n15085), .Z(n12840) );
  OAI21_X1 U15095 ( .B1(n12841), .B2(n12859), .A(n12840), .ZN(P3_U3444) );
  MUX2_X1 U15096 ( .A(n12843), .B(n12842), .S(n15086), .Z(n12846) );
  NAND2_X1 U15097 ( .A1(n12844), .A2(n12872), .ZN(n12845) );
  OAI211_X1 U15098 ( .C1(n12867), .C2(n12847), .A(n12846), .B(n12845), .ZN(
        P3_U3441) );
  MUX2_X1 U15099 ( .A(n12849), .B(n12848), .S(n15085), .Z(n12853) );
  AOI22_X1 U15100 ( .A1(n12851), .A2(n12872), .B1(n12870), .B2(n12850), .ZN(
        n12852) );
  NAND2_X1 U15101 ( .A1(n12853), .A2(n12852), .ZN(P3_U3438) );
  INV_X1 U15102 ( .A(P3_REG0_REG_15__SCAN_IN), .ZN(n12855) );
  MUX2_X1 U15103 ( .A(n12855), .B(n12854), .S(n15085), .Z(n12858) );
  NAND2_X1 U15104 ( .A1(n12856), .A2(n12870), .ZN(n12857) );
  OAI211_X1 U15105 ( .C1(n12860), .C2(n12859), .A(n12858), .B(n12857), .ZN(
        P3_U3435) );
  MUX2_X1 U15106 ( .A(n12862), .B(n12861), .S(n15085), .Z(n12865) );
  NAND2_X1 U15107 ( .A1(n12863), .A2(n12872), .ZN(n12864) );
  OAI211_X1 U15108 ( .C1(n12867), .C2(n12866), .A(n12865), .B(n12864), .ZN(
        P3_U3432) );
  INV_X1 U15109 ( .A(P3_REG0_REG_13__SCAN_IN), .ZN(n12869) );
  MUX2_X1 U15110 ( .A(n12869), .B(n12868), .S(n15085), .Z(n12875) );
  AOI22_X1 U15111 ( .A1(n12873), .A2(n12872), .B1(n12871), .B2(n12870), .ZN(
        n12874) );
  NAND2_X1 U15112 ( .A1(n12875), .A2(n12874), .ZN(P3_U3429) );
  NAND4_X1 U15113 ( .A1(n12877), .A2(P3_IR_REG_31__SCAN_IN), .A3(
        P3_STATE_REG_SCAN_IN), .A4(n9378), .ZN(n12879) );
  OAI22_X1 U15114 ( .A1(n12876), .A2(n12879), .B1(n12878), .B2(n11338), .ZN(
        n12880) );
  AOI21_X1 U15115 ( .B1(n12882), .B2(n12881), .A(n12880), .ZN(n12883) );
  INV_X1 U15116 ( .A(n12883), .ZN(P3_U3264) );
  INV_X1 U15117 ( .A(n12884), .ZN(n12885) );
  XNOR2_X1 U15118 ( .A(n13412), .B(n6528), .ZN(n12888) );
  NAND2_X1 U15119 ( .A1(n13035), .A2(n12940), .ZN(n12887) );
  XNOR2_X1 U15120 ( .A(n12888), .B(n12887), .ZN(n13004) );
  INV_X1 U15121 ( .A(n12887), .ZN(n12889) );
  AND2_X1 U15122 ( .A1(n13034), .A2(n13326), .ZN(n12891) );
  XNOR2_X1 U15123 ( .A(n13402), .B(n6528), .ZN(n12893) );
  AND2_X1 U15124 ( .A1(n13033), .A2(n13326), .ZN(n12892) );
  NOR2_X1 U15125 ( .A1(n12893), .A2(n12892), .ZN(n12983) );
  NAND2_X1 U15126 ( .A1(n12893), .A2(n12892), .ZN(n12984) );
  XNOR2_X1 U15127 ( .A(n13459), .B(n6528), .ZN(n12894) );
  NAND2_X1 U15128 ( .A1(n13032), .A2(n12940), .ZN(n12895) );
  XNOR2_X1 U15129 ( .A(n12894), .B(n12895), .ZN(n12955) );
  INV_X1 U15130 ( .A(n12895), .ZN(n12896) );
  XNOR2_X1 U15131 ( .A(n13263), .B(n6528), .ZN(n12898) );
  XNOR2_X1 U15132 ( .A(n12899), .B(n12898), .ZN(n12995) );
  NAND2_X1 U15133 ( .A1(n13031), .A2(n13326), .ZN(n12994) );
  AND2_X1 U15134 ( .A1(n12899), .A2(n12898), .ZN(n12900) );
  XNOR2_X1 U15135 ( .A(n13385), .B(n6528), .ZN(n12901) );
  NAND2_X1 U15136 ( .A1(n13030), .A2(n13326), .ZN(n12925) );
  INV_X1 U15137 ( .A(n12901), .ZN(n12903) );
  XNOR2_X1 U15138 ( .A(n13233), .B(n6541), .ZN(n12905) );
  NAND2_X1 U15139 ( .A1(n13029), .A2(n12940), .ZN(n12904) );
  NOR2_X1 U15140 ( .A1(n12905), .A2(n12904), .ZN(n12906) );
  AOI21_X1 U15141 ( .B1(n12905), .B2(n12904), .A(n12906), .ZN(n12975) );
  INV_X1 U15142 ( .A(n12906), .ZN(n12907) );
  XNOR2_X1 U15143 ( .A(n13375), .B(n6540), .ZN(n12909) );
  NAND2_X1 U15144 ( .A1(n13028), .A2(n13326), .ZN(n12908) );
  NOR2_X1 U15145 ( .A1(n12909), .A2(n12908), .ZN(n12910) );
  AOI21_X1 U15146 ( .B1(n12909), .B2(n12908), .A(n12910), .ZN(n12965) );
  INV_X1 U15147 ( .A(n12910), .ZN(n12911) );
  NAND2_X1 U15148 ( .A1(n13027), .A2(n13326), .ZN(n12912) );
  XNOR2_X1 U15149 ( .A(n13205), .B(n6528), .ZN(n12914) );
  XOR2_X1 U15150 ( .A(n12912), .B(n12914), .Z(n13013) );
  INV_X1 U15151 ( .A(n12912), .ZN(n12913) );
  XNOR2_X1 U15152 ( .A(n13187), .B(n6540), .ZN(n12917) );
  NAND2_X1 U15153 ( .A1(n13026), .A2(n9445), .ZN(n12916) );
  NOR2_X1 U15154 ( .A1(n12917), .A2(n12916), .ZN(n12937) );
  AOI21_X1 U15155 ( .B1(n12917), .B2(n12916), .A(n12937), .ZN(n12918) );
  OAI211_X1 U15156 ( .C1(n12919), .C2(n12918), .A(n12939), .B(n12973), .ZN(
        n12923) );
  INV_X1 U15157 ( .A(n12920), .ZN(n13188) );
  AOI22_X1 U15158 ( .A1(n14336), .A2(n13025), .B1(n13027), .B2(n14334), .ZN(
        n13184) );
  OAI22_X1 U15159 ( .A1(n14343), .A2(n13184), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n15265), .ZN(n12921) );
  AOI21_X1 U15160 ( .B1(n13188), .B2(n13000), .A(n12921), .ZN(n12922) );
  OAI211_X1 U15161 ( .C1(n13442), .C2(n14340), .A(n12923), .B(n12922), .ZN(
        P2_U3186) );
  XOR2_X1 U15162 ( .A(n12925), .B(n12924), .Z(n12930) );
  AOI22_X1 U15163 ( .A1(n13031), .A2(n14334), .B1(n14336), .B2(n13029), .ZN(
        n13241) );
  INV_X1 U15164 ( .A(n12926), .ZN(n13244) );
  AOI22_X1 U15165 ( .A1(n13000), .A2(n13244), .B1(P2_REG3_REG_23__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12927) );
  OAI21_X1 U15166 ( .B1(n13241), .B2(n14343), .A(n12927), .ZN(n12928) );
  AOI21_X1 U15167 ( .B1(n13385), .B2(n13019), .A(n12928), .ZN(n12929) );
  OAI21_X1 U15168 ( .B1(n12930), .B2(n14342), .A(n12929), .ZN(P2_U3188) );
  OAI21_X1 U15169 ( .B1(n6693), .B2(n6564), .A(n12931), .ZN(n12932) );
  NAND2_X1 U15170 ( .A1(n12932), .A2(n12973), .ZN(n12936) );
  INV_X1 U15171 ( .A(n13313), .ZN(n12934) );
  AOI22_X1 U15172 ( .A1(n13033), .A2(n14336), .B1(n14334), .B2(n13035), .ZN(
        n13304) );
  NAND2_X1 U15173 ( .A1(P2_U3088), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n13148)
         );
  OAI21_X1 U15174 ( .B1(n13304), .B2(n14343), .A(n13148), .ZN(n12933) );
  AOI21_X1 U15175 ( .B1(n12934), .B2(n13000), .A(n12933), .ZN(n12935) );
  OAI211_X1 U15176 ( .C1(n8168), .C2(n14340), .A(n12936), .B(n12935), .ZN(
        P2_U3191) );
  INV_X1 U15177 ( .A(n12937), .ZN(n12938) );
  NAND2_X1 U15178 ( .A1(n12939), .A2(n12938), .ZN(n12945) );
  NAND2_X1 U15179 ( .A1(n13025), .A2(n9445), .ZN(n12941) );
  XNOR2_X1 U15180 ( .A(n6528), .B(n12941), .ZN(n12943) );
  XNOR2_X1 U15181 ( .A(n13356), .B(n12943), .ZN(n12944) );
  XNOR2_X1 U15182 ( .A(n12945), .B(n12944), .ZN(n12953) );
  OAI22_X1 U15183 ( .A1(n12949), .A2(n12948), .B1(n12947), .B2(n12946), .ZN(
        n13172) );
  AOI22_X1 U15184 ( .A1(n13016), .A2(n13172), .B1(P2_REG3_REG_28__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12950) );
  OAI21_X1 U15185 ( .B1(n13166), .B2(n14348), .A(n12950), .ZN(n12951) );
  AOI21_X1 U15186 ( .B1(n13356), .B2(n13019), .A(n12951), .ZN(n12952) );
  OAI21_X1 U15187 ( .B1(n12953), .B2(n14342), .A(n12952), .ZN(P2_U3192) );
  OAI211_X1 U15188 ( .C1(n12956), .C2(n12955), .A(n12954), .B(n12973), .ZN(
        n12963) );
  NAND2_X1 U15189 ( .A1(n13031), .A2(n14336), .ZN(n12958) );
  NAND2_X1 U15190 ( .A1(n13033), .A2(n14334), .ZN(n12957) );
  NAND2_X1 U15191 ( .A1(n12958), .A2(n12957), .ZN(n13273) );
  INV_X1 U15192 ( .A(n13277), .ZN(n12960) );
  INV_X1 U15193 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n12959) );
  OAI22_X1 U15194 ( .A1(n12960), .A2(n14348), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n12959), .ZN(n12961) );
  AOI21_X1 U15195 ( .B1(n13273), .B2(n13016), .A(n12961), .ZN(n12962) );
  OAI211_X1 U15196 ( .C1(n6797), .C2(n14340), .A(n12963), .B(n12962), .ZN(
        P2_U3195) );
  OAI211_X1 U15197 ( .C1(n12966), .C2(n12965), .A(n12964), .B(n12973), .ZN(
        n12972) );
  INV_X1 U15198 ( .A(n12967), .ZN(n13217) );
  NAND2_X1 U15199 ( .A1(n13029), .A2(n14334), .ZN(n12969) );
  NAND2_X1 U15200 ( .A1(n13027), .A2(n14336), .ZN(n12968) );
  AND2_X1 U15201 ( .A1(n12969), .A2(n12968), .ZN(n13213) );
  OAI22_X1 U15202 ( .A1(n14343), .A2(n13213), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n15148), .ZN(n12970) );
  AOI21_X1 U15203 ( .B1(n13217), .B2(n13000), .A(n12970), .ZN(n12971) );
  OAI211_X1 U15204 ( .C1(n13220), .C2(n14340), .A(n12972), .B(n12971), .ZN(
        P2_U3197) );
  OAI211_X1 U15205 ( .C1(n12976), .C2(n12975), .A(n12974), .B(n12973), .ZN(
        n12982) );
  NAND2_X1 U15206 ( .A1(n13030), .A2(n14334), .ZN(n12978) );
  NAND2_X1 U15207 ( .A1(n13028), .A2(n14336), .ZN(n12977) );
  NAND2_X1 U15208 ( .A1(n12978), .A2(n12977), .ZN(n13226) );
  AOI22_X1 U15209 ( .A1(n13016), .A2(n13226), .B1(P2_REG3_REG_24__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12979) );
  OAI21_X1 U15210 ( .B1(n13231), .B2(n14348), .A(n12979), .ZN(n12980) );
  AOI21_X1 U15211 ( .B1(n13233), .B2(n13019), .A(n12980), .ZN(n12981) );
  NAND2_X1 U15212 ( .A1(n12982), .A2(n12981), .ZN(P2_U3201) );
  INV_X1 U15213 ( .A(n12983), .ZN(n12985) );
  NAND2_X1 U15214 ( .A1(n12985), .A2(n12984), .ZN(n12986) );
  XNOR2_X1 U15215 ( .A(n12987), .B(n12986), .ZN(n12992) );
  AOI22_X1 U15216 ( .A1(n13032), .A2(n14336), .B1(n14334), .B2(n13034), .ZN(
        n13290) );
  INV_X1 U15217 ( .A(n13290), .ZN(n12988) );
  AOI22_X1 U15218 ( .A1(n12988), .A2(n13016), .B1(P2_REG3_REG_20__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12989) );
  OAI21_X1 U15219 ( .B1(n13295), .B2(n14348), .A(n12989), .ZN(n12990) );
  AOI21_X1 U15220 ( .B1(n13402), .B2(n13019), .A(n12990), .ZN(n12991) );
  OAI21_X1 U15221 ( .B1(n12992), .B2(n14342), .A(n12991), .ZN(P2_U3205) );
  AOI211_X1 U15222 ( .C1(n12995), .C2(n12994), .A(n14342), .B(n12993), .ZN(
        n12996) );
  INV_X1 U15223 ( .A(n12996), .ZN(n13003) );
  INV_X1 U15224 ( .A(n13261), .ZN(n13001) );
  AND2_X1 U15225 ( .A1(n13030), .A2(n14336), .ZN(n12997) );
  AOI21_X1 U15226 ( .B1(n13032), .B2(n14334), .A(n12997), .ZN(n13257) );
  OAI22_X1 U15227 ( .A1(n13257), .A2(n14343), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n12998), .ZN(n12999) );
  AOI21_X1 U15228 ( .B1(n13001), .B2(n13000), .A(n12999), .ZN(n13002) );
  OAI211_X1 U15229 ( .C1(n13456), .C2(n14340), .A(n13003), .B(n13002), .ZN(
        P2_U3207) );
  XNOR2_X1 U15230 ( .A(n13005), .B(n13004), .ZN(n13011) );
  NOR2_X1 U15231 ( .A1(n14348), .A2(n13324), .ZN(n13009) );
  AND2_X1 U15232 ( .A1(n13036), .A2(n14334), .ZN(n13006) );
  AOI21_X1 U15233 ( .B1(n13034), .B2(n14336), .A(n13006), .ZN(n13337) );
  OAI21_X1 U15234 ( .B1(n13337), .B2(n14343), .A(n13007), .ZN(n13008) );
  AOI211_X1 U15235 ( .C1(n13412), .C2(n13019), .A(n13009), .B(n13008), .ZN(
        n13010) );
  OAI21_X1 U15236 ( .B1(n13011), .B2(n14342), .A(n13010), .ZN(P2_U3210) );
  AOI21_X1 U15237 ( .B1(n13013), .B2(n13012), .A(n6621), .ZN(n13021) );
  NAND2_X1 U15238 ( .A1(n13028), .A2(n14334), .ZN(n13015) );
  NAND2_X1 U15239 ( .A1(n13026), .A2(n14336), .ZN(n13014) );
  NAND2_X1 U15240 ( .A1(n13015), .A2(n13014), .ZN(n13198) );
  AOI22_X1 U15241 ( .A1(n13016), .A2(n13198), .B1(P2_REG3_REG_26__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13017) );
  OAI21_X1 U15242 ( .B1(n13203), .B2(n14348), .A(n13017), .ZN(n13018) );
  AOI21_X1 U15243 ( .B1(n13205), .B2(n13019), .A(n13018), .ZN(n13020) );
  OAI21_X1 U15244 ( .B1(n13021), .B2(n14342), .A(n13020), .ZN(P2_U3212) );
  INV_X2 U15245 ( .A(P2_U3947), .ZN(n13043) );
  MUX2_X1 U15246 ( .A(n13022), .B(P2_DATAO_REG_31__SCAN_IN), .S(n13043), .Z(
        P2_U3562) );
  MUX2_X1 U15247 ( .A(n13023), .B(P2_DATAO_REG_30__SCAN_IN), .S(n13043), .Z(
        P2_U3561) );
  MUX2_X1 U15248 ( .A(n13024), .B(P2_DATAO_REG_29__SCAN_IN), .S(n13043), .Z(
        P2_U3560) );
  MUX2_X1 U15249 ( .A(n13025), .B(P2_DATAO_REG_28__SCAN_IN), .S(n13043), .Z(
        P2_U3559) );
  MUX2_X1 U15250 ( .A(n13026), .B(P2_DATAO_REG_27__SCAN_IN), .S(n13043), .Z(
        P2_U3558) );
  MUX2_X1 U15251 ( .A(n13027), .B(P2_DATAO_REG_26__SCAN_IN), .S(n13043), .Z(
        P2_U3557) );
  MUX2_X1 U15252 ( .A(n13028), .B(P2_DATAO_REG_25__SCAN_IN), .S(n13043), .Z(
        P2_U3556) );
  MUX2_X1 U15253 ( .A(n13029), .B(P2_DATAO_REG_24__SCAN_IN), .S(n13043), .Z(
        P2_U3555) );
  MUX2_X1 U15254 ( .A(n13030), .B(P2_DATAO_REG_23__SCAN_IN), .S(n13043), .Z(
        P2_U3554) );
  MUX2_X1 U15255 ( .A(n13031), .B(P2_DATAO_REG_22__SCAN_IN), .S(n13043), .Z(
        P2_U3553) );
  MUX2_X1 U15256 ( .A(n13032), .B(P2_DATAO_REG_21__SCAN_IN), .S(n13043), .Z(
        P2_U3552) );
  MUX2_X1 U15257 ( .A(n13033), .B(P2_DATAO_REG_20__SCAN_IN), .S(n13043), .Z(
        P2_U3551) );
  MUX2_X1 U15258 ( .A(n13034), .B(P2_DATAO_REG_19__SCAN_IN), .S(n13043), .Z(
        P2_U3550) );
  MUX2_X1 U15259 ( .A(n13035), .B(P2_DATAO_REG_18__SCAN_IN), .S(n13043), .Z(
        P2_U3549) );
  MUX2_X1 U15260 ( .A(n13036), .B(P2_DATAO_REG_17__SCAN_IN), .S(n13043), .Z(
        P2_U3548) );
  MUX2_X1 U15261 ( .A(n13037), .B(P2_DATAO_REG_16__SCAN_IN), .S(n13043), .Z(
        P2_U3547) );
  MUX2_X1 U15262 ( .A(n14337), .B(P2_DATAO_REG_15__SCAN_IN), .S(n13043), .Z(
        P2_U3546) );
  MUX2_X1 U15263 ( .A(n13038), .B(P2_DATAO_REG_14__SCAN_IN), .S(n13043), .Z(
        P2_U3545) );
  MUX2_X1 U15264 ( .A(n14335), .B(P2_DATAO_REG_13__SCAN_IN), .S(n13043), .Z(
        P2_U3544) );
  MUX2_X1 U15265 ( .A(n13039), .B(P2_DATAO_REG_12__SCAN_IN), .S(n13043), .Z(
        P2_U3543) );
  MUX2_X1 U15266 ( .A(n13040), .B(P2_DATAO_REG_11__SCAN_IN), .S(n13043), .Z(
        P2_U3542) );
  MUX2_X1 U15267 ( .A(n13041), .B(P2_DATAO_REG_10__SCAN_IN), .S(n13043), .Z(
        P2_U3541) );
  MUX2_X1 U15268 ( .A(n13042), .B(P2_DATAO_REG_9__SCAN_IN), .S(n13043), .Z(
        P2_U3540) );
  MUX2_X1 U15269 ( .A(n13044), .B(P2_DATAO_REG_8__SCAN_IN), .S(n13043), .Z(
        P2_U3539) );
  MUX2_X1 U15270 ( .A(n13045), .B(P2_DATAO_REG_7__SCAN_IN), .S(n13043), .Z(
        P2_U3538) );
  MUX2_X1 U15271 ( .A(n13046), .B(P2_DATAO_REG_6__SCAN_IN), .S(n13043), .Z(
        P2_U3537) );
  MUX2_X1 U15272 ( .A(n13047), .B(P2_DATAO_REG_5__SCAN_IN), .S(n13043), .Z(
        P2_U3536) );
  MUX2_X1 U15273 ( .A(n13048), .B(P2_DATAO_REG_4__SCAN_IN), .S(n13043), .Z(
        P2_U3535) );
  MUX2_X1 U15274 ( .A(n13049), .B(P2_DATAO_REG_3__SCAN_IN), .S(n13043), .Z(
        P2_U3534) );
  MUX2_X1 U15275 ( .A(n13050), .B(P2_DATAO_REG_2__SCAN_IN), .S(n13043), .Z(
        P2_U3533) );
  MUX2_X1 U15276 ( .A(n13051), .B(P2_DATAO_REG_1__SCAN_IN), .S(n13043), .Z(
        P2_U3532) );
  MUX2_X1 U15277 ( .A(n11928), .B(P2_DATAO_REG_0__SCAN_IN), .S(n13043), .Z(
        P2_U3531) );
  OAI211_X1 U15278 ( .C1(n13054), .C2(n13053), .A(n14756), .B(n13052), .ZN(
        n13063) );
  OAI211_X1 U15279 ( .C1(n13057), .C2(n13056), .A(n14759), .B(n13055), .ZN(
        n13062) );
  INV_X1 U15280 ( .A(n13058), .ZN(n13059) );
  AOI22_X1 U15281 ( .A1(n14754), .A2(n13059), .B1(P2_REG3_REG_1__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13061) );
  NAND2_X1 U15282 ( .A1(n14752), .A2(P2_ADDR_REG_1__SCAN_IN), .ZN(n13060) );
  NAND4_X1 U15283 ( .A1(n13063), .A2(n13062), .A3(n13061), .A4(n13060), .ZN(
        P2_U3215) );
  OAI211_X1 U15284 ( .C1(n13065), .C2(n13064), .A(n14756), .B(n13078), .ZN(
        n13072) );
  OAI211_X1 U15285 ( .C1(n13067), .C2(n13066), .A(n14759), .B(n13084), .ZN(
        n13071) );
  AOI22_X1 U15286 ( .A1(n14754), .A2(n13068), .B1(P2_U3088), .B2(
        P2_REG3_REG_2__SCAN_IN), .ZN(n13070) );
  NAND2_X1 U15287 ( .A1(n14752), .A2(P2_ADDR_REG_2__SCAN_IN), .ZN(n13069) );
  NAND4_X1 U15288 ( .A1(n13072), .A2(n13071), .A3(n13070), .A4(n13069), .ZN(
        P2_U3216) );
  OAI21_X1 U15289 ( .B1(n14739), .B2(n13074), .A(n13073), .ZN(n13075) );
  AOI21_X1 U15290 ( .B1(n14752), .B2(P2_ADDR_REG_3__SCAN_IN), .A(n13075), .ZN(
        n13088) );
  MUX2_X1 U15291 ( .A(n9301), .B(P2_REG2_REG_3__SCAN_IN), .S(n13081), .Z(
        n13076) );
  NAND3_X1 U15292 ( .A1(n13078), .A2(n13077), .A3(n13076), .ZN(n13079) );
  NAND3_X1 U15293 ( .A1(n14756), .A2(n13080), .A3(n13079), .ZN(n13087) );
  MUX2_X1 U15294 ( .A(n7623), .B(P2_REG1_REG_3__SCAN_IN), .S(n13081), .Z(
        n13082) );
  NAND3_X1 U15295 ( .A1(n13084), .A2(n13083), .A3(n13082), .ZN(n13085) );
  NAND3_X1 U15296 ( .A1(n14759), .A2(n14663), .A3(n13085), .ZN(n13086) );
  NAND3_X1 U15297 ( .A1(n13088), .A2(n13087), .A3(n13086), .ZN(P2_U3217) );
  OAI21_X1 U15298 ( .B1(n14739), .B2(n13090), .A(n13089), .ZN(n13091) );
  AOI21_X1 U15299 ( .B1(n14752), .B2(P2_ADDR_REG_7__SCAN_IN), .A(n13091), .ZN(
        n13103) );
  MUX2_X1 U15300 ( .A(n10182), .B(P2_REG2_REG_7__SCAN_IN), .S(n13096), .Z(
        n13092) );
  NAND3_X1 U15301 ( .A1(n13094), .A2(n13093), .A3(n13092), .ZN(n13095) );
  NAND3_X1 U15302 ( .A1(n14756), .A2(n13108), .A3(n13095), .ZN(n13102) );
  MUX2_X1 U15303 ( .A(n9333), .B(P2_REG1_REG_7__SCAN_IN), .S(n13096), .Z(
        n13097) );
  NAND3_X1 U15304 ( .A1(n13099), .A2(n13098), .A3(n13097), .ZN(n13100) );
  NAND3_X1 U15305 ( .A1(n14759), .A2(n13114), .A3(n13100), .ZN(n13101) );
  NAND3_X1 U15306 ( .A1(n13103), .A2(n13102), .A3(n13101), .ZN(P2_U3221) );
  NOR2_X1 U15307 ( .A1(n14736), .A2(n7040), .ZN(n13104) );
  AOI211_X1 U15308 ( .C1(n14754), .C2(n13111), .A(n13105), .B(n13104), .ZN(
        n13119) );
  MUX2_X1 U15309 ( .A(n10474), .B(P2_REG2_REG_8__SCAN_IN), .S(n13111), .Z(
        n13106) );
  NAND3_X1 U15310 ( .A1(n13108), .A2(n13107), .A3(n13106), .ZN(n13109) );
  NAND3_X1 U15311 ( .A1(n14756), .A2(n13110), .A3(n13109), .ZN(n13118) );
  MUX2_X1 U15312 ( .A(n9336), .B(P2_REG1_REG_8__SCAN_IN), .S(n13111), .Z(
        n13112) );
  NAND3_X1 U15313 ( .A1(n13114), .A2(n13113), .A3(n13112), .ZN(n13115) );
  NAND3_X1 U15314 ( .A1(n14759), .A2(n13116), .A3(n13115), .ZN(n13117) );
  NAND3_X1 U15315 ( .A1(n13119), .A2(n13118), .A3(n13117), .ZN(P2_U3222) );
  OAI211_X1 U15316 ( .C1(n13122), .C2(n13121), .A(n14756), .B(n13120), .ZN(
        n13131) );
  OAI21_X1 U15317 ( .B1(n14739), .B2(n13124), .A(n13123), .ZN(n13125) );
  AOI21_X1 U15318 ( .B1(n14752), .B2(P2_ADDR_REG_17__SCAN_IN), .A(n13125), 
        .ZN(n13130) );
  OAI211_X1 U15319 ( .C1(n13128), .C2(n13127), .A(n14759), .B(n13126), .ZN(
        n13129) );
  NAND3_X1 U15320 ( .A1(n13131), .A2(n13130), .A3(n13129), .ZN(P2_U3231) );
  NOR2_X1 U15321 ( .A1(n13133), .A2(n13132), .ZN(n13134) );
  XNOR2_X1 U15322 ( .A(n13134), .B(P2_REG2_REG_19__SCAN_IN), .ZN(n13143) );
  INV_X1 U15323 ( .A(n13143), .ZN(n13141) );
  NAND2_X1 U15324 ( .A1(n13136), .A2(n13135), .ZN(n13137) );
  NAND2_X1 U15325 ( .A1(n13138), .A2(n13137), .ZN(n13139) );
  XNOR2_X1 U15326 ( .A(n13139), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n13142) );
  NAND2_X1 U15327 ( .A1(n13142), .A2(n14759), .ZN(n13140) );
  OAI211_X1 U15328 ( .C1(n13141), .C2(n14745), .A(n14739), .B(n13140), .ZN(
        n13146) );
  INV_X1 U15329 ( .A(n14759), .ZN(n14711) );
  OAI22_X1 U15330 ( .A1(n13143), .A2(n14745), .B1(n13142), .B2(n14711), .ZN(
        n13145) );
  MUX2_X1 U15331 ( .A(n13146), .B(n13145), .S(n13144), .Z(n13147) );
  INV_X1 U15332 ( .A(n13147), .ZN(n13149) );
  OAI211_X1 U15333 ( .C1(n7477), .C2(n14736), .A(n13149), .B(n13148), .ZN(
        P2_U3233) );
  NAND2_X1 U15334 ( .A1(n13150), .A2(n13316), .ZN(n13153) );
  INV_X1 U15335 ( .A(n13151), .ZN(n13346) );
  NOR2_X1 U15336 ( .A1(n14367), .A2(n13346), .ZN(n13157) );
  AOI21_X1 U15337 ( .B1(n14367), .B2(P2_REG2_REG_31__SCAN_IN), .A(n13157), 
        .ZN(n13152) );
  OAI211_X1 U15338 ( .C1(n6806), .C2(n13311), .A(n13153), .B(n13152), .ZN(
        P2_U3234) );
  OAI211_X1 U15339 ( .C1(n13436), .C2(n13155), .A(n9550), .B(n13154), .ZN(
        n13347) );
  NOR2_X1 U15340 ( .A1(n13281), .A2(n13156), .ZN(n13158) );
  AOI211_X1 U15341 ( .C1(n13159), .C2(n14355), .A(n13158), .B(n13157), .ZN(
        n13160) );
  OAI21_X1 U15342 ( .B1(n13347), .B2(n13330), .A(n13160), .ZN(P2_U3235) );
  XNOR2_X1 U15343 ( .A(n13162), .B(n13161), .ZN(n13355) );
  AOI22_X1 U15344 ( .A1(n13356), .A2(n14355), .B1(n14367), .B2(
        P2_REG2_REG_28__SCAN_IN), .ZN(n13178) );
  INV_X1 U15345 ( .A(n13164), .ZN(n13165) );
  AOI211_X1 U15346 ( .C1(n13356), .C2(n13186), .A(n9445), .B(n13165), .ZN(
        n13358) );
  INV_X1 U15347 ( .A(n13358), .ZN(n13168) );
  OAI22_X1 U15348 ( .A1(n13168), .A2(n13167), .B1(n13323), .B2(n13166), .ZN(
        n13176) );
  NAND2_X1 U15349 ( .A1(n13169), .A2(n13335), .ZN(n13175) );
  AOI21_X1 U15350 ( .B1(n13180), .B2(n13171), .A(n13170), .ZN(n13174) );
  INV_X1 U15351 ( .A(n13172), .ZN(n13173) );
  OAI21_X1 U15352 ( .B1(n13175), .B2(n13174), .A(n13173), .ZN(n13360) );
  OAI21_X1 U15353 ( .B1(n13176), .B2(n13360), .A(n13281), .ZN(n13177) );
  OAI211_X1 U15354 ( .C1(n13355), .C2(n13342), .A(n13178), .B(n13177), .ZN(
        P2_U3237) );
  XOR2_X1 U15355 ( .A(n13181), .B(n13179), .Z(n13365) );
  INV_X1 U15356 ( .A(n13365), .ZN(n13193) );
  OAI21_X1 U15357 ( .B1(n13182), .B2(n13181), .A(n13180), .ZN(n13183) );
  NAND2_X1 U15358 ( .A1(n13183), .A2(n13335), .ZN(n13185) );
  NAND2_X1 U15359 ( .A1(n13185), .A2(n13184), .ZN(n13363) );
  AOI211_X1 U15360 ( .C1(n13187), .C2(n13201), .A(n13326), .B(n13163), .ZN(
        n13364) );
  NAND2_X1 U15361 ( .A1(n13364), .A2(n14362), .ZN(n13190) );
  AOI22_X1 U15362 ( .A1(n14367), .A2(P2_REG2_REG_27__SCAN_IN), .B1(n14354), 
        .B2(n13188), .ZN(n13189) );
  OAI211_X1 U15363 ( .C1(n13442), .C2(n13311), .A(n13190), .B(n13189), .ZN(
        n13191) );
  AOI21_X1 U15364 ( .B1(n13363), .B2(n13281), .A(n13191), .ZN(n13192) );
  OAI21_X1 U15365 ( .B1(n13193), .B2(n13342), .A(n13192), .ZN(P2_U3238) );
  INV_X1 U15366 ( .A(n13196), .ZN(n13194) );
  XNOR2_X1 U15367 ( .A(n13195), .B(n13194), .ZN(n13370) );
  XNOR2_X1 U15368 ( .A(n13197), .B(n13196), .ZN(n13199) );
  AOI21_X1 U15369 ( .B1(n13199), .B2(n13335), .A(n13198), .ZN(n13369) );
  INV_X1 U15370 ( .A(n13369), .ZN(n13208) );
  NAND2_X1 U15371 ( .A1(n13216), .A2(n13205), .ZN(n13200) );
  NAND3_X1 U15372 ( .A1(n13201), .A2(n9550), .A3(n13200), .ZN(n13368) );
  NAND2_X1 U15373 ( .A1(n14367), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n13202) );
  OAI21_X1 U15374 ( .B1(n13323), .B2(n13203), .A(n13202), .ZN(n13204) );
  AOI21_X1 U15375 ( .B1(n13205), .B2(n14355), .A(n13204), .ZN(n13206) );
  OAI21_X1 U15376 ( .B1(n13368), .B2(n13330), .A(n13206), .ZN(n13207) );
  AOI21_X1 U15377 ( .B1(n13208), .B2(n13281), .A(n13207), .ZN(n13209) );
  OAI21_X1 U15378 ( .B1(n13370), .B2(n13342), .A(n13209), .ZN(P2_U3239) );
  XNOR2_X1 U15379 ( .A(n13210), .B(n13211), .ZN(n13377) );
  XNOR2_X1 U15380 ( .A(n13212), .B(n13211), .ZN(n13214) );
  OAI21_X1 U15381 ( .B1(n13214), .B2(n14351), .A(n13213), .ZN(n13373) );
  OR2_X1 U15382 ( .A1(n13220), .A2(n13228), .ZN(n13215) );
  AND3_X1 U15383 ( .A1(n13216), .A2(n13215), .A3(n9550), .ZN(n13374) );
  NAND2_X1 U15384 ( .A1(n13374), .A2(n14362), .ZN(n13219) );
  AOI22_X1 U15385 ( .A1(n14367), .A2(P2_REG2_REG_25__SCAN_IN), .B1(n14354), 
        .B2(n13217), .ZN(n13218) );
  OAI211_X1 U15386 ( .C1(n13220), .C2(n13311), .A(n13219), .B(n13218), .ZN(
        n13221) );
  AOI21_X1 U15387 ( .B1(n13373), .B2(n13281), .A(n13221), .ZN(n13222) );
  OAI21_X1 U15388 ( .B1(n13377), .B2(n13342), .A(n13222), .ZN(P2_U3240) );
  XNOR2_X1 U15389 ( .A(n13223), .B(n13224), .ZN(n13380) );
  XNOR2_X1 U15390 ( .A(n13225), .B(n13224), .ZN(n13227) );
  AOI21_X1 U15391 ( .B1(n13227), .B2(n13335), .A(n13226), .ZN(n13379) );
  INV_X1 U15392 ( .A(n13379), .ZN(n13236) );
  AND2_X1 U15393 ( .A1(n7436), .A2(n13233), .ZN(n13229) );
  OR3_X1 U15394 ( .A1(n13229), .A2(n13228), .A3(n9445), .ZN(n13378) );
  NAND2_X1 U15395 ( .A1(n14367), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n13230) );
  OAI21_X1 U15396 ( .B1(n13323), .B2(n13231), .A(n13230), .ZN(n13232) );
  AOI21_X1 U15397 ( .B1(n13233), .B2(n14355), .A(n13232), .ZN(n13234) );
  OAI21_X1 U15398 ( .B1(n13378), .B2(n13330), .A(n13234), .ZN(n13235) );
  AOI21_X1 U15399 ( .B1(n13236), .B2(n13281), .A(n13235), .ZN(n13237) );
  OAI21_X1 U15400 ( .B1(n13342), .B2(n13380), .A(n13237), .ZN(P2_U3241) );
  XOR2_X1 U15401 ( .A(n13239), .B(n13238), .Z(n13387) );
  XNOR2_X1 U15402 ( .A(n13240), .B(n13239), .ZN(n13242) );
  OAI21_X1 U15403 ( .B1(n13242), .B2(n14351), .A(n13241), .ZN(n13383) );
  AOI21_X1 U15404 ( .B1(n13259), .B2(n13385), .A(n13326), .ZN(n13243) );
  AND2_X1 U15405 ( .A1(n13243), .A2(n7436), .ZN(n13384) );
  NAND2_X1 U15406 ( .A1(n13384), .A2(n14362), .ZN(n13246) );
  AOI22_X1 U15407 ( .A1(n14367), .A2(P2_REG2_REG_23__SCAN_IN), .B1(n14354), 
        .B2(n13244), .ZN(n13245) );
  OAI211_X1 U15408 ( .C1(n13247), .C2(n13311), .A(n13246), .B(n13245), .ZN(
        n13248) );
  AOI21_X1 U15409 ( .B1(n13383), .B2(n13281), .A(n13248), .ZN(n13249) );
  OAI21_X1 U15410 ( .B1(n13387), .B2(n13342), .A(n13249), .ZN(P2_U3242) );
  NAND2_X1 U15411 ( .A1(n13251), .A2(n13250), .ZN(n13252) );
  NAND2_X1 U15412 ( .A1(n13253), .A2(n13252), .ZN(n13390) );
  NAND2_X1 U15413 ( .A1(n13254), .A2(n7960), .ZN(n13255) );
  NAND3_X1 U15414 ( .A1(n13256), .A2(n13335), .A3(n13255), .ZN(n13258) );
  INV_X1 U15415 ( .A(n13389), .ZN(n13266) );
  OAI211_X1 U15416 ( .C1(n6575), .C2(n13456), .A(n9550), .B(n13259), .ZN(
        n13388) );
  OAI22_X1 U15417 ( .A1(n13261), .A2(n13323), .B1(n13260), .B2(n13281), .ZN(
        n13262) );
  AOI21_X1 U15418 ( .B1(n13263), .B2(n14355), .A(n13262), .ZN(n13264) );
  OAI21_X1 U15419 ( .B1(n13388), .B2(n13330), .A(n13264), .ZN(n13265) );
  AOI21_X1 U15420 ( .B1(n13266), .B2(n13281), .A(n13265), .ZN(n13267) );
  OAI21_X1 U15421 ( .B1(n13342), .B2(n13390), .A(n13267), .ZN(P2_U3243) );
  XNOR2_X1 U15422 ( .A(n13268), .B(n13270), .ZN(n13393) );
  INV_X1 U15423 ( .A(n13393), .ZN(n13284) );
  NAND3_X1 U15424 ( .A1(n13286), .A2(n13270), .A3(n13269), .ZN(n13271) );
  NAND2_X1 U15425 ( .A1(n13272), .A2(n13271), .ZN(n13274) );
  AOI21_X1 U15426 ( .B1(n13274), .B2(n13335), .A(n13273), .ZN(n13395) );
  INV_X1 U15427 ( .A(n13395), .ZN(n13282) );
  NAND2_X1 U15428 ( .A1(n13292), .A2(n13459), .ZN(n13275) );
  NAND2_X1 U15429 ( .A1(n13275), .A2(n9550), .ZN(n13276) );
  OR2_X1 U15430 ( .A1(n6575), .A2(n13276), .ZN(n13394) );
  AOI22_X1 U15431 ( .A1(n13277), .A2(n14354), .B1(P2_REG2_REG_21__SCAN_IN), 
        .B2(n14367), .ZN(n13279) );
  NAND2_X1 U15432 ( .A1(n13459), .A2(n14355), .ZN(n13278) );
  OAI211_X1 U15433 ( .C1(n13394), .C2(n13330), .A(n13279), .B(n13278), .ZN(
        n13280) );
  AOI21_X1 U15434 ( .B1(n13282), .B2(n13281), .A(n13280), .ZN(n13283) );
  OAI21_X1 U15435 ( .B1(n13342), .B2(n13284), .A(n13283), .ZN(P2_U3244) );
  XNOR2_X1 U15436 ( .A(n13285), .B(n13289), .ZN(n13404) );
  INV_X1 U15437 ( .A(n13286), .ZN(n13287) );
  AOI21_X1 U15438 ( .B1(n13289), .B2(n13288), .A(n13287), .ZN(n13291) );
  OAI21_X1 U15439 ( .B1(n13291), .B2(n14351), .A(n13290), .ZN(n13400) );
  AOI21_X1 U15440 ( .B1(n13309), .B2(n13402), .A(n13326), .ZN(n13293) );
  AND2_X1 U15441 ( .A1(n13293), .A2(n13292), .ZN(n13401) );
  NAND2_X1 U15442 ( .A1(n13401), .A2(n14362), .ZN(n13298) );
  OAI22_X1 U15443 ( .A1(n13295), .A2(n13323), .B1(n13294), .B2(n13281), .ZN(
        n13296) );
  AOI21_X1 U15444 ( .B1(n13402), .B2(n14355), .A(n13296), .ZN(n13297) );
  NAND2_X1 U15445 ( .A1(n13298), .A2(n13297), .ZN(n13299) );
  AOI21_X1 U15446 ( .B1(n13400), .B2(n13281), .A(n13299), .ZN(n13300) );
  OAI21_X1 U15447 ( .B1(n13342), .B2(n13404), .A(n13300), .ZN(P2_U3245) );
  XNOR2_X1 U15448 ( .A(n13301), .B(n13302), .ZN(n13405) );
  XNOR2_X1 U15449 ( .A(n13303), .B(n13302), .ZN(n13305) );
  OAI21_X1 U15450 ( .B1(n13305), .B2(n14351), .A(n13304), .ZN(n13306) );
  AOI21_X1 U15451 ( .B1(n13307), .B2(n13405), .A(n13306), .ZN(n13409) );
  INV_X1 U15452 ( .A(n13308), .ZN(n13328) );
  INV_X1 U15453 ( .A(n13309), .ZN(n13310) );
  AOI21_X1 U15454 ( .B1(n13406), .B2(n13328), .A(n13310), .ZN(n13407) );
  NOR2_X1 U15455 ( .A1(n8168), .A2(n13311), .ZN(n13315) );
  OAI22_X1 U15456 ( .A1(n13313), .A2(n13323), .B1(n13281), .B2(n13312), .ZN(
        n13314) );
  AOI211_X1 U15457 ( .C1(n13407), .C2(n13316), .A(n13315), .B(n13314), .ZN(
        n13319) );
  NAND2_X1 U15458 ( .A1(n13405), .A2(n13317), .ZN(n13318) );
  OAI211_X1 U15459 ( .C1(n13409), .C2(n14367), .A(n13319), .B(n13318), .ZN(
        P2_U3246) );
  OR2_X1 U15460 ( .A1(n13320), .A2(n13334), .ZN(n13321) );
  NAND2_X1 U15461 ( .A1(n13322), .A2(n13321), .ZN(n13411) );
  INV_X1 U15462 ( .A(n13411), .ZN(n13341) );
  INV_X1 U15463 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n13325) );
  OAI22_X1 U15464 ( .A1(n13281), .A2(n13325), .B1(n13324), .B2(n13323), .ZN(
        n13332) );
  AOI21_X1 U15465 ( .B1(n6523), .B2(n13327), .A(n13326), .ZN(n13329) );
  NAND2_X1 U15466 ( .A1(n13329), .A2(n13328), .ZN(n13414) );
  NOR2_X1 U15467 ( .A1(n13414), .A2(n13330), .ZN(n13331) );
  AOI211_X1 U15468 ( .C1(n14355), .C2(n6523), .A(n13332), .B(n13331), .ZN(
        n13340) );
  XNOR2_X1 U15469 ( .A(n13334), .B(n13333), .ZN(n13336) );
  NAND2_X1 U15470 ( .A1(n13336), .A2(n13335), .ZN(n13338) );
  NAND2_X1 U15471 ( .A1(n13338), .A2(n13337), .ZN(n13416) );
  NAND2_X1 U15472 ( .A1(n13416), .A2(n13281), .ZN(n13339) );
  OAI211_X1 U15473 ( .C1(n13342), .C2(n13341), .A(n13340), .B(n13339), .ZN(
        P2_U3247) );
  INV_X1 U15474 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n13344) );
  MUX2_X1 U15475 ( .A(n13344), .B(n13343), .S(n14829), .Z(n13345) );
  OAI21_X1 U15476 ( .B1(n6806), .B2(n13423), .A(n13345), .ZN(P2_U3530) );
  AND2_X1 U15477 ( .A1(n13347), .A2(n13346), .ZN(n13433) );
  MUX2_X1 U15478 ( .A(n13348), .B(n13433), .S(n14829), .Z(n13349) );
  OAI21_X1 U15479 ( .B1(n13436), .B2(n13423), .A(n13349), .ZN(P2_U3529) );
  AOI21_X1 U15480 ( .B1(n14810), .B2(n13351), .A(n13350), .ZN(n13352) );
  OAI211_X1 U15481 ( .C1(n13354), .C2(n14791), .A(n13353), .B(n13352), .ZN(
        n13437) );
  MUX2_X1 U15482 ( .A(P2_REG1_REG_29__SCAN_IN), .B(n13437), .S(n14829), .Z(
        P2_U3528) );
  MUX2_X1 U15483 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n13438), .S(n14829), .Z(
        P2_U3527) );
  MUX2_X1 U15484 ( .A(n13366), .B(n13439), .S(n14829), .Z(n13367) );
  OAI21_X1 U15485 ( .B1(n13442), .B2(n13423), .A(n13367), .ZN(P2_U3526) );
  OAI211_X1 U15486 ( .C1(n13370), .C2(n14791), .A(n13369), .B(n13368), .ZN(
        n13443) );
  MUX2_X1 U15487 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n13443), .S(n14829), .Z(
        n13371) );
  INV_X1 U15488 ( .A(n13371), .ZN(n13372) );
  OAI21_X1 U15489 ( .B1(n13446), .B2(n13423), .A(n13372), .ZN(P2_U3525) );
  AOI211_X1 U15490 ( .C1(n14810), .C2(n13375), .A(n13374), .B(n13373), .ZN(
        n13376) );
  OAI21_X1 U15491 ( .B1(n14791), .B2(n13377), .A(n13376), .ZN(n13447) );
  MUX2_X1 U15492 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n13447), .S(n14829), .Z(
        P2_U3524) );
  OAI211_X1 U15493 ( .C1(n14791), .C2(n13380), .A(n13379), .B(n13378), .ZN(
        n13448) );
  MUX2_X1 U15494 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n13448), .S(n14829), .Z(
        n13381) );
  INV_X1 U15495 ( .A(n13381), .ZN(n13382) );
  OAI21_X1 U15496 ( .B1(n13451), .B2(n13423), .A(n13382), .ZN(P2_U3523) );
  AOI211_X1 U15497 ( .C1(n14810), .C2(n13385), .A(n13384), .B(n13383), .ZN(
        n13386) );
  OAI21_X1 U15498 ( .B1(n14791), .B2(n13387), .A(n13386), .ZN(n13452) );
  MUX2_X1 U15499 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n13452), .S(n14829), .Z(
        P2_U3522) );
  OAI211_X1 U15500 ( .C1(n13390), .C2(n14791), .A(n13389), .B(n13388), .ZN(
        n13453) );
  MUX2_X1 U15501 ( .A(n13453), .B(P2_REG1_REG_22__SCAN_IN), .S(n14827), .Z(
        n13391) );
  INV_X1 U15502 ( .A(n13391), .ZN(n13392) );
  OAI21_X1 U15503 ( .B1(n13456), .B2(n13423), .A(n13392), .ZN(P2_U3521) );
  NAND2_X1 U15504 ( .A1(n13393), .A2(n14378), .ZN(n13396) );
  NAND3_X1 U15505 ( .A1(n13396), .A2(n13395), .A3(n13394), .ZN(n13457) );
  MUX2_X1 U15506 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n13457), .S(n14829), .Z(
        n13397) );
  AOI21_X1 U15507 ( .B1(n13398), .B2(n13459), .A(n13397), .ZN(n13399) );
  INV_X1 U15508 ( .A(n13399), .ZN(P2_U3520) );
  AOI211_X1 U15509 ( .C1(n14810), .C2(n13402), .A(n13401), .B(n13400), .ZN(
        n13403) );
  OAI21_X1 U15510 ( .B1(n14791), .B2(n13404), .A(n13403), .ZN(n13462) );
  MUX2_X1 U15511 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n13462), .S(n14829), .Z(
        P2_U3519) );
  INV_X1 U15512 ( .A(n13405), .ZN(n13410) );
  AOI22_X1 U15513 ( .A1(n13407), .A2(n9550), .B1(n14810), .B2(n13406), .ZN(
        n13408) );
  OAI211_X1 U15514 ( .C1(n14803), .C2(n13410), .A(n13409), .B(n13408), .ZN(
        n13463) );
  MUX2_X1 U15515 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n13463), .S(n14829), .Z(
        P2_U3518) );
  AND2_X1 U15516 ( .A1(n13411), .A2(n14378), .ZN(n13417) );
  NAND2_X1 U15517 ( .A1(n13412), .A2(n14810), .ZN(n13413) );
  NAND2_X1 U15518 ( .A1(n13414), .A2(n13413), .ZN(n13415) );
  MUX2_X1 U15519 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n13464), .S(n14829), .Z(
        P2_U3517) );
  AOI211_X1 U15520 ( .C1(n13420), .C2(n14378), .A(n13419), .B(n13418), .ZN(
        n13465) );
  MUX2_X1 U15521 ( .A(n13421), .B(n13465), .S(n14829), .Z(n13422) );
  OAI21_X1 U15522 ( .B1(n13469), .B2(n13423), .A(n13422), .ZN(P2_U3516) );
  NAND3_X1 U15523 ( .A1(n13425), .A2(n14378), .A3(n13424), .ZN(n13429) );
  NAND2_X1 U15524 ( .A1(n13426), .A2(n14810), .ZN(n13427) );
  NAND3_X1 U15525 ( .A1(n13429), .A2(n13428), .A3(n13427), .ZN(n13430) );
  NOR2_X1 U15526 ( .A1(n13431), .A2(n13430), .ZN(n13470) );
  MUX2_X1 U15527 ( .A(n15259), .B(n13470), .S(n14829), .Z(n13432) );
  INV_X1 U15528 ( .A(n13432), .ZN(P2_U3515) );
  MUX2_X1 U15529 ( .A(n13434), .B(n13433), .S(n14821), .Z(n13435) );
  OAI21_X1 U15530 ( .B1(n13436), .B2(n13468), .A(n13435), .ZN(P2_U3497) );
  MUX2_X1 U15531 ( .A(P2_REG0_REG_29__SCAN_IN), .B(n13437), .S(n14821), .Z(
        P2_U3496) );
  MUX2_X1 U15532 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n13438), .S(n14821), .Z(
        P2_U3495) );
  MUX2_X1 U15533 ( .A(n13440), .B(n13439), .S(n14821), .Z(n13441) );
  OAI21_X1 U15534 ( .B1(n13442), .B2(n13468), .A(n13441), .ZN(P2_U3494) );
  MUX2_X1 U15535 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n13443), .S(n14821), .Z(
        n13444) );
  INV_X1 U15536 ( .A(n13444), .ZN(n13445) );
  OAI21_X1 U15537 ( .B1(n13446), .B2(n13468), .A(n13445), .ZN(P2_U3493) );
  MUX2_X1 U15538 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n13447), .S(n14821), .Z(
        P2_U3492) );
  MUX2_X1 U15539 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n13448), .S(n14821), .Z(
        n13449) );
  INV_X1 U15540 ( .A(n13449), .ZN(n13450) );
  OAI21_X1 U15541 ( .B1(n13451), .B2(n13468), .A(n13450), .ZN(P2_U3491) );
  MUX2_X1 U15542 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n13452), .S(n14821), .Z(
        P2_U3490) );
  MUX2_X1 U15543 ( .A(n13453), .B(P2_REG0_REG_22__SCAN_IN), .S(n14819), .Z(
        n13454) );
  INV_X1 U15544 ( .A(n13454), .ZN(n13455) );
  OAI21_X1 U15545 ( .B1(n13456), .B2(n13468), .A(n13455), .ZN(P2_U3489) );
  MUX2_X1 U15546 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n13457), .S(n14821), .Z(
        n13458) );
  AOI21_X1 U15547 ( .B1(n13460), .B2(n13459), .A(n13458), .ZN(n13461) );
  INV_X1 U15548 ( .A(n13461), .ZN(P2_U3488) );
  MUX2_X1 U15549 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n13462), .S(n14821), .Z(
        P2_U3487) );
  MUX2_X1 U15550 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n13463), .S(n14821), .Z(
        P2_U3486) );
  MUX2_X1 U15551 ( .A(n13464), .B(P2_REG0_REG_18__SCAN_IN), .S(n14819), .Z(
        P2_U3484) );
  INV_X1 U15552 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n13466) );
  MUX2_X1 U15553 ( .A(n13466), .B(n13465), .S(n14821), .Z(n13467) );
  OAI21_X1 U15554 ( .B1(n13469), .B2(n13468), .A(n13467), .ZN(P2_U3481) );
  INV_X1 U15555 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n13471) );
  MUX2_X1 U15556 ( .A(n13471), .B(n13470), .S(n14821), .Z(n13472) );
  INV_X1 U15557 ( .A(n13472), .ZN(P2_U3478) );
  INV_X1 U15558 ( .A(n8795), .ZN(n14262) );
  NOR4_X1 U15559 ( .A1(n13474), .A2(P2_IR_REG_30__SCAN_IN), .A3(n13473), .A4(
        P2_U3088), .ZN(n13475) );
  AOI21_X1 U15560 ( .B1(P1_DATAO_REG_31__SCAN_IN), .B2(n13480), .A(n13475), 
        .ZN(n13476) );
  OAI21_X1 U15561 ( .B1(n14262), .B2(n6534), .A(n13476), .ZN(P2_U3296) );
  OAI222_X1 U15562 ( .A1(n6534), .A2(n13478), .B1(P2_U3088), .B2(n7470), .C1(
        n13477), .C2(n11904), .ZN(P2_U3298) );
  AOI21_X1 U15563 ( .B1(n13480), .B2(P1_DATAO_REG_28__SCAN_IN), .A(n13479), 
        .ZN(n13481) );
  OAI21_X1 U15564 ( .B1(n13482), .B2(n6534), .A(n13481), .ZN(P2_U3299) );
  INV_X1 U15565 ( .A(n13483), .ZN(n14263) );
  OAI222_X1 U15566 ( .A1(n11904), .A2(n13485), .B1(n6534), .B2(n14263), .C1(
        n13484), .C2(P2_U3088), .ZN(P2_U3300) );
  INV_X1 U15567 ( .A(n13486), .ZN(n14268) );
  OAI222_X1 U15568 ( .A1(n13488), .A2(P2_U3088), .B1(n6534), .B2(n14268), .C1(
        n13487), .C2(n11904), .ZN(P2_U3301) );
  INV_X1 U15569 ( .A(n13489), .ZN(n13490) );
  MUX2_X1 U15570 ( .A(n13490), .B(n15206), .S(P2_STATE_REG_SCAN_IN), .Z(
        P2_U3327) );
  INV_X1 U15571 ( .A(n13956), .ZN(n14151) );
  NAND2_X1 U15572 ( .A1(n13956), .A2(n13640), .ZN(n13492) );
  NAND2_X1 U15573 ( .A1(n13910), .A2(n6536), .ZN(n13491) );
  NAND2_X1 U15574 ( .A1(n13492), .A2(n13491), .ZN(n13493) );
  XNOR2_X1 U15575 ( .A(n13493), .B(n13637), .ZN(n13497) );
  NAND2_X1 U15576 ( .A1(n13956), .A2(n6536), .ZN(n13495) );
  NAND2_X1 U15577 ( .A1(n13910), .A2(n13636), .ZN(n13494) );
  NAND2_X1 U15578 ( .A1(n13495), .A2(n13494), .ZN(n13496) );
  NOR2_X1 U15579 ( .A1(n13497), .A2(n13496), .ZN(n13634) );
  AOI21_X1 U15580 ( .B1(n13497), .B2(n13496), .A(n13634), .ZN(n13611) );
  INV_X1 U15581 ( .A(n13500), .ZN(n13501) );
  INV_X1 U15582 ( .A(n14392), .ZN(n13514) );
  NAND2_X1 U15583 ( .A1(n14405), .A2(n13640), .ZN(n13504) );
  NAND2_X1 U15584 ( .A1(n13760), .A2(n6536), .ZN(n13503) );
  NAND2_X1 U15585 ( .A1(n13504), .A2(n13503), .ZN(n13505) );
  XNOR2_X1 U15586 ( .A(n13505), .B(n13591), .ZN(n13508) );
  NOR2_X1 U15587 ( .A1(n13506), .A2(n13548), .ZN(n13507) );
  AOI21_X1 U15588 ( .B1(n14405), .B2(n6536), .A(n13507), .ZN(n13509) );
  NAND2_X1 U15589 ( .A1(n13508), .A2(n13509), .ZN(n13515) );
  INV_X1 U15590 ( .A(n13508), .ZN(n13511) );
  INV_X1 U15591 ( .A(n13509), .ZN(n13510) );
  NAND2_X1 U15592 ( .A1(n13511), .A2(n13510), .ZN(n13512) );
  NAND2_X1 U15593 ( .A1(n13515), .A2(n13512), .ZN(n14391) );
  AOI22_X1 U15594 ( .A1(n13754), .A2(n13640), .B1(n6536), .B2(n13759), .ZN(
        n13516) );
  XOR2_X1 U15595 ( .A(n13637), .B(n13516), .Z(n13518) );
  OAI22_X1 U15596 ( .A1(n6967), .A2(n13549), .B1(n13517), .B2(n13548), .ZN(
        n13745) );
  NAND2_X1 U15597 ( .A1(n13890), .A2(n13640), .ZN(n13520) );
  NAND2_X1 U15598 ( .A1(n14106), .A2(n6536), .ZN(n13519) );
  NAND2_X1 U15599 ( .A1(n13520), .A2(n13519), .ZN(n13521) );
  XNOR2_X1 U15600 ( .A(n13521), .B(n13637), .ZN(n13525) );
  NAND2_X1 U15601 ( .A1(n13890), .A2(n6536), .ZN(n13523) );
  NAND2_X1 U15602 ( .A1(n14106), .A2(n13636), .ZN(n13522) );
  NAND2_X1 U15603 ( .A1(n13523), .A2(n13522), .ZN(n13524) );
  NOR2_X1 U15604 ( .A1(n13525), .A2(n13524), .ZN(n13526) );
  AOI21_X1 U15605 ( .B1(n13525), .B2(n13524), .A(n13526), .ZN(n13681) );
  INV_X1 U15606 ( .A(n13526), .ZN(n13691) );
  NAND2_X1 U15607 ( .A1(n14218), .A2(n13640), .ZN(n13528) );
  NAND2_X1 U15608 ( .A1(n14088), .A2(n6536), .ZN(n13527) );
  NAND2_X1 U15609 ( .A1(n13528), .A2(n13527), .ZN(n13529) );
  XNOR2_X1 U15610 ( .A(n13529), .B(n13591), .ZN(n13531) );
  AND2_X1 U15611 ( .A1(n14088), .A2(n13636), .ZN(n13530) );
  AOI21_X1 U15612 ( .B1(n14218), .B2(n6536), .A(n13530), .ZN(n13532) );
  NAND2_X1 U15613 ( .A1(n13531), .A2(n13532), .ZN(n13536) );
  INV_X1 U15614 ( .A(n13531), .ZN(n13534) );
  INV_X1 U15615 ( .A(n13532), .ZN(n13533) );
  NAND2_X1 U15616 ( .A1(n13534), .A2(n13533), .ZN(n13535) );
  NAND2_X1 U15617 ( .A1(n13536), .A2(n13535), .ZN(n13690) );
  INV_X1 U15618 ( .A(n13536), .ZN(n13537) );
  AOI22_X1 U15619 ( .A1(n14096), .A2(n6536), .B1(n13636), .B2(n14109), .ZN(
        n13542) );
  NAND2_X1 U15620 ( .A1(n14096), .A2(n13640), .ZN(n13539) );
  NAND2_X1 U15621 ( .A1(n14109), .A2(n6536), .ZN(n13538) );
  NAND2_X1 U15622 ( .A1(n13539), .A2(n13538), .ZN(n13540) );
  XNOR2_X1 U15623 ( .A(n13540), .B(n13637), .ZN(n13541) );
  XOR2_X1 U15624 ( .A(n13542), .B(n13541), .Z(n13724) );
  INV_X1 U15625 ( .A(n13541), .ZN(n13543) );
  OAI22_X1 U15626 ( .A1(n14079), .A2(n13549), .B1(n14210), .B2(n13548), .ZN(
        n13546) );
  OAI22_X1 U15627 ( .A1(n14079), .A2(n9939), .B1(n14210), .B2(n13549), .ZN(
        n13544) );
  XNOR2_X1 U15628 ( .A(n13544), .B(n13637), .ZN(n13545) );
  XOR2_X1 U15629 ( .A(n13546), .B(n13545), .Z(n13628) );
  NAND2_X1 U15630 ( .A1(n13629), .A2(n13628), .ZN(n13627) );
  NAND2_X1 U15631 ( .A1(n13627), .A2(n13547), .ZN(n13709) );
  OAI22_X1 U15632 ( .A1(n14061), .A2(n13549), .B1(n14074), .B2(n13548), .ZN(
        n13551) );
  OAI22_X1 U15633 ( .A1(n14061), .A2(n9939), .B1(n14074), .B2(n13549), .ZN(
        n13550) );
  XNOR2_X1 U15634 ( .A(n13550), .B(n13637), .ZN(n13552) );
  XOR2_X1 U15635 ( .A(n13551), .B(n13552), .Z(n13708) );
  NAND2_X1 U15636 ( .A1(n14190), .A2(n13640), .ZN(n13555) );
  NAND2_X1 U15637 ( .A1(n14025), .A2(n6536), .ZN(n13554) );
  NAND2_X1 U15638 ( .A1(n13555), .A2(n13554), .ZN(n13556) );
  XNOR2_X1 U15639 ( .A(n13556), .B(n13591), .ZN(n13559) );
  INV_X1 U15640 ( .A(n13559), .ZN(n13561) );
  AND2_X1 U15641 ( .A1(n14025), .A2(n13636), .ZN(n13557) );
  AOI21_X1 U15642 ( .B1(n14190), .B2(n6536), .A(n13557), .ZN(n13558) );
  INV_X1 U15643 ( .A(n13558), .ZN(n13560) );
  AOI21_X1 U15644 ( .B1(n13561), .B2(n13560), .A(n13562), .ZN(n13650) );
  INV_X1 U15645 ( .A(n13562), .ZN(n13715) );
  NAND2_X1 U15646 ( .A1(n14186), .A2(n13640), .ZN(n13564) );
  NAND2_X1 U15647 ( .A1(n13900), .A2(n6536), .ZN(n13563) );
  NAND2_X1 U15648 ( .A1(n13564), .A2(n13563), .ZN(n13565) );
  XNOR2_X1 U15649 ( .A(n13565), .B(n13591), .ZN(n13568) );
  AND2_X1 U15650 ( .A1(n13900), .A2(n13636), .ZN(n13566) );
  AOI21_X1 U15651 ( .B1(n14186), .B2(n6536), .A(n13566), .ZN(n13567) );
  NAND2_X1 U15652 ( .A1(n13568), .A2(n13567), .ZN(n13569) );
  OAI21_X1 U15653 ( .B1(n13568), .B2(n13567), .A(n13569), .ZN(n13714) );
  INV_X1 U15654 ( .A(n13569), .ZN(n13620) );
  NAND2_X1 U15655 ( .A1(n14181), .A2(n13640), .ZN(n13571) );
  NAND2_X1 U15656 ( .A1(n14026), .A2(n6536), .ZN(n13570) );
  NAND2_X1 U15657 ( .A1(n13571), .A2(n13570), .ZN(n13572) );
  XNOR2_X1 U15658 ( .A(n13572), .B(n13591), .ZN(n13574) );
  AND2_X1 U15659 ( .A1(n14026), .A2(n13636), .ZN(n13573) );
  AOI21_X1 U15660 ( .B1(n14181), .B2(n6536), .A(n13573), .ZN(n13575) );
  NAND2_X1 U15661 ( .A1(n13574), .A2(n13575), .ZN(n13701) );
  INV_X1 U15662 ( .A(n13574), .ZN(n13577) );
  INV_X1 U15663 ( .A(n13575), .ZN(n13576) );
  NAND2_X1 U15664 ( .A1(n13577), .A2(n13576), .ZN(n13578) );
  NAND2_X1 U15665 ( .A1(n14176), .A2(n13640), .ZN(n13580) );
  NAND2_X1 U15666 ( .A1(n13980), .A2(n6536), .ZN(n13579) );
  NAND2_X1 U15667 ( .A1(n13580), .A2(n13579), .ZN(n13581) );
  XNOR2_X1 U15668 ( .A(n13581), .B(n13591), .ZN(n13583) );
  AND2_X1 U15669 ( .A1(n13980), .A2(n13636), .ZN(n13582) );
  AOI21_X1 U15670 ( .B1(n14176), .B2(n6536), .A(n13582), .ZN(n13584) );
  NAND2_X1 U15671 ( .A1(n13583), .A2(n13584), .ZN(n13588) );
  INV_X1 U15672 ( .A(n13583), .ZN(n13586) );
  INV_X1 U15673 ( .A(n13584), .ZN(n13585) );
  NAND2_X1 U15674 ( .A1(n13586), .A2(n13585), .ZN(n13587) );
  NAND2_X1 U15675 ( .A1(n13588), .A2(n13587), .ZN(n13700) );
  INV_X1 U15676 ( .A(n13588), .ZN(n13672) );
  NAND2_X1 U15677 ( .A1(n14168), .A2(n13640), .ZN(n13590) );
  NAND2_X1 U15678 ( .A1(n13907), .A2(n6536), .ZN(n13589) );
  NAND2_X1 U15679 ( .A1(n13590), .A2(n13589), .ZN(n13592) );
  XNOR2_X1 U15680 ( .A(n13592), .B(n13591), .ZN(n13594) );
  AND2_X1 U15681 ( .A1(n13907), .A2(n13636), .ZN(n13593) );
  AOI21_X1 U15682 ( .B1(n14168), .B2(n6536), .A(n13593), .ZN(n13595) );
  NAND2_X1 U15683 ( .A1(n13594), .A2(n13595), .ZN(n13599) );
  INV_X1 U15684 ( .A(n13594), .ZN(n13597) );
  INV_X1 U15685 ( .A(n13595), .ZN(n13596) );
  NAND2_X1 U15686 ( .A1(n13597), .A2(n13596), .ZN(n13598) );
  NAND2_X1 U15687 ( .A1(n14162), .A2(n13640), .ZN(n13601) );
  NAND2_X1 U15688 ( .A1(n13979), .A2(n6536), .ZN(n13600) );
  NAND2_X1 U15689 ( .A1(n13601), .A2(n13600), .ZN(n13602) );
  XNOR2_X1 U15690 ( .A(n13602), .B(n13637), .ZN(n13607) );
  NAND2_X1 U15691 ( .A1(n14162), .A2(n6536), .ZN(n13605) );
  NAND2_X1 U15692 ( .A1(n13979), .A2(n13603), .ZN(n13604) );
  NAND2_X1 U15693 ( .A1(n13605), .A2(n13604), .ZN(n13606) );
  NOR2_X1 U15694 ( .A1(n13607), .A2(n13606), .ZN(n13608) );
  AOI21_X1 U15695 ( .B1(n13607), .B2(n13606), .A(n13608), .ZN(n13733) );
  INV_X1 U15696 ( .A(n13608), .ZN(n13609) );
  OAI21_X1 U15697 ( .B1(n13611), .B2(n13610), .A(n13635), .ZN(n13612) );
  INV_X1 U15698 ( .A(n13945), .ZN(n13886) );
  OAI22_X1 U15699 ( .A1(n13748), .A2(n13886), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13613), .ZN(n13615) );
  NOR2_X1 U15700 ( .A1(n14401), .A2(n13954), .ZN(n13614) );
  AOI211_X1 U15701 ( .C1(n13750), .C2(n13979), .A(n13615), .B(n13614), .ZN(
        n13616) );
  INV_X1 U15702 ( .A(n14181), .ZN(n14018) );
  INV_X1 U15703 ( .A(n13617), .ZN(n13622) );
  NOR3_X1 U15704 ( .A1(n13618), .A2(n13620), .A3(n13619), .ZN(n13621) );
  OAI21_X1 U15705 ( .B1(n13622), .B2(n13621), .A(n14395), .ZN(n13626) );
  INV_X1 U15706 ( .A(n13900), .ZN(n13876) );
  OAI22_X1 U15707 ( .A1(n13876), .A2(n14561), .B1(n13881), .B2(n14581), .ZN(
        n14011) );
  INV_X1 U15708 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n13623) );
  OAI22_X1 U15709 ( .A1(n14401), .A2(n14015), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13623), .ZN(n13624) );
  AOI21_X1 U15710 ( .B1(n14011), .B2(n14397), .A(n13624), .ZN(n13625) );
  OAI211_X1 U15711 ( .C1(n14018), .C2(n13743), .A(n13626), .B(n13625), .ZN(
        P1_U3216) );
  OAI211_X1 U15712 ( .C1(n13629), .C2(n13628), .A(n13627), .B(n14395), .ZN(
        n13633) );
  NAND2_X1 U15713 ( .A1(n13750), .A2(n14109), .ZN(n13630) );
  NAND2_X1 U15714 ( .A1(P1_U3086), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n13850)
         );
  OAI211_X1 U15715 ( .C1(n14074), .C2(n13748), .A(n13630), .B(n13850), .ZN(
        n13631) );
  AOI21_X1 U15716 ( .B1(n14072), .B2(n13740), .A(n13631), .ZN(n13632) );
  OAI211_X1 U15717 ( .C1(n14079), .C2(n13743), .A(n13633), .B(n13632), .ZN(
        P1_U3219) );
  AOI22_X1 U15718 ( .A1(n14143), .A2(n6536), .B1(n13636), .B2(n13945), .ZN(
        n13638) );
  XNOR2_X1 U15719 ( .A(n13638), .B(n13637), .ZN(n13642) );
  AOI22_X1 U15720 ( .A1(n14143), .A2(n13640), .B1(n6536), .B2(n13945), .ZN(
        n13641) );
  XNOR2_X1 U15721 ( .A(n13642), .B(n13641), .ZN(n13643) );
  NAND2_X1 U15722 ( .A1(n13910), .A2(n14107), .ZN(n13645) );
  NAND2_X1 U15723 ( .A1(n13758), .A2(n14108), .ZN(n13644) );
  NAND2_X1 U15724 ( .A1(n13645), .A2(n13644), .ZN(n13929) );
  AOI22_X1 U15725 ( .A1(n14397), .A2(n13929), .B1(P1_REG3_REG_28__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13646) );
  OAI21_X1 U15726 ( .B1(n14401), .B2(n13931), .A(n13646), .ZN(n13647) );
  AOI21_X1 U15727 ( .B1(n14143), .B2(n14398), .A(n13647), .ZN(n13648) );
  OAI21_X1 U15728 ( .B1(n13649), .B2(n13756), .A(n13648), .ZN(P1_U3220) );
  INV_X1 U15729 ( .A(n14190), .ZN(n14045) );
  OAI21_X1 U15730 ( .B1(n13651), .B2(n13650), .A(n13716), .ZN(n13652) );
  NAND2_X1 U15731 ( .A1(n13652), .A2(n14395), .ZN(n13657) );
  OAI22_X1 U15732 ( .A1(n13876), .A2(n14581), .B1(n14074), .B2(n14561), .ZN(
        n14040) );
  INV_X1 U15733 ( .A(n14043), .ZN(n13654) );
  OAI22_X1 U15734 ( .A1(n13654), .A2(n14401), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13653), .ZN(n13655) );
  AOI21_X1 U15735 ( .B1(n14040), .B2(n14397), .A(n13655), .ZN(n13656) );
  OAI211_X1 U15736 ( .C1(n14045), .C2(n13743), .A(n13657), .B(n13656), .ZN(
        P1_U3223) );
  NAND2_X1 U15737 ( .A1(P1_REG3_REG_12__SCAN_IN), .A2(P1_U3086), .ZN(n14467)
         );
  NAND2_X1 U15738 ( .A1(n14397), .A2(n13658), .ZN(n13659) );
  OAI211_X1 U15739 ( .C1(n14401), .C2(n13660), .A(n14467), .B(n13659), .ZN(
        n13666) );
  INV_X1 U15740 ( .A(n13661), .ZN(n13662) );
  AOI211_X1 U15741 ( .C1(n13664), .C2(n13663), .A(n13756), .B(n13662), .ZN(
        n13665) );
  AOI211_X1 U15742 ( .C1(n13667), .C2(n14398), .A(n13666), .B(n13665), .ZN(
        n13668) );
  INV_X1 U15743 ( .A(n13668), .ZN(P1_U3224) );
  INV_X1 U15744 ( .A(n14168), .ZN(n13987) );
  INV_X1 U15745 ( .A(n13669), .ZN(n13674) );
  NOR3_X1 U15746 ( .A1(n13670), .A2(n13672), .A3(n13671), .ZN(n13673) );
  OAI21_X1 U15747 ( .B1(n13674), .B2(n13673), .A(n14395), .ZN(n13679) );
  INV_X1 U15748 ( .A(n13675), .ZN(n13985) );
  AOI22_X1 U15749 ( .A1(n13718), .A2(n13979), .B1(P1_REG3_REG_25__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13676) );
  OAI21_X1 U15750 ( .B1(n13720), .B2(n13881), .A(n13676), .ZN(n13677) );
  AOI21_X1 U15751 ( .B1(n13985), .B2(n13740), .A(n13677), .ZN(n13678) );
  OAI211_X1 U15752 ( .C1(n13987), .C2(n13743), .A(n13679), .B(n13678), .ZN(
        P1_U3225) );
  OAI21_X1 U15753 ( .B1(n13681), .B2(n13680), .A(n13692), .ZN(n13682) );
  NAND2_X1 U15754 ( .A1(n13682), .A2(n14395), .ZN(n13689) );
  OAI21_X1 U15755 ( .B1(n13748), .B2(n13684), .A(n13683), .ZN(n13687) );
  NOR2_X1 U15756 ( .A1(n14401), .A2(n13685), .ZN(n13686) );
  AOI211_X1 U15757 ( .C1(n13750), .C2(n13759), .A(n13687), .B(n13686), .ZN(
        n13688) );
  OAI211_X1 U15758 ( .C1(n14223), .C2(n13743), .A(n13689), .B(n13688), .ZN(
        P1_U3226) );
  INV_X1 U15759 ( .A(n14218), .ZN(n14120) );
  AND3_X1 U15760 ( .A1(n13692), .A2(n13691), .A3(n13690), .ZN(n13693) );
  OAI21_X1 U15761 ( .B1(n13694), .B2(n13693), .A(n14395), .ZN(n13699) );
  INV_X1 U15762 ( .A(n14109), .ZN(n14073) );
  OAI21_X1 U15763 ( .B1(n14073), .B2(n13748), .A(n13695), .ZN(n13697) );
  NOR2_X1 U15764 ( .A1(n14401), .A2(n14116), .ZN(n13696) );
  AOI211_X1 U15765 ( .C1(n13750), .C2(n14106), .A(n13697), .B(n13696), .ZN(
        n13698) );
  OAI211_X1 U15766 ( .C1(n14120), .C2(n13743), .A(n13699), .B(n13698), .ZN(
        P1_U3228) );
  AND3_X1 U15767 ( .A1(n13617), .A2(n13701), .A3(n13700), .ZN(n13702) );
  OAI21_X1 U15768 ( .B1(n13670), .B2(n13702), .A(n14395), .ZN(n13707) );
  INV_X1 U15769 ( .A(n13703), .ZN(n14001) );
  AOI22_X1 U15770 ( .A1(n14107), .A2(n14026), .B1(n13907), .B2(n14108), .ZN(
        n13995) );
  INV_X1 U15771 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n13704) );
  OAI22_X1 U15772 ( .A1(n13995), .A2(n13738), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13704), .ZN(n13705) );
  AOI21_X1 U15773 ( .B1(n14001), .B2(n13740), .A(n13705), .ZN(n13706) );
  OAI211_X1 U15774 ( .C1(n6982), .C2(n13743), .A(n13707), .B(n13706), .ZN(
        P1_U3229) );
  XNOR2_X1 U15775 ( .A(n13709), .B(n13708), .ZN(n13713) );
  INV_X1 U15776 ( .A(n14025), .ZN(n13874) );
  OAI22_X1 U15777 ( .A1(n13874), .A2(n14581), .B1(n14210), .B2(n14561), .ZN(
        n14196) );
  AOI22_X1 U15778 ( .A1(n14196), .A2(n14397), .B1(P1_REG3_REG_20__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13710) );
  OAI21_X1 U15779 ( .B1(n14057), .B2(n14401), .A(n13710), .ZN(n13711) );
  AOI21_X1 U15780 ( .B1(n14197), .B2(n14398), .A(n13711), .ZN(n13712) );
  OAI21_X1 U15781 ( .B1(n13713), .B2(n13756), .A(n13712), .ZN(P1_U3233) );
  AND3_X1 U15782 ( .A1(n13716), .A2(n13715), .A3(n13714), .ZN(n13717) );
  OAI21_X1 U15783 ( .B1(n13618), .B2(n13717), .A(n14395), .ZN(n13723) );
  AOI22_X1 U15784 ( .A1(n13718), .A2(n14026), .B1(P1_REG3_REG_22__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13719) );
  OAI21_X1 U15785 ( .B1(n13720), .B2(n13874), .A(n13719), .ZN(n13721) );
  AOI21_X1 U15786 ( .B1(n14031), .B2(n13740), .A(n13721), .ZN(n13722) );
  OAI211_X1 U15787 ( .C1(n13743), .C2(n14033), .A(n13723), .B(n13722), .ZN(
        P1_U3235) );
  AOI21_X1 U15788 ( .B1(n13725), .B2(n13724), .A(n6686), .ZN(n13730) );
  NAND2_X1 U15789 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n13827)
         );
  OAI21_X1 U15790 ( .B1(n14210), .B2(n13748), .A(n13827), .ZN(n13726) );
  AOI21_X1 U15791 ( .B1(n13750), .B2(n14088), .A(n13726), .ZN(n13727) );
  OAI21_X1 U15792 ( .B1(n14092), .B2(n14401), .A(n13727), .ZN(n13728) );
  AOI21_X1 U15793 ( .B1(n14096), .B2(n14398), .A(n13728), .ZN(n13729) );
  OAI21_X1 U15794 ( .B1(n13730), .B2(n13756), .A(n13729), .ZN(P1_U3238) );
  INV_X1 U15795 ( .A(n14162), .ZN(n13744) );
  OAI21_X1 U15796 ( .B1(n13733), .B2(n13732), .A(n13731), .ZN(n13734) );
  NAND2_X1 U15797 ( .A1(n13734), .A2(n14395), .ZN(n13742) );
  INV_X1 U15798 ( .A(n13735), .ZN(n13970) );
  NAND2_X1 U15799 ( .A1(n13907), .A2(n14107), .ZN(n13737) );
  NAND2_X1 U15800 ( .A1(n13910), .A2(n14108), .ZN(n13736) );
  AND2_X1 U15801 ( .A1(n13737), .A2(n13736), .ZN(n14159) );
  OAI22_X1 U15802 ( .A1(n13738), .A2(n14159), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n15274), .ZN(n13739) );
  AOI21_X1 U15803 ( .B1(n13970), .B2(n13740), .A(n13739), .ZN(n13741) );
  OAI211_X1 U15804 ( .C1(n13744), .C2(n13743), .A(n13742), .B(n13741), .ZN(
        P1_U3240) );
  XNOR2_X1 U15805 ( .A(n13746), .B(n13745), .ZN(n13757) );
  OAI22_X1 U15806 ( .A1(n13748), .A2(n13864), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13747), .ZN(n13749) );
  AOI21_X1 U15807 ( .B1(n13750), .B2(n13760), .A(n13749), .ZN(n13751) );
  OAI21_X1 U15808 ( .B1(n13752), .B2(n14401), .A(n13751), .ZN(n13753) );
  AOI21_X1 U15809 ( .B1(n13754), .B2(n14398), .A(n13753), .ZN(n13755) );
  OAI21_X1 U15810 ( .B1(n13757), .B2(n13756), .A(n13755), .ZN(P1_U3241) );
  MUX2_X1 U15811 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(n13855), .S(P1_U4016), .Z(
        P1_U3591) );
  MUX2_X1 U15812 ( .A(n13919), .B(P1_DATAO_REG_30__SCAN_IN), .S(n13773), .Z(
        P1_U3590) );
  MUX2_X1 U15813 ( .A(n13758), .B(P1_DATAO_REG_29__SCAN_IN), .S(n13773), .Z(
        P1_U3589) );
  MUX2_X1 U15814 ( .A(n13945), .B(P1_DATAO_REG_28__SCAN_IN), .S(n13773), .Z(
        P1_U3588) );
  MUX2_X1 U15815 ( .A(n13910), .B(P1_DATAO_REG_27__SCAN_IN), .S(n13773), .Z(
        P1_U3587) );
  MUX2_X1 U15816 ( .A(n13979), .B(P1_DATAO_REG_26__SCAN_IN), .S(n13773), .Z(
        P1_U3586) );
  MUX2_X1 U15817 ( .A(n13907), .B(P1_DATAO_REG_25__SCAN_IN), .S(n13773), .Z(
        P1_U3585) );
  MUX2_X1 U15818 ( .A(n13980), .B(P1_DATAO_REG_24__SCAN_IN), .S(n13773), .Z(
        P1_U3584) );
  MUX2_X1 U15819 ( .A(n14026), .B(P1_DATAO_REG_23__SCAN_IN), .S(n13773), .Z(
        P1_U3583) );
  MUX2_X1 U15820 ( .A(n13900), .B(P1_DATAO_REG_22__SCAN_IN), .S(n13773), .Z(
        P1_U3582) );
  MUX2_X1 U15821 ( .A(n14025), .B(P1_DATAO_REG_21__SCAN_IN), .S(n13773), .Z(
        P1_U3581) );
  MUX2_X1 U15822 ( .A(n13872), .B(P1_DATAO_REG_20__SCAN_IN), .S(n13773), .Z(
        P1_U3580) );
  INV_X1 U15823 ( .A(n14210), .ZN(n13895) );
  MUX2_X1 U15824 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n13895), .S(P1_U4016), .Z(
        P1_U3579) );
  MUX2_X1 U15825 ( .A(n14109), .B(P1_DATAO_REG_18__SCAN_IN), .S(n13773), .Z(
        P1_U3578) );
  MUX2_X1 U15826 ( .A(n14088), .B(P1_DATAO_REG_17__SCAN_IN), .S(n13773), .Z(
        P1_U3577) );
  MUX2_X1 U15827 ( .A(n14106), .B(P1_DATAO_REG_16__SCAN_IN), .S(n13773), .Z(
        P1_U3576) );
  MUX2_X1 U15828 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n13759), .S(P1_U4016), .Z(
        P1_U3575) );
  MUX2_X1 U15829 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n13760), .S(P1_U4016), .Z(
        P1_U3574) );
  MUX2_X1 U15830 ( .A(n13761), .B(P1_DATAO_REG_13__SCAN_IN), .S(n13773), .Z(
        P1_U3573) );
  MUX2_X1 U15831 ( .A(n13762), .B(P1_DATAO_REG_12__SCAN_IN), .S(n13773), .Z(
        P1_U3572) );
  MUX2_X1 U15832 ( .A(n13763), .B(P1_DATAO_REG_11__SCAN_IN), .S(n13773), .Z(
        P1_U3571) );
  MUX2_X1 U15833 ( .A(n13764), .B(P1_DATAO_REG_10__SCAN_IN), .S(n13773), .Z(
        P1_U3570) );
  MUX2_X1 U15834 ( .A(n13765), .B(P1_DATAO_REG_9__SCAN_IN), .S(n13773), .Z(
        P1_U3569) );
  MUX2_X1 U15835 ( .A(n13766), .B(P1_DATAO_REG_8__SCAN_IN), .S(n13773), .Z(
        P1_U3568) );
  MUX2_X1 U15836 ( .A(n13767), .B(P1_DATAO_REG_7__SCAN_IN), .S(n13773), .Z(
        P1_U3567) );
  MUX2_X1 U15837 ( .A(n13768), .B(P1_DATAO_REG_6__SCAN_IN), .S(n13773), .Z(
        P1_U3566) );
  MUX2_X1 U15838 ( .A(n13769), .B(P1_DATAO_REG_5__SCAN_IN), .S(n13773), .Z(
        P1_U3565) );
  MUX2_X1 U15839 ( .A(n8944), .B(P1_DATAO_REG_4__SCAN_IN), .S(n13773), .Z(
        P1_U3564) );
  MUX2_X1 U15840 ( .A(n13771), .B(P1_DATAO_REG_3__SCAN_IN), .S(n13773), .Z(
        P1_U3563) );
  MUX2_X1 U15841 ( .A(n13772), .B(P1_DATAO_REG_2__SCAN_IN), .S(n13773), .Z(
        P1_U3562) );
  MUX2_X1 U15842 ( .A(n14556), .B(P1_DATAO_REG_1__SCAN_IN), .S(n13773), .Z(
        P1_U3561) );
  MUX2_X1 U15843 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(n8344), .S(P1_U4016), .Z(
        P1_U3560) );
  INV_X1 U15844 ( .A(n13774), .ZN(n13777) );
  OAI211_X1 U15845 ( .C1(n13777), .C2(n13776), .A(n14478), .B(n13775), .ZN(
        n13786) );
  AOI22_X1 U15846 ( .A1(n14472), .A2(P1_ADDR_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(P1_U3086), .ZN(n13785) );
  INV_X1 U15847 ( .A(n13778), .ZN(n13779) );
  NAND2_X1 U15848 ( .A1(n14476), .A2(n13779), .ZN(n13784) );
  OAI211_X1 U15849 ( .C1(n13782), .C2(n13781), .A(n14483), .B(n13780), .ZN(
        n13783) );
  NAND4_X1 U15850 ( .A1(n13786), .A2(n13785), .A3(n13784), .A4(n13783), .ZN(
        P1_U3244) );
  AOI22_X1 U15851 ( .A1(n14472), .A2(P1_ADDR_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(P1_U3086), .ZN(n13800) );
  INV_X1 U15852 ( .A(n13787), .ZN(n13790) );
  MUX2_X1 U15853 ( .A(n8371), .B(P1_REG1_REG_2__SCAN_IN), .S(n13797), .Z(
        n13789) );
  INV_X1 U15854 ( .A(n13811), .ZN(n13788) );
  AOI211_X1 U15855 ( .C1(n13790), .C2(n13789), .A(n13788), .B(n14459), .ZN(
        n13796) );
  INV_X1 U15856 ( .A(n13791), .ZN(n13794) );
  MUX2_X1 U15857 ( .A(n15232), .B(P1_REG2_REG_2__SCAN_IN), .S(n13797), .Z(
        n13793) );
  INV_X1 U15858 ( .A(n13805), .ZN(n13792) );
  AOI211_X1 U15859 ( .C1(n13794), .C2(n13793), .A(n13792), .B(n14464), .ZN(
        n13795) );
  NOR2_X1 U15860 ( .A1(n13796), .A2(n13795), .ZN(n13799) );
  NAND2_X1 U15861 ( .A1(n14476), .A2(n13797), .ZN(n13798) );
  NAND4_X1 U15862 ( .A1(n13801), .A2(n13800), .A3(n13799), .A4(n13798), .ZN(
        P1_U3245) );
  INV_X1 U15863 ( .A(n13802), .ZN(n13807) );
  NAND3_X1 U15864 ( .A1(n13805), .A2(n13804), .A3(n13803), .ZN(n13806) );
  NAND3_X1 U15865 ( .A1(n14478), .A2(n13807), .A3(n13806), .ZN(n13817) );
  AOI22_X1 U15866 ( .A1(n14472), .A2(P1_ADDR_REG_3__SCAN_IN), .B1(
        P1_REG3_REG_3__SCAN_IN), .B2(P1_U3086), .ZN(n13816) );
  NAND2_X1 U15867 ( .A1(n14476), .A2(n13808), .ZN(n13815) );
  MUX2_X1 U15868 ( .A(n8385), .B(P1_REG1_REG_3__SCAN_IN), .S(n13808), .Z(
        n13809) );
  NAND3_X1 U15869 ( .A1(n13811), .A2(n13810), .A3(n13809), .ZN(n13812) );
  NAND3_X1 U15870 ( .A1(n14483), .A2(n13813), .A3(n13812), .ZN(n13814) );
  NAND4_X1 U15871 ( .A1(n13817), .A2(n13816), .A3(n13815), .A4(n13814), .ZN(
        P1_U3246) );
  INV_X1 U15872 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n13819) );
  OAI21_X1 U15873 ( .B1(n13819), .B2(n13821), .A(n13818), .ZN(n13838) );
  XNOR2_X1 U15874 ( .A(n13838), .B(n13831), .ZN(n13820) );
  NAND2_X1 U15875 ( .A1(P1_REG2_REG_18__SCAN_IN), .A2(n13820), .ZN(n13841) );
  OAI211_X1 U15876 ( .C1(n13820), .C2(P1_REG2_REG_18__SCAN_IN), .A(n14478), 
        .B(n13841), .ZN(n13830) );
  INV_X1 U15877 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n13822) );
  XNOR2_X1 U15878 ( .A(n13831), .B(n13833), .ZN(n13825) );
  NAND2_X1 U15879 ( .A1(P1_REG1_REG_18__SCAN_IN), .A2(n13825), .ZN(n13835) );
  OAI211_X1 U15880 ( .C1(P1_REG1_REG_18__SCAN_IN), .C2(n13825), .A(n14483), 
        .B(n13835), .ZN(n13826) );
  NAND2_X1 U15881 ( .A1(n13827), .A2(n13826), .ZN(n13828) );
  AOI21_X1 U15882 ( .B1(n14472), .B2(P1_ADDR_REG_18__SCAN_IN), .A(n13828), 
        .ZN(n13829) );
  OAI211_X1 U15883 ( .C1(n13832), .C2(n13831), .A(n13830), .B(n13829), .ZN(
        P1_U3261) );
  NAND2_X1 U15884 ( .A1(n13839), .A2(n13833), .ZN(n13834) );
  NAND2_X1 U15885 ( .A1(n13835), .A2(n13834), .ZN(n13837) );
  INV_X1 U15886 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n13836) );
  XNOR2_X1 U15887 ( .A(n13837), .B(n13836), .ZN(n13846) );
  INV_X1 U15888 ( .A(n13846), .ZN(n13844) );
  NAND2_X1 U15889 ( .A1(n13839), .A2(n13838), .ZN(n13840) );
  NAND2_X1 U15890 ( .A1(n13841), .A2(n13840), .ZN(n13842) );
  XOR2_X1 U15891 ( .A(P1_REG2_REG_19__SCAN_IN), .B(n13842), .Z(n13845) );
  NOR2_X1 U15892 ( .A1(n13845), .A2(n14464), .ZN(n13843) );
  AOI211_X1 U15893 ( .C1(n14483), .C2(n13844), .A(n14476), .B(n13843), .ZN(
        n13849) );
  AOI22_X1 U15894 ( .A1(n13846), .A2(n14483), .B1(n14478), .B2(n13845), .ZN(
        n13848) );
  MUX2_X1 U15895 ( .A(n13849), .B(n13848), .S(n13847), .Z(n13851) );
  OAI211_X1 U15896 ( .C1(n13852), .C2(n14469), .A(n13851), .B(n13850), .ZN(
        P1_U3262) );
  INV_X1 U15897 ( .A(n14136), .ZN(n13917) );
  OR2_X2 U15898 ( .A1(n13984), .A2(n14162), .ZN(n13968) );
  OR2_X2 U15899 ( .A1(n13956), .A2(n13968), .ZN(n13952) );
  NOR2_X2 U15900 ( .A1(n14143), .A2(n13952), .ZN(n13930) );
  NAND2_X1 U15901 ( .A1(n13917), .A2(n13930), .ZN(n13916) );
  NAND2_X1 U15902 ( .A1(n14127), .A2(n14099), .ZN(n13857) );
  INV_X1 U15903 ( .A(P1_B_REG_SCAN_IN), .ZN(n13853) );
  NOR2_X1 U15904 ( .A1(n14264), .A2(n13853), .ZN(n13854) );
  NOR2_X1 U15905 ( .A1(n14581), .A2(n13854), .ZN(n13918) );
  NAND2_X1 U15906 ( .A1(n13855), .A2(n13918), .ZN(n14132) );
  NOR2_X1 U15907 ( .A1(n6531), .A2(n14132), .ZN(n13859) );
  AOI21_X1 U15908 ( .B1(n6531), .B2(P1_REG2_REG_31__SCAN_IN), .A(n13859), .ZN(
        n13856) );
  OAI211_X1 U15909 ( .C1(n14128), .C2(n14119), .A(n13857), .B(n13856), .ZN(
        P1_U3263) );
  XNOR2_X1 U15910 ( .A(n14134), .B(n13916), .ZN(n13858) );
  NAND2_X1 U15911 ( .A1(n13858), .A2(n14546), .ZN(n14133) );
  NAND2_X1 U15912 ( .A1(n6531), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n13861) );
  INV_X1 U15913 ( .A(n13859), .ZN(n13860) );
  OAI211_X1 U15914 ( .C1(n14134), .C2(n14119), .A(n13861), .B(n13860), .ZN(
        n13862) );
  INV_X1 U15915 ( .A(n13862), .ZN(n13863) );
  OAI21_X1 U15916 ( .B1(n14133), .B2(n13959), .A(n13863), .ZN(P1_U3264) );
  INV_X1 U15917 ( .A(n13910), .ZN(n13885) );
  NAND2_X1 U15918 ( .A1(n14104), .A2(n13867), .ZN(n14087) );
  NOR2_X1 U15919 ( .A1(n14096), .A2(n14073), .ZN(n13868) );
  NAND2_X1 U15920 ( .A1(n14054), .A2(n13871), .ZN(n14053) );
  NAND2_X1 U15921 ( .A1(n14061), .A2(n13872), .ZN(n13873) );
  OR2_X1 U15922 ( .A1(n14190), .A2(n13874), .ZN(n13875) );
  NAND2_X1 U15923 ( .A1(n14186), .A2(n13876), .ZN(n13877) );
  INV_X1 U15924 ( .A(n13903), .ZN(n14020) );
  NAND2_X1 U15925 ( .A1(n14181), .A2(n13879), .ZN(n13880) );
  INV_X1 U15926 ( .A(n13907), .ZN(n13882) );
  NAND2_X1 U15927 ( .A1(n14168), .A2(n13882), .ZN(n13883) );
  INV_X1 U15928 ( .A(n13948), .ZN(n13884) );
  INV_X1 U15929 ( .A(n14143), .ZN(n13934) );
  XNOR2_X1 U15930 ( .A(n13887), .B(n13913), .ZN(n14140) );
  NAND2_X1 U15931 ( .A1(n13890), .A2(n14106), .ZN(n13888) );
  NAND2_X1 U15932 ( .A1(n13889), .A2(n13888), .ZN(n13892) );
  OR2_X1 U15933 ( .A1(n13890), .A2(n14106), .ZN(n13891) );
  NAND2_X1 U15934 ( .A1(n14096), .A2(n14109), .ZN(n13894) );
  INV_X1 U15935 ( .A(n14096), .ZN(n14211) );
  OR2_X1 U15936 ( .A1(n14203), .A2(n13895), .ZN(n13896) );
  INV_X1 U15937 ( .A(n13896), .ZN(n13897) );
  OR2_X1 U15938 ( .A1(n14061), .A2(n14074), .ZN(n13898) );
  OR2_X1 U15939 ( .A1(n14186), .A2(n13900), .ZN(n13901) );
  NAND2_X1 U15940 ( .A1(n13902), .A2(n13901), .ZN(n14019) );
  OR2_X1 U15941 ( .A1(n14181), .A2(n14026), .ZN(n13904) );
  OR2_X1 U15942 ( .A1(n14176), .A2(n13980), .ZN(n13905) );
  NAND2_X1 U15943 ( .A1(n14168), .A2(n13907), .ZN(n13908) );
  NAND2_X1 U15944 ( .A1(n14167), .A2(n13908), .ZN(n13964) );
  NAND2_X1 U15945 ( .A1(n14162), .A2(n13979), .ZN(n13909) );
  OR2_X1 U15946 ( .A1(n13956), .A2(n13910), .ZN(n13911) );
  NAND2_X1 U15947 ( .A1(n13938), .A2(n13912), .ZN(n13915) );
  XNOR2_X1 U15948 ( .A(n13915), .B(n13914), .ZN(n14135) );
  NAND2_X1 U15949 ( .A1(n13919), .A2(n13918), .ZN(n14137) );
  OAI22_X1 U15950 ( .A1(n13921), .A2(n14137), .B1(n13920), .B2(n14542), .ZN(
        n13924) );
  NAND2_X1 U15951 ( .A1(n13945), .A2(n14107), .ZN(n14138) );
  NAND2_X1 U15952 ( .A1(n6531), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n13922) );
  OAI21_X1 U15953 ( .B1(n6531), .B2(n14138), .A(n13922), .ZN(n13923) );
  AOI211_X1 U15954 ( .C1(n14136), .C2(n14566), .A(n13924), .B(n13923), .ZN(
        n13925) );
  OAI21_X1 U15955 ( .B1(n14139), .B2(n13959), .A(n13925), .ZN(n13926) );
  AOI21_X1 U15956 ( .B1(n14135), .B2(n14083), .A(n13926), .ZN(n13927) );
  OAI21_X1 U15957 ( .B1(n14140), .B2(n14085), .A(n13927), .ZN(P1_U3356) );
  AOI211_X1 U15958 ( .C1(n14143), .C2(n13952), .A(n14572), .B(n13930), .ZN(
        n14142) );
  INV_X1 U15959 ( .A(n13931), .ZN(n13932) );
  AOI22_X1 U15960 ( .A1(n6531), .A2(P1_REG2_REG_28__SCAN_IN), .B1(n13932), 
        .B2(n14567), .ZN(n13933) );
  OAI21_X1 U15961 ( .B1(n13934), .B2(n14119), .A(n13933), .ZN(n13935) );
  AOI21_X1 U15962 ( .B1(n14142), .B2(n14574), .A(n13935), .ZN(n13940) );
  NAND2_X1 U15963 ( .A1(n13937), .A2(n13936), .ZN(n14141) );
  NAND3_X1 U15964 ( .A1(n13938), .A2(n14083), .A3(n14141), .ZN(n13939) );
  OAI211_X1 U15965 ( .C1(n14149), .C2(n6531), .A(n13940), .B(n13939), .ZN(
        P1_U3265) );
  NOR2_X1 U15966 ( .A1(n13948), .A2(n7294), .ZN(n13942) );
  AND2_X1 U15967 ( .A1(n13965), .A2(n13942), .ZN(n13943) );
  OAI21_X1 U15968 ( .B1(n13944), .B2(n13943), .A(n14497), .ZN(n13947) );
  AOI22_X1 U15969 ( .A1(n14107), .A2(n13979), .B1(n13945), .B2(n14108), .ZN(
        n13946) );
  AND2_X2 U15970 ( .A1(n13947), .A2(n13946), .ZN(n14155) );
  NAND2_X1 U15971 ( .A1(n13949), .A2(n13948), .ZN(n13950) );
  NAND2_X1 U15972 ( .A1(n13951), .A2(n13950), .ZN(n14153) );
  AOI21_X1 U15973 ( .B1(n13956), .B2(n13968), .A(n14572), .ZN(n13953) );
  NAND2_X1 U15974 ( .A1(n13953), .A2(n13952), .ZN(n14150) );
  INV_X1 U15975 ( .A(n13954), .ZN(n13955) );
  AOI22_X1 U15976 ( .A1(n6531), .A2(P1_REG2_REG_27__SCAN_IN), .B1(n13955), 
        .B2(n14567), .ZN(n13958) );
  NAND2_X1 U15977 ( .A1(n13956), .A2(n14566), .ZN(n13957) );
  OAI211_X1 U15978 ( .C1(n14150), .C2(n13959), .A(n13958), .B(n13957), .ZN(
        n13960) );
  AOI21_X1 U15979 ( .B1(n14153), .B2(n14083), .A(n13960), .ZN(n13961) );
  OAI21_X1 U15980 ( .B1(n14155), .B2(n6531), .A(n13961), .ZN(P1_U3266) );
  OAI21_X1 U15981 ( .B1(n13964), .B2(n13963), .A(n13962), .ZN(n14165) );
  OAI21_X1 U15982 ( .B1(n13966), .B2(n6740), .A(n13965), .ZN(n14158) );
  NAND2_X1 U15983 ( .A1(n14158), .A2(n13967), .ZN(n13975) );
  AOI21_X1 U15984 ( .B1(n13984), .B2(n14162), .A(n14572), .ZN(n13969) );
  AND2_X1 U15985 ( .A1(n13969), .A2(n13968), .ZN(n14160) );
  NAND2_X1 U15986 ( .A1(n14162), .A2(n14566), .ZN(n13972) );
  AOI22_X1 U15987 ( .A1(n6531), .A2(P1_REG2_REG_26__SCAN_IN), .B1(n13970), 
        .B2(n14567), .ZN(n13971) );
  OAI211_X1 U15988 ( .C1(n6531), .C2(n14159), .A(n13972), .B(n13971), .ZN(
        n13973) );
  AOI21_X1 U15989 ( .B1(n14160), .B2(n14574), .A(n13973), .ZN(n13974) );
  OAI211_X1 U15990 ( .C1(n14165), .C2(n14123), .A(n13975), .B(n13974), .ZN(
        P1_U3267) );
  OAI21_X1 U15991 ( .B1(n13977), .B2(n13989), .A(n13976), .ZN(n13978) );
  NAND2_X1 U15992 ( .A1(n13978), .A2(n14497), .ZN(n13982) );
  AOI22_X1 U15993 ( .A1(n14107), .A2(n13980), .B1(n13979), .B2(n14108), .ZN(
        n13981) );
  NAND2_X1 U15994 ( .A1(n13982), .A2(n13981), .ZN(n14173) );
  INV_X1 U15995 ( .A(n14173), .ZN(n13993) );
  OR2_X1 U15996 ( .A1(n13987), .A2(n6591), .ZN(n13983) );
  AND2_X1 U15997 ( .A1(n13984), .A2(n13983), .ZN(n14169) );
  AOI22_X1 U15998 ( .A1(n6531), .A2(P1_REG2_REG_25__SCAN_IN), .B1(n13985), 
        .B2(n14567), .ZN(n13986) );
  OAI21_X1 U15999 ( .B1(n13987), .B2(n14119), .A(n13986), .ZN(n13988) );
  AOI21_X1 U16000 ( .B1(n14169), .B2(n14099), .A(n13988), .ZN(n13992) );
  NAND2_X1 U16001 ( .A1(n13990), .A2(n13989), .ZN(n14166) );
  NAND3_X1 U16002 ( .A1(n14167), .A2(n14166), .A3(n14083), .ZN(n13991) );
  OAI211_X1 U16003 ( .C1(n13993), .C2(n6531), .A(n13992), .B(n13991), .ZN(
        P1_U3268) );
  XNOR2_X1 U16004 ( .A(n13994), .B(n13998), .ZN(n14003) );
  INV_X1 U16005 ( .A(n14493), .ZN(n14596) );
  INV_X1 U16006 ( .A(n13995), .ZN(n14000) );
  AOI211_X1 U16007 ( .C1(n13998), .C2(n13997), .A(n14560), .B(n13996), .ZN(
        n13999) );
  AOI211_X1 U16008 ( .C1(n14176), .C2(n14013), .A(n14572), .B(n6591), .ZN(
        n14175) );
  AOI22_X1 U16009 ( .A1(n6531), .A2(P1_REG2_REG_24__SCAN_IN), .B1(n14001), 
        .B2(n14567), .ZN(n14002) );
  OAI21_X1 U16010 ( .B1(n6982), .B2(n14119), .A(n14002), .ZN(n14007) );
  INV_X1 U16011 ( .A(n14003), .ZN(n14179) );
  INV_X1 U16012 ( .A(n14004), .ZN(n14005) );
  NAND2_X1 U16013 ( .A1(n14543), .A2(n14005), .ZN(n14502) );
  NOR2_X1 U16014 ( .A1(n14179), .A2(n14502), .ZN(n14006) );
  AOI211_X1 U16015 ( .C1(n14175), .C2(n14574), .A(n14007), .B(n14006), .ZN(
        n14008) );
  OAI21_X1 U16016 ( .B1(n14178), .B2(n6531), .A(n14008), .ZN(P1_U3269) );
  OAI21_X1 U16017 ( .B1(n14010), .B2(n14020), .A(n14009), .ZN(n14012) );
  AOI21_X1 U16018 ( .B1(n14012), .B2(n14497), .A(n14011), .ZN(n14183) );
  INV_X1 U16019 ( .A(n14013), .ZN(n14014) );
  AOI211_X1 U16020 ( .C1(n14181), .C2(n14028), .A(n14572), .B(n14014), .ZN(
        n14180) );
  INV_X1 U16021 ( .A(n14015), .ZN(n14016) );
  AOI22_X1 U16022 ( .A1(n6531), .A2(P1_REG2_REG_23__SCAN_IN), .B1(n14016), 
        .B2(n14567), .ZN(n14017) );
  OAI21_X1 U16023 ( .B1(n14018), .B2(n14119), .A(n14017), .ZN(n14022) );
  XNOR2_X1 U16024 ( .A(n14019), .B(n14020), .ZN(n14184) );
  NOR2_X1 U16025 ( .A1(n14184), .A2(n14123), .ZN(n14021) );
  AOI211_X1 U16026 ( .C1(n14180), .C2(n14574), .A(n14022), .B(n14021), .ZN(
        n14023) );
  OAI21_X1 U16027 ( .B1(n6531), .B2(n14183), .A(n14023), .ZN(P1_U3270) );
  XNOR2_X1 U16028 ( .A(n14024), .B(n14034), .ZN(n14027) );
  AOI222_X1 U16029 ( .A1(n14497), .A2(n14027), .B1(n14026), .B2(n14108), .C1(
        n14025), .C2(n14107), .ZN(n14188) );
  INV_X1 U16030 ( .A(n14042), .ZN(n14030) );
  INV_X1 U16031 ( .A(n14028), .ZN(n14029) );
  AOI211_X1 U16032 ( .C1(n14186), .C2(n14030), .A(n14572), .B(n14029), .ZN(
        n14185) );
  AOI22_X1 U16033 ( .A1(n14031), .A2(n14567), .B1(P1_REG2_REG_22__SCAN_IN), 
        .B2(n6531), .ZN(n14032) );
  OAI21_X1 U16034 ( .B1(n14033), .B2(n14119), .A(n14032), .ZN(n14037) );
  XOR2_X1 U16035 ( .A(n14035), .B(n14034), .Z(n14189) );
  NOR2_X1 U16036 ( .A1(n14189), .A2(n14123), .ZN(n14036) );
  AOI211_X1 U16037 ( .C1(n14185), .C2(n14574), .A(n14037), .B(n14036), .ZN(
        n14038) );
  OAI21_X1 U16038 ( .B1(n6531), .B2(n14188), .A(n14038), .ZN(P1_U3271) );
  XOR2_X1 U16039 ( .A(n14039), .B(n14049), .Z(n14041) );
  AOI21_X1 U16040 ( .B1(n14041), .B2(n14497), .A(n14040), .ZN(n14193) );
  AOI21_X1 U16041 ( .B1(n14190), .B2(n14055), .A(n14042), .ZN(n14191) );
  AOI22_X1 U16042 ( .A1(n14043), .A2(n14567), .B1(n6531), .B2(
        P1_REG2_REG_21__SCAN_IN), .ZN(n14044) );
  OAI21_X1 U16043 ( .B1(n14045), .B2(n14119), .A(n14044), .ZN(n14051) );
  INV_X1 U16044 ( .A(n14046), .ZN(n14047) );
  AOI21_X1 U16045 ( .B1(n14049), .B2(n14048), .A(n14047), .ZN(n14194) );
  NOR2_X1 U16046 ( .A1(n14194), .A2(n14123), .ZN(n14050) );
  AOI211_X1 U16047 ( .C1(n14191), .C2(n14099), .A(n14051), .B(n14050), .ZN(
        n14052) );
  OAI21_X1 U16048 ( .B1(n6531), .B2(n14193), .A(n14052), .ZN(P1_U3272) );
  OAI21_X1 U16049 ( .B1(n14054), .B2(n13871), .A(n14053), .ZN(n14201) );
  AOI21_X1 U16050 ( .B1(n14077), .B2(n14197), .A(n14572), .ZN(n14056) );
  AND2_X1 U16051 ( .A1(n14056), .A2(n14055), .ZN(n14195) );
  INV_X1 U16052 ( .A(n14057), .ZN(n14058) );
  AOI22_X1 U16053 ( .A1(P1_REG2_REG_20__SCAN_IN), .A2(n6531), .B1(n14058), 
        .B2(n14567), .ZN(n14060) );
  NAND2_X1 U16054 ( .A1(n14196), .A2(n14543), .ZN(n14059) );
  OAI211_X1 U16055 ( .C1(n14061), .C2(n14119), .A(n14060), .B(n14059), .ZN(
        n14062) );
  AOI21_X1 U16056 ( .B1(n14195), .B2(n14574), .A(n14062), .ZN(n14067) );
  OR2_X1 U16057 ( .A1(n14064), .A2(n14063), .ZN(n14198) );
  NAND3_X1 U16058 ( .A1(n14198), .A2(n14083), .A3(n14065), .ZN(n14066) );
  OAI211_X1 U16059 ( .C1(n14201), .C2(n14085), .A(n14067), .B(n14066), .ZN(
        P1_U3273) );
  XNOR2_X1 U16060 ( .A(n14069), .B(n14068), .ZN(n14209) );
  XNOR2_X1 U16061 ( .A(n14071), .B(n14070), .ZN(n14207) );
  AOI22_X1 U16062 ( .A1(n6531), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n14072), 
        .B2(n14567), .ZN(n14076) );
  OAI22_X1 U16063 ( .A1(n14074), .A2(n14581), .B1(n14073), .B2(n14561), .ZN(
        n14202) );
  NAND2_X1 U16064 ( .A1(n14202), .A2(n14543), .ZN(n14075) );
  OAI211_X1 U16065 ( .C1(n14079), .C2(n14119), .A(n14076), .B(n14075), .ZN(
        n14082) );
  INV_X1 U16066 ( .A(n14098), .ZN(n14078) );
  OAI21_X1 U16067 ( .B1(n14079), .B2(n14078), .A(n14077), .ZN(n14205) );
  NOR2_X1 U16068 ( .A1(n14205), .A2(n14080), .ZN(n14081) );
  AOI211_X1 U16069 ( .C1(n14083), .C2(n14207), .A(n14082), .B(n14081), .ZN(
        n14084) );
  OAI21_X1 U16070 ( .B1(n14209), .B2(n14085), .A(n14084), .ZN(P1_U3274) );
  XNOR2_X1 U16071 ( .A(n14087), .B(n14086), .ZN(n14089) );
  AOI22_X1 U16072 ( .A1(n14089), .A2(n14497), .B1(n14107), .B2(n14088), .ZN(
        n14215) );
  XNOR2_X1 U16073 ( .A(n14091), .B(n14090), .ZN(n14216) );
  NOR2_X1 U16074 ( .A1(n14542), .A2(n14092), .ZN(n14093) );
  AOI21_X1 U16075 ( .B1(n6531), .B2(P1_REG2_REG_18__SCAN_IN), .A(n14093), .ZN(
        n14094) );
  OAI21_X1 U16076 ( .B1(n14570), .B2(n14210), .A(n14094), .ZN(n14095) );
  AOI21_X1 U16077 ( .B1(n14096), .B2(n14566), .A(n14095), .ZN(n14101) );
  NAND2_X1 U16078 ( .A1(n14096), .A2(n14113), .ZN(n14097) );
  AND2_X1 U16079 ( .A1(n14098), .A2(n14097), .ZN(n14213) );
  NAND2_X1 U16080 ( .A1(n14213), .A2(n14099), .ZN(n14100) );
  OAI211_X1 U16081 ( .C1(n14216), .C2(n14123), .A(n14101), .B(n14100), .ZN(
        n14102) );
  INV_X1 U16082 ( .A(n14102), .ZN(n14103) );
  OAI21_X1 U16083 ( .B1(n14215), .B2(n6531), .A(n14103), .ZN(P1_U3275) );
  OAI211_X1 U16084 ( .C1(n14105), .C2(n14121), .A(n14104), .B(n14497), .ZN(
        n14111) );
  AOI22_X1 U16085 ( .A1(n14109), .A2(n14108), .B1(n14107), .B2(n14106), .ZN(
        n14110) );
  AND2_X1 U16086 ( .A1(n14111), .A2(n14110), .ZN(n14219) );
  INV_X1 U16087 ( .A(n14112), .ZN(n14115) );
  INV_X1 U16088 ( .A(n14113), .ZN(n14114) );
  AOI211_X1 U16089 ( .C1(n14218), .C2(n14115), .A(n14572), .B(n14114), .ZN(
        n14217) );
  INV_X1 U16090 ( .A(n14116), .ZN(n14117) );
  AOI22_X1 U16091 ( .A1(n6531), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n14117), 
        .B2(n14567), .ZN(n14118) );
  OAI21_X1 U16092 ( .B1(n14120), .B2(n14119), .A(n14118), .ZN(n14125) );
  XNOR2_X1 U16093 ( .A(n14122), .B(n14121), .ZN(n14221) );
  NOR2_X1 U16094 ( .A1(n14221), .A2(n14123), .ZN(n14124) );
  AOI211_X1 U16095 ( .C1(n14217), .C2(n14574), .A(n14125), .B(n14124), .ZN(
        n14126) );
  OAI21_X1 U16096 ( .B1(n6531), .B2(n14219), .A(n14126), .ZN(P1_U3276) );
  OAI21_X1 U16097 ( .B1(n14128), .B2(n14638), .A(n14132), .ZN(n14129) );
  INV_X1 U16098 ( .A(n14129), .ZN(n14130) );
  NAND2_X1 U16099 ( .A1(n14131), .A2(n14130), .ZN(n14235) );
  MUX2_X1 U16100 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n14235), .S(n14658), .Z(
        P1_U3559) );
  OAI211_X1 U16101 ( .C1(n14134), .C2(n14638), .A(n14133), .B(n14132), .ZN(
        n14236) );
  MUX2_X1 U16102 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n14236), .S(n14658), .Z(
        P1_U3558) );
  MUX2_X1 U16103 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n14237), .S(n14658), .Z(
        P1_U3557) );
  NAND2_X1 U16104 ( .A1(n14141), .A2(n14641), .ZN(n14145) );
  AOI21_X1 U16105 ( .B1(n14143), .B2(n14607), .A(n14142), .ZN(n14144) );
  OAI21_X1 U16106 ( .B1(n14146), .B2(n14145), .A(n14144), .ZN(n14147) );
  NAND2_X1 U16107 ( .A1(n14149), .A2(n14148), .ZN(n14238) );
  MUX2_X1 U16108 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n14238), .S(n14658), .Z(
        P1_U3556) );
  INV_X1 U16109 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n14156) );
  OAI21_X1 U16110 ( .B1(n14151), .B2(n14638), .A(n14150), .ZN(n14152) );
  AOI21_X1 U16111 ( .B1(n14153), .B2(n14641), .A(n14152), .ZN(n14154) );
  MUX2_X1 U16112 ( .A(n14156), .B(n14239), .S(n14658), .Z(n14157) );
  INV_X1 U16113 ( .A(n14157), .ZN(P1_U3555) );
  NAND2_X1 U16114 ( .A1(n14158), .A2(n14497), .ZN(n14164) );
  INV_X1 U16115 ( .A(n14159), .ZN(n14161) );
  AOI211_X1 U16116 ( .C1(n14162), .C2(n14607), .A(n14161), .B(n14160), .ZN(
        n14163) );
  OAI211_X1 U16117 ( .C1(n14611), .C2(n14165), .A(n14164), .B(n14163), .ZN(
        n14241) );
  MUX2_X1 U16118 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n14241), .S(n14658), .Z(
        P1_U3554) );
  NAND3_X1 U16119 ( .A1(n14167), .A2(n14166), .A3(n14641), .ZN(n14171) );
  AOI22_X1 U16120 ( .A1(n14169), .A2(n14546), .B1(n14168), .B2(n14607), .ZN(
        n14170) );
  NAND2_X1 U16121 ( .A1(n14171), .A2(n14170), .ZN(n14172) );
  NOR2_X1 U16122 ( .A1(n14173), .A2(n14172), .ZN(n14242) );
  MUX2_X1 U16123 ( .A(n15337), .B(n14242), .S(n14658), .Z(n14174) );
  INV_X1 U16124 ( .A(n14174), .ZN(P1_U3553) );
  AOI21_X1 U16125 ( .B1(n14176), .B2(n14607), .A(n14175), .ZN(n14177) );
  OAI211_X1 U16126 ( .C1(n14592), .C2(n14179), .A(n14178), .B(n14177), .ZN(
        n14245) );
  MUX2_X1 U16127 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n14245), .S(n14658), .Z(
        P1_U3552) );
  AOI21_X1 U16128 ( .B1(n14181), .B2(n14607), .A(n14180), .ZN(n14182) );
  OAI211_X1 U16129 ( .C1(n14611), .C2(n14184), .A(n14183), .B(n14182), .ZN(
        n14246) );
  MUX2_X1 U16130 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n14246), .S(n14658), .Z(
        P1_U3551) );
  AOI21_X1 U16131 ( .B1(n14186), .B2(n14607), .A(n14185), .ZN(n14187) );
  OAI211_X1 U16132 ( .C1(n14611), .C2(n14189), .A(n14188), .B(n14187), .ZN(
        n14247) );
  MUX2_X1 U16133 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n14247), .S(n14658), .Z(
        P1_U3550) );
  AOI22_X1 U16134 ( .A1(n14191), .A2(n14546), .B1(n14190), .B2(n14607), .ZN(
        n14192) );
  OAI211_X1 U16135 ( .C1(n14194), .C2(n14611), .A(n14193), .B(n14192), .ZN(
        n14248) );
  MUX2_X1 U16136 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n14248), .S(n14658), .Z(
        P1_U3549) );
  AOI211_X1 U16137 ( .C1(n14197), .C2(n14607), .A(n14196), .B(n14195), .ZN(
        n14200) );
  NAND3_X1 U16138 ( .A1(n14198), .A2(n14065), .A3(n14641), .ZN(n14199) );
  OAI211_X1 U16139 ( .C1(n14201), .C2(n14560), .A(n14200), .B(n14199), .ZN(
        n14249) );
  MUX2_X1 U16140 ( .A(n14249), .B(P1_REG1_REG_20__SCAN_IN), .S(n14655), .Z(
        P1_U3548) );
  AOI21_X1 U16141 ( .B1(n14203), .B2(n14607), .A(n14202), .ZN(n14204) );
  OAI21_X1 U16142 ( .B1(n14205), .B2(n14572), .A(n14204), .ZN(n14206) );
  AOI21_X1 U16143 ( .B1(n14207), .B2(n14641), .A(n14206), .ZN(n14208) );
  OAI21_X1 U16144 ( .B1(n14209), .B2(n14560), .A(n14208), .ZN(n14250) );
  MUX2_X1 U16145 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n14250), .S(n14658), .Z(
        P1_U3547) );
  OAI22_X1 U16146 ( .A1(n14211), .A2(n14638), .B1(n14210), .B2(n14581), .ZN(
        n14212) );
  AOI21_X1 U16147 ( .B1(n14546), .B2(n14213), .A(n14212), .ZN(n14214) );
  OAI211_X1 U16148 ( .C1(n14611), .C2(n14216), .A(n14215), .B(n14214), .ZN(
        n14251) );
  MUX2_X1 U16149 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n14251), .S(n14658), .Z(
        P1_U3546) );
  AOI21_X1 U16150 ( .B1(n14218), .B2(n14607), .A(n14217), .ZN(n14220) );
  OAI211_X1 U16151 ( .C1(n14611), .C2(n14221), .A(n14220), .B(n14219), .ZN(
        n14252) );
  MUX2_X1 U16152 ( .A(n14252), .B(P1_REG1_REG_17__SCAN_IN), .S(n14655), .Z(
        P1_U3545) );
  OAI21_X1 U16153 ( .B1(n14223), .B2(n14638), .A(n14222), .ZN(n14225) );
  AOI211_X1 U16154 ( .C1(n14226), .C2(n14641), .A(n14225), .B(n14224), .ZN(
        n14227) );
  OAI21_X1 U16155 ( .B1(n14560), .B2(n14228), .A(n14227), .ZN(n14253) );
  MUX2_X1 U16156 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n14253), .S(n14658), .Z(
        P1_U3544) );
  OAI21_X1 U16157 ( .B1(n6967), .B2(n14638), .A(n14229), .ZN(n14230) );
  AOI21_X1 U16158 ( .B1(n14231), .B2(n14641), .A(n14230), .ZN(n14232) );
  AND2_X1 U16159 ( .A1(n14233), .A2(n14232), .ZN(n14254) );
  MUX2_X1 U16160 ( .A(n15145), .B(n14254), .S(n14658), .Z(n14234) );
  INV_X1 U16161 ( .A(n14234), .ZN(P1_U3543) );
  MUX2_X1 U16162 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n14235), .S(n14645), .Z(
        P1_U3527) );
  MUX2_X1 U16163 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n14236), .S(n14645), .Z(
        P1_U3526) );
  MUX2_X1 U16164 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n14238), .S(n14645), .Z(
        P1_U3524) );
  MUX2_X1 U16165 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n14240), .S(n14645), .Z(
        P1_U3523) );
  MUX2_X1 U16166 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n14241), .S(n14645), .Z(
        P1_U3522) );
  INV_X1 U16167 ( .A(P1_REG0_REG_25__SCAN_IN), .ZN(n14243) );
  MUX2_X1 U16168 ( .A(n14243), .B(n14242), .S(n14645), .Z(n14244) );
  INV_X1 U16169 ( .A(n14244), .ZN(P1_U3521) );
  MUX2_X1 U16170 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n14245), .S(n14645), .Z(
        P1_U3520) );
  MUX2_X1 U16171 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n14246), .S(n14645), .Z(
        P1_U3519) );
  MUX2_X1 U16172 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n14247), .S(n14645), .Z(
        P1_U3518) );
  MUX2_X1 U16173 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n14248), .S(n14645), .Z(
        P1_U3517) );
  MUX2_X1 U16174 ( .A(n14249), .B(P1_REG0_REG_20__SCAN_IN), .S(n14643), .Z(
        P1_U3516) );
  MUX2_X1 U16175 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n14250), .S(n14645), .Z(
        P1_U3515) );
  MUX2_X1 U16176 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n14251), .S(n14645), .Z(
        P1_U3513) );
  MUX2_X1 U16177 ( .A(n14252), .B(P1_REG0_REG_17__SCAN_IN), .S(n14643), .Z(
        P1_U3510) );
  MUX2_X1 U16178 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n14253), .S(n14645), .Z(
        P1_U3507) );
  MUX2_X1 U16179 ( .A(n14255), .B(n14254), .S(n14645), .Z(n14256) );
  INV_X1 U16180 ( .A(n14256), .ZN(P1_U3504) );
  NOR4_X1 U16181 ( .A1(n14257), .A2(P1_IR_REG_30__SCAN_IN), .A3(P1_U3086), 
        .A4(n14258), .ZN(n14259) );
  AOI21_X1 U16182 ( .B1(P2_DATAO_REG_31__SCAN_IN), .B2(n14260), .A(n14259), 
        .ZN(n14261) );
  OAI21_X1 U16183 ( .B1(n14262), .B2(n6535), .A(n14261), .ZN(P1_U3324) );
  INV_X1 U16184 ( .A(n14265), .ZN(n14269) );
  OAI222_X1 U16185 ( .A1(n14269), .A2(P1_U3086), .B1(n6535), .B2(n14268), .C1(
        n14267), .C2(n14266), .ZN(P1_U3329) );
  MUX2_X1 U16186 ( .A(n14271), .B(n14270), .S(P1_U3086), .Z(P1_U3333) );
  INV_X1 U16187 ( .A(n14272), .ZN(n14273) );
  MUX2_X1 U16188 ( .A(n14273), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  INV_X1 U16189 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n15242) );
  XNOR2_X1 U16190 ( .A(n14275), .B(n15242), .ZN(SUB_1596_U62) );
  AOI21_X1 U16191 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(
        P3_WR_REG_SCAN_IN), .ZN(n14276) );
  OAI21_X1 U16192 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(n14276), 
        .ZN(U28) );
  AOI21_X1 U16193 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(
        P3_RD_REG_SCAN_IN), .ZN(n14277) );
  OAI21_X1 U16194 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(n14277), 
        .ZN(U29) );
  OAI222_X1 U16195 ( .A1(n14282), .A2(n14281), .B1(n14282), .B2(n14280), .C1(
        n14279), .C2(n14278), .ZN(SUB_1596_U61) );
  AOI21_X1 U16196 ( .B1(n14285), .B2(n14284), .A(n14283), .ZN(SUB_1596_U57) );
  OAI21_X1 U16197 ( .B1(n14288), .B2(n14287), .A(n14286), .ZN(n14289) );
  XNOR2_X1 U16198 ( .A(n14289), .B(P2_ADDR_REG_8__SCAN_IN), .ZN(SUB_1596_U55)
         );
  OAI222_X1 U16199 ( .A1(n14703), .A2(n14293), .B1(n14703), .B2(n14292), .C1(
        n14291), .C2(n14290), .ZN(SUB_1596_U54) );
  OAI222_X1 U16200 ( .A1(n14298), .A2(n14297), .B1(n14298), .B2(n14296), .C1(
        n14295), .C2(n14294), .ZN(SUB_1596_U70) );
  AOI21_X1 U16201 ( .B1(n14301), .B2(n14300), .A(n14299), .ZN(n14302) );
  XOR2_X1 U16202 ( .A(P2_ADDR_REG_17__SCAN_IN), .B(n14302), .Z(SUB_1596_U63)
         );
  XNOR2_X1 U16203 ( .A(n14303), .B(n14308), .ZN(n14305) );
  AOI222_X1 U16204 ( .A1(n15046), .A2(n14305), .B1(n14984), .B2(n15041), .C1(
        n14304), .C2(n15038), .ZN(n14325) );
  AOI22_X1 U16205 ( .A1(n15052), .A2(P3_REG2_REG_12__SCAN_IN), .B1(n15055), 
        .B2(n14306), .ZN(n14312) );
  XNOR2_X1 U16206 ( .A(n14307), .B(n14308), .ZN(n14328) );
  NOR2_X1 U16207 ( .A1(n14309), .A2(n15018), .ZN(n14327) );
  AOI22_X1 U16208 ( .A1(n14328), .A2(n14310), .B1(n14991), .B2(n14327), .ZN(
        n14311) );
  OAI211_X1 U16209 ( .C1(n15052), .C2(n14325), .A(n14312), .B(n14311), .ZN(
        P3_U3221) );
  INV_X1 U16210 ( .A(n15010), .ZN(n15033) );
  INV_X1 U16211 ( .A(n14313), .ZN(n14979) );
  OAI21_X1 U16212 ( .B1(n14979), .B2(n14314), .A(n14317), .ZN(n14316) );
  NAND2_X1 U16213 ( .A1(n14316), .A2(n14315), .ZN(n14331) );
  XNOR2_X1 U16214 ( .A(n14318), .B(n14317), .ZN(n14319) );
  OAI222_X1 U16215 ( .A1(n15029), .A2(n15393), .B1(n15031), .B2(n14320), .C1(
        n14319), .C2(n15027), .ZN(n14329) );
  AOI21_X1 U16216 ( .B1(n15033), .B2(n14331), .A(n14329), .ZN(n14324) );
  NOR2_X1 U16217 ( .A1(n14321), .A2(n15018), .ZN(n14330) );
  INV_X1 U16218 ( .A(n15394), .ZN(n14322) );
  AOI22_X1 U16219 ( .A1(n14991), .A2(n14330), .B1(n15055), .B2(n14322), .ZN(
        n14323) );
  OAI221_X1 U16220 ( .B1(n15052), .B2(n14324), .C1(n15057), .C2(n10584), .A(
        n14323), .ZN(P3_U3222) );
  INV_X1 U16221 ( .A(n14325), .ZN(n14326) );
  AOI211_X1 U16222 ( .C1(n14328), .C2(n15083), .A(n14327), .B(n14326), .ZN(
        n14332) );
  AOI22_X1 U16223 ( .A1(n15096), .A2(n14332), .B1(n11129), .B2(n15094), .ZN(
        P3_U3471) );
  AOI211_X1 U16224 ( .C1(n15083), .C2(n14331), .A(n14330), .B(n14329), .ZN(
        n14333) );
  AOI22_X1 U16225 ( .A1(n15096), .A2(n14333), .B1(n10582), .B2(n15094), .ZN(
        P3_U3470) );
  AOI22_X1 U16226 ( .A1(n15086), .A2(n11078), .B1(n14332), .B2(n15085), .ZN(
        P3_U3426) );
  AOI22_X1 U16227 ( .A1(n15086), .A2(n10585), .B1(n14333), .B2(n15085), .ZN(
        P3_U3423) );
  AOI22_X1 U16228 ( .A1(n14337), .A2(n14336), .B1(n14335), .B2(n14334), .ZN(
        n14350) );
  AOI21_X1 U16229 ( .B1(n14339), .B2(n14338), .A(n6683), .ZN(n14341) );
  OAI222_X1 U16230 ( .A1(n14343), .A2(n14350), .B1(n14342), .B2(n14341), .C1(
        n14340), .C2(n8167), .ZN(n14344) );
  INV_X1 U16231 ( .A(n14344), .ZN(n14346) );
  OAI211_X1 U16232 ( .C1(n14348), .C2(n14347), .A(n14346), .B(n14345), .ZN(
        P2_U3187) );
  XOR2_X1 U16233 ( .A(n14349), .B(n14358), .Z(n14352) );
  OAI21_X1 U16234 ( .B1(n14352), .B2(n14351), .A(n14350), .ZN(n14369) );
  INV_X1 U16235 ( .A(n14369), .ZN(n14366) );
  AOI222_X1 U16236 ( .A1(n14356), .A2(n14355), .B1(P2_REG2_REG_14__SCAN_IN), 
        .B2(n14367), .C1(n14354), .C2(n14353), .ZN(n14365) );
  XOR2_X1 U16237 ( .A(n14358), .B(n14357), .Z(n14371) );
  OAI211_X1 U16238 ( .C1(n8167), .C2(n10990), .A(n9550), .B(n14360), .ZN(
        n14368) );
  INV_X1 U16239 ( .A(n14368), .ZN(n14361) );
  AOI22_X1 U16240 ( .A1(n14371), .A2(n14363), .B1(n14362), .B2(n14361), .ZN(
        n14364) );
  OAI211_X1 U16241 ( .C1(n14367), .C2(n14366), .A(n14365), .B(n14364), .ZN(
        P2_U3251) );
  OAI21_X1 U16242 ( .B1(n8167), .B2(n14806), .A(n14368), .ZN(n14370) );
  AOI211_X1 U16243 ( .C1(n14378), .C2(n14371), .A(n14370), .B(n14369), .ZN(
        n14387) );
  AOI22_X1 U16244 ( .A1(n14829), .A2(n14387), .B1(n14372), .B2(n14827), .ZN(
        P2_U3513) );
  OAI21_X1 U16245 ( .B1(n14374), .B2(n14806), .A(n14373), .ZN(n14376) );
  AOI211_X1 U16246 ( .C1(n14378), .C2(n14377), .A(n14376), .B(n14375), .ZN(
        n14389) );
  AOI22_X1 U16247 ( .A1(n14829), .A2(n14389), .B1(n10153), .B2(n14827), .ZN(
        P2_U3512) );
  INV_X1 U16248 ( .A(n14803), .ZN(n14815) );
  NAND2_X1 U16249 ( .A1(n14379), .A2(n14810), .ZN(n14380) );
  NAND2_X1 U16250 ( .A1(n14381), .A2(n14380), .ZN(n14382) );
  AOI21_X1 U16251 ( .B1(n14383), .B2(n14815), .A(n14382), .ZN(n14384) );
  AOI22_X1 U16252 ( .A1(n14829), .A2(n14390), .B1(n14386), .B2(n14827), .ZN(
        P2_U3511) );
  AOI22_X1 U16253 ( .A1(n14821), .A2(n14387), .B1(n7829), .B2(n14819), .ZN(
        P2_U3472) );
  INV_X1 U16254 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n14388) );
  AOI22_X1 U16255 ( .A1(n14821), .A2(n14389), .B1(n14388), .B2(n14819), .ZN(
        P2_U3469) );
  AOI22_X1 U16256 ( .A1(n14821), .A2(n14390), .B1(n7797), .B2(n14819), .ZN(
        P2_U3466) );
  NAND2_X1 U16257 ( .A1(n14392), .A2(n14391), .ZN(n14393) );
  NAND2_X1 U16258 ( .A1(n14394), .A2(n14393), .ZN(n14396) );
  AOI222_X1 U16259 ( .A1(n14398), .A2(n14405), .B1(n14404), .B2(n14397), .C1(
        n14396), .C2(n14395), .ZN(n14400) );
  OAI211_X1 U16260 ( .C1(n14402), .C2(n14401), .A(n14400), .B(n14399), .ZN(
        P1_U3215) );
  AOI211_X1 U16261 ( .C1(n14405), .C2(n14607), .A(n14404), .B(n14403), .ZN(
        n14406) );
  OAI21_X1 U16262 ( .B1(n14611), .B2(n14407), .A(n14406), .ZN(n14408) );
  AOI21_X1 U16263 ( .B1(n14497), .B2(n14409), .A(n14408), .ZN(n14417) );
  AOI22_X1 U16264 ( .A1(n14658), .A2(n14417), .B1(n8554), .B2(n14655), .ZN(
        P1_U3542) );
  OAI21_X1 U16265 ( .B1(n14411), .B2(n14638), .A(n14410), .ZN(n14413) );
  AOI211_X1 U16266 ( .C1(n14414), .C2(n14641), .A(n14413), .B(n14412), .ZN(
        n14419) );
  AOI22_X1 U16267 ( .A1(n14658), .A2(n14419), .B1(n14415), .B2(n14655), .ZN(
        P1_U3539) );
  INV_X1 U16268 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n14416) );
  AOI22_X1 U16269 ( .A1(n14645), .A2(n14417), .B1(n14416), .B2(n14643), .ZN(
        P1_U3501) );
  INV_X1 U16270 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n14418) );
  AOI22_X1 U16271 ( .A1(n14645), .A2(n14419), .B1(n14418), .B2(n14643), .ZN(
        P1_U3492) );
  OAI21_X1 U16272 ( .B1(n14422), .B2(n14421), .A(n14420), .ZN(n14423) );
  XNOR2_X1 U16273 ( .A(n14423), .B(P2_ADDR_REG_11__SCAN_IN), .ZN(SUB_1596_U69)
         );
  OAI21_X1 U16274 ( .B1(n14425), .B2(n15365), .A(n14424), .ZN(SUB_1596_U68) );
  AOI21_X1 U16275 ( .B1(n14428), .B2(n14427), .A(n14426), .ZN(n14429) );
  XOR2_X1 U16276 ( .A(P2_ADDR_REG_13__SCAN_IN), .B(n14429), .Z(SUB_1596_U67)
         );
  OAI21_X1 U16277 ( .B1(n14432), .B2(n14431), .A(n14430), .ZN(n14433) );
  XNOR2_X1 U16278 ( .A(n14433), .B(P2_ADDR_REG_14__SCAN_IN), .ZN(SUB_1596_U66)
         );
  AOI21_X1 U16279 ( .B1(n14436), .B2(n14435), .A(n14434), .ZN(n14437) );
  XOR2_X1 U16280 ( .A(P2_ADDR_REG_15__SCAN_IN), .B(n14437), .Z(SUB_1596_U65)
         );
  AOI21_X1 U16281 ( .B1(n14440), .B2(n14439), .A(n14438), .ZN(n14441) );
  XOR2_X1 U16282 ( .A(P2_ADDR_REG_16__SCAN_IN), .B(n14441), .Z(SUB_1596_U64)
         );
  NOR2_X1 U16283 ( .A1(n14442), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n14444) );
  OR2_X1 U16284 ( .A1(n14443), .A2(n14444), .ZN(n14447) );
  INV_X1 U16285 ( .A(n14444), .ZN(n14446) );
  MUX2_X1 U16286 ( .A(n14447), .B(n14446), .S(n14445), .Z(n14449) );
  NAND2_X1 U16287 ( .A1(n14449), .A2(n14448), .ZN(n14451) );
  AOI22_X1 U16288 ( .A1(n14472), .A2(P1_ADDR_REG_0__SCAN_IN), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(P1_U3086), .ZN(n14450) );
  OAI21_X1 U16289 ( .B1(n14452), .B2(n14451), .A(n14450), .ZN(P1_U3243) );
  AOI21_X1 U16290 ( .B1(n14455), .B2(n14454), .A(n14453), .ZN(n14465) );
  AOI21_X1 U16291 ( .B1(n14458), .B2(n14457), .A(n14456), .ZN(n14460) );
  OR2_X1 U16292 ( .A1(n14460), .A2(n14459), .ZN(n14463) );
  NAND2_X1 U16293 ( .A1(n14476), .A2(n14461), .ZN(n14462) );
  OAI211_X1 U16294 ( .C1(n14465), .C2(n14464), .A(n14463), .B(n14462), .ZN(
        n14466) );
  INV_X1 U16295 ( .A(n14466), .ZN(n14468) );
  OAI211_X1 U16296 ( .C1(n14470), .C2(n14469), .A(n14468), .B(n14467), .ZN(
        P1_U3255) );
  INV_X1 U16297 ( .A(n14471), .ZN(n14477) );
  NAND2_X1 U16298 ( .A1(n14472), .A2(P1_ADDR_REG_13__SCAN_IN), .ZN(n14474) );
  NAND2_X1 U16299 ( .A1(n14474), .A2(n14473), .ZN(n14475) );
  AOI21_X1 U16300 ( .B1(n14477), .B2(n14476), .A(n14475), .ZN(n14488) );
  OAI211_X1 U16301 ( .C1(n14481), .C2(n14480), .A(n14479), .B(n14478), .ZN(
        n14487) );
  OAI211_X1 U16302 ( .C1(n14485), .C2(n14484), .A(n14483), .B(n14482), .ZN(
        n14486) );
  NAND3_X1 U16303 ( .A1(n14488), .A2(n14487), .A3(n14486), .ZN(P1_U3256) );
  OAI21_X1 U16304 ( .B1(n14490), .B2(n14491), .A(n14489), .ZN(n14496) );
  XNOR2_X1 U16305 ( .A(n14492), .B(n14491), .ZN(n14501) );
  NOR2_X1 U16306 ( .A1(n14501), .A2(n14493), .ZN(n14494) );
  AOI211_X1 U16307 ( .C1(n14497), .C2(n14496), .A(n14495), .B(n14494), .ZN(
        n14629) );
  INV_X1 U16308 ( .A(n14498), .ZN(n14499) );
  AOI222_X1 U16309 ( .A1(n14500), .A2(n14566), .B1(P1_REG2_REG_9__SCAN_IN), 
        .B2(n6531), .C1(n14567), .C2(n14499), .ZN(n14507) );
  INV_X1 U16310 ( .A(n14501), .ZN(n14632) );
  INV_X1 U16311 ( .A(n14502), .ZN(n14575) );
  OAI211_X1 U16312 ( .C1(n14628), .C2(n14504), .A(n14546), .B(n14503), .ZN(
        n14627) );
  INV_X1 U16313 ( .A(n14627), .ZN(n14505) );
  AOI22_X1 U16314 ( .A1(n14632), .A2(n14575), .B1(n14574), .B2(n14505), .ZN(
        n14506) );
  OAI211_X1 U16315 ( .C1(n6531), .C2(n14629), .A(n14507), .B(n14506), .ZN(
        P1_U3284) );
  XNOR2_X1 U16316 ( .A(n14508), .B(n14512), .ZN(n14625) );
  INV_X1 U16317 ( .A(n14509), .ZN(n14510) );
  AOI211_X1 U16318 ( .C1(n14512), .C2(n14511), .A(n14560), .B(n14510), .ZN(
        n14513) );
  AOI211_X1 U16319 ( .C1(n14596), .C2(n14625), .A(n14514), .B(n14513), .ZN(
        n14622) );
  INV_X1 U16320 ( .A(n14515), .ZN(n14516) );
  AOI222_X1 U16321 ( .A1(n14517), .A2(n14566), .B1(P1_REG2_REG_7__SCAN_IN), 
        .B2(n6531), .C1(n14567), .C2(n14516), .ZN(n14522) );
  OAI211_X1 U16322 ( .C1(n14621), .C2(n14519), .A(n14546), .B(n14518), .ZN(
        n14620) );
  INV_X1 U16323 ( .A(n14620), .ZN(n14520) );
  AOI22_X1 U16324 ( .A1(n14625), .A2(n14575), .B1(n14574), .B2(n14520), .ZN(
        n14521) );
  OAI211_X1 U16325 ( .C1(n6531), .C2(n14622), .A(n14522), .B(n14521), .ZN(
        P1_U3286) );
  XNOR2_X1 U16326 ( .A(n14523), .B(n14524), .ZN(n14619) );
  NOR2_X1 U16327 ( .A1(n14525), .A2(n14560), .ZN(n14526) );
  AOI211_X1 U16328 ( .C1(n14596), .C2(n14619), .A(n14527), .B(n14526), .ZN(
        n14616) );
  INV_X1 U16329 ( .A(n14528), .ZN(n14529) );
  AOI222_X1 U16330 ( .A1(n14530), .A2(n14566), .B1(P1_REG2_REG_5__SCAN_IN), 
        .B2(n6531), .C1(n14567), .C2(n14529), .ZN(n14535) );
  OAI211_X1 U16331 ( .C1(n14615), .C2(n14532), .A(n14546), .B(n14531), .ZN(
        n14614) );
  INV_X1 U16332 ( .A(n14614), .ZN(n14533) );
  AOI22_X1 U16333 ( .A1(n14619), .A2(n14575), .B1(n14574), .B2(n14533), .ZN(
        n14534) );
  OAI211_X1 U16334 ( .C1(n6531), .C2(n14616), .A(n14535), .B(n14534), .ZN(
        P1_U3288) );
  XNOR2_X1 U16335 ( .A(n14536), .B(n14538), .ZN(n14603) );
  XNOR2_X1 U16336 ( .A(n14537), .B(n14538), .ZN(n14540) );
  OAI21_X1 U16337 ( .B1(n14540), .B2(n14560), .A(n14539), .ZN(n14541) );
  AOI21_X1 U16338 ( .B1(n14596), .B2(n14603), .A(n14541), .ZN(n14600) );
  OAI22_X1 U16339 ( .A1(n14543), .A2(n9116), .B1(P1_REG3_REG_3__SCAN_IN), .B2(
        n14542), .ZN(n14544) );
  AOI21_X1 U16340 ( .B1(n14566), .B2(n14545), .A(n14544), .ZN(n14551) );
  OAI211_X1 U16341 ( .C1(n14599), .C2(n14548), .A(n14547), .B(n14546), .ZN(
        n14598) );
  INV_X1 U16342 ( .A(n14598), .ZN(n14549) );
  AOI22_X1 U16343 ( .A1(n14603), .A2(n14575), .B1(n14574), .B2(n14549), .ZN(
        n14550) );
  OAI211_X1 U16344 ( .C1(n6531), .C2(n14600), .A(n14551), .B(n14550), .ZN(
        P1_U3290) );
  XNOR2_X1 U16345 ( .A(n14557), .B(n14552), .ZN(n14585) );
  NAND2_X1 U16346 ( .A1(n14553), .A2(n6539), .ZN(n14554) );
  NAND2_X1 U16347 ( .A1(n14555), .A2(n14554), .ZN(n14573) );
  XNOR2_X1 U16348 ( .A(n14573), .B(n14556), .ZN(n14559) );
  NAND2_X1 U16349 ( .A1(n14557), .A2(n14561), .ZN(n14558) );
  MUX2_X1 U16350 ( .A(n14559), .B(n14558), .S(n8344), .Z(n14564) );
  INV_X1 U16351 ( .A(n8344), .ZN(n14562) );
  OAI21_X1 U16352 ( .B1(n14562), .B2(n14561), .A(n14560), .ZN(n14563) );
  AOI22_X1 U16353 ( .A1(n14596), .A2(n14585), .B1(n14564), .B2(n14563), .ZN(
        n14587) );
  NAND2_X1 U16354 ( .A1(n14566), .A2(n6539), .ZN(n14569) );
  AOI22_X1 U16355 ( .A1(n6531), .A2(P1_REG2_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(n14567), .ZN(n14568) );
  OAI211_X1 U16356 ( .C1(n14570), .C2(n14582), .A(n14569), .B(n14568), .ZN(
        n14571) );
  INV_X1 U16357 ( .A(n14571), .ZN(n14577) );
  NOR2_X1 U16358 ( .A1(n14573), .A2(n14572), .ZN(n14584) );
  AOI22_X1 U16359 ( .A1(n14575), .A2(n14585), .B1(n14574), .B2(n14584), .ZN(
        n14576) );
  OAI211_X1 U16360 ( .C1(n6531), .C2(n14587), .A(n14577), .B(n14576), .ZN(
        P1_U3292) );
  AND2_X1 U16361 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n14579), .ZN(P1_U3294) );
  AND2_X1 U16362 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n14579), .ZN(P1_U3295) );
  AND2_X1 U16363 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n14579), .ZN(P1_U3296) );
  INV_X1 U16364 ( .A(n14579), .ZN(n14578) );
  INV_X1 U16365 ( .A(P1_D_REG_28__SCAN_IN), .ZN(n15185) );
  NOR2_X1 U16366 ( .A1(n14578), .A2(n15185), .ZN(P1_U3297) );
  AND2_X1 U16367 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n14579), .ZN(P1_U3298) );
  AND2_X1 U16368 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n14579), .ZN(P1_U3299) );
  AND2_X1 U16369 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n14579), .ZN(P1_U3300) );
  AND2_X1 U16370 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n14579), .ZN(P1_U3301) );
  AND2_X1 U16371 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n14579), .ZN(P1_U3302) );
  AND2_X1 U16372 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n14579), .ZN(P1_U3303) );
  AND2_X1 U16373 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n14579), .ZN(P1_U3304) );
  AND2_X1 U16374 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n14579), .ZN(P1_U3305) );
  AND2_X1 U16375 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n14579), .ZN(P1_U3306) );
  INV_X1 U16376 ( .A(P1_D_REG_18__SCAN_IN), .ZN(n15157) );
  NOR2_X1 U16377 ( .A1(n14578), .A2(n15157), .ZN(P1_U3307) );
  AND2_X1 U16378 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n14579), .ZN(P1_U3308) );
  AND2_X1 U16379 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n14579), .ZN(P1_U3309) );
  AND2_X1 U16380 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n14579), .ZN(P1_U3310) );
  AND2_X1 U16381 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n14579), .ZN(P1_U3311) );
  AND2_X1 U16382 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n14579), .ZN(P1_U3312) );
  AND2_X1 U16383 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n14579), .ZN(P1_U3313) );
  INV_X1 U16384 ( .A(P1_D_REG_11__SCAN_IN), .ZN(n15369) );
  NOR2_X1 U16385 ( .A1(n14578), .A2(n15369), .ZN(P1_U3314) );
  AND2_X1 U16386 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n14579), .ZN(P1_U3315) );
  AND2_X1 U16387 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n14579), .ZN(P1_U3316) );
  AND2_X1 U16388 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n14579), .ZN(P1_U3317) );
  AND2_X1 U16389 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n14579), .ZN(P1_U3318) );
  AND2_X1 U16390 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n14579), .ZN(P1_U3319) );
  AND2_X1 U16391 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n14579), .ZN(P1_U3320) );
  AND2_X1 U16392 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n14579), .ZN(P1_U3321) );
  AND2_X1 U16393 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n14579), .ZN(P1_U3322) );
  AND2_X1 U16394 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n14579), .ZN(P1_U3323) );
  INV_X1 U16395 ( .A(n14592), .ZN(n14633) );
  OAI22_X1 U16396 ( .A1(n14582), .A2(n14581), .B1(n14580), .B2(n14638), .ZN(
        n14583) );
  AOI211_X1 U16397 ( .C1(n14585), .C2(n14633), .A(n14584), .B(n14583), .ZN(
        n14586) );
  AND2_X1 U16398 ( .A1(n14587), .A2(n14586), .ZN(n14646) );
  INV_X1 U16399 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n15167) );
  AOI22_X1 U16400 ( .A1(n14645), .A2(n14646), .B1(n15167), .B2(n14643), .ZN(
        P1_U3462) );
  AOI21_X1 U16401 ( .B1(n14589), .B2(n14607), .A(n14588), .ZN(n14590) );
  OAI211_X1 U16402 ( .C1(n14593), .C2(n14592), .A(n14591), .B(n14590), .ZN(
        n14594) );
  AOI21_X1 U16403 ( .B1(n14596), .B2(n14595), .A(n14594), .ZN(n14647) );
  INV_X1 U16404 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n14597) );
  AOI22_X1 U16405 ( .A1(n14645), .A2(n14647), .B1(n14597), .B2(n14643), .ZN(
        P1_U3465) );
  OAI21_X1 U16406 ( .B1(n14599), .B2(n14638), .A(n14598), .ZN(n14602) );
  INV_X1 U16407 ( .A(n14600), .ZN(n14601) );
  AOI211_X1 U16408 ( .C1(n14633), .C2(n14603), .A(n14602), .B(n14601), .ZN(
        n14648) );
  INV_X1 U16409 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n14604) );
  AOI22_X1 U16410 ( .A1(n14645), .A2(n14648), .B1(n14604), .B2(n14643), .ZN(
        P1_U3468) );
  AOI211_X1 U16411 ( .C1(n14608), .C2(n14607), .A(n14606), .B(n14605), .ZN(
        n14609) );
  OAI21_X1 U16412 ( .B1(n14611), .B2(n14610), .A(n14609), .ZN(n14612) );
  INV_X1 U16413 ( .A(n14612), .ZN(n14649) );
  INV_X1 U16414 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n14613) );
  AOI22_X1 U16415 ( .A1(n14645), .A2(n14649), .B1(n14613), .B2(n14643), .ZN(
        P1_U3471) );
  OAI21_X1 U16416 ( .B1(n14615), .B2(n14638), .A(n14614), .ZN(n14618) );
  INV_X1 U16417 ( .A(n14616), .ZN(n14617) );
  AOI211_X1 U16418 ( .C1(n14633), .C2(n14619), .A(n14618), .B(n14617), .ZN(
        n14650) );
  INV_X1 U16419 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n15160) );
  AOI22_X1 U16420 ( .A1(n14645), .A2(n14650), .B1(n15160), .B2(n14643), .ZN(
        P1_U3474) );
  OAI21_X1 U16421 ( .B1(n14621), .B2(n14638), .A(n14620), .ZN(n14624) );
  INV_X1 U16422 ( .A(n14622), .ZN(n14623) );
  AOI211_X1 U16423 ( .C1(n14633), .C2(n14625), .A(n14624), .B(n14623), .ZN(
        n14652) );
  INV_X1 U16424 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n14626) );
  AOI22_X1 U16425 ( .A1(n14645), .A2(n14652), .B1(n14626), .B2(n14643), .ZN(
        P1_U3480) );
  OAI21_X1 U16426 ( .B1(n14628), .B2(n14638), .A(n14627), .ZN(n14631) );
  INV_X1 U16427 ( .A(n14629), .ZN(n14630) );
  AOI211_X1 U16428 ( .C1(n14633), .C2(n14632), .A(n14631), .B(n14630), .ZN(
        n14654) );
  INV_X1 U16429 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n14634) );
  AOI22_X1 U16430 ( .A1(n14645), .A2(n14654), .B1(n14634), .B2(n14643), .ZN(
        P1_U3486) );
  INV_X1 U16431 ( .A(n14635), .ZN(n14639) );
  OAI211_X1 U16432 ( .C1(n14639), .C2(n14638), .A(n14637), .B(n14636), .ZN(
        n14640) );
  AOI21_X1 U16433 ( .B1(n14642), .B2(n14641), .A(n14640), .ZN(n14657) );
  INV_X1 U16434 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n14644) );
  AOI22_X1 U16435 ( .A1(n14645), .A2(n14657), .B1(n14644), .B2(n14643), .ZN(
        P1_U3489) );
  AOI22_X1 U16436 ( .A1(n14658), .A2(n14646), .B1(n8358), .B2(n14655), .ZN(
        P1_U3529) );
  AOI22_X1 U16437 ( .A1(n14658), .A2(n14647), .B1(n8371), .B2(n14655), .ZN(
        P1_U3530) );
  AOI22_X1 U16438 ( .A1(n14658), .A2(n14648), .B1(n8385), .B2(n14655), .ZN(
        P1_U3531) );
  AOI22_X1 U16439 ( .A1(n14658), .A2(n14649), .B1(n9103), .B2(n14655), .ZN(
        P1_U3532) );
  AOI22_X1 U16440 ( .A1(n14658), .A2(n14650), .B1(n9107), .B2(n14655), .ZN(
        P1_U3533) );
  AOI22_X1 U16441 ( .A1(n14658), .A2(n14652), .B1(n14651), .B2(n14655), .ZN(
        P1_U3535) );
  AOI22_X1 U16442 ( .A1(n14658), .A2(n14654), .B1(n14653), .B2(n14655), .ZN(
        P1_U3537) );
  AOI22_X1 U16443 ( .A1(n14658), .A2(n14657), .B1(n14656), .B2(n14655), .ZN(
        P1_U3538) );
  NOR2_X1 U16444 ( .A1(n14752), .A2(P2_U3947), .ZN(P2_U3087) );
  INV_X1 U16445 ( .A(n14659), .ZN(n14667) );
  MUX2_X1 U16446 ( .A(P2_REG1_REG_4__SCAN_IN), .B(n9325), .S(n14660), .Z(
        n14661) );
  NAND3_X1 U16447 ( .A1(n14663), .A2(n14662), .A3(n14661), .ZN(n14664) );
  AND3_X1 U16448 ( .A1(n14759), .A2(n14665), .A3(n14664), .ZN(n14666) );
  AOI211_X1 U16449 ( .C1(n14754), .C2(n14668), .A(n14667), .B(n14666), .ZN(
        n14672) );
  OAI211_X1 U16450 ( .C1(n14670), .C2(n14669), .A(n14756), .B(n14676), .ZN(
        n14671) );
  OAI211_X1 U16451 ( .C1(n14736), .C2(n15156), .A(n14672), .B(n14671), .ZN(
        P2_U3218) );
  INV_X1 U16452 ( .A(n14673), .ZN(n14680) );
  MUX2_X1 U16453 ( .A(n10171), .B(P2_REG2_REG_5__SCAN_IN), .S(n14681), .Z(
        n14674) );
  NAND3_X1 U16454 ( .A1(n14676), .A2(n14675), .A3(n14674), .ZN(n14677) );
  AND3_X1 U16455 ( .A1(n14756), .A2(n14678), .A3(n14677), .ZN(n14679) );
  AOI211_X1 U16456 ( .C1(n14754), .C2(n14681), .A(n14680), .B(n14679), .ZN(
        n14686) );
  OAI211_X1 U16457 ( .C1(n14684), .C2(n14683), .A(n14759), .B(n14682), .ZN(
        n14685) );
  OAI211_X1 U16458 ( .C1(n14736), .C2(n15411), .A(n14686), .B(n14685), .ZN(
        P2_U3219) );
  NAND2_X1 U16459 ( .A1(n14688), .A2(n14687), .ZN(n14689) );
  NAND2_X1 U16460 ( .A1(n14690), .A2(n14689), .ZN(n14691) );
  NAND2_X1 U16461 ( .A1(n14691), .A2(n14756), .ZN(n14698) );
  NAND2_X1 U16462 ( .A1(n14693), .A2(n14692), .ZN(n14694) );
  NAND2_X1 U16463 ( .A1(n14695), .A2(n14694), .ZN(n14696) );
  NAND2_X1 U16464 ( .A1(n14696), .A2(n14759), .ZN(n14697) );
  OAI211_X1 U16465 ( .C1(n14739), .C2(n14699), .A(n14698), .B(n14697), .ZN(
        n14700) );
  INV_X1 U16466 ( .A(n14700), .ZN(n14702) );
  OAI211_X1 U16467 ( .C1(n14703), .C2(n14736), .A(n14702), .B(n14701), .ZN(
        P2_U3223) );
  NOR2_X1 U16468 ( .A1(n14739), .A2(n14704), .ZN(n14705) );
  AOI211_X1 U16469 ( .C1(n14752), .C2(P2_ADDR_REG_10__SCAN_IN), .A(n14706), 
        .B(n14705), .ZN(n14718) );
  AOI21_X1 U16470 ( .B1(n14708), .B2(n14707), .A(n14745), .ZN(n14710) );
  NAND2_X1 U16471 ( .A1(n14710), .A2(n14709), .ZN(n14717) );
  AOI21_X1 U16472 ( .B1(n14713), .B2(n14712), .A(n14711), .ZN(n14715) );
  NAND2_X1 U16473 ( .A1(n14715), .A2(n14714), .ZN(n14716) );
  NAND3_X1 U16474 ( .A1(n14718), .A2(n14717), .A3(n14716), .ZN(P2_U3224) );
  NOR2_X1 U16475 ( .A1(n14720), .A2(n14719), .ZN(n14721) );
  OAI21_X1 U16476 ( .B1(n14722), .B2(n14721), .A(n14759), .ZN(n14731) );
  INV_X1 U16477 ( .A(n14723), .ZN(n14725) );
  NAND3_X1 U16478 ( .A1(n14726), .A2(n14725), .A3(n14724), .ZN(n14727) );
  NAND2_X1 U16479 ( .A1(n14728), .A2(n14727), .ZN(n14729) );
  NAND2_X1 U16480 ( .A1(n14729), .A2(n14756), .ZN(n14730) );
  OAI211_X1 U16481 ( .C1(n14739), .C2(n14732), .A(n14731), .B(n14730), .ZN(
        n14733) );
  INV_X1 U16482 ( .A(n14733), .ZN(n14735) );
  OAI211_X1 U16483 ( .C1(n15365), .C2(n14736), .A(n14735), .B(n14734), .ZN(
        P2_U3226) );
  OAI21_X1 U16484 ( .B1(n14739), .B2(n14738), .A(n14737), .ZN(n14740) );
  AOI21_X1 U16485 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(n14752), .A(n14740), 
        .ZN(n14751) );
  OAI211_X1 U16486 ( .C1(n14743), .C2(n14742), .A(n14741), .B(n14759), .ZN(
        n14750) );
  AOI211_X1 U16487 ( .C1(n14747), .C2(n14746), .A(n14745), .B(n14744), .ZN(
        n14748) );
  INV_X1 U16488 ( .A(n14748), .ZN(n14749) );
  NAND3_X1 U16489 ( .A1(n14751), .A2(n14750), .A3(n14749), .ZN(P2_U3227) );
  AOI22_X1 U16490 ( .A1(n14752), .A2(P2_ADDR_REG_15__SCAN_IN), .B1(
        P2_REG3_REG_15__SCAN_IN), .B2(P2_U3088), .ZN(n14764) );
  NAND2_X1 U16491 ( .A1(n14754), .A2(n14753), .ZN(n14763) );
  OAI211_X1 U16492 ( .C1(P2_REG2_REG_15__SCAN_IN), .C2(n14757), .A(n14756), 
        .B(n14755), .ZN(n14762) );
  OAI211_X1 U16493 ( .C1(n14760), .C2(P2_REG1_REG_15__SCAN_IN), .A(n14759), 
        .B(n14758), .ZN(n14761) );
  NAND4_X1 U16494 ( .A1(n14764), .A2(n14763), .A3(n14762), .A4(n14761), .ZN(
        P2_U3229) );
  NOR2_X1 U16495 ( .A1(n14770), .A2(n14765), .ZN(n14766) );
  AND2_X1 U16496 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n14767), .ZN(P2_U3266) );
  AND2_X1 U16497 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n14767), .ZN(P2_U3267) );
  AND2_X1 U16498 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n14767), .ZN(P2_U3268) );
  INV_X1 U16499 ( .A(P2_D_REG_28__SCAN_IN), .ZN(n15184) );
  NOR2_X1 U16500 ( .A1(n14766), .A2(n15184), .ZN(P2_U3269) );
  AND2_X1 U16501 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n14767), .ZN(P2_U3270) );
  AND2_X1 U16502 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n14767), .ZN(P2_U3271) );
  INV_X1 U16503 ( .A(P2_D_REG_25__SCAN_IN), .ZN(n15236) );
  NOR2_X1 U16504 ( .A1(n14766), .A2(n15236), .ZN(P2_U3272) );
  AND2_X1 U16505 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n14767), .ZN(P2_U3273) );
  AND2_X1 U16506 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n14767), .ZN(P2_U3274) );
  AND2_X1 U16507 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n14767), .ZN(P2_U3275) );
  AND2_X1 U16508 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n14767), .ZN(P2_U3276) );
  AND2_X1 U16509 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n14767), .ZN(P2_U3277) );
  AND2_X1 U16510 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n14767), .ZN(P2_U3278) );
  INV_X1 U16511 ( .A(P2_D_REG_18__SCAN_IN), .ZN(n15201) );
  NOR2_X1 U16512 ( .A1(n14766), .A2(n15201), .ZN(P2_U3279) );
  AND2_X1 U16513 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n14767), .ZN(P2_U3280) );
  AND2_X1 U16514 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n14767), .ZN(P2_U3281) );
  AND2_X1 U16515 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n14767), .ZN(P2_U3282) );
  AND2_X1 U16516 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n14767), .ZN(P2_U3283) );
  AND2_X1 U16517 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n14767), .ZN(P2_U3284) );
  AND2_X1 U16518 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n14767), .ZN(P2_U3285) );
  AND2_X1 U16519 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n14767), .ZN(P2_U3286) );
  INV_X1 U16520 ( .A(P2_D_REG_10__SCAN_IN), .ZN(n15309) );
  NOR2_X1 U16521 ( .A1(n14766), .A2(n15309), .ZN(P2_U3287) );
  AND2_X1 U16522 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n14767), .ZN(P2_U3288) );
  AND2_X1 U16523 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n14767), .ZN(P2_U3289) );
  INV_X1 U16524 ( .A(P2_D_REG_7__SCAN_IN), .ZN(n15214) );
  NOR2_X1 U16525 ( .A1(n14766), .A2(n15214), .ZN(P2_U3290) );
  AND2_X1 U16526 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n14767), .ZN(P2_U3291) );
  AND2_X1 U16527 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n14767), .ZN(P2_U3292) );
  AND2_X1 U16528 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n14767), .ZN(P2_U3293) );
  AND2_X1 U16529 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n14767), .ZN(P2_U3294) );
  AND2_X1 U16530 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n14767), .ZN(P2_U3295) );
  AOI22_X1 U16531 ( .A1(n14773), .A2(n14769), .B1(n14768), .B2(n14770), .ZN(
        P2_U3416) );
  AOI22_X1 U16532 ( .A1(n14773), .A2(n14772), .B1(n14771), .B2(n14770), .ZN(
        P2_U3417) );
  INV_X1 U16533 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n14774) );
  AOI22_X1 U16534 ( .A1(n14821), .A2(n14775), .B1(n14774), .B2(n14819), .ZN(
        P2_U3430) );
  AOI21_X1 U16535 ( .B1(n6538), .B2(n14803), .A(n14776), .ZN(n14780) );
  OAI211_X1 U16536 ( .C1(n6795), .C2(n14806), .A(n14778), .B(n14777), .ZN(
        n14779) );
  NOR2_X1 U16537 ( .A1(n14780), .A2(n14779), .ZN(n14822) );
  AOI22_X1 U16538 ( .A1(n14821), .A2(n14822), .B1(n7673), .B2(n14819), .ZN(
        P2_U3445) );
  AOI21_X1 U16539 ( .B1(n14810), .B2(n14782), .A(n14781), .ZN(n14783) );
  OAI211_X1 U16540 ( .C1(n14785), .C2(n14803), .A(n14784), .B(n14783), .ZN(
        n14786) );
  INV_X1 U16541 ( .A(n14786), .ZN(n14823) );
  AOI22_X1 U16542 ( .A1(n14821), .A2(n14823), .B1(n7689), .B2(n14819), .ZN(
        P2_U3448) );
  AOI21_X1 U16543 ( .B1(n14810), .B2(n14788), .A(n14787), .ZN(n14789) );
  OAI211_X1 U16544 ( .C1(n14792), .C2(n14791), .A(n14790), .B(n14789), .ZN(
        n14793) );
  INV_X1 U16545 ( .A(n14793), .ZN(n14824) );
  AOI22_X1 U16546 ( .A1(n14821), .A2(n14824), .B1(n7707), .B2(n14819), .ZN(
        P2_U3451) );
  OR2_X1 U16547 ( .A1(n14794), .A2(n14803), .ZN(n14801) );
  OR2_X1 U16548 ( .A1(n14794), .A2(n6538), .ZN(n14800) );
  NAND2_X1 U16549 ( .A1(n14795), .A2(n14810), .ZN(n14796) );
  AND2_X1 U16550 ( .A1(n14797), .A2(n14796), .ZN(n14798) );
  AND4_X1 U16551 ( .A1(n14801), .A2(n14800), .A3(n14799), .A4(n14798), .ZN(
        n14825) );
  AOI22_X1 U16552 ( .A1(n14821), .A2(n14825), .B1(n7723), .B2(n14819), .ZN(
        P2_U3454) );
  AOI21_X1 U16553 ( .B1(n6538), .B2(n14803), .A(n14802), .ZN(n14809) );
  OAI211_X1 U16554 ( .C1(n14807), .C2(n14806), .A(n14805), .B(n14804), .ZN(
        n14808) );
  NOR2_X1 U16555 ( .A1(n14809), .A2(n14808), .ZN(n14826) );
  AOI22_X1 U16556 ( .A1(n14821), .A2(n14826), .B1(n7744), .B2(n14819), .ZN(
        P2_U3457) );
  NAND2_X1 U16557 ( .A1(n14811), .A2(n14810), .ZN(n14812) );
  NAND2_X1 U16558 ( .A1(n14813), .A2(n14812), .ZN(n14814) );
  AOI21_X1 U16559 ( .B1(n14816), .B2(n14815), .A(n14814), .ZN(n14817) );
  AND2_X1 U16560 ( .A1(n14818), .A2(n14817), .ZN(n14828) );
  INV_X1 U16561 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n14820) );
  AOI22_X1 U16562 ( .A1(n14821), .A2(n14828), .B1(n14820), .B2(n14819), .ZN(
        P2_U3460) );
  AOI22_X1 U16563 ( .A1(n14829), .A2(n14822), .B1(n9329), .B2(n14827), .ZN(
        P2_U3504) );
  AOI22_X1 U16564 ( .A1(n14829), .A2(n14823), .B1(n9330), .B2(n14827), .ZN(
        P2_U3505) );
  AOI22_X1 U16565 ( .A1(n14829), .A2(n14824), .B1(n9333), .B2(n14827), .ZN(
        P2_U3506) );
  AOI22_X1 U16566 ( .A1(n14829), .A2(n14825), .B1(n9336), .B2(n14827), .ZN(
        P2_U3507) );
  AOI22_X1 U16567 ( .A1(n14829), .A2(n14826), .B1(n9340), .B2(n14827), .ZN(
        P2_U3508) );
  AOI22_X1 U16568 ( .A1(n14829), .A2(n14828), .B1(n7756), .B2(n14827), .ZN(
        P2_U3509) );
  NOR2_X1 U16569 ( .A1(P3_U3897), .A2(n14969), .ZN(P3_U3150) );
  NOR2_X1 U16570 ( .A1(n14830), .A2(P3_REG2_REG_3__SCAN_IN), .ZN(n14832) );
  NOR2_X1 U16571 ( .A1(n14832), .A2(n14831), .ZN(n14848) );
  OAI21_X1 U16572 ( .B1(n14834), .B2(n8211), .A(n14833), .ZN(n14841) );
  OR3_X1 U16573 ( .A1(n14837), .A2(n14836), .A3(n14835), .ZN(n14839) );
  AOI21_X1 U16574 ( .B1(n14854), .B2(n14839), .A(n14838), .ZN(n14840) );
  AOI211_X1 U16575 ( .C1(n14843), .C2(n14842), .A(n14841), .B(n14840), .ZN(
        n14847) );
  XNOR2_X1 U16576 ( .A(n14844), .B(P3_REG1_REG_3__SCAN_IN), .ZN(n14845) );
  NAND2_X1 U16577 ( .A1(n14973), .A2(n14845), .ZN(n14846) );
  OAI211_X1 U16578 ( .C1(n14848), .C2(n14977), .A(n14847), .B(n14846), .ZN(
        P3_U3185) );
  AOI21_X1 U16579 ( .B1(n14851), .B2(n14850), .A(n14849), .ZN(n14866) );
  AND3_X1 U16580 ( .A1(n14854), .A2(n14853), .A3(n14852), .ZN(n14855) );
  OAI21_X1 U16581 ( .B1(n14871), .B2(n14855), .A(n14961), .ZN(n14856) );
  OAI21_X1 U16582 ( .B1(n14966), .B2(n14857), .A(n14856), .ZN(n14858) );
  AOI211_X1 U16583 ( .C1(P3_ADDR_REG_4__SCAN_IN), .C2(n14969), .A(n14859), .B(
        n14858), .ZN(n14865) );
  OAI21_X1 U16584 ( .B1(n14862), .B2(n14861), .A(n14860), .ZN(n14863) );
  NAND2_X1 U16585 ( .A1(n14973), .A2(n14863), .ZN(n14864) );
  OAI211_X1 U16586 ( .C1(n14866), .C2(n14977), .A(n14865), .B(n14864), .ZN(
        P3_U3186) );
  AOI21_X1 U16587 ( .B1(n10928), .B2(n14868), .A(n14867), .ZN(n14883) );
  INV_X1 U16588 ( .A(n14890), .ZN(n14873) );
  NOR3_X1 U16589 ( .A1(n14871), .A2(n14870), .A3(n14869), .ZN(n14872) );
  OAI21_X1 U16590 ( .B1(n14873), .B2(n14872), .A(n14961), .ZN(n14874) );
  OAI21_X1 U16591 ( .B1(n14966), .B2(n14875), .A(n14874), .ZN(n14876) );
  AOI211_X1 U16592 ( .C1(P3_ADDR_REG_5__SCAN_IN), .C2(n14969), .A(n14877), .B(
        n14876), .ZN(n14882) );
  OAI21_X1 U16593 ( .B1(P3_REG1_REG_5__SCAN_IN), .B2(n14879), .A(n14878), .ZN(
        n14880) );
  NAND2_X1 U16594 ( .A1(n14973), .A2(n14880), .ZN(n14881) );
  OAI211_X1 U16595 ( .C1(n14883), .C2(n14977), .A(n14882), .B(n14881), .ZN(
        P3_U3187) );
  INV_X1 U16596 ( .A(n14884), .ZN(n14885) );
  AOI21_X1 U16597 ( .B1(n14887), .B2(n14886), .A(n14885), .ZN(n14902) );
  AND3_X1 U16598 ( .A1(n14890), .A2(n14889), .A3(n14888), .ZN(n14891) );
  OAI21_X1 U16599 ( .B1(n14907), .B2(n14891), .A(n14961), .ZN(n14892) );
  OAI21_X1 U16600 ( .B1(n14966), .B2(n14893), .A(n14892), .ZN(n14894) );
  AOI211_X1 U16601 ( .C1(P3_ADDR_REG_6__SCAN_IN), .C2(n14969), .A(n14895), .B(
        n14894), .ZN(n14901) );
  OAI21_X1 U16602 ( .B1(n14898), .B2(n14897), .A(n14896), .ZN(n14899) );
  NAND2_X1 U16603 ( .A1(n14973), .A2(n14899), .ZN(n14900) );
  OAI211_X1 U16604 ( .C1(n14902), .C2(n14977), .A(n14901), .B(n14900), .ZN(
        P3_U3188) );
  AOI21_X1 U16605 ( .B1(n10940), .B2(n14904), .A(n14903), .ZN(n14919) );
  INV_X1 U16606 ( .A(n14925), .ZN(n14909) );
  NOR3_X1 U16607 ( .A1(n14907), .A2(n14906), .A3(n14905), .ZN(n14908) );
  OAI21_X1 U16608 ( .B1(n14909), .B2(n14908), .A(n14961), .ZN(n14910) );
  OAI21_X1 U16609 ( .B1(n14966), .B2(n14911), .A(n14910), .ZN(n14912) );
  AOI211_X1 U16610 ( .C1(P3_ADDR_REG_7__SCAN_IN), .C2(n14969), .A(n14913), .B(
        n14912), .ZN(n14918) );
  OAI21_X1 U16611 ( .B1(P3_REG1_REG_7__SCAN_IN), .B2(n14915), .A(n14914), .ZN(
        n14916) );
  NAND2_X1 U16612 ( .A1(n14916), .A2(n14973), .ZN(n14917) );
  OAI211_X1 U16613 ( .C1(n14919), .C2(n14977), .A(n14918), .B(n14917), .ZN(
        P3_U3189) );
  AOI21_X1 U16614 ( .B1(n14922), .B2(n14921), .A(n14920), .ZN(n14937) );
  AND3_X1 U16615 ( .A1(n14925), .A2(n14924), .A3(n14923), .ZN(n14926) );
  OAI21_X1 U16616 ( .B1(n14942), .B2(n14926), .A(n14961), .ZN(n14927) );
  OAI21_X1 U16617 ( .B1(n14966), .B2(n14928), .A(n14927), .ZN(n14929) );
  AOI211_X1 U16618 ( .C1(P3_ADDR_REG_8__SCAN_IN), .C2(n14969), .A(n14930), .B(
        n14929), .ZN(n14936) );
  OAI21_X1 U16619 ( .B1(n14933), .B2(n14932), .A(n14931), .ZN(n14934) );
  NAND2_X1 U16620 ( .A1(n14934), .A2(n14973), .ZN(n14935) );
  OAI211_X1 U16621 ( .C1(n14937), .C2(n14977), .A(n14936), .B(n14935), .ZN(
        P3_U3190) );
  AOI21_X1 U16622 ( .B1(n10953), .B2(n14939), .A(n14938), .ZN(n14954) );
  INV_X1 U16623 ( .A(n14960), .ZN(n14944) );
  NOR3_X1 U16624 ( .A1(n14942), .A2(n14941), .A3(n14940), .ZN(n14943) );
  OAI21_X1 U16625 ( .B1(n14944), .B2(n14943), .A(n14961), .ZN(n14945) );
  OAI21_X1 U16626 ( .B1(n14966), .B2(n14946), .A(n14945), .ZN(n14947) );
  AOI211_X1 U16627 ( .C1(P3_ADDR_REG_9__SCAN_IN), .C2(n14969), .A(n14948), .B(
        n14947), .ZN(n14953) );
  OAI21_X1 U16628 ( .B1(P3_REG1_REG_9__SCAN_IN), .B2(n14950), .A(n14949), .ZN(
        n14951) );
  NAND2_X1 U16629 ( .A1(n14951), .A2(n14973), .ZN(n14952) );
  OAI211_X1 U16630 ( .C1(n14954), .C2(n14977), .A(n14953), .B(n14952), .ZN(
        P3_U3191) );
  AOI21_X1 U16631 ( .B1(n14957), .B2(n14956), .A(n14955), .ZN(n14978) );
  AND3_X1 U16632 ( .A1(n14960), .A2(n14959), .A3(n14958), .ZN(n14962) );
  OAI21_X1 U16633 ( .B1(n14963), .B2(n14962), .A(n14961), .ZN(n14964) );
  OAI21_X1 U16634 ( .B1(n14966), .B2(n14965), .A(n14964), .ZN(n14967) );
  AOI211_X1 U16635 ( .C1(P3_ADDR_REG_10__SCAN_IN), .C2(n14969), .A(n14968), 
        .B(n14967), .ZN(n14976) );
  OAI21_X1 U16636 ( .B1(n14972), .B2(n14971), .A(n14970), .ZN(n14974) );
  NAND2_X1 U16637 ( .A1(n14974), .A2(n14973), .ZN(n14975) );
  OAI211_X1 U16638 ( .C1(n14978), .C2(n14977), .A(n14976), .B(n14975), .ZN(
        P3_U3192) );
  AOI21_X1 U16639 ( .B1(n14982), .B2(n14980), .A(n14979), .ZN(n15084) );
  OAI211_X1 U16640 ( .C1(n14983), .C2(n14982), .A(n14981), .B(n15046), .ZN(
        n14987) );
  AOI22_X1 U16641 ( .A1(n15041), .A2(n14985), .B1(n14984), .B2(n15038), .ZN(
        n14986) );
  NAND2_X1 U16642 ( .A1(n14987), .A2(n14986), .ZN(n15081) );
  AOI21_X1 U16643 ( .B1(n15084), .B2(n15033), .A(n15081), .ZN(n14993) );
  AND2_X1 U16644 ( .A1(n14988), .A2(n15049), .ZN(n15082) );
  NOR2_X1 U16645 ( .A1(n15020), .A2(n14989), .ZN(n14990) );
  AOI21_X1 U16646 ( .B1(n14991), .B2(n15082), .A(n14990), .ZN(n14992) );
  OAI221_X1 U16647 ( .B1(n15052), .B2(n14993), .C1(n15057), .C2(n10959), .A(
        n14992), .ZN(P3_U3223) );
  OAI21_X1 U16648 ( .B1(n15010), .B2(n14995), .A(n14994), .ZN(n14998) );
  AOI222_X1 U16649 ( .A1(n15057), .A2(n14998), .B1(n14997), .B2(n15055), .C1(
        n14996), .C2(n15014), .ZN(n14999) );
  OAI21_X1 U16650 ( .B1(n15057), .B2(n10946), .A(n14999), .ZN(P3_U3225) );
  OAI21_X1 U16651 ( .B1(n15001), .B2(n15010), .A(n15000), .ZN(n15002) );
  MUX2_X1 U16652 ( .A(P3_REG2_REG_7__SCAN_IN), .B(n15002), .S(n15057), .Z(
        n15003) );
  AOI21_X1 U16653 ( .B1(n15014), .B2(n15004), .A(n15003), .ZN(n15005) );
  OAI21_X1 U16654 ( .B1(n15006), .B2(n15020), .A(n15005), .ZN(P3_U3226) );
  INV_X1 U16655 ( .A(n15007), .ZN(n15009) );
  OAI21_X1 U16656 ( .B1(n15010), .B2(n15009), .A(n15008), .ZN(n15011) );
  MUX2_X1 U16657 ( .A(P3_REG2_REG_6__SCAN_IN), .B(n15011), .S(n15057), .Z(
        n15012) );
  AOI21_X1 U16658 ( .B1(n15014), .B2(n15013), .A(n15012), .ZN(n15015) );
  OAI21_X1 U16659 ( .B1(n15016), .B2(n15020), .A(n15015), .ZN(P3_U3227) );
  OAI21_X1 U16660 ( .B1(n15017), .B2(n15025), .A(n11683), .ZN(n15066) );
  NOR2_X1 U16661 ( .A1(n15019), .A2(n15018), .ZN(n15065) );
  INV_X1 U16662 ( .A(n15065), .ZN(n15023) );
  OAI22_X1 U16663 ( .A1(n15023), .A2(n15022), .B1(n15021), .B2(n15020), .ZN(
        n15032) );
  XNOR2_X1 U16664 ( .A(n15024), .B(n15025), .ZN(n15026) );
  OAI222_X1 U16665 ( .A1(n15031), .A2(n15030), .B1(n15029), .B2(n15028), .C1(
        n15027), .C2(n15026), .ZN(n15064) );
  AOI211_X1 U16666 ( .C1(n15033), .C2(n15066), .A(n15032), .B(n15064), .ZN(
        n15034) );
  AOI22_X1 U16667 ( .A1(n15052), .A2(n10045), .B1(n15034), .B2(n15057), .ZN(
        P3_U3231) );
  XNOR2_X1 U16668 ( .A(n10097), .B(n15035), .ZN(n15045) );
  AND2_X1 U16669 ( .A1(n15037), .A2(n15036), .ZN(n15047) );
  AOI22_X1 U16670 ( .A1(n15041), .A2(n15040), .B1(n15039), .B2(n15038), .ZN(
        n15042) );
  OAI21_X1 U16671 ( .B1(n15047), .B2(n15043), .A(n15042), .ZN(n15044) );
  AOI21_X1 U16672 ( .B1(n15046), .B2(n15045), .A(n15044), .ZN(n15059) );
  INV_X1 U16673 ( .A(n15047), .ZN(n15062) );
  AND2_X1 U16674 ( .A1(n15049), .A2(n15048), .ZN(n15061) );
  AOI22_X1 U16675 ( .A1(n15062), .A2(n15051), .B1(n15061), .B2(n15050), .ZN(
        n15053) );
  AOI21_X1 U16676 ( .B1(n15059), .B2(n15053), .A(n15052), .ZN(n15054) );
  AOI21_X1 U16677 ( .B1(P3_REG3_REG_1__SCAN_IN), .B2(n15055), .A(n15054), .ZN(
        n15056) );
  OAI21_X1 U16678 ( .B1(n9739), .B2(n15057), .A(n15056), .ZN(P3_U3232) );
  INV_X1 U16679 ( .A(n15058), .ZN(n15063) );
  INV_X1 U16680 ( .A(n15059), .ZN(n15060) );
  AOI211_X1 U16681 ( .C1(n15063), .C2(n15062), .A(n15061), .B(n15060), .ZN(
        n15088) );
  AOI22_X1 U16682 ( .A1(n15086), .A2(n9737), .B1(n15088), .B2(n15085), .ZN(
        P3_U3393) );
  AOI211_X1 U16683 ( .C1(n15083), .C2(n15066), .A(n15065), .B(n15064), .ZN(
        n15089) );
  AOI22_X1 U16684 ( .A1(n15086), .A2(n9392), .B1(n15089), .B2(n15085), .ZN(
        P3_U3396) );
  INV_X1 U16685 ( .A(P3_REG0_REG_3__SCAN_IN), .ZN(n15070) );
  AOI211_X1 U16686 ( .C1(n15069), .C2(n15083), .A(n15068), .B(n15067), .ZN(
        n15090) );
  AOI22_X1 U16687 ( .A1(n15086), .A2(n15070), .B1(n15090), .B2(n15085), .ZN(
        P3_U3399) );
  INV_X1 U16688 ( .A(n15071), .ZN(n15073) );
  AOI211_X1 U16689 ( .C1(n15083), .C2(n15074), .A(n15073), .B(n15072), .ZN(
        n15091) );
  AOI22_X1 U16690 ( .A1(n15086), .A2(n10011), .B1(n15091), .B2(n15085), .ZN(
        P3_U3402) );
  INV_X1 U16691 ( .A(P3_REG0_REG_5__SCAN_IN), .ZN(n15324) );
  AOI211_X1 U16692 ( .C1(n15077), .C2(n15083), .A(n15076), .B(n15075), .ZN(
        n15092) );
  AOI22_X1 U16693 ( .A1(n15086), .A2(n15324), .B1(n15092), .B2(n15085), .ZN(
        P3_U3405) );
  AOI211_X1 U16694 ( .C1(n15080), .C2(n15083), .A(n15079), .B(n15078), .ZN(
        n15093) );
  AOI22_X1 U16695 ( .A1(n15086), .A2(n10561), .B1(n15093), .B2(n15085), .ZN(
        P3_U3417) );
  AOI211_X1 U16696 ( .C1(n15084), .C2(n15083), .A(n15082), .B(n15081), .ZN(
        n15095) );
  AOI22_X1 U16697 ( .A1(n15086), .A2(n10569), .B1(n15095), .B2(n15085), .ZN(
        P3_U3420) );
  INV_X1 U16698 ( .A(P3_REG1_REG_1__SCAN_IN), .ZN(n15087) );
  AOI22_X1 U16699 ( .A1(n15096), .A2(n15088), .B1(n15087), .B2(n15094), .ZN(
        P3_U3460) );
  AOI22_X1 U16700 ( .A1(n15096), .A2(n15089), .B1(n10044), .B2(n15094), .ZN(
        P3_U3461) );
  AOI22_X1 U16701 ( .A1(n15096), .A2(n15090), .B1(n10914), .B2(n15094), .ZN(
        P3_U3462) );
  AOI22_X1 U16702 ( .A1(n15096), .A2(n15091), .B1(n10920), .B2(n15094), .ZN(
        P3_U3463) );
  AOI22_X1 U16703 ( .A1(n15096), .A2(n15092), .B1(n10927), .B2(n15094), .ZN(
        P3_U3464) );
  AOI22_X1 U16704 ( .A1(n15096), .A2(n15093), .B1(n10952), .B2(n15094), .ZN(
        P3_U3468) );
  AOI22_X1 U16705 ( .A1(n15096), .A2(n15095), .B1(n10958), .B2(n15094), .ZN(
        P3_U3469) );
  NOR4_X1 U16706 ( .A1(n7353), .A2(P2_DATAO_REG_0__SCAN_IN), .A3(
        P3_IR_REG_30__SCAN_IN), .A4(P3_D_REG_0__SCAN_IN), .ZN(n15097) );
  NAND3_X1 U16707 ( .A1(n15097), .A2(P3_D_REG_15__SCAN_IN), .A3(
        P3_D_REG_6__SCAN_IN), .ZN(n15107) );
  NOR4_X1 U16708 ( .A1(P1_DATAO_REG_25__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .A3(P3_ADDR_REG_4__SCAN_IN), .A4(n15297), .ZN(n15103) );
  NAND4_X1 U16709 ( .A1(P3_IR_REG_15__SCAN_IN), .A2(P3_REG3_REG_7__SCAN_IN), 
        .A3(n9700), .A4(n15216), .ZN(n15101) );
  NAND4_X1 U16710 ( .A1(P3_REG3_REG_10__SCAN_IN), .A2(P3_REG3_REG_9__SCAN_IN), 
        .A3(P1_ADDR_REG_5__SCAN_IN), .A4(P3_ADDR_REG_6__SCAN_IN), .ZN(n15100)
         );
  NAND4_X1 U16711 ( .A1(P3_REG2_REG_5__SCAN_IN), .A2(P3_REG0_REG_5__SCAN_IN), 
        .A3(P3_REG0_REG_1__SCAN_IN), .A4(SI_1_), .ZN(n15099) );
  NAND4_X1 U16712 ( .A1(P1_RD_REG_SCAN_IN), .A2(P3_REG0_REG_9__SCAN_IN), .A3(
        n15278), .A4(n10939), .ZN(n15098) );
  NOR4_X1 U16713 ( .A1(n15101), .A2(n15100), .A3(n15099), .A4(n15098), .ZN(
        n15102) );
  NAND4_X1 U16714 ( .A1(n15105), .A2(n15104), .A3(n15103), .A4(n15102), .ZN(
        n15106) );
  NOR4_X1 U16715 ( .A1(P1_DATAO_REG_11__SCAN_IN), .A2(n9378), .A3(n15107), 
        .A4(n15106), .ZN(n15139) );
  NAND4_X1 U16716 ( .A1(P2_DATAO_REG_27__SCAN_IN), .A2(
        P2_DATAO_REG_20__SCAN_IN), .A3(P1_DATAO_REG_13__SCAN_IN), .A4(SI_31_), 
        .ZN(n15111) );
  NAND4_X1 U16717 ( .A1(P2_REG3_REG_26__SCAN_IN), .A2(P2_REG3_REG_17__SCAN_IN), 
        .A3(P2_REG2_REG_19__SCAN_IN), .A4(P2_REG2_REG_31__SCAN_IN), .ZN(n15110) );
  NAND4_X1 U16718 ( .A1(P2_DATAO_REG_23__SCAN_IN), .A2(P2_REG3_REG_1__SCAN_IN), 
        .A3(P1_REG3_REG_26__SCAN_IN), .A4(P2_ADDR_REG_18__SCAN_IN), .ZN(n15109) );
  NAND4_X1 U16719 ( .A1(P3_REG3_REG_19__SCAN_IN), .A2(P3_REG3_REG_17__SCAN_IN), 
        .A3(SI_27_), .A4(SI_23_), .ZN(n15108) );
  NOR4_X1 U16720 ( .A1(n15111), .A2(n15110), .A3(n15109), .A4(n15108), .ZN(
        n15138) );
  NAND4_X1 U16721 ( .A1(P1_D_REG_28__SCAN_IN), .A2(P1_D_REG_11__SCAN_IN), .A3(
        P1_REG0_REG_20__SCAN_IN), .A4(P1_REG2_REG_8__SCAN_IN), .ZN(n15115) );
  NAND4_X1 U16722 ( .A1(P1_D_REG_18__SCAN_IN), .A2(P1_REG1_REG_25__SCAN_IN), 
        .A3(P1_REG1_REG_22__SCAN_IN), .A4(P1_REG0_REG_19__SCAN_IN), .ZN(n15114) );
  NAND4_X1 U16723 ( .A1(P2_REG2_REG_16__SCAN_IN), .A2(P1_REG3_REG_22__SCAN_IN), 
        .A3(P1_REG3_REG_19__SCAN_IN), .A4(P1_REG1_REG_15__SCAN_IN), .ZN(n15113) );
  NAND4_X1 U16724 ( .A1(P2_DATAO_REG_24__SCAN_IN), .A2(P1_REG1_REG_18__SCAN_IN), .A3(P1_REG1_REG_14__SCAN_IN), .A4(P1_REG0_REG_12__SCAN_IN), .ZN(n15112) );
  NOR4_X1 U16725 ( .A1(n15115), .A2(n15114), .A3(n15113), .A4(n15112), .ZN(
        n15137) );
  NOR4_X1 U16726 ( .A1(P1_IR_REG_29__SCAN_IN), .A2(P1_REG2_REG_25__SCAN_IN), 
        .A3(P1_REG0_REG_21__SCAN_IN), .A4(P1_REG0_REG_30__SCAN_IN), .ZN(n15119) );
  NOR4_X1 U16727 ( .A1(n15206), .A2(P2_REG2_REG_10__SCAN_IN), .A3(
        P2_REG3_REG_2__SCAN_IN), .A4(P1_IR_REG_24__SCAN_IN), .ZN(n15118) );
  NOR4_X1 U16728 ( .A1(SI_19_), .A2(P1_REG2_REG_12__SCAN_IN), .A3(
        P2_ADDR_REG_8__SCAN_IN), .A4(P2_ADDR_REG_12__SCAN_IN), .ZN(n15117) );
  NOR4_X1 U16729 ( .A1(P1_IR_REG_2__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .A3(
        P1_REG0_REG_5__SCAN_IN), .A4(P1_REG2_REG_2__SCAN_IN), .ZN(n15116) );
  NAND4_X1 U16730 ( .A1(n15119), .A2(n15118), .A3(n15117), .A4(n15116), .ZN(
        n15135) );
  NOR4_X1 U16731 ( .A1(P2_REG3_REG_27__SCAN_IN), .A2(P1_IR_REG_8__SCAN_IN), 
        .A3(P1_IR_REG_5__SCAN_IN), .A4(P3_DATAO_REG_21__SCAN_IN), .ZN(n15123)
         );
  NOR4_X1 U16732 ( .A1(P1_DATAO_REG_16__SCAN_IN), .A2(P3_REG2_REG_0__SCAN_IN), 
        .A3(P3_DATAO_REG_23__SCAN_IN), .A4(n15296), .ZN(n15122) );
  NOR4_X1 U16733 ( .A1(SI_12_), .A2(P2_REG1_REG_6__SCAN_IN), .A3(
        P2_REG2_REG_7__SCAN_IN), .A4(P2_REG0_REG_7__SCAN_IN), .ZN(n15121) );
  NOR4_X1 U16734 ( .A1(P2_D_REG_10__SCAN_IN), .A2(P2_REG1_REG_22__SCAN_IN), 
        .A3(P2_REG0_REG_21__SCAN_IN), .A4(P2_REG0_REG_25__SCAN_IN), .ZN(n15120) );
  NAND4_X1 U16735 ( .A1(n15123), .A2(n15122), .A3(n15121), .A4(n15120), .ZN(
        n15134) );
  NAND4_X1 U16736 ( .A1(P2_REG1_REG_28__SCAN_IN), .A2(P2_REG0_REG_28__SCAN_IN), 
        .A3(P1_D_REG_0__SCAN_IN), .A4(P1_REG0_REG_1__SCAN_IN), .ZN(n15127) );
  NAND4_X1 U16737 ( .A1(P1_IR_REG_23__SCAN_IN), .A2(P3_DATAO_REG_19__SCAN_IN), 
        .A3(P3_DATAO_REG_31__SCAN_IN), .A4(P3_DATAO_REG_2__SCAN_IN), .ZN(
        n15126) );
  NAND4_X1 U16738 ( .A1(P2_REG2_REG_1__SCAN_IN), .A2(P2_REG1_REG_7__SCAN_IN), 
        .A3(P1_REG1_REG_29__SCAN_IN), .A4(P1_REG1_REG_30__SCAN_IN), .ZN(n15125) );
  NAND4_X1 U16739 ( .A1(P2_D_REG_18__SCAN_IN), .A2(P2_D_REG_7__SCAN_IN), .A3(
        P2_REG0_REG_19__SCAN_IN), .A4(P2_REG0_REG_12__SCAN_IN), .ZN(n15124) );
  OR4_X1 U16740 ( .A1(n15127), .A2(n15126), .A3(n15125), .A4(n15124), .ZN(
        n15133) );
  NOR4_X1 U16741 ( .A1(P2_DATAO_REG_31__SCAN_IN), .A2(P1_DATAO_REG_15__SCAN_IN), .A3(P2_REG3_REG_25__SCAN_IN), .A4(P2_REG2_REG_24__SCAN_IN), .ZN(n15131) );
  NOR4_X1 U16742 ( .A1(P2_REG2_REG_22__SCAN_IN), .A2(P2_REG1_REG_18__SCAN_IN), 
        .A3(P2_REG1_REG_16__SCAN_IN), .A4(P1_REG2_REG_30__SCAN_IN), .ZN(n15130) );
  NOR4_X1 U16743 ( .A1(n15257), .A2(n15198), .A3(n15310), .A4(
        P3_WR_REG_SCAN_IN), .ZN(n15129) );
  NOR4_X1 U16744 ( .A1(P3_REG1_REG_23__SCAN_IN), .A2(P3_REG2_REG_21__SCAN_IN), 
        .A3(P3_REG0_REG_18__SCAN_IN), .A4(P3_ADDR_REG_18__SCAN_IN), .ZN(n15128) );
  NAND4_X1 U16745 ( .A1(n15131), .A2(n15130), .A3(n15129), .A4(n15128), .ZN(
        n15132) );
  NOR4_X1 U16746 ( .A1(n15135), .A2(n15134), .A3(n15133), .A4(n15132), .ZN(
        n15136) );
  NAND4_X1 U16747 ( .A1(n15139), .A2(n15138), .A3(n15137), .A4(n15136), .ZN(
        n15406) );
  AOI22_X1 U16748 ( .A1(n9330), .A2(keyinput30), .B1(n10939), .B2(keyinput7), 
        .ZN(n15140) );
  OAI221_X1 U16749 ( .B1(n9330), .B2(keyinput30), .C1(n10939), .C2(keyinput7), 
        .A(n15140), .ZN(n15152) );
  INV_X1 U16750 ( .A(P1_REG2_REG_30__SCAN_IN), .ZN(n15143) );
  AOI22_X1 U16751 ( .A1(n15143), .A2(keyinput0), .B1(keyinput123), .B2(n15142), 
        .ZN(n15141) );
  OAI221_X1 U16752 ( .B1(n15143), .B2(keyinput0), .C1(n15142), .C2(keyinput123), .A(n15141), .ZN(n15151) );
  AOI22_X1 U16753 ( .A1(n15146), .A2(keyinput112), .B1(n15145), .B2(keyinput44), .ZN(n15144) );
  OAI221_X1 U16754 ( .B1(n15146), .B2(keyinput112), .C1(n15145), .C2(
        keyinput44), .A(n15144), .ZN(n15150) );
  AOI22_X1 U16755 ( .A1(n7578), .A2(keyinput98), .B1(n15148), .B2(keyinput105), 
        .ZN(n15147) );
  OAI221_X1 U16756 ( .B1(n7578), .B2(keyinput98), .C1(n15148), .C2(keyinput105), .A(n15147), .ZN(n15149) );
  NOR4_X1 U16757 ( .A1(n15152), .A2(n15151), .A3(n15150), .A4(n15149), .ZN(
        n15196) );
  AOI22_X1 U16758 ( .A1(n7797), .A2(keyinput17), .B1(n15154), .B2(keyinput59), 
        .ZN(n15153) );
  OAI221_X1 U16759 ( .B1(n7797), .B2(keyinput17), .C1(n15154), .C2(keyinput59), 
        .A(n15153), .ZN(n15165) );
  AOI22_X1 U16760 ( .A1(n15157), .A2(keyinput36), .B1(keyinput61), .B2(n15156), 
        .ZN(n15155) );
  OAI221_X1 U16761 ( .B1(n15157), .B2(keyinput36), .C1(n15156), .C2(keyinput61), .A(n15155), .ZN(n15164) );
  AOI22_X1 U16762 ( .A1(n15160), .A2(keyinput104), .B1(keyinput122), .B2(
        n15159), .ZN(n15158) );
  OAI221_X1 U16763 ( .B1(n15160), .B2(keyinput104), .C1(n15159), .C2(
        keyinput122), .A(n15158), .ZN(n15163) );
  AOI22_X1 U16764 ( .A1(n10561), .A2(keyinput21), .B1(keyinput64), .B2(n10182), 
        .ZN(n15161) );
  OAI221_X1 U16765 ( .B1(n10561), .B2(keyinput21), .C1(n10182), .C2(keyinput64), .A(n15161), .ZN(n15162) );
  NOR4_X1 U16766 ( .A1(n15165), .A2(n15164), .A3(n15163), .A4(n15162), .ZN(
        n15195) );
  AOI22_X1 U16767 ( .A1(n15167), .A2(keyinput62), .B1(keyinput60), .B2(n8198), 
        .ZN(n15166) );
  OAI221_X1 U16768 ( .B1(n15167), .B2(keyinput62), .C1(n8198), .C2(keyinput60), 
        .A(n15166), .ZN(n15178) );
  AOI22_X1 U16769 ( .A1(n11409), .A2(keyinput93), .B1(n12877), .B2(keyinput37), 
        .ZN(n15168) );
  OAI221_X1 U16770 ( .B1(n11409), .B2(keyinput93), .C1(n12877), .C2(keyinput37), .A(n15168), .ZN(n15177) );
  AOI22_X1 U16771 ( .A1(n15171), .A2(keyinput72), .B1(n15170), .B2(keyinput73), 
        .ZN(n15169) );
  OAI221_X1 U16772 ( .B1(n15171), .B2(keyinput72), .C1(n15170), .C2(keyinput73), .A(n15169), .ZN(n15176) );
  AOI22_X1 U16773 ( .A1(n15174), .A2(keyinput78), .B1(keyinput40), .B2(n15173), 
        .ZN(n15172) );
  OAI221_X1 U16774 ( .B1(n15174), .B2(keyinput78), .C1(n15173), .C2(keyinput40), .A(n15172), .ZN(n15175) );
  NOR4_X1 U16775 ( .A1(n15178), .A2(n15177), .A3(n15176), .A4(n15175), .ZN(
        n15194) );
  AOI22_X1 U16776 ( .A1(n15181), .A2(keyinput46), .B1(keyinput39), .B2(n15180), 
        .ZN(n15179) );
  OAI221_X1 U16777 ( .B1(n15181), .B2(keyinput46), .C1(n15180), .C2(keyinput39), .A(n15179), .ZN(n15192) );
  AOI22_X1 U16778 ( .A1(n10865), .A2(keyinput103), .B1(n9333), .B2(keyinput102), .ZN(n15182) );
  OAI221_X1 U16779 ( .B1(n10865), .B2(keyinput103), .C1(n9333), .C2(
        keyinput102), .A(n15182), .ZN(n15191) );
  AOI22_X1 U16780 ( .A1(n15185), .A2(keyinput27), .B1(n15184), .B2(keyinput25), 
        .ZN(n15183) );
  OAI221_X1 U16781 ( .B1(n15185), .B2(keyinput27), .C1(n15184), .C2(keyinput25), .A(n15183), .ZN(n15190) );
  AOI22_X1 U16782 ( .A1(n15188), .A2(keyinput53), .B1(keyinput29), .B2(n15187), 
        .ZN(n15186) );
  OAI221_X1 U16783 ( .B1(n15188), .B2(keyinput53), .C1(n15187), .C2(keyinput29), .A(n15186), .ZN(n15189) );
  NOR4_X1 U16784 ( .A1(n15192), .A2(n15191), .A3(n15190), .A4(n15189), .ZN(
        n15193) );
  NAND4_X1 U16785 ( .A1(n15196), .A2(n15195), .A3(n15194), .A4(n15193), .ZN(
        n15384) );
  AOI22_X1 U16786 ( .A1(n15199), .A2(keyinput70), .B1(keyinput81), .B2(n15198), 
        .ZN(n15197) );
  OAI221_X1 U16787 ( .B1(n15199), .B2(keyinput70), .C1(n15198), .C2(keyinput81), .A(n15197), .ZN(n15212) );
  AOI22_X1 U16788 ( .A1(n15202), .A2(keyinput14), .B1(keyinput16), .B2(n15201), 
        .ZN(n15200) );
  OAI221_X1 U16789 ( .B1(n15202), .B2(keyinput14), .C1(n15201), .C2(keyinput16), .A(n15200), .ZN(n15211) );
  AOI22_X1 U16790 ( .A1(n15205), .A2(keyinput118), .B1(n15204), .B2(keyinput26), .ZN(n15203) );
  OAI221_X1 U16791 ( .B1(n15205), .B2(keyinput118), .C1(n15204), .C2(
        keyinput26), .A(n15203), .ZN(n15210) );
  XNOR2_X1 U16792 ( .A(n15206), .B(keyinput69), .ZN(n15208) );
  XNOR2_X1 U16793 ( .A(P1_IR_REG_5__SCAN_IN), .B(keyinput89), .ZN(n15207) );
  NAND2_X1 U16794 ( .A1(n15208), .A2(n15207), .ZN(n15209) );
  NOR4_X1 U16795 ( .A1(n15212), .A2(n15211), .A3(n15210), .A4(n15209), .ZN(
        n15254) );
  AOI22_X1 U16796 ( .A1(n10425), .A2(keyinput45), .B1(n15214), .B2(keyinput2), 
        .ZN(n15213) );
  OAI221_X1 U16797 ( .B1(n10425), .B2(keyinput45), .C1(n15214), .C2(keyinput2), 
        .A(n15213), .ZN(n15225) );
  AOI22_X1 U16798 ( .A1(n15217), .A2(keyinput56), .B1(keyinput71), .B2(n15216), 
        .ZN(n15215) );
  OAI221_X1 U16799 ( .B1(n15217), .B2(keyinput56), .C1(n15216), .C2(keyinput71), .A(n15215), .ZN(n15224) );
  INV_X1 U16800 ( .A(P3_WR_REG_SCAN_IN), .ZN(n15219) );
  AOI22_X1 U16801 ( .A1(n15219), .A2(keyinput106), .B1(n9700), .B2(keyinput48), 
        .ZN(n15218) );
  OAI221_X1 U16802 ( .B1(n15219), .B2(keyinput106), .C1(n9700), .C2(keyinput48), .A(n15218), .ZN(n15223) );
  AOI22_X1 U16803 ( .A1(n7368), .A2(keyinput125), .B1(keyinput20), .B2(n15221), 
        .ZN(n15220) );
  OAI221_X1 U16804 ( .B1(n7368), .B2(keyinput125), .C1(n15221), .C2(keyinput20), .A(n15220), .ZN(n15222) );
  NOR4_X1 U16805 ( .A1(n15225), .A2(n15224), .A3(n15223), .A4(n15222), .ZN(
        n15253) );
  AOI22_X1 U16806 ( .A1(n15227), .A2(keyinput33), .B1(keyinput109), .B2(n8309), 
        .ZN(n15226) );
  OAI221_X1 U16807 ( .B1(n15227), .B2(keyinput33), .C1(n8309), .C2(keyinput109), .A(n15226), .ZN(n15240) );
  AOI22_X1 U16808 ( .A1(n15230), .A2(keyinput47), .B1(n15229), .B2(keyinput127), .ZN(n15228) );
  OAI221_X1 U16809 ( .B1(n15230), .B2(keyinput47), .C1(n15229), .C2(
        keyinput127), .A(n15228), .ZN(n15239) );
  AOI22_X1 U16810 ( .A1(n15233), .A2(keyinput41), .B1(keyinput94), .B2(n15232), 
        .ZN(n15231) );
  OAI221_X1 U16811 ( .B1(n15233), .B2(keyinput41), .C1(n15232), .C2(keyinput94), .A(n15231), .ZN(n15238) );
  AOI22_X1 U16812 ( .A1(n15236), .A2(keyinput1), .B1(keyinput113), .B2(n15235), 
        .ZN(n15234) );
  OAI221_X1 U16813 ( .B1(n15236), .B2(keyinput1), .C1(n15235), .C2(keyinput113), .A(n15234), .ZN(n15237) );
  NOR4_X1 U16814 ( .A1(n15240), .A2(n15239), .A3(n15238), .A4(n15237), .ZN(
        n15252) );
  AOI22_X1 U16815 ( .A1(n10364), .A2(keyinput110), .B1(keyinput107), .B2(
        n15242), .ZN(n15241) );
  OAI221_X1 U16816 ( .B1(n10364), .B2(keyinput110), .C1(n15242), .C2(
        keyinput107), .A(n15241), .ZN(n15250) );
  AOI22_X1 U16817 ( .A1(n10928), .A2(keyinput86), .B1(n10557), .B2(keyinput101), .ZN(n15243) );
  OAI221_X1 U16818 ( .B1(n10928), .B2(keyinput86), .C1(n10557), .C2(
        keyinput101), .A(n15243), .ZN(n15249) );
  XNOR2_X1 U16819 ( .A(P2_REG1_REG_18__SCAN_IN), .B(keyinput19), .ZN(n15247)
         );
  XNOR2_X1 U16820 ( .A(P3_IR_REG_15__SCAN_IN), .B(keyinput83), .ZN(n15246) );
  XNOR2_X1 U16821 ( .A(P2_REG0_REG_25__SCAN_IN), .B(keyinput121), .ZN(n15245)
         );
  XNOR2_X1 U16822 ( .A(P1_IR_REG_24__SCAN_IN), .B(keyinput68), .ZN(n15244) );
  NAND4_X1 U16823 ( .A1(n15247), .A2(n15246), .A3(n15245), .A4(n15244), .ZN(
        n15248) );
  NOR3_X1 U16824 ( .A1(n15250), .A2(n15249), .A3(n15248), .ZN(n15251) );
  NAND4_X1 U16825 ( .A1(n15254), .A2(n15253), .A3(n15252), .A4(n15251), .ZN(
        n15383) );
  INV_X1 U16826 ( .A(P1_REG2_REG_25__SCAN_IN), .ZN(n15256) );
  AOI22_X1 U16827 ( .A1(n15257), .A2(keyinput65), .B1(n15256), .B2(keyinput92), 
        .ZN(n15255) );
  OAI221_X1 U16828 ( .B1(n15257), .B2(keyinput65), .C1(n15256), .C2(keyinput92), .A(n15255), .ZN(n15269) );
  AOI22_X1 U16829 ( .A1(n15260), .A2(keyinput9), .B1(keyinput13), .B2(n15259), 
        .ZN(n15258) );
  OAI221_X1 U16830 ( .B1(n15260), .B2(keyinput9), .C1(n15259), .C2(keyinput13), 
        .A(n15258), .ZN(n15268) );
  AOI22_X1 U16831 ( .A1(n15263), .A2(keyinput42), .B1(keyinput116), .B2(n15262), .ZN(n15261) );
  OAI221_X1 U16832 ( .B1(n15263), .B2(keyinput42), .C1(n15262), .C2(
        keyinput116), .A(n15261), .ZN(n15267) );
  AOI22_X1 U16833 ( .A1(n15265), .A2(keyinput49), .B1(keyinput35), .B2(n7707), 
        .ZN(n15264) );
  OAI221_X1 U16834 ( .B1(n15265), .B2(keyinput49), .C1(n7707), .C2(keyinput35), 
        .A(n15264), .ZN(n15266) );
  NOR4_X1 U16835 ( .A1(n15269), .A2(n15268), .A3(n15267), .A4(n15266), .ZN(
        n15319) );
  AOI22_X1 U16836 ( .A1(n15272), .A2(keyinput34), .B1(keyinput79), .B2(n15271), 
        .ZN(n15270) );
  OAI221_X1 U16837 ( .B1(n15272), .B2(keyinput34), .C1(n15271), .C2(keyinput79), .A(n15270), .ZN(n15285) );
  AOI22_X1 U16838 ( .A1(n15275), .A2(keyinput114), .B1(keyinput124), .B2(
        n15274), .ZN(n15273) );
  OAI221_X1 U16839 ( .B1(n15275), .B2(keyinput114), .C1(n15274), .C2(
        keyinput124), .A(n15273), .ZN(n15284) );
  AOI22_X1 U16840 ( .A1(n15278), .A2(keyinput11), .B1(keyinput82), .B2(n15277), 
        .ZN(n15276) );
  OAI221_X1 U16841 ( .B1(n15278), .B2(keyinput11), .C1(n15277), .C2(keyinput82), .A(n15276), .ZN(n15283) );
  AOI22_X1 U16842 ( .A1(n15281), .A2(keyinput74), .B1(n15280), .B2(keyinput8), 
        .ZN(n15279) );
  OAI221_X1 U16843 ( .B1(n15281), .B2(keyinput74), .C1(n15280), .C2(keyinput8), 
        .A(n15279), .ZN(n15282) );
  NOR4_X1 U16844 ( .A1(n15285), .A2(n15284), .A3(n15283), .A4(n15282), .ZN(
        n15318) );
  INV_X1 U16845 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n15287) );
  AOI22_X1 U16846 ( .A1(n15288), .A2(keyinput5), .B1(keyinput54), .B2(n15287), 
        .ZN(n15286) );
  OAI221_X1 U16847 ( .B1(n15288), .B2(keyinput5), .C1(n15287), .C2(keyinput54), 
        .A(n15286), .ZN(n15301) );
  AOI22_X1 U16848 ( .A1(n15291), .A2(keyinput15), .B1(keyinput75), .B2(n15290), 
        .ZN(n15289) );
  OAI221_X1 U16849 ( .B1(n15291), .B2(keyinput15), .C1(n15290), .C2(keyinput75), .A(n15289), .ZN(n15300) );
  AOI22_X1 U16850 ( .A1(n15294), .A2(keyinput18), .B1(n15293), .B2(keyinput80), 
        .ZN(n15292) );
  OAI221_X1 U16851 ( .B1(n15294), .B2(keyinput18), .C1(n15293), .C2(keyinput80), .A(n15292), .ZN(n15299) );
  AOI22_X1 U16852 ( .A1(n15297), .A2(keyinput91), .B1(keyinput10), .B2(n15296), 
        .ZN(n15295) );
  OAI221_X1 U16853 ( .B1(n15297), .B2(keyinput91), .C1(n15296), .C2(keyinput10), .A(n15295), .ZN(n15298) );
  NOR4_X1 U16854 ( .A1(n15301), .A2(n15300), .A3(n15299), .A4(n15298), .ZN(
        n15317) );
  AOI22_X1 U16855 ( .A1(n15303), .A2(keyinput96), .B1(n12606), .B2(keyinput66), 
        .ZN(n15302) );
  OAI221_X1 U16856 ( .B1(n15303), .B2(keyinput96), .C1(n12606), .C2(keyinput66), .A(n15302), .ZN(n15307) );
  XNOR2_X1 U16857 ( .A(n15304), .B(keyinput108), .ZN(n15306) );
  XNOR2_X1 U16858 ( .A(n7040), .B(keyinput50), .ZN(n15305) );
  OR3_X1 U16859 ( .A1(n15307), .A2(n15306), .A3(n15305), .ZN(n15315) );
  AOI22_X1 U16860 ( .A1(n15310), .A2(keyinput22), .B1(n15309), .B2(keyinput4), 
        .ZN(n15308) );
  OAI221_X1 U16861 ( .B1(n15310), .B2(keyinput22), .C1(n15309), .C2(keyinput4), 
        .A(n15308), .ZN(n15314) );
  AOI22_X1 U16862 ( .A1(n15312), .A2(keyinput12), .B1(keyinput120), .B2(n7979), 
        .ZN(n15311) );
  OAI221_X1 U16863 ( .B1(n15312), .B2(keyinput12), .C1(n7979), .C2(keyinput120), .A(n15311), .ZN(n15313) );
  NOR3_X1 U16864 ( .A1(n15315), .A2(n15314), .A3(n15313), .ZN(n15316) );
  NAND4_X1 U16865 ( .A1(n15319), .A2(n15318), .A3(n15317), .A4(n15316), .ZN(
        n15382) );
  INV_X1 U16866 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n15321) );
  AOI22_X1 U16867 ( .A1(n15322), .A2(keyinput28), .B1(keyinput55), .B2(n15321), 
        .ZN(n15320) );
  OAI221_X1 U16868 ( .B1(n15322), .B2(keyinput28), .C1(n15321), .C2(keyinput55), .A(n15320), .ZN(n15334) );
  AOI22_X1 U16869 ( .A1(n15325), .A2(keyinput6), .B1(keyinput32), .B2(n15324), 
        .ZN(n15323) );
  OAI221_X1 U16870 ( .B1(n15325), .B2(keyinput6), .C1(n15324), .C2(keyinput32), 
        .A(n15323), .ZN(n15333) );
  AOI22_X1 U16871 ( .A1(n8321), .A2(keyinput111), .B1(keyinput43), .B2(n15327), 
        .ZN(n15326) );
  OAI221_X1 U16872 ( .B1(n8321), .B2(keyinput111), .C1(n15327), .C2(keyinput43), .A(n15326), .ZN(n15332) );
  AOI22_X1 U16873 ( .A1(n15330), .A2(keyinput58), .B1(keyinput38), .B2(n15329), 
        .ZN(n15328) );
  OAI221_X1 U16874 ( .B1(n15330), .B2(keyinput58), .C1(n15329), .C2(keyinput38), .A(n15328), .ZN(n15331) );
  NOR4_X1 U16875 ( .A1(n15334), .A2(n15333), .A3(n15332), .A4(n15331), .ZN(
        n15380) );
  AOI22_X1 U16876 ( .A1(n15337), .A2(keyinput100), .B1(keyinput31), .B2(n15336), .ZN(n15335) );
  OAI221_X1 U16877 ( .B1(n15337), .B2(keyinput100), .C1(n15336), .C2(
        keyinput31), .A(n15335), .ZN(n15340) );
  XNOR2_X1 U16878 ( .A(n15338), .B(keyinput3), .ZN(n15339) );
  NOR2_X1 U16879 ( .A1(n15340), .A2(n15339), .ZN(n15351) );
  INV_X1 U16880 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n15342) );
  AOI22_X1 U16881 ( .A1(n13312), .A2(keyinput115), .B1(keyinput23), .B2(n15342), .ZN(n15341) );
  OAI221_X1 U16882 ( .B1(n13312), .B2(keyinput115), .C1(n15342), .C2(
        keyinput23), .A(n15341), .ZN(n15343) );
  INV_X1 U16883 ( .A(n15343), .ZN(n15350) );
  AOI22_X1 U16884 ( .A1(n15346), .A2(keyinput119), .B1(n15345), .B2(keyinput76), .ZN(n15344) );
  OAI221_X1 U16885 ( .B1(n15346), .B2(keyinput119), .C1(n15345), .C2(
        keyinput76), .A(n15344), .ZN(n15347) );
  INV_X1 U16886 ( .A(n15347), .ZN(n15349) );
  XNOR2_X1 U16887 ( .A(P1_IR_REG_8__SCAN_IN), .B(keyinput87), .ZN(n15348) );
  AND4_X1 U16888 ( .A1(n15351), .A2(n15350), .A3(n15349), .A4(n15348), .ZN(
        n15379) );
  AOI22_X1 U16889 ( .A1(n15353), .A2(keyinput95), .B1(keyinput77), .B2(n8554), 
        .ZN(n15352) );
  OAI221_X1 U16890 ( .B1(n15353), .B2(keyinput95), .C1(n8554), .C2(keyinput77), 
        .A(n15352), .ZN(n15363) );
  INV_X1 U16891 ( .A(P1_RD_REG_SCAN_IN), .ZN(n15356) );
  AOI22_X1 U16892 ( .A1(n15356), .A2(keyinput99), .B1(keyinput84), .B2(n15355), 
        .ZN(n15354) );
  OAI221_X1 U16893 ( .B1(n15356), .B2(keyinput99), .C1(n15355), .C2(keyinput84), .A(n15354), .ZN(n15362) );
  XOR2_X1 U16894 ( .A(n9378), .B(keyinput63), .Z(n15360) );
  XNOR2_X1 U16895 ( .A(P2_REG0_REG_19__SCAN_IN), .B(keyinput85), .ZN(n15359)
         );
  XNOR2_X1 U16896 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(keyinput51), .ZN(n15358)
         );
  XNOR2_X1 U16897 ( .A(P1_IR_REG_23__SCAN_IN), .B(keyinput97), .ZN(n15357) );
  NAND4_X1 U16898 ( .A1(n15360), .A2(n15359), .A3(n15358), .A4(n15357), .ZN(
        n15361) );
  NOR3_X1 U16899 ( .A1(n15363), .A2(n15362), .A3(n15361), .ZN(n15378) );
  AOI22_X1 U16900 ( .A1(n15365), .A2(keyinput52), .B1(n12878), .B2(keyinput88), 
        .ZN(n15364) );
  OAI221_X1 U16901 ( .B1(n15365), .B2(keyinput52), .C1(n12878), .C2(keyinput88), .A(n15364), .ZN(n15376) );
  AOI22_X1 U16902 ( .A1(n15367), .A2(keyinput117), .B1(keyinput67), .B2(n13260), .ZN(n15366) );
  OAI221_X1 U16903 ( .B1(n15367), .B2(keyinput117), .C1(n13260), .C2(
        keyinput67), .A(n15366), .ZN(n15375) );
  AOI22_X1 U16904 ( .A1(n15370), .A2(keyinput24), .B1(n15369), .B2(keyinput90), 
        .ZN(n15368) );
  OAI221_X1 U16905 ( .B1(n15370), .B2(keyinput24), .C1(n15369), .C2(keyinput90), .A(n15368), .ZN(n15374) );
  AOI22_X1 U16906 ( .A1(n15372), .A2(keyinput126), .B1(n9737), .B2(keyinput57), 
        .ZN(n15371) );
  OAI221_X1 U16907 ( .B1(n15372), .B2(keyinput126), .C1(n9737), .C2(keyinput57), .A(n15371), .ZN(n15373) );
  NOR4_X1 U16908 ( .A1(n15376), .A2(n15375), .A3(n15374), .A4(n15373), .ZN(
        n15377) );
  NAND4_X1 U16909 ( .A1(n15380), .A2(n15379), .A3(n15378), .A4(n15377), .ZN(
        n15381) );
  NOR4_X1 U16910 ( .A1(n15384), .A2(n15383), .A3(n15382), .A4(n15381), .ZN(
        n15404) );
  AOI21_X1 U16911 ( .B1(n15387), .B2(n15386), .A(n15385), .ZN(n15402) );
  NAND2_X1 U16912 ( .A1(n15389), .A2(n15388), .ZN(n15391) );
  OAI211_X1 U16913 ( .C1(n15393), .C2(n15392), .A(n15391), .B(n15390), .ZN(
        n15397) );
  NOR2_X1 U16914 ( .A1(n15395), .A2(n15394), .ZN(n15396) );
  AOI211_X1 U16915 ( .C1(n15399), .C2(n15398), .A(n15397), .B(n15396), .ZN(
        n15400) );
  OAI21_X1 U16916 ( .B1(n15402), .B2(n15401), .A(n15400), .ZN(n15403) );
  XOR2_X1 U16917 ( .A(n15404), .B(n15403), .Z(n15405) );
  XNOR2_X1 U16918 ( .A(n15406), .B(n15405), .ZN(P3_U3176) );
  OAI21_X1 U16919 ( .B1(n15409), .B2(n15408), .A(n15407), .ZN(SUB_1596_U59) );
  OAI21_X1 U16920 ( .B1(n15412), .B2(n15411), .A(n15410), .ZN(SUB_1596_U58) );
  XOR2_X1 U16921 ( .A(P2_ADDR_REG_0__SCAN_IN), .B(n15413), .Z(SUB_1596_U53) );
  AOI21_X1 U16922 ( .B1(n15416), .B2(n15415), .A(n15414), .ZN(SUB_1596_U56) );
  OAI21_X1 U16923 ( .B1(n15419), .B2(n15418), .A(n15417), .ZN(SUB_1596_U60) );
  AOI21_X1 U16924 ( .B1(n15422), .B2(n15421), .A(n15420), .ZN(SUB_1596_U5) );
  BUF_X1 U7355 ( .A(n11946), .Z(n6524) );
  CLKBUF_X1 U7367 ( .A(n12915), .Z(n6540) );
  CLKBUF_X1 U7378 ( .A(n9738), .Z(n11438) );
  CLKBUF_X2 U7628 ( .A(n9740), .Z(n6530) );
  NAND2_X2 U9187 ( .A1(n7793), .A2(n7792), .ZN(n14379) );
endmodule

