

module b21_C_2inp_gates_syn ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, 
        P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, 
        P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, 
        P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, 
        P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, 
        P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, 
        P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, 
        P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, 
        P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, 
        P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, 
        P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, 
        P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, 
        P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, 
        P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, 
        P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, 
        P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, 
        P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, 
        P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, 
        P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, 
        P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, 
        P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, 
        P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, 
        P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, 
        P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, 
        P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, 
        ADD_1071_U57, ADD_1071_U58, ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, 
        ADD_1071_U62, ADD_1071_U63, ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, 
        ADD_1071_U50, ADD_1071_U51, ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, 
        ADD_1071_U5, ADD_1071_U46, U126, U123, P1_U3353, P1_U3352, P1_U3351, 
        P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, 
        P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, 
        P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, 
        P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, 
        P1_U3322, P1_U3440, P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, 
        P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, 
        P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, 
        P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, 
        P1_U3296, P1_U3295, P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, 
        P1_U3460, P1_U3463, P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, 
        P1_U3481, P1_U3484, P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, 
        P1_U3502, P1_U3505, P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, 
        P1_U3514, P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, 
        P1_U3521, P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, 
        P1_U3528, P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, 
        P1_U3535, P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, 
        P1_U3542, P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, 
        P1_U3549, P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, 
        P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, 
        P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, 
        P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, 
        P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, 
        P1_U3355, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, 
        P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, 
        P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, 
        P1_U3242, P1_U3241, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, 
        P1_U3560, P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, 
        P1_U3567, P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, 
        P1_U3574, P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, 
        P1_U3581, P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, 
        P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, 
        P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, 
        P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, 
        P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, 
        P1_U3211, P1_U3084, P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, 
        P2_U3355, P2_U3354, P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, 
        P2_U3348, P2_U3347, P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, 
        P2_U3341, P2_U3340, P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, 
        P2_U3334, P2_U3333, P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, 
        P2_U3327, P2_U3437, P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, 
        P2_U3322, P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, 
        P2_U3315, P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, 
        P2_U3308, P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, 
        P2_U3301, P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, 
        P2_U3457, P2_U3460, P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, 
        P2_U3478, P2_U3481, P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, 
        P2_U3499, P2_U3502, P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, 
        P2_U3511, P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, 
        P2_U3518, P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, 
        P2_U3525, P2_U3526, P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, 
        P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, 
        P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, 
        P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, 
        P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, 
        P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, 
        P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, 
        P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, 
        P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, 
        P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, 
        P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, 
        P2_U3246, P2_U3245, P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, 
        P2_U3557, P2_U3558, P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, 
        P2_U3564, P2_U3565, P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, 
        P2_U3571, P2_U3572, P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, 
        P2_U3578, P2_U3579, P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, 
        P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, 
        P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, 
        P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, 
        P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, 
        P2_U3215, P2_U3152, P2_U3151, P2_U3966, keyinput63, keyinput62, 
        keyinput61, keyinput60, keyinput59, keyinput58, keyinput57, keyinput56, 
        keyinput55, keyinput54, keyinput53, keyinput52, keyinput51, keyinput50, 
        keyinput49, keyinput48, keyinput47, keyinput46, keyinput45, keyinput44, 
        keyinput43, keyinput42, keyinput41, keyinput40, keyinput39, keyinput38, 
        keyinput37, keyinput36, keyinput35, keyinput34, keyinput33, keyinput32, 
        keyinput31, keyinput30, keyinput29, keyinput28, keyinput27, keyinput26, 
        keyinput25, keyinput24, keyinput23, keyinput22, keyinput21, keyinput20, 
        keyinput19, keyinput18, keyinput17, keyinput16, keyinput15, keyinput14, 
        keyinput13, keyinput12, keyinput11, keyinput10, keyinput9, keyinput8, 
        keyinput7, keyinput6, keyinput5, keyinput4, keyinput3, keyinput2, 
        keyinput1, keyinput0 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN,
         P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN,
         P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN,
         P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN,
         P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN,
         P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN,
         P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN,
         P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN,
         P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN,
         P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN,
         P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN,
         P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN,
         P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN,
         P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN,
         P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN,
         P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN,
         P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN,
         P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN,
         P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN,
         P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN,
         P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN,
         P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, keyinput63, keyinput62, keyinput61,
         keyinput60, keyinput59, keyinput58, keyinput57, keyinput56,
         keyinput55, keyinput54, keyinput53, keyinput52, keyinput51,
         keyinput50, keyinput49, keyinput48, keyinput47, keyinput46,
         keyinput45, keyinput44, keyinput43, keyinput42, keyinput41,
         keyinput40, keyinput39, keyinput38, keyinput37, keyinput36,
         keyinput35, keyinput34, keyinput33, keyinput32, keyinput31,
         keyinput30, keyinput29, keyinput28, keyinput27, keyinput26,
         keyinput25, keyinput24, keyinput23, keyinput22, keyinput21,
         keyinput20, keyinput19, keyinput18, keyinput17, keyinput16,
         keyinput15, keyinput14, keyinput13, keyinput12, keyinput11,
         keyinput10, keyinput9, keyinput8, keyinput7, keyinput6, keyinput5,
         keyinput4, keyinput3, keyinput2, keyinput1, keyinput0;
  output ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, ADD_1071_U57, ADD_1071_U58,
         ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, ADD_1071_U62, ADD_1071_U63,
         ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, ADD_1071_U50, ADD_1071_U51,
         ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, ADD_1071_U5, ADD_1071_U46,
         U126, U123, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349,
         P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342,
         P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335,
         P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328,
         P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, P1_U3322, P1_U3440,
         P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316,
         P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309,
         P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302,
         P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295,
         P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, P1_U3460, P1_U3463,
         P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, P1_U3481, P1_U3484,
         P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, P1_U3502, P1_U3505,
         P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515,
         P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522,
         P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529,
         P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536,
         P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543,
         P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550,
         P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, P1_U3290, P1_U3289,
         P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282,
         P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275,
         P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268,
         P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, P1_U3355, P1_U3262,
         P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255,
         P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248,
         P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3242, P1_U3241,
         P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561,
         P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568,
         P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575,
         P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582,
         P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, P1_U3239, P1_U3238,
         P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231,
         P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224,
         P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217,
         P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, P1_U3084,
         P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, P2_U3355, P2_U3354,
         P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, P2_U3348, P2_U3347,
         P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, P2_U3341, P2_U3340,
         P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, P2_U3334, P2_U3333,
         P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, P2_U3327, P2_U3437,
         P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321,
         P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314,
         P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307,
         P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300,
         P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, P2_U3457, P2_U3460,
         P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481,
         P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, P2_U3499, P2_U3502,
         P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512,
         P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519,
         P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526,
         P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, P2_U3532, P2_U3533,
         P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540,
         P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547,
         P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, P2_U3295, P2_U3294,
         P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287,
         P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280,
         P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273,
         P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266,
         P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259,
         P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252,
         P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245,
         P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558,
         P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, P2_U3564, P2_U3565,
         P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, P2_U3571, P2_U3572,
         P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, P2_U3578, P2_U3579,
         P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, P2_U3243, P2_U3242,
         P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235,
         P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228,
         P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221,
         P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3152,
         P2_U3151, P2_U3966;
  wire   n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271,
         n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281,
         n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291,
         n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301,
         n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311,
         n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321,
         n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331,
         n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341,
         n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351,
         n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361,
         n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371,
         n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381,
         n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391,
         n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401,
         n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411,
         n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421,
         n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431,
         n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441,
         n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451,
         n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461,
         n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471,
         n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481,
         n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491,
         n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501,
         n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511,
         n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521,
         n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531,
         n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541,
         n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551,
         n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561,
         n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571,
         n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581,
         n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591,
         n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601,
         n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611,
         n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621,
         n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631,
         n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641,
         n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651,
         n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661,
         n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671,
         n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681,
         n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691,
         n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701,
         n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711,
         n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721,
         n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731,
         n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741,
         n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751,
         n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761,
         n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771,
         n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781,
         n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791,
         n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801,
         n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811,
         n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821,
         n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831,
         n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841,
         n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851,
         n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861,
         n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871,
         n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881,
         n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891,
         n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901,
         n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911,
         n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921,
         n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931,
         n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941,
         n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951,
         n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961,
         n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971,
         n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981,
         n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991,
         n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001,
         n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011,
         n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021,
         n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031,
         n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041,
         n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051,
         n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061,
         n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071,
         n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081,
         n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091,
         n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101,
         n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111,
         n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121,
         n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131,
         n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141,
         n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151,
         n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161,
         n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171,
         n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181,
         n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191,
         n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201,
         n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211,
         n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221,
         n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231,
         n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241,
         n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251,
         n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261,
         n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271,
         n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281,
         n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291,
         n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301,
         n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311,
         n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321,
         n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331,
         n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341,
         n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351,
         n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361,
         n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371,
         n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381,
         n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391,
         n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401,
         n5402, n5403, n5404, n5405, n5407, n5408, n5409, n5410, n5411, n5412,
         n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422,
         n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432,
         n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442,
         n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452,
         n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462,
         n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472,
         n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482,
         n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492,
         n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502,
         n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512,
         n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522,
         n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532,
         n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542,
         n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552,
         n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562,
         n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572,
         n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582,
         n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592,
         n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602,
         n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612,
         n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622,
         n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632,
         n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642,
         n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652,
         n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662,
         n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672,
         n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682,
         n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692,
         n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702,
         n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712,
         n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722,
         n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732,
         n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742,
         n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752,
         n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762,
         n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772,
         n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782,
         n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792,
         n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802,
         n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812,
         n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822,
         n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832,
         n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842,
         n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852,
         n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862,
         n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872,
         n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882,
         n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892,
         n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902,
         n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912,
         n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922,
         n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932,
         n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942,
         n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952,
         n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962,
         n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972,
         n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982,
         n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992,
         n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002,
         n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012,
         n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022,
         n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032,
         n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042,
         n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052,
         n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062,
         n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072,
         n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082,
         n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092,
         n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102,
         n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112,
         n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122,
         n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132,
         n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142,
         n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152,
         n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162,
         n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172,
         n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182,
         n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192,
         n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202,
         n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212,
         n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222,
         n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232,
         n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242,
         n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252,
         n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262,
         n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272,
         n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282,
         n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292,
         n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302,
         n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312,
         n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322,
         n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332,
         n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342,
         n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352,
         n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362,
         n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372,
         n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382,
         n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392,
         n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402,
         n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412,
         n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422,
         n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432,
         n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442,
         n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452,
         n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462,
         n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472,
         n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482,
         n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492,
         n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502,
         n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512,
         n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522,
         n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532,
         n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542,
         n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552,
         n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562,
         n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572,
         n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582,
         n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592,
         n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602,
         n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612,
         n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622,
         n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632,
         n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642,
         n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652,
         n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662,
         n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672,
         n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682,
         n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692,
         n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702,
         n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712,
         n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722,
         n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732,
         n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742,
         n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752,
         n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762,
         n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772,
         n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782,
         n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792,
         n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802,
         n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812,
         n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822,
         n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832,
         n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842,
         n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852,
         n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862,
         n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872,
         n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882,
         n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892,
         n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902,
         n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912,
         n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922,
         n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932,
         n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942,
         n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952,
         n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962,
         n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972,
         n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982,
         n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992,
         n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002,
         n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012,
         n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022,
         n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032,
         n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042,
         n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052,
         n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062,
         n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072,
         n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082,
         n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092,
         n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102,
         n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112,
         n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122,
         n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132,
         n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142,
         n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152,
         n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162,
         n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172,
         n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182,
         n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192,
         n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202,
         n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212,
         n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222,
         n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232,
         n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242,
         n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252,
         n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262,
         n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272,
         n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282,
         n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292,
         n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302,
         n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312,
         n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322,
         n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332,
         n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342,
         n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352,
         n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362,
         n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372,
         n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382,
         n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392,
         n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402,
         n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412,
         n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422,
         n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432,
         n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442,
         n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452,
         n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462,
         n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472,
         n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482,
         n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492,
         n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502,
         n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512,
         n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522,
         n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532,
         n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542,
         n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552,
         n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562,
         n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572,
         n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582,
         n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592,
         n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602,
         n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612,
         n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622,
         n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632,
         n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642,
         n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652,
         n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662,
         n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672,
         n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682,
         n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692,
         n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702,
         n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712,
         n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722,
         n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732,
         n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742,
         n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752,
         n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762,
         n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772,
         n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782,
         n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792,
         n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802,
         n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812,
         n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822,
         n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832,
         n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842,
         n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852,
         n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862,
         n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872,
         n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882,
         n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892,
         n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902,
         n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912,
         n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922,
         n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932,
         n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942,
         n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952,
         n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962,
         n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972,
         n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982,
         n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992,
         n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002,
         n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012,
         n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022,
         n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032,
         n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042,
         n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052,
         n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062,
         n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072,
         n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082,
         n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092,
         n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102,
         n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112,
         n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122,
         n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132,
         n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142,
         n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152,
         n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162,
         n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172,
         n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182,
         n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192,
         n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202,
         n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212,
         n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222,
         n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232,
         n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242,
         n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252,
         n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262,
         n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272,
         n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282,
         n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292,
         n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302,
         n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312,
         n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322,
         n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332,
         n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342,
         n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352,
         n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362,
         n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372,
         n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382,
         n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392,
         n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402,
         n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412,
         n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422,
         n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432,
         n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442,
         n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452,
         n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462,
         n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472,
         n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482,
         n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492,
         n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502,
         n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512,
         n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522,
         n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532,
         n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542,
         n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552,
         n8553, n8554, n8555, n8556, n8557, n8558, n8560, n8561, n8562, n8563,
         n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573,
         n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583,
         n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593,
         n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603,
         n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613,
         n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623,
         n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633,
         n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643,
         n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653,
         n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663,
         n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673,
         n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683,
         n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693,
         n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703,
         n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713,
         n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723,
         n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733,
         n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743,
         n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753,
         n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763,
         n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773,
         n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783,
         n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793,
         n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803,
         n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813,
         n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823,
         n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833,
         n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843,
         n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853,
         n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863,
         n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873,
         n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883,
         n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893,
         n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903,
         n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913,
         n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923,
         n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933,
         n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943,
         n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953,
         n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963,
         n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973,
         n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983,
         n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993,
         n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003,
         n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013,
         n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023,
         n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033,
         n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043,
         n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053,
         n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063,
         n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073,
         n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083,
         n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093,
         n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103,
         n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113,
         n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123,
         n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133,
         n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143,
         n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153,
         n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163,
         n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173,
         n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183,
         n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193,
         n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203,
         n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213,
         n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223,
         n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233,
         n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243,
         n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253,
         n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263,
         n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273,
         n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283,
         n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293,
         n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303,
         n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313,
         n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323,
         n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333,
         n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343,
         n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353,
         n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363,
         n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373,
         n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383,
         n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393,
         n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403,
         n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413,
         n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423,
         n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433,
         n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443,
         n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453,
         n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463,
         n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473,
         n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483,
         n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493,
         n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503,
         n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513,
         n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523,
         n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533,
         n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543,
         n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553,
         n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563,
         n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573,
         n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583,
         n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593,
         n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603,
         n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613,
         n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623,
         n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633,
         n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643,
         n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653,
         n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663,
         n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673,
         n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683,
         n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693,
         n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703,
         n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713,
         n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723,
         n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733,
         n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743,
         n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753,
         n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763,
         n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773,
         n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783,
         n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793,
         n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803,
         n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813,
         n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823,
         n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833,
         n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843,
         n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853,
         n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863,
         n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873,
         n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883,
         n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893,
         n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903,
         n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913,
         n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923,
         n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933,
         n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943,
         n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953,
         n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963,
         n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973,
         n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983,
         n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993,
         n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001, n10002,
         n10003, n10004, n10005, n10006, n10007, n10008, n10009, n10010,
         n10011, n10012, n10013, n10014, n10015, n10016, n10017, n10018,
         n10019, n10020, n10021, n10022, n10023, n10024, n10025, n10026,
         n10027, n10028, n10029;

  NAND2_X2 U4767 ( .A1(n6596), .A2(P2_U3152), .ZN(n8049) );
  XNOR2_X1 U4768 ( .A(n8455), .B(n8453), .ZN(n8454) );
  NAND2_X1 U4769 ( .A1(n8346), .A2(n4274), .ZN(n8277) );
  NAND2_X1 U4770 ( .A1(n4507), .A2(n6505), .ZN(n8621) );
  NAND2_X1 U4771 ( .A1(n6197), .A2(n6196), .ZN(n9304) );
  NOR2_X1 U4772 ( .A1(n4550), .A2(n7683), .ZN(n9245) );
  OAI21_X1 U4773 ( .B1(n5316), .B2(n5315), .A(n5314), .ZN(n5331) );
  INV_X2 U4774 ( .A(n5641), .ZN(n6866) );
  INV_X1 U4775 ( .A(n5912), .ZN(n6213) );
  AND4_X1 U4776 ( .A1(n4939), .A2(n4938), .A3(n4937), .A4(n4936), .ZN(n6954)
         );
  INV_X1 U4777 ( .A(n6541), .ZN(n6536) );
  AND4_X1 U4779 ( .A1(n4917), .A2(n4916), .A3(n4915), .A4(n4914), .ZN(n7116)
         );
  AND4_X1 U4780 ( .A1(n4848), .A2(n4847), .A3(n4846), .A4(n4845), .ZN(n7117)
         );
  OAI21_X1 U4781 ( .B1(n5251), .B2(n4735), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n4861) );
  OAI211_X1 U4783 ( .C1(n4990), .C2(n6599), .A(n4904), .B(n4903), .ZN(n7123)
         );
  INV_X2 U4784 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n8552) );
  OAI21_X1 U4785 ( .B1(n8359), .B2(n4676), .A(n4674), .ZN(n5591) );
  NOR2_X1 U4786 ( .A1(P2_IR_REG_3__SCAN_IN), .A2(P2_IR_REG_2__SCAN_IN), .ZN(
        n4811) );
  INV_X2 U4787 ( .A(n6500), .ZN(n6370) );
  AND2_X1 U4788 ( .A1(n8346), .A2(n4502), .ZN(n8315) );
  INV_X2 U4789 ( .A(n6520), .ZN(n6544) );
  OAI21_X1 U4790 ( .B1(n9254), .B2(n4275), .A(n4324), .ZN(n9240) );
  NOR2_X2 U4791 ( .A1(n8366), .A2(n8486), .ZN(n8346) );
  INV_X1 U4792 ( .A(n6986), .ZN(n7052) );
  CLKBUF_X2 U4793 ( .A(n5957), .Z(n8718) );
  AOI21_X1 U4796 ( .B1(n4628), .B2(n4632), .A(n4326), .ZN(n4626) );
  NAND2_X1 U4797 ( .A1(n5394), .A2(n5393), .ZN(n8486) );
  INV_X1 U4798 ( .A(n7436), .ZN(n7156) );
  AND4_X1 U4799 ( .A1(n4989), .A2(n4988), .A3(n4987), .A4(n4986), .ZN(n8084)
         );
  INV_X1 U4800 ( .A(n6587), .ZN(n6586) );
  INV_X1 U4801 ( .A(n8949), .ZN(n6846) );
  AND2_X2 U4802 ( .A1(n9386), .A2(n9390), .ZN(n6223) );
  NAND2_X1 U4803 ( .A1(n6251), .A2(n5874), .ZN(n6587) );
  NAND2_X1 U4804 ( .A1(n5044), .A2(n5043), .ZN(n5062) );
  INV_X1 U4805 ( .A(n7123), .ZN(n6875) );
  AOI211_X1 U4806 ( .C1(n8471), .C2(n8450), .A(n8303), .B(n8302), .ZN(n8304)
         );
  XNOR2_X1 U4807 ( .A(n4861), .B(n4860), .ZN(n5645) );
  INV_X2 U4808 ( .A(n9609), .ZN(n9597) );
  NAND2_X1 U4809 ( .A1(n5432), .A2(n5431), .ZN(n8481) );
  NOR2_X2 U4810 ( .A1(n6846), .A2(n6311), .ZN(n6836) );
  INV_X1 U4811 ( .A(n6596), .ZN(n4262) );
  INV_X4 U4812 ( .A(n6596), .ZN(n6597) );
  NAND2_X2 U4813 ( .A1(n7544), .A2(n6414), .ZN(n7628) );
  NAND2_X2 U4814 ( .A1(n4776), .A2(n4333), .ZN(n7544) );
  OAI21_X2 U4815 ( .B1(n7497), .B2(n8836), .A(n8894), .ZN(n7425) );
  OAI21_X2 U4816 ( .B1(n5062), .B2(n5061), .A(n5063), .ZN(n5079) );
  XNOR2_X2 U4817 ( .A(n5867), .B(P1_IR_REG_26__SCAN_IN), .ZN(n6251) );
  NOR2_X2 U4818 ( .A1(n4949), .A2(P2_IR_REG_4__SCAN_IN), .ZN(n4971) );
  XNOR2_X2 U4819 ( .A(n5425), .B(n5420), .ZN(n7641) );
  XNOR2_X2 U4820 ( .A(n4837), .B(P2_IR_REG_30__SCAN_IN), .ZN(n8034) );
  XNOR2_X1 U4821 ( .A(n4897), .B(n4873), .ZN(n4896) );
  NAND2_X1 U4822 ( .A1(n4872), .A2(n4883), .ZN(n4897) );
  AND2_X1 U4823 ( .A1(n9386), .A2(n5899), .ZN(n6628) );
  AOI21_X1 U4824 ( .B1(n8168), .B2(n4395), .A(n4318), .ZN(n5418) );
  NAND2_X1 U4825 ( .A1(n5591), .A2(n5757), .ZN(n8310) );
  XNOR2_X1 U4826 ( .A(n5415), .B(n5413), .ZN(n8169) );
  NAND2_X1 U4827 ( .A1(n4519), .A2(n4518), .ZN(n8642) );
  NAND2_X1 U4828 ( .A1(n7788), .A2(n7789), .ZN(n5584) );
  NAND3_X1 U4829 ( .A1(n7370), .A2(n7368), .A3(n7369), .ZN(n7367) );
  NAND2_X1 U4830 ( .A1(n8139), .A2(n8087), .ZN(n5675) );
  NAND2_X1 U4831 ( .A1(n8084), .A2(n7156), .ZN(n5671) );
  NAND2_X1 U4832 ( .A1(n8247), .A2(n6875), .ZN(n5658) );
  INV_X1 U4833 ( .A(n6779), .ZN(n6867) );
  INV_X1 U4834 ( .A(n9725), .ZN(n7039) );
  INV_X1 U4835 ( .A(n6822), .ZN(n8824) );
  NAND2_X1 U4836 ( .A1(n8816), .A2(n9248), .ZN(n8814) );
  NOR2_X1 U4837 ( .A1(n6314), .A2(n6825), .ZN(n6823) );
  INV_X2 U4838 ( .A(n8666), .ZN(n6838) );
  INV_X1 U4839 ( .A(n5785), .ZN(n5749) );
  INV_X2 U4840 ( .A(n5645), .ZN(n5295) );
  INV_X1 U4841 ( .A(n5926), .ZN(n6014) );
  NOR2_X1 U4842 ( .A1(P1_IR_REG_17__SCAN_IN), .A2(P1_IR_REG_16__SCAN_IN), .ZN(
        n5863) );
  INV_X1 U4843 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n5861) );
  OR2_X1 U4844 ( .A1(n6580), .A2(n6551), .ZN(n6573) );
  AND2_X1 U4845 ( .A1(n4783), .A2(n4782), .ZN(n8686) );
  AND2_X1 U4846 ( .A1(n4700), .A2(n4278), .ZN(n8070) );
  NAND2_X1 U4847 ( .A1(n6499), .A2(n6498), .ZN(n8652) );
  AND2_X1 U4848 ( .A1(n4630), .A2(n4329), .ZN(n4628) );
  INV_X1 U4849 ( .A(n4675), .ZN(n4674) );
  OR2_X1 U4850 ( .A1(n8353), .A2(n4809), .ZN(n4806) );
  AND2_X1 U4851 ( .A1(n4361), .A2(n4359), .ZN(n9051) );
  AOI21_X1 U4852 ( .B1(n8422), .B2(n4295), .A(n4788), .ZN(n8373) );
  INV_X1 U4853 ( .A(n4808), .ZN(n4807) );
  OAI21_X1 U4854 ( .B1(n4809), .B2(n8357), .A(n8060), .ZN(n4808) );
  OR2_X1 U4855 ( .A1(n9047), .A2(n9510), .ZN(n4361) );
  AOI21_X1 U4856 ( .B1(n7811), .B2(n5246), .A(n5245), .ZN(n7797) );
  NAND2_X1 U4857 ( .A1(n7582), .A2(n5707), .ZN(n7662) );
  AND2_X1 U4858 ( .A1(n9246), .A2(n4335), .ZN(n9166) );
  NAND2_X1 U4859 ( .A1(n9697), .A2(n7553), .ZN(n9696) );
  NAND2_X1 U4860 ( .A1(n7367), .A2(n6395), .ZN(n7386) );
  NAND2_X1 U4861 ( .A1(n5335), .A2(n5334), .ZN(n8502) );
  OR2_X1 U4862 ( .A1(n8927), .A2(n9253), .ZN(n4275) );
  NAND2_X1 U4863 ( .A1(n5273), .A2(n5272), .ZN(n8519) );
  NAND2_X1 U4864 ( .A1(n6113), .A2(n6112), .ZN(n9347) );
  NAND2_X1 U4865 ( .A1(n6376), .A2(n6375), .ZN(n7369) );
  OR2_X1 U4866 ( .A1(n6284), .A2(n8840), .ZN(n7674) );
  NAND2_X1 U4867 ( .A1(n6063), .A2(n6062), .ZN(n7691) );
  NAND2_X1 U4868 ( .A1(n8740), .A2(n8749), .ZN(n8840) );
  NAND2_X1 U4869 ( .A1(n4490), .A2(n4489), .ZN(n9699) );
  NAND2_X1 U4870 ( .A1(n6078), .A2(n6077), .ZN(n7648) );
  OR2_X1 U4871 ( .A1(n7078), .A2(n7075), .ZN(n6386) );
  NAND2_X2 U4872 ( .A1(n6049), .A2(n6048), .ZN(n9358) );
  INV_X1 U4873 ( .A(n9698), .ZN(n4490) );
  OAI21_X1 U4874 ( .B1(n7177), .B2(n4285), .A(n4656), .ZN(n7496) );
  OAI21_X1 U4875 ( .B1(n6907), .B2(n4666), .A(n5686), .ZN(n4665) );
  OR2_X1 U4876 ( .A1(n4667), .A2(n4668), .ZN(n4666) );
  NAND2_X2 U4877 ( .A1(n7188), .A2(n9613), .ZN(n9609) );
  NAND2_X1 U4878 ( .A1(n5648), .A2(n5663), .ZN(n6956) );
  NAND2_X1 U4879 ( .A1(n6954), .A2(n9725), .ZN(n5790) );
  AND4_X1 U4880 ( .A1(n5011), .A2(n5010), .A3(n5009), .A4(n5008), .ZN(n8139)
         );
  OAI211_X1 U4881 ( .C1(n4990), .C2(n6606), .A(n4976), .B(n4975), .ZN(n6986)
         );
  AOI21_X1 U4882 ( .B1(n6370), .B2(n6311), .A(n6315), .ZN(n6316) );
  INV_X4 U4883 ( .A(n6522), .ZN(n6377) );
  NAND2_X2 U4884 ( .A1(n7028), .A2(n4876), .ZN(n5433) );
  NAND3_X1 U4885 ( .A1(n4579), .A2(n4580), .A3(n4995), .ZN(n5014) );
  INV_X1 U4886 ( .A(n4913), .ZN(n4933) );
  INV_X1 U4887 ( .A(n6309), .ZN(n8997) );
  CLKBUF_X1 U4888 ( .A(n6309), .Z(n8816) );
  AND2_X1 U4889 ( .A1(n4844), .A2(n8557), .ZN(n4913) );
  AND2_X1 U4890 ( .A1(n7090), .A2(n6587), .ZN(n6320) );
  AND2_X1 U4891 ( .A1(n4844), .A2(n4843), .ZN(n4935) );
  OAI211_X1 U4892 ( .C1(n6014), .C2(n6599), .A(n5929), .B(n5928), .ZN(n8666)
         );
  CLKBUF_X1 U4893 ( .A(n6304), .Z(n8951) );
  INV_X1 U4894 ( .A(n4843), .ZN(n8557) );
  AND2_X1 U4895 ( .A1(n6590), .A2(n6597), .ZN(n5926) );
  AND2_X1 U4896 ( .A1(n6590), .A2(n6596), .ZN(n5957) );
  NAND2_X1 U4897 ( .A1(n5856), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5859) );
  NAND2_X1 U4898 ( .A1(n4841), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4837) );
  XNOR2_X1 U4899 ( .A(n5860), .B(n5861), .ZN(n8987) );
  XNOR2_X1 U4900 ( .A(n5886), .B(P1_IR_REG_30__SCAN_IN), .ZN(n9386) );
  NOR2_X1 U4901 ( .A1(n5060), .A2(n4320), .ZN(n5211) );
  OR2_X1 U4902 ( .A1(n5889), .A2(n9380), .ZN(n5886) );
  OR2_X1 U4903 ( .A1(n5894), .A2(n9380), .ZN(n4544) );
  OR2_X1 U4904 ( .A1(n6074), .A2(n4819), .ZN(n5880) );
  NOR2_X1 U4905 ( .A1(n5871), .A2(n4434), .ZN(n5894) );
  NAND2_X2 U4906 ( .A1(n6597), .A2(P1_U3084), .ZN(n6951) );
  NAND2_X1 U4907 ( .A1(n4436), .A2(n4435), .ZN(n4434) );
  NAND2_X1 U4908 ( .A1(n6072), .A2(n5866), .ZN(n5871) );
  NAND2_X1 U4909 ( .A1(n4818), .A2(n5872), .ZN(n4785) );
  AND4_X1 U4910 ( .A1(n6016), .A2(n5851), .A3(n5850), .A4(n5849), .ZN(n5852)
         );
  NAND2_X1 U4911 ( .A1(n5848), .A2(n4775), .ZN(n4774) );
  AND4_X1 U4912 ( .A1(n5176), .A2(n4854), .A3(n4731), .A4(n4851), .ZN(n4830)
         );
  INV_X1 U4913 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n5875) );
  INV_X1 U4914 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n9857) );
  INV_X1 U4915 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n4761) );
  NOR2_X1 U4916 ( .A1(P1_IR_REG_7__SCAN_IN), .A2(P1_IR_REG_11__SCAN_IN), .ZN(
        n5851) );
  NOR2_X1 U4917 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(P1_IR_REG_10__SCAN_IN), .ZN(
        n5850) );
  NOR2_X1 U4918 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_12__SCAN_IN), .ZN(
        n5849) );
  NOR2_X1 U4919 ( .A1(P2_IR_REG_7__SCAN_IN), .A2(P2_IR_REG_6__SCAN_IN), .ZN(
        n4849) );
  NOR2_X1 U4920 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(P1_IR_REG_2__SCAN_IN), .ZN(
        n5847) );
  INV_X1 U4921 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n4851) );
  INV_X1 U4922 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n5179) );
  INV_X1 U4923 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n5176) );
  NOR2_X1 U4924 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(P1_IR_REG_6__SCAN_IN), .ZN(
        n6016) );
  INV_X1 U4925 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n4854) );
  INV_X1 U4926 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n5848) );
  INV_X1 U4927 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n4856) );
  INV_X1 U4928 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n9847) );
  INV_X1 U4929 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n5881) );
  INV_X1 U4930 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n4760) );
  INV_X4 U4931 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3152) );
  INV_X1 U4932 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n6085) );
  INV_X1 U4933 ( .A(n4933), .ZN(n5475) );
  OR2_X1 U4934 ( .A1(n7118), .A2(n6962), .ZN(n7034) );
  NOR3_X2 U4935 ( .A1(n7665), .A2(n4499), .A3(n8519), .ZN(n4497) );
  XNOR2_X2 U4936 ( .A(n5445), .B(n5444), .ZN(n7722) );
  NOR2_X2 U4937 ( .A1(n9144), .A2(n9310), .ZN(n9136) );
  NAND3_X2 U4938 ( .A1(n5908), .A2(n5907), .A3(n4451), .ZN(n6321) );
  AOI21_X2 U4939 ( .B1(n9359), .B2(n9284), .A(n9283), .ZN(n9285) );
  AND4_X2 U4940 ( .A1(n4894), .A2(n4893), .A3(n4892), .A4(n4891), .ZN(n5576)
         );
  INV_X1 U4941 ( .A(n5575), .ZN(n7462) );
  OAI211_X2 U4942 ( .C1(n4990), .C2(n6603), .A(n4875), .B(n4874), .ZN(n5575)
         );
  AND2_X2 U4943 ( .A1(n6245), .A2(n9083), .ZN(n9060) );
  XNOR2_X2 U4944 ( .A(n4544), .B(n5896), .ZN(n5909) );
  OR2_X1 U4945 ( .A1(n6199), .A2(n6198), .ZN(n6210) );
  INV_X1 U4946 ( .A(n4923), .ZN(n5023) );
  AOI21_X1 U4947 ( .B1(n4716), .B2(n4718), .A(n4715), .ZN(n4714) );
  INV_X1 U4948 ( .A(n8201), .ZN(n4715) );
  NAND2_X1 U4949 ( .A1(n4804), .A2(n4301), .ZN(n4803) );
  INV_X2 U4950 ( .A(n5023), .ZN(n5634) );
  INV_X1 U4951 ( .A(n4264), .ZN(n6226) );
  NAND2_X1 U4952 ( .A1(n4433), .A2(n4432), .ZN(n8745) );
  NAND2_X1 U4953 ( .A1(n8738), .A2(n4445), .ZN(n4433) );
  NAND2_X1 U4954 ( .A1(n8737), .A2(n8814), .ZN(n4432) );
  NAND2_X1 U4955 ( .A1(n4419), .A2(n4423), .ZN(n4418) );
  INV_X1 U4956 ( .A(n4407), .ZN(n4406) );
  NAND2_X1 U4957 ( .A1(n8811), .A2(n8809), .ZN(n4443) );
  NOR2_X1 U4958 ( .A1(P1_IR_REG_27__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), .ZN(
        n5895) );
  AND2_X1 U4959 ( .A1(n5078), .A2(n4713), .ZN(n4719) );
  INV_X1 U4960 ( .A(n8109), .ZN(n4713) );
  OR2_X1 U4961 ( .A1(n8509), .A2(n8154), .ZN(n5738) );
  AND2_X1 U4962 ( .A1(n5807), .A2(n4685), .ZN(n4681) );
  NOR2_X1 U4963 ( .A1(n5580), .A2(n4690), .ZN(n4689) );
  INV_X1 U4964 ( .A(n5804), .ZN(n4690) );
  AND2_X1 U4965 ( .A1(n7201), .A2(n7199), .ZN(n4802) );
  INV_X1 U4966 ( .A(n7407), .ZN(n7201) );
  OR2_X1 U4967 ( .A1(n8460), .A2(n6758), .ZN(n5777) );
  NOR2_X1 U4968 ( .A1(n8530), .A2(n7820), .ZN(n4500) );
  INV_X1 U4969 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n4392) );
  INV_X1 U4970 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n4831) );
  NAND2_X1 U4971 ( .A1(n4853), .A2(n4731), .ZN(n4730) );
  INV_X1 U4972 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n5090) );
  AND2_X1 U4973 ( .A1(n4973), .A2(n4849), .ZN(n5051) );
  INV_X1 U4974 ( .A(n8582), .ZN(n4526) );
  NOR2_X1 U4975 ( .A1(n9124), .A2(n4634), .ZN(n4633) );
  INV_X1 U4976 ( .A(n4636), .ZN(n4634) );
  INV_X1 U4977 ( .A(n8851), .ZN(n4639) );
  INV_X1 U4978 ( .A(n4621), .ZN(n4619) );
  OR2_X1 U4979 ( .A1(n6152), .A2(n8591), .ZN(n6163) );
  OR2_X1 U4980 ( .A1(n4552), .A2(n4553), .ZN(n4550) );
  OR2_X1 U4981 ( .A1(n7648), .A2(n9264), .ZN(n4552) );
  OR2_X1 U4982 ( .A1(n9264), .A2(n9243), .ZN(n8925) );
  NAND2_X1 U4983 ( .A1(n5601), .A2(n5600), .ZN(n5612) );
  NAND2_X1 U4984 ( .A1(n5597), .A2(n5596), .ZN(n5601) );
  NAND2_X1 U4985 ( .A1(n4585), .A2(n4586), .ZN(n5487) );
  INV_X1 U4986 ( .A(n4587), .ZN(n4586) );
  OAI21_X1 U4987 ( .B1(n4589), .B2(n4588), .A(n5463), .ZN(n4587) );
  INV_X1 U4988 ( .A(n5423), .ZN(n4593) );
  OAI21_X1 U4989 ( .B1(n4607), .B2(n4606), .A(n4349), .ZN(n4605) );
  INV_X1 U4990 ( .A(n5288), .ZN(n4606) );
  INV_X1 U4991 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n4775) );
  AND2_X1 U4992 ( .A1(n7229), .A2(n5077), .ZN(n5078) );
  OR2_X1 U4993 ( .A1(n5231), .A2(n5230), .ZN(n5233) );
  OR2_X1 U4994 ( .A1(n5829), .A2(n9715), .ZN(n5641) );
  NAND2_X1 U4995 ( .A1(n8080), .A2(n5025), .ZN(n8133) );
  NAND2_X1 U4996 ( .A1(n5506), .A2(n5645), .ZN(n5829) );
  NOR2_X1 U4997 ( .A1(n8005), .A2(n8004), .ZN(n8003) );
  OR2_X1 U4998 ( .A1(n8486), .A2(n8362), .ZN(n5752) );
  AOI21_X1 U4999 ( .B1(n8373), .B2(n8382), .A(n8058), .ZN(n8353) );
  AND2_X1 U5000 ( .A1(n8353), .A2(n8357), .ZN(n8355) );
  OR2_X1 U5001 ( .A1(n8526), .A2(n7828), .ZN(n5721) );
  NAND2_X1 U5002 ( .A1(n8053), .A2(n8052), .ZN(n8435) );
  AOI21_X1 U5003 ( .B1(n4671), .B2(n4673), .A(n4313), .ZN(n4670) );
  AND2_X1 U5004 ( .A1(n7783), .A2(n5710), .ZN(n7759) );
  NAND2_X1 U5005 ( .A1(n9696), .A2(n4311), .ZN(n7578) );
  NAND2_X1 U5006 ( .A1(n5636), .A2(n5635), .ZN(n8453) );
  AND3_X1 U5007 ( .A1(n4973), .A2(n4833), .A3(n4297), .ZN(n5508) );
  XNOR2_X1 U5008 ( .A(n4863), .B(P2_IR_REG_21__SCAN_IN), .ZN(n5821) );
  NAND2_X1 U5009 ( .A1(n4289), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4863) );
  NAND2_X1 U5010 ( .A1(n5211), .A2(n4855), .ZN(n5251) );
  NAND2_X1 U5011 ( .A1(n5845), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n6222) );
  INV_X1 U5012 ( .A(n6223), .ZN(n6212) );
  AND4_X1 U5013 ( .A1(n5925), .A2(n5924), .A3(n5923), .A4(n5922), .ZN(n7104)
         );
  OR2_X1 U5014 ( .A1(n5855), .A2(n5854), .ZN(n4819) );
  AND2_X1 U5015 ( .A1(n5904), .A2(n5903), .ZN(n9096) );
  INV_X1 U5016 ( .A(n9143), .ZN(n6301) );
  NAND2_X1 U5017 ( .A1(n7092), .A2(n6269), .ZN(n6991) );
  NAND2_X1 U5018 ( .A1(n5890), .A2(n9381), .ZN(n5899) );
  NAND2_X1 U5019 ( .A1(n8723), .A2(n8814), .ZN(n4447) );
  OAI21_X1 U5020 ( .B1(n8722), .B2(n4446), .A(n4445), .ZN(n4444) );
  OAI21_X1 U5021 ( .B1(n4431), .B2(n8747), .A(n4430), .ZN(n4429) );
  AND2_X1 U5022 ( .A1(n8746), .A2(n8835), .ZN(n4430) );
  AOI21_X1 U5023 ( .B1(n8745), .B2(n8744), .A(n8743), .ZN(n4431) );
  NOR2_X1 U5024 ( .A1(n4428), .A2(n4427), .ZN(n4426) );
  INV_X1 U5025 ( .A(n8748), .ZN(n4427) );
  INV_X1 U5026 ( .A(n8749), .ZN(n4428) );
  NAND2_X1 U5027 ( .A1(n8791), .A2(n9176), .ZN(n4424) );
  OAI21_X1 U5028 ( .B1(n8780), .B2(n4449), .A(n4448), .ZN(n8782) );
  NAND2_X1 U5029 ( .A1(n8778), .A2(n8880), .ZN(n4449) );
  NOR2_X1 U5030 ( .A1(n8823), .A2(n8814), .ZN(n4448) );
  AOI21_X1 U5031 ( .B1(n4416), .B2(n4415), .A(n8814), .ZN(n4414) );
  INV_X1 U5032 ( .A(n4419), .ZN(n4415) );
  NOR2_X1 U5033 ( .A1(n5349), .A2(n4408), .ZN(n4407) );
  INV_X1 U5034 ( .A(n5313), .ZN(n4408) );
  AOI21_X1 U5035 ( .B1(n4698), .B2(n8281), .A(n5618), .ZN(n4697) );
  INV_X1 U5036 ( .A(n5675), .ZN(n4668) );
  INV_X1 U5037 ( .A(n5671), .ZN(n4667) );
  INV_X1 U5038 ( .A(n6276), .ZN(n4658) );
  INV_X1 U5039 ( .A(n9211), .ZN(n4455) );
  OAI21_X1 U5040 ( .B1(n5612), .B2(n5611), .A(n5610), .ZN(n5629) );
  AND2_X1 U5041 ( .A1(n4739), .A2(n5198), .ZN(n4738) );
  AND2_X1 U5042 ( .A1(n4738), .A2(n4602), .ZN(n4601) );
  NAND2_X1 U5043 ( .A1(n4603), .A2(n5130), .ZN(n4602) );
  INV_X1 U5044 ( .A(n5126), .ZN(n4603) );
  NAND2_X1 U5045 ( .A1(n4601), .A2(n4604), .ZN(n4598) );
  INV_X1 U5046 ( .A(n5130), .ZN(n4604) );
  INV_X1 U5047 ( .A(n4583), .ZN(n4582) );
  OAI21_X1 U5048 ( .B1(n4965), .B2(n4584), .A(n4991), .ZN(n4583) );
  INV_X1 U5049 ( .A(n4969), .ZN(n4584) );
  INV_X1 U5050 ( .A(P1_RD_REG_SCAN_IN), .ZN(n4759) );
  INV_X1 U5051 ( .A(n7743), .ZN(n4728) );
  NOR2_X1 U5052 ( .A1(n7619), .A2(n4727), .ZN(n4726) );
  INV_X1 U5053 ( .A(n5150), .ZN(n4727) );
  XNOR2_X1 U5054 ( .A(n8142), .B(n5433), .ZN(n5074) );
  NOR2_X1 U5055 ( .A1(n4724), .A2(n4400), .ZN(n4398) );
  INV_X1 U5056 ( .A(n4401), .ZN(n4400) );
  INV_X1 U5057 ( .A(n4726), .ZN(n4722) );
  NOR2_X1 U5058 ( .A1(n8123), .A2(n4410), .ZN(n4409) );
  INV_X1 U5059 ( .A(n5281), .ZN(n4410) );
  OR2_X1 U5060 ( .A1(n8466), .A2(n8299), .ZN(n8064) );
  INV_X1 U5061 ( .A(n5752), .ZN(n4676) );
  OR2_X1 U5062 ( .A1(n8481), .A2(n8313), .ZN(n5757) );
  INV_X1 U5063 ( .A(n8057), .ZN(n4789) );
  OR2_X1 U5064 ( .A1(n8497), .A2(n8361), .ZN(n8356) );
  NAND2_X1 U5065 ( .A1(n7793), .A2(n4500), .ZN(n4499) );
  AND2_X1 U5066 ( .A1(n5807), .A2(n5806), .ZN(n9690) );
  NOR2_X1 U5067 ( .A1(n7436), .A2(n8084), .ZN(n4799) );
  OAI21_X1 U5068 ( .B1(n7156), .B2(n8243), .A(n6905), .ZN(n4801) );
  NOR2_X1 U5069 ( .A1(n4798), .A2(n4799), .ZN(n4796) );
  NAND2_X1 U5070 ( .A1(n5658), .A2(n6955), .ZN(n4812) );
  AND2_X1 U5071 ( .A1(n5830), .A2(n5821), .ZN(n5567) );
  AND2_X1 U5072 ( .A1(n4297), .A2(n4834), .ZN(n4814) );
  INV_X1 U5073 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n4834) );
  AND2_X1 U5074 ( .A1(n4827), .A2(n4849), .ZN(n4829) );
  INV_X1 U5075 ( .A(n6419), .ZN(n4517) );
  INV_X1 U5076 ( .A(n4770), .ZN(n4515) );
  OAI22_X1 U5077 ( .A1(n6522), .A2(n6992), .B1(n9650), .B2(n6500), .ZN(n6340)
         );
  AND2_X1 U5078 ( .A1(n4766), .A2(n6492), .ZN(n4765) );
  INV_X1 U5079 ( .A(n4538), .ZN(n4537) );
  NAND2_X1 U5080 ( .A1(n8612), .A2(n4539), .ZN(n4538) );
  INV_X1 U5081 ( .A(n6455), .ZN(n4539) );
  OR2_X1 U5082 ( .A1(n9293), .A2(n9107), .ZN(n8869) );
  OR2_X1 U5083 ( .A1(n9288), .A2(n9096), .ZN(n8865) );
  NOR2_X1 U5084 ( .A1(n8890), .A2(n4465), .ZN(n4464) );
  OR2_X1 U5085 ( .A1(n9320), .A2(n9152), .ZN(n8822) );
  NOR2_X1 U5086 ( .A1(n4620), .A2(n4617), .ZN(n4616) );
  INV_X1 U5087 ( .A(n4623), .ZN(n4617) );
  INV_X1 U5088 ( .A(n9186), .ZN(n4620) );
  NAND2_X1 U5089 ( .A1(n4328), .A2(n4266), .ZN(n4621) );
  NAND2_X1 U5090 ( .A1(n5841), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n6135) );
  INV_X1 U5091 ( .A(n6125), .ZN(n5841) );
  OR2_X1 U5092 ( .A1(n6114), .A2(n8614), .ZN(n6125) );
  NOR2_X1 U5093 ( .A1(n6282), .A2(n6287), .ZN(n4644) );
  NOR2_X1 U5094 ( .A1(n8704), .A2(n9435), .ZN(n4643) );
  INV_X1 U5095 ( .A(n7673), .ZN(n4368) );
  AND2_X1 U5096 ( .A1(n9260), .A2(n4751), .ZN(n4750) );
  NAND2_X1 U5097 ( .A1(n6088), .A2(n6014), .ZN(n4751) );
  NAND2_X1 U5098 ( .A1(n5839), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n6090) );
  INV_X1 U5099 ( .A(n6079), .ZN(n5839) );
  OR2_X1 U5100 ( .A1(n9358), .A2(n7698), .ZN(n8740) );
  NAND2_X1 U5101 ( .A1(n8997), .A2(n9049), .ZN(n6816) );
  AND2_X1 U5102 ( .A1(n4548), .A2(n9214), .ZN(n9176) );
  XNOR2_X1 U5103 ( .A(n5629), .B(n5628), .ZN(n5627) );
  INV_X1 U5104 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n5896) );
  INV_X1 U5105 ( .A(n5895), .ZN(n4530) );
  INV_X1 U5106 ( .A(n4785), .ZN(n4436) );
  AND2_X1 U5107 ( .A1(n5866), .A2(n4533), .ZN(n4532) );
  NOR2_X1 U5108 ( .A1(n4785), .A2(n5895), .ZN(n4533) );
  AND2_X1 U5109 ( .A1(n5463), .A2(n5451), .ZN(n5461) );
  AOI21_X1 U5110 ( .B1(n5424), .B2(n4592), .A(n4590), .ZN(n4589) );
  INV_X1 U5111 ( .A(n5443), .ZN(n4590) );
  OAI21_X1 U5112 ( .B1(n5379), .B2(n5378), .A(n5377), .ZN(n5389) );
  INV_X1 U5113 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n5876) );
  AND2_X1 U5114 ( .A1(n5332), .A2(n5321), .ZN(n5330) );
  AND2_X1 U5115 ( .A1(n5266), .A2(n5249), .ZN(n4607) );
  INV_X1 U5116 ( .A(n5152), .ZN(n4743) );
  OR2_X1 U5117 ( .A1(n6042), .A2(P1_IR_REG_11__SCAN_IN), .ZN(n6043) );
  NAND2_X1 U5118 ( .A1(n4600), .A2(n5130), .ZN(n5153) );
  NAND2_X1 U5119 ( .A1(n8191), .A2(n5376), .ZN(n5415) );
  NAND2_X1 U5120 ( .A1(n8093), .A2(n5485), .ZN(n5548) );
  NAND2_X1 U5121 ( .A1(n4397), .A2(n4396), .ZN(n7229) );
  INV_X1 U5122 ( .A(n7227), .ZN(n4397) );
  NAND2_X1 U5123 ( .A1(n8133), .A2(n5072), .ZN(n7230) );
  AOI21_X1 U5124 ( .B1(n4719), .B2(n4717), .A(n4323), .ZN(n4716) );
  INV_X1 U5125 ( .A(n5072), .ZN(n4717) );
  INV_X1 U5126 ( .A(n4719), .ZN(n4718) );
  NAND2_X1 U5127 ( .A1(n5003), .A2(n5002), .ZN(n8080) );
  AND2_X1 U5128 ( .A1(n8216), .A2(n4705), .ZN(n4704) );
  NAND2_X1 U5129 ( .A1(n4279), .A2(n4706), .ZN(n4705) );
  INV_X1 U5130 ( .A(n4708), .ZN(n4706) );
  INV_X1 U5131 ( .A(n4279), .ZN(n4707) );
  MUX2_X1 U5132 ( .A(n5787), .B(n5786), .S(n5785), .Z(n5788) );
  AND4_X1 U5133 ( .A1(n5237), .A2(n5236), .A3(n5235), .A4(n5234), .ZN(n7840)
         );
  AND4_X1 U5134 ( .A1(n4964), .A2(n4963), .A3(n4962), .A4(n4961), .ZN(n6978)
         );
  NOR2_X1 U5135 ( .A1(n8003), .A2(n4291), .ZN(n7992) );
  OR2_X1 U5136 ( .A1(n7992), .A2(n7991), .ZN(n4476) );
  NOR2_X1 U5137 ( .A1(n7975), .A2(n4340), .ZN(n7967) );
  OR2_X1 U5138 ( .A1(n7967), .A2(n7966), .ZN(n4482) );
  OR2_X1 U5139 ( .A1(n7933), .A2(n7932), .ZN(n4480) );
  AND2_X1 U5140 ( .A1(n4480), .A2(n4479), .ZN(n7922) );
  NAND2_X1 U5141 ( .A1(n7351), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n4479) );
  OR2_X1 U5142 ( .A1(n7922), .A2(n7921), .ZN(n4478) );
  NOR2_X1 U5143 ( .A1(n7908), .A2(n4356), .ZN(n7899) );
  NOR2_X1 U5144 ( .A1(n7899), .A2(n7900), .ZN(n7898) );
  NOR2_X1 U5145 ( .A1(n4852), .A2(P2_IR_REG_9__SCAN_IN), .ZN(n4853) );
  INV_X1 U5146 ( .A(n8459), .ZN(n8269) );
  OR2_X1 U5147 ( .A1(n8477), .A2(n8300), .ZN(n8062) );
  AND2_X1 U5148 ( .A1(n8367), .A2(n8232), .ZN(n8059) );
  NAND2_X1 U5149 ( .A1(n8344), .A2(n4810), .ZN(n4809) );
  INV_X1 U5150 ( .A(n8059), .ZN(n4810) );
  NAND2_X1 U5151 ( .A1(n8359), .A2(n4267), .ZN(n8341) );
  NAND2_X1 U5152 ( .A1(n4504), .A2(n4503), .ZN(n8366) );
  AND4_X1 U5153 ( .A1(n5402), .A2(n5401), .A3(n5400), .A4(n5399), .ZN(n8362)
         );
  AND4_X1 U5154 ( .A1(n5410), .A2(n5409), .A3(n5408), .A4(n5407), .ZN(n8383)
         );
  NAND2_X1 U5155 ( .A1(n8412), .A2(n8396), .ZN(n8391) );
  AOI21_X1 U5156 ( .B1(n4791), .B2(n8056), .A(n4309), .ZN(n4790) );
  NOR2_X1 U5157 ( .A1(n8418), .A2(n4792), .ZN(n4791) );
  INV_X1 U5158 ( .A(n4794), .ZN(n4792) );
  OR2_X1 U5159 ( .A1(n8515), .A2(n8446), .ZN(n4794) );
  OR2_X1 U5160 ( .A1(n8422), .A2(n8056), .ZN(n4793) );
  AND2_X1 U5161 ( .A1(n5738), .A2(n5739), .ZN(n8418) );
  INV_X1 U5162 ( .A(n4679), .ZN(n4678) );
  OAI21_X1 U5163 ( .B1(n4284), .B2(n4680), .A(n8424), .ZN(n4679) );
  INV_X1 U5164 ( .A(n5726), .ZN(n4680) );
  AND2_X1 U5165 ( .A1(n5725), .A2(n8408), .ZN(n8424) );
  NAND2_X1 U5166 ( .A1(n5584), .A2(n4284), .ZN(n8442) );
  NOR2_X1 U5167 ( .A1(n7665), .A2(n4499), .ZN(n8436) );
  OR2_X1 U5168 ( .A1(n5255), .A2(n7885), .ZN(n5302) );
  AND2_X1 U5169 ( .A1(n5721), .A2(n5719), .ZN(n7789) );
  NAND2_X1 U5170 ( .A1(n7662), .A2(n7661), .ZN(n7660) );
  AND2_X1 U5171 ( .A1(n7849), .A2(n5567), .ZN(n8443) );
  INV_X1 U5172 ( .A(n9756), .ZN(n8445) );
  NAND2_X1 U5173 ( .A1(n7578), .A2(n4286), .ZN(n7659) );
  AOI21_X1 U5174 ( .B1(n4689), .B2(n4687), .A(n4686), .ZN(n4685) );
  INV_X1 U5175 ( .A(n4689), .ZN(n4688) );
  AND2_X1 U5176 ( .A1(n7552), .A2(n7551), .ZN(n9697) );
  INV_X1 U5177 ( .A(n9690), .ZN(n7553) );
  AND4_X1 U5178 ( .A1(n5104), .A2(n5103), .A3(n5102), .A4(n5101), .ZN(n9757)
         );
  NAND2_X1 U5179 ( .A1(n4385), .A2(n4384), .ZN(n7205) );
  OAI21_X1 U5180 ( .B1(n9749), .B2(n4386), .A(n7203), .ZN(n4384) );
  INV_X1 U5181 ( .A(n7202), .ZN(n4386) );
  NAND2_X1 U5182 ( .A1(n7200), .A2(n4802), .ZN(n7404) );
  INV_X1 U5183 ( .A(n8443), .ZN(n9758) );
  AND2_X1 U5184 ( .A1(n5652), .A2(n5794), .ZN(n4662) );
  NAND2_X1 U5185 ( .A1(n4662), .A2(n7112), .ZN(n7114) );
  NAND2_X1 U5186 ( .A1(n6769), .A2(n6770), .ZN(n6874) );
  OR2_X1 U5187 ( .A1(n9741), .A2(n5821), .ZN(n6762) );
  NAND2_X1 U5188 ( .A1(n5560), .A2(n5567), .ZN(n9756) );
  INV_X1 U5189 ( .A(n9693), .ZN(n9753) );
  NAND2_X1 U5190 ( .A1(n6778), .A2(n6777), .ZN(n9693) );
  NAND2_X1 U5191 ( .A1(n5606), .A2(n5605), .ZN(n8460) );
  INV_X1 U5192 ( .A(n9726), .ZN(n9788) );
  INV_X1 U5193 ( .A(n6766), .ZN(n9715) );
  OR2_X1 U5194 ( .A1(n6687), .A2(n5525), .ZN(n9707) );
  AND2_X1 U5195 ( .A1(n7779), .A2(n5528), .ZN(n9708) );
  NAND2_X1 U5196 ( .A1(n4842), .A2(n4841), .ZN(n4843) );
  NAND2_X1 U5197 ( .A1(n4394), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4393) );
  NAND2_X1 U5198 ( .A1(n5517), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5524) );
  AOI21_X1 U5199 ( .B1(n5251), .B2(P2_IR_REG_31__SCAN_IN), .A(n4733), .ZN(
        n4732) );
  NAND2_X1 U5200 ( .A1(n4734), .A2(n4860), .ZN(n4733) );
  NAND2_X1 U5201 ( .A1(n4735), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4734) );
  INV_X1 U5202 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n4832) );
  INV_X1 U5203 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n4711) );
  OR2_X1 U5204 ( .A1(n6163), .A2(n8655), .ZN(n6175) );
  NAND2_X1 U5205 ( .A1(n8697), .A2(n8698), .ZN(n4777) );
  OR2_X1 U5206 ( .A1(n6090), .A2(n6089), .ZN(n6099) );
  NAND2_X1 U5207 ( .A1(n4541), .A2(n4777), .ZN(n8604) );
  AND2_X1 U5208 ( .A1(n8696), .A2(n8606), .ZN(n4541) );
  NAND2_X1 U5209 ( .A1(n8574), .A2(n8575), .ZN(n8622) );
  INV_X1 U5210 ( .A(n4508), .ZN(n4507) );
  NAND2_X1 U5211 ( .A1(n8662), .A2(n4506), .ZN(n8631) );
  AND2_X1 U5212 ( .A1(n6856), .A2(n6339), .ZN(n4506) );
  OR2_X1 U5213 ( .A1(n4521), .A2(n4524), .ZN(n4520) );
  NOR2_X1 U5214 ( .A1(n4526), .A2(n4522), .ZN(n4521) );
  INV_X1 U5215 ( .A(n8672), .ZN(n4522) );
  NOR2_X1 U5216 ( .A1(n7693), .A2(n4771), .ZN(n4770) );
  INV_X1 U5217 ( .A(n6422), .ZN(n4771) );
  NAND2_X1 U5218 ( .A1(n7628), .A2(n6419), .ZN(n4772) );
  NAND2_X1 U5219 ( .A1(n7386), .A2(n7384), .ZN(n4776) );
  AOI21_X1 U5220 ( .B1(n4782), .B2(n6517), .A(n8685), .ZN(n4780) );
  INV_X1 U5221 ( .A(n8597), .ZN(n4782) );
  NAND2_X1 U5222 ( .A1(n4438), .A2(n4437), .ZN(n8819) );
  AND2_X1 U5223 ( .A1(n4334), .A2(n4441), .ZN(n4437) );
  NAND2_X1 U5224 ( .A1(n9057), .A2(n9055), .ZN(n4822) );
  AND2_X1 U5225 ( .A1(n8987), .A2(n9049), .ZN(n6817) );
  OR2_X1 U5226 ( .A1(n9525), .A2(n9524), .ZN(n4565) );
  AOI21_X1 U5227 ( .B1(P1_REG1_REG_8__SCAN_IN), .B2(n9516), .A(n9511), .ZN(
        n9530) );
  AND2_X1 U5228 ( .A1(n4565), .A2(n4564), .ZN(n6725) );
  NAND2_X1 U5229 ( .A1(n9528), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n4564) );
  OR2_X1 U5230 ( .A1(n6725), .A2(n6724), .ZN(n4563) );
  XNOR2_X1 U5231 ( .A(n7595), .B(n7599), .ZN(n9551) );
  OAI21_X1 U5232 ( .B1(n9554), .B2(P1_REG1_REG_14__SCAN_IN), .A(n9555), .ZN(
        n7709) );
  OR2_X1 U5233 ( .A1(n7598), .A2(n7597), .ZN(n4569) );
  OR2_X1 U5234 ( .A1(n6222), .A2(n5846), .ZN(n6248) );
  NOR2_X1 U5235 ( .A1(n9093), .A2(n8868), .ZN(n4745) );
  NAND2_X1 U5236 ( .A1(n4459), .A2(n4457), .ZN(n9104) );
  AOI21_X1 U5237 ( .B1(n4461), .B2(n4463), .A(n4458), .ZN(n4457) );
  INV_X1 U5238 ( .A(n8797), .ZN(n4458) );
  AOI21_X1 U5239 ( .B1(n4633), .B2(n4631), .A(n4322), .ZN(n4630) );
  INV_X1 U5240 ( .A(n4283), .ZN(n4631) );
  INV_X1 U5241 ( .A(n4633), .ZN(n4632) );
  AND2_X1 U5242 ( .A1(n4462), .A2(n9124), .ZN(n4461) );
  OR2_X1 U5243 ( .A1(n4464), .A2(n4463), .ZN(n4462) );
  NAND2_X1 U5244 ( .A1(n9155), .A2(n4464), .ZN(n4460) );
  NAND2_X1 U5245 ( .A1(n4327), .A2(n4639), .ZN(n4636) );
  AND2_X1 U5246 ( .A1(n8873), .A2(n8797), .ZN(n9124) );
  OR2_X1 U5247 ( .A1(n8851), .A2(n4296), .ZN(n9132) );
  AOI21_X1 U5248 ( .B1(n9160), .B2(n6299), .A(n6298), .ZN(n9143) );
  AND2_X1 U5249 ( .A1(n9320), .A2(n9179), .ZN(n6298) );
  INV_X1 U5250 ( .A(n9150), .ZN(n6183) );
  NAND2_X1 U5251 ( .A1(n9212), .A2(n9211), .ZN(n6139) );
  NAND2_X1 U5252 ( .A1(n9246), .A2(n4549), .ZN(n9205) );
  AND2_X1 U5253 ( .A1(n8880), .A2(n8891), .ZN(n9211) );
  NAND2_X1 U5254 ( .A1(n6295), .A2(n6294), .ZN(n9204) );
  OAI21_X1 U5255 ( .B1(n9240), .B2(n8772), .A(n8774), .ZN(n9229) );
  OR2_X1 U5256 ( .A1(n8772), .A2(n8769), .ZN(n9241) );
  NAND2_X1 U5257 ( .A1(n6098), .A2(n6097), .ZN(n9264) );
  NAND2_X1 U5258 ( .A1(n6071), .A2(n8752), .ZN(n9254) );
  NAND2_X1 U5259 ( .A1(n7177), .A2(n4268), .ZN(n7242) );
  NAND2_X1 U5260 ( .A1(n4473), .A2(n5977), .ZN(n7180) );
  AND2_X1 U5261 ( .A1(n4474), .A2(n5976), .ZN(n4473) );
  INV_X1 U5262 ( .A(n7183), .ZN(n4474) );
  AND4_X1 U5263 ( .A1(n5945), .A2(n5944), .A3(n5943), .A4(n5942), .ZN(n7103)
         );
  AND2_X1 U5264 ( .A1(n8902), .A2(n8724), .ZN(n7063) );
  NAND2_X1 U5265 ( .A1(n6991), .A2(n8828), .ZN(n6990) );
  OR2_X1 U5266 ( .A1(n6588), .A2(n8993), .ZN(n9586) );
  NAND2_X1 U5267 ( .A1(n6833), .A2(n6268), .ZN(n4612) );
  NAND2_X1 U5268 ( .A1(n5957), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n4511) );
  OR2_X1 U5269 ( .A1(n6014), .A2(n6605), .ZN(n4510) );
  NAND2_X1 U5270 ( .A1(n4614), .A2(n6267), .ZN(n6835) );
  INV_X1 U5271 ( .A(n6833), .ZN(n4614) );
  NAND2_X1 U5272 ( .A1(n5920), .A2(n5919), .ZN(n8956) );
  INV_X1 U5273 ( .A(n8825), .ZN(n6267) );
  INV_X1 U5274 ( .A(n9586), .ZN(n9231) );
  XNOR2_X1 U5275 ( .A(n6321), .B(n8949), .ZN(n6822) );
  NAND2_X1 U5276 ( .A1(n8716), .A2(n8715), .ZN(n9276) );
  AOI21_X1 U5277 ( .B1(n4470), .B2(n9590), .A(n4748), .ZN(n9286) );
  OAI22_X1 U5278 ( .A1(n9096), .A2(n6241), .B1(n6243), .B2(n6242), .ZN(n4748)
         );
  XNOR2_X1 U5279 ( .A(n4749), .B(n8856), .ZN(n4470) );
  AND2_X1 U5280 ( .A1(n9288), .A2(n9002), .ZN(n6302) );
  NAND2_X1 U5281 ( .A1(n6208), .A2(n6207), .ZN(n9300) );
  NAND2_X1 U5282 ( .A1(n6186), .A2(n6185), .ZN(n9310) );
  INV_X1 U5283 ( .A(n9149), .ZN(n9313) );
  INV_X1 U5284 ( .A(n9269), .ZN(n4654) );
  INV_X1 U5285 ( .A(n9270), .ZN(n4655) );
  OR2_X1 U5286 ( .A1(n7094), .A2(n8942), .ZN(n9664) );
  NAND2_X1 U5287 ( .A1(n8816), .A2(n8861), .ZN(n7094) );
  XNOR2_X1 U5288 ( .A(n5627), .B(SI_30_), .ZN(n8717) );
  XNOR2_X1 U5289 ( .A(n5597), .B(n5596), .ZN(n7846) );
  INV_X1 U5290 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n5853) );
  INV_X1 U5291 ( .A(n5946), .ZN(n4773) );
  CLKBUF_X1 U5292 ( .A(n5960), .Z(n5961) );
  NAND2_X1 U5293 ( .A1(n4945), .A2(n4370), .ZN(n4369) );
  INV_X1 U5294 ( .A(n4946), .ZN(n4370) );
  AND4_X1 U5295 ( .A1(n5168), .A2(n5167), .A3(n5166), .A4(n5165), .ZN(n7746)
         );
  AND2_X1 U5296 ( .A1(n4886), .A2(n6868), .ZN(n8042) );
  NAND2_X1 U5297 ( .A1(n8041), .A2(n8042), .ZN(n8040) );
  AND4_X1 U5298 ( .A1(n5329), .A2(n5328), .A3(n5327), .A4(n5326), .ZN(n8154)
         );
  NAND2_X1 U5299 ( .A1(n5216), .A2(n5215), .ZN(n8530) );
  NAND2_X1 U5300 ( .A1(n5254), .A2(n5253), .ZN(n8526) );
  AND4_X1 U5301 ( .A1(n5144), .A2(n5143), .A3(n5142), .A4(n5141), .ZN(n8204)
         );
  NAND2_X1 U5302 ( .A1(n5229), .A2(n5228), .ZN(n7820) );
  INV_X1 U5303 ( .A(n7840), .ZN(n8234) );
  NAND2_X1 U5304 ( .A1(n8029), .A2(n9679), .ZN(n4486) );
  AOI21_X1 U5305 ( .B1(n4270), .B2(n8028), .A(n4485), .ZN(n4484) );
  NAND2_X1 U5306 ( .A1(n8030), .A2(n5295), .ZN(n4485) );
  NAND2_X1 U5307 ( .A1(n8274), .A2(n4377), .ZN(n4375) );
  NOR2_X1 U5308 ( .A1(n8071), .A2(n4379), .ZN(n4377) );
  OR2_X1 U5309 ( .A1(n8274), .A2(n4380), .ZN(n4376) );
  INV_X1 U5310 ( .A(n8071), .ZN(n4380) );
  OR2_X1 U5311 ( .A1(n8355), .A2(n8354), .ZN(n8491) );
  NAND2_X1 U5312 ( .A1(n9808), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n4381) );
  NOR2_X1 U5313 ( .A1(n4282), .A2(n4496), .ZN(n4495) );
  INV_X1 U5314 ( .A(n8457), .ZN(n4496) );
  AND4_X1 U5315 ( .A1(n5971), .A2(n5970), .A3(n5969), .A4(n5968), .ZN(n7185)
         );
  NAND2_X1 U5316 ( .A1(n6134), .A2(n6133), .ZN(n9334) );
  INV_X1 U5317 ( .A(n8688), .ZN(n6574) );
  AND4_X1 U5318 ( .A1(n5984), .A2(n5983), .A3(n5982), .A4(n5981), .ZN(n7307)
         );
  NAND2_X1 U5319 ( .A1(n4769), .A2(n8644), .ZN(n8590) );
  NAND2_X1 U5320 ( .A1(n8642), .A2(n8643), .ZN(n4769) );
  AND2_X1 U5321 ( .A1(n6182), .A2(n6181), .ZN(n9164) );
  AND4_X1 U5322 ( .A1(n6001), .A2(n6000), .A3(n5999), .A4(n5998), .ZN(n9588)
         );
  AND2_X1 U5323 ( .A1(n6159), .A2(n6158), .ZN(n9165) );
  INV_X1 U5324 ( .A(n9173), .ZN(n9320) );
  AND2_X1 U5325 ( .A1(n6206), .A2(n6205), .ZN(n9135) );
  NAND2_X1 U5326 ( .A1(n6218), .A2(n6217), .ZN(n9126) );
  NAND2_X1 U5327 ( .A1(n6195), .A2(n6194), .ZN(n9125) );
  OR2_X1 U5328 ( .A1(n8625), .A2(n6212), .ZN(n6195) );
  AOI21_X1 U5329 ( .B1(n9478), .B2(P1_REG1_REG_5__SCAN_IN), .A(n9473), .ZN(
        n9493) );
  NOR2_X1 U5330 ( .A1(n9485), .A2(n4343), .ZN(n9503) );
  NAND2_X1 U5331 ( .A1(n9503), .A2(n9504), .ZN(n9502) );
  NAND2_X1 U5332 ( .A1(n6234), .A2(n6233), .ZN(n9284) );
  OR2_X1 U5333 ( .A1(n9287), .A2(n9271), .ZN(n6307) );
  AND2_X1 U5334 ( .A1(n9609), .A2(n6845), .ZN(n9605) );
  NAND2_X1 U5335 ( .A1(n4447), .A2(n4444), .ZN(n8732) );
  NAND2_X1 U5336 ( .A1(n4429), .A2(n4426), .ZN(n8750) );
  AOI21_X1 U5337 ( .B1(n4422), .B2(n4421), .A(n4420), .ZN(n4419) );
  INV_X1 U5338 ( .A(n8791), .ZN(n4421) );
  INV_X1 U5339 ( .A(n8821), .ZN(n4420) );
  INV_X1 U5340 ( .A(n8782), .ZN(n8781) );
  AOI21_X1 U5341 ( .B1(n8777), .B2(n8776), .A(n8775), .ZN(n8780) );
  AND2_X1 U5342 ( .A1(n8298), .A2(n5594), .ZN(n4694) );
  NOR2_X1 U5343 ( .A1(n4699), .A2(n4696), .ZN(n4695) );
  INV_X1 U5344 ( .A(n5594), .ZN(n4696) );
  OR2_X1 U5345 ( .A1(n4833), .A2(n8552), .ZN(n4390) );
  NOR2_X1 U5346 ( .A1(n4768), .A2(n4764), .ZN(n4763) );
  INV_X1 U5347 ( .A(n8643), .ZN(n4764) );
  INV_X1 U5348 ( .A(n8589), .ZN(n4768) );
  NAND2_X1 U5349 ( .A1(n8589), .A2(n4767), .ZN(n4766) );
  INV_X1 U5350 ( .A(n8644), .ZN(n4767) );
  AOI21_X1 U5351 ( .B1(n4414), .B2(n4417), .A(n4465), .ZN(n4412) );
  OR2_X1 U5352 ( .A1(n8789), .A2(n4417), .ZN(n4413) );
  INV_X1 U5353 ( .A(n5461), .ZN(n4588) );
  INV_X1 U5354 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n5290) );
  AOI21_X1 U5355 ( .B1(n4407), .B2(n4405), .A(n4314), .ZN(n4404) );
  OR2_X1 U5356 ( .A1(n4710), .A2(n4406), .ZN(n4403) );
  INV_X1 U5357 ( .A(n4409), .ZN(n4405) );
  NOR2_X1 U5358 ( .A1(n8265), .A2(n8264), .ZN(n5783) );
  MUX2_X1 U5359 ( .A(n5817), .B(n5818), .S(n5785), .Z(n5781) );
  NOR2_X1 U5360 ( .A1(n8481), .A2(n8477), .ZN(n4502) );
  OR2_X1 U5361 ( .A1(n8486), .A2(n8231), .ZN(n8060) );
  INV_X1 U5362 ( .A(n4672), .ZN(n4671) );
  OAI21_X1 U5363 ( .B1(n7661), .B2(n4673), .A(n5583), .ZN(n4672) );
  INV_X1 U5364 ( .A(n5582), .ZN(n4673) );
  NAND2_X1 U5365 ( .A1(n7757), .A2(n4805), .ZN(n4804) );
  INV_X1 U5366 ( .A(n7658), .ZN(n4805) );
  INV_X1 U5367 ( .A(SI_15_), .ZN(n9921) );
  INV_X1 U5368 ( .A(SI_9_), .ZN(n9908) );
  AOI21_X1 U5369 ( .B1(n4664), .B2(n4663), .A(n4665), .ZN(n7406) );
  INV_X1 U5370 ( .A(n4666), .ZN(n4663) );
  NAND2_X1 U5371 ( .A1(n8282), .A2(n5769), .ZN(n4700) );
  AND2_X1 U5372 ( .A1(n9764), .A2(n9767), .ZN(n9766) );
  AND2_X1 U5373 ( .A1(n7462), .A2(n4505), .ZN(n7119) );
  OR2_X1 U5374 ( .A1(P2_IR_REG_27__SCAN_IN), .A2(P2_IR_REG_26__SCAN_IN), .ZN(
        n4864) );
  INV_X1 U5375 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n4394) );
  NAND2_X1 U5376 ( .A1(n4390), .A2(n4388), .ZN(n4387) );
  AND2_X1 U5377 ( .A1(n8552), .A2(P2_IR_REG_27__SCAN_IN), .ZN(n4388) );
  NAND2_X1 U5378 ( .A1(n4509), .A2(n8652), .ZN(n4508) );
  NAND2_X1 U5379 ( .A1(n8651), .A2(n8654), .ZN(n4509) );
  NAND2_X1 U5380 ( .A1(n6335), .A2(n6334), .ZN(n6336) );
  NOR2_X1 U5381 ( .A1(n4443), .A2(n4290), .ZN(n4439) );
  AOI21_X1 U5382 ( .B1(n4272), .B2(n4299), .A(n8810), .ZN(n4440) );
  INV_X1 U5383 ( .A(n4442), .ZN(n4441) );
  OAI21_X1 U5384 ( .B1(n4272), .B2(n8814), .A(n8813), .ZN(n4442) );
  INV_X1 U5385 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n6064) );
  NOR2_X1 U5386 ( .A1(n7594), .A2(n4571), .ZN(n7595) );
  AND2_X1 U5387 ( .A1(n7601), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n4571) );
  AND2_X1 U5388 ( .A1(n4266), .A2(n6297), .ZN(n4623) );
  NOR2_X1 U5389 ( .A1(n9339), .A2(n9334), .ZN(n4549) );
  NAND2_X1 U5390 ( .A1(n9269), .A2(n6292), .ZN(n4653) );
  INV_X1 U5391 ( .A(n6292), .ZN(n4650) );
  NAND2_X1 U5392 ( .A1(n6923), .A2(n8714), .ZN(n4754) );
  OR2_X1 U5393 ( .A1(n7691), .A2(n8695), .ZN(n4553) );
  AND2_X1 U5394 ( .A1(n7691), .A2(n9009), .ZN(n6285) );
  NAND2_X1 U5395 ( .A1(n5837), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n6051) );
  INV_X1 U5396 ( .A(n6034), .ZN(n5837) );
  INV_X1 U5397 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n6021) );
  INV_X1 U5398 ( .A(n4657), .ZN(n4656) );
  OAI21_X1 U5399 ( .B1(n4268), .B2(n4285), .A(n6277), .ZN(n4657) );
  OR2_X1 U5400 ( .A1(n6007), .A2(n6006), .ZN(n6022) );
  INV_X1 U5401 ( .A(n4746), .ZN(n4456) );
  NAND2_X1 U5402 ( .A1(n4746), .A2(n4455), .ZN(n4454) );
  NOR2_X1 U5403 ( .A1(n8823), .A2(n4747), .ZN(n4746) );
  NAND2_X1 U5404 ( .A1(n5896), .A2(n4435), .ZN(n4784) );
  AND2_X1 U5405 ( .A1(n5488), .A2(n5469), .ZN(n5486) );
  AND2_X1 U5406 ( .A1(n5390), .A2(n5385), .ZN(n5388) );
  AND2_X1 U5407 ( .A1(n4598), .A2(n4737), .ZN(n4597) );
  AOI21_X1 U5408 ( .B1(n4271), .B2(n4738), .A(n4348), .ZN(n4737) );
  AOI21_X1 U5409 ( .B1(n5173), .B2(n4741), .A(n4740), .ZN(n4739) );
  INV_X1 U5410 ( .A(n5175), .ZN(n4740) );
  INV_X1 U5411 ( .A(n5151), .ZN(n4741) );
  NAND2_X1 U5412 ( .A1(n4582), .A2(n4584), .ZN(n4580) );
  NAND2_X1 U5413 ( .A1(n4966), .A2(n4582), .ZN(n4579) );
  AND2_X2 U5414 ( .A1(n4758), .A2(n4756), .ZN(n6596) );
  INV_X1 U5415 ( .A(P2_RD_REG_SCAN_IN), .ZN(n4757) );
  OR2_X1 U5416 ( .A1(n5454), .A2(n8219), .ZN(n5473) );
  NAND2_X1 U5417 ( .A1(n7615), .A2(n4726), .ZN(n4725) );
  NAND2_X1 U5418 ( .A1(n7824), .A2(n7823), .ZN(n4710) );
  NOR2_X1 U5419 ( .A1(n7612), .A2(n4402), .ZN(n4401) );
  INV_X1 U5420 ( .A(n5123), .ZN(n4402) );
  OR2_X1 U5421 ( .A1(n8172), .A2(n8171), .ZN(n4395) );
  NAND2_X1 U5422 ( .A1(n4399), .A2(n4720), .ZN(n7811) );
  AOI21_X1 U5423 ( .B1(n4723), .B2(n4722), .A(n4721), .ZN(n4720) );
  INV_X1 U5424 ( .A(n5197), .ZN(n4721) );
  NOR2_X1 U5425 ( .A1(n5415), .A2(n5414), .ZN(n8168) );
  OR2_X1 U5426 ( .A1(n8135), .A2(n5076), .ZN(n7227) );
  NAND2_X1 U5427 ( .A1(n4710), .A2(n4409), .ZN(n8121) );
  OR2_X1 U5428 ( .A1(n5324), .A2(n9926), .ZN(n5367) );
  AND2_X1 U5429 ( .A1(n6760), .A2(n6759), .ZN(n7027) );
  OR2_X1 U5430 ( .A1(n8159), .A2(n4709), .ZN(n4708) );
  INV_X1 U5431 ( .A(n8158), .ZN(n4709) );
  NAND2_X1 U5432 ( .A1(n4862), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5516) );
  NOR2_X1 U5433 ( .A1(n6695), .A2(n6696), .ZN(n7339) );
  AND2_X1 U5434 ( .A1(n4476), .A2(n4475), .ZN(n7977) );
  NAND2_X1 U5435 ( .A1(n7342), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n4475) );
  AND2_X1 U5436 ( .A1(n4482), .A2(n4481), .ZN(n7956) );
  NAND2_X1 U5437 ( .A1(n7345), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n4481) );
  NOR2_X1 U5438 ( .A1(n7956), .A2(n7955), .ZN(n7954) );
  AND2_X1 U5439 ( .A1(n4478), .A2(n4477), .ZN(n7910) );
  NAND2_X1 U5440 ( .A1(n7353), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n4477) );
  INV_X1 U5441 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n8203) );
  NOR2_X1 U5442 ( .A1(n7898), .A2(n4354), .ZN(n7360) );
  NAND2_X1 U5443 ( .A1(n7360), .A2(n7359), .ZN(n7449) );
  NOR2_X1 U5444 ( .A1(n5060), .A2(n4730), .ZN(n5158) );
  NOR2_X1 U5445 ( .A1(n7873), .A2(n7874), .ZN(n8251) );
  NAND2_X1 U5446 ( .A1(n8251), .A2(n8250), .ZN(n8249) );
  NAND2_X1 U5447 ( .A1(n8249), .A2(n4471), .ZN(n7888) );
  OR2_X1 U5448 ( .A1(n8258), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n4471) );
  NOR2_X1 U5449 ( .A1(n7888), .A2(n7887), .ZN(n7886) );
  INV_X1 U5450 ( .A(n8064), .ZN(n4379) );
  NAND2_X1 U5451 ( .A1(n8308), .A2(n5760), .ZN(n8297) );
  NAND2_X1 U5452 ( .A1(n8346), .A2(n4269), .ZN(n8291) );
  OAI21_X1 U5453 ( .B1(n4267), .B2(n4676), .A(n5814), .ZN(n4675) );
  AND2_X1 U5454 ( .A1(n5481), .A2(n5480), .ZN(n8314) );
  NAND2_X1 U5455 ( .A1(n5761), .A2(n5760), .ZN(n8311) );
  OR2_X1 U5456 ( .A1(n8481), .A2(n8230), .ZN(n8061) );
  NAND2_X1 U5457 ( .A1(n8306), .A2(n8311), .ZN(n8305) );
  AND2_X1 U5458 ( .A1(n8346), .A2(n8331), .ZN(n8326) );
  AND4_X1 U5459 ( .A1(n5372), .A2(n5371), .A3(n5370), .A4(n5369), .ZN(n8361)
         );
  OAI21_X1 U5460 ( .B1(n4790), .B2(n4789), .A(n4317), .ZN(n4788) );
  INV_X1 U5461 ( .A(n5233), .ZN(n5217) );
  AND2_X1 U5462 ( .A1(n4683), .A2(n5806), .ZN(n4682) );
  INV_X1 U5463 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n5138) );
  NAND2_X1 U5464 ( .A1(n9766), .A2(n9772), .ZN(n7260) );
  AND2_X1 U5465 ( .A1(n5804), .A2(n5803), .ZN(n7209) );
  AND4_X1 U5466 ( .A1(n5119), .A2(n5118), .A3(n5117), .A4(n5116), .ZN(n8112)
         );
  AND2_X1 U5467 ( .A1(n9751), .A2(n5676), .ZN(n7407) );
  AND4_X1 U5468 ( .A1(n5059), .A2(n5058), .A3(n5057), .A4(n5056), .ZN(n8138)
         );
  AND4_X1 U5469 ( .A1(n5038), .A2(n5037), .A3(n5036), .A4(n5035), .ZN(n9759)
         );
  NAND2_X1 U5470 ( .A1(n4795), .A2(n4797), .ZN(n7198) );
  OR2_X1 U5471 ( .A1(n4800), .A2(n4799), .ZN(n4797) );
  INV_X1 U5472 ( .A(n4801), .ZN(n4800) );
  NAND2_X1 U5473 ( .A1(n5578), .A2(n6907), .ZN(n6912) );
  AND2_X1 U5474 ( .A1(n7033), .A2(n7052), .ZN(n6916) );
  NAND2_X1 U5475 ( .A1(n6958), .A2(n4659), .ZN(n6883) );
  AND2_X1 U5476 ( .A1(n5790), .A2(n5648), .ZN(n4659) );
  NOR2_X2 U5477 ( .A1(n7034), .A2(n9725), .ZN(n7033) );
  NAND2_X1 U5478 ( .A1(n7119), .A2(n6875), .ZN(n7118) );
  AND2_X1 U5479 ( .A1(n7419), .A2(n7380), .ZN(n6766) );
  NAND2_X1 U5480 ( .A1(n4700), .A2(n4698), .ZN(n8069) );
  AND2_X1 U5481 ( .A1(n5777), .A2(n5776), .ZN(n8071) );
  NAND2_X1 U5482 ( .A1(n5471), .A2(n5470), .ZN(n8470) );
  NAND2_X1 U5483 ( .A1(n5362), .A2(n5361), .ZN(n8497) );
  INV_X1 U5484 ( .A(n4500), .ZN(n4498) );
  NAND2_X1 U5485 ( .A1(n7404), .A2(n7202), .ZN(n9750) );
  AND2_X1 U5486 ( .A1(n5829), .A2(n6766), .ZN(n9726) );
  NAND2_X1 U5487 ( .A1(n5514), .A2(n5513), .ZN(n5529) );
  NAND2_X1 U5488 ( .A1(n4292), .A2(n4833), .ZN(n5513) );
  NAND2_X1 U5489 ( .A1(n4867), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5512) );
  XNOR2_X1 U5490 ( .A(n5524), .B(n5523), .ZN(n5826) );
  NAND2_X1 U5491 ( .A1(n4856), .A2(n4736), .ZN(n4735) );
  INV_X1 U5492 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n4860) );
  OAI21_X1 U5493 ( .B1(n5251), .B2(P2_IR_REG_17__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5271) );
  AND2_X1 U5494 ( .A1(n5110), .A2(n5092), .ZN(n7355) );
  AOI21_X1 U5495 ( .B1(n4515), .B2(n4514), .A(n4293), .ZN(n4512) );
  INV_X1 U5496 ( .A(n4353), .ZN(n4514) );
  NAND2_X1 U5497 ( .A1(n5843), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n6188) );
  NAND2_X1 U5498 ( .A1(n6343), .A2(n6344), .ZN(n6856) );
  INV_X1 U5499 ( .A(n6099), .ZN(n5840) );
  NAND2_X1 U5500 ( .A1(n8631), .A2(n6350), .ZN(n8632) );
  XNOR2_X1 U5501 ( .A(n6338), .B(n6336), .ZN(n8664) );
  NAND2_X1 U5502 ( .A1(n8661), .A2(n8664), .ZN(n8662) );
  AOI21_X1 U5503 ( .B1(n6447), .B2(n4304), .A(n4536), .ZN(n4535) );
  NOR2_X1 U5504 ( .A1(n4540), .A2(n4537), .ZN(n4536) );
  AND2_X1 U5505 ( .A1(n8612), .A2(n8606), .ZN(n4540) );
  NAND2_X1 U5506 ( .A1(n5891), .A2(n4450), .ZN(n4453) );
  AND2_X1 U5507 ( .A1(n5899), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n4450) );
  NAND2_X1 U5508 ( .A1(n6672), .A2(n6807), .ZN(n6671) );
  NAND2_X1 U5509 ( .A1(n6650), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n4364) );
  AOI21_X1 U5510 ( .B1(P1_REG1_REG_3__SCAN_IN), .B2(n6719), .A(n6708), .ZN(
        n9462) );
  NAND2_X1 U5511 ( .A1(n9538), .A2(n9539), .ZN(n9537) );
  AND2_X1 U5512 ( .A1(n4563), .A2(n4562), .ZN(n9541) );
  NAND2_X1 U5513 ( .A1(n6942), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n4562) );
  NAND2_X1 U5514 ( .A1(n9537), .A2(n4363), .ZN(n6936) );
  OR2_X1 U5515 ( .A1(n9536), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n4363) );
  NAND2_X1 U5516 ( .A1(n7006), .A2(n7007), .ZN(n7600) );
  AND2_X1 U5517 ( .A1(n8865), .A2(n8804), .ZN(n9069) );
  NAND2_X1 U5518 ( .A1(n4555), .A2(n4554), .ZN(n9089) );
  AND2_X1 U5519 ( .A1(n6230), .A2(n6229), .ZN(n9107) );
  AND2_X1 U5520 ( .A1(n6210), .A2(n6200), .ZN(n9119) );
  NAND2_X1 U5521 ( .A1(n9136), .A2(n9121), .ZN(n9116) );
  AND2_X1 U5522 ( .A1(n6170), .A2(n6169), .ZN(n9152) );
  OR2_X1 U5523 ( .A1(n9167), .A2(n9313), .ZN(n9144) );
  NAND2_X1 U5524 ( .A1(n9177), .A2(n8791), .ZN(n9162) );
  NAND2_X1 U5525 ( .A1(n4615), .A2(n4618), .ZN(n9160) );
  AOI21_X1 U5526 ( .B1(n4619), .B2(n9186), .A(n4315), .ZN(n4618) );
  NAND2_X1 U5527 ( .A1(n4622), .A2(n4621), .ZN(n9187) );
  NAND2_X1 U5528 ( .A1(n9204), .A2(n4623), .ZN(n4622) );
  AND2_X1 U5529 ( .A1(n9245), .A2(n6244), .ZN(n9246) );
  NAND2_X1 U5530 ( .A1(n9246), .A2(n9227), .ZN(n9221) );
  OAI21_X1 U5531 ( .B1(n9270), .B2(n4651), .A(n4649), .ZN(n9220) );
  INV_X1 U5532 ( .A(n4652), .ZN(n4651) );
  AOI21_X1 U5533 ( .B1(n4652), .B2(n4650), .A(n4308), .ZN(n4649) );
  AND2_X1 U5534 ( .A1(n4653), .A2(n6293), .ZN(n4652) );
  AND3_X1 U5535 ( .A1(n6131), .A2(n6130), .A3(n6129), .ZN(n9244) );
  OR2_X1 U5536 ( .A1(n9255), .A2(n8927), .ZN(n4488) );
  AND2_X1 U5537 ( .A1(n8925), .A2(n6291), .ZN(n9269) );
  NAND2_X1 U5538 ( .A1(n4755), .A2(n8920), .ZN(n9255) );
  INV_X1 U5539 ( .A(n7727), .ZN(n4755) );
  NAND2_X1 U5540 ( .A1(n4754), .A2(n6088), .ZN(n8695) );
  NAND2_X1 U5541 ( .A1(n4641), .A2(n4367), .ZN(n7725) );
  AOI21_X1 U5542 ( .B1(n6286), .B2(n4644), .A(n4643), .ZN(n4641) );
  INV_X1 U5543 ( .A(n6287), .ZN(n4645) );
  AND2_X1 U5544 ( .A1(n8924), .A2(n8920), .ZN(n8846) );
  NAND2_X1 U5545 ( .A1(n6059), .A2(n8753), .ZN(n7677) );
  INV_X1 U5546 ( .A(n9008), .ZN(n8704) );
  AND2_X1 U5547 ( .A1(n8755), .A2(n8752), .ZN(n8842) );
  NAND2_X1 U5548 ( .A1(n6032), .A2(n6031), .ZN(n7428) );
  OR2_X1 U5549 ( .A1(n7503), .A2(n7428), .ZN(n7489) );
  AND4_X1 U5550 ( .A1(n6056), .A2(n6055), .A3(n6054), .A4(n6053), .ZN(n7698)
         );
  NAND2_X1 U5551 ( .A1(n9581), .A2(n9395), .ZN(n7503) );
  AND2_X1 U5552 ( .A1(n9579), .A2(n9663), .ZN(n9581) );
  NAND2_X1 U5553 ( .A1(n7242), .A2(n6276), .ZN(n9578) );
  NOR2_X1 U5554 ( .A1(n7246), .A2(n7267), .ZN(n9579) );
  NAND2_X1 U5555 ( .A1(n4547), .A2(n7192), .ZN(n7246) );
  AND2_X1 U5556 ( .A1(n7060), .A2(n6272), .ZN(n7135) );
  NAND2_X1 U5557 ( .A1(n7135), .A2(n8729), .ZN(n7134) );
  AND2_X1 U5558 ( .A1(n7064), .A2(n9657), .ZN(n7141) );
  AND2_X1 U5559 ( .A1(n4545), .A2(n8636), .ZN(n7064) );
  NOR2_X1 U5560 ( .A1(n7096), .A2(n7100), .ZN(n4545) );
  AND4_X1 U5561 ( .A1(n5934), .A2(n5933), .A3(n5932), .A4(n5931), .ZN(n6992)
         );
  NAND2_X1 U5562 ( .A1(n4546), .A2(n9650), .ZN(n7098) );
  INV_X1 U5563 ( .A(n7096), .ZN(n4546) );
  AND2_X1 U5564 ( .A1(n8954), .A2(n8959), .ZN(n8825) );
  AND2_X1 U5565 ( .A1(n6562), .A2(n6520), .ZN(n6844) );
  AND3_X2 U5566 ( .A1(n4647), .A2(n4646), .A3(n4273), .ZN(n8949) );
  NAND2_X1 U5567 ( .A1(n5926), .A2(n5910), .ZN(n4646) );
  NAND2_X1 U5568 ( .A1(n5957), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n4647) );
  OR2_X1 U5569 ( .A1(n8814), .A2(n8942), .ZN(n7145) );
  AND2_X1 U5570 ( .A1(n6737), .A2(n8990), .ZN(n9359) );
  XNOR2_X1 U5571 ( .A(n4609), .B(n5632), .ZN(n8551) );
  OAI21_X1 U5572 ( .B1(n5627), .B2(n5626), .A(n5630), .ZN(n4609) );
  XNOR2_X1 U5573 ( .A(n5612), .B(n5604), .ZN(n8555) );
  NAND2_X1 U5574 ( .A1(n4543), .A2(n4542), .ZN(n6805) );
  NAND2_X1 U5575 ( .A1(n4531), .A2(n4529), .ZN(n4542) );
  NAND2_X1 U5576 ( .A1(n4530), .A2(n4312), .ZN(n4529) );
  XNOR2_X1 U5577 ( .A(n5487), .B(n5486), .ZN(n7805) );
  OAI21_X1 U5578 ( .B1(n4595), .B2(n4591), .A(n4589), .ZN(n5462) );
  NAND2_X1 U5579 ( .A1(n4595), .A2(n5420), .ZN(n4594) );
  NAND2_X1 U5580 ( .A1(n5857), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5858) );
  NAND2_X1 U5581 ( .A1(n4596), .A2(n5332), .ZN(n5350) );
  NAND2_X1 U5582 ( .A1(n4608), .A2(n4607), .ZN(n5289) );
  NAND2_X1 U5583 ( .A1(n4608), .A2(n5249), .ZN(n5267) );
  XNOR2_X1 U5584 ( .A(n5225), .B(n5224), .ZN(n6923) );
  NAND2_X1 U5585 ( .A1(n4742), .A2(n5151), .ZN(n5174) );
  NAND2_X1 U5586 ( .A1(n4744), .A2(n4743), .ZN(n4742) );
  AND2_X1 U5587 ( .A1(n6047), .A2(n6060), .ZN(n7011) );
  XNOR2_X1 U5588 ( .A(n5125), .B(n5126), .ZN(n6637) );
  NAND2_X1 U5589 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), .ZN(
        n4556) );
  AOI21_X1 U5590 ( .B1(n4704), .B2(n4707), .A(n5460), .ZN(n4702) );
  NAND2_X1 U5591 ( .A1(n4725), .A2(n4287), .ZN(n7742) );
  NAND2_X1 U5592 ( .A1(n7230), .A2(n5078), .ZN(n8108) );
  NAND2_X1 U5593 ( .A1(n4710), .A2(n5281), .ZN(n8124) );
  OR2_X1 U5594 ( .A1(n5548), .A2(n5542), .ZN(n5552) );
  NAND2_X1 U5595 ( .A1(n5548), .A2(n5547), .ZN(n5551) );
  NAND2_X1 U5596 ( .A1(n5124), .A2(n5123), .ZN(n7613) );
  NAND2_X1 U5597 ( .A1(n5124), .A2(n4401), .ZN(n7615) );
  NAND2_X1 U5598 ( .A1(n8121), .A2(n5313), .ZN(n8183) );
  NAND2_X1 U5599 ( .A1(n5323), .A2(n5322), .ZN(n8509) );
  NAND2_X1 U5600 ( .A1(n7615), .A2(n5150), .ZN(n7620) );
  OAI21_X1 U5601 ( .B1(n8133), .B2(n4718), .A(n4716), .ZN(n8200) );
  OR2_X1 U5602 ( .A1(n6979), .A2(n9756), .ZN(n8221) );
  AND2_X1 U5603 ( .A1(n8040), .A2(n4890), .ZN(n6898) );
  NAND2_X1 U5604 ( .A1(n4703), .A2(n4279), .ZN(n8217) );
  NAND2_X1 U5605 ( .A1(n8161), .A2(n4708), .ZN(n4703) );
  OAI21_X1 U5606 ( .B1(n8161), .B2(n4707), .A(n4704), .ZN(n8215) );
  INV_X1 U5607 ( .A(n8189), .ZN(n8214) );
  AND4_X1 U5608 ( .A1(n5191), .A2(n5190), .A3(n5189), .A4(n5188), .ZN(n7818)
         );
  OR2_X1 U5609 ( .A1(n6979), .A2(n9758), .ZN(n8220) );
  NAND2_X1 U5610 ( .A1(n7461), .A2(n5540), .ZN(n8207) );
  XNOR2_X1 U5611 ( .A(n5516), .B(P2_IR_REG_22__SCAN_IN), .ZN(n5830) );
  OR2_X1 U5612 ( .A1(n5643), .A2(n5642), .ZN(n4575) );
  AND2_X1 U5613 ( .A1(n5559), .A2(n5558), .ZN(n6758) );
  NAND2_X1 U5614 ( .A1(n5503), .A2(n5502), .ZN(n8299) );
  OR2_X1 U5615 ( .A1(n5564), .A2(n5553), .ZN(n5503) );
  XNOR2_X1 U5616 ( .A(n4487), .B(P2_IR_REG_1__SCAN_IN), .ZN(n7340) );
  NAND2_X1 U5617 ( .A1(n9689), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4487) );
  INV_X1 U5618 ( .A(n4476), .ZN(n7990) );
  INV_X1 U5619 ( .A(n4482), .ZN(n7965) );
  INV_X1 U5620 ( .A(n4480), .ZN(n7931) );
  INV_X1 U5621 ( .A(n4478), .ZN(n7920) );
  INV_X1 U5622 ( .A(n4853), .ZN(n4729) );
  AND2_X1 U5623 ( .A1(n5181), .A2(n5226), .ZN(n7768) );
  AND2_X1 U5624 ( .A1(n5614), .A2(n5613), .ZN(n8459) );
  AOI21_X1 U5625 ( .B1(n8461), .B2(n8450), .A(n8077), .ZN(n4366) );
  NAND2_X1 U5626 ( .A1(n8071), .A2(n4379), .ZN(n4378) );
  NAND2_X1 U5627 ( .A1(n8341), .A2(n5752), .ZN(n8333) );
  NOR2_X1 U5628 ( .A1(n8355), .A2(n8059), .ZN(n8345) );
  OR2_X1 U5629 ( .A1(n8355), .A2(n4809), .ZN(n8343) );
  NAND2_X1 U5630 ( .A1(n8359), .A2(n5748), .ZN(n8339) );
  NAND2_X1 U5631 ( .A1(n4787), .A2(n4790), .ZN(n8390) );
  NAND2_X1 U5632 ( .A1(n8422), .A2(n4791), .ZN(n4787) );
  NAND2_X1 U5633 ( .A1(n4793), .A2(n4791), .ZN(n8508) );
  NAND2_X1 U5634 ( .A1(n4793), .A2(n4794), .ZN(n8419) );
  NAND2_X1 U5635 ( .A1(n8442), .A2(n5726), .ZN(n8423) );
  NAND2_X1 U5636 ( .A1(n5298), .A2(n5297), .ZN(n8515) );
  AND2_X1 U5637 ( .A1(n5584), .A2(n5721), .ZN(n4823) );
  NAND2_X1 U5638 ( .A1(n7784), .A2(n7783), .ZN(n7787) );
  NAND2_X1 U5639 ( .A1(n7660), .A2(n5582), .ZN(n7752) );
  NAND2_X1 U5640 ( .A1(n7659), .A2(n7658), .ZN(n7758) );
  AND2_X1 U5641 ( .A1(n7578), .A2(n7577), .ZN(n7580) );
  NAND2_X1 U5642 ( .A1(n9696), .A2(n7554), .ZN(n7556) );
  OAI21_X1 U5643 ( .B1(n7208), .B2(n4688), .A(n4685), .ZN(n9691) );
  NAND2_X1 U5644 ( .A1(n4691), .A2(n5804), .ZN(n7258) );
  NAND2_X1 U5645 ( .A1(n7208), .A2(n5803), .ZN(n4691) );
  NAND2_X1 U5646 ( .A1(n6906), .A2(n6905), .ZN(n7167) );
  NAND2_X1 U5647 ( .A1(n6958), .A2(n5648), .ZN(n4660) );
  NOR2_X1 U5648 ( .A1(n4662), .A2(n7112), .ZN(n4661) );
  NAND2_X1 U5649 ( .A1(n6874), .A2(n4813), .ZN(n7113) );
  OR2_X1 U5650 ( .A1(n6762), .A2(n9707), .ZN(n7461) );
  INV_X1 U5651 ( .A(n9999), .ZN(n8450) );
  NAND2_X1 U5652 ( .A1(n9794), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n4494) );
  OR2_X1 U5653 ( .A1(n8491), .A2(n9731), .ZN(n8496) );
  AND2_X1 U5654 ( .A1(n5826), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9714) );
  INV_X1 U5655 ( .A(n9709), .ZN(n9712) );
  INV_X1 U5656 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n4836) );
  NAND2_X1 U5657 ( .A1(n5511), .A2(n4867), .ZN(n7763) );
  INV_X1 U5658 ( .A(n5510), .ZN(n5511) );
  XNOR2_X1 U5659 ( .A(n5520), .B(n5519), .ZN(n7656) );
  INV_X1 U5660 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n5519) );
  INV_X1 U5661 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n7421) );
  INV_X1 U5662 ( .A(n5830), .ZN(n7419) );
  INV_X1 U5663 ( .A(n5821), .ZN(n7380) );
  INV_X1 U5664 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n9870) );
  INV_X1 U5665 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n7378) );
  INV_X1 U5666 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n4858) );
  NAND2_X1 U5667 ( .A1(n4857), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4859) );
  INV_X1 U5668 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n8050) );
  INV_X1 U5669 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n6972) );
  INV_X1 U5670 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n9884) );
  INV_X1 U5671 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n9887) );
  INV_X1 U5672 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n6684) );
  INV_X1 U5673 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n6640) );
  INV_X1 U5674 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n6635) );
  INV_X1 U5675 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n6625) );
  INV_X1 U5676 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n6607) );
  INV_X1 U5677 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n6600) );
  BUF_X1 U5678 ( .A(P2_IR_REG_0__SCAN_IN), .Z(n9689) );
  NAND2_X1 U5679 ( .A1(n6020), .A2(n6019), .ZN(n7505) );
  NAND2_X1 U5680 ( .A1(n8662), .A2(n6339), .ZN(n6858) );
  NAND2_X1 U5681 ( .A1(n4523), .A2(n8672), .ZN(n4528) );
  OR2_X1 U5682 ( .A1(n8675), .A2(n8673), .ZN(n4523) );
  AND2_X1 U5683 ( .A1(n6552), .A2(n8700), .ZN(n6553) );
  CLKBUF_X1 U5684 ( .A(n6747), .Z(n6748) );
  INV_X1 U5685 ( .A(n4783), .ZN(n8598) );
  AND4_X1 U5686 ( .A1(n6095), .A2(n6094), .A3(n6093), .A4(n6092), .ZN(n9260)
         );
  AND2_X1 U5687 ( .A1(n8696), .A2(n4777), .ZN(n8605) );
  NAND2_X1 U5688 ( .A1(n8604), .A2(n6455), .ZN(n8613) );
  AOI21_X1 U5689 ( .B1(n4521), .B2(n8673), .A(n4288), .ZN(n4518) );
  NAND2_X1 U5690 ( .A1(n4772), .A2(n4770), .ZN(n7695) );
  AND4_X1 U5691 ( .A1(n6027), .A2(n6026), .A3(n6025), .A4(n6024), .ZN(n9587)
         );
  NAND2_X1 U5692 ( .A1(n4776), .A2(n7383), .ZN(n7543) );
  NAND2_X1 U5693 ( .A1(n6555), .A2(n9613), .ZN(n8680) );
  AND4_X1 U5694 ( .A1(n5956), .A2(n5955), .A3(n5954), .A4(n5953), .ZN(n7294)
         );
  INV_X1 U5695 ( .A(n8690), .ZN(n8707) );
  NAND2_X1 U5696 ( .A1(n6557), .A2(n8993), .ZN(n8705) );
  NOR2_X1 U5697 ( .A1(n8684), .A2(n4779), .ZN(n4778) );
  INV_X1 U5698 ( .A(n4780), .ZN(n4779) );
  INV_X1 U5699 ( .A(n8682), .ZN(n8700) );
  INV_X1 U5700 ( .A(n8676), .ZN(n8710) );
  NAND2_X1 U5701 ( .A1(n8819), .A2(n8817), .ZN(n8818) );
  INV_X1 U5702 ( .A(n6817), .ZN(n8990) );
  INV_X1 U5703 ( .A(n9135), .ZN(n9004) );
  INV_X1 U5704 ( .A(n7294), .ZN(n9017) );
  INV_X1 U5705 ( .A(n7104), .ZN(n9020) );
  AND2_X1 U5706 ( .A1(n5914), .A2(n5913), .ZN(n5917) );
  NAND2_X1 U5707 ( .A1(n6791), .A2(n6792), .ZN(n6790) );
  NAND2_X1 U5708 ( .A1(n6719), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n4560) );
  NAND2_X1 U5709 ( .A1(n4294), .A2(n9465), .ZN(n9464) );
  NAND2_X1 U5710 ( .A1(n9464), .A2(n4557), .ZN(n9481) );
  NAND2_X1 U5711 ( .A1(n4559), .A2(n4558), .ZN(n4557) );
  INV_X1 U5712 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n4558) );
  INV_X1 U5713 ( .A(n9470), .ZN(n4559) );
  NAND2_X1 U5714 ( .A1(n9502), .A2(n4341), .ZN(n9518) );
  NAND2_X1 U5715 ( .A1(n9518), .A2(n9519), .ZN(n9517) );
  INV_X1 U5716 ( .A(n4565), .ZN(n9523) );
  INV_X1 U5717 ( .A(n4563), .ZN(n6941) );
  NOR2_X1 U5718 ( .A1(n7015), .A2(n7014), .ZN(n7594) );
  NOR2_X1 U5719 ( .A1(n7010), .A2(n4572), .ZN(n7015) );
  AND2_X1 U5720 ( .A1(n7011), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n4572) );
  NAND2_X1 U5721 ( .A1(n7600), .A2(n4362), .ZN(n9557) );
  OR2_X1 U5722 ( .A1(n7601), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n4362) );
  INV_X1 U5723 ( .A(n4569), .ZN(n7705) );
  NOR2_X1 U5724 ( .A1(n7712), .A2(n7711), .ZN(n7715) );
  OAI21_X1 U5725 ( .B1(n7598), .B2(n4567), .A(n4566), .ZN(n9022) );
  NAND2_X1 U5726 ( .A1(n4570), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n4567) );
  NAND2_X1 U5727 ( .A1(n7706), .A2(n4570), .ZN(n4566) );
  INV_X1 U5728 ( .A(n7708), .ZN(n4570) );
  INV_X1 U5729 ( .A(n7706), .ZN(n4568) );
  INV_X1 U5730 ( .A(n9543), .ZN(n9563) );
  AOI21_X1 U5731 ( .B1(n9042), .B2(P1_REG1_REG_17__SCAN_IN), .A(n9041), .ZN(
        n9571) );
  XNOR2_X1 U5732 ( .A(n5882), .B(n5881), .ZN(n9049) );
  INV_X1 U5733 ( .A(n9510), .ZN(n9574) );
  AOI21_X1 U5734 ( .B1(n9046), .B2(n9543), .A(n4360), .ZN(n4359) );
  NAND2_X1 U5735 ( .A1(n8720), .A2(n8719), .ZN(n9279) );
  NAND2_X1 U5736 ( .A1(n6232), .A2(n6231), .ZN(n9288) );
  NAND2_X1 U5737 ( .A1(n6219), .A2(n8867), .ZN(n9094) );
  NAND2_X1 U5738 ( .A1(n4630), .A2(n4629), .ZN(n9103) );
  OR2_X1 U5739 ( .A1(n6301), .A2(n4632), .ZN(n4629) );
  NAND2_X1 U5740 ( .A1(n4460), .A2(n8794), .ZN(n9123) );
  NAND2_X1 U5741 ( .A1(n4635), .A2(n4636), .ZN(n9115) );
  NAND2_X1 U5742 ( .A1(n6301), .A2(n4283), .ZN(n4635) );
  NAND2_X1 U5743 ( .A1(n9155), .A2(n8887), .ZN(n9133) );
  AND2_X1 U5744 ( .A1(n4637), .A2(n4640), .ZN(n9131) );
  NAND2_X1 U5745 ( .A1(n6301), .A2(n6300), .ZN(n4637) );
  AND2_X1 U5746 ( .A1(n6173), .A2(n6172), .ZN(n9149) );
  INV_X1 U5747 ( .A(n9613), .ZN(n9595) );
  AND2_X1 U5748 ( .A1(n6162), .A2(n6161), .ZN(n9173) );
  NAND2_X1 U5749 ( .A1(n9187), .A2(n9186), .ZN(n9188) );
  NAND2_X1 U5750 ( .A1(n6139), .A2(n8891), .ZN(n9198) );
  AND2_X1 U5751 ( .A1(n4624), .A2(n4625), .ZN(n9193) );
  NAND2_X1 U5752 ( .A1(n9204), .A2(n6297), .ZN(n4624) );
  NAND2_X1 U5753 ( .A1(n9268), .A2(n6292), .ZN(n9239) );
  NAND2_X1 U5754 ( .A1(n4642), .A2(n6286), .ZN(n7644) );
  NAND2_X1 U5755 ( .A1(n7673), .A2(n6282), .ZN(n4642) );
  NAND2_X1 U5756 ( .A1(n7180), .A2(n8734), .ZN(n7244) );
  AND2_X1 U5757 ( .A1(n7177), .A2(n6274), .ZN(n7243) );
  NAND2_X1 U5758 ( .A1(n5977), .A2(n5976), .ZN(n7182) );
  NAND2_X1 U5759 ( .A1(n9609), .A2(n6844), .ZN(n9271) );
  NAND2_X1 U5760 ( .A1(n6990), .A2(n6270), .ZN(n7062) );
  INV_X1 U5761 ( .A(n9605), .ZN(n9599) );
  NAND2_X1 U5762 ( .A1(n6835), .A2(n6268), .ZN(n7093) );
  AND3_X1 U5763 ( .A1(n6587), .A2(P1_STATE_REG_SCAN_IN), .A3(n7572), .ZN(n9649) );
  INV_X1 U5764 ( .A(n5899), .ZN(n9390) );
  NAND2_X1 U5765 ( .A1(n5870), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5867) );
  INV_X1 U5766 ( .A(n8987), .ZN(n8942) );
  INV_X1 U5767 ( .A(n9049), .ZN(n9248) );
  INV_X1 U5768 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n6925) );
  INV_X1 U5769 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n6745) );
  OR2_X1 U5770 ( .A1(n6076), .A2(n6075), .ZN(n7599) );
  INV_X1 U5771 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n6733) );
  INV_X1 U5772 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n6638) );
  XNOR2_X1 U5773 ( .A(n5062), .B(n5050), .ZN(n6619) );
  AND2_X1 U5774 ( .A1(n6002), .A2(n5993), .ZN(n9516) );
  NOR2_X1 U5775 ( .A1(n6597), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9383) );
  XNOR2_X1 U5776 ( .A(n5972), .B(P1_IR_REG_6__SCAN_IN), .ZN(n9490) );
  NAND2_X1 U5777 ( .A1(n4581), .A2(n4969), .ZN(n4992) );
  NAND2_X1 U5778 ( .A1(n4966), .A2(n4965), .ZN(n4581) );
  AND2_X1 U5779 ( .A1(n5963), .A2(n5962), .ZN(n9478) );
  XNOR2_X1 U5780 ( .A(n4922), .B(n4946), .ZN(n6605) );
  NOR2_X1 U5781 ( .A1(n7535), .A2(n10021), .ZN(n9840) );
  AOI21_X1 U5782 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(P1_ADDR_REG_10__SCAN_IN), 
        .A(n9838), .ZN(n9837) );
  NOR2_X1 U5783 ( .A1(n9837), .A2(n9836), .ZN(n9835) );
  AOI21_X1 U5784 ( .B1(P2_ADDR_REG_11__SCAN_IN), .B2(P1_ADDR_REG_11__SCAN_IN), 
        .A(n9835), .ZN(n9834) );
  OAI21_X1 U5785 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(P1_ADDR_REG_12__SCAN_IN), 
        .A(n9832), .ZN(n9830) );
  OAI21_X1 U5786 ( .B1(n8031), .B2(n5295), .A(n4483), .ZN(n8032) );
  NAND2_X1 U5787 ( .A1(n4486), .A2(n4484), .ZN(n4483) );
  OAI21_X1 U5788 ( .B1(n8454), .B2(n9780), .A(n4495), .ZN(n8535) );
  AOI21_X1 U5789 ( .B1(n4383), .B2(n4372), .A(n4371), .ZN(P2_U3549) );
  AND2_X1 U5790 ( .A1(n4381), .A2(n9808), .ZN(n4371) );
  NAND2_X1 U5791 ( .A1(n8462), .A2(n4381), .ZN(n4373) );
  OAI21_X1 U5792 ( .B1(n8454), .B2(n4493), .A(n4491), .ZN(P2_U3519) );
  NAND2_X1 U5793 ( .A1(n9796), .A2(n9727), .ZN(n4493) );
  INV_X1 U5794 ( .A(n4492), .ZN(n4491) );
  OAI21_X1 U5795 ( .B1(n4495), .B2(n9794), .A(n4494), .ZN(n4492) );
  AND2_X1 U5796 ( .A1(n6307), .A2(n6306), .ZN(n4824) );
  NAND2_X1 U5797 ( .A1(n9365), .A2(n9672), .ZN(n4467) );
  INV_X1 U5798 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n4466) );
  AND2_X1 U5799 ( .A1(n5891), .A2(n5899), .ZN(n4265) );
  OR2_X1 U5800 ( .A1(n9329), .A2(n9214), .ZN(n4266) );
  INV_X2 U5801 ( .A(n5030), .ZN(n4982) );
  NAND3_X1 U5802 ( .A1(n5917), .A2(n5916), .A3(n5915), .ZN(n6314) );
  AND2_X1 U5803 ( .A1(n4677), .A2(n5748), .ZN(n4267) );
  AND2_X1 U5804 ( .A1(n6275), .A2(n6274), .ZN(n4268) );
  AND2_X1 U5805 ( .A1(n4502), .A2(n8296), .ZN(n4269) );
  XNOR2_X1 U5806 ( .A(P2_REG2_REG_19__SCAN_IN), .B(n8021), .ZN(n4270) );
  NAND2_X1 U5807 ( .A1(n5173), .A2(n4743), .ZN(n4271) );
  NAND2_X1 U5808 ( .A1(n9276), .A2(n8721), .ZN(n4272) );
  OR2_X1 U5809 ( .A1(n6590), .A2(n4648), .ZN(n4273) );
  AND2_X1 U5810 ( .A1(n8064), .A2(n5595), .ZN(n8281) );
  NAND2_X1 U5811 ( .A1(n4773), .A2(n5848), .ZN(n5958) );
  OR2_X1 U5812 ( .A1(n9313), .A2(n9164), .ZN(n8887) );
  INV_X1 U5813 ( .A(n8887), .ZN(n4465) );
  AND2_X1 U5814 ( .A1(n4269), .A2(n4501), .ZN(n4274) );
  AND2_X1 U5815 ( .A1(n9329), .A2(n8592), .ZN(n8823) );
  AND2_X1 U5816 ( .A1(n4549), .A2(n4548), .ZN(n4276) );
  AND2_X1 U5817 ( .A1(n4378), .A2(n9793), .ZN(n4277) );
  XNOR2_X1 U5818 ( .A(n4859), .B(n4858), .ZN(n5506) );
  INV_X1 U5819 ( .A(n8890), .ZN(n4425) );
  INV_X1 U5820 ( .A(n6522), .ZN(n6510) );
  INV_X1 U5821 ( .A(n7648), .ZN(n9435) );
  XNOR2_X1 U5822 ( .A(n4556), .B(P1_IR_REG_1__SCAN_IN), .ZN(n6651) );
  NAND2_X1 U5823 ( .A1(n6864), .A2(n7462), .ZN(n5794) );
  NOR2_X1 U5824 ( .A1(n5887), .A2(P1_IR_REG_29__SCAN_IN), .ZN(n5889) );
  OR2_X1 U5825 ( .A1(n8466), .A2(n8097), .ZN(n4278) );
  OR2_X1 U5826 ( .A1(n5442), .A2(n8158), .ZN(n4279) );
  OR2_X1 U5827 ( .A1(n4974), .A2(n4973), .ZN(n4280) );
  AND4_X1 U5828 ( .A1(n4821), .A2(n4830), .A3(n4829), .A4(n4828), .ZN(n4281)
         );
  AND2_X1 U5829 ( .A1(n8453), .A2(n9726), .ZN(n4282) );
  AND2_X1 U5830 ( .A1(n4639), .A2(n6300), .ZN(n4283) );
  NAND2_X1 U5831 ( .A1(n8071), .A2(n4278), .ZN(n4699) );
  AND2_X1 U5832 ( .A1(n4825), .A2(n5721), .ZN(n4284) );
  OR2_X1 U5833 ( .A1(n6278), .A2(n4658), .ZN(n4285) );
  AND2_X1 U5834 ( .A1(n7579), .A2(n7577), .ZN(n4286) );
  OR2_X1 U5835 ( .A1(n5172), .A2(n5171), .ZN(n4287) );
  NAND2_X1 U5836 ( .A1(n4973), .A2(n4833), .ZN(n4862) );
  AND2_X1 U5837 ( .A1(n6475), .A2(n6474), .ZN(n4288) );
  INV_X1 U5838 ( .A(n7232), .ZN(n4396) );
  NAND2_X1 U5839 ( .A1(n4973), .A2(n4281), .ZN(n4289) );
  OR3_X1 U5840 ( .A1(n9071), .A2(n8935), .A3(n8802), .ZN(n4290) );
  AND2_X1 U5841 ( .A1(n8008), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n4291) );
  OAI211_X1 U5842 ( .C1(n6014), .C2(n6601), .A(n5949), .B(n5948), .ZN(n6996)
         );
  INV_X1 U5843 ( .A(n4417), .ZN(n4416) );
  NAND2_X1 U5844 ( .A1(n4418), .A2(n4425), .ZN(n4417) );
  AND3_X1 U5845 ( .A1(n4973), .A2(n4814), .A3(n4392), .ZN(n4292) );
  INV_X1 U5846 ( .A(n8794), .ZN(n4463) );
  INV_X1 U5847 ( .A(n5803), .ZN(n4687) );
  XOR2_X1 U5848 ( .A(n6434), .B(n6544), .Z(n4293) );
  AND2_X1 U5849 ( .A1(n4561), .A2(n4560), .ZN(n4294) );
  INV_X1 U5850 ( .A(n8344), .ZN(n4677) );
  NAND2_X1 U5851 ( .A1(n6141), .A2(n6140), .ZN(n9329) );
  INV_X1 U5852 ( .A(n9329), .ZN(n4548) );
  OR2_X1 U5853 ( .A1(n9386), .A2(n5899), .ZN(n5912) );
  AND2_X1 U5854 ( .A1(n4791), .A2(n8057), .ZN(n4295) );
  AND2_X1 U5855 ( .A1(n9310), .A2(n9125), .ZN(n4296) );
  NOR3_X1 U5856 ( .A1(P2_IR_REG_23__SCAN_IN), .A2(P2_IR_REG_22__SCAN_IN), .A3(
        P2_IR_REG_24__SCAN_IN), .ZN(n4297) );
  NAND2_X1 U5857 ( .A1(n4508), .A2(n6504), .ZN(n8574) );
  INV_X1 U5858 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n4855) );
  AND2_X1 U5859 ( .A1(n6790), .A2(n4364), .ZN(n4298) );
  INV_X1 U5860 ( .A(n7045), .ZN(n4505) );
  OAI21_X1 U5861 ( .B1(n6923), .B2(n4753), .A(n4750), .ZN(n8920) );
  OR2_X1 U5862 ( .A1(n8805), .A2(n8856), .ZN(n4299) );
  NAND2_X1 U5863 ( .A1(n6123), .A2(n6122), .ZN(n9339) );
  AND2_X1 U5864 ( .A1(n9329), .A2(n9214), .ZN(n4300) );
  OR2_X1 U5865 ( .A1(n7820), .A2(n8234), .ZN(n4301) );
  NOR2_X1 U5866 ( .A1(n7691), .A2(n9009), .ZN(n4302) );
  AND2_X1 U5867 ( .A1(n6139), .A2(n4746), .ZN(n4303) );
  AND2_X1 U5868 ( .A1(n4538), .A2(n6446), .ZN(n4304) );
  AND2_X1 U5869 ( .A1(n4697), .A2(n4693), .ZN(n4305) );
  INV_X1 U5870 ( .A(n4555), .ZN(n9108) );
  NOR2_X1 U5871 ( .A1(n9300), .A2(n9116), .ZN(n4555) );
  AND2_X1 U5872 ( .A1(n7785), .A2(n7783), .ZN(n4306) );
  AND2_X1 U5873 ( .A1(n4413), .A2(n4414), .ZN(n4307) );
  INV_X1 U5874 ( .A(n6268), .ZN(n4613) );
  NAND2_X1 U5875 ( .A1(n5453), .A2(n5452), .ZN(n8477) );
  AND2_X1 U5876 ( .A1(n9347), .A2(n9234), .ZN(n4308) );
  INV_X1 U5877 ( .A(n4504), .ZN(n8374) );
  NOR2_X1 U5878 ( .A1(n8391), .A2(n8497), .ZN(n4504) );
  AND2_X1 U5879 ( .A1(n8509), .A2(n8426), .ZN(n4309) );
  NOR2_X1 U5880 ( .A1(n8269), .A2(n5637), .ZN(n4310) );
  AND2_X1 U5881 ( .A1(n7555), .A2(n7554), .ZN(n4311) );
  NAND2_X1 U5882 ( .A1(n6151), .A2(n6150), .ZN(n9324) );
  OR2_X1 U5883 ( .A1(n4435), .A2(n9380), .ZN(n4312) );
  INV_X1 U5884 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n4435) );
  AND3_X1 U5885 ( .A1(n4999), .A2(n4998), .A3(n4997), .ZN(n7436) );
  INV_X1 U5886 ( .A(n8853), .ZN(n9093) );
  AND2_X1 U5887 ( .A1(n8869), .A2(n8803), .ZN(n8853) );
  INV_X1 U5888 ( .A(n4724), .ZN(n4723) );
  NAND2_X1 U5889 ( .A1(n4287), .A2(n4728), .ZN(n4724) );
  NOR2_X1 U5890 ( .A1(n8530), .A2(n7801), .ZN(n4313) );
  NOR2_X1 U5891 ( .A1(n5348), .A2(n5347), .ZN(n4314) );
  NOR2_X1 U5892 ( .A1(n9182), .A2(n9165), .ZN(n4315) );
  INV_X1 U5893 ( .A(n4423), .ZN(n4422) );
  NAND2_X1 U5894 ( .A1(n8878), .A2(n4424), .ZN(n4423) );
  NAND3_X1 U5895 ( .A1(n5179), .A2(n5176), .A3(n4854), .ZN(n4316) );
  NAND2_X1 U5896 ( .A1(n8502), .A2(n8410), .ZN(n4317) );
  NOR2_X1 U5897 ( .A1(n5417), .A2(n5416), .ZN(n4318) );
  OR2_X1 U5898 ( .A1(n5871), .A2(P1_IR_REG_24__SCAN_IN), .ZN(n4319) );
  OR2_X1 U5899 ( .A1(n4730), .A2(n4316), .ZN(n4320) );
  AND2_X1 U5900 ( .A1(n8742), .A2(n8744), .ZN(n8832) );
  AND2_X1 U5901 ( .A1(n5054), .A2(n5053), .ZN(n4321) );
  NOR2_X1 U5902 ( .A1(n9304), .A2(n9004), .ZN(n4322) );
  NOR2_X1 U5903 ( .A1(n5106), .A2(n5105), .ZN(n4323) );
  AND2_X1 U5904 ( .A1(n4488), .A2(n8925), .ZN(n4324) );
  AND2_X1 U5905 ( .A1(n4286), .A2(n7757), .ZN(n4325) );
  NOR2_X1 U5906 ( .A1(n9112), .A2(n9095), .ZN(n4326) );
  AND2_X1 U5907 ( .A1(n5175), .A2(n5157), .ZN(n5173) );
  OR2_X1 U5908 ( .A1(n4638), .A2(n4296), .ZN(n4327) );
  OR2_X1 U5909 ( .A1(n6296), .A2(n4300), .ZN(n4328) );
  INV_X1 U5910 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n4731) );
  OR2_X1 U5911 ( .A1(n9300), .A2(n9126), .ZN(n4329) );
  AND2_X1 U5912 ( .A1(n6160), .A2(n4454), .ZN(n4330) );
  AND2_X1 U5913 ( .A1(n6271), .A2(n6270), .ZN(n4331) );
  AND2_X1 U5914 ( .A1(n4538), .A2(n8698), .ZN(n4332) );
  AND2_X1 U5915 ( .A1(n6409), .A2(n7383), .ZN(n4333) );
  OR2_X1 U5916 ( .A1(n4440), .A2(n4443), .ZN(n4334) );
  AND2_X1 U5917 ( .A1(n4276), .A2(n9182), .ZN(n4335) );
  INV_X1 U5918 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n4736) );
  AND2_X1 U5919 ( .A1(n4272), .A2(n4439), .ZN(n4336) );
  AND2_X1 U5920 ( .A1(n4802), .A2(n7203), .ZN(n4337) );
  INV_X1 U5921 ( .A(n4699), .ZN(n4698) );
  NOR2_X1 U5922 ( .A1(n4785), .A2(n4784), .ZN(n4338) );
  INV_X1 U5923 ( .A(n6522), .ZN(n6538) );
  INV_X1 U5924 ( .A(n4912), .ZN(n5030) );
  NAND2_X1 U5925 ( .A1(n5493), .A2(n5492), .ZN(n8466) );
  INV_X1 U5926 ( .A(n8466), .ZN(n4501) );
  INV_X1 U5927 ( .A(n8814), .ZN(n4445) );
  NAND2_X1 U5928 ( .A1(n4655), .A2(n4654), .ZN(n9268) );
  AND2_X1 U5929 ( .A1(n9246), .A2(n4276), .ZN(n4339) );
  NAND2_X1 U5930 ( .A1(n6221), .A2(n6220), .ZN(n9293) );
  INV_X1 U5931 ( .A(n9293), .ZN(n4554) );
  AND2_X1 U5932 ( .A1(n7982), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n4340) );
  OR2_X1 U5933 ( .A1(n9498), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n4341) );
  OAI21_X1 U5934 ( .B1(n8435), .B2(n8055), .A(n8054), .ZN(n8422) );
  INV_X1 U5935 ( .A(n8891), .ZN(n4747) );
  OR2_X1 U5936 ( .A1(n7665), .A2(n7820), .ZN(n4342) );
  AND2_X1 U5937 ( .A1(n9490), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n4343) );
  NAND2_X1 U5938 ( .A1(n5387), .A2(n5386), .ZN(n8367) );
  INV_X1 U5939 ( .A(n8367), .ZN(n4503) );
  OR3_X1 U5940 ( .A1(n7683), .A2(n7648), .A3(n7691), .ZN(n4344) );
  NAND2_X1 U5941 ( .A1(n4772), .A2(n6422), .ZN(n7692) );
  OR2_X1 U5942 ( .A1(n7665), .A2(n4498), .ZN(n4345) );
  NAND2_X1 U5943 ( .A1(n6447), .A2(n6446), .ZN(n8696) );
  AND2_X1 U5944 ( .A1(n4569), .A2(n4568), .ZN(n4346) );
  NAND2_X1 U5945 ( .A1(n7784), .A2(n4306), .ZN(n8053) );
  AND2_X1 U5946 ( .A1(n4725), .A2(n4723), .ZN(n4347) );
  INV_X1 U5947 ( .A(n4551), .ZN(n9261) );
  NOR3_X1 U5948 ( .A1(n7683), .A2(n4553), .A3(n7648), .ZN(n4551) );
  AND2_X1 U5949 ( .A1(n5200), .A2(SI_14_), .ZN(n4348) );
  OR2_X1 U5950 ( .A1(n5287), .A2(n5286), .ZN(n4349) );
  AND2_X1 U5951 ( .A1(n5351), .A2(n5332), .ZN(n4350) );
  AND2_X1 U5952 ( .A1(n5247), .A2(n5288), .ZN(n4351) );
  OR2_X1 U5953 ( .A1(n5060), .A2(n4729), .ZN(n4352) );
  INV_X1 U5954 ( .A(n4640), .ZN(n4638) );
  INV_X1 U5955 ( .A(n6296), .ZN(n4625) );
  AND2_X2 U5956 ( .A1(n6786), .A2(n6785), .ZN(n9796) );
  AND2_X1 U5957 ( .A1(n6431), .A2(n6430), .ZN(n4353) );
  NAND2_X1 U5958 ( .A1(n6912), .A2(n5671), .ZN(n7168) );
  AND2_X1 U5959 ( .A1(n7357), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n4354) );
  NAND2_X1 U5960 ( .A1(n5137), .A2(n5136), .ZN(n9786) );
  INV_X1 U5961 ( .A(n9786), .ZN(n4489) );
  OR2_X1 U5962 ( .A1(n9672), .A2(n4466), .ZN(n4355) );
  INV_X1 U5963 ( .A(n7187), .ZN(n4547) );
  NAND2_X1 U5964 ( .A1(n7200), .A2(n7199), .ZN(n7402) );
  AND2_X1 U5965 ( .A1(n7355), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n4356) );
  INV_X1 U5966 ( .A(n4592), .ZN(n4591) );
  NOR2_X1 U5967 ( .A1(n5444), .A2(n4593), .ZN(n4592) );
  NOR2_X1 U5968 ( .A1(n7115), .A2(n4661), .ZN(n4357) );
  AND2_X1 U5969 ( .A1(n4592), .A2(n5461), .ZN(n4358) );
  INV_X1 U5970 ( .A(n9727), .ZN(n9780) );
  INV_X1 U5971 ( .A(n9045), .ZN(n4360) );
  INV_X1 U5972 ( .A(n8901), .ZN(n4446) );
  NAND2_X1 U5973 ( .A1(n6656), .A2(n6657), .ZN(n4561) );
  INV_X1 U5974 ( .A(n6651), .ZN(n4648) );
  NOR2_X2 U5975 ( .A1(n4867), .A2(n4835), .ZN(n4838) );
  NAND2_X2 U5976 ( .A1(n4391), .A2(n4833), .ZN(n4867) );
  NAND2_X2 U5977 ( .A1(n5113), .A2(n5112), .ZN(n8208) );
  INV_X1 U5978 ( .A(n5802), .ZN(n4686) );
  NAND2_X1 U5979 ( .A1(n4382), .A2(n4383), .ZN(n8537) );
  NAND2_X1 U5980 ( .A1(n4682), .A2(n4684), .ZN(n7559) );
  INV_X1 U5981 ( .A(n4365), .ZN(n8078) );
  OAI21_X1 U5982 ( .B1(n8463), .B2(n10001), .A(n4366), .ZN(n4365) );
  INV_X1 U5983 ( .A(n5153), .ZN(n4744) );
  NAND3_X1 U5984 ( .A1(n6286), .A2(n4645), .A3(n4368), .ZN(n4367) );
  NAND2_X1 U5985 ( .A1(n6301), .A2(n4628), .ZN(n4627) );
  NAND2_X1 U5986 ( .A1(n4467), .A2(n4355), .ZN(P1_U3520) );
  XNOR2_X2 U5987 ( .A(n5174), .B(n5173), .ZN(n6730) );
  INV_X1 U5988 ( .A(n4469), .ZN(n4468) );
  NOR2_X1 U5989 ( .A1(n9067), .A2(n6302), .ZN(n6303) );
  NAND2_X1 U5990 ( .A1(n4599), .A2(n4597), .ZN(n5225) );
  NAND2_X2 U5991 ( .A1(n5391), .A2(n5390), .ZN(n5425) );
  NAND2_X1 U5992 ( .A1(n5331), .A2(n5330), .ZN(n4596) );
  AND2_X2 U5993 ( .A1(n4947), .A2(n4369), .ZN(n4966) );
  NAND2_X1 U5994 ( .A1(n9286), .A2(n4468), .ZN(n9365) );
  NAND2_X1 U5995 ( .A1(n4594), .A2(n5423), .ZN(n5445) );
  NAND2_X1 U5996 ( .A1(n5355), .A2(n5354), .ZN(n5379) );
  MUX2_X1 U5997 ( .A(n4921), .B(n6604), .S(n6596), .Z(n4940) );
  NAND2_X1 U5998 ( .A1(n4627), .A2(n4626), .ZN(n9088) );
  OAI21_X1 U5999 ( .B1(n9287), .B2(n9426), .A(n9285), .ZN(n4469) );
  NOR2_X1 U6000 ( .A1(n9068), .A2(n9069), .ZN(n9067) );
  AND2_X1 U6001 ( .A1(n8463), .A2(n8462), .ZN(n4382) );
  NOR2_X1 U6002 ( .A1(n4374), .A2(n4373), .ZN(n4372) );
  INV_X1 U6003 ( .A(n8463), .ZN(n4374) );
  NAND3_X1 U6004 ( .A1(n4376), .A2(n4277), .A3(n4375), .ZN(n4383) );
  NAND3_X1 U6005 ( .A1(n4376), .A2(n4378), .A3(n4375), .ZN(n8464) );
  NAND2_X1 U6006 ( .A1(n4337), .A2(n7200), .ZN(n4385) );
  NAND3_X1 U6007 ( .A1(n4389), .A2(n4393), .A3(n4387), .ZN(n4870) );
  NAND3_X1 U6008 ( .A1(n4292), .A2(n4390), .A3(P2_IR_REG_27__SCAN_IN), .ZN(
        n4389) );
  AND2_X2 U6009 ( .A1(n4973), .A2(n4814), .ZN(n4391) );
  INV_X2 U6010 ( .A(n4990), .ZN(n5633) );
  NAND2_X2 U6011 ( .A1(n4885), .A2(n6596), .ZN(n4990) );
  NAND2_X2 U6012 ( .A1(n5828), .A2(n5560), .ZN(n4885) );
  NAND2_X1 U6013 ( .A1(n6611), .A2(n5633), .ZN(n5022) );
  NAND2_X1 U6014 ( .A1(n4398), .A2(n5124), .ZN(n4399) );
  NAND2_X1 U6015 ( .A1(n4403), .A2(n4404), .ZN(n5375) );
  OAI21_X2 U6016 ( .B1(n6619), .B2(n4990), .A(n4321), .ZN(n8142) );
  NAND2_X1 U6017 ( .A1(n4411), .A2(n4412), .ZN(n8786) );
  NAND2_X1 U6018 ( .A1(n8789), .A2(n4414), .ZN(n4411) );
  NAND2_X1 U6019 ( .A1(n8806), .A2(n4336), .ZN(n4438) );
  NAND2_X1 U6020 ( .A1(n8722), .A2(n8908), .ZN(n8723) );
  NAND2_X1 U6021 ( .A1(n5940), .A2(n8957), .ZN(n8722) );
  INV_X1 U6022 ( .A(n5912), .ZN(n5921) );
  INV_X1 U6023 ( .A(n4452), .ZN(n4451) );
  OAI21_X1 U6024 ( .B1(n5912), .B2(n6829), .A(n4453), .ZN(n4452) );
  OAI21_X1 U6025 ( .B1(n9212), .B2(n4456), .A(n4330), .ZN(n9177) );
  NAND2_X1 U6026 ( .A1(n9155), .A2(n4461), .ZN(n4459) );
  OAI21_X1 U6027 ( .B1(n9155), .B2(n4463), .A(n4461), .ZN(n9122) );
  NAND3_X1 U6028 ( .A1(n8832), .A2(n8734), .A3(n7180), .ZN(n4472) );
  NAND2_X1 U6029 ( .A1(n4472), .A2(n8742), .ZN(n9585) );
  MUX2_X1 U6030 ( .A(n6693), .B(P2_REG1_REG_1__SCAN_IN), .S(n7340), .Z(n6695)
         );
  NAND3_X1 U6031 ( .A1(n6072), .A2(n4338), .A3(n5866), .ZN(n5887) );
  OR2_X2 U6032 ( .A1(n7260), .A2(n8208), .ZN(n9698) );
  NAND2_X1 U6033 ( .A1(n8268), .A2(n8459), .ZN(n8455) );
  INV_X1 U6034 ( .A(n4497), .ZN(n8437) );
  NOR2_X2 U6035 ( .A1(n8428), .A2(n8509), .ZN(n8412) );
  NOR2_X2 U6036 ( .A1(n4867), .A2(n4864), .ZN(n4868) );
  AOI21_X2 U6037 ( .B1(n8622), .B2(n8621), .A(n8620), .ZN(n8624) );
  INV_X1 U6038 ( .A(n7100), .ZN(n9650) );
  NAND3_X1 U6039 ( .A1(n5939), .A2(n4511), .A3(n4510), .ZN(n7100) );
  NAND2_X1 U6040 ( .A1(n4513), .A2(n4512), .ZN(n8561) );
  NAND2_X1 U6041 ( .A1(n4516), .A2(n7628), .ZN(n4513) );
  AOI21_X1 U6042 ( .B1(n4770), .B2(n4517), .A(n4353), .ZN(n4516) );
  OAI21_X1 U6043 ( .B1(n7628), .B2(n4515), .A(n4516), .ZN(n6437) );
  NAND2_X1 U6044 ( .A1(n8675), .A2(n4520), .ZN(n4519) );
  NAND2_X1 U6045 ( .A1(n8675), .A2(n8673), .ZN(n4527) );
  NOR2_X1 U6046 ( .A1(n4526), .A2(n4525), .ZN(n4524) );
  INV_X1 U6047 ( .A(n8673), .ZN(n4525) );
  NAND2_X1 U6048 ( .A1(n4528), .A2(n4527), .ZN(n8583) );
  NAND2_X1 U6049 ( .A1(n6072), .A2(n4532), .ZN(n4531) );
  AND2_X2 U6050 ( .A1(n5960), .A2(n5852), .ZN(n6072) );
  NAND2_X1 U6051 ( .A1(n8697), .A2(n4332), .ZN(n4534) );
  NAND2_X1 U6052 ( .A1(n4535), .A2(n4534), .ZN(n6464) );
  NAND2_X2 U6053 ( .A1(n5909), .A2(n6805), .ZN(n6590) );
  INV_X1 U6054 ( .A(n5894), .ZN(n4543) );
  NAND2_X1 U6055 ( .A1(n6838), .A2(n6836), .ZN(n7096) );
  NOR2_X1 U6056 ( .A1(n7683), .A2(n7691), .ZN(n7684) );
  MUX2_X1 U6057 ( .A(P1_REG2_REG_1__SCAN_IN), .B(n6855), .S(n6651), .Z(n6672)
         );
  XNOR2_X1 U6058 ( .A(n7704), .B(n7710), .ZN(n7598) );
  AOI21_X1 U6059 ( .B1(n5789), .B2(n5788), .A(n5820), .ZN(n5825) );
  NAND2_X1 U6060 ( .A1(n4573), .A2(n5833), .ZN(P2_U3244) );
  NAND2_X1 U6061 ( .A1(n4574), .A2(n5827), .ZN(n4573) );
  NAND3_X1 U6062 ( .A1(n4578), .A2(n4576), .A3(n4575), .ZN(n4574) );
  NAND2_X1 U6063 ( .A1(n5825), .A2(n4577), .ZN(n4576) );
  AND2_X1 U6064 ( .A1(n6777), .A2(n9715), .ZN(n4577) );
  NAND2_X1 U6065 ( .A1(n5824), .A2(n5823), .ZN(n4578) );
  INV_X1 U6066 ( .A(n5425), .ZN(n4595) );
  NAND2_X1 U6067 ( .A1(n5425), .A2(n4358), .ZN(n4585) );
  NAND2_X1 U6068 ( .A1(n4596), .A2(n4350), .ZN(n5355) );
  NAND2_X1 U6069 ( .A1(n5127), .A2(n4601), .ZN(n4599) );
  NAND2_X1 U6070 ( .A1(n5127), .A2(n5126), .ZN(n4600) );
  AOI21_X1 U6071 ( .B1(n5248), .B2(n4351), .A(n4605), .ZN(n5316) );
  NAND2_X1 U6072 ( .A1(n5248), .A2(n5247), .ZN(n4608) );
  NAND2_X1 U6073 ( .A1(n5017), .A2(n5016), .ZN(n5041) );
  NAND2_X1 U6074 ( .A1(n5489), .A2(n5488), .ZN(n5597) );
  OR2_X2 U6075 ( .A1(n7170), .A2(n8087), .ZN(n7412) );
  NAND2_X1 U6076 ( .A1(n4698), .A2(n4694), .ZN(n4693) );
  NAND2_X1 U6077 ( .A1(n5487), .A2(n5486), .ZN(n5489) );
  NAND2_X1 U6078 ( .A1(n5079), .A2(n4820), .ZN(n5081) );
  NAND2_X1 U6079 ( .A1(n9098), .A2(n8869), .ZN(n9072) );
  NOR2_X1 U6080 ( .A1(n9073), .A2(n8807), .ZN(n4749) );
  NOR2_X2 U6081 ( .A1(n7412), .A2(n8142), .ZN(n9764) );
  NOR2_X2 U6082 ( .A1(n9699), .A2(n7587), .ZN(n7588) );
  INV_X1 U6083 ( .A(n4610), .ZN(n4611) );
  OAI21_X1 U6084 ( .B1(n6267), .B2(n4613), .A(n7102), .ZN(n4610) );
  NAND2_X1 U6085 ( .A1(n4612), .A2(n4611), .ZN(n7092) );
  NAND2_X1 U6086 ( .A1(n9204), .A2(n4616), .ZN(n4615) );
  NAND2_X1 U6087 ( .A1(n9313), .A2(n9005), .ZN(n4640) );
  NAND2_X1 U6088 ( .A1(n7725), .A2(n8695), .ZN(n6288) );
  INV_X2 U6089 ( .A(n6590), .ZN(n6132) );
  NAND2_X1 U6090 ( .A1(n6990), .A2(n4331), .ZN(n7060) );
  XNOR2_X1 U6091 ( .A(n4660), .B(n7030), .ZN(n7032) );
  INV_X1 U6092 ( .A(n5578), .ZN(n4664) );
  NAND2_X1 U6093 ( .A1(n7662), .A2(n4671), .ZN(n4669) );
  NAND2_X1 U6094 ( .A1(n4669), .A2(n4670), .ZN(n7788) );
  OAI21_X2 U6095 ( .B1(n5584), .B2(n4680), .A(n4678), .ZN(n8407) );
  NAND2_X1 U6096 ( .A1(n7208), .A2(n4681), .ZN(n4684) );
  NAND3_X1 U6097 ( .A1(n5807), .A2(n4685), .A3(n4688), .ZN(n4683) );
  OAI21_X1 U6098 ( .B1(n8297), .B2(n8298), .A(n5594), .ZN(n8282) );
  NAND2_X1 U6099 ( .A1(n4692), .A2(n4305), .ZN(n5625) );
  NAND2_X1 U6100 ( .A1(n8297), .A2(n4695), .ZN(n4692) );
  NAND2_X1 U6101 ( .A1(n6898), .A2(n6897), .ZN(n6896) );
  XNOR2_X1 U6102 ( .A(n4889), .B(n4887), .ZN(n8041) );
  NAND2_X1 U6103 ( .A1(n8161), .A2(n4704), .ZN(n4701) );
  NAND2_X1 U6104 ( .A1(n4701), .A2(n4702), .ZN(n8095) );
  NAND2_X1 U6105 ( .A1(n4901), .A2(n4711), .ZN(n4925) );
  NAND2_X1 U6106 ( .A1(n8133), .A2(n4716), .ZN(n4712) );
  NAND2_X1 U6107 ( .A1(n4714), .A2(n4712), .ZN(n5124) );
  INV_X1 U6108 ( .A(n4732), .ZN(n4857) );
  OAI21_X1 U6109 ( .B1(n5153), .B2(n4271), .A(n4739), .ZN(n5201) );
  NAND2_X1 U6110 ( .A1(n6219), .A2(n4745), .ZN(n9098) );
  NAND2_X1 U6111 ( .A1(n4754), .A2(n4752), .ZN(n8924) );
  NOR2_X1 U6112 ( .A1(n9260), .A2(n4753), .ZN(n4752) );
  INV_X1 U6113 ( .A(n6088), .ZN(n4753) );
  NAND3_X1 U6114 ( .A1(n4757), .A2(P2_ADDR_REG_19__SCAN_IN), .A3(
        P1_ADDR_REG_19__SCAN_IN), .ZN(n4756) );
  NAND3_X1 U6115 ( .A1(n4761), .A2(n4760), .A3(n4759), .ZN(n4758) );
  NAND2_X1 U6116 ( .A1(n8642), .A2(n4763), .ZN(n4762) );
  NAND2_X1 U6117 ( .A1(n4762), .A2(n4765), .ZN(n6496) );
  NOR2_X2 U6118 ( .A1(n5946), .A2(n4774), .ZN(n5960) );
  NAND2_X1 U6119 ( .A1(n8624), .A2(n4782), .ZN(n4781) );
  OR2_X1 U6120 ( .A1(n8624), .A2(n6517), .ZN(n4783) );
  NAND2_X2 U6121 ( .A1(n4781), .A2(n4778), .ZN(n8688) );
  NAND3_X1 U6122 ( .A1(n4786), .A2(n6331), .A3(n6332), .ZN(n6747) );
  NAND2_X1 U6123 ( .A1(n6328), .A2(n6327), .ZN(n6332) );
  NAND2_X1 U6124 ( .A1(n6326), .A2(n6325), .ZN(n4786) );
  NAND2_X1 U6125 ( .A1(n4786), .A2(n6332), .ZN(n6746) );
  NAND2_X1 U6126 ( .A1(n6880), .A2(n4796), .ZN(n4795) );
  NAND2_X1 U6127 ( .A1(n6880), .A2(n6884), .ZN(n6906) );
  INV_X1 U6128 ( .A(n6884), .ZN(n4798) );
  AOI21_X1 U6129 ( .B1(n7578), .B2(n4325), .A(n4803), .ZN(n7760) );
  NAND2_X1 U6130 ( .A1(n4806), .A2(n4807), .ZN(n8324) );
  NAND2_X1 U6131 ( .A1(n4901), .A2(n4811), .ZN(n4949) );
  NOR2_X4 U6132 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n4901) );
  INV_X1 U6133 ( .A(n4812), .ZN(n7112) );
  NAND3_X1 U6134 ( .A1(n6874), .A2(n4813), .A3(n4812), .ZN(n6877) );
  NAND2_X1 U6135 ( .A1(n5575), .A2(n6864), .ZN(n4813) );
  INV_X2 U6136 ( .A(n5433), .ZN(n5504) );
  OR2_X1 U6137 ( .A1(n5912), .A2(n5911), .ZN(n5914) );
  NAND2_X1 U6138 ( .A1(n6867), .A2(n7045), .ZN(n6776) );
  OR2_X2 U6139 ( .A1(n8437), .A2(n8515), .ZN(n8428) );
  NAND2_X1 U6140 ( .A1(n6803), .A2(n6319), .ZN(n6328) );
  NAND2_X2 U6141 ( .A1(n6367), .A2(n6366), .ZN(n7078) );
  CLKBUF_X1 U6142 ( .A(n8662), .Z(n8663) );
  AND2_X1 U6143 ( .A1(n6779), .A2(n7045), .ZN(n6770) );
  NAND2_X2 U6144 ( .A1(n8632), .A2(n6354), .ZN(n7285) );
  INV_X1 U6145 ( .A(n9706), .ZN(n7564) );
  OR2_X1 U6146 ( .A1(n4554), .A2(n8713), .ZN(n4815) );
  AND2_X1 U6147 ( .A1(n8815), .A2(n8993), .ZN(n9233) );
  AND2_X1 U6148 ( .A1(n5108), .A2(n5086), .ZN(n4816) );
  NAND2_X1 U6149 ( .A1(n5906), .A2(n5905), .ZN(n9590) );
  AND2_X1 U6150 ( .A1(n8815), .A2(n9248), .ZN(n4817) );
  AND2_X1 U6151 ( .A1(n5885), .A2(n5884), .ZN(n4818) );
  AND2_X1 U6152 ( .A1(n5080), .A2(n5067), .ZN(n4820) );
  AND4_X1 U6153 ( .A1(n5179), .A2(n4736), .A3(n4856), .A4(n4855), .ZN(n4821)
         );
  NAND2_X1 U6154 ( .A1(n7564), .A2(n7029), .ZN(n8452) );
  INV_X1 U6155 ( .A(n7117), .ZN(n6864) );
  AND2_X1 U6156 ( .A1(n5724), .A2(n5726), .ZN(n4825) );
  NOR2_X1 U6157 ( .A1(n6285), .A2(n7674), .ZN(n4826) );
  INV_X2 U6158 ( .A(n9670), .ZN(n9672) );
  INV_X1 U6159 ( .A(n9676), .ZN(n9362) );
  INV_X1 U6160 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n5884) );
  NAND2_X1 U6161 ( .A1(n4310), .A2(n5623), .ZN(n5624) );
  INV_X1 U6162 ( .A(n8311), .ZN(n5592) );
  OR2_X1 U6163 ( .A1(n4864), .A2(P2_IR_REG_28__SCAN_IN), .ZN(n4835) );
  INV_X1 U6164 ( .A(n6750), .ZN(n6331) );
  INV_X1 U6165 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n5206) );
  INV_X1 U6166 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n9926) );
  NAND2_X1 U6167 ( .A1(n5593), .A2(n5592), .ZN(n8308) );
  INV_X1 U6168 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n5515) );
  INV_X1 U6169 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n4850) );
  INV_X1 U6170 ( .A(n6175), .ZN(n5843) );
  INV_X1 U6171 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n6089) );
  INV_X1 U6172 ( .A(n6142), .ZN(n5842) );
  INV_X1 U6173 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n6006) );
  OR2_X1 U6174 ( .A1(n6022), .A2(n6021), .ZN(n6034) );
  INV_X1 U6175 ( .A(n9069), .ZN(n9071) );
  NAND2_X1 U6176 ( .A1(n6013), .A2(n8835), .ZN(n7497) );
  INV_X1 U6177 ( .A(n7063), .ZN(n6271) );
  INV_X1 U6178 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n5885) );
  INV_X1 U6179 ( .A(SI_16_), .ZN(n5207) );
  INV_X1 U6180 ( .A(SI_13_), .ZN(n5154) );
  AND2_X1 U6181 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(P2_REG3_REG_9__SCAN_IN), 
        .ZN(n5098) );
  INV_X1 U6182 ( .A(n7154), .ZN(n5002) );
  AND2_X1 U6183 ( .A1(n5641), .A2(n6778), .ZN(n5642) );
  OR2_X1 U6184 ( .A1(n5437), .A2(n5436), .ZN(n5454) );
  INV_X1 U6185 ( .A(n4280), .ZN(n7345) );
  OR2_X1 U6186 ( .A1(n8470), .A2(n8229), .ZN(n8063) );
  AND2_X1 U6187 ( .A1(n5689), .A2(n5678), .ZN(n9749) );
  NAND2_X1 U6188 ( .A1(n5576), .A2(n7123), .ZN(n6955) );
  INV_X1 U6189 ( .A(n9707), .ZN(n6759) );
  INV_X1 U6190 ( .A(n6210), .ZN(n5845) );
  AND2_X1 U6191 ( .A1(n5898), .A2(n6248), .ZN(n9078) );
  NAND2_X1 U6192 ( .A1(n5842), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n6152) );
  OR2_X1 U6193 ( .A1(n6065), .A2(n6064), .ZN(n6079) );
  INV_X1 U6194 ( .A(n7090), .ZN(n6305) );
  NOR2_X1 U6195 ( .A1(n4826), .A2(n4302), .ZN(n6286) );
  NAND2_X1 U6196 ( .A1(n8997), .A2(n8951), .ZN(n6588) );
  INV_X1 U6197 ( .A(n8951), .ZN(n8861) );
  INV_X1 U6198 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n5872) );
  OR2_X1 U6199 ( .A1(n6029), .A2(P1_IR_REG_10__SCAN_IN), .ZN(n6042) );
  OR2_X1 U6200 ( .A1(n5403), .A2(n8102), .ZN(n5405) );
  OR2_X1 U6201 ( .A1(n5546), .A2(n5545), .ZN(n5547) );
  OR2_X1 U6202 ( .A1(n5114), .A2(n8203), .ZN(n5139) );
  INV_X1 U6203 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n7885) );
  XNOR2_X1 U6204 ( .A(n8470), .B(n8314), .ZN(n8298) );
  OR2_X1 U6205 ( .A1(n5139), .A2(n5138), .ZN(n5163) );
  NAND2_X1 U6206 ( .A1(n8074), .A2(n8073), .ZN(n8075) );
  AND2_X1 U6207 ( .A1(n5506), .A2(n6766), .ZN(n9727) );
  NAND2_X1 U6208 ( .A1(n6774), .A2(n6773), .ZN(n7563) );
  NAND2_X1 U6209 ( .A1(n5506), .A2(n5507), .ZN(n9741) );
  INV_X1 U6210 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n5523) );
  INV_X1 U6211 ( .A(n9126), .ZN(n9095) );
  INV_X1 U6212 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n8584) );
  AND2_X1 U6213 ( .A1(n6532), .A2(n6531), .ZN(n6575) );
  NAND2_X1 U6214 ( .A1(n5840), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n6114) );
  INV_X1 U6215 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n8614) );
  OAI211_X1 U6216 ( .C1(n8819), .C2(n4817), .A(n4822), .B(n8818), .ZN(n8820)
         );
  OR2_X1 U6217 ( .A1(n6135), .A2(n8584), .ZN(n6142) );
  NAND2_X1 U6218 ( .A1(n9149), .A2(n9164), .ZN(n6300) );
  INV_X1 U6219 ( .A(n9011), .ZN(n7634) );
  INV_X1 U6220 ( .A(n8832), .ZN(n6275) );
  INV_X1 U6221 ( .A(n9664), .ZN(n9340) );
  AND2_X1 U6222 ( .A1(n6819), .A2(n6818), .ZN(n9593) );
  OR2_X1 U6223 ( .A1(n9664), .A2(n9049), .ZN(n6735) );
  AND2_X1 U6224 ( .A1(n5249), .A2(n5210), .ZN(n5247) );
  INV_X1 U6225 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n9380) );
  AND2_X1 U6226 ( .A1(n5496), .A2(n5474), .ZN(n8294) );
  INV_X1 U6227 ( .A(n8221), .ZN(n8195) );
  AND2_X1 U6228 ( .A1(n5569), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8224) );
  INV_X1 U6229 ( .A(n7575), .ZN(n5827) );
  AND3_X1 U6230 ( .A1(n5441), .A2(n5440), .A3(n5439), .ZN(n8313) );
  AND4_X1 U6231 ( .A1(n5260), .A2(n5259), .A3(n5258), .A4(n5257), .ZN(n7828)
         );
  AND2_X1 U6232 ( .A1(n6700), .A2(n8072), .ZN(n8028) );
  NAND2_X1 U6233 ( .A1(n6694), .A2(n5828), .ZN(n9682) );
  INV_X1 U6234 ( .A(n9682), .ZN(n9679) );
  INV_X1 U6235 ( .A(n7461), .ZN(n9993) );
  INV_X1 U6236 ( .A(n7120), .ZN(n9702) );
  INV_X1 U6237 ( .A(n8415), .ZN(n9996) );
  AOI21_X1 U6238 ( .B1(n9708), .B2(n9711), .A(n9710), .ZN(n7025) );
  AND2_X1 U6239 ( .A1(n7563), .A2(n9741), .ZN(n9731) );
  INV_X1 U6240 ( .A(n9731), .ZN(n9793) );
  AND3_X1 U6241 ( .A1(n7027), .A2(n6765), .A3(n6764), .ZN(n6786) );
  AND2_X1 U6242 ( .A1(n6597), .A2(P2_U3152), .ZN(n8556) );
  INV_X1 U6243 ( .A(n8820), .ZN(n8946) );
  OR2_X1 U6244 ( .A1(n8689), .A2(n6212), .ZN(n6218) );
  AND4_X1 U6245 ( .A1(n6104), .A2(n6103), .A3(n6102), .A4(n6101), .ZN(n9243)
         );
  AND2_X1 U6246 ( .A1(n6655), .A2(n8992), .ZN(n9543) );
  INV_X1 U6247 ( .A(n7599), .ZN(n9554) );
  OR2_X1 U6248 ( .A1(n6654), .A2(n8992), .ZN(n9510) );
  INV_X1 U6249 ( .A(n9279), .ZN(n9061) );
  AND2_X1 U6250 ( .A1(n9609), .A2(n7095), .ZN(n9604) );
  AND2_X1 U6251 ( .A1(n9609), .A2(n7091), .ZN(n9583) );
  AND3_X1 U6252 ( .A1(n6813), .A2(n6812), .A3(n9649), .ZN(n6814) );
  AND2_X1 U6253 ( .A1(n9593), .A2(n7145), .ZN(n9426) );
  AND3_X1 U6254 ( .A1(n6812), .A2(n9643), .A3(n6263), .ZN(n6736) );
  INV_X1 U6255 ( .A(n7145), .ZN(n9669) );
  XNOR2_X1 U6256 ( .A(n5879), .B(n9857), .ZN(n7572) );
  AND2_X1 U6257 ( .A1(n6120), .A2(n6111), .ZN(n9042) );
  AND2_X1 U6258 ( .A1(n5522), .A2(n5521), .ZN(n6687) );
  INV_X1 U6259 ( .A(n5572), .ZN(n5573) );
  OR2_X1 U6260 ( .A1(n5549), .A2(n9726), .ZN(n8189) );
  INV_X1 U6261 ( .A(n8154), .ZN(n8426) );
  INV_X1 U6262 ( .A(n7828), .ZN(n8444) );
  OR2_X1 U6263 ( .A1(n7120), .A2(n9780), .ZN(n9999) );
  INV_X1 U6264 ( .A(n7564), .ZN(n10001) );
  AND2_X1 U6265 ( .A1(n7035), .A2(n7461), .ZN(n9706) );
  INV_X1 U6266 ( .A(n9810), .ZN(n9808) );
  AND2_X2 U6267 ( .A1(n6786), .A2(n7025), .ZN(n9810) );
  INV_X1 U6268 ( .A(n9796), .ZN(n9794) );
  NOR2_X1 U6269 ( .A1(n9708), .A2(n9707), .ZN(n9709) );
  INV_X1 U6270 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n9978) );
  INV_X1 U6271 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n6731) );
  AND2_X1 U6272 ( .A1(n6586), .A2(n7572), .ZN(n6641) );
  NAND2_X1 U6273 ( .A1(n6580), .A2(n6553), .ZN(n6572) );
  OR2_X1 U6274 ( .A1(n6556), .A2(n6560), .ZN(n8682) );
  INV_X1 U6275 ( .A(n7143), .ZN(n7299) );
  INV_X1 U6276 ( .A(n9096), .ZN(n9002) );
  INV_X1 U6277 ( .A(n9152), .ZN(n9179) );
  INV_X1 U6278 ( .A(n7307), .ZN(n9015) );
  OR2_X1 U6279 ( .A1(P1_U3083), .A2(n6641), .ZN(n9561) );
  OR2_X1 U6280 ( .A1(n9664), .A2(n5883), .ZN(n9613) );
  INV_X1 U6281 ( .A(n9440), .ZN(n9676) );
  AND2_X1 U6282 ( .A1(n6815), .A2(n6814), .ZN(n9440) );
  OR3_X1 U6283 ( .A1(n9355), .A2(n9354), .A3(n9353), .ZN(n9378) );
  NAND2_X1 U6284 ( .A1(n6815), .A2(n6736), .ZN(n9670) );
  INV_X1 U6285 ( .A(n9649), .ZN(n9645) );
  INV_X1 U6286 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n6949) );
  INV_X1 U6287 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n6686) );
  INV_X1 U6288 ( .A(n9383), .ZN(n7085) );
  NOR2_X1 U6289 ( .A1(n9840), .A2(n9839), .ZN(n9838) );
  AND2_X1 U6290 ( .A1(n6687), .A2(n9714), .ZN(P2_U3966) );
  AND2_X1 U6291 ( .A1(n6641), .A2(P1_STATE_REG_SCAN_IN), .ZN(P1_U4006) );
  NOR2_X1 U6292 ( .A1(P2_IR_REG_10__SCAN_IN), .A2(P2_IR_REG_9__SCAN_IN), .ZN(
        n4827) );
  NOR3_X1 U6293 ( .A1(P2_IR_REG_8__SCAN_IN), .A2(P2_IR_REG_20__SCAN_IN), .A3(
        P2_IR_REG_19__SCAN_IN), .ZN(n4828) );
  AND2_X2 U6294 ( .A1(n4281), .A2(n4831), .ZN(n4833) );
  AND2_X2 U6295 ( .A1(n4971), .A2(n4832), .ZN(n4973) );
  NAND2_X1 U6296 ( .A1(n4838), .A2(n4836), .ZN(n4841) );
  INV_X1 U6297 ( .A(n4838), .ZN(n4839) );
  NAND2_X1 U6298 ( .A1(n4839), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4840) );
  MUX2_X1 U6299 ( .A(P2_IR_REG_31__SCAN_IN), .B(n4840), .S(
        P2_IR_REG_29__SCAN_IN), .Z(n4842) );
  AND2_X4 U6300 ( .A1(n8034), .A2(n8557), .ZN(n5398) );
  NAND2_X1 U6301 ( .A1(n5398), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n4848) );
  AND2_X2 U6302 ( .A1(n8034), .A2(n4843), .ZN(n4912) );
  NAND2_X1 U6303 ( .A1(n4912), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n4847) );
  INV_X1 U6304 ( .A(n8034), .ZN(n4844) );
  NAND2_X1 U6305 ( .A1(n4913), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n4846) );
  NAND2_X1 U6306 ( .A1(n4935), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n4845) );
  NAND2_X1 U6307 ( .A1(n5051), .A2(n4850), .ZN(n5060) );
  NAND2_X1 U6308 ( .A1(n5090), .A2(n4851), .ZN(n4852) );
  OR2_X1 U6309 ( .A1(n7117), .A2(n6866), .ZN(n4889) );
  OR2_X2 U6310 ( .A1(n4868), .A2(n8552), .ZN(n4866) );
  INV_X1 U6311 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n4865) );
  XNOR2_X2 U6312 ( .A(n4866), .B(n4865), .ZN(n5560) );
  INV_X1 U6313 ( .A(n4868), .ZN(n4869) );
  NAND2_X1 U6314 ( .A1(n4870), .A2(n4869), .ZN(n5828) );
  NAND3_X1 U6315 ( .A1(n4262), .A2(SI_0_), .A3(P2_DATAO_REG_0__SCAN_IN), .ZN(
        n4872) );
  AND2_X1 U6316 ( .A1(SI_0_), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n4871) );
  NAND2_X1 U6317 ( .A1(n6596), .A2(n4871), .ZN(n4883) );
  INV_X1 U6318 ( .A(SI_1_), .ZN(n4873) );
  MUX2_X1 U6319 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .S(n4262), .Z(n4895) );
  XNOR2_X1 U6320 ( .A(n4896), .B(n4895), .ZN(n6603) );
  AND2_X2 U6321 ( .A1(n4885), .A2(n6597), .ZN(n4923) );
  NAND2_X1 U6322 ( .A1(n4923), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n4875) );
  INV_X1 U6323 ( .A(n4885), .ZN(n4924) );
  NAND2_X1 U6324 ( .A1(n4924), .A2(n7340), .ZN(n4874) );
  NAND2_X1 U6325 ( .A1(n5506), .A2(n5821), .ZN(n7028) );
  NAND2_X1 U6326 ( .A1(n5295), .A2(n5830), .ZN(n6777) );
  NAND3_X1 U6327 ( .A1(n6777), .A2(n7380), .A3(n9715), .ZN(n4876) );
  XNOR2_X1 U6328 ( .A(n5575), .B(n5433), .ZN(n4887) );
  NAND2_X1 U6329 ( .A1(n5398), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n4880) );
  NAND2_X1 U6330 ( .A1(n4912), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n4879) );
  NAND2_X1 U6331 ( .A1(n4913), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n4878) );
  NAND2_X1 U6332 ( .A1(n4935), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n4877) );
  NAND4_X1 U6333 ( .A1(n4880), .A2(n4879), .A3(n4878), .A4(n4877), .ZN(n6779)
         );
  NAND2_X1 U6334 ( .A1(n6596), .A2(SI_0_), .ZN(n4882) );
  INV_X1 U6335 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n4881) );
  NAND2_X1 U6336 ( .A1(n4882), .A2(n4881), .ZN(n4884) );
  AND2_X1 U6337 ( .A1(n4884), .A2(n4883), .ZN(n8560) );
  MUX2_X1 U6338 ( .A(n9689), .B(n8560), .S(n4885), .Z(n7045) );
  NAND2_X1 U6339 ( .A1(n6770), .A2(n5641), .ZN(n6868) );
  NAND2_X1 U6340 ( .A1(n5504), .A2(n4505), .ZN(n4886) );
  INV_X1 U6341 ( .A(n4887), .ZN(n4888) );
  NAND2_X1 U6342 ( .A1(n4889), .A2(n4888), .ZN(n4890) );
  NAND2_X1 U6343 ( .A1(n5398), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n4894) );
  NAND2_X1 U6344 ( .A1(n4912), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n4893) );
  NAND2_X1 U6345 ( .A1(n4913), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n4892) );
  NAND2_X1 U6346 ( .A1(n4935), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n4891) );
  NOR2_X1 U6347 ( .A1(n5576), .A2(n6866), .ZN(n4905) );
  NAND2_X1 U6348 ( .A1(n4896), .A2(n4895), .ZN(n4899) );
  NAND2_X1 U6349 ( .A1(n4897), .A2(SI_1_), .ZN(n4898) );
  NAND2_X1 U6350 ( .A1(n4899), .A2(n4898), .ZN(n4919) );
  MUX2_X1 U6351 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(P2_DATAO_REG_2__SCAN_IN), 
        .S(n4262), .Z(n4920) );
  INV_X1 U6352 ( .A(SI_2_), .ZN(n4900) );
  XNOR2_X1 U6353 ( .A(n4920), .B(n4900), .ZN(n4918) );
  XNOR2_X1 U6354 ( .A(n4918), .B(n4919), .ZN(n6599) );
  NAND2_X1 U6355 ( .A1(n4923), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n4904) );
  OR2_X1 U6356 ( .A1(n4901), .A2(n8552), .ZN(n4902) );
  XNOR2_X1 U6357 ( .A(n4902), .B(P2_IR_REG_2__SCAN_IN), .ZN(n8008) );
  NAND2_X1 U6358 ( .A1(n4924), .A2(n8008), .ZN(n4903) );
  XNOR2_X1 U6359 ( .A(n7123), .B(n5433), .ZN(n4906) );
  NAND2_X1 U6360 ( .A1(n4905), .A2(n4906), .ZN(n4910) );
  INV_X1 U6361 ( .A(n4905), .ZN(n4908) );
  INV_X1 U6362 ( .A(n4906), .ZN(n4907) );
  NAND2_X1 U6363 ( .A1(n4908), .A2(n4907), .ZN(n4909) );
  AND2_X1 U6364 ( .A1(n4910), .A2(n4909), .ZN(n6897) );
  NAND2_X1 U6365 ( .A1(n6896), .A2(n4910), .ZN(n6929) );
  INV_X1 U6366 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n4911) );
  NAND2_X1 U6367 ( .A1(n5398), .A2(n4911), .ZN(n4917) );
  NAND2_X1 U6368 ( .A1(n4912), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n4916) );
  NAND2_X1 U6369 ( .A1(n4913), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n4915) );
  NAND2_X1 U6370 ( .A1(n4935), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n4914) );
  OR2_X1 U6371 ( .A1(n7116), .A2(n6866), .ZN(n4929) );
  NAND2_X1 U6372 ( .A1(n4919), .A2(n4918), .ZN(n4944) );
  NAND2_X1 U6373 ( .A1(n4920), .A2(SI_2_), .ZN(n4942) );
  NAND2_X1 U6374 ( .A1(n4944), .A2(n4942), .ZN(n4922) );
  INV_X1 U6375 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n6604) );
  INV_X1 U6376 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n4921) );
  XNOR2_X1 U6377 ( .A(n4940), .B(SI_3_), .ZN(n4946) );
  NAND2_X1 U6378 ( .A1(n4923), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n4928) );
  CLKBUF_X3 U6379 ( .A(n4924), .Z(n5296) );
  NAND2_X1 U6380 ( .A1(n4925), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4926) );
  XNOR2_X1 U6381 ( .A(n4926), .B(P2_IR_REG_3__SCAN_IN), .ZN(n7342) );
  NAND2_X1 U6382 ( .A1(n5296), .A2(n7342), .ZN(n4927) );
  OAI211_X2 U6383 ( .C1(n4990), .C2(n6605), .A(n4928), .B(n4927), .ZN(n6962)
         );
  XNOR2_X1 U6384 ( .A(n6962), .B(n5433), .ZN(n4930) );
  XNOR2_X1 U6385 ( .A(n4929), .B(n4930), .ZN(n6928) );
  NAND2_X1 U6386 ( .A1(n6929), .A2(n6928), .ZN(n6927) );
  INV_X1 U6387 ( .A(n4929), .ZN(n4931) );
  NAND2_X1 U6388 ( .A1(n4931), .A2(n4930), .ZN(n4932) );
  NAND2_X1 U6389 ( .A1(n6927), .A2(n4932), .ZN(n6976) );
  NAND2_X1 U6390 ( .A1(n4982), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n4939) );
  INV_X2 U6391 ( .A(n4933), .ZN(n5619) );
  NAND2_X1 U6392 ( .A1(n5619), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n4938) );
  INV_X1 U6393 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n4934) );
  XNOR2_X1 U6394 ( .A(n4934), .B(P2_REG3_REG_3__SCAN_IN), .ZN(n7037) );
  NAND2_X1 U6395 ( .A1(n5398), .A2(n7037), .ZN(n4937) );
  NAND2_X1 U6396 ( .A1(n5554), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n4936) );
  OR2_X1 U6397 ( .A1(n6954), .A2(n6866), .ZN(n4953) );
  INV_X1 U6398 ( .A(n4940), .ZN(n4941) );
  NAND2_X1 U6399 ( .A1(n4941), .A2(SI_3_), .ZN(n4945) );
  AND2_X1 U6400 ( .A1(n4942), .A2(n4945), .ZN(n4943) );
  NAND2_X1 U6401 ( .A1(n4944), .A2(n4943), .ZN(n4947) );
  INV_X1 U6402 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n4948) );
  MUX2_X1 U6403 ( .A(n6600), .B(n4948), .S(n4262), .Z(n4967) );
  XNOR2_X1 U6404 ( .A(n4967), .B(SI_4_), .ZN(n4965) );
  XNOR2_X1 U6405 ( .A(n4966), .B(n4965), .ZN(n6601) );
  NAND2_X1 U6406 ( .A1(n5634), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n4952) );
  NAND2_X1 U6407 ( .A1(n4949), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4950) );
  XNOR2_X1 U6408 ( .A(n4950), .B(P2_IR_REG_4__SCAN_IN), .ZN(n7982) );
  NAND2_X1 U6409 ( .A1(n5296), .A2(n7982), .ZN(n4951) );
  OAI211_X2 U6410 ( .C1(n4990), .C2(n6601), .A(n4952), .B(n4951), .ZN(n9725)
         );
  XNOR2_X1 U6411 ( .A(n5504), .B(n9725), .ZN(n4954) );
  NAND2_X1 U6412 ( .A1(n4953), .A2(n4954), .ZN(n6974) );
  NAND2_X1 U6413 ( .A1(n6976), .A2(n6974), .ZN(n4957) );
  INV_X1 U6414 ( .A(n4953), .ZN(n4956) );
  INV_X1 U6415 ( .A(n4954), .ZN(n4955) );
  NAND2_X1 U6416 ( .A1(n4956), .A2(n4955), .ZN(n6975) );
  NAND2_X1 U6417 ( .A1(n4957), .A2(n6975), .ZN(n6984) );
  NAND2_X1 U6418 ( .A1(n4982), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n4964) );
  NAND2_X1 U6419 ( .A1(n5619), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n4963) );
  NAND3_X1 U6420 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .A3(P2_REG3_REG_5__SCAN_IN), .ZN(n4984) );
  INV_X1 U6421 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n4959) );
  NAND2_X1 U6422 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n4958) );
  NAND2_X1 U6423 ( .A1(n4959), .A2(n4958), .ZN(n4960) );
  AND2_X1 U6424 ( .A1(n4984), .A2(n4960), .ZN(n7050) );
  NAND2_X1 U6425 ( .A1(n5398), .A2(n7050), .ZN(n4962) );
  NAND2_X1 U6426 ( .A1(n5554), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n4961) );
  OR2_X1 U6427 ( .A1(n6978), .A2(n6866), .ZN(n4977) );
  INV_X1 U6428 ( .A(n4967), .ZN(n4968) );
  NAND2_X1 U6429 ( .A1(n4968), .A2(SI_4_), .ZN(n4969) );
  INV_X1 U6430 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n4970) );
  MUX2_X1 U6431 ( .A(n6607), .B(n4970), .S(n6597), .Z(n4993) );
  XNOR2_X1 U6432 ( .A(n4993), .B(SI_5_), .ZN(n4991) );
  XNOR2_X1 U6433 ( .A(n4992), .B(n4991), .ZN(n6606) );
  NAND2_X1 U6434 ( .A1(n5634), .A2(P1_DATAO_REG_5__SCAN_IN), .ZN(n4976) );
  NOR2_X1 U6435 ( .A1(n4971), .A2(n8552), .ZN(n4972) );
  MUX2_X1 U6436 ( .A(n8552), .B(n4972), .S(P2_IR_REG_5__SCAN_IN), .Z(n4974) );
  INV_X1 U6437 ( .A(n4973), .ZN(n5018) );
  NAND2_X1 U6438 ( .A1(n5296), .A2(n7345), .ZN(n4975) );
  XNOR2_X1 U6439 ( .A(n6986), .B(n5433), .ZN(n4978) );
  XNOR2_X1 U6440 ( .A(n4977), .B(n4978), .ZN(n6983) );
  NAND2_X1 U6441 ( .A1(n6984), .A2(n6983), .ZN(n4981) );
  INV_X1 U6442 ( .A(n4977), .ZN(n4979) );
  NAND2_X1 U6443 ( .A1(n4979), .A2(n4978), .ZN(n4980) );
  NAND2_X1 U6444 ( .A1(n4981), .A2(n4980), .ZN(n7153) );
  INV_X1 U6445 ( .A(n7153), .ZN(n5003) );
  NAND2_X1 U6446 ( .A1(n5554), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n4989) );
  NAND2_X1 U6447 ( .A1(n4982), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n4988) );
  INV_X1 U6448 ( .A(n4984), .ZN(n4983) );
  NAND2_X1 U6449 ( .A1(n4983), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5006) );
  INV_X1 U6450 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n7953) );
  NAND2_X1 U6451 ( .A1(n4984), .A2(n7953), .ZN(n4985) );
  AND2_X1 U6452 ( .A1(n5006), .A2(n4985), .ZN(n7434) );
  NAND2_X1 U6453 ( .A1(n5398), .A2(n7434), .ZN(n4987) );
  NAND2_X1 U6454 ( .A1(n5475), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n4986) );
  OR2_X1 U6455 ( .A1(n8084), .A2(n6866), .ZN(n5001) );
  INV_X1 U6456 ( .A(n4993), .ZN(n4994) );
  NAND2_X1 U6457 ( .A1(n4994), .A2(SI_5_), .ZN(n4995) );
  MUX2_X1 U6458 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .S(n6597), .Z(n5015) );
  XNOR2_X1 U6459 ( .A(n5015), .B(SI_6_), .ZN(n5012) );
  XNOR2_X1 U6460 ( .A(n5014), .B(n5012), .ZN(n6608) );
  NAND2_X1 U6461 ( .A1(n5633), .A2(n6608), .ZN(n4999) );
  NAND2_X1 U6462 ( .A1(n5634), .A2(P1_DATAO_REG_6__SCAN_IN), .ZN(n4998) );
  NAND2_X1 U6463 ( .A1(n5018), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4996) );
  XNOR2_X1 U6464 ( .A(n4996), .B(P2_IR_REG_6__SCAN_IN), .ZN(n7347) );
  NAND2_X1 U6465 ( .A1(n5296), .A2(n7347), .ZN(n4997) );
  XNOR2_X1 U6466 ( .A(n7436), .B(n5433), .ZN(n5000) );
  NAND2_X1 U6467 ( .A1(n5001), .A2(n5000), .ZN(n8079) );
  OAI21_X1 U6468 ( .B1(n5001), .B2(n5000), .A(n8079), .ZN(n7154) );
  NAND2_X1 U6469 ( .A1(n4982), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n5011) );
  NAND2_X1 U6470 ( .A1(n5554), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n5010) );
  INV_X1 U6471 ( .A(n5006), .ZN(n5004) );
  NAND2_X1 U6472 ( .A1(n5004), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n5033) );
  INV_X1 U6473 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n5005) );
  NAND2_X1 U6474 ( .A1(n5006), .A2(n5005), .ZN(n5007) );
  AND2_X1 U6475 ( .A1(n5033), .A2(n5007), .ZN(n8088) );
  NAND2_X1 U6476 ( .A1(n5398), .A2(n8088), .ZN(n5009) );
  NAND2_X1 U6477 ( .A1(n5619), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n5008) );
  OR2_X1 U6478 ( .A1(n8139), .A2(n6866), .ZN(n5026) );
  INV_X1 U6479 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n9965) );
  INV_X1 U6480 ( .A(n5012), .ZN(n5013) );
  NAND2_X1 U6481 ( .A1(n5014), .A2(n5013), .ZN(n5017) );
  NAND2_X1 U6482 ( .A1(n5015), .A2(SI_6_), .ZN(n5016) );
  MUX2_X1 U6483 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .S(n6597), .Z(n5042) );
  XNOR2_X1 U6484 ( .A(n5042), .B(SI_7_), .ZN(n5039) );
  XNOR2_X1 U6485 ( .A(n5041), .B(n5039), .ZN(n6611) );
  OR2_X1 U6486 ( .A1(n5018), .A2(P2_IR_REG_6__SCAN_IN), .ZN(n5019) );
  NAND2_X1 U6487 ( .A1(n5019), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5020) );
  XNOR2_X1 U6488 ( .A(n5020), .B(P2_IR_REG_7__SCAN_IN), .ZN(n7349) );
  NAND2_X1 U6489 ( .A1(n5296), .A2(n7349), .ZN(n5021) );
  OAI211_X1 U6490 ( .C1(n5023), .C2(n9965), .A(n5022), .B(n5021), .ZN(n8087)
         );
  XNOR2_X1 U6491 ( .A(n5504), .B(n8087), .ZN(n5027) );
  XNOR2_X1 U6492 ( .A(n5026), .B(n5027), .ZN(n8082) );
  INV_X1 U6493 ( .A(n8082), .ZN(n5024) );
  AND2_X1 U6494 ( .A1(n5024), .A2(n8079), .ZN(n5025) );
  INV_X1 U6495 ( .A(n5026), .ZN(n5029) );
  INV_X1 U6496 ( .A(n5027), .ZN(n5028) );
  NAND2_X1 U6497 ( .A1(n5029), .A2(n5028), .ZN(n8132) );
  NAND2_X1 U6498 ( .A1(n5554), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n5038) );
  NAND2_X1 U6499 ( .A1(n4982), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n5037) );
  INV_X1 U6500 ( .A(n5033), .ZN(n5031) );
  NAND2_X1 U6501 ( .A1(n5031), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n5097) );
  INV_X1 U6502 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n5032) );
  NAND2_X1 U6503 ( .A1(n5033), .A2(n5032), .ZN(n5034) );
  AND2_X1 U6504 ( .A1(n5097), .A2(n5034), .ZN(n8143) );
  NAND2_X1 U6505 ( .A1(n5398), .A2(n8143), .ZN(n5036) );
  NAND2_X1 U6506 ( .A1(n5619), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n5035) );
  OR2_X1 U6507 ( .A1(n9759), .A2(n6866), .ZN(n5075) );
  INV_X1 U6508 ( .A(n5075), .ZN(n5055) );
  INV_X1 U6509 ( .A(n5039), .ZN(n5040) );
  NAND2_X1 U6510 ( .A1(n5041), .A2(n5040), .ZN(n5044) );
  NAND2_X1 U6511 ( .A1(n5042), .A2(SI_7_), .ZN(n5043) );
  INV_X1 U6512 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n6620) );
  INV_X1 U6513 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n5045) );
  MUX2_X1 U6514 ( .A(n6620), .B(n5045), .S(n6597), .Z(n5047) );
  INV_X1 U6515 ( .A(SI_8_), .ZN(n5046) );
  NAND2_X1 U6516 ( .A1(n5047), .A2(n5046), .ZN(n5063) );
  INV_X1 U6517 ( .A(n5047), .ZN(n5048) );
  NAND2_X1 U6518 ( .A1(n5048), .A2(SI_8_), .ZN(n5049) );
  NAND2_X1 U6519 ( .A1(n5063), .A2(n5049), .ZN(n5061) );
  INV_X1 U6520 ( .A(n5061), .ZN(n5050) );
  NAND2_X1 U6521 ( .A1(n5634), .A2(P1_DATAO_REG_8__SCAN_IN), .ZN(n5054) );
  OR2_X1 U6522 ( .A1(n5051), .A2(n8552), .ZN(n5052) );
  XNOR2_X1 U6523 ( .A(n5052), .B(P2_IR_REG_8__SCAN_IN), .ZN(n7351) );
  NAND2_X1 U6524 ( .A1(n5296), .A2(n7351), .ZN(n5053) );
  NAND2_X1 U6525 ( .A1(n5055), .A2(n5074), .ZN(n5073) );
  AND2_X1 U6526 ( .A1(n8132), .A2(n5073), .ZN(n7226) );
  NAND2_X1 U6527 ( .A1(n4982), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n5059) );
  NAND2_X1 U6528 ( .A1(n5619), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n5058) );
  XNOR2_X1 U6529 ( .A(n5097), .B(P2_REG3_REG_9__SCAN_IN), .ZN(n9994) );
  NAND2_X1 U6530 ( .A1(n5398), .A2(n9994), .ZN(n5057) );
  NAND2_X1 U6531 ( .A1(n5554), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n5056) );
  OR2_X1 U6532 ( .A1(n8138), .A2(n6866), .ZN(n5071) );
  NAND2_X1 U6533 ( .A1(n5060), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5088) );
  XNOR2_X1 U6534 ( .A(n5088), .B(P2_IR_REG_9__SCAN_IN), .ZN(n7353) );
  INV_X1 U6535 ( .A(n7353), .ZN(n7930) );
  INV_X1 U6536 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n5064) );
  MUX2_X1 U6537 ( .A(n6625), .B(n5064), .S(n6597), .Z(n5065) );
  NAND2_X1 U6538 ( .A1(n5065), .A2(n9908), .ZN(n5080) );
  INV_X1 U6539 ( .A(n5065), .ZN(n5066) );
  NAND2_X1 U6540 ( .A1(n5066), .A2(SI_9_), .ZN(n5067) );
  XNOR2_X1 U6541 ( .A(n5079), .B(n4820), .ZN(n6622) );
  NAND2_X1 U6542 ( .A1(n6622), .A2(n5633), .ZN(n5069) );
  NAND2_X1 U6543 ( .A1(n5634), .A2(P1_DATAO_REG_9__SCAN_IN), .ZN(n5068) );
  OAI211_X1 U6544 ( .C1(n4885), .C2(n7930), .A(n5069), .B(n5068), .ZN(n9995)
         );
  XNOR2_X1 U6545 ( .A(n9995), .B(n5504), .ZN(n5070) );
  NAND2_X1 U6546 ( .A1(n5071), .A2(n5070), .ZN(n5077) );
  OAI21_X1 U6547 ( .B1(n5071), .B2(n5070), .A(n5077), .ZN(n7232) );
  AND2_X1 U6548 ( .A1(n7226), .A2(n4396), .ZN(n5072) );
  INV_X1 U6549 ( .A(n5073), .ZN(n5076) );
  XNOR2_X1 U6550 ( .A(n5075), .B(n5074), .ZN(n8135) );
  NAND2_X1 U6551 ( .A1(n5081), .A2(n5080), .ZN(n5107) );
  INV_X1 U6552 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n5082) );
  MUX2_X1 U6553 ( .A(n6635), .B(n5082), .S(n6597), .Z(n5084) );
  INV_X1 U6554 ( .A(SI_10_), .ZN(n5083) );
  NAND2_X1 U6555 ( .A1(n5084), .A2(n5083), .ZN(n5108) );
  INV_X1 U6556 ( .A(n5084), .ZN(n5085) );
  NAND2_X1 U6557 ( .A1(n5085), .A2(SI_10_), .ZN(n5086) );
  XNOR2_X1 U6558 ( .A(n5107), .B(n4816), .ZN(n6626) );
  NAND2_X1 U6559 ( .A1(n6626), .A2(n5633), .ZN(n5094) );
  INV_X1 U6560 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n5087) );
  NAND2_X1 U6561 ( .A1(n5088), .A2(n5087), .ZN(n5089) );
  NAND2_X1 U6562 ( .A1(n5089), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5091) );
  NAND2_X1 U6563 ( .A1(n5091), .A2(n5090), .ZN(n5110) );
  OR2_X1 U6564 ( .A1(n5091), .A2(n5090), .ZN(n5092) );
  AOI22_X1 U6565 ( .A1(n5634), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n5296), .B2(
        n7355), .ZN(n5093) );
  NAND2_X1 U6566 ( .A1(n5094), .A2(n5093), .ZN(n8115) );
  XNOR2_X1 U6567 ( .A(n8115), .B(n5504), .ZN(n5106) );
  NAND2_X1 U6568 ( .A1(n4982), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n5104) );
  NAND2_X1 U6569 ( .A1(n5619), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n5103) );
  INV_X1 U6570 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n5096) );
  INV_X1 U6571 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n5095) );
  OAI21_X1 U6572 ( .B1(n5097), .B2(n5096), .A(n5095), .ZN(n5100) );
  INV_X1 U6573 ( .A(n5097), .ZN(n5099) );
  NAND2_X1 U6574 ( .A1(n5099), .A2(n5098), .ZN(n5114) );
  AND2_X1 U6575 ( .A1(n5100), .A2(n5114), .ZN(n8116) );
  NAND2_X1 U6576 ( .A1(n5398), .A2(n8116), .ZN(n5102) );
  NAND2_X1 U6577 ( .A1(n5554), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n5101) );
  OR2_X1 U6578 ( .A1(n9757), .A2(n6866), .ZN(n5105) );
  XNOR2_X1 U6579 ( .A(n5106), .B(n5105), .ZN(n8109) );
  NAND2_X1 U6580 ( .A1(n5107), .A2(n4816), .ZN(n5109) );
  NAND2_X1 U6581 ( .A1(n5109), .A2(n5108), .ZN(n5125) );
  MUX2_X1 U6582 ( .A(n6640), .B(n6638), .S(n6597), .Z(n5128) );
  XNOR2_X1 U6583 ( .A(n5128), .B(SI_11_), .ZN(n5126) );
  NAND2_X1 U6584 ( .A1(n6637), .A2(n5633), .ZN(n5113) );
  NAND2_X1 U6585 ( .A1(n5110), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5111) );
  XNOR2_X1 U6586 ( .A(n5111), .B(P2_IR_REG_11__SCAN_IN), .ZN(n7357) );
  AOI22_X1 U6587 ( .A1(n5634), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n5296), .B2(
        n7357), .ZN(n5112) );
  XNOR2_X1 U6588 ( .A(n8208), .B(n5504), .ZN(n5120) );
  NAND2_X1 U6589 ( .A1(n4982), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n5119) );
  NAND2_X1 U6590 ( .A1(n5554), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n5118) );
  NAND2_X1 U6591 ( .A1(n5114), .A2(n8203), .ZN(n5115) );
  AND2_X1 U6592 ( .A1(n5139), .A2(n5115), .ZN(n8209) );
  NAND2_X1 U6593 ( .A1(n5398), .A2(n8209), .ZN(n5117) );
  NAND2_X1 U6594 ( .A1(n5619), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n5116) );
  NOR2_X1 U6595 ( .A1(n8112), .A2(n6866), .ZN(n5121) );
  XNOR2_X1 U6596 ( .A(n5120), .B(n5121), .ZN(n8201) );
  INV_X1 U6597 ( .A(n5120), .ZN(n5122) );
  NAND2_X1 U6598 ( .A1(n5122), .A2(n5121), .ZN(n5123) );
  INV_X1 U6599 ( .A(n5125), .ZN(n5127) );
  INV_X1 U6600 ( .A(n5128), .ZN(n5129) );
  NAND2_X1 U6601 ( .A1(n5129), .A2(SI_11_), .ZN(n5130) );
  MUX2_X1 U6602 ( .A(n6684), .B(n6686), .S(n6597), .Z(n5132) );
  INV_X1 U6603 ( .A(SI_12_), .ZN(n5131) );
  NAND2_X1 U6604 ( .A1(n5132), .A2(n5131), .ZN(n5151) );
  INV_X1 U6605 ( .A(n5132), .ZN(n5133) );
  NAND2_X1 U6606 ( .A1(n5133), .A2(SI_12_), .ZN(n5134) );
  NAND2_X1 U6607 ( .A1(n5151), .A2(n5134), .ZN(n5152) );
  XNOR2_X1 U6608 ( .A(n5153), .B(n5152), .ZN(n6683) );
  NAND2_X1 U6609 ( .A1(n6683), .A2(n5633), .ZN(n5137) );
  NAND2_X1 U6610 ( .A1(n4352), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5135) );
  XNOR2_X1 U6611 ( .A(n5135), .B(P2_IR_REG_12__SCAN_IN), .ZN(n7450) );
  AOI22_X1 U6612 ( .A1(n5634), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n5296), .B2(
        n7450), .ZN(n5136) );
  XNOR2_X1 U6613 ( .A(n9786), .B(n5504), .ZN(n5145) );
  NAND2_X1 U6614 ( .A1(n4982), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n5144) );
  NAND2_X1 U6615 ( .A1(n5554), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n5143) );
  NAND2_X1 U6616 ( .A1(n5139), .A2(n5138), .ZN(n5140) );
  AND2_X1 U6617 ( .A1(n5163), .A2(n5140), .ZN(n9695) );
  NAND2_X1 U6618 ( .A1(n5398), .A2(n9695), .ZN(n5142) );
  NAND2_X1 U6619 ( .A1(n5619), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n5141) );
  OR2_X1 U6620 ( .A1(n8204), .A2(n6866), .ZN(n5146) );
  NAND2_X1 U6621 ( .A1(n5145), .A2(n5146), .ZN(n5150) );
  INV_X1 U6622 ( .A(n5145), .ZN(n5148) );
  INV_X1 U6623 ( .A(n5146), .ZN(n5147) );
  NAND2_X1 U6624 ( .A1(n5148), .A2(n5147), .ZN(n5149) );
  NAND2_X1 U6625 ( .A1(n5150), .A2(n5149), .ZN(n7612) );
  MUX2_X1 U6626 ( .A(n6731), .B(n6733), .S(n6597), .Z(n5155) );
  NAND2_X1 U6627 ( .A1(n5155), .A2(n5154), .ZN(n5175) );
  INV_X1 U6628 ( .A(n5155), .ZN(n5156) );
  NAND2_X1 U6629 ( .A1(n5156), .A2(SI_13_), .ZN(n5157) );
  NAND2_X1 U6630 ( .A1(n6730), .A2(n5633), .ZN(n5160) );
  OR2_X1 U6631 ( .A1(n5158), .A2(n8552), .ZN(n5177) );
  XNOR2_X1 U6632 ( .A(n5177), .B(P2_IR_REG_13__SCAN_IN), .ZN(n7475) );
  AOI22_X1 U6633 ( .A1(n5634), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n5296), .B2(
        n7475), .ZN(n5159) );
  NAND2_X2 U6634 ( .A1(n5160), .A2(n5159), .ZN(n7587) );
  XNOR2_X1 U6635 ( .A(n7587), .B(n5433), .ZN(n5169) );
  NAND2_X1 U6636 ( .A1(n5554), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n5168) );
  NAND2_X1 U6637 ( .A1(n4982), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n5167) );
  INV_X1 U6638 ( .A(n5163), .ZN(n5161) );
  NAND2_X1 U6639 ( .A1(n5161), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n5186) );
  INV_X1 U6640 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n5162) );
  NAND2_X1 U6641 ( .A1(n5163), .A2(n5162), .ZN(n5164) );
  AND2_X1 U6642 ( .A1(n5186), .A2(n5164), .ZN(n7625) );
  NAND2_X1 U6643 ( .A1(n5398), .A2(n7625), .ZN(n5166) );
  NAND2_X1 U6644 ( .A1(n5619), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n5165) );
  NOR2_X1 U6645 ( .A1(n7746), .A2(n6866), .ZN(n5170) );
  XNOR2_X1 U6646 ( .A(n5169), .B(n5170), .ZN(n7619) );
  INV_X1 U6647 ( .A(n5169), .ZN(n5172) );
  INV_X1 U6648 ( .A(n5170), .ZN(n5171) );
  MUX2_X1 U6649 ( .A(n9887), .B(n6745), .S(n6597), .Z(n5199) );
  XNOR2_X1 U6650 ( .A(n5199), .B(SI_14_), .ZN(n5198) );
  XNOR2_X1 U6651 ( .A(n5201), .B(n5198), .ZN(n6743) );
  NAND2_X1 U6652 ( .A1(n6743), .A2(n5633), .ZN(n5183) );
  NAND2_X1 U6653 ( .A1(n5177), .A2(n5176), .ZN(n5178) );
  NAND2_X1 U6654 ( .A1(n5178), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5180) );
  OR2_X1 U6655 ( .A1(n5180), .A2(n5179), .ZN(n5181) );
  NAND2_X1 U6656 ( .A1(n5180), .A2(n5179), .ZN(n5226) );
  AOI22_X1 U6657 ( .A1(n5634), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n5296), .B2(
        n7768), .ZN(n5182) );
  NAND2_X1 U6658 ( .A1(n5183), .A2(n5182), .ZN(n7657) );
  XNOR2_X1 U6659 ( .A(n7657), .B(n5504), .ZN(n5192) );
  INV_X1 U6660 ( .A(n5186), .ZN(n5184) );
  NAND2_X1 U6661 ( .A1(n5184), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n5231) );
  INV_X1 U6662 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n5185) );
  NAND2_X1 U6663 ( .A1(n5186), .A2(n5185), .ZN(n5187) );
  AND2_X1 U6664 ( .A1(n5231), .A2(n5187), .ZN(n7749) );
  NAND2_X1 U6665 ( .A1(n5398), .A2(n7749), .ZN(n5191) );
  NAND2_X1 U6666 ( .A1(n4982), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n5190) );
  NAND2_X1 U6667 ( .A1(n5619), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n5189) );
  NAND2_X1 U6668 ( .A1(n5554), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n5188) );
  OR2_X1 U6669 ( .A1(n7818), .A2(n6866), .ZN(n5193) );
  NAND2_X1 U6670 ( .A1(n5192), .A2(n5193), .ZN(n5197) );
  INV_X1 U6671 ( .A(n5192), .ZN(n5195) );
  INV_X1 U6672 ( .A(n5193), .ZN(n5194) );
  NAND2_X1 U6673 ( .A1(n5195), .A2(n5194), .ZN(n5196) );
  NAND2_X1 U6674 ( .A1(n5197), .A2(n5196), .ZN(n7743) );
  INV_X1 U6675 ( .A(n5199), .ZN(n5200) );
  MUX2_X1 U6676 ( .A(n9884), .B(n6925), .S(n6597), .Z(n5202) );
  NAND2_X1 U6677 ( .A1(n5202), .A2(n9921), .ZN(n5205) );
  INV_X1 U6678 ( .A(n5202), .ZN(n5203) );
  NAND2_X1 U6679 ( .A1(n5203), .A2(SI_15_), .ZN(n5204) );
  NAND2_X1 U6680 ( .A1(n5205), .A2(n5204), .ZN(n5224) );
  OAI21_X2 U6681 ( .B1(n5225), .B2(n5224), .A(n5205), .ZN(n5248) );
  MUX2_X1 U6682 ( .A(n5206), .B(n6949), .S(n6597), .Z(n5208) );
  NAND2_X1 U6683 ( .A1(n5208), .A2(n5207), .ZN(n5249) );
  INV_X1 U6684 ( .A(n5208), .ZN(n5209) );
  NAND2_X1 U6685 ( .A1(n5209), .A2(SI_16_), .ZN(n5210) );
  XNOR2_X1 U6686 ( .A(n5248), .B(n5247), .ZN(n6894) );
  NAND2_X1 U6687 ( .A1(n6894), .A2(n5633), .ZN(n5216) );
  NOR2_X1 U6688 ( .A1(n5211), .A2(n8552), .ZN(n5212) );
  MUX2_X1 U6689 ( .A(n8552), .B(n5212), .S(P2_IR_REG_16__SCAN_IN), .Z(n5213)
         );
  INV_X1 U6690 ( .A(n5213), .ZN(n5214) );
  AND2_X1 U6691 ( .A1(n5214), .A2(n5251), .ZN(n8258) );
  AOI22_X1 U6692 ( .A1(n5634), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n5296), .B2(
        n8258), .ZN(n5215) );
  XNOR2_X1 U6693 ( .A(n8530), .B(n5433), .ZN(n5240) );
  NAND2_X1 U6694 ( .A1(n4982), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n5223) );
  NAND2_X1 U6695 ( .A1(n5619), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n5222) );
  INV_X1 U6696 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n5230) );
  NAND2_X1 U6697 ( .A1(n5217), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n5255) );
  INV_X1 U6698 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n5218) );
  NAND2_X1 U6699 ( .A1(n5233), .A2(n5218), .ZN(n5219) );
  AND2_X1 U6700 ( .A1(n5255), .A2(n5219), .ZN(n7842) );
  NAND2_X1 U6701 ( .A1(n5398), .A2(n7842), .ZN(n5221) );
  NAND2_X1 U6702 ( .A1(n5554), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n5220) );
  NAND4_X1 U6703 ( .A1(n5223), .A2(n5222), .A3(n5221), .A4(n5220), .ZN(n8233)
         );
  AND2_X1 U6704 ( .A1(n8233), .A2(n5641), .ZN(n5241) );
  NAND2_X1 U6705 ( .A1(n5240), .A2(n5241), .ZN(n7836) );
  NAND2_X1 U6706 ( .A1(n6923), .A2(n5633), .ZN(n5229) );
  NAND2_X1 U6707 ( .A1(n5226), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5227) );
  XNOR2_X1 U6708 ( .A(n5227), .B(P2_IR_REG_15__SCAN_IN), .ZN(n7864) );
  AOI22_X1 U6709 ( .A1(n5634), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n5296), .B2(
        n7864), .ZN(n5228) );
  XNOR2_X1 U6710 ( .A(n7820), .B(n5504), .ZN(n7810) );
  INV_X1 U6711 ( .A(n7810), .ZN(n5238) );
  NAND2_X1 U6712 ( .A1(n5554), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n5237) );
  NAND2_X1 U6713 ( .A1(n4982), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n5236) );
  NAND2_X1 U6714 ( .A1(n5231), .A2(n5230), .ZN(n5232) );
  AND2_X1 U6715 ( .A1(n5233), .A2(n5232), .ZN(n7815) );
  NAND2_X1 U6716 ( .A1(n5398), .A2(n7815), .ZN(n5235) );
  NAND2_X1 U6717 ( .A1(n5619), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n5234) );
  OR2_X1 U6718 ( .A1(n7840), .A2(n6866), .ZN(n7813) );
  INV_X1 U6719 ( .A(n7813), .ZN(n7833) );
  NAND2_X1 U6720 ( .A1(n5238), .A2(n7833), .ZN(n5239) );
  AND2_X1 U6721 ( .A1(n7836), .A2(n5239), .ZN(n5246) );
  NAND3_X1 U6722 ( .A1(n7836), .A2(n7810), .A3(n7813), .ZN(n5244) );
  INV_X1 U6723 ( .A(n5240), .ZN(n5243) );
  INV_X1 U6724 ( .A(n5241), .ZN(n5242) );
  NAND2_X1 U6725 ( .A1(n5243), .A2(n5242), .ZN(n7835) );
  NAND2_X1 U6726 ( .A1(n5244), .A2(n7835), .ZN(n5245) );
  INV_X1 U6727 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n5250) );
  MUX2_X1 U6728 ( .A(n6972), .B(n5250), .S(n6597), .Z(n5268) );
  XNOR2_X1 U6729 ( .A(n5268), .B(SI_17_), .ZN(n5266) );
  XNOR2_X1 U6730 ( .A(n5267), .B(n5266), .ZN(n6970) );
  NAND2_X1 U6731 ( .A1(n6970), .A2(n5633), .ZN(n5254) );
  NAND2_X1 U6732 ( .A1(n5251), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5252) );
  XNOR2_X1 U6733 ( .A(n5252), .B(P2_IR_REG_17__SCAN_IN), .ZN(n7875) );
  AOI22_X1 U6734 ( .A1(n5634), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n5296), .B2(
        n7875), .ZN(n5253) );
  XNOR2_X1 U6735 ( .A(n8526), .B(n5504), .ZN(n5261) );
  NAND2_X1 U6736 ( .A1(n4982), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n5260) );
  NAND2_X1 U6737 ( .A1(n5554), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n5259) );
  NAND2_X1 U6738 ( .A1(n5255), .A2(n7885), .ZN(n5256) );
  AND2_X1 U6739 ( .A1(n5302), .A2(n5256), .ZN(n7798) );
  NAND2_X1 U6740 ( .A1(n5398), .A2(n7798), .ZN(n5258) );
  NAND2_X1 U6741 ( .A1(n5475), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n5257) );
  NOR2_X1 U6742 ( .A1(n7828), .A2(n6866), .ZN(n5262) );
  XNOR2_X1 U6743 ( .A(n5261), .B(n5262), .ZN(n7796) );
  NAND2_X1 U6744 ( .A1(n7797), .A2(n7796), .ZN(n5265) );
  INV_X1 U6745 ( .A(n5261), .ZN(n5263) );
  NAND2_X1 U6746 ( .A1(n5263), .A2(n5262), .ZN(n5264) );
  NAND2_X1 U6747 ( .A1(n5265), .A2(n5264), .ZN(n7824) );
  INV_X1 U6748 ( .A(n5268), .ZN(n5269) );
  NAND2_X1 U6749 ( .A1(n5269), .A2(SI_17_), .ZN(n5283) );
  NAND2_X1 U6750 ( .A1(n5289), .A2(n5283), .ZN(n5270) );
  MUX2_X1 U6751 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .S(n6597), .Z(n5282) );
  XNOR2_X1 U6752 ( .A(n5282), .B(SI_18_), .ZN(n5285) );
  XNOR2_X1 U6753 ( .A(n5270), .B(n5285), .ZN(n7084) );
  NAND2_X1 U6754 ( .A1(n7084), .A2(n5633), .ZN(n5273) );
  XNOR2_X1 U6755 ( .A(n5271), .B(P2_IR_REG_18__SCAN_IN), .ZN(n8022) );
  AOI22_X1 U6756 ( .A1(n5634), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n5296), .B2(
        n8022), .ZN(n5272) );
  XNOR2_X1 U6757 ( .A(n8519), .B(n5433), .ZN(n5280) );
  NAND2_X1 U6758 ( .A1(n4982), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n5277) );
  NAND2_X1 U6759 ( .A1(n5619), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n5276) );
  XNOR2_X1 U6760 ( .A(n5302), .B(P2_REG3_REG_18__SCAN_IN), .ZN(n8439) );
  NAND2_X1 U6761 ( .A1(n5398), .A2(n8439), .ZN(n5275) );
  NAND2_X1 U6762 ( .A1(n5554), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n5274) );
  NAND4_X1 U6763 ( .A1(n5277), .A2(n5276), .A3(n5275), .A4(n5274), .ZN(n8425)
         );
  NAND2_X1 U6764 ( .A1(n8425), .A2(n5641), .ZN(n5278) );
  XNOR2_X1 U6765 ( .A(n5280), .B(n5278), .ZN(n7823) );
  INV_X1 U6766 ( .A(n5278), .ZN(n5279) );
  NAND2_X1 U6767 ( .A1(n5280), .A2(n5279), .ZN(n5281) );
  NAND2_X1 U6768 ( .A1(n5282), .A2(SI_18_), .ZN(n5284) );
  AND2_X1 U6769 ( .A1(n5283), .A2(n5284), .ZN(n5288) );
  INV_X1 U6770 ( .A(n5284), .ZN(n5287) );
  INV_X1 U6771 ( .A(n5285), .ZN(n5286) );
  MUX2_X1 U6772 ( .A(n8050), .B(n5290), .S(n4262), .Z(n5292) );
  INV_X1 U6773 ( .A(SI_19_), .ZN(n5291) );
  NAND2_X1 U6774 ( .A1(n5292), .A2(n5291), .ZN(n5314) );
  INV_X1 U6775 ( .A(n5292), .ZN(n5293) );
  NAND2_X1 U6776 ( .A1(n5293), .A2(SI_19_), .ZN(n5294) );
  NAND2_X1 U6777 ( .A1(n5314), .A2(n5294), .ZN(n5315) );
  XNOR2_X1 U6778 ( .A(n5316), .B(n5315), .ZN(n7088) );
  NAND2_X1 U6779 ( .A1(n7088), .A2(n5633), .ZN(n5298) );
  AOI22_X1 U6780 ( .A1(n5634), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n5296), .B2(
        n5295), .ZN(n5297) );
  XNOR2_X1 U6781 ( .A(n8515), .B(n5504), .ZN(n5308) );
  NAND2_X1 U6782 ( .A1(n5554), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n5307) );
  NAND2_X1 U6783 ( .A1(n4982), .A2(P2_REG2_REG_19__SCAN_IN), .ZN(n5306) );
  INV_X1 U6784 ( .A(n5302), .ZN(n5300) );
  AND2_X1 U6785 ( .A1(P2_REG3_REG_19__SCAN_IN), .A2(P2_REG3_REG_18__SCAN_IN), 
        .ZN(n5299) );
  NAND2_X1 U6786 ( .A1(n5300), .A2(n5299), .ZN(n5324) );
  INV_X1 U6787 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n7825) );
  INV_X1 U6788 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n5301) );
  OAI21_X1 U6789 ( .B1(n5302), .B2(n7825), .A(n5301), .ZN(n5303) );
  AND2_X1 U6790 ( .A1(n5324), .A2(n5303), .ZN(n8430) );
  NAND2_X1 U6791 ( .A1(n5398), .A2(n8430), .ZN(n5305) );
  NAND2_X1 U6792 ( .A1(n5619), .A2(P2_REG1_REG_19__SCAN_IN), .ZN(n5304) );
  NAND4_X1 U6793 ( .A1(n5307), .A2(n5306), .A3(n5305), .A4(n5304), .ZN(n8446)
         );
  NAND2_X1 U6794 ( .A1(n8446), .A2(n5641), .ZN(n5309) );
  NAND2_X1 U6795 ( .A1(n5308), .A2(n5309), .ZN(n5313) );
  INV_X1 U6796 ( .A(n5308), .ZN(n5311) );
  INV_X1 U6797 ( .A(n5309), .ZN(n5310) );
  NAND2_X1 U6798 ( .A1(n5311), .A2(n5310), .ZN(n5312) );
  NAND2_X1 U6799 ( .A1(n5313), .A2(n5312), .ZN(n8123) );
  INV_X1 U6800 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n5317) );
  MUX2_X1 U6801 ( .A(n7378), .B(n5317), .S(n6597), .Z(n5319) );
  INV_X1 U6802 ( .A(SI_20_), .ZN(n5318) );
  NAND2_X1 U6803 ( .A1(n5319), .A2(n5318), .ZN(n5332) );
  INV_X1 U6804 ( .A(n5319), .ZN(n5320) );
  NAND2_X1 U6805 ( .A1(n5320), .A2(SI_20_), .ZN(n5321) );
  XNOR2_X1 U6806 ( .A(n5331), .B(n5330), .ZN(n7195) );
  NAND2_X1 U6807 ( .A1(n7195), .A2(n5633), .ZN(n5323) );
  NAND2_X1 U6808 ( .A1(n5634), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n5322) );
  XNOR2_X1 U6809 ( .A(n8509), .B(n5433), .ZN(n5345) );
  NAND2_X1 U6810 ( .A1(n5554), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n5329) );
  NAND2_X1 U6811 ( .A1(n4982), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n5328) );
  NAND2_X1 U6812 ( .A1(n5324), .A2(n9926), .ZN(n5325) );
  AND2_X1 U6813 ( .A1(n5367), .A2(n5325), .ZN(n8413) );
  NAND2_X1 U6814 ( .A1(n5398), .A2(n8413), .ZN(n5327) );
  NAND2_X1 U6815 ( .A1(n5475), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n5326) );
  NOR2_X1 U6816 ( .A1(n8154), .A2(n6866), .ZN(n5344) );
  XNOR2_X1 U6817 ( .A(n5345), .B(n5344), .ZN(n8182) );
  INV_X1 U6818 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n5333) );
  MUX2_X1 U6819 ( .A(n9870), .B(n5333), .S(n6597), .Z(n5352) );
  XNOR2_X1 U6820 ( .A(n5352), .B(SI_21_), .ZN(n5351) );
  XNOR2_X1 U6821 ( .A(n5350), .B(n5351), .ZN(n7275) );
  NAND2_X1 U6822 ( .A1(n7275), .A2(n5633), .ZN(n5335) );
  NAND2_X1 U6823 ( .A1(n5634), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n5334) );
  XNOR2_X1 U6824 ( .A(n8502), .B(n5433), .ZN(n5342) );
  NAND2_X1 U6825 ( .A1(n4982), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n5339) );
  NAND2_X1 U6826 ( .A1(n5619), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n5338) );
  XNOR2_X1 U6827 ( .A(n5367), .B(P2_REG3_REG_21__SCAN_IN), .ZN(n8394) );
  NAND2_X1 U6828 ( .A1(n5398), .A2(n8394), .ZN(n5337) );
  NAND2_X1 U6829 ( .A1(n5554), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n5336) );
  NAND4_X1 U6830 ( .A1(n5339), .A2(n5338), .A3(n5337), .A4(n5336), .ZN(n8410)
         );
  NAND2_X1 U6831 ( .A1(n8410), .A2(n5641), .ZN(n5341) );
  INV_X1 U6832 ( .A(n5341), .ZN(n5340) );
  NAND2_X1 U6833 ( .A1(n5342), .A2(n5340), .ZN(n5346) );
  INV_X1 U6834 ( .A(n5346), .ZN(n5343) );
  XNOR2_X1 U6835 ( .A(n5342), .B(n5341), .ZN(n8150) );
  NOR2_X1 U6836 ( .A1(n5343), .A2(n8150), .ZN(n5348) );
  OR2_X1 U6837 ( .A1(n8182), .A2(n5348), .ZN(n5349) );
  NAND2_X1 U6838 ( .A1(n5345), .A2(n5344), .ZN(n8148) );
  AND2_X1 U6839 ( .A1(n8148), .A2(n5346), .ZN(n5347) );
  INV_X1 U6840 ( .A(n5352), .ZN(n5353) );
  NAND2_X1 U6841 ( .A1(n5353), .A2(SI_21_), .ZN(n5354) );
  INV_X1 U6842 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n5356) );
  MUX2_X1 U6843 ( .A(n7421), .B(n5356), .S(n6597), .Z(n5358) );
  INV_X1 U6844 ( .A(SI_22_), .ZN(n5357) );
  NAND2_X1 U6845 ( .A1(n5358), .A2(n5357), .ZN(n5377) );
  INV_X1 U6846 ( .A(n5358), .ZN(n5359) );
  NAND2_X1 U6847 ( .A1(n5359), .A2(SI_22_), .ZN(n5360) );
  NAND2_X1 U6848 ( .A1(n5377), .A2(n5360), .ZN(n5378) );
  XNOR2_X1 U6849 ( .A(n5379), .B(n5378), .ZN(n7381) );
  NAND2_X1 U6850 ( .A1(n7381), .A2(n5633), .ZN(n5362) );
  NAND2_X1 U6851 ( .A1(n5634), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n5361) );
  XNOR2_X1 U6852 ( .A(n8497), .B(n5504), .ZN(n5373) );
  XNOR2_X1 U6853 ( .A(n5375), .B(n5373), .ZN(n8193) );
  NAND2_X1 U6854 ( .A1(n4912), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n5372) );
  NAND2_X1 U6855 ( .A1(n5554), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n5371) );
  INV_X1 U6856 ( .A(n5367), .ZN(n5364) );
  AND2_X1 U6857 ( .A1(P2_REG3_REG_21__SCAN_IN), .A2(P2_REG3_REG_22__SCAN_IN), 
        .ZN(n5363) );
  NAND2_X1 U6858 ( .A1(n5364), .A2(n5363), .ZN(n5403) );
  INV_X1 U6859 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n5366) );
  INV_X1 U6860 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n5365) );
  OAI21_X1 U6861 ( .B1(n5367), .B2(n5366), .A(n5365), .ZN(n5368) );
  AND2_X1 U6862 ( .A1(n5403), .A2(n5368), .ZN(n8375) );
  NAND2_X1 U6863 ( .A1(n5398), .A2(n8375), .ZN(n5370) );
  NAND2_X1 U6864 ( .A1(n5475), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n5369) );
  OR2_X1 U6865 ( .A1(n8361), .A2(n6866), .ZN(n8192) );
  NAND2_X1 U6866 ( .A1(n8193), .A2(n8192), .ZN(n8191) );
  INV_X1 U6867 ( .A(n5373), .ZN(n5374) );
  OR2_X1 U6868 ( .A1(n5375), .A2(n5374), .ZN(n5376) );
  INV_X1 U6869 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n5381) );
  INV_X1 U6870 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n5380) );
  MUX2_X1 U6871 ( .A(n5381), .B(n5380), .S(n6597), .Z(n5383) );
  INV_X1 U6872 ( .A(SI_23_), .ZN(n5382) );
  NAND2_X1 U6873 ( .A1(n5383), .A2(n5382), .ZN(n5390) );
  INV_X1 U6874 ( .A(n5383), .ZN(n5384) );
  NAND2_X1 U6875 ( .A1(n5384), .A2(SI_23_), .ZN(n5385) );
  XNOR2_X1 U6876 ( .A(n5389), .B(n5388), .ZN(n7571) );
  NAND2_X1 U6877 ( .A1(n7571), .A2(n5633), .ZN(n5387) );
  NAND2_X1 U6878 ( .A1(n5634), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n5386) );
  XNOR2_X1 U6879 ( .A(n8367), .B(n5433), .ZN(n5413) );
  NAND2_X1 U6880 ( .A1(n5389), .A2(n5388), .ZN(n5391) );
  INV_X1 U6881 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n7654) );
  INV_X1 U6882 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n5392) );
  MUX2_X1 U6883 ( .A(n7654), .B(n5392), .S(n6597), .Z(n5421) );
  XNOR2_X1 U6884 ( .A(n5421), .B(SI_24_), .ZN(n5420) );
  NAND2_X1 U6885 ( .A1(n7641), .A2(n5633), .ZN(n5394) );
  NAND2_X1 U6886 ( .A1(n5634), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n5393) );
  XNOR2_X1 U6887 ( .A(n8486), .B(n5433), .ZN(n8172) );
  INV_X1 U6888 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n8102) );
  INV_X1 U6889 ( .A(n5405), .ZN(n5395) );
  NAND2_X1 U6890 ( .A1(n5395), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n5437) );
  INV_X1 U6891 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n5396) );
  NAND2_X1 U6892 ( .A1(n5405), .A2(n5396), .ZN(n5397) );
  AND2_X1 U6893 ( .A1(n5437), .A2(n5397), .ZN(n8347) );
  NAND2_X1 U6894 ( .A1(n8347), .A2(n5398), .ZN(n5402) );
  NAND2_X1 U6895 ( .A1(n4912), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n5401) );
  NAND2_X1 U6896 ( .A1(n5554), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n5400) );
  NAND2_X1 U6897 ( .A1(n5619), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n5399) );
  INV_X1 U6898 ( .A(n8362), .ZN(n8231) );
  NAND2_X1 U6899 ( .A1(n4982), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n5410) );
  NAND2_X1 U6900 ( .A1(n5554), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n5409) );
  NAND2_X1 U6901 ( .A1(n5403), .A2(n8102), .ZN(n5404) );
  AND2_X1 U6902 ( .A1(n5405), .A2(n5404), .ZN(n8368) );
  NAND2_X1 U6903 ( .A1(n5398), .A2(n8368), .ZN(n5408) );
  NAND2_X1 U6904 ( .A1(n5619), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n5407) );
  NOR2_X1 U6905 ( .A1(n8383), .A2(n6866), .ZN(n8170) );
  OAI21_X1 U6906 ( .B1(n8172), .B2(n8231), .A(n8170), .ZN(n5411) );
  INV_X1 U6907 ( .A(n5411), .ZN(n5412) );
  NAND2_X1 U6908 ( .A1(n8169), .A2(n5412), .ZN(n5419) );
  NOR2_X1 U6909 ( .A1(n8362), .A2(n6866), .ZN(n8171) );
  INV_X1 U6910 ( .A(n5413), .ZN(n5414) );
  INV_X1 U6911 ( .A(n8172), .ZN(n5417) );
  INV_X1 U6912 ( .A(n8171), .ZN(n5416) );
  NAND2_X2 U6913 ( .A1(n5419), .A2(n5418), .ZN(n8161) );
  INV_X1 U6914 ( .A(n5420), .ZN(n5424) );
  INV_X1 U6915 ( .A(n5421), .ZN(n5422) );
  NAND2_X1 U6916 ( .A1(n5422), .A2(SI_24_), .ZN(n5423) );
  INV_X1 U6917 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n7765) );
  INV_X1 U6918 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n5426) );
  MUX2_X1 U6919 ( .A(n7765), .B(n5426), .S(n4262), .Z(n5428) );
  INV_X1 U6920 ( .A(SI_25_), .ZN(n5427) );
  NAND2_X1 U6921 ( .A1(n5428), .A2(n5427), .ZN(n5443) );
  INV_X1 U6922 ( .A(n5428), .ZN(n5429) );
  NAND2_X1 U6923 ( .A1(n5429), .A2(SI_25_), .ZN(n5430) );
  NAND2_X1 U6924 ( .A1(n5443), .A2(n5430), .ZN(n5444) );
  NAND2_X1 U6925 ( .A1(n7722), .A2(n5633), .ZN(n5432) );
  NAND2_X1 U6926 ( .A1(n5634), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n5431) );
  XNOR2_X1 U6927 ( .A(n8481), .B(n5433), .ZN(n8159) );
  NAND2_X1 U6928 ( .A1(n5554), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n5435) );
  NAND2_X1 U6929 ( .A1(n4912), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n5434) );
  AND2_X1 U6930 ( .A1(n5435), .A2(n5434), .ZN(n5441) );
  INV_X1 U6931 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n5436) );
  NAND2_X1 U6932 ( .A1(n5437), .A2(n5436), .ZN(n5438) );
  NAND2_X1 U6933 ( .A1(n5454), .A2(n5438), .ZN(n8328) );
  INV_X1 U6934 ( .A(n5398), .ZN(n5553) );
  OR2_X1 U6935 ( .A1(n8328), .A2(n5553), .ZN(n5440) );
  NAND2_X1 U6936 ( .A1(n5475), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n5439) );
  INV_X1 U6937 ( .A(n8313), .ZN(n8230) );
  NAND2_X1 U6938 ( .A1(n8230), .A2(n5641), .ZN(n8158) );
  INV_X1 U6939 ( .A(n8159), .ZN(n5442) );
  INV_X1 U6940 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n5447) );
  INV_X1 U6941 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n5446) );
  MUX2_X1 U6942 ( .A(n5447), .B(n5446), .S(n6597), .Z(n5449) );
  INV_X1 U6943 ( .A(SI_26_), .ZN(n5448) );
  NAND2_X1 U6944 ( .A1(n5449), .A2(n5448), .ZN(n5463) );
  INV_X1 U6945 ( .A(n5449), .ZN(n5450) );
  NAND2_X1 U6946 ( .A1(n5450), .A2(SI_26_), .ZN(n5451) );
  XNOR2_X1 U6947 ( .A(n5462), .B(n5461), .ZN(n7778) );
  NAND2_X1 U6948 ( .A1(n7778), .A2(n5633), .ZN(n5453) );
  NAND2_X1 U6949 ( .A1(n5634), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n5452) );
  XNOR2_X1 U6950 ( .A(n8477), .B(n5504), .ZN(n5459) );
  INV_X1 U6951 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n8219) );
  NAND2_X1 U6952 ( .A1(n5454), .A2(n8219), .ZN(n5455) );
  NAND2_X1 U6953 ( .A1(n5473), .A2(n5455), .ZN(n8218) );
  AOI22_X1 U6954 ( .A1(n4982), .A2(P2_REG2_REG_26__SCAN_IN), .B1(n5554), .B2(
        P2_REG0_REG_26__SCAN_IN), .ZN(n5457) );
  NAND2_X1 U6955 ( .A1(n5619), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n5456) );
  OAI211_X1 U6956 ( .C1(n8218), .C2(n5553), .A(n5457), .B(n5456), .ZN(n8300)
         );
  NAND2_X1 U6957 ( .A1(n8300), .A2(n5641), .ZN(n5458) );
  NOR2_X1 U6958 ( .A1(n5459), .A2(n5458), .ZN(n5460) );
  AOI21_X1 U6959 ( .B1(n5459), .B2(n5458), .A(n5460), .ZN(n8216) );
  INV_X1 U6960 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n5465) );
  INV_X1 U6961 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n5464) );
  MUX2_X1 U6962 ( .A(n5465), .B(n5464), .S(n6597), .Z(n5467) );
  INV_X1 U6963 ( .A(SI_27_), .ZN(n5466) );
  NAND2_X1 U6964 ( .A1(n5467), .A2(n5466), .ZN(n5488) );
  INV_X1 U6965 ( .A(n5467), .ZN(n5468) );
  NAND2_X1 U6966 ( .A1(n5468), .A2(SI_27_), .ZN(n5469) );
  NAND2_X1 U6967 ( .A1(n7805), .A2(n5633), .ZN(n5471) );
  NAND2_X1 U6968 ( .A1(n5634), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n5470) );
  XNOR2_X1 U6969 ( .A(n8470), .B(n5504), .ZN(n5483) );
  INV_X1 U6970 ( .A(n5473), .ZN(n5472) );
  NAND2_X1 U6971 ( .A1(n5472), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n5496) );
  INV_X1 U6972 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n9973) );
  NAND2_X1 U6973 ( .A1(n5473), .A2(n9973), .ZN(n5474) );
  NAND2_X1 U6974 ( .A1(n8294), .A2(n5398), .ZN(n5481) );
  INV_X1 U6975 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n5478) );
  NAND2_X1 U6976 ( .A1(n4912), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n5477) );
  NAND2_X1 U6977 ( .A1(n5554), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n5476) );
  OAI211_X1 U6978 ( .C1(n5478), .C2(n4933), .A(n5477), .B(n5476), .ZN(n5479)
         );
  INV_X1 U6979 ( .A(n5479), .ZN(n5480) );
  OR2_X1 U6980 ( .A1(n8314), .A2(n6866), .ZN(n5482) );
  NOR2_X1 U6981 ( .A1(n5483), .A2(n5482), .ZN(n5484) );
  AOI21_X1 U6982 ( .B1(n5483), .B2(n5482), .A(n5484), .ZN(n8094) );
  NAND2_X1 U6983 ( .A1(n8095), .A2(n8094), .ZN(n8093) );
  INV_X1 U6984 ( .A(n5484), .ZN(n5485) );
  INV_X1 U6985 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n5491) );
  INV_X1 U6986 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n5490) );
  MUX2_X1 U6987 ( .A(n5491), .B(n5490), .S(n6597), .Z(n5599) );
  XNOR2_X1 U6988 ( .A(n5599), .B(SI_28_), .ZN(n5596) );
  NAND2_X1 U6989 ( .A1(n7846), .A2(n5633), .ZN(n5493) );
  NAND2_X1 U6990 ( .A1(n5634), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n5492) );
  INV_X1 U6991 ( .A(n5496), .ZN(n5494) );
  NAND2_X1 U6992 ( .A1(n5494), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n8065) );
  INV_X1 U6993 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n5495) );
  NAND2_X1 U6994 ( .A1(n5496), .A2(n5495), .ZN(n5497) );
  NAND2_X1 U6995 ( .A1(n8065), .A2(n5497), .ZN(n5564) );
  INV_X1 U6996 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n5500) );
  NAND2_X1 U6997 ( .A1(n5554), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n5499) );
  NAND2_X1 U6998 ( .A1(n4912), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n5498) );
  OAI211_X1 U6999 ( .C1(n5500), .C2(n4933), .A(n5499), .B(n5498), .ZN(n5501)
         );
  INV_X1 U7000 ( .A(n5501), .ZN(n5502) );
  NAND2_X1 U7001 ( .A1(n8299), .A2(n5641), .ZN(n5505) );
  XNOR2_X1 U7002 ( .A(n5505), .B(n5504), .ZN(n5543) );
  INV_X1 U7003 ( .A(n5543), .ZN(n5544) );
  AND2_X1 U7004 ( .A1(n5295), .A2(n7419), .ZN(n5507) );
  NOR2_X1 U7005 ( .A1(n5508), .A2(n8552), .ZN(n5509) );
  MUX2_X1 U7006 ( .A(n8552), .B(n5509), .S(P2_IR_REG_25__SCAN_IN), .Z(n5510)
         );
  MUX2_X1 U7007 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5512), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n5514) );
  NOR2_X1 U7008 ( .A1(n7763), .A2(n5529), .ZN(n5522) );
  NAND2_X1 U7009 ( .A1(n5516), .A2(n5515), .ZN(n5517) );
  NAND2_X1 U7010 ( .A1(n5524), .A2(n5523), .ZN(n5518) );
  NAND2_X1 U7011 ( .A1(n5518), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5520) );
  INV_X1 U7012 ( .A(n7656), .ZN(n5521) );
  INV_X1 U7013 ( .A(n9714), .ZN(n5525) );
  INV_X1 U7014 ( .A(n5529), .ZN(n7779) );
  INV_X1 U7015 ( .A(P2_B_REG_SCAN_IN), .ZN(n5526) );
  XOR2_X1 U7016 ( .A(n7656), .B(n5526), .Z(n5527) );
  NAND2_X1 U7017 ( .A1(n7763), .A2(n5527), .ZN(n5528) );
  INV_X1 U7018 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n9711) );
  AND2_X1 U7019 ( .A1(n7656), .A2(n5529), .ZN(n9710) );
  AND2_X1 U7020 ( .A1(n7763), .A2(n5529), .ZN(n9713) );
  AOI21_X1 U7021 ( .B1(n9708), .B2(n9978), .A(n9713), .ZN(n6763) );
  NOR4_X1 U7022 ( .A1(P2_D_REG_17__SCAN_IN), .A2(P2_D_REG_18__SCAN_IN), .A3(
        P2_D_REG_19__SCAN_IN), .A4(P2_D_REG_20__SCAN_IN), .ZN(n5533) );
  NOR4_X1 U7023 ( .A1(P2_D_REG_15__SCAN_IN), .A2(P2_D_REG_12__SCAN_IN), .A3(
        P2_D_REG_14__SCAN_IN), .A4(P2_D_REG_16__SCAN_IN), .ZN(n5532) );
  NOR4_X1 U7024 ( .A1(P2_D_REG_26__SCAN_IN), .A2(P2_D_REG_27__SCAN_IN), .A3(
        P2_D_REG_28__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n5531) );
  NOR4_X1 U7025 ( .A1(P2_D_REG_21__SCAN_IN), .A2(P2_D_REG_23__SCAN_IN), .A3(
        P2_D_REG_24__SCAN_IN), .A4(P2_D_REG_25__SCAN_IN), .ZN(n5530) );
  NAND4_X1 U7026 ( .A1(n5533), .A2(n5532), .A3(n5531), .A4(n5530), .ZN(n5538)
         );
  NOR2_X1 U7027 ( .A1(P2_D_REG_11__SCAN_IN), .A2(P2_D_REG_22__SCAN_IN), .ZN(
        n9968) );
  NOR4_X1 U7028 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        P2_D_REG_13__SCAN_IN), .A4(P2_D_REG_2__SCAN_IN), .ZN(n5536) );
  NOR4_X1 U7029 ( .A1(P2_D_REG_7__SCAN_IN), .A2(P2_D_REG_8__SCAN_IN), .A3(
        P2_D_REG_9__SCAN_IN), .A4(P2_D_REG_10__SCAN_IN), .ZN(n5535) );
  NOR4_X1 U7030 ( .A1(P2_D_REG_3__SCAN_IN), .A2(P2_D_REG_4__SCAN_IN), .A3(
        P2_D_REG_5__SCAN_IN), .A4(P2_D_REG_6__SCAN_IN), .ZN(n5534) );
  NAND4_X1 U7031 ( .A1(n9968), .A2(n5536), .A3(n5535), .A4(n5534), .ZN(n5537)
         );
  OAI21_X1 U7032 ( .B1(n5538), .B2(n5537), .A(n9708), .ZN(n6761) );
  NAND2_X1 U7033 ( .A1(n6763), .A2(n6761), .ZN(n7024) );
  INV_X1 U7034 ( .A(n7024), .ZN(n5539) );
  AND2_X1 U7035 ( .A1(n7025), .A2(n5539), .ZN(n5565) );
  AND2_X1 U7036 ( .A1(n5565), .A2(n6759), .ZN(n5563) );
  NOR2_X1 U7037 ( .A1(n5506), .A2(n9715), .ZN(n7036) );
  NAND2_X1 U7038 ( .A1(n5563), .A2(n7036), .ZN(n5540) );
  NOR3_X1 U7039 ( .A1(n4501), .A2(n8207), .A3(n5544), .ZN(n5541) );
  AOI21_X1 U7040 ( .B1(n4501), .B2(n5544), .A(n5541), .ZN(n5542) );
  NOR3_X1 U7041 ( .A1(n4501), .A2(n5543), .A3(n8207), .ZN(n5546) );
  NOR2_X1 U7042 ( .A1(n8466), .A2(n5544), .ZN(n5545) );
  INV_X1 U7043 ( .A(n8207), .ZN(n8227) );
  INV_X1 U7044 ( .A(n5567), .ZN(n6772) );
  NAND2_X1 U7045 ( .A1(n5563), .A2(n6772), .ZN(n5549) );
  OAI21_X1 U7046 ( .B1(n4501), .B2(n8227), .A(n8189), .ZN(n5550) );
  NAND3_X1 U7047 ( .A1(n5552), .A2(n5551), .A3(n5550), .ZN(n5574) );
  OR2_X1 U7048 ( .A1(n8065), .A2(n5553), .ZN(n5559) );
  INV_X1 U7049 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n9938) );
  NAND2_X1 U7050 ( .A1(n4982), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n5556) );
  NAND2_X1 U7051 ( .A1(n5554), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n5555) );
  OAI211_X1 U7052 ( .C1(n9938), .C2(n4933), .A(n5556), .B(n5555), .ZN(n5557)
         );
  INV_X1 U7053 ( .A(n5557), .ZN(n5558) );
  INV_X1 U7054 ( .A(n5560), .ZN(n7849) );
  OR2_X1 U7055 ( .A1(n8314), .A2(n9758), .ZN(n5561) );
  OAI21_X1 U7056 ( .B1(n6758), .B2(n9756), .A(n5561), .ZN(n8283) );
  INV_X1 U7057 ( .A(n8283), .ZN(n5571) );
  INV_X1 U7058 ( .A(n5829), .ZN(n5562) );
  NAND2_X1 U7059 ( .A1(n5563), .A2(n5562), .ZN(n6979) );
  INV_X1 U7060 ( .A(n5564), .ZN(n8279) );
  INV_X1 U7061 ( .A(n5565), .ZN(n5566) );
  NAND2_X1 U7062 ( .A1(n6762), .A2(n5566), .ZN(n6865) );
  INV_X1 U7063 ( .A(n6687), .ZN(n5568) );
  NAND2_X1 U7064 ( .A1(n5829), .A2(n5567), .ZN(n6760) );
  NAND4_X1 U7065 ( .A1(n6865), .A2(n5568), .A3(n5826), .A4(n6760), .ZN(n5569)
         );
  AOI22_X1 U7066 ( .A1(n8279), .A2(n8224), .B1(P2_REG3_REG_28__SCAN_IN), .B2(
        P2_U3152), .ZN(n5570) );
  OAI21_X1 U7067 ( .B1(n5571), .B2(n6979), .A(n5570), .ZN(n5572) );
  NAND2_X1 U7068 ( .A1(n5574), .A2(n5573), .ZN(P2_U3222) );
  NAND2_X1 U7069 ( .A1(n7117), .A2(n5575), .ZN(n5793) );
  NAND2_X1 U7070 ( .A1(n5793), .A2(n6776), .ZN(n5652) );
  INV_X1 U7071 ( .A(n5576), .ZN(n8247) );
  NAND2_X1 U7072 ( .A1(n7114), .A2(n6955), .ZN(n5577) );
  NAND2_X1 U7073 ( .A1(n7116), .A2(n6962), .ZN(n5648) );
  INV_X1 U7074 ( .A(n7116), .ZN(n8246) );
  INV_X1 U7075 ( .A(n6962), .ZN(n7397) );
  NAND2_X1 U7076 ( .A1(n8246), .A2(n7397), .ZN(n5663) );
  INV_X1 U7077 ( .A(n6956), .ZN(n5796) );
  NAND2_X1 U7078 ( .A1(n5577), .A2(n5796), .ZN(n6958) );
  INV_X1 U7079 ( .A(n6978), .ZN(n8244) );
  NAND2_X1 U7080 ( .A1(n8244), .A2(n7052), .ZN(n5791) );
  INV_X1 U7081 ( .A(n6954), .ZN(n8245) );
  NAND2_X1 U7082 ( .A1(n8245), .A2(n7039), .ZN(n6882) );
  AND2_X1 U7083 ( .A1(n5791), .A2(n6882), .ZN(n5664) );
  NAND2_X1 U7084 ( .A1(n6883), .A2(n5664), .ZN(n6910) );
  NAND2_X1 U7085 ( .A1(n6978), .A2(n6986), .ZN(n6908) );
  NAND2_X1 U7086 ( .A1(n6910), .A2(n6908), .ZN(n5578) );
  INV_X1 U7087 ( .A(n8084), .ZN(n8243) );
  XNOR2_X1 U7088 ( .A(n8243), .B(n7156), .ZN(n6907) );
  INV_X1 U7089 ( .A(n8139), .ZN(n8242) );
  INV_X1 U7090 ( .A(n8087), .ZN(n9735) );
  NAND2_X1 U7091 ( .A1(n8242), .A2(n9735), .ZN(n5686) );
  NAND2_X1 U7092 ( .A1(n9759), .A2(n8142), .ZN(n9751) );
  INV_X1 U7093 ( .A(n9759), .ZN(n8241) );
  INV_X1 U7094 ( .A(n8142), .ZN(n9743) );
  NAND2_X1 U7095 ( .A1(n8241), .A2(n9743), .ZN(n5676) );
  NAND2_X1 U7096 ( .A1(n7406), .A2(n7407), .ZN(n7405) );
  NAND2_X1 U7097 ( .A1(n7405), .A2(n9751), .ZN(n5579) );
  NAND2_X1 U7098 ( .A1(n8138), .A2(n9995), .ZN(n5689) );
  INV_X1 U7099 ( .A(n8138), .ZN(n8240) );
  INV_X1 U7100 ( .A(n9995), .ZN(n9767) );
  NAND2_X1 U7101 ( .A1(n8240), .A2(n9767), .ZN(n5678) );
  NAND2_X1 U7102 ( .A1(n5579), .A2(n9749), .ZN(n9755) );
  NAND2_X1 U7103 ( .A1(n9755), .A2(n5689), .ZN(n7208) );
  INV_X1 U7104 ( .A(n8115), .ZN(n9772) );
  INV_X1 U7105 ( .A(n9757), .ZN(n8239) );
  NAND2_X1 U7106 ( .A1(n9772), .A2(n8239), .ZN(n5803) );
  NAND2_X1 U7107 ( .A1(n9757), .A2(n8115), .ZN(n5804) );
  NAND2_X1 U7108 ( .A1(n8208), .A2(n8112), .ZN(n5801) );
  INV_X1 U7109 ( .A(n5801), .ZN(n5580) );
  OR2_X1 U7110 ( .A1(n8112), .A2(n8208), .ZN(n5802) );
  OR2_X1 U7111 ( .A1(n9786), .A2(n8204), .ZN(n5807) );
  INV_X1 U7112 ( .A(n5807), .ZN(n5698) );
  NAND2_X1 U7113 ( .A1(n9786), .A2(n8204), .ZN(n5806) );
  OR2_X1 U7114 ( .A1(n7587), .A2(n7746), .ZN(n5703) );
  NAND2_X1 U7115 ( .A1(n7587), .A2(n7746), .ZN(n5702) );
  AND2_X2 U7116 ( .A1(n5703), .A2(n5702), .ZN(n7558) );
  NAND2_X1 U7117 ( .A1(n7559), .A2(n7558), .ZN(n5581) );
  NAND2_X1 U7118 ( .A1(n5581), .A2(n5702), .ZN(n7581) );
  OR2_X1 U7119 ( .A1(n7657), .A2(n7818), .ZN(n5707) );
  NAND2_X1 U7120 ( .A1(n7657), .A2(n7818), .ZN(n5706) );
  NAND2_X1 U7121 ( .A1(n5707), .A2(n5706), .ZN(n7579) );
  OR2_X2 U7122 ( .A1(n7581), .A2(n7579), .ZN(n7582) );
  XNOR2_X1 U7123 ( .A(n7820), .B(n7840), .ZN(n7757) );
  INV_X1 U7124 ( .A(n7757), .ZN(n7661) );
  INV_X1 U7125 ( .A(n7820), .ZN(n9401) );
  NAND2_X1 U7126 ( .A1(n9401), .A2(n8234), .ZN(n5582) );
  INV_X1 U7127 ( .A(n8233), .ZN(n7801) );
  NAND2_X1 U7128 ( .A1(n8530), .A2(n7801), .ZN(n5583) );
  NAND2_X1 U7129 ( .A1(n8526), .A2(n7828), .ZN(n5719) );
  INV_X1 U7130 ( .A(n8425), .ZN(n8127) );
  OR2_X1 U7131 ( .A1(n8519), .A2(n8127), .ZN(n5724) );
  NAND2_X1 U7132 ( .A1(n8519), .A2(n8127), .ZN(n5726) );
  INV_X1 U7133 ( .A(n8446), .ZN(n8186) );
  OR2_X1 U7134 ( .A1(n8515), .A2(n8186), .ZN(n5725) );
  NAND2_X1 U7135 ( .A1(n8515), .A2(n8186), .ZN(n8408) );
  NAND2_X1 U7136 ( .A1(n8509), .A2(n8154), .ZN(n5739) );
  INV_X1 U7137 ( .A(n8418), .ZN(n5585) );
  INV_X1 U7138 ( .A(n8408), .ZN(n5735) );
  NOR2_X1 U7139 ( .A1(n5585), .A2(n5735), .ZN(n5586) );
  NAND2_X1 U7140 ( .A1(n8407), .A2(n5586), .ZN(n5587) );
  NAND2_X1 U7141 ( .A1(n5587), .A2(n5738), .ZN(n8397) );
  INV_X1 U7142 ( .A(n8410), .ZN(n8384) );
  OR2_X1 U7143 ( .A1(n8502), .A2(n8384), .ZN(n5742) );
  NAND2_X1 U7144 ( .A1(n8502), .A2(n8384), .ZN(n8378) );
  NAND2_X1 U7145 ( .A1(n5742), .A2(n8378), .ZN(n8398) );
  OR2_X2 U7146 ( .A1(n8397), .A2(n8398), .ZN(n8399) );
  NAND2_X1 U7147 ( .A1(n8497), .A2(n8361), .ZN(n5733) );
  NAND2_X1 U7148 ( .A1(n8356), .A2(n5733), .ZN(n8382) );
  INV_X1 U7149 ( .A(n8378), .ZN(n5588) );
  NOR2_X1 U7150 ( .A1(n8382), .A2(n5588), .ZN(n5589) );
  NAND2_X2 U7151 ( .A1(n8399), .A2(n5589), .ZN(n8379) );
  OR2_X1 U7152 ( .A1(n8367), .A2(n8383), .ZN(n5750) );
  NAND2_X1 U7153 ( .A1(n8367), .A2(n8383), .ZN(n5748) );
  NAND2_X1 U7154 ( .A1(n5750), .A2(n5748), .ZN(n8357) );
  INV_X1 U7155 ( .A(n8356), .ZN(n5729) );
  NOR2_X1 U7156 ( .A1(n8357), .A2(n5729), .ZN(n5590) );
  NAND2_X2 U7157 ( .A1(n8379), .A2(n5590), .ZN(n8359) );
  NAND2_X1 U7158 ( .A1(n8486), .A2(n8362), .ZN(n5754) );
  NAND2_X1 U7159 ( .A1(n5752), .A2(n5754), .ZN(n8344) );
  NAND2_X1 U7160 ( .A1(n8481), .A2(n8313), .ZN(n5759) );
  NAND2_X1 U7161 ( .A1(n5757), .A2(n5759), .ZN(n8332) );
  INV_X1 U7162 ( .A(n8332), .ZN(n5814) );
  INV_X1 U7163 ( .A(n8310), .ZN(n5593) );
  INV_X1 U7164 ( .A(n8300), .ZN(n8096) );
  OR2_X1 U7165 ( .A1(n8477), .A2(n8096), .ZN(n5761) );
  NAND2_X1 U7166 ( .A1(n8477), .A2(n8096), .ZN(n5760) );
  OR2_X1 U7167 ( .A1(n8470), .A2(n8314), .ZN(n5594) );
  NAND2_X1 U7168 ( .A1(n8466), .A2(n8299), .ZN(n5595) );
  INV_X1 U7169 ( .A(n8281), .ZN(n5769) );
  INV_X1 U7170 ( .A(n8299), .ZN(n8097) );
  INV_X1 U7171 ( .A(SI_28_), .ZN(n5598) );
  NAND2_X1 U7172 ( .A1(n5599), .A2(n5598), .ZN(n5600) );
  INV_X1 U7173 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n5603) );
  INV_X1 U7174 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n5602) );
  MUX2_X1 U7175 ( .A(n5603), .B(n5602), .S(n6597), .Z(n5608) );
  XNOR2_X1 U7176 ( .A(n5608), .B(SI_29_), .ZN(n5604) );
  NAND2_X1 U7177 ( .A1(n8555), .A2(n5633), .ZN(n5606) );
  NAND2_X1 U7178 ( .A1(n5634), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n5605) );
  NAND2_X1 U7179 ( .A1(n8460), .A2(n6758), .ZN(n5776) );
  INV_X1 U7180 ( .A(SI_29_), .ZN(n5607) );
  AND2_X1 U7181 ( .A1(n5608), .A2(n5607), .ZN(n5611) );
  INV_X1 U7182 ( .A(n5608), .ZN(n5609) );
  NAND2_X1 U7183 ( .A1(n5609), .A2(SI_29_), .ZN(n5610) );
  MUX2_X1 U7184 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(P2_DATAO_REG_30__SCAN_IN), 
        .S(n6597), .Z(n5628) );
  NAND2_X1 U7185 ( .A1(n8717), .A2(n5633), .ZN(n5614) );
  NAND2_X1 U7186 ( .A1(n5634), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n5613) );
  NAND2_X1 U7187 ( .A1(n5475), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n5617) );
  NAND2_X1 U7188 ( .A1(n5554), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n5616) );
  NAND2_X1 U7189 ( .A1(n4912), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n5615) );
  AND3_X1 U7190 ( .A1(n5617), .A2(n5616), .A3(n5615), .ZN(n5638) );
  NAND2_X1 U7191 ( .A1(n5638), .A2(n5821), .ZN(n5623) );
  OAI21_X1 U7192 ( .B1(n8459), .B2(n5623), .A(n5776), .ZN(n5618) );
  INV_X1 U7193 ( .A(P2_REG2_REG_30__SCAN_IN), .ZN(n5622) );
  NAND2_X1 U7194 ( .A1(n5554), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n5621) );
  NAND2_X1 U7195 ( .A1(n5619), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n5620) );
  OAI211_X1 U7196 ( .C1(n5030), .C2(n5622), .A(n5621), .B(n5620), .ZN(n8228)
         );
  INV_X1 U7197 ( .A(n8228), .ZN(n5637) );
  NAND2_X1 U7198 ( .A1(n5625), .A2(n5624), .ZN(n5639) );
  INV_X1 U7199 ( .A(SI_30_), .ZN(n5626) );
  NAND2_X1 U7200 ( .A1(n5629), .A2(n5628), .ZN(n5630) );
  MUX2_X1 U7201 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(P2_DATAO_REG_31__SCAN_IN), 
        .S(n6597), .Z(n5631) );
  XNOR2_X1 U7202 ( .A(n5631), .B(SI_31_), .ZN(n5632) );
  NAND2_X1 U7203 ( .A1(n8551), .A2(n5633), .ZN(n5636) );
  NAND2_X1 U7204 ( .A1(n5634), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(n5635) );
  NOR2_X1 U7205 ( .A1(n8453), .A2(n5638), .ZN(n5784) );
  AND2_X1 U7206 ( .A1(n8269), .A2(n5637), .ZN(n5644) );
  NOR2_X1 U7207 ( .A1(n5784), .A2(n5644), .ZN(n5817) );
  INV_X1 U7208 ( .A(n8453), .ZN(n8265) );
  INV_X1 U7209 ( .A(n5638), .ZN(n8264) );
  AOI21_X1 U7210 ( .B1(n5639), .B2(n5817), .A(n5783), .ZN(n5640) );
  XNOR2_X1 U7211 ( .A(n5640), .B(n5295), .ZN(n5643) );
  INV_X1 U7212 ( .A(n5506), .ZN(n5820) );
  NAND2_X1 U7213 ( .A1(n5820), .A2(n5821), .ZN(n6778) );
  INV_X1 U7214 ( .A(n5644), .ZN(n5780) );
  OR2_X1 U7215 ( .A1(n5830), .A2(n7380), .ZN(n5646) );
  OR2_X1 U7216 ( .A1(n5645), .A2(n5646), .ZN(n5785) );
  AND2_X1 U7217 ( .A1(n5801), .A2(n5804), .ZN(n5685) );
  AND2_X1 U7218 ( .A1(n6908), .A2(n5790), .ZN(n5647) );
  MUX2_X1 U7219 ( .A(n5664), .B(n5647), .S(n5749), .Z(n5662) );
  NAND2_X1 U7220 ( .A1(n5790), .A2(n5648), .ZN(n5650) );
  NAND2_X1 U7221 ( .A1(n6908), .A2(n5671), .ZN(n5649) );
  AOI21_X1 U7222 ( .B1(n5662), .B2(n5650), .A(n5649), .ZN(n5656) );
  NAND2_X1 U7223 ( .A1(n6779), .A2(n4505), .ZN(n5792) );
  AND2_X1 U7224 ( .A1(n5792), .A2(n5821), .ZN(n5651) );
  OAI211_X1 U7225 ( .C1(n5652), .C2(n5651), .A(n5658), .B(n5794), .ZN(n5653)
         );
  NAND3_X1 U7226 ( .A1(n5653), .A2(n6955), .A3(n5785), .ZN(n5654) );
  NAND3_X1 U7227 ( .A1(n5662), .A2(n5796), .A3(n5654), .ZN(n5655) );
  OAI21_X1 U7228 ( .B1(n5656), .B2(n5749), .A(n5655), .ZN(n5661) );
  OR2_X1 U7229 ( .A1(n8084), .A2(n7156), .ZN(n5666) );
  NAND2_X1 U7230 ( .A1(n5794), .A2(n5792), .ZN(n5657) );
  NAND3_X1 U7231 ( .A1(n6955), .A2(n5793), .A3(n5657), .ZN(n5659) );
  NAND3_X1 U7232 ( .A1(n5659), .A2(n5749), .A3(n5658), .ZN(n5660) );
  NAND3_X1 U7233 ( .A1(n5661), .A2(n5666), .A3(n5660), .ZN(n5670) );
  INV_X1 U7234 ( .A(n5662), .ZN(n5665) );
  AOI22_X1 U7235 ( .A1(n5665), .A2(n5791), .B1(n5664), .B2(n5663), .ZN(n5668)
         );
  INV_X1 U7236 ( .A(n5666), .ZN(n5667) );
  OAI21_X1 U7237 ( .B1(n5668), .B2(n5667), .A(n5749), .ZN(n5669) );
  NAND2_X1 U7238 ( .A1(n5670), .A2(n5669), .ZN(n5674) );
  NOR2_X1 U7239 ( .A1(n5671), .A2(n5785), .ZN(n5672) );
  NAND2_X1 U7240 ( .A1(n5675), .A2(n5686), .ZN(n7197) );
  NOR2_X1 U7241 ( .A1(n5672), .A2(n7197), .ZN(n5673) );
  NAND2_X1 U7242 ( .A1(n5674), .A2(n5673), .ZN(n5687) );
  NAND3_X1 U7243 ( .A1(n5687), .A2(n7407), .A3(n5675), .ZN(n5677) );
  NAND3_X1 U7244 ( .A1(n5677), .A2(n5678), .A3(n5676), .ZN(n5683) );
  INV_X1 U7245 ( .A(n5678), .ZN(n5680) );
  NAND2_X1 U7246 ( .A1(n5804), .A2(n5689), .ZN(n5679) );
  MUX2_X1 U7247 ( .A(n5680), .B(n5679), .S(n5785), .Z(n5681) );
  NOR2_X1 U7248 ( .A1(n5681), .A2(n4687), .ZN(n5690) );
  NAND2_X1 U7249 ( .A1(n5802), .A2(n5803), .ZN(n5682) );
  AOI21_X1 U7250 ( .B1(n5683), .B2(n5690), .A(n5682), .ZN(n5684) );
  MUX2_X1 U7251 ( .A(n5685), .B(n5684), .S(n5785), .Z(n5697) );
  NAND3_X1 U7252 ( .A1(n5687), .A2(n7407), .A3(n5686), .ZN(n5688) );
  AOI21_X1 U7253 ( .B1(n5688), .B2(n9751), .A(n5785), .ZN(n5692) );
  INV_X1 U7254 ( .A(n5689), .ZN(n5691) );
  OAI21_X1 U7255 ( .B1(n5692), .B2(n5691), .A(n5690), .ZN(n5696) );
  NAND2_X1 U7256 ( .A1(n5807), .A2(n5802), .ZN(n5694) );
  NAND2_X1 U7257 ( .A1(n5806), .A2(n5801), .ZN(n5693) );
  MUX2_X1 U7258 ( .A(n5694), .B(n5693), .S(n5785), .Z(n5695) );
  AOI21_X1 U7259 ( .B1(n5697), .B2(n5696), .A(n5695), .ZN(n5701) );
  INV_X1 U7260 ( .A(n5806), .ZN(n5699) );
  MUX2_X1 U7261 ( .A(n5699), .B(n5698), .S(n5785), .Z(n5700) );
  OAI21_X1 U7262 ( .B1(n5701), .B2(n5700), .A(n7558), .ZN(n5705) );
  INV_X1 U7263 ( .A(n7579), .ZN(n7583) );
  MUX2_X1 U7264 ( .A(n5703), .B(n5702), .S(n5749), .Z(n5704) );
  NAND3_X1 U7265 ( .A1(n5705), .A2(n7583), .A3(n5704), .ZN(n5709) );
  MUX2_X1 U7266 ( .A(n5707), .B(n5706), .S(n5785), .Z(n5708) );
  NAND3_X1 U7267 ( .A1(n5709), .A2(n7661), .A3(n5708), .ZN(n5715) );
  NAND2_X1 U7268 ( .A1(n8530), .A2(n8233), .ZN(n7783) );
  OR2_X1 U7269 ( .A1(n8530), .A2(n8233), .ZN(n5710) );
  INV_X1 U7270 ( .A(n7759), .ZN(n5714) );
  OR2_X1 U7271 ( .A1(n7840), .A2(n5749), .ZN(n5712) );
  NAND2_X1 U7272 ( .A1(n7840), .A2(n5749), .ZN(n5711) );
  MUX2_X1 U7273 ( .A(n5712), .B(n5711), .S(n7820), .Z(n5713) );
  NAND3_X1 U7274 ( .A1(n5715), .A2(n5714), .A3(n5713), .ZN(n5718) );
  MUX2_X1 U7275 ( .A(n8233), .B(n8530), .S(n5785), .Z(n5716) );
  NAND2_X1 U7276 ( .A1(n5716), .A2(n7783), .ZN(n5717) );
  NAND3_X1 U7277 ( .A1(n5718), .A2(n7789), .A3(n5717), .ZN(n5723) );
  AND2_X1 U7278 ( .A1(n5726), .A2(n5719), .ZN(n5720) );
  MUX2_X1 U7279 ( .A(n5721), .B(n5720), .S(n5749), .Z(n5722) );
  NAND2_X1 U7280 ( .A1(n5723), .A2(n5722), .ZN(n5737) );
  NAND2_X1 U7281 ( .A1(n5725), .A2(n5724), .ZN(n5734) );
  AOI21_X1 U7282 ( .B1(n5737), .B2(n5726), .A(n5734), .ZN(n5728) );
  NAND2_X1 U7283 ( .A1(n5739), .A2(n8408), .ZN(n5727) );
  OAI211_X1 U7284 ( .C1(n5728), .C2(n5727), .A(n5738), .B(n5742), .ZN(n5731)
         );
  AND2_X1 U7285 ( .A1(n5733), .A2(n8378), .ZN(n5730) );
  AOI21_X1 U7286 ( .B1(n5731), .B2(n5730), .A(n5729), .ZN(n5732) );
  MUX2_X1 U7287 ( .A(n5733), .B(n5732), .S(n5785), .Z(n5746) );
  INV_X1 U7288 ( .A(n8357), .ZN(n5745) );
  INV_X1 U7289 ( .A(n5734), .ZN(n5736) );
  AOI21_X1 U7290 ( .B1(n5737), .B2(n5736), .A(n5735), .ZN(n5741) );
  INV_X1 U7291 ( .A(n5738), .ZN(n5740) );
  OAI211_X1 U7292 ( .C1(n5741), .C2(n5740), .A(n8378), .B(n5739), .ZN(n5743)
         );
  NAND4_X1 U7293 ( .A1(n5743), .A2(n5749), .A3(n8356), .A4(n5742), .ZN(n5744)
         );
  NAND3_X1 U7294 ( .A1(n5746), .A2(n5745), .A3(n5744), .ZN(n5747) );
  OAI211_X1 U7295 ( .C1(n5749), .C2(n5748), .A(n5747), .B(n5754), .ZN(n5753)
         );
  AOI21_X1 U7296 ( .B1(n5752), .B2(n5750), .A(n5785), .ZN(n5751) );
  AOI21_X1 U7297 ( .B1(n5753), .B2(n5752), .A(n5751), .ZN(n5756) );
  OAI21_X1 U7298 ( .B1(n5754), .B2(n5785), .A(n5814), .ZN(n5755) );
  OR3_X1 U7299 ( .A1(n5756), .A2(n8311), .A3(n5755), .ZN(n5766) );
  NAND2_X1 U7300 ( .A1(n5761), .A2(n5757), .ZN(n5758) );
  NAND2_X1 U7301 ( .A1(n5758), .A2(n5760), .ZN(n5764) );
  NAND2_X1 U7302 ( .A1(n5760), .A2(n5759), .ZN(n5762) );
  NAND2_X1 U7303 ( .A1(n5762), .A2(n5761), .ZN(n5763) );
  MUX2_X1 U7304 ( .A(n5764), .B(n5763), .S(n5785), .Z(n5765) );
  AOI21_X1 U7305 ( .B1(n5766), .B2(n5765), .A(n8298), .ZN(n5771) );
  NOR2_X1 U7306 ( .A1(n8314), .A2(n5785), .ZN(n5768) );
  AND2_X1 U7307 ( .A1(n8314), .A2(n5785), .ZN(n5767) );
  MUX2_X1 U7308 ( .A(n5768), .B(n5767), .S(n8470), .Z(n5770) );
  OAI21_X1 U7309 ( .B1(n5771), .B2(n5770), .A(n5769), .ZN(n5774) );
  OR3_X1 U7310 ( .A1(n8466), .A2(n8097), .A3(n5785), .ZN(n5773) );
  NAND3_X1 U7311 ( .A1(n8466), .A2(n8097), .A3(n5785), .ZN(n5772) );
  NAND3_X1 U7312 ( .A1(n5774), .A2(n5773), .A3(n5772), .ZN(n5775) );
  NAND2_X1 U7313 ( .A1(n5775), .A2(n8071), .ZN(n5779) );
  MUX2_X1 U7314 ( .A(n5777), .B(n5776), .S(n5785), .Z(n5778) );
  NAND3_X1 U7315 ( .A1(n5780), .A2(n5779), .A3(n5778), .ZN(n5782) );
  NOR2_X1 U7316 ( .A1(n5783), .A2(n4310), .ZN(n5818) );
  OAI21_X1 U7317 ( .B1(n4310), .B2(n5782), .A(n5781), .ZN(n5789) );
  INV_X1 U7318 ( .A(n5783), .ZN(n5787) );
  INV_X1 U7319 ( .A(n5784), .ZN(n5786) );
  INV_X1 U7320 ( .A(n5825), .ZN(n5824) );
  NAND2_X1 U7321 ( .A1(n5790), .A2(n6882), .ZN(n7021) );
  INV_X1 U7322 ( .A(n7021), .ZN(n7030) );
  NAND2_X1 U7323 ( .A1(n6908), .A2(n5791), .ZN(n6884) );
  AND2_X1 U7324 ( .A1(n6776), .A2(n5792), .ZN(n9716) );
  NAND4_X1 U7325 ( .A1(n7112), .A2(n7030), .A3(n4798), .A4(n9716), .ZN(n5798)
         );
  NAND2_X1 U7326 ( .A1(n5794), .A2(n5793), .ZN(n6769) );
  INV_X1 U7327 ( .A(n6769), .ZN(n5795) );
  NAND3_X1 U7328 ( .A1(n5796), .A2(n5795), .A3(n5820), .ZN(n5797) );
  NOR2_X1 U7329 ( .A1(n5798), .A2(n5797), .ZN(n5800) );
  INV_X1 U7330 ( .A(n7197), .ZN(n5799) );
  NAND4_X1 U7331 ( .A1(n5800), .A2(n5799), .A3(n7407), .A4(n6907), .ZN(n5805)
         );
  NAND2_X1 U7332 ( .A1(n5802), .A2(n5801), .ZN(n7257) );
  INV_X1 U7333 ( .A(n7209), .ZN(n7204) );
  INV_X1 U7334 ( .A(n9749), .ZN(n9752) );
  NOR4_X1 U7335 ( .A1(n5805), .A2(n7257), .A3(n7204), .A4(n9752), .ZN(n5808)
         );
  NAND4_X1 U7336 ( .A1(n5808), .A2(n7583), .A3(n7558), .A4(n9690), .ZN(n5809)
         );
  NOR3_X1 U7337 ( .A1(n7759), .A2(n7757), .A3(n5809), .ZN(n5810) );
  AND4_X1 U7338 ( .A1(n8424), .A2(n7789), .A3(n4825), .A4(n5810), .ZN(n5811)
         );
  NAND2_X1 U7339 ( .A1(n8418), .A2(n5811), .ZN(n5812) );
  NOR4_X1 U7340 ( .A1(n8357), .A2(n8382), .A3(n8398), .A4(n5812), .ZN(n5813)
         );
  NAND3_X1 U7341 ( .A1(n5814), .A2(n4677), .A3(n5813), .ZN(n5815) );
  NOR4_X1 U7342 ( .A1(n8281), .A2(n8298), .A3(n8311), .A4(n5815), .ZN(n5816)
         );
  NAND4_X1 U7343 ( .A1(n5818), .A2(n8071), .A3(n5817), .A4(n5816), .ZN(n5819)
         );
  XNOR2_X1 U7344 ( .A(n5819), .B(n5645), .ZN(n5822) );
  OAI22_X1 U7345 ( .A1(n5822), .A2(n5821), .B1(n5820), .B2(n6777), .ZN(n5823)
         );
  OR2_X1 U7346 ( .A1(n5826), .A2(P2_U3152), .ZN(n7575) );
  NOR4_X1 U7347 ( .A1(n5829), .A2(n9758), .A3(n9707), .A4(n5828), .ZN(n5832)
         );
  OAI21_X1 U7348 ( .B1(n7575), .B2(n5830), .A(P2_B_REG_SCAN_IN), .ZN(n5831) );
  OR2_X1 U7349 ( .A1(n5832), .A2(n5831), .ZN(n5833) );
  NAND3_X1 U7350 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .A3(P1_REG3_REG_5__SCAN_IN), .ZN(n5966) );
  INV_X1 U7351 ( .A(n5966), .ZN(n5834) );
  NAND2_X1 U7352 ( .A1(n5834), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n5979) );
  INV_X1 U7353 ( .A(n5979), .ZN(n5835) );
  NAND2_X1 U7354 ( .A1(n5835), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n5996) );
  INV_X1 U7355 ( .A(n5996), .ZN(n5836) );
  NAND2_X1 U7356 ( .A1(n5836), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n6007) );
  INV_X1 U7357 ( .A(n6051), .ZN(n5838) );
  NAND2_X1 U7358 ( .A1(n5838), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n6065) );
  INV_X1 U7359 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n8591) );
  INV_X1 U7360 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n8655) );
  INV_X1 U7361 ( .A(n6188), .ZN(n5844) );
  NAND2_X1 U7362 ( .A1(n5844), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n6199) );
  INV_X1 U7363 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n6198) );
  NAND2_X1 U7364 ( .A1(P1_REG3_REG_27__SCAN_IN), .A2(P1_REG3_REG_28__SCAN_IN), 
        .ZN(n5846) );
  NOR2_X2 U7365 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5927) );
  NAND2_X1 U7366 ( .A1(n5927), .A2(n5847), .ZN(n5946) );
  NAND2_X1 U7367 ( .A1(n6072), .A2(n5853), .ZN(n6074) );
  NAND2_X1 U7368 ( .A1(n9847), .A2(n6085), .ZN(n5855) );
  INV_X1 U7369 ( .A(n5863), .ZN(n5854) );
  NOR2_X2 U7370 ( .A1(n5880), .A2(P1_IR_REG_19__SCAN_IN), .ZN(n5877) );
  OR2_X2 U7371 ( .A1(n5877), .A2(n9380), .ZN(n5860) );
  NAND2_X1 U7372 ( .A1(n5860), .A2(n5861), .ZN(n5856) );
  NAND2_X1 U7373 ( .A1(n5859), .A2(n5875), .ZN(n5857) );
  XNOR2_X1 U7374 ( .A(n5858), .B(n5876), .ZN(n6309) );
  XNOR2_X1 U7375 ( .A(n5859), .B(P1_IR_REG_21__SCAN_IN), .ZN(n6304) );
  NOR2_X1 U7376 ( .A1(P1_IR_REG_14__SCAN_IN), .A2(P1_IR_REG_22__SCAN_IN), .ZN(
        n5862) );
  NAND4_X1 U7377 ( .A1(n5863), .A2(n5862), .A3(n5861), .A4(n6085), .ZN(n5865)
         );
  NAND4_X1 U7378 ( .A1(n9847), .A2(n9857), .A3(n5875), .A4(n5881), .ZN(n5864)
         );
  NOR2_X1 U7379 ( .A1(n5865), .A2(n5864), .ZN(n5866) );
  NAND2_X1 U7380 ( .A1(n4319), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5868) );
  NAND2_X1 U7381 ( .A1(n5868), .A2(n5885), .ZN(n5870) );
  OR2_X1 U7382 ( .A1(n5868), .A2(n5885), .ZN(n5869) );
  NAND2_X1 U7383 ( .A1(n5870), .A2(n5869), .ZN(n6264) );
  NAND2_X1 U7384 ( .A1(n5871), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5873) );
  XNOR2_X1 U7385 ( .A(n5873), .B(n5872), .ZN(n6249) );
  NOR2_X1 U7386 ( .A1(n6264), .A2(n6249), .ZN(n5874) );
  NAND4_X1 U7387 ( .A1(n5877), .A2(n5861), .A3(n5876), .A4(n5875), .ZN(n5878)
         );
  NAND2_X1 U7388 ( .A1(n5878), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5879) );
  NAND2_X1 U7389 ( .A1(n5880), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5882) );
  NAND2_X1 U7390 ( .A1(n9649), .A2(n9248), .ZN(n5883) );
  NAND2_X1 U7391 ( .A1(n5887), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5888) );
  MUX2_X1 U7392 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5888), .S(
        P1_IR_REG_29__SCAN_IN), .Z(n5890) );
  INV_X1 U7393 ( .A(n5889), .ZN(n9381) );
  INV_X1 U7394 ( .A(P1_REG2_REG_30__SCAN_IN), .ZN(n9062) );
  NAND2_X1 U7395 ( .A1(n6213), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n5893) );
  INV_X1 U7396 ( .A(n9386), .ZN(n5891) );
  NAND2_X1 U7397 ( .A1(n6629), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n5892) );
  OAI211_X1 U7398 ( .C1(n6226), .C2(n9062), .A(n5893), .B(n5892), .ZN(n9001)
         );
  INV_X1 U7399 ( .A(n9001), .ZN(n6243) );
  INV_X1 U7400 ( .A(n6805), .ZN(n8992) );
  INV_X1 U7401 ( .A(n5909), .ZN(n8993) );
  AOI21_X1 U7402 ( .B1(n8992), .B2(P1_B_REG_SCAN_IN), .A(n9586), .ZN(n9056) );
  INV_X1 U7403 ( .A(n9056), .ZN(n6242) );
  INV_X1 U7404 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n6581) );
  INV_X1 U7405 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n5897) );
  OAI21_X1 U7406 ( .B1(n6222), .B2(n6581), .A(n5897), .ZN(n5898) );
  NAND2_X1 U7407 ( .A1(n9078), .A2(n6223), .ZN(n5904) );
  INV_X1 U7408 ( .A(P1_REG2_REG_28__SCAN_IN), .ZN(n9080) );
  NAND2_X1 U7409 ( .A1(n6629), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n5901) );
  NAND2_X1 U7410 ( .A1(n6213), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n5900) );
  OAI211_X1 U7411 ( .C1(n9080), .C2(n6226), .A(n5901), .B(n5900), .ZN(n5902)
         );
  INV_X1 U7412 ( .A(n5902), .ZN(n5903) );
  INV_X1 U7413 ( .A(n6588), .ZN(n8815) );
  INV_X1 U7414 ( .A(n9233), .ZN(n6241) );
  NAND2_X1 U7415 ( .A1(n8997), .A2(n9248), .ZN(n5906) );
  NAND2_X1 U7416 ( .A1(n8951), .A2(n8942), .ZN(n5905) );
  INV_X1 U7417 ( .A(n9590), .ZN(n6240) );
  NAND2_X1 U7418 ( .A1(n6223), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n5908) );
  NAND2_X1 U7419 ( .A1(n6628), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n5907) );
  INV_X1 U7420 ( .A(n6603), .ZN(n5910) );
  INV_X1 U7421 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n5911) );
  NAND2_X1 U7422 ( .A1(n4265), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n5913) );
  NAND2_X1 U7423 ( .A1(n6223), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n5916) );
  NAND2_X1 U7424 ( .A1(n4264), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n5915) );
  NAND2_X1 U7425 ( .A1(n6597), .A2(SI_0_), .ZN(n5918) );
  XNOR2_X1 U7426 ( .A(n5918), .B(P2_DATAO_REG_0__SCAN_IN), .ZN(n9393) );
  MUX2_X1 U7427 ( .A(P1_IR_REG_0__SCAN_IN), .B(n9393), .S(n6590), .Z(n6311) );
  INV_X1 U7428 ( .A(n6311), .ZN(n6825) );
  NAND2_X1 U7429 ( .A1(n8824), .A2(n6823), .ZN(n5920) );
  INV_X1 U7430 ( .A(n6321), .ZN(n8039) );
  NAND2_X1 U7431 ( .A1(n8039), .A2(n6846), .ZN(n5919) );
  NAND2_X1 U7432 ( .A1(n6223), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n5925) );
  NAND2_X1 U7433 ( .A1(n5921), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n5924) );
  NAND2_X1 U7434 ( .A1(n4263), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n5923) );
  NAND2_X1 U7435 ( .A1(n4265), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n5922) );
  NAND2_X1 U7436 ( .A1(n5957), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n5929) );
  OR2_X1 U7437 ( .A1(n5927), .A2(n9380), .ZN(n5936) );
  XNOR2_X1 U7438 ( .A(n5936), .B(P1_IR_REG_2__SCAN_IN), .ZN(n6650) );
  NAND2_X1 U7439 ( .A1(n6132), .A2(n6650), .ZN(n5928) );
  NAND2_X1 U7440 ( .A1(n7104), .A2(n8666), .ZN(n8954) );
  NAND2_X1 U7441 ( .A1(n9020), .A2(n6838), .ZN(n8959) );
  NAND2_X1 U7442 ( .A1(n8956), .A2(n8825), .ZN(n5930) );
  NAND2_X1 U7443 ( .A1(n5930), .A2(n8954), .ZN(n8911) );
  INV_X1 U7444 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n7099) );
  NAND2_X1 U7445 ( .A1(n6223), .A2(n7099), .ZN(n5934) );
  NAND2_X1 U7446 ( .A1(n5921), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n5933) );
  NAND2_X1 U7447 ( .A1(n4264), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n5932) );
  NAND2_X1 U7448 ( .A1(n4265), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n5931) );
  INV_X1 U7449 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n5935) );
  NAND2_X1 U7450 ( .A1(n5936), .A2(n5935), .ZN(n5937) );
  NAND2_X1 U7451 ( .A1(n5937), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5938) );
  XNOR2_X1 U7452 ( .A(n5938), .B(P1_IR_REG_3__SCAN_IN), .ZN(n6719) );
  NAND2_X1 U7453 ( .A1(n6132), .A2(n6719), .ZN(n5939) );
  NAND2_X1 U7454 ( .A1(n6992), .A2(n7100), .ZN(n8957) );
  INV_X1 U7455 ( .A(n6992), .ZN(n9019) );
  NAND2_X1 U7456 ( .A1(n9019), .A2(n9650), .ZN(n8907) );
  NAND2_X1 U7457 ( .A1(n8957), .A2(n8907), .ZN(n7102) );
  INV_X1 U7458 ( .A(n7102), .ZN(n8826) );
  NAND2_X1 U7459 ( .A1(n8911), .A2(n8826), .ZN(n5940) );
  NAND2_X1 U7460 ( .A1(n5921), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n5945) );
  NAND2_X1 U7461 ( .A1(n4265), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n5944) );
  INV_X1 U7462 ( .A(P1_REG3_REG_4__SCAN_IN), .ZN(n5941) );
  XNOR2_X1 U7463 ( .A(n5941), .B(P1_REG3_REG_3__SCAN_IN), .ZN(n8638) );
  NAND2_X1 U7464 ( .A1(n6223), .A2(n8638), .ZN(n5943) );
  NAND2_X1 U7465 ( .A1(n4263), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n5942) );
  INV_X1 U7466 ( .A(n7103), .ZN(n9018) );
  NAND2_X1 U7467 ( .A1(n5957), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n5949) );
  NAND2_X1 U7468 ( .A1(n5946), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5947) );
  XNOR2_X1 U7469 ( .A(n5947), .B(P1_IR_REG_4__SCAN_IN), .ZN(n9470) );
  NAND2_X1 U7470 ( .A1(n6132), .A2(n9470), .ZN(n5948) );
  INV_X1 U7471 ( .A(n6996), .ZN(n8636) );
  NAND2_X1 U7472 ( .A1(n9018), .A2(n8636), .ZN(n8908) );
  NAND2_X1 U7473 ( .A1(n5921), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n5956) );
  NAND2_X1 U7474 ( .A1(n4265), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n5955) );
  INV_X1 U7475 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n5951) );
  NAND2_X1 U7476 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .ZN(n5950) );
  NAND2_X1 U7477 ( .A1(n5951), .A2(n5950), .ZN(n5952) );
  AND2_X1 U7478 ( .A1(n5966), .A2(n5952), .ZN(n7129) );
  NAND2_X1 U7479 ( .A1(n6223), .A2(n7129), .ZN(n5954) );
  NAND2_X1 U7480 ( .A1(n4263), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n5953) );
  NAND2_X1 U7481 ( .A1(n8718), .A2(P2_DATAO_REG_5__SCAN_IN), .ZN(n5965) );
  NAND2_X1 U7482 ( .A1(n5958), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5959) );
  MUX2_X1 U7483 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5959), .S(
        P1_IR_REG_5__SCAN_IN), .Z(n5963) );
  INV_X1 U7484 ( .A(n5961), .ZN(n5962) );
  NAND2_X1 U7485 ( .A1(n6132), .A2(n9478), .ZN(n5964) );
  OAI211_X1 U7486 ( .C1(n6014), .C2(n6606), .A(n5965), .B(n5964), .ZN(n7069)
         );
  NAND2_X1 U7487 ( .A1(n7294), .A2(n7069), .ZN(n8902) );
  NAND2_X1 U7488 ( .A1(n7103), .A2(n6996), .ZN(n8901) );
  NAND2_X1 U7489 ( .A1(n8902), .A2(n8901), .ZN(n8725) );
  NAND2_X1 U7490 ( .A1(n6213), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n5971) );
  NAND2_X1 U7491 ( .A1(n4265), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n5970) );
  INV_X1 U7492 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n7292) );
  NAND2_X1 U7493 ( .A1(n5966), .A2(n7292), .ZN(n5967) );
  AND2_X1 U7494 ( .A1(n5979), .A2(n5967), .ZN(n7293) );
  NAND2_X1 U7495 ( .A1(n6223), .A2(n7293), .ZN(n5969) );
  NAND2_X1 U7496 ( .A1(n4264), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n5968) );
  OR2_X1 U7497 ( .A1(n5961), .A2(n9380), .ZN(n5972) );
  AOI22_X1 U7498 ( .A1(n8718), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n6132), .B2(
        n9490), .ZN(n5974) );
  INV_X2 U7499 ( .A(n6014), .ZN(n8714) );
  NAND2_X1 U7500 ( .A1(n6608), .A2(n8714), .ZN(n5973) );
  NAND2_X1 U7501 ( .A1(n5974), .A2(n5973), .ZN(n7143) );
  NAND2_X1 U7502 ( .A1(n7185), .A2(n7143), .ZN(n8903) );
  INV_X1 U7503 ( .A(n8903), .ZN(n5975) );
  NOR2_X1 U7504 ( .A1(n8725), .A2(n5975), .ZN(n8964) );
  NAND2_X1 U7505 ( .A1(n8723), .A2(n8964), .ZN(n5977) );
  INV_X1 U7506 ( .A(n7069), .ZN(n9657) );
  NAND2_X1 U7507 ( .A1(n9017), .A2(n9657), .ZN(n8724) );
  INV_X1 U7508 ( .A(n8724), .ZN(n8728) );
  NAND2_X1 U7509 ( .A1(n8903), .A2(n8728), .ZN(n8962) );
  INV_X1 U7510 ( .A(n7185), .ZN(n9016) );
  NAND2_X1 U7511 ( .A1(n9016), .A2(n7299), .ZN(n8733) );
  AND2_X1 U7512 ( .A1(n8962), .A2(n8733), .ZN(n5976) );
  NAND2_X1 U7513 ( .A1(n5921), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n5984) );
  NAND2_X1 U7514 ( .A1(n4263), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n5983) );
  INV_X1 U7515 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n5978) );
  NAND2_X1 U7516 ( .A1(n5979), .A2(n5978), .ZN(n5980) );
  AND2_X1 U7517 ( .A1(n5996), .A2(n5980), .ZN(n7189) );
  NAND2_X1 U7518 ( .A1(n6223), .A2(n7189), .ZN(n5982) );
  NAND2_X1 U7519 ( .A1(n4265), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n5981) );
  NAND2_X1 U7520 ( .A1(n6611), .A2(n8714), .ZN(n5988) );
  INV_X1 U7521 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n5985) );
  NAND2_X1 U7522 ( .A1(n5961), .A2(n5985), .ZN(n5986) );
  NAND2_X1 U7523 ( .A1(n5986), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5989) );
  XNOR2_X1 U7524 ( .A(n5989), .B(P1_IR_REG_7__SCAN_IN), .ZN(n9498) );
  AOI22_X1 U7525 ( .A1(n8718), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n6132), .B2(
        n9498), .ZN(n5987) );
  NAND2_X1 U7526 ( .A1(n5988), .A2(n5987), .ZN(n7221) );
  NAND2_X1 U7527 ( .A1(n7307), .A2(n7221), .ZN(n8734) );
  INV_X1 U7528 ( .A(n7221), .ZN(n7192) );
  NAND2_X1 U7529 ( .A1(n7192), .A2(n9015), .ZN(n8735) );
  NAND2_X1 U7530 ( .A1(n8734), .A2(n8735), .ZN(n7183) );
  OR2_X1 U7531 ( .A1(n6619), .A2(n6014), .ZN(n5995) );
  INV_X1 U7532 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n9889) );
  NAND2_X1 U7533 ( .A1(n5989), .A2(n9889), .ZN(n5990) );
  NAND2_X1 U7534 ( .A1(n5990), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5992) );
  INV_X1 U7535 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n5991) );
  NAND2_X1 U7536 ( .A1(n5992), .A2(n5991), .ZN(n6002) );
  OR2_X1 U7537 ( .A1(n5992), .A2(n5991), .ZN(n5993) );
  AOI22_X1 U7538 ( .A1(n8718), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n6132), .B2(
        n9516), .ZN(n5994) );
  NAND2_X1 U7539 ( .A1(n5995), .A2(n5994), .ZN(n7267) );
  NAND2_X1 U7540 ( .A1(n6629), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n6001) );
  NAND2_X1 U7541 ( .A1(n5921), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n6000) );
  INV_X1 U7542 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n7305) );
  NAND2_X1 U7543 ( .A1(n5996), .A2(n7305), .ZN(n5997) );
  AND2_X1 U7544 ( .A1(n6007), .A2(n5997), .ZN(n7306) );
  NAND2_X1 U7545 ( .A1(n6223), .A2(n7306), .ZN(n5999) );
  NAND2_X1 U7546 ( .A1(n4264), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n5998) );
  OR2_X1 U7547 ( .A1(n7267), .A2(n9588), .ZN(n8742) );
  NAND2_X1 U7548 ( .A1(n7267), .A2(n9588), .ZN(n8744) );
  NAND2_X1 U7549 ( .A1(n6622), .A2(n8714), .ZN(n6005) );
  NAND2_X1 U7550 ( .A1(n6002), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6003) );
  XNOR2_X1 U7551 ( .A(n6003), .B(P1_IR_REG_9__SCAN_IN), .ZN(n9528) );
  AOI22_X1 U7552 ( .A1(n8718), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n6132), .B2(
        n9528), .ZN(n6004) );
  NAND2_X1 U7553 ( .A1(n6005), .A2(n6004), .ZN(n6382) );
  NAND2_X1 U7554 ( .A1(n6007), .A2(n6006), .ZN(n6008) );
  AND2_X1 U7555 ( .A1(n6022), .A2(n6008), .ZN(n9596) );
  NAND2_X1 U7556 ( .A1(n6223), .A2(n9596), .ZN(n6012) );
  NAND2_X1 U7557 ( .A1(n6213), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n6011) );
  NAND2_X1 U7558 ( .A1(n4263), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n6010) );
  NAND2_X1 U7559 ( .A1(n6629), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n6009) );
  NAND4_X1 U7560 ( .A1(n6012), .A2(n6011), .A3(n6010), .A4(n6009), .ZN(n9013)
         );
  INV_X1 U7561 ( .A(n9013), .ZN(n7498) );
  NAND2_X1 U7562 ( .A1(n6382), .A2(n7498), .ZN(n8834) );
  NAND2_X1 U7563 ( .A1(n9585), .A2(n8834), .ZN(n6013) );
  OR2_X1 U7564 ( .A1(n6382), .A2(n7498), .ZN(n8835) );
  NAND2_X1 U7565 ( .A1(n6626), .A2(n8714), .ZN(n6020) );
  NOR2_X1 U7566 ( .A1(P1_IR_REG_7__SCAN_IN), .A2(P1_IR_REG_9__SCAN_IN), .ZN(
        n6015) );
  AND2_X1 U7567 ( .A1(n6016), .A2(n6015), .ZN(n6017) );
  NAND2_X1 U7568 ( .A1(n5961), .A2(n6017), .ZN(n6029) );
  NAND2_X1 U7569 ( .A1(n6029), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6018) );
  XNOR2_X1 U7570 ( .A(n6018), .B(P1_IR_REG_10__SCAN_IN), .ZN(n6942) );
  AOI22_X1 U7571 ( .A1(n8718), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n6132), .B2(
        n6942), .ZN(n6019) );
  NAND2_X1 U7572 ( .A1(n6213), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n6027) );
  NAND2_X1 U7573 ( .A1(n4264), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n6026) );
  NAND2_X1 U7574 ( .A1(n6022), .A2(n6021), .ZN(n6023) );
  AND2_X1 U7575 ( .A1(n6034), .A2(n6023), .ZN(n7504) );
  NAND2_X1 U7576 ( .A1(n6223), .A2(n7504), .ZN(n6025) );
  NAND2_X1 U7577 ( .A1(n6629), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n6024) );
  XNOR2_X1 U7578 ( .A(n7505), .B(n9587), .ZN(n8836) );
  OR2_X1 U7579 ( .A1(n7505), .A2(n9587), .ZN(n8746) );
  INV_X1 U7580 ( .A(n8834), .ZN(n8747) );
  NAND2_X1 U7581 ( .A1(n8746), .A2(n8747), .ZN(n6028) );
  NAND2_X1 U7582 ( .A1(n7505), .A2(n9587), .ZN(n8748) );
  AND2_X1 U7583 ( .A1(n6028), .A2(n8748), .ZN(n8894) );
  NAND2_X1 U7584 ( .A1(n6637), .A2(n8714), .ZN(n6032) );
  NAND2_X1 U7585 ( .A1(n6042), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6030) );
  XNOR2_X1 U7586 ( .A(n6030), .B(P1_IR_REG_11__SCAN_IN), .ZN(n9536) );
  AOI22_X1 U7587 ( .A1(n8718), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n6132), .B2(
        n9536), .ZN(n6031) );
  NAND2_X1 U7588 ( .A1(n6629), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n6039) );
  NAND2_X1 U7589 ( .A1(n6213), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n6038) );
  INV_X1 U7590 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n6033) );
  NAND2_X1 U7591 ( .A1(n6034), .A2(n6033), .ZN(n6035) );
  AND2_X1 U7592 ( .A1(n6051), .A2(n6035), .ZN(n7546) );
  NAND2_X1 U7593 ( .A1(n6223), .A2(n7546), .ZN(n6037) );
  NAND2_X1 U7594 ( .A1(n4263), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n6036) );
  NAND4_X1 U7595 ( .A1(n6039), .A2(n6038), .A3(n6037), .A4(n6036), .ZN(n9011)
         );
  OR2_X1 U7596 ( .A1(n7428), .A2(n7634), .ZN(n6040) );
  NAND2_X1 U7597 ( .A1(n7425), .A2(n6040), .ZN(n6041) );
  NAND2_X1 U7598 ( .A1(n7428), .A2(n7634), .ZN(n6057) );
  NAND2_X1 U7599 ( .A1(n6041), .A2(n6057), .ZN(n7486) );
  NAND2_X1 U7600 ( .A1(n6683), .A2(n8714), .ZN(n6049) );
  NAND2_X1 U7601 ( .A1(n6043), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6046) );
  INV_X1 U7602 ( .A(n6046), .ZN(n6044) );
  NAND2_X1 U7603 ( .A1(n6044), .A2(P1_IR_REG_12__SCAN_IN), .ZN(n6047) );
  INV_X1 U7604 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n6045) );
  NAND2_X1 U7605 ( .A1(n6046), .A2(n6045), .ZN(n6060) );
  AOI22_X1 U7606 ( .A1(n8718), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n6132), .B2(
        n7011), .ZN(n6048) );
  NAND2_X1 U7607 ( .A1(n6629), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n6056) );
  NAND2_X1 U7608 ( .A1(n6213), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n6055) );
  INV_X1 U7609 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n6050) );
  NAND2_X1 U7610 ( .A1(n6051), .A2(n6050), .ZN(n6052) );
  AND2_X1 U7611 ( .A1(n6065), .A2(n6052), .ZN(n7633) );
  NAND2_X1 U7612 ( .A1(n6223), .A2(n7633), .ZN(n6054) );
  NAND2_X1 U7613 ( .A1(n4264), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n6053) );
  NAND2_X1 U7614 ( .A1(n9358), .A2(n7698), .ZN(n8749) );
  XNOR2_X1 U7615 ( .A(n7428), .B(n7634), .ZN(n8839) );
  OR2_X1 U7616 ( .A1(n8840), .A2(n8839), .ZN(n6058) );
  NAND2_X1 U7617 ( .A1(n8749), .A2(n6057), .ZN(n8896) );
  NAND2_X1 U7618 ( .A1(n8896), .A2(n8740), .ZN(n8753) );
  NAND2_X1 U7619 ( .A1(n6058), .A2(n8753), .ZN(n8756) );
  NAND2_X1 U7620 ( .A1(n7486), .A2(n8756), .ZN(n6059) );
  NAND2_X1 U7621 ( .A1(n6730), .A2(n8714), .ZN(n6063) );
  NAND2_X1 U7622 ( .A1(n6060), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6061) );
  XNOR2_X1 U7623 ( .A(n6061), .B(P1_IR_REG_13__SCAN_IN), .ZN(n7601) );
  AOI22_X1 U7624 ( .A1(n8718), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n6132), .B2(
        n7601), .ZN(n6062) );
  NAND2_X1 U7625 ( .A1(n6213), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n6070) );
  NAND2_X1 U7626 ( .A1(n6629), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n6069) );
  NAND2_X1 U7627 ( .A1(n6065), .A2(n6064), .ZN(n6066) );
  AND2_X1 U7628 ( .A1(n6079), .A2(n6066), .ZN(n7681) );
  NAND2_X1 U7629 ( .A1(n6223), .A2(n7681), .ZN(n6068) );
  NAND2_X1 U7630 ( .A1(n4263), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n6067) );
  NAND4_X1 U7631 ( .A1(n6070), .A2(n6069), .A3(n6068), .A4(n6067), .ZN(n9009)
         );
  INV_X1 U7632 ( .A(n9009), .ZN(n8568) );
  OR2_X1 U7633 ( .A1(n7691), .A2(n8568), .ZN(n8755) );
  NAND2_X1 U7634 ( .A1(n7691), .A2(n8568), .ZN(n8752) );
  NAND2_X1 U7635 ( .A1(n7677), .A2(n8842), .ZN(n6071) );
  NAND2_X1 U7636 ( .A1(n6743), .A2(n8714), .ZN(n6078) );
  NOR2_X1 U7637 ( .A1(n6072), .A2(n9380), .ZN(n6073) );
  MUX2_X1 U7638 ( .A(n9380), .B(n6073), .S(P1_IR_REG_14__SCAN_IN), .Z(n6076)
         );
  INV_X1 U7639 ( .A(n6074), .ZN(n6075) );
  AOI22_X1 U7640 ( .A1(n8718), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n6132), .B2(
        n9554), .ZN(n6077) );
  NAND2_X1 U7641 ( .A1(n6213), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n6084) );
  NAND2_X1 U7642 ( .A1(n4264), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n6083) );
  INV_X1 U7643 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n8566) );
  NAND2_X1 U7644 ( .A1(n6079), .A2(n8566), .ZN(n6080) );
  AND2_X1 U7645 ( .A1(n6090), .A2(n6080), .ZN(n8567) );
  NAND2_X1 U7646 ( .A1(n6223), .A2(n8567), .ZN(n6082) );
  NAND2_X1 U7647 ( .A1(n6629), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n6081) );
  NAND4_X1 U7648 ( .A1(n6084), .A2(n6083), .A3(n6082), .A4(n6081), .ZN(n9008)
         );
  OR2_X1 U7649 ( .A1(n7648), .A2(n8704), .ZN(n8763) );
  NAND2_X1 U7650 ( .A1(n7648), .A2(n8704), .ZN(n8761) );
  NAND2_X1 U7651 ( .A1(n8763), .A2(n8761), .ZN(n8844) );
  NAND2_X1 U7652 ( .A1(n6074), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6086) );
  XNOR2_X1 U7653 ( .A(n6086), .B(n6085), .ZN(n7710) );
  INV_X1 U7654 ( .A(n7710), .ZN(n6087) );
  AOI22_X1 U7655 ( .A1(n8718), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n6132), .B2(
        n6087), .ZN(n6088) );
  NAND2_X1 U7656 ( .A1(n6213), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n6095) );
  NAND2_X1 U7657 ( .A1(n6629), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n6094) );
  NAND2_X1 U7658 ( .A1(n6090), .A2(n6089), .ZN(n6091) );
  AND2_X1 U7659 ( .A1(n6099), .A2(n6091), .ZN(n8703) );
  NAND2_X1 U7660 ( .A1(n6223), .A2(n8703), .ZN(n6093) );
  NAND2_X1 U7661 ( .A1(n4263), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n6092) );
  INV_X1 U7662 ( .A(n8920), .ZN(n6105) );
  OR2_X1 U7663 ( .A1(n8844), .A2(n6105), .ZN(n9253) );
  NAND2_X1 U7664 ( .A1(n6894), .A2(n8714), .ZN(n6098) );
  OR2_X1 U7665 ( .A1(n6074), .A2(P1_IR_REG_15__SCAN_IN), .ZN(n6096) );
  NAND2_X1 U7666 ( .A1(n6096), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6107) );
  XNOR2_X1 U7667 ( .A(n6107), .B(P1_IR_REG_16__SCAN_IN), .ZN(n9027) );
  AOI22_X1 U7668 ( .A1(n8718), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n6132), .B2(
        n9027), .ZN(n6097) );
  NAND2_X1 U7669 ( .A1(n6213), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n6104) );
  NAND2_X1 U7670 ( .A1(n4264), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n6103) );
  INV_X1 U7671 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n9951) );
  NAND2_X1 U7672 ( .A1(n6099), .A2(n9951), .ZN(n6100) );
  AND2_X1 U7673 ( .A1(n6114), .A2(n6100), .ZN(n9263) );
  NAND2_X1 U7674 ( .A1(n6223), .A2(n9263), .ZN(n6102) );
  NAND2_X1 U7675 ( .A1(n6629), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n6101) );
  NAND2_X1 U7676 ( .A1(n9264), .A2(n9243), .ZN(n6291) );
  INV_X1 U7677 ( .A(n6291), .ZN(n8927) );
  AND2_X1 U7678 ( .A1(n8846), .A2(n8763), .ZN(n7727) );
  NAND2_X1 U7679 ( .A1(n6970), .A2(n8714), .ZN(n6113) );
  INV_X1 U7680 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n6106) );
  NAND2_X1 U7681 ( .A1(n6107), .A2(n6106), .ZN(n6108) );
  NAND2_X1 U7682 ( .A1(n6108), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6110) );
  INV_X1 U7683 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n6109) );
  NAND2_X1 U7684 ( .A1(n6110), .A2(n6109), .ZN(n6120) );
  OR2_X1 U7685 ( .A1(n6110), .A2(n6109), .ZN(n6111) );
  AOI22_X1 U7686 ( .A1(n8718), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n6132), .B2(
        n9042), .ZN(n6112) );
  NAND2_X1 U7687 ( .A1(n6213), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n6119) );
  NAND2_X1 U7688 ( .A1(n6114), .A2(n8614), .ZN(n6115) );
  AND2_X1 U7689 ( .A1(n6125), .A2(n6115), .ZN(n8615) );
  NAND2_X1 U7690 ( .A1(n8615), .A2(n6223), .ZN(n6118) );
  NAND2_X1 U7691 ( .A1(n6629), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n6117) );
  NAND2_X1 U7692 ( .A1(n4263), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n6116) );
  NAND4_X1 U7693 ( .A1(n6119), .A2(n6118), .A3(n6117), .A4(n6116), .ZN(n9234)
         );
  INV_X1 U7694 ( .A(n9234), .ZN(n9259) );
  NOR2_X1 U7695 ( .A1(n9347), .A2(n9259), .ZN(n8772) );
  NAND2_X1 U7696 ( .A1(n9347), .A2(n9259), .ZN(n8774) );
  NAND2_X1 U7697 ( .A1(n7084), .A2(n8714), .ZN(n6123) );
  NAND2_X1 U7698 ( .A1(n6120), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6121) );
  XNOR2_X1 U7699 ( .A(n6121), .B(P1_IR_REG_18__SCAN_IN), .ZN(n9569) );
  AOI22_X1 U7700 ( .A1(n8718), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n6132), .B2(
        n9569), .ZN(n6122) );
  INV_X1 U7701 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n6124) );
  NAND2_X1 U7702 ( .A1(n6125), .A2(n6124), .ZN(n6126) );
  NAND2_X1 U7703 ( .A1(n6135), .A2(n6126), .ZN(n9224) );
  OR2_X1 U7704 ( .A1(n9224), .A2(n6212), .ZN(n6131) );
  NAND2_X1 U7705 ( .A1(n6213), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n6128) );
  NAND2_X1 U7706 ( .A1(n4264), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n6127) );
  AND2_X1 U7707 ( .A1(n6128), .A2(n6127), .ZN(n6130) );
  NAND2_X1 U7708 ( .A1(n6629), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n6129) );
  OR2_X1 U7709 ( .A1(n9339), .A2(n9244), .ZN(n8778) );
  NAND2_X1 U7710 ( .A1(n9339), .A2(n9244), .ZN(n8779) );
  NAND2_X1 U7711 ( .A1(n8778), .A2(n8779), .ZN(n9219) );
  INV_X1 U7712 ( .A(n9219), .ZN(n9230) );
  NAND2_X1 U7713 ( .A1(n9229), .A2(n9230), .ZN(n9228) );
  NAND2_X1 U7714 ( .A1(n9228), .A2(n8779), .ZN(n9212) );
  NAND2_X1 U7715 ( .A1(n7088), .A2(n8714), .ZN(n6134) );
  AOI22_X1 U7716 ( .A1(n8718), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n9248), .B2(
        n6132), .ZN(n6133) );
  NAND2_X1 U7717 ( .A1(n6135), .A2(n8584), .ZN(n6136) );
  NAND2_X1 U7718 ( .A1(n6142), .A2(n6136), .ZN(n9207) );
  AOI22_X1 U7719 ( .A1(n6629), .A2(P1_REG0_REG_19__SCAN_IN), .B1(n6213), .B2(
        P1_REG1_REG_19__SCAN_IN), .ZN(n6138) );
  NAND2_X1 U7720 ( .A1(n4263), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n6137) );
  OAI211_X1 U7721 ( .C1(n9207), .C2(n6212), .A(n6138), .B(n6137), .ZN(n9232)
         );
  INV_X1 U7722 ( .A(n9232), .ZN(n8677) );
  OR2_X1 U7723 ( .A1(n9334), .A2(n8677), .ZN(n8880) );
  NAND2_X1 U7724 ( .A1(n9334), .A2(n8677), .ZN(n8891) );
  NAND2_X1 U7725 ( .A1(n7195), .A2(n8714), .ZN(n6141) );
  NAND2_X1 U7726 ( .A1(n8718), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n6140) );
  INV_X1 U7727 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n8646) );
  NAND2_X1 U7728 ( .A1(n6142), .A2(n8646), .ZN(n6143) );
  NAND2_X1 U7729 ( .A1(n6152), .A2(n6143), .ZN(n9194) );
  OR2_X1 U7730 ( .A1(n9194), .A2(n6212), .ZN(n6149) );
  INV_X1 U7731 ( .A(P1_REG2_REG_20__SCAN_IN), .ZN(n6146) );
  NAND2_X1 U7732 ( .A1(n6629), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n6145) );
  NAND2_X1 U7733 ( .A1(n6213), .A2(P1_REG1_REG_20__SCAN_IN), .ZN(n6144) );
  OAI211_X1 U7734 ( .C1(n6146), .C2(n6226), .A(n6145), .B(n6144), .ZN(n6147)
         );
  INV_X1 U7735 ( .A(n6147), .ZN(n6148) );
  NAND2_X1 U7736 ( .A1(n6149), .A2(n6148), .ZN(n9214) );
  INV_X1 U7737 ( .A(n9214), .ZN(n8592) );
  NAND2_X1 U7738 ( .A1(n7275), .A2(n8714), .ZN(n6151) );
  NAND2_X1 U7739 ( .A1(n8718), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n6150) );
  NAND2_X1 U7740 ( .A1(n6152), .A2(n8591), .ZN(n6153) );
  NAND2_X1 U7741 ( .A1(n6163), .A2(n6153), .ZN(n9183) );
  OR2_X1 U7742 ( .A1(n9183), .A2(n6212), .ZN(n6159) );
  INV_X1 U7743 ( .A(P1_REG2_REG_21__SCAN_IN), .ZN(n6156) );
  NAND2_X1 U7744 ( .A1(n6213), .A2(P1_REG1_REG_21__SCAN_IN), .ZN(n6155) );
  NAND2_X1 U7745 ( .A1(n6629), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n6154) );
  OAI211_X1 U7746 ( .C1(n6226), .C2(n6156), .A(n6155), .B(n6154), .ZN(n6157)
         );
  INV_X1 U7747 ( .A(n6157), .ZN(n6158) );
  OR2_X1 U7748 ( .A1(n9324), .A2(n9165), .ZN(n8790) );
  NAND2_X1 U7749 ( .A1(n9324), .A2(n9165), .ZN(n8791) );
  NAND2_X1 U7750 ( .A1(n8790), .A2(n8791), .ZN(n9186) );
  NOR2_X1 U7751 ( .A1(n9186), .A2(n9176), .ZN(n6160) );
  NAND2_X1 U7752 ( .A1(n7381), .A2(n8714), .ZN(n6162) );
  NAND2_X1 U7753 ( .A1(n8718), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n6161) );
  NAND2_X1 U7754 ( .A1(n6163), .A2(n8655), .ZN(n6164) );
  NAND2_X1 U7755 ( .A1(n6175), .A2(n6164), .ZN(n8656) );
  INV_X1 U7756 ( .A(n8656), .ZN(n9170) );
  NAND2_X1 U7757 ( .A1(n9170), .A2(n6223), .ZN(n6170) );
  INV_X1 U7758 ( .A(P1_REG2_REG_22__SCAN_IN), .ZN(n6167) );
  NAND2_X1 U7759 ( .A1(n6213), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n6166) );
  NAND2_X1 U7760 ( .A1(n6629), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n6165) );
  OAI211_X1 U7761 ( .C1(n6226), .C2(n6167), .A(n6166), .B(n6165), .ZN(n6168)
         );
  INV_X1 U7762 ( .A(n6168), .ZN(n6169) );
  NAND2_X1 U7763 ( .A1(n9162), .A2(n8822), .ZN(n6171) );
  NAND2_X1 U7764 ( .A1(n9320), .A2(n9152), .ZN(n8821) );
  NAND2_X1 U7765 ( .A1(n6171), .A2(n8821), .ZN(n9151) );
  INV_X1 U7766 ( .A(n9151), .ZN(n6184) );
  NAND2_X1 U7767 ( .A1(n7571), .A2(n8714), .ZN(n6173) );
  NAND2_X1 U7768 ( .A1(n8718), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n6172) );
  INV_X1 U7769 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n6174) );
  NAND2_X1 U7770 ( .A1(n6175), .A2(n6174), .ZN(n6176) );
  NAND2_X1 U7771 ( .A1(n6188), .A2(n6176), .ZN(n9146) );
  OR2_X1 U7772 ( .A1(n9146), .A2(n6212), .ZN(n6182) );
  INV_X1 U7773 ( .A(P1_REG2_REG_23__SCAN_IN), .ZN(n6179) );
  NAND2_X1 U7774 ( .A1(n6629), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n6178) );
  NAND2_X1 U7775 ( .A1(n6213), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n6177) );
  OAI211_X1 U7776 ( .C1(n6179), .C2(n6226), .A(n6178), .B(n6177), .ZN(n6180)
         );
  INV_X1 U7777 ( .A(n6180), .ZN(n6181) );
  NAND2_X1 U7778 ( .A1(n9313), .A2(n9164), .ZN(n8973) );
  NAND2_X1 U7779 ( .A1(n8887), .A2(n8973), .ZN(n9150) );
  NAND2_X2 U7780 ( .A1(n6184), .A2(n6183), .ZN(n9155) );
  NAND2_X1 U7781 ( .A1(n7641), .A2(n8714), .ZN(n6186) );
  NAND2_X1 U7782 ( .A1(n8718), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n6185) );
  INV_X1 U7783 ( .A(n9310), .ZN(n9140) );
  INV_X1 U7784 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n6187) );
  NAND2_X1 U7785 ( .A1(n6188), .A2(n6187), .ZN(n6189) );
  NAND2_X1 U7786 ( .A1(n6199), .A2(n6189), .ZN(n8625) );
  INV_X1 U7787 ( .A(P1_REG2_REG_24__SCAN_IN), .ZN(n6192) );
  NAND2_X1 U7788 ( .A1(n6629), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n6191) );
  NAND2_X1 U7789 ( .A1(n6213), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n6190) );
  OAI211_X1 U7790 ( .C1(n6192), .C2(n6226), .A(n6191), .B(n6190), .ZN(n6193)
         );
  INV_X1 U7791 ( .A(n6193), .ZN(n6194) );
  AND2_X1 U7792 ( .A1(n9140), .A2(n9125), .ZN(n8890) );
  INV_X1 U7793 ( .A(n9125), .ZN(n9153) );
  NAND2_X1 U7794 ( .A1(n9310), .A2(n9153), .ZN(n8794) );
  NAND2_X1 U7795 ( .A1(n7722), .A2(n8714), .ZN(n6197) );
  NAND2_X1 U7796 ( .A1(n8718), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n6196) );
  NAND2_X1 U7797 ( .A1(n6199), .A2(n6198), .ZN(n6200) );
  NAND2_X1 U7798 ( .A1(n9119), .A2(n6223), .ZN(n6206) );
  INV_X1 U7799 ( .A(P1_REG2_REG_25__SCAN_IN), .ZN(n6203) );
  NAND2_X1 U7800 ( .A1(n6629), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n6202) );
  NAND2_X1 U7801 ( .A1(n6213), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n6201) );
  OAI211_X1 U7802 ( .C1(n6203), .C2(n6226), .A(n6202), .B(n6201), .ZN(n6204)
         );
  INV_X1 U7803 ( .A(n6204), .ZN(n6205) );
  OR2_X1 U7804 ( .A1(n9304), .A2(n9135), .ZN(n8873) );
  NAND2_X1 U7805 ( .A1(n9304), .A2(n9135), .ZN(n8797) );
  NAND2_X1 U7806 ( .A1(n7778), .A2(n8714), .ZN(n6208) );
  NAND2_X1 U7807 ( .A1(n8718), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n6207) );
  INV_X1 U7808 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n6209) );
  NAND2_X1 U7809 ( .A1(n6210), .A2(n6209), .ZN(n6211) );
  NAND2_X1 U7810 ( .A1(n6222), .A2(n6211), .ZN(n8689) );
  INV_X1 U7811 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n9937) );
  NAND2_X1 U7812 ( .A1(n4263), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n6215) );
  NAND2_X1 U7813 ( .A1(n6629), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n6214) );
  OAI211_X1 U7814 ( .C1(n5912), .C2(n9937), .A(n6215), .B(n6214), .ZN(n6216)
         );
  INV_X1 U7815 ( .A(n6216), .ZN(n6217) );
  XNOR2_X1 U7816 ( .A(n9300), .B(n9126), .ZN(n9105) );
  NAND2_X1 U7817 ( .A1(n9104), .A2(n9105), .ZN(n6219) );
  NAND2_X1 U7818 ( .A1(n9300), .A2(n9095), .ZN(n8867) );
  NAND2_X1 U7819 ( .A1(n7805), .A2(n8714), .ZN(n6221) );
  NAND2_X1 U7820 ( .A1(n8718), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n6220) );
  XNOR2_X1 U7821 ( .A(n6222), .B(P1_REG3_REG_27__SCAN_IN), .ZN(n9091) );
  NAND2_X1 U7822 ( .A1(n9091), .A2(n6223), .ZN(n6230) );
  INV_X1 U7823 ( .A(P1_REG2_REG_27__SCAN_IN), .ZN(n6227) );
  NAND2_X1 U7824 ( .A1(n6629), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n6225) );
  NAND2_X1 U7825 ( .A1(n6213), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n6224) );
  OAI211_X1 U7826 ( .C1(n6227), .C2(n6226), .A(n6225), .B(n6224), .ZN(n6228)
         );
  INV_X1 U7827 ( .A(n6228), .ZN(n6229) );
  NAND2_X1 U7828 ( .A1(n9293), .A2(n9107), .ZN(n8803) );
  NAND2_X1 U7829 ( .A1(n7846), .A2(n8714), .ZN(n6232) );
  NAND2_X1 U7830 ( .A1(n8718), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n6231) );
  NAND2_X1 U7831 ( .A1(n9288), .A2(n9096), .ZN(n8804) );
  NOR2_X1 U7832 ( .A1(n9072), .A2(n9071), .ZN(n9073) );
  INV_X1 U7833 ( .A(n8804), .ZN(n8807) );
  NAND2_X1 U7834 ( .A1(n8555), .A2(n8714), .ZN(n6234) );
  NAND2_X1 U7835 ( .A1(n8718), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n6233) );
  INV_X1 U7836 ( .A(n6248), .ZN(n6239) );
  INV_X1 U7837 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n6237) );
  NAND2_X1 U7838 ( .A1(n6629), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n6236) );
  NAND2_X1 U7839 ( .A1(n4264), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n6235) );
  OAI211_X1 U7840 ( .C1(n6237), .C2(n5912), .A(n6236), .B(n6235), .ZN(n6238)
         );
  AOI21_X1 U7841 ( .B1(n6239), .B2(n6223), .A(n6238), .ZN(n9075) );
  OR2_X1 U7842 ( .A1(n9284), .A2(n9075), .ZN(n8866) );
  NAND2_X1 U7843 ( .A1(n9284), .A2(n9075), .ZN(n8863) );
  NAND2_X1 U7844 ( .A1(n8866), .A2(n8863), .ZN(n8856) );
  INV_X1 U7845 ( .A(n9304), .ZN(n9121) );
  NAND2_X1 U7846 ( .A1(n7141), .A2(n7299), .ZN(n7187) );
  INV_X1 U7847 ( .A(n6382), .ZN(n9663) );
  INV_X1 U7848 ( .A(n7505), .ZN(n9395) );
  OR2_X2 U7849 ( .A1(n7489), .A2(n9358), .ZN(n7683) );
  INV_X1 U7850 ( .A(n9347), .ZN(n6244) );
  INV_X1 U7851 ( .A(n9339), .ZN(n9227) );
  INV_X1 U7852 ( .A(n9324), .ZN(n9182) );
  NAND2_X1 U7853 ( .A1(n9166), .A2(n9173), .ZN(n9167) );
  NOR2_X2 U7854 ( .A1(n9288), .A2(n9089), .ZN(n9083) );
  INV_X1 U7855 ( .A(n9083), .ZN(n6246) );
  INV_X1 U7856 ( .A(n9284), .ZN(n6245) );
  AOI211_X1 U7857 ( .C1(n9284), .C2(n6246), .A(n9664), .B(n9060), .ZN(n9283)
         );
  NAND2_X1 U7858 ( .A1(n9283), .A2(n9049), .ZN(n6247) );
  OAI211_X1 U7859 ( .C1(n6248), .C2(n9613), .A(n9286), .B(n6247), .ZN(n6265)
         );
  OR2_X1 U7860 ( .A1(n6588), .A2(n6817), .ZN(n6812) );
  NAND2_X1 U7861 ( .A1(n6264), .A2(P1_B_REG_SCAN_IN), .ZN(n6250) );
  INV_X1 U7862 ( .A(n6249), .ZN(n7642) );
  MUX2_X1 U7863 ( .A(n6250), .B(P1_B_REG_SCAN_IN), .S(n7642), .Z(n6252) );
  NAND2_X1 U7864 ( .A1(n6252), .A2(n6251), .ZN(n9614) );
  OAI22_X1 U7865 ( .A1(n9614), .A2(P1_D_REG_0__SCAN_IN), .B1(n6251), .B2(n7642), .ZN(n6550) );
  AND2_X1 U7866 ( .A1(n6550), .A2(n9649), .ZN(n9643) );
  NOR4_X1 U7867 ( .A1(P1_D_REG_14__SCAN_IN), .A2(P1_D_REG_16__SCAN_IN), .A3(
        P1_D_REG_17__SCAN_IN), .A4(P1_D_REG_18__SCAN_IN), .ZN(n6256) );
  NOR4_X1 U7868 ( .A1(P1_D_REG_11__SCAN_IN), .A2(P1_D_REG_12__SCAN_IN), .A3(
        P1_D_REG_15__SCAN_IN), .A4(P1_D_REG_13__SCAN_IN), .ZN(n6255) );
  NOR4_X1 U7869 ( .A1(P1_D_REG_24__SCAN_IN), .A2(P1_D_REG_25__SCAN_IN), .A3(
        P1_D_REG_26__SCAN_IN), .A4(P1_D_REG_27__SCAN_IN), .ZN(n6254) );
  NOR4_X1 U7870 ( .A1(P1_D_REG_19__SCAN_IN), .A2(P1_D_REG_23__SCAN_IN), .A3(
        P1_D_REG_20__SCAN_IN), .A4(P1_D_REG_21__SCAN_IN), .ZN(n6253) );
  NAND4_X1 U7871 ( .A1(n6256), .A2(n6255), .A3(n6254), .A4(n6253), .ZN(n6261)
         );
  NOR2_X1 U7872 ( .A1(P1_D_REG_28__SCAN_IN), .A2(P1_D_REG_29__SCAN_IN), .ZN(
        n9970) );
  NOR4_X1 U7873 ( .A1(P1_D_REG_30__SCAN_IN), .A2(P1_D_REG_31__SCAN_IN), .A3(
        P1_D_REG_22__SCAN_IN), .A4(P1_D_REG_7__SCAN_IN), .ZN(n6259) );
  NOR4_X1 U7874 ( .A1(P1_D_REG_6__SCAN_IN), .A2(P1_D_REG_8__SCAN_IN), .A3(
        P1_D_REG_9__SCAN_IN), .A4(P1_D_REG_10__SCAN_IN), .ZN(n6258) );
  NOR4_X1 U7875 ( .A1(P1_D_REG_2__SCAN_IN), .A2(P1_D_REG_3__SCAN_IN), .A3(
        P1_D_REG_4__SCAN_IN), .A4(P1_D_REG_5__SCAN_IN), .ZN(n6257) );
  NAND4_X1 U7876 ( .A1(n9970), .A2(n6259), .A3(n6258), .A4(n6257), .ZN(n6260)
         );
  NOR2_X1 U7877 ( .A1(n6261), .A2(n6260), .ZN(n6262) );
  NOR2_X1 U7878 ( .A1(n9614), .A2(n6262), .ZN(n6549) );
  INV_X1 U7879 ( .A(n6549), .ZN(n6263) );
  INV_X1 U7880 ( .A(n6264), .ZN(n7723) );
  OAI22_X1 U7881 ( .A1(n9614), .A2(P1_D_REG_1__SCAN_IN), .B1(n6251), .B2(n7723), .ZN(n6734) );
  INV_X1 U7882 ( .A(n6734), .ZN(n9646) );
  NAND2_X1 U7883 ( .A1(n6736), .A2(n9646), .ZN(n7188) );
  NAND2_X1 U7884 ( .A1(n6265), .A2(n9609), .ZN(n6308) );
  AND2_X1 U7885 ( .A1(n6314), .A2(n6311), .ZN(n6821) );
  NAND2_X1 U7886 ( .A1(n6822), .A2(n6821), .ZN(n6820) );
  NAND2_X1 U7887 ( .A1(n6321), .A2(n6846), .ZN(n6266) );
  NAND2_X1 U7888 ( .A1(n6820), .A2(n6266), .ZN(n6833) );
  NAND2_X1 U7889 ( .A1(n7104), .A2(n6838), .ZN(n6268) );
  NAND2_X1 U7890 ( .A1(n6992), .A2(n9650), .ZN(n6269) );
  NAND2_X1 U7891 ( .A1(n8901), .A2(n8908), .ZN(n8828) );
  NAND2_X1 U7892 ( .A1(n7103), .A2(n8636), .ZN(n6270) );
  NAND2_X1 U7893 ( .A1(n9017), .A2(n7069), .ZN(n6272) );
  NAND2_X1 U7894 ( .A1(n8903), .A2(n8733), .ZN(n8729) );
  NAND2_X1 U7895 ( .A1(n7185), .A2(n7299), .ZN(n6273) );
  NAND2_X1 U7896 ( .A1(n7134), .A2(n6273), .ZN(n7178) );
  NAND2_X1 U7897 ( .A1(n7178), .A2(n7183), .ZN(n7177) );
  NAND2_X1 U7898 ( .A1(n7307), .A2(n7192), .ZN(n6274) );
  INV_X1 U7899 ( .A(n9588), .ZN(n9014) );
  NAND2_X1 U7900 ( .A1(n7267), .A2(n9014), .ZN(n6276) );
  AND2_X1 U7901 ( .A1(n6382), .A2(n9013), .ZN(n6278) );
  OR2_X1 U7902 ( .A1(n6382), .A2(n9013), .ZN(n6277) );
  NAND2_X1 U7903 ( .A1(n7496), .A2(n8836), .ZN(n7423) );
  OR2_X1 U7904 ( .A1(n7428), .A2(n9011), .ZN(n6279) );
  INV_X1 U7905 ( .A(n9587), .ZN(n9012) );
  OR2_X1 U7906 ( .A1(n7505), .A2(n9012), .ZN(n7422) );
  AND2_X1 U7907 ( .A1(n6279), .A2(n7422), .ZN(n6280) );
  NAND2_X1 U7908 ( .A1(n7423), .A2(n6280), .ZN(n7673) );
  NAND2_X1 U7909 ( .A1(n7428), .A2(n9011), .ZN(n7484) );
  INV_X1 U7910 ( .A(n7698), .ZN(n9010) );
  NAND2_X1 U7911 ( .A1(n9358), .A2(n9010), .ZN(n6283) );
  AND2_X1 U7912 ( .A1(n7484), .A2(n6283), .ZN(n7672) );
  INV_X1 U7913 ( .A(n6285), .ZN(n6281) );
  AND2_X1 U7914 ( .A1(n7672), .A2(n6281), .ZN(n6282) );
  INV_X1 U7915 ( .A(n6283), .ZN(n6284) );
  NOR2_X1 U7916 ( .A1(n7648), .A2(n9008), .ZN(n6287) );
  NAND2_X1 U7917 ( .A1(n6288), .A2(n9260), .ZN(n6290) );
  OR2_X1 U7918 ( .A1(n7725), .A2(n8695), .ZN(n6289) );
  NAND2_X1 U7919 ( .A1(n6290), .A2(n6289), .ZN(n9270) );
  INV_X1 U7920 ( .A(n9243), .ZN(n9006) );
  NAND2_X1 U7921 ( .A1(n9264), .A2(n9006), .ZN(n6292) );
  OR2_X1 U7922 ( .A1(n9347), .A2(n9234), .ZN(n6293) );
  NAND2_X1 U7923 ( .A1(n9220), .A2(n9219), .ZN(n6295) );
  INV_X1 U7924 ( .A(n9244), .ZN(n9213) );
  NAND2_X1 U7925 ( .A1(n9339), .A2(n9213), .ZN(n6294) );
  OR2_X1 U7926 ( .A1(n9334), .A2(n9232), .ZN(n6297) );
  AND2_X1 U7927 ( .A1(n9334), .A2(n9232), .ZN(n6296) );
  NAND2_X1 U7928 ( .A1(n9173), .A2(n9152), .ZN(n6299) );
  INV_X1 U7929 ( .A(n9164), .ZN(n9005) );
  NOR2_X1 U7930 ( .A1(n9310), .A2(n9125), .ZN(n8851) );
  INV_X1 U7931 ( .A(n9300), .ZN(n9112) );
  INV_X1 U7932 ( .A(n9107), .ZN(n9003) );
  OAI22_X1 U7933 ( .A1(n9088), .A2(n8853), .B1(n9003), .B2(n9293), .ZN(n9068)
         );
  XOR2_X1 U7934 ( .A(n8856), .B(n6303), .Z(n9287) );
  AND2_X2 U7935 ( .A1(n6304), .A2(n8987), .ZN(n7090) );
  OR2_X1 U7936 ( .A1(n6816), .A2(n6305), .ZN(n6562) );
  NAND2_X4 U7937 ( .A1(n6816), .A2(n6305), .ZN(n6520) );
  NOR2_X1 U7938 ( .A1(n7094), .A2(n8987), .ZN(n6845) );
  AOI22_X1 U7939 ( .A1(n9284), .A2(n9605), .B1(P1_REG2_REG_29__SCAN_IN), .B2(
        n9597), .ZN(n6306) );
  NAND2_X1 U7940 ( .A1(n6308), .A2(n4824), .ZN(P1_U3355) );
  INV_X2 U7941 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3084) );
  OR2_X4 U7942 ( .A1(n6586), .A2(n7090), .ZN(n6500) );
  AND2_X1 U7943 ( .A1(n6309), .A2(n6817), .ZN(n6310) );
  NOR2_X4 U7944 ( .A1(n6500), .A2(n6310), .ZN(n6541) );
  AOI22_X1 U7945 ( .A1(n6311), .A2(n6320), .B1(P1_IR_REG_0__SCAN_IN), .B2(
        n6586), .ZN(n6312) );
  INV_X1 U7946 ( .A(n6312), .ZN(n6313) );
  AOI21_X1 U7947 ( .B1(n6314), .B2(n6541), .A(n6313), .ZN(n6804) );
  NAND2_X1 U7948 ( .A1(n6314), .A2(n6320), .ZN(n6317) );
  AND2_X1 U7949 ( .A1(n6586), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n6315) );
  NAND2_X1 U7950 ( .A1(n6317), .A2(n6316), .ZN(n6802) );
  NAND2_X1 U7951 ( .A1(n6804), .A2(n6802), .ZN(n6803) );
  INV_X1 U7952 ( .A(n6520), .ZN(n6318) );
  OR2_X1 U7953 ( .A1(n6802), .A2(n6318), .ZN(n6319) );
  INV_X1 U7954 ( .A(n6328), .ZN(n6326) );
  INV_X2 U7955 ( .A(n6320), .ZN(n6522) );
  NAND2_X1 U7956 ( .A1(n6321), .A2(n6377), .ZN(n6323) );
  NAND2_X1 U7957 ( .A1(n6846), .A2(n6370), .ZN(n6322) );
  NAND2_X1 U7958 ( .A1(n6323), .A2(n6322), .ZN(n6324) );
  XNOR2_X1 U7959 ( .A(n6324), .B(n6318), .ZN(n6327) );
  INV_X1 U7960 ( .A(n6327), .ZN(n6325) );
  NAND2_X1 U7961 ( .A1(n6321), .A2(n6541), .ZN(n6330) );
  NAND2_X1 U7962 ( .A1(n6846), .A2(n6377), .ZN(n6329) );
  NAND2_X1 U7963 ( .A1(n6330), .A2(n6329), .ZN(n6750) );
  NAND2_X1 U7964 ( .A1(n6747), .A2(n6332), .ZN(n8661) );
  OAI22_X1 U7965 ( .A1(n7104), .A2(n6522), .B1(n6838), .B2(n6500), .ZN(n6333)
         );
  XNOR2_X1 U7966 ( .A(n6333), .B(n6544), .ZN(n6338) );
  OR2_X1 U7967 ( .A1(n7104), .A2(n6536), .ZN(n6335) );
  NAND2_X1 U7968 ( .A1(n8666), .A2(n6377), .ZN(n6334) );
  INV_X1 U7969 ( .A(n6336), .ZN(n6337) );
  NAND2_X1 U7970 ( .A1(n6338), .A2(n6337), .ZN(n6339) );
  XNOR2_X1 U7971 ( .A(n6340), .B(n6544), .ZN(n6343) );
  OR2_X1 U7972 ( .A1(n6992), .A2(n6536), .ZN(n6342) );
  NAND2_X1 U7973 ( .A1(n7100), .A2(n6377), .ZN(n6341) );
  AND2_X1 U7974 ( .A1(n6342), .A2(n6341), .ZN(n6344) );
  INV_X1 U7975 ( .A(n6343), .ZN(n6346) );
  INV_X1 U7976 ( .A(n6344), .ZN(n6345) );
  NAND2_X1 U7977 ( .A1(n6346), .A2(n6345), .ZN(n8630) );
  OAI22_X1 U7978 ( .A1(n7103), .A2(n6522), .B1(n8636), .B2(n6500), .ZN(n6347)
         );
  XNOR2_X1 U7979 ( .A(n6347), .B(n6544), .ZN(n6353) );
  OR2_X1 U7980 ( .A1(n7103), .A2(n6536), .ZN(n6349) );
  NAND2_X1 U7981 ( .A1(n6996), .A2(n6377), .ZN(n6348) );
  NAND2_X1 U7982 ( .A1(n6349), .A2(n6348), .ZN(n6351) );
  XNOR2_X1 U7983 ( .A(n6353), .B(n6351), .ZN(n8634) );
  AND2_X1 U7984 ( .A1(n8630), .A2(n8634), .ZN(n6350) );
  INV_X1 U7985 ( .A(n6351), .ZN(n6352) );
  NAND2_X1 U7986 ( .A1(n6353), .A2(n6352), .ZN(n6354) );
  OR2_X1 U7987 ( .A1(n7294), .A2(n6536), .ZN(n6356) );
  NAND2_X1 U7988 ( .A1(n7069), .A2(n6377), .ZN(n6355) );
  NAND2_X1 U7989 ( .A1(n6356), .A2(n6355), .ZN(n7127) );
  OAI22_X1 U7990 ( .A1(n7294), .A2(n6522), .B1(n9657), .B2(n6500), .ZN(n6357)
         );
  XNOR2_X1 U7991 ( .A(n6357), .B(n6520), .ZN(n6362) );
  OAI22_X1 U7992 ( .A1(n7185), .A2(n6522), .B1(n7299), .B2(n6500), .ZN(n6358)
         );
  XNOR2_X1 U7993 ( .A(n6358), .B(n6520), .ZN(n7288) );
  OR2_X1 U7994 ( .A1(n7185), .A2(n6536), .ZN(n6360) );
  NAND2_X1 U7995 ( .A1(n7143), .A2(n6377), .ZN(n6359) );
  NAND2_X1 U7996 ( .A1(n6360), .A2(n6359), .ZN(n7287) );
  AOI22_X1 U7997 ( .A1(n7127), .A2(n6362), .B1(n7288), .B2(n7287), .ZN(n6361)
         );
  NAND2_X1 U7998 ( .A1(n7285), .A2(n6361), .ZN(n6367) );
  OAI21_X1 U7999 ( .B1(n6362), .B2(n7127), .A(n7287), .ZN(n6365) );
  INV_X1 U8000 ( .A(n7288), .ZN(n6364) );
  INV_X1 U8001 ( .A(n6362), .ZN(n7286) );
  NOR2_X1 U8002 ( .A1(n7127), .A2(n7287), .ZN(n6363) );
  AOI22_X1 U8003 ( .A1(n6365), .A2(n6364), .B1(n7286), .B2(n6363), .ZN(n6366)
         );
  OR2_X1 U8004 ( .A1(n7307), .A2(n6536), .ZN(n6369) );
  NAND2_X1 U8005 ( .A1(n7221), .A2(n6377), .ZN(n6368) );
  AND2_X1 U8006 ( .A1(n6369), .A2(n6368), .ZN(n7075) );
  NAND2_X1 U8007 ( .A1(n7221), .A2(n6370), .ZN(n6371) );
  OAI21_X1 U8008 ( .B1(n7307), .B2(n6522), .A(n6371), .ZN(n6372) );
  XNOR2_X1 U8009 ( .A(n6372), .B(n6544), .ZN(n6383) );
  NAND2_X1 U8010 ( .A1(n6386), .A2(n6383), .ZN(n6376) );
  NAND2_X1 U8011 ( .A1(n7078), .A2(n7075), .ZN(n6384) );
  NAND2_X1 U8012 ( .A1(n7267), .A2(n6377), .ZN(n6374) );
  OR2_X1 U8013 ( .A1(n9588), .A2(n6536), .ZN(n6373) );
  NAND2_X1 U8014 ( .A1(n6374), .A2(n6373), .ZN(n6385) );
  AND2_X1 U8015 ( .A1(n6384), .A2(n6385), .ZN(n6375) );
  NAND2_X1 U8016 ( .A1(n6382), .A2(n6370), .ZN(n6379) );
  NAND2_X1 U8017 ( .A1(n9013), .A2(n6377), .ZN(n6378) );
  NAND2_X1 U8018 ( .A1(n6379), .A2(n6378), .ZN(n6380) );
  XNOR2_X1 U8019 ( .A(n6380), .B(n6520), .ZN(n6392) );
  AND2_X1 U8020 ( .A1(n9013), .A2(n6541), .ZN(n6381) );
  AOI21_X1 U8021 ( .B1(n6382), .B2(n6510), .A(n6381), .ZN(n6393) );
  XNOR2_X1 U8022 ( .A(n6392), .B(n6393), .ZN(n7368) );
  INV_X1 U8023 ( .A(n6383), .ZN(n7076) );
  NAND2_X1 U8024 ( .A1(n6384), .A2(n7076), .ZN(n6388) );
  INV_X1 U8025 ( .A(n6385), .ZN(n6387) );
  NAND3_X1 U8026 ( .A1(n6388), .A2(n6387), .A3(n6386), .ZN(n7301) );
  NAND2_X1 U8027 ( .A1(n7267), .A2(n6370), .ZN(n6390) );
  OR2_X1 U8028 ( .A1(n9588), .A2(n6522), .ZN(n6389) );
  NAND2_X1 U8029 ( .A1(n6390), .A2(n6389), .ZN(n6391) );
  XNOR2_X1 U8030 ( .A(n6391), .B(n6520), .ZN(n7300) );
  NAND2_X1 U8031 ( .A1(n7301), .A2(n7300), .ZN(n7370) );
  INV_X1 U8032 ( .A(n6392), .ZN(n6394) );
  NAND2_X1 U8033 ( .A1(n6394), .A2(n6393), .ZN(n6395) );
  NAND2_X1 U8034 ( .A1(n7505), .A2(n6370), .ZN(n6397) );
  OR2_X1 U8035 ( .A1(n9587), .A2(n6522), .ZN(n6396) );
  NAND2_X1 U8036 ( .A1(n6397), .A2(n6396), .ZN(n6398) );
  XNOR2_X1 U8037 ( .A(n6398), .B(n6520), .ZN(n6401) );
  NAND2_X1 U8038 ( .A1(n7505), .A2(n6538), .ZN(n6400) );
  OR2_X1 U8039 ( .A1(n9587), .A2(n6536), .ZN(n6399) );
  NAND2_X1 U8040 ( .A1(n6400), .A2(n6399), .ZN(n6402) );
  NAND2_X1 U8041 ( .A1(n6401), .A2(n6402), .ZN(n7384) );
  INV_X1 U8042 ( .A(n6401), .ZN(n6404) );
  INV_X1 U8043 ( .A(n6402), .ZN(n6403) );
  NAND2_X1 U8044 ( .A1(n6404), .A2(n6403), .ZN(n7383) );
  NAND2_X1 U8045 ( .A1(n7428), .A2(n6370), .ZN(n6406) );
  NAND2_X1 U8046 ( .A1(n9011), .A2(n6538), .ZN(n6405) );
  NAND2_X1 U8047 ( .A1(n6406), .A2(n6405), .ZN(n6407) );
  XNOR2_X1 U8048 ( .A(n6407), .B(n6544), .ZN(n6410) );
  AND2_X1 U8049 ( .A1(n9011), .A2(n6541), .ZN(n6408) );
  AOI21_X1 U8050 ( .B1(n7428), .B2(n6510), .A(n6408), .ZN(n6411) );
  XNOR2_X1 U8051 ( .A(n6410), .B(n6411), .ZN(n7542) );
  INV_X1 U8052 ( .A(n7542), .ZN(n6409) );
  INV_X1 U8053 ( .A(n6410), .ZN(n6413) );
  INV_X1 U8054 ( .A(n6411), .ZN(n6412) );
  NAND2_X1 U8055 ( .A1(n6413), .A2(n6412), .ZN(n6414) );
  NAND2_X1 U8056 ( .A1(n9358), .A2(n6370), .ZN(n6416) );
  OR2_X1 U8057 ( .A1(n7698), .A2(n6522), .ZN(n6415) );
  NAND2_X1 U8058 ( .A1(n6416), .A2(n6415), .ZN(n6417) );
  XNOR2_X1 U8059 ( .A(n6417), .B(n6544), .ZN(n7630) );
  NOR2_X1 U8060 ( .A1(n7698), .A2(n6536), .ZN(n6418) );
  AOI21_X1 U8061 ( .B1(n9358), .B2(n6538), .A(n6418), .ZN(n6420) );
  NAND2_X1 U8062 ( .A1(n7630), .A2(n6420), .ZN(n6419) );
  INV_X1 U8063 ( .A(n7630), .ZN(n6421) );
  INV_X1 U8064 ( .A(n6420), .ZN(n7629) );
  NAND2_X1 U8065 ( .A1(n6421), .A2(n7629), .ZN(n6422) );
  NAND2_X1 U8066 ( .A1(n7691), .A2(n6370), .ZN(n6424) );
  NAND2_X1 U8067 ( .A1(n9009), .A2(n6538), .ZN(n6423) );
  NAND2_X1 U8068 ( .A1(n6424), .A2(n6423), .ZN(n6425) );
  XNOR2_X1 U8069 ( .A(n6425), .B(n6520), .ZN(n6428) );
  NAND2_X1 U8070 ( .A1(n7691), .A2(n6538), .ZN(n6427) );
  NAND2_X1 U8071 ( .A1(n9009), .A2(n6541), .ZN(n6426) );
  NAND2_X1 U8072 ( .A1(n6427), .A2(n6426), .ZN(n6429) );
  AND2_X1 U8073 ( .A1(n6428), .A2(n6429), .ZN(n7693) );
  INV_X1 U8074 ( .A(n6428), .ZN(n6431) );
  INV_X1 U8075 ( .A(n6429), .ZN(n6430) );
  NAND2_X1 U8076 ( .A1(n7648), .A2(n6370), .ZN(n6433) );
  NAND2_X1 U8077 ( .A1(n9008), .A2(n6538), .ZN(n6432) );
  NAND2_X1 U8078 ( .A1(n6433), .A2(n6432), .ZN(n6434) );
  NAND2_X1 U8079 ( .A1(n7648), .A2(n6538), .ZN(n6436) );
  NAND2_X1 U8080 ( .A1(n9008), .A2(n6541), .ZN(n6435) );
  NAND2_X1 U8081 ( .A1(n6436), .A2(n6435), .ZN(n8563) );
  NAND2_X1 U8082 ( .A1(n8561), .A2(n8563), .ZN(n6444) );
  INV_X1 U8083 ( .A(n6437), .ZN(n6438) );
  NAND2_X1 U8084 ( .A1(n6438), .A2(n4293), .ZN(n8562) );
  NAND2_X1 U8085 ( .A1(n8695), .A2(n6370), .ZN(n6440) );
  OR2_X1 U8086 ( .A1(n9260), .A2(n6522), .ZN(n6439) );
  NAND2_X1 U8087 ( .A1(n6440), .A2(n6439), .ZN(n6441) );
  XNOR2_X1 U8088 ( .A(n6441), .B(n6544), .ZN(n6445) );
  NAND3_X1 U8089 ( .A1(n6444), .A2(n8562), .A3(n6445), .ZN(n8697) );
  NAND2_X1 U8090 ( .A1(n8695), .A2(n6538), .ZN(n6443) );
  OR2_X1 U8091 ( .A1(n9260), .A2(n6536), .ZN(n6442) );
  NAND2_X1 U8092 ( .A1(n6443), .A2(n6442), .ZN(n8698) );
  NAND2_X1 U8093 ( .A1(n6444), .A2(n8562), .ZN(n6447) );
  INV_X1 U8094 ( .A(n6445), .ZN(n6446) );
  NAND2_X1 U8095 ( .A1(n9264), .A2(n6370), .ZN(n6449) );
  OR2_X1 U8096 ( .A1(n9243), .A2(n6522), .ZN(n6448) );
  NAND2_X1 U8097 ( .A1(n6449), .A2(n6448), .ZN(n6450) );
  XNOR2_X1 U8098 ( .A(n6450), .B(n6520), .ZN(n6452) );
  NOR2_X1 U8099 ( .A1(n9243), .A2(n6536), .ZN(n6451) );
  AOI21_X1 U8100 ( .B1(n9264), .B2(n6510), .A(n6451), .ZN(n6453) );
  XNOR2_X1 U8101 ( .A(n6452), .B(n6453), .ZN(n8606) );
  INV_X1 U8102 ( .A(n6452), .ZN(n6454) );
  NAND2_X1 U8103 ( .A1(n6454), .A2(n6453), .ZN(n6455) );
  NAND2_X1 U8104 ( .A1(n9347), .A2(n6370), .ZN(n6457) );
  NAND2_X1 U8105 ( .A1(n9234), .A2(n6538), .ZN(n6456) );
  NAND2_X1 U8106 ( .A1(n6457), .A2(n6456), .ZN(n6458) );
  XNOR2_X1 U8107 ( .A(n6458), .B(n6520), .ZN(n6460) );
  AND2_X1 U8108 ( .A1(n9234), .A2(n6541), .ZN(n6459) );
  AOI21_X1 U8109 ( .B1(n9347), .B2(n6538), .A(n6459), .ZN(n6461) );
  XNOR2_X1 U8110 ( .A(n6460), .B(n6461), .ZN(n8612) );
  INV_X1 U8111 ( .A(n6460), .ZN(n6462) );
  NAND2_X1 U8112 ( .A1(n6462), .A2(n6461), .ZN(n6463) );
  NAND2_X1 U8113 ( .A1(n6464), .A2(n6463), .ZN(n8675) );
  NAND2_X1 U8114 ( .A1(n9339), .A2(n6370), .ZN(n6466) );
  NAND2_X1 U8115 ( .A1(n9213), .A2(n6538), .ZN(n6465) );
  NAND2_X1 U8116 ( .A1(n6466), .A2(n6465), .ZN(n6467) );
  XNOR2_X1 U8117 ( .A(n6467), .B(n6544), .ZN(n8673) );
  NOR2_X1 U8118 ( .A1(n9244), .A2(n6536), .ZN(n6468) );
  AOI21_X1 U8119 ( .B1(n9339), .B2(n6510), .A(n6468), .ZN(n8672) );
  NAND2_X1 U8120 ( .A1(n9334), .A2(n6370), .ZN(n6470) );
  NAND2_X1 U8121 ( .A1(n9232), .A2(n6538), .ZN(n6469) );
  NAND2_X1 U8122 ( .A1(n6470), .A2(n6469), .ZN(n6471) );
  XNOR2_X1 U8123 ( .A(n6471), .B(n6520), .ZN(n6473) );
  AND2_X1 U8124 ( .A1(n9232), .A2(n6541), .ZN(n6472) );
  AOI21_X1 U8125 ( .B1(n9334), .B2(n6538), .A(n6472), .ZN(n6474) );
  XNOR2_X1 U8126 ( .A(n6473), .B(n6474), .ZN(n8582) );
  INV_X1 U8127 ( .A(n6473), .ZN(n6475) );
  NAND2_X1 U8128 ( .A1(n9329), .A2(n6370), .ZN(n6477) );
  NAND2_X1 U8129 ( .A1(n9214), .A2(n6538), .ZN(n6476) );
  NAND2_X1 U8130 ( .A1(n6477), .A2(n6476), .ZN(n6478) );
  XNOR2_X1 U8131 ( .A(n6478), .B(n6520), .ZN(n6481) );
  NAND2_X1 U8132 ( .A1(n9329), .A2(n6538), .ZN(n6480) );
  NAND2_X1 U8133 ( .A1(n9214), .A2(n6541), .ZN(n6479) );
  NAND2_X1 U8134 ( .A1(n6480), .A2(n6479), .ZN(n6482) );
  NAND2_X1 U8135 ( .A1(n6481), .A2(n6482), .ZN(n8643) );
  INV_X1 U8136 ( .A(n6481), .ZN(n6484) );
  INV_X1 U8137 ( .A(n6482), .ZN(n6483) );
  NAND2_X1 U8138 ( .A1(n6484), .A2(n6483), .ZN(n8644) );
  NAND2_X1 U8139 ( .A1(n9324), .A2(n6370), .ZN(n6486) );
  INV_X1 U8140 ( .A(n9165), .ZN(n9199) );
  NAND2_X1 U8141 ( .A1(n9199), .A2(n6538), .ZN(n6485) );
  NAND2_X1 U8142 ( .A1(n6486), .A2(n6485), .ZN(n6487) );
  XNOR2_X1 U8143 ( .A(n6487), .B(n6520), .ZN(n6489) );
  NOR2_X1 U8144 ( .A1(n9165), .A2(n6536), .ZN(n6488) );
  AOI21_X1 U8145 ( .B1(n9324), .B2(n6510), .A(n6488), .ZN(n6490) );
  XNOR2_X1 U8146 ( .A(n6489), .B(n6490), .ZN(n8589) );
  INV_X1 U8147 ( .A(n6489), .ZN(n6491) );
  NAND2_X1 U8148 ( .A1(n6491), .A2(n6490), .ZN(n6492) );
  OR2_X1 U8149 ( .A1(n9173), .A2(n6522), .ZN(n6494) );
  NAND2_X1 U8150 ( .A1(n9179), .A2(n6541), .ZN(n6493) );
  AND2_X1 U8151 ( .A1(n6494), .A2(n6493), .ZN(n6497) );
  NAND2_X1 U8152 ( .A1(n6496), .A2(n6497), .ZN(n8651) );
  OAI22_X1 U8153 ( .A1(n9173), .A2(n6500), .B1(n9152), .B2(n6522), .ZN(n6495)
         );
  XNOR2_X1 U8154 ( .A(n6495), .B(n6520), .ZN(n8654) );
  INV_X1 U8155 ( .A(n6496), .ZN(n6499) );
  INV_X1 U8156 ( .A(n6497), .ZN(n6498) );
  OAI22_X1 U8157 ( .A1(n9149), .A2(n6500), .B1(n9164), .B2(n6522), .ZN(n6501)
         );
  XNOR2_X1 U8158 ( .A(n6501), .B(n6520), .ZN(n6504) );
  OR2_X1 U8159 ( .A1(n9149), .A2(n6522), .ZN(n6503) );
  NAND2_X1 U8160 ( .A1(n9005), .A2(n6541), .ZN(n6502) );
  AND2_X1 U8161 ( .A1(n6503), .A2(n6502), .ZN(n8575) );
  INV_X1 U8162 ( .A(n6504), .ZN(n6505) );
  NAND2_X1 U8163 ( .A1(n9310), .A2(n6370), .ZN(n6507) );
  NAND2_X1 U8164 ( .A1(n9125), .A2(n6538), .ZN(n6506) );
  NAND2_X1 U8165 ( .A1(n6507), .A2(n6506), .ZN(n6508) );
  XNOR2_X1 U8166 ( .A(n6508), .B(n6544), .ZN(n6511) );
  AND2_X1 U8167 ( .A1(n9125), .A2(n6541), .ZN(n6509) );
  AOI21_X1 U8168 ( .B1(n9310), .B2(n6510), .A(n6509), .ZN(n6512) );
  NAND2_X1 U8169 ( .A1(n6511), .A2(n6512), .ZN(n6516) );
  INV_X1 U8170 ( .A(n6511), .ZN(n6514) );
  INV_X1 U8171 ( .A(n6512), .ZN(n6513) );
  NAND2_X1 U8172 ( .A1(n6514), .A2(n6513), .ZN(n6515) );
  NAND2_X1 U8173 ( .A1(n6516), .A2(n6515), .ZN(n8620) );
  INV_X1 U8174 ( .A(n6516), .ZN(n6517) );
  NAND2_X1 U8175 ( .A1(n9304), .A2(n6370), .ZN(n6519) );
  NAND2_X1 U8176 ( .A1(n9004), .A2(n6538), .ZN(n6518) );
  NAND2_X1 U8177 ( .A1(n6519), .A2(n6518), .ZN(n6521) );
  XNOR2_X1 U8178 ( .A(n6521), .B(n6520), .ZN(n6524) );
  OAI22_X1 U8179 ( .A1(n9121), .A2(n6522), .B1(n9135), .B2(n6536), .ZN(n6523)
         );
  XNOR2_X1 U8180 ( .A(n6524), .B(n6523), .ZN(n8597) );
  NOR2_X1 U8181 ( .A1(n6524), .A2(n6523), .ZN(n8685) );
  NAND2_X1 U8182 ( .A1(n9300), .A2(n6370), .ZN(n6526) );
  NAND2_X1 U8183 ( .A1(n9126), .A2(n6538), .ZN(n6525) );
  NAND2_X1 U8184 ( .A1(n6526), .A2(n6525), .ZN(n6527) );
  XNOR2_X1 U8185 ( .A(n6527), .B(n6544), .ZN(n6529) );
  AND2_X1 U8186 ( .A1(n9126), .A2(n6541), .ZN(n6528) );
  AOI21_X1 U8187 ( .B1(n9300), .B2(n6538), .A(n6528), .ZN(n6530) );
  XNOR2_X1 U8188 ( .A(n6529), .B(n6530), .ZN(n8684) );
  INV_X1 U8189 ( .A(n6529), .ZN(n6532) );
  INV_X1 U8190 ( .A(n6530), .ZN(n6531) );
  NAND2_X1 U8191 ( .A1(n9293), .A2(n6370), .ZN(n6534) );
  OR2_X1 U8192 ( .A1(n9107), .A2(n6522), .ZN(n6533) );
  NAND2_X1 U8193 ( .A1(n6534), .A2(n6533), .ZN(n6535) );
  XNOR2_X1 U8194 ( .A(n6535), .B(n6544), .ZN(n6540) );
  NOR2_X1 U8195 ( .A1(n9107), .A2(n6536), .ZN(n6537) );
  AOI21_X1 U8196 ( .B1(n9293), .B2(n6538), .A(n6537), .ZN(n6539) );
  NAND2_X1 U8197 ( .A1(n6540), .A2(n6539), .ZN(n6567) );
  OAI21_X1 U8198 ( .B1(n6540), .B2(n6539), .A(n6567), .ZN(n6576) );
  NOR3_X4 U8199 ( .A1(n6574), .A2(n6575), .A3(n6576), .ZN(n6580) );
  NAND2_X1 U8200 ( .A1(n9288), .A2(n6538), .ZN(n6543) );
  NAND2_X1 U8201 ( .A1(n9002), .A2(n6541), .ZN(n6542) );
  NAND2_X1 U8202 ( .A1(n6543), .A2(n6542), .ZN(n6545) );
  XNOR2_X1 U8203 ( .A(n6545), .B(n6544), .ZN(n6548) );
  NAND2_X1 U8204 ( .A1(n9288), .A2(n6370), .ZN(n6546) );
  OAI21_X1 U8205 ( .B1(n9096), .B2(n6522), .A(n6546), .ZN(n6547) );
  XNOR2_X1 U8206 ( .A(n6548), .B(n6547), .ZN(n6552) );
  INV_X1 U8207 ( .A(n6552), .ZN(n6568) );
  NOR2_X1 U8208 ( .A1(n6550), .A2(n6549), .ZN(n6813) );
  NAND2_X1 U8209 ( .A1(n6813), .A2(n9646), .ZN(n6751) );
  OR2_X1 U8210 ( .A1(n6751), .A2(n9645), .ZN(n6556) );
  INV_X1 U8211 ( .A(n7094), .ZN(n6737) );
  OR2_X1 U8212 ( .A1(n9359), .A2(n8815), .ZN(n6560) );
  NAND3_X1 U8213 ( .A1(n6568), .A2(n8700), .A3(n6567), .ZN(n6551) );
  INV_X1 U8214 ( .A(n6845), .ZN(n6554) );
  OR2_X1 U8215 ( .A1(n6556), .A2(n6554), .ZN(n6555) );
  NOR2_X1 U8216 ( .A1(n6556), .A2(n6562), .ZN(n6557) );
  NAND2_X1 U8217 ( .A1(n6557), .A2(n5909), .ZN(n8676) );
  INV_X1 U8218 ( .A(n8705), .ZN(n8668) );
  NAND2_X1 U8219 ( .A1(n9003), .A2(n8668), .ZN(n6566) );
  INV_X1 U8220 ( .A(n6751), .ZN(n6559) );
  AND3_X1 U8221 ( .A1(n6812), .A2(n6587), .A3(n7572), .ZN(n6558) );
  OAI21_X1 U8222 ( .B1(n6560), .B2(n6559), .A(n6558), .ZN(n6561) );
  NAND2_X1 U8223 ( .A1(n6561), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6564) );
  INV_X1 U8224 ( .A(n6562), .ZN(n8994) );
  OR2_X1 U8225 ( .A1(n8994), .A2(n6845), .ZN(n6563) );
  NAND3_X1 U8226 ( .A1(n6563), .A2(n9649), .A3(n6751), .ZN(n6753) );
  NAND2_X1 U8227 ( .A1(n6564), .A2(n6753), .ZN(n8690) );
  AOI22_X1 U8228 ( .A1(n9078), .A2(n8690), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3084), .ZN(n6565) );
  OAI211_X1 U8229 ( .C1(n9075), .C2(n8676), .A(n6566), .B(n6565), .ZN(n6570)
         );
  NOR3_X1 U8230 ( .A1(n6568), .A2(n8682), .A3(n6567), .ZN(n6569) );
  AOI211_X1 U8231 ( .C1(n9288), .C2(n8680), .A(n6570), .B(n6569), .ZN(n6571)
         );
  NAND3_X1 U8232 ( .A1(n6573), .A2(n6572), .A3(n6571), .ZN(P1_U3218) );
  INV_X1 U8233 ( .A(n6575), .ZN(n6578) );
  INV_X1 U8234 ( .A(n6576), .ZN(n6577) );
  AOI21_X1 U8235 ( .B1(n8688), .B2(n6578), .A(n6577), .ZN(n6579) );
  OAI21_X1 U8236 ( .B1(n6580), .B2(n6579), .A(n8700), .ZN(n6585) );
  OAI22_X1 U8237 ( .A1(n9095), .A2(n8705), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n6581), .ZN(n6583) );
  NOR2_X1 U8238 ( .A1(n9096), .A2(n8676), .ZN(n6582) );
  AOI211_X1 U8239 ( .C1(n9091), .C2(n8690), .A(n6583), .B(n6582), .ZN(n6584)
         );
  INV_X1 U8240 ( .A(n8680), .ZN(n8713) );
  NAND3_X1 U8241 ( .A1(n6585), .A2(n6584), .A3(n4815), .ZN(P1_U3212) );
  NAND2_X1 U8242 ( .A1(n6588), .A2(n6587), .ZN(n6589) );
  NAND2_X1 U8243 ( .A1(n6589), .A2(n7572), .ZN(n6646) );
  NAND2_X1 U8244 ( .A1(n6646), .A2(n6590), .ZN(n6666) );
  NAND2_X1 U8245 ( .A1(n6666), .A2(P1_STATE_REG_SCAN_IN), .ZN(P1_U3083) );
  INV_X1 U8246 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n6591) );
  INV_X1 U8247 ( .A(n6650), .ZN(n6797) );
  OAI222_X1 U8248 ( .A1(n7085), .A2(n6591), .B1(n6951), .B2(n6599), .C1(
        P1_U3084), .C2(n6797), .ZN(P1_U3351) );
  INV_X1 U8249 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n6592) );
  OAI222_X1 U8250 ( .A1(n7085), .A2(n6592), .B1(n6951), .B2(n6603), .C1(
        P1_U3084), .C2(n4648), .ZN(P1_U3352) );
  CLKBUF_X1 U8251 ( .A(n9383), .Z(n9389) );
  AOI22_X1 U8252 ( .A1(P2_DATAO_REG_4__SCAN_IN), .A2(n9389), .B1(n9470), .B2(
        P1_STATE_REG_SCAN_IN), .ZN(n6593) );
  OAI21_X1 U8253 ( .B1(n6601), .B2(n6951), .A(n6593), .ZN(P1_U3349) );
  AOI22_X1 U8254 ( .A1(n9478), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_5__SCAN_IN), .B2(n9389), .ZN(n6594) );
  OAI21_X1 U8255 ( .B1(n6606), .B2(n6951), .A(n6594), .ZN(P1_U3348) );
  AOI22_X1 U8256 ( .A1(n6719), .A2(P1_STATE_REG_SCAN_IN), .B1(n9389), .B2(
        P2_DATAO_REG_3__SCAN_IN), .ZN(n6595) );
  OAI21_X1 U8257 ( .B1(n6605), .B2(n6951), .A(n6595), .ZN(P1_U3350) );
  INV_X1 U8258 ( .A(n8008), .ZN(n8017) );
  INV_X1 U8259 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n6598) );
  INV_X1 U8260 ( .A(n8556), .ZN(n8051) );
  OAI222_X1 U8261 ( .A1(P2_U3152), .A2(n8017), .B1(n8049), .B2(n6599), .C1(
        n6598), .C2(n8051), .ZN(P2_U3356) );
  INV_X1 U8262 ( .A(n7982), .ZN(n7989) );
  OAI222_X1 U8263 ( .A1(P2_U3152), .A2(n7989), .B1(n8049), .B2(n6601), .C1(
        n6600), .C2(n8051), .ZN(P2_U3354) );
  INV_X1 U8264 ( .A(n7340), .ZN(n7324) );
  INV_X1 U8265 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n6602) );
  OAI222_X1 U8266 ( .A1(P2_U3152), .A2(n7324), .B1(n8049), .B2(n6603), .C1(
        n6602), .C2(n8051), .ZN(P2_U3357) );
  INV_X1 U8267 ( .A(n7342), .ZN(n8001) );
  OAI222_X1 U8268 ( .A1(P2_U3152), .A2(n8001), .B1(n8049), .B2(n6605), .C1(
        n6604), .C2(n8051), .ZN(P2_U3355) );
  OAI222_X1 U8269 ( .A1(n8051), .A2(n6607), .B1(n8049), .B2(n6606), .C1(
        P2_U3152), .C2(n4280), .ZN(P2_U3353) );
  INV_X1 U8270 ( .A(n6608), .ZN(n6610) );
  AOI22_X1 U8271 ( .A1(n9490), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_6__SCAN_IN), .B2(n9389), .ZN(n6609) );
  OAI21_X1 U8272 ( .B1(n6610), .B2(n6951), .A(n6609), .ZN(P1_U3347) );
  INV_X1 U8273 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n9902) );
  INV_X1 U8274 ( .A(n7347), .ZN(n7964) );
  OAI222_X1 U8275 ( .A1(n8051), .A2(n9902), .B1(n8049), .B2(n6610), .C1(
        P2_U3152), .C2(n7964), .ZN(P2_U3352) );
  INV_X1 U8276 ( .A(n6611), .ZN(n6616) );
  AOI22_X1 U8277 ( .A1(n9498), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_7__SCAN_IN), .B2(n9389), .ZN(n6612) );
  OAI21_X1 U8278 ( .B1(n6616), .B2(n6951), .A(n6612), .ZN(P1_U3346) );
  INV_X1 U8279 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n6614) );
  NAND2_X1 U8280 ( .A1(n6779), .A2(P2_U3966), .ZN(n6613) );
  OAI21_X1 U8281 ( .B1(n6614), .B2(P2_U3966), .A(n6613), .ZN(P2_U3552) );
  AOI22_X1 U8282 ( .A1(n9516), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(n9383), .ZN(n6615) );
  OAI21_X1 U8283 ( .B1(n6619), .B2(n6951), .A(n6615), .ZN(P1_U3345) );
  INV_X1 U8284 ( .A(n7349), .ZN(n7952) );
  OAI222_X1 U8285 ( .A1(n8051), .A2(n9965), .B1(n8049), .B2(n6616), .C1(
        P2_U3152), .C2(n7952), .ZN(P2_U3351) );
  OAI21_X1 U8286 ( .B1(n9707), .B2(n6772), .A(n4885), .ZN(n6618) );
  NAND2_X1 U8287 ( .A1(n9707), .A2(n7575), .ZN(n6617) );
  NAND2_X1 U8288 ( .A1(n6618), .A2(n6617), .ZN(n8033) );
  INV_X1 U8289 ( .A(n8033), .ZN(n9681) );
  NOR2_X1 U8290 ( .A1(n9681), .A2(P2_U3966), .ZN(P2_U3151) );
  INV_X1 U8291 ( .A(n7351), .ZN(n7941) );
  OAI222_X1 U8292 ( .A1(n8051), .A2(n6620), .B1(n8049), .B2(n6619), .C1(
        P2_U3152), .C2(n7941), .ZN(P2_U3350) );
  INV_X1 U8293 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n9859) );
  NAND2_X1 U8294 ( .A1(n8264), .A2(P2_U3966), .ZN(n6621) );
  OAI21_X1 U8295 ( .B1(n9859), .B2(P2_U3966), .A(n6621), .ZN(P2_U3583) );
  INV_X1 U8296 ( .A(n6622), .ZN(n6624) );
  AOI22_X1 U8297 ( .A1(n9528), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_9__SCAN_IN), .B2(n9383), .ZN(n6623) );
  OAI21_X1 U8298 ( .B1(n6624), .B2(n6951), .A(n6623), .ZN(P1_U3344) );
  OAI222_X1 U8299 ( .A1(n8051), .A2(n6625), .B1(n8049), .B2(n6624), .C1(n7930), 
        .C2(P2_U3152), .ZN(P2_U3349) );
  INV_X1 U8300 ( .A(n6626), .ZN(n6636) );
  AOI22_X1 U8301 ( .A1(n6942), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n9383), .ZN(n6627) );
  OAI21_X1 U8302 ( .B1(n6636), .B2(n6951), .A(n6627), .ZN(P1_U3343) );
  INV_X1 U8303 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n6634) );
  NAND2_X1 U8304 ( .A1(n6213), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n6632) );
  NAND2_X1 U8305 ( .A1(n4263), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n6631) );
  NAND2_X1 U8306 ( .A1(n6629), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n6630) );
  NAND3_X1 U8307 ( .A1(n6632), .A2(n6631), .A3(n6630), .ZN(n9055) );
  NAND2_X1 U8308 ( .A1(n9055), .A2(P1_U4006), .ZN(n6633) );
  OAI21_X1 U8309 ( .B1(P1_U4006), .B2(n6634), .A(n6633), .ZN(P1_U3586) );
  INV_X1 U8310 ( .A(n7355), .ZN(n7918) );
  OAI222_X1 U8311 ( .A1(P2_U3152), .A2(n7918), .B1(n8049), .B2(n6636), .C1(
        n6635), .C2(n8051), .ZN(P2_U3348) );
  INV_X1 U8312 ( .A(n6637), .ZN(n6639) );
  INV_X1 U8313 ( .A(n9536), .ZN(n6940) );
  OAI222_X1 U8314 ( .A1(n7085), .A2(n6638), .B1(n6951), .B2(n6639), .C1(n6940), 
        .C2(P1_U3084), .ZN(P1_U3342) );
  INV_X1 U8315 ( .A(n7357), .ZN(n7907) );
  OAI222_X1 U8316 ( .A1(n8051), .A2(n6640), .B1(n8049), .B2(n6639), .C1(n7907), 
        .C2(P2_U3152), .ZN(P2_U3347) );
  INV_X1 U8317 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n6660) );
  NOR2_X1 U8318 ( .A1(n6805), .A2(P1_U3084), .ZN(n7806) );
  AND2_X1 U8319 ( .A1(n7806), .A2(n5909), .ZN(n6642) );
  NAND2_X1 U8320 ( .A1(n6646), .A2(n6642), .ZN(n9045) );
  AND2_X1 U8321 ( .A1(P1_U3084), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n6860) );
  INV_X1 U8322 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n6904) );
  MUX2_X1 U8323 ( .A(P1_REG1_REG_2__SCAN_IN), .B(n6904), .S(n6650), .Z(n6792)
         );
  INV_X1 U8324 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n6829) );
  MUX2_X1 U8325 ( .A(P1_REG1_REG_1__SCAN_IN), .B(n6829), .S(n6651), .Z(n6675)
         );
  NAND2_X1 U8326 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), 
        .ZN(n6679) );
  INV_X1 U8327 ( .A(n6679), .ZN(n6643) );
  NAND2_X1 U8328 ( .A1(n6675), .A2(n6643), .ZN(n6676) );
  NAND2_X1 U8329 ( .A1(n6651), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n6644) );
  NAND2_X1 U8330 ( .A1(n6676), .A2(n6644), .ZN(n6791) );
  INV_X1 U8331 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n6645) );
  MUX2_X1 U8332 ( .A(n6645), .B(P1_REG1_REG_3__SCAN_IN), .S(n6719), .Z(n6647)
         );
  NOR2_X1 U8333 ( .A1(n4298), .A2(n6647), .ZN(n6708) );
  NOR2_X1 U8334 ( .A1(n5909), .A2(P1_U3084), .ZN(n7847) );
  NAND2_X1 U8335 ( .A1(n6646), .A2(n7847), .ZN(n6654) );
  AOI211_X1 U8336 ( .C1(n4298), .C2(n6647), .A(n6708), .B(n9510), .ZN(n6648)
         );
  AOI211_X1 U8337 ( .C1(n4360), .C2(n6719), .A(n6860), .B(n6648), .ZN(n6659)
         );
  INV_X1 U8338 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n6649) );
  MUX2_X1 U8339 ( .A(P1_REG2_REG_3__SCAN_IN), .B(n6649), .S(n6719), .Z(n6657)
         );
  INV_X1 U8340 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n6653) );
  MUX2_X1 U8341 ( .A(P1_REG2_REG_2__SCAN_IN), .B(n6653), .S(n6650), .Z(n6795)
         );
  INV_X1 U8342 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n6855) );
  AND2_X1 U8343 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(
        n6807) );
  NAND2_X1 U8344 ( .A1(n6651), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n6652) );
  NAND2_X1 U8345 ( .A1(n6671), .A2(n6652), .ZN(n6794) );
  NAND2_X1 U8346 ( .A1(n6795), .A2(n6794), .ZN(n6793) );
  OAI21_X1 U8347 ( .B1(n6653), .B2(n6797), .A(n6793), .ZN(n6656) );
  INV_X1 U8348 ( .A(n6654), .ZN(n6655) );
  OAI211_X1 U8349 ( .C1(n6657), .C2(n6656), .A(n9543), .B(n4561), .ZN(n6658)
         );
  OAI211_X1 U8350 ( .C1(n6660), .C2(n9561), .A(n6659), .B(n6658), .ZN(P1_U3244) );
  INV_X1 U8351 ( .A(n9561), .ZN(n9573) );
  INV_X1 U8352 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n9612) );
  NAND3_X1 U8353 ( .A1(n9574), .A2(P1_IR_REG_0__SCAN_IN), .A3(n5911), .ZN(
        n6668) );
  OR2_X1 U8354 ( .A1(n6805), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n6661) );
  AOI21_X1 U8355 ( .B1(n8993), .B2(n6661), .A(P1_IR_REG_0__SCAN_IN), .ZN(n6808) );
  AOI21_X1 U8356 ( .B1(P1_IR_REG_0__SCAN_IN), .B2(P1_REG2_REG_0__SCAN_IN), .A(
        n6805), .ZN(n6664) );
  NOR2_X1 U8357 ( .A1(n5911), .A2(P1_IR_REG_0__SCAN_IN), .ZN(n6662) );
  OR2_X1 U8358 ( .A1(n5909), .A2(n6662), .ZN(n6663) );
  OAI21_X1 U8359 ( .B1(n6664), .B2(n6663), .A(P1_STATE_REG_SCAN_IN), .ZN(n6665) );
  OR3_X1 U8360 ( .A1(n6666), .A2(n6808), .A3(n6665), .ZN(n6667) );
  OAI211_X1 U8361 ( .C1(P1_STATE_REG_SCAN_IN), .C2(n9612), .A(n6668), .B(n6667), .ZN(n6669) );
  AOI21_X1 U8362 ( .B1(n9573), .B2(P1_ADDR_REG_0__SCAN_IN), .A(n6669), .ZN(
        n6670) );
  INV_X1 U8363 ( .A(n6670), .ZN(P1_U3241) );
  OAI211_X1 U8364 ( .C1(n6672), .C2(n6807), .A(n9543), .B(n6671), .ZN(n6674)
         );
  NAND2_X1 U8365 ( .A1(P1_U3084), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n6673) );
  OAI211_X1 U8366 ( .C1(n9045), .C2(n4648), .A(n6674), .B(n6673), .ZN(n6681)
         );
  INV_X1 U8367 ( .A(n6675), .ZN(n6678) );
  INV_X1 U8368 ( .A(n6676), .ZN(n6677) );
  AOI211_X1 U8369 ( .C1(n6679), .C2(n6678), .A(n6677), .B(n9510), .ZN(n6680)
         );
  AOI211_X1 U8370 ( .C1(P1_ADDR_REG_1__SCAN_IN), .C2(n9573), .A(n6681), .B(
        n6680), .ZN(n6682) );
  INV_X1 U8371 ( .A(n6682), .ZN(P1_U3242) );
  INV_X1 U8372 ( .A(n6683), .ZN(n6685) );
  INV_X1 U8373 ( .A(n7450), .ZN(n7314) );
  OAI222_X1 U8374 ( .A1(n8051), .A2(n6684), .B1(n8049), .B2(n6685), .C1(
        P2_U3152), .C2(n7314), .ZN(P2_U3346) );
  INV_X1 U8375 ( .A(n7011), .ZN(n6939) );
  OAI222_X1 U8376 ( .A1(n7085), .A2(n6686), .B1(n6951), .B2(n6685), .C1(
        P1_U3084), .C2(n6939), .ZN(P1_U3341) );
  NAND2_X1 U8377 ( .A1(n4885), .A2(n6772), .ZN(n6691) );
  NAND2_X1 U8378 ( .A1(n6687), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6688) );
  NAND2_X1 U8379 ( .A1(n6688), .A2(n7575), .ZN(n6689) );
  NAND2_X1 U8380 ( .A1(n6689), .A2(n7849), .ZN(n6690) );
  OAI21_X1 U8381 ( .B1(n9707), .B2(n6691), .A(n6690), .ZN(n6694) );
  OR2_X1 U8382 ( .A1(n6694), .A2(P2_U3966), .ZN(n6700) );
  NOR2_X1 U8383 ( .A1(n5828), .A2(n7575), .ZN(n6692) );
  OAI21_X2 U8384 ( .B1(n6700), .B2(n6692), .A(n5560), .ZN(n8030) );
  INV_X1 U8385 ( .A(n8030), .ZN(n9684) );
  INV_X1 U8386 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n9815) );
  INV_X1 U8387 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n9907) );
  OAI22_X1 U8388 ( .A1(n8033), .A2(n9815), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9907), .ZN(n6698) );
  NAND2_X1 U8389 ( .A1(n9689), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n6696) );
  INV_X1 U8390 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n6693) );
  AOI211_X1 U8391 ( .C1(n6696), .C2(n6695), .A(n7339), .B(n9682), .ZN(n6697)
         );
  AOI211_X1 U8392 ( .C1(n9684), .C2(n7340), .A(n6698), .B(n6697), .ZN(n6704)
         );
  AND2_X1 U8393 ( .A1(n9689), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n6702) );
  INV_X1 U8394 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n6699) );
  MUX2_X1 U8395 ( .A(P2_REG2_REG_1__SCAN_IN), .B(n6699), .S(n7340), .Z(n6701)
         );
  INV_X1 U8396 ( .A(n5828), .ZN(n8072) );
  NAND2_X1 U8397 ( .A1(n8028), .A2(n7849), .ZN(n8027) );
  INV_X1 U8398 ( .A(n8027), .ZN(n9680) );
  NAND3_X1 U8399 ( .A1(n6701), .A2(P2_REG2_REG_0__SCAN_IN), .A3(n9689), .ZN(
        n8011) );
  OAI211_X1 U8400 ( .C1(n6702), .C2(n6701), .A(n9680), .B(n8011), .ZN(n6703)
         );
  NAND2_X1 U8401 ( .A1(n6704), .A2(n6703), .ZN(P2_U3246) );
  INV_X1 U8402 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n6729) );
  NAND2_X1 U8403 ( .A1(n9516), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n6705) );
  OAI21_X1 U8404 ( .B1(n9516), .B2(P1_REG1_REG_8__SCAN_IN), .A(n6705), .ZN(
        n9512) );
  NOR2_X1 U8405 ( .A1(P1_REG1_REG_7__SCAN_IN), .A2(n9498), .ZN(n6706) );
  AOI21_X1 U8406 ( .B1(n9498), .B2(P1_REG1_REG_7__SCAN_IN), .A(n6706), .ZN(
        n9501) );
  NAND2_X1 U8407 ( .A1(P1_REG1_REG_5__SCAN_IN), .A2(n9478), .ZN(n6707) );
  OAI21_X1 U8408 ( .B1(n9478), .B2(P1_REG1_REG_5__SCAN_IN), .A(n6707), .ZN(
        n9474) );
  NOR2_X1 U8409 ( .A1(n9470), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n6709) );
  AOI21_X1 U8410 ( .B1(n9470), .B2(P1_REG1_REG_4__SCAN_IN), .A(n6709), .ZN(
        n9463) );
  NAND2_X1 U8411 ( .A1(n9462), .A2(n9463), .ZN(n9461) );
  OAI21_X1 U8412 ( .B1(n9470), .B2(P1_REG1_REG_4__SCAN_IN), .A(n9461), .ZN(
        n9475) );
  NOR2_X1 U8413 ( .A1(n9474), .A2(n9475), .ZN(n9473) );
  NOR2_X1 U8414 ( .A1(n9490), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n6710) );
  AOI21_X1 U8415 ( .B1(P1_REG1_REG_6__SCAN_IN), .B2(n9490), .A(n6710), .ZN(
        n9492) );
  NAND2_X1 U8416 ( .A1(n9493), .A2(n9492), .ZN(n9491) );
  OAI21_X1 U8417 ( .B1(n9490), .B2(P1_REG1_REG_6__SCAN_IN), .A(n9491), .ZN(
        n9500) );
  NAND2_X1 U8418 ( .A1(n9501), .A2(n9500), .ZN(n9499) );
  OAI21_X1 U8419 ( .B1(P1_REG1_REG_7__SCAN_IN), .B2(n9498), .A(n9499), .ZN(
        n9513) );
  NOR2_X1 U8420 ( .A1(n9512), .A2(n9513), .ZN(n9511) );
  NOR2_X1 U8421 ( .A1(n9528), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n6711) );
  AOI21_X1 U8422 ( .B1(P1_REG1_REG_9__SCAN_IN), .B2(n9528), .A(n6711), .ZN(
        n9531) );
  NAND2_X1 U8423 ( .A1(n9530), .A2(n9531), .ZN(n9529) );
  OAI21_X1 U8424 ( .B1(P1_REG1_REG_9__SCAN_IN), .B2(n9528), .A(n9529), .ZN(
        n6714) );
  INV_X1 U8425 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n6712) );
  MUX2_X1 U8426 ( .A(P1_REG1_REG_10__SCAN_IN), .B(n6712), .S(n6942), .Z(n6713)
         );
  NAND2_X1 U8427 ( .A1(n6713), .A2(n6714), .ZN(n6935) );
  OAI21_X1 U8428 ( .B1(n6714), .B2(n6713), .A(n6935), .ZN(n6715) );
  NAND2_X1 U8429 ( .A1(n6715), .A2(n9574), .ZN(n6728) );
  AND2_X1 U8430 ( .A1(P1_U3084), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n7389) );
  NOR2_X1 U8431 ( .A1(n9516), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n6716) );
  AOI21_X1 U8432 ( .B1(P1_REG2_REG_8__SCAN_IN), .B2(n9516), .A(n6716), .ZN(
        n9519) );
  NOR2_X1 U8433 ( .A1(P1_REG2_REG_7__SCAN_IN), .A2(n9498), .ZN(n6717) );
  AOI21_X1 U8434 ( .B1(n9498), .B2(P1_REG2_REG_7__SCAN_IN), .A(n6717), .ZN(
        n9504) );
  NOR2_X1 U8435 ( .A1(P1_REG2_REG_5__SCAN_IN), .A2(n9478), .ZN(n6718) );
  AOI21_X1 U8436 ( .B1(n9478), .B2(P1_REG2_REG_5__SCAN_IN), .A(n6718), .ZN(
        n9480) );
  NOR2_X1 U8437 ( .A1(n9470), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n6720) );
  AOI21_X1 U8438 ( .B1(n9470), .B2(P1_REG2_REG_4__SCAN_IN), .A(n6720), .ZN(
        n9465) );
  NAND2_X1 U8439 ( .A1(n9480), .A2(n9481), .ZN(n9479) );
  OAI21_X1 U8440 ( .B1(P1_REG2_REG_5__SCAN_IN), .B2(n9478), .A(n9479), .ZN(
        n9487) );
  NAND2_X1 U8441 ( .A1(n9490), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n6721) );
  OAI21_X1 U8442 ( .B1(n9490), .B2(P1_REG2_REG_6__SCAN_IN), .A(n6721), .ZN(
        n9486) );
  NOR2_X1 U8443 ( .A1(n9487), .A2(n9486), .ZN(n9485) );
  OAI21_X1 U8444 ( .B1(P1_REG2_REG_8__SCAN_IN), .B2(n9516), .A(n9517), .ZN(
        n9525) );
  NAND2_X1 U8445 ( .A1(n9528), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n6722) );
  OAI21_X1 U8446 ( .B1(n9528), .B2(P1_REG2_REG_9__SCAN_IN), .A(n6722), .ZN(
        n9524) );
  INV_X1 U8447 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n6723) );
  MUX2_X1 U8448 ( .A(n6723), .B(P1_REG2_REG_10__SCAN_IN), .S(n6942), .Z(n6724)
         );
  AOI211_X1 U8449 ( .C1(n6725), .C2(n6724), .A(n6941), .B(n9563), .ZN(n6726)
         );
  AOI211_X1 U8450 ( .C1(n4360), .C2(n6942), .A(n7389), .B(n6726), .ZN(n6727)
         );
  OAI211_X1 U8451 ( .C1(n9561), .C2(n6729), .A(n6728), .B(n6727), .ZN(P1_U3251) );
  INV_X1 U8452 ( .A(n6730), .ZN(n6732) );
  INV_X1 U8453 ( .A(n7475), .ZN(n7448) );
  OAI222_X1 U8454 ( .A1(n8051), .A2(n6731), .B1(n8049), .B2(n6732), .C1(n7448), 
        .C2(P2_U3152), .ZN(P2_U3345) );
  INV_X1 U8455 ( .A(n7601), .ZN(n7009) );
  OAI222_X1 U8456 ( .A1(n7085), .A2(n6733), .B1(n6951), .B2(n6732), .C1(n7009), 
        .C2(P1_U3084), .ZN(P1_U3340) );
  AND2_X1 U8457 ( .A1(n6735), .A2(n6734), .ZN(n6815) );
  INV_X1 U8458 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n6742) );
  AND2_X1 U8459 ( .A1(n6314), .A2(n6825), .ZN(n8948) );
  NOR2_X1 U8460 ( .A1(n6823), .A2(n8948), .ZN(n8827) );
  OR3_X1 U8461 ( .A1(n8827), .A2(n6737), .A3(n8994), .ZN(n6739) );
  NAND2_X1 U8462 ( .A1(n6321), .A2(n9231), .ZN(n6738) );
  NAND2_X1 U8463 ( .A1(n6739), .A2(n6738), .ZN(n9603) );
  INV_X1 U8464 ( .A(n9603), .ZN(n6740) );
  OAI21_X1 U8465 ( .B1(n6825), .B2(n7094), .A(n6740), .ZN(n6872) );
  NAND2_X1 U8466 ( .A1(n6872), .A2(n9672), .ZN(n6741) );
  OAI21_X1 U8467 ( .B1(n9672), .B2(n6742), .A(n6741), .ZN(P1_U3454) );
  INV_X1 U8468 ( .A(n6743), .ZN(n6744) );
  INV_X1 U8469 ( .A(n7768), .ZN(n7473) );
  OAI222_X1 U8470 ( .A1(n8051), .A2(n9887), .B1(n8049), .B2(n6744), .C1(n7473), 
        .C2(P2_U3152), .ZN(P2_U3344) );
  OAI222_X1 U8471 ( .A1(n7085), .A2(n6745), .B1(n6951), .B2(n6744), .C1(n7599), 
        .C2(P1_U3084), .ZN(P1_U3339) );
  INV_X1 U8472 ( .A(n6748), .ZN(n6749) );
  AOI21_X1 U8473 ( .B1(n6750), .B2(n6746), .A(n6749), .ZN(n6756) );
  INV_X1 U8474 ( .A(n9359), .ZN(n9662) );
  NAND2_X1 U8475 ( .A1(n9662), .A2(n6751), .ZN(n6752) );
  NAND4_X1 U8476 ( .A1(n6753), .A2(n9649), .A3(n6812), .A4(n6752), .ZN(n8667)
         );
  AOI22_X1 U8477 ( .A1(n8667), .A2(P1_REG3_REG_1__SCAN_IN), .B1(n8680), .B2(
        n6846), .ZN(n6755) );
  AOI22_X1 U8478 ( .A1(n8668), .A2(n6314), .B1(n8710), .B2(n9020), .ZN(n6754)
         );
  OAI211_X1 U8479 ( .C1(n6756), .C2(n8682), .A(n6755), .B(n6754), .ZN(P1_U3220) );
  INV_X2 U8480 ( .A(P2_U3966), .ZN(n8248) );
  NAND2_X1 U8481 ( .A1(P2_DATAO_REG_29__SCAN_IN), .A2(n8248), .ZN(n6757) );
  OAI21_X1 U8482 ( .B1(n6758), .B2(n8248), .A(n6757), .ZN(P2_U3581) );
  AND2_X1 U8483 ( .A1(n6762), .A2(n6761), .ZN(n6765) );
  INV_X1 U8484 ( .A(n6763), .ZN(n6764) );
  NAND2_X1 U8485 ( .A1(n5575), .A2(n7045), .ZN(n6767) );
  NAND2_X1 U8486 ( .A1(n6767), .A2(n9727), .ZN(n6768) );
  NOR2_X1 U8487 ( .A1(n7119), .A2(n6768), .ZN(n7459) );
  OR2_X1 U8488 ( .A1(n6770), .A2(n6769), .ZN(n6771) );
  NAND2_X1 U8489 ( .A1(n6874), .A2(n6771), .ZN(n7463) );
  NAND2_X1 U8490 ( .A1(n7028), .A2(n7419), .ZN(n6774) );
  AND2_X1 U8491 ( .A1(n5645), .A2(n6772), .ZN(n6773) );
  NOR2_X1 U8492 ( .A1(n7463), .A2(n9731), .ZN(n6775) );
  AOI211_X1 U8493 ( .C1(n9726), .C2(n5575), .A(n7459), .B(n6775), .ZN(n6783)
         );
  XNOR2_X1 U8494 ( .A(n6769), .B(n6776), .ZN(n6782) );
  OR2_X1 U8495 ( .A1(n5576), .A2(n9756), .ZN(n6781) );
  NAND2_X1 U8496 ( .A1(n6779), .A2(n8443), .ZN(n6780) );
  NAND2_X1 U8497 ( .A1(n6781), .A2(n6780), .ZN(n8045) );
  AOI21_X1 U8498 ( .B1(n6782), .B2(n9693), .A(n8045), .ZN(n7467) );
  NAND2_X1 U8499 ( .A1(n6783), .A2(n7467), .ZN(n6787) );
  NAND2_X1 U8500 ( .A1(n6787), .A2(n9810), .ZN(n6784) );
  OAI21_X1 U8501 ( .B1(n9810), .B2(n6693), .A(n6784), .ZN(P2_U3521) );
  INV_X1 U8502 ( .A(n7025), .ZN(n6785) );
  INV_X1 U8503 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n6789) );
  NAND2_X1 U8504 ( .A1(n6787), .A2(n9796), .ZN(n6788) );
  OAI21_X1 U8505 ( .B1(n9796), .B2(n6789), .A(n6788), .ZN(P2_U3454) );
  OAI21_X1 U8506 ( .B1(n6792), .B2(n6791), .A(n6790), .ZN(n6801) );
  OAI211_X1 U8507 ( .C1(n6795), .C2(n6794), .A(n9543), .B(n6793), .ZN(n6800)
         );
  INV_X1 U8508 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n6796) );
  OAI22_X1 U8509 ( .A1(n9045), .A2(n6797), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n6796), .ZN(n6798) );
  INV_X1 U8510 ( .A(n6798), .ZN(n6799) );
  OAI211_X1 U8511 ( .C1(n6801), .C2(n9510), .A(n6800), .B(n6799), .ZN(n6810)
         );
  OAI21_X1 U8512 ( .B1(n6804), .B2(n6802), .A(n6803), .ZN(n8036) );
  INV_X1 U8513 ( .A(n8036), .ZN(n6806) );
  MUX2_X1 U8514 ( .A(n6807), .B(n6806), .S(n6805), .Z(n6809) );
  INV_X2 U8515 ( .A(P1_U4006), .ZN(n9021) );
  AOI211_X1 U8516 ( .C1(n6809), .C2(n8993), .A(n6808), .B(n9021), .ZN(n9468)
         );
  AOI211_X1 U8517 ( .C1(n9573), .C2(P1_ADDR_REG_2__SCAN_IN), .A(n6810), .B(
        n9468), .ZN(n6811) );
  INV_X1 U8518 ( .A(n6811), .ZN(P1_U3243) );
  OR2_X1 U8519 ( .A1(n6816), .A2(n7090), .ZN(n6819) );
  NAND3_X1 U8520 ( .A1(n8816), .A2(n8951), .A3(n6817), .ZN(n6818) );
  OAI21_X1 U8521 ( .B1(n6822), .B2(n6821), .A(n6820), .ZN(n6849) );
  XNOR2_X1 U8522 ( .A(n8824), .B(n6823), .ZN(n6824) );
  AOI222_X1 U8523 ( .A1(n9590), .A2(n6824), .B1(n9020), .B2(n9231), .C1(n6314), 
        .C2(n9233), .ZN(n6848) );
  OAI21_X1 U8524 ( .B1(n8949), .B2(n6825), .A(n9340), .ZN(n6826) );
  NOR2_X1 U8525 ( .A1(n6826), .A2(n6836), .ZN(n6852) );
  AOI21_X1 U8526 ( .B1(n9359), .B2(n6846), .A(n6852), .ZN(n6827) );
  OAI211_X1 U8527 ( .C1(n9426), .C2(n6849), .A(n6848), .B(n6827), .ZN(n6830)
         );
  NAND2_X1 U8528 ( .A1(n6830), .A2(n9440), .ZN(n6828) );
  OAI21_X1 U8529 ( .B1(n9362), .B2(n6829), .A(n6828), .ZN(P1_U3524) );
  INV_X1 U8530 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n6832) );
  NAND2_X1 U8531 ( .A1(n6830), .A2(n9672), .ZN(n6831) );
  OAI21_X1 U8532 ( .B1(n9672), .B2(n6832), .A(n6831), .ZN(P1_U3457) );
  NAND2_X1 U8533 ( .A1(n6833), .A2(n8825), .ZN(n6834) );
  NAND2_X1 U8534 ( .A1(n6835), .A2(n6834), .ZN(n7853) );
  OR2_X1 U8535 ( .A1(n6836), .A2(n6838), .ZN(n6837) );
  NAND2_X1 U8536 ( .A1(n7096), .A2(n6837), .ZN(n7856) );
  OAI22_X1 U8537 ( .A1(n7856), .A2(n9664), .B1(n6838), .B2(n9662), .ZN(n6842)
         );
  XNOR2_X1 U8538 ( .A(n6267), .B(n8956), .ZN(n6841) );
  INV_X1 U8539 ( .A(n9593), .ZN(n7726) );
  NAND2_X1 U8540 ( .A1(n7853), .A2(n7726), .ZN(n6840) );
  AOI22_X1 U8541 ( .A1(n9019), .A2(n9231), .B1(n9233), .B2(n6321), .ZN(n6839)
         );
  OAI211_X1 U8542 ( .C1(n6841), .C2(n6240), .A(n6840), .B(n6839), .ZN(n7852)
         );
  AOI211_X1 U8543 ( .C1(n9669), .C2(n7853), .A(n6842), .B(n7852), .ZN(n6902)
         );
  NAND2_X1 U8544 ( .A1(n9670), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n6843) );
  OAI21_X1 U8545 ( .B1(n6902), .B2(n9670), .A(n6843), .ZN(P1_U3460) );
  INV_X1 U8546 ( .A(n6844), .ZN(n6850) );
  AOI22_X1 U8547 ( .A1(n9595), .A2(P1_REG3_REG_1__SCAN_IN), .B1(n6846), .B2(
        n6845), .ZN(n6847) );
  OAI211_X1 U8548 ( .C1(n6850), .C2(n6849), .A(n6848), .B(n6847), .ZN(n6851)
         );
  NAND2_X1 U8549 ( .A1(n6851), .A2(n9609), .ZN(n6854) );
  AND2_X1 U8550 ( .A1(n9609), .A2(n9049), .ZN(n9169) );
  NAND2_X1 U8551 ( .A1(n9169), .A2(n6852), .ZN(n6853) );
  OAI211_X1 U8552 ( .C1(n6855), .C2(n9609), .A(n6854), .B(n6853), .ZN(P1_U3290) );
  NAND2_X1 U8553 ( .A1(n6856), .A2(n8630), .ZN(n6857) );
  XNOR2_X1 U8554 ( .A(n6858), .B(n6857), .ZN(n6863) );
  AOI22_X1 U8555 ( .A1(n8668), .A2(n9020), .B1(n8710), .B2(n9018), .ZN(n6862)
         );
  NOR2_X1 U8556 ( .A1(n8713), .A2(n9650), .ZN(n6859) );
  AOI211_X1 U8557 ( .C1(n7099), .C2(n8690), .A(n6860), .B(n6859), .ZN(n6861)
         );
  OAI211_X1 U8558 ( .C1(n6863), .C2(n8682), .A(n6862), .B(n6861), .ZN(P1_U3216) );
  NAND2_X1 U8559 ( .A1(n7027), .A2(n6865), .ZN(n8044) );
  AOI22_X1 U8560 ( .A1(n6864), .A2(n8195), .B1(n8044), .B2(
        P2_REG3_REG_0__SCAN_IN), .ZN(n6871) );
  OAI21_X1 U8561 ( .B1(n6867), .B2(n6866), .A(n4505), .ZN(n6869) );
  NAND3_X1 U8562 ( .A1(n6869), .A2(n6868), .A3(n8214), .ZN(n6870) );
  OAI211_X1 U8563 ( .C1(n8227), .C2(n4505), .A(n6871), .B(n6870), .ZN(P2_U3234) );
  NAND2_X1 U8564 ( .A1(n6872), .A2(n9440), .ZN(n6873) );
  OAI21_X1 U8565 ( .B1(n9440), .B2(n5911), .A(n6873), .ZN(P1_U3523) );
  INV_X1 U8566 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n6890) );
  NAND2_X1 U8567 ( .A1(n5576), .A2(n6875), .ZN(n6876) );
  NAND2_X1 U8568 ( .A1(n6877), .A2(n6876), .ZN(n6953) );
  NAND2_X1 U8569 ( .A1(n6953), .A2(n6956), .ZN(n6952) );
  NAND2_X1 U8570 ( .A1(n7116), .A2(n7397), .ZN(n6878) );
  NAND2_X1 U8571 ( .A1(n6952), .A2(n6878), .ZN(n7022) );
  NAND2_X1 U8572 ( .A1(n7022), .A2(n7021), .ZN(n7020) );
  NAND2_X1 U8573 ( .A1(n6954), .A2(n7039), .ZN(n6879) );
  NAND2_X1 U8574 ( .A1(n7020), .A2(n6879), .ZN(n6880) );
  OAI21_X1 U8575 ( .B1(n6880), .B2(n6884), .A(n6906), .ZN(n6881) );
  INV_X1 U8576 ( .A(n6881), .ZN(n7057) );
  NAND2_X1 U8577 ( .A1(n6883), .A2(n6882), .ZN(n6885) );
  XNOR2_X1 U8578 ( .A(n6885), .B(n6884), .ZN(n6886) );
  OAI22_X1 U8579 ( .A1(n6954), .A2(n9758), .B1(n8084), .B2(n9756), .ZN(n6985)
         );
  AOI21_X1 U8580 ( .B1(n6886), .B2(n9693), .A(n6985), .ZN(n7049) );
  INV_X1 U8581 ( .A(n7033), .ZN(n6887) );
  AOI211_X1 U8582 ( .C1(n6986), .C2(n6887), .A(n9780), .B(n6916), .ZN(n7054)
         );
  AOI21_X1 U8583 ( .B1(n9726), .B2(n6986), .A(n7054), .ZN(n6888) );
  OAI211_X1 U8584 ( .C1(n7057), .C2(n9731), .A(n7049), .B(n6888), .ZN(n6891)
         );
  NAND2_X1 U8585 ( .A1(n6891), .A2(n9796), .ZN(n6889) );
  OAI21_X1 U8586 ( .B1(n9796), .B2(n6890), .A(n6889), .ZN(P2_U3466) );
  INV_X1 U8587 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n6893) );
  NAND2_X1 U8588 ( .A1(n6891), .A2(n9810), .ZN(n6892) );
  OAI21_X1 U8589 ( .B1(n9810), .B2(n6893), .A(n6892), .ZN(P2_U3525) );
  INV_X1 U8590 ( .A(n6894), .ZN(n6950) );
  AOI22_X1 U8591 ( .A1(n8258), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_16__SCAN_IN), .B2(n8556), .ZN(n6895) );
  OAI21_X1 U8592 ( .B1(n6950), .B2(n8049), .A(n6895), .ZN(P2_U3342) );
  OAI211_X1 U8593 ( .C1(n6898), .C2(n6897), .A(n6896), .B(n8214), .ZN(n6901)
         );
  OAI22_X1 U8594 ( .A1(n7116), .A2(n8221), .B1(n7117), .B2(n8220), .ZN(n6899)
         );
  AOI21_X1 U8595 ( .B1(P2_REG3_REG_2__SCAN_IN), .B2(n8044), .A(n6899), .ZN(
        n6900) );
  OAI211_X1 U8596 ( .C1(n6875), .C2(n8227), .A(n6901), .B(n6900), .ZN(P2_U3239) );
  OR2_X1 U8597 ( .A1(n6902), .A2(n9676), .ZN(n6903) );
  OAI21_X1 U8598 ( .B1(n9362), .B2(n6904), .A(n6903), .ZN(P1_U3525) );
  INV_X1 U8599 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n9848) );
  NAND2_X1 U8600 ( .A1(n6978), .A2(n7052), .ZN(n6905) );
  XNOR2_X1 U8601 ( .A(n7167), .B(n6907), .ZN(n7442) );
  INV_X1 U8602 ( .A(n6907), .ZN(n6909) );
  NAND3_X1 U8603 ( .A1(n6910), .A2(n6909), .A3(n6908), .ZN(n6911) );
  AOI21_X1 U8604 ( .B1(n6912), .B2(n6911), .A(n9753), .ZN(n6915) );
  OR2_X1 U8605 ( .A1(n8139), .A2(n9756), .ZN(n6914) );
  OR2_X1 U8606 ( .A1(n6978), .A2(n9758), .ZN(n6913) );
  NAND2_X1 U8607 ( .A1(n6914), .A2(n6913), .ZN(n7155) );
  NOR2_X1 U8608 ( .A1(n6915), .A2(n7155), .ZN(n7437) );
  INV_X1 U8609 ( .A(n6916), .ZN(n6917) );
  NAND2_X1 U8610 ( .A1(n6916), .A2(n7436), .ZN(n7170) );
  INV_X1 U8611 ( .A(n7170), .ZN(n7171) );
  AOI211_X1 U8612 ( .C1(n7156), .C2(n6917), .A(n9780), .B(n7171), .ZN(n7440)
         );
  AOI21_X1 U8613 ( .B1(n9726), .B2(n7156), .A(n7440), .ZN(n6918) );
  OAI211_X1 U8614 ( .C1(n7442), .C2(n9731), .A(n7437), .B(n6918), .ZN(n6920)
         );
  NAND2_X1 U8615 ( .A1(n6920), .A2(n9796), .ZN(n6919) );
  OAI21_X1 U8616 ( .B1(n9796), .B2(n9848), .A(n6919), .ZN(P2_U3469) );
  INV_X1 U8617 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n6922) );
  NAND2_X1 U8618 ( .A1(n6920), .A2(n9810), .ZN(n6921) );
  OAI21_X1 U8619 ( .B1(n9810), .B2(n6922), .A(n6921), .ZN(P2_U3526) );
  INV_X1 U8620 ( .A(n6923), .ZN(n6924) );
  INV_X1 U8621 ( .A(n7864), .ZN(n7872) );
  OAI222_X1 U8622 ( .A1(n8051), .A2(n9884), .B1(n8049), .B2(n6924), .C1(
        P2_U3152), .C2(n7872), .ZN(P2_U3343) );
  OAI222_X1 U8623 ( .A1(n7085), .A2(n6925), .B1(n6951), .B2(n6924), .C1(
        P1_U3084), .C2(n7710), .ZN(P1_U3338) );
  NAND2_X1 U8624 ( .A1(n9021), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n6926) );
  OAI21_X1 U8625 ( .B1(n9075), .B2(n9021), .A(n6926), .ZN(P1_U3584) );
  INV_X1 U8626 ( .A(n8224), .ZN(n8177) );
  OAI211_X1 U8627 ( .C1(n6929), .C2(n6928), .A(n6927), .B(n8214), .ZN(n6933)
         );
  NOR2_X1 U8628 ( .A1(n5576), .A2(n8220), .ZN(n6931) );
  OAI22_X1 U8629 ( .A1(n6954), .A2(n8221), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n4911), .ZN(n6930) );
  AOI211_X1 U8630 ( .C1(n6962), .C2(n8207), .A(n6931), .B(n6930), .ZN(n6932)
         );
  OAI211_X1 U8631 ( .C1(P2_REG3_REG_3__SCAN_IN), .C2(n8177), .A(n6933), .B(
        n6932), .ZN(P2_U3220) );
  INV_X1 U8632 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n6934) );
  MUX2_X1 U8633 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n6934), .S(n7011), .Z(n6937)
         );
  INV_X1 U8634 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n9452) );
  AOI22_X1 U8635 ( .A1(n9536), .A2(P1_REG1_REG_11__SCAN_IN), .B1(n9452), .B2(
        n6940), .ZN(n9539) );
  OAI21_X1 U8636 ( .B1(P1_REG1_REG_10__SCAN_IN), .B2(n6942), .A(n6935), .ZN(
        n9538) );
  NAND2_X1 U8637 ( .A1(n6936), .A2(n6937), .ZN(n7005) );
  OAI21_X1 U8638 ( .B1(n6937), .B2(n6936), .A(n7005), .ZN(n6947) );
  NAND2_X1 U8639 ( .A1(n9573), .A2(P1_ADDR_REG_12__SCAN_IN), .ZN(n6938) );
  NAND2_X1 U8640 ( .A1(P1_U3084), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n7632) );
  OAI211_X1 U8641 ( .C1(n9045), .C2(n6939), .A(n6938), .B(n7632), .ZN(n6946)
         );
  XNOR2_X1 U8642 ( .A(n7011), .B(P1_REG2_REG_12__SCAN_IN), .ZN(n6944) );
  INV_X1 U8643 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n9844) );
  AOI22_X1 U8644 ( .A1(n9536), .A2(P1_REG2_REG_11__SCAN_IN), .B1(n9844), .B2(
        n6940), .ZN(n9542) );
  NAND2_X1 U8645 ( .A1(n9542), .A2(n9541), .ZN(n9540) );
  OAI21_X1 U8646 ( .B1(P1_REG2_REG_11__SCAN_IN), .B2(n9536), .A(n9540), .ZN(
        n6943) );
  NOR2_X1 U8647 ( .A1(n6943), .A2(n6944), .ZN(n7010) );
  AOI211_X1 U8648 ( .C1(n6944), .C2(n6943), .A(n9563), .B(n7010), .ZN(n6945)
         );
  AOI211_X1 U8649 ( .C1(n9574), .C2(n6947), .A(n6946), .B(n6945), .ZN(n6948)
         );
  INV_X1 U8650 ( .A(n6948), .ZN(P1_U3253) );
  INV_X1 U8651 ( .A(n9027), .ZN(n7718) );
  OAI222_X1 U8652 ( .A1(P1_U3084), .A2(n7718), .B1(n6951), .B2(n6950), .C1(
        n6949), .C2(n7085), .ZN(P1_U3337) );
  INV_X1 U8653 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n6966) );
  OAI21_X1 U8654 ( .B1(n6953), .B2(n6956), .A(n6952), .ZN(n7399) );
  INV_X1 U8655 ( .A(n7399), .ZN(n6964) );
  INV_X1 U8656 ( .A(n7563), .ZN(n9763) );
  OAI22_X1 U8657 ( .A1(n6954), .A2(n9756), .B1(n5576), .B2(n9758), .ZN(n6960)
         );
  NAND3_X1 U8658 ( .A1(n7114), .A2(n6956), .A3(n6955), .ZN(n6957) );
  AOI21_X1 U8659 ( .B1(n6958), .B2(n6957), .A(n9753), .ZN(n6959) );
  AOI211_X1 U8660 ( .C1(n9763), .C2(n7399), .A(n6960), .B(n6959), .ZN(n7401)
         );
  INV_X1 U8661 ( .A(n7034), .ZN(n6961) );
  AOI21_X1 U8662 ( .B1(n6962), .B2(n7118), .A(n6961), .ZN(n7395) );
  AOI22_X1 U8663 ( .A1(n7395), .A2(n9727), .B1(n9726), .B2(n6962), .ZN(n6963)
         );
  OAI211_X1 U8664 ( .C1(n6964), .C2(n9741), .A(n7401), .B(n6963), .ZN(n6967)
         );
  NAND2_X1 U8665 ( .A1(n6967), .A2(n9810), .ZN(n6965) );
  OAI21_X1 U8666 ( .B1(n9810), .B2(n6966), .A(n6965), .ZN(P2_U3523) );
  INV_X1 U8667 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n6969) );
  NAND2_X1 U8668 ( .A1(n6967), .A2(n9796), .ZN(n6968) );
  OAI21_X1 U8669 ( .B1(n9796), .B2(n6969), .A(n6968), .ZN(P2_U3460) );
  INV_X1 U8670 ( .A(n6970), .ZN(n6973) );
  AOI22_X1 U8671 ( .A1(n9042), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n9383), .ZN(n6971) );
  OAI21_X1 U8672 ( .B1(n6973), .B2(n6951), .A(n6971), .ZN(P1_U3336) );
  INV_X1 U8673 ( .A(n7875), .ZN(n7893) );
  OAI222_X1 U8674 ( .A1(P2_U3152), .A2(n7893), .B1(n8049), .B2(n6973), .C1(
        n6972), .C2(n8051), .ZN(P2_U3341) );
  NAND2_X1 U8675 ( .A1(n6975), .A2(n6974), .ZN(n6977) );
  XOR2_X1 U8676 ( .A(n6977), .B(n6976), .Z(n6982) );
  OAI22_X1 U8677 ( .A1(n7116), .A2(n9758), .B1(n6978), .B2(n9756), .ZN(n7031)
         );
  INV_X1 U8678 ( .A(n6979), .ZN(n8175) );
  AOI22_X1 U8679 ( .A1(n7031), .A2(n8175), .B1(P2_REG3_REG_4__SCAN_IN), .B2(
        P2_U3152), .ZN(n6981) );
  AOI22_X1 U8680 ( .A1(n8224), .A2(n7037), .B1(n9725), .B2(n8207), .ZN(n6980)
         );
  OAI211_X1 U8681 ( .C1(n6982), .C2(n8189), .A(n6981), .B(n6980), .ZN(P2_U3232) );
  XNOR2_X1 U8682 ( .A(n6984), .B(n6983), .ZN(n6989) );
  AOI22_X1 U8683 ( .A1(n6985), .A2(n8175), .B1(P2_REG3_REG_5__SCAN_IN), .B2(
        P2_U3152), .ZN(n6988) );
  AOI22_X1 U8684 ( .A1(n8224), .A2(n7050), .B1(n6986), .B2(n8207), .ZN(n6987)
         );
  OAI211_X1 U8685 ( .C1(n6989), .C2(n8189), .A(n6988), .B(n6987), .ZN(P2_U3229) );
  INV_X1 U8686 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n7000) );
  OAI21_X1 U8687 ( .B1(n6991), .B2(n8828), .A(n6990), .ZN(n7281) );
  INV_X1 U8688 ( .A(n7281), .ZN(n6998) );
  OAI22_X1 U8689 ( .A1(n6992), .A2(n6241), .B1(n7294), .B2(n9586), .ZN(n6995)
         );
  XNOR2_X1 U8690 ( .A(n8722), .B(n8828), .ZN(n6993) );
  NOR2_X1 U8691 ( .A1(n6993), .A2(n6240), .ZN(n6994) );
  AOI211_X1 U8692 ( .C1(n7726), .C2(n7281), .A(n6995), .B(n6994), .ZN(n7283)
         );
  AOI21_X1 U8693 ( .B1(n6996), .B2(n7098), .A(n7064), .ZN(n7277) );
  AOI22_X1 U8694 ( .A1(n7277), .A2(n9340), .B1(n9359), .B2(n6996), .ZN(n6997)
         );
  OAI211_X1 U8695 ( .C1(n6998), .C2(n7145), .A(n7283), .B(n6997), .ZN(n7001)
         );
  NAND2_X1 U8696 ( .A1(n7001), .A2(n9362), .ZN(n6999) );
  OAI21_X1 U8697 ( .B1(n9440), .B2(n7000), .A(n6999), .ZN(P1_U3527) );
  INV_X1 U8698 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n7003) );
  NAND2_X1 U8699 ( .A1(n7001), .A2(n9672), .ZN(n7002) );
  OAI21_X1 U8700 ( .B1(n9672), .B2(n7003), .A(n7002), .ZN(P1_U3466) );
  INV_X1 U8701 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n7004) );
  MUX2_X1 U8702 ( .A(P1_REG1_REG_13__SCAN_IN), .B(n7004), .S(n7601), .Z(n7007)
         );
  OAI21_X1 U8703 ( .B1(n7011), .B2(P1_REG1_REG_12__SCAN_IN), .A(n7005), .ZN(
        n7006) );
  OAI21_X1 U8704 ( .B1(n7007), .B2(n7006), .A(n7600), .ZN(n7018) );
  NAND2_X1 U8705 ( .A1(n9573), .A2(P1_ADDR_REG_13__SCAN_IN), .ZN(n7008) );
  NAND2_X1 U8706 ( .A1(P1_U3084), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n7697) );
  OAI211_X1 U8707 ( .C1(n9045), .C2(n7009), .A(n7008), .B(n7697), .ZN(n7017)
         );
  OR2_X1 U8708 ( .A1(n7601), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n7013) );
  NAND2_X1 U8709 ( .A1(P1_REG2_REG_13__SCAN_IN), .A2(n7601), .ZN(n7012) );
  NAND2_X1 U8710 ( .A1(n7013), .A2(n7012), .ZN(n7014) );
  AOI211_X1 U8711 ( .C1(n7015), .C2(n7014), .A(n9563), .B(n7594), .ZN(n7016)
         );
  AOI211_X1 U8712 ( .C1(n9574), .C2(n7018), .A(n7017), .B(n7016), .ZN(n7019)
         );
  INV_X1 U8713 ( .A(n7019), .ZN(P1_U3254) );
  OAI21_X1 U8714 ( .B1(n7022), .B2(n7021), .A(n7020), .ZN(n7023) );
  INV_X1 U8715 ( .A(n7023), .ZN(n9732) );
  NOR2_X1 U8716 ( .A1(n7025), .A2(n7024), .ZN(n7026) );
  NAND2_X1 U8717 ( .A1(n7027), .A2(n7026), .ZN(n7035) );
  OR2_X1 U8718 ( .A1(n7028), .A2(n5645), .ZN(n7206) );
  NAND2_X1 U8719 ( .A1(n7563), .A2(n7206), .ZN(n7029) );
  INV_X1 U8720 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n7327) );
  AOI21_X1 U8721 ( .B1(n7032), .B2(n9693), .A(n7031), .ZN(n9730) );
  MUX2_X1 U8722 ( .A(n7327), .B(n9730), .S(n7564), .Z(n7042) );
  AOI21_X1 U8723 ( .B1(n9725), .B2(n7034), .A(n7033), .ZN(n9728) );
  OR2_X1 U8724 ( .A1(n7035), .A2(n5295), .ZN(n7120) );
  NAND2_X1 U8725 ( .A1(n7564), .A2(n7036), .ZN(n8415) );
  INV_X1 U8726 ( .A(n7037), .ZN(n7038) );
  OAI22_X1 U8727 ( .A1(n8415), .A2(n7039), .B1(n7461), .B2(n7038), .ZN(n7040)
         );
  AOI21_X1 U8728 ( .B1(n9728), .B2(n8450), .A(n7040), .ZN(n7041) );
  OAI211_X1 U8729 ( .C1(n9732), .C2(n8452), .A(n7042), .B(n7041), .ZN(P2_U3292) );
  OAI22_X1 U8730 ( .A1(n9716), .A2(n9753), .B1(n7117), .B2(n9756), .ZN(n9718)
         );
  INV_X1 U8731 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n7043) );
  INV_X1 U8732 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n9933) );
  OAI22_X1 U8733 ( .A1(n7564), .A2(n7043), .B1(n9933), .B2(n7461), .ZN(n7044)
         );
  AOI21_X1 U8734 ( .B1(n9718), .B2(n7564), .A(n7044), .ZN(n7047) );
  OAI21_X1 U8735 ( .B1(n9996), .B2(n8450), .A(n7045), .ZN(n7046) );
  OAI211_X1 U8736 ( .C1(n9716), .C2(n8452), .A(n7047), .B(n7046), .ZN(P2_U3296) );
  INV_X1 U8737 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n7048) );
  MUX2_X1 U8738 ( .A(n7049), .B(n7048), .S(n9706), .Z(n7056) );
  INV_X1 U8739 ( .A(n7050), .ZN(n7051) );
  OAI22_X1 U8740 ( .A1(n8415), .A2(n7052), .B1(n7461), .B2(n7051), .ZN(n7053)
         );
  AOI21_X1 U8741 ( .B1(n7054), .B2(n9702), .A(n7053), .ZN(n7055) );
  OAI211_X1 U8742 ( .C1(n7057), .C2(n8452), .A(n7056), .B(n7055), .ZN(P2_U3291) );
  NOR2_X1 U8743 ( .A1(n7063), .A2(n4446), .ZN(n7058) );
  AOI21_X1 U8744 ( .B1(n8723), .B2(n8901), .A(n6271), .ZN(n7136) );
  AOI21_X1 U8745 ( .B1(n7058), .B2(n8723), .A(n7136), .ZN(n7059) );
  OAI222_X1 U8746 ( .A1(n9586), .A2(n7185), .B1(n6241), .B2(n7103), .C1(n6240), 
        .C2(n7059), .ZN(n9658) );
  INV_X1 U8747 ( .A(n9658), .ZN(n7074) );
  INV_X1 U8748 ( .A(n7060), .ZN(n7061) );
  AOI21_X1 U8749 ( .B1(n7063), .B2(n7062), .A(n7061), .ZN(n9661) );
  INV_X1 U8750 ( .A(n9271), .ZN(n9189) );
  OAI21_X1 U8751 ( .B1(n7064), .B2(n9657), .A(n9340), .ZN(n7065) );
  OR2_X1 U8752 ( .A1(n7065), .A2(n7141), .ZN(n9656) );
  INV_X1 U8753 ( .A(n9169), .ZN(n7071) );
  INV_X1 U8754 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n7067) );
  INV_X1 U8755 ( .A(n7129), .ZN(n7066) );
  OAI22_X1 U8756 ( .A1(n9609), .A2(n7067), .B1(n7066), .B2(n9613), .ZN(n7068)
         );
  AOI21_X1 U8757 ( .B1(n9605), .B2(n7069), .A(n7068), .ZN(n7070) );
  OAI21_X1 U8758 ( .B1(n9656), .B2(n7071), .A(n7070), .ZN(n7072) );
  AOI21_X1 U8759 ( .B1(n9661), .B2(n9189), .A(n7072), .ZN(n7073) );
  OAI21_X1 U8760 ( .B1(n7074), .B2(n9597), .A(n7073), .ZN(P1_U3286) );
  XNOR2_X1 U8761 ( .A(n7076), .B(n7075), .ZN(n7077) );
  XNOR2_X1 U8762 ( .A(n7078), .B(n7077), .ZN(n7079) );
  NAND2_X1 U8763 ( .A1(n7079), .A2(n8700), .ZN(n7083) );
  AND2_X1 U8764 ( .A1(P1_U3084), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n9497) );
  INV_X1 U8765 ( .A(n7189), .ZN(n7080) );
  OAI22_X1 U8766 ( .A1(n8707), .A2(n7080), .B1(n8705), .B2(n7185), .ZN(n7081)
         );
  AOI211_X1 U8767 ( .C1(n8710), .C2(n9014), .A(n9497), .B(n7081), .ZN(n7082)
         );
  OAI211_X1 U8768 ( .C1(n7192), .C2(n8713), .A(n7083), .B(n7082), .ZN(P1_U3211) );
  INV_X1 U8769 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n9935) );
  INV_X1 U8770 ( .A(n7084), .ZN(n7086) );
  INV_X1 U8771 ( .A(n9569), .ZN(n9040) );
  OAI222_X1 U8772 ( .A1(n7085), .A2(n9935), .B1(n6951), .B2(n7086), .C1(
        P1_U3084), .C2(n9040), .ZN(P1_U3335) );
  INV_X1 U8773 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n7087) );
  INV_X1 U8774 ( .A(n8022), .ZN(n7881) );
  OAI222_X1 U8775 ( .A1(n8051), .A2(n7087), .B1(n8049), .B2(n7086), .C1(
        P2_U3152), .C2(n7881), .ZN(P2_U3340) );
  INV_X1 U8776 ( .A(n7088), .ZN(n8048) );
  AOI22_X1 U8777 ( .A1(n9248), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_19__SCAN_IN), .B2(n9389), .ZN(n7089) );
  OAI21_X1 U8778 ( .B1(n8048), .B2(n6951), .A(n7089), .ZN(P1_U3334) );
  AND2_X1 U8779 ( .A1(n7090), .A2(n9248), .ZN(n7091) );
  OAI21_X1 U8780 ( .B1(n7093), .B2(n7102), .A(n7092), .ZN(n9654) );
  NOR2_X1 U8781 ( .A1(n7094), .A2(n8990), .ZN(n7095) );
  INV_X1 U8782 ( .A(n9604), .ZN(n9066) );
  NAND2_X1 U8783 ( .A1(n7096), .A2(n7100), .ZN(n7097) );
  NAND2_X1 U8784 ( .A1(n7098), .A2(n7097), .ZN(n9651) );
  AOI22_X1 U8785 ( .A1(n9605), .A2(n7100), .B1(n9595), .B2(n7099), .ZN(n7101)
         );
  OAI21_X1 U8786 ( .B1(n9066), .B2(n9651), .A(n7101), .ZN(n7110) );
  XNOR2_X1 U8787 ( .A(n8911), .B(n7102), .ZN(n7108) );
  NAND2_X1 U8788 ( .A1(n9654), .A2(n7726), .ZN(n7107) );
  OAI22_X1 U8789 ( .A1(n7104), .A2(n6241), .B1(n7103), .B2(n9586), .ZN(n7105)
         );
  INV_X1 U8790 ( .A(n7105), .ZN(n7106) );
  OAI211_X1 U8791 ( .C1(n6240), .C2(n7108), .A(n7107), .B(n7106), .ZN(n9652)
         );
  MUX2_X1 U8792 ( .A(n9652), .B(P1_REG2_REG_3__SCAN_IN), .S(n9597), .Z(n7109)
         );
  AOI211_X1 U8793 ( .C1(n9583), .C2(n9654), .A(n7110), .B(n7109), .ZN(n7111)
         );
  INV_X1 U8794 ( .A(n7111), .ZN(P1_U3288) );
  XNOR2_X1 U8795 ( .A(n7113), .B(n7112), .ZN(n9723) );
  INV_X1 U8796 ( .A(n9723), .ZN(n7126) );
  INV_X1 U8797 ( .A(n7114), .ZN(n7115) );
  OAI222_X1 U8798 ( .A1(n9758), .A2(n7117), .B1(n9756), .B2(n7116), .C1(n9753), 
        .C2(n4357), .ZN(n9721) );
  NAND2_X1 U8799 ( .A1(n9721), .A2(n7564), .ZN(n7125) );
  OAI211_X1 U8800 ( .C1(n7119), .C2(n6875), .A(n7118), .B(n9727), .ZN(n9720)
         );
  INV_X1 U8801 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n8002) );
  OAI22_X1 U8802 ( .A1(n9720), .A2(n7120), .B1(n8002), .B2(n7461), .ZN(n7122)
         );
  INV_X1 U8803 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n9883) );
  NOR2_X1 U8804 ( .A1(n7564), .A2(n9883), .ZN(n7121) );
  AOI211_X1 U8805 ( .C1(n9996), .C2(n7123), .A(n7122), .B(n7121), .ZN(n7124)
         );
  OAI211_X1 U8806 ( .C1(n7126), .C2(n8452), .A(n7125), .B(n7124), .ZN(P2_U3294) );
  XNOR2_X1 U8807 ( .A(n7285), .B(n7286), .ZN(n7128) );
  NOR2_X1 U8808 ( .A1(n7128), .A2(n7127), .ZN(n7284) );
  AOI21_X1 U8809 ( .B1(n7128), .B2(n7127), .A(n7284), .ZN(n7133) );
  AOI22_X1 U8810 ( .A1(n8668), .A2(n9018), .B1(n7129), .B2(n8690), .ZN(n7132)
         );
  AND2_X1 U8811 ( .A1(P1_U3084), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n9477) );
  NOR2_X1 U8812 ( .A1(n8713), .A2(n9657), .ZN(n7130) );
  AOI211_X1 U8813 ( .C1(n8710), .C2(n9016), .A(n9477), .B(n7130), .ZN(n7131)
         );
  OAI211_X1 U8814 ( .C1(n7133), .C2(n8682), .A(n7132), .B(n7131), .ZN(P1_U3225) );
  INV_X1 U8815 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n7148) );
  OAI21_X1 U8816 ( .B1(n7135), .B2(n8729), .A(n7134), .ZN(n7164) );
  INV_X1 U8817 ( .A(n7164), .ZN(n7146) );
  INV_X1 U8818 ( .A(n8902), .ZN(n8727) );
  NOR2_X1 U8819 ( .A1(n7136), .A2(n8727), .ZN(n7137) );
  XOR2_X1 U8820 ( .A(n8729), .B(n7137), .Z(n7139) );
  AOI22_X1 U8821 ( .A1(n9233), .A2(n9017), .B1(n9015), .B2(n9231), .ZN(n7138)
         );
  OAI21_X1 U8822 ( .B1(n7139), .B2(n6240), .A(n7138), .ZN(n7140) );
  AOI21_X1 U8823 ( .B1(n7726), .B2(n7164), .A(n7140), .ZN(n7166) );
  INV_X1 U8824 ( .A(n7141), .ZN(n7142) );
  AOI21_X1 U8825 ( .B1(n7143), .B2(n7142), .A(n4547), .ZN(n7160) );
  AOI22_X1 U8826 ( .A1(n7160), .A2(n9340), .B1(n9359), .B2(n7143), .ZN(n7144)
         );
  OAI211_X1 U8827 ( .C1(n7146), .C2(n7145), .A(n7166), .B(n7144), .ZN(n7149)
         );
  NAND2_X1 U8828 ( .A1(n7149), .A2(n9440), .ZN(n7147) );
  OAI21_X1 U8829 ( .B1(n9440), .B2(n7148), .A(n7147), .ZN(P1_U3529) );
  INV_X1 U8830 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n7151) );
  NAND2_X1 U8831 ( .A1(n7149), .A2(n9672), .ZN(n7150) );
  OAI21_X1 U8832 ( .B1(n9672), .B2(n7151), .A(n7150), .ZN(P1_U3472) );
  INV_X1 U8833 ( .A(n8080), .ZN(n7152) );
  AOI21_X1 U8834 ( .B1(n7154), .B2(n7153), .A(n7152), .ZN(n7159) );
  AOI22_X1 U8835 ( .A1(n7155), .A2(n8175), .B1(P2_REG3_REG_6__SCAN_IN), .B2(
        P2_U3152), .ZN(n7158) );
  AOI22_X1 U8836 ( .A1(n8224), .A2(n7434), .B1(n7156), .B2(n8207), .ZN(n7157)
         );
  OAI211_X1 U8837 ( .C1(n7159), .C2(n8189), .A(n7158), .B(n7157), .ZN(P2_U3241) );
  NAND2_X1 U8838 ( .A1(n7160), .A2(n9604), .ZN(n7162) );
  AOI22_X1 U8839 ( .A1(n9597), .A2(P1_REG2_REG_6__SCAN_IN), .B1(n7293), .B2(
        n9595), .ZN(n7161) );
  OAI211_X1 U8840 ( .C1(n7299), .C2(n9599), .A(n7162), .B(n7161), .ZN(n7163)
         );
  AOI21_X1 U8841 ( .B1(n7164), .B2(n9583), .A(n7163), .ZN(n7165) );
  OAI21_X1 U8842 ( .B1(n7166), .B2(n9597), .A(n7165), .ZN(P1_U3285) );
  XNOR2_X1 U8843 ( .A(n7198), .B(n7197), .ZN(n9739) );
  INV_X1 U8844 ( .A(n9739), .ZN(n7176) );
  XNOR2_X1 U8845 ( .A(n7168), .B(n7197), .ZN(n7169) );
  OAI222_X1 U8846 ( .A1(n9756), .A2(n9759), .B1(n9758), .B2(n8084), .C1(n7169), 
        .C2(n9753), .ZN(n9737) );
  OAI21_X1 U8847 ( .B1(n7171), .B2(n9735), .A(n7412), .ZN(n9736) );
  AOI22_X1 U8848 ( .A1(n9706), .A2(P2_REG2_REG_7__SCAN_IN), .B1(n8088), .B2(
        n9993), .ZN(n7173) );
  NAND2_X1 U8849 ( .A1(n9996), .A2(n8087), .ZN(n7172) );
  OAI211_X1 U8850 ( .C1(n9736), .C2(n9999), .A(n7173), .B(n7172), .ZN(n7174)
         );
  AOI21_X1 U8851 ( .B1(n9737), .B2(n7564), .A(n7174), .ZN(n7175) );
  OAI21_X1 U8852 ( .B1(n7176), .B2(n8452), .A(n7175), .ZN(P2_U3289) );
  OAI21_X1 U8853 ( .B1(n7178), .B2(n7183), .A(n7177), .ZN(n7179) );
  INV_X1 U8854 ( .A(n7179), .ZN(n7223) );
  INV_X1 U8855 ( .A(n7180), .ZN(n7181) );
  AOI21_X1 U8856 ( .B1(n7183), .B2(n7182), .A(n7181), .ZN(n7184) );
  OAI222_X1 U8857 ( .A1(n9586), .A2(n9588), .B1(n6241), .B2(n7185), .C1(n6240), 
        .C2(n7184), .ZN(n7219) );
  INV_X1 U8858 ( .A(n7246), .ZN(n7186) );
  AOI211_X1 U8859 ( .C1(n7221), .C2(n7187), .A(n9664), .B(n7186), .ZN(n7220)
         );
  OR2_X1 U8860 ( .A1(n7188), .A2(n9248), .ZN(n9267) );
  INV_X1 U8861 ( .A(n9267), .ZN(n7490) );
  NAND2_X1 U8862 ( .A1(n7220), .A2(n7490), .ZN(n7191) );
  AOI22_X1 U8863 ( .A1(n9597), .A2(P1_REG2_REG_7__SCAN_IN), .B1(n7189), .B2(
        n9595), .ZN(n7190) );
  OAI211_X1 U8864 ( .C1(n7192), .C2(n9599), .A(n7191), .B(n7190), .ZN(n7193)
         );
  AOI21_X1 U8865 ( .B1(n7219), .B2(n9609), .A(n7193), .ZN(n7194) );
  OAI21_X1 U8866 ( .B1(n7223), .B2(n9271), .A(n7194), .ZN(P1_U3284) );
  INV_X1 U8867 ( .A(n7195), .ZN(n7377) );
  AOI22_X1 U8868 ( .A1(n8942), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_20__SCAN_IN), .B2(n9383), .ZN(n7196) );
  OAI21_X1 U8869 ( .B1(n7377), .B2(n6951), .A(n7196), .ZN(P1_U3333) );
  NAND2_X1 U8870 ( .A1(n7198), .A2(n7197), .ZN(n7200) );
  NAND2_X1 U8871 ( .A1(n8139), .A2(n9735), .ZN(n7199) );
  NAND2_X1 U8872 ( .A1(n8241), .A2(n8142), .ZN(n7202) );
  NAND2_X1 U8873 ( .A1(n8138), .A2(n9767), .ZN(n7203) );
  NAND2_X1 U8874 ( .A1(n7205), .A2(n7204), .ZN(n7254) );
  OAI21_X1 U8875 ( .B1(n7205), .B2(n7204), .A(n7254), .ZN(n9771) );
  INV_X1 U8876 ( .A(n7206), .ZN(n7207) );
  NAND2_X1 U8877 ( .A1(n7564), .A2(n7207), .ZN(n7570) );
  XNOR2_X1 U8878 ( .A(n7208), .B(n7209), .ZN(n7211) );
  OAI22_X1 U8879 ( .A1(n8138), .A2(n9758), .B1(n8112), .B2(n9756), .ZN(n7210)
         );
  AOI21_X1 U8880 ( .B1(n7211), .B2(n9693), .A(n7210), .ZN(n7212) );
  OAI21_X1 U8881 ( .B1(n9771), .B2(n7563), .A(n7212), .ZN(n9774) );
  NAND2_X1 U8882 ( .A1(n9774), .A2(n7564), .ZN(n7218) );
  INV_X1 U8883 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n7214) );
  INV_X1 U8884 ( .A(n8116), .ZN(n7213) );
  OAI22_X1 U8885 ( .A1(n7564), .A2(n7214), .B1(n7213), .B2(n7461), .ZN(n7216)
         );
  OAI21_X1 U8886 ( .B1(n9766), .B2(n9772), .A(n7260), .ZN(n9773) );
  NOR2_X1 U8887 ( .A1(n9773), .A2(n9999), .ZN(n7215) );
  AOI211_X1 U8888 ( .C1(n9996), .C2(n8115), .A(n7216), .B(n7215), .ZN(n7217)
         );
  OAI211_X1 U8889 ( .C1(n9771), .C2(n7570), .A(n7218), .B(n7217), .ZN(P2_U3286) );
  INV_X1 U8890 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n7225) );
  AOI211_X1 U8891 ( .C1(n9359), .C2(n7221), .A(n7220), .B(n7219), .ZN(n7222)
         );
  OAI21_X1 U8892 ( .B1(n9426), .B2(n7223), .A(n7222), .ZN(n7239) );
  NAND2_X1 U8893 ( .A1(n7239), .A2(n9440), .ZN(n7224) );
  OAI21_X1 U8894 ( .B1(n9362), .B2(n7225), .A(n7224), .ZN(P1_U3530) );
  NAND2_X1 U8895 ( .A1(n8133), .A2(n7226), .ZN(n7228) );
  AND2_X1 U8896 ( .A1(n7228), .A2(n7227), .ZN(n7233) );
  NAND2_X1 U8897 ( .A1(n7230), .A2(n7229), .ZN(n7231) );
  AOI21_X1 U8898 ( .B1(n7233), .B2(n7232), .A(n7231), .ZN(n7238) );
  NOR2_X1 U8899 ( .A1(n8227), .A2(n9767), .ZN(n7236) );
  NAND2_X1 U8900 ( .A1(n8239), .A2(n8195), .ZN(n7234) );
  NAND2_X1 U8901 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(P2_U3152), .ZN(n7919) );
  OAI211_X1 U8902 ( .C1(n9759), .C2(n8220), .A(n7234), .B(n7919), .ZN(n7235)
         );
  AOI211_X1 U8903 ( .C1(n8224), .C2(n9994), .A(n7236), .B(n7235), .ZN(n7237)
         );
  OAI21_X1 U8904 ( .B1(n7238), .B2(n8189), .A(n7237), .ZN(P2_U3233) );
  INV_X1 U8905 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n7241) );
  NAND2_X1 U8906 ( .A1(n7239), .A2(n9672), .ZN(n7240) );
  OAI21_X1 U8907 ( .B1(n9672), .B2(n7241), .A(n7240), .ZN(P1_U3475) );
  INV_X1 U8908 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n7249) );
  OAI21_X1 U8909 ( .B1(n7243), .B2(n6275), .A(n7242), .ZN(n7274) );
  XNOR2_X1 U8910 ( .A(n7244), .B(n8832), .ZN(n7245) );
  AOI222_X1 U8911 ( .A1(n9590), .A2(n7245), .B1(n9013), .B2(n9231), .C1(n9015), 
        .C2(n9233), .ZN(n7269) );
  AOI21_X1 U8912 ( .B1(n7267), .B2(n7246), .A(n9579), .ZN(n7272) );
  AOI22_X1 U8913 ( .A1(n7272), .A2(n9340), .B1(n9359), .B2(n7267), .ZN(n7247)
         );
  OAI211_X1 U8914 ( .C1(n7274), .C2(n9426), .A(n7269), .B(n7247), .ZN(n7250)
         );
  NAND2_X1 U8915 ( .A1(n7250), .A2(n9440), .ZN(n7248) );
  OAI21_X1 U8916 ( .B1(n9362), .B2(n7249), .A(n7248), .ZN(P1_U3531) );
  INV_X1 U8917 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n7252) );
  NAND2_X1 U8918 ( .A1(n7250), .A2(n9672), .ZN(n7251) );
  OAI21_X1 U8919 ( .B1(n9672), .B2(n7252), .A(n7251), .ZN(P1_U3478) );
  NAND2_X1 U8920 ( .A1(n8239), .A2(n8115), .ZN(n7253) );
  NAND2_X1 U8921 ( .A1(n7254), .A2(n7253), .ZN(n7255) );
  NAND2_X1 U8922 ( .A1(n7255), .A2(n7257), .ZN(n7552) );
  OR2_X1 U8923 ( .A1(n7255), .A2(n7257), .ZN(n7256) );
  AND2_X1 U8924 ( .A1(n7552), .A2(n7256), .ZN(n9784) );
  INV_X1 U8925 ( .A(n9784), .ZN(n7266) );
  XNOR2_X1 U8926 ( .A(n7258), .B(n7257), .ZN(n7259) );
  OAI222_X1 U8927 ( .A1(n9756), .A2(n8204), .B1(n9758), .B2(n9757), .C1(n7259), 
        .C2(n9753), .ZN(n9782) );
  INV_X1 U8928 ( .A(n7260), .ZN(n7261) );
  INV_X1 U8929 ( .A(n8208), .ZN(n9779) );
  OAI21_X1 U8930 ( .B1(n7261), .B2(n9779), .A(n9698), .ZN(n9781) );
  AOI22_X1 U8931 ( .A1(n9706), .A2(P2_REG2_REG_11__SCAN_IN), .B1(n8209), .B2(
        n9993), .ZN(n7263) );
  NAND2_X1 U8932 ( .A1(n9996), .A2(n8208), .ZN(n7262) );
  OAI211_X1 U8933 ( .C1(n9781), .C2(n9999), .A(n7263), .B(n7262), .ZN(n7264)
         );
  AOI21_X1 U8934 ( .B1(n9782), .B2(n7564), .A(n7264), .ZN(n7265) );
  OAI21_X1 U8935 ( .B1(n8452), .B2(n7266), .A(n7265), .ZN(P2_U3285) );
  INV_X1 U8936 ( .A(n7267), .ZN(n7312) );
  AOI22_X1 U8937 ( .A1(n9597), .A2(P1_REG2_REG_8__SCAN_IN), .B1(n7306), .B2(
        n9595), .ZN(n7268) );
  OAI21_X1 U8938 ( .B1(n9599), .B2(n7312), .A(n7268), .ZN(n7271) );
  NOR2_X1 U8939 ( .A1(n7269), .A2(n9597), .ZN(n7270) );
  AOI211_X1 U8940 ( .C1(n7272), .C2(n9604), .A(n7271), .B(n7270), .ZN(n7273)
         );
  OAI21_X1 U8941 ( .B1(n9271), .B2(n7274), .A(n7273), .ZN(P1_U3283) );
  INV_X1 U8942 ( .A(n7275), .ZN(n7379) );
  AOI22_X1 U8943 ( .A1(n8951), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_21__SCAN_IN), .B2(n9389), .ZN(n7276) );
  OAI21_X1 U8944 ( .B1(n7379), .B2(n6951), .A(n7276), .ZN(P1_U3332) );
  NAND2_X1 U8945 ( .A1(n7277), .A2(n9604), .ZN(n7279) );
  AOI22_X1 U8946 ( .A1(n9597), .A2(P1_REG2_REG_4__SCAN_IN), .B1(n8638), .B2(
        n9595), .ZN(n7278) );
  OAI211_X1 U8947 ( .C1(n8636), .C2(n9599), .A(n7279), .B(n7278), .ZN(n7280)
         );
  AOI21_X1 U8948 ( .B1(n7281), .B2(n9583), .A(n7280), .ZN(n7282) );
  OAI21_X1 U8949 ( .B1(n7283), .B2(n9597), .A(n7282), .ZN(P1_U3287) );
  AOI21_X1 U8950 ( .B1(n7286), .B2(n7285), .A(n7284), .ZN(n7290) );
  XNOR2_X1 U8951 ( .A(n7288), .B(n7287), .ZN(n7289) );
  XNOR2_X1 U8952 ( .A(n7290), .B(n7289), .ZN(n7291) );
  NAND2_X1 U8953 ( .A1(n7291), .A2(n8700), .ZN(n7298) );
  NOR2_X1 U8954 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7292), .ZN(n9489) );
  INV_X1 U8955 ( .A(n7293), .ZN(n7295) );
  OAI22_X1 U8956 ( .A1(n8707), .A2(n7295), .B1(n8705), .B2(n7294), .ZN(n7296)
         );
  AOI211_X1 U8957 ( .C1(n8710), .C2(n9015), .A(n9489), .B(n7296), .ZN(n7297)
         );
  OAI211_X1 U8958 ( .C1(n7299), .C2(n8713), .A(n7298), .B(n7297), .ZN(P1_U3237) );
  INV_X1 U8959 ( .A(n7369), .ZN(n7304) );
  AOI21_X1 U8960 ( .B1(n7369), .B2(n7301), .A(n7300), .ZN(n7302) );
  NOR2_X1 U8961 ( .A1(n7302), .A2(n8682), .ZN(n7303) );
  OAI21_X1 U8962 ( .B1(n7304), .B2(n7370), .A(n7303), .ZN(n7311) );
  NOR2_X1 U8963 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7305), .ZN(n9515) );
  INV_X1 U8964 ( .A(n7306), .ZN(n7308) );
  OAI22_X1 U8965 ( .A1(n8707), .A2(n7308), .B1(n8705), .B2(n7307), .ZN(n7309)
         );
  AOI211_X1 U8966 ( .C1(n8710), .C2(n9013), .A(n9515), .B(n7309), .ZN(n7310)
         );
  OAI211_X1 U8967 ( .C1(n7312), .C2(n8713), .A(n7311), .B(n7310), .ZN(P1_U3219) );
  INV_X1 U8968 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n7315) );
  NOR2_X1 U8969 ( .A1(n7450), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n7444) );
  INV_X1 U8970 ( .A(n7444), .ZN(n7313) );
  OAI21_X1 U8971 ( .B1(n7315), .B2(n7314), .A(n7313), .ZN(n7338) );
  INV_X1 U8972 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n7336) );
  NAND2_X1 U8973 ( .A1(n7355), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n7335) );
  MUX2_X1 U8974 ( .A(P2_REG2_REG_10__SCAN_IN), .B(n7214), .S(n7355), .Z(n7914)
         );
  NAND2_X1 U8975 ( .A1(n7353), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n7334) );
  INV_X1 U8976 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n7316) );
  MUX2_X1 U8977 ( .A(n7316), .B(P2_REG2_REG_9__SCAN_IN), .S(n7353), .Z(n7317)
         );
  INV_X1 U8978 ( .A(n7317), .ZN(n7926) );
  NAND2_X1 U8979 ( .A1(n7351), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n7333) );
  INV_X1 U8980 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n7318) );
  MUX2_X1 U8981 ( .A(n7318), .B(P2_REG2_REG_8__SCAN_IN), .S(n7351), .Z(n7319)
         );
  INV_X1 U8982 ( .A(n7319), .ZN(n7937) );
  NAND2_X1 U8983 ( .A1(n7349), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n7332) );
  INV_X1 U8984 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n7320) );
  MUX2_X1 U8985 ( .A(n7320), .B(P2_REG2_REG_7__SCAN_IN), .S(n7349), .Z(n7321)
         );
  INV_X1 U8986 ( .A(n7321), .ZN(n7948) );
  NAND2_X1 U8987 ( .A1(n7347), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n7331) );
  INV_X1 U8988 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n7322) );
  MUX2_X1 U8989 ( .A(P2_REG2_REG_6__SCAN_IN), .B(n7322), .S(n7347), .Z(n7960)
         );
  NAND2_X1 U8990 ( .A1(n7345), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n7330) );
  MUX2_X1 U8991 ( .A(P2_REG2_REG_5__SCAN_IN), .B(n7048), .S(n4280), .Z(n7323)
         );
  INV_X1 U8992 ( .A(n7323), .ZN(n7971) );
  INV_X1 U8993 ( .A(n8011), .ZN(n7326) );
  NOR2_X1 U8994 ( .A1(n7324), .A2(n6699), .ZN(n8009) );
  MUX2_X1 U8995 ( .A(P2_REG2_REG_2__SCAN_IN), .B(n9883), .S(n8008), .Z(n7325)
         );
  OAI21_X1 U8996 ( .B1(n7326), .B2(n8009), .A(n7325), .ZN(n8014) );
  NAND2_X1 U8997 ( .A1(n8008), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n7996) );
  INV_X1 U8998 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n7393) );
  MUX2_X1 U8999 ( .A(n7393), .B(P2_REG2_REG_3__SCAN_IN), .S(n7342), .Z(n7995)
         );
  AOI21_X1 U9000 ( .B1(n8014), .B2(n7996), .A(n7995), .ZN(n7980) );
  NOR2_X1 U9001 ( .A1(n8001), .A2(n7393), .ZN(n7981) );
  MUX2_X1 U9002 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n7327), .S(n7982), .Z(n7328)
         );
  OAI21_X1 U9003 ( .B1(n7980), .B2(n7981), .A(n7328), .ZN(n7986) );
  NAND2_X1 U9004 ( .A1(n7982), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n7329) );
  NAND2_X1 U9005 ( .A1(n7986), .A2(n7329), .ZN(n7972) );
  NAND2_X1 U9006 ( .A1(n7971), .A2(n7972), .ZN(n7970) );
  NAND2_X1 U9007 ( .A1(n7330), .A2(n7970), .ZN(n7961) );
  NAND2_X1 U9008 ( .A1(n7960), .A2(n7961), .ZN(n7959) );
  NAND2_X1 U9009 ( .A1(n7331), .A2(n7959), .ZN(n7949) );
  NAND2_X1 U9010 ( .A1(n7948), .A2(n7949), .ZN(n7947) );
  NAND2_X1 U9011 ( .A1(n7332), .A2(n7947), .ZN(n7938) );
  NAND2_X1 U9012 ( .A1(n7937), .A2(n7938), .ZN(n7936) );
  NAND2_X1 U9013 ( .A1(n7333), .A2(n7936), .ZN(n7927) );
  NAND2_X1 U9014 ( .A1(n7926), .A2(n7927), .ZN(n7925) );
  NAND2_X1 U9015 ( .A1(n7334), .A2(n7925), .ZN(n7915) );
  NAND2_X1 U9016 ( .A1(n7914), .A2(n7915), .ZN(n7913) );
  NAND2_X1 U9017 ( .A1(n7335), .A2(n7913), .ZN(n7896) );
  MUX2_X1 U9018 ( .A(n7336), .B(P2_REG2_REG_11__SCAN_IN), .S(n7357), .Z(n7895)
         );
  NOR2_X1 U9019 ( .A1(n7896), .A2(n7895), .ZN(n7894) );
  AOI21_X1 U9020 ( .B1(n7907), .B2(n7336), .A(n7894), .ZN(n7337) );
  NOR2_X1 U9021 ( .A1(n7337), .A2(n7338), .ZN(n7443) );
  AOI21_X1 U9022 ( .B1(n7338), .B2(n7337), .A(n7443), .ZN(n7366) );
  INV_X1 U9023 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n7363) );
  AOI21_X1 U9024 ( .B1(P2_REG1_REG_1__SCAN_IN), .B2(n7340), .A(n7339), .ZN(
        n8005) );
  INV_X1 U9025 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n7341) );
  MUX2_X1 U9026 ( .A(n7341), .B(P2_REG1_REG_2__SCAN_IN), .S(n8008), .Z(n8004)
         );
  MUX2_X1 U9027 ( .A(n6966), .B(P2_REG1_REG_3__SCAN_IN), .S(n7342), .Z(n7991)
         );
  NAND2_X1 U9028 ( .A1(n7982), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n7343) );
  OAI21_X1 U9029 ( .B1(n7982), .B2(P2_REG1_REG_4__SCAN_IN), .A(n7343), .ZN(
        n7976) );
  NOR2_X1 U9030 ( .A1(n7977), .A2(n7976), .ZN(n7975) );
  NAND2_X1 U9031 ( .A1(n7345), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n7344) );
  OAI21_X1 U9032 ( .B1(n7345), .B2(P2_REG1_REG_5__SCAN_IN), .A(n7344), .ZN(
        n7966) );
  NAND2_X1 U9033 ( .A1(n7347), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n7346) );
  OAI21_X1 U9034 ( .B1(n7347), .B2(P2_REG1_REG_6__SCAN_IN), .A(n7346), .ZN(
        n7955) );
  AOI21_X1 U9035 ( .B1(n7347), .B2(P2_REG1_REG_6__SCAN_IN), .A(n7954), .ZN(
        n7944) );
  NAND2_X1 U9036 ( .A1(n7349), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n7348) );
  OAI21_X1 U9037 ( .B1(n7349), .B2(P2_REG1_REG_7__SCAN_IN), .A(n7348), .ZN(
        n7943) );
  NOR2_X1 U9038 ( .A1(n7944), .A2(n7943), .ZN(n7942) );
  AOI21_X1 U9039 ( .B1(n7349), .B2(P2_REG1_REG_7__SCAN_IN), .A(n7942), .ZN(
        n7933) );
  INV_X1 U9040 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n7350) );
  MUX2_X1 U9041 ( .A(n7350), .B(P2_REG1_REG_8__SCAN_IN), .S(n7351), .Z(n7932)
         );
  INV_X1 U9042 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n7352) );
  MUX2_X1 U9043 ( .A(n7352), .B(P2_REG1_REG_9__SCAN_IN), .S(n7353), .Z(n7921)
         );
  INV_X1 U9044 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n7354) );
  MUX2_X1 U9045 ( .A(n7354), .B(P2_REG1_REG_10__SCAN_IN), .S(n7355), .Z(n7909)
         );
  NOR2_X1 U9046 ( .A1(n7910), .A2(n7909), .ZN(n7908) );
  INV_X1 U9047 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n7356) );
  MUX2_X1 U9048 ( .A(n7356), .B(P2_REG1_REG_11__SCAN_IN), .S(n7357), .Z(n7900)
         );
  INV_X1 U9049 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n7358) );
  MUX2_X1 U9050 ( .A(P2_REG1_REG_12__SCAN_IN), .B(n7358), .S(n7450), .Z(n7359)
         );
  OAI21_X1 U9051 ( .B1(n7360), .B2(n7359), .A(n7449), .ZN(n7361) );
  NAND2_X1 U9052 ( .A1(n9679), .A2(n7361), .ZN(n7362) );
  NAND2_X1 U9053 ( .A1(P2_U3152), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n7609) );
  OAI211_X1 U9054 ( .C1(n8033), .C2(n7363), .A(n7362), .B(n7609), .ZN(n7364)
         );
  AOI21_X1 U9055 ( .B1(n9684), .B2(n7450), .A(n7364), .ZN(n7365) );
  OAI21_X1 U9056 ( .B1(n7366), .B2(n8027), .A(n7365), .ZN(P2_U3257) );
  INV_X1 U9057 ( .A(n7367), .ZN(n7372) );
  AOI21_X1 U9058 ( .B1(n7370), .B2(n7369), .A(n7368), .ZN(n7371) );
  OAI21_X1 U9059 ( .B1(n7372), .B2(n7371), .A(n8700), .ZN(n7376) );
  AND2_X1 U9060 ( .A1(P1_U3084), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n9527) );
  INV_X1 U9061 ( .A(n9596), .ZN(n7373) );
  OAI22_X1 U9062 ( .A1(n8707), .A2(n7373), .B1(n8705), .B2(n9588), .ZN(n7374)
         );
  AOI211_X1 U9063 ( .C1(n8710), .C2(n9012), .A(n9527), .B(n7374), .ZN(n7375)
         );
  OAI211_X1 U9064 ( .C1(n9663), .C2(n8713), .A(n7376), .B(n7375), .ZN(P1_U3229) );
  OAI222_X1 U9065 ( .A1(n8051), .A2(n7378), .B1(P2_U3152), .B2(n5506), .C1(
        n8049), .C2(n7377), .ZN(P2_U3338) );
  OAI222_X1 U9066 ( .A1(n8051), .A2(n9870), .B1(P2_U3152), .B2(n7380), .C1(
        n8049), .C2(n7379), .ZN(P2_U3337) );
  INV_X1 U9067 ( .A(n7381), .ZN(n7420) );
  AOI22_X1 U9068 ( .A1(n8997), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_22__SCAN_IN), .B2(n9383), .ZN(n7382) );
  OAI21_X1 U9069 ( .B1(n7420), .B2(n6951), .A(n7382), .ZN(P1_U3331) );
  NAND2_X1 U9070 ( .A1(n7384), .A2(n7383), .ZN(n7385) );
  XNOR2_X1 U9071 ( .A(n7386), .B(n7385), .ZN(n7392) );
  INV_X1 U9072 ( .A(n7504), .ZN(n7387) );
  OAI22_X1 U9073 ( .A1(n8707), .A2(n7387), .B1(n8705), .B2(n7498), .ZN(n7388)
         );
  AOI211_X1 U9074 ( .C1(n8710), .C2(n9011), .A(n7389), .B(n7388), .ZN(n7391)
         );
  NAND2_X1 U9075 ( .A1(n7505), .A2(n8680), .ZN(n7390) );
  OAI211_X1 U9076 ( .C1(n7392), .C2(n8682), .A(n7391), .B(n7390), .ZN(P1_U3215) );
  INV_X1 U9077 ( .A(n7570), .ZN(n10005) );
  OAI22_X1 U9078 ( .A1(n7564), .A2(n7393), .B1(P2_REG3_REG_3__SCAN_IN), .B2(
        n7461), .ZN(n7394) );
  AOI21_X1 U9079 ( .B1(n7395), .B2(n8450), .A(n7394), .ZN(n7396) );
  OAI21_X1 U9080 ( .B1(n7397), .B2(n8415), .A(n7396), .ZN(n7398) );
  AOI21_X1 U9081 ( .B1(n7399), .B2(n10005), .A(n7398), .ZN(n7400) );
  OAI21_X1 U9082 ( .B1(n7401), .B2(n10001), .A(n7400), .ZN(P2_U3293) );
  NAND2_X1 U9083 ( .A1(n7402), .A2(n7407), .ZN(n7403) );
  NAND2_X1 U9084 ( .A1(n7404), .A2(n7403), .ZN(n9742) );
  OR2_X1 U9085 ( .A1(n9742), .A2(n7563), .ZN(n7411) );
  OAI21_X1 U9086 ( .B1(n7407), .B2(n7406), .A(n7405), .ZN(n7409) );
  OAI22_X1 U9087 ( .A1(n8139), .A2(n9758), .B1(n8138), .B2(n9756), .ZN(n7408)
         );
  AOI21_X1 U9088 ( .B1(n7409), .B2(n9693), .A(n7408), .ZN(n7410) );
  NAND2_X1 U9089 ( .A1(n7411), .A2(n7410), .ZN(n9747) );
  NAND2_X1 U9090 ( .A1(n9747), .A2(n7564), .ZN(n7418) );
  AND2_X1 U9091 ( .A1(n7412), .A2(n8142), .ZN(n7413) );
  OR2_X1 U9092 ( .A1(n7413), .A2(n9764), .ZN(n9744) );
  INV_X1 U9093 ( .A(n9744), .ZN(n7416) );
  AOI22_X1 U9094 ( .A1(n10001), .A2(P2_REG2_REG_8__SCAN_IN), .B1(n8143), .B2(
        n9993), .ZN(n7414) );
  OAI21_X1 U9095 ( .B1(n8415), .B2(n9743), .A(n7414), .ZN(n7415) );
  AOI21_X1 U9096 ( .B1(n7416), .B2(n8450), .A(n7415), .ZN(n7417) );
  OAI211_X1 U9097 ( .C1(n9742), .C2(n7570), .A(n7418), .B(n7417), .ZN(P2_U3288) );
  OAI222_X1 U9098 ( .A1(n8051), .A2(n7421), .B1(n8049), .B2(n7420), .C1(n7419), 
        .C2(P2_U3152), .ZN(P2_U3336) );
  NAND2_X1 U9099 ( .A1(n7423), .A2(n7422), .ZN(n7424) );
  XNOR2_X1 U9100 ( .A(n7424), .B(n8839), .ZN(n9451) );
  INV_X1 U9101 ( .A(n9451), .ZN(n7433) );
  XNOR2_X1 U9102 ( .A(n7425), .B(n8839), .ZN(n7426) );
  OAI222_X1 U9103 ( .A1(n9586), .A2(n7698), .B1(n6241), .B2(n9587), .C1(n6240), 
        .C2(n7426), .ZN(n9449) );
  INV_X1 U9104 ( .A(n7503), .ZN(n7427) );
  INV_X1 U9105 ( .A(n7428), .ZN(n9447) );
  OAI21_X1 U9106 ( .B1(n7427), .B2(n9447), .A(n7489), .ZN(n9448) );
  AOI22_X1 U9107 ( .A1(n9597), .A2(P1_REG2_REG_11__SCAN_IN), .B1(n7546), .B2(
        n9595), .ZN(n7430) );
  NAND2_X1 U9108 ( .A1(n7428), .A2(n9605), .ZN(n7429) );
  OAI211_X1 U9109 ( .C1(n9448), .C2(n9066), .A(n7430), .B(n7429), .ZN(n7431)
         );
  AOI21_X1 U9110 ( .B1(n9449), .B2(n9609), .A(n7431), .ZN(n7432) );
  OAI21_X1 U9111 ( .B1(n7433), .B2(n9271), .A(n7432), .ZN(P1_U3280) );
  AOI22_X1 U9112 ( .A1(n10001), .A2(P2_REG2_REG_6__SCAN_IN), .B1(n7434), .B2(
        n9993), .ZN(n7435) );
  OAI21_X1 U9113 ( .B1(n8415), .B2(n7436), .A(n7435), .ZN(n7439) );
  NOR2_X1 U9114 ( .A1(n7437), .A2(n10001), .ZN(n7438) );
  AOI211_X1 U9115 ( .C1(n7440), .C2(n9702), .A(n7439), .B(n7438), .ZN(n7441)
         );
  OAI21_X1 U9116 ( .B1(n8452), .B2(n7442), .A(n7441), .ZN(P2_U3290) );
  NOR2_X1 U9117 ( .A1(n7444), .A2(n7443), .ZN(n7447) );
  INV_X1 U9118 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n7445) );
  AOI22_X1 U9119 ( .A1(n7475), .A2(n7445), .B1(P2_REG2_REG_13__SCAN_IN), .B2(
        n7448), .ZN(n7446) );
  NOR2_X1 U9120 ( .A1(n7447), .A2(n7446), .ZN(n7468) );
  AOI21_X1 U9121 ( .B1(n7447), .B2(n7446), .A(n7468), .ZN(n7458) );
  INV_X1 U9122 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n7455) );
  INV_X1 U9123 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n9419) );
  AOI22_X1 U9124 ( .A1(n7475), .A2(P2_REG1_REG_13__SCAN_IN), .B1(n9419), .B2(
        n7448), .ZN(n7452) );
  OAI21_X1 U9125 ( .B1(n7450), .B2(P2_REG1_REG_12__SCAN_IN), .A(n7449), .ZN(
        n7451) );
  NAND2_X1 U9126 ( .A1(n7452), .A2(n7451), .ZN(n7474) );
  OAI21_X1 U9127 ( .B1(n7452), .B2(n7451), .A(n7474), .ZN(n7453) );
  NAND2_X1 U9128 ( .A1(n9679), .A2(n7453), .ZN(n7454) );
  NAND2_X1 U9129 ( .A1(P2_U3152), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n7621) );
  OAI211_X1 U9130 ( .C1(n8033), .C2(n7455), .A(n7454), .B(n7621), .ZN(n7456)
         );
  AOI21_X1 U9131 ( .B1(n9684), .B2(n7475), .A(n7456), .ZN(n7457) );
  OAI21_X1 U9132 ( .B1(n7458), .B2(n8027), .A(n7457), .ZN(P2_U3258) );
  NAND2_X1 U9133 ( .A1(n9702), .A2(n7459), .ZN(n7460) );
  OAI21_X1 U9134 ( .B1(n9907), .B2(n7461), .A(n7460), .ZN(n7465) );
  OAI22_X1 U9135 ( .A1(n7463), .A2(n8452), .B1(n7462), .B2(n8415), .ZN(n7464)
         );
  AOI211_X1 U9136 ( .C1(n10001), .C2(P2_REG2_REG_1__SCAN_IN), .A(n7465), .B(
        n7464), .ZN(n7466) );
  OAI21_X1 U9137 ( .B1(n9706), .B2(n7467), .A(n7466), .ZN(P2_U3295) );
  NOR2_X1 U9138 ( .A1(n7475), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n7469) );
  NOR2_X1 U9139 ( .A1(n7469), .A2(n7468), .ZN(n7472) );
  INV_X1 U9140 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n7470) );
  AOI22_X1 U9141 ( .A1(n7768), .A2(n7470), .B1(P2_REG2_REG_14__SCAN_IN), .B2(
        n7473), .ZN(n7471) );
  NOR2_X1 U9142 ( .A1(n7472), .A2(n7471), .ZN(n7769) );
  AOI21_X1 U9143 ( .B1(n7472), .B2(n7471), .A(n7769), .ZN(n7483) );
  INV_X1 U9144 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n9412) );
  AOI22_X1 U9145 ( .A1(n7768), .A2(P2_REG1_REG_14__SCAN_IN), .B1(n9412), .B2(
        n7473), .ZN(n7477) );
  OAI21_X1 U9146 ( .B1(n7475), .B2(P2_REG1_REG_13__SCAN_IN), .A(n7474), .ZN(
        n7476) );
  NAND2_X1 U9147 ( .A1(n7477), .A2(n7476), .ZN(n7766) );
  OAI21_X1 U9148 ( .B1(n7477), .B2(n7476), .A(n7766), .ZN(n7478) );
  NAND2_X1 U9149 ( .A1(n7478), .A2(n9679), .ZN(n7482) );
  INV_X1 U9150 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n7479) );
  NAND2_X1 U9151 ( .A1(P2_U3152), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n7744) );
  OAI21_X1 U9152 ( .B1(n8033), .B2(n7479), .A(n7744), .ZN(n7480) );
  AOI21_X1 U9153 ( .B1(n9684), .B2(n7768), .A(n7480), .ZN(n7481) );
  OAI211_X1 U9154 ( .C1(n7483), .C2(n8027), .A(n7482), .B(n7481), .ZN(P2_U3259) );
  NAND2_X1 U9155 ( .A1(n7673), .A2(n7484), .ZN(n7485) );
  XNOR2_X1 U9156 ( .A(n7485), .B(n8840), .ZN(n9361) );
  XNOR2_X1 U9157 ( .A(n7486), .B(n8840), .ZN(n7487) );
  OAI222_X1 U9158 ( .A1(n9586), .A2(n8568), .B1(n6241), .B2(n7634), .C1(n7487), 
        .C2(n6240), .ZN(n9356) );
  INV_X1 U9159 ( .A(n9358), .ZN(n7493) );
  INV_X1 U9160 ( .A(n7683), .ZN(n7488) );
  AOI211_X1 U9161 ( .C1(n9358), .C2(n7489), .A(n9664), .B(n7488), .ZN(n9357)
         );
  NAND2_X1 U9162 ( .A1(n9357), .A2(n7490), .ZN(n7492) );
  AOI22_X1 U9163 ( .A1(n9597), .A2(P1_REG2_REG_12__SCAN_IN), .B1(n7633), .B2(
        n9595), .ZN(n7491) );
  OAI211_X1 U9164 ( .C1(n7493), .C2(n9599), .A(n7492), .B(n7491), .ZN(n7494)
         );
  AOI21_X1 U9165 ( .B1(n9356), .B2(n9609), .A(n7494), .ZN(n7495) );
  OAI21_X1 U9166 ( .B1(n9361), .B2(n9271), .A(n7495), .ZN(P1_U3279) );
  XOR2_X1 U9167 ( .A(n7496), .B(n8836), .Z(n7502) );
  XNOR2_X1 U9168 ( .A(n7497), .B(n8836), .ZN(n7500) );
  OAI22_X1 U9169 ( .A1(n7498), .A2(n6241), .B1(n7634), .B2(n9586), .ZN(n7499)
         );
  AOI21_X1 U9170 ( .B1(n7500), .B2(n9590), .A(n7499), .ZN(n7501) );
  OAI21_X1 U9171 ( .B1(n7502), .B2(n9593), .A(n7501), .ZN(n9396) );
  INV_X1 U9172 ( .A(n9396), .ZN(n7510) );
  INV_X1 U9173 ( .A(n7502), .ZN(n9398) );
  OAI211_X1 U9174 ( .C1(n9581), .C2(n9395), .A(n9340), .B(n7503), .ZN(n9394)
         );
  AOI22_X1 U9175 ( .A1(n9597), .A2(P1_REG2_REG_10__SCAN_IN), .B1(n7504), .B2(
        n9595), .ZN(n7507) );
  NAND2_X1 U9176 ( .A1(n7505), .A2(n9605), .ZN(n7506) );
  OAI211_X1 U9177 ( .C1(n9394), .C2(n9267), .A(n7507), .B(n7506), .ZN(n7508)
         );
  AOI21_X1 U9178 ( .B1(n9398), .B2(n9583), .A(n7508), .ZN(n7509) );
  OAI21_X1 U9179 ( .B1(n7510), .B2(n9597), .A(n7509), .ZN(P1_U3281) );
  INV_X1 U9180 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n10019) );
  NOR2_X1 U9181 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n7511) );
  AOI21_X1 U9182 ( .B1(P1_ADDR_REG_17__SCAN_IN), .B2(P2_ADDR_REG_17__SCAN_IN), 
        .A(n7511), .ZN(n9819) );
  NOR2_X1 U9183 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n7512) );
  AOI21_X1 U9184 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(P2_ADDR_REG_16__SCAN_IN), 
        .A(n7512), .ZN(n9822) );
  NOR2_X1 U9185 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n7513) );
  AOI21_X1 U9186 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(P2_ADDR_REG_15__SCAN_IN), 
        .A(n7513), .ZN(n9825) );
  NOR2_X1 U9187 ( .A1(P1_ADDR_REG_14__SCAN_IN), .A2(P2_ADDR_REG_14__SCAN_IN), 
        .ZN(n7514) );
  AOI21_X1 U9188 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(P1_ADDR_REG_14__SCAN_IN), 
        .A(n7514), .ZN(n9828) );
  NOR2_X1 U9189 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n7515) );
  AOI21_X1 U9190 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(P2_ADDR_REG_13__SCAN_IN), 
        .A(n7515), .ZN(n9831) );
  NOR2_X1 U9191 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n7522) );
  INV_X1 U9192 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n7516) );
  INV_X1 U9193 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n9947) );
  AOI22_X1 U9194 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(n7516), .B1(
        P2_ADDR_REG_4__SCAN_IN), .B2(n9947), .ZN(n10029) );
  NAND2_X1 U9195 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n7520) );
  XOR2_X1 U9196 ( .A(P1_ADDR_REG_3__SCAN_IN), .B(P2_ADDR_REG_3__SCAN_IN), .Z(
        n10027) );
  NAND2_X1 U9197 ( .A1(P2_ADDR_REG_2__SCAN_IN), .A2(P1_ADDR_REG_2__SCAN_IN), 
        .ZN(n7518) );
  XOR2_X1 U9198 ( .A(P2_ADDR_REG_2__SCAN_IN), .B(P1_ADDR_REG_2__SCAN_IN), .Z(
        n10025) );
  AOI21_X1 U9199 ( .B1(P1_ADDR_REG_0__SCAN_IN), .B2(P2_ADDR_REG_0__SCAN_IN), 
        .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n9811) );
  NAND3_X1 U9200 ( .A1(P2_ADDR_REG_0__SCAN_IN), .A2(P1_ADDR_REG_0__SCAN_IN), 
        .A3(P1_ADDR_REG_1__SCAN_IN), .ZN(n9813) );
  OAI21_X1 U9201 ( .B1(n9811), .B2(n9815), .A(n9813), .ZN(n10024) );
  NAND2_X1 U9202 ( .A1(n10025), .A2(n10024), .ZN(n7517) );
  NAND2_X1 U9203 ( .A1(n7518), .A2(n7517), .ZN(n10026) );
  NAND2_X1 U9204 ( .A1(n10027), .A2(n10026), .ZN(n7519) );
  NAND2_X1 U9205 ( .A1(n7520), .A2(n7519), .ZN(n10028) );
  NOR2_X1 U9206 ( .A1(n10029), .A2(n10028), .ZN(n7521) );
  NOR2_X1 U9207 ( .A1(n7522), .A2(n7521), .ZN(n7523) );
  NOR2_X1 U9208 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n7523), .ZN(n10013) );
  AND2_X1 U9209 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n7523), .ZN(n10014) );
  NOR2_X1 U9210 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n10014), .ZN(n7524) );
  NOR2_X1 U9211 ( .A1(n10013), .A2(n7524), .ZN(n7525) );
  NAND2_X1 U9212 ( .A1(n7525), .A2(P1_ADDR_REG_6__SCAN_IN), .ZN(n7527) );
  XOR2_X1 U9213 ( .A(n7525), .B(P1_ADDR_REG_6__SCAN_IN), .Z(n10012) );
  NAND2_X1 U9214 ( .A1(n10012), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n7526) );
  NAND2_X1 U9215 ( .A1(n7527), .A2(n7526), .ZN(n7528) );
  NAND2_X1 U9216 ( .A1(P1_ADDR_REG_7__SCAN_IN), .A2(n7528), .ZN(n7530) );
  INV_X1 U9217 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n9509) );
  XNOR2_X1 U9218 ( .A(n9509), .B(n7528), .ZN(n10016) );
  NAND2_X1 U9219 ( .A1(n10016), .A2(P2_ADDR_REG_7__SCAN_IN), .ZN(n7529) );
  NAND2_X1 U9220 ( .A1(n7530), .A2(n7529), .ZN(n7531) );
  NAND2_X1 U9221 ( .A1(P1_ADDR_REG_8__SCAN_IN), .A2(n7531), .ZN(n7533) );
  XOR2_X1 U9222 ( .A(P1_ADDR_REG_8__SCAN_IN), .B(n7531), .Z(n10011) );
  NAND2_X1 U9223 ( .A1(n10011), .A2(P2_ADDR_REG_8__SCAN_IN), .ZN(n7532) );
  NAND2_X1 U9224 ( .A1(n7533), .A2(n7532), .ZN(n7534) );
  AND2_X1 U9225 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(n7534), .ZN(n7535) );
  INV_X1 U9226 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n10023) );
  XNOR2_X1 U9227 ( .A(P2_ADDR_REG_9__SCAN_IN), .B(n7534), .ZN(n10022) );
  NOR2_X1 U9228 ( .A1(n10023), .A2(n10022), .ZN(n10021) );
  NAND2_X1 U9229 ( .A1(P1_ADDR_REG_10__SCAN_IN), .A2(P2_ADDR_REG_10__SCAN_IN), 
        .ZN(n7536) );
  OAI21_X1 U9230 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(P2_ADDR_REG_10__SCAN_IN), 
        .A(n7536), .ZN(n9839) );
  NAND2_X1 U9231 ( .A1(P1_ADDR_REG_11__SCAN_IN), .A2(P2_ADDR_REG_11__SCAN_IN), 
        .ZN(n7537) );
  OAI21_X1 U9232 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(P2_ADDR_REG_11__SCAN_IN), 
        .A(n7537), .ZN(n9836) );
  NOR2_X1 U9233 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n7538) );
  AOI21_X1 U9234 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(P2_ADDR_REG_12__SCAN_IN), 
        .A(n7538), .ZN(n9833) );
  NAND2_X1 U9235 ( .A1(n9834), .A2(n9833), .ZN(n9832) );
  NAND2_X1 U9236 ( .A1(n9831), .A2(n9830), .ZN(n9829) );
  OAI21_X1 U9237 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(P1_ADDR_REG_13__SCAN_IN), 
        .A(n9829), .ZN(n9827) );
  NAND2_X1 U9238 ( .A1(n9828), .A2(n9827), .ZN(n9826) );
  OAI21_X1 U9239 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(P2_ADDR_REG_14__SCAN_IN), 
        .A(n9826), .ZN(n9824) );
  NAND2_X1 U9240 ( .A1(n9825), .A2(n9824), .ZN(n9823) );
  OAI21_X1 U9241 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(P1_ADDR_REG_15__SCAN_IN), 
        .A(n9823), .ZN(n9821) );
  NAND2_X1 U9242 ( .A1(n9822), .A2(n9821), .ZN(n9820) );
  OAI21_X1 U9243 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(P1_ADDR_REG_16__SCAN_IN), 
        .A(n9820), .ZN(n9818) );
  NAND2_X1 U9244 ( .A1(n9819), .A2(n9818), .ZN(n9817) );
  OAI21_X1 U9245 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(P1_ADDR_REG_17__SCAN_IN), 
        .A(n9817), .ZN(n10018) );
  NOR2_X1 U9246 ( .A1(n10019), .A2(n10018), .ZN(n7539) );
  NAND2_X1 U9247 ( .A1(n10019), .A2(n10018), .ZN(n10017) );
  OAI21_X1 U9248 ( .B1(P1_ADDR_REG_18__SCAN_IN), .B2(n7539), .A(n10017), .ZN(
        n7541) );
  XNOR2_X1 U9249 ( .A(n4761), .B(P2_ADDR_REG_19__SCAN_IN), .ZN(n7540) );
  XNOR2_X1 U9250 ( .A(n7541), .B(n7540), .ZN(ADD_1071_U4) );
  AOI21_X1 U9251 ( .B1(n7543), .B2(n7542), .A(n8682), .ZN(n7545) );
  NAND2_X1 U9252 ( .A1(n7545), .A2(n7544), .ZN(n7550) );
  NOR2_X1 U9253 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6033), .ZN(n9535) );
  INV_X1 U9254 ( .A(n7546), .ZN(n7547) );
  OAI22_X1 U9255 ( .A1(n8707), .A2(n7547), .B1(n8705), .B2(n9587), .ZN(n7548)
         );
  AOI211_X1 U9256 ( .C1(n8710), .C2(n9010), .A(n9535), .B(n7548), .ZN(n7549)
         );
  OAI211_X1 U9257 ( .C1(n9447), .C2(n8713), .A(n7550), .B(n7549), .ZN(P1_U3234) );
  INV_X1 U9258 ( .A(n8112), .ZN(n8238) );
  NAND2_X1 U9259 ( .A1(n8208), .A2(n8238), .ZN(n7551) );
  INV_X1 U9260 ( .A(n8204), .ZN(n8237) );
  OR2_X1 U9261 ( .A1(n9786), .A2(n8237), .ZN(n7554) );
  INV_X1 U9262 ( .A(n7558), .ZN(n7555) );
  NAND2_X1 U9263 ( .A1(n7556), .A2(n7558), .ZN(n7557) );
  NAND2_X1 U9264 ( .A1(n7578), .A2(n7557), .ZN(n9413) );
  XNOR2_X1 U9265 ( .A(n7559), .B(n7558), .ZN(n7561) );
  OAI22_X1 U9266 ( .A1(n8204), .A2(n9758), .B1(n7818), .B2(n9756), .ZN(n7560)
         );
  AOI21_X1 U9267 ( .B1(n7561), .B2(n9693), .A(n7560), .ZN(n7562) );
  OAI21_X1 U9268 ( .B1(n9413), .B2(n7563), .A(n7562), .ZN(n9416) );
  NAND2_X1 U9269 ( .A1(n9416), .A2(n7564), .ZN(n7569) );
  XNOR2_X1 U9270 ( .A(n9699), .B(n7587), .ZN(n9415) );
  INV_X1 U9271 ( .A(n9415), .ZN(n7567) );
  INV_X1 U9272 ( .A(n7587), .ZN(n9414) );
  AOI22_X1 U9273 ( .A1(n9706), .A2(P2_REG2_REG_13__SCAN_IN), .B1(n7625), .B2(
        n9993), .ZN(n7565) );
  OAI21_X1 U9274 ( .B1(n9414), .B2(n8415), .A(n7565), .ZN(n7566) );
  AOI21_X1 U9275 ( .B1(n7567), .B2(n8450), .A(n7566), .ZN(n7568) );
  OAI211_X1 U9276 ( .C1(n9413), .C2(n7570), .A(n7569), .B(n7568), .ZN(P2_U3283) );
  INV_X1 U9277 ( .A(n7571), .ZN(n7576) );
  OR2_X1 U9278 ( .A1(n7572), .A2(P1_U3084), .ZN(n8996) );
  INV_X1 U9279 ( .A(n8996), .ZN(n8988) );
  AOI21_X1 U9280 ( .B1(P2_DATAO_REG_23__SCAN_IN), .B2(n9383), .A(n8988), .ZN(
        n7573) );
  OAI21_X1 U9281 ( .B1(n7576), .B2(n6951), .A(n7573), .ZN(P1_U3330) );
  NAND2_X1 U9282 ( .A1(n8556), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n7574) );
  OAI211_X1 U9283 ( .C1(n7576), .C2(n8049), .A(n7575), .B(n7574), .ZN(P2_U3335) );
  INV_X1 U9284 ( .A(n7746), .ZN(n8236) );
  NAND2_X1 U9285 ( .A1(n7587), .A2(n8236), .ZN(n7577) );
  OAI21_X1 U9286 ( .B1(n7580), .B2(n7579), .A(n7659), .ZN(n9411) );
  INV_X1 U9287 ( .A(n9411), .ZN(n7593) );
  INV_X1 U9288 ( .A(n7581), .ZN(n7584) );
  OAI211_X1 U9289 ( .C1(n7584), .C2(n7583), .A(n7582), .B(n9693), .ZN(n7586)
         );
  AOI22_X1 U9290 ( .A1(n8445), .A2(n8234), .B1(n8236), .B2(n8443), .ZN(n7585)
         );
  NAND2_X1 U9291 ( .A1(n7586), .A2(n7585), .ZN(n9410) );
  INV_X1 U9292 ( .A(n7657), .ZN(n9407) );
  NAND2_X1 U9293 ( .A1(n7588), .A2(n9407), .ZN(n7665) );
  OAI21_X1 U9294 ( .B1(n7588), .B2(n9407), .A(n7665), .ZN(n9408) );
  AOI22_X1 U9295 ( .A1(n9706), .A2(P2_REG2_REG_14__SCAN_IN), .B1(n7749), .B2(
        n9993), .ZN(n7590) );
  NAND2_X1 U9296 ( .A1(n7657), .A2(n9996), .ZN(n7589) );
  OAI211_X1 U9297 ( .C1(n9408), .C2(n9999), .A(n7590), .B(n7589), .ZN(n7591)
         );
  AOI21_X1 U9298 ( .B1(n9410), .B2(n7564), .A(n7591), .ZN(n7592) );
  OAI21_X1 U9299 ( .B1(n7593), .B2(n8452), .A(n7592), .ZN(P2_U3282) );
  NOR2_X1 U9300 ( .A1(n7595), .A2(n7599), .ZN(n7596) );
  INV_X1 U9301 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n9550) );
  NOR2_X1 U9302 ( .A1(n9550), .A2(n9551), .ZN(n9549) );
  NOR2_X1 U9303 ( .A1(n7596), .A2(n9549), .ZN(n7704) );
  INV_X1 U9304 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n7597) );
  AOI211_X1 U9305 ( .C1(n7598), .C2(n7597), .A(n7705), .B(n9563), .ZN(n7607)
         );
  INV_X1 U9306 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n9439) );
  AOI22_X1 U9307 ( .A1(n9554), .A2(P1_REG1_REG_14__SCAN_IN), .B1(n9439), .B2(
        n7599), .ZN(n9556) );
  NAND2_X1 U9308 ( .A1(n9556), .A2(n9557), .ZN(n9555) );
  XNOR2_X1 U9309 ( .A(n7709), .B(n7710), .ZN(n7603) );
  INV_X1 U9310 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n7602) );
  NOR2_X1 U9311 ( .A1(n7602), .A2(n7603), .ZN(n7711) );
  AOI211_X1 U9312 ( .C1(n7603), .C2(n7602), .A(n7711), .B(n9510), .ZN(n7606)
         );
  NAND2_X1 U9313 ( .A1(n9573), .A2(P1_ADDR_REG_15__SCAN_IN), .ZN(n7604) );
  NAND2_X1 U9314 ( .A1(P1_U3084), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n8702) );
  OAI211_X1 U9315 ( .C1(n9045), .C2(n7710), .A(n7604), .B(n8702), .ZN(n7605)
         );
  OR3_X1 U9316 ( .A1(n7607), .A2(n7606), .A3(n7605), .ZN(P1_U3256) );
  INV_X1 U9317 ( .A(n9695), .ZN(n7611) );
  OR2_X1 U9318 ( .A1(n8112), .A2(n9758), .ZN(n7608) );
  OAI21_X1 U9319 ( .B1(n7746), .B2(n9756), .A(n7608), .ZN(n9692) );
  NAND2_X1 U9320 ( .A1(n9692), .A2(n8175), .ZN(n7610) );
  OAI211_X1 U9321 ( .C1(n8177), .C2(n7611), .A(n7610), .B(n7609), .ZN(n7617)
         );
  NAND2_X1 U9322 ( .A1(n7613), .A2(n7612), .ZN(n7614) );
  AOI21_X1 U9323 ( .B1(n7615), .B2(n7614), .A(n8189), .ZN(n7616) );
  AOI211_X1 U9324 ( .C1(n9786), .C2(n8207), .A(n7617), .B(n7616), .ZN(n7618)
         );
  INV_X1 U9325 ( .A(n7618), .ZN(P2_U3226) );
  XNOR2_X1 U9326 ( .A(n7620), .B(n7619), .ZN(n7627) );
  INV_X1 U9327 ( .A(n7818), .ZN(n8235) );
  NAND2_X1 U9328 ( .A1(n8235), .A2(n8195), .ZN(n7622) );
  OAI211_X1 U9329 ( .C1(n8204), .C2(n8220), .A(n7622), .B(n7621), .ZN(n7624)
         );
  NOR2_X1 U9330 ( .A1(n9414), .A2(n8227), .ZN(n7623) );
  AOI211_X1 U9331 ( .C1(n8224), .C2(n7625), .A(n7624), .B(n7623), .ZN(n7626)
         );
  OAI21_X1 U9332 ( .B1(n7627), .B2(n8189), .A(n7626), .ZN(P2_U3236) );
  XNOR2_X1 U9333 ( .A(n7630), .B(n7629), .ZN(n7631) );
  XNOR2_X1 U9334 ( .A(n7628), .B(n7631), .ZN(n7640) );
  INV_X1 U9335 ( .A(n7632), .ZN(n7637) );
  INV_X1 U9336 ( .A(n7633), .ZN(n7635) );
  OAI22_X1 U9337 ( .A1(n8707), .A2(n7635), .B1(n8705), .B2(n7634), .ZN(n7636)
         );
  AOI211_X1 U9338 ( .C1(n8710), .C2(n9009), .A(n7637), .B(n7636), .ZN(n7639)
         );
  NAND2_X1 U9339 ( .A1(n9358), .A2(n8680), .ZN(n7638) );
  OAI211_X1 U9340 ( .C1(n7640), .C2(n8682), .A(n7639), .B(n7638), .ZN(P1_U3222) );
  INV_X1 U9341 ( .A(n7641), .ZN(n7655) );
  AOI22_X1 U9342 ( .A1(n7642), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_24__SCAN_IN), .B2(n9383), .ZN(n7643) );
  OAI21_X1 U9343 ( .B1(n7655), .B2(n6951), .A(n7643), .ZN(P1_U3329) );
  XNOR2_X1 U9344 ( .A(n7644), .B(n8844), .ZN(n9438) );
  INV_X1 U9345 ( .A(n9438), .ZN(n7653) );
  OR2_X1 U9346 ( .A1(n9254), .A2(n8844), .ZN(n7728) );
  NAND2_X1 U9347 ( .A1(n9254), .A2(n8844), .ZN(n7645) );
  NAND3_X1 U9348 ( .A1(n7728), .A2(n9590), .A3(n7645), .ZN(n7647) );
  INV_X1 U9349 ( .A(n9260), .ZN(n9007) );
  AOI22_X1 U9350 ( .A1(n9007), .A2(n9231), .B1(n9233), .B2(n9009), .ZN(n7646)
         );
  NAND2_X1 U9351 ( .A1(n7647), .A2(n7646), .ZN(n9437) );
  OAI211_X1 U9352 ( .C1(n7684), .C2(n9435), .A(n4344), .B(n9340), .ZN(n9434)
         );
  AOI22_X1 U9353 ( .A1(n9597), .A2(P1_REG2_REG_14__SCAN_IN), .B1(n8567), .B2(
        n9595), .ZN(n7650) );
  NAND2_X1 U9354 ( .A1(n7648), .A2(n9605), .ZN(n7649) );
  OAI211_X1 U9355 ( .C1(n9434), .C2(n9267), .A(n7650), .B(n7649), .ZN(n7651)
         );
  AOI21_X1 U9356 ( .B1(n9437), .B2(n9609), .A(n7651), .ZN(n7652) );
  OAI21_X1 U9357 ( .B1(n7653), .B2(n9271), .A(n7652), .ZN(P1_U3277) );
  OAI222_X1 U9358 ( .A1(P2_U3152), .A2(n7656), .B1(n8049), .B2(n7655), .C1(
        n7654), .C2(n8051), .ZN(P2_U3334) );
  OR2_X1 U9359 ( .A1(n7657), .A2(n8235), .ZN(n7658) );
  XNOR2_X1 U9360 ( .A(n7758), .B(n7757), .ZN(n9405) );
  INV_X1 U9361 ( .A(n9405), .ZN(n7671) );
  OAI211_X1 U9362 ( .C1(n7662), .C2(n7661), .A(n7660), .B(n9693), .ZN(n7664)
         );
  AOI22_X1 U9363 ( .A1(n8235), .A2(n8443), .B1(n8445), .B2(n8233), .ZN(n7663)
         );
  NAND2_X1 U9364 ( .A1(n7664), .A2(n7663), .ZN(n9404) );
  INV_X1 U9365 ( .A(n7665), .ZN(n7666) );
  OAI21_X1 U9366 ( .B1(n7666), .B2(n9401), .A(n4342), .ZN(n9402) );
  AOI22_X1 U9367 ( .A1(n9706), .A2(P2_REG2_REG_15__SCAN_IN), .B1(n7815), .B2(
        n9993), .ZN(n7668) );
  NAND2_X1 U9368 ( .A1(n7820), .A2(n9996), .ZN(n7667) );
  OAI211_X1 U9369 ( .C1(n9402), .C2(n9999), .A(n7668), .B(n7667), .ZN(n7669)
         );
  AOI21_X1 U9370 ( .B1(n9404), .B2(n7564), .A(n7669), .ZN(n7670) );
  OAI21_X1 U9371 ( .B1(n7671), .B2(n8452), .A(n7670), .ZN(P2_U3281) );
  NAND2_X1 U9372 ( .A1(n7673), .A2(n7672), .ZN(n7675) );
  AND2_X1 U9373 ( .A1(n7675), .A2(n7674), .ZN(n7676) );
  XOR2_X1 U9374 ( .A(n8842), .B(n7676), .Z(n9441) );
  INV_X1 U9375 ( .A(n9583), .ZN(n7690) );
  XNOR2_X1 U9376 ( .A(n7677), .B(n8842), .ZN(n7679) );
  OAI22_X1 U9377 ( .A1(n8704), .A2(n9586), .B1(n7698), .B2(n6241), .ZN(n7678)
         );
  AOI21_X1 U9378 ( .B1(n7679), .B2(n9590), .A(n7678), .ZN(n7680) );
  OAI21_X1 U9379 ( .B1(n9441), .B2(n9593), .A(n7680), .ZN(n9444) );
  NAND2_X1 U9380 ( .A1(n9444), .A2(n9609), .ZN(n7689) );
  INV_X1 U9381 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n7682) );
  INV_X1 U9382 ( .A(n7681), .ZN(n7699) );
  OAI22_X1 U9383 ( .A1(n9609), .A2(n7682), .B1(n7699), .B2(n9613), .ZN(n7687)
         );
  AND2_X1 U9384 ( .A1(n7683), .A2(n7691), .ZN(n7685) );
  OR2_X1 U9385 ( .A1(n7685), .A2(n7684), .ZN(n9443) );
  NOR2_X1 U9386 ( .A1(n9443), .A2(n9066), .ZN(n7686) );
  AOI211_X1 U9387 ( .C1(n9605), .C2(n7691), .A(n7687), .B(n7686), .ZN(n7688)
         );
  OAI211_X1 U9388 ( .C1(n9441), .C2(n7690), .A(n7689), .B(n7688), .ZN(P1_U3278) );
  INV_X1 U9389 ( .A(n7691), .ZN(n9442) );
  OAI21_X1 U9390 ( .B1(n4353), .B2(n7693), .A(n7692), .ZN(n7694) );
  OAI21_X1 U9391 ( .B1(n7695), .B2(n4353), .A(n7694), .ZN(n7696) );
  NAND2_X1 U9392 ( .A1(n7696), .A2(n8700), .ZN(n7703) );
  INV_X1 U9393 ( .A(n7697), .ZN(n7701) );
  OAI22_X1 U9394 ( .A1(n8707), .A2(n7699), .B1(n8705), .B2(n7698), .ZN(n7700)
         );
  AOI211_X1 U9395 ( .C1(n8710), .C2(n9008), .A(n7701), .B(n7700), .ZN(n7702)
         );
  OAI211_X1 U9396 ( .C1(n9442), .C2(n8713), .A(n7703), .B(n7702), .ZN(P1_U3232) );
  NOR2_X1 U9397 ( .A1(n7704), .A2(n7710), .ZN(n7706) );
  NAND2_X1 U9398 ( .A1(P1_REG2_REG_16__SCAN_IN), .A2(n9027), .ZN(n7707) );
  OAI21_X1 U9399 ( .B1(n9027), .B2(P1_REG2_REG_16__SCAN_IN), .A(n7707), .ZN(
        n7708) );
  AOI211_X1 U9400 ( .C1(n4346), .C2(n7708), .A(n9022), .B(n9563), .ZN(n7721)
         );
  NOR2_X1 U9401 ( .A1(n7710), .A2(n7709), .ZN(n7712) );
  INV_X1 U9402 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n9433) );
  NOR2_X1 U9403 ( .A1(n9027), .A2(n9433), .ZN(n7713) );
  AOI21_X1 U9404 ( .B1(n9027), .B2(n9433), .A(n7713), .ZN(n7714) );
  NOR2_X1 U9405 ( .A1(n7715), .A2(n7714), .ZN(n9026) );
  AOI211_X1 U9406 ( .C1(n7715), .C2(n7714), .A(n9026), .B(n9510), .ZN(n7720)
         );
  NAND2_X1 U9407 ( .A1(n9573), .A2(P1_ADDR_REG_16__SCAN_IN), .ZN(n7717) );
  NAND2_X1 U9408 ( .A1(P1_REG3_REG_16__SCAN_IN), .A2(P1_U3084), .ZN(n7716) );
  OAI211_X1 U9409 ( .C1(n9045), .C2(n7718), .A(n7717), .B(n7716), .ZN(n7719)
         );
  OR3_X1 U9410 ( .A1(n7721), .A2(n7720), .A3(n7719), .ZN(P1_U3257) );
  INV_X1 U9411 ( .A(n7722), .ZN(n7764) );
  AOI22_X1 U9412 ( .A1(n7723), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_25__SCAN_IN), .B2(n9389), .ZN(n7724) );
  OAI21_X1 U9413 ( .B1(n7764), .B2(n6951), .A(n7724), .ZN(P1_U3328) );
  XNOR2_X1 U9414 ( .A(n7725), .B(n8846), .ZN(n9350) );
  NAND2_X1 U9415 ( .A1(n9350), .A2(n7726), .ZN(n7735) );
  AND2_X1 U9416 ( .A1(n7728), .A2(n8763), .ZN(n7730) );
  NAND2_X1 U9417 ( .A1(n7728), .A2(n7727), .ZN(n7729) );
  OAI21_X1 U9418 ( .B1(n7730), .B2(n8846), .A(n7729), .ZN(n7733) );
  NAND2_X1 U9419 ( .A1(n9008), .A2(n9233), .ZN(n7731) );
  OAI21_X1 U9420 ( .B1(n9243), .B2(n9586), .A(n7731), .ZN(n7732) );
  AOI21_X1 U9421 ( .B1(n7733), .B2(n9590), .A(n7732), .ZN(n7734) );
  NAND2_X1 U9422 ( .A1(n7735), .A2(n7734), .ZN(n9354) );
  INV_X1 U9423 ( .A(n9354), .ZN(n7741) );
  NAND2_X1 U9424 ( .A1(n4344), .A2(n8695), .ZN(n7736) );
  NAND2_X1 U9425 ( .A1(n9261), .A2(n7736), .ZN(n9352) );
  AOI22_X1 U9426 ( .A1(n9597), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n8703), .B2(
        n9595), .ZN(n7738) );
  NAND2_X1 U9427 ( .A1(n8695), .A2(n9605), .ZN(n7737) );
  OAI211_X1 U9428 ( .C1(n9352), .C2(n9066), .A(n7738), .B(n7737), .ZN(n7739)
         );
  AOI21_X1 U9429 ( .B1(n9350), .B2(n9583), .A(n7739), .ZN(n7740) );
  OAI21_X1 U9430 ( .B1(n7741), .B2(n9597), .A(n7740), .ZN(P1_U3276) );
  AOI21_X1 U9431 ( .B1(n7743), .B2(n7742), .A(n4347), .ZN(n7751) );
  NAND2_X1 U9432 ( .A1(n8234), .A2(n8195), .ZN(n7745) );
  OAI211_X1 U9433 ( .C1(n7746), .C2(n8220), .A(n7745), .B(n7744), .ZN(n7748)
         );
  NOR2_X1 U9434 ( .A1(n9407), .A2(n8227), .ZN(n7747) );
  AOI211_X1 U9435 ( .C1(n8224), .C2(n7749), .A(n7748), .B(n7747), .ZN(n7750)
         );
  OAI21_X1 U9436 ( .B1(n7751), .B2(n8189), .A(n7750), .ZN(P2_U3217) );
  XNOR2_X1 U9437 ( .A(n7752), .B(n7759), .ZN(n7753) );
  AOI222_X1 U9438 ( .A1(n9693), .A2(n7753), .B1(n8444), .B2(n8445), .C1(n8234), 
        .C2(n8443), .ZN(n8533) );
  XOR2_X1 U9439 ( .A(n8530), .B(n4342), .Z(n8531) );
  INV_X1 U9440 ( .A(n8530), .ZN(n7755) );
  AOI22_X1 U9441 ( .A1(n10001), .A2(P2_REG2_REG_16__SCAN_IN), .B1(n7842), .B2(
        n9993), .ZN(n7754) );
  OAI21_X1 U9442 ( .B1(n7755), .B2(n8415), .A(n7754), .ZN(n7756) );
  AOI21_X1 U9443 ( .B1(n8531), .B2(n8450), .A(n7756), .ZN(n7762) );
  OR2_X1 U9444 ( .A1(n7760), .A2(n7759), .ZN(n8529) );
  NAND2_X1 U9445 ( .A1(n7760), .A2(n7759), .ZN(n7784) );
  INV_X1 U9446 ( .A(n8452), .ZN(n9703) );
  NAND3_X1 U9447 ( .A1(n8529), .A2(n7784), .A3(n9703), .ZN(n7761) );
  OAI211_X1 U9448 ( .C1(n8533), .C2(n9706), .A(n7762), .B(n7761), .ZN(P2_U3280) );
  OAI222_X1 U9449 ( .A1(n8051), .A2(n7765), .B1(n8049), .B2(n7764), .C1(
        P2_U3152), .C2(n7763), .ZN(P2_U3333) );
  OAI21_X1 U9450 ( .B1(n7768), .B2(P2_REG1_REG_14__SCAN_IN), .A(n7766), .ZN(
        n7871) );
  XNOR2_X1 U9451 ( .A(n7871), .B(n7872), .ZN(n7767) );
  INV_X1 U9452 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n9406) );
  NOR2_X1 U9453 ( .A1(n9406), .A2(n7767), .ZN(n7873) );
  AOI211_X1 U9454 ( .C1(n7767), .C2(n9406), .A(n7873), .B(n9682), .ZN(n7777)
         );
  NOR2_X1 U9455 ( .A1(n7768), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n7770) );
  NOR2_X1 U9456 ( .A1(n7770), .A2(n7769), .ZN(n7863) );
  XNOR2_X1 U9457 ( .A(n7863), .B(n7864), .ZN(n7771) );
  NOR2_X1 U9458 ( .A1(P2_REG2_REG_15__SCAN_IN), .A2(n7771), .ZN(n7865) );
  AOI21_X1 U9459 ( .B1(n7771), .B2(P2_REG2_REG_15__SCAN_IN), .A(n7865), .ZN(
        n7772) );
  NOR2_X1 U9460 ( .A1(n7772), .A2(n8027), .ZN(n7776) );
  AND2_X1 U9461 ( .A1(P2_U3152), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n7773) );
  AOI21_X1 U9462 ( .B1(n9681), .B2(P2_ADDR_REG_15__SCAN_IN), .A(n7773), .ZN(
        n7774) );
  OAI21_X1 U9463 ( .B1(n8030), .B2(n7872), .A(n7774), .ZN(n7775) );
  OR3_X1 U9464 ( .A1(n7777), .A2(n7776), .A3(n7775), .ZN(P2_U3260) );
  INV_X1 U9465 ( .A(n7778), .ZN(n7782) );
  AOI22_X1 U9466 ( .A1(n7779), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_26__SCAN_IN), .B2(n8556), .ZN(n7780) );
  OAI21_X1 U9467 ( .B1(n7782), .B2(n8049), .A(n7780), .ZN(P2_U3332) );
  AOI22_X1 U9468 ( .A1(n6251), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_26__SCAN_IN), .B2(n9389), .ZN(n7781) );
  OAI21_X1 U9469 ( .B1(n7782), .B2(n6951), .A(n7781), .ZN(P1_U3327) );
  INV_X1 U9470 ( .A(n7789), .ZN(n7785) );
  INV_X1 U9471 ( .A(n8053), .ZN(n7786) );
  AOI21_X1 U9472 ( .B1(n7789), .B2(n7787), .A(n7786), .ZN(n8528) );
  XNOR2_X1 U9473 ( .A(n7788), .B(n7789), .ZN(n7790) );
  OAI222_X1 U9474 ( .A1(n9756), .A2(n8127), .B1(n9758), .B2(n7801), .C1(n9753), 
        .C2(n7790), .ZN(n8524) );
  INV_X1 U9475 ( .A(n8526), .ZN(n7793) );
  AOI211_X1 U9476 ( .C1(n8526), .C2(n4345), .A(n9780), .B(n8436), .ZN(n8525)
         );
  NAND2_X1 U9477 ( .A1(n8525), .A2(n9702), .ZN(n7792) );
  AOI22_X1 U9478 ( .A1(n10001), .A2(P2_REG2_REG_17__SCAN_IN), .B1(n7798), .B2(
        n9993), .ZN(n7791) );
  OAI211_X1 U9479 ( .C1(n7793), .C2(n8415), .A(n7792), .B(n7791), .ZN(n7794)
         );
  AOI21_X1 U9480 ( .B1(n8524), .B2(n7564), .A(n7794), .ZN(n7795) );
  OAI21_X1 U9481 ( .B1(n8528), .B2(n8452), .A(n7795), .ZN(P2_U3279) );
  XNOR2_X1 U9482 ( .A(n7797), .B(n7796), .ZN(n7804) );
  AOI22_X1 U9483 ( .A1(n8195), .A2(n8425), .B1(P2_REG3_REG_17__SCAN_IN), .B2(
        P2_U3152), .ZN(n7800) );
  NAND2_X1 U9484 ( .A1(n8224), .A2(n7798), .ZN(n7799) );
  OAI211_X1 U9485 ( .C1(n7801), .C2(n8220), .A(n7800), .B(n7799), .ZN(n7802)
         );
  AOI21_X1 U9486 ( .B1(n8526), .B2(n8207), .A(n7802), .ZN(n7803) );
  OAI21_X1 U9487 ( .B1(n7804), .B2(n8189), .A(n7803), .ZN(P2_U3230) );
  INV_X1 U9488 ( .A(n7805), .ZN(n7809) );
  AOI21_X1 U9489 ( .B1(n9389), .B2(P2_DATAO_REG_27__SCAN_IN), .A(n7806), .ZN(
        n7807) );
  OAI21_X1 U9490 ( .B1(n7809), .B2(n6951), .A(n7807), .ZN(P1_U3326) );
  AOI22_X1 U9491 ( .A1(n8072), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_27__SCAN_IN), .B2(n8556), .ZN(n7808) );
  OAI21_X1 U9492 ( .B1(n7809), .B2(n8049), .A(n7808), .ZN(P2_U3331) );
  NOR2_X1 U9493 ( .A1(n7811), .A2(n7810), .ZN(n7834) );
  INV_X1 U9494 ( .A(n7834), .ZN(n7812) );
  NAND2_X1 U9495 ( .A1(n7811), .A2(n7810), .ZN(n7832) );
  NAND2_X1 U9496 ( .A1(n7812), .A2(n7832), .ZN(n7814) );
  XNOR2_X1 U9497 ( .A(n7814), .B(n7813), .ZN(n7822) );
  AOI22_X1 U9498 ( .A1(n8195), .A2(n8233), .B1(P2_REG3_REG_15__SCAN_IN), .B2(
        P2_U3152), .ZN(n7817) );
  NAND2_X1 U9499 ( .A1(n8224), .A2(n7815), .ZN(n7816) );
  OAI211_X1 U9500 ( .C1(n7818), .C2(n8220), .A(n7817), .B(n7816), .ZN(n7819)
         );
  AOI21_X1 U9501 ( .B1(n7820), .B2(n8207), .A(n7819), .ZN(n7821) );
  OAI21_X1 U9502 ( .B1(n7822), .B2(n8189), .A(n7821), .ZN(P2_U3243) );
  XNOR2_X1 U9503 ( .A(n7824), .B(n7823), .ZN(n7831) );
  NOR2_X1 U9504 ( .A1(n7825), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7877) );
  AOI21_X1 U9505 ( .B1(n8195), .B2(n8446), .A(n7877), .ZN(n7827) );
  NAND2_X1 U9506 ( .A1(n8224), .A2(n8439), .ZN(n7826) );
  OAI211_X1 U9507 ( .C1(n7828), .C2(n8220), .A(n7827), .B(n7826), .ZN(n7829)
         );
  AOI21_X1 U9508 ( .B1(n8519), .B2(n8207), .A(n7829), .ZN(n7830) );
  OAI21_X1 U9509 ( .B1(n7831), .B2(n8189), .A(n7830), .ZN(P2_U3240) );
  OAI21_X1 U9510 ( .B1(n7834), .B2(n7833), .A(n7832), .ZN(n7838) );
  NAND2_X1 U9511 ( .A1(n7836), .A2(n7835), .ZN(n7837) );
  XNOR2_X1 U9512 ( .A(n7838), .B(n7837), .ZN(n7845) );
  NAND2_X1 U9513 ( .A1(n8444), .A2(n8195), .ZN(n7839) );
  NAND2_X1 U9514 ( .A1(P2_REG3_REG_16__SCAN_IN), .A2(P2_U3152), .ZN(n8253) );
  OAI211_X1 U9515 ( .C1(n7840), .C2(n8220), .A(n7839), .B(n8253), .ZN(n7841)
         );
  AOI21_X1 U9516 ( .B1(n7842), .B2(n8224), .A(n7841), .ZN(n7844) );
  NAND2_X1 U9517 ( .A1(n8530), .A2(n8207), .ZN(n7843) );
  OAI211_X1 U9518 ( .C1(n7845), .C2(n8189), .A(n7844), .B(n7843), .ZN(P2_U3228) );
  INV_X1 U9519 ( .A(n7846), .ZN(n7851) );
  AOI21_X1 U9520 ( .B1(n9389), .B2(P2_DATAO_REG_28__SCAN_IN), .A(n7847), .ZN(
        n7848) );
  OAI21_X1 U9521 ( .B1(n7851), .B2(n6951), .A(n7848), .ZN(P1_U3325) );
  AOI22_X1 U9522 ( .A1(n7849), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_28__SCAN_IN), .B2(n8556), .ZN(n7850) );
  OAI21_X1 U9523 ( .B1(n7851), .B2(n8049), .A(n7850), .ZN(P2_U3330) );
  MUX2_X1 U9524 ( .A(n7852), .B(P1_REG2_REG_2__SCAN_IN), .S(n9597), .Z(n7858)
         );
  NAND2_X1 U9525 ( .A1(n7853), .A2(n9583), .ZN(n7855) );
  AOI22_X1 U9526 ( .A1(n9605), .A2(n8666), .B1(n9595), .B2(
        P1_REG3_REG_2__SCAN_IN), .ZN(n7854) );
  OAI211_X1 U9527 ( .C1(n9066), .C2(n7856), .A(n7855), .B(n7854), .ZN(n7857)
         );
  OR2_X1 U9528 ( .A1(n7858), .A2(n7857), .ZN(P1_U3289) );
  NAND2_X1 U9529 ( .A1(n7875), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n7868) );
  INV_X1 U9530 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n7859) );
  MUX2_X1 U9531 ( .A(n7859), .B(P2_REG2_REG_17__SCAN_IN), .S(n7875), .Z(n7860)
         );
  INV_X1 U9532 ( .A(n7860), .ZN(n7883) );
  NAND2_X1 U9533 ( .A1(n8258), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n7867) );
  INV_X1 U9534 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n7861) );
  MUX2_X1 U9535 ( .A(n7861), .B(P2_REG2_REG_16__SCAN_IN), .S(n8258), .Z(n7862)
         );
  INV_X1 U9536 ( .A(n7862), .ZN(n8256) );
  NOR2_X1 U9537 ( .A1(n7864), .A2(n7863), .ZN(n7866) );
  NOR2_X1 U9538 ( .A1(n7866), .A2(n7865), .ZN(n8257) );
  NAND2_X1 U9539 ( .A1(n8256), .A2(n8257), .ZN(n8255) );
  NAND2_X1 U9540 ( .A1(n7867), .A2(n8255), .ZN(n7884) );
  NAND2_X1 U9541 ( .A1(n7883), .A2(n7884), .ZN(n7882) );
  NAND2_X1 U9542 ( .A1(n7868), .A2(n7882), .ZN(n8018) );
  XOR2_X1 U9543 ( .A(n8022), .B(n8018), .Z(n7869) );
  NAND2_X1 U9544 ( .A1(P2_REG2_REG_18__SCAN_IN), .A2(n7869), .ZN(n8019) );
  OAI211_X1 U9545 ( .C1(n7869), .C2(P2_REG2_REG_18__SCAN_IN), .A(n9680), .B(
        n8019), .ZN(n7880) );
  INV_X1 U9546 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n7870) );
  XNOR2_X1 U9547 ( .A(n8022), .B(n7870), .ZN(n8025) );
  XNOR2_X1 U9548 ( .A(n7875), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n7887) );
  XOR2_X1 U9549 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n8258), .Z(n8250) );
  NOR2_X1 U9550 ( .A1(n7872), .A2(n7871), .ZN(n7874) );
  AOI21_X1 U9551 ( .B1(P2_REG1_REG_17__SCAN_IN), .B2(n7875), .A(n7886), .ZN(
        n8024) );
  XNOR2_X1 U9552 ( .A(n8025), .B(n8024), .ZN(n7878) );
  NOR2_X1 U9553 ( .A1(n8033), .A2(n10019), .ZN(n7876) );
  AOI211_X1 U9554 ( .C1(n9679), .C2(n7878), .A(n7877), .B(n7876), .ZN(n7879)
         );
  OAI211_X1 U9555 ( .C1(n8030), .C2(n7881), .A(n7880), .B(n7879), .ZN(P2_U3263) );
  OAI211_X1 U9556 ( .C1(n7884), .C2(n7883), .A(n9680), .B(n7882), .ZN(n7892)
         );
  NOR2_X1 U9557 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7885), .ZN(n7890) );
  AOI211_X1 U9558 ( .C1(n7888), .C2(n7887), .A(n7886), .B(n9682), .ZN(n7889)
         );
  AOI211_X1 U9559 ( .C1(n9681), .C2(P2_ADDR_REG_17__SCAN_IN), .A(n7890), .B(
        n7889), .ZN(n7891) );
  OAI211_X1 U9560 ( .C1(n8030), .C2(n7893), .A(n7892), .B(n7891), .ZN(P2_U3262) );
  AOI21_X1 U9561 ( .B1(n7896), .B2(n7895), .A(n7894), .ZN(n7897) );
  OR2_X1 U9562 ( .A1(n7897), .A2(n8027), .ZN(n7906) );
  AOI21_X1 U9563 ( .B1(n7900), .B2(n7899), .A(n7898), .ZN(n7904) );
  INV_X1 U9564 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n7902) );
  OR2_X1 U9565 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8203), .ZN(n7901) );
  OAI21_X1 U9566 ( .B1(n8033), .B2(n7902), .A(n7901), .ZN(n7903) );
  AOI21_X1 U9567 ( .B1(n9679), .B2(n7904), .A(n7903), .ZN(n7905) );
  OAI211_X1 U9568 ( .C1(n8030), .C2(n7907), .A(n7906), .B(n7905), .ZN(P2_U3256) );
  NAND2_X1 U9569 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(P2_U3152), .ZN(n8111) );
  INV_X1 U9570 ( .A(n8111), .ZN(n7912) );
  AOI211_X1 U9571 ( .C1(n7910), .C2(n7909), .A(n7908), .B(n9682), .ZN(n7911)
         );
  AOI211_X1 U9572 ( .C1(n9681), .C2(P2_ADDR_REG_10__SCAN_IN), .A(n7912), .B(
        n7911), .ZN(n7917) );
  OAI211_X1 U9573 ( .C1(n7915), .C2(n7914), .A(n9680), .B(n7913), .ZN(n7916)
         );
  OAI211_X1 U9574 ( .C1(n8030), .C2(n7918), .A(n7917), .B(n7916), .ZN(P2_U3255) );
  INV_X1 U9575 ( .A(n7919), .ZN(n7924) );
  AOI211_X1 U9576 ( .C1(n7922), .C2(n7921), .A(n7920), .B(n9682), .ZN(n7923)
         );
  AOI211_X1 U9577 ( .C1(n9681), .C2(P2_ADDR_REG_9__SCAN_IN), .A(n7924), .B(
        n7923), .ZN(n7929) );
  OAI211_X1 U9578 ( .C1(n7927), .C2(n7926), .A(n9680), .B(n7925), .ZN(n7928)
         );
  OAI211_X1 U9579 ( .C1(n8030), .C2(n7930), .A(n7929), .B(n7928), .ZN(P2_U3254) );
  NAND2_X1 U9580 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(P2_U3152), .ZN(n8137) );
  INV_X1 U9581 ( .A(n8137), .ZN(n7935) );
  AOI211_X1 U9582 ( .C1(n7933), .C2(n7932), .A(n7931), .B(n9682), .ZN(n7934)
         );
  AOI211_X1 U9583 ( .C1(n9681), .C2(P2_ADDR_REG_8__SCAN_IN), .A(n7935), .B(
        n7934), .ZN(n7940) );
  OAI211_X1 U9584 ( .C1(n7938), .C2(n7937), .A(n9680), .B(n7936), .ZN(n7939)
         );
  OAI211_X1 U9585 ( .C1(n8030), .C2(n7941), .A(n7940), .B(n7939), .ZN(P2_U3253) );
  NOR2_X1 U9586 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n5005), .ZN(n7946) );
  AOI211_X1 U9587 ( .C1(n7944), .C2(n7943), .A(n7942), .B(n9682), .ZN(n7945)
         );
  AOI211_X1 U9588 ( .C1(n9681), .C2(P2_ADDR_REG_7__SCAN_IN), .A(n7946), .B(
        n7945), .ZN(n7951) );
  OAI211_X1 U9589 ( .C1(n7949), .C2(n7948), .A(n9680), .B(n7947), .ZN(n7950)
         );
  OAI211_X1 U9590 ( .C1(n8030), .C2(n7952), .A(n7951), .B(n7950), .ZN(P2_U3252) );
  NOR2_X1 U9591 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7953), .ZN(n7958) );
  AOI211_X1 U9592 ( .C1(n7956), .C2(n7955), .A(n7954), .B(n9682), .ZN(n7957)
         );
  AOI211_X1 U9593 ( .C1(n9681), .C2(P2_ADDR_REG_6__SCAN_IN), .A(n7958), .B(
        n7957), .ZN(n7963) );
  OAI211_X1 U9594 ( .C1(n7961), .C2(n7960), .A(n9680), .B(n7959), .ZN(n7962)
         );
  OAI211_X1 U9595 ( .C1(n8030), .C2(n7964), .A(n7963), .B(n7962), .ZN(P2_U3251) );
  AND2_X1 U9596 ( .A1(P2_U3152), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n7969) );
  AOI211_X1 U9597 ( .C1(n7967), .C2(n7966), .A(n7965), .B(n9682), .ZN(n7968)
         );
  AOI211_X1 U9598 ( .C1(n9681), .C2(P2_ADDR_REG_5__SCAN_IN), .A(n7969), .B(
        n7968), .ZN(n7974) );
  OAI211_X1 U9599 ( .C1(n7972), .C2(n7971), .A(n9680), .B(n7970), .ZN(n7973)
         );
  OAI211_X1 U9600 ( .C1(n8030), .C2(n4280), .A(n7974), .B(n7973), .ZN(P2_U3250) );
  AND2_X1 U9601 ( .A1(P2_U3152), .A2(P2_REG3_REG_4__SCAN_IN), .ZN(n7979) );
  AOI211_X1 U9602 ( .C1(n7977), .C2(n7976), .A(n7975), .B(n9682), .ZN(n7978)
         );
  AOI211_X1 U9603 ( .C1(n9681), .C2(P2_ADDR_REG_4__SCAN_IN), .A(n7979), .B(
        n7978), .ZN(n7988) );
  INV_X1 U9604 ( .A(n7980), .ZN(n7998) );
  INV_X1 U9605 ( .A(n7981), .ZN(n7984) );
  MUX2_X1 U9606 ( .A(n7327), .B(P2_REG2_REG_4__SCAN_IN), .S(n7982), .Z(n7983)
         );
  NAND3_X1 U9607 ( .A1(n7998), .A2(n7984), .A3(n7983), .ZN(n7985) );
  NAND3_X1 U9608 ( .A1(n9680), .A2(n7986), .A3(n7985), .ZN(n7987) );
  OAI211_X1 U9609 ( .C1(n8030), .C2(n7989), .A(n7988), .B(n7987), .ZN(P2_U3249) );
  NOR2_X1 U9610 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n4911), .ZN(n7994) );
  AOI211_X1 U9611 ( .C1(n7992), .C2(n7991), .A(n7990), .B(n9682), .ZN(n7993)
         );
  AOI211_X1 U9612 ( .C1(n9681), .C2(P2_ADDR_REG_3__SCAN_IN), .A(n7994), .B(
        n7993), .ZN(n8000) );
  NAND3_X1 U9613 ( .A1(n8014), .A2(n7996), .A3(n7995), .ZN(n7997) );
  NAND3_X1 U9614 ( .A1(n9680), .A2(n7998), .A3(n7997), .ZN(n7999) );
  OAI211_X1 U9615 ( .C1(n8030), .C2(n8001), .A(n8000), .B(n7999), .ZN(P2_U3248) );
  NOR2_X1 U9616 ( .A1(n8002), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8007) );
  AOI211_X1 U9617 ( .C1(n8005), .C2(n8004), .A(n8003), .B(n9682), .ZN(n8006)
         );
  AOI211_X1 U9618 ( .C1(n9681), .C2(P2_ADDR_REG_2__SCAN_IN), .A(n8007), .B(
        n8006), .ZN(n8016) );
  MUX2_X1 U9619 ( .A(n9883), .B(P2_REG2_REG_2__SCAN_IN), .S(n8008), .Z(n8012)
         );
  INV_X1 U9620 ( .A(n8009), .ZN(n8010) );
  NAND3_X1 U9621 ( .A1(n8012), .A2(n8011), .A3(n8010), .ZN(n8013) );
  NAND3_X1 U9622 ( .A1(n9680), .A2(n8014), .A3(n8013), .ZN(n8015) );
  OAI211_X1 U9623 ( .C1(n8030), .C2(n8017), .A(n8016), .B(n8015), .ZN(P2_U3247) );
  NAND2_X1 U9624 ( .A1(n8018), .A2(n8022), .ZN(n8020) );
  NAND2_X1 U9625 ( .A1(n8020), .A2(n8019), .ZN(n8021) );
  NOR2_X1 U9626 ( .A1(n8022), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n8023) );
  AOI21_X1 U9627 ( .B1(n8025), .B2(n8024), .A(n8023), .ZN(n8026) );
  XNOR2_X1 U9628 ( .A(n8026), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n8029) );
  OAI22_X1 U9629 ( .A1(n4270), .A2(n8027), .B1(n8029), .B2(n9682), .ZN(n8031)
         );
  INV_X1 U9630 ( .A(n8028), .ZN(n9683) );
  NAND2_X1 U9631 ( .A1(P2_U3152), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n8125) );
  OAI211_X1 U9632 ( .C1(n4760), .C2(n8033), .A(n8032), .B(n8125), .ZN(P2_U3264) );
  INV_X1 U9633 ( .A(n8717), .ZN(n9388) );
  AOI22_X1 U9634 ( .A1(n8034), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_30__SCAN_IN), .B2(n8556), .ZN(n8035) );
  OAI21_X1 U9635 ( .B1(n9388), .B2(n8049), .A(n8035), .ZN(P2_U3328) );
  NAND2_X1 U9636 ( .A1(n8036), .A2(n8700), .ZN(n8038) );
  AOI22_X1 U9637 ( .A1(n8667), .A2(P1_REG3_REG_0__SCAN_IN), .B1(n8680), .B2(
        n6311), .ZN(n8037) );
  OAI211_X1 U9638 ( .C1(n8039), .C2(n8676), .A(n8038), .B(n8037), .ZN(P1_U3230) );
  OAI21_X1 U9639 ( .B1(n8042), .B2(n8041), .A(n8040), .ZN(n8043) );
  NAND2_X1 U9640 ( .A1(n8043), .A2(n8214), .ZN(n8047) );
  AOI22_X1 U9641 ( .A1(n8045), .A2(n8175), .B1(n8044), .B2(
        P2_REG3_REG_1__SCAN_IN), .ZN(n8046) );
  OAI211_X1 U9642 ( .C1(n7462), .C2(n8227), .A(n8047), .B(n8046), .ZN(P2_U3224) );
  OAI222_X1 U9643 ( .A1(n8051), .A2(n8050), .B1(n8049), .B2(n8048), .C1(n5645), 
        .C2(P2_U3152), .ZN(P2_U3339) );
  OR2_X1 U9644 ( .A1(n8526), .A2(n8444), .ZN(n8052) );
  NOR2_X1 U9645 ( .A1(n8519), .A2(n8425), .ZN(n8055) );
  NAND2_X1 U9646 ( .A1(n8519), .A2(n8425), .ZN(n8054) );
  AND2_X1 U9647 ( .A1(n8515), .A2(n8446), .ZN(n8056) );
  OR2_X1 U9648 ( .A1(n8502), .A2(n8410), .ZN(n8057) );
  INV_X1 U9649 ( .A(n8361), .ZN(n8402) );
  NOR2_X1 U9650 ( .A1(n8497), .A2(n8402), .ZN(n8058) );
  INV_X1 U9651 ( .A(n8383), .ZN(n8232) );
  NAND2_X1 U9652 ( .A1(n8324), .A2(n8332), .ZN(n8323) );
  NAND2_X1 U9653 ( .A1(n8323), .A2(n8061), .ZN(n8306) );
  NAND2_X1 U9654 ( .A1(n8305), .A2(n8062), .ZN(n8289) );
  NAND2_X1 U9655 ( .A1(n8289), .A2(n8298), .ZN(n8288) );
  INV_X1 U9656 ( .A(n8314), .ZN(n8229) );
  NAND2_X1 U9657 ( .A1(n8288), .A2(n8063), .ZN(n8275) );
  NAND2_X1 U9658 ( .A1(n8275), .A2(n8281), .ZN(n8274) );
  INV_X1 U9659 ( .A(n8519), .ZN(n8441) );
  INV_X1 U9660 ( .A(n8502), .ZN(n8396) );
  INV_X1 U9661 ( .A(n8481), .ZN(n8331) );
  INV_X1 U9662 ( .A(n8477), .ZN(n8320) );
  INV_X1 U9663 ( .A(n8470), .ZN(n8296) );
  NOR2_X2 U9664 ( .A1(n8277), .A2(n8460), .ZN(n8268) );
  AOI21_X1 U9665 ( .B1(n8460), .B2(n8277), .A(n8268), .ZN(n8461) );
  INV_X1 U9666 ( .A(n8460), .ZN(n8068) );
  INV_X1 U9667 ( .A(n8065), .ZN(n8066) );
  AOI22_X1 U9668 ( .A1(n8066), .A2(n9993), .B1(n10001), .B2(
        P2_REG2_REG_29__SCAN_IN), .ZN(n8067) );
  OAI21_X1 U9669 ( .B1(n8068), .B2(n8415), .A(n8067), .ZN(n8077) );
  OAI21_X1 U9670 ( .B1(n8071), .B2(n8070), .A(n8069), .ZN(n8076) );
  NAND2_X1 U9671 ( .A1(n8299), .A2(n8443), .ZN(n8074) );
  AOI21_X1 U9672 ( .B1(n8072), .B2(P2_B_REG_SCAN_IN), .A(n9756), .ZN(n8263) );
  NAND2_X1 U9673 ( .A1(n8228), .A2(n8263), .ZN(n8073) );
  AOI21_X2 U9674 ( .B1(n8076), .B2(n9693), .A(n8075), .ZN(n8463) );
  OAI21_X1 U9675 ( .B1(n8464), .B2(n8452), .A(n8078), .ZN(P2_U3267) );
  NAND2_X1 U9676 ( .A1(n8080), .A2(n8079), .ZN(n8081) );
  XOR2_X1 U9677 ( .A(n8082), .B(n8081), .Z(n8083) );
  NAND2_X1 U9678 ( .A1(n8083), .A2(n8214), .ZN(n8092) );
  OAI22_X1 U9679 ( .A1(n9759), .A2(n8221), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n5005), .ZN(n8086) );
  NOR2_X1 U9680 ( .A1(n8084), .A2(n8220), .ZN(n8085) );
  NOR2_X1 U9681 ( .A1(n8086), .A2(n8085), .ZN(n8091) );
  NAND2_X1 U9682 ( .A1(n8207), .A2(n8087), .ZN(n8090) );
  NAND2_X1 U9683 ( .A1(n8224), .A2(n8088), .ZN(n8089) );
  NAND4_X1 U9684 ( .A1(n8092), .A2(n8091), .A3(n8090), .A4(n8089), .ZN(
        P2_U3215) );
  OAI211_X1 U9685 ( .C1(n8095), .C2(n8094), .A(n8093), .B(n8214), .ZN(n8101)
         );
  OAI22_X1 U9686 ( .A1(n8096), .A2(n8220), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9973), .ZN(n8099) );
  NOR2_X1 U9687 ( .A1(n8097), .A2(n8221), .ZN(n8098) );
  AOI211_X1 U9688 ( .C1(n8224), .C2(n8294), .A(n8099), .B(n8098), .ZN(n8100)
         );
  OAI211_X1 U9689 ( .C1(n8296), .C2(n8227), .A(n8101), .B(n8100), .ZN(P2_U3216) );
  XNOR2_X1 U9690 ( .A(n8169), .B(n8170), .ZN(n8107) );
  NOR2_X1 U9691 ( .A1(n8361), .A2(n8220), .ZN(n8104) );
  OAI22_X1 U9692 ( .A1(n8362), .A2(n8221), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8102), .ZN(n8103) );
  AOI211_X1 U9693 ( .C1(n8224), .C2(n8368), .A(n8104), .B(n8103), .ZN(n8106)
         );
  NAND2_X1 U9694 ( .A1(n8367), .A2(n8207), .ZN(n8105) );
  OAI211_X1 U9695 ( .C1(n8107), .C2(n8189), .A(n8106), .B(n8105), .ZN(P2_U3218) );
  XOR2_X1 U9696 ( .A(n8109), .B(n8108), .Z(n8110) );
  NAND2_X1 U9697 ( .A1(n8110), .A2(n8214), .ZN(n8120) );
  OAI21_X1 U9698 ( .B1(n8112), .B2(n8221), .A(n8111), .ZN(n8114) );
  NOR2_X1 U9699 ( .A1(n8138), .A2(n8220), .ZN(n8113) );
  NOR2_X1 U9700 ( .A1(n8114), .A2(n8113), .ZN(n8119) );
  NAND2_X1 U9701 ( .A1(n8207), .A2(n8115), .ZN(n8118) );
  NAND2_X1 U9702 ( .A1(n8224), .A2(n8116), .ZN(n8117) );
  NAND4_X1 U9703 ( .A1(n8120), .A2(n8119), .A3(n8118), .A4(n8117), .ZN(
        P2_U3219) );
  INV_X1 U9704 ( .A(n8121), .ZN(n8122) );
  AOI21_X1 U9705 ( .B1(n8124), .B2(n8123), .A(n8122), .ZN(n8131) );
  NAND2_X1 U9706 ( .A1(n8426), .A2(n8195), .ZN(n8126) );
  OAI211_X1 U9707 ( .C1(n8127), .C2(n8220), .A(n8126), .B(n8125), .ZN(n8128)
         );
  AOI21_X1 U9708 ( .B1(n8430), .B2(n8224), .A(n8128), .ZN(n8130) );
  NAND2_X1 U9709 ( .A1(n8515), .A2(n8207), .ZN(n8129) );
  OAI211_X1 U9710 ( .C1(n8131), .C2(n8189), .A(n8130), .B(n8129), .ZN(P2_U3221) );
  NAND2_X1 U9711 ( .A1(n8133), .A2(n8132), .ZN(n8134) );
  XOR2_X1 U9712 ( .A(n8135), .B(n8134), .Z(n8136) );
  NAND2_X1 U9713 ( .A1(n8136), .A2(n8214), .ZN(n8147) );
  OAI21_X1 U9714 ( .B1(n8138), .B2(n8221), .A(n8137), .ZN(n8141) );
  NOR2_X1 U9715 ( .A1(n8139), .A2(n8220), .ZN(n8140) );
  NOR2_X1 U9716 ( .A1(n8141), .A2(n8140), .ZN(n8146) );
  NAND2_X1 U9717 ( .A1(n8207), .A2(n8142), .ZN(n8145) );
  NAND2_X1 U9718 ( .A1(n8224), .A2(n8143), .ZN(n8144) );
  NAND4_X1 U9719 ( .A1(n8147), .A2(n8146), .A3(n8145), .A4(n8144), .ZN(
        P2_U3223) );
  OR2_X1 U9720 ( .A1(n8183), .A2(n8182), .ZN(n8149) );
  NAND2_X1 U9721 ( .A1(n8149), .A2(n8148), .ZN(n8151) );
  XNOR2_X1 U9722 ( .A(n8151), .B(n8150), .ZN(n8157) );
  AOI22_X1 U9723 ( .A1(n8402), .A2(n8195), .B1(P2_REG3_REG_21__SCAN_IN), .B2(
        P2_U3152), .ZN(n8153) );
  NAND2_X1 U9724 ( .A1(n8224), .A2(n8394), .ZN(n8152) );
  OAI211_X1 U9725 ( .C1(n8154), .C2(n8220), .A(n8153), .B(n8152), .ZN(n8155)
         );
  AOI21_X1 U9726 ( .B1(n8502), .B2(n8207), .A(n8155), .ZN(n8156) );
  OAI21_X1 U9727 ( .B1(n8157), .B2(n8189), .A(n8156), .ZN(P2_U3225) );
  XNOR2_X1 U9728 ( .A(n8159), .B(n8158), .ZN(n8160) );
  XNOR2_X1 U9729 ( .A(n8161), .B(n8160), .ZN(n8167) );
  NAND2_X1 U9730 ( .A1(n8300), .A2(n8445), .ZN(n8163) );
  OR2_X1 U9731 ( .A1(n8362), .A2(n9758), .ZN(n8162) );
  NAND2_X1 U9732 ( .A1(n8163), .A2(n8162), .ZN(n8334) );
  AOI22_X1 U9733 ( .A1(n8334), .A2(n8175), .B1(P2_REG3_REG_25__SCAN_IN), .B2(
        P2_U3152), .ZN(n8164) );
  OAI21_X1 U9734 ( .B1(n8328), .B2(n8177), .A(n8164), .ZN(n8165) );
  AOI21_X1 U9735 ( .B1(n8481), .B2(n8207), .A(n8165), .ZN(n8166) );
  OAI21_X1 U9736 ( .B1(n8167), .B2(n8189), .A(n8166), .ZN(P2_U3227) );
  AOI21_X1 U9737 ( .B1(n8170), .B2(n8169), .A(n8168), .ZN(n8174) );
  XNOR2_X1 U9738 ( .A(n8172), .B(n8171), .ZN(n8173) );
  XNOR2_X1 U9739 ( .A(n8174), .B(n8173), .ZN(n8181) );
  INV_X1 U9740 ( .A(n8347), .ZN(n8178) );
  OAI22_X1 U9741 ( .A1(n8313), .A2(n9756), .B1(n8383), .B2(n9758), .ZN(n8340)
         );
  AOI22_X1 U9742 ( .A1(n8340), .A2(n8175), .B1(P2_REG3_REG_24__SCAN_IN), .B2(
        P2_U3152), .ZN(n8176) );
  OAI21_X1 U9743 ( .B1(n8178), .B2(n8177), .A(n8176), .ZN(n8179) );
  AOI21_X1 U9744 ( .B1(n8486), .B2(n8207), .A(n8179), .ZN(n8180) );
  OAI21_X1 U9745 ( .B1(n8181), .B2(n8189), .A(n8180), .ZN(P2_U3231) );
  XNOR2_X1 U9746 ( .A(n8183), .B(n8182), .ZN(n8190) );
  AOI22_X1 U9747 ( .A1(n8195), .A2(n8410), .B1(P2_REG3_REG_20__SCAN_IN), .B2(
        P2_U3152), .ZN(n8185) );
  NAND2_X1 U9748 ( .A1(n8224), .A2(n8413), .ZN(n8184) );
  OAI211_X1 U9749 ( .C1(n8186), .C2(n8220), .A(n8185), .B(n8184), .ZN(n8187)
         );
  AOI21_X1 U9750 ( .B1(n8509), .B2(n8207), .A(n8187), .ZN(n8188) );
  OAI21_X1 U9751 ( .B1(n8190), .B2(n8189), .A(n8188), .ZN(P2_U3235) );
  INV_X1 U9752 ( .A(n8497), .ZN(n8377) );
  OAI21_X1 U9753 ( .B1(n8193), .B2(n8192), .A(n8191), .ZN(n8194) );
  NAND2_X1 U9754 ( .A1(n8194), .A2(n8214), .ZN(n8199) );
  AOI22_X1 U9755 ( .A1(n8232), .A2(n8195), .B1(P2_REG3_REG_22__SCAN_IN), .B2(
        P2_U3152), .ZN(n8196) );
  OAI21_X1 U9756 ( .B1(n8384), .B2(n8220), .A(n8196), .ZN(n8197) );
  AOI21_X1 U9757 ( .B1(n8375), .B2(n8224), .A(n8197), .ZN(n8198) );
  OAI211_X1 U9758 ( .C1(n8377), .C2(n8227), .A(n8199), .B(n8198), .ZN(P2_U3237) );
  XOR2_X1 U9759 ( .A(n8201), .B(n8200), .Z(n8202) );
  NAND2_X1 U9760 ( .A1(n8202), .A2(n8214), .ZN(n8213) );
  OAI22_X1 U9761 ( .A1(n8204), .A2(n8221), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8203), .ZN(n8206) );
  NOR2_X1 U9762 ( .A1(n9757), .A2(n8220), .ZN(n8205) );
  NOR2_X1 U9763 ( .A1(n8206), .A2(n8205), .ZN(n8212) );
  NAND2_X1 U9764 ( .A1(n8208), .A2(n8207), .ZN(n8211) );
  NAND2_X1 U9765 ( .A1(n8224), .A2(n8209), .ZN(n8210) );
  NAND4_X1 U9766 ( .A1(n8213), .A2(n8212), .A3(n8211), .A4(n8210), .ZN(
        P2_U3238) );
  OAI211_X1 U9767 ( .C1(n8217), .C2(n8216), .A(n8215), .B(n8214), .ZN(n8226)
         );
  INV_X1 U9768 ( .A(n8218), .ZN(n8317) );
  OAI22_X1 U9769 ( .A1(n8313), .A2(n8220), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8219), .ZN(n8223) );
  NOR2_X1 U9770 ( .A1(n8314), .A2(n8221), .ZN(n8222) );
  AOI211_X1 U9771 ( .C1(n8224), .C2(n8317), .A(n8223), .B(n8222), .ZN(n8225)
         );
  OAI211_X1 U9772 ( .C1(n8320), .C2(n8227), .A(n8226), .B(n8225), .ZN(P2_U3242) );
  MUX2_X1 U9773 ( .A(n8228), .B(P2_DATAO_REG_30__SCAN_IN), .S(n8248), .Z(
        P2_U3582) );
  MUX2_X1 U9774 ( .A(n8299), .B(P2_DATAO_REG_28__SCAN_IN), .S(n8248), .Z(
        P2_U3580) );
  MUX2_X1 U9775 ( .A(n8229), .B(P2_DATAO_REG_27__SCAN_IN), .S(n8248), .Z(
        P2_U3579) );
  MUX2_X1 U9776 ( .A(n8300), .B(P2_DATAO_REG_26__SCAN_IN), .S(n8248), .Z(
        P2_U3578) );
  MUX2_X1 U9777 ( .A(n8230), .B(P2_DATAO_REG_25__SCAN_IN), .S(n8248), .Z(
        P2_U3577) );
  MUX2_X1 U9778 ( .A(n8231), .B(P2_DATAO_REG_24__SCAN_IN), .S(n8248), .Z(
        P2_U3576) );
  MUX2_X1 U9779 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(n8232), .S(P2_U3966), .Z(
        P2_U3575) );
  MUX2_X1 U9780 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n8402), .S(P2_U3966), .Z(
        P2_U3574) );
  MUX2_X1 U9781 ( .A(n8410), .B(P2_DATAO_REG_21__SCAN_IN), .S(n8248), .Z(
        P2_U3573) );
  MUX2_X1 U9782 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n8426), .S(P2_U3966), .Z(
        P2_U3572) );
  MUX2_X1 U9783 ( .A(n8446), .B(P2_DATAO_REG_19__SCAN_IN), .S(n8248), .Z(
        P2_U3571) );
  MUX2_X1 U9784 ( .A(n8425), .B(P2_DATAO_REG_18__SCAN_IN), .S(n8248), .Z(
        P2_U3570) );
  MUX2_X1 U9785 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n8444), .S(P2_U3966), .Z(
        P2_U3569) );
  MUX2_X1 U9786 ( .A(n8233), .B(P2_DATAO_REG_16__SCAN_IN), .S(n8248), .Z(
        P2_U3568) );
  MUX2_X1 U9787 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(n8234), .S(P2_U3966), .Z(
        P2_U3567) );
  MUX2_X1 U9788 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(n8235), .S(P2_U3966), .Z(
        P2_U3566) );
  MUX2_X1 U9789 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(n8236), .S(P2_U3966), .Z(
        P2_U3565) );
  MUX2_X1 U9790 ( .A(n8237), .B(P2_DATAO_REG_12__SCAN_IN), .S(n8248), .Z(
        P2_U3564) );
  MUX2_X1 U9791 ( .A(n8238), .B(P2_DATAO_REG_11__SCAN_IN), .S(n8248), .Z(
        P2_U3563) );
  MUX2_X1 U9792 ( .A(n8239), .B(P2_DATAO_REG_10__SCAN_IN), .S(n8248), .Z(
        P2_U3562) );
  MUX2_X1 U9793 ( .A(n8240), .B(P2_DATAO_REG_9__SCAN_IN), .S(n8248), .Z(
        P2_U3561) );
  MUX2_X1 U9794 ( .A(n8241), .B(P2_DATAO_REG_8__SCAN_IN), .S(n8248), .Z(
        P2_U3560) );
  MUX2_X1 U9795 ( .A(n8242), .B(P2_DATAO_REG_7__SCAN_IN), .S(n8248), .Z(
        P2_U3559) );
  MUX2_X1 U9796 ( .A(n8243), .B(P2_DATAO_REG_6__SCAN_IN), .S(n8248), .Z(
        P2_U3558) );
  MUX2_X1 U9797 ( .A(n8244), .B(P2_DATAO_REG_5__SCAN_IN), .S(n8248), .Z(
        P2_U3557) );
  MUX2_X1 U9798 ( .A(n8245), .B(P2_DATAO_REG_4__SCAN_IN), .S(n8248), .Z(
        P2_U3556) );
  MUX2_X1 U9799 ( .A(n8246), .B(P2_DATAO_REG_3__SCAN_IN), .S(n8248), .Z(
        P2_U3555) );
  MUX2_X1 U9800 ( .A(n8247), .B(P2_DATAO_REG_2__SCAN_IN), .S(n8248), .Z(
        P2_U3554) );
  MUX2_X1 U9801 ( .A(n6864), .B(P2_DATAO_REG_1__SCAN_IN), .S(n8248), .Z(
        P2_U3553) );
  OAI21_X1 U9802 ( .B1(n8251), .B2(n8250), .A(n8249), .ZN(n8252) );
  NAND2_X1 U9803 ( .A1(n8252), .A2(n9679), .ZN(n8262) );
  INV_X1 U9804 ( .A(n8253), .ZN(n8254) );
  AOI21_X1 U9805 ( .B1(n9681), .B2(P2_ADDR_REG_16__SCAN_IN), .A(n8254), .ZN(
        n8261) );
  OAI211_X1 U9806 ( .C1(n8257), .C2(n8256), .A(n9680), .B(n8255), .ZN(n8260)
         );
  NAND2_X1 U9807 ( .A1(n9684), .A2(n8258), .ZN(n8259) );
  NAND4_X1 U9808 ( .A1(n8262), .A2(n8261), .A3(n8260), .A4(n8259), .ZN(
        P2_U3261) );
  NAND2_X1 U9809 ( .A1(n8264), .A2(n8263), .ZN(n8457) );
  NOR2_X1 U9810 ( .A1(n8457), .A2(n10001), .ZN(n8271) );
  NOR2_X1 U9811 ( .A1(n8265), .A2(n8415), .ZN(n8266) );
  AOI211_X1 U9812 ( .C1(P2_REG2_REG_31__SCAN_IN), .C2(n9706), .A(n8271), .B(
        n8266), .ZN(n8267) );
  OAI21_X1 U9813 ( .B1(n9999), .B2(n8454), .A(n8267), .ZN(P2_U3265) );
  INV_X1 U9814 ( .A(n8268), .ZN(n8270) );
  NAND2_X1 U9815 ( .A1(n8270), .A2(n8269), .ZN(n8456) );
  NAND3_X1 U9816 ( .A1(n8456), .A2(n8450), .A3(n8455), .ZN(n8273) );
  AOI21_X1 U9817 ( .B1(n9706), .B2(P2_REG2_REG_30__SCAN_IN), .A(n8271), .ZN(
        n8272) );
  OAI211_X1 U9818 ( .C1(n8459), .C2(n8415), .A(n8273), .B(n8272), .ZN(P2_U3266) );
  OAI21_X1 U9819 ( .B1(n8275), .B2(n8281), .A(n8274), .ZN(n8276) );
  INV_X1 U9820 ( .A(n8276), .ZN(n8469) );
  INV_X1 U9821 ( .A(n8277), .ZN(n8278) );
  AOI211_X1 U9822 ( .C1(n8466), .C2(n8291), .A(n9780), .B(n8278), .ZN(n8465)
         );
  AOI22_X1 U9823 ( .A1(n8279), .A2(n9993), .B1(P2_REG2_REG_28__SCAN_IN), .B2(
        n10001), .ZN(n8280) );
  OAI21_X1 U9824 ( .B1(n4501), .B2(n8415), .A(n8280), .ZN(n8286) );
  XNOR2_X1 U9825 ( .A(n8282), .B(n8281), .ZN(n8284) );
  AOI21_X1 U9826 ( .B1(n8284), .B2(n9693), .A(n8283), .ZN(n8468) );
  NOR2_X1 U9827 ( .A1(n8468), .A2(n10001), .ZN(n8285) );
  AOI211_X1 U9828 ( .C1(n8465), .C2(n9702), .A(n8286), .B(n8285), .ZN(n8287)
         );
  OAI21_X1 U9829 ( .B1(n8469), .B2(n8452), .A(n8287), .ZN(P2_U3268) );
  OAI21_X1 U9830 ( .B1(n8289), .B2(n8298), .A(n8288), .ZN(n8290) );
  INV_X1 U9831 ( .A(n8290), .ZN(n8474) );
  INV_X1 U9832 ( .A(n8315), .ZN(n8293) );
  INV_X1 U9833 ( .A(n8291), .ZN(n8292) );
  AOI21_X1 U9834 ( .B1(n8470), .B2(n8293), .A(n8292), .ZN(n8471) );
  AOI22_X1 U9835 ( .A1(P2_REG2_REG_27__SCAN_IN), .A2(n10001), .B1(n8294), .B2(
        n9993), .ZN(n8295) );
  OAI21_X1 U9836 ( .B1(n8296), .B2(n8415), .A(n8295), .ZN(n8303) );
  XOR2_X1 U9837 ( .A(n8298), .B(n8297), .Z(n8301) );
  AOI222_X1 U9838 ( .A1(n9693), .A2(n8301), .B1(n8300), .B2(n8443), .C1(n8299), 
        .C2(n8445), .ZN(n8473) );
  NOR2_X1 U9839 ( .A1(n8473), .A2(n10001), .ZN(n8302) );
  OAI21_X1 U9840 ( .B1(n8474), .B2(n8452), .A(n8304), .ZN(P2_U3269) );
  OAI21_X1 U9841 ( .B1(n8306), .B2(n8311), .A(n8305), .ZN(n8307) );
  INV_X1 U9842 ( .A(n8307), .ZN(n8479) );
  INV_X1 U9843 ( .A(n8308), .ZN(n8309) );
  AOI21_X1 U9844 ( .B1(n8311), .B2(n8310), .A(n8309), .ZN(n8312) );
  OAI222_X1 U9845 ( .A1(n9756), .A2(n8314), .B1(n9758), .B2(n8313), .C1(n9753), 
        .C2(n8312), .ZN(n8475) );
  INV_X1 U9846 ( .A(n8326), .ZN(n8316) );
  AOI211_X1 U9847 ( .C1(n8477), .C2(n8316), .A(n9780), .B(n8315), .ZN(n8476)
         );
  NAND2_X1 U9848 ( .A1(n8476), .A2(n9702), .ZN(n8319) );
  AOI22_X1 U9849 ( .A1(n9706), .A2(P2_REG2_REG_26__SCAN_IN), .B1(n8317), .B2(
        n9993), .ZN(n8318) );
  OAI211_X1 U9850 ( .C1(n8320), .C2(n8415), .A(n8319), .B(n8318), .ZN(n8321)
         );
  AOI21_X1 U9851 ( .B1(n8475), .B2(n7564), .A(n8321), .ZN(n8322) );
  OAI21_X1 U9852 ( .B1(n8479), .B2(n8452), .A(n8322), .ZN(P2_U3270) );
  OAI21_X1 U9853 ( .B1(n8324), .B2(n8332), .A(n8323), .ZN(n8325) );
  INV_X1 U9854 ( .A(n8325), .ZN(n8484) );
  INV_X1 U9855 ( .A(n8346), .ZN(n8327) );
  AOI211_X1 U9856 ( .C1(n8481), .C2(n8327), .A(n9780), .B(n8326), .ZN(n8480)
         );
  INV_X1 U9857 ( .A(n8328), .ZN(n8329) );
  AOI22_X1 U9858 ( .A1(n10001), .A2(P2_REG2_REG_25__SCAN_IN), .B1(n8329), .B2(
        n9993), .ZN(n8330) );
  OAI21_X1 U9859 ( .B1(n8331), .B2(n8415), .A(n8330), .ZN(n8337) );
  XNOR2_X1 U9860 ( .A(n8333), .B(n8332), .ZN(n8335) );
  AOI21_X1 U9861 ( .B1(n8335), .B2(n9693), .A(n8334), .ZN(n8483) );
  NOR2_X1 U9862 ( .A1(n8483), .A2(n10001), .ZN(n8336) );
  AOI211_X1 U9863 ( .C1(n9702), .C2(n8480), .A(n8337), .B(n8336), .ZN(n8338)
         );
  OAI21_X1 U9864 ( .B1(n8484), .B2(n8452), .A(n8338), .ZN(P2_U3271) );
  AOI21_X1 U9865 ( .B1(n8339), .B2(n8344), .A(n9753), .ZN(n8342) );
  AOI21_X1 U9866 ( .B1(n8342), .B2(n8341), .A(n8340), .ZN(n8489) );
  OAI21_X1 U9867 ( .B1(n8345), .B2(n8344), .A(n8343), .ZN(n8485) );
  NAND2_X1 U9868 ( .A1(n8485), .A2(n9703), .ZN(n8352) );
  AOI21_X1 U9869 ( .B1(n8486), .B2(n8366), .A(n8346), .ZN(n8487) );
  INV_X1 U9870 ( .A(n8486), .ZN(n8349) );
  AOI22_X1 U9871 ( .A1(n9706), .A2(P2_REG2_REG_24__SCAN_IN), .B1(n8347), .B2(
        n9993), .ZN(n8348) );
  OAI21_X1 U9872 ( .B1(n8349), .B2(n8415), .A(n8348), .ZN(n8350) );
  AOI21_X1 U9873 ( .B1(n8487), .B2(n8450), .A(n8350), .ZN(n8351) );
  OAI211_X1 U9874 ( .C1(n10001), .C2(n8489), .A(n8352), .B(n8351), .ZN(
        P2_U3272) );
  NOR2_X1 U9875 ( .A1(n8353), .A2(n8357), .ZN(n8354) );
  NAND2_X1 U9876 ( .A1(n8379), .A2(n8356), .ZN(n8358) );
  NAND2_X1 U9877 ( .A1(n8358), .A2(n8357), .ZN(n8360) );
  AOI21_X1 U9878 ( .B1(n8360), .B2(n8359), .A(n9753), .ZN(n8364) );
  OAI22_X1 U9879 ( .A1(n8362), .A2(n9756), .B1(n8361), .B2(n9758), .ZN(n8363)
         );
  OR2_X1 U9880 ( .A1(n8364), .A2(n8363), .ZN(n8494) );
  NAND2_X1 U9881 ( .A1(n8374), .A2(n8367), .ZN(n8365) );
  NAND2_X1 U9882 ( .A1(n8366), .A2(n8365), .ZN(n8492) );
  NOR2_X1 U9883 ( .A1(n8492), .A2(n9999), .ZN(n8371) );
  AOI22_X1 U9884 ( .A1(n10001), .A2(P2_REG2_REG_23__SCAN_IN), .B1(n8368), .B2(
        n9993), .ZN(n8369) );
  OAI21_X1 U9885 ( .B1(n4503), .B2(n8415), .A(n8369), .ZN(n8370) );
  AOI211_X1 U9886 ( .C1(n8494), .C2(n7564), .A(n8371), .B(n8370), .ZN(n8372)
         );
  OAI21_X1 U9887 ( .B1(n8491), .B2(n8452), .A(n8372), .ZN(P2_U3273) );
  XOR2_X1 U9888 ( .A(n8382), .B(n8373), .Z(n8501) );
  AOI21_X1 U9889 ( .B1(n8497), .B2(n8391), .A(n4504), .ZN(n8498) );
  AOI22_X1 U9890 ( .A1(n10001), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n8375), .B2(
        n9993), .ZN(n8376) );
  OAI21_X1 U9891 ( .B1(n8377), .B2(n8415), .A(n8376), .ZN(n8388) );
  NAND2_X1 U9892 ( .A1(n8399), .A2(n8378), .ZN(n8381) );
  INV_X1 U9893 ( .A(n8379), .ZN(n8380) );
  AOI211_X1 U9894 ( .C1(n8382), .C2(n8381), .A(n9753), .B(n8380), .ZN(n8386)
         );
  OAI22_X1 U9895 ( .A1(n8384), .A2(n9758), .B1(n8383), .B2(n9756), .ZN(n8385)
         );
  NOR2_X1 U9896 ( .A1(n8386), .A2(n8385), .ZN(n8500) );
  NOR2_X1 U9897 ( .A1(n8500), .A2(n9706), .ZN(n8387) );
  AOI211_X1 U9898 ( .C1(n8498), .C2(n8450), .A(n8388), .B(n8387), .ZN(n8389)
         );
  OAI21_X1 U9899 ( .B1(n8452), .B2(n8501), .A(n8389), .ZN(P2_U3274) );
  XNOR2_X1 U9900 ( .A(n8390), .B(n8398), .ZN(n8506) );
  INV_X1 U9901 ( .A(n8412), .ZN(n8393) );
  INV_X1 U9902 ( .A(n8391), .ZN(n8392) );
  AOI21_X1 U9903 ( .B1(n8502), .B2(n8393), .A(n8392), .ZN(n8503) );
  AOI22_X1 U9904 ( .A1(n10001), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n8394), .B2(
        n9993), .ZN(n8395) );
  OAI21_X1 U9905 ( .B1(n8396), .B2(n8415), .A(n8395), .ZN(n8405) );
  INV_X1 U9906 ( .A(n8397), .ZN(n8401) );
  INV_X1 U9907 ( .A(n8398), .ZN(n8400) );
  OAI21_X1 U9908 ( .B1(n8401), .B2(n8400), .A(n8399), .ZN(n8403) );
  AOI222_X1 U9909 ( .A1(n9693), .A2(n8403), .B1(n8402), .B2(n8445), .C1(n8426), 
        .C2(n8443), .ZN(n8505) );
  NOR2_X1 U9910 ( .A1(n8505), .A2(n9706), .ZN(n8404) );
  AOI211_X1 U9911 ( .C1(n8503), .C2(n8450), .A(n8405), .B(n8404), .ZN(n8406)
         );
  OAI21_X1 U9912 ( .B1(n8452), .B2(n8506), .A(n8406), .ZN(P2_U3275) );
  NAND2_X1 U9913 ( .A1(n8407), .A2(n8408), .ZN(n8409) );
  XNOR2_X1 U9914 ( .A(n8409), .B(n8418), .ZN(n8411) );
  AOI222_X1 U9915 ( .A1(n9693), .A2(n8411), .B1(n8410), .B2(n8445), .C1(n8446), 
        .C2(n8443), .ZN(n8512) );
  AOI21_X1 U9916 ( .B1(n8509), .B2(n8428), .A(n8412), .ZN(n8510) );
  INV_X1 U9917 ( .A(n8509), .ZN(n8416) );
  AOI22_X1 U9918 ( .A1(n10001), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n8413), .B2(
        n9993), .ZN(n8414) );
  OAI21_X1 U9919 ( .B1(n8416), .B2(n8415), .A(n8414), .ZN(n8417) );
  AOI21_X1 U9920 ( .B1(n8510), .B2(n8450), .A(n8417), .ZN(n8421) );
  NAND2_X1 U9921 ( .A1(n8419), .A2(n8418), .ZN(n8507) );
  NAND3_X1 U9922 ( .A1(n8508), .A2(n8507), .A3(n9703), .ZN(n8420) );
  OAI211_X1 U9923 ( .C1(n8512), .C2(n9706), .A(n8421), .B(n8420), .ZN(P2_U3276) );
  XOR2_X1 U9924 ( .A(n8422), .B(n8424), .Z(n8518) );
  OAI21_X1 U9925 ( .B1(n8424), .B2(n8423), .A(n8407), .ZN(n8427) );
  AOI222_X1 U9926 ( .A1(n9693), .A2(n8427), .B1(n8426), .B2(n8445), .C1(n8425), 
        .C2(n8443), .ZN(n8517) );
  INV_X1 U9927 ( .A(n8428), .ZN(n8429) );
  AOI211_X1 U9928 ( .C1(n8515), .C2(n8437), .A(n9780), .B(n8429), .ZN(n8514)
         );
  AOI22_X1 U9929 ( .A1(n8514), .A2(n5645), .B1(n9993), .B2(n8430), .ZN(n8431)
         );
  AOI21_X1 U9930 ( .B1(n8517), .B2(n8431), .A(n9706), .ZN(n8432) );
  INV_X1 U9931 ( .A(n8432), .ZN(n8434) );
  AOI22_X1 U9932 ( .A1(n8515), .A2(n9996), .B1(n9706), .B2(
        P2_REG2_REG_19__SCAN_IN), .ZN(n8433) );
  OAI211_X1 U9933 ( .C1(n8518), .C2(n8452), .A(n8434), .B(n8433), .ZN(P2_U3277) );
  XNOR2_X1 U9934 ( .A(n8435), .B(n4825), .ZN(n8523) );
  INV_X1 U9935 ( .A(n8436), .ZN(n8438) );
  AOI21_X1 U9936 ( .B1(n8519), .B2(n8438), .A(n4497), .ZN(n8520) );
  AOI22_X1 U9937 ( .A1(n10001), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n8439), .B2(
        n9993), .ZN(n8440) );
  OAI21_X1 U9938 ( .B1(n8441), .B2(n8415), .A(n8440), .ZN(n8449) );
  OAI21_X1 U9939 ( .B1(n4823), .B2(n4825), .A(n8442), .ZN(n8447) );
  AOI222_X1 U9940 ( .A1(n9693), .A2(n8447), .B1(n8446), .B2(n8445), .C1(n8444), 
        .C2(n8443), .ZN(n8522) );
  NOR2_X1 U9941 ( .A1(n8522), .A2(n9706), .ZN(n8448) );
  AOI211_X1 U9942 ( .C1(n8520), .C2(n8450), .A(n8449), .B(n8448), .ZN(n8451)
         );
  OAI21_X1 U9943 ( .B1(n8523), .B2(n8452), .A(n8451), .ZN(P2_U3278) );
  MUX2_X1 U9944 ( .A(P2_REG1_REG_31__SCAN_IN), .B(n8535), .S(n9810), .Z(
        P2_U3551) );
  NAND3_X1 U9945 ( .A1(n8456), .A2(n9727), .A3(n8455), .ZN(n8458) );
  OAI211_X1 U9946 ( .C1(n8459), .C2(n9788), .A(n8458), .B(n8457), .ZN(n8536)
         );
  MUX2_X1 U9947 ( .A(P2_REG1_REG_30__SCAN_IN), .B(n8536), .S(n9810), .Z(
        P2_U3550) );
  AOI22_X1 U9948 ( .A1(n8461), .A2(n9727), .B1(n9726), .B2(n8460), .ZN(n8462)
         );
  AOI21_X1 U9949 ( .B1(n9726), .B2(n8466), .A(n8465), .ZN(n8467) );
  OAI211_X1 U9950 ( .C1(n8469), .C2(n9731), .A(n8468), .B(n8467), .ZN(n8538)
         );
  MUX2_X1 U9951 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n8538), .S(n9810), .Z(
        P2_U3548) );
  AOI22_X1 U9952 ( .A1(n8471), .A2(n9727), .B1(n9726), .B2(n8470), .ZN(n8472)
         );
  OAI211_X1 U9953 ( .C1(n8474), .C2(n9731), .A(n8473), .B(n8472), .ZN(n8539)
         );
  MUX2_X1 U9954 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n8539), .S(n9810), .Z(
        P2_U3547) );
  AOI211_X1 U9955 ( .C1(n9726), .C2(n8477), .A(n8476), .B(n8475), .ZN(n8478)
         );
  OAI21_X1 U9956 ( .B1(n8479), .B2(n9731), .A(n8478), .ZN(n8540) );
  MUX2_X1 U9957 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n8540), .S(n9810), .Z(
        P2_U3546) );
  AOI21_X1 U9958 ( .B1(n9726), .B2(n8481), .A(n8480), .ZN(n8482) );
  OAI211_X1 U9959 ( .C1(n8484), .C2(n9731), .A(n8483), .B(n8482), .ZN(n8541)
         );
  MUX2_X1 U9960 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n8541), .S(n9810), .Z(
        P2_U3545) );
  INV_X1 U9961 ( .A(n8485), .ZN(n8490) );
  AOI22_X1 U9962 ( .A1(n8487), .A2(n9727), .B1(n9726), .B2(n8486), .ZN(n8488)
         );
  OAI211_X1 U9963 ( .C1(n8490), .C2(n9731), .A(n8489), .B(n8488), .ZN(n8542)
         );
  MUX2_X1 U9964 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n8542), .S(n9810), .Z(
        P2_U3544) );
  OAI22_X1 U9965 ( .A1(n8492), .A2(n9780), .B1(n4503), .B2(n9788), .ZN(n8493)
         );
  NOR2_X1 U9966 ( .A1(n8494), .A2(n8493), .ZN(n8495) );
  NAND2_X1 U9967 ( .A1(n8496), .A2(n8495), .ZN(n8543) );
  MUX2_X1 U9968 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n8543), .S(n9810), .Z(
        P2_U3543) );
  AOI22_X1 U9969 ( .A1(n8498), .A2(n9727), .B1(n9726), .B2(n8497), .ZN(n8499)
         );
  OAI211_X1 U9970 ( .C1(n8501), .C2(n9731), .A(n8500), .B(n8499), .ZN(n8544)
         );
  MUX2_X1 U9971 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n8544), .S(n9810), .Z(
        P2_U3542) );
  AOI22_X1 U9972 ( .A1(n8503), .A2(n9727), .B1(n9726), .B2(n8502), .ZN(n8504)
         );
  OAI211_X1 U9973 ( .C1(n8506), .C2(n9731), .A(n8505), .B(n8504), .ZN(n8545)
         );
  MUX2_X1 U9974 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n8545), .S(n9810), .Z(
        P2_U3541) );
  NAND3_X1 U9975 ( .A1(n8508), .A2(n9793), .A3(n8507), .ZN(n8513) );
  AOI22_X1 U9976 ( .A1(n8510), .A2(n9727), .B1(n9726), .B2(n8509), .ZN(n8511)
         );
  NAND3_X1 U9977 ( .A1(n8513), .A2(n8512), .A3(n8511), .ZN(n8546) );
  MUX2_X1 U9978 ( .A(n8546), .B(P2_REG1_REG_20__SCAN_IN), .S(n9808), .Z(
        P2_U3540) );
  AOI21_X1 U9979 ( .B1(n9726), .B2(n8515), .A(n8514), .ZN(n8516) );
  OAI211_X1 U9980 ( .C1(n8518), .C2(n9731), .A(n8517), .B(n8516), .ZN(n8547)
         );
  MUX2_X1 U9981 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n8547), .S(n9810), .Z(
        P2_U3539) );
  AOI22_X1 U9982 ( .A1(n8520), .A2(n9727), .B1(n9726), .B2(n8519), .ZN(n8521)
         );
  OAI211_X1 U9983 ( .C1(n8523), .C2(n9731), .A(n8522), .B(n8521), .ZN(n8548)
         );
  MUX2_X1 U9984 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n8548), .S(n9810), .Z(
        P2_U3538) );
  AOI211_X1 U9985 ( .C1(n9726), .C2(n8526), .A(n8525), .B(n8524), .ZN(n8527)
         );
  OAI21_X1 U9986 ( .B1(n8528), .B2(n9731), .A(n8527), .ZN(n8549) );
  MUX2_X1 U9987 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n8549), .S(n9810), .Z(
        P2_U3537) );
  NAND3_X1 U9988 ( .A1(n8529), .A2(n9793), .A3(n7784), .ZN(n8534) );
  AOI22_X1 U9989 ( .A1(n8531), .A2(n9727), .B1(n9726), .B2(n8530), .ZN(n8532)
         );
  NAND3_X1 U9990 ( .A1(n8534), .A2(n8533), .A3(n8532), .ZN(n8550) );
  MUX2_X1 U9991 ( .A(n8550), .B(P2_REG1_REG_16__SCAN_IN), .S(n9808), .Z(
        P2_U3536) );
  MUX2_X1 U9992 ( .A(P2_REG0_REG_30__SCAN_IN), .B(n8536), .S(n9796), .Z(
        P2_U3518) );
  MUX2_X1 U9993 ( .A(P2_REG0_REG_29__SCAN_IN), .B(n8537), .S(n9796), .Z(
        P2_U3517) );
  MUX2_X1 U9994 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n8538), .S(n9796), .Z(
        P2_U3516) );
  MUX2_X1 U9995 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n8539), .S(n9796), .Z(
        P2_U3515) );
  MUX2_X1 U9996 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n8540), .S(n9796), .Z(
        P2_U3514) );
  MUX2_X1 U9997 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n8541), .S(n9796), .Z(
        P2_U3513) );
  MUX2_X1 U9998 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n8542), .S(n9796), .Z(
        P2_U3512) );
  MUX2_X1 U9999 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n8543), .S(n9796), .Z(
        P2_U3511) );
  MUX2_X1 U10000 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n8544), .S(n9796), .Z(
        P2_U3510) );
  MUX2_X1 U10001 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n8545), .S(n9796), .Z(
        P2_U3509) );
  MUX2_X1 U10002 ( .A(n8546), .B(P2_REG0_REG_20__SCAN_IN), .S(n9794), .Z(
        P2_U3508) );
  MUX2_X1 U10003 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n8547), .S(n9796), .Z(
        P2_U3507) );
  MUX2_X1 U10004 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n8548), .S(n9796), .Z(
        P2_U3505) );
  MUX2_X1 U10005 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n8549), .S(n9796), .Z(
        P2_U3502) );
  MUX2_X1 U10006 ( .A(n8550), .B(P2_REG0_REG_16__SCAN_IN), .S(n9794), .Z(
        P2_U3499) );
  INV_X1 U10007 ( .A(n8551), .ZN(n9385) );
  NOR4_X1 U10008 ( .A1(n4841), .A2(P2_IR_REG_30__SCAN_IN), .A3(n8552), .A4(
        P2_U3152), .ZN(n8553) );
  AOI21_X1 U10009 ( .B1(n8556), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n8553), .ZN(
        n8554) );
  OAI21_X1 U10010 ( .B1(n9385), .B2(n8049), .A(n8554), .ZN(P2_U3327) );
  INV_X1 U10011 ( .A(n8555), .ZN(n9392) );
  AOI22_X1 U10012 ( .A1(n8557), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_29__SCAN_IN), .B2(n8556), .ZN(n8558) );
  OAI21_X1 U10013 ( .B1(n9392), .B2(n8049), .A(n8558), .ZN(P2_U3329) );
  MUX2_X1 U10014 ( .A(n8560), .B(n9689), .S(P2_STATE_REG_SCAN_IN), .Z(P2_U3358) );
  NAND2_X1 U10015 ( .A1(n8562), .A2(n8561), .ZN(n8564) );
  XNOR2_X1 U10016 ( .A(n8564), .B(n8563), .ZN(n8565) );
  NAND2_X1 U10017 ( .A1(n8565), .A2(n8700), .ZN(n8572) );
  NOR2_X1 U10018 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n8566), .ZN(n9553) );
  INV_X1 U10019 ( .A(n8567), .ZN(n8569) );
  OAI22_X1 U10020 ( .A1(n8707), .A2(n8569), .B1(n8705), .B2(n8568), .ZN(n8570)
         );
  AOI211_X1 U10021 ( .C1(n8710), .C2(n9007), .A(n9553), .B(n8570), .ZN(n8571)
         );
  OAI211_X1 U10022 ( .C1(n9435), .C2(n8713), .A(n8572), .B(n8571), .ZN(
        P1_U3213) );
  INV_X1 U10023 ( .A(n8621), .ZN(n8573) );
  NOR2_X1 U10024 ( .A1(n8622), .A2(n8573), .ZN(n8577) );
  AOI21_X1 U10025 ( .B1(n8574), .B2(n8621), .A(n8575), .ZN(n8576) );
  OAI21_X1 U10026 ( .B1(n8577), .B2(n8576), .A(n8700), .ZN(n8581) );
  AOI22_X1 U10027 ( .A1(n9179), .A2(n8668), .B1(P1_REG3_REG_23__SCAN_IN), .B2(
        P1_U3084), .ZN(n8578) );
  OAI21_X1 U10028 ( .B1(n8707), .B2(n9146), .A(n8578), .ZN(n8579) );
  AOI21_X1 U10029 ( .B1(n8710), .B2(n9125), .A(n8579), .ZN(n8580) );
  OAI211_X1 U10030 ( .C1(n9149), .C2(n8713), .A(n8581), .B(n8580), .ZN(
        P1_U3214) );
  XOR2_X1 U10031 ( .A(n8583), .B(n8582), .Z(n8588) );
  OAI22_X1 U10032 ( .A1(n8592), .A2(n8676), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8584), .ZN(n8586) );
  OAI22_X1 U10033 ( .A1(n8707), .A2(n9207), .B1(n8705), .B2(n9244), .ZN(n8585)
         );
  AOI211_X1 U10034 ( .C1(n9334), .C2(n8680), .A(n8586), .B(n8585), .ZN(n8587)
         );
  OAI21_X1 U10035 ( .B1(n8588), .B2(n8682), .A(n8587), .ZN(P1_U3217) );
  XOR2_X1 U10036 ( .A(n8590), .B(n8589), .Z(n8596) );
  OAI22_X1 U10037 ( .A1(n8592), .A2(n8705), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8591), .ZN(n8594) );
  OAI22_X1 U10038 ( .A1(n9152), .A2(n8676), .B1(n8707), .B2(n9183), .ZN(n8593)
         );
  AOI211_X1 U10039 ( .C1(n9324), .C2(n8680), .A(n8594), .B(n8593), .ZN(n8595)
         );
  OAI21_X1 U10040 ( .B1(n8596), .B2(n8682), .A(n8595), .ZN(P1_U3221) );
  AOI21_X1 U10041 ( .B1(n8598), .B2(n8597), .A(n8686), .ZN(n8603) );
  NAND2_X1 U10042 ( .A1(n9126), .A2(n8710), .ZN(n8600) );
  AOI22_X1 U10043 ( .A1(n9119), .A2(n8690), .B1(P1_REG3_REG_25__SCAN_IN), .B2(
        P1_U3084), .ZN(n8599) );
  OAI211_X1 U10044 ( .C1(n9153), .C2(n8705), .A(n8600), .B(n8599), .ZN(n8601)
         );
  AOI21_X1 U10045 ( .B1(n9304), .B2(n8680), .A(n8601), .ZN(n8602) );
  OAI21_X1 U10046 ( .B1(n8603), .B2(n8682), .A(n8602), .ZN(P1_U3223) );
  INV_X1 U10047 ( .A(n9264), .ZN(n9429) );
  OAI21_X1 U10048 ( .B1(n8606), .B2(n8605), .A(n8604), .ZN(n8607) );
  NAND2_X1 U10049 ( .A1(n8607), .A2(n8700), .ZN(n8611) );
  NOR2_X1 U10050 ( .A1(n8705), .A2(n9260), .ZN(n8609) );
  OAI22_X1 U10051 ( .A1(n8676), .A2(n9259), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9951), .ZN(n8608) );
  AOI211_X1 U10052 ( .C1(n9263), .C2(n8690), .A(n8609), .B(n8608), .ZN(n8610)
         );
  OAI211_X1 U10053 ( .C1(n9429), .C2(n8713), .A(n8611), .B(n8610), .ZN(
        P1_U3224) );
  XOR2_X1 U10054 ( .A(n8613), .B(n8612), .Z(n8619) );
  OAI22_X1 U10055 ( .A1(n8705), .A2(n9243), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8614), .ZN(n8617) );
  INV_X1 U10056 ( .A(n8615), .ZN(n9247) );
  OAI22_X1 U10057 ( .A1(n8707), .A2(n9247), .B1(n8676), .B2(n9244), .ZN(n8616)
         );
  AOI211_X1 U10058 ( .C1(n9347), .C2(n8680), .A(n8617), .B(n8616), .ZN(n8618)
         );
  OAI21_X1 U10059 ( .B1(n8619), .B2(n8682), .A(n8618), .ZN(P1_U3226) );
  AND3_X1 U10060 ( .A1(n8622), .A2(n8621), .A3(n8620), .ZN(n8623) );
  OAI21_X1 U10061 ( .B1(n8624), .B2(n8623), .A(n8700), .ZN(n8629) );
  INV_X1 U10062 ( .A(n8625), .ZN(n9137) );
  AOI22_X1 U10063 ( .A1(n9137), .A2(n8690), .B1(P1_REG3_REG_24__SCAN_IN), .B2(
        P1_U3084), .ZN(n8626) );
  OAI21_X1 U10064 ( .B1(n9164), .B2(n8705), .A(n8626), .ZN(n8627) );
  AOI21_X1 U10065 ( .B1(n9004), .B2(n8710), .A(n8627), .ZN(n8628) );
  OAI211_X1 U10066 ( .C1(n9140), .C2(n8713), .A(n8629), .B(n8628), .ZN(
        P1_U3227) );
  AND2_X1 U10067 ( .A1(n8631), .A2(n8630), .ZN(n8633) );
  OAI21_X1 U10068 ( .B1(n8634), .B2(n8633), .A(n8632), .ZN(n8635) );
  NAND2_X1 U10069 ( .A1(n8635), .A2(n8700), .ZN(n8641) );
  AOI22_X1 U10070 ( .A1(n8668), .A2(n9019), .B1(n8710), .B2(n9017), .ZN(n8640)
         );
  AND2_X1 U10071 ( .A1(P1_U3084), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n9469) );
  NOR2_X1 U10072 ( .A1(n8713), .A2(n8636), .ZN(n8637) );
  AOI211_X1 U10073 ( .C1(n8638), .C2(n8690), .A(n9469), .B(n8637), .ZN(n8639)
         );
  NAND3_X1 U10074 ( .A1(n8641), .A2(n8640), .A3(n8639), .ZN(P1_U3228) );
  NAND2_X1 U10075 ( .A1(n8644), .A2(n8643), .ZN(n8645) );
  XNOR2_X1 U10076 ( .A(n8642), .B(n8645), .ZN(n8650) );
  OAI22_X1 U10077 ( .A1(n9165), .A2(n8676), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8646), .ZN(n8648) );
  OAI22_X1 U10078 ( .A1(n8707), .A2(n9194), .B1(n8677), .B2(n8705), .ZN(n8647)
         );
  AOI211_X1 U10079 ( .C1(n9329), .C2(n8680), .A(n8648), .B(n8647), .ZN(n8649)
         );
  OAI21_X1 U10080 ( .B1(n8650), .B2(n8682), .A(n8649), .ZN(P1_U3231) );
  NAND2_X1 U10081 ( .A1(n8652), .A2(n8651), .ZN(n8653) );
  XOR2_X1 U10082 ( .A(n8654), .B(n8653), .Z(n8660) );
  OAI22_X1 U10083 ( .A1(n9165), .A2(n8705), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8655), .ZN(n8658) );
  OAI22_X1 U10084 ( .A1(n9164), .A2(n8676), .B1(n8707), .B2(n8656), .ZN(n8657)
         );
  AOI211_X1 U10085 ( .C1(n9320), .C2(n8680), .A(n8658), .B(n8657), .ZN(n8659)
         );
  OAI21_X1 U10086 ( .B1(n8660), .B2(n8682), .A(n8659), .ZN(P1_U3233) );
  OAI21_X1 U10087 ( .B1(n8664), .B2(n8661), .A(n8663), .ZN(n8665) );
  NAND2_X1 U10088 ( .A1(n8665), .A2(n8700), .ZN(n8671) );
  AOI22_X1 U10089 ( .A1(n8667), .A2(P1_REG3_REG_2__SCAN_IN), .B1(n8680), .B2(
        n8666), .ZN(n8670) );
  AOI22_X1 U10090 ( .A1(n8668), .A2(n6321), .B1(n8710), .B2(n9019), .ZN(n8669)
         );
  NAND3_X1 U10091 ( .A1(n8671), .A2(n8670), .A3(n8669), .ZN(P1_U3235) );
  XNOR2_X1 U10092 ( .A(n8673), .B(n8672), .ZN(n8674) );
  XNOR2_X1 U10093 ( .A(n8675), .B(n8674), .ZN(n8683) );
  NAND2_X1 U10094 ( .A1(P1_U3084), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n9562) );
  OAI21_X1 U10095 ( .B1(n8677), .B2(n8676), .A(n9562), .ZN(n8679) );
  OAI22_X1 U10096 ( .A1(n8707), .A2(n9224), .B1(n8705), .B2(n9259), .ZN(n8678)
         );
  AOI211_X1 U10097 ( .C1(n9339), .C2(n8680), .A(n8679), .B(n8678), .ZN(n8681)
         );
  OAI21_X1 U10098 ( .B1(n8683), .B2(n8682), .A(n8681), .ZN(P1_U3236) );
  OAI21_X1 U10099 ( .B1(n8686), .B2(n8685), .A(n8684), .ZN(n8687) );
  NAND3_X1 U10100 ( .A1(n8688), .A2(n8700), .A3(n8687), .ZN(n8694) );
  INV_X1 U10101 ( .A(n8689), .ZN(n9109) );
  AOI22_X1 U10102 ( .A1(n9109), .A2(n8690), .B1(P1_REG3_REG_26__SCAN_IN), .B2(
        P1_U3084), .ZN(n8691) );
  OAI21_X1 U10103 ( .B1(n9135), .B2(n8705), .A(n8691), .ZN(n8692) );
  AOI21_X1 U10104 ( .B1(n9003), .B2(n8710), .A(n8692), .ZN(n8693) );
  OAI211_X1 U10105 ( .C1(n9112), .C2(n8713), .A(n8694), .B(n8693), .ZN(
        P1_U3238) );
  INV_X1 U10106 ( .A(n8695), .ZN(n9351) );
  NAND2_X1 U10107 ( .A1(n8696), .A2(n8697), .ZN(n8699) );
  XNOR2_X1 U10108 ( .A(n8699), .B(n8698), .ZN(n8701) );
  NAND2_X1 U10109 ( .A1(n8701), .A2(n8700), .ZN(n8712) );
  INV_X1 U10110 ( .A(n8702), .ZN(n8709) );
  INV_X1 U10111 ( .A(n8703), .ZN(n8706) );
  OAI22_X1 U10112 ( .A1(n8707), .A2(n8706), .B1(n8705), .B2(n8704), .ZN(n8708)
         );
  AOI211_X1 U10113 ( .C1(n8710), .C2(n9006), .A(n8709), .B(n8708), .ZN(n8711)
         );
  OAI211_X1 U10114 ( .C1(n9351), .C2(n8713), .A(n8712), .B(n8711), .ZN(
        P1_U3239) );
  NAND2_X1 U10115 ( .A1(n8551), .A2(n8714), .ZN(n8716) );
  NAND2_X1 U10116 ( .A1(n8718), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(n8715) );
  NAND2_X1 U10117 ( .A1(n8717), .A2(n8714), .ZN(n8720) );
  NAND2_X1 U10118 ( .A1(n8718), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n8719) );
  OR2_X1 U10119 ( .A1(n9279), .A2(n6243), .ZN(n8858) );
  NAND2_X1 U10120 ( .A1(n8858), .A2(n9055), .ZN(n8721) );
  NAND2_X1 U10121 ( .A1(n8724), .A2(n8908), .ZN(n8900) );
  MUX2_X1 U10122 ( .A(n8900), .B(n8725), .S(n8814), .Z(n8726) );
  INV_X1 U10123 ( .A(n8726), .ZN(n8731) );
  MUX2_X1 U10124 ( .A(n8728), .B(n8727), .S(n4445), .Z(n8730) );
  AOI211_X1 U10125 ( .C1(n8732), .C2(n8731), .A(n8730), .B(n8729), .ZN(n8736)
         );
  NAND2_X1 U10126 ( .A1(n8735), .A2(n8733), .ZN(n8963) );
  AND2_X1 U10127 ( .A1(n8744), .A2(n8734), .ZN(n8897) );
  OAI21_X1 U10128 ( .B1(n8736), .B2(n8963), .A(n8897), .ZN(n8738) );
  NAND2_X1 U10129 ( .A1(n8734), .A2(n8903), .ZN(n8830) );
  OAI21_X1 U10130 ( .B1(n8736), .B2(n8830), .A(n8735), .ZN(n8737) );
  INV_X1 U10131 ( .A(n8745), .ZN(n8739) );
  NAND3_X1 U10132 ( .A1(n8746), .A2(n8742), .A3(n8835), .ZN(n8916) );
  OAI21_X1 U10133 ( .B1(n8739), .B2(n8916), .A(n8894), .ZN(n8741) );
  NAND2_X1 U10134 ( .A1(n8741), .A2(n8740), .ZN(n8751) );
  INV_X1 U10135 ( .A(n8742), .ZN(n8743) );
  MUX2_X1 U10136 ( .A(n8751), .B(n8750), .S(n8814), .Z(n8760) );
  NAND2_X1 U10137 ( .A1(n8761), .A2(n8752), .ZN(n8893) );
  INV_X1 U10138 ( .A(n8753), .ZN(n8754) );
  NOR2_X1 U10139 ( .A1(n8893), .A2(n8754), .ZN(n8758) );
  NAND2_X1 U10140 ( .A1(n8763), .A2(n8755), .ZN(n8762) );
  INV_X1 U10141 ( .A(n8756), .ZN(n8757) );
  NOR2_X1 U10142 ( .A1(n8762), .A2(n8757), .ZN(n8914) );
  MUX2_X1 U10143 ( .A(n8758), .B(n8914), .S(n8814), .Z(n8759) );
  OAI21_X1 U10144 ( .B1(n8760), .B2(n8839), .A(n8759), .ZN(n8766) );
  NAND2_X1 U10145 ( .A1(n8762), .A2(n8761), .ZN(n8764) );
  NAND2_X1 U10146 ( .A1(n8893), .A2(n8763), .ZN(n8919) );
  MUX2_X1 U10147 ( .A(n8764), .B(n8919), .S(n8814), .Z(n8765) );
  NAND3_X1 U10148 ( .A1(n8766), .A2(n8846), .A3(n8765), .ZN(n8768) );
  MUX2_X1 U10149 ( .A(n8920), .B(n8924), .S(n8814), .Z(n8767) );
  NAND3_X1 U10150 ( .A1(n8768), .A2(n9269), .A3(n8767), .ZN(n8777) );
  INV_X1 U10151 ( .A(n8774), .ZN(n8769) );
  INV_X1 U10152 ( .A(n8925), .ZN(n8770) );
  MUX2_X1 U10153 ( .A(n8770), .B(n8927), .S(n8814), .Z(n8771) );
  NOR2_X1 U10154 ( .A1(n9241), .A2(n8771), .ZN(n8776) );
  INV_X1 U10155 ( .A(n8772), .ZN(n8773) );
  NAND2_X1 U10156 ( .A1(n8773), .A2(n8778), .ZN(n8879) );
  NAND2_X1 U10157 ( .A1(n8779), .A2(n8774), .ZN(n8928) );
  MUX2_X1 U10158 ( .A(n8879), .B(n8928), .S(n4445), .Z(n8775) );
  NAND2_X1 U10159 ( .A1(n8781), .A2(n8891), .ZN(n8785) );
  INV_X1 U10160 ( .A(n9176), .ZN(n8881) );
  NAND3_X1 U10161 ( .A1(n8881), .A2(n8814), .A3(n8880), .ZN(n8784) );
  NAND2_X1 U10162 ( .A1(n8891), .A2(n8779), .ZN(n8882) );
  NOR2_X1 U10163 ( .A1(n8780), .A2(n8882), .ZN(n8783) );
  AOI22_X1 U10164 ( .A1(n8785), .A2(n8784), .B1(n8783), .B2(n8782), .ZN(n8789)
         );
  AND2_X1 U10165 ( .A1(n8822), .A2(n8790), .ZN(n8878) );
  AND2_X1 U10166 ( .A1(n8797), .A2(n8794), .ZN(n8931) );
  OAI211_X1 U10167 ( .C1(n8890), .C2(n8973), .A(n8786), .B(n8931), .ZN(n8788)
         );
  OAI21_X1 U10168 ( .B1(n4463), .B2(n8887), .A(n8873), .ZN(n8787) );
  MUX2_X1 U10169 ( .A(n8788), .B(n8787), .S(n8814), .Z(n8800) );
  NAND2_X1 U10170 ( .A1(n8789), .A2(n8878), .ZN(n8795) );
  NAND2_X1 U10171 ( .A1(n8790), .A2(n8823), .ZN(n8792) );
  AND2_X1 U10172 ( .A1(n8792), .A2(n8791), .ZN(n8793) );
  NAND2_X1 U10173 ( .A1(n8821), .A2(n8793), .ZN(n8892) );
  NAND2_X1 U10174 ( .A1(n8892), .A2(n8822), .ZN(n8884) );
  NAND4_X1 U10175 ( .A1(n8795), .A2(n6183), .A3(n8794), .A4(n8884), .ZN(n8796)
         );
  AOI21_X1 U10176 ( .B1(n4425), .B2(n8796), .A(n4307), .ZN(n8799) );
  MUX2_X1 U10177 ( .A(n8873), .B(n8797), .S(n8814), .Z(n8798) );
  OAI211_X1 U10178 ( .C1(n8800), .C2(n8799), .A(n9105), .B(n8798), .ZN(n8806)
         );
  INV_X1 U10179 ( .A(n8869), .ZN(n8935) );
  NAND2_X1 U10180 ( .A1(n8803), .A2(n8867), .ZN(n8801) );
  NOR2_X1 U10181 ( .A1(n9300), .A2(n9095), .ZN(n8872) );
  MUX2_X1 U10182 ( .A(n8801), .B(n8872), .S(n8814), .Z(n8802) );
  NAND2_X1 U10183 ( .A1(n8804), .A2(n8803), .ZN(n8871) );
  AND3_X1 U10184 ( .A1(n8871), .A2(n8814), .A3(n8865), .ZN(n8805) );
  AOI211_X1 U10185 ( .C1(n8865), .C2(n8869), .A(n8814), .B(n8807), .ZN(n8810)
         );
  NAND2_X1 U10186 ( .A1(n9055), .A2(n9001), .ZN(n8808) );
  NAND2_X1 U10187 ( .A1(n9279), .A2(n8808), .ZN(n8811) );
  MUX2_X1 U10188 ( .A(n8863), .B(n8866), .S(n8814), .Z(n8809) );
  INV_X1 U10189 ( .A(n9055), .ZN(n8937) );
  NAND2_X1 U10190 ( .A1(n9276), .A2(n8937), .ZN(n8859) );
  INV_X1 U10191 ( .A(n8811), .ZN(n8812) );
  NAND3_X1 U10192 ( .A1(n8859), .A2(n8812), .A3(n8814), .ZN(n8813) );
  INV_X1 U10193 ( .A(n9276), .ZN(n9057) );
  NAND2_X1 U10194 ( .A1(n8816), .A2(n8951), .ZN(n8817) );
  NAND2_X1 U10195 ( .A1(n8822), .A2(n8821), .ZN(n9161) );
  NOR2_X1 U10196 ( .A1(n9176), .A2(n8823), .ZN(n9197) );
  NAND4_X1 U10197 ( .A1(n8827), .A2(n8826), .A3(n8825), .A4(n8824), .ZN(n8829)
         );
  NOR3_X1 U10198 ( .A1(n8829), .A2(n6271), .A3(n8828), .ZN(n8833) );
  INV_X1 U10199 ( .A(n8830), .ZN(n8831) );
  INV_X1 U10200 ( .A(n8963), .ZN(n8910) );
  NAND4_X1 U10201 ( .A1(n8833), .A2(n8832), .A3(n8831), .A4(n8910), .ZN(n8837)
         );
  NAND2_X1 U10202 ( .A1(n8835), .A2(n8834), .ZN(n9584) );
  OR3_X1 U10203 ( .A1(n8837), .A2(n8836), .A3(n9584), .ZN(n8838) );
  NOR3_X1 U10204 ( .A1(n8840), .A2(n8839), .A3(n8838), .ZN(n8841) );
  NAND2_X1 U10205 ( .A1(n8842), .A2(n8841), .ZN(n8843) );
  NOR2_X1 U10206 ( .A1(n8844), .A2(n8843), .ZN(n8845) );
  NAND3_X1 U10207 ( .A1(n9269), .A2(n8846), .A3(n8845), .ZN(n8847) );
  NOR2_X1 U10208 ( .A1(n9241), .A2(n8847), .ZN(n8848) );
  NAND4_X1 U10209 ( .A1(n9197), .A2(n9230), .A3(n9211), .A4(n8848), .ZN(n8849)
         );
  OR3_X1 U10210 ( .A1(n9161), .A2(n9186), .A3(n8849), .ZN(n8850) );
  NOR2_X1 U10211 ( .A1(n9150), .A2(n8850), .ZN(n8852) );
  AND4_X1 U10212 ( .A1(n8853), .A2(n9124), .A3(n8852), .A4(n9132), .ZN(n8854)
         );
  NAND3_X1 U10213 ( .A1(n9069), .A2(n8854), .A3(n9105), .ZN(n8855) );
  NOR2_X1 U10214 ( .A1(n8856), .A2(n8855), .ZN(n8857) );
  NAND2_X1 U10215 ( .A1(n9279), .A2(n6243), .ZN(n8864) );
  NAND3_X1 U10216 ( .A1(n4822), .A2(n8857), .A3(n8864), .ZN(n8860) );
  NAND2_X1 U10217 ( .A1(n8859), .A2(n8858), .ZN(n8984) );
  OR2_X1 U10218 ( .A1(n8860), .A2(n8984), .ZN(n8862) );
  NAND2_X1 U10219 ( .A1(n8862), .A2(n8861), .ZN(n8944) );
  AND2_X1 U10220 ( .A1(n8864), .A2(n8863), .ZN(n8947) );
  AND2_X1 U10221 ( .A1(n8866), .A2(n8865), .ZN(n8877) );
  INV_X1 U10222 ( .A(n8867), .ZN(n8868) );
  AND2_X1 U10223 ( .A1(n8869), .A2(n8868), .ZN(n8870) );
  OR2_X1 U10224 ( .A1(n8871), .A2(n8870), .ZN(n8933) );
  INV_X1 U10225 ( .A(n8872), .ZN(n8874) );
  AND2_X1 U10226 ( .A1(n8874), .A2(n8873), .ZN(n8875) );
  OR2_X1 U10227 ( .A1(n8933), .A2(n8875), .ZN(n8876) );
  AND2_X1 U10228 ( .A1(n8877), .A2(n8876), .ZN(n8981) );
  INV_X1 U10229 ( .A(n8878), .ZN(n8886) );
  INV_X1 U10230 ( .A(n8879), .ZN(n8883) );
  OAI211_X1 U10231 ( .C1(n8883), .C2(n8882), .A(n8881), .B(n8880), .ZN(n8885)
         );
  OAI211_X1 U10232 ( .C1(n8886), .C2(n8885), .A(n8884), .B(n8973), .ZN(n8888)
         );
  NAND2_X1 U10233 ( .A1(n8888), .A2(n8887), .ZN(n8889) );
  NOR2_X1 U10234 ( .A1(n8890), .A2(n8889), .ZN(n8977) );
  NOR2_X1 U10235 ( .A1(n8892), .A2(n4747), .ZN(n8974) );
  INV_X1 U10236 ( .A(n8893), .ZN(n8898) );
  INV_X1 U10237 ( .A(n8894), .ZN(n8895) );
  NOR2_X1 U10238 ( .A1(n8896), .A2(n8895), .ZN(n8915) );
  NAND4_X1 U10239 ( .A1(n8920), .A2(n8898), .A3(n8897), .A4(n8915), .ZN(n8899)
         );
  OR3_X1 U10240 ( .A1(n8928), .A2(n8927), .A3(n8899), .ZN(n8971) );
  INV_X1 U10241 ( .A(n8900), .ZN(n8906) );
  NAND2_X1 U10242 ( .A1(n8901), .A2(n8957), .ZN(n8905) );
  NAND2_X1 U10243 ( .A1(n8903), .A2(n8902), .ZN(n8904) );
  AOI21_X1 U10244 ( .B1(n8906), .B2(n8905), .A(n8904), .ZN(n8913) );
  AND2_X1 U10245 ( .A1(n8908), .A2(n8907), .ZN(n8909) );
  AND3_X1 U10246 ( .A1(n8910), .A2(n8909), .A3(n8962), .ZN(n8961) );
  NAND2_X1 U10247 ( .A1(n8911), .A2(n8961), .ZN(n8912) );
  OAI21_X1 U10248 ( .B1(n8913), .B2(n8963), .A(n8912), .ZN(n8929) );
  INV_X1 U10249 ( .A(n8914), .ZN(n8922) );
  INV_X1 U10250 ( .A(n8915), .ZN(n8918) );
  INV_X1 U10251 ( .A(n8916), .ZN(n8917) );
  NOR2_X1 U10252 ( .A1(n8918), .A2(n8917), .ZN(n8921) );
  OAI211_X1 U10253 ( .C1(n8922), .C2(n8921), .A(n8920), .B(n8919), .ZN(n8923)
         );
  AND3_X1 U10254 ( .A1(n8925), .A2(n8924), .A3(n8923), .ZN(n8926) );
  OR3_X1 U10255 ( .A1(n8928), .A2(n8927), .A3(n8926), .ZN(n8969) );
  OAI21_X1 U10256 ( .B1(n8971), .B2(n8929), .A(n8969), .ZN(n8930) );
  NAND3_X1 U10257 ( .A1(n8974), .A2(n8973), .A3(n8930), .ZN(n8932) );
  INV_X1 U10258 ( .A(n8931), .ZN(n8975) );
  AOI21_X1 U10259 ( .B1(n8977), .B2(n8932), .A(n8975), .ZN(n8934) );
  INV_X1 U10260 ( .A(n8933), .ZN(n8978) );
  OAI21_X1 U10261 ( .B1(n8935), .B2(n8934), .A(n8978), .ZN(n8936) );
  AOI22_X1 U10262 ( .A1(n9279), .A2(n8937), .B1(n8981), .B2(n8936), .ZN(n8938)
         );
  NAND2_X1 U10263 ( .A1(n8947), .A2(n8938), .ZN(n8939) );
  NAND2_X1 U10264 ( .A1(n8939), .A2(n4272), .ZN(n8940) );
  NAND3_X1 U10265 ( .A1(n8940), .A2(n8951), .A3(n4822), .ZN(n8941) );
  NAND3_X1 U10266 ( .A1(n8944), .A2(n9049), .A3(n8941), .ZN(n8943) );
  OAI211_X1 U10267 ( .C1(n8944), .C2(n9049), .A(n8943), .B(n8942), .ZN(n8945)
         );
  NOR2_X1 U10268 ( .A1(n8946), .A2(n8945), .ZN(n9000) );
  INV_X1 U10269 ( .A(n8947), .ZN(n8983) );
  INV_X1 U10270 ( .A(n8948), .ZN(n8952) );
  NAND2_X1 U10271 ( .A1(n6321), .A2(n8949), .ZN(n8950) );
  NAND3_X1 U10272 ( .A1(n8952), .A2(n8951), .A3(n8950), .ZN(n8953) );
  NAND2_X1 U10273 ( .A1(n8954), .A2(n8953), .ZN(n8955) );
  OR2_X1 U10274 ( .A1(n8956), .A2(n8955), .ZN(n8960) );
  INV_X1 U10275 ( .A(n8957), .ZN(n8958) );
  AOI21_X1 U10276 ( .B1(n8960), .B2(n8959), .A(n8958), .ZN(n8968) );
  INV_X1 U10277 ( .A(n8961), .ZN(n8967) );
  INV_X1 U10278 ( .A(n8962), .ZN(n8965) );
  OR3_X1 U10279 ( .A1(n8965), .A2(n8964), .A3(n8963), .ZN(n8966) );
  OAI21_X1 U10280 ( .B1(n8968), .B2(n8967), .A(n8966), .ZN(n8970) );
  OAI21_X1 U10281 ( .B1(n8971), .B2(n8970), .A(n8969), .ZN(n8972) );
  NAND3_X1 U10282 ( .A1(n8974), .A2(n8973), .A3(n8972), .ZN(n8976) );
  AOI21_X1 U10283 ( .B1(n8977), .B2(n8976), .A(n8975), .ZN(n8979) );
  OAI21_X1 U10284 ( .B1(n8979), .B2(n9093), .A(n8978), .ZN(n8980) );
  AND2_X1 U10285 ( .A1(n8981), .A2(n8980), .ZN(n8982) );
  NOR2_X1 U10286 ( .A1(n8983), .A2(n8982), .ZN(n8985) );
  OR2_X1 U10287 ( .A1(n8985), .A2(n8984), .ZN(n8986) );
  NAND2_X1 U10288 ( .A1(n8986), .A2(n4822), .ZN(n8991) );
  NAND3_X1 U10289 ( .A1(n8991), .A2(n9248), .A3(n8987), .ZN(n8989) );
  OAI211_X1 U10290 ( .C1(n8991), .C2(n8990), .A(n8989), .B(n8988), .ZN(n8999)
         );
  NAND4_X1 U10291 ( .A1(n8994), .A2(n8993), .A3(n8992), .A4(n9649), .ZN(n8995)
         );
  OAI211_X1 U10292 ( .C1(n8997), .C2(n8996), .A(n8995), .B(P1_B_REG_SCAN_IN), 
        .ZN(n8998) );
  OAI21_X1 U10293 ( .B1(n9000), .B2(n8999), .A(n8998), .ZN(P1_U3240) );
  MUX2_X1 U10294 ( .A(n9001), .B(P1_DATAO_REG_30__SCAN_IN), .S(n9021), .Z(
        P1_U3585) );
  MUX2_X1 U10295 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n9002), .S(P1_U4006), .Z(
        P1_U3583) );
  MUX2_X1 U10296 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n9003), .S(P1_U4006), .Z(
        P1_U3582) );
  MUX2_X1 U10297 ( .A(n9126), .B(P1_DATAO_REG_26__SCAN_IN), .S(n9021), .Z(
        P1_U3581) );
  MUX2_X1 U10298 ( .A(n9004), .B(P1_DATAO_REG_25__SCAN_IN), .S(n9021), .Z(
        P1_U3580) );
  MUX2_X1 U10299 ( .A(n9125), .B(P1_DATAO_REG_24__SCAN_IN), .S(n9021), .Z(
        P1_U3579) );
  MUX2_X1 U10300 ( .A(n9005), .B(P1_DATAO_REG_23__SCAN_IN), .S(n9021), .Z(
        P1_U3578) );
  MUX2_X1 U10301 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n9179), .S(P1_U4006), .Z(
        P1_U3577) );
  MUX2_X1 U10302 ( .A(n9199), .B(P1_DATAO_REG_21__SCAN_IN), .S(n9021), .Z(
        P1_U3576) );
  MUX2_X1 U10303 ( .A(n9214), .B(P1_DATAO_REG_20__SCAN_IN), .S(n9021), .Z(
        P1_U3575) );
  MUX2_X1 U10304 ( .A(n9232), .B(P1_DATAO_REG_19__SCAN_IN), .S(n9021), .Z(
        P1_U3574) );
  MUX2_X1 U10305 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n9213), .S(P1_U4006), .Z(
        P1_U3573) );
  MUX2_X1 U10306 ( .A(n9234), .B(P1_DATAO_REG_17__SCAN_IN), .S(n9021), .Z(
        P1_U3572) );
  MUX2_X1 U10307 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n9006), .S(P1_U4006), .Z(
        P1_U3571) );
  MUX2_X1 U10308 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n9007), .S(P1_U4006), .Z(
        P1_U3570) );
  MUX2_X1 U10309 ( .A(n9008), .B(P1_DATAO_REG_14__SCAN_IN), .S(n9021), .Z(
        P1_U3569) );
  MUX2_X1 U10310 ( .A(n9009), .B(P1_DATAO_REG_13__SCAN_IN), .S(n9021), .Z(
        P1_U3568) );
  MUX2_X1 U10311 ( .A(n9010), .B(P1_DATAO_REG_12__SCAN_IN), .S(n9021), .Z(
        P1_U3567) );
  MUX2_X1 U10312 ( .A(n9011), .B(P1_DATAO_REG_11__SCAN_IN), .S(n9021), .Z(
        P1_U3566) );
  MUX2_X1 U10313 ( .A(n9012), .B(P1_DATAO_REG_10__SCAN_IN), .S(n9021), .Z(
        P1_U3565) );
  MUX2_X1 U10314 ( .A(n9013), .B(P1_DATAO_REG_9__SCAN_IN), .S(n9021), .Z(
        P1_U3564) );
  MUX2_X1 U10315 ( .A(n9014), .B(P1_DATAO_REG_8__SCAN_IN), .S(n9021), .Z(
        P1_U3563) );
  MUX2_X1 U10316 ( .A(n9015), .B(P1_DATAO_REG_7__SCAN_IN), .S(n9021), .Z(
        P1_U3562) );
  MUX2_X1 U10317 ( .A(n9016), .B(P1_DATAO_REG_6__SCAN_IN), .S(n9021), .Z(
        P1_U3561) );
  MUX2_X1 U10318 ( .A(n9017), .B(P1_DATAO_REG_5__SCAN_IN), .S(n9021), .Z(
        P1_U3560) );
  MUX2_X1 U10319 ( .A(n9018), .B(P1_DATAO_REG_4__SCAN_IN), .S(n9021), .Z(
        P1_U3559) );
  MUX2_X1 U10320 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n9019), .S(P1_U4006), .Z(
        P1_U3558) );
  MUX2_X1 U10321 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n9020), .S(P1_U4006), .Z(
        P1_U3557) );
  MUX2_X1 U10322 ( .A(n6321), .B(P1_DATAO_REG_1__SCAN_IN), .S(n9021), .Z(
        P1_U3556) );
  MUX2_X1 U10323 ( .A(n6314), .B(P1_DATAO_REG_0__SCAN_IN), .S(n9021), .Z(
        P1_U3555) );
  INV_X1 U10324 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n9036) );
  AOI21_X1 U10325 ( .B1(n9027), .B2(P1_REG2_REG_16__SCAN_IN), .A(n9022), .ZN(
        n9025) );
  INV_X1 U10326 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n9842) );
  NOR2_X1 U10327 ( .A1(n9042), .A2(n9842), .ZN(n9023) );
  AOI21_X1 U10328 ( .B1(n9042), .B2(n9842), .A(n9023), .ZN(n9024) );
  NOR2_X1 U10329 ( .A1(n9025), .A2(n9024), .ZN(n9037) );
  AOI211_X1 U10330 ( .C1(n9025), .C2(n9024), .A(n9037), .B(n9563), .ZN(n9034)
         );
  AOI21_X1 U10331 ( .B1(n9027), .B2(P1_REG1_REG_16__SCAN_IN), .A(n9026), .ZN(
        n9029) );
  XNOR2_X1 U10332 ( .A(n9042), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n9028) );
  NOR2_X1 U10333 ( .A1(n9029), .A2(n9028), .ZN(n9041) );
  AOI211_X1 U10334 ( .C1(n9029), .C2(n9028), .A(n9041), .B(n9510), .ZN(n9033)
         );
  INV_X1 U10335 ( .A(n9042), .ZN(n9031) );
  NAND2_X1 U10336 ( .A1(P1_REG3_REG_17__SCAN_IN), .A2(P1_U3084), .ZN(n9030) );
  OAI21_X1 U10337 ( .B1(n9045), .B2(n9031), .A(n9030), .ZN(n9032) );
  NOR3_X1 U10338 ( .A1(n9034), .A2(n9033), .A3(n9032), .ZN(n9035) );
  OAI21_X1 U10339 ( .B1(n9561), .B2(n9036), .A(n9035), .ZN(P1_U3258) );
  AOI21_X1 U10340 ( .B1(n9042), .B2(P1_REG2_REG_17__SCAN_IN), .A(n9037), .ZN(
        n9566) );
  NAND2_X1 U10341 ( .A1(n9569), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n9038) );
  OAI21_X1 U10342 ( .B1(n9569), .B2(P1_REG2_REG_18__SCAN_IN), .A(n9038), .ZN(
        n9565) );
  NOR2_X1 U10343 ( .A1(n9566), .A2(n9565), .ZN(n9564) );
  AOI21_X1 U10344 ( .B1(P1_REG2_REG_18__SCAN_IN), .B2(n9569), .A(n9564), .ZN(
        n9039) );
  XNOR2_X1 U10345 ( .A(P1_REG2_REG_19__SCAN_IN), .B(n9039), .ZN(n9048) );
  INV_X1 U10346 ( .A(n9048), .ZN(n9046) );
  INV_X1 U10347 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n9875) );
  AOI22_X1 U10348 ( .A1(n9569), .A2(P1_REG1_REG_18__SCAN_IN), .B1(n9875), .B2(
        n9040), .ZN(n9572) );
  NAND2_X1 U10349 ( .A1(n9572), .A2(n9571), .ZN(n9570) );
  OAI21_X1 U10350 ( .B1(n9569), .B2(P1_REG1_REG_18__SCAN_IN), .A(n9570), .ZN(
        n9044) );
  INV_X1 U10351 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n9043) );
  XOR2_X1 U10352 ( .A(n9044), .B(n9043), .Z(n9047) );
  AOI22_X1 U10353 ( .A1(n9048), .A2(n9543), .B1(n9574), .B2(n9047), .ZN(n9050)
         );
  MUX2_X1 U10354 ( .A(n9051), .B(n9050), .S(n9049), .Z(n9053) );
  NAND2_X1 U10355 ( .A1(P1_REG3_REG_19__SCAN_IN), .A2(P1_U3084), .ZN(n9052) );
  OAI211_X1 U10356 ( .C1(n4761), .C2(n9561), .A(n9053), .B(n9052), .ZN(
        P1_U3260) );
  NAND2_X1 U10357 ( .A1(n9061), .A2(n9060), .ZN(n9054) );
  XNOR2_X1 U10358 ( .A(n9054), .B(n9276), .ZN(n9278) );
  NAND2_X1 U10359 ( .A1(n9056), .A2(n9055), .ZN(n9281) );
  NOR2_X1 U10360 ( .A1(n9597), .A2(n9281), .ZN(n9063) );
  NOR2_X1 U10361 ( .A1(n9057), .A2(n9599), .ZN(n9058) );
  AOI211_X1 U10362 ( .C1(n9597), .C2(P1_REG2_REG_31__SCAN_IN), .A(n9063), .B(
        n9058), .ZN(n9059) );
  OAI21_X1 U10363 ( .B1(n9278), .B2(n9066), .A(n9059), .ZN(P1_U3261) );
  XNOR2_X1 U10364 ( .A(n9061), .B(n9060), .ZN(n9282) );
  NOR2_X1 U10365 ( .A1(n9609), .A2(n9062), .ZN(n9064) );
  AOI211_X1 U10366 ( .C1(n9279), .C2(n9605), .A(n9064), .B(n9063), .ZN(n9065)
         );
  OAI21_X1 U10367 ( .B1(n9282), .B2(n9066), .A(n9065), .ZN(P1_U3262) );
  AOI21_X1 U10368 ( .B1(n9069), .B2(n9068), .A(n9067), .ZN(n9070) );
  INV_X1 U10369 ( .A(n9070), .ZN(n9292) );
  AND2_X1 U10370 ( .A1(n9072), .A2(n9071), .ZN(n9074) );
  OR2_X1 U10371 ( .A1(n9074), .A2(n9073), .ZN(n9077) );
  OAI22_X1 U10372 ( .A1(n9107), .A2(n6241), .B1(n9075), .B2(n9586), .ZN(n9076)
         );
  AOI21_X1 U10373 ( .B1(n9077), .B2(n9590), .A(n9076), .ZN(n9291) );
  NAND2_X1 U10374 ( .A1(n9078), .A2(n9595), .ZN(n9079) );
  OAI21_X1 U10375 ( .B1(n9609), .B2(n9080), .A(n9079), .ZN(n9081) );
  AOI21_X1 U10376 ( .B1(n9288), .B2(n9605), .A(n9081), .ZN(n9085) );
  AND2_X1 U10377 ( .A1(n9089), .A2(n9288), .ZN(n9082) );
  NOR2_X1 U10378 ( .A1(n9083), .A2(n9082), .ZN(n9289) );
  NAND2_X1 U10379 ( .A1(n9289), .A2(n9604), .ZN(n9084) );
  OAI211_X1 U10380 ( .C1(n9291), .C2(n9597), .A(n9085), .B(n9084), .ZN(n9086)
         );
  INV_X1 U10381 ( .A(n9086), .ZN(n9087) );
  OAI21_X1 U10382 ( .B1(n9292), .B2(n9271), .A(n9087), .ZN(P1_U3263) );
  XNOR2_X1 U10383 ( .A(n9088), .B(n9093), .ZN(n9297) );
  INV_X1 U10384 ( .A(n9089), .ZN(n9090) );
  AOI21_X1 U10385 ( .B1(n9293), .B2(n9108), .A(n9090), .ZN(n9294) );
  AOI22_X1 U10386 ( .A1(n9091), .A2(n9595), .B1(P1_REG2_REG_27__SCAN_IN), .B2(
        n9597), .ZN(n9092) );
  OAI21_X1 U10387 ( .B1(n4554), .B2(n9599), .A(n9092), .ZN(n9101) );
  AOI21_X1 U10388 ( .B1(n9094), .B2(n9093), .A(n6240), .ZN(n9099) );
  OAI22_X1 U10389 ( .A1(n9096), .A2(n9586), .B1(n9095), .B2(n6241), .ZN(n9097)
         );
  AOI21_X1 U10390 ( .B1(n9099), .B2(n9098), .A(n9097), .ZN(n9296) );
  NOR2_X1 U10391 ( .A1(n9296), .A2(n9597), .ZN(n9100) );
  AOI211_X1 U10392 ( .C1(n9604), .C2(n9294), .A(n9101), .B(n9100), .ZN(n9102)
         );
  OAI21_X1 U10393 ( .B1(n9297), .B2(n9271), .A(n9102), .ZN(P1_U3264) );
  XNOR2_X1 U10394 ( .A(n9103), .B(n9105), .ZN(n9302) );
  XOR2_X1 U10395 ( .A(n9105), .B(n9104), .Z(n9106) );
  OAI222_X1 U10396 ( .A1(n9586), .A2(n9107), .B1(n6241), .B2(n9135), .C1(n6240), .C2(n9106), .ZN(n9298) );
  AOI211_X1 U10397 ( .C1(n9300), .C2(n9116), .A(n9664), .B(n4555), .ZN(n9299)
         );
  NAND2_X1 U10398 ( .A1(n9299), .A2(n9169), .ZN(n9111) );
  AOI22_X1 U10399 ( .A1(n9109), .A2(n9595), .B1(P1_REG2_REG_26__SCAN_IN), .B2(
        n9597), .ZN(n9110) );
  OAI211_X1 U10400 ( .C1(n9112), .C2(n9599), .A(n9111), .B(n9110), .ZN(n9113)
         );
  AOI21_X1 U10401 ( .B1(n9298), .B2(n9609), .A(n9113), .ZN(n9114) );
  OAI21_X1 U10402 ( .B1(n9302), .B2(n9271), .A(n9114), .ZN(P1_U3265) );
  XOR2_X1 U10403 ( .A(n9124), .B(n9115), .Z(n9307) );
  INV_X1 U10404 ( .A(n9136), .ZN(n9118) );
  INV_X1 U10405 ( .A(n9116), .ZN(n9117) );
  AOI211_X1 U10406 ( .C1(n9304), .C2(n9118), .A(n9664), .B(n9117), .ZN(n9303)
         );
  AOI22_X1 U10407 ( .A1(n9119), .A2(n9595), .B1(P1_REG2_REG_25__SCAN_IN), .B2(
        n9597), .ZN(n9120) );
  OAI21_X1 U10408 ( .B1(n9121), .B2(n9599), .A(n9120), .ZN(n9129) );
  OAI21_X1 U10409 ( .B1(n9124), .B2(n9123), .A(n9122), .ZN(n9127) );
  AOI222_X1 U10410 ( .A1(n9590), .A2(n9127), .B1(n9126), .B2(n9231), .C1(n9125), .C2(n9233), .ZN(n9306) );
  NOR2_X1 U10411 ( .A1(n9306), .A2(n9597), .ZN(n9128) );
  AOI211_X1 U10412 ( .C1(n9169), .C2(n9303), .A(n9129), .B(n9128), .ZN(n9130)
         );
  OAI21_X1 U10413 ( .B1(n9307), .B2(n9271), .A(n9130), .ZN(P1_U3266) );
  XNOR2_X1 U10414 ( .A(n9131), .B(n9132), .ZN(n9312) );
  XNOR2_X1 U10415 ( .A(n9133), .B(n9132), .ZN(n9134) );
  OAI222_X1 U10416 ( .A1(n9586), .A2(n9135), .B1(n6241), .B2(n9164), .C1(n9134), .C2(n6240), .ZN(n9308) );
  AOI211_X1 U10417 ( .C1(n9310), .C2(n9144), .A(n9664), .B(n9136), .ZN(n9309)
         );
  NAND2_X1 U10418 ( .A1(n9309), .A2(n9169), .ZN(n9139) );
  AOI22_X1 U10419 ( .A1(n9137), .A2(n9595), .B1(P1_REG2_REG_24__SCAN_IN), .B2(
        n9597), .ZN(n9138) );
  OAI211_X1 U10420 ( .C1(n9140), .C2(n9599), .A(n9139), .B(n9138), .ZN(n9141)
         );
  AOI21_X1 U10421 ( .B1(n9308), .B2(n9609), .A(n9141), .ZN(n9142) );
  OAI21_X1 U10422 ( .B1(n9312), .B2(n9271), .A(n9142), .ZN(P1_U3267) );
  XNOR2_X1 U10423 ( .A(n9143), .B(n6183), .ZN(n9317) );
  INV_X1 U10424 ( .A(n9144), .ZN(n9145) );
  AOI21_X1 U10425 ( .B1(n9313), .B2(n9167), .A(n9145), .ZN(n9314) );
  INV_X1 U10426 ( .A(n9146), .ZN(n9147) );
  AOI22_X1 U10427 ( .A1(n9147), .A2(n9595), .B1(P1_REG2_REG_23__SCAN_IN), .B2(
        n9597), .ZN(n9148) );
  OAI21_X1 U10428 ( .B1(n9149), .B2(n9599), .A(n9148), .ZN(n9158) );
  AOI21_X1 U10429 ( .B1(n9151), .B2(n9150), .A(n6240), .ZN(n9156) );
  OAI22_X1 U10430 ( .A1(n9153), .A2(n9586), .B1(n9152), .B2(n6241), .ZN(n9154)
         );
  AOI21_X1 U10431 ( .B1(n9156), .B2(n9155), .A(n9154), .ZN(n9316) );
  NOR2_X1 U10432 ( .A1(n9316), .A2(n9597), .ZN(n9157) );
  AOI211_X1 U10433 ( .C1(n9314), .C2(n9604), .A(n9158), .B(n9157), .ZN(n9159)
         );
  OAI21_X1 U10434 ( .B1(n9317), .B2(n9271), .A(n9159), .ZN(P1_U3268) );
  XNOR2_X1 U10435 ( .A(n9160), .B(n9161), .ZN(n9322) );
  XNOR2_X1 U10436 ( .A(n9162), .B(n9161), .ZN(n9163) );
  OAI222_X1 U10437 ( .A1(n6241), .A2(n9165), .B1(n9586), .B2(n9164), .C1(n9163), .C2(n6240), .ZN(n9318) );
  INV_X1 U10438 ( .A(n9166), .ZN(n9181) );
  INV_X1 U10439 ( .A(n9167), .ZN(n9168) );
  AOI211_X1 U10440 ( .C1(n9320), .C2(n9181), .A(n9664), .B(n9168), .ZN(n9319)
         );
  NAND2_X1 U10441 ( .A1(n9319), .A2(n9169), .ZN(n9172) );
  AOI22_X1 U10442 ( .A1(n9170), .A2(n9595), .B1(P1_REG2_REG_22__SCAN_IN), .B2(
        n9597), .ZN(n9171) );
  OAI211_X1 U10443 ( .C1(n9173), .C2(n9599), .A(n9172), .B(n9171), .ZN(n9174)
         );
  AOI21_X1 U10444 ( .B1(n9318), .B2(n9609), .A(n9174), .ZN(n9175) );
  OAI21_X1 U10445 ( .B1(n9322), .B2(n9271), .A(n9175), .ZN(P1_U3269) );
  OAI21_X1 U10446 ( .B1(n4303), .B2(n9176), .A(n9186), .ZN(n9178) );
  NAND2_X1 U10447 ( .A1(n9178), .A2(n9177), .ZN(n9180) );
  AOI222_X1 U10448 ( .A1(n9590), .A2(n9180), .B1(n9214), .B2(n9233), .C1(n9179), .C2(n9231), .ZN(n9327) );
  INV_X1 U10449 ( .A(n9327), .ZN(n9185) );
  OAI211_X1 U10450 ( .C1(n9182), .C2(n4339), .A(n9181), .B(n9340), .ZN(n9325)
         );
  OAI22_X1 U10451 ( .A1(n9325), .A2(n9248), .B1(n9613), .B2(n9183), .ZN(n9184)
         );
  OAI21_X1 U10452 ( .B1(n9185), .B2(n9184), .A(n9609), .ZN(n9192) );
  AOI22_X1 U10453 ( .A1(n9324), .A2(n9605), .B1(n9597), .B2(
        P1_REG2_REG_21__SCAN_IN), .ZN(n9191) );
  OR2_X1 U10454 ( .A1(n9187), .A2(n9186), .ZN(n9323) );
  NAND3_X1 U10455 ( .A1(n9323), .A2(n9188), .A3(n9189), .ZN(n9190) );
  NAND3_X1 U10456 ( .A1(n9192), .A2(n9191), .A3(n9190), .ZN(P1_U3270) );
  XNOR2_X1 U10457 ( .A(n9193), .B(n9197), .ZN(n9333) );
  AOI21_X1 U10458 ( .B1(n9329), .B2(n9205), .A(n4339), .ZN(n9330) );
  INV_X1 U10459 ( .A(n9194), .ZN(n9195) );
  AOI22_X1 U10460 ( .A1(n9597), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n9195), .B2(
        n9595), .ZN(n9196) );
  OAI21_X1 U10461 ( .B1(n4548), .B2(n9599), .A(n9196), .ZN(n9202) );
  XNOR2_X1 U10462 ( .A(n9198), .B(n9197), .ZN(n9200) );
  AOI222_X1 U10463 ( .A1(n9590), .A2(n9200), .B1(n9199), .B2(n9231), .C1(n9232), .C2(n9233), .ZN(n9332) );
  NOR2_X1 U10464 ( .A1(n9332), .A2(n9597), .ZN(n9201) );
  AOI211_X1 U10465 ( .C1(n9330), .C2(n9604), .A(n9202), .B(n9201), .ZN(n9203)
         );
  OAI21_X1 U10466 ( .B1(n9271), .B2(n9333), .A(n9203), .ZN(P1_U3271) );
  XOR2_X1 U10467 ( .A(n9211), .B(n9204), .Z(n9338) );
  INV_X1 U10468 ( .A(n9205), .ZN(n9206) );
  AOI21_X1 U10469 ( .B1(n9334), .B2(n9221), .A(n9206), .ZN(n9335) );
  INV_X1 U10470 ( .A(n9334), .ZN(n9210) );
  INV_X1 U10471 ( .A(n9207), .ZN(n9208) );
  AOI22_X1 U10472 ( .A1(n9597), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n9208), .B2(
        n9595), .ZN(n9209) );
  OAI21_X1 U10473 ( .B1(n9210), .B2(n9599), .A(n9209), .ZN(n9217) );
  XNOR2_X1 U10474 ( .A(n9212), .B(n9211), .ZN(n9215) );
  AOI222_X1 U10475 ( .A1(n9590), .A2(n9215), .B1(n9214), .B2(n9231), .C1(n9213), .C2(n9233), .ZN(n9337) );
  NOR2_X1 U10476 ( .A1(n9337), .A2(n9597), .ZN(n9216) );
  AOI211_X1 U10477 ( .C1(n9335), .C2(n9604), .A(n9217), .B(n9216), .ZN(n9218)
         );
  OAI21_X1 U10478 ( .B1(n9271), .B2(n9338), .A(n9218), .ZN(P1_U3272) );
  XNOR2_X1 U10479 ( .A(n9220), .B(n9219), .ZN(n9344) );
  INV_X1 U10480 ( .A(n9246), .ZN(n9223) );
  INV_X1 U10481 ( .A(n9221), .ZN(n9222) );
  AOI21_X1 U10482 ( .B1(n9339), .B2(n9223), .A(n9222), .ZN(n9341) );
  INV_X1 U10483 ( .A(n9224), .ZN(n9225) );
  AOI22_X1 U10484 ( .A1(n9597), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n9225), .B2(
        n9595), .ZN(n9226) );
  OAI21_X1 U10485 ( .B1(n9227), .B2(n9599), .A(n9226), .ZN(n9237) );
  OAI21_X1 U10486 ( .B1(n9230), .B2(n9229), .A(n9228), .ZN(n9235) );
  AOI222_X1 U10487 ( .A1(n9590), .A2(n9235), .B1(n9234), .B2(n9233), .C1(n9232), .C2(n9231), .ZN(n9343) );
  NOR2_X1 U10488 ( .A1(n9343), .A2(n9597), .ZN(n9236) );
  AOI211_X1 U10489 ( .C1(n9341), .C2(n9604), .A(n9237), .B(n9236), .ZN(n9238)
         );
  OAI21_X1 U10490 ( .B1(n9271), .B2(n9344), .A(n9238), .ZN(P1_U3273) );
  XNOR2_X1 U10491 ( .A(n9239), .B(n9241), .ZN(n9349) );
  AOI22_X1 U10492 ( .A1(n9347), .A2(n9605), .B1(n9597), .B2(
        P1_REG2_REG_17__SCAN_IN), .ZN(n9252) );
  XOR2_X1 U10493 ( .A(n9241), .B(n9240), .Z(n9242) );
  OAI222_X1 U10494 ( .A1(n9586), .A2(n9244), .B1(n6241), .B2(n9243), .C1(n6240), .C2(n9242), .ZN(n9345) );
  INV_X1 U10495 ( .A(n9245), .ZN(n9262) );
  AOI211_X1 U10496 ( .C1(n9347), .C2(n9262), .A(n9664), .B(n9246), .ZN(n9346)
         );
  INV_X1 U10497 ( .A(n9346), .ZN(n9249) );
  OAI22_X1 U10498 ( .A1(n9249), .A2(n9248), .B1(n9613), .B2(n9247), .ZN(n9250)
         );
  OAI21_X1 U10499 ( .B1(n9345), .B2(n9250), .A(n9609), .ZN(n9251) );
  OAI211_X1 U10500 ( .C1(n9349), .C2(n9271), .A(n9252), .B(n9251), .ZN(
        P1_U3274) );
  OR2_X1 U10501 ( .A1(n9254), .A2(n9253), .ZN(n9256) );
  AND2_X1 U10502 ( .A1(n9256), .A2(n9255), .ZN(n9257) );
  XOR2_X1 U10503 ( .A(n9269), .B(n9257), .Z(n9258) );
  OAI222_X1 U10504 ( .A1(n6241), .A2(n9260), .B1(n9586), .B2(n9259), .C1(n9258), .C2(n6240), .ZN(n9430) );
  OAI211_X1 U10505 ( .C1(n9429), .C2(n4551), .A(n9262), .B(n9340), .ZN(n9428)
         );
  AOI22_X1 U10506 ( .A1(n9597), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n9263), .B2(
        n9595), .ZN(n9266) );
  NAND2_X1 U10507 ( .A1(n9264), .A2(n9605), .ZN(n9265) );
  OAI211_X1 U10508 ( .C1(n9428), .C2(n9267), .A(n9266), .B(n9265), .ZN(n9274)
         );
  INV_X1 U10509 ( .A(n9268), .ZN(n9272) );
  AND2_X1 U10510 ( .A1(n9270), .A2(n9269), .ZN(n9427) );
  NOR3_X1 U10511 ( .A1(n9272), .A2(n9427), .A3(n9271), .ZN(n9273) );
  AOI211_X1 U10512 ( .C1(n9609), .C2(n9430), .A(n9274), .B(n9273), .ZN(n9275)
         );
  INV_X1 U10513 ( .A(n9275), .ZN(P1_U3275) );
  NAND2_X1 U10514 ( .A1(n9276), .A2(n9359), .ZN(n9277) );
  OAI211_X1 U10515 ( .C1(n9278), .C2(n9664), .A(n9277), .B(n9281), .ZN(n9363)
         );
  MUX2_X1 U10516 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n9363), .S(n9362), .Z(
        P1_U3554) );
  NAND2_X1 U10517 ( .A1(n9279), .A2(n9359), .ZN(n9280) );
  OAI211_X1 U10518 ( .C1(n9282), .C2(n9664), .A(n9281), .B(n9280), .ZN(n9364)
         );
  MUX2_X1 U10519 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n9364), .S(n9440), .Z(
        P1_U3553) );
  MUX2_X1 U10520 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n9365), .S(n9440), .Z(
        P1_U3552) );
  AOI22_X1 U10521 ( .A1(n9289), .A2(n9340), .B1(n9359), .B2(n9288), .ZN(n9290)
         );
  OAI211_X1 U10522 ( .C1(n9292), .C2(n9426), .A(n9291), .B(n9290), .ZN(n9366)
         );
  MUX2_X1 U10523 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n9366), .S(n9440), .Z(
        P1_U3551) );
  AOI22_X1 U10524 ( .A1(n9294), .A2(n9340), .B1(n9359), .B2(n9293), .ZN(n9295)
         );
  OAI211_X1 U10525 ( .C1(n9297), .C2(n9426), .A(n9296), .B(n9295), .ZN(n9367)
         );
  MUX2_X1 U10526 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n9367), .S(n9440), .Z(
        P1_U3550) );
  AOI211_X1 U10527 ( .C1(n9359), .C2(n9300), .A(n9299), .B(n9298), .ZN(n9301)
         );
  OAI21_X1 U10528 ( .B1(n9302), .B2(n9426), .A(n9301), .ZN(n9368) );
  MUX2_X1 U10529 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n9368), .S(n9440), .Z(
        P1_U3549) );
  AOI21_X1 U10530 ( .B1(n9359), .B2(n9304), .A(n9303), .ZN(n9305) );
  OAI211_X1 U10531 ( .C1(n9307), .C2(n9426), .A(n9306), .B(n9305), .ZN(n9369)
         );
  MUX2_X1 U10532 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n9369), .S(n9440), .Z(
        P1_U3548) );
  AOI211_X1 U10533 ( .C1(n9359), .C2(n9310), .A(n9309), .B(n9308), .ZN(n9311)
         );
  OAI21_X1 U10534 ( .B1(n9312), .B2(n9426), .A(n9311), .ZN(n9370) );
  MUX2_X1 U10535 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n9370), .S(n9440), .Z(
        P1_U3547) );
  AOI22_X1 U10536 ( .A1(n9314), .A2(n9340), .B1(n9359), .B2(n9313), .ZN(n9315)
         );
  OAI211_X1 U10537 ( .C1(n9317), .C2(n9426), .A(n9316), .B(n9315), .ZN(n9371)
         );
  MUX2_X1 U10538 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n9371), .S(n9440), .Z(
        P1_U3546) );
  AOI211_X1 U10539 ( .C1(n9359), .C2(n9320), .A(n9319), .B(n9318), .ZN(n9321)
         );
  OAI21_X1 U10540 ( .B1(n9322), .B2(n9426), .A(n9321), .ZN(n9372) );
  MUX2_X1 U10541 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n9372), .S(n9440), .Z(
        P1_U3545) );
  INV_X1 U10542 ( .A(n9426), .ZN(n9660) );
  NAND3_X1 U10543 ( .A1(n9323), .A2(n9188), .A3(n9660), .ZN(n9328) );
  NAND2_X1 U10544 ( .A1(n9324), .A2(n9359), .ZN(n9326) );
  NAND4_X1 U10545 ( .A1(n9328), .A2(n9327), .A3(n9326), .A4(n9325), .ZN(n9373)
         );
  MUX2_X1 U10546 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n9373), .S(n9362), .Z(
        P1_U3544) );
  AOI22_X1 U10547 ( .A1(n9330), .A2(n9340), .B1(n9359), .B2(n9329), .ZN(n9331)
         );
  OAI211_X1 U10548 ( .C1(n9333), .C2(n9426), .A(n9332), .B(n9331), .ZN(n9374)
         );
  MUX2_X1 U10549 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n9374), .S(n9362), .Z(
        P1_U3543) );
  AOI22_X1 U10550 ( .A1(n9335), .A2(n9340), .B1(n9359), .B2(n9334), .ZN(n9336)
         );
  OAI211_X1 U10551 ( .C1(n9338), .C2(n9426), .A(n9337), .B(n9336), .ZN(n9375)
         );
  MUX2_X1 U10552 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n9375), .S(n9362), .Z(
        P1_U3542) );
  AOI22_X1 U10553 ( .A1(n9341), .A2(n9340), .B1(n9359), .B2(n9339), .ZN(n9342)
         );
  OAI211_X1 U10554 ( .C1(n9344), .C2(n9426), .A(n9343), .B(n9342), .ZN(n9376)
         );
  MUX2_X1 U10555 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n9376), .S(n9362), .Z(
        P1_U3541) );
  AOI211_X1 U10556 ( .C1(n9359), .C2(n9347), .A(n9346), .B(n9345), .ZN(n9348)
         );
  OAI21_X1 U10557 ( .B1(n9426), .B2(n9349), .A(n9348), .ZN(n9377) );
  MUX2_X1 U10558 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n9377), .S(n9362), .Z(
        P1_U3540) );
  AND2_X1 U10559 ( .A1(n9350), .A2(n9669), .ZN(n9355) );
  OAI22_X1 U10560 ( .A1(n9352), .A2(n9664), .B1(n9351), .B2(n9662), .ZN(n9353)
         );
  MUX2_X1 U10561 ( .A(P1_REG1_REG_15__SCAN_IN), .B(n9378), .S(n9362), .Z(
        P1_U3538) );
  AOI211_X1 U10562 ( .C1(n9359), .C2(n9358), .A(n9357), .B(n9356), .ZN(n9360)
         );
  OAI21_X1 U10563 ( .B1(n9426), .B2(n9361), .A(n9360), .ZN(n9379) );
  MUX2_X1 U10564 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n9379), .S(n9362), .Z(
        P1_U3535) );
  MUX2_X1 U10565 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n9363), .S(n9672), .Z(
        P1_U3522) );
  MUX2_X1 U10566 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n9364), .S(n9672), .Z(
        P1_U3521) );
  MUX2_X1 U10567 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n9366), .S(n9672), .Z(
        P1_U3519) );
  MUX2_X1 U10568 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n9367), .S(n9672), .Z(
        P1_U3518) );
  MUX2_X1 U10569 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n9368), .S(n9672), .Z(
        P1_U3517) );
  MUX2_X1 U10570 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n9369), .S(n9672), .Z(
        P1_U3516) );
  MUX2_X1 U10571 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n9370), .S(n9672), .Z(
        P1_U3515) );
  MUX2_X1 U10572 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n9371), .S(n9672), .Z(
        P1_U3514) );
  MUX2_X1 U10573 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n9372), .S(n9672), .Z(
        P1_U3513) );
  MUX2_X1 U10574 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n9373), .S(n9672), .Z(
        P1_U3512) );
  MUX2_X1 U10575 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n9374), .S(n9672), .Z(
        P1_U3511) );
  MUX2_X1 U10576 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n9375), .S(n9672), .Z(
        P1_U3510) );
  MUX2_X1 U10577 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n9376), .S(n9672), .Z(
        P1_U3508) );
  MUX2_X1 U10578 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n9377), .S(n9672), .Z(
        P1_U3505) );
  MUX2_X1 U10579 ( .A(n9378), .B(P1_REG0_REG_15__SCAN_IN), .S(n9670), .Z(
        P1_U3499) );
  MUX2_X1 U10580 ( .A(P1_REG0_REG_12__SCAN_IN), .B(n9379), .S(n9672), .Z(
        P1_U3490) );
  NOR4_X1 U10581 ( .A1(n9381), .A2(P1_IR_REG_30__SCAN_IN), .A3(n9380), .A4(
        P1_U3084), .ZN(n9382) );
  AOI21_X1 U10582 ( .B1(n9383), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n9382), .ZN(
        n9384) );
  OAI21_X1 U10583 ( .B1(n9385), .B2(n6951), .A(n9384), .ZN(P1_U3322) );
  AOI22_X1 U10584 ( .A1(n9386), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_30__SCAN_IN), .B2(n9389), .ZN(n9387) );
  OAI21_X1 U10585 ( .B1(n9388), .B2(n6951), .A(n9387), .ZN(P1_U3323) );
  AOI22_X1 U10586 ( .A1(n9390), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_29__SCAN_IN), .B2(n9389), .ZN(n9391) );
  OAI21_X1 U10587 ( .B1(n9392), .B2(n6951), .A(n9391), .ZN(P1_U3324) );
  MUX2_X1 U10588 ( .A(n9393), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3353) );
  OAI21_X1 U10589 ( .B1(n9395), .B2(n9662), .A(n9394), .ZN(n9397) );
  AOI211_X1 U10590 ( .C1(n9669), .C2(n9398), .A(n9397), .B(n9396), .ZN(n9400)
         );
  INV_X1 U10591 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n9399) );
  AOI22_X1 U10592 ( .A1(n9672), .A2(n9400), .B1(n9399), .B2(n9670), .ZN(
        P1_U3484) );
  AOI22_X1 U10593 ( .A1(n9440), .A2(n9400), .B1(n6712), .B2(n9676), .ZN(
        P1_U3533) );
  OAI22_X1 U10594 ( .A1(n9402), .A2(n9780), .B1(n9401), .B2(n9788), .ZN(n9403)
         );
  AOI211_X1 U10595 ( .C1(n9405), .C2(n9793), .A(n9404), .B(n9403), .ZN(n9421)
         );
  AOI22_X1 U10596 ( .A1(n9810), .A2(n9421), .B1(n9406), .B2(n9808), .ZN(
        P2_U3535) );
  OAI22_X1 U10597 ( .A1(n9408), .A2(n9780), .B1(n9407), .B2(n9788), .ZN(n9409)
         );
  AOI211_X1 U10598 ( .C1(n9411), .C2(n9793), .A(n9410), .B(n9409), .ZN(n9423)
         );
  AOI22_X1 U10599 ( .A1(n9810), .A2(n9423), .B1(n9412), .B2(n9808), .ZN(
        P2_U3534) );
  INV_X1 U10600 ( .A(n9741), .ZN(n9777) );
  INV_X1 U10601 ( .A(n9413), .ZN(n9418) );
  OAI22_X1 U10602 ( .A1(n9415), .A2(n9780), .B1(n9414), .B2(n9788), .ZN(n9417)
         );
  AOI211_X1 U10603 ( .C1(n9777), .C2(n9418), .A(n9417), .B(n9416), .ZN(n9425)
         );
  AOI22_X1 U10604 ( .A1(n9810), .A2(n9425), .B1(n9419), .B2(n9808), .ZN(
        P2_U3533) );
  INV_X1 U10605 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n9420) );
  AOI22_X1 U10606 ( .A1(n9796), .A2(n9421), .B1(n9420), .B2(n9794), .ZN(
        P2_U3496) );
  INV_X1 U10607 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n9422) );
  AOI22_X1 U10608 ( .A1(n9796), .A2(n9423), .B1(n9422), .B2(n9794), .ZN(
        P2_U3493) );
  INV_X1 U10609 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n9424) );
  AOI22_X1 U10610 ( .A1(n9796), .A2(n9425), .B1(n9424), .B2(n9794), .ZN(
        P2_U3490) );
  NOR2_X1 U10611 ( .A1(n9427), .A2(n9426), .ZN(n9432) );
  OAI21_X1 U10612 ( .B1(n9429), .B2(n9662), .A(n9428), .ZN(n9431) );
  AOI211_X1 U10613 ( .C1(n9432), .C2(n9268), .A(n9431), .B(n9430), .ZN(n9454)
         );
  AOI22_X1 U10614 ( .A1(n9440), .A2(n9454), .B1(n9433), .B2(n9676), .ZN(
        P1_U3539) );
  OAI21_X1 U10615 ( .B1(n9435), .B2(n9662), .A(n9434), .ZN(n9436) );
  AOI211_X1 U10616 ( .C1(n9438), .C2(n9660), .A(n9437), .B(n9436), .ZN(n9456)
         );
  AOI22_X1 U10617 ( .A1(n9440), .A2(n9456), .B1(n9439), .B2(n9676), .ZN(
        P1_U3537) );
  INV_X1 U10618 ( .A(n9441), .ZN(n9446) );
  OAI22_X1 U10619 ( .A1(n9443), .A2(n9664), .B1(n9442), .B2(n9662), .ZN(n9445)
         );
  AOI211_X1 U10620 ( .C1(n9669), .C2(n9446), .A(n9445), .B(n9444), .ZN(n9458)
         );
  AOI22_X1 U10621 ( .A1(n9440), .A2(n9458), .B1(n7004), .B2(n9676), .ZN(
        P1_U3536) );
  OAI22_X1 U10622 ( .A1(n9448), .A2(n9664), .B1(n9447), .B2(n9662), .ZN(n9450)
         );
  AOI211_X1 U10623 ( .C1(n9451), .C2(n9660), .A(n9450), .B(n9449), .ZN(n9460)
         );
  AOI22_X1 U10624 ( .A1(n9362), .A2(n9460), .B1(n9452), .B2(n9676), .ZN(
        P1_U3534) );
  INV_X1 U10625 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n9453) );
  AOI22_X1 U10626 ( .A1(n9672), .A2(n9454), .B1(n9453), .B2(n9670), .ZN(
        P1_U3502) );
  INV_X1 U10627 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n9455) );
  AOI22_X1 U10628 ( .A1(n9672), .A2(n9456), .B1(n9455), .B2(n9670), .ZN(
        P1_U3496) );
  INV_X1 U10629 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n9457) );
  AOI22_X1 U10630 ( .A1(n9672), .A2(n9458), .B1(n9457), .B2(n9670), .ZN(
        P1_U3493) );
  INV_X1 U10631 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n9459) );
  AOI22_X1 U10632 ( .A1(n9672), .A2(n9460), .B1(n9459), .B2(n9670), .ZN(
        P1_U3487) );
  INV_X1 U10633 ( .A(P1_WR_REG_SCAN_IN), .ZN(n9890) );
  XOR2_X1 U10634 ( .A(n9890), .B(P2_WR_REG_SCAN_IN), .Z(U123) );
  INV_X1 U10635 ( .A(P2_RD_REG_SCAN_IN), .ZN(n9939) );
  XOR2_X1 U10636 ( .A(P1_RD_REG_SCAN_IN), .B(n9939), .Z(U126) );
  OAI21_X1 U10637 ( .B1(n9463), .B2(n9462), .A(n9461), .ZN(n9467) );
  OAI21_X1 U10638 ( .B1(n4294), .B2(n9465), .A(n9464), .ZN(n9466) );
  AOI22_X1 U10639 ( .A1(n9574), .A2(n9467), .B1(n9543), .B2(n9466), .ZN(n9472)
         );
  AOI211_X1 U10640 ( .C1(n4360), .C2(n9470), .A(n9469), .B(n9468), .ZN(n9471)
         );
  OAI211_X1 U10641 ( .C1(n9947), .C2(n9561), .A(n9472), .B(n9471), .ZN(
        P1_U3245) );
  INV_X1 U10642 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n9905) );
  AOI211_X1 U10643 ( .C1(n9475), .C2(n9474), .A(n9473), .B(n9510), .ZN(n9476)
         );
  AOI211_X1 U10644 ( .C1(n4360), .C2(n9478), .A(n9477), .B(n9476), .ZN(n9484)
         );
  OAI21_X1 U10645 ( .B1(n9481), .B2(n9480), .A(n9479), .ZN(n9482) );
  NAND2_X1 U10646 ( .A1(n9543), .A2(n9482), .ZN(n9483) );
  OAI211_X1 U10647 ( .C1(n9561), .C2(n9905), .A(n9484), .B(n9483), .ZN(
        P1_U3246) );
  AOI211_X1 U10648 ( .C1(n9487), .C2(n9486), .A(n9485), .B(n9563), .ZN(n9488)
         );
  AOI211_X1 U10649 ( .C1(n4360), .C2(n9490), .A(n9489), .B(n9488), .ZN(n9496)
         );
  OAI21_X1 U10650 ( .B1(n9493), .B2(n9492), .A(n9491), .ZN(n9494) );
  AOI22_X1 U10651 ( .A1(n9573), .A2(P1_ADDR_REG_6__SCAN_IN), .B1(n9574), .B2(
        n9494), .ZN(n9495) );
  NAND2_X1 U10652 ( .A1(n9496), .A2(n9495), .ZN(P1_U3247) );
  AOI21_X1 U10653 ( .B1(n4360), .B2(n9498), .A(n9497), .ZN(n9508) );
  OAI21_X1 U10654 ( .B1(n9501), .B2(n9500), .A(n9499), .ZN(n9506) );
  OAI21_X1 U10655 ( .B1(n9504), .B2(n9503), .A(n9502), .ZN(n9505) );
  AOI22_X1 U10656 ( .A1(n9506), .A2(n9574), .B1(n9505), .B2(n9543), .ZN(n9507)
         );
  OAI211_X1 U10657 ( .C1(n9561), .C2(n9509), .A(n9508), .B(n9507), .ZN(
        P1_U3248) );
  AOI211_X1 U10658 ( .C1(n9513), .C2(n9512), .A(n9511), .B(n9510), .ZN(n9514)
         );
  AOI211_X1 U10659 ( .C1(n4360), .C2(n9516), .A(n9515), .B(n9514), .ZN(n9522)
         );
  OAI21_X1 U10660 ( .B1(n9519), .B2(n9518), .A(n9517), .ZN(n9520) );
  AOI22_X1 U10661 ( .A1(n9520), .A2(n9543), .B1(n9573), .B2(
        P1_ADDR_REG_8__SCAN_IN), .ZN(n9521) );
  NAND2_X1 U10662 ( .A1(n9522), .A2(n9521), .ZN(P1_U3249) );
  AOI211_X1 U10663 ( .C1(n9525), .C2(n9524), .A(n9523), .B(n9563), .ZN(n9526)
         );
  AOI211_X1 U10664 ( .C1(n4360), .C2(n9528), .A(n9527), .B(n9526), .ZN(n9534)
         );
  OAI21_X1 U10665 ( .B1(n9531), .B2(n9530), .A(n9529), .ZN(n9532) );
  NAND2_X1 U10666 ( .A1(n9532), .A2(n9574), .ZN(n9533) );
  OAI211_X1 U10667 ( .C1(n10023), .C2(n9561), .A(n9534), .B(n9533), .ZN(
        P1_U3250) );
  INV_X1 U10668 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n9548) );
  AOI21_X1 U10669 ( .B1(n4360), .B2(n9536), .A(n9535), .ZN(n9547) );
  OAI21_X1 U10670 ( .B1(n9539), .B2(n9538), .A(n9537), .ZN(n9545) );
  OAI21_X1 U10671 ( .B1(n9542), .B2(n9541), .A(n9540), .ZN(n9544) );
  AOI22_X1 U10672 ( .A1(n9545), .A2(n9574), .B1(n9544), .B2(n9543), .ZN(n9546)
         );
  OAI211_X1 U10673 ( .C1(n9561), .C2(n9548), .A(n9547), .B(n9546), .ZN(
        P1_U3252) );
  INV_X1 U10674 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n9966) );
  AOI211_X1 U10675 ( .C1(n9551), .C2(n9550), .A(n9549), .B(n9563), .ZN(n9552)
         );
  AOI211_X1 U10676 ( .C1(n4360), .C2(n9554), .A(n9553), .B(n9552), .ZN(n9560)
         );
  OAI21_X1 U10677 ( .B1(n9557), .B2(n9556), .A(n9555), .ZN(n9558) );
  NAND2_X1 U10678 ( .A1(n9558), .A2(n9574), .ZN(n9559) );
  OAI211_X1 U10679 ( .C1(n9561), .C2(n9966), .A(n9560), .B(n9559), .ZN(
        P1_U3255) );
  INV_X1 U10680 ( .A(n9562), .ZN(n9568) );
  AOI211_X1 U10681 ( .C1(n9566), .C2(n9565), .A(n9564), .B(n9563), .ZN(n9567)
         );
  AOI211_X1 U10682 ( .C1(n9569), .C2(n4360), .A(n9568), .B(n9567), .ZN(n9577)
         );
  OAI21_X1 U10683 ( .B1(n9572), .B2(n9571), .A(n9570), .ZN(n9575) );
  AOI22_X1 U10684 ( .A1(n9575), .A2(n9574), .B1(n9573), .B2(
        P1_ADDR_REG_18__SCAN_IN), .ZN(n9576) );
  NAND2_X1 U10685 ( .A1(n9577), .A2(n9576), .ZN(P1_U3259) );
  XNOR2_X1 U10686 ( .A(n9578), .B(n9584), .ZN(n9594) );
  INV_X1 U10687 ( .A(n9594), .ZN(n9668) );
  NOR2_X1 U10688 ( .A1(n9579), .A2(n9663), .ZN(n9580) );
  OR2_X1 U10689 ( .A1(n9581), .A2(n9580), .ZN(n9665) );
  INV_X1 U10690 ( .A(n9665), .ZN(n9582) );
  AOI22_X1 U10691 ( .A1(n9668), .A2(n9583), .B1(n9604), .B2(n9582), .ZN(n9602)
         );
  XNOR2_X1 U10692 ( .A(n9585), .B(n9584), .ZN(n9591) );
  OAI22_X1 U10693 ( .A1(n9588), .A2(n6241), .B1(n9587), .B2(n9586), .ZN(n9589)
         );
  AOI21_X1 U10694 ( .B1(n9591), .B2(n9590), .A(n9589), .ZN(n9592) );
  OAI21_X1 U10695 ( .B1(n9594), .B2(n9593), .A(n9592), .ZN(n9666) );
  AOI22_X1 U10696 ( .A1(n9597), .A2(P1_REG2_REG_9__SCAN_IN), .B1(n9596), .B2(
        n9595), .ZN(n9598) );
  OAI21_X1 U10697 ( .B1(n9663), .B2(n9599), .A(n9598), .ZN(n9600) );
  AOI21_X1 U10698 ( .B1(n9666), .B2(n9609), .A(n9600), .ZN(n9601) );
  NAND2_X1 U10699 ( .A1(n9602), .A2(n9601), .ZN(P1_U3282) );
  INV_X1 U10700 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n9608) );
  NAND2_X1 U10701 ( .A1(n9603), .A2(n9609), .ZN(n9607) );
  OAI21_X1 U10702 ( .B1(n9605), .B2(n9604), .A(n6311), .ZN(n9606) );
  OAI211_X1 U10703 ( .C1(n9609), .C2(n9608), .A(n9607), .B(n9606), .ZN(n9610)
         );
  INV_X1 U10704 ( .A(n9610), .ZN(n9611) );
  OAI21_X1 U10705 ( .B1(n9613), .B2(n9612), .A(n9611), .ZN(P1_U3291) );
  INV_X1 U10706 ( .A(n9614), .ZN(n9615) );
  NOR2_X4 U10707 ( .A1(n9645), .A2(n9615), .ZN(n9642) );
  INV_X1 U10708 ( .A(P1_D_REG_31__SCAN_IN), .ZN(n9616) );
  NOR2_X1 U10709 ( .A1(n9642), .A2(n9616), .ZN(P1_U3292) );
  INV_X1 U10710 ( .A(P1_D_REG_30__SCAN_IN), .ZN(n9617) );
  NOR2_X1 U10711 ( .A1(n9642), .A2(n9617), .ZN(P1_U3293) );
  INV_X1 U10712 ( .A(P1_D_REG_29__SCAN_IN), .ZN(n9918) );
  NOR2_X1 U10713 ( .A1(n9642), .A2(n9918), .ZN(P1_U3294) );
  INV_X1 U10714 ( .A(P1_D_REG_28__SCAN_IN), .ZN(n9917) );
  NOR2_X1 U10715 ( .A1(n9642), .A2(n9917), .ZN(P1_U3295) );
  INV_X1 U10716 ( .A(P1_D_REG_27__SCAN_IN), .ZN(n9618) );
  NOR2_X1 U10717 ( .A1(n9642), .A2(n9618), .ZN(P1_U3296) );
  INV_X1 U10718 ( .A(P1_D_REG_26__SCAN_IN), .ZN(n9619) );
  NOR2_X1 U10719 ( .A1(n9642), .A2(n9619), .ZN(P1_U3297) );
  INV_X1 U10720 ( .A(P1_D_REG_25__SCAN_IN), .ZN(n9620) );
  NOR2_X1 U10721 ( .A1(n9642), .A2(n9620), .ZN(P1_U3298) );
  INV_X1 U10722 ( .A(P1_D_REG_24__SCAN_IN), .ZN(n9621) );
  NOR2_X1 U10723 ( .A1(n9642), .A2(n9621), .ZN(P1_U3299) );
  INV_X1 U10724 ( .A(P1_D_REG_23__SCAN_IN), .ZN(n9622) );
  NOR2_X1 U10725 ( .A1(n9642), .A2(n9622), .ZN(P1_U3300) );
  INV_X1 U10726 ( .A(P1_D_REG_22__SCAN_IN), .ZN(n9845) );
  NOR2_X1 U10727 ( .A1(n9642), .A2(n9845), .ZN(P1_U3301) );
  INV_X1 U10728 ( .A(P1_D_REG_21__SCAN_IN), .ZN(n9623) );
  NOR2_X1 U10729 ( .A1(n9642), .A2(n9623), .ZN(P1_U3302) );
  INV_X1 U10730 ( .A(P1_D_REG_20__SCAN_IN), .ZN(n9624) );
  NOR2_X1 U10731 ( .A1(n9642), .A2(n9624), .ZN(P1_U3303) );
  INV_X1 U10732 ( .A(P1_D_REG_19__SCAN_IN), .ZN(n9625) );
  NOR2_X1 U10733 ( .A1(n9642), .A2(n9625), .ZN(P1_U3304) );
  INV_X1 U10734 ( .A(P1_D_REG_18__SCAN_IN), .ZN(n9626) );
  NOR2_X1 U10735 ( .A1(n9642), .A2(n9626), .ZN(P1_U3305) );
  INV_X1 U10736 ( .A(P1_D_REG_17__SCAN_IN), .ZN(n9627) );
  NOR2_X1 U10737 ( .A1(n9642), .A2(n9627), .ZN(P1_U3306) );
  INV_X1 U10738 ( .A(P1_D_REG_16__SCAN_IN), .ZN(n9628) );
  NOR2_X1 U10739 ( .A1(n9642), .A2(n9628), .ZN(P1_U3307) );
  INV_X1 U10740 ( .A(P1_D_REG_15__SCAN_IN), .ZN(n9629) );
  NOR2_X1 U10741 ( .A1(n9642), .A2(n9629), .ZN(P1_U3308) );
  INV_X1 U10742 ( .A(P1_D_REG_14__SCAN_IN), .ZN(n9630) );
  NOR2_X1 U10743 ( .A1(n9642), .A2(n9630), .ZN(P1_U3309) );
  INV_X1 U10744 ( .A(P1_D_REG_13__SCAN_IN), .ZN(n9631) );
  NOR2_X1 U10745 ( .A1(n9642), .A2(n9631), .ZN(P1_U3310) );
  INV_X1 U10746 ( .A(P1_D_REG_12__SCAN_IN), .ZN(n9632) );
  NOR2_X1 U10747 ( .A1(n9642), .A2(n9632), .ZN(P1_U3311) );
  INV_X1 U10748 ( .A(P1_D_REG_11__SCAN_IN), .ZN(n9633) );
  NOR2_X1 U10749 ( .A1(n9642), .A2(n9633), .ZN(P1_U3312) );
  INV_X1 U10750 ( .A(P1_D_REG_10__SCAN_IN), .ZN(n9634) );
  NOR2_X1 U10751 ( .A1(n9642), .A2(n9634), .ZN(P1_U3313) );
  INV_X1 U10752 ( .A(P1_D_REG_9__SCAN_IN), .ZN(n9635) );
  NOR2_X1 U10753 ( .A1(n9642), .A2(n9635), .ZN(P1_U3314) );
  INV_X1 U10754 ( .A(P1_D_REG_8__SCAN_IN), .ZN(n9636) );
  NOR2_X1 U10755 ( .A1(n9642), .A2(n9636), .ZN(P1_U3315) );
  INV_X1 U10756 ( .A(P1_D_REG_7__SCAN_IN), .ZN(n9911) );
  NOR2_X1 U10757 ( .A1(n9642), .A2(n9911), .ZN(P1_U3316) );
  INV_X1 U10758 ( .A(P1_D_REG_6__SCAN_IN), .ZN(n9637) );
  NOR2_X1 U10759 ( .A1(n9642), .A2(n9637), .ZN(P1_U3317) );
  INV_X1 U10760 ( .A(P1_D_REG_5__SCAN_IN), .ZN(n9638) );
  NOR2_X1 U10761 ( .A1(n9642), .A2(n9638), .ZN(P1_U3318) );
  INV_X1 U10762 ( .A(P1_D_REG_4__SCAN_IN), .ZN(n9639) );
  NOR2_X1 U10763 ( .A1(n9642), .A2(n9639), .ZN(P1_U3319) );
  INV_X1 U10764 ( .A(P1_D_REG_3__SCAN_IN), .ZN(n9640) );
  NOR2_X1 U10765 ( .A1(n9642), .A2(n9640), .ZN(P1_U3320) );
  INV_X1 U10766 ( .A(P1_D_REG_2__SCAN_IN), .ZN(n9641) );
  NOR2_X1 U10767 ( .A1(n9642), .A2(n9641), .ZN(P1_U3321) );
  INV_X1 U10768 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n9644) );
  AOI21_X1 U10769 ( .B1(n9645), .B2(n9644), .A(n9643), .ZN(P1_U3440) );
  INV_X1 U10770 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n9648) );
  NAND2_X1 U10771 ( .A1(n9646), .A2(n9649), .ZN(n9647) );
  OAI21_X1 U10772 ( .B1(n9649), .B2(n9648), .A(n9647), .ZN(P1_U3441) );
  OAI22_X1 U10773 ( .A1(n9651), .A2(n9664), .B1(n9650), .B2(n9662), .ZN(n9653)
         );
  AOI211_X1 U10774 ( .C1(n9669), .C2(n9654), .A(n9653), .B(n9652), .ZN(n9673)
         );
  INV_X1 U10775 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n9655) );
  AOI22_X1 U10776 ( .A1(n9672), .A2(n9673), .B1(n9655), .B2(n9670), .ZN(
        P1_U3463) );
  OAI21_X1 U10777 ( .B1(n9657), .B2(n9662), .A(n9656), .ZN(n9659) );
  AOI211_X1 U10778 ( .C1(n9661), .C2(n9660), .A(n9659), .B(n9658), .ZN(n9675)
         );
  INV_X1 U10779 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n9924) );
  AOI22_X1 U10780 ( .A1(n9672), .A2(n9675), .B1(n9924), .B2(n9670), .ZN(
        P1_U3469) );
  OAI22_X1 U10781 ( .A1(n9665), .A2(n9664), .B1(n9663), .B2(n9662), .ZN(n9667)
         );
  AOI211_X1 U10782 ( .C1(n9669), .C2(n9668), .A(n9667), .B(n9666), .ZN(n9678)
         );
  INV_X1 U10783 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n9671) );
  AOI22_X1 U10784 ( .A1(n9672), .A2(n9678), .B1(n9671), .B2(n9670), .ZN(
        P1_U3481) );
  AOI22_X1 U10785 ( .A1(n9362), .A2(n9673), .B1(n6645), .B2(n9676), .ZN(
        P1_U3526) );
  INV_X1 U10786 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n9674) );
  AOI22_X1 U10787 ( .A1(n9362), .A2(n9675), .B1(n9674), .B2(n9676), .ZN(
        P1_U3528) );
  INV_X1 U10788 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n9677) );
  AOI22_X1 U10789 ( .A1(n9362), .A2(n9678), .B1(n9677), .B2(n9676), .ZN(
        P1_U3532) );
  AOI22_X1 U10790 ( .A1(n9680), .A2(P2_REG2_REG_0__SCAN_IN), .B1(
        P2_REG1_REG_0__SCAN_IN), .B2(n9679), .ZN(n9688) );
  AOI22_X1 U10791 ( .A1(n9681), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3152), .ZN(n9687) );
  OAI22_X1 U10792 ( .A1(n9683), .A2(P2_REG2_REG_0__SCAN_IN), .B1(
        P2_REG1_REG_0__SCAN_IN), .B2(n9682), .ZN(n9685) );
  OAI21_X1 U10793 ( .B1(n9685), .B2(n9684), .A(n9689), .ZN(n9686) );
  OAI211_X1 U10794 ( .C1(n9689), .C2(n9688), .A(n9687), .B(n9686), .ZN(
        P2_U3245) );
  XNOR2_X1 U10795 ( .A(n9691), .B(n7553), .ZN(n9694) );
  AOI21_X1 U10796 ( .B1(n9694), .B2(n9693), .A(n9692), .ZN(n9789) );
  AOI222_X1 U10797 ( .A1(n9786), .A2(n9996), .B1(P2_REG2_REG_12__SCAN_IN), 
        .B2(n9706), .C1(n9993), .C2(n9695), .ZN(n9705) );
  OAI21_X1 U10798 ( .B1(n9697), .B2(n7553), .A(n9696), .ZN(n9792) );
  AOI21_X1 U10799 ( .B1(n9698), .B2(n9786), .A(n9780), .ZN(n9700) );
  NAND2_X1 U10800 ( .A1(n9700), .A2(n9699), .ZN(n9787) );
  INV_X1 U10801 ( .A(n9787), .ZN(n9701) );
  AOI22_X1 U10802 ( .A1(n9792), .A2(n9703), .B1(n9702), .B2(n9701), .ZN(n9704)
         );
  OAI211_X1 U10803 ( .C1(n9706), .C2(n9789), .A(n9705), .B(n9704), .ZN(
        P2_U3284) );
  AND2_X1 U10804 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n9712), .ZN(P2_U3297) );
  AND2_X1 U10805 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n9712), .ZN(P2_U3298) );
  AND2_X1 U10806 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n9712), .ZN(P2_U3299) );
  AND2_X1 U10807 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n9712), .ZN(P2_U3300) );
  AND2_X1 U10808 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n9712), .ZN(P2_U3301) );
  AND2_X1 U10809 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n9712), .ZN(P2_U3302) );
  AND2_X1 U10810 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n9712), .ZN(P2_U3303) );
  AND2_X1 U10811 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n9712), .ZN(P2_U3304) );
  AND2_X1 U10812 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n9712), .ZN(P2_U3305) );
  INV_X1 U10813 ( .A(P2_D_REG_22__SCAN_IN), .ZN(n9949) );
  NOR2_X1 U10814 ( .A1(n9709), .A2(n9949), .ZN(P2_U3306) );
  AND2_X1 U10815 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n9712), .ZN(P2_U3307) );
  AND2_X1 U10816 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n9712), .ZN(P2_U3308) );
  AND2_X1 U10817 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n9712), .ZN(P2_U3309) );
  AND2_X1 U10818 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n9712), .ZN(P2_U3310) );
  AND2_X1 U10819 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n9712), .ZN(P2_U3311) );
  AND2_X1 U10820 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n9712), .ZN(P2_U3312) );
  AND2_X1 U10821 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n9712), .ZN(P2_U3313) );
  AND2_X1 U10822 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n9712), .ZN(P2_U3314) );
  INV_X1 U10823 ( .A(P2_D_REG_13__SCAN_IN), .ZN(n9903) );
  NOR2_X1 U10824 ( .A1(n9709), .A2(n9903), .ZN(P2_U3315) );
  AND2_X1 U10825 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n9712), .ZN(P2_U3316) );
  INV_X1 U10826 ( .A(P2_D_REG_11__SCAN_IN), .ZN(n9886) );
  NOR2_X1 U10827 ( .A1(n9709), .A2(n9886), .ZN(P2_U3317) );
  AND2_X1 U10828 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n9712), .ZN(P2_U3318) );
  AND2_X1 U10829 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n9712), .ZN(P2_U3319) );
  AND2_X1 U10830 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n9712), .ZN(P2_U3320) );
  AND2_X1 U10831 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n9712), .ZN(P2_U3321) );
  AND2_X1 U10832 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n9712), .ZN(P2_U3322) );
  AND2_X1 U10833 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n9712), .ZN(P2_U3323) );
  AND2_X1 U10834 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n9712), .ZN(P2_U3324) );
  AND2_X1 U10835 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n9712), .ZN(P2_U3325) );
  AND2_X1 U10836 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n9712), .ZN(P2_U3326) );
  AOI22_X1 U10837 ( .A1(n9711), .A2(n9712), .B1(n9714), .B2(n9710), .ZN(
        P2_U3437) );
  AOI22_X1 U10838 ( .A1(n9714), .A2(n9713), .B1(n9978), .B2(n9712), .ZN(
        P2_U3438) );
  OAI22_X1 U10839 ( .A1(n9716), .A2(n9731), .B1(n9715), .B2(n4505), .ZN(n9717)
         );
  NOR2_X1 U10840 ( .A1(n9718), .A2(n9717), .ZN(n9798) );
  INV_X1 U10841 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n9719) );
  AOI22_X1 U10842 ( .A1(n9796), .A2(n9798), .B1(n9719), .B2(n9794), .ZN(
        P2_U3451) );
  OAI21_X1 U10843 ( .B1(n6875), .B2(n9788), .A(n9720), .ZN(n9722) );
  AOI211_X1 U10844 ( .C1(n9723), .C2(n9793), .A(n9722), .B(n9721), .ZN(n9799)
         );
  INV_X1 U10845 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n9724) );
  AOI22_X1 U10846 ( .A1(n9796), .A2(n9799), .B1(n9724), .B2(n9794), .ZN(
        P2_U3457) );
  AOI22_X1 U10847 ( .A1(n9728), .A2(n9727), .B1(n9726), .B2(n9725), .ZN(n9729)
         );
  OAI211_X1 U10848 ( .C1(n9732), .C2(n9731), .A(n9730), .B(n9729), .ZN(n9733)
         );
  INV_X1 U10849 ( .A(n9733), .ZN(n9801) );
  INV_X1 U10850 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n9734) );
  AOI22_X1 U10851 ( .A1(n9796), .A2(n9801), .B1(n9734), .B2(n9794), .ZN(
        P2_U3463) );
  OAI22_X1 U10852 ( .A1(n9736), .A2(n9780), .B1(n9735), .B2(n9788), .ZN(n9738)
         );
  AOI211_X1 U10853 ( .C1(n9793), .C2(n9739), .A(n9738), .B(n9737), .ZN(n9803)
         );
  INV_X1 U10854 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n9740) );
  AOI22_X1 U10855 ( .A1(n9796), .A2(n9803), .B1(n9740), .B2(n9794), .ZN(
        P2_U3472) );
  NOR2_X1 U10856 ( .A1(n9742), .A2(n9741), .ZN(n9746) );
  OAI22_X1 U10857 ( .A1(n9744), .A2(n9780), .B1(n9743), .B2(n9788), .ZN(n9745)
         );
  NOR3_X1 U10858 ( .A1(n9747), .A2(n9746), .A3(n9745), .ZN(n9804) );
  INV_X1 U10859 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n9748) );
  AOI22_X1 U10860 ( .A1(n9796), .A2(n9804), .B1(n9748), .B2(n9794), .ZN(
        P2_U3475) );
  XNOR2_X1 U10861 ( .A(n9750), .B(n9749), .ZN(n10006) );
  NAND3_X1 U10862 ( .A1(n7405), .A2(n9752), .A3(n9751), .ZN(n9754) );
  AOI21_X1 U10863 ( .B1(n9755), .B2(n9754), .A(n9753), .ZN(n9761) );
  OAI22_X1 U10864 ( .A1(n9759), .A2(n9758), .B1(n9757), .B2(n9756), .ZN(n9760)
         );
  OR2_X1 U10865 ( .A1(n9761), .A2(n9760), .ZN(n9762) );
  AOI21_X1 U10866 ( .B1(n10006), .B2(n9763), .A(n9762), .ZN(n10002) );
  NOR2_X1 U10867 ( .A1(n9764), .A2(n9767), .ZN(n9765) );
  OR2_X1 U10868 ( .A1(n9766), .A2(n9765), .ZN(n10000) );
  OAI22_X1 U10869 ( .A1(n10000), .A2(n9780), .B1(n9767), .B2(n9788), .ZN(n9768) );
  AOI21_X1 U10870 ( .B1(n10006), .B2(n9777), .A(n9768), .ZN(n9769) );
  AND2_X1 U10871 ( .A1(n10002), .A2(n9769), .ZN(n9805) );
  INV_X1 U10872 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n9770) );
  AOI22_X1 U10873 ( .A1(n9796), .A2(n9805), .B1(n9770), .B2(n9794), .ZN(
        P2_U3478) );
  INV_X1 U10874 ( .A(n9771), .ZN(n9776) );
  OAI22_X1 U10875 ( .A1(n9773), .A2(n9780), .B1(n9772), .B2(n9788), .ZN(n9775)
         );
  AOI211_X1 U10876 ( .C1(n9777), .C2(n9776), .A(n9775), .B(n9774), .ZN(n9806)
         );
  INV_X1 U10877 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n9778) );
  AOI22_X1 U10878 ( .A1(n9796), .A2(n9806), .B1(n9778), .B2(n9794), .ZN(
        P2_U3481) );
  OAI22_X1 U10879 ( .A1(n9781), .A2(n9780), .B1(n9779), .B2(n9788), .ZN(n9783)
         );
  AOI211_X1 U10880 ( .C1(n9784), .C2(n9793), .A(n9783), .B(n9782), .ZN(n9807)
         );
  INV_X1 U10881 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n9785) );
  AOI22_X1 U10882 ( .A1(n9796), .A2(n9807), .B1(n9785), .B2(n9794), .ZN(
        P2_U3484) );
  OAI21_X1 U10883 ( .B1(n4489), .B2(n9788), .A(n9787), .ZN(n9791) );
  INV_X1 U10884 ( .A(n9789), .ZN(n9790) );
  AOI211_X1 U10885 ( .C1(n9793), .C2(n9792), .A(n9791), .B(n9790), .ZN(n9809)
         );
  INV_X1 U10886 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n9795) );
  AOI22_X1 U10887 ( .A1(n9796), .A2(n9809), .B1(n9795), .B2(n9794), .ZN(
        P2_U3487) );
  INV_X1 U10888 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n9797) );
  AOI22_X1 U10889 ( .A1(n9810), .A2(n9798), .B1(n9797), .B2(n9808), .ZN(
        P2_U3520) );
  AOI22_X1 U10890 ( .A1(n9810), .A2(n9799), .B1(n7341), .B2(n9808), .ZN(
        P2_U3522) );
  INV_X1 U10891 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n9800) );
  AOI22_X1 U10892 ( .A1(n9810), .A2(n9801), .B1(n9800), .B2(n9808), .ZN(
        P2_U3524) );
  INV_X1 U10893 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n9802) );
  AOI22_X1 U10894 ( .A1(n9810), .A2(n9803), .B1(n9802), .B2(n9808), .ZN(
        P2_U3527) );
  AOI22_X1 U10895 ( .A1(n9810), .A2(n9804), .B1(n7350), .B2(n9808), .ZN(
        P2_U3528) );
  AOI22_X1 U10896 ( .A1(n9810), .A2(n9805), .B1(n7352), .B2(n9808), .ZN(
        P2_U3529) );
  AOI22_X1 U10897 ( .A1(n9810), .A2(n9806), .B1(n7354), .B2(n9808), .ZN(
        P2_U3530) );
  AOI22_X1 U10898 ( .A1(n9810), .A2(n9807), .B1(n7356), .B2(n9808), .ZN(
        P2_U3531) );
  AOI22_X1 U10899 ( .A1(n9810), .A2(n9809), .B1(n7358), .B2(n9808), .ZN(
        P2_U3532) );
  INV_X1 U10900 ( .A(n9811), .ZN(n9812) );
  NAND2_X1 U10901 ( .A1(n9813), .A2(n9812), .ZN(n9814) );
  XOR2_X1 U10902 ( .A(n9815), .B(n9814), .Z(ADD_1071_U5) );
  INV_X1 U10903 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n9816) );
  INV_X1 U10904 ( .A(P2_ADDR_REG_0__SCAN_IN), .ZN(n9849) );
  AOI22_X1 U10905 ( .A1(P2_ADDR_REG_0__SCAN_IN), .A2(P1_ADDR_REG_0__SCAN_IN), 
        .B1(n9816), .B2(n9849), .ZN(ADD_1071_U46) );
  OAI21_X1 U10906 ( .B1(n9819), .B2(n9818), .A(n9817), .ZN(ADD_1071_U56) );
  OAI21_X1 U10907 ( .B1(n9822), .B2(n9821), .A(n9820), .ZN(ADD_1071_U57) );
  OAI21_X1 U10908 ( .B1(n9825), .B2(n9824), .A(n9823), .ZN(ADD_1071_U58) );
  OAI21_X1 U10909 ( .B1(n9828), .B2(n9827), .A(n9826), .ZN(ADD_1071_U59) );
  OAI21_X1 U10910 ( .B1(n9831), .B2(n9830), .A(n9829), .ZN(ADD_1071_U60) );
  OAI21_X1 U10911 ( .B1(n9834), .B2(n9833), .A(n9832), .ZN(ADD_1071_U61) );
  AOI21_X1 U10912 ( .B1(n9837), .B2(n9836), .A(n9835), .ZN(ADD_1071_U62) );
  AOI21_X1 U10913 ( .B1(n9840), .B2(n9839), .A(n9838), .ZN(ADD_1071_U63) );
  AOI22_X1 U10914 ( .A1(n9842), .A2(keyinput49), .B1(keyinput0), .B2(n7356), 
        .ZN(n9841) );
  OAI221_X1 U10915 ( .B1(n9842), .B2(keyinput49), .C1(n7356), .C2(keyinput0), 
        .A(n9841), .ZN(n9855) );
  AOI22_X1 U10916 ( .A1(n9845), .A2(keyinput40), .B1(keyinput28), .B2(n9844), 
        .ZN(n9843) );
  OAI221_X1 U10917 ( .B1(n9845), .B2(keyinput40), .C1(n9844), .C2(keyinput28), 
        .A(n9843), .ZN(n9854) );
  AOI22_X1 U10918 ( .A1(n9848), .A2(keyinput22), .B1(n9847), .B2(keyinput50), 
        .ZN(n9846) );
  OAI221_X1 U10919 ( .B1(n9848), .B2(keyinput22), .C1(n9847), .C2(keyinput50), 
        .A(n9846), .ZN(n9853) );
  XOR2_X1 U10920 ( .A(n9849), .B(keyinput14), .Z(n9851) );
  XNOR2_X1 U10921 ( .A(P1_IR_REG_12__SCAN_IN), .B(keyinput59), .ZN(n9850) );
  NAND2_X1 U10922 ( .A1(n9851), .A2(n9850), .ZN(n9852) );
  NOR4_X1 U10923 ( .A1(n9855), .A2(n9854), .A3(n9853), .A4(n9852), .ZN(n9900)
         );
  AOI22_X1 U10924 ( .A1(n9973), .A2(keyinput46), .B1(n9857), .B2(keyinput19), 
        .ZN(n9856) );
  OAI221_X1 U10925 ( .B1(n9973), .B2(keyinput46), .C1(n9857), .C2(keyinput19), 
        .A(n9856), .ZN(n9868) );
  INV_X1 U10926 ( .A(SI_6_), .ZN(n9860) );
  AOI22_X1 U10927 ( .A1(n9860), .A2(keyinput42), .B1(keyinput7), .B2(n9859), 
        .ZN(n9858) );
  OAI221_X1 U10928 ( .B1(n9860), .B2(keyinput42), .C1(n9859), .C2(keyinput7), 
        .A(n9858), .ZN(n9867) );
  INV_X1 U10929 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n9862) );
  INV_X1 U10930 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n9972) );
  AOI22_X1 U10931 ( .A1(n9862), .A2(keyinput32), .B1(n9972), .B2(keyinput8), 
        .ZN(n9861) );
  OAI221_X1 U10932 ( .B1(n9862), .B2(keyinput32), .C1(n9972), .C2(keyinput8), 
        .A(n9861), .ZN(n9866) );
  INV_X1 U10933 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n9864) );
  AOI22_X1 U10934 ( .A1(n9864), .A2(keyinput48), .B1(keyinput58), .B2(n5622), 
        .ZN(n9863) );
  OAI221_X1 U10935 ( .B1(n9864), .B2(keyinput48), .C1(n5622), .C2(keyinput58), 
        .A(n9863), .ZN(n9865) );
  NOR4_X1 U10936 ( .A1(n9868), .A2(n9867), .A3(n9866), .A4(n9865), .ZN(n9899)
         );
  AOI22_X1 U10937 ( .A1(n9870), .A2(keyinput24), .B1(keyinput29), .B2(n6033), 
        .ZN(n9869) );
  OAI221_X1 U10938 ( .B1(n9870), .B2(keyinput24), .C1(n6033), .C2(keyinput29), 
        .A(n9869), .ZN(n9881) );
  INV_X1 U10939 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n9872) );
  AOI22_X1 U10940 ( .A1(n9872), .A2(keyinput52), .B1(n6723), .B2(keyinput55), 
        .ZN(n9871) );
  OAI221_X1 U10941 ( .B1(n9872), .B2(keyinput52), .C1(n6723), .C2(keyinput55), 
        .A(n9871), .ZN(n9880) );
  INV_X1 U10942 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n9874) );
  AOI22_X1 U10943 ( .A1(n9875), .A2(keyinput53), .B1(keyinput34), .B2(n9874), 
        .ZN(n9873) );
  OAI221_X1 U10944 ( .B1(n9875), .B2(keyinput53), .C1(n9874), .C2(keyinput34), 
        .A(n9873), .ZN(n9879) );
  XNOR2_X1 U10945 ( .A(P2_IR_REG_12__SCAN_IN), .B(keyinput35), .ZN(n9877) );
  XNOR2_X1 U10946 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(keyinput57), .ZN(n9876)
         );
  NAND2_X1 U10947 ( .A1(n9877), .A2(n9876), .ZN(n9878) );
  NOR4_X1 U10948 ( .A1(n9881), .A2(n9880), .A3(n9879), .A4(n9878), .ZN(n9898)
         );
  AOI22_X1 U10949 ( .A1(n9884), .A2(keyinput62), .B1(keyinput36), .B2(n9883), 
        .ZN(n9882) );
  OAI221_X1 U10950 ( .B1(n9884), .B2(keyinput62), .C1(n9883), .C2(keyinput36), 
        .A(n9882), .ZN(n9896) );
  AOI22_X1 U10951 ( .A1(n9887), .A2(keyinput17), .B1(keyinput2), .B2(n9886), 
        .ZN(n9885) );
  OAI221_X1 U10952 ( .B1(n9887), .B2(keyinput17), .C1(n9886), .C2(keyinput2), 
        .A(n9885), .ZN(n9895) );
  AOI22_X1 U10953 ( .A1(n9890), .A2(keyinput51), .B1(n9889), .B2(keyinput38), 
        .ZN(n9888) );
  OAI221_X1 U10954 ( .B1(n9890), .B2(keyinput51), .C1(n9889), .C2(keyinput38), 
        .A(n9888), .ZN(n9894) );
  XNOR2_X1 U10955 ( .A(P1_REG2_REG_24__SCAN_IN), .B(keyinput56), .ZN(n9892) );
  XNOR2_X1 U10956 ( .A(SI_2_), .B(keyinput61), .ZN(n9891) );
  NAND2_X1 U10957 ( .A1(n9892), .A2(n9891), .ZN(n9893) );
  NOR4_X1 U10958 ( .A1(n9896), .A2(n9895), .A3(n9894), .A4(n9893), .ZN(n9897)
         );
  NAND4_X1 U10959 ( .A1(n9900), .A2(n9899), .A3(n9898), .A4(n9897), .ZN(n9964)
         );
  AOI22_X1 U10960 ( .A1(n9903), .A2(keyinput31), .B1(n9902), .B2(keyinput43), 
        .ZN(n9901) );
  OAI221_X1 U10961 ( .B1(n9903), .B2(keyinput31), .C1(n9902), .C2(keyinput43), 
        .A(n9901), .ZN(n9915) );
  AOI22_X1 U10962 ( .A1(n9965), .A2(keyinput44), .B1(keyinput39), .B2(n9905), 
        .ZN(n9904) );
  OAI221_X1 U10963 ( .B1(n9965), .B2(keyinput44), .C1(n9905), .C2(keyinput39), 
        .A(n9904), .ZN(n9914) );
  AOI22_X1 U10964 ( .A1(n9908), .A2(keyinput54), .B1(keyinput12), .B2(n9907), 
        .ZN(n9906) );
  OAI221_X1 U10965 ( .B1(n9908), .B2(keyinput54), .C1(n9907), .C2(keyinput12), 
        .A(n9906), .ZN(n9913) );
  INV_X1 U10966 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n9910) );
  AOI22_X1 U10967 ( .A1(n9911), .A2(keyinput18), .B1(keyinput47), .B2(n9910), 
        .ZN(n9909) );
  OAI221_X1 U10968 ( .B1(n9911), .B2(keyinput18), .C1(n9910), .C2(keyinput47), 
        .A(n9909), .ZN(n9912) );
  NOR4_X1 U10969 ( .A1(n9915), .A2(n9914), .A3(n9913), .A4(n9912), .ZN(n9962)
         );
  AOI22_X1 U10970 ( .A1(n9918), .A2(keyinput10), .B1(n9917), .B2(keyinput60), 
        .ZN(n9916) );
  OAI221_X1 U10971 ( .B1(n9918), .B2(keyinput10), .C1(n9917), .C2(keyinput60), 
        .A(n9916), .ZN(n9930) );
  INV_X1 U10972 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n9920) );
  AOI22_X1 U10973 ( .A1(n9921), .A2(keyinput63), .B1(keyinput16), .B2(n9920), 
        .ZN(n9919) );
  OAI221_X1 U10974 ( .B1(n9921), .B2(keyinput63), .C1(n9920), .C2(keyinput16), 
        .A(n9919), .ZN(n9929) );
  INV_X1 U10975 ( .A(SI_21_), .ZN(n9923) );
  AOI22_X1 U10976 ( .A1(n9924), .A2(keyinput21), .B1(n9923), .B2(keyinput27), 
        .ZN(n9922) );
  OAI221_X1 U10977 ( .B1(n9924), .B2(keyinput21), .C1(n9923), .C2(keyinput27), 
        .A(n9922), .ZN(n9928) );
  AOI22_X1 U10978 ( .A1(n9966), .A2(keyinput4), .B1(n9926), .B2(keyinput20), 
        .ZN(n9925) );
  OAI221_X1 U10979 ( .B1(n9966), .B2(keyinput4), .C1(n9926), .C2(keyinput20), 
        .A(n9925), .ZN(n9927) );
  NOR4_X1 U10980 ( .A1(n9930), .A2(n9929), .A3(n9928), .A4(n9927), .ZN(n9961)
         );
  INV_X1 U10981 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n9932) );
  AOI22_X1 U10982 ( .A1(n9933), .A2(keyinput33), .B1(keyinput1), .B2(n9932), 
        .ZN(n9931) );
  OAI221_X1 U10983 ( .B1(n9933), .B2(keyinput33), .C1(n9932), .C2(keyinput1), 
        .A(n9931), .ZN(n9945) );
  AOI22_X1 U10984 ( .A1(n9978), .A2(keyinput26), .B1(n9935), .B2(keyinput30), 
        .ZN(n9934) );
  OAI221_X1 U10985 ( .B1(n9978), .B2(keyinput26), .C1(n9935), .C2(keyinput30), 
        .A(n9934), .ZN(n9944) );
  AOI22_X1 U10986 ( .A1(n9938), .A2(keyinput3), .B1(n9937), .B2(keyinput15), 
        .ZN(n9936) );
  OAI221_X1 U10987 ( .B1(n9938), .B2(keyinput3), .C1(n9937), .C2(keyinput15), 
        .A(n9936), .ZN(n9943) );
  XOR2_X1 U10988 ( .A(n9939), .B(keyinput11), .Z(n9941) );
  XNOR2_X1 U10989 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(keyinput13), .ZN(n9940) );
  NAND2_X1 U10990 ( .A1(n9941), .A2(n9940), .ZN(n9942) );
  NOR4_X1 U10991 ( .A1(n9945), .A2(n9944), .A3(n9943), .A4(n9942), .ZN(n9960)
         );
  AOI22_X1 U10992 ( .A1(n9947), .A2(keyinput25), .B1(n7350), .B2(keyinput6), 
        .ZN(n9946) );
  OAI221_X1 U10993 ( .B1(n9947), .B2(keyinput25), .C1(n7350), .C2(keyinput6), 
        .A(n9946), .ZN(n9958) );
  AOI22_X1 U10994 ( .A1(n9949), .A2(keyinput37), .B1(keyinput45), .B2(n7455), 
        .ZN(n9948) );
  OAI221_X1 U10995 ( .B1(n9949), .B2(keyinput37), .C1(n7455), .C2(keyinput45), 
        .A(n9948), .ZN(n9957) );
  AOI22_X1 U10996 ( .A1(n8584), .A2(keyinput23), .B1(keyinput5), .B2(n9951), 
        .ZN(n9950) );
  OAI221_X1 U10997 ( .B1(n8584), .B2(keyinput23), .C1(n9951), .C2(keyinput5), 
        .A(n9950), .ZN(n9956) );
  INV_X1 U10998 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n9952) );
  XOR2_X1 U10999 ( .A(n9952), .B(keyinput9), .Z(n9954) );
  XNOR2_X1 U11000 ( .A(P2_IR_REG_1__SCAN_IN), .B(keyinput41), .ZN(n9953) );
  NAND2_X1 U11001 ( .A1(n9954), .A2(n9953), .ZN(n9955) );
  NOR4_X1 U11002 ( .A1(n9958), .A2(n9957), .A3(n9956), .A4(n9955), .ZN(n9959)
         );
  NAND4_X1 U11003 ( .A1(n9962), .A2(n9961), .A3(n9960), .A4(n9959), .ZN(n9963)
         );
  NOR2_X1 U11004 ( .A1(n9964), .A2(n9963), .ZN(n10010) );
  NAND4_X1 U11005 ( .A1(P1_DATAO_REG_6__SCAN_IN), .A2(SI_6_), .A3(
        P1_DATAO_REG_3__SCAN_IN), .A4(n9965), .ZN(n9992) );
  NOR4_X1 U11006 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .A3(P1_ADDR_REG_5__SCAN_IN), .A4(n9966), .ZN(n9971) );
  NOR2_X1 U11007 ( .A1(P2_RD_REG_SCAN_IN), .A2(n7455), .ZN(n9967) );
  AND4_X1 U11008 ( .A1(n9968), .A2(P2_IR_REG_1__SCAN_IN), .A3(n9967), .A4(
        n4731), .ZN(n9969) );
  NAND3_X1 U11009 ( .A1(n9971), .A2(n9970), .A3(n9969), .ZN(n9991) );
  NOR4_X1 U11010 ( .A1(SI_15_), .A2(P2_REG0_REG_26__SCAN_IN), .A3(
        P2_REG0_REG_19__SCAN_IN), .A4(P2_REG1_REG_11__SCAN_IN), .ZN(n9977) );
  NOR4_X1 U11011 ( .A1(P1_DATAO_REG_21__SCAN_IN), .A2(P1_REG3_REG_16__SCAN_IN), 
        .A3(P1_REG0_REG_2__SCAN_IN), .A4(P1_REG0_REG_31__SCAN_IN), .ZN(n9976)
         );
  NOR4_X1 U11012 ( .A1(P1_REG3_REG_19__SCAN_IN), .A2(P1_REG3_REG_11__SCAN_IN), 
        .A3(P1_REG2_REG_11__SCAN_IN), .A4(P2_DATAO_REG_31__SCAN_IN), .ZN(n9975) );
  NOR4_X1 U11013 ( .A1(P1_REG2_REG_10__SCAN_IN), .A2(P2_REG2_REG_30__SCAN_IN), 
        .A3(n9973), .A4(n9972), .ZN(n9974) );
  NAND4_X1 U11014 ( .A1(n9977), .A2(n9976), .A3(n9975), .A4(n9974), .ZN(n9990)
         );
  NOR4_X1 U11015 ( .A1(P1_IR_REG_23__SCAN_IN), .A2(P2_DATAO_REG_18__SCAN_IN), 
        .A3(P1_DATAO_REG_17__SCAN_IN), .A4(n9978), .ZN(n9988) );
  NOR4_X1 U11016 ( .A1(P1_IR_REG_12__SCAN_IN), .A2(SI_21_), .A3(
        P2_REG1_REG_29__SCAN_IN), .A4(P2_REG0_REG_31__SCAN_IN), .ZN(n9987) );
  NAND2_X1 U11017 ( .A1(SI_9_), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n9980) );
  NAND4_X1 U11018 ( .A1(P2_D_REG_13__SCAN_IN), .A2(P2_REG2_REG_2__SCAN_IN), 
        .A3(P2_REG3_REG_1__SCAN_IN), .A4(P2_REG3_REG_0__SCAN_IN), .ZN(n9979)
         );
  NOR4_X1 U11019 ( .A1(SI_2_), .A2(P2_REG1_REG_8__SCAN_IN), .A3(n9980), .A4(
        n9979), .ZN(n9986) );
  NAND4_X1 U11020 ( .A1(P1_IR_REG_18__SCAN_IN), .A2(P1_D_REG_22__SCAN_IN), 
        .A3(P1_DATAO_REG_15__SCAN_IN), .A4(P1_REG2_REG_17__SCAN_IN), .ZN(n9984) );
  NAND4_X1 U11021 ( .A1(P1_IR_REG_7__SCAN_IN), .A2(P1_DATAO_REG_14__SCAN_IN), 
        .A3(P1_REG2_REG_24__SCAN_IN), .A4(P1_WR_REG_SCAN_IN), .ZN(n9983) );
  NAND4_X1 U11022 ( .A1(P1_D_REG_7__SCAN_IN), .A2(P1_REG1_REG_18__SCAN_IN), 
        .A3(P1_REG0_REG_5__SCAN_IN), .A4(P2_REG3_REG_20__SCAN_IN), .ZN(n9982)
         );
  NAND4_X1 U11023 ( .A1(P1_REG1_REG_26__SCAN_IN), .A2(P2_REG0_REG_25__SCAN_IN), 
        .A3(P2_REG2_REG_21__SCAN_IN), .A4(P2_REG0_REG_24__SCAN_IN), .ZN(n9981)
         );
  NOR4_X1 U11024 ( .A1(n9984), .A2(n9983), .A3(n9982), .A4(n9981), .ZN(n9985)
         );
  NAND4_X1 U11025 ( .A1(n9988), .A2(n9987), .A3(n9986), .A4(n9985), .ZN(n9989)
         );
  NOR4_X1 U11026 ( .A1(n9992), .A2(n9991), .A3(n9990), .A4(n9989), .ZN(n10008)
         );
  AOI22_X1 U11027 ( .A1(n10001), .A2(P2_REG2_REG_9__SCAN_IN), .B1(n9994), .B2(
        n9993), .ZN(n9998) );
  NAND2_X1 U11028 ( .A1(n9996), .A2(n9995), .ZN(n9997) );
  OAI211_X1 U11029 ( .C1(n10000), .C2(n9999), .A(n9998), .B(n9997), .ZN(n10004) );
  NOR2_X1 U11030 ( .A1(n10002), .A2(n10001), .ZN(n10003) );
  AOI211_X1 U11031 ( .C1(n10006), .C2(n10005), .A(n10004), .B(n10003), .ZN(
        n10007) );
  XOR2_X1 U11032 ( .A(n10008), .B(n10007), .Z(n10009) );
  XNOR2_X1 U11033 ( .A(n10010), .B(n10009), .ZN(P2_U3287) );
  XOR2_X1 U11034 ( .A(n10011), .B(P2_ADDR_REG_8__SCAN_IN), .Z(ADD_1071_U48) );
  XOR2_X1 U11035 ( .A(n10012), .B(P2_ADDR_REG_6__SCAN_IN), .Z(ADD_1071_U50) );
  NOR2_X1 U11036 ( .A1(n10014), .A2(n10013), .ZN(n10015) );
  XOR2_X1 U11037 ( .A(n10015), .B(P1_ADDR_REG_5__SCAN_IN), .Z(ADD_1071_U51) );
  XOR2_X1 U11038 ( .A(n10016), .B(P2_ADDR_REG_7__SCAN_IN), .Z(ADD_1071_U49) );
  OAI21_X1 U11039 ( .B1(n10019), .B2(n10018), .A(n10017), .ZN(n10020) );
  XNOR2_X1 U11040 ( .A(n10020), .B(P1_ADDR_REG_18__SCAN_IN), .ZN(ADD_1071_U55)
         );
  AOI21_X1 U11041 ( .B1(n10023), .B2(n10022), .A(n10021), .ZN(ADD_1071_U47) );
  XOR2_X1 U11042 ( .A(n10025), .B(n10024), .Z(ADD_1071_U54) );
  XOR2_X1 U11043 ( .A(n10027), .B(n10026), .Z(ADD_1071_U53) );
  XNOR2_X1 U11044 ( .A(n10029), .B(n10028), .ZN(ADD_1071_U52) );
  CLKBUF_X1 U4782 ( .A(n6628), .Z(n4263) );
  BUF_X2 U4778 ( .A(n4935), .Z(n5554) );
  CLKBUF_X1 U4794 ( .A(n4265), .Z(n6629) );
  CLKBUF_X1 U4795 ( .A(n6628), .Z(n4264) );
endmodule

